module aes_core(clk, rst, ld, done, key, text_in, text_out);
input clk, rst, ld;
input [127:0] key, text_in;
output done;
output [127:0] text_out;
wire clk, rst, ld;
wire [127:0] key, text_in;
wire done;
wire [127:0] text_out;
wire dcnt[0] , dcnt[1] , dcnt[2] , dcnt[3] , ld_r, n_0, n_2, n_9;
wire n_14, n_15, n_18, n_21, n_22, n_26, n_62, n_63;
wire n_68, n_77, n_89, n_95, n_97, n_98, n_100, n_101;
wire n_106, n_107, n_109, n_111, n_112, n_123, n_124, n_129;
wire n_135, n_141, n_152, n_153, n_160, n_162, n_164, n_165;
wire n_167, n_171, n_176, n_177, n_178, n_183, n_187, n_191;
wire n_194, n_196, n_199, n_205, n_207, n_208, n_209, n_213;
wire n_214, n_218, n_221, n_228, n_229, n_230, n_234, n_238;
wire n_243, n_245, n_250, n_251, n_255, n_263, n_264, n_267;
wire n_271, n_273, n_274, n_276, n_277, n_279, n_280, n_282;
wire n_285, n_288, n_290, n_294, n_295, n_296, n_300, n_303;
wire n_305, n_310, n_315, n_319, n_320, n_328, n_330, n_332;
wire n_338, n_341, n_342, n_343, n_344, n_348, n_352, n_357;
wire n_360, n_362, n_367, n_370, n_377, n_378, n_379, n_380;
wire n_381, n_383, n_384, n_386, n_393, n_398, n_399, n_400;
wire n_408, n_424, n_427, n_430, n_434, n_435, n_437, n_440;
wire n_441, n_454, n_457, n_459, n_462, n_463, n_464, n_469;
wire n_470, n_473, n_474, n_477, n_479, n_481, n_482, n_485;
wire n_487, n_488, n_490, n_493, n_494, n_497, n_503, n_508;
wire n_509, n_510, n_514, n_519, n_523, n_525, n_527, n_528;
wire n_529, n_530, n_532, n_537, n_538, n_540, n_541, n_544;
wire n_546, n_547, n_557, n_561, n_563, n_569, n_571, n_575;
wire n_578, n_579, n_581, n_583, n_584, n_587, n_591, n_596;
wire n_600, n_606, n_607, n_612, n_619, n_622, n_623, n_624;
wire n_627, n_629, n_630, n_631, n_632, n_636, n_638, n_645;
wire n_646, n_654, n_656, n_663, n_664, n_665, n_668, n_669;
wire n_671, n_672, n_673, n_674, n_677, n_684, n_688, n_698;
wire n_706, n_709, n_713, n_714, n_718, n_719, n_720, n_730;
wire n_731, n_732, n_735, n_736, n_744, n_748, n_749, n_751;
wire n_753, n_755, n_759, n_764, n_767, n_770, n_772, n_773;
wire n_775, n_778, n_783, n_788, n_789, n_790, n_791, n_795;
wire n_801, n_802, n_803, n_804, n_805, n_807, n_818, n_819;
wire n_821, n_825, n_826, n_827, n_828, n_829, n_833, n_834;
wire n_844, n_849, n_850, n_853, n_862, n_867, n_868, n_869;
wire n_870, n_871, n_872, n_875, n_877, n_880, n_881, n_883;
wire n_884, n_894, n_896, n_897, n_899, n_900, n_901, n_902;
wire n_903, n_908, n_912, n_913, n_916, n_917, n_919, n_920;
wire n_925, n_926, n_931, n_932, n_933, n_941, n_959, n_960;
wire n_962, n_964, n_967, n_968, n_969, n_972, n_974, n_975;
wire n_976, n_977, n_980, n_981, n_982, n_983, n_986, n_988;
wire n_989, n_993, n_995, n_997, n_999, n_1000, n_1002, n_1003;
wire n_1004, n_1005, n_1006, n_1008, n_1010, n_1012, n_1014, n_1015;
wire n_1016, n_1018, n_1019, n_1020, n_1036, n_1037, n_1038, n_1039;
wire n_1040, n_1041, n_1043, n_1044, n_1046, n_1050, n_1051, n_1053;
wire n_1057, n_1063, n_1064, n_1065, n_1069, n_1072, n_1073, n_1074;
wire n_1075, n_1079, n_1080, n_1081, n_1082, n_1083, n_1085, n_1087;
wire n_1088, n_1098, n_1102, n_1103, n_1104, n_1106, n_1109, n_1110;
wire n_1113, n_1118, n_1120, n_1124, n_1125, n_1127, n_1129, n_1132;
wire n_1134, n_1135, n_1138, n_1140, n_1142, n_1147, n_1153, n_1155;
wire n_1157, n_1158, n_1163, n_1164, n_1165, n_1166, n_1173, n_1176;
wire n_1177, n_1185, n_1186, n_1191, n_1196, n_1198, n_1201, n_1204;
wire n_1205, n_1206, n_1212, n_1213, n_1217, n_1220, n_1221, n_1223;
wire n_1224, n_1226, n_1227, n_1228, n_1229, n_1230, n_1233, n_1235;
wire n_1236, n_1237, n_1238, n_1239, n_1241, n_1242, n_1243, n_1244;
wire n_1246, n_1248, n_1251, n_1252, n_1253, n_1255, n_1256, n_1258;
wire n_1260, n_1261, n_1263, n_1264, n_1266, n_1267, n_1268, n_1270;
wire n_1271, n_1272, n_1273, n_1278, n_1281, n_1282, n_1283, n_1284;
wire n_1285, n_1289, n_1291, n_1292, n_1294, n_1295, n_1296, n_1297;
wire n_1298, n_1302, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310;
wire n_1312, n_1313, n_1315, n_1316, n_1318, n_1319, n_1321, n_1324;
wire n_1325, n_1331, n_1332, n_1333, n_1335, n_1336, n_1339, n_1340;
wire n_1341, n_1347, n_1350, n_1353, n_1358, n_1361, n_1363, n_1365;
wire n_1368, n_1370, n_1371, n_1373, n_1376, n_1377, n_1378, n_1384;
wire n_1385, n_1386, n_1387, n_1389, n_1390, n_1395, n_1396, n_1397;
wire n_1402, n_1409, n_1416, n_1417, n_1423, n_1424, n_1427, n_1428;
wire n_1429, n_1430, n_1431, n_1441, n_1443, n_1447, n_1448, n_1456;
wire n_1457, n_1460, n_1461, n_1473, n_1477, n_1480, n_1483, n_1484;
wire n_1488, n_1491, n_1493, n_1494, n_1497, n_1500, n_1501, n_1502;
wire n_1503, n_1505, n_1507, n_1508, n_1509, n_1512, n_1513, n_1516;
wire n_1522, n_1525, n_1526, n_1528, n_1530, n_1531, n_1534, n_1538;
wire n_1539, n_1540, n_1541, n_1542, n_1544, n_1546, n_1547, n_1548;
wire n_1551, n_1552, n_1553, n_1555, n_1556, n_1558, n_1560, n_1562;
wire n_1564, n_1565, n_1568, n_1569, n_1570, n_1571, n_1572, n_1576;
wire n_1578, n_1581, n_1582, n_1584, n_1585, n_1588, n_1589, n_1591;
wire n_1593, n_1594, n_1599, n_1600, n_1601, n_1603, n_1606, n_1608;
wire n_1609, n_1610, n_1614, n_1615, n_1616, n_1618, n_1620, n_1621;
wire n_1626, n_1627, n_1628, n_1630, n_1632, n_1633, n_1634, n_1636;
wire n_1637, n_1641, n_1642, n_1644, n_1645, n_1647, n_1648, n_1651;
wire n_1653, n_1656, n_1658, n_1666, n_1667, n_1668, n_1671, n_1674;
wire n_1675, n_1678, n_1679, n_1683, n_1685, n_1686, n_1688, n_1691;
wire n_1693, n_1694, n_1695, n_1698, n_1699, n_1701, n_1706, n_1707;
wire n_1711, n_1712, n_1717, n_1724, n_1727, n_1731, n_1734, n_1735;
wire n_1736, n_1737, n_1739, n_1741, n_1742, n_1743, n_1744, n_1745;
wire n_1746, n_1747, n_1748, n_1749, n_1750, n_1752, n_1756, n_1758;
wire n_1760, n_1763, n_1768, n_1769, n_1770, n_1771, n_1772, n_1775;
wire n_1777, n_1779, n_1781, n_1782, n_1784, n_1786, n_1788, n_1789;
wire n_1791, n_1792, n_1797, n_1798, n_1805, n_1806, n_1807, n_1809;
wire n_1811, n_1813, n_1816, n_1817, n_1818, n_1819, n_1821, n_1822;
wire n_1823, n_1825, n_1827, n_1830, n_1833, n_1835, n_1837, n_1839;
wire n_1840, n_1842, n_1843, n_1845, n_1850, n_1851, n_1852, n_1854;
wire n_1858, n_1868, n_1874, n_1883, n_1886, n_1887, n_1888, n_1890;
wire n_1891, n_1895, n_1897, n_1899, n_1902, n_1904, n_1905, n_1907;
wire n_1911, n_1914, n_1915, n_1916, n_1918, n_1920, n_1921, n_1923;
wire n_1925, n_1928, n_1929, n_1930, n_1933, n_1934, n_1936, n_1938;
wire n_1939, n_1941, n_1942, n_1943, n_1946, n_1947, n_1954, n_1955;
wire n_1956, n_1958, n_1959, n_1960, n_1961, n_1963, n_1965, n_1968;
wire n_1969, n_1970, n_1971, n_1972, n_1982, n_1983, n_1984, n_1985;
wire n_1986, n_1987, n_1988, n_1989, n_1991, n_1993, n_1995, n_1996;
wire n_1997, n_1998, n_2001, n_2004, n_2007, n_2008, n_2009, n_2010;
wire n_2013, n_2017, n_2021, n_2022, n_2024, n_2025, n_2026, n_2035;
wire n_2040, n_2042, n_2043, n_2044, n_2047, n_2048, n_2049, n_2051;
wire n_2052, n_2053, n_2055, n_2060, n_2062, n_2063, n_2066, n_2067;
wire n_2069, n_2070, n_2071, n_2074, n_2076, n_2078, n_2079, n_2081;
wire n_2084, n_2085, n_2086, n_2089, n_2090, n_2091, n_2092, n_2093;
wire n_2094, n_2095, n_2096, n_2099, n_2100, n_2102, n_2105, n_2107;
wire n_2109, n_2111, n_2112, n_2113, n_2119, n_2121, n_2124, n_2125;
wire n_2128, n_2131, n_2135, n_2137, n_2140, n_2145, n_2146, n_2148;
wire n_2150, n_2151, n_2152, n_2153, n_2158, n_2160, n_2162, n_2164;
wire n_2168, n_2170, n_2173, n_2174, n_2175, n_2176, n_2180, n_2181;
wire n_2183, n_2185, n_2187, n_2191, n_2198, n_2201, n_2204, n_2206;
wire n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216;
wire n_2217, n_2218, n_2220, n_2227, n_2228, n_2229, n_2231, n_2234;
wire n_2235, n_2236, n_2237, n_2239, n_2241, n_2244, n_2247, n_2249;
wire n_2251, n_2253, n_2254, n_2259, n_2260, n_2265, n_2266, n_2267;
wire n_2276, n_2278, n_2279, n_2281, n_2286, n_2289, n_2290, n_2291;
wire n_2292, n_2295, n_2297, n_2298, n_2301, n_2302, n_2303, n_2304;
wire n_2305, n_2306, n_2307, n_2311, n_2318, n_2319, n_2320, n_2322;
wire n_2323, n_2324, n_2327, n_2329, n_2330, n_2331, n_2332, n_2333;
wire n_2334, n_2335, n_2336, n_2337, n_2342, n_2343, n_2344, n_2345;
wire n_2346, n_2349, n_2350, n_2351, n_2352, n_2353, n_2356, n_2357;
wire n_2359, n_2360, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367;
wire n_2368, n_2369, n_2372, n_2373, n_2374, n_2376, n_2380, n_2382;
wire n_2383, n_2384, n_2385, n_2386, n_2387, n_2390, n_2392, n_2393;
wire n_2394, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402;
wire n_2403, n_2404, n_2405, n_2406, n_2408, n_2409, n_2412, n_2413;
wire n_2415, n_2416, n_2417, n_2418, n_2420, n_2422, n_2423, n_2424;
wire n_2425, n_2426, n_2429, n_2430, n_2431, n_2433, n_2434, n_2435;
wire n_2436, n_2437, n_2438, n_2440, n_2441, n_2444, n_2446, n_2447;
wire n_2450, n_2452, n_2455, n_2456, n_2457, n_2459, n_2460, n_2461;
wire n_2462, n_2464, n_2466, n_2467, n_2468, n_2469, n_2470, n_2479;
wire n_2480, n_2481, n_2483, n_2484, n_2485, n_2487, n_2488, n_2492;
wire n_2494, n_2496, n_2502, n_2503, n_2505, n_2509, n_2510, n_2511;
wire n_2513, n_2514, n_2515, n_2516, n_2519, n_2521, n_2522, n_2524;
wire n_2526, n_2527, n_2530, n_2532, n_2534, n_2536, n_2537, n_2540;
wire n_2541, n_2543, n_2544, n_2547, n_2548, n_2550, n_2552, n_2555;
wire n_2556, n_2559, n_2560, n_2561, n_2563, n_2565, n_2568, n_2569;
wire n_2570, n_2573, n_2574, n_2575, n_2577, n_2580, n_2583, n_2585;
wire n_2586, n_2587, n_2588, n_2590, n_2591, n_2592, n_2594, n_2595;
wire n_2596, n_2598, n_2603, n_2604, n_2605, n_2606, n_2608, n_2609;
wire n_2611, n_2612, n_2613, n_2616, n_2617, n_2621, n_2623, n_2625;
wire n_2627, n_2628, n_2632, n_2633, n_2635, n_2636, n_2638, n_2639;
wire n_2640, n_2641, n_2643, n_2645, n_2646, n_2647, n_2648, n_2650;
wire n_2654, n_2655, n_2656, n_2658, n_2660, n_2662, n_2663, n_2664;
wire n_2665, n_2671, n_2672, n_2674, n_2676, n_2678, n_2680, n_2681;
wire n_2682, n_2683, n_2684, n_2687, n_2691, n_2692, n_2693, n_2694;
wire n_2695, n_2696, n_2699, n_2700, n_2701, n_2702, n_2704, n_2705;
wire n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2713, n_2714;
wire n_2715, n_2716, n_2718, n_2719, n_2720, n_2723, n_2724, n_2732;
wire n_2733, n_2738, n_2739, n_2741, n_2742, n_2743, n_2744, n_2745;
wire n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755;
wire n_2757, n_2760, n_2766, n_2768, n_2769, n_2770, n_2771, n_2772;
wire n_2774, n_2775, n_2777, n_2779, n_2781, n_2785, n_2787, n_2792;
wire n_2794, n_2795, n_2796, n_2798, n_2800, n_2803, n_2804, n_2805;
wire n_2807, n_2809, n_2810, n_2811, n_2818, n_2819, n_2820, n_2821;
wire n_2823, n_2824, n_2826, n_2827, n_2829, n_2830, n_2831, n_2834;
wire n_2835, n_2837, n_2838, n_2839, n_2843, n_2846, n_2848, n_2849;
wire n_2850, n_2852, n_2856, n_2859, n_2861, n_2862, n_2864, n_2865;
wire n_2868, n_2870, n_2872, n_2873, n_2875, n_2878, n_2880, n_2881;
wire n_2883, n_2884, n_2885, n_2886, n_2888, n_2889, n_2890, n_2891;
wire n_2892, n_2894, n_2895, n_2900, n_2901, n_2902, n_2905, n_2908;
wire n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2916, n_2917;
wire n_2918, n_2919, n_2921, n_2923, n_2924, n_2925, n_2926, n_2927;
wire n_2929, n_2930, n_2931, n_2933, n_2934, n_2935, n_2937, n_2938;
wire n_2943, n_2945, n_2950, n_2952, n_2954, n_2958, n_2959, n_2960;
wire n_2962, n_2968, n_2969, n_2972, n_2973, n_2978, n_2981, n_2983;
wire n_2988, n_2989, n_2990, n_2991, n_2993, n_2994, n_2999, n_3000;
wire n_3001, n_3002, n_3003, n_3005, n_3010, n_3013, n_3014, n_3016;
wire n_3017, n_3018, n_3020, n_3021, n_3022, n_3023, n_3024, n_3029;
wire n_3030, n_3032, n_3033, n_3034, n_3038, n_3039, n_3040, n_3041;
wire n_3044, n_3045, n_3046, n_3047, n_3049, n_3050, n_3052, n_3053;
wire n_3055, n_3059, n_3060, n_3065, n_3067, n_3069, n_3070, n_3071;
wire n_3073, n_3076, n_3077, n_3079, n_3080, n_3081, n_3082, n_3083;
wire n_3084, n_3085, n_3086, n_3087, n_3089, n_3091, n_3093, n_3096;
wire n_3097, n_3101, n_3102, n_3104, n_3105, n_3106, n_3107, n_3108;
wire n_3112, n_3119, n_3121, n_3122, n_3125, n_3126, n_3128, n_3130;
wire n_3131, n_3132, n_3133, n_3134, n_3135, n_3138, n_3141, n_3142;
wire n_3144, n_3145, n_3147, n_3148, n_3149, n_3150, n_3153, n_3157;
wire n_3159, n_3160, n_3161, n_3162, n_3163, n_3165, n_3166, n_3167;
wire n_3168, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176;
wire n_3177, n_3180, n_3183, n_3184, n_3186, n_3187, n_3192, n_3193;
wire n_3195, n_3197, n_3198, n_3199, n_3201, n_3202, n_3203, n_3204;
wire n_3206, n_3208, n_3209, n_3210, n_3212, n_3213, n_3214, n_3216;
wire n_3218, n_3219, n_3220, n_3221, n_3223, n_3224, n_3225, n_3226;
wire n_3227, n_3228, n_3230, n_3231, n_3232, n_3234, n_3235, n_3236;
wire n_3237, n_3240, n_3241, n_3242, n_3244, n_3245, n_3246, n_3247;
wire n_3248, n_3250, n_3251, n_3252, n_3253, n_3254, n_3256, n_3257;
wire n_3258, n_3260, n_3261, n_3264, n_3266, n_3267, n_3268, n_3269;
wire n_3270, n_3273, n_3276, n_3277, n_3279, n_3281, n_3282, n_3283;
wire n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291;
wire n_3292, n_3294, n_3295, n_3296, n_3297, n_3300, n_3301, n_3302;
wire n_3303, n_3304, n_3305, n_3306, n_3307, n_3310, n_3312, n_3314;
wire n_3316, n_3317, n_3318, n_3319, n_3322, n_3323, n_3326, n_3327;
wire n_3328, n_3329, n_3330, n_3331, n_3332, n_3334, n_3336, n_3338;
wire n_3339, n_3340, n_3341, n_3342, n_3343, n_3345, n_3346, n_3347;
wire n_3348, n_3349, n_3350, n_3353, n_3354, n_3358, n_3359, n_3362;
wire n_3364, n_3365, n_3366, n_3367, n_3372, n_3373, n_3375, n_3380;
wire n_3381, n_3384, n_3385, n_3386, n_3388, n_3390, n_3391, n_3393;
wire n_3394, n_3395, n_3396, n_3398, n_3399, n_3401, n_3402, n_3403;
wire n_3404, n_3405, n_3406, n_3407, n_3409, n_3410, n_3411, n_3417;
wire n_3418, n_3419, n_3420, n_3421, n_3422, n_3425, n_3427, n_3429;
wire n_3433, n_3437, n_3438, n_3443, n_3444, n_3445, n_3448, n_3449;
wire n_3454, n_3455, n_3456, n_3457, n_3459, n_3460, n_3461, n_3463;
wire n_3464, n_3465, n_3466, n_3467, n_3469, n_3471, n_3473, n_3475;
wire n_3480, n_3482, n_3483, n_3485, n_3488, n_3489, n_3491, n_3493;
wire n_3494, n_3495, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503;
wire n_3504, n_3505, n_3506, n_3511, n_3512, n_3513, n_3514, n_3517;
wire n_3518, n_3519, n_3521, n_3522, n_3530, n_3532, n_3533, n_3534;
wire n_3535, n_3536, n_3538, n_3541, n_3543, n_3545, n_3546, n_3551;
wire n_3552, n_3557, n_3559, n_3560, n_3562, n_3565, n_3566, n_3567;
wire n_3569, n_3571, n_3573, n_3574, n_3575, n_3577, n_3579, n_3581;
wire n_3582, n_3585, n_3587, n_3588, n_3589, n_3590, n_3594, n_3597;
wire n_3599, n_3600, n_3601, n_3603, n_3604, n_3605, n_3609, n_3610;
wire n_3612, n_3613, n_3615, n_3616, n_3617, n_3619, n_3621, n_3622;
wire n_3624, n_3625, n_3626, n_3630, n_3631, n_3632, n_3633, n_3634;
wire n_3636, n_3639, n_3640, n_3642, n_3643, n_3644, n_3646, n_3650;
wire n_3651, n_3652, n_3653, n_3654, n_3656, n_3660, n_3663, n_3664;
wire n_3666, n_3667, n_3668, n_3669, n_3671, n_3672, n_3673, n_3676;
wire n_3677, n_3678, n_3679, n_3680, n_3682, n_3683, n_3686, n_3687;
wire n_3689, n_3691, n_3692, n_3694, n_3695, n_3696, n_3697, n_3698;
wire n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706;
wire n_3707, n_3710, n_3711, n_3714, n_3715, n_3716, n_3717, n_3718;
wire n_3721, n_3722, n_3723, n_3724, n_3725, n_3726, n_3728, n_3729;
wire n_3732, n_3735, n_3736, n_3739, n_3743, n_3746, n_3748, n_3749;
wire n_3753, n_3754, n_3755, n_3756, n_3758, n_3760, n_3764, n_3765;
wire n_3768, n_3769, n_3770, n_3771, n_3772, n_3774, n_3776, n_3777;
wire n_3778, n_3783, n_3785, n_3787, n_3791, n_3796, n_3797, n_3799;
wire n_3800, n_3802, n_3804, n_3805, n_3806, n_3807, n_3809, n_3811;
wire n_3812, n_3813, n_3814, n_3816, n_3817, n_3818, n_3820, n_3823;
wire n_3824, n_3825, n_3827, n_3829, n_3830, n_3831, n_3833, n_3834;
wire n_3835, n_3836, n_3837, n_3840, n_3841, n_3842, n_3844, n_3845;
wire n_3849, n_3851, n_3852, n_3858, n_3859, n_3861, n_3862, n_3865;
wire n_3867, n_3868, n_3869, n_3870, n_3871, n_3874, n_3883, n_3886;
wire n_3887, n_3888, n_3890, n_3891, n_3893, n_3895, n_3896, n_3900;
wire n_3903, n_3907, n_3909, n_3910, n_3911, n_3913, n_3915, n_3916;
wire n_3917, n_3918, n_3920, n_3921, n_3922, n_3923, n_3924, n_3925;
wire n_3926, n_3927, n_3929, n_3930, n_3931, n_3932, n_3933, n_3936;
wire n_3938, n_3940, n_3942, n_3943, n_3945, n_3948, n_3954, n_3955;
wire n_3959, n_3963, n_3964, n_3965, n_3966, n_3967, n_3972, n_3973;
wire n_3975, n_3979, n_3980, n_3981, n_3982, n_3984, n_3987, n_3989;
wire n_3990, n_3991, n_3992, n_3993, n_3997, n_3999, n_4000, n_4001;
wire n_4002, n_4003, n_4004, n_4006, n_4007, n_4009, n_4012, n_4014;
wire n_4015, n_4017, n_4018, n_4019, n_4021, n_4022, n_4023, n_4025;
wire n_4026, n_4027, n_4028, n_4030, n_4034, n_4036, n_4037, n_4038;
wire n_4039, n_4042, n_4043, n_4045, n_4046, n_4048, n_4049, n_4051;
wire n_4055, n_4060, n_4070, n_4071, n_4072, n_4073, n_4076, n_4077;
wire n_4079, n_4080, n_4082, n_4083, n_4084, n_4093, n_4094, n_4095;
wire n_4098, n_4099, n_4100, n_4102, n_4103, n_4104, n_4105, n_4106;
wire n_4107, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, n_4114;
wire n_4115, n_4117, n_4122, n_4123, n_4124, n_4126, n_4127, n_4128;
wire n_4129, n_4130, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137;
wire n_4138, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, n_4146;
wire n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4154, n_4155;
wire n_4157, n_4158, n_4159, n_4162, n_4163, n_4164, n_4165, n_4166;
wire n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174;
wire n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, n_4184;
wire n_4185, n_4187, n_4188, n_4189, n_4190, n_4191, n_4194, n_4195;
wire n_4196, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205;
wire n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, n_4213;
wire n_4214, n_4215, n_4216, n_4217, n_4219, n_4220, n_4221, n_4222;
wire n_4223, n_4224, n_4225, n_4227, n_4228, n_4229, n_4232, n_4233;
wire n_4234, n_4235, n_4238, n_4241, n_4242, n_4243, n_4245, n_4246;
wire n_4247, n_4248, n_4249, n_4250, n_4251, n_4253, n_4255, n_4256;
wire n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4264, n_4265;
wire n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273;
wire n_4274, n_4275, n_4276, n_4277, n_4279, n_4280, n_4281, n_4282;
wire n_4283, n_4285, n_4286, n_4289, n_4290, n_4291, n_4292, n_4293;
wire n_4295, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4304;
wire n_4307, n_4308, n_4309, n_4310, n_4312, n_4314, n_4315, n_4316;
wire n_4318, n_4319, n_4320, n_4321, n_4323, n_4325, n_4326, n_4327;
wire n_4328, n_4329, n_4330, n_4331, n_4332, n_4334, n_4335, n_4339;
wire n_4340, n_4342, n_4343, n_4344, n_4345, n_4346, n_4349, n_4350;
wire n_4353, n_4354, n_4356, n_4357, n_4358, n_4359, n_4363, n_4364;
wire n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372;
wire n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380;
wire n_4381, n_4382, n_4384, n_4385, n_4386, n_4388, n_4389, n_4390;
wire n_4391, n_4392, n_4393, n_4394, n_4396, n_4397, n_4400, n_4401;
wire n_4402, n_4403, n_4404, n_4405, n_4406, n_4407, n_4408, n_4410;
wire n_4412, n_4413, n_4414, n_4416, n_4417, n_4418, n_4419, n_4420;
wire n_4421, n_4422, n_4423, n_4424, n_4426, n_4427, n_4428, n_4429;
wire n_4430, n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439;
wire n_4441, n_4444, n_4447, n_4450, n_4451, n_4452, n_4453, n_4454;
wire n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462;
wire n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4470, n_4471;
wire n_4475, n_4476, n_4477, n_4478, n_4480, n_4481, n_4482, n_4483;
wire n_4484, n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492;
wire n_4493, n_4496, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504;
wire n_4505, n_4507, n_4509, n_4511, n_4512, n_4513, n_4514, n_4516;
wire n_4517, n_4518, n_4519, n_4520, n_4521, n_4522, n_4523, n_4525;
wire n_4526, n_4529, n_4533, n_4534, n_4536, n_4537, n_4539, n_4540;
wire n_4543, n_4544, n_4546, n_4547, n_4548, n_4549, n_4550, n_4552;
wire n_4553, n_4554, n_4555, n_4557, n_4558, n_4559, n_4561, n_4562;
wire n_4563, n_4565, n_4567, n_4568, n_4569, n_4570, n_4572, n_4573;
wire n_4575, n_4581, n_4582, n_4585, n_4586, n_4588, n_4590, n_4592;
wire n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600;
wire n_4601, n_4602, n_4604, n_4605, n_4606, n_4607, n_4611, n_4612;
wire n_4613, n_4614, n_4618, n_4619, n_4622, n_4625, n_4626, n_4627;
wire n_4632, n_4634, n_4635, n_4636, n_4638, n_4639, n_4640, n_4642;
wire n_4643, n_4644, n_4646, n_4647, n_4650, n_4653, n_4655, n_4658;
wire n_4659, n_4663, n_4664, n_4665, n_4666, n_4668, n_4669, n_4671;
wire n_4672, n_4675, n_4676, n_4678, n_4679, n_4681, n_4682, n_4684;
wire n_4685, n_4687, n_4688, n_4689, n_4691, n_4692, n_4694, n_4695;
wire n_4697, n_4699, n_4700, n_4701, n_4703, n_4704, n_4705, n_4706;
wire n_4708, n_4709, n_4712, n_4713, n_4714, n_4715, n_4718, n_4721;
wire n_4722, n_4724, n_4726, n_4727, n_4728, n_4730, n_4731, n_4732;
wire n_4736, n_4738, n_4739, n_4740, n_4741, n_4743, n_4744, n_4745;
wire n_4748, n_4750, n_4752, n_4753, n_4754, n_4755, n_4757, n_4758;
wire n_4760, n_4761, n_4762, n_4764, n_4767, n_4769, n_4770, n_4771;
wire n_4772, n_4773, n_4776, n_4777, n_4778, n_4782, n_4783, n_4784;
wire n_4786, n_4787, n_4788, n_4789, n_4792, n_4796, n_4798, n_4800;
wire n_4801, n_4802, n_4803, n_4804, n_4807, n_4811, n_4814, n_4819;
wire n_4820, n_4824, n_4825, n_4827, n_4828, n_4829, n_4830, n_4832;
wire n_4833, n_4835, n_4836, n_4837, n_4838, n_4839, n_4841, n_4842;
wire n_4844, n_4845, n_4846, n_4847, n_4848, n_4849, n_4850, n_4851;
wire n_4852, n_4853, n_4855, n_4856, n_4857, n_4859, n_4860, n_4861;
wire n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4872;
wire n_4875, n_4878, n_4881, n_4882, n_4883, n_4884, n_4886, n_4887;
wire n_4891, n_4893, n_4894, n_4897, n_4898, n_4899, n_4900, n_4901;
wire n_4902, n_4903, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909;
wire n_4911, n_4912, n_4914, n_4915, n_4916, n_4919, n_4920, n_4922;
wire n_4923, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930, n_4934;
wire n_4938, n_4939, n_4941, n_4943, n_4945, n_4947, n_4950, n_4951;
wire n_4955, n_4957, n_4960, n_4961, n_4962, n_4963, n_4965, n_4966;
wire n_4967, n_4969, n_4970, n_4973, n_4974, n_4976, n_4977, n_4978;
wire n_4979, n_4980, n_4981, n_4983, n_4984, n_4986, n_4987, n_4988;
wire n_4989, n_4993, n_4994, n_4997, n_5004, n_5005, n_5006, n_5007;
wire n_5008, n_5009, n_5010, n_5011, n_5012, n_5013, n_5014, n_5015;
wire n_5017, n_5018, n_5019, n_5020, n_5021, n_5024, n_5025, n_5030;
wire n_5032, n_5033, n_5034, n_5037, n_5038, n_5040, n_5042, n_5044;
wire n_5047, n_5048, n_5052, n_5053, n_5054, n_5058, n_5061, n_5064;
wire n_5066, n_5068, n_5072, n_5073, n_5074, n_5077, n_5079, n_5085;
wire n_5086, n_5091, n_5093, n_5096, n_5099, n_5101, n_5102, n_5103;
wire n_5104, n_5105, n_5108, n_5111, n_5112, n_5114, n_5117, n_5118;
wire n_5119, n_5120, n_5122, n_5123, n_5124, n_5126, n_5128, n_5129;
wire n_5130, n_5131, n_5134, n_5135, n_5136, n_5137, n_5138, n_5140;
wire n_5143, n_5144, n_5145, n_5146, n_5147, n_5148, n_5149, n_5150;
wire n_5151, n_5152, n_5153, n_5154, n_5155, n_5156, n_5159, n_5160;
wire n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167, n_5168;
wire n_5169, n_5170, n_5171, n_5172, n_5174, n_5175, n_5176, n_5177;
wire n_5178, n_5179, n_5180, n_5181, n_5182, n_5186, n_5187, n_5188;
wire n_5191, n_5193, n_5194, n_5196, n_5197, n_5198, n_5201, n_5202;
wire n_5203, n_5204, n_5205, n_5206, n_5208, n_5210, n_5211, n_5212;
wire n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219, n_5221;
wire n_5222, n_5224, n_5225, n_5226, n_5227, n_5228, n_5229, n_5230;
wire n_5231, n_5232, n_5233, n_5236, n_5237, n_5239, n_5240, n_5242;
wire n_5243, n_5247, n_5250, n_5251, n_5252, n_5253, n_5255, n_5257;
wire n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, n_5269;
wire n_5271, n_5272, n_5273, n_5276, n_5278, n_5280, n_5282, n_5285;
wire n_5288, n_5289, n_5290, n_5294, n_5295, n_5296, n_5297, n_5298;
wire n_5299, n_5301, n_5303, n_5304, n_5305, n_5306, n_5307, n_5309;
wire n_5310, n_5311, n_5312, n_5313, n_5315, n_5316, n_5317, n_5318;
wire n_5319, n_5322, n_5323, n_5324, n_5326, n_5327, n_5329, n_5330;
wire n_5331, n_5333, n_5334, n_5337, n_5340, n_5341, n_5343, n_5344;
wire n_5345, n_5346, n_5347, n_5349, n_5350, n_5352, n_5354, n_5355;
wire n_5357, n_5358, n_5360, n_5363, n_5365, n_5366, n_5367, n_5368;
wire n_5369, n_5370, n_5371, n_5373, n_5374, n_5375, n_5378, n_5380;
wire n_5381, n_5382, n_5383, n_5385, n_5386, n_5387, n_5388, n_5389;
wire n_5393, n_5394, n_5396, n_5397, n_5398, n_5399, n_5400, n_5402;
wire n_5403, n_5404, n_5405, n_5406, n_5408, n_5410, n_5411, n_5413;
wire n_5414, n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421;
wire n_5422, n_5423, n_5424, n_5425, n_5427, n_5428, n_5430, n_5435;
wire n_5436, n_5437, n_5439, n_5440, n_5441, n_5442, n_5443, n_5444;
wire n_5446, n_5447, n_5448, n_5450, n_5452, n_5453, n_5454, n_5455;
wire n_5456, n_5457, n_5458, n_5460, n_5462, n_5463, n_5467, n_5468;
wire n_5469, n_5470, n_5471, n_5472, n_5474, n_5475, n_5476, n_5477;
wire n_5481, n_5483, n_5484, n_5485, n_5487, n_5490, n_5491, n_5492;
wire n_5493, n_5494, n_5495, n_5496, n_5499, n_5502, n_5503, n_5504;
wire n_5505, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512, n_5513;
wire n_5514, n_5516, n_5517, n_5521, n_5522, n_5525, n_5527, n_5528;
wire n_5529, n_5530, n_5531, n_5532, n_5536, n_5537, n_5538, n_5540;
wire n_5541, n_5542, n_5543, n_5544, n_5545, n_5546, n_5547, n_5548;
wire n_5550, n_5552, n_5554, n_5555, n_5558, n_5559, n_5560, n_5563;
wire n_5564, n_5567, n_5568, n_5569, n_5571, n_5574, n_5575, n_5576;
wire n_5578, n_5580, n_5581, n_5585, n_5586, n_5588, n_5589, n_5590;
wire n_5591, n_5593, n_5594, n_5595, n_5599, n_5600, n_5601, n_5602;
wire n_5603, n_5605, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612;
wire n_5613, n_5614, n_5616, n_5617, n_5618, n_5619, n_5620, n_5621;
wire n_5625, n_5626, n_5628, n_5629, n_5630, n_5631, n_5634, n_5638;
wire n_5641, n_5642, n_5643, n_5644, n_5645, n_5646, n_5648, n_5650;
wire n_5652, n_5653, n_5654, n_5656, n_5657, n_5659, n_5660, n_5661;
wire n_5662, n_5663, n_5664, n_5665, n_5667, n_5668, n_5670, n_5671;
wire n_5674, n_5675, n_5677, n_5678, n_5680, n_5681, n_5682, n_5684;
wire n_5685, n_5686, n_5687, n_5688, n_5689, n_5690, n_5691, n_5692;
wire n_5693, n_5694, n_5697, n_5700, n_5704, n_5705, n_5706, n_5707;
wire n_5708, n_5709, n_5711, n_5712, n_5714, n_5715, n_5716, n_5717;
wire n_5719, n_5721, n_5722, n_5723, n_5724, n_5725, n_5726, n_5728;
wire n_5730, n_5731, n_5733, n_5734, n_5735, n_5736, n_5738, n_5740;
wire n_5741, n_5742, n_5743, n_5744, n_5745, n_5747, n_5749, n_5750;
wire n_5751, n_5752, n_5753, n_5755, n_5757, n_5759, n_5760, n_5761;
wire n_5762, n_5763, n_5764, n_5765, n_5766, n_5767, n_5768, n_5769;
wire n_5770, n_5771, n_5772, n_5774, n_5775, n_5776, n_5777, n_5778;
wire n_5779, n_5780, n_5781, n_5783, n_5784, n_5786, n_5787, n_5788;
wire n_5789, n_5791, n_5792, n_5795, n_5796, n_5798, n_5799, n_5800;
wire n_5801, n_5802, n_5803, n_5804, n_5805, n_5806, n_5807, n_5808;
wire n_5809, n_5810, n_5812, n_5813, n_5816, n_5817, n_5818, n_5819;
wire n_5820, n_5822, n_5823, n_5826, n_5827, n_5828, n_5829, n_5832;
wire n_5833, n_5834, n_5835, n_5837, n_5838, n_5839, n_5841, n_5842;
wire n_5843, n_5845, n_5846, n_5848, n_5850, n_5851, n_5852, n_5853;
wire n_5854, n_5855, n_5856, n_5857, n_5859, n_5860, n_5861, n_5862;
wire n_5864, n_5866, n_5867, n_5868, n_5870, n_5871, n_5872, n_5874;
wire n_5875, n_5878, n_5881, n_5882, n_5884, n_5885, n_5886, n_5887;
wire n_5888, n_5891, n_5892, n_5893, n_5894, n_5895, n_5896, n_5897;
wire n_5906, n_5907, n_5910, n_5911, n_5912, n_5913, n_5914, n_5915;
wire n_5917, n_5918, n_5921, n_5922, n_5923, n_5924, n_5925, n_5926;
wire n_5928, n_5929, n_5930, n_5931, n_5932, n_5934, n_5935, n_5936;
wire n_5937, n_5938, n_5939, n_5941, n_5942, n_5943, n_5944, n_5945;
wire n_5946, n_5947, n_5949, n_5950, n_5951, n_5953, n_5955, n_5956;
wire n_5957, n_5958, n_5960, n_5961, n_5963, n_5966, n_5967, n_5968;
wire n_5969, n_5970, n_5971, n_5972, n_5973, n_5974, n_5975, n_5976;
wire n_5978, n_5979, n_5981, n_5982, n_5983, n_5984, n_5985, n_5986;
wire n_5988, n_5989, n_5990, n_5991, n_5992, n_5994, n_5996, n_5997;
wire n_5998, n_6000, n_6001, n_6003, n_6004, n_6005, n_6006, n_6007;
wire n_6008, n_6009, n_6010, n_6011, n_6012, n_6015, n_6018, n_6020;
wire n_6021, n_6022, n_6023, n_6024, n_6025, n_6026, n_6027, n_6028;
wire n_6031, n_6032, n_6033, n_6034, n_6035, n_6036, n_6038, n_6040;
wire n_6041, n_6042, n_6043, n_6044, n_6045, n_6046, n_6047, n_6048;
wire n_6050, n_6051, n_6052, n_6053, n_6055, n_6056, n_6057, n_6058;
wire n_6059, n_6060, n_6062, n_6063, n_6064, n_6065, n_6066, n_6067;
wire n_6068, n_6069, n_6072, n_6074, n_6076, n_6077, n_6078, n_6079;
wire n_6080, n_6081, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087;
wire n_6088, n_6092, n_6093, n_6094, n_6096, n_6097, n_6099, n_6102;
wire n_6104, n_6105, n_6106, n_6107, n_6108, n_6111, n_6113, n_6114;
wire n_6117, n_6119, n_6121, n_6122, n_6126, n_6127, n_6128, n_6131;
wire n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6140;
wire n_6141, n_6142, n_6144, n_6145, n_6148, n_6149, n_6151, n_6153;
wire n_6154, n_6155, n_6158, n_6162, n_6164, n_6166, n_6167, n_6169;
wire n_6170, n_6171, n_6173, n_6179, n_6181, n_6183, n_6184, n_6185;
wire n_6188, n_6189, n_6191, n_6194, n_6197, n_6198, n_6200, n_6202;
wire n_6204, n_6205, n_6206, n_6207, n_6209, n_6210, n_6211, n_6212;
wire n_6213, n_6216, n_6217, n_6218, n_6219, n_6220, n_6222, n_6223;
wire n_6226, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232, n_6233;
wire n_6234, n_6235, n_6237, n_6238, n_6239, n_6243, n_6244, n_6245;
wire n_6246, n_6247, n_6248, n_6249, n_6250, n_6252, n_6254, n_6255;
wire n_6256, n_6258, n_6260, n_6261, n_6265, n_6266, n_6268, n_6269;
wire n_6270, n_6274, n_6275, n_6276, n_6277, n_6278, n_6279, n_6280;
wire n_6281, n_6282, n_6283, n_6285, n_6286, n_6287, n_6289, n_6291;
wire n_6293, n_6294, n_6295, n_6298, n_6301, n_6302, n_6303, n_6304;
wire n_6306, n_6308, n_6310, n_6312, n_6313, n_6314, n_6315, n_6319;
wire n_6325, n_6327, n_6328, n_6329, n_6330, n_6332, n_6333, n_6334;
wire n_6335, n_6336, n_6337, n_6338, n_6339, n_6341, n_6342, n_6344;
wire n_6346, n_6347, n_6350, n_6352, n_6353, n_6354, n_6355, n_6356;
wire n_6358, n_6361, n_6363, n_6364, n_6365, n_6366, n_6368, n_6369;
wire n_6370, n_6371, n_6372, n_6373, n_6374, n_6375, n_6376, n_6377;
wire n_6384, n_6386, n_6390, n_6391, n_6392, n_6393, n_6394, n_6396;
wire n_6397, n_6398, n_6399, n_6400, n_6401, n_6402, n_6404, n_6405;
wire n_6406, n_6407, n_6408, n_6409, n_6413, n_6414, n_6415, n_6416;
wire n_6417, n_6418, n_6419, n_6420, n_6421, n_6422, n_6423, n_6425;
wire n_6426, n_6427, n_6428, n_6429, n_6431, n_6432, n_6434, n_6435;
wire n_6436, n_6437, n_6438, n_6439, n_6440, n_6441, n_6442, n_6443;
wire n_6444, n_6445, n_6446, n_6447, n_6448, n_6449, n_6450, n_6451;
wire n_6452, n_6453, n_6457, n_6458, n_6459, n_6461, n_6462, n_6463;
wire n_6464, n_6468, n_6469, n_6470, n_6475, n_6476, n_6477, n_6478;
wire n_6479, n_6480, n_6482, n_6486, n_6488, n_6489, n_6490, n_6491;
wire n_6492, n_6493, n_6494, n_6495, n_6496, n_6497, n_6498, n_6499;
wire n_6500, n_6505, n_6510, n_6511, n_6512, n_6515, n_6516, n_6521;
wire n_6522, n_6523, n_6527, n_6528, n_6529, n_6530, n_6531, n_6532;
wire n_6533, n_6534, n_6535, n_6536, n_6537, n_6539, n_6540, n_6542;
wire n_6544, n_6545, n_6546, n_6547, n_6548, n_6549, n_6551, n_6553;
wire n_6554, n_6555, n_6556, n_6557, n_6558, n_6563, n_6564, n_6565;
wire n_6567, n_6569, n_6571, n_6573, n_6574, n_6575, n_6577, n_6578;
wire n_6579, n_6580, n_6581, n_6582, n_6583, n_6584, n_6586, n_6587;
wire n_6588, n_6589, n_6590, n_6592, n_6593, n_6594, n_6595, n_6597;
wire n_6598, n_6599, n_6600, n_6601, n_6603, n_6604, n_6606, n_6607;
wire n_6609, n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616;
wire n_6618, n_6619, n_6620, n_6621, n_6623, n_6624, n_6627, n_6633;
wire n_6634, n_6635, n_6636, n_6637, n_6639, n_6640, n_6641, n_6644;
wire n_6645, n_6647, n_6648, n_6652, n_6653, n_6654, n_6655, n_6656;
wire n_6657, n_6659, n_6660, n_6661, n_6665, n_6669, n_6670, n_6671;
wire n_6672, n_6673, n_6674, n_6676, n_6677, n_6678, n_6679, n_6680;
wire n_6681, n_6684, n_6685, n_6687, n_6688, n_6689, n_6692, n_6694;
wire n_6696, n_6697, n_6698, n_6699, n_6700, n_6701, n_6703, n_6705;
wire n_6706, n_6709, n_6711, n_6712, n_6713, n_6714, n_6715, n_6716;
wire n_6717, n_6720, n_6721, n_6723, n_6724, n_6725, n_6727, n_6728;
wire n_6730, n_6731, n_6732, n_6733, n_6734, n_6735, n_6738, n_6739;
wire n_6740, n_6742, n_6743, n_6744, n_6745, n_6746, n_6747, n_6748;
wire n_6749, n_6750, n_6751, n_6753, n_6754, n_6755, n_6756, n_6758;
wire n_6759, n_6760, n_6762, n_6764, n_6766, n_6767, n_6768, n_6769;
wire n_6772, n_6773, n_6774, n_6775, n_6779, n_6780, n_6783, n_6784;
wire n_6785, n_6790, n_6791, n_6794, n_6797, n_6801, n_6802, n_6803;
wire n_6804, n_6805, n_6806, n_6808, n_6809, n_6810, n_6811, n_6812;
wire n_6813, n_6814, n_6815, n_6816, n_6817, n_6818, n_6819, n_6821;
wire n_6822, n_6823, n_6824, n_6825, n_6827, n_6828, n_6829, n_6830;
wire n_6831, n_6833, n_6834, n_6835, n_6836, n_6837, n_6838, n_6840;
wire n_6841, n_6842, n_6843, n_6844, n_6846, n_6847, n_6848, n_6849;
wire n_6850, n_6851, n_6853, n_6855, n_6856, n_6857, n_6858, n_6861;
wire n_6862, n_6863, n_6865, n_6866, n_6868, n_6870, n_6871, n_6872;
wire n_6873, n_6874, n_6875, n_6877, n_6878, n_6879, n_6880, n_6882;
wire n_6884, n_6885, n_6887, n_6888, n_6889, n_6890, n_6891, n_6892;
wire n_6895, n_6896, n_6897, n_6898, n_6900, n_6901, n_6902, n_6903;
wire n_6904, n_6905, n_6906, n_6907, n_6908, n_6910, n_6911, n_6913;
wire n_6914, n_6915, n_6916, n_6918, n_6919, n_6920, n_6921, n_6922;
wire n_6923, n_6924, n_6926, n_6927, n_6928, n_6929, n_6930, n_6931;
wire n_6933, n_6934, n_6935, n_6937, n_6938, n_6939, n_6940, n_6941;
wire n_6942, n_6943, n_6944, n_6945, n_6946, n_6947, n_6948, n_6950;
wire n_6951, n_6952, n_6953, n_6955, n_6956, n_6957, n_6958, n_6960;
wire n_6961, n_6962, n_6963, n_6964, n_6965, n_6966, n_6967, n_6968;
wire n_6969, n_6970, n_6971, n_6972, n_6974, n_6976, n_6977, n_6978;
wire n_6979, n_6980, n_6982, n_6983, n_6985, n_6986, n_6987, n_6988;
wire n_6989, n_6990, n_6991, n_6992, n_6993, n_6994, n_6995, n_6996;
wire n_6997, n_6999, n_7000, n_7002, n_7003, n_7004, n_7005, n_7006;
wire n_7008, n_7011, n_7013, n_7014, n_7015, n_7016, n_7018, n_7020;
wire n_7022, n_7023, n_7025, n_7026, n_7027, n_7028, n_7030, n_7031;
wire n_7032, n_7033, n_7035, n_7036, n_7038, n_7039, n_7040, n_7041;
wire n_7042, n_7043, n_7044, n_7046, n_7047, n_7048, n_7050, n_7051;
wire n_7052, n_7053, n_7056, n_7058, n_7059, n_7061, n_7062, n_7063;
wire n_7064, n_7065, n_7066, n_7067, n_7068, n_7069, n_7071, n_7072;
wire n_7073, n_7075, n_7076, n_7077, n_7079, n_7081, n_7082, n_7083;
wire n_7084, n_7085, n_7086, n_7088, n_7089, n_7090, n_7091, n_7093;
wire n_7095, n_7096, n_7098, n_7099, n_7100, n_7101, n_7102, n_7104;
wire n_7106, n_7108, n_7109, n_7110, n_7112, n_7113, n_7114, n_7115;
wire n_7116, n_7117, n_7119, n_7120, n_7121, n_7123, n_7124, n_7125;
wire n_7126, n_7127, n_7128, n_7130, n_7131, n_7132, n_7136, n_7137;
wire n_7138, n_7139, n_7140, n_7141, n_7142, n_7143, n_7144, n_7145;
wire n_7146, n_7147, n_7152, n_7153, n_7155, n_7157, n_7158, n_7159;
wire n_7160, n_7161, n_7162, n_7163, n_7164, n_7165, n_7166, n_7167;
wire n_7168, n_7169, n_7170, n_7171, n_7172, n_7173, n_7175, n_7176;
wire n_7177, n_7178, n_7180, n_7181, n_7182, n_7183, n_7184, n_7185;
wire n_7187, n_7188, n_7190, n_7191, n_7192, n_7193, n_7194, n_7195;
wire n_7196, n_7197, n_7198, n_7199, n_7201, n_7202, n_7203, n_7204;
wire n_7205, n_7206, n_7207, n_7208, n_7209, n_7210, n_7211, n_7212;
wire n_7213, n_7214, n_7215, n_7216, n_7217, n_7218, n_7219, n_7220;
wire n_7221, n_7222, n_7226, n_7227, n_7228, n_7230, n_7232, n_7233;
wire n_7235, n_7237, n_7238, n_7239, n_7240, n_7241, n_7242, n_7243;
wire n_7244, n_7245, n_7247, n_7249, n_7250, n_7252, n_7253, n_7255;
wire n_7256, n_7257, n_7258, n_7259, n_7260, n_7262, n_7263, n_7264;
wire n_7266, n_7267, n_7269, n_7272, n_7274, n_7275, n_7276, n_7278;
wire n_7282, n_7283, n_7286, n_7288, n_7290, n_7291, n_7292, n_7293;
wire n_7294, n_7296, n_7297, n_7298, n_7299, n_7301, n_7302, n_7303;
wire n_7305, n_7306, n_7307, n_7308, n_7309, n_7310, n_7312, n_7315;
wire n_7316, n_7317, n_7318, n_7319, n_7320, n_7321, n_7322, n_7324;
wire n_7325, n_7326, n_7327, n_7328, n_7329, n_7330, n_7331, n_7332;
wire n_7333, n_7334, n_7336, n_7337, n_7339, n_7340, n_7343, n_7344;
wire n_7345, n_7346, n_7347, n_7348, n_7349, n_7350, n_7351, n_7352;
wire n_7353, n_7354, n_7355, n_7357, n_7358, n_7359, n_7362, n_7363;
wire n_7365, n_7366, n_7367, n_7368, n_7369, n_7370, n_7371, n_7372;
wire n_7373, n_7376, n_7377, n_7378, n_7380, n_7381, n_7382, n_7383;
wire n_7384, n_7385, n_7386, n_7388, n_7389, n_7390, n_7391, n_7393;
wire n_7394, n_7395, n_7397, n_7399, n_7403, n_7404, n_7406, n_7407;
wire n_7408, n_7409, n_7410, n_7411, n_7412, n_7414, n_7415, n_7416;
wire n_7417, n_7418, n_7419, n_7420, n_7421, n_7422, n_7424, n_7427;
wire n_7428, n_7429, n_7430, n_7432, n_7433, n_7434, n_7436, n_7437;
wire n_7438, n_7440, n_7441, n_7443, n_7444, n_7446, n_7447, n_7448;
wire n_7450, n_7452, n_7453, n_7454, n_7455, n_7456, n_7457, n_7458;
wire n_7459, n_7461, n_7463, n_7464, n_7466, n_7467, n_7469, n_7470;
wire n_7471, n_7472, n_7473, n_7476, n_7477, n_7478, n_7479, n_7480;
wire n_7481, n_7482, n_7483, n_7485, n_7486, n_7487, n_7488, n_7489;
wire n_7490, n_7492, n_7494, n_7495, n_7496, n_7497, n_7498, n_7499;
wire n_7503, n_7504, n_7505, n_7506, n_7507, n_7509, n_7511, n_7512;
wire n_7513, n_7517, n_7518, n_7519, n_7520, n_7521, n_7522, n_7523;
wire n_7524, n_7526, n_7527, n_7528, n_7529, n_7531, n_7532, n_7534;
wire n_7535, n_7536, n_7537, n_7540, n_7541, n_7542, n_7543, n_7544;
wire n_7545, n_7546, n_7547, n_7548, n_7549, n_7550, n_7551, n_7552;
wire n_7553, n_7554, n_7555, n_7556, n_7557, n_7558, n_7559, n_7563;
wire n_7564, n_7565, n_7566, n_7567, n_7568, n_7569, n_7572, n_7573;
wire n_7574, n_7576, n_7577, n_7578, n_7579, n_7583, n_7584, n_7585;
wire n_7586, n_7590, n_7591, n_7592, n_7593, n_7594, n_7595, n_7596;
wire n_7597, n_7598, n_7599, n_7600, n_7601, n_7602, n_7603, n_7605;
wire n_7606, n_7607, n_7608, n_7609, n_7610, n_7614, n_7615, n_7616;
wire n_7617, n_7618, n_7619, n_7620, n_7623, n_7624, n_7625, n_7626;
wire n_7628, n_7629, n_7630, n_7631, n_7632, n_7634, n_7635, n_7636;
wire n_7637, n_7639, n_7640, n_7641, n_7642, n_7644, n_7645, n_7649;
wire n_7650, n_7653, n_7656, n_7658, n_7659, n_7661, n_7662, n_7663;
wire n_7664, n_7665, n_7666, n_7667, n_7668, n_7671, n_7672, n_7673;
wire n_7674, n_7675, n_7676, n_7678, n_7679, n_7680, n_7682, n_7683;
wire n_7685, n_7686, n_7687, n_7688, n_7690, n_7694, n_7696, n_7698;
wire n_7700, n_7701, n_7702, n_7703, n_7705, n_7708, n_7709, n_7710;
wire n_7711, n_7712, n_7713, n_7714, n_7717, n_7718, n_7719, n_7721;
wire n_7722, n_7723, n_7724, n_7725, n_7726, n_7727, n_7728, n_7730;
wire n_7732, n_7733, n_7734, n_7739, n_7741, n_7742, n_7744, n_7745;
wire n_7746, n_7748, n_7753, n_7755, n_7756, n_7757, n_7758, n_7759;
wire n_7763, n_7767, n_7769, n_7770, n_7771, n_7775, n_7776, n_7777;
wire n_7778, n_7782, n_7783, n_7784, n_7785, n_7786, n_7787, n_7789;
wire n_7792, n_7794, n_7795, n_7796, n_7797, n_7798, n_7799, n_7800;
wire n_7802, n_7803, n_7804, n_7805, n_7806, n_7807, n_7808, n_7810;
wire n_7811, n_7812, n_7813, n_7814, n_7815, n_7816, n_7818, n_7820;
wire n_7821, n_7822, n_7823, n_7824, n_7826, n_7828, n_7830, n_7831;
wire n_7832, n_7833, n_7834, n_7835, n_7837, n_7840, n_7841, n_7843;
wire n_7844, n_7845, n_7846, n_7847, n_7849, n_7851, n_7853, n_7854;
wire n_7858, n_7859, n_7860, n_7862, n_7864, n_7865, n_7867, n_7868;
wire n_7870, n_7871, n_7874, n_7875, n_7876, n_7877, n_7878, n_7879;
wire n_7881, n_7882, n_7883, n_7885, n_7887, n_7888, n_7889, n_7890;
wire n_7892, n_7893, n_7894, n_7895, n_7898, n_7899, n_7900, n_7902;
wire n_7903, n_7904, n_7905, n_7906, n_7910, n_7911, n_7912, n_7913;
wire n_7917, n_7919, n_7921, n_7923, n_7925, n_7927, n_7928, n_7929;
wire n_7930, n_7931, n_7932, n_7933, n_7934, n_7935, n_7936, n_7937;
wire n_7938, n_7939, n_7940, n_7942, n_7943, n_7944, n_7945, n_7946;
wire n_7947, n_7948, n_7950, n_7952, n_7953, n_7954, n_7955, n_7956;
wire n_7957, n_7959, n_7961, n_7963, n_7964, n_7965, n_7966, n_7967;
wire n_7968, n_7969, n_7971, n_7973, n_7974, n_7975, n_7976, n_7978;
wire n_7979, n_7981, n_7982, n_7983, n_7984, n_7985, n_7992, n_7995;
wire n_7996, n_7997, n_7999, n_8000, n_8001, n_8003, n_8006, n_8007;
wire n_8008, n_8009, n_8010, n_8012, n_8013, n_8014, n_8015, n_8016;
wire n_8017, n_8018, n_8019, n_8020, n_8021, n_8022, n_8023, n_8024;
wire n_8025, n_8026, n_8029, n_8030, n_8034, n_8035, n_8036, n_8037;
wire n_8038, n_8039, n_8047, n_8048, n_8049, n_8052, n_8059, n_8062;
wire n_8063, n_8064, n_8068, n_8069, n_8070, n_8071, n_8073, n_8075;
wire n_8076, n_8077, n_8078, n_8079, n_8080, n_8083, n_8085, n_8086;
wire n_8088, n_8089, n_8090, n_8091, n_8092, n_8093, n_8094, n_8095;
wire n_8096, n_8097, n_8098, n_8099, n_8100, n_8101, n_8103, n_8104;
wire n_8105, n_8106, n_8107, n_8108, n_8109, n_8110, n_8111, n_8112;
wire n_8113, n_8114, n_8115, n_8116, n_8117, n_8118, n_8119, n_8120;
wire n_8121, n_8123, n_8124, n_8125, n_8126, n_8127, n_8128, n_8129;
wire n_8130, n_8132, n_8135, n_8137, n_8138, n_8139, n_8140, n_8141;
wire n_8142, n_8143, n_8144, n_8145, n_8146, n_8148, n_8149, n_8152;
wire n_8154, n_8155, n_8157, n_8159, n_8161, n_8163, n_8164, n_8165;
wire n_8166, n_8167, n_8169, n_8170, n_8171, n_8172, n_8173, n_8174;
wire n_8176, n_8177, n_8181, n_8183, n_8184, n_8185, n_8186, n_8187;
wire n_8188, n_8189, n_8191, n_8192, n_8193, n_8194, n_8195, n_8197;
wire n_8198, n_8199, n_8201, n_8202, n_8203, n_8205, n_8206, n_8209;
wire n_8210, n_8212, n_8213, n_8215, n_8216, n_8217, n_8218, n_8219;
wire n_8221, n_8222, n_8223, n_8224, n_8227, n_8228, n_8229, n_8231;
wire n_8233, n_8234, n_8235, n_8239, n_8240, n_8243, n_8244, n_8245;
wire n_8246, n_8247, n_8249, n_8250, n_8251, n_8253, n_8254, n_8255;
wire n_8256, n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8264;
wire n_8265, n_8266, n_8267, n_8268, n_8269, n_8272, n_8273, n_8274;
wire n_8275, n_8276, n_8277, n_8282, n_8283, n_8284, n_8285, n_8286;
wire n_8287, n_8288, n_8289, n_8290, n_8291, n_8292, n_8293, n_8294;
wire n_8295, n_8296, n_8297, n_8298, n_8299, n_8300, n_8301, n_8302;
wire n_8306, n_8308, n_8309, n_8314, n_8317, n_8318, n_8319, n_8320;
wire n_8321, n_8322, n_8323, n_8324, n_8325, n_8326, n_8328, n_8329;
wire n_8330, n_8331, n_8333, n_8334, n_8335, n_8336, n_8337, n_8338;
wire n_8339, n_8341, n_8342, n_8343, n_8344, n_8345, n_8346, n_8347;
wire n_8348, n_8349, n_8351, n_8353, n_8354, n_8355, n_8356, n_8357;
wire n_8358, n_8360, n_8361, n_8362, n_8363, n_8364, n_8366, n_8367;
wire n_8368, n_8370, n_8371, n_8375, n_8377, n_8378, n_8379, n_8380;
wire n_8381, n_8382, n_8383, n_8384, n_8386, n_8388, n_8389, n_8390;
wire n_8391, n_8392, n_8393, n_8395, n_8396, n_8397, n_8398, n_8399;
wire n_8402, n_8403, n_8404, n_8405, n_8406, n_8408, n_8411, n_8412;
wire n_8414, n_8415, n_8417, n_8418, n_8419, n_8420, n_8421, n_8422;
wire n_8423, n_8424, n_8425, n_8426, n_8427, n_8428, n_8429, n_8431;
wire n_8433, n_8435, n_8436, n_8437, n_8438, n_8439, n_8441, n_8442;
wire n_8443, n_8444, n_8445, n_8447, n_8448, n_8449, n_8451, n_8452;
wire n_8454, n_8456, n_8458, n_8459, n_8460, n_8462, n_8464, n_8465;
wire n_8466, n_8467, n_8469, n_8470, n_8471, n_8472, n_8473, n_8477;
wire n_8478, n_8480, n_8481, n_8482, n_8483, n_8484, n_8486, n_8487;
wire n_8488, n_8489, n_8490, n_8491, n_8492, n_8493, n_8495, n_8496;
wire n_8497, n_8498, n_8499, n_8500, n_8502, n_8503, n_8504, n_8505;
wire n_8507, n_8508, n_8510, n_8511, n_8513, n_8514, n_8515, n_8516;
wire n_8518, n_8519, n_8520, n_8521, n_8522, n_8523, n_8524, n_8525;
wire n_8526, n_8527, n_8529, n_8532, n_8534, n_8535, n_8536, n_8537;
wire n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544, n_8545;
wire n_8546, n_8548, n_8549, n_8550, n_8552, n_8553, n_8554, n_8555;
wire n_8556, n_8557, n_8559, n_8560, n_8561, n_8564, n_8565, n_8566;
wire n_8567, n_8568, n_8569, n_8570, n_8571, n_8572, n_8573, n_8576;
wire n_8580, n_8581, n_8583, n_8584, n_8585, n_8586, n_8587, n_8588;
wire n_8590, n_8592, n_8593, n_8595, n_8597, n_8598, n_8600, n_8603;
wire n_8604, n_8605, n_8607, n_8608, n_8610, n_8611, n_8612, n_8613;
wire n_8614, n_8615, n_8619, n_8620, n_8621, n_8627, n_8628, n_8629;
wire n_8632, n_8633, n_8634, n_8635, n_8636, n_8637, n_8638, n_8640;
wire n_8641, n_8642, n_8643, n_8644, n_8645, n_8648, n_8649, n_8650;
wire n_8652, n_8654, n_8655, n_8657, n_8658, n_8660, n_8661, n_8662;
wire n_8663, n_8664, n_8665, n_8666, n_8667, n_8668, n_8669, n_8670;
wire n_8671, n_8672, n_8673, n_8674, n_8675, n_8678, n_8679, n_8680;
wire n_8681, n_8682, n_8683, n_8684, n_8685, n_8686, n_8687, n_8688;
wire n_8690, n_8691, n_8695, n_8696, n_8699, n_8700, n_8701, n_8702;
wire n_8703, n_8704, n_8706, n_8707, n_8708, n_8709, n_8711, n_8712;
wire n_8713, n_8714, n_8715, n_8719, n_8720, n_8721, n_8723, n_8724;
wire n_8725, n_8726, n_8729, n_8730, n_8734, n_8735, n_8736, n_8737;
wire n_8742, n_8743, n_8744, n_8745, n_8746, n_8747, n_8748, n_8749;
wire n_8755, n_8756, n_8757, n_8759, n_8760, n_8763, n_8768, n_8769;
wire n_8770, n_8772, n_8774, n_8775, n_8777, n_8778, n_8779, n_8780;
wire n_8784, n_8788, n_8791, n_8793, n_8794, n_8795, n_8797, n_8799;
wire n_8800, n_8801, n_8803, n_8805, n_8806, n_8808, n_8809, n_8810;
wire n_8811, n_8812, n_8813, n_8814, n_8815, n_8816, n_8817, n_8818;
wire n_8820, n_8821, n_8822, n_8823, n_8824, n_8827, n_8828, n_8830;
wire n_8833, n_8834, n_8835, n_8837, n_8839, n_8840, n_8842, n_8844;
wire n_8845, n_8846, n_8847, n_8848, n_8849, n_8850, n_8851, n_8852;
wire n_8855, n_8856, n_8857, n_8858, n_8859, n_8860, n_8861, n_8862;
wire n_8863, n_8865, n_8866, n_8867, n_8868, n_8870, n_8871, n_8872;
wire n_8874, n_8875, n_8876, n_8877, n_8878, n_8879, n_8880, n_8881;
wire n_8883, n_8884, n_8885, n_8887, n_8888, n_8889, n_8890, n_8891;
wire n_8892, n_8894, n_8895, n_8896, n_8897, n_8898, n_8900, n_8901;
wire n_8902, n_8903, n_8904, n_8905, n_8907, n_8908, n_8909, n_8910;
wire n_8911, n_8912, n_8913, n_8914, n_8915, n_8916, n_8917, n_8918;
wire n_8921, n_8922, n_8924, n_8925, n_8927, n_8928, n_8929, n_8931;
wire n_8932, n_8933, n_8934, n_8935, n_8936, n_8937, n_8939, n_8940;
wire n_8941, n_8942, n_8943, n_8944, n_8945, n_8946, n_8948, n_8951;
wire n_8952, n_8954, n_8956, n_8958, n_8959, n_8962, n_8963, n_8966;
wire n_8968, n_8969, n_8970, n_8971, n_8972, n_8973, n_8974, n_8976;
wire n_8977, n_8978, n_8979, n_8980, n_8983, n_8984, n_8986, n_8990;
wire n_8992, n_8995, n_8996, n_8997, n_9000, n_9003, n_9004, n_9005;
wire n_9006, n_9008, n_9013, n_9015, n_9016, n_9017, n_9018, n_9020;
wire n_9021, n_9023, n_9024, n_9026, n_9028, n_9029, n_9032, n_9033;
wire n_9034, n_9035, n_9037, n_9038, n_9039, n_9040, n_9041, n_9043;
wire n_9044, n_9045, n_9046, n_9047, n_9048, n_9050, n_9051, n_9053;
wire n_9054, n_9056, n_9057, n_9058, n_9060, n_9061, n_9064, n_9066;
wire n_9068, n_9069, n_9071, n_9073, n_9074, n_9075, n_9077, n_9078;
wire n_9079, n_9081, n_9082, n_9084, n_9085, n_9088, n_9089, n_9091;
wire n_9092, n_9093, n_9094, n_9095, n_9096, n_9098, n_9099, n_9101;
wire n_9103, n_9105, n_9106, n_9107, n_9108, n_9111, n_9112, n_9113;
wire n_9114, n_9115, n_9116, n_9118, n_9123, n_9124, n_9125, n_9126;
wire n_9127, n_9129, n_9130, n_9132, n_9133, n_9134, n_9135, n_9136;
wire n_9138, n_9139, n_9140, n_9142, n_9143, n_9144, n_9145, n_9146;
wire n_9149, n_9152, n_9155, n_9156, n_9157, n_9158, n_9159, n_9160;
wire n_9161, n_9162, n_9163, n_9164, n_9165, n_9166, n_9167, n_9169;
wire n_9170, n_9171, n_9172, n_9173, n_9174, n_9175, n_9176, n_9179;
wire n_9180, n_9181, n_9182, n_9183, n_9184, n_9186, n_9187, n_9188;
wire n_9189, n_9190, n_9191, n_9192, n_9193, n_9195, n_9196, n_9197;
wire n_9198, n_9199, n_9200, n_9201, n_9202, n_9203, n_9204, n_9205;
wire n_9207, n_9208, n_9209, n_9210, n_9211, n_9212, n_9213, n_9214;
wire n_9215, n_9217, n_9219, n_9220, n_9221, n_9222, n_9225, n_9226;
wire n_9227, n_9228, n_9229, n_9230, n_9232, n_9233, n_9234, n_9235;
wire n_9236, n_9237, n_9238, n_9241, n_9242, n_9243, n_9244, n_9245;
wire n_9246, n_9247, n_9249, n_9250, n_9251, n_9253, n_9254, n_9255;
wire n_9257, n_9258, n_9260, n_9261, n_9262, n_9264, n_9265, n_9268;
wire n_9269, n_9272, n_9273, n_9274, n_9276, n_9278, n_9279, n_9281;
wire n_9282, n_9283, n_9284, n_9285, n_9286, n_9288, n_9289, n_9290;
wire n_9291, n_9293, n_9294, n_9295, n_9296, n_9297, n_9298, n_9299;
wire n_9300, n_9301, n_9303, n_9304, n_9305, n_9306, n_9307, n_9308;
wire n_9309, n_9310, n_9311, n_9312, n_9313, n_9314, n_9315, n_9316;
wire n_9317, n_9318, n_9319, n_9320, n_9321, n_9322, n_9323, n_9325;
wire n_9326, n_9327, n_9328, n_9329, n_9330, n_9331, n_9332, n_9333;
wire n_9334, n_9335, n_9336, n_9337, n_9338, n_9340, n_9341, n_9342;
wire n_9343, n_9344, n_9345, n_9346, n_9348, n_9349, n_9350, n_9351;
wire n_9352, n_9353, n_9354, n_9355, n_9356, n_9357, n_9361, n_9362;
wire n_9363, n_9364, n_9365, n_9366, n_9368, n_9369, n_9370, n_9371;
wire n_9372, n_9374, n_9375, n_9377, n_9380, n_9382, n_9384, n_9385;
wire n_9386, n_9387, n_9388, n_9389, n_9390, n_9392, n_9394, n_9395;
wire n_9397, n_9399, n_9402, n_9403, n_9404, n_9405, n_9406, n_9407;
wire n_9409, n_9410, n_9414, n_9415, n_9416, n_9417, n_9418, n_9419;
wire n_9420, n_9424, n_9425, n_9426, n_9428, n_9429, n_9430, n_9431;
wire n_9433, n_9435, n_9436, n_9437, n_9439, n_9440, n_9442, n_9444;
wire n_9445, n_9446, n_9449, n_9450, n_9451, n_9456, n_9457, n_9459;
wire n_9460, n_9462, n_9463, n_9464, n_9465, n_9466, n_9467, n_9469;
wire n_9471, n_9472, n_9473, n_9474, n_9475, n_9477, n_9479, n_9480;
wire n_9481, n_9482, n_9483, n_9486, n_9487, n_9489, n_9491, n_9495;
wire n_9497, n_9500, n_9501, n_9502, n_9504, n_9505, n_9508, n_9509;
wire n_9510, n_9511, n_9513, n_9514, n_9515, n_9522, n_9523, n_9524;
wire n_9525, n_9526, n_9527, n_9528, n_9529, n_9530, n_9531, n_9532;
wire n_9534, n_9537, n_9538, n_9539, n_9541, n_9543, n_9545, n_9547;
wire n_9548, n_9549, n_9550, n_9552, n_9553, n_9555, n_9556, n_9557;
wire n_9558, n_9559, n_9560, n_9561, n_9562, n_9564, n_9565, n_9566;
wire n_9567, n_9568, n_9569, n_9572, n_9573, n_9574, n_9575, n_9576;
wire n_9577, n_9579, n_9580, n_9581, n_9582, n_9584, n_9585, n_9586;
wire n_9587, n_9588, n_9590, n_9592, n_9593, n_9594, n_9595, n_9596;
wire n_9597, n_9599, n_9601, n_9602, n_9604, n_9605, n_9607, n_9609;
wire n_9610, n_9612, n_9614, n_9615, n_9617, n_9619, n_9621, n_9624;
wire n_9625, n_9626, n_9627, n_9628, n_9629, n_9632, n_9635, n_9636;
wire n_9637, n_9638, n_9639, n_9640, n_9641, n_9644, n_9645, n_9646;
wire n_9647, n_9648, n_9649, n_9650, n_9651, n_9654, n_9656, n_9660;
wire n_9661, n_9665, n_9668, n_9669, n_9672, n_9673, n_9674, n_9675;
wire n_9676, n_9681, n_9682, n_9683, n_9685, n_9686, n_9688, n_9690;
wire n_9691, n_9692, n_9693, n_9694, n_9695, n_9696, n_9697, n_9698;
wire n_9699, n_9700, n_9701, n_9702, n_9703, n_9704, n_9705, n_9706;
wire n_9707, n_9708, n_9709, n_9710, n_9711, n_9712, n_9713, n_9714;
wire n_9715, n_9716, n_9717, n_9718, n_9719, n_9720, n_9721, n_9722;
wire n_9726, n_9727, n_9729, n_9730, n_9732, n_9734, n_9735, n_9736;
wire n_9737, n_9738, n_9739, n_9742, n_9743, n_9745, n_9746, n_9748;
wire n_9750, n_9753, n_9754, n_9755, n_9756, n_9759, n_9762, n_9763;
wire n_9764, n_9765, n_9767, n_9769, n_9772, n_9773, n_9774, n_9775;
wire n_9779, n_9781, n_9782, n_9783, n_9784, n_9785, n_9786, n_9787;
wire n_9789, n_9790, n_9791, n_9792, n_9793, n_9794, n_9795, n_9796;
wire n_9797, n_9798, n_9799, n_9800, n_9801, n_9802, n_9803, n_9804;
wire n_9805, n_9807, n_9808, n_9809, n_9810, n_9811, n_9814, n_9815;
wire n_9817, n_9818, n_9819, n_9820, n_9821, n_9823, n_9825, n_9827;
wire n_9828, n_9829, n_9830, n_9831, n_9832, n_9834, n_9835, n_9837;
wire n_9838, n_9841, n_9842, n_9843, n_9844, n_9845, n_9846, n_9847;
wire n_9848, n_9849, n_9850, n_9852, n_9856, n_9858, n_9860, n_9863;
wire n_9864, n_9866, n_9868, n_9869, n_9870, n_9871, n_9872, n_9873;
wire n_9874, n_9875, n_9876, n_9878, n_9879, n_9882, n_9883, n_9884;
wire n_9885, n_9889, n_9891, n_9892, n_9893, n_9894, n_9896, n_9897;
wire n_9899, n_9900, n_9901, n_9903, n_9904, n_9905, n_9906, n_9907;
wire n_9908, n_9909, n_9910, n_9911, n_9912, n_9913, n_9914, n_9915;
wire n_9916, n_9917, n_9918, n_9920, n_9921, n_9922, n_9923, n_9924;
wire n_9927, n_9928, n_9929, n_9930, n_9931, n_9933, n_9935, n_9936;
wire n_9937, n_9938, n_9939, n_9940, n_9942, n_9943, n_9944, n_9946;
wire n_9947, n_9948, n_9949, n_9950, n_9951, n_9952, n_9953, n_9955;
wire n_9956, n_9957, n_9958, n_9959, n_9960, n_9961, n_9962, n_9963;
wire n_9965, n_9966, n_9968, n_9970, n_9976, n_9977, n_9978, n_9979;
wire n_9980, n_9981, n_9982, n_9987, n_9988, n_9990, n_9991, n_9992;
wire n_9993, n_9995, n_9996, n_9997, n_9999, n_10000, n_10003,n_10005;
wire n_10008, n_10012, n_10014, n_10017, n_10018, n_10020, n_10023,n_10025;
wire n_10026, n_10027, n_10028, n_10029, n_10030, n_10031, n_10034,n_10035;
wire n_10036, n_10037, n_10038, n_10041, n_10043, n_10044, n_10046,n_10048;
wire n_10049, n_10050, n_10051, n_10052, n_10053, n_10057, n_10058,n_10060;
wire n_10061, n_10062, n_10063, n_10065, n_10069, n_10071, n_10072,n_10074;
wire n_10077, n_10078, n_10079, n_10081, n_10082, n_10083, n_10084,n_10085;
wire n_10087, n_10088, n_10089, n_10090, n_10091, n_10093, n_10094,n_10095;
wire n_10096, n_10098, n_10099, n_10100, n_10101, n_10102, n_10104,n_10105;
wire n_10108, n_10109, n_10110, n_10112, n_10115, n_10119, n_10121,n_10122;
wire n_10124, n_10125, n_10126, n_10127, n_10129, n_10130, n_10131,n_10133;
wire n_10134, n_10135, n_10136, n_10137, n_10138, n_10139, n_10140,n_10141;
wire n_10142, n_10144, n_10146, n_10147, n_10149, n_10150, n_10152,n_10154;
wire n_10156, n_10157, n_10158, n_10160, n_10162, n_10163, n_10164,n_10165;
wire n_10166, n_10170, n_10171, n_10172, n_10174, n_10175, n_10177,n_10179;
wire n_10180, n_10181, n_10182, n_10183, n_10185, n_10188, n_10191,n_10192;
wire n_10193, n_10194, n_10195, n_10197, n_10198, n_10199, n_10201,n_10202;
wire n_10203, n_10204, n_10206, n_10207, n_10208, n_10209, n_10212,n_10213;
wire n_10215, n_10216, n_10217, n_10218, n_10220, n_10221, n_10222,n_10223;
wire n_10226, n_10227, n_10229, n_10231, n_10232, n_10235, n_10237,n_10238;
wire n_10239, n_10241, n_10242, n_10243, n_10245, n_10248, n_10249,n_10250;
wire n_10251, n_10252, n_10253, n_10254, n_10255, n_10258, n_10260,n_10263;
wire n_10264, n_10265, n_10266, n_10267, n_10268, n_10269, n_10272,n_10273;
wire n_10277, n_10278, n_10279, n_10283, n_10284, n_10285, n_10286,n_10287;
wire n_10288, n_10289, n_10290, n_10292, n_10294, n_10295, n_10296,n_10297;
wire n_10299, n_10302, n_10304, n_10305, n_10306, n_10307, n_10309,n_10311;
wire n_10312, n_10313, n_10314, n_10315, n_10316, n_10317, n_10318,n_10319;
wire n_10320, n_10321, n_10322, n_10323, n_10324, n_10326, n_10327,n_10328;
wire n_10329, n_10331, n_10332, n_10333, n_10334, n_10336, n_10337,n_10338;
wire n_10339, n_10341, n_10342, n_10344, n_10345, n_10346, n_10347,n_10348;
wire n_10350, n_10351, n_10353, n_10354, n_10355, n_10356, n_10357,n_10358;
wire n_10359, n_10361, n_10362, n_10366, n_10367, n_10369, n_10370,n_10372;
wire n_10373, n_10374, n_10376, n_10377, n_10380, n_10381, n_10382,n_10383;
wire n_10384, n_10385, n_10387, n_10389, n_10390, n_10391, n_10392,n_10393;
wire n_10395, n_10396, n_10397, n_10398, n_10400, n_10401, n_10402,n_10405;
wire n_10407, n_10408, n_10410, n_10411, n_10413, n_10414, n_10415,n_10417;
wire n_10418, n_10421, n_10424, n_10425, n_10429, n_10431, n_10432,n_10434;
wire n_10436, n_10437, n_10438, n_10440, n_10441, n_10443, n_10444,n_10445;
wire n_10447, n_10448, n_10449, n_10451, n_10452, n_10453, n_10454,n_10455;
wire n_10456, n_10457, n_10460, n_10462, n_10463, n_10465, n_10466,n_10467;
wire n_10469, n_10471, n_10472, n_10474, n_10475, n_10476, n_10478,n_10480;
wire n_10481, n_10483, n_10484, n_10485, n_10486, n_10488, n_10489,n_10492;
wire n_10493, n_10495, n_10496, n_10498, n_10501, n_10502, n_10506,n_10507;
wire n_10508, n_10509, n_10510, n_10512, n_10513, n_10514, n_10515,n_10516;
wire n_10518, n_10519, n_10520, n_10521, n_10522, n_10523, n_10524,n_10531;
wire n_10535, n_10537, n_10539, n_10542, n_10543, n_10546, n_10547,n_10548;
wire n_10549, n_10550, n_10551, n_10552, n_10556, n_10561, n_10562,n_10565;
wire n_10566, n_10569, n_10573, n_10574, n_10575, n_10580, n_10581,n_10585;
wire n_10586, n_10589, n_10590, n_10595, n_10598, n_10599, n_10600,n_10603;
wire n_10604, n_10605, n_10607, n_10608, n_10609, n_10610, n_10613,n_10616;
wire n_10618, n_10619, n_10621, n_10622, n_10629, n_10630, n_10631,n_10632;
wire n_10633, n_10634, n_10635, n_10637, n_10638, n_10640, n_10644,n_10645;
wire n_10646, n_10653, n_10654, n_10655, n_10656, n_10657, n_10658,n_10659;
wire n_10660, n_10661, n_10662, n_10663, n_10664, n_10665, n_10667,n_10668;
wire n_10669, n_10670, n_10671, n_10672, n_10673, n_10674, n_10675,n_10676;
wire n_10677, n_10678, n_10679, n_10680, n_10681, n_10682, n_10683,n_10685;
wire n_10686, n_10687, n_10688, n_10690, n_10691, n_10692, n_10693,n_10694;
wire n_10696, n_10697, n_10698, n_10699, n_10700, n_10701, n_10702,n_10703;
wire n_10704, n_10705, n_10706, n_10707, n_10708, n_10710, n_10711,n_10712;
wire n_10713, n_10714, n_10716, n_10717, n_10718, n_10719, n_10720,n_10721;
wire n_10723, n_10724, n_10725, n_10726, n_10727, n_10728, n_10729,n_10730;
wire n_10731, n_10732, n_10733, n_10734, n_10735, n_10737, n_10738,n_10740;
wire n_10741, n_10742, n_10743, n_10744, n_10745, n_10746, n_10747,n_10748;
wire n_10749, n_10750, n_10751, n_10752, n_10754, n_10756, n_10757,n_10758;
wire n_10759, n_10760, n_10761, n_10763, n_10765, n_10767, n_10768,n_10769;
wire n_10770, n_10771, n_10774, n_10775, n_10776, n_10777, n_10778,n_10779;
wire n_10780, n_10781, n_10782, n_10783, n_10784, n_10785, n_10786,n_10788;
wire n_10789, n_10790, n_10791, n_10792, n_10794, n_10795, n_10796,n_10797;
wire n_10798, n_10799, n_10801, n_10802, n_10804, n_10805, n_10806,n_10807;
wire n_10809, n_10810, n_10812, n_10815, n_10816, n_10817, n_10818,n_10819;
wire n_10820, n_10821, n_10822, n_10823, n_10824, n_10825, n_10826,n_10827;
wire n_10828, n_10829, n_10830, n_10831, n_10832, n_10833, n_10834,n_10835;
wire n_10836, n_10837, n_10838, n_10839, n_10840, n_10841, n_10842,n_10843;
wire n_10844, n_10845, n_10846, n_10847, n_10849, n_10850, n_10851,n_10853;
wire n_10854, n_10855, n_10856, n_10857, n_10858, n_10859, n_10860,n_10861;
wire n_10862, n_10863, n_10864, n_10865, n_10866, n_10867, n_10868,n_10869;
wire n_10870, n_10871, n_10873, n_10874, n_10876, n_10878, n_10879,n_10880;
wire n_10881, n_10882, n_10883, n_10885, n_10887, n_10888, n_10889,n_10890;
wire n_10891, n_10892, n_10893, n_10894, n_10896, n_10897, n_10900,n_10901;
wire n_10902, n_10903, n_10904, n_10905, n_10906, n_10907, n_10909,n_10910;
wire n_10911, n_10912, n_10913, n_10914, n_10915, n_10916, n_10917,n_10918;
wire n_10919, n_10920, n_10921, n_10922, n_10923, n_10924, n_10926,n_10927;
wire n_10928, n_10930, n_10931, n_10932, n_10933, n_10934, n_10935,n_10936;
wire n_10937, n_10938, n_10939, n_10940, n_10941, n_10943, n_10945,n_10947;
wire n_10948, n_10949, n_10950, n_10952, n_10954, n_10955, n_10956,n_10957;
wire n_10959, n_10960, n_10961, n_10962, n_10964, n_10967, n_10968,n_10969;
wire n_10971, n_10972, n_10974, n_10975, n_10976, n_10977, n_10978,n_10979;
wire n_10980, n_10982, n_10983, n_10984, n_10985, n_10986, n_10987,n_10988;
wire n_10991, n_10992, n_10993, n_10994, n_10995, n_10996, n_10997,n_10998;
wire n_10999, n_11000, n_11001, n_11002, n_11003, n_11004, n_11005,n_11006;
wire n_11007, n_11008, n_11010, n_11011, n_11012, n_11013, n_11014,n_11015;
wire n_11017, n_11019, n_11020, n_11021, n_11022, n_11023, n_11024,n_11025;
wire n_11027, n_11028, n_11029, n_11030, n_11031, n_11032, n_11033,n_11034;
wire n_11035, n_11036, n_11039, n_11040, n_11041, n_11042, n_11043,n_11045;
wire n_11046, n_11047, n_11049, n_11050, n_11051, n_11052, n_11053,n_11056;
wire n_11057, n_11059, n_11060, n_11061, n_11062, n_11063, n_11064,n_11065;
wire n_11066, n_11067, n_11068, n_11071, n_11072, n_11073, n_11074,n_11075;
wire n_11076, n_11077, n_11078, n_11079, n_11080, n_11081, n_11083,n_11084;
wire n_11085, n_11086, n_11087, n_11088, n_11089, n_11091, n_11092,n_11094;
wire n_11095, n_11096, n_11097, n_11098, n_11099, n_11100, n_11102,n_11103;
wire n_11104, n_11105, n_11106, n_11107, n_11108, n_11109, n_11110,n_11111;
wire n_11112, n_11113, n_11114, n_11115, n_11116, n_11117, n_11118,n_11119;
wire n_11120, n_11122, n_11123, n_11124, n_11125, n_11126, n_11127,n_11131;
wire n_11132, n_11133, n_11134, n_11135, n_11137, n_11138, n_11139,n_11141;
wire n_11142, n_11143, n_11144, n_11145, n_11146, n_11150, n_11151,n_11152;
wire n_11154, n_11155, n_11156, n_11157, n_11158, n_11159, n_11161,n_11162;
wire n_11163, n_11165, n_11167, n_11168, n_11171, n_11172, n_11173,n_11175;
wire n_11177, n_11178, n_11179, n_11181, n_11182, n_11183, n_11184,n_11185;
wire n_11186, n_11188, n_11189, n_11190, n_11191, n_11192, n_11193,n_11194;
wire n_11195, n_11196, n_11197, n_11198, n_11199, n_11200, n_11203,n_11204;
wire n_11206, n_11207, n_11208, n_11209, n_11211, n_11213, n_11214,n_11215;
wire n_11217, n_11219, n_11220, n_11221, n_11222, n_11223, n_11224,n_11227;
wire n_11228, n_11230, n_11231, n_11233, n_11234, n_11235, n_11237,n_11238;
wire n_11240, n_11241, n_11242, n_11244, n_11246, n_11247, n_11249,n_11250;
wire n_11251, n_11253, n_11254, n_11255, n_11256, n_11257, n_11258,n_11259;
wire n_11260, n_11261, n_11262, n_11263, n_11264, n_11266, n_11267,n_11271;
wire n_11272, n_11273, n_11275, n_11276, n_11277, n_11278, n_11279,n_11280;
wire n_11281, n_11282, n_11284, n_11285, n_11286, n_11287, n_11288,n_11290;
wire n_11291, n_11292, n_11295, n_11296, n_11298, n_11299, n_11300,n_11302;
wire n_11303, n_11304, n_11305, n_11307, n_11309, n_11311, n_11312,n_11313;
wire n_11315, n_11316, n_11317, n_11318, n_11319, n_11321, n_11322,n_11323;
wire n_11324, n_11325, n_11326, n_11327, n_11328, n_11329, n_11330,n_11331;
wire n_11332, n_11333, n_11334, n_11336, n_11337, n_11338, n_11339,n_11340;
wire n_11342, n_11345, n_11346, n_11348, n_11349, n_11350, n_11351,n_11353;
wire n_11354, n_11356, n_11358, n_11359, n_11361, n_11362, n_11363,n_11365;
wire n_11366, n_11367, n_11368, n_11369, n_11371, n_11373, n_11374,n_11375;
wire n_11377, n_11378, n_11379, n_11380, n_11381, n_11383, n_11384,n_11385;
wire n_11386, n_11387, n_11388, n_11389, n_11390, n_11391, n_11393,n_11394;
wire n_11395, n_11397, n_11400, n_11401, n_11404, n_11406, n_11407,n_11409;
wire n_11411, n_11412, n_11413, n_11414, n_11416, n_11417, n_11418,n_11419;
wire n_11420, n_11421, n_11422, n_11423, n_11424, n_11425, n_11426,n_11428;
wire n_11431, n_11432, n_11433, n_11434, n_11435, n_11436, n_11437,n_11438;
wire n_11439, n_11440, n_11445, n_11447, n_11448, n_11449, n_11450,n_11451;
wire n_11452, n_11453, n_11454, n_11456, n_11457, n_11460, n_11461,n_11462;
wire n_11463, n_11464, n_11465, n_11466, n_11468, n_11469, n_11470,n_11471;
wire n_11473, n_11474, n_11476, n_11478, n_11480, n_11483, n_11484,n_11485;
wire n_11486, n_11487, n_11488, n_11489, n_11490, n_11491, n_11492,n_11493;
wire n_11494, n_11495, n_11496, n_11498, n_11499, n_11500, n_11501,n_11502;
wire n_11503, n_11504, n_11505, n_11506, n_11507, n_11508, n_11509,n_11510;
wire n_11511, n_11512, n_11513, n_11514, n_11515, n_11516, n_11517,n_11518;
wire n_11519, n_11520, n_11521, n_11522, n_11523, n_11524, n_11525,n_11527;
wire n_11528, n_11529, n_11530, n_11531, n_11532, n_11533, n_11534,n_11535;
wire n_11538, n_11539, n_11540, n_11542, n_11543, n_11544, n_11545,n_11546;
wire n_11547, n_11549, n_11550, n_11551, n_11553, n_11554, n_11555,n_11556;
wire n_11557, n_11558, n_11559, n_11560, n_11561, n_11562, n_11563,n_11564;
wire n_11565, n_11566, n_11567, n_11568, n_11569, n_11570, n_11572,n_11573;
wire n_11574, n_11575, n_11576, n_11577, n_11578, n_11579, n_11580,n_11581;
wire n_11582, n_11583, n_11584, n_11585, n_11586, n_11587, n_11589,n_11590;
wire n_11592, n_11593, n_11594, n_11596, n_11597, n_11598, n_11599,n_11600;
wire n_11601, n_11602, n_11603, n_11604, n_11606, n_11608, n_11609,n_11611;
wire n_11612, n_11613, n_11614, n_11615, n_11616, n_11617, n_11618,n_11620;
wire n_11621, n_11623, n_11624, n_11625, n_11626, n_11627, n_11628,n_11632;
wire n_11636, n_11641, n_11642, n_11643, n_11647, n_11648, n_11649,n_11650;
wire n_11655, n_11656, n_11658, n_11660, n_11661, n_11662, n_11663,n_11664;
wire n_11666, n_11667, n_11668, n_11669, n_11670, n_11671, n_11672,n_11674;
wire n_11676, n_11677, n_11678, n_11681, n_11682, n_11683, n_11685,n_11686;
wire n_11687, n_11689, n_11690, n_11694, n_11696, n_11698, n_11699,n_11700;
wire n_11701, n_11705, n_11707, n_11709, n_11710, n_11712, n_11713,n_11714;
wire n_11715, n_11716, n_11718, n_11725, n_11727, n_11728, n_11729,n_11730;
wire n_11731, n_11732, n_11733, n_11734, n_11735, n_11738, n_11739,n_11740;
wire n_11741, n_11742, n_11743, n_11744, n_11745, n_11746, n_11749,n_11750;
wire n_11752, n_11753, n_11756, n_11758, n_11760, n_11762, n_11764,n_11768;
wire n_11772, n_11773, n_11774, n_11776, n_11777, n_11778, n_11782,n_11784;
wire n_11787, n_11791, n_11792, n_11795, n_11798, n_11799, n_11800,n_11801;
wire n_11802, n_11805, n_11808, n_11810, n_11811, n_11812, n_11815,n_11816;
wire n_11817, n_11818, n_11819, n_11820, n_11821, n_11823, n_11827,n_11831;
wire n_11833, n_11834, n_11835, n_11836, n_11837, n_11839, n_11842,n_11843;
wire n_11845, n_11848, n_11849, n_11850, n_11851, n_11853, n_11854,n_11856;
wire n_11857, n_11858, n_11860, n_11861, n_11862, n_11864, n_11865,n_11871;
wire n_11875, n_11876, n_11877, n_11878, n_11880, n_11882, n_11883,n_11884;
wire n_11885, n_11886, n_11887, n_11888, n_11889, n_11893, n_11895,n_11897;
wire n_11898, n_11900, n_11901, n_11902, n_11909, n_11914, n_11916,n_11917;
wire n_11918, n_11920, n_11921, n_11923, n_11924, n_11925, n_11927,n_11929;
wire n_11931, n_11932, n_11934, n_11936, n_11940, n_11945, n_11946,n_11948;
wire n_11949, n_11951, n_11953, n_11956, n_11957, n_11958, n_11963,n_11965;
wire n_11967, n_11972, n_11975, n_11976, n_11977, n_11978, n_11980,n_11981;
wire n_11984, n_11985, n_11988, n_11989, n_11990, n_11993, n_11994,n_11996;
wire n_11998, n_11999, n_12001, n_12006, n_12009, n_12012, n_12013,n_12014;
wire n_12015, n_12019, n_12020, n_12021, n_12023, n_12024, n_12025,n_12026;
wire n_12027, n_12028, n_12029, n_12032, n_12036, n_12042, n_12043,n_12049;
wire n_12052, n_12054, n_12055, n_12056, n_12057, n_12058, n_12059,n_12060;
wire n_12061, n_12063, n_12067, n_12068, n_12070, n_12071, n_12072,n_12073;
wire n_12075, n_12077, n_12078, n_12079, n_12081, n_12082, n_12085,n_12091;
wire n_12093, n_12095, n_12096, n_12098, n_12099, n_12100, n_12102,n_12105;
wire n_12106, n_12108, n_12112, n_12113, n_12114, n_12115, n_12116,n_12117;
wire n_12118, n_12119, n_12120, n_12121, n_12122, n_12123, n_12124,n_12125;
wire n_12126, n_12127, n_12128, n_12129, n_12130, n_12132, n_12133,n_12134;
wire n_12135, n_12136, n_12137, n_12138, n_12139, n_12140, n_12141,n_12143;
wire n_12144, n_12145, n_12146, n_12148, n_12149, n_12150, n_12152,n_12153;
wire n_12154, n_12155, n_12156, n_12158, n_12159, n_12160, n_12161,n_12162;
wire n_12163, n_12165, n_12166, n_12167, n_12168, n_12169, n_12170,n_12172;
wire n_12173, n_12174, n_12175, n_12176, n_12177, n_12178, n_12180,n_12181;
wire n_12182, n_12183, n_12185, n_12186, n_12187, n_12188, n_12189,n_12190;
wire n_12191, n_12192, n_12193, n_12194, n_12195, n_12197, n_12198,n_12199;
wire n_12200, n_12202, n_12203, n_12204, n_12205, n_12206, n_12207,n_12208;
wire n_12209, n_12210, n_12211, n_12212, n_12213, n_12214, n_12215,n_12216;
wire n_12217, n_12219, n_12220, n_12221, n_12222, n_12223, n_12224,n_12225;
wire n_12226, n_12227, n_12228, n_12230, n_12231, n_12233, n_12234,n_12235;
wire n_12237, n_12238, n_12239, n_12242, n_12243, n_12244, n_12245,n_12246;
wire n_12247, n_12248, n_12249, n_12250, n_12251, n_12252, n_12253,n_12254;
wire n_12255, n_12256, n_12257, n_12258, n_12260, n_12261, n_12263,n_12264;
wire n_12265, n_12266, n_12267, n_12268, n_12270, n_12271, n_12272,n_12274;
wire n_12275, n_12276, n_12277, n_12278, n_12279, n_12280, n_12281,n_12282;
wire n_12285, n_12286, n_12288, n_12289, n_12290, n_12291, n_12292,n_12293;
wire n_12294, n_12296, n_12298, n_12299, n_12300, n_12301, n_12302,n_12303;
wire n_12305, n_12306, n_12307, n_12308, n_12309, n_12310, n_12312,n_12313;
wire n_12314, n_12315, n_12316, n_12317, n_12319, n_12320, n_12321,n_12322;
wire n_12323, n_12324, n_12325, n_12326, n_12327, n_12328, n_12329,n_12330;
wire n_12331, n_12333, n_12334, n_12335, n_12336, n_12337, n_12338,n_12339;
wire n_12340, n_12341, n_12342, n_12344, n_12345, n_12346, n_12347,n_12348;
wire n_12349, n_12350, n_12351, n_12352, n_12353, n_12354, n_12355,n_12356;
wire n_12358, n_12359, n_12360, n_12361, n_12362, n_12363, n_12364,n_12365;
wire n_12366, n_12368, n_12369, n_12370, n_12371, n_12372, n_12373,n_12374;
wire n_12375, n_12376, n_12377, n_12378, n_12379, n_12380, n_12381,n_12382;
wire n_12383, n_12384, n_12385, n_12386, n_12387, n_12389, n_12390,n_12392;
wire n_12393, n_12395, n_12396, n_12397, n_12399, n_12400, n_12402,n_12403;
wire n_12404, n_12405, n_12406, n_12408, n_12409, n_12410, n_12411,n_12412;
wire n_12413, n_12414, n_12416, n_12417, n_12418, n_12420, n_12421,n_12422;
wire n_12423, n_12424, n_12425, n_12426, n_12427, n_12428, n_12429,n_12430;
wire n_12432, n_12433, n_12435, n_12436, n_12437, n_12438, n_12439,n_12440;
wire n_12441, n_12443, n_12444, n_12445, n_12446, n_12447, n_12448,n_12449;
wire n_12450, n_12451, n_12452, n_12457, n_12459, n_12460, n_12461,n_12462;
wire n_12463, n_12465, n_12466, n_12467, n_12468, n_12469, n_12470,n_12471;
wire n_12472, n_12473, n_12474, n_12475, n_12476, n_12477, n_12478,n_12479;
wire n_12480, n_12481, n_12483, n_12484, n_12485, n_12486, n_12487,n_12488;
wire n_12493, n_12494, n_12495, n_12496, n_12497, n_12498, n_12499,n_12500;
wire n_12501, n_12502, n_12503, n_12504, n_12505, n_12506, n_12507,n_12508;
wire n_12509, n_12510, n_12512, n_12513, n_12514, n_12515, n_12516,n_12517;
wire n_12518, n_12520, n_12521, n_12524, n_12526, n_12527, n_12528,n_12529;
wire n_12530, n_12531, n_12532, n_12533, n_12534, n_12535, n_12536,n_12538;
wire n_12541, n_12542, n_12544, n_12545, n_12546, n_12548, n_12549,n_12550;
wire n_12553, n_12555, n_12556, n_12558, n_12559, n_12560, n_12561,n_12562;
wire n_12563, n_12564, n_12565, n_12566, n_12567, n_12568, n_12569,n_12570;
wire n_12571, n_12572, n_12573, n_12576, n_12578, n_12580, n_12581,n_12582;
wire n_12584, n_12586, n_12587, n_12588, n_12589, n_12591, n_12592,n_12593;
wire n_12594, n_12596, n_12597, n_12598, n_12599, n_12601, n_12603,n_12604;
wire n_12605, n_12607, n_12609, n_12610, n_12612, n_12613, n_12614,n_12617;
wire n_12620, n_12624, n_12625, n_12626, n_12627, n_12628, n_12629,n_12630;
wire n_12631, n_12632, n_12633, n_12634, n_12635, n_12636, n_12637,n_12638;
wire n_12639, n_12640, n_12641, n_12642, n_12643, n_12644, n_12645,n_12646;
wire n_12647, n_12648, n_12649, n_12650, n_12652, n_12653, n_12654,n_12655;
wire n_12656, n_12657, n_12658, n_12660, n_12661, n_12662, n_12663,n_12664;
wire n_12665, n_12666, n_12667, n_12668, n_12669, n_12670, n_12671,n_12672;
wire n_12673, n_12674, n_12675, n_12676, n_12677, n_12678, n_12680,n_12681;
wire n_12682, n_12686, n_12688, n_12691, n_12692, n_12694, n_12695,n_12696;
wire n_12697, n_12698, n_12699, n_12701, n_12702, n_12703, n_12705,n_12706;
wire n_12707, n_12708, n_12709, n_12710, n_12712, n_12713, n_12714,n_12715;
wire n_12716, n_12717, n_12718, n_12719, n_12720, n_12721, n_12722,n_12723;
wire n_12724, n_12725, n_12727, n_12728, n_12730, n_12731, n_12732,n_12733;
wire n_12734, n_12735, n_12736, n_12737, n_12738, n_12739, n_12740,n_12741;
wire n_12742, n_12745, n_12746, n_12747, n_12748, n_12749, n_12750,n_12751;
wire n_12752, n_12753, n_12754, n_12755, n_12756, n_12759, n_12760,n_12761;
wire n_12762, n_12763, n_12765, n_12767, n_12768, n_12769, n_12771,n_12772;
wire n_12773, n_12774, n_12775, n_12776, n_12777, n_12778, n_12779,n_12780;
wire n_12781, n_12782, n_12783, n_12784, n_12785, n_12786, n_12787,n_12788;
wire n_12789, n_12792, n_12794, n_12795, n_12796, n_12797, n_12798,n_12800;
wire n_12801, n_12802, n_12803, n_12804, n_12805, n_12806, n_12807,n_12810;
wire n_12811, n_12813, n_12814, n_12815, n_12816, n_12817, n_12818,n_12819;
wire n_12822, n_12823, n_12824, n_12825, n_12827, n_12828, n_12829,n_12830;
wire n_12831, n_12833, n_12834, n_12835, n_12836, n_12838, n_12840,n_12843;
wire n_12844, n_12845, n_12846, n_12847, n_12848, n_12849, n_12850,n_12851;
wire n_12852, n_12853, n_12854, n_12855, n_12856, n_12857, n_12858,n_12859;
wire n_12860, n_12861, n_12862, n_12864, n_12865, n_12868, n_12869,n_12870;
wire n_12871, n_12872, n_12873, n_12875, n_12877, n_12879, n_12880,n_12881;
wire n_12882, n_12883, n_12884, n_12885, n_12886, n_12887, n_12890,n_12892;
wire n_12893, n_12894, n_12895, n_12896, n_12898, n_12900, n_12902,n_12903;
wire n_12906, n_12907, n_12909, n_12910, n_12911, n_12912, n_12914,n_12916;
wire n_12917, n_12918, n_12919, n_12920, n_12922, n_12923, n_12924,n_12925;
wire n_12926, n_12928, n_12929, n_12930, n_12931, n_12932, n_12934,n_12935;
wire n_12937, n_12938, n_12939, n_12941, n_12943, n_12944, n_12945,n_12946;
wire n_12950, n_12952, n_12953, n_12955, n_12957, n_12958, n_12959,n_12960;
wire n_12963, n_12964, n_12965, n_12966, n_12968, n_12969, n_12970,n_12971;
wire n_12972, n_12973, n_12974, n_12977, n_12979, n_12980, n_12981,n_12983;
wire n_12984, n_12985, n_12986, n_12987, n_12988, n_12989, n_12990,n_12991;
wire n_12993, n_12994, n_12995, n_12996, n_12997, n_12998, n_13000,n_13002;
wire n_13003, n_13004, n_13005, n_13006, n_13008, n_13010, n_13011,n_13012;
wire n_13013, n_13015, n_13016, n_13018, n_13019, n_13020, n_13022,n_13023;
wire n_13025, n_13026, n_13027, n_13028, n_13030, n_13031, n_13032,n_13033;
wire n_13034, n_13035, n_13036, n_13037, n_13039, n_13040, n_13042,n_13043;
wire n_13044, n_13046, n_13047, n_13050, n_13051, n_13052, n_13053,n_13054;
wire n_13055, n_13056, n_13058, n_13060, n_13062, n_13063, n_13064,n_13065;
wire n_13066, n_13067, n_13068, n_13069, n_13071, n_13072, n_13073,n_13074;
wire n_13076, n_13077, n_13079, n_13080, n_13081, n_13082, n_13083,n_13084;
wire n_13087, n_13090, n_13092, n_13093, n_13094, n_13095, n_13097,n_13098;
wire n_13101, n_13102, n_13104, n_13105, n_13107, n_13108, n_13109,n_13110;
wire n_13113, n_13114, n_13115, n_13116, n_13117, n_13118, n_13119,n_13120;
wire n_13121, n_13122, n_13123, n_13124, n_13125, n_13126, n_13127,n_13128;
wire n_13129, n_13130, n_13132, n_13133, n_13134, n_13135, n_13136,n_13137;
wire n_13138, n_13139, n_13140, n_13141, n_13142, n_13143, n_13144,n_13145;
wire n_13146, n_13147, n_13148, n_13149, n_13151, n_13152, n_13153,n_13154;
wire n_13156, n_13157, n_13158, n_13159, n_13160, n_13162, n_13163,n_13164;
wire n_13165, n_13166, n_13167, n_13168, n_13169, n_13170, n_13171,n_13172;
wire n_13173, n_13174, n_13175, n_13176, n_13177, n_13178, n_13179,n_13180;
wire n_13181, n_13182, n_13183, n_13184, n_13185, n_13186, n_13187,n_13188;
wire n_13189, n_13190, n_13191, n_13192, n_13193, n_13194, n_13195,n_13196;
wire n_13197, n_13198, n_13199, n_13200, n_13201, n_13202, n_13203,n_13204;
wire n_13205, n_13206, n_13207, n_13208, n_13209, n_13210, n_13211,n_13212;
wire n_13213, n_13214, n_13216, n_13217, n_13218, n_13219, n_13220,n_13221;
wire n_13222, n_13223, n_13225, n_13226, n_13227, n_13229, n_13230,n_13231;
wire n_13232, n_13233, n_13234, n_13235, n_13236, n_13237, n_13239,n_13240;
wire n_13241, n_13242, n_13243, n_13244, n_13246, n_13247, n_13248,n_13249;
wire n_13250, n_13252, n_13253, n_13254, n_13255, n_13256, n_13257,n_13258;
wire n_13259, n_13260, n_13261, n_13262, n_13263, n_13265, n_13267,n_13268;
wire n_13269, n_13270, n_13271, n_13272, n_13274, n_13275, n_13276,n_13277;
wire n_13278, n_13279, n_13280, n_13281, n_13282, n_13283, n_13285,n_13288;
wire n_13290, n_13291, n_13293, n_13294, n_13295, n_13296, n_13298,n_13299;
wire n_13300, n_13301, n_13302, n_13303, n_13305, n_13306, n_13307,n_13308;
wire n_13309, n_13310, n_13311, n_13312, n_13313, n_13314, n_13315,n_13316;
wire n_13317, n_13318, n_13319, n_13320, n_13321, n_13322, n_13323,n_13324;
wire n_13325, n_13326, n_13327, n_13328, n_13329, n_13330, n_13331,n_13332;
wire n_13333, n_13334, n_13335, n_13336, n_13337, n_13340, n_13341,n_13342;
wire n_13344, n_13345, n_13346, n_13347, n_13348, n_13349, n_13350,n_13351;
wire n_13352, n_13355, n_13356, n_13357, n_13358, n_13359, n_13360,n_13361;
wire n_13362, n_13363, n_13364, n_13365, n_13366, n_13367, n_13368,n_13369;
wire n_13370, n_13371, n_13372, n_13373, n_13374, n_13375, n_13376,n_13378;
wire n_13379, n_13380, n_13381, n_13382, n_13383, n_13384, n_13385,n_13387;
wire n_13388, n_13389, n_13390, n_13393, n_13395, n_13396, n_13397,n_13398;
wire n_13399, n_13402, n_13403, n_13404, n_13405, n_13407, n_13408,n_13410;
wire n_13411, n_13412, n_13414, n_13415, n_13416, n_13417, n_13418,n_13419;
wire n_13420, n_13421, n_13422, n_13423, n_13424, n_13425, n_13426,n_13427;
wire n_13428, n_13429, n_13430, n_13431, n_13432, n_13433, n_13434,n_13435;
wire n_13436, n_13437, n_13438, n_13440, n_13441, n_13442, n_13443,n_13444;
wire n_13445, n_13446, n_13447, n_13448, n_13449, n_13450, n_13451,n_13452;
wire n_13454, n_13455, n_13457, n_13458, n_13460, n_13461, n_13462,n_13463;
wire n_13465, n_13466, n_13467, n_13468, n_13469, n_13470, n_13471,n_13472;
wire n_13473, n_13474, n_13475, n_13476, n_13477, n_13479, n_13481,n_13482;
wire n_13483, n_13484, n_13485, n_13487, n_13488, n_13489, n_13490,n_13491;
wire n_13492, n_13493, n_13495, n_13496, n_13497, n_13498, n_13499,n_13502;
wire n_13503, n_13504, n_13505, n_13506, n_13507, n_13508, n_13510,n_13511;
wire n_13512, n_13513, n_13514, n_13515, n_13516, n_13517, n_13518,n_13519;
wire n_13520, n_13521, n_13522, n_13524, n_13525, n_13526, n_13527,n_13528;
wire n_13530, n_13531, n_13532, n_13534, n_13535, n_13536, n_13537,n_13538;
wire n_13539, n_13542, n_13543, n_13544, n_13546, n_13547, n_13548,n_13549;
wire n_13550, n_13551, n_13552, n_13553, n_13554, n_13555, n_13556,n_13557;
wire n_13559, n_13560, n_13561, n_13562, n_13563, n_13564, n_13565,n_13566;
wire n_13567, n_13568, n_13569, n_13570, n_13571, n_13572, n_13573,n_13574;
wire n_13575, n_13576, n_13578, n_13579, n_13581, n_13582, n_13584,n_13585;
wire n_13587, n_13588, n_13589, n_13590, n_13592, n_13593, n_13594,n_13595;
wire n_13596, n_13598, n_13602, n_13603, n_13604, n_13605, n_13606,n_13607;
wire n_13608, n_13609, n_13610, n_13611, n_13612, n_13613, n_13614,n_13616;
wire n_13617, n_13618, n_13619, n_13621, n_13622, n_13623, n_13624,n_13625;
wire n_13626, n_13628, n_13630, n_13632, n_13633, n_13635, n_13636,n_13637;
wire n_13638, n_13640, n_13642, n_13644, n_13645, n_13646, n_13647,n_13649;
wire n_13651, n_13652, n_13654, n_13655, n_13656, n_13657, n_13659,n_13660;
wire n_13661, n_13663, n_13664, n_13665, n_13666, n_13667, n_13668,n_13670;
wire n_13671, n_13672, n_13674, n_13675, n_13676, n_13677, n_13678,n_13679;
wire n_13680, n_13681, n_13682, n_13684, n_13685, n_13686, n_13688,n_13690;
wire n_13694, n_13695, n_13696, n_13697, n_13698, n_13699, n_13700,n_13701;
wire n_13702, n_13703, n_13704, n_13705, n_13706, n_13708, n_13709,n_13710;
wire n_13711, n_13712, n_13713, n_13714, n_13716, n_13717, n_13719,n_13720;
wire n_13721, n_13722, n_13723, n_13724, n_13725, n_13726, n_13727,n_13728;
wire n_13729, n_13730, n_13731, n_13732, n_13733, n_13734, n_13735,n_13736;
wire n_13738, n_13739, n_13740, n_13741, n_13742, n_13743, n_13744,n_13745;
wire n_13748, n_13749, n_13750, n_13751, n_13752, n_13753, n_13754,n_13756;
wire n_13758, n_13759, n_13760, n_13761, n_13762, n_13763, n_13764,n_13765;
wire n_13766, n_13767, n_13768, n_13769, n_13770, n_13771, n_13772,n_13773;
wire n_13774, n_13775, n_13776, n_13777, n_13778, n_13781, n_13782,n_13783;
wire n_13784, n_13786, n_13787, n_13791, n_13795, n_13797, n_13798,n_13799;
wire n_13800, n_13801, n_13802, n_13803, n_13804, n_13805, n_13806,n_13807;
wire n_13809, n_13810, n_13811, n_13812, n_13813, n_13814, n_13815,n_13816;
wire n_13817, n_13818, n_13819, n_13820, n_13822, n_13825, n_13826,n_13827;
wire n_13828, n_13830, n_13834, n_13835, n_13837, n_13838, n_13839,n_13842;
wire n_13843, n_13846, n_13847, n_13848, n_13849, n_13851, n_13852,n_13853;
wire n_13855, n_13857, n_13858, n_13864, n_13871, n_13872, n_13873,n_13875;
wire n_13879, n_13880, n_13881, n_13882, n_13884, n_13885, n_13886,n_13895;
wire n_13896, n_13898, n_13899, n_13900, n_13907, n_13909, n_13910,n_13912;
wire n_13914, n_13915, n_13917, n_13920, n_13921, n_13926, n_13927,n_13928;
wire n_13931, n_13932, n_13935, n_13936, n_13939, n_13940, n_13942,n_13946;
wire n_13947, n_13949, n_13950, n_13951, n_13952, n_13953, n_13954,n_13955;
wire n_13956, n_13957, n_13958, n_13959, n_13960, n_13961, n_13962,n_13963;
wire n_13964, n_13965, n_13966, n_13967, n_13970, n_13971, n_13972,n_13973;
wire n_13974, n_13975, n_13976, n_13977, n_13979, n_13980, n_13982,n_13984;
wire n_13985, n_13986, n_13987, n_13988, n_13989, n_13990, n_13991,n_13992;
wire n_13993, n_13994, n_13995, n_13996, n_13997, n_13998, n_13999,n_14000;
wire n_14001, n_14002, n_14003, n_14004, n_14005, n_14006, n_14007,n_14008;
wire n_14009, n_14010, n_14011, n_14012, n_14013, n_14014, n_14015,n_14017;
wire n_14019, n_14020, n_14021, n_14025, n_14026, n_14027, n_14028,n_14029;
wire n_14031, n_14032, n_14033, n_14034, n_14036, n_14037, n_14038,n_14039;
wire n_14040, n_14041, n_14042, n_14043, n_14044, n_14045, n_14046,n_14047;
wire n_14048, n_14049, n_14050, n_14051, n_14052, n_14053, n_14054,n_14055;
wire n_14056, n_14058, n_14059, n_14060, n_14061, n_14063, n_14064,n_14066;
wire n_14067, n_14068, n_14069, n_14070, n_14074, n_14075, n_14076,n_14077;
wire n_14078, n_14079, n_14080, n_14081, n_14082, n_14084, n_14085,n_14086;
wire n_14087, n_14088, n_14093, n_14094, n_14095, n_14096, n_14097,n_14098;
wire n_14099, n_14100, n_14101, n_14102, n_14105, n_14106, n_14107,n_14108;
wire n_14110, n_14111, n_14112, n_14113, n_14114, n_14115, n_14116,n_14120;
wire n_14121, n_14122, n_14123, n_14125, n_14126, n_14127, n_14128,n_14129;
wire n_14130, n_14131, n_14132, n_14133, n_14134, n_14135, n_14137,n_14138;
wire n_14139, n_14140, n_14141, n_14142, n_14143, n_14145, n_14146,n_14147;
wire n_14148, n_14149, n_14150, n_14151, n_14152, n_14153, n_14154,n_14155;
wire n_14156, n_14157, n_14158, n_14159, n_14160, n_14161, n_14164,n_14165;
wire n_14167, n_14169, n_14170, n_14171, n_14173, n_14175, n_14176,n_14177;
wire n_14179, n_14180, n_14181, n_14182, n_14183, n_14184, n_14185,n_14186;
wire n_14187, n_14188, n_14189, n_14190, n_14191, n_14192, n_14193,n_14194;
wire n_14195, n_14196, n_14198, n_14200, n_14201, n_14202, n_14203,n_14204;
wire n_14205, n_14206, n_14207, n_14208, n_14209, n_14210, n_14213,n_14214;
wire n_14216, n_14217, n_14219, n_14220, n_14221, n_14222, n_14223,n_14225;
wire n_14226, n_14227, n_14228, n_14230, n_14231, n_14232, n_14233,n_14235;
wire n_14236, n_14237, n_14239, n_14240, n_14241, n_14242, n_14243,n_14244;
wire n_14245, n_14246, n_14247, n_14250, n_14251, n_14252, n_14253,n_14254;
wire n_14257, n_14258, n_14259, n_14261, n_14262, n_14263, n_14264,n_14265;
wire n_14266, n_14267, n_14268, n_14269, n_14270, n_14271, n_14272,n_14273;
wire n_14274, n_14275, n_14276, n_14277, n_14279, n_14281, n_14283,n_14284;
wire n_14285, n_14286, n_14288, n_14289, n_14290, n_14291, n_14292,n_14293;
wire n_14294, n_14295, n_14296, n_14297, n_14298, n_14299, n_14301,n_14303;
wire n_14304, n_14306, n_14307, n_14308, n_14309, n_14310, n_14313,n_14314;
wire n_14315, n_14316, n_14317, n_14318, n_14319, n_14320, n_14321,n_14322;
wire n_14323, n_14324, n_14325, n_14326, n_14327, n_14328, n_14329,n_14330;
wire n_14331, n_14332, n_14333, n_14334, n_14336, n_14337, n_14338,n_14340;
wire n_14341, n_14342, n_14343, n_14344, n_14345, n_14346, n_14348,n_14349;
wire n_14350, n_14351, n_14353, n_14354, n_14356, n_14357, n_14358,n_14360;
wire n_14361, n_14362, n_14364, n_14365, n_14366, n_14367, n_14368,n_14369;
wire n_14370, n_14371, n_14372, n_14374, n_14376, n_14377, n_14378,n_14379;
wire n_14380, n_14381, n_14382, n_14383, n_14384, n_14385, n_14386,n_14387;
wire n_14388, n_14390, n_14391, n_14392, n_14393, n_14394, n_14395,n_14396;
wire n_14397, n_14398, n_14399, n_14400, n_14401, n_14402, n_14403,n_14405;
wire n_14406, n_14407, n_14408, n_14409, n_14412, n_14413, n_14414,n_14415;
wire n_14416, n_14417, n_14418, n_14419, n_14420, n_14421, n_14422,n_14424;
wire n_14425, n_14426, n_14427, n_14428, n_14429, n_14430, n_14431,n_14433;
wire n_14434, n_14435, n_14436, n_14437, n_14438, n_14439, n_14440,n_14442;
wire n_14443, n_14444, n_14447, n_14448, n_14450, n_14451, n_14452,n_14454;
wire n_14455, n_14458, n_14459, n_14460, n_14461, n_14462, n_14463,n_14464;
wire n_14466, n_14467, n_14468, n_14469, n_14470, n_14471, n_14472,n_14473;
wire n_14474, n_14475, n_14477, n_14478, n_14479, n_14481, n_14482,n_14483;
wire n_14484, n_14486, n_14487, n_14488, n_14489, n_14490, n_14491,n_14492;
wire n_14493, n_14495, n_14497, n_14498, n_14499, n_14500, n_14501,n_14502;
wire n_14503, n_14505, n_14506, n_14508, n_14510, n_14511, n_14512,n_14513;
wire n_14514, n_14516, n_14517, n_14518, n_14519, n_14520, n_14521,n_14522;
wire n_14523, n_14524, n_14525, n_14526, n_14527, n_14528, n_14529,n_14531;
wire n_14532, n_14533, n_14534, n_14535, n_14536, n_14537, n_14538,n_14540;
wire n_14542, n_14543, n_14544, n_14545, n_14546, n_14547, n_14548,n_14549;
wire n_14551, n_14553, n_14554, n_14555, n_14556, n_14557, n_14558,n_14559;
wire n_14560, n_14561, n_14562, n_14564, n_14565, n_14567, n_14568,n_14569;
wire n_14570, n_14571, n_14573, n_14574, n_14575, n_14577, n_14579,n_14580;
wire n_14581, n_14582, n_14583, n_14585, n_14587, n_14588, n_14589,n_14590;
wire n_14592, n_14593, n_14594, n_14596, n_14597, n_14598, n_14600,n_14601;
wire n_14603, n_14604, n_14605, n_14607, n_14608, n_14610, n_14611,n_14613;
wire n_14615, n_14616, n_14617, n_14619, n_14621, n_14623, n_14624,n_14625;
wire n_14626, n_14627, n_14628, n_14630, n_14633, n_14635, n_14636,n_14637;
wire n_14638, n_14639, n_14640, n_14641, n_14642, n_14643, n_14644,n_14646;
wire n_14647, n_14648, n_14649, n_14650, n_14652, n_14653, n_14655,n_14656;
wire n_14657, n_14658, n_14659, n_14660, n_14661, n_14662, n_14663,n_14666;
wire n_14667, n_14668, n_14669, n_14670, n_14671, n_14672, n_14673,n_14674;
wire n_14675, n_14676, n_14677, n_14678, n_14679, n_14680, n_14681,n_14682;
wire n_14687, n_14689, n_14690, n_14691, n_14692, n_14694, n_14695,n_14696;
wire n_14697, n_14698, n_14700, n_14701, n_14702, n_14704, n_14705,n_14706;
wire n_14707, n_14708, n_14709, n_14712, n_14714, n_14718, n_14719,n_14721;
wire n_14722, n_14723, n_14724, n_14725, n_14726, n_14727, n_14728,n_14729;
wire n_14730, n_14731, n_14734, n_14735, n_14736, n_14737, n_14738,n_14739;
wire n_14740, n_14741, n_14742, n_14743, n_14744, n_14745, n_14746,n_14747;
wire n_14748, n_14749, n_14751, n_14752, n_14754, n_14755, n_14756,n_14757;
wire n_14758, n_14759, n_14760, n_14761, n_14762, n_14763, n_14764,n_14765;
wire n_14766, n_14767, n_14768, n_14769, n_14770, n_14771, n_14772,n_14773;
wire n_14774, n_14776, n_14777, n_14778, n_14779, n_14781, n_14782,n_14783;
wire n_14784, n_14785, n_14786, n_14787, n_14788, n_14789, n_14790,n_14791;
wire n_14792, n_14793, n_14794, n_14795, n_14796, n_14797, n_14798,n_14800;
wire n_14801, n_14802, n_14803, n_14804, n_14805, n_14806, n_14807,n_14808;
wire n_14809, n_14812, n_14813, n_14814, n_14815, n_14816, n_14818,n_14819;
wire n_14821, n_14822, n_14823, n_14824, n_14825, n_14826, n_14827,n_14828;
wire n_14831, n_14832, n_14833, n_14834, n_14835, n_14836, n_14837,n_14839;
wire n_14840, n_14841, n_14842, n_14843, n_14845, n_14846, n_14848,n_14849;
wire n_14850, n_14851, n_14852, n_14853, n_14854, n_14855, n_14856,n_14857;
wire n_14858, n_14859, n_14860, n_14861, n_14862, n_14863, n_14864,n_14865;
wire n_14866, n_14867, n_14868, n_14869, n_14870, n_14872, n_14873,n_14874;
wire n_14875, n_14877, n_14878, n_14879, n_14880, n_14881, n_14882,n_14883;
wire n_14884, n_14885, n_14886, n_14887, n_14888, n_14889, n_14890,n_14892;
wire n_14893, n_14894, n_14895, n_14897, n_14898, n_14899, n_14900,n_14901;
wire n_14902, n_14903, n_14904, n_14905, n_14907, n_14908, n_14909,n_14911;
wire n_14912, n_14913, n_14914, n_14915, n_14917, n_14918, n_14919,n_14921;
wire n_14922, n_14923, n_14925, n_14926, n_14927, n_14928, n_14929,n_14930;
wire n_14931, n_14932, n_14933, n_14934, n_14935, n_14936, n_14937,n_14938;
wire n_14939, n_14940, n_14941, n_14942, n_14943, n_14944, n_14945,n_14946;
wire n_14947, n_14948, n_14949, n_14950, n_14951, n_14952, n_14953,n_14954;
wire n_14955, n_14956, n_14957, n_14958, n_14959, n_14960, n_14961,n_14962;
wire n_14963, n_14964, n_14965, n_14966, n_14967, n_14969, n_14970,n_14972;
wire n_14974, n_14975, n_14976, n_14977, n_14978, n_14979, n_14980,n_14981;
wire n_14983, n_14984, n_14985, n_14986, n_14988, n_14989, n_14990,n_14991;
wire n_14992, n_14993, n_14995, n_14996, n_14997, n_14998, n_14999,n_15000;
wire n_15001, n_15002, n_15003, n_15006, n_15007, n_15008, n_15009,n_15010;
wire n_15011, n_15012, n_15013, n_15014, n_15015, n_15016, n_15018,n_15019;
wire n_15020, n_15021, n_15024, n_15026, n_15027, n_15028, n_15029,n_15033;
wire n_15034, n_15035, n_15036, n_15037, n_15038, n_15039, n_15040,n_15041;
wire n_15042, n_15044, n_15045, n_15046, n_15047, n_15048, n_15050,n_15051;
wire n_15052, n_15053, n_15054, n_15055, n_15056, n_15057, n_15059,n_15061;
wire n_15062, n_15063, n_15064, n_15065, n_15066, n_15067, n_15068,n_15069;
wire n_15070, n_15071, n_15072, n_15073, n_15074, n_15075, n_15076,n_15077;
wire n_15078, n_15079, n_15080, n_15081, n_15082, n_15084, n_15085,n_15086;
wire n_15087, n_15089, n_15090, n_15091, n_15092, n_15094, n_15095,n_15096;
wire n_15098, n_15099, n_15100, n_15101, n_15102, n_15103, n_15104,n_15105;
wire n_15106, n_15107, n_15108, n_15109, n_15110, n_15111, n_15112,n_15113;
wire n_15114, n_15115, n_15116, n_15117, n_15118, n_15119, n_15121,n_15122;
wire n_15123, n_15124, n_15125, n_15126, n_15127, n_15128, n_15129,n_15130;
wire n_15131, n_15132, n_15133, n_15135, n_15136, n_15137, n_15138,n_15139;
wire n_15140, n_15141, n_15142, n_15143, n_15145, n_15146, n_15147,n_15149;
wire n_15151, n_15152, n_15153, n_15154, n_15156, n_15157, n_15159,n_15160;
wire n_15161, n_15163, n_15165, n_15166, n_15168, n_15170, n_15171,n_15172;
wire n_15173, n_15174, n_15175, n_15176, n_15177, n_15178, n_15179,n_15180;
wire n_15181, n_15182, n_15183, n_15184, n_15185, n_15186, n_15187,n_15188;
wire n_15189, n_15190, n_15192, n_15194, n_15195, n_15196, n_15197,n_15199;
wire n_15200, n_15204, n_15205, n_15206, n_15207, n_15208, n_15209,n_15210;
wire n_15211, n_15212, n_15214, n_15216, n_15217, n_15218, n_15219,n_15221;
wire n_15222, n_15223, n_15224, n_15225, n_15226, n_15227, n_15228,n_15229;
wire n_15230, n_15231, n_15232, n_15233, n_15234, n_15235, n_15236,n_15237;
wire n_15238, n_15239, n_15240, n_15241, n_15242, n_15243, n_15244,n_15245;
wire n_15246, n_15247, n_15248, n_15250, n_15252, n_15254, n_15255,n_15256;
wire n_15257, n_15258, n_15259, n_15260, n_15261, n_15262, n_15263,n_15265;
wire n_15266, n_15267, n_15268, n_15269, n_15272, n_15274, n_15275,n_15276;
wire n_15277, n_15278, n_15279, n_15280, n_15281, n_15282, n_15283,n_15284;
wire n_15285, n_15286, n_15287, n_15288, n_15289, n_15291, n_15292,n_15293;
wire n_15294, n_15296, n_15297, n_15298, n_15299, n_15300, n_15301,n_15302;
wire n_15303, n_15304, n_15305, n_15306, n_15307, n_15308, n_15309,n_15310;
wire n_15311, n_15312, n_15313, n_15314, n_15315, n_15316, n_15317,n_15318;
wire n_15319, n_15320, n_15321, n_15322, n_15323, n_15324, n_15325,n_15326;
wire n_15327, n_15328, n_15329, n_15330, n_15332, n_15333, n_15337,n_15339;
wire n_15340, n_15341, n_15342, n_15343, n_15344, n_15345, n_15346,n_15347;
wire n_15348, n_15349, n_15350, n_15351, n_15352, n_15353, n_15354,n_15355;
wire n_15356, n_15357, n_15358, n_15359, n_15360, n_15362, n_15363,n_15365;
wire n_15367, n_15368, n_15370, n_15371, n_15372, n_15374, n_15376,n_15378;
wire n_15379, n_15381, n_15384, n_15386, n_15387, n_15388, n_15389,n_15390;
wire n_15392, n_15393, n_15395, n_15396, n_15397, n_15399, n_15400,n_15402;
wire n_15403, n_15404, n_15411, n_15412, n_15413, n_15414, n_15415,n_15416;
wire n_15418, n_15419, n_15420, n_15421, n_15423, n_15424, n_15425,n_15426;
wire n_15427, n_15428, n_15430, n_15431, n_15432, n_15433, n_15434,n_15435;
wire n_15437, n_15439, n_15440, n_15441, n_15442, n_15443, n_15444,n_15445;
wire n_15447, n_15448, n_15450, n_15451, n_15452, n_15453, n_15456,n_15457;
wire n_15458, n_15460, n_15461, n_15462, n_15463, n_15464, n_15465,n_15466;
wire n_15468, n_15469, n_15472, n_15473, n_15474, n_15475, n_15477,n_15478;
wire n_15479, n_15480, n_15481, n_15482, n_15483, n_15484, n_15485,n_15486;
wire n_15487, n_15488, n_15489, n_15490, n_15491, n_15492, n_15493,n_15495;
wire n_15496, n_15497, n_15498, n_15499, n_15501, n_15502, n_15503,n_15505;
wire n_15506, n_15507, n_15508, n_15509, n_15511, n_15512, n_15513,n_15514;
wire n_15515, n_15516, n_15518, n_15519, n_15522, n_15523, n_15524,n_15527;
wire n_15528, n_15529, n_15530, n_15531, n_15532, n_15533, n_15534,n_15535;
wire n_15536, n_15537, n_15538, n_15539, n_15540, n_15541, n_15542,n_15543;
wire n_15544, n_15545, n_15547, n_15549, n_15551, n_15552, n_15553,n_15554;
wire n_15555, n_15556, n_15557, n_15558, n_15559, n_15561, n_15563,n_15564;
wire n_15566, n_15567, n_15568, n_15569, n_15570, n_15571, n_15572,n_15573;
wire n_15574, n_15575, n_15576, n_15578, n_15579, n_15580, n_15581,n_15582;
wire n_15583, n_15584, n_15585, n_15586, n_15587, n_15588, n_15589,n_15590;
wire n_15591, n_15592, n_15593, n_15595, n_15596, n_15597, n_15598,n_15599;
wire n_15600, n_15601, n_15602, n_15603, n_15604, n_15605, n_15606,n_15608;
wire n_15609, n_15610, n_15611, n_15612, n_15614, n_15615, n_15616,n_15617;
wire n_15620, n_15621, n_15623, n_15625, n_15626, n_15627, n_15628,n_15629;
wire n_15630, n_15631, n_15633, n_15635, n_15636, n_15637, n_15638,n_15640;
wire n_15641, n_15642, n_15644, n_15645, n_15647, n_15648, n_15649,n_15650;
wire n_15652, n_15655, n_15656, n_15657, n_15658, n_15659, n_15660,n_15661;
wire n_15663, n_15667, n_15669, n_15670, n_15673, n_15674, n_15675,n_15676;
wire n_15677, n_15678, n_15680, n_15681, n_15682, n_15683, n_15685,n_15686;
wire n_15687, n_15688, n_15689, n_15690, n_15691, n_15692, n_15693,n_15694;
wire n_15697, n_15698, n_15699, n_15700, n_15701, n_15702, n_15703,n_15704;
wire n_15705, n_15706, n_15707, n_15708, n_15709, n_15710, n_15711,n_15712;
wire n_15713, n_15714, n_15715, n_15717, n_15720, n_15721, n_15722,n_15723;
wire n_15724, n_15725, n_15726, n_15727, n_15729, n_15730, n_15731,n_15732;
wire n_15733, n_15734, n_15735, n_15738, n_15741, n_15742, n_15743,n_15745;
wire n_15748, n_15750, n_15751, n_15752, n_15754, n_15758, n_15759,n_15761;
wire n_15762, n_15764, n_15765, n_15766, n_15767, n_15768, n_15770,n_15773;
wire n_15774, n_15775, n_15776, n_15777, n_15780, n_15781, n_15784,n_15786;
wire n_15788, n_15789, n_15791, n_15792, n_15794, n_15795, n_15796,n_15797;
wire n_15798, n_15799, n_15800, n_15801, n_15802, n_15811, n_15812,n_15813;
wire n_15814, n_15816, n_15817, n_15818, n_15819, n_15821, n_15822,n_15824;
wire n_15825, n_15826, n_15829, n_15830, n_15833, n_15834, n_15835,n_15836;
wire n_15837, n_15838, n_15845, n_15846, n_15847, n_15848, n_15849,n_15850;
wire n_15851, n_15852, n_15853, n_15854, n_15855, n_15856, n_15857,n_15858;
wire n_15859, n_15860, n_15861, n_15862, n_15863, n_15864, n_15865,n_15866;
wire n_15867, n_15868, n_15869, n_15870, n_15871, n_15873, n_15874,n_15875;
wire n_15877, n_15878, n_15879, n_15880, n_15881, n_15882, n_15883,n_15884;
wire n_15886, n_15887, n_15888, n_15890, n_15891, n_15892, n_15893,n_15894;
wire n_15895, n_15896, n_15897, n_15898, n_15900, n_15901, n_15902,n_15903;
wire n_15906, n_15908, n_15909, n_15910, n_15912, n_15913, n_15914,n_15916;
wire n_15917, n_15918, n_15919, n_15920, n_15922, n_15923, n_15924,n_15926;
wire n_15927, n_15930, n_15931, n_15932, n_15934, n_15935, n_15936,n_15937;
wire n_15939, n_15940, n_15941, n_15942, n_15943, n_15944, n_15945,n_15947;
wire n_15948, n_15949, n_15950, n_15951, n_15952, n_15953, n_15954,n_15955;
wire n_15956, n_15958, n_15960, n_15961, n_15963, n_15964, n_15965,n_15966;
wire n_15967, n_15968, n_15969, n_15970, n_15972, n_15976, n_15977,n_15979;
wire n_15982, n_15983, n_15984, n_15985, n_15986, n_15987, n_15988,n_15990;
wire n_15991, n_15992, n_15993, n_15994, n_15996, n_15997, n_15998,n_15999;
wire n_16000, n_16002, n_16003, n_16004, n_16005, n_16006, n_16007,n_16008;
wire n_16009, n_16010, n_16013, n_16014, n_16016, n_16017, n_16018,n_16019;
wire n_16020, n_16022, n_16023, n_16024, n_16027, n_16030, n_16031,n_16032;
wire n_16034, n_16037, n_16038, n_16039, n_16040, n_16041, n_16044,n_16045;
wire n_16046, n_16048, n_16049, n_16050, n_16051, n_16052, n_16053,n_16054;
wire n_16055, n_16057, n_16058, n_16059, n_16061, n_16063, n_16064,n_16065;
wire n_16067, n_16068, n_16069, n_16070, n_16071, n_16072, n_16073,n_16074;
wire n_16075, n_16076, n_16077, n_16078, n_16079, n_16080, n_16081,n_16082;
wire n_16083, n_16084, n_16086, n_16087, n_16089, n_16090, n_16091,n_16092;
wire n_16093, n_16094, n_16095, n_16096, n_16097, n_16098, n_16100,n_16101;
wire n_16102, n_16103, n_16104, n_16106, n_16108, n_16110, n_16111,n_16112;
wire n_16113, n_16115, n_16116, n_16118, n_16119, n_16121, n_16123,n_16124;
wire n_16125, n_16126, n_16127, n_16128, n_16129, n_16130, n_16131,n_16132;
wire n_16133, n_16134, n_16135, n_16137, n_16138, n_16139, n_16140,n_16141;
wire n_16142, n_16143, n_16144, n_16146, n_16149, n_16151, n_16153,n_16154;
wire n_16157, n_16159, n_16161, n_16162, n_16163, n_16164, n_16168,n_16169;
wire n_16172, n_16174, n_16175, n_16176, n_16177, n_16182, n_16183,n_16184;
wire n_16185, n_16186, n_16187, n_16188, n_16195, n_16196, n_16197,n_16198;
wire n_16199, n_16200, n_16204, n_16207, n_16208, n_16209, n_16210,n_16213;
wire n_16215, n_16217, n_16221, n_16223, n_16224, n_16225, n_16226,n_16228;
wire n_16229, n_16236, n_16237, n_16238, n_16240, n_16245, n_16246,n_16249;
wire n_16250, n_16251, n_16253, n_16254, n_16257, n_16259, n_16262,n_16263;
wire n_16264, n_16265, n_16266, n_16267, n_16268, n_16271, n_16272,n_16275;
wire n_16278, n_16279, n_16280, n_16281, n_16282, n_16283, n_16284,n_16285;
wire n_16286, n_16287, n_16288, n_16289, n_16290, n_16291, n_16292,n_16293;
wire n_16294, n_16296, n_16297, n_16298, n_16299, n_16300, n_16301,n_16302;
wire n_16304, n_16306, n_16308, n_16309, n_16310, n_16312, n_16313,n_16314;
wire n_16315, n_16316, n_16317, n_16318, n_16319, n_16320, n_16321,n_16322;
wire n_16323, n_16324, n_16325, n_16326, n_16327, n_16328, n_16329,n_16330;
wire n_16331, n_16332, n_16333, n_16334, n_16336, n_16337, n_16338,n_16339;
wire n_16340, n_16341, n_16342, n_16343, n_16345, n_16346, n_16347,n_16348;
wire n_16349, n_16351, n_16352, n_16354, n_16355, n_16356, n_16357,n_16358;
wire n_16359, n_16360, n_16361, n_16362, n_16364, n_16365, n_16366,n_16367;
wire n_16368, n_16369, n_16371, n_16372, n_16373, n_16374, n_16375,n_16376;
wire n_16377, n_16378, n_16379, n_16380, n_16381, n_16382, n_16383,n_16384;
wire n_16385, n_16386, n_16387, n_16388, n_16389, n_16390, n_16391,n_16392;
wire n_16393, n_16394, n_16395, n_16396, n_16397, n_16398, n_16399,n_16400;
wire n_16401, n_16402, n_16403, n_16404, n_16405, n_16406, n_16407,n_16408;
wire n_16409, n_16410, n_16411, n_16412, n_16413, n_16414, n_16415,n_16416;
wire n_16417, n_16419, n_16420, n_16421, n_16422, n_16423, n_16424,n_16425;
wire n_16426, n_16427, n_16428, n_16429, n_16430, n_16431, n_16432,n_16433;
wire n_16434, n_16435, n_16436, n_16437, n_16439, n_16440, n_16441,n_16442;
wire n_16443, n_16444, n_16445, n_16446, n_16447, n_16448, n_16449,n_16450;
wire n_16452, n_16453, n_16454, n_16455, n_16456, n_16457, n_16459,n_16460;
wire n_16461, n_16462, n_16463, n_16464, n_16465, n_16466, n_16467,n_16468;
wire n_16469, n_16470, n_16471, n_16472, n_16473, n_16474, n_16476,n_16477;
wire n_16478, n_16479, n_16480, n_16481, n_16482, n_16484, n_16485,n_16486;
wire n_16487, n_16488, n_16489, n_16490, n_16491, n_16492, n_16493,n_16494;
wire n_16495, n_16496, n_16497, n_16499, n_16500, n_16501, n_16502,n_16503;
wire n_16504, n_16505, n_16506, n_16507, n_16508, n_16509, n_16510,n_16511;
wire n_16512, n_16513, n_16514, n_16515, n_16517, n_16518, n_16519,n_16520;
wire n_16522, n_16523, n_16524, n_16525, n_16526, n_16527, n_16528,n_16529;
wire n_16530, n_16532, n_16533, n_16534, n_16535, n_16536, n_16537,n_16538;
wire n_16539, n_16540, n_16541, n_16542, n_16543, n_16544, n_16545,n_16548;
wire n_16549, n_16550, n_16551, n_16552, n_16553, n_16554, n_16555,n_16557;
wire n_16558, n_16559, n_16560, n_16561, n_16563, n_16564, n_16565,n_16567;
wire n_16568, n_16569, n_16570, n_16571, n_16572, n_16573, n_16574,n_16575;
wire n_16576, n_16577, n_16578, n_16579, n_16580, n_16581, n_16582,n_16583;
wire n_16584, n_16586, n_16587, n_16588, n_16589, n_16590, n_16592,n_16593;
wire n_16594, n_16595, n_16596, n_16597, n_16599, n_16600, n_16601,n_16602;
wire n_16603, n_16604, n_16605, n_16606, n_16607, n_16608, n_16610,n_16611;
wire n_16612, n_16614, n_16616, n_16617, n_16618, n_16621, n_16622,n_16623;
wire n_16624, n_16625, n_16629, n_16630, n_16633, n_16634, n_16635,n_16636;
wire n_16637, n_16638, n_16639, n_16640, n_16641, n_16642, n_16644,n_16645;
wire n_16646, n_16647, n_16648, n_16649, n_16650, n_16651, n_16652,n_16653;
wire n_16655, n_16656, n_16657, n_16658, n_16659, n_16660, n_16661,n_16663;
wire n_16664, n_16665, n_16666, n_16668, n_16669, n_16670, n_16671,n_16672;
wire n_16673, n_16674, n_16675, n_16676, n_16678, n_16679, n_16680,n_16681;
wire n_16682, n_16683, n_16684, n_16685, n_16686, n_16687, n_16688,n_16689;
wire n_16690, n_16693, n_16694, n_16695, n_16696, n_16700, n_16701,n_16703;
wire n_16704, n_16705, n_16706, n_16707, n_16708, n_16709, n_16711,n_16712;
wire n_16713, n_16714, n_16715, n_16716, n_16717, n_16718, n_16719,n_16720;
wire n_16721, n_16722, n_16724, n_16725, n_16726, n_16727, n_16728,n_16730;
wire n_16731, n_16732, n_16733, n_16737, n_16738, n_16739, n_16740,n_16742;
wire n_16744, n_16745, n_16746, n_16748, n_16749, n_16751, n_16752,n_16753;
wire n_16754, n_16756, n_16757, n_16758, n_16759, n_16761, n_16762,n_16763;
wire n_16764, n_16765, n_16766, n_16767, n_16768, n_16769, n_16772,n_16773;
wire n_16774, n_16775, n_16776, n_16777, n_16778, n_16780, n_16781,n_16782;
wire n_16784, n_16785, n_16786, n_16787, n_16788, n_16789, n_16790,n_16791;
wire n_16792, n_16793, n_16794, n_16796, n_16797, n_16798, n_16800,n_16801;
wire n_16802, n_16805, n_16806, n_16807, n_16808, n_16809, n_16810,n_16811;
wire n_16812, n_16813, n_16816, n_16817, n_16818, n_16820, n_16822,n_16823;
wire n_16825, n_16826, n_16827, n_16828, n_16829, n_16830, n_16832,n_16833;
wire n_16834, n_16835, n_16836, n_16837, n_16840, n_16841, n_16842,n_16843;
wire n_16844, n_16845, n_16848, n_16849, n_16850, n_16851, n_16852,n_16853;
wire n_16854, n_16855, n_16856, n_16857, n_16858, n_16859, n_16860,n_16861;
wire n_16862, n_16863, n_16864, n_16865, n_16867, n_16868, n_16871,n_16873;
wire n_16874, n_16875, n_16877, n_16878, n_16879, n_16880, n_16882,n_16883;
wire n_16884, n_16889, n_16890, n_16891, n_16892, n_16893, n_16894,n_16895;
wire n_16896, n_16897, n_16898, n_16902, n_16903, n_16904, n_16905,n_16906;
wire n_16907, n_16908, n_16909, n_16910, n_16911, n_16912, n_16913,n_16916;
wire n_16917, n_16918, n_16919, n_16920, n_16921, n_16922, n_16924,n_16925;
wire n_16926, n_16927, n_16928, n_16929, n_16931, n_16933, n_16934,n_16935;
wire n_16936, n_16937, n_16938, n_16939, n_16940, n_16941, n_16942,n_16943;
wire n_16944, n_16945, n_16946, n_16947, n_16948, n_16949, n_16950,n_16951;
wire n_16952, n_16954, n_16955, n_16956, n_16958, n_16959, n_16960,n_16962;
wire n_16963, n_16964, n_16965, n_16966, n_16967, n_16968, n_16969,n_16970;
wire n_16972, n_16973, n_16974, n_16976, n_16977, n_16978, n_16979,n_16980;
wire n_16981, n_16982, n_16984, n_16985, n_16986, n_16987, n_16988,n_16989;
wire n_16990, n_16991, n_16992, n_16993, n_16994, n_16995, n_16996,n_16997;
wire n_16998, n_16999, n_17000, n_17001, n_17002, n_17003, n_17004,n_17005;
wire n_17006, n_17007, n_17009, n_17010, n_17011, n_17012, n_17013,n_17014;
wire n_17015, n_17016, n_17017, n_17018, n_17019, n_17020, n_17021,n_17022;
wire n_17023, n_17024, n_17025, n_17026, n_17028, n_17029, n_17030,n_17031;
wire n_17032, n_17033, n_17034, n_17035, n_17036, n_17037, n_17038,n_17039;
wire n_17040, n_17041, n_17042, n_17043, n_17045, n_17046, n_17047,n_17048;
wire n_17049, n_17050, n_17053, n_17054, n_17057, n_17058, n_17059,n_17060;
wire n_17061, n_17062, n_17063, n_17064, n_17065, n_17067, n_17068,n_17069;
wire n_17070, n_17071, n_17072, n_17073, n_17074, n_17076, n_17077,n_17078;
wire n_17080, n_17081, n_17082, n_17083, n_17084, n_17085, n_17086,n_17088;
wire n_17089, n_17090, n_17091, n_17092, n_17093, n_17094, n_17095,n_17096;
wire n_17097, n_17098, n_17099, n_17100, n_17101, n_17102, n_17103,n_17104;
wire n_17105, n_17106, n_17107, n_17108, n_17110, n_17111, n_17112,n_17113;
wire n_17114, n_17115, n_17116, n_17118, n_17119, n_17121, n_17122,n_17123;
wire n_17124, n_17125, n_17126, n_17127, n_17128, n_17129, n_17130,n_17131;
wire n_17133, n_17134, n_17136, n_17137, n_17138, n_17139, n_17140,n_17141;
wire n_17142, n_17143, n_17145, n_17146, n_17147, n_17150, n_17151,n_17152;
wire n_17153, n_17154, n_17155, n_17156, n_17157, n_17158, n_17159,n_17161;
wire n_17162, n_17164, n_17165, n_17167, n_17169, n_17170, n_17172,n_17173;
wire n_17174, n_17175, n_17176, n_17177, n_17178, n_17179, n_17180,n_17181;
wire n_17182, n_17183, n_17184, n_17185, n_17186, n_17187, n_17188,n_17189;
wire n_17191, n_17192, n_17193, n_17195, n_17196, n_17197, n_17198,n_17199;
wire n_17201, n_17203, n_17205, n_17207, n_17208, n_17209, n_17210,n_17211;
wire n_17212, n_17213, n_17214, n_17215, n_17216, n_17217, n_17218,n_17219;
wire n_17220, n_17221, n_17222, n_17223, n_17224, n_17226, n_17227,n_17228;
wire n_17229, n_17230, n_17231, n_17232, n_17233, n_17234, n_17235,n_17236;
wire n_17237, n_17238, n_17239, n_17240, n_17242, n_17243, n_17244,n_17245;
wire n_17246, n_17247, n_17249, n_17250, n_17251, n_17253, n_17254,n_17255;
wire n_17257, n_17258, n_17259, n_17260, n_17261, n_17262, n_17263,n_17265;
wire n_17266, n_17268, n_17269, n_17270, n_17271, n_17272, n_17274,n_17275;
wire n_17277, n_17279, n_17281, n_17283, n_17284, n_17285, n_17286,n_17287;
wire n_17288, n_17289, n_17290, n_17291, n_17292, n_17293, n_17294,n_17295;
wire n_17296, n_17297, n_17298, n_17299, n_17301, n_17302, n_17303,n_17304;
wire n_17305, n_17306, n_17307, n_17308, n_17309, n_17310, n_17311,n_17312;
wire n_17313, n_17314, n_17315, n_17316, n_17317, n_17318, n_17319,n_17320;
wire n_17321, n_17322, n_17323, n_17324, n_17325, n_17326, n_17327,n_17328;
wire n_17329, n_17330, n_17331, n_17332, n_17333, n_17335, n_17337,n_17339;
wire n_17340, n_17341, n_17342, n_17343, n_17344, n_17345, n_17346,n_17347;
wire n_17348, n_17349, n_17350, n_17351, n_17353, n_17354, n_17356,n_17357;
wire n_17358, n_17359, n_17360, n_17361, n_17362, n_17363, n_17364,n_17365;
wire n_17366, n_17367, n_17369, n_17372, n_17373, n_17374, n_17375,n_17376;
wire n_17377, n_17380, n_17381, n_17382, n_17383, n_17384, n_17385,n_17386;
wire n_17387, n_17388, n_17389, n_17390, n_17392, n_17393, n_17395,n_17396;
wire n_17397, n_17399, n_17400, n_17402, n_17404, n_17405, n_17406,n_17408;
wire n_17409, n_17410, n_17411, n_17412, n_17413, n_17414, n_17415,n_17416;
wire n_17417, n_17418, n_17419, n_17421, n_17422, n_17423, n_17424,n_17425;
wire n_17426, n_17427, n_17429, n_17430, n_17431, n_17435, n_17437,n_17438;
wire n_17439, n_17442, n_17443, n_17444, n_17445, n_17446, n_17447,n_17448;
wire n_17449, n_17450, n_17451, n_17453, n_17454, n_17455, n_17456,n_17457;
wire n_17458, n_17459, n_17461, n_17462, n_17465, n_17467, n_17470,n_17472;
wire n_17473, n_17474, n_17477, n_17479, n_17480, n_17481, n_17482,n_17483;
wire n_17484, n_17485, n_17486, n_17487, n_17489, n_17491, n_17493,n_17494;
wire n_17495, n_17496, n_17498, n_17499, n_17500, n_17501, n_17503,n_17504;
wire n_17505, n_17506, n_17507, n_17508, n_17509, n_17510, n_17511,n_17512;
wire n_17514, n_17516, n_17517, n_17519, n_17521, n_17522, n_17523,n_17525;
wire n_17526, n_17527, n_17528, n_17530, n_17531, n_17532, n_17533,n_17535;
wire n_17537, n_17538, n_17539, n_17540, n_17541, n_17542, n_17543,n_17544;
wire n_17545, n_17546, n_17547, n_17548, n_17549, n_17551, n_17552,n_17554;
wire n_17555, n_17556, n_17557, n_17558, n_17559, n_17560, n_17561,n_17562;
wire n_17563, n_17564, n_17565, n_17567, n_17568, n_17569, n_17571,n_17572;
wire n_17573, n_17575, n_17576, n_17577, n_17578, n_17579, n_17580,n_17582;
wire n_17584, n_17585, n_17586, n_17587, n_17588, n_17589, n_17590,n_17591;
wire n_17592, n_17593, n_17594, n_17595, n_17596, n_17597, n_17598,n_17599;
wire n_17600, n_17601, n_17602, n_17604, n_17605, n_17606, n_17607,n_17608;
wire n_17609, n_17610, n_17611, n_17616, n_17617, n_17618, n_17619,n_17620;
wire n_17621, n_17622, n_17623, n_17624, n_17625, n_17626, n_17628,n_17629;
wire n_17630, n_17632, n_17633, n_17634, n_17635, n_17636, n_17638,n_17640;
wire n_17641, n_17642, n_17643, n_17645, n_17646, n_17647, n_17649,n_17650;
wire n_17651, n_17652, n_17653, n_17655, n_17657, n_17658, n_17659,n_17660;
wire n_17665, n_17667, n_17668, n_17669, n_17672, n_17675, n_17676,n_17677;
wire n_17678, n_17679, n_17680, n_17681, n_17682, n_17683, n_17684,n_17685;
wire n_17686, n_17687, n_17688, n_17689, n_17690, n_17691, n_17692,n_17693;
wire n_17694, n_17695, n_17697, n_17698, n_17700, n_17701, n_17702,n_17703;
wire n_17704, n_17705, n_17706, n_17707, n_17708, n_17710, n_17712,n_17713;
wire n_17714, n_17715, n_17716, n_17717, n_17718, n_17719, n_17720,n_17721;
wire n_17722, n_17723, n_17724, n_17725, n_17726, n_17727, n_17728,n_17729;
wire n_17730, n_17731, n_17732, n_17733, n_17734, n_17735, n_17736,n_17737;
wire n_17738, n_17739, n_17740, n_17741, n_17742, n_17743, n_17744,n_17745;
wire n_17746, n_17747, n_17748, n_17749, n_17750, n_17752, n_17753,n_17754;
wire n_17755, n_17756, n_17757, n_17758, n_17759, n_17760, n_17761,n_17762;
wire n_17763, n_17764, n_17765, n_17768, n_17770, n_17771, n_17772,n_17773;
wire n_17774, n_17775, n_17776, n_17777, n_17781, n_17782, n_17783,n_17785;
wire n_17786, n_17787, n_17788, n_17789, n_17790, n_17791, n_17792,n_17793;
wire n_17794, n_17795, n_17796, n_17797, n_17798, n_17799, n_17801,n_17802;
wire n_17803, n_17804, n_17805, n_17806, n_17807, n_17808, n_17809,n_17811;
wire n_17812, n_17813, n_17814, n_17815, n_17816, n_17817, n_17818,n_17819;
wire n_17820, n_17821, n_17822, n_17823, n_17824, n_17825, n_17827,n_17828;
wire n_17830, n_17831, n_17832, n_17833, n_17834, n_17835, n_17836,n_17837;
wire n_17838, n_17839, n_17840, n_17841, n_17842, n_17843, n_17844,n_17845;
wire n_17846, n_17847, n_17848, n_17849, n_17850, n_17851, n_17852,n_17854;
wire n_17856, n_17858, n_17860, n_17861, n_17862, n_17863, n_17864,n_17865;
wire n_17866, n_17867, n_17868, n_17869, n_17872, n_17875, n_17877,n_17879;
wire n_17880, n_17881, n_17882, n_17883, n_17884, n_17886, n_17887,n_17888;
wire n_17889, n_17890, n_17893, n_17894, n_17896, n_17897, n_17898,n_17899;
wire n_17900, n_17901, n_17902, n_17904, n_17906, n_17907, n_17908,n_17910;
wire n_17911, n_17912, n_17914, n_17915, n_17916, n_17918, n_17919,n_17920;
wire n_17921, n_17922, n_17923, n_17924, n_17925, n_17926, n_17927,n_17928;
wire n_17929, n_17930, n_17931, n_17932, n_17933, n_17934, n_17935,n_17936;
wire n_17937, n_17938, n_17939, n_17940, n_17942, n_17943, n_17944,n_17948;
wire n_17950, n_17951, n_17954, n_17955, n_17956, n_17958, n_17960,n_17961;
wire n_17962, n_17963, n_17966, n_17968, n_17969, n_17970, n_17972,n_17973;
wire n_17974, n_17975, n_17977, n_17978, n_17979, n_17980, n_17981,n_17982;
wire n_17983, n_17984, n_17985, n_17986, n_17987, n_17989, n_17990,n_17991;
wire n_17992, n_17993, n_17995, n_17996, n_17997, n_17998, n_17999,n_18000;
wire n_18001, n_18002, n_18003, n_18004, n_18005, n_18007, n_18009,n_18010;
wire n_18011, n_18012, n_18013, n_18014, n_18016, n_18017, n_18018,n_18019;
wire n_18021, n_18023, n_18024, n_18026, n_18027, n_18028, n_18032,n_18033;
wire n_18035, n_18036, n_18037, n_18038, n_18039, n_18040, n_18041,n_18042;
wire n_18043, n_18044, n_18045, n_18046, n_18047, n_18048, n_18049,n_18050;
wire n_18051, n_18052, n_18053, n_18054, n_18057, n_18058, n_18059,n_18060;
wire n_18061, n_18062, n_18063, n_18064, n_18065, n_18066, n_18067,n_18068;
wire n_18069, n_18070, n_18071, n_18073, n_18074, n_18080, n_18081,n_18082;
wire n_18083, n_18084, n_18085, n_18086, n_18087, n_18088, n_18089,n_18090;
wire n_18091, n_18092, n_18093, n_18094, n_18095, n_18096, n_18097,n_18098;
wire n_18099, n_18100, n_18101, n_18102, n_18103, n_18104, n_18105,n_18106;
wire n_18107, n_18108, n_18109, n_18110, n_18111, n_18112, n_18113,n_18114;
wire n_18115, n_18116, n_18117, n_18118, n_18119, n_18120, n_18121,n_18122;
wire n_18123, n_18125, n_18126, n_18127, n_18129, n_18130, n_18134,n_18136;
wire n_18137, n_18138, n_18140, n_18141, n_18142, n_18143, n_18145,n_18147;
wire n_18148, n_18150, n_18151, n_18152, n_18153, n_18154, n_18155,n_18156;
wire n_18157, n_18160, n_18161, n_18162, n_18163, n_18164, n_18168,n_18169;
wire n_18170, n_18172, n_18173, n_18174, n_18176, n_18177, n_18179,n_18181;
wire n_18182, n_18183, n_18184, n_18188, n_18189, n_18192, n_18193,n_18194;
wire n_18195, n_18196, n_18197, n_18199, n_18201, n_18202, n_18203,n_18204;
wire n_18205, n_18206, n_18207, n_18208, n_18209, n_18210, n_18211,n_18212;
wire n_18213, n_18214, n_18215, n_18216, n_18217, n_18219, n_18220,n_18221;
wire n_18224, n_18225, n_18227, n_18228, n_18229, n_18231, n_18232,n_18233;
wire n_18234, n_18235, n_18236, n_18237, n_18238, n_18239, n_18241,n_18242;
wire n_18243, n_18244, n_18245, n_18246, n_18248, n_18249, n_18250,n_18251;
wire n_18252, n_18253, n_18254, n_18255, n_18256, n_18257, n_18258,n_18259;
wire n_18260, n_18261, n_18262, n_18263, n_18264, n_18265, n_18266,n_18267;
wire n_18268, n_18269, n_18270, n_18271, n_18273, n_18274, n_18275,n_18276;
wire n_18277, n_18278, n_18279, n_18280, n_18281, n_18282, n_18283,n_18285;
wire n_18286, n_18287, n_18288, n_18289, n_18290, n_18292, n_18293,n_18294;
wire n_18295, n_18296, n_18297, n_18298, n_18300, n_18301, n_18302,n_18303;
wire n_18304, n_18307, n_18308, n_18309, n_18310, n_18311, n_18312,n_18313;
wire n_18314, n_18316, n_18319, n_18320, n_18321, n_18323, n_18324,n_18325;
wire n_18326, n_18328, n_18329, n_18330, n_18333, n_18334, n_18335,n_18336;
wire n_18337, n_18339, n_18340, n_18341, n_18342, n_18343, n_18344,n_18345;
wire n_18346, n_18347, n_18348, n_18350, n_18351, n_18352, n_18353,n_18354;
wire n_18355, n_18356, n_18357, n_18358, n_18359, n_18360, n_18361,n_18362;
wire n_18363, n_18365, n_18366, n_18367, n_18368, n_18369, n_18370,n_18372;
wire n_18374, n_18375, n_18376, n_18377, n_18379, n_18381, n_18382,n_18383;
wire n_18384, n_18385, n_18386, n_18387, n_18388, n_18390, n_18391,n_18392;
wire n_18393, n_18394, n_18396, n_18397, n_18398, n_18399, n_18400,n_18401;
wire n_18402, n_18403, n_18404, n_18405, n_18406, n_18407, n_18408,n_18409;
wire n_18410, n_18411, n_18412, n_18413, n_18414, n_18415, n_18417,n_18418;
wire n_18419, n_18420, n_18421, n_18422, n_18423, n_18424, n_18425,n_18429;
wire n_18430, n_18431, n_18432, n_18433, n_18434, n_18436, n_18437,n_18438;
wire n_18439, n_18440, n_18441, n_18442, n_18443, n_18445, n_18447,n_18449;
wire n_18450, n_18451, n_18453, n_18454, n_18455, n_18456, n_18457,n_18459;
wire n_18460, n_18462, n_18463, n_18464, n_18465, n_18466, n_18469,n_18470;
wire n_18472, n_18473, n_18474, n_18475, n_18478, n_18479, n_18480,n_18481;
wire n_18483, n_18485, n_18487, n_18488, n_18491, n_18494, n_18496,n_18497;
wire n_18500, n_18502, n_18503, n_18506, n_18508, n_18510, n_18511,n_18512;
wire n_18513, n_18514, n_18515, n_18516, n_18517, n_18518, n_18519,n_18520;
wire n_18521, n_18522, n_18523, n_18524, n_18529, n_18530, n_18533,n_18534;
wire n_18535, n_18536, n_18538, n_18539, n_18540, n_18541, n_18544,n_18545;
wire n_18546, n_18549, n_18551, n_18552, n_18553, n_18554, n_18555,n_18556;
wire n_18557, n_18558, n_18559, n_18561, n_18563, n_18565, n_18567,n_18568;
wire n_18569, n_18570, n_18571, n_18573, n_18574, n_18575, n_18576,n_18577;
wire n_18578, n_18579, n_18580, n_18581, n_18582, n_18583, n_18584,n_18585;
wire n_18586, n_18587, n_18588, n_18590, n_18591, n_18592, n_18593,n_18594;
wire n_18596, n_18597, n_18598, n_18599, n_18601, n_18602, n_18603,n_18604;
wire n_18605, n_18610, n_18611, n_18613, n_18614, n_18615, n_18616,n_18617;
wire n_18618, n_18619, n_18620, n_18621, n_18622, n_18624, n_18626,n_18627;
wire n_18630, n_18631, n_18632, n_18633, n_18634, n_18635, n_18636,n_18640;
wire n_18641, n_18642, n_18643, n_18644, n_18645, n_18647, n_18648,n_18649;
wire n_18651, n_18652, n_18653, n_18654, n_18655, n_18656, n_18658,n_18659;
wire n_18660, n_18661, n_18662, n_18663, n_18664, n_18665, n_18666,n_18668;
wire n_18669, n_18670, n_18671, n_18672, n_18673, n_18674, n_18675,n_18676;
wire n_18678, n_18679, n_18680, n_18681, n_18682, n_18683, n_18684,n_18685;
wire n_18686, n_18687, n_18688, n_18689, n_18690, n_18691, n_18692,n_18694;
wire n_18695, n_18696, n_18697, n_18698, n_18699, n_18700, n_18702,n_18703;
wire n_18704, n_18706, n_18707, n_18708, n_18709, n_18711, n_18712,n_18713;
wire n_18714, n_18715, n_18716, n_18718, n_18719, n_18721, n_18722,n_18723;
wire n_18724, n_18725, n_18728, n_18729, n_18731, n_18732, n_18734,n_18738;
wire n_18739, n_18740, n_18741, n_18744, n_18745, n_18746, n_18747,n_18748;
wire n_18749, n_18750, n_18751, n_18752, n_18753, n_18754, n_18755,n_18756;
wire n_18758, n_18759, n_18760, n_18761, n_18762, n_18763, n_18764,n_18765;
wire n_18766, n_18767, n_18768, n_18771, n_18772, n_18773, n_18774,n_18776;
wire n_18777, n_18778, n_18779, n_18780, n_18781, n_18782, n_18783,n_18784;
wire n_18785, n_18786, n_18788, n_18789, n_18790, n_18792, n_18793,n_18794;
wire n_18795, n_18796, n_18797, n_18799, n_18800, n_18801, n_18802,n_18803;
wire n_18804, n_18806, n_18807, n_18808, n_18809, n_18810, n_18811,n_18812;
wire n_18814, n_18815, n_18816, n_18817, n_18818, n_18819, n_18820,n_18821;
wire n_18822, n_18823, n_18825, n_18826, n_18827, n_18828, n_18829,n_18831;
wire n_18833, n_18834, n_18835, n_18836, n_18838, n_18839, n_18840,n_18841;
wire n_18842, n_18843, n_18844, n_18845, n_18846, n_18847, n_18848,n_18849;
wire n_18850, n_18852, n_18853, n_18854, n_18855, n_18856, n_18859,n_18860;
wire n_18861, n_18862, n_18864, n_18865, n_18866, n_18867, n_18868,n_18869;
wire n_18870, n_18871, n_18873, n_18875, n_18876, n_18878, n_18879,n_18880;
wire n_18881, n_18882, n_18883, n_18884, n_18886, n_18887, n_18888,n_18889;
wire n_18890, n_18891, n_18893, n_18895, n_18896, n_18898, n_18899,n_18900;
wire n_18901, n_18902, n_18903, n_18904, n_18905, n_18906, n_18907,n_18908;
wire n_18910, n_18911, n_18912, n_18913, n_18914, n_18915, n_18916,n_18918;
wire n_18920, n_18921, n_18922, n_18923, n_18925, n_18926, n_18927,n_18928;
wire n_18929, n_18930, n_18931, n_18932, n_18933, n_18934, n_18936,n_18937;
wire n_18938, n_18940, n_18941, n_18942, n_18943, n_18945, n_18946,n_18947;
wire n_18948, n_18949, n_18951, n_18952, n_18953, n_18954, n_18955,n_18957;
wire n_18958, n_18959, n_18960, n_18961, n_18963, n_18964, n_18965,n_18966;
wire n_18967, n_18968, n_18969, n_18970, n_18971, n_18972, n_18973,n_18974;
wire n_18975, n_18978, n_18979, n_18980, n_18982, n_18983, n_18986,n_18988;
wire n_18991, n_18992, n_18993, n_18994, n_18995, n_18996, n_18997,n_18998;
wire n_18999, n_19000, n_19001, n_19002, n_19003, n_19004, n_19006,n_19007;
wire n_19008, n_19009, n_19010, n_19011, n_19012, n_19013, n_19015,n_19016;
wire n_19018, n_19019, n_19020, n_19021, n_19022, n_19023, n_19024,n_19025;
wire n_19026, n_19027, n_19028, n_19030, n_19031, n_19032, n_19033,n_19035;
wire n_19036, n_19037, n_19038, n_19039, n_19040, n_19041, n_19042,n_19043;
wire n_19044, n_19045, n_19046, n_19047, n_19048, n_19049, n_19050,n_19051;
wire n_19052, n_19053, n_19055, n_19057, n_19058, n_19059, n_19060,n_19062;
wire n_19065, n_19068, n_19070, n_19071, n_19072, n_19075, n_19078,n_19079;
wire n_19081, n_19082, n_19083, n_19084, n_19085, n_19086, n_19090,n_19092;
wire n_19094, n_19095, n_19096, n_19097, n_19098, n_19100, n_19101,n_19102;
wire n_19103, n_19104, n_19105, n_19106, n_19107, n_19108, n_19109,n_19110;
wire n_19111, n_19112, n_19113, n_19114, n_19115, n_19116, n_19118,n_19121;
wire n_19123, n_19125, n_19126, n_19127, n_19129, n_19130, n_19131,n_19132;
wire n_19133, n_19134, n_19136, n_19137, n_19138, n_19142, n_19143,n_19144;
wire n_19145, n_19147, n_19148, n_19149, n_19150, n_19151, n_19152,n_19153;
wire n_19154, n_19156, n_19157, n_19158, n_19159, n_19160, n_19161,n_19162;
wire n_19164, n_19165, n_19166, n_19167, n_19168, n_19169, n_19170,n_19172;
wire n_19173, n_19174, n_19175, n_19177, n_19181, n_19182, n_19184,n_19186;
wire n_19187, n_19188, n_19189, n_19190, n_19191, n_19192, n_19194,n_19195;
wire n_19196, n_19198, n_19199, n_19200, n_19202, n_19203, n_19204,n_19205;
wire n_19207, n_19208, n_19210, n_19211, n_19212, n_19213, n_19216,n_19217;
wire n_19218, n_19219, n_19220, n_19221, n_19223, n_19224, n_19225,n_19226;
wire n_19227, n_19228, n_19230, n_19231, n_19232, n_19234, n_19236,n_19237;
wire n_19240, n_19241, n_19242, n_19243, n_19244, n_19245, n_19246,n_19247;
wire n_19248, n_19249, n_19250, n_19251, n_19252, n_19253, n_19255,n_19256;
wire n_19257, n_19258, n_19259, n_19260, n_19261, n_19263, n_19264,n_19266;
wire n_19267, n_19268, n_19270, n_19271, n_19272, n_19273, n_19274,n_19275;
wire n_19276, n_19279, n_19280, n_19281, n_19282, n_19284, n_19285,n_19286;
wire n_19287, n_19288, n_19290, n_19291, n_19292, n_19293, n_19294,n_19295;
wire n_19296, n_19297, n_19298, n_19299, n_19300, n_19301, n_19302,n_19304;
wire n_19307, n_19308, n_19309, n_19310, n_19311, n_19312, n_19313,n_19314;
wire n_19315, n_19318, n_19319, n_19320, n_19321, n_19322, n_19325,n_19327;
wire n_19328, n_19329, n_19330, n_19331, n_19332, n_19333, n_19334,n_19339;
wire n_19340, n_19341, n_19342, n_19344, n_19345, n_19347, n_19348,n_19349;
wire n_19350, n_19351, n_19352, n_19353, n_19354, n_19355, n_19356,n_19358;
wire n_19360, n_19361, n_19362, n_19363, n_19364, n_19365, n_19367,n_19368;
wire n_19369, n_19370, n_19371, n_19372, n_19373, n_19374, n_19375,n_19376;
wire n_19377, n_19379, n_19381, n_19383, n_19384, n_19385, n_19386,n_19388;
wire n_19389, n_19391, n_19392, n_19393, n_19394, n_19395, n_19397,n_19398;
wire n_19400, n_19401, n_19402, n_19404, n_19405, n_19406, n_19407,n_19408;
wire n_19410, n_19411, n_19413, n_19414, n_19415, n_19416, n_19417,n_19418;
wire n_19420, n_19421, n_19422, n_19423, n_19424, n_19427, n_19428,n_19429;
wire n_19430, n_19431, n_19432, n_19433, n_19434, n_19436, n_19438,n_19439;
wire n_19441, n_19442, n_19443, n_19444, n_19445, n_19446, n_19447,n_19448;
wire n_19450, n_19451, n_19452, n_19453, n_19454, n_19455, n_19456,n_19457;
wire n_19458, n_19459, n_19460, n_19461, n_19462, n_19463, n_19464,n_19465;
wire n_19466, n_19467, n_19469, n_19470, n_19471, n_19472, n_19473,n_19474;
wire n_19475, n_19476, n_19477, n_19479, n_19480, n_19481, n_19482,n_19484;
wire n_19485, n_19486, n_19487, n_19490, n_19491, n_19492, n_19495,n_19496;
wire n_19497, n_19498, n_19499, n_19500, n_19502, n_19503, n_19504,n_19508;
wire n_19510, n_19511, n_19515, n_19516, n_19517, n_19518, n_19520,n_19521;
wire n_19522, n_19524, n_19525, n_19526, n_19528, n_19529, n_19530,n_19531;
wire n_19532, n_19533, n_19534, n_19535, n_19536, n_19538, n_19539,n_19540;
wire n_19541, n_19542, n_19543, n_19544, n_19545, n_19547, n_19548,n_19549;
wire n_19550, n_19551, n_19552, n_19553, n_19554, n_19555, n_19556,n_19557;
wire n_19558, n_19559, n_19561, n_19564, n_19565, n_19566, n_19567,n_19568;
wire n_19569, n_19570, n_19571, n_19572, n_19573, n_19574, n_19575,n_19576;
wire n_19577, n_19578, n_19579, n_19580, n_19581, n_19582, n_19583,n_19585;
wire n_19586, n_19587, n_19588, n_19589, n_19590, n_19591, n_19592,n_19593;
wire n_19594, n_19595, n_19596, n_19597, n_19598, n_19599, n_19600,n_19602;
wire n_19604, n_19605, n_19607, n_19608, n_19609, n_19610, n_19611,n_19612;
wire n_19614, n_19617, n_19618, n_19619, n_19620, n_19621, n_19623,n_19626;
wire n_19628, n_19629, n_19630, n_19631, n_19632, n_19635, n_19637,n_19638;
wire n_19639, n_19640, n_19641, n_19643, n_19644, n_19645, n_19646,n_19648;
wire n_19649, n_19650, n_19651, n_19653, n_19654, n_19656, n_19658,n_19659;
wire n_19660, n_19661, n_19662, n_19663, n_19664, n_19665, n_19666,n_19667;
wire n_19669, n_19671, n_19673, n_19674, n_19676, n_19678, n_19679,n_19681;
wire n_19682, n_19683, n_19684, n_19686, n_19687, n_19688, n_19689,n_19690;
wire n_19692, n_19693, n_19696, n_19700, n_19701, n_19702, n_19703,n_19704;
wire n_19707, n_19708, n_19709, n_19710, n_19711, n_19712, n_19715,n_19716;
wire n_19717, n_19718, n_19719, n_19720, n_19721, n_19722, n_19723,n_19725;
wire n_19726, n_19727, n_19730, n_19731, n_19732, n_19735, n_19736,n_19737;
wire n_19738, n_19739, n_19740, n_19741, n_19742, n_19743, n_19746,n_19747;
wire n_19748, n_19749, n_19750, n_19751, n_19752, n_19753, n_19754,n_19755;
wire n_19756, n_19757, n_19759, n_19760, n_19761, n_19762, n_19764,n_19766;
wire n_19767, n_19770, n_19771, n_19773, n_19775, n_19776, n_19778,n_19779;
wire n_19780, n_19781, n_19782, n_19784, n_19786, n_19787, n_19788,n_19790;
wire n_19791, n_19793, n_19794, n_19795, n_19796, n_19797, n_19798,n_19799;
wire n_19800, n_19801, n_19802, n_19803, n_19805, n_19806, n_19807,n_19808;
wire n_19811, n_19812, n_19813, n_19814, n_19815, n_19816, n_19817,n_19818;
wire n_19819, n_19821, n_19822, n_19823, n_19825, n_19827, n_19828,n_19829;
wire n_19830, n_19831, n_19832, n_19833, n_19834, n_19835, n_19836,n_19838;
wire n_19839, n_19841, n_19842, n_19844, n_19845, n_19846, n_19847,n_19848;
wire n_19850, n_19851, n_19852, n_19853, n_19854, n_19855, n_19856,n_19857;
wire n_19860, n_19862, n_19863, n_19864, n_19866, n_19867, n_19868,n_19869;
wire n_19870, n_19872, n_19873, n_19875, n_19877, n_19878, n_19880,n_19881;
wire n_19882, n_19884, n_19885, n_19886, n_19887, n_19889, n_19893,n_19895;
wire n_19896, n_19897, n_19898, n_19900, n_19901, n_19902, n_19904,n_19905;
wire n_19908, n_19909, n_19910, n_19911, n_19914, n_19915, n_19917,n_19918;
wire n_19920, n_19921, n_19922, n_19923, n_19924, n_19925, n_19927,n_19928;
wire n_19929, n_19930, n_19931, n_19932, n_19933, n_19934, n_19935,n_19936;
wire n_19937, n_19938, n_19939, n_19940, n_19941, n_19942, n_19943,n_19944;
wire n_19945, n_19946, n_19947, n_19948, n_19949, n_19950, n_19951,n_19952;
wire n_19953, n_19954, n_19955, n_19956, n_19957, n_19958, n_19959,n_19960;
wire n_19961, n_19963, n_19964, n_19965, n_19966, n_19967, n_19968,n_19969;
wire n_19971, n_19974, n_19976, n_19979, n_19980, n_19981, n_19982,n_19983;
wire n_19985, n_19987, n_19989, n_19990, n_19991, n_19992, n_19993,n_19994;
wire n_19995, n_19996, n_19997, n_19998, n_19999, n_20000, n_20001,n_20002;
wire n_20003, n_20004, n_20005, n_20007, n_20008, n_20009, n_20010,n_20011;
wire n_20012, n_20013, n_20014, n_20015, n_20016, n_20017, n_20018,n_20019;
wire n_20020, n_20021, n_20022, n_20023, n_20024, n_20027, n_20029,n_20030;
wire n_20031, n_20033, n_20034, n_20036, n_20038, n_20039, n_20040,n_20041;
wire n_20042, n_20043, n_20044, n_20045, n_20046, n_20047, n_20049,n_20050;
wire n_20052, n_20053, n_20054, n_20055, n_20056, n_20057, n_20058,n_20059;
wire n_20060, n_20061, n_20062, n_20063, n_20064, n_20065, n_20066,n_20068;
wire n_20071, n_20072, n_20073, n_20074, n_20075, n_20077, n_20078,n_20079;
wire n_20080, n_20081, n_20082, n_20083, n_20084, n_20085, n_20087,n_20088;
wire n_20089, n_20091, n_20092, n_20093, n_20095, n_20096, n_20097,n_20098;
wire n_20099, n_20100, n_20101, n_20102, n_20103, n_20104, n_20105,n_20107;
wire n_20108, n_20109, n_20110, n_20111, n_20112, n_20113, n_20115,n_20116;
wire n_20117, n_20118, n_20119, n_20120, n_20121, n_20122, n_20123,n_20124;
wire n_20126, n_20127, n_20128, n_20130, n_20132, n_20133, n_20134,n_20135;
wire n_20137, n_20138, n_20140, n_20141, n_20143, n_20144, n_20145,n_20148;
wire n_20149, n_20150, n_20152, n_20153, n_20154, n_20155, n_20156,n_20157;
wire n_20158, n_20161, n_20162, n_20163, n_20164, n_20165, n_20166,n_20168;
wire n_20169, n_20171, n_20172, n_20173, n_20175, n_20176, n_20177,n_20178;
wire n_20179, n_20180, n_20181, n_20182, n_20183, n_20184, n_20185,n_20186;
wire n_20187, n_20188, n_20189, n_20190, n_20191, n_20192, n_20193,n_20195;
wire n_20197, n_20198, n_20199, n_20200, n_20202, n_20203, n_20204,n_20205;
wire n_20206, n_20208, n_20211, n_20212, n_20213, n_20214, n_20215,n_20216;
wire n_20217, n_20218, n_20219, n_20221, n_20222, n_20225, n_20226,n_20227;
wire n_20229, n_20230, n_20232, n_20233, n_20234, n_20236, n_20237,n_20239;
wire n_20240, n_20243, n_20245, n_20246, n_20247, n_20248, n_20250,n_20251;
wire n_20256, n_20257, n_20258, n_20259, n_20260, n_20261, n_20262,n_20263;
wire n_20264, n_20265, n_20266, n_20267, n_20268, n_20269, n_20270,n_20271;
wire n_20272, n_20273, n_20274, n_20275, n_20277, n_20278, n_20279,n_20281;
wire n_20282, n_20285, n_20286, n_20287, n_20288, n_20289, n_20290,n_20292;
wire n_20293, n_20294, n_20295, n_20297, n_20298, n_20299, n_20300,n_20301;
wire n_20302, n_20303, n_20304, n_20305, n_20306, n_20307, n_20308,n_20309;
wire n_20310, n_20311, n_20312, n_20313, n_20314, n_20315, n_20316,n_20317;
wire n_20318, n_20319, n_20322, n_20324, n_20325, n_20326, n_20327,n_20328;
wire n_20329, n_20331, n_20332, n_20333, n_20334, n_20335, n_20336,n_20337;
wire n_20338, n_20339, n_20340, n_20341, n_20343, n_20344, n_20346,n_20348;
wire n_20349, n_20351, n_20352, n_20353, n_20357, n_20358, n_20359,n_20360;
wire n_20361, n_20362, n_20363, n_20364, n_20365, n_20367, n_20369,n_20370;
wire n_20371, n_20372, n_20373, n_20374, n_20375, n_20378, n_20380,n_20382;
wire n_20383, n_20384, n_20385, n_20386, n_20387, n_20388, n_20389,n_20392;
wire n_20393, n_20394, n_20396, n_20397, n_20398, n_20399, n_20400,n_20401;
wire n_20403, n_20404, n_20405, n_20406, n_20407, n_20408, n_20410,n_20411;
wire n_20412, n_20416, n_20417, n_20418, n_20419, n_20422, n_20426,n_20428;
wire n_20429, n_20430, n_20431, n_20432, n_20435, n_20437, n_20438,n_20439;
wire n_20441, n_20442, n_20443, n_20444, n_20447, n_20448, n_20450,n_20451;
wire n_20452, n_20453, n_20454, n_20455, n_20456, n_20457, n_20458,n_20460;
wire n_20461, n_20462, n_20463, n_20464, n_20465, n_20466, n_20467,n_20468;
wire n_20469, n_20470, n_20471, n_20472, n_20473, n_20475, n_20476,n_20477;
wire n_20478, n_20480, n_20482, n_20483, n_20484, n_20485, n_20487,n_20488;
wire n_20489, n_20491, n_20493, n_20494, n_20495, n_20496, n_20498,n_20499;
wire n_20500, n_20501, n_20502, n_20503, n_20504, n_20505, n_20506,n_20508;
wire n_20509, n_20511, n_20512, n_20513, n_20515, n_20516, n_20517,n_20518;
wire n_20519, n_20520, n_20521, n_20522, n_20523, n_20524, n_20525,n_20526;
wire n_20527, n_20528, n_20529, n_20530, n_20532, n_20533, n_20534,n_20535;
wire n_20536, n_20537, n_20538, n_20539, n_20540, n_20541, n_20543,n_20544;
wire n_20546, n_20547, n_20548, n_20549, n_20550, n_20551, n_20552,n_20554;
wire n_20555, n_20557, n_20558, n_20560, n_20562, n_20563, n_20564,n_20565;
wire n_20566, n_20567, n_20568, n_20571, n_20572, n_20573, n_20574,n_20575;
wire n_20576, n_20577, n_20578, n_20579, n_20580, n_20581, n_20582,n_20583;
wire n_20584, n_20585, n_20587, n_20590, n_20591, n_20592, n_20593,n_20594;
wire n_20595, n_20596, n_20598, n_20600, n_20601, n_20602, n_20603,n_20604;
wire n_20605, n_20606, n_20607, n_20608, n_20609, n_20610, n_20611,n_20615;
wire n_20616, n_20617, n_20618, n_20619, n_20620, n_20621, n_20622,n_20623;
wire n_20624, n_20625, n_20626, n_20627, n_20628, n_20629, n_20631,n_20632;
wire n_20633, n_20634, n_20635, n_20637, n_20638, n_20639, n_20643,n_20644;
wire n_20645, n_20647, n_20648, n_20650, n_20651, n_20654, n_20656,n_20657;
wire n_20658, n_20659, n_20660, n_20661, n_20662, n_20663, n_20664,n_20667;
wire n_20668, n_20675, n_20677, n_20678, n_20679, n_20680, n_20682,n_20683;
wire n_20684, n_20685, n_20686, n_20688, n_20690, n_20693, n_20694,n_20695;
wire n_20698, n_20699, n_20701, n_20705, n_20706, n_20710, n_20711,n_20713;
wire n_20715, n_20716, n_20717, n_20719, n_20720, n_20721, n_20722,n_20723;
wire n_20724, n_20725, n_20728, n_20729, n_20730, n_20732, n_20733,n_20734;
wire n_20735, n_20737, n_20738, n_20739, n_20742, n_20743, n_20744,n_20745;
wire n_20746, n_20747, n_20748, n_20750, n_20752, n_20753, n_20754,n_20755;
wire n_20756, n_20757, n_20758, n_20759, n_20760, n_20761, n_20762,n_20764;
wire n_20765, n_20766, n_20767, n_20768, n_20770, n_20771, n_20772,n_20775;
wire n_20777, n_20778, n_20780, n_20781, n_20783, n_20784, n_20785,n_20786;
wire n_20791, n_20792, n_20794, n_20795, n_20796, n_20798, n_20802,n_20803;
wire n_20804, n_20805, n_20806, n_20808, n_20809, n_20810, n_20811,n_20814;
wire n_20815, n_20816, n_20818, n_20819, n_20820, n_20821, n_20823,n_20827;
wire n_20828, n_20830, n_20831, n_20832, n_20833, n_20834, n_20835,n_20836;
wire n_20837, n_20838, n_20840, n_20841, n_20842, n_20844, n_20847,n_20849;
wire n_20850, n_20851, n_20852, n_20853, n_20854, n_20855, n_20856,n_20857;
wire n_20858, n_20859, n_20860, n_20861, n_20862, n_20863, n_20864,n_20865;
wire n_20866, n_20867, n_20868, n_20869, n_20870, n_20874, n_20875,n_20878;
wire n_20879, n_20880, n_20882, n_20884, n_20886, n_20888, n_20889,n_20890;
wire n_20891, n_20893, n_20894, n_20896, n_20898, n_20899, n_20900,n_20901;
wire n_20902, n_20903, n_20904, n_20905, n_20906, n_20910, n_20911,n_20912;
wire n_20913, n_20914, n_20916, n_20918, n_20919, n_20921, n_20923,n_20924;
wire n_20925, n_20926, n_20927, n_20928, n_20929, n_20931, n_20932,n_20933;
wire n_20934, n_20935, n_20936, n_20937, n_20938, n_20939, n_20940,n_20941;
wire n_20943, n_20945, n_20946, n_20947, n_20948, n_20949, n_20950,n_20951;
wire n_20952, n_20953, n_20954, n_20955, n_20956, n_20957, n_20958,n_20962;
wire n_20964, n_20965, n_20966, n_20967, n_20968, n_20969, n_20970,n_20971;
wire n_20972, n_20974, n_20976, n_20978, n_20979, n_20980, n_20981,n_20982;
wire n_20984, n_20985, n_20986, n_20987, n_20988, n_20989, n_20990,n_20991;
wire n_20993, n_20994, n_20995, n_20997, n_21000, n_21002, n_21004,n_21005;
wire n_21006, n_21007, n_21008, n_21010, n_21012, n_21014, n_21015,n_21016;
wire n_21018, n_21020, n_21022, n_21023, n_21024, n_21025, n_21027,n_21029;
wire n_21031, n_21034, n_21035, n_21036, n_21037, n_21038, n_21040,n_21041;
wire n_21043, n_21046, n_21047, n_21048, n_21049, n_21050, n_21052,n_21053;
wire n_21054, n_21055, n_21056, n_21057, n_21060, n_21061, n_21065,n_21066;
wire n_21067, n_21068, n_21070, n_21071, n_21072, n_21073, n_21075,n_21076;
wire n_21077, n_21078, n_21079, n_21081, n_21082, n_21083, n_21085,n_21087;
wire n_21092, n_21093, n_21094, n_21095, n_21098, n_21100, n_21101,n_21104;
wire n_21106, n_21108, n_21110, n_21112, n_21113, n_21114, n_21116,n_21118;
wire n_21119, n_21120, n_21121, n_21122, n_21124, n_21125, n_21126,n_21127;
wire n_21128, n_21130, n_21131, n_21132, n_21133, n_21134, n_21135,n_21137;
wire n_21138, n_21139, n_21140, n_21141, n_21142, n_21145, n_21146,n_21147;
wire n_21148, n_21149, n_21150, n_21151, n_21152, n_21153, n_21154,n_21155;
wire n_21156, n_21157, n_21158, n_21159, n_21162, n_21163, n_21164,n_21165;
wire n_21168, n_21169, n_21172, n_21173, n_21174, n_21175, n_21177,n_21179;
wire n_21180, n_21181, n_21183, n_21184, n_21185, n_21186, n_21187,n_21188;
wire n_21189, n_21190, n_21191, n_21192, n_21194, n_21195, n_21196,n_21197;
wire n_21200, n_21201, n_21202, n_21205, n_21207, n_21208, n_21209,n_21210;
wire n_21211, n_21214, n_21215, n_21216, n_21217, n_21218, n_21219,n_21220;
wire n_21222, n_21225, n_21227, n_21228, n_21229, n_21230, n_21233,n_21235;
wire n_21236, n_21238, n_21239, n_21240, n_21241, n_21242, n_21243,n_21246;
wire n_21247, n_21248, n_21249, n_21252, n_21254, n_21256, n_21257,n_21258;
wire n_21259, n_21260, n_21261, n_21262, n_21263, n_21264, n_21265,n_21266;
wire n_21267, n_21268, n_21269, n_21270, n_21271, n_21272, n_21273,n_21274;
wire n_21275, n_21276, n_21278, n_21279, n_21283, n_21284, n_21286,n_21288;
wire n_21289, n_21290, n_21291, n_21292, n_21293, n_21294, n_21295,n_21297;
wire n_21298, n_21300, n_21303, n_21304, n_21306, n_21307, n_21308,n_21312;
wire n_21314, n_21315, n_21316, n_21317, n_21320, n_21323, n_21326,n_21327;
wire n_21328, n_21329, n_21331, n_21332, n_21333, n_21339, n_21340,n_21341;
wire n_21342, n_21343, n_21345, n_21346, n_21348, n_21349, n_21350,n_21352;
wire n_21353, n_21354, n_21355, n_21356, n_21357, n_21358, n_21360,n_21361;
wire n_21362, n_21363, n_21364, n_21366, n_21368, n_21369, n_21370,n_21371;
wire n_21372, n_21373, n_21374, n_21375, n_21376, n_21379, n_21381,n_21382;
wire n_21383, n_21384, n_21386, n_21388, n_21389, n_21390, n_21391,n_21392;
wire n_21393, n_21395, n_21396, n_21398, n_21399, n_21400, n_21404,n_21405;
wire n_21406, n_21409, n_21410, n_21411, n_21412, n_21413, n_21416,n_21417;
wire n_21419, n_21420, n_21422, n_21423, n_21426, n_21427, n_21429,n_21430;
wire n_21431, n_21432, n_21433, n_21434, n_21435, n_21436, n_21437,n_21438;
wire n_21439, n_21442, n_21445, n_21446, n_21447, n_21450, n_21451,n_21452;
wire n_21454, n_21455, n_21458, n_21460, n_21461, n_21462, n_21463,n_21464;
wire n_21465, n_21467, n_21469, n_21470, n_21471, n_21472, n_21473,n_21474;
wire n_21475, n_21476, n_21477, n_21478, n_21479, n_21481, n_21484,n_21485;
wire n_21486, n_21487, n_21492, n_21493, n_21494, n_21495, n_21498,n_21499;
wire n_21501, n_21504, n_21505, n_21506, n_21507, n_21509, n_21511,n_21513;
wire n_21516, n_21517, n_21518, n_21519, n_21520, n_21524, n_21526,n_21530;
wire n_21532, n_21533, n_21535, n_21538, n_21540, n_21549, n_21550,n_21552;
wire n_21553, n_21558, n_21563, n_21566, n_21567, n_21568, n_21569,n_21570;
wire n_21571, n_21573, n_21574, n_21576, n_21577, n_21579, n_21581,n_21583;
wire n_21585, n_21586, n_21587, n_21593, n_21594, n_21597, n_21598,n_21599;
wire n_21601, n_21603, n_21604, n_21605, n_21606, n_21607, n_21608,n_21609;
wire n_21611, n_21613, n_21614, n_21615, n_21616, n_21618, n_21620,n_21622;
wire n_21623, n_21624, n_21625, n_21626, n_21627, n_21629, n_21630,n_21631;
wire n_21632, n_21634, n_21635, n_21637, n_21638, n_21642, n_21647,n_21648;
wire n_21649, n_21651, n_21655, n_21656, n_21657, n_21658, n_21659,n_21660;
wire n_21661, n_21662, n_21663, n_21665, n_21666, n_21668, n_21671,n_21675;
wire n_21676, n_21677, n_21678, n_21680, n_21681, n_21682, n_21683,n_21684;
wire n_21686, n_21687, n_21688, n_21693, n_21694, n_21697, n_21699,n_21700;
wire n_21701, n_21704, n_21705, n_21706, n_21707, n_21708, n_21709,n_21711;
wire n_21712, n_21717, n_21718, n_21723, n_21724, n_21725, n_21727,n_21728;
wire n_21729, n_21730, n_21737, n_21738, n_21739, n_21742, n_21743,n_21747;
wire n_21750, n_21751, n_21754, n_21755, n_21756, n_21757, n_21758,n_21762;
wire n_21764, n_21765, n_21767, n_21769, n_21770, n_21772, n_21779,n_21781;
wire n_21782, n_21784, n_21785, n_21786, n_21792, n_21797, n_21798,n_21800;
wire n_21802, n_21803, n_21806, n_21808, n_21809, n_21810, n_21811,n_21812;
wire n_21813, n_21814, n_21815, n_21816, n_21820, n_21821, n_21822,n_21825;
wire n_21826, n_21827, n_21831, n_21832, n_21834, n_21835, n_21837,n_21839;
wire n_21842, n_21843, n_21844, n_21845, n_21846, n_21847, n_21848,n_21850;
wire n_21852, n_21853, n_21855, n_21857, n_21858, n_21859, n_21860,n_21861;
wire n_21863, n_21865, n_21867, n_21869, n_21870, n_21875, n_21889,n_21891;
wire n_21897, n_21899, n_21901, n_21905, n_21909, n_21910, n_21911,n_21915;
wire n_21917, n_21920, n_21922, n_21923, n_21924, n_21926, n_21927,n_21928;
wire n_21929, n_21930, n_21933, n_21937, n_21938, n_21939, n_21945,n_21954;
wire n_21955, n_21956, n_21959, n_21960, n_21963, n_21970, n_21974,n_21975;
wire n_21976, n_21977, n_21978, n_21979, n_21981, n_21982, n_21983,n_21984;
wire n_21986, n_21991, n_21992, n_21993, n_21995, n_21996, n_21999,n_22000;
wire n_22005, n_22007, n_22008, n_22013, n_22014, n_22015, n_22016,n_22017;
wire n_22020, n_22024, n_22027, n_22028, n_22029, n_22030, n_22033,n_22035;
wire n_22036, n_22041, n_22042, n_22044, n_22046, n_22047, n_22053,n_22054;
wire n_22055, n_22056, n_22057, n_22060, n_22062, n_22063, n_22064,n_22065;
wire n_22066, n_22067, n_22069, n_22070, n_22074, n_22075, n_22076,n_22077;
wire n_22078, n_22079, n_22082, n_22086, n_22089, n_22090, n_22091,n_22092;
wire n_22093, n_22094, n_22099, n_22101, n_22109, n_22111, n_22113,n_22117;
wire n_22118, n_22119, n_22126, n_22128, n_22143, n_22145, n_22146,n_22148;
wire n_22149, n_22150, n_22152, n_22154, n_22156, n_22160, n_22161,n_22163;
wire n_22164, n_22167, n_22168, n_22169, n_22173, n_22174, n_22175,n_22176;
wire n_22178, n_22179, n_22187, n_22189, n_22190, n_22195, n_22196,n_22197;
wire n_22200, n_22203, n_22214, n_22215, n_22218, n_22219, n_22221,n_22222;
wire n_22223, n_22224, n_22229, n_22231, n_22240, n_22246, n_22251,n_22252;
wire n_22259, n_22261, n_22266, n_22267, n_22268, n_22269, n_22270,n_22274;
wire n_22275, n_22277, n_22287, n_22288, n_22289, n_22292, n_22295,n_22297;
wire n_22298, n_22299, n_22301, n_22302, n_22311, n_22313, n_22317,n_22320;
wire n_22325, n_22327, n_22334, n_22339, n_22341, n_22343, n_22348,n_22349;
wire n_22353, n_22356, n_22357, n_22359, n_22361, n_22362, n_22363,n_22371;
wire n_22372, n_22377, n_22378, n_22381, n_22388, n_22389, n_22396,n_22403;
wire n_22405, n_22409, n_22412, n_22413, n_22414, n_22417, n_22418,n_22419;
wire n_22420, n_22422, n_22423, n_22424, n_22425, n_22427, n_22429,n_22431;
wire n_22432, n_22433, n_22434, n_22435, n_22437, n_22441, n_22442,n_22448;
wire n_22451, n_22455, n_22456, n_22462, n_22463, n_22465, n_22467,n_22471;
wire n_22480, n_22482, n_22483, n_22487, n_22488, n_22490, n_22493,n_22496;
wire n_22497, n_22498, n_22500, n_22501, n_22502, n_22503, n_22504,n_22505;
wire n_22507, n_22508, n_22509, n_22511, n_22517, n_22519, n_22521,n_22522;
wire n_22524, n_22525, n_22526, n_22527, n_22528, n_22529, n_22534,n_22535;
wire n_22536, n_22539, n_22546, n_22547, n_22548, n_22549, n_22550,n_22551;
wire n_22554, n_22555, n_22556, n_22557, n_22559, n_22560, n_22563,n_22564;
wire n_22565, n_22566, n_22567, n_22568, n_22569, n_22570, n_22571,n_22572;
wire n_22573, n_22576, n_22578, n_22579, n_22580, n_22581, n_22582,n_22583;
wire n_22584, n_22585, n_22586, n_22587, n_22588, n_22591, n_22592,n_22593;
wire n_22594, n_22595, n_22596, n_22597, n_22598, n_22600, n_22603,n_22605;
wire n_22608, n_22609, n_22618, n_22620, n_22621, n_22622, n_22625,n_22628;
wire n_22631, n_22632, n_22636, n_22638, n_22639, n_22640, n_22641,n_22642;
wire n_22643, n_22644, n_22646, n_22647, n_22648, n_22649, n_22650,n_22651;
wire n_22652, n_22653, n_22654, n_22655, n_22657, n_22660, n_22662,n_22663;
wire n_22665, n_22666, n_22668, n_22671, n_22674, n_22676, n_22678,n_22681;
wire n_22685, n_22686, n_22688, n_22689, n_22691, n_22692, n_22693,n_22694;
wire n_22695, n_22696, n_22697, n_22698, n_22699, n_22700, n_22701,n_22702;
wire n_22703, n_22704, n_22705, n_22708, n_22709, n_22710, n_22711,n_22712;
wire n_22713, n_22714, n_22715, n_22716, n_22717, n_22718, n_22719,n_22721;
wire n_22723, n_22724, n_22725, n_22726, n_22727, n_22728, n_22730,n_22734;
wire n_22735, n_22736, n_22737, n_22738, n_22743, n_22744, n_22745,n_22746;
wire n_22747, n_22748, n_22749, n_22750, n_22751, n_22752, n_22754,n_22755;
wire n_22757, n_22759, n_22762, n_22763, n_22764, n_22765, n_22766,n_22767;
wire n_22768, n_22769, n_22770, n_22772, n_22773, n_22774, n_22775,n_22777;
wire n_22778, n_22779, n_22780, n_22781, n_22782, n_22783, n_22784,n_22785;
wire n_22786, n_22787, n_22788, n_22789, n_22790, n_22793, n_22794,n_22795;
wire n_22796, n_22797, n_22798, n_22799, n_22800, n_22801, n_22802,n_22804;
wire n_22805, n_22807, n_22808, n_22810, n_22811, n_22812, n_22815,n_22816;
wire n_22817, n_22819, n_22820, n_22821, n_22824, n_22826, n_22828,n_22829;
wire n_22830, n_22831, n_22832, n_22833, n_22834, n_22840, n_22841,n_22842;
wire n_22844, n_22847, n_22848, n_22849, n_22851, n_22852, n_22853,n_22854;
wire n_22855, n_22856, n_22859, n_22863, n_22867, n_22868, n_22873,n_22875;
wire n_22876, n_22877, n_22878, n_22880, n_22881, n_22882, n_22886,n_22887;
wire n_22890, n_22891, n_22892, n_22895, n_22899, n_22902, n_22906,n_22909;
wire n_22911, n_22913, n_22914, n_22915, n_22917, n_22918, n_22921,n_22924;
wire n_22928, n_22929, n_22931, n_22932, n_22934, n_22935, n_22936,n_22937;
wire n_22939, n_22940, n_22941, n_22942, n_22943, n_22944, n_22945,n_22949;
wire n_22950, n_22952, n_22953, n_22954, n_22955, n_22956, n_22959,n_22962;
wire n_22963, n_22964, n_22965, n_22967, n_22968, n_22972, n_22973,n_22974;
wire n_22975, n_22976, n_22977, n_22978, n_22979, n_22980, n_22981,n_22982;
wire n_22984, n_22985, n_22986, n_22987, n_22988, n_22989, n_22991,n_22992;
wire n_22993, n_22994, n_22995, n_22996, n_22997, n_22998, n_22999,n_23000;
wire n_23001, n_23002, n_23003, n_23004, n_23005, n_23006, n_23007,n_23008;
wire n_23009, n_23010, n_23011, n_23012, n_23013, n_23014, n_23015,n_23016;
wire n_23017, n_23018, n_23019, n_23021, n_23022, n_23023, n_23024,n_23025;
wire n_23030, n_23031, n_23033, n_23034, n_23036, n_23037, n_23038,n_23039;
wire n_23042, n_23043, n_23044, n_23045, n_23047, n_23048, n_23049,n_23050;
wire n_23051, n_23052, n_23053, n_23054, n_23055, n_23056, n_23058,n_23060;
wire n_23061, n_23062, n_23064, n_23065, n_23066, n_23067, n_23068,n_23069;
wire n_23070, n_23071, n_23072, n_23073, n_23076, n_23077, n_23078,n_23079;
wire n_23080, n_23081, n_23082, n_23083, n_23084, n_23085, n_23086,n_23087;
wire n_23089, n_23090, n_23091, n_23092, n_23093, n_23094, n_23095,n_23096;
wire n_23098, n_23099, n_23100, n_23103, n_23105, n_23106, n_23107,n_23109;
wire n_23110, n_23111, n_23114, n_23115, n_23116, n_23117, n_23118,n_23119;
wire n_23120, n_23121, n_23122, n_23131, n_23135, n_23138, n_23139,n_23140;
wire n_23141, n_23143, n_23144, n_23145, n_23147, n_23154, n_23155,n_23156;
wire n_23157, n_23158, n_23159, n_23160, n_23161, n_23162, n_23163,n_23165;
wire n_23166, n_23167, n_23168, n_23169, n_23170, n_23171, n_23173,n_23174;
wire n_23176, n_23177, n_23179, n_23180, n_23181, n_23182, n_23183,n_23184;
wire n_23185, n_23187, n_23188, n_23189, n_23190, n_23191, n_23192,n_23193;
wire n_23195, n_23196, n_23198, n_23200, n_23202, n_23204, n_23205,n_23206;
wire n_23210, n_23211, n_23213, n_23215, n_23216, n_23217, n_23219,n_23221;
wire n_23222, n_23223, n_23224, n_23225, n_23226, n_23227, n_23228,n_23230;
wire n_23231, n_23232, n_23233, n_23234, n_23235, n_23236, n_23237,n_23238;
wire n_23239, n_23240, n_23241, n_23242, n_23244, n_23246, n_23247,n_23248;
wire n_23249, n_23250, n_23251, n_23252, n_23253, n_23254, n_23255,n_23256;
wire n_23257, n_23258, n_23259, n_23260, n_23261, n_23263, n_23264,n_23265;
wire n_23266, n_23267, n_23269, n_23270, n_23271, n_23274, n_23275,n_23276;
wire n_23277, n_23278, n_23279, n_23280, n_23281, n_23283, n_23284,n_23285;
wire n_23286, n_23287, n_23288, n_23289, n_23290, n_23291, n_23292,n_23294;
wire n_23295, n_23296, n_23297, n_23299, n_23301, n_23303, n_23304,n_23305;
wire n_23306, n_23307, n_23308, n_23309, n_23310, n_23311, n_23312,n_23313;
wire n_23314, n_23316, n_23317, n_23318, n_23319, n_23320, n_23322,n_23323;
wire n_23324, n_23326, n_23327, n_23328, n_23329, n_23330, n_23331,n_23332;
wire n_23333, n_23334, n_23335, n_23336, n_23337, n_23338, n_23340,n_23341;
wire n_23342, n_23343, n_23344, n_23345, n_23346, n_23347, n_23348,n_23350;
wire n_23351, n_23352, n_23353, n_23354, n_23355, n_23356, n_23357,n_23358;
wire n_23360, n_23361, n_23362, n_23363, n_23364, n_23366, n_23367,n_23369;
wire n_23373, n_23374, n_23375, n_23376, n_23377, n_23378, n_23379,n_23380;
wire n_23382, n_23383, n_23384, n_23385, n_23386, n_23387, n_23389,n_23390;
wire n_23391, n_23392, n_23393, n_23394, n_23395, n_23396, n_23397,n_23398;
wire n_23399, n_23400, n_23401, n_23402, n_23403, n_23405, n_23406,n_23407;
wire n_23408, n_23409, n_23410, n_23411, n_23412, n_23414, n_23415,n_23416;
wire n_23417, n_23418, n_23419, n_23422, n_23423, n_23424, n_23425,n_23429;
wire n_23431, n_23432, n_23434, n_23435, n_23440, n_23441, n_23442,n_23444;
wire n_23445, n_23446, n_23448, n_23451, n_23452, n_23454, n_23455,n_23456;
wire n_23457, n_23458, n_23468, n_23469, n_23470, n_23471, n_23472,n_23473;
wire n_23474, n_23475, n_23476, n_23480, n_23481, n_23482, n_23483,n_23484;
wire n_23485, n_23486, n_23487, n_23488, n_23489, n_23490, n_23491,n_23493;
wire n_23494, n_23495, n_23496, n_23497, n_23498, n_23499, n_23500,n_23501;
wire n_23502, n_23503, n_23507, n_23510, n_23512, n_23514, n_23515,n_23516;
wire n_23517, n_23518, n_23519, n_23522, n_23523, n_23525, n_23527,n_23528;
wire n_23531, n_23532, n_23533, n_23534, n_23535, n_23537, n_23539,n_23541;
wire n_23543, n_23544, n_23545, n_23546, n_23547, n_23548, n_23549,n_23550;
wire n_23551, n_23552, n_23553, n_23554, n_23555, n_23556, n_23557,n_23558;
wire n_23559, n_23560, n_23561, n_23562, n_23563, n_23564, n_23565,n_23566;
wire n_23567, n_23568, n_23569, n_23570, n_23571, n_23573, n_23574,n_23575;
wire n_23576, n_23577, n_23579, n_23580, n_23581, n_23583, n_23584,n_23585;
wire n_23586, n_23587, n_23588, n_23589, n_23590, n_23591, n_23592,n_23593;
wire n_23594, n_23595, n_23596, n_23597, n_23598, n_23599, n_23600,n_23601;
wire n_23602, n_23603, n_23604, n_23605, n_23606, n_23607, n_23609,n_23610;
wire n_23611, n_23613, n_23614, n_23615, n_23616, n_23617, n_23618,n_23619;
wire n_23620, n_23621, n_23622, n_23623, n_23625, n_23626, n_23627,n_23628;
wire n_23629, n_23630, n_23631, n_23633, n_23634, n_23635, n_23636,n_23637;
wire n_23638, n_23639, n_23640, n_23643, n_23644, n_23646, n_23649,n_23650;
wire n_23652, n_23653, n_23656, n_23657, n_23659, n_23661, n_23662,n_23663;
wire n_23664, n_23667, n_23668, n_23669, n_23670, n_23671, n_23673,n_23674;
wire n_23675, n_23676, n_23677, n_23678, n_23679, n_23680, n_23681,n_23683;
wire n_23684, n_23686, n_23687, n_23688, n_23689, n_23690, n_23692,n_23693;
wire n_23694, n_23695, n_23696, n_23697, n_23698, n_23700, n_23701,n_23702;
wire n_23703, n_23704, n_23706, n_23707, n_23708, n_23709, n_23710,n_23711;
wire n_23712, n_23713, n_23714, n_23715, n_23716, n_23718, n_23720,n_23722;
wire n_23723, n_23724, n_23725, n_23726, n_23727, n_23728, n_23729,n_23730;
wire n_23731, n_23732, n_23733, n_23734, n_23735, n_23736, n_23737,n_23738;
wire n_23739, n_23740, n_23741, n_23742, n_23743, n_23744, n_23745,n_23746;
wire n_23747, n_23748, n_23749, n_23751, n_23752, n_23753, n_23754,n_23755;
wire n_23756, n_23757, n_23758, n_23759, n_23760, n_23761, n_23762,n_23763;
wire n_23765, n_23766, n_23769, n_23770, n_23771, n_23772, n_23773,n_23774;
wire n_23775, n_23777, n_23778, n_23779, n_23780, n_23781, n_23782,n_23783;
wire n_23784, n_23785, n_23786, n_23788, n_23789, n_23790, n_23791,n_23792;
wire n_23793, n_23794, n_23795, n_23796, n_23797, n_23798, n_23802,n_23803;
wire n_23804, n_23805, n_23806, n_23809, n_23810, n_23811, n_23817,n_23819;
wire n_23820, n_23822, n_23824, n_23826, n_23827, n_23828, n_23829,n_23838;
wire n_23839, n_23840, n_23841, n_23842, n_23843, n_23844, n_23845,n_23846;
wire n_23847, n_23848, n_23849, n_23850, n_23851, n_23852, n_23853,n_23854;
wire n_23858, n_23859, n_23860, n_23861, n_23862, n_23863, n_23864,n_23865;
wire n_23866, n_23867, n_23868, n_23869, n_23871, n_23872, n_23873,n_23878;
wire n_23879, n_23880, n_23881, n_23882, n_23883, n_23884, n_23885,n_23886;
wire n_23887, n_23888, n_23889, n_23890, n_23891, n_23892, n_23893,n_23894;
wire n_23895, n_23896, n_23897, n_23898, n_23899, n_23900, n_23901,n_23902;
wire n_23903, n_23904, n_23905, n_23906, n_23907, n_23908, n_23909,n_23910;
wire n_23912, n_23914, n_23915, n_23916, n_23917, n_23918, n_23919,n_23920;
wire n_23921, n_23922, n_23923, n_23924, n_23925, n_23926, n_23927,n_23928;
wire n_23929, n_23930, n_23932, n_23933, n_23934, n_23935, n_23936,n_23937;
wire n_23938, n_23939, n_23940, n_23941, n_23942, n_23943, n_23945,n_23946;
wire n_23947, n_23948, n_23949, n_23950, n_23951, n_23952, n_23954,n_23955;
wire n_23956, n_23958, n_23959, n_23960, n_23962, n_23963, n_23964,n_23965;
wire n_23966, n_23967, n_23968, n_23971, n_23972, n_23975, n_23976,n_23977;
wire n_23978, n_23979, n_23980, n_23981, n_23982, n_23983, n_23984,n_23985;
wire n_23986, n_23987, n_23989, n_23990, n_23991, n_23992, n_23993,n_23994;
wire n_23996, n_23997, n_23998, n_23999, n_24000, n_24001, n_24002,n_24003;
wire n_24004, n_24005, n_24006, n_24007, n_24008, n_24009, n_24010,n_24011;
wire n_24012, n_24013, n_24014, n_24015, n_24016, n_24017, n_24019,n_24021;
wire n_24022, n_24023, n_24026, n_24027, n_24028, n_24029, n_24030,n_24031;
wire n_24032, n_24033, n_24034, n_24035, n_24036, n_24037, n_24038,n_24039;
wire n_24040, n_24041, n_24042, n_24043, n_24044, n_24045, n_24046,n_24047;
wire n_24048, n_24049, n_24050, n_24051, n_24052, n_24053, n_24054,n_24055;
wire n_24056, n_24057, n_24058, n_24059, n_24060, n_24062, n_24063,n_24064;
wire n_24065, n_24066, n_24067, n_24068, n_24069, n_24070, n_24071,n_24072;
wire n_24073, n_24075, n_24076, n_24077, n_24078, n_24079, n_24080,n_24082;
wire n_24083, n_24084, n_24085, n_24087, n_24088, n_24089, n_24090,n_24091;
wire n_24092, n_24093, n_24094, n_24095, n_24096, n_24097, n_24098,n_24099;
wire n_24100, n_24101, n_24102, n_24103, n_24104, n_24105, n_24108,n_24109;
wire n_24110, n_24111, n_24112, n_24113, n_24114, n_24115, n_24116,n_24118;
wire n_24120, n_24121, n_24122, n_24123, n_24124, n_24125, n_24126,n_24127;
wire n_24128, n_24129, n_24130, n_24131, n_24132, n_24133, n_24134,n_24135;
wire n_24136, n_24137, n_24138, n_24139, n_24140, n_24141, n_24142,n_24143;
wire n_24144, n_24145, n_24147, n_24148, n_24149, n_24150, n_24151,n_24152;
wire n_24153, n_24154, n_24155, n_24156, n_24157, n_24158, n_24159,n_24160;
wire n_24161, n_24163, n_24165, n_24166, n_24167, n_24168, n_24169,n_24170;
wire n_24171, n_24172, n_24173, n_24174, n_24175, n_24176, n_24177,n_24178;
wire n_24179, n_24180, n_24181, n_24182, n_24183, n_24184, n_24185,n_24186;
wire n_24187, n_24188, n_24189, n_24192, n_24193, n_24194, n_24195,n_24196;
wire n_24197, n_24198, n_24199, n_24200, n_24201, n_24202, n_24204,n_24205;
wire n_24206, n_24207, n_24208, n_24209, n_24210, n_24211, n_24212,n_24213;
wire n_24214, n_24215, n_24217, n_24218, n_24219, n_24220, n_24222,n_24223;
wire n_24224, n_24226, n_24227, n_24228, n_24229, n_24230, n_24231,n_24232;
wire n_24233, n_24234, n_24235, n_24236, n_24237, n_24238, n_24239,n_24240;
wire n_24241, n_24242, n_24243, n_24245, n_24247, n_24248, n_24249,n_24251;
wire n_24252, n_24253, n_24254, n_24255, n_24256, n_24257, n_24258,n_24259;
wire n_24260, n_24261, n_24262, n_24263, n_24264, n_24265, n_24266,n_24267;
wire n_24268, n_24269, n_24270, n_24271, n_24272, n_24273, n_24275,n_24276;
wire n_24277, n_24278, n_24279, n_24280, n_24281, n_24283, n_24284,n_24285;
wire n_24287, n_24288, n_24289, n_24293, n_24294, n_24295, n_24296,n_24297;
wire n_24298, n_24299, n_24300, n_24301, n_24302, n_24303, n_24304,n_24305;
wire n_24306, n_24307, n_24308, n_24309, n_24310, n_24311, n_24312,n_24313;
wire n_24314, n_24315, n_24316, n_24318, n_24319, n_24321, n_24322,n_24323;
wire n_24324, n_24325, n_24326, n_24327, n_24328, n_24329, n_24330,n_24331;
wire n_24332, n_24333, n_24335, n_24337, n_24338, n_24340, n_24341,n_24342;
wire n_24343, n_24344, n_24345, n_24346, n_24347, n_24349, n_24350,n_24351;
wire n_24352, n_24353, n_24355, n_24357, n_24358, n_24359, n_24360,n_24361;
wire n_24362, n_24363, n_24364, n_24365, n_24366, n_24367, n_24369,n_24370;
wire n_24371, n_24372, n_24373, n_24374, n_24375, n_24376, n_24378,n_24379;
wire n_24380, n_24381, n_24382, n_24383, n_24384, n_24385, n_24386,n_24387;
wire n_24390, n_24391, n_24392, n_24393, n_24394, n_24395, n_24396,n_24397;
wire n_24398, n_24400, n_24401, n_24402, n_24403, n_24404, n_24405,n_24406;
wire n_24407, n_24408, n_24409, n_24410, n_24411, n_24412, n_24413,n_24414;
wire n_24415, n_24416, n_24417, n_24418, n_24419, n_24420, n_24421,n_24422;
wire n_24423, n_24424, n_24425, n_24426, n_24427, n_24428, n_24430,n_24433;
wire n_24435, n_24436, n_24437, n_24438, n_24439, n_24440, n_24441,n_24442;
wire n_24443, n_24444, n_24445, n_24446, n_24447, n_24448, n_24449,n_24450;
wire n_24451, n_24452, n_24453, n_24454, n_24455, n_24456, n_24457,n_24458;
wire n_24459, n_24460, n_24461, n_24462, n_24463, n_24464, n_24465,n_24466;
wire n_24467, n_24468, n_24469, n_24471, n_24472, n_24473, n_24475,n_24476;
wire n_24478, n_24479, n_24480, n_24481, n_24482, n_24483, n_24484,n_24485;
wire n_24486, n_24487, n_24488, n_24489, n_24490, n_24491, n_24492,n_24496;
wire n_24497, n_24498, n_24501, n_24502, n_24505, n_24506, n_24507,n_24508;
wire n_24509, n_24510, n_24511, n_24512, n_24514, n_24515, n_24516,n_24517;
wire n_24518, n_24519, n_24520, n_24521, n_24522, n_24523, n_24524,n_24525;
wire n_24526, n_24527, n_24528, n_24529, n_24530, n_24532, n_24533,n_24534;
wire n_24535, n_24536, n_24537, n_24538, n_24539, n_24540, n_24541,n_24542;
wire n_24543, n_24544, n_24545, n_24547, n_24548, n_24549, n_24550,n_24551;
wire n_24552, n_24553, n_24554, n_24555, n_24556, n_24557, n_24558,n_24559;
wire n_24560, n_24561, n_24562, n_24563, n_24564, n_24565, n_24566,n_24568;
wire n_24570, n_24571, n_24573, n_24574, n_24575, n_24576, n_24577,n_24578;
wire n_24579, n_24580, n_24581, n_24582, n_24583, n_24584, n_24585,n_24586;
wire n_24587, n_24588, n_24589, n_24590, n_24591, n_24592, n_24593,n_24594;
wire n_24595, n_24596, n_24597, n_24598, n_24599, n_24600, n_24601,n_24602;
wire n_24603, n_24604, n_24605, n_24606, n_24607, n_24608, n_24609,n_24610;
wire n_24611, n_24612, n_24613, n_24614, n_24615, n_24616, n_24617,n_24618;
wire n_24619, n_24620, n_24621, n_24622, n_24623, n_24624, n_24625,n_24626;
wire n_24627, n_24628, n_24629, n_24630, n_24631, n_24632, n_24633,n_24634;
wire n_24635, n_24636, n_24637, n_24638, n_24639, n_24640, n_24641,n_24642;
wire n_24643, n_24644, n_24645, n_24646, n_24647, n_24648, n_24649,n_24650;
wire n_24651, n_24652, n_24653, n_24654, n_24655, n_24659, n_24660,n_24661;
wire n_24662, n_24666, n_24667, n_24668, n_24669, n_24670, n_24671,n_24672;
wire n_24673, n_24674, n_24675, n_24676, n_24677, n_24678, n_24679,n_24680;
wire n_24681, n_24682, n_24683, n_24684, n_24685, n_24686, n_24687,n_24688;
wire n_24689, n_24690, n_24691, n_24692, n_24693, n_24694, n_24695,n_24696;
wire n_24697, n_24698, n_24699, n_24700, n_24701, n_24702, n_24703,n_24704;
wire n_24705, n_24706, n_24707, n_24708, n_24709, n_24710, n_24711,n_24712;
wire n_24713, n_24714, n_24715, n_24717, n_24718, n_24719, n_24720,n_24721;
wire n_24722, n_24723, n_24724, n_24725, n_24726, n_24727, n_24728,n_24729;
wire n_24730, n_24731, n_24733, n_24734, n_24735, n_24736, n_24737,n_24738;
wire n_24739, n_24740, n_24741, n_24742, n_24743, n_24745, n_24746,n_24747;
wire n_24749, n_24750, n_24751, n_24752, n_24753, n_24754, n_24755,n_24756;
wire n_24757, n_24758, n_24759, n_24760, n_24761, n_24763, n_24764,n_24765;
wire n_24766, n_24768, n_24769, n_24770, n_24771, n_24772, n_24773,n_24775;
wire n_24776, n_24777, n_24778, n_24779, n_24780, n_24781, n_24782,n_24783;
wire n_24784, n_24785, n_24786, n_24787, n_24788, n_24789, n_24790,n_24791;
wire n_24792, n_24793, n_24794, n_24795, n_24796, n_24797, n_24798,n_24799;
wire n_24800, n_24801, n_24802, n_24804, n_24805, n_24806, n_24807,n_24808;
wire n_24809, n_24810, n_24811, n_24812, n_24813, n_24814, n_24815,n_24816;
wire n_24817, n_24818, n_24819, n_24820, n_24821, n_24822, n_24823,n_24824;
wire n_24825, n_24826, n_24827, n_24830, n_24831, n_24832, n_24833,n_24834;
wire n_24835, n_24836, n_24837, n_24838, n_24839, n_24840, n_24841,n_24842;
wire n_24843, n_24844, n_24845, n_24847, n_24848, n_24849, n_24850,n_24851;
wire n_24852, n_24853, n_24854, n_24855, n_24856, n_24857, n_24858,n_24859;
wire n_24860, n_24861, n_24862, n_24863, n_24864, n_24865, n_24866,n_24868;
wire n_24869, n_24870, n_24871, n_24872, n_24873, n_24874, n_24875,n_24876;
wire n_24877, n_24878, n_24879, n_24880, n_24881, n_24882, n_24883,n_24884;
wire n_24885, n_24886, n_24887, n_24888, n_24889, n_24890, n_24891,n_24892;
wire n_24893, n_24894, n_24895, n_24896, n_24897, n_24898, n_24899,n_24901;
wire n_24902, n_24903, n_24904, n_24905, n_24906, n_24907, n_24908,n_24909;
wire n_24910, n_24911, n_24912, n_24913, n_24914, n_24915, n_24916,n_24918;
wire n_24919, n_24920, n_24921, n_24922, n_24923, n_24924, n_24925,n_24926;
wire n_24927, n_24929, n_24930, n_24931, n_24932, n_24933, n_24934,n_24935;
wire n_24936, n_24937, n_24938, n_24939, n_24940, n_24941, n_24943,n_24944;
wire n_24945, n_24946, n_24947, n_24948, n_24949, n_24950, n_24951,n_24952;
wire n_24953, n_24954, n_24955, n_24956, n_24957, n_24958, n_24959,n_24960;
wire n_24961, n_24962, n_24963, n_24964, n_24965, n_24966, n_24967,n_24968;
wire n_24969, n_24972, n_24973, n_24974, n_24975, n_24976, n_24977,n_24978;
wire n_24979, n_24980, n_24981, n_24982, n_24983, n_24984, n_24985,n_24986;
wire n_24987, n_24988, n_24989, n_24990, n_24991, n_24992, n_24993,n_24994;
wire n_24995, n_24996, n_24997, n_24998, n_24999, n_25000, n_25001,n_25002;
wire n_25003, n_25004, n_25005, n_25006, n_25007, n_25008, n_25009,n_25010;
wire n_25011, n_25012, n_25013, n_25014, n_25015, n_25016, n_25017,n_25018;
wire n_25019, n_25020, n_25021, n_25022, n_25023, n_25024, n_25025,n_25026;
wire n_25027, n_25028, n_25029, n_25030, n_25031, n_25032, n_25033,n_25034;
wire n_25035, n_25039, n_25040, n_25041, n_25042, n_25043, n_25044,n_25045;
wire n_25046, n_25047, n_25049, n_25050, n_25051, n_25052, n_25053,n_25054;
wire n_25055, n_25056, n_25057, n_25058, n_25059, n_25060, n_25061,n_25062;
wire n_25063, n_25064, n_25065, n_25066, n_25067, n_25071, n_25072,n_25073;
wire n_25074, n_25075, n_25076, n_25077, n_25078, n_25079, n_25080,n_25081;
wire n_25082, n_25083, n_25084, n_25085, n_25086, n_25087, n_25088,n_25089;
wire n_25090, n_25091, n_25092, n_25093, n_25094, n_25095, n_25096,n_25097;
wire n_25098, n_25099, n_25100, n_25101, n_25102, n_25103, n_25104,n_25105;
wire n_25106, n_25107, n_25108, n_25109, n_25110, n_25111, n_25112,n_25113;
wire n_25114, n_25115, n_25116, n_25117, n_25118, n_25119, n_25120,n_25121;
wire n_25122, n_25123, n_25124, n_25125, n_25126, n_25127, n_25128,n_25129;
wire n_25130, n_25131, n_25132, n_25133, n_25134, n_25135, n_25136,n_25137;
wire n_25138, n_25139, n_25140, n_25141, n_25143, n_25144, n_25145,n_25146;
wire n_25147, n_25148, n_25149, n_25150, n_25151, n_25152, n_25153,n_25154;
wire n_25155, n_25156, n_25157, n_25159, n_25160, n_25161, n_25162,n_25163;
wire n_25164, n_25165, n_25167, n_25168, n_25169, n_25170, n_25171,n_25172;
wire n_25174, n_25175, n_25176, n_25177, n_25178, n_25179, n_25180,n_25181;
wire n_25182, n_25183, n_25184, n_25185, n_25187, n_25188, n_25191,n_25192;
wire n_25193, n_25194, n_25196, n_25197, n_25198, n_25200, n_25202,n_25203;
wire n_25204, n_25205, n_25206, n_25207, n_25208, n_25209, n_25210,n_25211;
wire n_25213, n_25214, n_25215, n_25216, n_25217, n_25218, n_25219,n_25220;
wire n_25221, n_25222, n_25223, n_25226, n_25227, n_25228, n_25229,n_25230;
wire n_25231, n_25232, n_25233, n_25234, n_25235, n_25236, n_25237,n_25238;
wire n_25239, n_25240, n_25241, n_25242, n_25243, n_25244, n_25245,n_25246;
wire n_25247, n_25248, n_25249, n_25250, n_25251, n_25252, n_25253,n_25254;
wire n_25255, n_25256, n_25262, n_25263, n_25264, n_25265, n_25267,n_25268;
wire n_25269, n_25271, n_25272, n_25273, n_25274, n_25275, n_25276,n_25277;
wire n_25278, n_25281, n_25282, n_25283, n_25285, n_25286, n_25288,n_25289;
wire n_25290, n_25291, n_25292, n_25293, n_25294, n_25295, n_25296,n_25297;
wire n_25298, n_25299, n_25300, n_25301, n_25302, n_25303, n_25304,n_25305;
wire n_25306, n_25307, n_25308, n_25309, n_25310, n_25311, n_25313,n_25314;
wire n_25315, n_25316, n_25317, n_25318, n_25319, n_25320, n_25321,n_25322;
wire n_25323, n_25324, n_25325, n_25327, n_25328, n_25329, n_25330,n_25331;
wire n_25332, n_25333, n_25334, n_25335, n_25336, n_25337, n_25338,n_25339;
wire n_25340, n_25341, n_25342, n_25343, n_25344, n_25345, n_25346,n_25347;
wire n_25348, n_25349, n_25350, n_25351, n_25352, n_25353, n_25354,n_25355;
wire n_25356, n_25357, n_25358, n_25359, n_25360, n_25361, n_25362,n_25364;
wire n_25365, n_25366, n_25367, n_25368, n_25369, n_25370, n_25371,n_25372;
wire n_25373, n_25374, n_25375, n_25376, n_25377, n_25378, n_25379,n_25380;
wire n_25381, n_25382, n_25383, n_25384, n_25385, n_25386, n_25387,n_25388;
wire n_25389, n_25390, n_25391, n_25392, n_25393, n_25394, n_25395,n_25396;
wire n_25397, n_25398, n_25399, n_25400, n_25401, n_25402, n_25403,n_25404;
wire n_25405, n_25406, n_25407, n_25408, n_25409, n_25410, n_25411,n_25412;
wire n_25414, n_25415, n_25416, n_25418, n_25419, n_25420, n_25421,n_25422;
wire n_25423, n_25424, n_25425, n_25426, n_25427, n_25428, n_25429,n_25430;
wire n_25431, n_25432, n_25433, n_25434, n_25435, n_25436, n_25437,n_25438;
wire n_25439, n_25440, n_25453, n_25454, n_25455, n_25456, n_25457,n_25460;
wire n_25463, n_25467, n_25468, n_25476, n_25477, n_25478, n_25481,n_25482;
wire n_25483, n_25484, n_25487, n_25488, n_25496, n_25497, n_25502,n_25503;
wire n_25504, n_25506, n_25507, n_25508, n_25511, n_25512, n_25515,n_25516;
wire n_25517, n_25518, n_25522, n_25523, n_25526, n_25535, n_25536,n_25537;
wire n_25542, n_25543, n_25546, n_25547, n_25550, n_25551, n_25563,n_25564;
wire n_25565, n_25571, n_25578, n_25579, n_25580, n_25581, n_25582,n_25583;
wire n_25584, n_25585, n_25589, n_25590, n_25591, n_25592, n_25596,n_25597;
wire n_25598, n_25599, n_25600, n_25601, n_25602, n_25603, n_25610,n_25611;
wire n_25612, n_25613, n_25614, n_25615, n_25616, n_25617, n_25618,n_25621;
wire n_25622, n_25623, n_25624, n_25626, n_25627, n_25628, n_25629,n_25631;
wire n_25632, n_25635, n_25636, n_25637, n_25638, n_25639, n_25640,n_25641;
wire n_25642, n_25643, n_25652, n_25653, n_25654, n_25659, n_25660,n_25664;
wire n_25665, n_25666, n_25667, n_25668, n_25669, n_25672, n_25673,n_25675;
wire n_25676, n_25677, n_25678, n_25679, n_25685, n_25686, n_25690,n_25691;
wire n_25695, n_25696, n_25697, n_25700, n_25701, n_25702, n_25703,n_25704;
wire n_25705, n_25706, n_25707, n_25708, n_25709, n_25710, n_25711,n_25714;
wire n_25715, n_25717, n_25718, n_25719, n_25720, n_25721, n_25722,n_25725;
wire n_25726, n_25727, n_25728, n_25729, n_25730, n_25731, n_25732,n_25733;
wire n_25734, n_25735, n_25736, n_25737, n_25738, n_25739, n_25741,n_25744;
wire n_25745, n_25746, n_25747, n_25758, n_25759, n_25760, n_25763,n_25768;
wire n_25769, n_25770, n_25771, n_25772, n_25773, n_25774, n_25775,n_25776;
wire n_25777, n_25780, n_25781, n_25782, n_25783, n_25785, n_25786,n_25787;
wire n_25788, n_25789, n_25790, n_25791, n_25796, n_25799, n_25800,n_25801;
wire n_25802, n_25803, n_25804, n_25806, n_25808, n_25809, n_25810,n_25811;
wire n_25812, n_25813, n_25816, n_25817, n_25820, n_25821, n_25822,n_25823;
wire n_25824, n_25825, n_25826, n_25827, n_25828, n_25833, n_25834,n_25837;
wire n_25838, n_25848, n_25850, n_25855, n_25856, n_25857, n_25858,n_25860;
wire n_25861, n_25862, n_25863, n_25864, n_25865, n_25866, n_25876,n_25877;
wire n_25878, n_25880, n_25881, n_25882, n_25883, n_25884, n_25885,n_25886;
wire n_25887, n_25888, n_25889, n_25890, n_25891, n_25893, n_25894,n_25895;
wire n_25896, n_25897, n_25898, n_25899, n_25901, n_25902, n_25907,n_25911;
wire n_25916, n_25917, n_25918, n_25919, n_25922, n_25923, n_25924,n_25925;
wire n_25926, n_25936, n_25937, n_25938, n_25939, n_25940, n_25941,n_25942;
wire n_25943, n_25944, n_25945, n_25946, n_25947, n_25948, n_25949,n_25950;
wire n_25951, n_25953, n_25954, n_25955, n_25956, n_25957, n_25958,n_25959;
wire n_25960, n_25961, n_25963, n_25965, n_25991, n_25992, n_25994,n_25995;
wire n_25996, n_25997, n_25998, n_25999, n_26000, n_26007, n_26011,n_26012;
wire n_26013, n_26015, n_26016, n_26017, n_26018, n_26019, n_26020,n_26021;
wire n_26022, n_26024, n_26025, n_26026, n_26027, n_26028, n_26029,n_26030;
wire n_26032, n_26033, n_26034, n_26035, n_26036, n_26037, n_26038,n_26039;
wire n_26040, n_26041, n_26042, n_26043, n_26044, n_26045, n_26047,n_26048;
wire n_26050, n_26051, n_26052, n_26053, n_26054, n_26055, n_26056,n_26057;
wire n_26058, n_26059, n_26060, n_26061, n_26062, n_26063, n_26064,n_26065;
wire n_26066, n_26068, n_26069, n_26070, n_26071, n_26073, n_26074,n_26075;
wire n_26076, n_26077, n_26078, n_26079, n_26080, n_26081, n_26083,n_26085;
wire n_26086, n_26087, n_26088, n_26089, n_26090, n_26091, n_26092,n_26093;
wire n_26094, n_26095, n_26096, n_26097, n_26098, n_26100, n_26101,n_26102;
wire n_26103, n_26104, n_26129, n_26130, n_26132, n_26133, n_26134,n_26135;
wire n_26137, n_26138, n_26139, n_26140, n_26142, n_26143, n_26144,n_26145;
wire n_26156, n_26159, n_26160, n_26162, n_26163, n_26164, n_26165,n_26166;
wire n_26167, n_26168, n_26169, n_26172, n_26173, n_26174, n_26175,n_26176;
wire n_26177, n_26178, n_26180, n_26185, n_26192, n_26194, n_26197,n_26198;
wire n_26199, n_26200, n_26201, n_26202, n_26203, n_26204, n_26211,n_26212;
wire n_26213, n_26214, n_26215, n_26216, n_26217, n_26218, n_26219,n_26220;
wire n_26221, n_26222, n_26223, n_26224, n_26225, n_26226, n_26227,n_26228;
wire n_26229, n_26230, n_26231, n_26232, n_26233, n_26234, n_26236,n_26237;
wire n_26238, n_26239, n_26240, n_26241, n_26242, n_26243, n_26244,n_26245;
wire n_26246, n_26247, n_26248, n_26249, n_26250, n_26251, n_26252,n_26253;
wire n_26261, n_26262, n_26263, n_26264, n_26266, n_26267, n_26268,n_26269;
wire n_26270, n_26271, n_26272, n_26273, n_26276, n_26277, n_26278,n_26279;
wire n_26281, n_26282, n_26284, n_26285, n_26286, n_26287, n_26297,n_26298;
wire n_26299, n_26300, n_26301, n_26302, n_26303, n_26306, n_26307,n_26308;
wire n_26309, n_26310, n_26311, n_26312, n_26313, n_26314, n_26315,n_26316;
wire n_26317, n_26318, n_26319, n_26322, n_26323, n_26324, n_26325,n_26326;
wire n_26327, n_26350, n_26356, n_26357, n_26358, n_26360, n_26361,n_26362;
wire n_26363, n_26364, n_26365, n_26366, n_26367, n_26368, n_26369,n_26370;
wire n_26371, n_26372, n_26374, n_26375, n_26376, n_26377, n_26379,n_26380;
wire n_26381, n_26382, n_26383, n_26384, n_26385, n_26386, n_26388,n_26393;
wire n_26394, n_26395, n_26396, n_26398, n_26399, n_26400, n_26401,n_26402;
wire n_26403, n_26404, n_26405, n_26406, n_26410, n_26411, n_26414,n_26416;
wire n_26417, n_26418, n_26419, n_26420, n_26421, n_26422, n_26423,n_26424;
wire n_26425, n_26426, n_26427, n_26428, n_26429, n_26430, n_26432,n_26433;
wire n_26434, n_26435, n_26436, n_26437, n_26438, n_26439, n_26440,n_26441;
wire n_26456, n_26457, n_26458, n_26461, n_26464, n_26465, n_26466,n_26467;
wire n_26468, n_26469, n_26470, n_26472, n_26473, n_26474, n_26476,n_26477;
wire n_26478, n_26479, n_26480, n_26481, n_26482, n_26483, n_26485,n_26486;
wire n_26488, n_26489, n_26490, n_26491, n_26492, n_26493, n_26494,n_26495;
wire n_26496, n_26497, n_26498, n_26499, n_26500, n_26501, n_26503,n_26504;
wire n_26505, n_26506, n_26507, n_26508, n_26509, n_26510, n_26511,n_26512;
wire n_26514, n_26515, n_26516, n_26517, n_26518, n_26519, n_26521,n_26522;
wire n_26523, n_26524, n_26525, n_26526, n_26527, n_26528, n_26529,n_26530;
wire n_26531, n_26532, n_26533, n_26534, n_26535, n_26536, n_26537,n_26539;
wire n_26540, n_26541, n_26542, n_26543, n_26546, n_26547, n_26549,n_26550;
wire n_26553, n_26555, n_26556, n_26597, n_26601, n_26602, n_26603,n_26613;
wire n_26614, n_26615, n_26616, n_26617, n_26618, n_26619, n_26621,n_26622;
wire n_26623, n_26624, n_26625, n_26627, n_26628, n_26629, n_26630,n_26631;
wire n_26632, n_26633, n_26634, n_26637, n_26638, n_26639, n_26640,n_26646;
wire n_26654, n_26657, n_26661, n_26662, n_26663, n_26665, n_26666,n_26667;
wire n_26668, n_26669, n_26670, n_26671, n_26672, n_26673, n_26674,n_26675;
wire n_26676, n_26677, n_26678, n_26679, n_26680, n_26682, n_26683,n_26684;
wire n_26685, n_26686, n_26687, n_26689, n_26690, n_26691, n_26692,n_26694;
wire n_26695, n_26696, n_26697, n_26698, n_26700, n_26701, n_26702,n_26703;
wire n_26704, n_26705, n_26706, n_26707, n_26708, n_26709, n_26710,n_26713;
wire n_26715, n_26716, n_26720, n_26721, n_26724, n_26725, n_26726,n_26727;
wire n_26728, n_26729, n_26730, n_26731, n_26732, n_26733, n_26734,n_26735;
wire n_26736, n_26737, n_26738, n_26739, n_26740, n_26741, n_26742,n_26743;
wire n_26744, n_26745, n_26746, n_26747, n_26748, n_26749, n_26750,n_26751;
wire n_26775, n_26776, n_26777, n_26778, n_26779, n_26780, n_26781,n_26782;
wire n_26783, n_26784, n_26786, n_26787, n_26788, n_26789, n_26790,n_26791;
wire n_26792, n_26795, n_26796, n_26797, n_26798, n_26799, n_26800,n_26801;
wire n_26802, n_26814, n_26815, n_26816, n_26817, n_26818, n_26819,n_26820;
wire n_26821, n_26822, n_26826, n_26827, n_26828, n_26829, n_26830,n_26831;
wire n_26832, n_26833, n_26834, n_26836, n_26837, n_26838, n_26839,n_26840;
wire n_26841, n_26842, n_26843, n_26844, n_26846, n_26848, n_26849,n_26850;
wire n_26851, n_26853, n_26854, n_26855, n_26858, n_26863, n_26864,n_26865;
wire n_26866, n_26867, n_26868, n_26869, n_26870, n_26871, n_26872,n_26873;
wire n_26874, n_26877, n_26878, n_26879, n_26880, n_26881, n_26882,n_26883;
wire n_26885, n_26887, n_26888, n_26889, n_26890, n_26891, n_26893,n_26894;
wire n_26895, n_26896, n_26897, n_26898, n_26899, n_26900, n_26901,n_26902;
wire n_26903, n_26904, n_26905, n_26906, n_26907, n_26908, n_26909,n_26910;
wire n_26911, n_26912, n_26913, n_26914, n_26915, n_26916, n_26918,n_26919;
wire n_26920, n_26921, n_26922, n_26923, n_26924, n_26926, n_26927,n_26928;
wire n_26929, n_26930, n_26931, n_26937, n_26938, n_26939, n_26940,n_26941;
wire n_26942, n_26943, n_26944, n_26945, n_26946, n_26947, n_26948,n_26949;
wire n_26950, n_26951, n_26952, n_26954, n_26955, n_26956, n_26957,n_26958;
wire n_26960, n_26961, n_26962, n_26963, n_26964, n_26965, n_26966,n_26967;
wire n_26969, n_26970, n_26971, n_26972, n_26973, n_26974, n_26975,n_26976;
wire n_26977, n_26978, n_26979, n_26980, n_26981, n_26982, n_26983,n_26984;
wire n_26985, n_26986, n_26987, n_26989, n_26990, n_26991, n_26992,n_26993;
wire n_26994, n_26995, n_26996, n_26997, n_26998, n_27000, n_27002,n_27003;
wire n_27004, n_27005, n_27007, n_27008, n_27009, n_27010, n_27011,n_27012;
wire n_27013, n_27014, n_27015, n_27018, n_27019, n_27020, n_27021,n_27022;
wire n_27023, n_27024, n_27025, n_27028, n_27029, n_27030, n_27031,n_27032;
wire n_27033, n_27034, n_27035, n_27036, n_27037, n_27038, n_27039,n_27040;
wire n_27041, n_27042, n_27043, n_27044, n_27045, n_27046, n_27047,n_27048;
wire n_27049, n_27051, n_27053, n_27054, n_27055, n_27056, n_27057,n_27058;
wire n_27059, n_27060, n_27061, n_27063, n_27065, n_27066, n_27067,n_27068;
wire n_27069, n_27070, n_27071, n_27072, n_27075, n_27076, n_27077,n_27080;
wire n_27081, n_27082, n_27083, n_27084, n_27085, n_27089, n_27090,n_27096;
wire n_27097, n_27098, n_27099, n_27100, n_27104, n_27105, n_27106,n_27107;
wire n_27108, n_27109, n_27111, n_27112, n_27113, n_27114, n_27116,n_27117;
wire n_27118, n_27119, n_27120, n_27121, n_27122, n_27124, n_27126,n_27127;
wire n_27128, n_27130, n_27131, n_27132, n_27133, n_27135, n_27136,n_27137;
wire n_27138, n_27139, n_27140, n_27141, n_27142, n_27143, n_27144,n_27145;
wire n_27147, n_27151, n_27152, n_27153, n_27154, n_27155, n_27156,n_27157;
wire n_27160, n_27161, n_27162, n_27177, n_27178, n_27179, n_27182,n_27185;
wire n_27186, n_27187, n_27188, n_27189, n_27190, n_27191, n_27192,n_27193;
wire n_27194, n_27195, n_27196, n_27197, n_27198, n_27199, n_27202,n_27203;
wire n_27204, n_27206, n_27207, n_27208, n_27209, n_27210, n_27211,n_27213;
wire n_27214, n_27215, n_27216, n_27217, n_27218, n_27219, n_27220,n_27222;
wire n_27223, n_27224, n_27225, n_27227, n_27228, n_27229, n_27230,n_27231;
wire n_27232, n_27233, n_27234, n_27235, n_27236, n_27237, n_27238,n_27239;
wire n_27240, n_27241, n_27242, n_27243, n_27244, n_27245, n_27246,n_27247;
wire n_27248, n_27260, n_27261, n_27262, n_27263, n_27264, n_27265,n_27266;
wire n_27267, n_27268, n_27269, n_27271, n_27272, n_27273, n_27282,n_27287;
wire n_27288, n_27289, n_27290, n_27294, n_27296, n_27297, n_27298,n_27300;
wire n_27301, n_27302, n_27303, n_27304, n_27305, n_27306, n_27307,n_27308;
wire n_27309, n_27310, n_27311, n_27312, n_27313, n_27314, n_27315,n_27316;
wire n_27317, n_27318, n_27319, n_27320, n_27321, n_27322, n_27323,n_27334;
wire n_27335, n_27336, n_27339, n_27340, n_27341, n_27342, n_27344,n_27345;
wire n_27346, n_27347, n_27348, n_27350, n_27351, n_27352, n_27353,n_27355;
wire n_27356, n_27357, n_27358, n_27359, n_27360, n_27361, n_27362,n_27363;
wire n_27364, n_27365, n_27366, n_27367, n_27368, n_27369, n_27370,n_27371;
wire n_27372, n_27373, n_27375, n_27377, n_27379, n_27380, n_27381,n_27382;
wire n_27384, n_27385, n_27386, n_27387, n_27388, n_27389, n_27390,n_27391;
wire n_27392, n_27393, n_27396, n_27397, n_27398, n_27399, n_27401,n_27403;
wire n_27405, n_27406, n_27407, n_27408, n_27409, n_27410, n_27411,n_27412;
wire n_27413, n_27418, n_27419, n_27420, n_27421, n_27422, n_27423,n_27424;
wire n_27425, n_27426, n_27427, n_27428, n_27429, n_27430, n_27431,n_27432;
wire n_27433, n_27434, n_27435, n_27436, n_27437, n_27438, n_27439,n_27440;
wire n_27441, n_27442, n_27444, n_27445, n_27446, n_27447, n_27448,n_27449;
wire n_27450, n_27451, n_27452, n_27453, n_27454, n_27455, n_27456,n_27457;
wire n_27458, n_27459, n_27460, n_27461, n_27462, n_27463, n_27464,n_27465;
wire n_27466, n_27467, n_27468, n_27470, n_27471, n_27472, n_27473,n_27474;
wire n_27475, n_27478, n_27479, n_27480, n_27481, n_27483, n_27485,n_27486;
wire n_27487, n_27488, n_27489, n_27490, n_27491, n_27492, n_27493,n_27494;
wire n_27495, n_27496, n_27500, n_27501, n_27502, n_27503, n_27504,n_27505;
wire n_27508, n_27509, n_27510, n_27513, n_27514, n_27515, n_27516,n_27517;
wire n_27518, n_27519, n_27520, n_27521, n_27522, n_27523, n_27524,n_27525;
wire n_27526, n_27527, n_27528, n_27529, n_27531, n_27532, n_27533,n_27534;
wire n_27535, n_27536, n_27537, n_27552, n_27553, n_27554, n_27556,n_27557;
wire n_27558, n_27559, n_27560, n_27561, n_27562, n_27563, n_27564,n_27565;
wire n_27566, n_27569, n_27570, n_27571, n_27572, n_27573, n_27574,n_27585;
wire n_27586, n_27587, n_27588, n_27589, n_27592, n_27593, n_27594,n_27595;
wire n_27596, n_27598, n_27599, n_27600, n_27601, n_27603, n_27604,n_27605;
wire n_27606, n_27607, n_27608, n_27609, n_27610, n_27611, n_27612,n_27614;
wire n_27615, n_27616, n_27617, n_27618, n_27619, n_27620, n_27622,n_27623;
wire n_27624, n_27627, n_27640, n_27641, n_27642, n_27643, n_27645,n_27646;
wire n_27650, n_27652, n_27655, n_27656, n_27657, n_27658, n_27659,n_27660;
wire n_27661, n_27663, n_27664, n_27665, n_27666, n_27668, n_27669,n_27671;
wire n_27672, n_27673, n_27674, n_27675, n_27676, n_27677, n_27678,n_27679;
wire n_27681, n_27682, n_27683, n_27684, n_27686, n_27687, n_27688,n_27690;
wire n_27691, n_27692, n_27693, n_27694, n_27695, n_27696, n_27697,n_27699;
wire n_27700, n_27701, n_27702, n_27703, n_27704, n_27705, n_27706,n_27707;
wire n_27708, n_27709, n_27710, n_27711, n_27712, n_27713, n_27714,n_27715;
wire n_27716, n_27717, n_27718, n_27720, n_27722, n_27723, n_27724,n_27725;
wire n_27726, n_27727, n_27728, n_27729, n_27730, n_27731, n_27732,n_27735;
wire n_27736, n_27737, n_27738, n_27739, n_27740, n_27741, n_27744,n_27745;
wire n_27746, n_27747, n_27751, n_27752, n_27753, n_27757, n_27778,n_27779;
wire n_27780, n_27781, n_27782, n_27783, n_27784, n_27785, n_27786,n_27787;
wire n_27788, n_27789, n_27790, n_27791, n_27792, n_27793, n_27794,n_27795;
wire n_27797, n_27798, n_27799, n_27800, n_27801, n_27802, n_27803,n_27804;
wire n_27805, n_27806, n_27807, n_27809, n_27810, n_27811, n_27812,n_27814;
wire n_27815, n_27816, n_27817, n_27819, n_27821, n_27822, n_27823,n_27825;
wire n_27826, n_27828, n_27829, n_27830, n_27831, n_27833, n_27834,n_27835;
wire n_27836, n_27840, n_27841, n_27842, n_27843, n_27844, n_27845,n_27846;
wire n_27847, n_27848, n_27849, n_27850, n_27851, n_27853, n_27854,n_27855;
wire n_27856, n_27872, n_27873, n_27874, n_27875, n_27876, n_27884,n_27885;
wire n_27886, n_27887, n_27889, n_27890, n_27891, n_27892, n_27893,n_27894;
wire n_27896, n_27897, n_27898, n_27899, n_27900, n_27901, n_27904,n_27905;
wire n_27906, n_27907, n_27908, n_27909, n_27910, n_27911, n_27912,n_27913;
wire n_27914, n_27915, n_27916, n_27917, n_27918, n_27919, n_27939,n_27940;
wire n_27941, n_27942, n_27943, n_27944, n_27945, n_27946, n_27947,n_27948;
wire n_27949, n_27950, n_27951, n_27952, n_27953, n_27954, n_27955,n_27956;
wire n_27957, n_27963, n_27964, n_27965, n_27966, n_27969, n_27970,n_27983;
wire n_27984, n_27985, n_27987, n_27988, n_27990, n_27991, n_28018,n_28019;
wire n_28020, n_28021, n_28022, n_28023, n_28024, n_28025, n_28026,n_28027;
wire n_28028, n_28029, n_28030, n_28031, n_28032, n_28035, n_28036,n_28037;
wire n_28038, n_28039, n_28040, n_28041, n_28042, n_28045, n_28046,n_28047;
wire n_28048, n_28049, n_28050, n_28051, n_28052, n_28053, n_28054,n_28055;
wire n_28057, n_28060, n_28061, n_28062, n_28063, n_28064, n_28065,n_28066;
wire n_28067, n_28068, n_28069, n_28070, n_28071, n_28072, n_28073,n_28074;
wire n_28075, n_28076, n_28077, n_28078, n_28079, n_28080, n_28109,n_28110;
wire n_28111, n_28112, n_28113, n_28114, n_28115, n_28116, n_28117,n_28118;
wire n_28119, n_28120, n_28121, n_28122, n_28123, n_28124, n_28125,n_28126;
wire n_28127, n_28128, n_28129, n_28130, n_28131, n_28132, n_28133,n_28134;
wire n_28135, n_28136, n_28137, n_28138, n_28141, n_28151, n_28152,n_28153;
wire n_28154, n_28156, n_28157, n_28158, n_28159, n_28160, n_28161,n_28162;
wire n_28163, n_28164, n_28165, n_28166, n_28167, n_28168, n_28169,n_28170;
wire n_28171, n_28172, n_28173, n_28174, n_28175, n_28176, n_28177,n_28178;
wire n_28179, n_28180, n_28181, n_28182, n_28183, n_28184, n_28185,n_28186;
wire n_28187, n_28188, n_28189, n_28192, n_28193, n_28194, n_28195,n_28196;
wire n_28197, n_28199, n_28200, n_28202, n_28203, n_28204, n_28205,n_28206;
wire n_28207, n_28209, n_28210, n_28211, n_28212, n_28213, n_28214,n_28217;
wire n_28218, n_28219, n_28220, n_28221, n_28222, n_28223, n_28224,n_28225;
wire n_28226, n_28239, n_28240, n_28242, n_28243, n_28245, n_28246,n_28247;
wire n_28248, n_28249, n_28250, n_28251, n_28252, n_28253, n_28254,n_28255;
wire n_28256, n_28257, n_28258, n_28259, n_28260, n_28261, n_28262,n_28263;
wire n_28264, n_28265, n_28266, n_28267, n_28268, n_28269, n_28270,n_28271;
wire n_28273, n_28274, n_28275, n_28276, n_28277, n_28278, n_28279,n_28280;
wire n_28283, n_28284, n_28285, n_28286, n_28287, n_28288, n_28310,n_28311;
wire n_28312, n_28313, n_28314, n_28315, n_28316, n_28317, n_28318,n_28319;
wire n_28320, n_28321, n_28322, n_28323, n_28324, n_28325, n_28326,n_28327;
wire n_28328, n_28329, n_28331, n_28332, n_28333, n_28336, n_28340,n_28341;
wire n_28344, n_28345, n_28346, n_28349, n_28350, n_28351, n_28357,n_28358;
wire n_28362, n_28364, n_28365, n_28373, n_28375, n_28380, n_28381,n_28398;
wire n_28402, n_28404, n_28407, n_28408, n_28410, n_28418, n_28419,n_28423;
wire n_28427, n_28433, n_28441, n_28444, n_28445, n_28447, n_28450,n_28452;
wire n_28459, n_28463, n_28464, n_28466, n_28469, n_28470, n_28472,n_28476;
wire n_28478, n_28480, n_28481, n_28482, n_28483, n_28484, n_28485,n_28487;
wire n_28488, n_28501, n_28502, n_28505, n_28506, n_28507, n_28508,n_28509;
wire n_28511, n_28540, n_28542, n_28547, n_28548, n_28549, n_28552,n_28553;
wire n_28556, n_28557, n_28558, n_28559, n_28560, n_28561, n_28562,n_28563;
wire n_28564, n_28566, n_28567, n_28568, n_28574, n_28575, n_28576,n_28577;
wire n_28578, n_28580, n_28581, n_28582, n_28583, n_28584, n_28585,n_28586;
wire n_28588, n_28589, n_28590, n_28591, n_28592, n_28593, n_28594,n_28595;
wire n_28596, n_28597, n_28598, n_28599, n_28601, n_28602, n_28603,n_28604;
wire n_28605, n_28606, n_28607, n_28609, n_28610, n_28611, n_28614,n_28615;
wire n_28616, n_28618, n_28619, n_28620, n_28631, n_28632, n_28642,n_28645;
wire n_28680, n_28686, n_28689, n_28692, n_28724, n_28725, n_28727,n_28728;
wire n_28733, n_28734, n_28742, n_28744, n_28749, n_28754, n_28757,n_28771;
wire n_28775, n_28776, n_28779, n_28780, n_28781, n_28785, n_28786,n_28787;
wire n_28792, n_28793, n_28796, n_28797, n_28798, n_28799, n_28800,n_28802;
wire n_28803, n_28804, n_28807, n_28809, n_28810, n_28812, n_28815,n_28816;
wire n_28820, n_28821, n_28822, n_28825, n_28826, n_28827, n_28829,n_28832;
wire n_28834, n_28836, n_28837, n_28838, n_28840, n_28841, n_28842,n_28843;
wire n_28845, n_28846, n_28847, n_28848, n_28849, n_28850, n_28851,n_28852;
wire n_28853, n_28854, n_28857, n_28858, n_28859, n_28860, n_28862,n_28865;
wire n_28866, n_28869, n_28870, n_28871, n_28872, n_28875, n_28877,n_28878;
wire n_28879, n_28880, n_28881, n_28882, n_28883, n_28884, n_28885,n_28886;
wire n_28887, n_28888, n_28889, n_28890, n_28892, n_28893, n_28894,n_28895;
wire n_28896, n_28897, n_28898, n_28899, n_28900, n_28901, n_28902,n_28903;
wire n_28904, n_28905, n_28907, n_28933, n_28986, n_28988, n_28991,n_28993;
wire n_28996, n_28998, n_29000, n_29002, n_29003, n_29005, n_29007,n_29014;
wire n_29018, n_29039, n_29048, n_29062, n_29065, n_29070, n_29074,n_29085;
wire n_29102, n_29106, n_29114, n_29115, n_29116, n_29119, n_29120,n_29121;
wire n_29122, n_29123, n_29124, n_29125, n_29126, n_29129, n_29130,n_29131;
wire n_29133, n_29134, n_29135, n_29136, n_29137, n_29139, n_29140,n_29142;
wire n_29143, n_29144, n_29145, n_29146, n_29147, n_29149, n_29150,n_29153;
wire n_29155, n_29158, n_29163, n_29166, n_29167, n_29171, n_29173,n_29176;
wire n_29177, n_29178, n_29179, n_29180, n_29181, n_29182, n_29185,n_29186;
wire n_29187, n_29188, n_29189, n_29190, n_29191, n_29192, n_29193,n_29195;
wire n_29196, n_29197, n_29198, n_29199, n_29200, n_29201, n_29202,n_29203;
wire n_29204, n_29205, n_29208, n_29210, n_29214, n_29215, n_29216,n_29217;
wire n_29221, n_29225, n_29228, n_29235, n_29244, n_29256, n_29262,n_29266;
wire n_29269, n_29275, n_29279, n_29286, n_29292, n_29297, n_29298,n_29300;
wire n_29301, n_29302, n_29303, n_29304, n_29305, n_29306, n_29307,n_29308;
wire n_29309, n_29310, n_29311, n_29312, n_29313, n_29314, n_29315,n_29316;
wire n_29317, n_29318, n_29319, n_29320, n_29321, n_29322, n_29323,n_29324;
wire n_29325, n_29326, n_29327, n_29329, n_29330, n_29331, n_29333,n_29336;
wire n_29337, n_29343, n_29347, n_29349, n_29350, n_29351, n_29353,n_29355;
wire n_29357, n_29358, n_29360, n_29363, n_29365, n_29366, n_29367,n_29368;
wire n_29369, n_29370, n_29371, n_29372, n_29373, n_29374, n_29375,n_29376;
wire n_29377, n_29378, n_29379, n_29380, n_29381, n_29382, n_29383,n_29384;
wire n_29385, n_29386, n_29387, n_29388, n_29389, n_29390, n_29391,n_29392;
wire n_29393, n_29395, n_29396, n_29397, n_29399, n_29400, n_29401,n_29402;
wire n_29403, n_29404, n_29405, n_29406, n_29407, n_29408, n_29409,n_29410;
wire n_29411, n_29412, n_29413, n_29414, n_29415, n_29416, n_29417,n_29418;
wire n_29419, n_29420, n_29421, n_29422, n_29423, n_29424, n_29425,n_29426;
wire n_29427, n_29428, n_29429, n_29430, n_29431, n_29432, n_29433,sa00[0] ;
wire sa00[1] , sa00[2] , sa00[3] , sa00[4] , sa00[5] , sa00[6], sa00[7] , sa01[0] ;
wire sa01[1] , sa01[2] , sa01[3] , sa01[4] , sa01[5] , sa01[6], sa01[7] , sa02[0] ;
wire sa02[4] , sa02[5] , sa02[6] , sa02[7] , sa03[0] , sa03[2], sa03[3] , sa03[4] ;
wire sa03[5] , sa03[6] , sa03[7] , sa10[0] , sa10[1] , sa10[2], sa10[3] , sa10[4] ;
wire sa10[5] , sa10[6] , sa10[7] , sa11[0] , sa11[1] , sa11[2], sa11[3] , sa11[4] ;
wire sa11[5] , sa11[6] , sa11[7] , sa12[0] , sa12[1] , sa12[2], sa12[3] , sa12[4] ;
wire sa12[5] , sa12[6] , sa12[7] , sa13[0] , sa13[1] , sa13[2], sa13[3] , sa13[4] ;
wire sa13[5] , sa13[6] , sa13[7] , sa20[0] , sa20[1] , sa20[2], sa20[3] , sa20[4] ;
wire sa20[5] , sa20[6] , sa20[7] , sa21[0] , sa21[1] , sa21[2], sa21[3] , sa21[4] ;
wire sa21[5] , sa21[6] , sa21[7] , sa22[0] , sa22[1] , sa22[2], sa22[3] , sa22[4] ;
wire sa22[5] , sa22[6] , sa22[7] , sa23[0] , sa23[1] , sa23[2], sa23[3] , sa23[4] ;
wire sa23[5] , sa23[6] , sa23[7] , sa30[0] , sa30[1] , sa30[2], sa30[3] , sa30[4] ;
wire sa30[5] , sa30[6] , sa30[7] , sa31[0] , sa31[1] , sa31[2], sa31[3] , sa31[4] ;
wire sa31[5] , sa31[6] , sa31[7] , sa32[0] , sa32[1] , sa32[2], sa32[3] , sa32[4] ;
wire sa32[5] , sa32[6] , sa32[7] , sa33[0] , sa33[1] , sa33[2], sa33[3] , sa33[4] ;
wire sa33[5] , sa33[6] , sa33[7] , text_in_r[0] , text_in_r[1] ,text_in_r[2] , text_in_r[3] , text_in_r[4] ;
wire text_in_r[5] , text_in_r[6] , text_in_r[7] , text_in_r[8] ,text_in_r[9] , text_in_r[10] , text_in_r[11] , text_in_r[12];
wire text_in_r[13] , text_in_r[14] , text_in_r[15] ,text_in_r[16] , text_in_r[17] , text_in_r[18] ,text_in_r[19] , text_in_r[20] ;
wire text_in_r[21] , text_in_r[22] , text_in_r[23] ,text_in_r[24] , text_in_r[25] , text_in_r[26] ,text_in_r[27] , text_in_r[28] ;
wire text_in_r[29] , text_in_r[30] , text_in_r[31] ,text_in_r[32] , text_in_r[33] , text_in_r[34] ,text_in_r[35] , text_in_r[36] ;
wire text_in_r[37] , text_in_r[38] , text_in_r[39] ,text_in_r[40] , text_in_r[41] , text_in_r[42] ,text_in_r[43] , text_in_r[44] ;
wire text_in_r[45] , text_in_r[46] , text_in_r[47] ,text_in_r[48] , text_in_r[49] , text_in_r[50] ,text_in_r[51] , text_in_r[52] ;
wire text_in_r[53] , text_in_r[54] , text_in_r[55] ,text_in_r[56] , text_in_r[57] , text_in_r[58] ,text_in_r[59] , text_in_r[60] ;
wire text_in_r[61] , text_in_r[62] , text_in_r[63] ,text_in_r[64] , text_in_r[65] , text_in_r[66] ,text_in_r[67] , text_in_r[68] ;
wire text_in_r[69] , text_in_r[70] , text_in_r[71] ,text_in_r[72] , text_in_r[73] , text_in_r[74] ,text_in_r[75] , text_in_r[76] ;
wire text_in_r[77] , text_in_r[78] , text_in_r[79] ,text_in_r[80] , text_in_r[81] , text_in_r[82] ,text_in_r[83] , text_in_r[84] ;
wire text_in_r[85] , text_in_r[86] , text_in_r[87] ,text_in_r[88] , text_in_r[89] , text_in_r[90] ,text_in_r[91] , text_in_r[92] ;
wire text_in_r[93] , text_in_r[94] , text_in_r[95] ,text_in_r[96] , text_in_r[97] , text_in_r[98] ,text_in_r[99] , text_in_r[100] ;
wire text_in_r[101] , text_in_r[102] , text_in_r[103] ,text_in_r[104] , text_in_r[105] , text_in_r[106] ,text_in_r[107] , text_in_r[108] ;
wire text_in_r[109] , text_in_r[110] , text_in_r[111] ,text_in_r[112] , text_in_r[113] , text_in_r[114] ,text_in_r[115] , text_in_r[116] ;
wire text_in_r[117] , text_in_r[118] , text_in_r[119] ,text_in_r[120] , text_in_r[121] , text_in_r[122] ,text_in_r[123] , text_in_r[124] ;
wire text_in_r[125] , text_in_r[126] , text_in_r[127] ,u0_r0_rcnt[0] , u0_r0_rcnt[1] , u0_r0_rcnt[2] ,u0_r0_rcnt[3] , u0_rcon_1053;
wire u0_rcon_1054, u0_rcon_1055, u0_rcon_1056, u0_rcon_1057,u0_rcon_1058, u0_rcon_1059, u0_rcon_1060, w0[0] ;
wire w0[1] , w0[2] , w0[3] , w0[4] , w0[6] , w0[7] , w0[8] ,w0[9] ;
wire w0[10] , w0[13] , w0[14] , w0[17] , w0[18] , w0[22] ,w0[25] , w0[26] ;
wire w0[28] , w0[30] , w0[31] , w1[0] , w1[1] , w1[3] , w1[4], w1[5] ;
wire w1[9] , w1[10] , w1[12] , w1[14] , w1[15] , w1[16] ,w1[17] , w1[18] ;
wire w1[20] , w1[23] , w1[24] , w1[25] , w1[27] , w1[31] ,w2[0] , w2[1] ;
wire w2[2] , w2[3] , w2[4] , w2[5] , w2[6] , w2[7] , w2[8] ,w2[9] ;
wire w2[10] , w2[11] , w2[12] , w2[13] , w2[14] , w2[15] ,w2[16] , w2[17] ;
wire w2[18] , w2[19] , w2[20] , w2[21] , w2[22] , w2[23] ,w2[24] , w2[25] ;
wire w2[26] , w2[27] , w2[28] , w2[30] , w2[31] , w3[0] ,w3[1] , w3[2] ;
wire w3[3] , w3[4] , w3[5] , w3[6] , w3[7] , w3[8] , w3[9] ,w3[10] ;
wire w3[11] , w3[12] , w3[13] , w3[14] , w3[15] , w3[16] ,w3[17] , w3[19] ;
wire w3[20] , w3[21] , w3[22] , w3[23] , w3[25] , w3[26] ,w3[28] , w3[29] ;
wire w3[30] , w3[31] ;
DFFX1 sa22_reg[4] (.CK (clk), .D (n_25439), .Q (sa22[4] ), .QN ());
DFFX1 sa02_reg[1] (.CK (clk), .D (n_25437), .Q (n_2204), .QN ());
DFFX1 sa01_reg[1] (.CK (clk), .D (n_25438), .Q (sa01[1] ), .QN ());
DFFX1 sa00_reg[1] (.CK (clk), .D (n_25436), .Q (sa00[1] ), .QN ());
DFFX1 sa03_reg[4] (.CK (clk), .D (n_25435), .Q (sa03[4] ), .QN ());
DFFX1 sa03_reg[3] (.CK (clk), .D (n_25423), .Q (sa03[3] ), .QN ());
DFFX1 sa33_reg[0] (.CK (clk), .D (n_25434), .Q (sa33[0] ), .QN ());
DFFX1 sa02_reg[4] (.CK (clk), .D (n_25433), .Q (sa02[4] ), .QN ());
DFFX1 sa12_reg[3] (.CK (clk), .D (n_25429), .Q (sa12[3] ), .QN ());
DFFX1 sa32_reg[3] (.CK (clk), .D (n_25427), .Q (sa32[3] ), .QN ());
SDFFSRX1 sa32_reg[0] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25378), .SE (n_25440), .SI (n_894), .Q (), .QN (sa32[0] ));
DFFX1 sa22_reg[3] (.CK (clk), .D (n_25430), .Q (sa22[3] ), .QN ());
SDFFSRX1 sa31_reg[0] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25350), .SE (n_25440), .SI (n_3393), .Q (sa31[0] ), .QN ());
DFFX1 sa02_reg[3] (.CK (clk), .D (n_25431), .Q (n_28933), .QN ());
DFFX1 sa20_reg[3] (.CK (clk), .D (n_25425), .Q (sa20[3] ), .QN ());
SDFFSRX1 sa30_reg[0] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25374), .SE (n_25440), .SI (n_884), .Q (sa30[0] ), .QN ());
DFFX1 sa00_reg[4] (.CK (clk), .D (n_25424), .Q (sa00[4] ), .QN ());
DFFX1 sa10_reg[0] (.CK (clk), .D (n_25421), .Q (sa10[0] ), .QN ());
DFFX1 sa03_reg[0] (.CK (clk), .D (n_25404), .Q (sa03[0] ), .QN ());
DFFX1 sa33_reg[3] (.CK (clk), .D (n_25406), .Q (sa33[3] ), .QN ());
DFFX1 sa13_reg[0] (.CK (clk), .D (n_25400), .Q (sa13[0] ), .QN ());
DFFSRX1 sa02_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25925), .Q (sa02[6] ), .QN ());
DFFX1 sa22_reg[5] (.CK (clk), .D (n_25414), .Q (sa22[5] ), .QN ());
DFFX1 sa13_reg[4] (.CK (clk), .D (n_25412), .Q (sa13[4] ), .QN ());
DFFX1 sa03_reg[1] (.CK (clk), .D (n_25390), .Q (n_908), .QN ());
DFFX1 sa32_reg[5] (.CK (clk), .D (n_25401), .Q (sa32[5] ), .QN ());
DFFX1 sa12_reg[1] (.CK (clk), .D (n_25399), .Q (sa12[1] ), .QN ());
DFFX1 sa13_reg[3] (.CK (clk), .D (n_25384), .Q (sa13[3] ), .QN ());
DFFX1 sa23_reg[3] (.CK (clk), .D (n_25419), .Q (sa23[3] ), .QN ());
DFFX1 sa02_reg[0] (.CK (clk), .D (n_25396), .Q (sa02[0] ), .QN ());
DFFX1 sa12_reg[0] (.CK (clk), .D (n_25394), .Q (sa12[0] ), .QN ());
DFFX1 sa21_reg[4] (.CK (clk), .D (n_25408), .Q (sa21[4] ), .QN ());
DFFX1 sa01_reg[4] (.CK (clk), .D (n_25411), .Q (sa01[4] ), .QN ());
DFFX1 sa31_reg[5] (.CK (clk), .D (n_25410), .Q (sa31[5] ), .QN ());
DFFX1 sa11_reg[1] (.CK (clk), .D (n_25405), .Q (sa11[1] ), .QN ());
DFFX1 sa21_reg[3] (.CK (clk), .D (n_25402), .Q (sa21[3] ), .QN ());
DFFX1 sa01_reg[0] (.CK (clk), .D (n_25397), .Q (sa01[0] ), .QN ());
DFFX1 sa21_reg[5] (.CK (clk), .D (n_25416), .Q (sa21[5] ), .QN ());
DFFX1 sa11_reg[0] (.CK (clk), .D (n_25398), .Q (sa11[0] ), .QN ());
DFFX1 sa10_reg[1] (.CK (clk), .D (n_25388), .Q (sa10[1] ), .QN ());
DFFX1 sa20_reg[1] (.CK (clk), .D (n_25387), .Q (sa20[1] ), .QN ());
DFFX1 sa00_reg[5] (.CK (clk), .D (n_25392), .Q (sa00[5] ), .QN ());
DFFSRX1 sa30_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25389), .Q (sa30[6] ), .QN ());
DFFX1 sa10_reg[3] (.CK (clk), .D (n_25385), .Q (sa10[3] ), .QN ());
DFFX1 sa00_reg[0] (.CK (clk), .D (n_25383), .Q (sa00[0] ), .QN ());
DFFSRX1 sa00_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25420), .Q (sa00[7] ), .QN ());
OAI21X1 g56961(.A0 (n_25349), .A1 (n_25432), .B0 (n_8395), .Y(n_25439));
OAI21X1 g57319(.A0 (n_25352), .A1 (n_25407), .B0 (n_8536), .Y(n_25438));
OAI21X1 g56974(.A0 (n_25348), .A1 (n_25426), .B0 (n_8665), .Y(n_25437));
OAI21X1 g57684(.A0 (n_25375), .A1 (n_25361), .B0 (n_8580), .Y(n_25436));
DFFSRX1 sa23_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25357), .Q (sa23[6] ), .QN ());
OAI21X1 g56632(.A0 (n_25296), .A1 (n_25415), .B0 (n_15789), .Y(n_25435));
DFFSRX1 sa13_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25365), .Q (sa13[6] ), .QN ());
DFFX1 sa13_reg[1] (.CK (clk), .D (n_25336), .Q (sa13[1] ), .QN ());
DFFX1 sa33_reg[4] (.CK (clk), .D (n_25345), .Q (sa33[4] ), .QN ());
DFFSRX1 sa23_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25346), .Q (sa23[7] ), .QN ());
DFFSRX1 sa33_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25347), .Q (sa33[7] ), .QN ());
DFFSRX1 sa03_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25379), .Q (sa03[6] ), .QN ());
OAI21X1 g56704(.A0 (n_25299), .A1 (ld_r), .B0 (n_8629), .Y (n_25434));
DFFX1 sa23_reg[0] (.CK (clk), .D (n_25354), .Q (sa23[0] ), .QN ());
DFFX1 sa02_reg[5] (.CK (clk), .D (n_25372), .Q (sa02[5] ), .QN ());
DFFSRX1 sa32_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25373), .Q (sa32[6] ), .QN ());
DFFSRX1 sa12_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25367), .Q (sa12[6] ), .QN ());
DFFSRX1 sa22_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25364), .Q (sa22[6] ), .QN ());
DFFX1 sa22_reg[1] (.CK (clk), .D (n_25360), .Q (sa22[1] ), .QN ());
DFFX1 sa12_reg[4] (.CK (clk), .D (n_25358), .Q (sa12[4] ), .QN ());
DFFX1 sa22_reg[0] (.CK (clk), .D (n_25351), .Q (sa22[0] ), .QN ());
DFFSRX1 sa01_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25369), .Q (sa01[6] ), .QN ());
DFFSRX1 sa11_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25368), .Q (sa11[6] ), .QN ());
DFFSRX1 sa31_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25366), .Q (sa31[6] ), .QN ());
DFFX1 sa01_reg[5] (.CK (clk), .D (n_25371), .Q (sa01[5] ), .QN ());
DFFX1 sa21_reg[1] (.CK (clk), .D (n_27892), .Q (sa21[1] ), .QN ());
DFFX1 sa11_reg[3] (.CK (clk), .D (n_25359), .Q (sa11[3] ), .QN ());
DFFX1 sa01_reg[3] (.CK (clk), .D (n_25362), .Q (sa01[3] ), .QN ());
DFFX1 sa21_reg[0] (.CK (clk), .D (n_25356), .Q (sa21[0] ), .QN ());
DFFX1 sa31_reg[3] (.CK (clk), .D (n_25355), .Q (sa31[3] ), .QN ());
DFFX1 sa10_reg[5] (.CK (clk), .D (n_25344), .Q (sa10[5] ), .QN ());
DFFX1 sa30_reg[5] (.CK (clk), .D (n_25342), .Q (sa30[5] ), .QN ());
DFFX1 sa20_reg[5] (.CK (clk), .D (n_25343), .Q (sa20[5] ), .QN ());
DFFX1 sa30_reg[1] (.CK (clk), .D (n_25340), .Q (sa30[1] ), .QN ());
DFFX1 sa00_reg[3] (.CK (clk), .D (n_25339), .Q (sa00[3] ), .QN ());
DFFX1 sa30_reg[4] (.CK (clk), .D (n_25338), .Q (sa30[4] ), .QN ());
DFFX1 sa10_reg[4] (.CK (clk), .D (n_25337), .Q (sa10[4] ), .QN ());
DFFSRX1 sa10_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25334), .Q (sa10[6] ), .QN ());
DFFX1 sa20_reg[0] (.CK (clk), .D (n_25333), .Q (sa20[0] ), .QN ());
DFFX1 sa30_reg[3] (.CK (clk), .D (n_25331), .Q (sa30[3] ), .QN ());
DFFX1 sa30_reg[2] (.CK (clk), .D (n_25380), .Q (sa30[2] ), .QN ());
DFFSRX1 sa00_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25381), .Q (sa00[6] ), .QN ());
DFFSRX1 sa20_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25377), .Q (sa20[6] ), .QN ());
DFFX1 sa20_reg[2] (.CK (clk), .D (n_25376), .Q (sa20[2] ), .QN ());
OAI21X1 g56959(.A0 (n_25292), .A1 (n_25432), .B0 (n_8711), .Y(n_25433));
OAI21X1 g56978(.A0 (n_25291), .A1 (n_25428), .B0 (n_8256), .Y(n_25431));
OAI21X1 g56980(.A0 (n_25289), .A1 (n_25395), .B0 (n_9794), .Y(n_25430));
OAI21X1 g56979(.A0 (n_25290), .A1 (n_25428), .B0 (n_8260), .Y(n_25429));
OAI21X1 g57010(.A0 (n_25288), .A1 (n_25426), .B0 (n_10235), .Y(n_25427));
OAI21X1 g57681(.A0 (n_25325), .A1 (n_25418), .B0 (n_8749), .Y(n_25425));
OAI21X1 g57685(.A0 (n_25324), .A1 (n_25422), .B0 (n_10041), .Y(n_25424));
OAI21X1 g56649(.A0 (n_25293), .A1 (n_25422), .B0 (n_19688), .Y(n_25423));
OAI21X1 g57687(.A0 (n_25323), .A1 (n_25382), .B0 (n_8345), .Y(n_25421));
NAND2X1 g57703(.A (n_25615), .B (n_25616), .Y (n_25420));
OAI21X1 g56652(.A0 (n_25231), .A1 (n_25418), .B0 (n_18515), .Y(n_25419));
DFFX1 sa03_reg[5] (.CK (clk), .D (n_25286), .Q (sa03[5] ), .QN ());
DFFX1 sa23_reg[4] (.CK (clk), .D (n_25306), .Q (sa23[4] ), .QN ());
DFFX1 sa33_reg[5] (.CK (clk), .D (n_25319), .Q (sa33[5] ), .QN ());
DFFX1 sa23_reg[5] (.CK (clk), .D (n_25315), .Q (sa23[5] ), .QN ());
DFFX1 sa33_reg[1] (.CK (clk), .D (n_25310), .Q (sa33[1] ), .QN ());
DFFX1 sa23_reg[1] (.CK (clk), .D (n_25321), .Q (sa23[1] ), .QN ());
DFFX1 sa33_reg[2] (.CK (clk), .D (n_25297), .Q (sa33[2] ), .QN ());
DFFX1 sa03_reg[2] (.CK (clk), .D (n_25314), .Q (sa03[2] ), .QN ());
DFFX1 sa23_reg[2] (.CK (clk), .D (n_25300), .Q (sa23[2] ), .QN ());
DFFSRX1 sa13_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25304), .Q (sa13[7] ), .QN ());
DFFSRX1 sa03_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25307), .Q (sa03[7] ), .QN ());
DFFX1 sa12_reg[5] (.CK (clk), .D (n_25316), .Q (sa12[5] ), .QN ());
DFFX1 sa32_reg[1] (.CK (clk), .D (n_25308), .Q (sa32[1] ), .QN ());
DFFSRX1 sa22_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25301), .Q (sa22[7] ), .QN ());
DFFSRX1 sa02_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25298), .Q (sa02[7] ), .QN ());
DFFSRX1 sa12_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25295), .Q (sa12[7] ), .QN ());
DFFSRX1 sa21_reg[6] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25317), .Q (sa21[6] ), .QN ());
DFFX1 sa11_reg[5] (.CK (clk), .D (n_25318), .Q (sa11[5] ), .QN ());
DFFX1 sa31_reg[1] (.CK (clk), .D (n_25313), .Q (sa31[1] ), .QN ());
DFFX1 sa11_reg[4] (.CK (clk), .D (n_25311), .Q (sa11[4] ), .QN ());
DFFX1 sa31_reg[2] (.CK (clk), .D (n_25309), .Q (sa31[2] ), .QN ());
DFFSRX1 sa01_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25303), .Q (sa01[7] ), .QN ());
DFFX1 sa21_reg[2] (.CK (clk), .D (n_25302), .Q (sa21[2] ), .QN ());
DFFX1 sa20_reg[4] (.CK (clk), .D (n_25285), .Q (sa20[4] ), .QN ());
DFFSRX1 sa20_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25328), .Q (sa20[7] ), .QN ());
DFFSRX1 sa10_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25330), .Q (sa10[7] ), .QN ());
DFFX1 sa30_reg[7] (.CK (clk), .D (n_25327), .Q (sa30[7] ), .QN ());
OAI21X1 g57266(.A0 (n_25254), .A1 (n_25415), .B0 (n_8159), .Y(n_25416));
OAI21X1 g56925(.A0 (n_25245), .A1 (ld_r), .B0 (n_8144), .Y (n_25414));
OAI21X1 g56633(.A0 (n_25240), .A1 (n_25386), .B0 (n_15720), .Y(n_25412));
OAI21X1 g57301(.A0 (n_25247), .A1 (n_25409), .B0 (n_8194), .Y(n_25411));
OAI21X1 g57303(.A0 (n_25248), .A1 (n_25409), .B0 (n_8123), .Y(n_25410));
OAI21X1 g57304(.A0 (n_25249), .A1 (n_25407), .B0 (n_8265), .Y(n_25408));
OAI21X1 g56667(.A0 (n_25263), .A1 (n_25403), .B0 (n_19720), .Y(n_25406));
OAI21X1 g57316(.A0 (n_25246), .A1 (n_25440), .B0 (n_8358), .Y(n_25405));
OAI21X1 g56668(.A0 (n_25267), .A1 (n_25403), .B0 (n_8199), .Y(n_25404));
OAI21X1 g57323(.A0 (n_25244), .A1 (n_25403), .B0 (n_10201), .Y(n_25402));
OAI21X1 g56958(.A0 (n_25237), .A1 (n_25432), .B0 (n_8484), .Y(n_25401));
OAI21X1 g56670(.A0 (n_25264), .A1 (n_25332), .B0 (n_8193), .Y(n_25400));
OAI21X1 g56972(.A0 (n_25236), .A1 (n_25428), .B0 (n_9197), .Y(n_25399));
OAI21X1 g57354(.A0 (n_25243), .A1 (n_25393), .B0 (n_8212), .Y(n_25398));
OAI21X1 g57357(.A0 (n_25242), .A1 (n_25391), .B0 (n_8429), .Y(n_25397));
OAI21X1 g57012(.A0 (n_25232), .A1 (n_25395), .B0 (n_8673), .Y(n_25396));
OAI21X1 g57013(.A0 (n_25233), .A1 (n_25393), .B0 (n_8202), .Y(n_25394));
OAI21X1 g57654(.A0 (n_25278), .A1 (n_25391), .B0 (n_8521), .Y(n_25392));
OAI21X1 g56646(.A0 (n_25235), .A1 (n_25422), .B0 (n_17389), .Y(n_25390));
NAND2X1 g57658(.A (n_25759), .B (n_25760), .Y (n_25389));
OAI21X1 g57676(.A0 (n_25272), .A1 (n_25341), .B0 (n_8229), .Y(n_25388));
OAI21X1 g57677(.A0 (n_25271), .A1 (n_25386), .B0 (n_8361), .Y(n_25387));
OAI21X1 g57680(.A0 (n_25268), .A1 (n_25418), .B0 (n_8628), .Y(n_25385));
OAI21X1 g56650(.A0 (n_25234), .A1 (n_25422), .B0 (n_20234), .Y(n_25384));
OAI21X1 g57686(.A0 (n_25265), .A1 (n_25382), .B0 (n_8299), .Y(n_25383));
NAND2X1 g57702(.A (n_8570), .B (n_25275), .Y (n_25381));
OAI21X1 g57701(.A0 (n_25217), .A1 (n_25335), .B0 (n_10090), .Y(n_25380));
NAND2X2 g56613(.A (n_13769), .B (n_25276), .Y (n_25379));
INVX1 g57122(.A (n_25329), .Y (n_25378));
NAND2X2 g57706(.A (n_7853), .B (n_25273), .Y (n_25377));
DFFX1 sa13_reg[5] (.CK (clk), .D (n_25262), .Q (sa13[5] ), .QN ());
DFFX1 sa33_reg[6] (.CK (clk), .D (n_25230), .Q (sa33[6] ), .QN ());
DFFX1 sa32_reg[2] (.CK (clk), .D (n_25252), .Q (sa32[2] ), .QN ());
DFFX1 sa02_reg[2] (.CK (clk), .D (n_25241), .Q (n_688), .QN ());
DFFX1 sa12_reg[2] (.CK (clk), .D (n_25239), .Q (sa12[2] ), .QN ());
DFFX1 sa22_reg[2] (.CK (clk), .D (n_25238), .Q (sa22[2] ), .QN ());
DFFX1 sa01_reg[2] (.CK (clk), .D (n_25253), .Q (sa01[2] ), .QN ());
DFFX1 sa11_reg[2] (.CK (clk), .D (n_25251), .Q (sa11[2] ), .QN ());
DFFSRX1 sa11_reg[7] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_25250), .Q (sa11[7] ), .QN ());
DFFX1 sa00_reg[2] (.CK (clk), .D (n_25282), .Q (sa00[2] ), .QN ());
DFFX1 u0_w_reg[2][19] (.CK (clk), .D (n_25277), .Q (w2[19] ), .QN());
DFFX1 sa10_reg[2] (.CK (clk), .D (n_25281), .Q (sa10[2] ), .QN ());
OAI21X1 g57767(.A0 (n_25211), .A1 (n_25353), .B0 (n_8183), .Y(n_25376));
MX2X1 g57780(.A (n_24728), .B (n_24727), .S0 (n_25205), .Y (n_25375));
INVX1 g57786(.A (n_25322), .Y (n_25374));
NAND2X2 g56919(.A (n_28317), .B (n_28318), .Y (n_25373));
OAI21X1 g56921(.A0 (n_25197), .A1 (n_25370), .B0 (n_8507), .Y(n_25372));
OAI21X1 g57262(.A0 (n_25203), .A1 (n_25370), .B0 (n_9545), .Y(n_25371));
NAND2X2 g57263(.A (n_25610), .B (n_25611), .Y (n_25369));
NAND2X1 g57264(.A (n_25772), .B (n_25773), .Y (n_25368));
NAND2X1 g56923(.A (n_8748), .B (n_25256), .Y (n_25367));
NAND2X2 g57268(.A (n_25600), .B (n_25601), .Y (n_25366));
NAND2X2 g56615(.A (n_29378), .B (n_29379), .Y (n_25365));
NAND2X1 g56926(.A (n_9742), .B (n_25255), .Y (n_25364));
OAI21X1 g57321(.A0 (n_25198), .A1 (n_25361), .B0 (n_8448), .Y(n_25362));
OAI21X1 g56957(.A0 (n_25191), .A1 (ld_r), .B0 (n_8149), .Y (n_25360));
OAI21X1 g57322(.A0 (n_25196), .A1 (n_25403), .B0 (n_9152), .Y(n_25359));
OAI21X1 g56960(.A0 (n_25188), .A1 (n_25432), .B0 (n_10974), .Y(n_25358));
NAND2X2 g56617(.A (n_25668), .B (n_25669), .Y (n_25357));
OAI21X1 g57358(.A0 (n_25192), .A1 (n_25386), .B0 (n_10093), .Y(n_25356));
OAI21X1 g57360(.A0 (n_25193), .A1 (n_25320), .B0 (n_10057), .Y(n_25355));
OAI21X1 g56675(.A0 (n_25215), .A1 (n_25353), .B0 (n_9289), .Y(n_25354));
MX2X1 g57382(.A (n_24678), .B (n_24677), .S0 (n_25206), .Y (n_25352));
OAI21X1 g57016(.A0 (n_25183), .A1 (n_25393), .B0 (n_8386), .Y(n_25351));
INVX1 g57466(.A (n_25294), .Y (n_25350));
MX2X1 g57018(.A (n_25209), .B (n_25210), .S0 (n_24633), .Y (n_25349));
MX2X1 g57039(.A (n_24621), .B (n_24620), .S0 (n_25207), .Y (n_25348));
NAND2X2 g56611(.A (n_25659), .B (n_25660), .Y (n_25347));
NAND2X2 g56647(.A (n_25675), .B (n_25676), .Y (n_25346));
OAI21X1 g56648(.A0 (n_25185), .A1 (n_25382), .B0 (n_15710), .Y(n_25345));
OAI21X1 g57655(.A0 (n_25228), .A1 (n_25391), .B0 (n_8608), .Y(n_25344));
OAI21X1 g57656(.A0 (n_25227), .A1 (n_25415), .B0 (n_8522), .Y(n_25343));
OAI21X1 g57657(.A0 (n_25229), .A1 (n_25341), .B0 (n_8734), .Y(n_25342));
OAI21X1 g57678(.A0 (n_25223), .A1 (n_25341), .B0 (n_8537), .Y(n_25340));
OAI21X1 g57679(.A0 (n_25222), .A1 (n_25305), .B0 (n_8721), .Y(n_25339));
OAI21X1 g57683(.A0 (n_25221), .A1 (n_25361), .B0 (n_9858), .Y(n_25338));
OAI21X1 g57688(.A0 (n_25220), .A1 (n_25382), .B0 (n_8384), .Y(n_25337));
OAI21X1 g56651(.A0 (n_25184), .A1 (n_25335), .B0 (n_11741), .Y(n_25336));
NAND2X2 g57689(.A (n_28561), .B (n_28562), .Y (n_25334));
OAI21X1 g57690(.A0 (n_25218), .A1 (n_25332), .B0 (n_10017), .Y(n_25333));
OAI21X1 g57691(.A0 (n_25219), .A1 (n_25332), .B0 (n_8135), .Y(n_25331));
NAND2X2 g57705(.A (n_25787), .B (n_25788), .Y (n_25330));
XOR2X1 g57123(.A (n_23523), .B (n_25153), .Y (n_25329));
NAND2X2 g57707(.A (n_25721), .B (n_25722), .Y (n_25328));
OAI21X1 g57708(.A0 (n_25168), .A1 (n_25418), .B0 (n_9549), .Y(n_25327));
NAND2X1 g57760(.A (n_25216), .B (n_25274), .Y (n_25615));
DFFX1 sa13_reg[2] (.CK (clk), .D (n_25202), .Q (sa13[2] ), .QN ());
DFFX1 sa32_reg[7] (.CK (clk), .D (n_25214), .Q (sa32[7] ), .QN ());
DFFX1 sa32_reg[4] (.CK (clk), .D (n_25200), .Q (sa32[4] ), .QN ());
DFFX1 sa31_reg[7] (.CK (clk), .D (n_25213), .Q (sa31[7] ), .QN ());
DFFX1 sa31_reg[4] (.CK (clk), .D (n_25204), .Q (sa31[4] ), .QN ());
DFFX1 sa21_reg[7] (.CK (clk), .D (n_25208), .Q (sa21[7] ), .QN ());
MX2X1 g57774(.A (n_24696), .B (n_24695), .S0 (n_25151), .Y (n_25325));
MX2X1 g57781(.A (n_28112), .B (n_25159), .S0 (n_24729), .Y (n_25324));
MX2X1 g57783(.A (n_24202), .B (n_24201), .S0 (n_25155), .Y (n_25323));
XOR2X1 g57787(.A (n_23487), .B (n_25149), .Y (n_25322));
OAI21X1 g56630(.A0 (n_25144), .A1 (n_25320), .B0 (n_11837), .Y(n_25321));
OAI21X1 g56631(.A0 (n_25133), .A1 (n_25320), .B0 (n_13817), .Y(n_25319));
OAI21X1 g57265(.A0 (n_25154), .A1 (n_25409), .B0 (n_8205), .Y(n_25318));
NAND2X1 g57267(.A (n_25704), .B (n_25705), .Y (n_25317));
OAI21X1 g56924(.A0 (n_25140), .A1 (n_25370), .B0 (n_8283), .Y(n_25316));
OAI21X1 g56616(.A0 (n_25177), .A1 (n_25407), .B0 (n_13847), .Y(n_25315));
OAI21X1 g56666(.A0 (n_25179), .A1 (n_25353), .B0 (n_18445), .Y(n_25314));
OAI21X1 g57300(.A0 (n_25145), .A1 (ld_r), .B0 (n_8126), .Y (n_25313));
OAI21X1 g57302(.A0 (n_25143), .A1 (n_25415), .B0 (n_8808), .Y(n_25311));
OAI21X1 g56634(.A0 (n_25137), .A1 (n_25341), .B0 (n_10227), .Y(n_25310));
OAI21X1 g57317(.A0 (n_25141), .A1 (n_25407), .B0 (n_8483), .Y(n_25309));
OAI21X1 g56956(.A0 (n_25132), .A1 (n_25426), .B0 (n_8777), .Y(n_25308));
NAND2X1 g56669(.A (n_29177), .B (n_29178), .Y (n_25307));
OAI21X1 g56635(.A0 (n_25134), .A1 (n_25305), .B0 (n_18346), .Y(n_25306));
NAND2X2 g56672(.A (n_25564), .B (n_25565), .Y (n_25304));
NAND2X1 g57353(.A (n_25602), .B (n_25603), .Y (n_25303));
OAI21X1 g57359(.A0 (n_25135), .A1 (n_25386), .B0 (n_8508), .Y(n_25302));
NAND2X1 g56976(.A (n_8143), .B (n_25194), .Y (n_25301));
OAI21X1 g56674(.A0 (n_25176), .A1 (n_25353), .B0 (n_19756), .Y(n_25300));
MX2X1 g56761(.A (n_23917), .B (n_23916), .S0 (n_25162), .Y (n_25299));
NAND2X1 g57011(.A (n_8357), .B (n_25187), .Y (n_25298));
OAI21X1 g56645(.A0 (n_25131), .A1 (n_25305), .B0 (n_18544), .Y(n_25297));
MX2X1 g56680(.A (n_25156), .B (n_25157), .S0 (n_24941), .Y (n_25296));
NAND2X2 g57015(.A (n_25730), .B (n_25731), .Y (n_25295));
XOR2X1 g57467(.A (n_23360), .B (n_25146), .Y (n_25294));
MX2X1 g56687(.A (n_24978), .B (n_24979), .S0 (n_25163), .Y (n_25293));
MX2X1 g57021(.A (n_25160), .B (n_25161), .S0 (n_24479), .Y (n_25292));
MX2X1 g57034(.A (n_24835), .B (n_24836), .S0 (n_25130), .Y (n_25291));
MX2X1 g57035(.A (n_24886), .B (n_24887), .S0 (n_25129), .Y (n_25290));
XOR2X1 g57036(.A (n_25150), .B (n_24622), .Y (n_25289));
MX2X1 g57061(.A (n_25181), .B (n_25182), .S0 (n_25009), .Y (n_25288));
NAND2X1 g57675(.A (n_25226), .B (n_25283), .Y (n_25759));
OAI21X1 g56612(.A0 (n_25178), .A1 (n_25409), .B0 (n_11681), .Y(n_25286));
OAI21X1 g57682(.A0 (n_25175), .A1 (n_25305), .B0 (n_9762), .Y(n_25285));
NAND2X1 g57699(.A (n_25283), .B (n_28604), .Y (n_28561));
OAI21X1 g57700(.A0 (n_25115), .A1 (n_25335), .B0 (n_8518), .Y(n_25282));
OAI21X1 g57704(.A0 (n_25107), .A1 (n_25335), .B0 (n_8593), .Y(n_25281));
NAND2X2 g56626(.A (n_25174), .B (n_25922), .Y (n_25659));
MX2X1 g57713(.A (n_25015), .B (n_25014), .S0 (n_25106), .Y (n_25278));
MX2X1 g57715(.A (n_25105), .B (key[51]), .S0 (n_25126), .Y (n_25277));
NAND2X2 g56627(.A (n_25167), .B (n_25283), .Y (n_25276));
DFFX1 u0_w_reg[3][29] (.CK (clk), .D (n_25180), .Q (w3[29] ), .QN());
DFFX1 u0_w_reg[0][19] (.CK (clk), .D (n_25172), .Q (n_24266), .QN());
DFFX1 u0_w_reg[1][19] (.CK (clk), .D (n_25171), .Q (), .QN (n_1385));
DFFX1 u0_w_reg[3][19] (.CK (clk), .D (n_25169), .Q (w3[19] ), .QN());
NAND2X1 g57759(.A (n_25164), .B (n_25274), .Y (n_25275));
NAND2X2 g57762(.A (n_25165), .B (n_25269), .Y (n_25273));
MX2X1 g57764(.A (n_25100), .B (n_25101), .S0 (n_24876), .Y (n_25272));
MX2X1 g57765(.A (n_24522), .B (n_24521), .S0 (n_25095), .Y (n_25271));
NAND2X2 g56628(.A (n_26998), .B (n_25269), .Y (n_29378));
XOR2X1 g57773(.A (n_24735), .B (n_25094), .Y (n_25268));
MX2X1 g56711(.A (n_24668), .B (n_24667), .S0 (n_25089), .Y (n_25267));
NAND2X1 g56629(.A (n_25170), .B (n_25274), .Y (n_25668));
MX2X1 g57782(.A (n_24206), .B (n_24205), .S0 (n_25084), .Y (n_25265));
MX2X1 g56712(.A (n_24660), .B (n_24659), .S0 (n_25088), .Y (n_25264));
MX2X1 g56720(.A (n_24674), .B (n_24675), .S0 (n_25077), .Y (n_25263));
OAI21X1 g56614(.A0 (n_25119), .A1 (ld_r), .B0 (n_13839), .Y(n_25262));
NAND2X2 g56665(.A (n_25128), .B (n_25922), .Y (n_25675));
NAND2X2 g57290(.A (n_25148), .B (n_25283), .Y (n_25610));
NAND2X1 g57291(.A (n_25147), .B (n_25269), .Y (n_25772));
NAND2X1 g57293(.A (n_25152), .B (n_25274), .Y (n_25600));
NAND2X1 g56936(.A (n_25139), .B (n_25922), .Y (n_28317));
NAND2X1 g56949(.A (n_25136), .B (n_25269), .Y (n_25256));
NAND2X1 g56950(.A (n_25138), .B (n_25283), .Y (n_25255));
MX2X1 g57326(.A (n_24694), .B (n_24693), .S0 (n_25109), .Y (n_25254));
OAI21X1 g57350(.A0 (n_25071), .A1 (n_25391), .B0 (n_8451), .Y(n_25253));
OAI21X1 g56973(.A0 (n_25066), .A1 (n_25428), .B0 (n_8526), .Y(n_25252));
OAI21X1 g57355(.A0 (n_25067), .A1 (n_25393), .B0 (n_8747), .Y(n_25251));
NAND2X1 g57356(.A (n_25824), .B (n_25825), .Y (n_25250));
MX2X1 g57361(.A (n_25090), .B (n_25091), .S0 (n_24691), .Y (n_25249));
MX2X1 g57363(.A (n_24832), .B (n_24833), .S0 (n_25111), .Y (n_25248));
MX2X1 g57364(.A (n_25085), .B (n_25086), .S0 (n_24539), .Y (n_25247));
MX2X1 g57374(.A (n_25099), .B (n_25098), .S0 (n_24827), .Y (n_25246));
MX2X1 g56982(.A (n_24642), .B (n_24641), .S0 (n_25108), .Y (n_25245));
XOR2X1 g57378(.A (n_25075), .B (n_24679), .Y (n_25244));
MX2X1 g57401(.A (n_24650), .B (n_24649), .S0 (n_25083), .Y (n_25243));
MX2X1 g57402(.A (n_24652), .B (n_24651), .S0 (n_25080), .Y (n_25242));
OAI21X1 g57008(.A0 (n_25064), .A1 (n_25395), .B0 (n_8678), .Y(n_25241));
MX2X1 g56679(.A (n_25018), .B (n_25017), .S0 (n_25116), .Y (n_25240));
OAI21X1 g57014(.A0 (n_25061), .A1 (n_25395), .B0 (n_8640), .Y(n_25239));
OAI21X1 g57017(.A0 (n_25063), .A1 (n_25370), .B0 (n_8408), .Y(n_25238));
MX2X1 g57019(.A (n_24801), .B (n_24802), .S0 (n_25113), .Y (n_25237));
MX2X1 g57031(.A (n_25097), .B (n_25096), .S0 (n_24794), .Y (n_25236));
MX2X1 g56685(.A (n_24587), .B (n_24586), .S0 (n_25087), .Y (n_25235));
MX2X1 g56689(.A (n_25093), .B (n_25092), .S0 (n_24743), .Y (n_25234));
MX2X1 g57059(.A (n_24789), .B (n_24788), .S0 (n_25082), .Y (n_25233));
MX2X1 g57060(.A (n_24783), .B (n_24782), .S0 (n_25081), .Y (n_25232));
XOR2X1 g56690(.A (n_24581), .B (n_25079), .Y (n_25231));
OAI21X1 g56610(.A0 (n_25118), .A1 (n_25320), .B0 (n_11713), .Y(n_25230));
MX2X1 g57714(.A (n_24725), .B (n_24726), .S0 (n_25044), .Y (n_25229));
MX2X1 g57717(.A (n_25042), .B (n_25043), .S0 (n_24923), .Y (n_25228));
MX2X1 g57718(.A (n_24759), .B (n_24758), .S0 (n_25041), .Y (n_25227));
MX2X1 g57719(.A (n_24964), .B (n_24965), .S0 (n_24592), .Y (n_25226));
DFFX1 u0_w_reg[2][21] (.CK (clk), .D (n_25127), .Q (w2[21] ), .QN());
DFFX1 u0_w_reg[0][27] (.CK (clk), .D (n_25125), .Q (n_2430), .QN ());
DFFX1 u0_w_reg[1][27] (.CK (clk), .D (n_25124), .Q (), .QN (w1[27]));
DFFX1 u0_w_reg[2][27] (.CK (clk), .D (n_25122), .Q (w2[27] ), .QN());
DFFX1 u0_w_reg[2][11] (.CK (clk), .D (n_25120), .Q (w2[11] ), .QN());
DFFX1 u0_w_reg[3][27] (.CK (clk), .D (n_25121), .Q (n_362), .QN ());
DFFX1 u0_w_reg[3][24] (.CK (clk), .D (n_25117), .Q (n_1138), .QN ());
NAND2X1 g57761(.A (n_25104), .B (n_25269), .Y (n_25787));
NAND2X1 g57763(.A (n_25110), .B (n_25283), .Y (n_25721));
MX2X1 g57766(.A (n_24878), .B (n_24877), .S0 (n_25025), .Y (n_25223));
XOR2X1 g57772(.A (n_24893), .B (n_24982), .Y (n_25222));
MX2X1 g57776(.A (n_24579), .B (n_24580), .S0 (n_25016), .Y (n_25221));
MX2X1 g57778(.A (n_25022), .B (n_25021), .S0 (n_25010), .Y (n_25220));
MX2X1 g57784(.A (n_25012), .B (n_25013), .S0 (n_25007), .Y (n_25219));
MX2X1 g57785(.A (n_24200), .B (n_24199), .S0 (n_25008), .Y (n_25218));
MX2X1 g57821(.A (n_24959), .B (n_24958), .S0 (n_24672), .Y (n_25217));
OAI21X1 g57838(.A0 (n_25102), .A1 (n_28336), .B0 (n_25103), .Y(n_25216));
MX2X1 g56719(.A (n_24654), .B (n_24653), .S0 (n_24966), .Y (n_25215));
OAI21X1 g56920(.A0 (n_24985), .A1 (ld_r), .B0 (n_8334), .Y (n_25214));
OAI21X1 g57269(.A0 (n_25011), .A1 (ld_r), .B0 (n_10050), .Y(n_25213));
NAND2X1 g57292(.A (n_25078), .B (n_25274), .Y (n_25704));
MX2X1 g58001(.A (n_24259), .B (n_24258), .S0 (n_24957), .Y (n_25211));
INVX1 g58005(.A (n_25209), .Y (n_25210));
OAI21X1 g57320(.A0 (n_24984), .A1 (n_25361), .B0 (n_8383), .Y(n_25208));
NAND2X1 g58017(.A (n_25074), .B (n_24997), .Y (n_25207));
NAND2X1 g58018(.A (n_25073), .B (n_24996), .Y (n_25206));
NAND2X1 g58021(.A (n_25072), .B (n_24995), .Y (n_25205));
OAI21X1 g57324(.A0 (n_24986), .A1 (n_25407), .B0 (n_8657), .Y(n_25204));
MX2X1 g57325(.A (n_24564), .B (n_23444), .S0 (n_24983), .Y (n_25203));
OAI21X1 g56671(.A0 (n_25051), .A1 (n_25332), .B0 (n_19036), .Y(n_25202));
OAI21X1 g56977(.A0 (n_24960), .A1 (n_25426), .B0 (n_8770), .Y(n_25200));
NAND2X1 g57373(.A (n_27876), .B (n_25283), .Y (n_25602));
MX2X1 g57376(.A (n_24980), .B (n_24981), .S0 (n_24968), .Y (n_25198));
MX2X1 g56981(.A (n_24576), .B (n_24577), .S0 (n_24956), .Y (n_25197));
MX2X1 g57377(.A (n_24890), .B (n_24891), .S0 (n_24967), .Y (n_25196));
NAND2X1 g56998(.A (n_25065), .B (n_25274), .Y (n_25194));
MX2X1 g57403(.A (n_24962), .B (n_24963), .S0 (n_24882), .Y (n_25193));
MX2X1 g57405(.A (n_24648), .B (n_24647), .S0 (n_24961), .Y (n_25192));
MX2X1 g57009(.A (n_24954), .B (n_24955), .S0 (n_24897), .Y (n_25191));
NAND2X2 g56683(.A (n_25112), .B (n_25283), .Y (n_25564));
NAND2X1 g56682(.A (n_25114), .B (n_25274), .Y (n_29177));
MX2X1 g57020(.A (n_25020), .B (n_25019), .S0 (n_24800), .Y (n_25188));
NAND2X1 g57029(.A (n_25062), .B (n_25274), .Y (n_25187));
NAND2X1 g57030(.A (n_25060), .B (n_25269), .Y (n_25730));
XOR2X1 g56686(.A (n_24574), .B (n_25029), .Y (n_25185));
MX2X1 g56688(.A (n_25023), .B (n_25024), .S0 (n_24585), .Y (n_25184));
MX2X1 g57063(.A (n_24787), .B (n_24786), .S0 (n_25055), .Y (n_25183));
INVX1 g57120(.A (n_25181), .Y (n_25182));
NAND2X1 g57711(.A (n_989), .B (n_25050), .Y (n_25180));
MX2X1 g56705(.A (n_24553), .B (n_24149), .S0 (n_24837), .Y (n_25179));
MX2X1 g56653(.A (n_24573), .B (n_28117), .S0 (n_24793), .Y (n_25178));
DFFX1 u0_w_reg[2][29] (.CK (clk), .D (n_25054), .Q (), .QN (n_1018));
DFFX1 u0_w_reg[0][29] (.CK (clk), .D (n_25056), .Q (n_497), .QN ());
DFFX1 u0_w_reg[2][5] (.CK (clk), .D (n_25053), .Q (w2[5] ), .QN ());
DFFX1 u0_w_reg[2][3] (.CK (clk), .D (n_25049), .Q (w2[3] ), .QN ());
MX2X1 g56654(.A (n_24628), .B (n_24627), .S0 (n_24922), .Y (n_25177));
MX2X1 g56709(.A (n_24520), .B (n_24519), .S0 (n_24812), .Y (n_25176));
MX2X1 g57775(.A (n_24838), .B (n_24839), .S0 (n_24885), .Y (n_25175));
OAI21X1 g56655(.A0 (n_25027), .A1 (n_25026), .B0 (n_25028), .Y(n_25174));
OAI21X1 g57788(.A0 (n_25046), .A1 (n_25045), .B0 (n_25047), .Y(n_28604));
MX2X1 g57835(.A (key[115]), .B (n_24826), .S0 (n_229), .Y (n_25172));
MX2X1 g57836(.A (key[83]), .B (n_24825), .S0 (n_229), .Y (n_25171));
OAI21X1 g56658(.A0 (n_25034), .A1 (n_25033), .B0 (n_25035), .Y(n_25170));
MX2X1 g57837(.A (key[19]), .B (n_24823), .S0 (n_360), .Y (n_25169));
MX2X1 g57840(.A (n_24830), .B (n_24831), .S0 (n_24819), .Y (n_25168));
OAI21X1 g56659(.A0 (n_25039), .A1 (n_24321), .B0 (n_25040), .Y(n_25167));
OAI21X1 g57868(.A0 (n_25031), .A1 (n_25030), .B0 (n_25032), .Y(n_25165));
MX2X1 g57877(.A (n_24754), .B (n_24752), .S0 (n_24820), .Y (n_25164));
MX2X1 g56733(.A (n_24805), .B (n_24804), .S0 (n_23709), .Y (n_25163));
NAND2X1 g58006(.A (n_24844), .B (n_24988), .Y (n_25209));
NAND2X1 g58011(.A (n_24989), .B (n_24848), .Y (n_25162));
INVX1 g58019(.A (n_25160), .Y (n_25161));
INVX1 g58022(.A (n_28112), .Y (n_25159));
INVX1 g58027(.A (n_25156), .Y (n_25157));
NAND2X1 g58030(.A (n_24994), .B (n_24862), .Y (n_25155));
MX2X1 g57328(.A (n_24932), .B (n_24933), .S0 (n_24692), .Y (n_25154));
NAND2X1 g58044(.A (n_24999), .B (n_24870), .Y (n_25153));
MX2X1 g57330(.A (n_24817), .B (n_24818), .S0 (n_24542), .Y (n_25152));
NAND2X1 g58048(.A (n_25001), .B (n_24875), .Y (n_25151));
NAND2X1 g58050(.A (n_25000), .B (n_24872), .Y (n_25150));
NAND2X1 g58051(.A (n_24993), .B (n_24854), .Y (n_25149));
OAI21X1 g57331(.A0 (n_25005), .A1 (n_28331), .B0 (n_25006), .Y(n_25148));
OAI21X1 g57332(.A0 (n_25003), .A1 (n_25002), .B0 (n_25004), .Y(n_25147));
NAND2X1 g58053(.A (n_24991), .B (n_24851), .Y (n_25146));
MX2X1 g57352(.A (n_24685), .B (n_24684), .S0 (n_24894), .Y (n_25145));
MX2X1 g56673(.A (n_24742), .B (n_24741), .S0 (n_24925), .Y (n_25144));
MX2X1 g57362(.A (n_24889), .B (n_24888), .S0 (n_24834), .Y (n_25143));
NAND2X1 g57372(.A (n_24969), .B (n_25269), .Y (n_25824));
MX2X1 g57375(.A (n_24814), .B (n_24813), .S0 (n_24676), .Y (n_25141));
MX2X1 g56984(.A (n_24930), .B (n_24931), .S0 (n_24635), .Y (n_25140));
MX2X1 g56985(.A (n_24821), .B (n_24822), .S0 (n_24638), .Y (n_25139));
OAI21X1 g56986(.A0 (n_24973), .A1 (n_24972), .B0 (n_24974), .Y(n_25138));
MX2X1 g56676(.A (n_24785), .B (n_24784), .S0 (n_24901), .Y (n_25137));
OAI21X1 g56988(.A0 (n_24976), .A1 (n_24975), .B0 (n_24977), .Y(n_25136));
MX2X1 g57395(.A (n_24661), .B (n_24662), .S0 (n_24811), .Y (n_25135));
MX2X1 g56677(.A (n_24884), .B (n_24883), .S0 (n_24781), .Y (n_25134));
MX2X1 g56678(.A (n_24945), .B (n_24946), .S0 (n_24934), .Y (n_25133));
MX2X1 g57007(.A (n_24626), .B (n_24625), .S0 (n_24902), .Y (n_25132));
MX2X1 g56684(.A (n_24816), .B (n_24815), .S0 (n_24892), .Y (n_25131));
MX2X1 g57078(.A (n_24810), .B (n_24809), .S0 (n_24426), .Y (n_25130));
MX2X1 g57079(.A (n_24634), .B (n_24987), .S0 (n_24204), .Y (n_25129));
OAI21X1 g56694(.A0 (n_25058), .A1 (n_25057), .B0 (n_25059), .Y(n_25128));
MX2X1 g57121(.A (n_23515), .B (n_23516), .S0 (n_24771), .Y (n_25181));
MX2X1 g57712(.A (n_24769), .B (key[53]), .S0 (n_25126), .Y (n_25127));
SDFFSRX1 u0_w_reg[1][29] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_24595), .SE (n_25052), .SI (key[93]), .Q (n_645), .QN ());
DFFX1 u0_w_reg[0][30] (.CK (clk), .D (n_24944), .Q (w0[30] ), .QN());
DFFX1 u0_w_reg[1][30] (.CK (clk), .D (n_24943), .Q (), .QN(n_22833));
DFFX1 u0_w_reg[3][30] (.CK (clk), .D (n_24939), .Q (w3[30] ), .QN());
DFFX1 u0_w_reg[0][21] (.CK (clk), .D (n_24938), .Q (n_24366), .QN());
DFFX1 u0_w_reg[1][21] (.CK (clk), .D (n_24936), .Q (), .QN(n_23397));
DFFX1 u0_w_reg[2][0] (.CK (clk), .D (n_24929), .Q (w2[0] ), .QN ());
DFFX1 u0_w_reg[2][10] (.CK (clk), .D (n_24927), .Q (w2[10] ), .QN());
DFFX1 u0_w_reg[2][14] (.CK (clk), .D (n_24924), .Q (w2[14] ), .QN());
DFFX1 u0_w_reg[2][30] (.CK (clk), .D (n_24940), .Q (w2[30] ), .QN());
DFFX1 u0_w_reg[2][16] (.CK (clk), .D (n_24926), .Q (w2[16] ), .QN());
DFFX1 u0_w_reg[2][8] (.CK (clk), .D (n_24916), .Q (w2[8] ), .QN ());
DFFX1 u0_w_reg[2][15] (.CK (clk), .D (n_24918), .Q (w2[15] ), .QN());
DFFX1 u0_w_reg[3][21] (.CK (clk), .D (n_24935), .Q (w3[21] ), .QN());
DFFX1 text_out_reg[12] (.CK (clk), .D (n_24947), .Q (text_out[12]),.QN ());
MX2X1 g57768(.A (n_24740), .B (key[123]), .S0 (n_25123), .Y(n_25125));
MX2X1 g57769(.A (n_24739), .B (key[91]), .S0 (n_25123), .Y (n_25124));
MX2X1 g57770(.A (n_24738), .B (key[59]), .S0 (n_25123), .Y (n_25122));
MX2X1 g57771(.A (n_24737), .B (key[27]), .S0 (n_698), .Y (n_25121));
MX2X1 g57779(.A (n_24730), .B (key[43]), .S0 (n_24937), .Y (n_25120));
MX2X1 g56656(.A (n_24760), .B (n_24761), .S0 (n_24451), .Y (n_25119));
MX2X1 g56657(.A (n_24671), .B (n_24670), .S0 (n_24455), .Y (n_25118));
NAND2X1 g57816(.A (n_1239), .B (n_24903), .Y (n_25117));
NAND2X1 g56716(.A (n_24914), .B (n_24756), .Y (n_25116));
MX2X1 g57820(.A (n_24699), .B (n_24840), .S0 (n_24690), .Y (n_25115));
MX2X1 g56717(.A (n_24096), .B (n_24094), .S0 (n_24680), .Y (n_25114));
NAND2X1 g57831(.A (n_24905), .B (n_24749), .Y (n_25113));
OAI21X1 g56718(.A0 (n_24920), .A1 (n_24919), .B0 (n_24921), .Y(n_25112));
NAND2X1 g57834(.A (n_24904), .B (n_24745), .Y (n_25111));
OAI21X1 g57839(.A0 (n_24907), .A1 (n_24906), .B0 (n_24908), .Y(n_25110));
NAND2X1 g57851(.A (n_24751), .B (n_24910), .Y (n_25109));
NAND2X1 g57852(.A (n_24750), .B (n_24909), .Y (n_25108));
MX2X1 g57853(.A (n_24689), .B (n_24688), .S0 (n_24452), .Y (n_25107));
MX2X1 g57862(.A (n_24617), .B (n_24618), .S0 (n_24346), .Y (n_25106));
XOR2X1 g57873(.A (n_1843), .B (n_24673), .Y (n_25105));
OAI21X1 g57875(.A0 (n_24912), .A1 (n_24911), .B0 (n_24913), .Y(n_25104));
NAND2X1 g57938(.A (n_25102), .B (n_28336), .Y (n_25103));
INVX1 g57953(.A (n_25100), .Y (n_25101));
INVX1 g57955(.A (n_25098), .Y (n_25099));
INVX1 g57957(.A (n_25096), .Y (n_25097));
NAND2X1 g57959(.A (n_24701), .B (n_24842), .Y (n_25095));
NAND2X1 g57973(.A (n_24703), .B (n_24843), .Y (n_25094));
INVX1 g57997(.A (n_25092), .Y (n_25093));
INVX1 g58003(.A (n_25090), .Y (n_25091));
NAND2X1 g58014(.A (n_24847), .B (n_24708), .Y (n_25089));
NAND2X1 g58016(.A (n_24707), .B (n_24845), .Y (n_25088));
NAND2X2 g58020(.A (n_24868), .B (n_24717), .Y (n_25160));
NAND2X1 g58024(.A (n_24866), .B (n_24715), .Y (n_25087));
INVX1 g58025(.A (n_25085), .Y (n_25086));
NAND2X2 g58028(.A (n_24864), .B (n_24712), .Y (n_25156));
NAND2X1 g58029(.A (n_24863), .B (n_24719), .Y (n_25084));
NAND2X1 g58031(.A (n_24861), .B (n_24711), .Y (n_25083));
NAND2X1 g58032(.A (n_24859), .B (n_24710), .Y (n_25082));
NAND2X1 g58033(.A (n_24857), .B (n_24709), .Y (n_25081));
NAND2X1 g58034(.A (n_24855), .B (n_24718), .Y (n_25080));
MX2X1 g58035(.A (n_24406), .B (n_24405), .S0 (n_25076), .Y (n_25079));
OAI21X1 g57329(.A0 (n_24880), .A1 (n_24879), .B0 (n_24881), .Y(n_25078));
MX2X1 g58046(.A (n_24505), .B (n_24212), .S0 (n_25076), .Y (n_25077));
NAND2X1 g58049(.A (n_24873), .B (n_24722), .Y (n_25075));
NAND2X1 g58125(.A (n_24998), .B (n_24953), .Y (n_25074));
NAND2X1 g58129(.A (n_24990), .B (n_24951), .Y (n_25073));
NAND2X1 g58133(.A (n_24992), .B (n_24949), .Y (n_25072));
MX2X1 g57393(.A (n_24899), .B (n_24898), .S0 (n_24669), .Y (n_25071));
MX2X1 g57404(.A (n_24687), .B (n_24686), .S0 (n_24655), .Y (n_25067));
MX2X1 g57032(.A (n_24644), .B (n_24643), .S0 (n_24619), .Y (n_25066));
OAI21X1 g57040(.A0 (n_24807), .A1 (n_24806), .B0 (n_24808), .Y(n_25065));
MX2X1 g57051(.A (n_24896), .B (n_24895), .S0 (n_24615), .Y (n_25064));
MX2X1 g57053(.A (n_24791), .B (n_24792), .S0 (n_24640), .Y (n_25063));
OAI21X1 g57058(.A0 (n_24795), .A1 (n_28775), .B0 (n_24796), .Y(n_25062));
MX2X1 g57062(.A (n_24537), .B (n_24536), .S0 (n_24790), .Y (n_25061));
OAI21X1 g57068(.A0 (n_24798), .A1 (n_24797), .B0 (n_24799), .Y(n_25060));
NAND2X1 g56703(.A (n_25058), .B (n_25057), .Y (n_25059));
MX2X1 g57709(.A (n_24596), .B (key[125]), .S0 (n_25123), .Y(n_25056));
MX2X1 g57124(.A (n_24184), .B (n_24183), .S0 (n_24467), .Y (n_25055));
MX2X1 g57710(.A (n_24594), .B (key[61]), .S0 (n_619), .Y (n_25054));
MX2X1 g57716(.A (n_24589), .B (key[37]), .S0 (ld), .Y (n_25053));
DFFX1 u0_w_reg[2][12] (.CK (clk), .D (n_24780), .Q (w2[12] ), .QN());
DFFX1 u0_w_reg[0][24] (.CK (clk), .D (n_24779), .Q (n_22981), .QN());
DFFX1 u0_w_reg[0][31] (.CK (clk), .D (n_24777), .Q (w0[31] ), .QN());
SDFFSRX1 u0_w_reg[1][24] (.RN (1'b1), .SN (1'b1), .CK (clk), .D(n_24372), .SE (n_25052), .SI (key[88]), .Q (w1[24] ), .QN ());
DFFX1 u0_w_reg[1][31] (.CK (clk), .D (n_24776), .Q (), .QN (w1[31]));
DFFX1 u0_w_reg[2][24] (.CK (clk), .D (n_24775), .Q (w2[24] ), .QN());
MX2X1 g56708(.A (n_24543), .B (n_24544), .S0 (n_24517), .Y (n_25051));
DFFX1 u0_w_reg[2][31] (.CK (clk), .D (n_24773), .Q (w2[31] ), .QN());
DFFX1 u0_w_reg[3][31] (.CK (clk), .D (n_24772), .Q (w3[31] ), .QN());
DFFX1 u0_w_reg[0][5] (.CK (clk), .D (n_24768), .Q (n_925), .QN ());
DFFX1 u0_w_reg[2][22] (.CK (clk), .D (n_24764), .Q (w2[22] ), .QN());
DFFX1 u0_w_reg[2][6] (.CK (clk), .D (n_24763), .Q (w2[6] ), .QN ());
DFFX1 u0_w_reg[3][5] (.CK (clk), .D (n_24765), .Q (w3[5] ), .QN ());
DFFX1 u0_w_reg[0][11] (.CK (clk), .D (n_24734), .Q (n_23363), .QN());
DFFX1 u0_w_reg[1][11] (.CK (clk), .D (n_24733), .Q (n_546), .QN ());
DFFX1 u0_w_reg[2][17] (.CK (clk), .D (n_24724), .Q (w2[17] ), .QN());
DFFX1 u0_w_reg[2][9] (.CK (clk), .D (n_24723), .Q (w2[9] ), .QN ());
DFFX1 u0_w_reg[3][11] (.CK (clk), .D (n_24731), .Q (w3[11] ), .QN());
DFFX1 text_out_reg[125] (.CK (clk), .D (n_24666), .Q(text_out[125]), .QN ());
DFFX1 text_out_reg[44] (.CK (clk), .D (n_24632), .Q (text_out[44]),.QN ());
NAND2X1 g57758(.A (n_24770), .B (n_360), .Y (n_25050));
MX2X1 g57777(.A (n_24563), .B (key[35]), .S0 (n_698), .Y (n_25049));
NAND2X1 g57803(.A (n_25046), .B (n_25045), .Y (n_25047));
NAND2X1 g57833(.A (n_24747), .B (n_24746), .Y (n_25044));
INVX1 g57844(.A (n_25042), .Y (n_25043));
NAND2X1 g57850(.A (n_24753), .B (n_24755), .Y (n_25041));
NAND2X1 g56661(.A (n_25039), .B (n_24394), .Y (n_25040));
NAND2X1 g56663(.A (n_25034), .B (n_25033), .Y (n_25035));
NAND2X1 g57929(.A (n_25031), .B (n_25030), .Y (n_25032));
MX2X1 g56732(.A (n_23908), .B (n_23907), .S0 (n_24480), .Y (n_25029));
NAND2X1 g56664(.A (n_25027), .B (n_25026), .Y (n_25028));
MX2X1 g57954(.A (n_24442), .B (n_24443), .S0 (n_26216), .Y (n_25100));
MX2X1 g57956(.A (n_24440), .B (n_24441), .S0 (n_24064), .Y (n_25098));
MX2X1 g57958(.A (n_24438), .B (n_24439), .S0 (n_24063), .Y (n_25096));
NAND2X1 g57962(.A (n_24697), .B (n_24698), .Y (n_25025));
INVX1 g57964(.A (n_25023), .Y (n_25024));
INVX1 g57987(.A (n_25021), .Y (n_25022));
INVX1 g57995(.A (n_25019), .Y (n_25020));
NAND2X1 g57998(.A (n_24558), .B (n_24706), .Y (n_25092));
INVX1 g57999(.A (n_25017), .Y (n_25018));
NAND2X1 g58004(.A (n_24557), .B (n_24705), .Y (n_25090));
MX2X1 g58009(.A (n_25015), .B (n_25014), .S0 (n_24478), .Y (n_25016));
NAND2X1 g58026(.A (n_24713), .B (n_24560), .Y (n_25085));
INVX1 g58038(.A (n_25012), .Y (n_25013));
XOR2X1 g57327(.A (n_24359), .B (n_24540), .Y (n_25011));
NAND2X1 g58041(.A (n_24720), .B (n_24561), .Y (n_25010));
MX2X1 g58045(.A (n_24301), .B (n_23919), .S0 (n_24871), .Y (n_25009));
MX2X1 g58047(.A (n_24610), .B (n_24609), .S0 (n_24471), .Y (n_25008));
MX2X1 g58052(.A (n_24645), .B (n_24509), .S0 (n_24874), .Y (n_25007));
NAND2X1 g57333(.A (n_28331), .B (n_25005), .Y (n_25006));
NAND2X1 g57334(.A (n_25003), .B (n_25002), .Y (n_25004));
NAND2X1 g58113(.A (n_24420), .B (n_24629), .Y (n_25001));
NAND2X1 g58117(.A (n_24193), .B (n_24624), .Y (n_25000));
NAND2X1 g58124(.A (n_24998), .B (n_24630), .Y (n_24999));
NAND2X1 g58126(.A (n_24869), .B (n_24952), .Y (n_24997));
NAND2X1 g58132(.A (n_24850), .B (n_24950), .Y (n_24996));
NAND2X1 g58136(.A (n_24853), .B (n_24948), .Y (n_24995));
DFFX1 u0_w_reg[1][5] (.CK (clk), .D (n_24766), .Q (), .QN (w1[5] ));
NAND2X1 g58144(.A (n_24700), .B (n_24637), .Y (n_24994));
NAND2X1 g58152(.A (n_24992), .B (n_24631), .Y (n_24993));
DFFX1 u0_w_reg[2][13] (.CK (clk), .D (n_24757), .Q (w2[13] ), .QN());
NAND2X1 g58155(.A (n_24990), .B (n_24623), .Y (n_24991));
NAND2X1 g58157(.A (n_24865), .B (n_24639), .Y (n_24989));
NAND2X1 g58172(.A (n_24987), .B (n_24577), .Y (n_24988));
XOR2X1 g57379(.A (n_24566), .B (n_24525), .Y (n_24986));
XOR2X1 g56983(.A (n_24362), .B (n_24488), .Y (n_24985));
MX2X1 g57383(.A (n_24523), .B (n_24524), .S0 (n_24538), .Y (n_24984));
MX2X1 g57384(.A (n_24453), .B (n_24454), .S0 (n_24123), .Y (n_24983));
NAND2X1 g58230(.A (n_24646), .B (n_24510), .Y (n_24982));
INVX1 g58233(.A (n_24980), .Y (n_24981));
INVX1 g58235(.A (n_24978), .Y (n_24979));
NAND2X1 g56990(.A (n_24976), .B (n_24975), .Y (n_24977));
NAND2X1 g56991(.A (n_24973), .B (n_24972), .Y (n_24974));
OAI21X1 g57410(.A0 (n_24682), .A1 (n_24681), .B0 (n_24683), .Y(n_24969));
MX2X1 g57419(.A (n_24486), .B (n_24485), .S0 (n_24298), .Y (n_24968));
MX2X1 g57420(.A (n_24483), .B (n_24704), .S0 (n_24072), .Y (n_24967));
MX2X1 g56770(.A (n_23945), .B (n_28564), .S0 (n_24464), .Y (n_24966));
INVX1 g58325(.A (n_24964), .Y (n_24965));
INVX1 g57463(.A (n_24962), .Y (n_24963));
MX2X1 g57465(.A (n_24048), .B (n_24047), .S0 (n_24469), .Y (n_24961));
XOR2X1 g57033(.A (n_24578), .B (n_24460), .Y (n_24960));
INVX1 g58433(.A (n_24958), .Y (n_24959));
NAND2X1 g58459(.A (n_24616), .B (n_24450), .Y (n_24957));
MX2X1 g57042(.A (n_24456), .B (n_24457), .S0 (n_23997), .Y (n_24956));
INVX1 g57064(.A (n_24954), .Y (n_24955));
INVX1 g58867(.A (n_24952), .Y (n_24953));
INVX1 g58872(.A (n_24950), .Y (n_24951));
INVX1 g58879(.A (n_24948), .Y (n_24949));
XOR2X1 g58913(.A (n_5306), .B (n_24169), .Y (n_24947));
DFFX1 u0_w_reg[1][3] (.CK (clk), .D (n_24570), .Q (w1[3] ), .QN ());
DFFX1 u0_w_reg[0][3] (.CK (clk), .D (n_24571), .Q (w0[3] ), .QN ());
DFFX1 u0_w_reg[3][3] (.CK (clk), .D (n_24568), .Q (w3[3] ), .QN ());
DFFX1 u0_w_reg[2][4] (.CK (clk), .D (n_24549), .Q (w2[4] ), .QN ());
DFFX1 u0_w_reg[1][28] (.CK (clk), .D (n_24547), .Q (), .QN (n_1308));
DFFX1 u0_w_reg[3][28] (.CK (clk), .D (n_24545), .Q (w3[28] ), .QN());
DFFX1 text_out_reg[93] (.CK (clk), .D (n_24515), .Q (text_out[93]),.QN ());
DFFX1 u0_w_reg[0][0] (.CK (clk), .D (n_24535), .Q (w0[0] ), .QN ());
DFFX1 text_out_reg[61] (.CK (clk), .D (n_24516), .Q (text_out[61]),.QN ());
DFFX1 u0_w_reg[0][16] (.CK (clk), .D (n_24534), .Q (n_424), .QN ());
DFFX1 u0_w_reg[1][0] (.CK (clk), .D (n_24533), .Q (), .QN (w1[0] ));
DFFX1 u0_w_reg[3][0] (.CK (clk), .D (n_24529), .Q (w3[0] ), .QN ());
DFFX1 u0_w_reg[1][16] (.CK (clk), .D (n_24532), .Q (), .QN (w1[16]));
DFFX1 u0_w_reg[3][16] (.CK (clk), .D (n_24528), .Q (w3[16] ), .QN());
DFFX1 text_out_reg[101] (.CK (clk), .D (n_24526), .Q(text_out[101]), .QN ());
DFFX1 text_out_reg[108] (.CK (clk), .D (n_24482), .Q(text_out[108]), .QN ());
DFFX1 text_out_reg[43] (.CK (clk), .D (n_24487), .Q (text_out[43]),.QN ());
DFFX1 text_out_reg[109] (.CK (clk), .D (n_24459), .Q(text_out[109]), .QN ());
DFFX1 text_out_reg[117] (.CK (clk), .D (n_24458), .Q(text_out[117]), .QN ());
DFFX1 text_out_reg[76] (.CK (clk), .D (n_24481), .Q (text_out[76]),.QN ());
DFFX1 text_out_reg[111] (.CK (clk), .D (n_24602), .Q(text_out[111]), .QN ());
DFFX1 text_out_reg[48] (.CK (clk), .D (n_24606), .Q (text_out[48]),.QN ());
DFFX1 text_out_reg[80] (.CK (clk), .D (n_24604), .Q (text_out[80]),.QN ());
DFFX1 text_out_reg[112] (.CK (clk), .D (n_24608), .Q(text_out[112]), .QN ());
DFFX1 text_out_reg[46] (.CK (clk), .D (n_24588), .Q (text_out[46]),.QN ());
DFFX1 text_out_reg[126] (.CK (clk), .D (n_24591), .Q(text_out[126]), .QN ());
DFFX1 text_out_reg[10] (.CK (clk), .D (n_24590), .Q (text_out[10]),.QN ());
INVX1 g56713(.A (n_24945), .Y (n_24946));
MX2X1 g57807(.A (n_24373), .B (key[126]), .S0 (n_24778), .Y(n_24944));
MX2X1 g57810(.A (n_24371), .B (key[94]), .S0 (n_24937), .Y (n_24943));
XOR2X1 g56715(.A (n_24134), .B (n_24430), .Y (n_24941));
MX2X1 g57814(.A (n_24370), .B (key[62]), .S0 (n_1914), .Y (n_24940));
MX2X1 g57818(.A (n_24369), .B (key[30]), .S0 (n_24937), .Y (n_24939));
MX2X1 g57822(.A (n_24367), .B (key[117]), .S0 (n_24937), .Y(n_24938));
MX2X1 g57823(.A (n_24365), .B (key[85]), .S0 (n_24937), .Y (n_24936));
MX2X1 g57824(.A (n_24363), .B (key[21]), .S0 (n_24915), .Y (n_24935));
NAND2X1 g57832(.A (n_24583), .B (n_24395), .Y (n_24934));
MX2X1 g57845(.A (n_23221), .B (n_28052), .S0 (n_24326), .Y (n_25042));
INVX1 g57846(.A (n_24932), .Y (n_24933));
INVX1 g57848(.A (n_24930), .Y (n_24931));
MX2X1 g57854(.A (n_24330), .B (key[32]), .S0 (n_619), .Y (n_24929));
MX2X1 g57855(.A (n_24331), .B (key[42]), .S0 (n_619), .Y (n_24927));
MX2X1 g57856(.A (n_24329), .B (key[48]), .S0 (n_619), .Y (n_24926));
NAND2X1 g56721(.A (n_24593), .B (n_24407), .Y (n_24925));
MX2X1 g57859(.A (n_24327), .B (key[46]), .S0 (n_24548), .Y (n_24924));
MX2X1 g57863(.A (n_23196), .B (n_23507), .S0 (n_24344), .Y (n_24923));
NAND2X1 g57869(.A (n_24584), .B (n_24396), .Y (n_24922));
NAND2X1 g56726(.A (n_24920), .B (n_24919), .Y (n_24921));
MX2X1 g57872(.A (n_24323), .B (key[47]), .S0 (n_619), .Y (n_24918));
MX2X1 g57874(.A (n_24322), .B (key[40]), .S0 (n_24915), .Y (n_24916));
NAND2X1 g56727(.A (n_24612), .B (n_24133), .Y (n_24914));
NAND2X1 g57928(.A (n_24912), .B (n_24911), .Y (n_24913));
NAND2X1 g57935(.A (n_23219), .B (n_24104), .Y (n_24910));
NAND2X1 g57937(.A (n_23537), .B (n_24514), .Y (n_24909));
NAND2X1 g57939(.A (n_24907), .B (n_24906), .Y (n_24908));
NAND2X1 g57940(.A (n_27488), .B (n_22596), .Y (n_24905));
NAND2X1 g57946(.A (n_24104), .B (n_22502), .Y (n_24904));
NAND2X1 g57948(.A (n_24541), .B (n_3721), .Y (n_24903));
NAND2X1 g57951(.A (n_24556), .B (n_24555), .Y (n_24902));
NAND2X1 g57952(.A (n_24554), .B (n_24552), .Y (n_24901));
MX2X1 g57961(.A (n_24896), .B (n_24895), .S0 (n_24858), .Y (n_24897));
NAND2X1 g57963(.A (n_24551), .B (n_24550), .Y (n_24894));
MX2X1 g57965(.A (n_24229), .B (n_24230), .S0 (n_23741), .Y (n_25023));
XOR2X1 g57972(.A (n_25518), .B (n_25517), .Y (n_24893));
MX2X1 g56737(.A (n_19433), .B (n_16480), .S0 (n_24270), .Y (n_24892));
MX2X1 g57988(.A (n_23739), .B (n_23738), .S0 (n_24297), .Y (n_25021));
INVX1 g57989(.A (n_24890), .Y (n_24891));
INVX1 g57991(.A (n_24888), .Y (n_24889));
INVX1 g57993(.A (n_24886), .Y (n_24887));
MX2X1 g57996(.A (n_24288), .B (n_24287), .S0 (n_24296), .Y (n_25019));
MX2X1 g58000(.A (n_24060), .B (n_24059), .S0 (n_24295), .Y (n_25017));
MX2X1 g58002(.A (n_25015), .B (n_25014), .S0 (n_24702), .Y (n_24885));
INVX1 g58007(.A (n_24883), .Y (n_24884));
NAND2X1 g58039(.A (n_24562), .B (n_24382), .Y (n_25012));
MX2X1 g58054(.A (n_24507), .B (n_24213), .S0 (n_24721), .Y (n_24882));
NAND2X1 g57335(.A (n_24880), .B (n_24879), .Y (n_24881));
INVX1 g58060(.A (n_24877), .Y (n_24878));
MX2X1 g58062(.A (n_23265), .B (n_23264), .S0 (n_24256), .Y (n_24876));
NAND2X1 g58114(.A (n_24419), .B (n_24874), .Y (n_24875));
NAND2X1 g58115(.A (n_24195), .B (n_24468), .Y (n_24873));
NAND2X1 g58118(.A (n_24192), .B (n_24871), .Y (n_24872));
NAND2X1 g58123(.A (n_24869), .B (n_24856), .Y (n_24870));
NAND2X1 g58130(.A (n_24502), .B (n_24030), .Y (n_24868));
NAND2X1 g58137(.A (n_24865), .B (n_24614), .Y (n_24866));
NAND2X1 g58141(.A (n_24498), .B (n_24026), .Y (n_24864));
NAND2X1 g58143(.A (n_24852), .B (n_24303), .Y (n_24863));
NAND2X1 g58145(.A (n_24841), .B (n_24636), .Y (n_24862));
NAND2X1 g58146(.A (n_25822), .B (n_24860), .Y (n_24861));
NAND2X1 g58148(.A (n_24858), .B (n_24492), .Y (n_24859));
NAND2X1 g58150(.A (n_24856), .B (n_23622), .Y (n_24857));
NAND2X1 g58151(.A (n_24083), .B (n_24849), .Y (n_24855));
NAND2X1 g58153(.A (n_24853), .B (n_24852), .Y (n_24854));
NAND2X1 g58156(.A (n_24850), .B (n_24849), .Y (n_24851));
NAND2X1 g58158(.A (n_24714), .B (n_26780), .Y (n_24848));
NAND2X1 g58159(.A (n_26780), .B (n_24310), .Y (n_24847));
NAND2X1 g58166(.A (n_24490), .B (n_23795), .Y (n_24845));
NAND2X1 g58171(.A (n_24634), .B (n_24576), .Y (n_24844));
NAND2X1 g58180(.A (n_24484), .B (n_23640), .Y (n_24843));
NAND2X1 g58182(.A (n_24841), .B (n_24840), .Y (n_24842));
INVX1 g58200(.A (n_24838), .Y (n_24839));
MX2X1 g56760(.A (n_24414), .B (n_24413), .S0 (n_23936), .Y (n_24837));
DFFX1 u0_w_reg[3][26] (.CK (clk), .D (n_24597), .Q (w3[26] ), .QN());
INVX1 g58231(.A (n_24835), .Y (n_24836));
NAND2X1 g58234(.A (n_24508), .B (n_24300), .Y (n_24980));
NAND2X2 g58236(.A (n_24506), .B (n_24299), .Y (n_24978));
NAND2X1 g57397(.A (n_24527), .B (n_24351), .Y (n_24834));
INVX1 g57398(.A (n_24832), .Y (n_24833));
XOR2X1 g58241(.A (n_24435), .B (n_23188), .Y (n_25102));
INVX1 g58246(.A (n_24830), .Y (n_24831));
NAND2X1 g57425(.A (n_24518), .B (n_24328), .Y (n_24827));
XOR2X1 g58287(.A (n_24266), .B (n_24824), .Y (n_24826));
XOR2X1 g58291(.A (n_1797), .B (n_24824), .Y (n_24825));
XOR2X1 g58296(.A (n_19345), .B (n_24824), .Y (n_24823));
DFFX1 u0_w_reg[1][26] (.CK (clk), .D (n_24600), .Q (), .QN(n_23053));
DFFX1 u0_w_reg[2][26] (.CK (clk), .D (n_24598), .Q (w2[26] ), .QN());
INVX1 g58312(.A (n_24821), .Y (n_24822));
MX2X1 g58319(.A (n_24397), .B (n_24398), .S0 (n_23898), .Y (n_24820));
NAND2X1 g58326(.A (n_24313), .B (n_24511), .Y (n_24964));
MX2X1 g58327(.A (n_2560), .B (w0[7] ), .S0 (n_24425), .Y (n_24819));
INVX1 g58328(.A (n_24817), .Y (n_24818));
MX2X1 g57464(.A (n_23354), .B (n_23355), .S0 (n_24284), .Y (n_24962));
INVX1 g58431(.A (n_24815), .Y (n_24816));
NAND2X1 g58434(.A (n_24445), .B (n_24234), .Y (n_24958));
INVX1 g58435(.A (n_24813), .Y (n_24814));
NAND2X1 g58438(.A (n_24446), .B (n_24237), .Y (n_24812));
NAND2X1 g58460(.A (n_24448), .B (n_24242), .Y (n_24811));
INVX1 g58512(.A (n_24809), .Y (n_24810));
NAND2X1 g57050(.A (n_24807), .B (n_24806), .Y (n_24808));
INVX1 g58519(.A (n_24804), .Y (n_24805));
INVX1 g57054(.A (n_24801), .Y (n_24802));
NAND2X1 g57057(.A (n_24461), .B (n_24262), .Y (n_24800));
DFFX1 u0_w_reg[0][26] (.CK (clk), .D (n_24601), .Q (w0[26] ), .QN());
NAND2X1 g57065(.A (n_24463), .B (n_24268), .Y (n_24954));
NAND2X1 g57071(.A (n_24798), .B (n_24797), .Y (n_24799));
NAND2X1 g57074(.A (n_24795), .B (n_28775), .Y (n_24796));
NAND2X1 g57084(.A (n_24447), .B (n_24238), .Y (n_24794));
XOR2X1 g56696(.A (n_25800), .B (n_25799), .Y (n_24793));
INVX1 g57125(.A (n_24791), .Y (n_24792));
MX2X1 g57127(.A (n_28822), .B (n_28820), .S0 (n_24187), .Y (n_24790));
OAI21X1 g58868(.A0 (n_24605), .A1 (n_24289), .B0 (n_24418), .Y(n_24952));
OAI21X1 g58873(.A0 (n_24603), .A1 (n_26634), .B0 (n_24417), .Y(n_24950));
INVX1 g57130(.A (n_24788), .Y (n_24789));
OAI21X1 g58880(.A0 (n_24607), .A1 (n_24496), .B0 (n_24416), .Y(n_24948));
INVX1 g57132(.A (n_24786), .Y (n_24787));
INVX1 g56706(.A (n_24784), .Y (n_24785));
INVX1 g57136(.A (n_24782), .Y (n_24783));
DFFX1 text_out_reg[0] (.CK (clk), .D (n_24324), .Q (text_out[0]),.QN ());
DFFX1 text_out_reg[4] (.CK (clk), .D (n_24360), .Q (text_out[4]),.QN ());
DFFX1 text_out_reg[6] (.CK (clk), .D (n_24385), .Q (text_out[6]),.QN ());
DFFX1 text_out_reg[32] (.CK (clk), .D (n_24437), .Q (text_out[32]),.QN ());
DFFX1 u0_w_reg[3][14] (.CK (clk), .D (n_24347), .Q (w3[14] ), .QN());
DFFX1 text_out_reg[64] (.CK (clk), .D (n_24318), .Q (text_out[64]),.QN ());
DFFX1 u0_w_reg[2][18] (.CK (clk), .D (n_24411), .Q (w2[18] ), .QN());
DFFX1 u0_w_reg[2][2] (.CK (clk), .D (n_24410), .Q (w2[2] ), .QN ());
DFFX1 u0_w_reg[2][23] (.CK (clk), .D (n_24387), .Q (w2[23] ), .QN());
DFFX1 u0_w_reg[2][20] (.CK (clk), .D (n_24376), .Q (w2[20] ), .QN());
DFFX1 u0_w_reg[2][28] (.CK (clk), .D (n_24374), .Q (w2[28] ), .QN());
DFFX1 u0_w_reg[0][10] (.CK (clk), .D (n_24357), .Q (w0[10] ), .QN());
DFFX1 u0_w_reg[0][13] (.CK (clk), .D (n_24343), .Q (w0[13] ), .QN());
DFFX1 u0_w_reg[0][15] (.CK (clk), .D (n_24342), .Q (n_23580), .QN());
DFFX1 u0_w_reg[0][8] (.CK (clk), .D (n_24341), .Q (w0[8] ), .QN ());
DFFX1 u0_w_reg[1][13] (.CK (clk), .D (n_24340), .Q (), .QN(n_23096));
DFFX1 u0_w_reg[1][14] (.CK (clk), .D (n_24349), .Q (w1[14] ), .QN());
DFFX1 u0_w_reg[1][15] (.CK (clk), .D (n_24338), .Q (w1[15] ), .QN());
DFFX1 u0_w_reg[1][10] (.CK (clk), .D (n_24355), .Q (w1[10] ), .QN());
DFFX1 u0_w_reg[1][8] (.CK (clk), .D (n_24337), .Q (n_23567), .QN ());
DFFX1 u0_w_reg[3][10] (.CK (clk), .D (n_24352), .Q (w3[10] ), .QN());
DFFX1 u0_w_reg[3][13] (.CK (clk), .D (n_24335), .Q (w3[13] ), .QN());
DFFX1 u0_w_reg[3][15] (.CK (clk), .D (n_24333), .Q (w3[15] ), .QN());
DFFX1 u0_w_reg[3][8] (.CK (clk), .D (n_24332), .Q (w3[8] ), .QN ());
DFFX1 text_out_reg[29] (.CK (clk), .D (n_24325), .Q (text_out[29]),.QN ());
DFFX1 text_out_reg[51] (.CK (clk), .D (n_24261), .Q (text_out[51]),.QN ());
DFFX1 text_out_reg[45] (.CK (clk), .D (n_24252), .Q (text_out[45]),.QN ());
DFFX1 text_out_reg[105] (.CK (clk), .D (n_24257), .Q(text_out[105]), .QN ());
DFFX1 text_out_reg[104] (.CK (clk), .D (n_24278), .Q(text_out[104]), .QN ());
DFFX1 text_out_reg[77] (.CK (clk), .D (n_24251), .Q (text_out[77]),.QN ());
DFFX1 text_out_reg[13] (.CK (clk), .D (n_24254), .Q (text_out[13]),.QN ());
DFFX1 text_out_reg[115] (.CK (clk), .D (n_24267), .Q(text_out[115]), .QN ());
DFFX1 text_out_reg[19] (.CK (clk), .D (n_24264), .Q (text_out[19]),.QN ());
DFFX1 text_out_reg[47] (.CK (clk), .D (n_24423), .Q (text_out[47]),.QN ());
DFFX1 text_out_reg[42] (.CK (clk), .D (n_24424), .Q (text_out[42]),.QN ());
DFFX1 text_out_reg[79] (.CK (clk), .D (n_24421), .Q (text_out[79]),.QN ());
DFFX1 text_out_reg[74] (.CK (clk), .D (n_24422), .Q (text_out[74]),.QN ());
DFFX1 text_out_reg[100] (.CK (clk), .D (n_24433), .Q(text_out[100]), .QN ());
DFFX1 text_out_reg[62] (.CK (clk), .D (n_24404), .Q (text_out[62]),.QN ());
DFFX1 text_out_reg[94] (.CK (clk), .D (n_24403), .Q (text_out[94]),.QN ());
DFFX1 text_out_reg[110] (.CK (clk), .D (n_24401), .Q(text_out[110]), .QN ());
DFFX1 text_out_reg[78] (.CK (clk), .D (n_24400), .Q (text_out[78]),.QN ());
DFFX1 text_out_reg[121] (.CK (clk), .D (n_24386), .Q(text_out[121]), .QN ());
DFFX1 text_out_reg[124] (.CK (clk), .D (n_24383), .Q(text_out[124]), .QN ());
XOR2X1 g56710(.A (n_24131), .B (n_23702), .Y (n_24781));
MX2X1 g57804(.A (n_24144), .B (key[44]), .S0 (n_24937), .Y (n_24780));
MX2X1 g57805(.A (n_24143), .B (key[120]), .S0 (n_24778), .Y(n_24779));
MX2X1 g56714(.A (n_4750), .B (n_790), .S0 (n_24135), .Y (n_24945));
MX2X1 g57808(.A (n_24142), .B (key[127]), .S0 (n_24599), .Y(n_24777));
MX2X1 g57811(.A (n_24141), .B (key[95]), .S0 (n_24937), .Y (n_24776));
MX2X1 g57812(.A (n_24140), .B (key[56]), .S0 (n_1914), .Y (n_24775));
MX2X1 g57815(.A (n_24139), .B (key[63]), .S0 (n_1914), .Y (n_24773));
MX2X1 g57819(.A (n_24138), .B (key[31]), .S0 (n_24937), .Y (n_24772));
NAND2X1 g57203(.A (n_24402), .B (n_24170), .Y (n_24771));
NAND2X1 g57828(.A (n_24393), .B (n_24391), .Y (n_24770));
XOR2X1 g57829(.A (n_1562), .B (n_24136), .Y (n_24769));
MX2X1 g57841(.A (n_24120), .B (key[101]), .S0 (ld), .Y (n_24768));
MX2X1 g57842(.A (n_24118), .B (key[69]), .S0 (ld), .Y (n_24766));
MX2X1 g57843(.A (n_24116), .B (key[5]), .S0 (n_25126), .Y (n_24765));
MX2X1 g57847(.A (n_23219), .B (n_28904), .S0 (n_24112), .Y (n_24932));
MX2X1 g57849(.A (n_23537), .B (n_27068), .S0 (n_24109), .Y (n_24930));
MX2X1 g57860(.A (n_24114), .B (key[54]), .S0 (n_1890), .Y (n_24764));
MX2X1 g57861(.A (n_24113), .B (key[38]), .S0 (n_1890), .Y (n_24763));
INVX1 g57864(.A (n_24760), .Y (n_24761));
INVX1 g57866(.A (n_24758), .Y (n_24759));
MX2X1 g57871(.A (n_24105), .B (key[45]), .S0 (n_619), .Y (n_24757));
NAND2X1 g56728(.A (n_24611), .B (n_24132), .Y (n_24756));
DFFX1 u0_w_reg[0][28] (.CK (clk), .D (n_24375), .Q (w0[28] ), .QN());
DFFX1 u0_w_reg[0][14] (.CK (clk), .D (n_24350), .Q (w0[14] ), .QN());
NAND2X1 g57932(.A (n_23221), .B (n_24754), .Y (n_24755));
NAND2X1 g57933(.A (n_23535), .B (n_24752), .Y (n_24753));
NAND2X1 g57934(.A (n_23534), .B (n_28332), .Y (n_24751));
NAND2X1 g57936(.A (n_23878), .B (n_27487), .Y (n_24750));
NAND2X1 g57941(.A (n_27487), .B (n_22840), .Y (n_24749));
NAND2X1 g57944(.A (n_24754), .B (n_23811), .Y (n_24747));
NAND2X1 g57945(.A (n_24752), .B (n_23099), .Y (n_24746));
NAND2X1 g57947(.A (n_28332), .B (n_22594), .Y (n_24745));
MX2X1 g56734(.A (n_23735), .B (n_24378), .S0 (n_23704), .Y (n_24743));
INVX1 g57966(.A (n_24741), .Y (n_24742));
XOR2X1 g57976(.A (u0_rcon_1056), .B (n_24058), .Y (n_24740));
XOR2X1 g57977(.A (n_1560), .B (n_24736), .Y (n_24739));
XOR2X1 g57978(.A (n_20309), .B (n_24053), .Y (n_24738));
XOR2X1 g57979(.A (n_18661), .B (n_24736), .Y (n_24737));
MX2X1 g57986(.A (n_24070), .B (n_24069), .S0 (n_24219), .Y (n_24735));
NAND2X1 g57990(.A (n_24381), .B (n_24153), .Y (n_24890));
MX2X1 g57992(.A (n_23737), .B (n_23736), .S0 (n_24068), .Y (n_24888));
NAND2X1 g57994(.A (n_24380), .B (n_24152), .Y (n_24886));
DFFX1 u0_w_reg[2][1] (.CK (clk), .D (n_24384), .Q (w2[1] ), .QN ());
NAND2X1 g58008(.A (n_24151), .B (n_24379), .Y (n_24883));
MX2X1 g58012(.A (key[107]), .B (n_24049), .S0 (n_360), .Y (n_24734));
MX2X1 g58013(.A (key[75]), .B (n_24046), .S0 (n_229), .Y (n_24733));
MX2X1 g58015(.A (key[11]), .B (n_24043), .S0 (n_360), .Y (n_24731));
DFFX1 u0_w_reg[2][7] (.CK (clk), .D (n_24415), .Q (w2[7] ), .QN ());
XOR2X1 g58037(.A (n_1556), .B (n_24044), .Y (n_24730));
XOR2X1 g58040(.A (n_24215), .B (n_23718), .Y (n_24729));
INVX1 g58042(.A (n_24727), .Y (n_24728));
INVX1 g58055(.A (n_24725), .Y (n_24726));
MX2X1 g58057(.A (n_24002), .B (key[49]), .S0 (n_25126), .Y (n_24724));
MX2X1 g58059(.A (n_24001), .B (key[41]), .S0 (n_619), .Y (n_24723));
MX2X1 g58061(.A (n_23484), .B (n_23485), .S0 (n_24005), .Y (n_24877));
XOR2X1 g58063(.A (n_23196), .B (n_24012), .Y (n_25045));
XOR2X1 g58064(.A (n_23683), .B (n_24009), .Y (n_25002));
XOR2X1 g58065(.A (n_23989), .B (n_24006), .Y (n_24975));
NAND2X1 g58116(.A (n_24194), .B (n_24721), .Y (n_24722));
NAND2X1 g58121(.A (n_24280), .B (n_24428), .Y (n_24720));
NAND3X1 g58127(.A (n_24085), .B (n_24476), .C (n_24475), .Y(n_24719));
NAND3X1 g58128(.A (n_24358), .B (n_24466), .C (n_24465), .Y(n_24718));
NAND2X1 g58131(.A (n_24501), .B (n_24575), .Y (n_24717));
NAND2X1 g58138(.A (n_24714), .B (n_24613), .Y (n_24715));
NAND2X1 g58139(.A (n_24294), .B (n_24027), .Y (n_24713));
NAND2X1 g58142(.A (n_24497), .B (n_26948), .Y (n_24712));
NAND2X1 g58147(.A (n_24272), .B (n_26637), .Y (n_24711));
NAND2X1 g58149(.A (n_24271), .B (n_24491), .Y (n_24710));
NAND3X1 g58154(.A (n_24361), .B (n_24473), .C (n_24472), .Y(n_24709));
NAND3X1 g58160(.A (n_24308), .B (n_26778), .C (n_26779), .Y(n_24708));
NAND2X1 g58165(.A (n_24489), .B (n_23384), .Y (n_24707));
NAND2X1 g58168(.A (n_24409), .B (n_24066), .Y (n_24706));
NAND2X1 g58169(.A (n_24704), .B (n_24565), .Y (n_24705));
NAND2X1 g58179(.A (n_28273), .B (n_24702), .Y (n_24703));
NAND2X1 g58181(.A (n_24700), .B (n_24699), .Y (n_24701));
DFFX1 text_out_reg[21] (.CK (clk), .D (n_24253), .Q (text_out[21]),.QN ());
NAND2X1 g58185(.A (n_24853), .B (n_24840), .Y (n_24698));
NAND2X1 g58186(.A (n_24992), .B (n_24699), .Y (n_24697));
INVX1 g58198(.A (n_24695), .Y (n_24696));
MX2X1 g58201(.A (n_23638), .B (n_23639), .S0 (n_24211), .Y (n_24838));
INVX1 g57380(.A (n_24693), .Y (n_24694));
MX2X1 g57385(.A (n_23683), .B (n_23195), .S0 (n_24122), .Y (n_24692));
XOR2X1 g57394(.A (n_23770), .B (n_24071), .Y (n_24691));
NAND2X2 g58232(.A (n_24302), .B (n_24079), .Y (n_24835));
MX2X1 g58237(.A (n_23470), .B (n_23471), .S0 (n_24222), .Y (n_24690));
NAND2X1 g58239(.A (n_24311), .B (n_24309), .Y (n_25027));
MX2X1 g57399(.A (w1[5] ), .B (n_23777), .S0 (n_24108), .Y (n_24832));
NAND2X1 g58245(.A (n_24307), .B (n_24305), .Y (n_25058));
NAND2X1 g58247(.A (n_24304), .B (n_24080), .Y (n_24830));
INVX1 g58249(.A (n_24688), .Y (n_24689));
INVX1 g58251(.A (n_24686), .Y (n_24687));
INVX1 g57408(.A (n_24684), .Y (n_24685));
NAND2X1 g57413(.A (n_24682), .B (n_24681), .Y (n_24683));
MX2X1 g56768(.A (n_24174), .B (n_24173), .S0 (n_23602), .Y (n_24680));
MX2X1 g57421(.A (n_24051), .B (n_24052), .S0 (n_23748), .Y (n_24679));
INVX1 g57423(.A (n_24677), .Y (n_24678));
MX2X1 g57426(.A (n_22778), .B (n_245), .S0 (n_24065), .Y (n_24676));
INVX1 g56771(.A (n_24674), .Y (n_24675));
XOR2X1 g58293(.A (n_2417), .B (n_24231), .Y (n_24673));
MX2X1 g58311(.A (w0[2] ), .B (n_2434), .S0 (n_24208), .Y (n_24672));
NAND2X1 g58313(.A (n_24100), .B (n_24314), .Y (n_24821));
INVX1 g58314(.A (n_24670), .Y (n_24671));
MX2X1 g57455(.A (n_24056), .B (n_24055), .S0 (n_24224), .Y (n_24669));
INVX1 g56777(.A (n_24667), .Y (n_24668));
NAND2X1 g58329(.A (n_24093), .B (n_24312), .Y (n_24817));
XOR2X1 g58330(.A (n_497), .B (n_23963), .Y (n_24666));
INVX1 g57468(.A (n_24661), .Y (n_24662));
INVX1 g56779(.A (n_24659), .Y (n_24660));
MX2X1 g57470(.A (n_23231), .B (n_24223), .S0 (n_24054), .Y (n_24655));
INVX1 g56781(.A (n_24653), .Y (n_24654));
INVX1 g57472(.A (n_24651), .Y (n_24652));
INVX1 g57474(.A (n_24649), .Y (n_24650));
INVX1 g57476(.A (n_24647), .Y (n_24648));
NAND2X1 g58417(.A (n_23853), .B (n_24645), .Y (n_24646));
INVX1 g58429(.A (n_24643), .Y (n_24644));
NAND2X1 g58432(.A (n_24239), .B (n_23964), .Y (n_24815));
NAND2X1 g58436(.A (n_24233), .B (n_23959), .Y (n_24813));
INVX1 g57037(.A (n_24641), .Y (n_24642));
NAND2X1 g58461(.A (n_24240), .B (n_23968), .Y (n_24640));
INVX1 g58463(.A (n_26780), .Y (n_24639));
MX2X1 g57041(.A (w2[6] ), .B (n_2437), .S0 (n_24000), .Y (n_24638));
INVX1 g58478(.A (n_24636), .Y (n_24637));
MX2X1 g57043(.A (n_23989), .B (n_23198), .S0 (n_23992), .Y (n_24635));
NAND2X1 g58513(.A (n_23980), .B (n_24247), .Y (n_24809));
NAND2X2 g58520(.A (n_23978), .B (n_24245), .Y (n_24804));
INVX1 g58527(.A (n_24634), .Y (n_24987));
XOR2X1 g57052(.A (n_28286), .B (n_28285), .Y (n_24633));
XOR2X1 g58532(.A (w2[12] ), .B (n_23878), .Y (n_24632));
MX2X1 g57055(.A (n_194), .B (w2[5] ), .S0 (n_23958), .Y (n_24801));
INVX1 g58576(.A (n_24852), .Y (n_24631));
INVX1 g58584(.A (n_24856), .Y (n_24630));
INVX1 g58587(.A (n_24874), .Y (n_24629));
INVX1 g56691(.A (n_24627), .Y (n_24628));
INVX1 g57066(.A (n_24625), .Y (n_24626));
INVX1 g58593(.A (n_24871), .Y (n_24624));
INVX1 g58595(.A (n_24849), .Y (n_24623));
NAND2X2 g58598(.A (n_25631), .B (n_25632), .Y (n_25076));
XOR2X1 g56693(.A (n_6352), .B (n_24163), .Y (n_25026));
NAND2X1 g58629(.A (n_24249), .B (n_23996), .Y (n_25030));
MX2X1 g57080(.A (n_24185), .B (n_24186), .S0 (n_23899), .Y (n_24622));
NAND2X1 g58631(.A (n_24248), .B (n_23990), .Y (n_24973));
INVX1 g57081(.A (n_24620), .Y (n_24621));
MX2X1 g57083(.A (w2[2] ), .B (n_1960), .S0 (n_24198), .Y (n_24619));
INVX1 g58647(.A (n_24617), .Y (n_24618));
DFFX1 text_out_reg[120] (.CK (clk), .D (n_24277), .Q(text_out[120]), .QN ());
XOR2X1 g56698(.A (n_23056), .B (n_24154), .Y (n_25033));
NAND2X1 g58767(.A (n_23514), .B (n_24412), .Y (n_24616));
XOR2X1 g56699(.A (n_24157), .B (n_23824), .Y (n_25039));
MX2X1 g57112(.A (n_24189), .B (n_24188), .S0 (n_24226), .Y (n_24615));
DFFX1 text_out_reg[16] (.CK (clk), .D (n_24209), .Q (text_out[16]),.QN ());
XOR2X1 g57119(.A (n_23202), .B (n_23937), .Y (n_24795));
MX2X1 g57126(.A (n_22911), .B (n_23584), .S0 (n_23862), .Y (n_24791));
NAND2X1 g57131(.A (n_24218), .B (n_23922), .Y (n_24788));
NAND2X1 g57133(.A (n_24217), .B (n_23918), .Y (n_24786));
INVX1 g58885(.A (n_24613), .Y (n_24614));
NAND2X1 g57137(.A (n_24214), .B (n_23925), .Y (n_24782));
INVX1 g58896(.A (n_24611), .Y (n_24612));
MX2X1 g56707(.A (n_23615), .B (n_23616), .S0 (n_23794), .Y (n_24784));
INVX1 g58928(.A (n_24609), .Y (n_24610));
DFFX1 text_out_reg[5] (.CK (clk), .D (n_24159), .Q (text_out[5]),.QN ());
DFFX1 text_out_reg[37] (.CK (clk), .D (n_23999), .Q (text_out[37]),.QN ());
DFFX1 text_out_reg[35] (.CK (clk), .D (n_24207), .Q (text_out[35]),.QN ());
DFFX1 text_out_reg[69] (.CK (clk), .D (n_24124), .Q (text_out[69]),.QN ());
DFFX1 text_out_reg[67] (.CK (clk), .D (n_24073), .Q (text_out[67]),.QN ());
DFFX1 u0_w_reg[2][25] (.CK (clk), .D (n_24166), .Q (w2[25] ), .QN());
DFFX1 u0_w_reg[1][25] (.CK (clk), .D (n_24167), .Q (), .QN (w1[25]));
DFFX1 u0_w_reg[0][12] (.CK (clk), .D (n_24148), .Q (n_23290), .QN());
DFFX1 u0_w_reg[3][12] (.CK (clk), .D (n_24145), .Q (w3[12] ), .QN());
DFFX1 u0_w_reg[0][22] (.CK (clk), .D (n_24130), .Q (w0[22] ), .QN());
DFFX1 u0_w_reg[0][6] (.CK (clk), .D (n_24129), .Q (w0[6] ), .QN ());
DFFX1 u0_w_reg[1][22] (.CK (clk), .D (n_24128), .Q (n_2440), .QN ());
DFFX1 u0_w_reg[1][6] (.CK (clk), .D (n_24127), .Q (n_23257), .QN ());
DFFX1 u0_w_reg[3][22] (.CK (clk), .D (n_24126), .Q (w3[22] ), .QN());
DFFX1 u0_w_reg[3][6] (.CK (clk), .D (n_24125), .Q (w3[6] ), .QN ());
DFFX1 text_out_reg[56] (.CK (clk), .D (n_24034), .Q (text_out[56]),.QN ());
DFFX1 u0_w_reg[0][17] (.CK (clk), .D (n_24023), .Q (w0[17] ), .QN());
DFFX1 text_out_reg[88] (.CK (clk), .D (n_24033), .Q (text_out[88]),.QN ());
DFFX1 u0_w_reg[0][9] (.CK (clk), .D (n_24022), .Q (w0[9] ), .QN ());
DFFX1 u0_w_reg[1][17] (.CK (clk), .D (n_24021), .Q (w1[17] ), .QN());
DFFX1 text_out_reg[53] (.CK (clk), .D (n_24004), .Q (text_out[53]),.QN ());
DFFX1 u0_w_reg[1][9] (.CK (clk), .D (n_24019), .Q (w1[9] ), .QN ());
DFFX1 u0_w_reg[3][17] (.CK (clk), .D (n_24017), .Q (w3[17] ), .QN());
DFFX1 u0_w_reg[3][9] (.CK (clk), .D (n_24016), .Q (w3[9] ), .QN ());
DFFX1 text_out_reg[85] (.CK (clk), .D (n_24003), .Q (text_out[85]),.QN ());
DFFX1 text_out_reg[83] (.CK (clk), .D (n_24015), .Q (text_out[83]),.QN ());
DFFX1 text_out_reg[24] (.CK (clk), .D (n_24035), .Q (text_out[24]),.QN ());
DFFX1 text_out_reg[75] (.CK (clk), .D (n_24050), .Q (text_out[75]),.QN ());
DFFX1 text_out_reg[123] (.CK (clk), .D (n_24036), .Q(text_out[123]), .QN ());
DFFX1 text_out_reg[73] (.CK (clk), .D (n_24013), .Q (text_out[73]),.QN ());
DFFX1 text_out_reg[106] (.CK (clk), .D (n_24197), .Q(text_out[106]), .QN ());
XOR2X1 g58934(.A (n_424), .B (n_24607), .Y (n_24608));
DFFX1 text_out_reg[82] (.CK (clk), .D (n_24180), .Q (text_out[82]),.QN ());
DFFX1 text_out_reg[30] (.CK (clk), .D (n_24171), .Q (text_out[30]),.QN ());
DFFX1 text_out_reg[23] (.CK (clk), .D (n_24175), .Q (text_out[23]),.QN ());
DFFX1 text_out_reg[18] (.CK (clk), .D (n_24181), .Q (text_out[18]),.QN ());
DFFX1 text_out_reg[114] (.CK (clk), .D (n_24182), .Q(text_out[114]), .QN ());
DFFX1 text_out_reg[57] (.CK (clk), .D (n_24161), .Q (text_out[57]),.QN ());
DFFX1 text_out_reg[89] (.CK (clk), .D (n_24160), .Q (text_out[89]),.QN ());
XOR2X1 g58936(.A (w2[16] ), .B (n_24605), .Y (n_24606));
DFFX1 text_out_reg[60] (.CK (clk), .D (n_24158), .Q (text_out[60]),.QN ());
XOR2X1 g58937(.A (n_23605), .B (n_24603), .Y (n_24604));
XOR2X1 g58995(.A (n_23580), .B (n_23820), .Y (n_24602));
MX2X1 g57806(.A (n_23793), .B (key[122]), .S0 (n_24778), .Y(n_24601));
MX2X1 g57809(.A (n_23792), .B (key[90]), .S0 (n_24599), .Y (n_24600));
MX2X1 g57813(.A (n_23790), .B (key[58]), .S0 (n_1914), .Y (n_24598));
MX2X1 g57817(.A (n_23789), .B (key[26]), .S0 (n_24599), .Y (n_24597));
MX2X1 g57825(.A (u0_rcon_1058), .B (n_18549), .S0 (n_23779), .Y(n_24596));
MX2X1 g57826(.A (n_24392), .B (n_24390), .S0 (n_4482), .Y (n_24595));
MX2X1 g57827(.A (n_20307), .B (n_20308), .S0 (n_23780), .Y (n_24594));
NAND2X1 g56725(.A (n_23696), .B (n_24099), .Y (n_24593));
MX2X1 g57865(.A (n_23819), .B (n_24169), .S0 (n_23772), .Y (n_24760));
MX2X1 g57867(.A (n_23452), .B (n_23451), .S0 (n_23786), .Y (n_24758));
MX2X1 g57870(.A (w0[6] ), .B (n_243), .S0 (n_23785), .Y (n_24592));
XOR2X1 g59308(.A (w0[30] ), .B (n_23803), .Y (n_24591));
XOR2X1 g59330(.A (n_13083), .B (n_24269), .Y (n_24590));
XOR2X1 g57876(.A (n_2633), .B (n_23778), .Y (n_24589));
XOR2X1 g59335(.A (w2[14] ), .B (n_24283), .Y (n_24588));
INVX1 g56729(.A (n_24586), .Y (n_24587));
MX2X1 g56731(.A (n_23947), .B (n_23946), .S0 (n_23698), .Y (n_24585));
NAND2X1 g57930(.A (n_23819), .B (n_24582), .Y (n_24584));
NAND2X1 g57942(.A (n_24582), .B (n_22500), .Y (n_24583));
NAND2X1 g57967(.A (n_23796), .B (n_24150), .Y (n_24741));
XOR2X1 g56735(.A (n_23920), .B (n_23703), .Y (n_24581));
INVX1 g57974(.A (n_24579), .Y (n_24580));
DFFX1 u0_w_reg[1][12] (.CK (clk), .D (n_24147), .Q (w1[12] ), .QN());
MX2X1 g57981(.A (n_24577), .B (n_24576), .S0 (n_24575), .Y (n_24578));
MX2X1 g57982(.A (n_28117), .B (n_24573), .S0 (n_26948), .Y (n_24574));
MX2X1 g57983(.A (key[99]), .B (n_23731), .S0 (n_360), .Y (n_24571));
MX2X1 g57984(.A (key[67]), .B (n_23732), .S0 (n_360), .Y (n_24570));
MX2X1 g57985(.A (key[3]), .B (n_23728), .S0 (n_360), .Y (n_24568));
MX2X1 g58010(.A (n_24565), .B (n_24564), .S0 (n_24559), .Y (n_24566));
DFFX1 u0_w_reg[3][25] (.CK (clk), .D (n_24165), .Q (w3[25] ), .QN());
DFFX1 u0_w_reg[0][25] (.CK (clk), .D (n_24168), .Q (w0[25] ), .QN());
XOR2X1 g58036(.A (n_1666), .B (n_23729), .Y (n_24563));
MX2X1 g58043(.A (n_23266), .B (n_23267), .S0 (n_23713), .Y (n_24727));
MX2X1 g58056(.A (n_925), .B (n_234), .S0 (n_23700), .Y (n_24725));
NAND2X1 g58120(.A (n_23482), .B (n_24042), .Y (n_24562));
NAND2X1 g58122(.A (n_24279), .B (n_24427), .Y (n_24561));
NAND2X1 g58140(.A (n_24293), .B (n_24559), .Y (n_24560));
NAND2X1 g58167(.A (n_24408), .B (n_24067), .Y (n_24558));
NAND2X1 g58170(.A (n_24281), .B (n_23135), .Y (n_24557));
NAND2X1 g58175(.A (n_24998), .B (n_24896), .Y (n_24556));
NAND2X1 g58176(.A (n_24869), .B (n_24895), .Y (n_24555));
NAND2X1 g58177(.A (n_24865), .B (n_24553), .Y (n_24554));
NAND2X1 g58178(.A (n_24714), .B (n_24149), .Y (n_24552));
NAND2X1 g58187(.A (n_24990), .B (n_24899), .Y (n_24551));
NAND2X1 g58188(.A (n_24850), .B (n_24898), .Y (n_24550));
MX2X1 g58192(.A (n_23949), .B (key[36]), .S0 (n_24548), .Y (n_24549));
MX2X1 g58195(.A (key[92]), .B (n_23943), .S0 (n_360), .Y (n_24547));
MX2X1 g58197(.A (key[28]), .B (n_23942), .S0 (n_360), .Y (n_24545));
NAND2X1 g58199(.A (n_23752), .B (n_24076), .Y (n_24695));
INVX1 g58203(.A (n_24543), .Y (n_24544));
MX2X1 g57381(.A (n_22824), .B (n_23081), .S0 (n_23784), .Y (n_24693));
MX2X1 g57387(.A (n_23257), .B (n_141), .S0 (n_23783), .Y (n_24542));
NAND2X1 g58219(.A (n_24077), .B (n_23753), .Y (n_24541));
XOR2X1 g57388(.A (n_28266), .B (n_28265), .Y (n_25005));
MX2X1 g57390(.A (n_22781), .B (n_97), .S0 (n_23781), .Y (n_24540));
XOR2X1 g57396(.A (n_23351), .B (n_23773), .Y (n_24539));
NAND2X1 g58242(.A (n_24089), .B (n_24087), .Y (n_24907));
NAND2X1 g58243(.A (n_24084), .B (n_23756), .Y (n_24538));
NAND2X1 g58244(.A (n_23755), .B (n_24082), .Y (n_24807));
MX2X1 g58250(.A (n_24449), .B (n_24255), .S0 (n_23924), .Y (n_24688));
MX2X1 g58252(.A (n_24241), .B (n_22939), .S0 (n_23923), .Y (n_24686));
INVX1 g58253(.A (n_24536), .Y (n_24537));
MX2X1 g58255(.A (key[96]), .B (n_23915), .S0 (n_229), .Y (n_24535));
MX2X1 g58257(.A (key[112]), .B (n_23914), .S0 (n_360), .Y (n_24534));
MX2X1 g58260(.A (key[64]), .B (n_23912), .S0 (n_229), .Y (n_24533));
MX2X1 g57409(.A (n_23356), .B (n_23357), .S0 (n_23769), .Y (n_24684));
MX2X1 g58262(.A (key[80]), .B (n_23910), .S0 (n_360), .Y (n_24532));
NAND2X1 g57414(.A (n_23061), .B (n_24102), .Y (n_24530));
MX2X1 g58265(.A (key[0]), .B (n_23906), .S0 (n_229), .Y (n_24529));
MX2X1 g58267(.A (key[16]), .B (n_23905), .S0 (n_229), .Y (n_24528));
NAND2X1 g57417(.A (n_23716), .B (n_24111), .Y (n_24527));
XOR2X1 g58270(.A (n_925), .B (n_24345), .Y (n_24526));
MX2X1 g57422(.A (n_23722), .B (n_23723), .S0 (n_23746), .Y (n_24525));
NAND2X1 g57424(.A (n_24115), .B (n_23775), .Y (n_24677));
MX2X1 g58283(.A (n_23000), .B (n_24345), .S0 (n_23895), .Y (n_25031));
MX2X1 g56772(.A (n_23610), .B (n_23611), .S0 (n_23940), .Y (n_24674));
INVX1 g57436(.A (n_24523), .Y (n_24524));
INVX1 g58298(.A (n_24521), .Y (n_24522));
INVX1 g56773(.A (n_24519), .Y (n_24520));
NAND2X1 g57451(.A (n_23385), .B (n_24011), .Y (n_24518));
MX2X1 g56775(.A (n_24269), .B (n_24172), .S0 (n_23926), .Y (n_24517));
NAND2X1 g58315(.A (n_24095), .B (n_24097), .Y (n_24670));
MX2X1 g58321(.A (n_24316), .B (n_22863), .S0 (n_23897), .Y (n_25046));
XOR2X1 g58332(.A (n_684), .B (n_28899), .Y (n_24516));
XOR2X1 g58333(.A (n_645), .B (n_23653), .Y (n_24515));
INVX1 g58337(.A (n_27487), .Y (n_24514));
NAND2X1 g56778(.A (n_24090), .B (n_23754), .Y (n_24667));
NAND2X1 g56780(.A (n_24078), .B (n_23751), .Y (n_24659));
MX2X1 g57469(.A (n_22576), .B (n_23378), .S0 (n_23727), .Y (n_24661));
NAND2X1 g57473(.A (n_24092), .B (n_23760), .Y (n_24651));
MX2X1 g58357(.A (n_24283), .B (n_23316), .S0 (n_23890), .Y (n_24797));
NAND2X1 g56782(.A (n_24075), .B (n_23749), .Y (n_24653));
NAND2X1 g57475(.A (n_24091), .B (n_23759), .Y (n_24649));
XOR2X1 g58358(.A (n_24512), .B (n_23889), .Y (n_24919));
NAND2X1 g57477(.A (n_24088), .B (n_23757), .Y (n_24647));
NAND2X1 g58395(.A (n_28333), .B (n_23963), .Y (n_24511));
NAND2X1 g58418(.A (n_23854), .B (n_24509), .Y (n_24510));
NAND2X1 g58421(.A (n_23851), .B (n_24507), .Y (n_24508));
NAND2X1 g58423(.A (n_23849), .B (n_24505), .Y (n_24506));
NAND2X1 g58430(.A (n_23966), .B (n_23659), .Y (n_24643));
MX2X1 g57038(.A (n_22967), .B (n_23278), .S0 (n_23681), .Y (n_24641));
INVX1 g58469(.A (n_24501), .Y (n_24502));
INVX1 g58476(.A (n_24497), .Y (n_24498));
OAI21X1 g58479(.A0 (n_26751), .A1 (n_24496), .B0 (n_23971), .Y(n_24636));
INVX1 g58483(.A (n_26637), .Y (n_25822));
INVX1 g58488(.A (n_24491), .Y (n_24492));
INVX1 g58493(.A (n_24489), .Y (n_24490));
MX2X1 g57045(.A (w2[7] ), .B (n_1769), .S0 (n_23680), .Y (n_24488));
XOR2X1 g58508(.A (w2[11] ), .B (n_23861), .Y (n_24487));
INVX1 g58517(.A (n_24485), .Y (n_24486));
INVX1 g58521(.A (n_24702), .Y (n_24484));
INVX1 g58523(.A (n_24704), .Y (n_24483));
NAND2X2 g58528(.A (n_23977), .B (n_23673), .Y (n_24634));
XOR2X1 g58531(.A (n_23290), .B (n_23535), .Y (n_24482));
XOR2X1 g58533(.A (w1[12] ), .B (n_23534), .Y (n_24481));
NAND2X1 g56811(.A (n_23972), .B (n_23661), .Y (n_24480));
XOR2X1 g57056(.A (n_29403), .B (n_29402), .Y (n_24479));
INVX1 g58567(.A (n_28110), .Y (n_24478));
NAND2X2 g58577(.A (n_24476), .B (n_24475), .Y (n_24852));
AOI21X1 g58579(.A0 (n_24462), .A1 (n_26217), .B0 (n_23982), .Y(n_24841));
NAND2X2 g58585(.A (n_24473), .B (n_24472), .Y (n_24856));
MX2X1 g58586(.A (n_23983), .B (n_24607), .S0 (n_26751), .Y (n_24471));
NAND2X2 g58588(.A (n_23976), .B (n_23671), .Y (n_24874));
MX2X1 g58589(.A (n_23984), .B (n_24603), .S0 (n_26638), .Y (n_24469));
INVX1 g58590(.A (n_24721), .Y (n_24468));
MX2X1 g58592(.A (n_23981), .B (n_24605), .S0 (n_27706), .Y (n_24467));
MX2X1 g56692(.A (n_27085), .B (n_23636), .S0 (n_23804), .Y (n_24627));
NAND2X2 g58594(.A (n_23975), .B (n_23668), .Y (n_24871));
MX2X1 g57067(.A (n_23517), .B (n_23518), .S0 (n_23939), .Y (n_24625));
NAND2X2 g58596(.A (n_24466), .B (n_24465), .Y (n_24849));
MX2X1 g58597(.A (n_23817), .B (n_24436), .S0 (n_27061), .Y (n_24464));
NAND2X1 g57072(.A (n_28603), .B (n_23574), .Y (n_24463));
MX2X1 g58609(.A (n_24462), .B (n_23820), .S0 (n_23189), .Y (n_24912));
NAND2X1 g57075(.A (n_24040), .B (n_24228), .Y (n_24461));
MX2X1 g57077(.A (n_23859), .B (n_23860), .S0 (n_23903), .Y (n_24460));
NAND2X1 g58630(.A (n_23993), .B (n_23684), .Y (n_24880));
NAND2X1 g58632(.A (n_23987), .B (n_23986), .Y (n_25034));
XOR2X1 g58634(.A (w0[13] ), .B (n_23507), .Y (n_24459));
XOR2X1 g58635(.A (n_24366), .B (n_23871), .Y (n_24458));
NAND2X1 g57082(.A (n_23650), .B (n_23960), .Y (n_24620));
INVX1 g58642(.A (n_24456), .Y (n_24457));
MX2X1 g56695(.A (n_1142), .B (n_2760), .S0 (n_23810), .Y (n_24455));
NAND2X1 g58648(.A (n_23690), .B (n_23998), .Y (n_24617));
INVX1 g58649(.A (n_24453), .Y (n_24454));
MX2X1 g58652(.A (n_23560), .B (n_23147), .S0 (n_26654), .Y (n_24452));
MX2X1 g56697(.A (n_23985), .B (n_23213), .S0 (n_23806), .Y (n_24451));
NAND2X1 g58768(.A (n_24449), .B (n_24444), .Y (n_24450));
NAND2X1 g58769(.A (n_22939), .B (n_24177), .Y (n_24448));
NAND2X1 g57108(.A (n_23891), .B (n_24008), .Y (n_24447));
NAND2X1 g58798(.A (n_22895), .B (n_24176), .Y (n_24446));
NAND2X1 g58801(.A (n_24444), .B (n_23955), .Y (n_24445));
INVX1 g58819(.A (n_24442), .Y (n_24443));
INVX1 g58821(.A (n_24440), .Y (n_24441));
INVX1 g58823(.A (n_24438), .Y (n_24439));
DFFX1 text_out_reg[41] (.CK (clk), .D (n_23695), .Q (text_out[41]),.QN ());
XOR2X1 g57129(.A (w2[0] ), .B (n_23541), .Y (n_24437));
OAI21X1 g58886(.A0 (n_24436), .A1 (n_24285), .B0 (n_23882), .Y(n_24613));
OAI21X1 g58895(.A0 (n_24273), .A1 (n_26218), .B0 (n_23880), .Y(n_24435));
AOI21X1 g58897(.A0 (n_27946), .A1 (n_26104), .B0 (n_23879), .Y(n_24611));
MX2X1 g57138(.A (n_23887), .B (n_23145), .S0 (n_23512), .Y (n_24798));
XOR2X1 g58910(.A (n_22881), .B (n_23452), .Y (n_24433));
INVX1 g58911(.A (n_24509), .Y (n_24645));
AOI21X1 g58924(.A0 (n_23883), .A1 (n_26104), .B0 (n_23884), .Y(n_24430));
DFFX1 text_out_reg[1] (.CK (clk), .D (n_23701), .Q (text_out[1]),.QN ());
DFFX1 text_out_reg[7] (.CK (clk), .D (n_23904), .Q (text_out[7]),.QN ());
DFFX1 text_out_reg[38] (.CK (clk), .D (n_23679), .Q (text_out[38]),.QN ());
DFFX1 text_out_reg[36] (.CK (clk), .D (n_23649), .Q (text_out[36]),.QN ());
DFFX1 text_out_reg[33] (.CK (clk), .D (n_23893), .Q (text_out[33]),.QN ());
DFFX1 text_out_reg[39] (.CK (clk), .D (n_23858), .Q (text_out[39]),.QN ());
INVX1 g58925(.A (n_24427), .Y (n_24428));
DFFX1 text_out_reg[68] (.CK (clk), .D (n_23774), .Q (text_out[68]),.QN ());
DFFX1 text_out_reg[70] (.CK (clk), .D (n_23782), .Q (text_out[70]),.QN ());
DFFX1 text_out_reg[71] (.CK (clk), .D (n_23724), .Q (text_out[71]),.QN ());
NAND2X2 g58929(.A (n_23886), .B (n_23555), .Y (n_24609));
DFFX1 text_out_reg[50] (.CK (clk), .D (n_23852), .Q (text_out[50]),.QN ());
DFFX1 text_out_reg[59] (.CK (clk), .D (n_23710), .Q (text_out[59]),.QN ());
DFFX1 text_out_reg[91] (.CK (clk), .D (n_23706), .Q (text_out[91]),.QN ());
DFFX1 text_out_reg[40] (.CK (clk), .D (n_23711), .Q (text_out[40]),.QN ());
DFFX1 text_out_reg[72] (.CK (clk), .D (n_23707), .Q (text_out[72]),.QN ());
DFFX1 u0_w_reg[0][4] (.CK (clk), .D (n_23952), .Q (w0[4] ), .QN ());
DFFX1 u0_w_reg[1][4] (.CK (clk), .D (n_23951), .Q (w1[4] ), .QN ());
DFFX1 u0_w_reg[3][4] (.CK (clk), .D (n_23950), .Q (w3[4] ), .QN ());
DFFX1 text_out_reg[9] (.CK (clk), .D (n_23948), .Q (text_out[9]),.QN ());
DFFX1 text_out_reg[31] (.CK (clk), .D (n_23894), .Q (text_out[31]),.QN ());
DFFX1 text_out_reg[102] (.CK (clk), .D (n_23901), .Q(text_out[102]), .QN ());
DFFX1 text_out_reg[55] (.CK (clk), .D (n_23840), .Q (text_out[55]),.QN ());
DFFX1 text_out_reg[54] (.CK (clk), .D (n_23827), .Q (text_out[54]),.QN ());
DFFX1 text_out_reg[90] (.CK (clk), .D (n_23839), .Q (text_out[90]),.QN ());
DFFX1 text_out_reg[119] (.CK (clk), .D (n_23842), .Q(text_out[119]), .QN ());
DFFX1 text_out_reg[22] (.CK (clk), .D (n_23828), .Q (text_out[22]),.QN ());
DFFX1 text_out_reg[103] (.CK (clk), .D (n_23838), .Q(text_out[103]), .QN ());
DFFX1 text_out_reg[15] (.CK (clk), .D (n_23841), .Q (text_out[15]),.QN ());
DFFX1 text_out_reg[14] (.CK (clk), .D (n_23829), .Q (text_out[14]),.QN ());
DFFX1 text_out_reg[92] (.CK (clk), .D (n_23797), .Q (text_out[92]),.QN ());
DFFX1 text_out_reg[116] (.CK (clk), .D (n_23809), .Q(text_out[116]), .QN ());
DFFX1 text_out_reg[66] (.CK (clk), .D (n_23734), .Q (text_out[66]),.QN ());
NAND2X1 g57164(.A (n_23885), .B (n_23550), .Y (n_24426));
OAI21X1 g58993(.A0 (n_23556), .A1 (n_24462), .B0 (n_23557), .Y(n_24425));
XOR2X1 g58998(.A (n_23184), .B (n_28821), .Y (n_24424));
XOR2X1 g58999(.A (w2[15] ), .B (n_23145), .Y (n_24423));
XOR2X1 g59002(.A (n_23047), .B (n_24223), .Y (n_24422));
XOR2X1 g59003(.A (w1[15] ), .B (n_23144), .Y (n_24421));
INVX1 g59020(.A (n_24419), .Y (n_24420));
NAND2X1 g59066(.A (n_23863), .B (n_23663), .Y (n_24418));
NAND2X1 g59068(.A (n_23865), .B (n_22442), .Y (n_24417));
NAND2X1 g59070(.A (n_23867), .B (n_26218), .Y (n_24416));
MX2X1 g57830(.A (n_23411), .B (key[39]), .S0 (n_24915), .Y (n_24415));
INVX1 g59264(.A (n_24413), .Y (n_24414));
INVX1 g59268(.A (n_24444), .Y (n_24412));
MX2X1 g57857(.A (n_23396), .B (key[50]), .S0 (n_24548), .Y (n_24411));
MX2X1 g57858(.A (n_23395), .B (key[34]), .S0 (n_24548), .Y (n_24410));
INVX1 g59287(.A (n_24408), .Y (n_24409));
NAND2X1 g56724(.A (n_23697), .B (n_24098), .Y (n_24407));
INVX1 g59289(.A (n_24405), .Y (n_24406));
XOR2X1 g59310(.A (w2[30] ), .B (n_23435), .Y (n_24404));
XOR2X1 g59311(.A (n_2587), .B (n_23432), .Y (n_24403));
NAND2X1 g57249(.A (n_26534), .B (n_23181), .Y (n_24402));
XOR2X1 g59331(.A (n_23599), .B (n_24316), .Y (n_24401));
XOR2X1 g59337(.A (w1[14] ), .B (n_24315), .Y (n_24400));
NAND2X1 g59343(.A (n_23469), .B (n_23822), .Y (n_25536));
MX2X1 g56730(.A (n_23633), .B (n_23634), .S0 (n_23338), .Y (n_24586));
INVX1 g59353(.A (n_24397), .Y (n_24398));
NAND2X1 g57931(.A (n_24394), .B (n_24169), .Y (n_24396));
NAND2X1 g57943(.A (n_24394), .B (n_22593), .Y (n_24395));
NAND2X1 g57949(.A (n_24392), .B (n_15851), .Y (n_24393));
NAND2X1 g57950(.A (n_24390), .B (n_15850), .Y (n_24391));
MX2X1 g57975(.A (n_23481), .B (n_23480), .S0 (n_23393), .Y (n_24579));
MX2X1 g57980(.A (n_23380), .B (key[55]), .S0 (n_1890), .Y (n_24387));
XOR2X1 g59596(.A (w0[25] ), .B (n_23107), .Y (n_24386));
DFFX1 text_out_reg[11] (.CK (clk), .D (n_23725), .Q (text_out[11]),.QN ());
DFFX1 text_out_reg[34] (.CK (clk), .D (n_23873), .Q (text_out[34]),.QN ());
XOR2X1 g56743(.A (n_1142), .B (n_24155), .Y (n_24385));
MX2X1 g58058(.A (n_23336), .B (key[33]), .S0 (ld), .Y (n_24384));
XOR2X1 g59837(.A (w0[28] ), .B (n_23099), .Y (n_24383));
NAND2X1 g58119(.A (n_23483), .B (n_24041), .Y (n_24382));
XOR2X1 g56747(.A (n_23358), .B (n_23593), .Y (n_25057));
NAND2X1 g58161(.A (n_23930), .B (n_23745), .Y (n_24381));
NAND2X1 g58163(.A (n_23928), .B (n_23743), .Y (n_24380));
NAND2X1 g58174(.A (n_24378), .B (n_28117), .Y (n_24379));
MX2X1 g58191(.A (n_23635), .B (key[52]), .S0 (n_24778), .Y (n_24376));
DFFX1 text_out_reg[27] (.CK (clk), .D (n_23712), .Q (text_out[27]),.QN ());
MX2X1 g58194(.A (n_23631), .B (key[124]), .S0 (n_619), .Y (n_24375));
MX2X1 g58196(.A (n_23627), .B (key[60]), .S0 (n_25126), .Y (n_24374));
MX2X1 g58204(.A (n_24236), .B (n_22895), .S0 (n_23618), .Y (n_24543));
XOR2X1 g58207(.A (u0_rcon_1059), .B (n_23597), .Y (n_24373));
XOR2X1 g58209(.A (n_2509), .B (n_23630), .Y (n_24372));
XOR2X1 g58213(.A (n_1606), .B (n_29188), .Y (n_24371));
XOR2X1 g57386(.A (n_23073), .B (n_23401), .Y (n_24879));
XOR2X1 g58217(.A (n_17375), .B (n_23592), .Y (n_24370));
XOR2X1 g58221(.A (n_13951), .B (n_29187), .Y (n_24369));
MX2X1 g57389(.A (n_24315), .B (n_23093), .S0 (n_23403), .Y (n_25003));
XOR2X1 g58223(.A (n_24366), .B (n_24364), .Y (n_24367));
XOR2X1 g58225(.A (n_2405), .B (n_24364), .Y (n_24365));
XOR2X1 g58228(.A (n_10653), .B (n_24364), .Y (n_24363));
MX2X1 g58238(.A (n_23434), .B (n_23435), .S0 (n_24361), .Y (n_24362));
XOR2X1 g56763(.A (n_3955), .B (n_23637), .Y (n_24360));
MX2X1 g58248(.A (n_23431), .B (n_23432), .S0 (n_24358), .Y (n_24359));
MX2X1 g58254(.A (n_23967), .B (n_22744), .S0 (n_23619), .Y (n_24536));
MX2X1 g58256(.A (key[106]), .B (n_23613), .S0 (n_229), .Y (n_24357));
MX2X1 g58261(.A (key[74]), .B (n_23609), .S0 (n_360), .Y (n_24355));
NAND2X1 g57415(.A (n_23062), .B (n_24101), .Y (n_24353));
MX2X1 g58266(.A (key[10]), .B (n_23604), .S0 (n_229), .Y (n_24352));
NAND2X1 g57418(.A (n_23715), .B (n_24110), .Y (n_24351));
MX2X1 g58271(.A (key[110]), .B (n_23600), .S0 (n_360), .Y (n_24350));
MX2X1 g58274(.A (key[78]), .B (n_23590), .S0 (n_360), .Y (n_24349));
MX2X1 g56769(.A (n_22621), .B (n_27946), .S0 (n_23598), .Y (n_24920));
MX2X1 g58277(.A (key[14]), .B (n_23591), .S0 (n_360), .Y (n_24347));
OAI21X1 g58280(.A0 (n_24345), .A1 (n_1019), .B0 (n_23766), .Y(n_24346));
OAI21X1 g58281(.A0 (n_24345), .A1 (n_23763), .B0 (n_23765), .Y(n_24344));
MX2X1 g58285(.A (key[109]), .B (n_23583), .S0 (n_360), .Y (n_24343));
MX2X1 g58286(.A (key[111]), .B (n_23581), .S0 (n_360), .Y (n_24342));
MX2X1 g58288(.A (key[104]), .B (n_23579), .S0 (n_229), .Y (n_24341));
MX2X1 g58289(.A (key[77]), .B (n_23577), .S0 (n_229), .Y (n_24340));
MX2X1 g58290(.A (key[79]), .B (n_23573), .S0 (n_229), .Y (n_24338));
MX2X1 g58292(.A (key[72]), .B (n_23571), .S0 (n_229), .Y (n_24337));
MX2X1 g58294(.A (key[13]), .B (n_23566), .S0 (n_229), .Y (n_24335));
MX2X1 g58295(.A (key[15]), .B (n_23565), .S0 (n_360), .Y (n_24333));
MX2X1 g57437(.A (n_23091), .B (n_22828), .S0 (n_23361), .Y (n_24523));
MX2X1 g58297(.A (key[8]), .B (n_23564), .S0 (n_229), .Y (n_24332));
NAND2X1 g58299(.A (n_23762), .B (n_23761), .Y (n_24521));
MX2X1 g56774(.A (n_28350), .B (n_28349), .S0 (n_23620), .Y (n_24519));
XOR2X1 g58306(.A (n_1833), .B (n_23607), .Y (n_24331));
XOR2X1 g58307(.A (n_606), .B (n_23603), .Y (n_24330));
XOR2X1 g58308(.A (n_2650), .B (n_23606), .Y (n_24329));
NAND2X1 g57452(.A (n_23386), .B (n_24010), .Y (n_24328));
XOR2X1 g58316(.A (n_1675), .B (n_23595), .Y (n_24327));
MX2X1 g58320(.A (n_22847), .B (n_23445), .S0 (n_24319), .Y (n_24326));
XOR2X1 g58331(.A (n_2959), .B (n_23308), .Y (n_24325));
XOR2X1 g56776(.A (n_22418), .B (n_29349), .Y (n_24324));
XOR2X1 g58341(.A (n_2010), .B (n_23569), .Y (n_24323));
XOR2X1 g58342(.A (n_1297), .B (n_23568), .Y (n_24322));
INVX1 g58343(.A (n_24582), .Y (n_24321));
MX2X1 g58353(.A (n_23531), .B (n_26510), .S0 (n_24319), .Y (n_24752));
XOR2X1 g57471(.A (n_1958), .B (n_27815), .Y (n_24318));
MX2X1 g58354(.A (n_26510), .B (n_23531), .S0 (n_24319), .Y (n_24754));
MX2X1 g58355(.A (n_24316), .B (n_22863), .S0 (n_23563), .Y (n_24911));
MX2X1 g58356(.A (n_24315), .B (n_23093), .S0 (n_23562), .Y (n_24681));
NAND2X1 g58391(.A (n_28776), .B (n_23656), .Y (n_24314));
NAND2X1 g58394(.A (n_23994), .B (n_23962), .Y (n_24313));
MX2X1 g57481(.A (n_23888), .B (n_23144), .S0 (n_23362), .Y (n_24682));
NAND2X1 g58396(.A (n_23475), .B (n_23653), .Y (n_24312));
NAND2X1 g58405(.A (n_23693), .B (n_24310), .Y (n_24311));
NAND2X1 g58406(.A (n_23120), .B (n_24308), .Y (n_24309));
NAND2X1 g58413(.A (n_24306), .B (n_24310), .Y (n_24307));
NAND2X1 g58414(.A (n_24512), .B (n_24308), .Y (n_24305));
NAND2X1 g58415(.A (n_23803), .B (n_24303), .Y (n_24304));
NAND2X1 g58419(.A (n_23502), .B (n_24301), .Y (n_24302));
NAND2X1 g58422(.A (n_23850), .B (n_24213), .Y (n_24300));
NAND2X1 g58424(.A (n_23848), .B (n_24212), .Y (n_24299));
NAND2X1 g57507(.A (n_23740), .B (n_23377), .Y (n_24298));
MX2X1 g58449(.A (n_23811), .B (n_23446), .S0 (n_24265), .Y (n_24297));
DFFX1 text_out_reg[2] (.CK (clk), .D (n_23938), .Q (text_out[2]),.QN ());
MX2X1 g58455(.A (n_22596), .B (n_22595), .S0 (n_24260), .Y (n_24296));
MX2X1 g58458(.A (n_22500), .B (n_28118), .S0 (n_24263), .Y (n_24295));
MX2X1 g58470(.A (n_24062), .B (n_23193), .S0 (n_24260), .Y (n_24501));
INVX1 g58474(.A (n_24293), .Y (n_24294));
MX2X1 g58477(.A (n_23499), .B (n_23498), .S0 (n_24263), .Y (n_24497));
OAI21X1 g58489(.A0 (n_27706), .A1 (n_24289), .B0 (n_23664), .Y(n_24491));
INVX1 g58491(.A (n_24287), .Y (n_24288));
OAI21X1 g58494(.A0 (n_27061), .A1 (n_24285), .B0 (n_23662), .Y(n_24489));
XOR2X1 g57044(.A (n_25563), .B (n_23269), .Y (n_24972));
NAND2X1 g57539(.A (n_23708), .B (n_23343), .Y (n_24284));
MX2X1 g57047(.A (n_24283), .B (n_23316), .S0 (n_23324), .Y (n_24976));
MX2X1 g58511(.A (n_23674), .B (n_25889), .S0 (n_24265), .Y (n_25518));
NAND2X1 g58518(.A (n_23678), .B (n_23677), .Y (n_24485));
NAND2X2 g58522(.A (n_23675), .B (n_23322), .Y (n_24702));
INVX2 g58524(.A (n_24281), .Y (n_24704));
INVX1 g58537(.A (n_24279), .Y (n_24280));
XOR2X1 g58550(.A (w0[8] ), .B (n_26217), .Y (n_24278));
XOR2X1 g58551(.A (n_22981), .B (n_26751), .Y (n_24277));
MX2X1 g58565(.A (n_24275), .B (n_24276), .S0 (n_26751), .Y (n_24853));
MX2X1 g58566(.A (n_24276), .B (n_24275), .S0 (n_26751), .Y (n_24992));
MX2X1 g58578(.A (n_24273), .B (n_24196), .S0 (n_26217), .Y (n_24700));
INVX1 g58580(.A (n_24272), .Y (n_24860));
INVX1 g58582(.A (n_24271), .Y (n_24858));
OAI21X1 g56817(.A0 (n_28350), .A1 (n_24269), .B0 (n_23686), .Y(n_24270));
NAND2X2 g58591(.A (n_23670), .B (n_23319), .Y (n_24721));
NAND2X1 g57073(.A (n_23575), .B (n_24220), .Y (n_24268));
XOR2X1 g58611(.A (n_24266), .B (n_24265), .Y (n_24267));
XOR2X1 g58612(.A (n_18792), .B (n_24263), .Y (n_24264));
NAND2X1 g57076(.A (n_24039), .B (n_24227), .Y (n_24262));
XOR2X1 g58613(.A (w2[19] ), .B (n_24260), .Y (n_24261));
INVX1 g58615(.A (n_24258), .Y (n_24259));
XOR2X1 g58617(.A (n_23169), .B (n_23514), .Y (n_24257));
OAI21X1 g58620(.A0 (n_24255), .A1 (n_24462), .B0 (n_23331), .Y(n_24256));
XOR2X1 g58636(.A (n_2239), .B (n_23527), .Y (n_24254));
XOR2X1 g58637(.A (n_6431), .B (n_23332), .Y (n_24253));
XOR2X1 g58638(.A (w2[13] ), .B (n_23198), .Y (n_24252));
XOR2X1 g58640(.A (n_764), .B (n_23195), .Y (n_24251));
NAND2X1 g58643(.A (n_23692), .B (n_23335), .Y (n_24456));
NAND2X1 g58650(.A (n_23689), .B (n_23334), .Y (n_24453));
NAND2X1 g58651(.A (n_23333), .B (n_23687), .Y (n_25800));
NAND2X1 g58692(.A (n_23507), .B (n_28336), .Y (n_24249));
NAND2X1 g58696(.A (n_23198), .B (n_28776), .Y (n_24248));
NAND2X1 g58723(.A (n_23667), .B (n_26534), .Y (n_24247));
NAND2X1 g58727(.A (n_24243), .B (n_28325), .Y (n_24245));
XOR2X1 g57095(.A (n_23010), .B (n_23510), .Y (n_24806));
NAND2X1 g58741(.A (n_24243), .B (n_22929), .Y (n_25631));
NAND2X1 g58770(.A (n_24241), .B (n_24232), .Y (n_24242));
NAND2X1 g58771(.A (n_22744), .B (n_23845), .Y (n_24240));
NAND2X1 g58775(.A (n_24235), .B (n_23956), .Y (n_24239));
NAND2X1 g57109(.A (n_23892), .B (n_24007), .Y (n_24238));
NAND2X1 g58799(.A (n_24236), .B (n_24235), .Y (n_24237));
NAND3X1 g58800(.A (n_23107), .B (n_24179), .C (n_24178), .Y(n_24234));
NAND2X1 g58802(.A (n_24232), .B (n_23111), .Y (n_24233));
CLKBUFX1 g58804(.A (n_24231), .Y (n_24824));
DFFX1 text_out_reg[28] (.CK (clk), .D (n_23798), .Q (text_out[28]),.QN ());
OAI21X1 g58820(.A0 (n_23867), .A1 (n_23955), .B0 (n_23868), .Y(n_24442));
OAI21X1 g58822(.A0 (n_23865), .A1 (n_23303), .B0 (n_23866), .Y(n_24440));
OAI21X1 g58824(.A0 (n_23863), .A1 (n_23305), .B0 (n_23864), .Y(n_24438));
INVX1 g58825(.A (n_24229), .Y (n_24230));
INVX1 g57116(.A (n_24227), .Y (n_24228));
DFFX1 text_out_reg[25] (.CK (clk), .D (n_23448), .Q (text_out[25]),.QN ());
DFFX1 u0_w_reg[3][7] (.CK (clk), .D (n_23412), .Q (w3[7] ), .QN ());
AOI22X1 g58864(.A0 (n_22674), .A1 (n_28822), .B0 (n_22644), .B1(n_28827), .Y (n_24226));
AOI22X1 g58865(.A0 (n_22798), .A1 (n_22906), .B0 (n_22868), .B1(n_24223), .Y (n_24224));
NAND2X1 g58866(.A (n_23533), .B (n_23532), .Y (n_24222));
INVX1 g57134(.A (n_24220), .Y (n_28603));
NAND2X1 g58890(.A (n_23539), .B (n_23222), .Y (n_24219));
NAND2X1 g57142(.A (n_23541), .B (n_2648), .Y (n_24218));
NAND2X2 g58912(.A (n_23554), .B (n_23227), .Y (n_24509));
NAND2X1 g57144(.A (n_23541), .B (n_1296), .Y (n_24217));
OAI21X1 g58917(.A0 (n_23552), .A1 (n_23551), .B0 (n_23553), .Y(n_24215));
NAND2X1 g57146(.A (n_23541), .B (n_1220), .Y (n_24214));
INVX1 g58919(.A (n_24213), .Y (n_24507));
DFFX1 text_out_reg[58] (.CK (clk), .D (n_23490), .Q (text_out[58]),.QN ());
INVX1 g58922(.A (n_24212), .Y (n_24505));
DFFX1 text_out_reg[122] (.CK (clk), .D (n_23493), .Q(text_out[122]), .QN ());
DFFX1 text_out_reg[3] (.CK (clk), .D (n_23345), .Q (text_out[3]),.QN ());
DFFX1 u0_w_reg[1][18] (.CK (clk), .D (n_23408), .Q (w1[18] ), .QN());
OAI21X1 g58926(.A0 (n_24210), .A1 (n_23547), .B0 (n_23548), .Y(n_24427));
DFFX1 text_out_reg[65] (.CK (clk), .D (n_23387), .Q (text_out[65]),.QN ());
DFFX1 u0_w_reg[1][7] (.CK (clk), .D (n_23414), .Q (n_22781), .QN ());
OAI21X1 g58927(.A0 (n_24210), .A1 (n_23545), .B0 (n_23546), .Y(n_24211));
DFFX1 u0_w_reg[0][2] (.CK (clk), .D (n_23409), .Q (w0[2] ), .QN ());
DFFX1 u0_w_reg[1][2] (.CK (clk), .D (n_23407), .Q (n_22778), .QN ());
DFFX1 u0_w_reg[3][18] (.CK (clk), .D (n_23406), .Q (n_267), .QN ());
DFFX1 u0_w_reg[3][2] (.CK (clk), .D (n_23405), .Q (w3[2] ), .QN ());
DFFX1 u0_w_reg[0][23] (.CK (clk), .D (n_23392), .Q (n_22717), .QN());
DFFX1 u0_w_reg[3][23] (.CK (clk), .D (n_23390), .Q (w3[23] ), .QN());
DFFX1 text_out_reg[107] (.CK (clk), .D (n_23364), .Q(text_out[107]), .QN ());
DFFX1 u0_w_reg[0][20] (.CK (clk), .D (n_23646), .Q (n_22653), .QN());
DFFX1 u0_w_reg[1][20] (.CK (clk), .D (n_23644), .Q (w1[20] ), .QN());
DFFX1 u0_w_reg[3][20] (.CK (clk), .D (n_23643), .Q (w3[20] ), .QN());
DFFX1 text_out_reg[97] (.CK (clk), .D (n_23614), .Q (text_out[97]),.QN ());
DFFX1 text_out_reg[63] (.CK (clk), .D (n_23586), .Q (text_out[63]),.QN ());
DFFX1 text_out_reg[96] (.CK (clk), .D (n_23601), .Q (text_out[96]),.QN ());
DFFX1 text_out_reg[113] (.CK (clk), .D (n_23621), .Q(text_out[113]), .QN ());
DFFX1 text_out_reg[127] (.CK (clk), .D (n_23587), .Q(text_out[127]), .QN ());
DFFX1 text_out_reg[118] (.CK (clk), .D (n_23474), .Q(text_out[118]), .QN ());
DFFX1 text_out_reg[26] (.CK (clk), .D (n_23491), .Q (text_out[26]),.QN ());
DFFX1 text_out_reg[98] (.CK (clk), .D (n_23472), .Q (text_out[98]),.QN ());
DFFX1 text_out_reg[52] (.CK (clk), .D (n_23441), .Q (text_out[52]),.QN ());
DFFX1 text_out_reg[84] (.CK (clk), .D (n_23440), .Q (text_out[84]),.QN ());
XOR2X1 g58935(.A (n_880), .B (n_24436), .Y (n_24209));
NAND2X1 g58967(.A (n_23558), .B (n_23228), .Y (n_24208));
XOR2X1 g57163(.A (w2[3] ), .B (n_23174), .Y (n_24207));
INVX1 g58968(.A (n_24205), .Y (n_24206));
MX2X1 g57165(.A (n_1842), .B (w2[19] ), .S0 (n_23174), .Y (n_24204));
AOI21X1 g57167(.A0 (n_23543), .A1 (n_23902), .B0 (n_23544), .Y(n_28285));
INVX1 g58986(.A (n_24201), .Y (n_24202));
INVX1 g58989(.A (n_24199), .Y (n_24200));
OAI21X1 g57168(.A0 (n_23584), .A1 (n_28820), .B0 (n_23559), .Y(n_24198));
XOR2X1 g58994(.A (w0[10] ), .B (n_23560), .Y (n_24197));
AOI21X1 g59021(.A0 (n_24196), .A1 (n_23560), .B0 (n_23561), .Y(n_24419));
INVX1 g59022(.A (n_24194), .Y (n_24195));
INVX1 g59024(.A (n_24192), .Y (n_24193));
INVX1 g57205(.A (n_24188), .Y (n_24189));
OAI21X1 g57207(.A0 (n_23872), .A1 (n_23494), .B0 (n_23495), .Y(n_24187));
INVX1 g57209(.A (n_24185), .Y (n_24186));
DFFX1 text_out_reg[95] (.CK (clk), .D (n_23585), .Q (text_out[95]),.QN ());
INVX1 g57221(.A (n_24183), .Y (n_24184));
XOR2X1 g59254(.A (w0[18] ), .B (n_23455), .Y (n_24182));
XOR2X1 g59257(.A (n_19310), .B (n_28799), .Y (n_24181));
XOR2X1 g59259(.A (w1[18] ), .B (n_22868), .Y (n_24180));
AOI22X1 g59265(.A0 (n_28800), .A1 (n_24172), .B0 (n_28798), .B1(n_23117), .Y (n_24413));
NAND2X2 g59269(.A (n_24179), .B (n_24178), .Y (n_24444));
INVX1 g59270(.A (n_24232), .Y (n_24177));
INVX1 g59274(.A (n_24235), .Y (n_24176));
XOR2X1 g59278(.A (n_3868), .B (n_23131), .Y (n_24175));
INVX1 g59285(.A (n_24173), .Y (n_24174));
OAI21X1 g59288(.A0 (n_23457), .A1 (n_23881), .B0 (n_23458), .Y(n_24408));
OAI21X1 g59290(.A0 (n_24172), .A1 (n_27946), .B0 (n_23456), .Y(n_24405));
XOR2X1 g59309(.A (n_5236), .B (n_23121), .Y (n_24171));
NAND2X1 g57250(.A (n_23979), .B (n_23869), .Y (n_24170));
DFFX1 u0_w_reg[0][7] (.CK (clk), .D (n_23415), .Q (w0[7] ), .QN ());
NAND2X1 g59354(.A (n_23159), .B (n_23468), .Y (n_24397));
DFFX1 u0_w_reg[0][18] (.CK (clk), .D (n_23410), .Q (w0[18] ), .QN());
MX2X1 g57968(.A (n_23072), .B (key[121]), .S0 (n_24915), .Y(n_24168));
MX2X1 g57969(.A (key[89]), .B (n_23071), .S0 (n_360), .Y (n_24167));
MX2X1 g57970(.A (n_23070), .B (key[57]), .S0 (n_1890), .Y (n_24166));
MX2X1 g57971(.A (key[25]), .B (n_23069), .S0 (n_360), .Y (n_24165));
OAI21X1 g56736(.A0 (n_24155), .A1 (n_27946), .B0 (n_23417), .Y(n_24163));
XOR2X1 g59598(.A (w2[25] ), .B (n_23115), .Y (n_24161));
XOR2X1 g59599(.A (n_153), .B (n_22842), .Y (n_24160));
XOR2X1 g56739(.A (n_4750), .B (n_23056), .Y (n_24159));
XOR2X1 g59839(.A (w2[28] ), .B (n_22840), .Y (n_24158));
OAI21X1 g56744(.A0 (n_23423), .A1 (n_3014), .B0 (n_23425), .Y(n_24157));
OAI21X1 g56745(.A0 (n_24155), .A1 (n_23422), .B0 (n_23424), .Y(n_24156));
OAI21X1 g56746(.A0 (n_24155), .A1 (n_23418), .B0 (n_23419), .Y(n_24154));
NAND2X1 g58162(.A (n_23929), .B (n_23744), .Y (n_24153));
NAND2X1 g58164(.A (n_23927), .B (n_23742), .Y (n_24152));
NAND2X1 g58173(.A (n_23735), .B (n_24573), .Y (n_24151));
NAND2X1 g58184(.A (n_23383), .B (n_24149), .Y (n_24150));
MX2X1 g58189(.A (n_23291), .B (key[108]), .S0 (n_3340), .Y (n_24148));
MX2X1 g58190(.A (n_23289), .B (key[76]), .S0 (n_3340), .Y (n_24147));
MX2X1 g58193(.A (n_23286), .B (key[12]), .S0 (ld), .Y (n_24145));
XOR2X1 g58202(.A (n_2894), .B (n_23287), .Y (n_24144));
XOR2X1 g58205(.A (u0_rcon_1053), .B (n_23271), .Y (n_24143));
XOR2X1 g58208(.A (u0_rcon_1060), .B (n_23285), .Y (n_24142));
XOR2X1 g58214(.A (n_1526), .B (n_24137), .Y (n_24141));
XOR2X1 g58215(.A (n_15448), .B (n_23263), .Y (n_24140));
XOR2X1 g58218(.A (n_17372), .B (n_23283), .Y (n_24139));
XOR2X1 g58222(.A (n_10655), .B (n_24137), .Y (n_24138));
MX2X1 g58227(.A (n_805), .B (n_23397), .S0 (n_23306), .Y (n_24136));
NAND2X1 g56762(.A (n_23389), .B (n_23065), .Y (n_24135));
NAND2X1 g56764(.A (n_23064), .B (n_23382), .Y (n_24134));
INVX1 g56765(.A (n_24132), .Y (n_24133));
NAND2X1 g56767(.A (n_23058), .B (n_23367), .Y (n_24131));
MX2X1 g58272(.A (n_23256), .B (key[118]), .S0 (n_24599), .Y(n_24130));
MX2X1 g58273(.A (key[102]), .B (n_23254), .S0 (n_360), .Y (n_24129));
MX2X1 g58275(.A (key[86]), .B (n_23252), .S0 (n_360), .Y (n_24128));
MX2X1 g58276(.A (key[70]), .B (n_23250), .S0 (n_229), .Y (n_24127));
MX2X1 g58278(.A (key[22]), .B (n_23248), .S0 (n_360), .Y (n_24126));
MX2X1 g58279(.A (key[6]), .B (n_23247), .S0 (n_229), .Y (n_24125));
XOR2X1 g57427(.A (w1[5] ), .B (n_23073), .Y (n_24124));
OAI21X1 g57428(.A0 (n_24121), .A1 (n_23399), .B0 (n_23400), .Y(n_24123));
OAI21X1 g57429(.A0 (n_24121), .A1 (n_23397), .B0 (n_23398), .Y(n_24122));
XOR2X1 g58302(.A (n_925), .B (n_22996), .Y (n_24120));
XOR2X1 g58303(.A (n_2450), .B (n_22996), .Y (n_24118));
XOR2X1 g58305(.A (n_12116), .B (n_22996), .Y (n_24116));
NAND2X1 g57453(.A (n_23066), .B (n_23347), .Y (n_24115));
XOR2X1 g58317(.A (n_1679), .B (n_23249), .Y (n_24114));
XOR2X1 g58318(.A (n_2438), .B (n_23258), .Y (n_24113));
MX2X1 g58322(.A (n_23350), .B (n_22875), .S0 (n_24103), .Y (n_24112));
INVX1 g57458(.A (n_24110), .Y (n_24111));
MX2X1 g58323(.A (n_23720), .B (n_25997), .S0 (n_28899), .Y (n_24109));
NAND2X1 g57461(.A (n_23076), .B (n_23394), .Y (n_24108));
XOR2X1 g58340(.A (n_2135), .B (n_23246), .Y (n_24105));
INVX2 g58345(.A (n_24394), .Y (n_24582));
MX2X1 g58352(.A (n_26423), .B (n_23215), .S0 (n_24103), .Y (n_24104));
INVX1 g57478(.A (n_24101), .Y (n_24102));
NAND2X1 g58390(.A (n_27522), .B (n_23657), .Y (n_24100));
INVX1 g56783(.A (n_24098), .Y (n_24099));
NAND2X1 g58392(.A (n_24096), .B (n_23771), .Y (n_24097));
NAND2X1 g58393(.A (n_24094), .B (n_23307), .Y (n_24095));
NAND2X1 g58397(.A (n_27872), .B (n_23652), .Y (n_24093));
NAND2X1 g57484(.A (n_27815), .B (n_23261), .Y (n_24092));
NAND2X1 g57486(.A (n_23369), .B (w1[16] ), .Y (n_24091));
NAND2X1 g56787(.A (n_29347), .B (n_2004), .Y (n_24090));
NAND2X1 g58407(.A (n_24316), .B (n_24303), .Y (n_24089));
NAND2X1 g57489(.A (n_23369), .B (n_112), .Y (n_24088));
NAND2X1 g58408(.A (n_22863), .B (n_24085), .Y (n_24087));
NAND2X1 g58409(.A (n_24083), .B (n_24315), .Y (n_24084));
NAND2X1 g58411(.A (n_23316), .B (n_23281), .Y (n_24082));
NAND2X1 g58416(.A (n_23802), .B (n_24085), .Y (n_24080));
NAND2X1 g58420(.A (n_23501), .B (n_23919), .Y (n_24079));
NAND2X1 g56789(.A (n_29347), .B (n_250), .Y (n_24078));
NAND2X1 g58425(.A (n_23628), .B (n_9157), .Y (n_24077));
NAND2X1 g58428(.A (n_23489), .B (n_23294), .Y (n_24076));
NAND2X1 g56791(.A (n_29350), .B (n_21708), .Y (n_24075));
XOR2X1 g57506(.A (w1[3] ), .B (n_23039), .Y (n_24073));
XOR2X1 g58441(.A (u0_rcon_1056), .B (n_24057), .Y (n_24736));
MX2X1 g57508(.A (n_1385), .B (n_2417), .S0 (n_23039), .Y (n_24072));
AOI21X1 g57510(.A0 (n_23374), .A1 (n_23747), .B0 (n_23375), .Y(n_24071));
INVX1 g58447(.A (n_24069), .Y (n_24070));
MX2X1 g58452(.A (n_22502), .B (n_22501), .S0 (n_24014), .Y (n_24068));
INVX1 g58456(.A (n_24066), .Y (n_24067));
OAI21X1 g57519(.A0 (n_23378), .A1 (n_24223), .B0 (n_23379), .Y(n_24065));
MX2X1 g58475(.A (n_23500), .B (n_26640), .S0 (n_23669), .Y (n_24293));
OAI21X1 g58485(.A0 (n_26967), .A1 (n_26634), .B0 (n_23314), .Y(n_24064));
OAI21X1 g58490(.A0 (n_24289), .A1 (n_28907), .B0 (n_23313), .Y(n_24063));
MX2X1 g58492(.A (n_23623), .B (n_24062), .S0 (n_26534), .Y (n_24287));
INVX1 g58498(.A (n_24059), .Y (n_24060));
XOR2X1 g58501(.A (n_2430), .B (n_24057), .Y (n_24058));
INVX1 g57541(.A (n_24055), .Y (n_24056));
OAI21X1 g57543(.A0 (n_23733), .A1 (n_23352), .B0 (n_23353), .Y(n_24054));
XOR2X1 g58505(.A (n_332), .B (n_24057), .Y (n_24053));
INVX1 g57545(.A (n_24051), .Y (n_24052));
XOR2X1 g58509(.A (n_546), .B (n_23676), .Y (n_24050));
XOR2X1 g58510(.A (n_23363), .B (n_24045), .Y (n_24049));
INVX1 g57550(.A (n_24047), .Y (n_24048));
XOR2X1 g58514(.A (n_2639), .B (n_24045), .Y (n_24046));
XOR2X1 g58515(.A (n_546), .B (n_24045), .Y (n_24044));
XOR2X1 g58516(.A (n_18669), .B (n_24045), .Y (n_24043));
NAND2X2 g58525(.A (n_23320), .B (n_23021), .Y (n_24281));
INVX1 g58529(.A (n_24041), .Y (n_24042));
MX2X1 g58538(.A (n_24196), .B (n_24273), .S0 (n_28052), .Y (n_24279));
INVX1 g58541(.A (n_24039), .Y (n_24040));
MX2X1 g58548(.A (n_24037), .B (n_24038), .S0 (n_27706), .Y (n_24869));
MX2X1 g58549(.A (n_24038), .B (n_24037), .S0 (n_27706), .Y (n_24998));
XOR2X1 g58552(.A (n_2430), .B (n_23206), .Y (n_24036));
XOR2X1 g58553(.A (n_1138), .B (n_27061), .Y (n_24035));
XOR2X1 g58556(.A (w2[24] ), .B (n_27706), .Y (n_24034));
XOR2X1 g58559(.A (w1[24] ), .B (n_26639), .Y (n_24033));
MX2X1 g58561(.A (n_24031), .B (n_24032), .S0 (n_26638), .Y (n_24850));
MX2X1 g58562(.A (n_24032), .B (n_24031), .S0 (n_26638), .Y (n_24990));
INVX1 g58563(.A (n_24575), .Y (n_24030));
MX2X1 g58570(.A (n_24028), .B (n_24029), .S0 (n_27061), .Y (n_24714));
MX2X1 g58571(.A (n_24029), .B (n_24028), .S0 (n_27061), .Y (n_24865));
INVX1 g58572(.A (n_24559), .Y (n_24027));
INVX1 g58574(.A (n_26948), .Y (n_24026));
AOI21X1 g58581(.A0 (n_23888), .A1 (n_26967), .B0 (n_23328), .Y(n_24272));
AOI21X1 g58583(.A0 (n_23887), .A1 (n_28907), .B0 (n_23327), .Y(n_24271));
MX2X1 g58600(.A (n_23173), .B (key[113]), .S0 (n_698), .Y (n_24023));
MX2X1 g58602(.A (key[105]), .B (n_23170), .S0 (n_360), .Y (n_24022));
MX2X1 g58603(.A (n_23168), .B (key[81]), .S0 (ld), .Y (n_24021));
MX2X1 g58605(.A (key[73]), .B (n_23167), .S0 (n_229), .Y (n_24019));
MX2X1 g58606(.A (n_23162), .B (key[17]), .S0 (ld), .Y (n_24017));
MX2X1 g58608(.A (key[9]), .B (n_23161), .S0 (n_229), .Y (n_24016));
XOR2X1 g58610(.A (n_29311), .B (n_23900), .Y (n_24906));
XOR2X1 g58614(.A (n_2417), .B (n_24014), .Y (n_24015));
MX2X1 g58616(.A (n_22663), .B (n_22662), .S0 (n_23160), .Y (n_24258));
XOR2X1 g58619(.A (w1[9] ), .B (n_22939), .Y (n_24013));
MX2X1 g58621(.A (n_23429), .B (n_23118), .S0 (n_26510), .Y (n_24012));
INVX1 g58622(.A (n_24010), .Y (n_24011));
MX2X1 g58624(.A (n_23119), .B (n_22851), .S0 (n_23688), .Y (n_24009));
INVX1 g58625(.A (n_24007), .Y (n_24008));
MX2X1 g58627(.A (n_23122), .B (n_22855), .S0 (n_26092), .Y (n_24006));
NAND2X1 g58633(.A (n_23036), .B (n_23330), .Y (n_24005));
XOR2X1 g58639(.A (w2[21] ), .B (n_23216), .Y (n_24004));
XOR2X1 g58641(.A (n_805), .B (n_23688), .Y (n_24003));
XOR2X1 g58644(.A (n_1564), .B (n_23179), .Y (n_24002));
XOR2X1 g58646(.A (n_1971), .B (n_23163), .Y (n_24001));
NAND2X1 g57085(.A (n_23312), .B (n_23317), .Y (n_24000));
XOR2X1 g57086(.A (n_194), .B (n_23269), .Y (n_23999));
NAND2X1 g58684(.A (n_23531), .B (n_27795), .Y (n_23998));
OAI21X1 g57087(.A0 (n_23991), .A1 (n_1018), .B0 (n_23311), .Y(n_23997));
NAND2X1 g58693(.A (n_23196), .B (n_23994), .Y (n_23996));
NAND2X1 g58694(.A (n_23195), .B (n_23476), .Y (n_23993));
OAI21X1 g57088(.A0 (n_23991), .A1 (n_23309), .B0 (n_23310), .Y(n_23992));
NAND2X1 g58697(.A (n_23989), .B (n_27522), .Y (n_23990));
NAND2X1 g58698(.A (n_23213), .B (n_24096), .Y (n_23987));
NAND2X1 g58699(.A (n_23985), .B (n_24094), .Y (n_23986));
NAND2X1 g58702(.A (n_23984), .B (n_26967), .Y (n_24465));
NAND2X1 g58709(.A (n_23983), .B (n_26217), .Y (n_24475));
OR2X1 g58712(.A (n_23983), .B (n_26217), .Y (n_24476));
NOR2X1 g58713(.A (n_24196), .B (n_26217), .Y (n_23982));
OR2X1 g58716(.A (n_28907), .B (n_23981), .Y (n_24473));
NAND2X1 g58717(.A (n_23981), .B (n_28907), .Y (n_24472));
OR2X1 g58718(.A (n_23984), .B (n_26967), .Y (n_24466));
DFFX1 u0_w_reg[3][1] (.CK (clk), .D (n_23337), .Q (w3[1] ), .QN ());
NAND2X1 g58722(.A (n_24260), .B (n_23979), .Y (n_23980));
NAND2X1 g58726(.A (n_24263), .B (n_22931), .Y (n_23978));
NAND2X1 g58732(.A (n_29133), .B (n_23519), .Y (n_23977));
NAND2X1 g58734(.A (n_24265), .B (n_23205), .Y (n_23976));
NAND2X1 g58738(.A (n_24260), .B (n_22941), .Y (n_23975));
NAND2X1 g58740(.A (n_24263), .B (n_23006), .Y (n_25632));
NAND2X1 g56837(.A (n_23819), .B (n_23344), .Y (n_23972));
NAND2X1 g58744(.A (n_26751), .B (n_26218), .Y (n_23971));
DFFX1 u0_w_reg[1][1] (.CK (clk), .D (n_23340), .Q (w1[1] ), .QN ());
DFFX1 text_out_reg[20] (.CK (clk), .D (n_23442), .Q (text_out[20]),.QN ());
DFFX1 u0_w_reg[1][23] (.CK (clk), .D (n_23391), .Q (w1[23] ), .QN());
NAND2X1 g58772(.A (n_23967), .B (n_23965), .Y (n_23968));
NAND2X1 g58773(.A (n_23965), .B (n_23114), .Y (n_23966));
NAND3X1 g58776(.A (n_22600), .B (n_23844), .C (n_23843), .Y(n_23964));
INVX2 g58794(.A (n_23962), .Y (n_23963));
NAND2X1 g57111(.A (n_23589), .B (n_23049), .Y (n_23960));
NAND3X1 g58803(.A (n_23110), .B (n_23847), .C (n_23846), .Y(n_23959));
NAND4X1 g58805(.A (n_28889), .B (n_28890), .C (n_18631), .D(n_21982), .Y (n_24231));
NAND2X1 g57113(.A (n_23165), .B (n_23617), .Y (n_23958));
DFFX1 u0_w_reg[0][1] (.CK (clk), .D (n_23341), .Q (w0[1] ), .QN ());
OAI21X1 g58826(.A0 (n_23956), .A1 (n_26781), .B0 (n_23525), .Y(n_24229));
OAI21X1 g57117(.A0 (n_23276), .A1 (n_23274), .B0 (n_23275), .Y(n_24227));
MX2X1 g58827(.A (n_22841), .B (n_23955), .S0 (n_23954), .Y (n_24840));
MX2X1 g58828(.A (n_23955), .B (n_23107), .S0 (n_23954), .Y (n_24699));
NAND2X1 g57118(.A (n_28895), .B (n_28896), .Y (n_28286));
MX2X1 g58830(.A (n_22882), .B (key[100]), .S0 (n_698), .Y (n_23952));
MX2X1 g58832(.A (n_22880), .B (key[68]), .S0 (n_25126), .Y (n_23951));
MX2X1 g58834(.A (n_22877), .B (key[4]), .S0 (n_25126), .Y (n_23950));
XOR2X1 g58843(.A (n_1544), .B (n_22878), .Y (n_23949));
XOR2X1 g58844(.A (n_20153), .B (n_22895), .Y (n_23948));
INVX1 g58852(.A (n_23946), .Y (n_23947));
INVX1 g56858(.A (n_28563), .Y (n_23945));
NAND2X2 g58923(.A (n_22972), .B (n_23225), .Y (n_24212));
XOR2X1 g58859(.A (n_2559), .B (n_23941), .Y (n_23943));
XOR2X1 g58862(.A (n_15854), .B (n_23941), .Y (n_23942));
NAND2X1 g56860(.A (n_23204), .B (n_23200), .Y (n_23940));
MX2X1 g57128(.A (n_26145), .B (n_22556), .S0 (n_27391), .Y (n_23939));
XOR2X1 g56861(.A (n_19433), .B (n_23935), .Y (n_23938));
OAI21X1 g58876(.A0 (n_23714), .A1 (n_23663), .B0 (n_23224), .Y(n_23937));
OAI21X1 g56862(.A0 (n_23935), .A1 (n_4582), .B0 (n_22968), .Y(n_23936));
NAND2X1 g58883(.A (n_23934), .B (n_23933), .Y (n_24308));
AND2X1 g58884(.A (n_23934), .B (n_23933), .Y (n_24310));
OAI21X1 g58889(.A0 (n_23348), .A1 (n_26634), .B0 (n_23223), .Y(n_23932));
MX2X1 g57135(.A (n_22727), .B (n_22725), .S0 (n_27391), .Y (n_24220));
INVX1 g58891(.A (n_23929), .Y (n_23930));
INVX1 g58893(.A (n_23927), .Y (n_23928));
OAI21X1 g56863(.A0 (n_23935), .A1 (n_13466), .B0 (n_22959), .Y(n_23926));
NAND2X1 g57141(.A (n_23921), .B (w2[24] ), .Y (n_23925));
MX2X1 g58906(.A (n_23454), .B (n_27384), .S0 (n_22668), .Y (n_23924));
MX2X1 g58907(.A (n_23139), .B (n_22867), .S0 (n_25739), .Y (n_23923));
NAND2X1 g57143(.A (n_23921), .B (w2[16] ), .Y (n_23922));
NAND2X1 g56865(.A (n_23211), .B (n_22943), .Y (n_23920));
INVX1 g58915(.A (n_23919), .Y (n_24301));
NAND2X1 g57145(.A (n_23921), .B (w2[8] ), .Y (n_23918));
NAND2X1 g58920(.A (n_23226), .B (n_22973), .Y (n_24213));
INVX1 g56866(.A (n_23916), .Y (n_23917));
DFFX1 text_out_reg[86] (.CK (clk), .D (n_23177), .Q (text_out[86]),.QN ());
XOR2X1 g58939(.A (w0[0] ), .B (n_22891), .Y (n_23915));
XOR2X1 g58941(.A (n_424), .B (n_23909), .Y (n_23914));
XOR2X1 g58946(.A (n_1959), .B (n_22891), .Y (n_23912));
XOR2X1 g58948(.A (n_2924), .B (n_23909), .Y (n_23910));
INVX1 g56872(.A (n_23907), .Y (n_23908));
XOR2X1 g58953(.A (n_6085), .B (n_22891), .Y (n_23906));
XOR2X1 g58955(.A (n_6088), .B (n_23909), .Y (n_23905));
XOR2X1 g56874(.A (n_6352), .B (n_22887), .Y (n_23904));
MX2X1 g57162(.A (n_23549), .B (n_23902), .S0 (n_27068), .Y (n_23903));
NAND2X1 g58969(.A (n_23244), .B (n_22982), .Y (n_24205));
XOR2X1 g58970(.A (n_243), .B (n_23900), .Y (n_23901));
MX2X1 g57166(.A (n_1555), .B (w2[11] ), .S0 (n_23902), .Y (n_23899));
OAI21X1 g58985(.A0 (n_23896), .A1 (n_23241), .B0 (n_23242), .Y(n_23898));
NAND2X1 g58987(.A (n_23240), .B (n_22980), .Y (n_24201));
OAI21X1 g58988(.A0 (n_23896), .A1 (n_23238), .B0 (n_23239), .Y(n_23897));
NAND2X1 g58990(.A (n_23237), .B (n_22978), .Y (n_24199));
OAI21X1 g58991(.A0 (n_23896), .A1 (n_23234), .B0 (n_23236), .Y(n_23895));
XOR2X1 g58997(.A (n_3667), .B (n_22902), .Y (n_23894));
XOR2X1 g57171(.A (w2[1] ), .B (n_23584), .Y (n_23893));
INVX1 g57172(.A (n_23891), .Y (n_23892));
MX2X1 g59018(.A (n_24038), .B (n_24037), .S0 (n_23826), .Y (n_23890));
MX2X1 g59019(.A (n_24029), .B (n_24028), .S0 (n_26135), .Y (n_23889));
AOI21X1 g59023(.A0 (n_23888), .A1 (n_23231), .B0 (n_23233), .Y(n_24194));
AOI21X1 g59025(.A0 (n_23887), .A1 (n_28826), .B0 (n_23230), .Y(n_24192));
NAND2X1 g59053(.A (n_24273), .B (n_23486), .Y (n_23886));
NAND2X1 g57188(.A (n_23174), .B (n_1270), .Y (n_23885));
NOR2X1 g59063(.A (n_23883), .B (n_26104), .Y (n_23884));
NAND2X1 g59073(.A (n_24436), .B (n_23881), .Y (n_23882));
NAND2X1 g59078(.A (n_24273), .B (n_23373), .Y (n_23880));
NOR2X1 g59079(.A (n_27946), .B (n_26104), .Y (n_23879));
XOR2X1 g57204(.A (w2[2] ), .B (n_23872), .Y (n_23873));
INVX1 g59116(.A (n_23531), .Y (n_23871));
OAI21X1 g57206(.A0 (n_23869), .A1 (n_23191), .B0 (n_23192), .Y(n_24188));
NAND2X1 g59139(.A (n_23867), .B (n_22598), .Y (n_23868));
NAND2X1 g59141(.A (n_23865), .B (n_22509), .Y (n_23866));
NAND2X1 g59142(.A (n_23863), .B (n_22511), .Y (n_23864));
OAI21X1 g57208(.A0 (n_23869), .A1 (n_23184), .B0 (n_23185), .Y(n_23862));
NAND2X1 g57210(.A (n_23183), .B (n_23180), .Y (n_24185));
INVX1 g59169(.A (n_23979), .Y (n_23861));
INVX1 g57216(.A (n_23859), .Y (n_23860));
XOR2X1 g57218(.A (n_1769), .B (n_23543), .Y (n_23858));
NAND2X1 g57222(.A (n_23190), .B (n_23187), .Y (n_24183));
INVX1 g59211(.A (n_24263), .Y (n_24243));
INVX1 g59255(.A (n_23853), .Y (n_23854));
XOR2X1 g59258(.A (w2[18] ), .B (n_22644), .Y (n_23852));
INVX1 g59262(.A (n_23850), .Y (n_23851));
INVX1 g59266(.A (n_23848), .Y (n_23849));
NAND2X2 g59271(.A (n_23847), .B (n_23846), .Y (n_24232));
INVX1 g59272(.A (n_23965), .Y (n_23845));
NAND2X2 g59275(.A (n_23844), .B (n_23843), .Y (n_24235));
XOR2X1 g59276(.A (n_22717), .B (n_23503), .Y (n_23842));
XOR2X1 g59277(.A (n_6335), .B (n_22621), .Y (n_23841));
XOR2X1 g59279(.A (w2[23] ), .B (n_22859), .Y (n_23840));
NAND2X1 g59286(.A (n_23141), .B (n_23140), .Y (n_24173));
XOR2X1 g59294(.A (n_2412), .B (n_22867), .Y (n_23839));
XOR2X1 g59295(.A (n_2560), .B (n_22853), .Y (n_23838));
XOR2X1 g59333(.A (n_5305), .B (n_24306), .Y (n_23829));
XOR2X1 g59334(.A (n_5231), .B (n_22856), .Y (n_23828));
XOR2X1 g59336(.A (w2[22] ), .B (n_23826), .Y (n_23827));
NAND2X1 g59355(.A (n_23158), .B (n_23154), .Y (n_28266));
NAND2X1 g59356(.A (n_23157), .B (n_23156), .Y (n_23824));
NAND2X1 g59367(.A (n_27525), .B (n_27806), .Y (n_23822));
DFFX1 text_out_reg[81] (.CK (clk), .D (n_23280), .Q (text_out[81]),.QN ());
INVX2 g59450(.A (n_24462), .Y (n_23820));
INVX2 g59481(.A (n_23819), .Y (n_24169));
INVX1 g59550(.A (n_26781), .Y (n_23817));
INVX2 g59571(.A (n_23983), .Y (n_24607));
INVX2 g59577(.A (n_23981), .Y (n_24605));
INVX2 g59582(.A (n_23984), .Y (n_24603));
MX2X1 g59616(.A (n_23811), .B (n_23446), .S0 (n_23445), .Y (n_25015));
NAND2X1 g56738(.A (n_23109), .B (n_23106), .Y (n_23810));
XOR2X1 g59625(.A (n_22653), .B (n_22848), .Y (n_23809));
OAI21X1 g56740(.A0 (n_23805), .A1 (n_3888), .B0 (n_23105), .Y(n_25799));
DFFX1 text_out_reg[99] (.CK (clk), .D (n_23299), .Q (text_out[99]),.QN ());
OAI21X1 g56741(.A0 (n_23805), .A1 (n_9467), .B0 (n_23103), .Y(n_23806));
OAI21X1 g56742(.A0 (n_25950), .A1 (n_3038), .B0 (n_23100), .Y(n_23804));
INVX1 g59812(.A (n_23802), .Y (n_23803));
XOR2X1 g59838(.A (n_2838), .B (n_22593), .Y (n_23798));
XOR2X1 g59840(.A (n_398), .B (n_22594), .Y (n_23797));
NAND2X1 g58183(.A (n_23795), .B (n_23301), .Y (n_23796));
MX2X1 g56759(.A (n_22539), .B (n_22755), .S0 (n_29353), .Y (n_23794));
XOR2X1 g58206(.A (u0_rcon_1055), .B (n_22987), .Y (n_23793));
XOR2X1 g58210(.A (n_2086), .B (n_23788), .Y (n_23792));
MX2X1 g58211(.A (n_18549), .B (u0_rcon_1058), .S0 (n_23791), .Y(n_24390));
XOR2X1 g58212(.A (u0_rcon_1058), .B (n_23791), .Y (n_24392));
XOR2X1 g58216(.A (n_20310), .B (n_22786), .Y (n_23790));
XOR2X1 g58220(.A (n_15852), .B (n_23788), .Y (n_23789));
OAI21X1 g56766(.A0 (n_27085), .A1 (n_13679), .B0 (n_23060), .Y(n_24132));
OAI21X1 g58282(.A0 (n_26232), .A1 (n_23087), .B0 (n_23089), .Y(n_23786));
NAND2X1 g58284(.A (n_23086), .B (n_23085), .Y (n_23785));
OAI21X1 g57430(.A0 (n_26871), .A1 (n_23096), .B0 (n_23098), .Y(n_23784));
NAND2X1 g57431(.A (n_23095), .B (n_23094), .Y (n_23783));
XOR2X1 g57432(.A (n_23257), .B (n_22828), .Y (n_23782));
NAND2X1 g57438(.A (n_23090), .B (n_23092), .Y (n_23781));
XOR2X1 g58300(.A (n_645), .B (n_23791), .Y (n_23780));
XOR2X1 g58301(.A (n_497), .B (n_23791), .Y (n_23779));
MX2X1 g58304(.A (n_23777), .B (w1[5] ), .S0 (n_22996), .Y (n_23778));
NAND2X1 g57454(.A (n_23067), .B (n_23346), .Y (n_23775));
XOR2X1 g57456(.A (w1[4] ), .B (n_22824), .Y (n_23774));
NAND2X1 g57457(.A (n_23084), .B (n_23082), .Y (n_23773));
OAI21X1 g57459(.A0 (n_23083), .A1 (n_23079), .B0 (n_23080), .Y(n_24110));
MX2X1 g58324(.A (n_23883), .B (n_28119), .S0 (n_23771), .Y (n_23772));
NAND2X1 g57460(.A (n_23078), .B (n_23077), .Y (n_23770));
MX2X1 g58346(.A (n_22955), .B (n_22956), .S0 (n_23771), .Y (n_24394));
MX2X1 g57479(.A (n_22582), .B (n_22586), .S0 (n_27815), .Y (n_24101));
MX2X1 g57480(.A (n_26522), .B (n_22738), .S0 (n_27815), .Y (n_23769));
MX2X1 g56784(.A (n_23210), .B (n_22962), .S0 (n_29353), .Y (n_24098));
NAND2X1 g58398(.A (n_26232), .B (n_1019), .Y (n_23766));
NAND2X1 g58399(.A (n_26232), .B (n_23763), .Y (n_23765));
NAND2X1 g58400(.A (n_25737), .B (n_23259), .Y (n_23762));
NAND2X1 g58401(.A (n_23260), .B (n_23292), .Y (n_23761));
NAND2X1 g57485(.A (n_23758), .B (w1[24] ), .Y (n_23760));
NAND2X1 g57487(.A (n_23758), .B (n_23605), .Y (n_23759));
NAND2X1 g57488(.A (n_23758), .B (n_23567), .Y (n_23757));
NAND2X1 g58410(.A (n_23093), .B (n_24358), .Y (n_23756));
NAND2X1 g58412(.A (n_24283), .B (n_23622), .Y (n_23755));
NAND2X1 g56788(.A (n_29351), .B (n_1138), .Y (n_23754));
NAND2X1 g58426(.A (n_23629), .B (n_9156), .Y (n_23753));
NAND2X1 g58427(.A (n_23488), .B (n_23295), .Y (n_23752));
NAND2X1 g56790(.A (n_29351), .B (n_880), .Y (n_23751));
NAND2X1 g56792(.A (n_29351), .B (w3[8] ), .Y (n_23749));
MX2X1 g57509(.A (n_1072), .B (n_546), .S0 (n_23747), .Y (n_23748));
NAND2X1 g58448(.A (n_23012), .B (n_23014), .Y (n_24069));
MX2X1 g57511(.A (n_23376), .B (n_23747), .S0 (n_28903), .Y (n_23746));
INVX1 g58450(.A (n_23744), .Y (n_23745));
INVX1 g58453(.A (n_23742), .Y (n_23743));
NAND2X1 g58457(.A (n_23007), .B (n_22793), .Y (n_24066));
OAI21X1 g58468(.A0 (n_25965), .A1 (n_24285), .B0 (n_23008), .Y(n_23741));
NAND2X1 g57524(.A (n_23039), .B (w1[27] ), .Y (n_23740));
INVX1 g58481(.A (n_23738), .Y (n_23739));
INVX1 g58486(.A (n_23736), .Y (n_23737));
INVX2 g58496(.A (n_23735), .Y (n_24378));
NAND2X1 g58499(.A (n_23017), .B (n_23015), .Y (n_24059));
XOR2X1 g57540(.A (n_22778), .B (n_23733), .Y (n_23734));
XOR2X1 g58500(.A (n_2229), .B (n_23730), .Y (n_23732));
XOR2X1 g58502(.A (w0[3] ), .B (n_23730), .Y (n_23731));
OAI21X1 g57542(.A0 (n_23726), .A1 (n_23053), .B0 (n_23054), .Y(n_24055));
XOR2X1 g58503(.A (w1[3] ), .B (n_23730), .Y (n_23729));
XOR2X1 g58504(.A (n_19905), .B (n_23730), .Y (n_23728));
OAI21X1 g57544(.A0 (n_23726), .A1 (n_23047), .B0 (n_23048), .Y(n_23727));
XOR2X1 g58507(.A (n_3943), .B (n_22932), .Y (n_23725));
NAND2X1 g57546(.A (n_23045), .B (n_23042), .Y (n_24051));
XOR2X1 g57547(.A (n_97), .B (n_23374), .Y (n_23724));
NAND2X1 g57551(.A (n_23052), .B (n_23051), .Y (n_24047));
NAND2X1 g58530(.A (n_23019), .B (n_23018), .Y (n_24041));
INVX1 g57558(.A (n_23722), .Y (n_23723));
MX2X1 g58534(.A (n_23720), .B (n_22608), .S0 (n_27068), .Y (n_29402));
MX2X1 g58535(.A (n_22847), .B (n_23445), .S0 (n_28052), .Y (n_23718));
INVX1 g58539(.A (n_23715), .Y (n_23716));
MX2X1 g58542(.A (n_23887), .B (n_23714), .S0 (n_27068), .Y (n_24039));
OAI21X1 g58547(.A0 (n_26081), .A1 (n_23023), .B0 (n_23024), .Y(n_23713));
XOR2X1 g58554(.A (n_1626), .B (n_22929), .Y (n_23712));
XOR2X1 g58555(.A (w2[8] ), .B (n_28905), .Y (n_23711));
XOR2X1 g58557(.A (w2[27] ), .B (n_22942), .Y (n_23710));
NAND2X1 g56813(.A (n_23009), .B (n_23005), .Y (n_23709));
NAND2X1 g57580(.A (n_23676), .B (n_23043), .Y (n_23708));
XOR2X1 g58558(.A (n_23567), .B (n_26967), .Y (n_23707));
XOR2X1 g58560(.A (n_332), .B (n_22935), .Y (n_23706));
NAND2X1 g56814(.A (n_23003), .B (n_22999), .Y (n_23704));
NAND2X2 g58564(.A (n_23034), .B (n_22811), .Y (n_24575));
NAND2X1 g56815(.A (n_22997), .B (n_22998), .Y (n_23703));
NAND2X2 g58573(.A (n_23030), .B (n_22808), .Y (n_24559));
NAND2X1 g56816(.A (n_22993), .B (n_22995), .Y (n_23702));
XOR2X1 g56818(.A (w3[1] ), .B (n_28350), .Y (n_23701));
MX2X1 g58599(.A (n_23196), .B (n_27795), .S0 (n_24210), .Y (n_23700));
NAND2X1 g56820(.A (n_22805), .B (n_23022), .Y (n_23698));
INVX1 g56821(.A (n_23696), .Y (n_23697));
XOR2X1 g58618(.A (w2[9] ), .B (n_22744), .Y (n_23695));
OAI21X1 g58623(.A0 (n_22939), .A1 (n_23888), .B0 (n_23038), .Y(n_24010));
OAI21X1 g58626(.A0 (n_22744), .A1 (n_23887), .B0 (n_23037), .Y(n_24007));
MX2X1 g58628(.A (n_23693), .B (n_22854), .S0 (n_23332), .Y (n_23694));
NAND2X1 g58681(.A (n_26092), .B (n_22924), .Y (n_23692));
NAND2X1 g58683(.A (n_26510), .B (n_23196), .Y (n_23690));
NAND2X1 g58685(.A (n_23688), .B (n_22921), .Y (n_23689));
NAND2X1 g58688(.A (n_23528), .B (n_26327), .Y (n_23687));
NAND2X1 g56831(.A (n_28350), .B (n_23116), .Y (n_23686));
NAND2X1 g58695(.A (n_23683), .B (n_27872), .Y (n_23684));
OAI21X1 g57089(.A0 (n_25899), .A1 (n_23001), .B0 (n_23002), .Y(n_23681));
NAND2X1 g57090(.A (n_23016), .B (n_23011), .Y (n_23680));
XOR2X1 g57091(.A (w2[6] ), .B (n_22985), .Y (n_23679));
NAND2X1 g58724(.A (n_24014), .B (n_23342), .Y (n_23678));
NAND2X1 g58725(.A (n_23318), .B (n_23676), .Y (n_23677));
NAND2X1 g58728(.A (n_24273), .B (n_23674), .Y (n_23675));
NAND2X1 g58733(.A (n_23326), .B (n_26534), .Y (n_23673));
NAND2X1 g58735(.A (n_23522), .B (n_23031), .Y (n_23671));
NAND2X1 g58736(.A (n_23669), .B (n_22934), .Y (n_23670));
NAND2X1 g58739(.A (n_23667), .B (n_27364), .Y (n_23668));
NAND2X1 g58748(.A (n_27706), .B (n_23663), .Y (n_23664));
NAND2X1 g58750(.A (n_27061), .B (n_23881), .Y (n_23662));
NAND2X1 g56838(.A (n_23004), .B (n_26104), .Y (n_23661));
NAND3X1 g58774(.A (n_23115), .B (n_23497), .C (n_23496), .Y(n_23659));
INVX1 g58778(.A (n_23657), .Y (n_23656));
INVX1 g58790(.A (n_23652), .Y (n_23653));
INVX1 g58796(.A (n_24319), .Y (n_23962));
NAND2X1 g57110(.A (n_23588), .B (n_23050), .Y (n_23650));
XOR2X1 g57114(.A (w2[4] ), .B (n_22967), .Y (n_23649));
INVX1 g58816(.A (n_24149), .Y (n_24553));
NAND2X1 g57115(.A (n_23277), .B (n_23279), .Y (n_29403));
MX2X1 g58829(.A (key[116]), .B (n_22654), .S0 (n_229), .Y (n_23646));
MX2X1 g58831(.A (key[84]), .B (n_22646), .S0 (n_229), .Y (n_23644));
MX2X1 g58833(.A (key[20]), .B (n_22648), .S0 (n_229), .Y (n_23643));
OAI21X1 g58836(.A0 (n_23297), .A1 (n_22964), .B0 (n_22965), .Y(n_25517));
INVX1 g58837(.A (n_23640), .Y (n_28273));
INVX1 g58841(.A (n_23638), .Y (n_23639));
INVX1 g56852(.A (n_23636), .Y (n_23637));
XOR2X1 g58848(.A (n_1982), .B (n_22650), .Y (n_23635));
INVX1 g58850(.A (n_23633), .Y (n_23634));
OAI21X1 g58853(.A0 (n_22949), .A1 (n_27946), .B0 (n_22950), .Y(n_23946));
XOR2X1 g58854(.A (u0_rcon_1057), .B (n_22652), .Y (n_23631));
INVX1 g58855(.A (n_23629), .Y (n_23630));
INVX1 g58856(.A (n_23629), .Y (n_23628));
XOR2X1 g58861(.A (n_20322), .B (n_22647), .Y (n_23627));
INVX2 g58869(.A (n_24358), .Y (n_24083));
NAND2X1 g58887(.A (n_23626), .B (n_23625), .Y (n_24085));
AND2X1 g58888(.A (n_23626), .B (n_23625), .Y (n_24303));
AOI22X1 g58892(.A0 (n_26634), .A1 (n_22906), .B0 (n_26640), .B1(n_29200), .Y (n_23929));
AOI22X1 g58894(.A0 (n_23663), .A1 (n_28826), .B0 (n_23623), .B1(n_28825), .Y (n_23927));
INVX1 g58899(.A (n_23622), .Y (n_24361));
XOR2X1 g58902(.A (w0[17] ), .B (n_23954), .Y (n_23621));
OAI21X1 g56864(.A0 (n_26680), .A1 (n_13083), .B0 (n_22952), .Y(n_23620));
MX2X1 g58908(.A (n_22899), .B (n_22642), .S0 (n_22488), .Y (n_23619));
MX2X1 g58909(.A (n_23138), .B (n_22631), .S0 (n_22483), .Y (n_23618));
NAND2X2 g58916(.A (n_22975), .B (n_22974), .Y (n_23919));
OAI22X1 g56867(.A0 (n_22886), .A1 (n_21687), .B0 (n_22994), .B1(n_22418), .Y (n_23916));
DFFX1 text_out_reg[87] (.CK (clk), .D (n_22915), .Q (text_out[87]),.QN ());
NAND2X1 g57148(.A (n_22924), .B (n_26986), .Y (n_23617));
DFFX1 text_out_reg[17] (.CK (clk), .D (n_22989), .Q (text_out[17]),.QN ());
INVX1 g56868(.A (n_23615), .Y (n_23616));
XOR2X1 g58938(.A (n_22704), .B (n_22663), .Y (n_23614));
XOR2X1 g58940(.A (w0[10] ), .B (n_29210), .Y (n_23613));
INVX1 g56870(.A (n_23610), .Y (n_23611));
XOR2X1 g58947(.A (n_1618), .B (n_29210), .Y (n_23609));
XOR2X1 g58950(.A (w1[10] ), .B (n_29210), .Y (n_23607));
XOR2X1 g58951(.A (n_23605), .B (n_22890), .Y (n_23606));
NAND2X1 g56873(.A (n_25789), .B (n_25790), .Y (n_23907));
XOR2X1 g58954(.A (n_19900), .B (n_29210), .Y (n_23604));
MX2X1 g58958(.A (n_1958), .B (w1[0] ), .S0 (n_22891), .Y (n_23603));
NAND2X1 g56875(.A (n_22759), .B (n_22963), .Y (n_23602));
XOR2X1 g58972(.A (w0[0] ), .B (n_22671), .Y (n_23601));
XOR2X1 g58973(.A (n_23599), .B (n_23594), .Y (n_23600));
NAND2X1 g56876(.A (n_22754), .B (n_22953), .Y (n_23598));
XOR2X1 g58975(.A (w0[30] ), .B (n_23596), .Y (n_23597));
XOR2X1 g58979(.A (w1[14] ), .B (n_23594), .Y (n_23595));
NAND2X1 g56877(.A (n_22736), .B (n_22940), .Y (n_23593));
XOR2X1 g58981(.A (n_2587), .B (n_23596), .Y (n_23592));
XOR2X1 g58982(.A (n_13954), .B (n_23594), .Y (n_23591));
XOR2X1 g58992(.A (n_2131), .B (n_23594), .Y (n_23590));
INVX1 g57169(.A (n_23588), .Y (n_23589));
XOR2X1 g58996(.A (w0[31] ), .B (n_22678), .Y (n_23587));
XOR2X1 g59000(.A (w2[31] ), .B (n_22676), .Y (n_23586));
XOR2X1 g59004(.A (n_338), .B (n_22681), .Y (n_23585));
OAI21X1 g57173(.A0 (n_23584), .A1 (n_22976), .B0 (n_22977), .Y(n_23891));
XOR2X1 g59005(.A (w0[13] ), .B (n_23576), .Y (n_23583));
XOR2X1 g59006(.A (n_23580), .B (n_27741), .Y (n_23581));
XOR2X1 g59007(.A (w0[8] ), .B (n_23570), .Y (n_23579));
XOR2X1 g59008(.A (n_2913), .B (n_23576), .Y (n_23577));
INVX1 g57174(.A (n_23574), .Y (n_23575));
XOR2X1 g59009(.A (n_1683), .B (n_27741), .Y (n_23573));
XOR2X1 g59010(.A (n_2693), .B (n_23570), .Y (n_23571));
XOR2X1 g59011(.A (w1[15] ), .B (n_27741), .Y (n_23569));
XOR2X1 g59012(.A (n_23567), .B (n_23570), .Y (n_23568));
XOR2X1 g59013(.A (n_15849), .B (n_23576), .Y (n_23566));
XOR2X1 g59014(.A (n_12114), .B (n_27741), .Y (n_23565));
XOR2X1 g59015(.A (n_6083), .B (n_23570), .Y (n_23564));
MX2X1 g59016(.A (n_24276), .B (n_24275), .S0 (n_23473), .Y (n_23563));
MX2X1 g59017(.A (n_24032), .B (n_24031), .S0 (n_23176), .Y (n_23562));
NOR2X1 g59045(.A (n_24196), .B (n_23560), .Y (n_23561));
NAND2X1 g57184(.A (n_23584), .B (n_28820), .Y (n_23559));
NAND2X1 g59049(.A (n_22984), .B (n_27323), .Y (n_23558));
NAND2X1 g59051(.A (n_23556), .B (n_24196), .Y (n_23557));
NAND2X1 g59052(.A (n_24196), .B (n_22697), .Y (n_23555));
NAND2X1 g59054(.A (n_24276), .B (n_22873), .Y (n_23554));
NAND2X1 g59058(.A (n_23552), .B (n_23551), .Y (n_23553));
NAND2X1 g57189(.A (n_23549), .B (w2[27] ), .Y (n_23550));
NAND2X1 g59064(.A (n_24210), .B (n_23547), .Y (n_23548));
NAND2X1 g59065(.A (n_23552), .B (n_23545), .Y (n_23546));
NOR2X1 g57190(.A (n_23543), .B (n_23902), .Y (n_23544));
INVX1 g57192(.A (n_23921), .Y (n_23541));
NAND2X1 g59076(.A (n_22620), .B (n_27323), .Y (n_23539));
INVX1 g59082(.A (n_23537), .Y (n_23878));
NAND2X1 g59098(.A (n_23455), .B (n_23147), .Y (n_23533));
NAND2X1 g59099(.A (n_23013), .B (n_23560), .Y (n_23532));
INVX2 g59115(.A (n_26510), .Y (n_23531));
INVX1 g59131(.A (n_23985), .Y (n_23527));
NAND2X1 g59143(.A (n_26781), .B (n_22505), .Y (n_23525));
INVX4 g59158(.A (n_23667), .Y (n_24260));
MX2X1 g57211(.A (n_23543), .B (n_23182), .S0 (w2[0] ), .Y (n_23523));
INVX4 g59162(.A (n_23522), .Y (n_24265));
INVX1 g59167(.A (n_26534), .Y (n_23519));
INVX1 g59170(.A (n_26534), .Y (n_23979));
INVX1 g57212(.A (n_23517), .Y (n_23518));
INVX1 g57214(.A (n_23515), .Y (n_23516));
NAND2X1 g57217(.A (n_22721), .B (n_22918), .Y (n_23859));
INVX1 g59193(.A (n_24449), .Y (n_23514));
NAND2X1 g57220(.A (n_22711), .B (n_22914), .Y (n_23512));
NAND2X1 g57223(.A (n_22710), .B (n_22913), .Y (n_23510));
MX2X1 g59256(.A (n_23503), .B (n_26218), .S0 (n_22622), .Y (n_23853));
INVX1 g59260(.A (n_23501), .Y (n_23502));
MX2X1 g59263(.A (n_23500), .B (n_26640), .S0 (n_22640), .Y (n_23850));
MX2X1 g59267(.A (n_23499), .B (n_23498), .S0 (n_28796), .Y (n_23848));
NAND2X2 g59273(.A (n_23497), .B (n_23496), .Y (n_23965));
NAND2X1 g57239(.A (n_23872), .B (n_23494), .Y (n_23495));
XOR2X1 g59291(.A (w0[26] ), .B (n_27385), .Y (n_23493));
XOR2X1 g59292(.A (n_16978), .B (n_22632), .Y (n_23491));
XOR2X1 g59293(.A (w2[26] ), .B (n_22643), .Y (n_23490));
INVX1 g59298(.A (n_23488), .Y (n_23489));
MX2X1 g59301(.A (n_23486), .B (n_22852), .S0 (w0[0] ), .Y (n_23487));
INVX1 g59302(.A (n_23484), .Y (n_23485));
INVX1 g59304(.A (n_23482), .Y (n_23483));
INVX1 g59306(.A (n_23480), .Y (n_23481));
MX2X1 g59317(.A (n_26135), .B (n_23155), .S0 (n_23693), .Y (n_24094));
MX2X1 g59318(.A (n_23155), .B (n_26135), .S0 (n_23693), .Y (n_24096));
INVX1 g59321(.A (n_27872), .Y (n_23476));
INVX1 g59322(.A (n_27872), .Y (n_23475));
MX2X1 g59328(.A (n_26481), .B (n_22618), .S0 (n_26225), .Y (n_23994));
XOR2X1 g59332(.A (n_23255), .B (n_23473), .Y (n_23474));
XOR2X1 g59339(.A (n_2434), .B (n_29002), .Y (n_23472));
INVX1 g59360(.A (n_23470), .Y (n_23471));
NAND2X1 g59366(.A (n_23826), .B (n_23316), .Y (n_23469));
NAND2X1 g59373(.A (n_22618), .B (n_26252), .Y (n_23468));
INVX2 g59451(.A (n_24273), .Y (n_24462));
DFFX1 text_out_reg[49] (.CK (clk), .D (n_22988), .Q (text_out[49]),.QN ());
NAND2X1 g59461(.A (n_23457), .B (n_23499), .Y (n_23458));
NAND2X1 g59462(.A (n_24172), .B (n_23416), .Y (n_23456));
NAND2X2 g59471(.A (n_23454), .B (n_23455), .Y (n_24179));
INVX4 g59483(.A (n_26104), .Y (n_23819));
INVX1 g59525(.A (n_23451), .Y (n_23452));
INVX4 g59573(.A (n_23867), .Y (n_23983));
INVX2 g59579(.A (n_23863), .Y (n_23981));
INVX4 g59584(.A (n_23865), .Y (n_23984));
XOR2X1 g59597(.A (n_21552), .B (n_22600), .Y (n_23448));
INVX2 g59612(.A (n_24577), .Y (n_24576));
MX2X1 g59615(.A (n_23446), .B (n_23811), .S0 (n_23445), .Y (n_25014));
INVX1 g59617(.A (n_24564), .Y (n_23444));
XOR2X1 g59626(.A (n_530), .B (n_22603), .Y (n_23442));
XOR2X1 g59627(.A (w2[20] ), .B (n_22608), .Y (n_23441));
XOR2X1 g59628(.A (w1[20] ), .B (n_22605), .Y (n_23440));
DFFX1 text_out_reg[8] (.CK (clk), .D (n_22826), .Q (text_out[8]),.QN ());
INVX1 g59785(.A (n_23434), .Y (n_23435));
INVX1 g59806(.A (n_23431), .Y (n_23432));
INVX1 g59814(.A (n_23429), .Y (n_23802));
NAND2X1 g56753(.A (n_27034), .B (n_3014), .Y (n_23425));
NAND2X1 g56755(.A (n_23423), .B (n_23422), .Y (n_23424));
NAND2X1 g56757(.A (n_23423), .B (n_23418), .Y (n_23419));
NAND2X1 g56758(.A (n_23423), .B (n_23416), .Y (n_23417));
MX2X1 g58224(.A (key[103]), .B (n_22785), .S0 (n_229), .Y (n_23415));
MX2X1 g58226(.A (key[71]), .B (n_22784), .S0 (n_229), .Y (n_23414));
MX2X1 g58229(.A (key[7]), .B (n_22780), .S0 (n_360), .Y (n_23412));
XOR2X1 g58240(.A (n_1770), .B (n_22782), .Y (n_23411));
MX2X1 g58258(.A (key[114]), .B (n_22777), .S0 (n_229), .Y (n_23410));
MX2X1 g58259(.A (key[98]), .B (n_22775), .S0 (n_229), .Y (n_23409));
MX2X1 g58263(.A (key[82]), .B (n_22768), .S0 (n_360), .Y (n_23408));
MX2X1 g58264(.A (key[66]), .B (n_22773), .S0 (n_229), .Y (n_23407));
MX2X1 g58268(.A (key[18]), .B (n_22770), .S0 (n_229), .Y (n_23406));
MX2X1 g58269(.A (key[2]), .B (n_22769), .S0 (n_229), .Y (n_23405));
OAI21X1 g57433(.A0 (n_23402), .A1 (n_22833), .B0 (n_22834), .Y(n_28265));
OAI21X1 g57434(.A0 (n_23402), .A1 (n_22831), .B0 (n_22832), .Y(n_23403));
OAI21X1 g57435(.A0 (n_23402), .A1 (n_22829), .B0 (n_22830), .Y(n_23401));
NAND2X1 g57441(.A (n_24121), .B (n_23399), .Y (n_23400));
NAND2X1 g57443(.A (n_24121), .B (n_23397), .Y (n_23398));
XOR2X1 g58309(.A (n_2770), .B (n_22772), .Y (n_23396));
XOR2X1 g58310(.A (n_1724), .B (n_22779), .Y (n_23395));
NAND2X1 g57496(.A (n_22921), .B (n_23083), .Y (n_23394));
MX2X1 g58437(.A (n_22746), .B (n_23296), .S0 (n_28052), .Y (n_23393));
MX2X1 g58444(.A (key[119]), .B (n_22718), .S0 (n_229), .Y (n_23392));
MX2X1 g58445(.A (key[87]), .B (n_22716), .S0 (n_229), .Y (n_23391));
MX2X1 g58446(.A (key[23]), .B (n_22712), .S0 (n_229), .Y (n_23390));
NAND2X1 g56793(.A (n_26327), .B (n_22992), .Y (n_23389));
NAND2X1 g58451(.A (n_22800), .B (n_22799), .Y (n_23744));
NAND2X1 g58454(.A (n_22797), .B (n_22796), .Y (n_23742));
XOR2X1 g57512(.A (w1[1] ), .B (n_23378), .Y (n_23387));
INVX1 g57515(.A (n_23385), .Y (n_23386));
INVX1 g58465(.A (n_23795), .Y (n_23384));
INVX1 g58466(.A (n_23795), .Y (n_23383));
NAND2X1 g56796(.A (n_23366), .B (n_2838), .Y (n_23382));
XOR2X1 g58473(.A (n_2175), .B (n_22714), .Y (n_23380));
NAND2X1 g57523(.A (n_23378), .B (n_29200), .Y (n_23379));
NAND2X1 g57525(.A (n_23376), .B (n_332), .Y (n_23377));
NOR2X1 g57526(.A (n_23374), .B (n_23747), .Y (n_23375));
MX2X1 g58482(.A (n_26213), .B (n_23373), .S0 (n_25889), .Y (n_23738));
INVX1 g57529(.A (n_23758), .Y (n_23369));
MX2X1 g58487(.A (n_26640), .B (n_22442), .S0 (n_26743), .Y (n_23736));
NAND2X1 g56799(.A (n_23366), .B (n_5306), .Y (n_23367));
NAND2X2 g58497(.A (n_22801), .B (n_22802), .Y (n_23735));
XOR2X1 g58506(.A (n_23363), .B (n_25889), .Y (n_23364));
NAND2X1 g57549(.A (n_22585), .B (n_22820), .Y (n_23362));
NAND2X1 g57552(.A (n_22584), .B (n_22817), .Y (n_23361));
MX2X1 g57553(.A (n_23374), .B (n_23044), .S0 (n_1958), .Y (n_23360));
INVX1 g57554(.A (n_23356), .Y (n_23357));
INVX1 g57556(.A (n_23354), .Y (n_23355));
NAND2X1 g57559(.A (n_22578), .B (n_22816), .Y (n_23722));
NAND2X1 g57563(.A (n_23733), .B (n_23352), .Y (n_23353));
MX2X1 g58536(.A (n_23350), .B (n_22605), .S0 (n_28903), .Y (n_23351));
MX2X1 g58540(.A (n_23888), .B (n_23348), .S0 (n_28904), .Y (n_23715));
INVX1 g58545(.A (n_23346), .Y (n_23347));
XOR2X1 g56812(.A (n_14878), .B (n_23344), .Y (n_23345));
NAND2X1 g57579(.A (n_23342), .B (n_23726), .Y (n_23343));
MX2X1 g58601(.A (n_22705), .B (key[97]), .S0 (ld), .Y (n_23341));
MX2X1 g58604(.A (n_22703), .B (key[65]), .S0 (n_698), .Y (n_23340));
NAND2X1 g56819(.A (n_22812), .B (n_22573), .Y (n_23338));
MX2X1 g58607(.A (n_22700), .B (key[1]), .S0 (n_698), .Y (n_23337));
OAI21X1 g56822(.A0 (n_28344), .A1 (n_933), .B0 (n_22804), .Y(n_23696));
XOR2X1 g58645(.A (n_1936), .B (n_22701), .Y (n_23336));
NAND2X1 g58682(.A (n_23217), .B (n_26929), .Y (n_23335));
NAND2X1 g58686(.A (n_23215), .B (n_27121), .Y (n_23334));
NAND2X1 g58687(.A (n_23332), .B (n_22954), .Y (n_23333));
NAND2X1 g58689(.A (n_24255), .B (n_24196), .Y (n_23331));
NAND2X1 g58700(.A (n_22937), .B (n_26691), .Y (n_23330));
NAND2X1 g58705(.A (n_28847), .B (n_26062), .Y (n_23329));
NOR2X1 g58714(.A (n_23232), .B (n_26967), .Y (n_23328));
NOR2X1 g58715(.A (n_23326), .B (n_28907), .Y (n_23327));
OAI21X1 g57092(.A0 (n_23323), .A1 (n_22794), .B0 (n_22795), .Y(n_25537));
OAI21X1 g57093(.A0 (n_23323), .A1 (n_22789), .B0 (n_22790), .Y(n_23324));
NAND2X1 g58729(.A (n_23143), .B (n_25889), .Y (n_23322));
OAI21X1 g57094(.A0 (n_23323), .A1 (n_22787), .B0 (n_22788), .Y(n_25563));
NAND2X1 g58730(.A (n_27005), .B (n_22936), .Y (n_23320));
NAND2X1 g58737(.A (n_23318), .B (n_27574), .Y (n_23319));
NAND2X1 g57098(.A (n_23316), .B (n_25899), .Y (n_23317));
NAND2X1 g58747(.A (n_26967), .B (n_23500), .Y (n_23314));
NAND2X1 g58749(.A (n_28907), .B (n_24062), .Y (n_23313));
OR2X1 g57099(.A (n_23316), .B (n_25899), .Y (n_23312));
NAND2X1 g57102(.A (n_23991), .B (n_1018), .Y (n_23311));
NAND2X1 g57104(.A (n_23991), .B (n_23309), .Y (n_23310));
INVX1 g58779(.A (n_28899), .Y (n_23657));
INVX1 g58787(.A (n_23307), .Y (n_23308));
INVX1 g58792(.A (n_24103), .Y (n_23652));
NAND2X2 g58797(.A (n_26832), .B (n_21419), .Y (n_24319));
CLKBUFX1 g58806(.A (n_23306), .Y (n_24364));
MX2X1 g58811(.A (n_22844), .B (n_23305), .S0 (n_23304), .Y (n_24895));
MX2X1 g58812(.A (n_23305), .B (n_22844), .S0 (n_23304), .Y (n_24896));
MX2X1 g58813(.A (n_22842), .B (n_23303), .S0 (n_25739), .Y (n_24898));
MX2X1 g58814(.A (n_23303), .B (n_22842), .S0 (n_25739), .Y (n_24899));
INVX2 g58817(.A (n_23301), .Y (n_24149));
XOR2X1 g58835(.A (w0[3] ), .B (n_23297), .Y (n_23299));
OAI21X1 g58838(.A0 (n_23296), .A1 (n_22750), .B0 (n_22751), .Y(n_23640));
INVX1 g58839(.A (n_23294), .Y (n_23295));
NAND2X2 g58842(.A (n_22749), .B (n_22747), .Y (n_23638));
INVX1 g56853(.A (n_27085), .Y (n_23636));
INVX1 g58930(.A (n_23292), .Y (n_25737));
XOR2X1 g58845(.A (n_23290), .B (n_23288), .Y (n_23291));
XOR2X1 g58846(.A (n_1786), .B (n_23288), .Y (n_23289));
XOR2X1 g58847(.A (w1[12] ), .B (n_23288), .Y (n_23287));
XOR2X1 g58849(.A (n_18663), .B (n_23288), .Y (n_23286));
NAND2X1 g58851(.A (n_22757), .B (n_22560), .Y (n_23633));
MX2X1 g58857(.A (n_13279), .B (u0_rcon_1053), .S0 (n_23270), .Y(n_23629));
XOR2X1 g58860(.A (u0_rcon_1060), .B (n_23284), .Y (n_24137));
INVX2 g58870(.A (n_22991), .Y (n_24358));
XOR2X1 g58874(.A (w0[31] ), .B (n_23284), .Y (n_23285));
XOR2X1 g58878(.A (n_338), .B (n_23284), .Y (n_23283));
INVX1 g58900(.A (n_23281), .Y (n_23622));
XOR2X1 g58905(.A (w1[17] ), .B (n_25738), .Y (n_23280));
NAND2X1 g57150(.A (n_23278), .B (w2[28] ), .Y (n_23279));
NAND2X1 g57149(.A (n_23276), .B (n_1428), .Y (n_23277));
NAND2X1 g57151(.A (n_23276), .B (n_23274), .Y (n_23275));
NAND2X1 g56869(.A (n_22767), .B (n_22566), .Y (n_23615));
NAND2X1 g57152(.A (n_23276), .B (n_1004), .Y (n_28896));
NAND2X1 g57153(.A (n_23278), .B (w2[12] ), .Y (n_28895));
MX2X1 g58943(.A (n_22981), .B (n_1318), .S0 (n_23270), .Y (n_23271));
INVX2 g57154(.A (n_23991), .Y (n_23269));
NAND2X1 g56871(.A (n_22765), .B (n_22563), .Y (n_23610));
INVX1 g58959(.A (n_23266), .Y (n_23267));
INVX1 g58962(.A (n_23264), .Y (n_23265));
MX2X1 g58964(.A (w1[24] ), .B (n_23261), .S0 (n_23270), .Y(n_23263));
INVX1 g58965(.A (n_23259), .Y (n_23260));
XOR2X1 g58971(.A (n_23257), .B (n_23253), .Y (n_23258));
XOR2X1 g58974(.A (n_23255), .B (n_23251), .Y (n_23256));
XOR2X1 g58976(.A (w0[6] ), .B (n_23253), .Y (n_23254));
XOR2X1 g58977(.A (n_1916), .B (n_23251), .Y (n_23252));
XOR2X1 g58978(.A (n_2422), .B (n_23253), .Y (n_23250));
XOR2X1 g58980(.A (n_2440), .B (n_23251), .Y (n_23249));
XOR2X1 g58983(.A (n_13950), .B (n_23251), .Y (n_23248));
XOR2X1 g58984(.A (n_9155), .B (n_23253), .Y (n_23247));
OAI21X1 g57170(.A0 (n_29326), .A1 (n_9), .B0 (n_22766), .Y (n_23588));
XOR2X1 g59001(.A (n_764), .B (n_22655), .Y (n_23246));
OAI21X1 g57175(.A0 (n_29326), .A1 (n_22762), .B0 (n_22763), .Y(n_23574));
NAND2X1 g59034(.A (n_22671), .B (n_1318), .Y (n_23244));
NAND2X1 g59037(.A (n_23235), .B (n_23241), .Y (n_23242));
NAND2X1 g59038(.A (n_22671), .B (n_221), .Y (n_23240));
NAND2X1 g59041(.A (n_23235), .B (n_23238), .Y (n_23239));
NAND2X1 g59042(.A (n_22671), .B (n_2692), .Y (n_23237));
NAND2X1 g59046(.A (n_23235), .B (n_23234), .Y (n_23236));
NOR2X1 g59047(.A (n_23232), .B (n_23231), .Y (n_23233));
NOR2X1 g59048(.A (n_23326), .B (n_28826), .Y (n_23230));
NAND2X1 g59050(.A (n_22662), .B (n_23560), .Y (n_23228));
NAND2X1 g59055(.A (n_24275), .B (n_27384), .Y (n_23227));
NAND2X1 g59059(.A (n_26316), .B (n_22638), .Y (n_23226));
NAND2X1 g59062(.A (n_23025), .B (n_27043), .Y (n_23225));
NAND2X1 g59069(.A (n_23714), .B (n_24062), .Y (n_23224));
NAND2X1 g59071(.A (n_23499), .B (n_26944), .Y (n_23934));
NAND2X1 g59072(.A (n_23025), .B (n_27018), .Y (n_23933));
NAND2X1 g59075(.A (n_23348), .B (n_23500), .Y (n_23223));
NAND2X1 g59077(.A (n_24496), .B (n_23560), .Y (n_23222));
INVX1 g57195(.A (n_27391), .Y (n_23921));
INVX1 g59084(.A (n_27068), .Y (n_23537));
INVX1 g59088(.A (n_23221), .Y (n_23535));
INVX1 g59094(.A (n_23219), .Y (n_23534));
INVX1 g59107(.A (n_23217), .Y (n_23216));
INVX2 g59122(.A (n_23215), .Y (n_23688));
INVX1 g59127(.A (n_23332), .Y (n_23528));
INVX2 g59133(.A (n_23213), .Y (n_23985));
NAND2X1 g56897(.A (n_23210), .B (n_22876), .Y (n_23211));
NAND2X2 g59157(.A (n_22666), .B (n_21927), .Y (n_24045));
INVX2 g59160(.A (n_22945), .Y (n_23667));
INVX2 g59165(.A (n_22944), .Y (n_23522));
NAND2X1 g57213(.A (n_22728), .B (n_22726), .Y (n_23517));
NAND2X1 g57215(.A (n_22723), .B (n_22724), .Y (n_23515));
NAND2X1 g59178(.A (n_22665), .B (n_22341), .Y (n_24057));
INVX1 g59188(.A (n_23205), .Y (n_23206));
INVX2 g59195(.A (n_24255), .Y (n_24449));
NAND2X1 g56901(.A (n_28325), .B (n_22876), .Y (n_23204));
INVX1 g59198(.A (n_23318), .Y (n_24014));
INVX1 g59199(.A (n_23318), .Y (n_23669));
NAND2X1 g57219(.A (n_22719), .B (n_22713), .Y (n_23202));
INVX2 g59203(.A (n_23342), .Y (n_23676));
NAND2X1 g56902(.A (n_22931), .B (n_26680), .Y (n_23200));
INVX2 g59232(.A (n_23198), .Y (n_23989));
INVX1 g59242(.A (n_23196), .Y (n_23507));
INVX2 g59248(.A (n_23195), .Y (n_23683));
MX2X1 g59261(.A (n_24062), .B (n_23193), .S0 (n_22526), .Y (n_23501));
NAND2X1 g57236(.A (n_23869), .B (n_23191), .Y (n_23192));
NAND2X1 g57242(.A (n_23182), .B (n_23887), .Y (n_23190));
NAND2X1 g59296(.A (n_22698), .B (n_22696), .Y (n_23189));
NAND2X1 g59297(.A (n_22695), .B (n_22694), .Y (n_23188));
NAND2X1 g57243(.A (n_22917), .B (n_23714), .Y (n_23187));
NAND2X1 g59299(.A (n_22692), .B (n_22691), .Y (n_23488));
NAND2X1 g59300(.A (n_22689), .B (n_22688), .Y (n_29311));
NAND2X2 g59303(.A (n_25727), .B (n_25728), .Y (n_23484));
NAND2X1 g57244(.A (n_23869), .B (n_23184), .Y (n_23185));
NAND2X1 g59305(.A (n_22686), .B (n_22685), .Y (n_23482));
NAND2X2 g59307(.A (n_25714), .B (n_25715), .Y (n_23480));
NAND2X1 g57245(.A (n_23182), .B (n_23181), .Y (n_23183));
NAND2X1 g57246(.A (n_22917), .B (n_23869), .Y (n_23180));
XOR2X1 g59329(.A (w1[17] ), .B (n_23171), .Y (n_23179));
XOR2X1 g59338(.A (n_2440), .B (n_23176), .Y (n_23177));
INVX2 g57258(.A (n_23549), .Y (n_23174));
XOR2X1 g59340(.A (w0[17] ), .B (n_23171), .Y (n_23173));
XOR2X1 g59344(.A (n_23169), .B (n_23166), .Y (n_23170));
XOR2X1 g59345(.A (n_2406), .B (n_23171), .Y (n_23168));
XOR2X1 g59347(.A (n_2425), .B (n_23166), .Y (n_23167));
NAND2X1 g57147(.A (n_26929), .B (n_26987), .Y (n_23165));
XOR2X1 g59349(.A (w1[9] ), .B (n_23166), .Y (n_23163));
XOR2X1 g59350(.A (n_10654), .B (n_23171), .Y (n_23162));
XOR2X1 g59352(.A (n_13953), .B (n_23166), .Y (n_23161));
NAND2X1 g59359(.A (n_22548), .B (n_22699), .Y (n_23160));
OAI21X1 g59361(.A0 (n_29003), .A1 (n_22546), .B0 (n_22547), .Y(n_23470));
NAND2X1 g59368(.A (n_23473), .B (n_22625), .Y (n_23159));
NAND2X1 g59369(.A (n_23176), .B (n_23093), .Y (n_23158));
NAND2X1 g59370(.A (n_22628), .B (n_26135), .Y (n_23157));
NAND2X1 g59371(.A (n_23155), .B (n_25866), .Y (n_23156));
NAND2X1 g59372(.A (n_26306), .B (n_26055), .Y (n_23154));
INVX4 g59448(.A (n_23143), .Y (n_24273));
NAND2X1 g59469(.A (n_23498), .B (n_23416), .Y (n_23141));
NAND2X1 g59470(.A (n_23881), .B (n_27945), .Y (n_23140));
NAND2X1 g59472(.A (n_23013), .B (n_27384), .Y (n_24178));
NAND2X1 g59473(.A (n_22641), .B (n_23139), .Y (n_23847));
NAND2X1 g59477(.A (n_28796), .B (n_23138), .Y (n_23844));
INVX1 g59527(.A (n_23552), .Y (n_23451));
NOR2X1 g59541(.A (n_16907), .B (n_22609), .Y (n_28889));
CLKBUFX3 g59553(.A (n_26781), .Y (n_24436));
CLKBUFX3 g59574(.A (n_27196), .Y (n_23867));
CLKBUFX3 g59585(.A (n_26433), .Y (n_23865));
MX2X1 g59614(.A (n_22504), .B (n_22503), .S0 (n_25997), .Y (n_24577));
INVX1 g59618(.A (n_24565), .Y (n_24564));
INVX1 g59619(.A (n_24565), .Y (n_23135));
INVX2 g59622(.A (n_28117), .Y (n_24573));
INVX1 g59662(.A (n_23316), .Y (n_24283));
INVX1 g59680(.A (n_24285), .Y (n_23131));
INVX1 g59787(.A (n_23122), .Y (n_23434));
INVX1 g59791(.A (n_23120), .Y (n_23121));
INVX1 g59808(.A (n_23119), .Y (n_23431));
INVX1 g59815(.A (n_23118), .Y (n_23429));
INVX1 g59821(.A (n_23457), .Y (n_23117));
INVX1 g59825(.A (n_24172), .Y (n_24269));
INVX1 g59826(.A (n_24172), .Y (n_23116));
INVX1 g59906(.A (n_23114), .Y (n_23115));
INVX1 g59919(.A (n_23111), .Y (n_23110));
OR2X1 g56750(.A (n_22628), .B (n_25950), .Y (n_23109));
NAND2X1 g56751(.A (n_24512), .B (n_25950), .Y (n_23106));
NAND2X1 g56752(.A (n_25950), .B (n_3888), .Y (n_23105));
NAND2X1 g56754(.A (n_25950), .B (n_9467), .Y (n_23103));
NAND2X1 g56756(.A (n_25950), .B (n_3038), .Y (n_23100));
NAND2X1 g57445(.A (n_26871), .B (n_23096), .Y (n_23098));
OR2X1 g57447(.A (n_23093), .B (n_26871), .Y (n_23095));
NAND2X1 g57448(.A (n_23093), .B (n_26871), .Y (n_23094));
NAND2X1 g57449(.A (n_23091), .B (n_23348), .Y (n_23092));
NAND2X1 g57450(.A (n_23402), .B (n_23888), .Y (n_23090));
NAND2X1 g58402(.A (n_26232), .B (n_23087), .Y (n_23089));
OR2X1 g58403(.A (n_22625), .B (n_26232), .Y (n_23086));
NAND2X1 g58404(.A (n_22863), .B (n_26232), .Y (n_23085));
NAND2X1 g57490(.A (n_23083), .B (n_1308), .Y (n_23084));
NAND2X1 g57491(.A (n_23081), .B (n_398), .Y (n_23082));
NAND2X1 g57492(.A (n_23083), .B (n_23079), .Y (n_23080));
NAND2X1 g57493(.A (n_23083), .B (n_1005), .Y (n_23078));
NAND2X1 g57494(.A (n_23081), .B (w1[12] ), .Y (n_23077));
NAND2X1 g57495(.A (n_27121), .B (n_26404), .Y (n_23076));
INVX2 g57498(.A (n_24121), .Y (n_23073));
XOR2X1 g58439(.A (u0_rcon_1054), .B (n_22551), .Y (n_23072));
XOR2X1 g58440(.A (n_3208), .B (n_23068), .Y (n_23071));
XOR2X1 g58442(.A (n_18555), .B (n_22549), .Y (n_23070));
XOR2X1 g58443(.A (n_15856), .B (n_23068), .Y (n_23069));
INVX1 g57513(.A (n_23066), .Y (n_23067));
NAND2X1 g56794(.A (n_22752), .B (n_27085), .Y (n_23065));
OAI21X1 g57516(.A0 (n_23378), .A1 (n_22591), .B0 (n_22592), .Y(n_23385));
NAND2X1 g56795(.A (n_27085), .B (n_15473), .Y (n_23064));
INVX1 g57517(.A (n_23061), .Y (n_23062));
OAI21X1 g58467(.A0 (n_26775), .A1 (n_23416), .B0 (n_22571), .Y(n_23795));
NAND2X1 g56797(.A (n_27085), .B (n_13679), .Y (n_23060));
INVX1 g57531(.A (n_27815), .Y (n_23758));
NAND2X1 g56798(.A (n_27085), .B (n_3301), .Y (n_23058));
INVX2 g56801(.A (n_23805), .Y (n_23056));
NAND2X1 g57548(.A (n_22588), .B (n_22587), .Y (n_23055));
NAND2X1 g57555(.A (n_22583), .B (n_22581), .Y (n_23356));
INVX1 g56806(.A (n_24155), .Y (n_23358));
NAND2X1 g57557(.A (n_22580), .B (n_22579), .Y (n_23354));
NAND2X1 g57560(.A (n_23726), .B (n_23053), .Y (n_23054));
NAND2X1 g57566(.A (n_23044), .B (n_23888), .Y (n_23052));
NAND2X1 g57567(.A (n_22819), .B (n_23348), .Y (n_23051));
INVX1 g58543(.A (n_23049), .Y (n_23050));
NAND2X1 g57568(.A (n_23726), .B (n_23047), .Y (n_23048));
OAI21X1 g58546(.A0 (n_26522), .A1 (n_25741), .B0 (n_22572), .Y(n_23346));
NAND2X1 g57569(.A (n_23044), .B (n_23043), .Y (n_23045));
NAND2X1 g57570(.A (n_22819), .B (n_23726), .Y (n_23042));
INVX2 g57588(.A (n_23376), .Y (n_23039));
NAND2X1 g58690(.A (n_22737), .B (n_23232), .Y (n_23038));
NAND2X1 g58691(.A (n_22555), .B (n_23326), .Y (n_23037));
NAND2X1 g58701(.A (n_26081), .B (n_22979), .Y (n_23036));
NAND2X1 g58703(.A (n_29135), .B (n_22743), .Y (n_23034));
NAND2X1 g58706(.A (n_24275), .B (n_23031), .Y (n_23033));
NAND2X1 g58707(.A (n_26317), .B (n_22734), .Y (n_23030));
NAND2X1 g58721(.A (n_26081), .B (n_23023), .Y (n_23024));
NAND2X1 g56835(.A (n_28349), .B (n_19532), .Y (n_23022));
NAND2X1 g58731(.A (n_23232), .B (n_26743), .Y (n_23021));
NAND2X1 g58742(.A (n_25889), .B (n_29005), .Y (n_23019));
NAND2X1 g58743(.A (n_23674), .B (n_29007), .Y (n_23018));
OR2X1 g58753(.A (n_22636), .B (n_28325), .Y (n_23017));
NAND2X1 g57100(.A (n_23323), .B (n_23887), .Y (n_23016));
NAND2X1 g58754(.A (n_23881), .B (n_28325), .Y (n_23015));
NAND2X1 g58757(.A (n_23013), .B (n_23031), .Y (n_23014));
OR2X1 g58758(.A (n_23013), .B (n_23031), .Y (n_23012));
NAND2X1 g57101(.A (n_23010), .B (n_23714), .Y (n_23011));
NAND2X1 g56839(.A (n_23344), .B (n_5817), .Y (n_23009));
NAND2X1 g58764(.A (n_26775), .B (n_23499), .Y (n_23008));
NAND2X1 g58765(.A (n_28796), .B (n_23006), .Y (n_23007));
NAND2X1 g56840(.A (n_23004), .B (n_1626), .Y (n_23005));
NAND2X1 g56841(.A (n_23344), .B (n_11312), .Y (n_23003));
NAND2X1 g57106(.A (n_25899), .B (n_23001), .Y (n_23002));
INVX2 g58784(.A (n_23000), .Y (n_24345));
INVX1 g58788(.A (n_23771), .Y (n_23307));
NAND2X1 g56842(.A (n_23004), .B (n_18792), .Y (n_22999));
NAND2X2 g58793(.A (n_26631), .B (n_21106), .Y (n_24103));
NAND2X1 g56843(.A (n_23004), .B (n_3943), .Y (n_22998));
NAND2X1 g56844(.A (n_23344), .B (n_7410), .Y (n_22997));
OR4X1 g58807(.A (n_17301), .B (n_14646), .C (n_22016), .D (n_22463),.Y (n_23306));
NAND2X1 g56845(.A (n_22994), .B (n_23344), .Y (n_22995));
NAND2X1 g56846(.A (n_23210), .B (n_23004), .Y (n_22993));
MX2X1 g58818(.A (n_22505), .B (n_22507), .S0 (n_26441), .Y (n_23301));
OR4X1 g56851(.A (n_21587), .B (n_21922), .C (n_13000), .D (n_22420),.Y (n_29353));
OAI21X1 g58840(.A0 (n_23296), .A1 (n_22557), .B0 (n_22559), .Y(n_23294));
INVX1 g56855(.A (n_27085), .Y (n_22992));
INVX1 g56856(.A (n_27085), .Y (n_23366));
XOR2X1 g58858(.A (u0_rcon_1055), .B (n_22986), .Y (n_23788));
MX2X1 g58871(.A (n_22441), .B (n_26640), .S0 (n_26317), .Y (n_22991));
MX2X1 g58901(.A (n_22471), .B (n_22519), .S0 (n_29135), .Y (n_23281));
XOR2X1 g58903(.A (n_19532), .B (n_22483), .Y (n_22989));
XOR2X1 g58904(.A (w2[17] ), .B (n_23304), .Y (n_22988));
XOR2X1 g58944(.A (w0[26] ), .B (n_22986), .Y (n_22987));
CLKBUFX3 g57156(.A (n_25899), .Y (n_23991));
INVX1 g57158(.A (n_23010), .Y (n_22985));
OAI21X1 g58960(.A0 (n_28287), .A1 (n_22569), .B0 (n_22570), .Y(n_23266));
OAI21X1 g58963(.A0 (n_22984), .A1 (n_22567), .B0 (n_22568), .Y(n_23264));
OAI21X1 g58966(.A0 (n_28287), .A1 (n_22564), .B0 (n_22565), .Y(n_23259));
NAND2X1 g59035(.A (n_22979), .B (n_22981), .Y (n_22982));
NAND2X1 g59039(.A (n_22979), .B (n_424), .Y (n_22980));
NAND2X1 g59043(.A (n_22979), .B (w0[8] ), .Y (n_22978));
NAND2X1 g57186(.A (n_23584), .B (n_22976), .Y (n_22977));
NAND2X1 g59056(.A (n_29135), .B (n_22524), .Y (n_22975));
NAND2X1 g59057(.A (n_22810), .B (n_27666), .Y (n_22974));
NAND2X1 g59060(.A (n_22807), .B (n_28211), .Y (n_22973));
NAND2X1 g59061(.A (n_26944), .B (n_22522), .Y (n_22972));
NAND2X1 g59067(.A (n_24275), .B (n_26213), .Y (n_23625));
NAND2X1 g56889(.A (n_22529), .B (n_3955), .Y (n_25789));
NAND2X1 g59074(.A (n_26062), .B (n_23373), .Y (n_23626));
NAND2X1 g56890(.A (n_26680), .B (n_4582), .Y (n_22968));
INVX1 g59090(.A (n_28052), .Y (n_23221));
INVX1 g59096(.A (n_28904), .Y (n_23219));
INVX1 g57198(.A (n_23278), .Y (n_22967));
NAND2X1 g59102(.A (n_23297), .B (n_22964), .Y (n_22965));
NAND2X1 g56892(.A (n_22962), .B (n_3667), .Y (n_22963));
INVX1 g59108(.A (n_26092), .Y (n_23217));
NAND2X1 g56893(.A (n_26680), .B (n_13466), .Y (n_22959));
INVX2 g59124(.A (n_26423), .Y (n_23215));
CLKBUFX3 g59128(.A (n_22956), .Y (n_23332));
INVX1 g59129(.A (n_22956), .Y (n_22955));
INVX2 g59135(.A (n_22954), .Y (n_23213));
NAND2X1 g56895(.A (n_22962), .B (n_3868), .Y (n_22953));
NAND2X1 g56896(.A (n_26680), .B (n_13083), .Y (n_22952));
NAND2X1 g59144(.A (n_22949), .B (n_23416), .Y (n_22950));
NAND2X2 g59145(.A (n_22528), .B (n_19621), .Y (n_28907));
OR4X1 g59161(.A (n_20754), .B (n_21535), .C (n_28129), .D (n_22429),.Y (n_22945));
OR4X1 g59166(.A (n_20753), .B (n_21751), .C (n_22197), .D (n_27051),.Y (n_22944));
NAND2X1 g56898(.A (n_27948), .B (n_26680), .Y (n_22943));
INVX1 g59173(.A (n_22941), .Y (n_22942));
NAND2X1 g56899(.A (n_22962), .B (n_1616), .Y (n_22940));
INVX1 g59182(.A (n_22939), .Y (n_24241));
INVX1 g59187(.A (n_23031), .Y (n_28847));
INVX1 g59189(.A (n_23031), .Y (n_23205));
NAND2X1 g59191(.A (n_22534), .B (n_22066), .Y (n_23730));
INVX1 g59192(.A (n_26081), .Y (n_22937));
CLKBUFX3 g59196(.A (n_26081), .Y (n_24255));
INVX2 g59200(.A (n_22735), .Y (n_23318));
INVX1 g59202(.A (n_26743), .Y (n_22936));
INVX2 g59205(.A (n_26743), .Y (n_23342));
INVX1 g59208(.A (n_22934), .Y (n_22935));
OR4X1 g59215(.A (n_20396), .B (n_21530), .C (n_28178), .D (n_22427),.Y (n_24263));
INVX1 g59216(.A (n_22931), .Y (n_22932));
INVX1 g59221(.A (n_23006), .Y (n_22929));
NAND2X1 g56904(.A (n_22962), .B (n_27945), .Y (n_22928));
CLKBUFX3 g59234(.A (n_26929), .Y (n_23198));
INVX1 g59236(.A (n_26929), .Y (n_22924));
INVX2 g59243(.A (n_27794), .Y (n_23196));
CLKBUFX3 g59250(.A (n_27121), .Y (n_23195));
INVX1 g59252(.A (n_27121), .Y (n_22921));
NAND2X1 g57234(.A (n_22917), .B (w2[4] ), .Y (n_22918));
XOR2X1 g59280(.A (w1[23] ), .B (n_28883), .Y (n_22915));
NAND2X1 g57241(.A (n_22917), .B (w2[23] ), .Y (n_22914));
NAND2X1 g57248(.A (n_22917), .B (w2[15] ), .Y (n_22913));
INVX2 g57259(.A (n_22909), .Y (n_23549));
CLKBUFX3 g57260(.A (n_22909), .Y (n_23902));
INVX2 g59406(.A (n_23231), .Y (n_24223));
INVX2 g59413(.A (n_23560), .Y (n_23147));
INVX1 g59425(.A (n_23887), .Y (n_23145));
INVX1 g59429(.A (n_24028), .Y (n_22902));
INVX1 g59431(.A (n_23025), .Y (n_24029));
INVX1 g59443(.A (n_23888), .Y (n_23144));
INVX4 g59447(.A (n_26242), .Y (n_24196));
INVX2 g59454(.A (n_26241), .Y (n_23143));
NAND2X1 g59474(.A (n_22798), .B (n_28211), .Y (n_23846));
NAND2X1 g59475(.A (n_22527), .B (n_22899), .Y (n_23497));
NAND2X1 g59478(.A (n_28797), .B (n_27043), .Y (n_23843));
INVX2 g59500(.A (n_24236), .Y (n_22895));
INVX2 g57295(.A (n_23181), .Y (n_23872));
INVX2 g59528(.A (n_22892), .Y (n_23552));
INVX2 g59529(.A (n_22892), .Y (n_24210));
CLKBUFX1 g59539(.A (n_22890), .Y (n_23909));
INVX1 g59563(.A (n_23556), .Y (n_23900));
INVX1 g56941(.A (n_22886), .Y (n_22887));
XOR2X1 g59602(.A (n_22881), .B (n_29216), .Y (n_22882));
XOR2X1 g59603(.A (n_1984), .B (n_29216), .Y (n_22880));
XOR2X1 g59605(.A (w1[4] ), .B (n_29217), .Y (n_22878));
XOR2X1 g59607(.A (n_15853), .B (n_29216), .Y (n_22877));
OAI21X1 g59610(.A0 (n_22651), .A1 (u0_rcon_1057), .B0 (n_22517), .Y(n_23941));
INVX1 g56951(.A (n_22876), .Y (n_23935));
MX2X1 g59620(.A (n_22456), .B (n_22455), .S0 (n_22875), .Y (n_24565));
INVX2 g59629(.A (n_27384), .Y (n_23454));
INVX1 g59630(.A (n_27384), .Y (n_22873));
INVX2 g59663(.A (n_27806), .Y (n_23316));
INVX2 g59675(.A (n_23139), .Y (n_22867));
INVX2 g59681(.A (n_23498), .Y (n_24285));
INVX1 g59702(.A (n_24512), .Y (n_24306));
INVX1 g59709(.A (n_22863), .Y (n_24316));
INVX1 g59718(.A (n_23093), .Y (n_24315));
INVX1 g59752(.A (n_24289), .Y (n_22859));
INVX1 g59761(.A (n_27525), .Y (n_23826));
INVX1 g59773(.A (n_23155), .Y (n_22856));
INVX1 g59788(.A (n_22855), .Y (n_23122));
INVX1 g59792(.A (n_23693), .Y (n_23120));
INVX1 g59793(.A (n_23693), .Y (n_22854));
INVX1 g59800(.A (n_22852), .Y (n_22853));
INVX1 g59809(.A (n_22851), .Y (n_23119));
INVX1 g59816(.A (n_26225), .Y (n_23118));
INVX2 g59822(.A (n_22849), .Y (n_23457));
INVX2 g59827(.A (n_22849), .Y (n_24172));
INVX1 g59872(.A (n_22847), .Y (n_22848));
INVX1 g59908(.A (n_22844), .Y (n_23114));
MX2X1 g58931(.A (n_22745), .B (n_22748), .S0 (n_26691), .Y (n_23292));
INVX1 g59920(.A (n_22842), .Y (n_23111));
INVX2 g59938(.A (n_23955), .Y (n_23107));
INVX1 g59939(.A (n_23955), .Y (n_22841));
INVX1 g60019(.A (n_23811), .Y (n_23099));
NAND2X1 g57442(.A (n_23402), .B (n_22833), .Y (n_22834));
NAND2X1 g57444(.A (n_23402), .B (n_22831), .Y (n_22832));
NAND2X1 g57446(.A (n_23402), .B (n_22829), .Y (n_22830));
CLKBUFX3 g57499(.A (n_26871), .Y (n_24121));
INVX1 g57501(.A (n_23091), .Y (n_22828));
OAI21X1 g57514(.A0 (n_26978), .A1 (w1[25] ), .B0 (n_22498), .Y(n_23066));
XOR2X1 g58462(.A (w3[8] ), .B (n_25965), .Y (n_22826));
OAI21X1 g57518(.A0 (n_26978), .A1 (n_22496), .B0 (n_22497), .Y(n_23061));
INVX1 g57534(.A (n_23081), .Y (n_22824));
CLKBUFX3 g56802(.A (n_25950), .Y (n_23805));
INVX2 g56807(.A (n_22821), .Y (n_24155));
INVX2 g56808(.A (n_22821), .Y (n_23423));
NAND2X1 g57564(.A (n_22819), .B (w1[23] ), .Y (n_22820));
OAI21X1 g58544(.A0 (n_26145), .A1 (n_22487), .B0 (n_22493), .Y(n_23049));
NAND2X1 g57572(.A (n_22819), .B (w1[15] ), .Y (n_22817));
NAND2X1 g57578(.A (n_22819), .B (w1[4] ), .Y (n_22816));
INVX2 g57589(.A (n_22815), .Y (n_23376));
CLKBUFX3 g57590(.A (n_22815), .Y (n_23747));
INVX2 g57605(.A (n_23043), .Y (n_23733));
NAND2X1 g56832(.A (n_28346), .B (n_124), .Y (n_22812));
NAND2X1 g58704(.A (n_22810), .B (n_27364), .Y (n_22811));
NAND2X1 g58708(.A (n_22807), .B (n_27574), .Y (n_22808));
NAND2X1 g56834(.A (n_28350), .B (n_19908), .Y (n_22805));
NAND2X1 g56836(.A (n_26287), .B (n_933), .Y (n_22804));
NAND2X1 g58751(.A (n_23416), .B (n_28324), .Y (n_22802));
OR2X1 g58752(.A (n_22437), .B (n_28324), .Y (n_22801));
OR2X1 g58759(.A (n_22639), .B (n_27574), .Y (n_22800));
NAND2X1 g58760(.A (n_22798), .B (n_27574), .Y (n_22799));
OR2X1 g58761(.A (n_22525), .B (n_27364), .Y (n_22797));
NAND2X1 g58762(.A (n_22674), .B (n_27364), .Y (n_22796));
NAND2X1 g57103(.A (n_23323), .B (n_22794), .Y (n_22795));
NAND2X1 g58766(.A (n_28797), .B (n_26949), .Y (n_22793));
NAND2X1 g57105(.A (n_23323), .B (n_22789), .Y (n_22790));
NAND2X1 g57107(.A (n_23323), .B (n_22787), .Y (n_22788));
INVX1 g58785(.A (n_26232), .Y (n_23000));
NAND2X2 g58789(.A (n_22554), .B (n_20305), .Y (n_23771));
XOR2X1 g58933(.A (n_2412), .B (n_22986), .Y (n_22786));
OR4X1 g58808(.A (n_18366), .B (n_13054), .C (n_21814), .D (n_22434),.Y (n_23791));
OR4X1 g58810(.A (n_18356), .B (n_19355), .C (n_21813), .D (n_22433),.Y (n_22996));
XOR2X1 g58875(.A (w0[7] ), .B (n_22783), .Y (n_22785));
XOR2X1 g58877(.A (n_2561), .B (n_22783), .Y (n_22784));
XOR2X1 g58881(.A (n_22781), .B (n_22783), .Y (n_22782));
XOR2X1 g58882(.A (n_12117), .B (n_22783), .Y (n_22780));
XOR2X1 g58932(.A (n_22778), .B (n_22774), .Y (n_22779));
XOR2X1 g58942(.A (w0[18] ), .B (n_28483), .Y (n_22777));
XOR2X1 g58945(.A (w0[2] ), .B (n_22774), .Y (n_22775));
XOR2X1 g58949(.A (n_2435), .B (n_22774), .Y (n_22773));
XOR2X1 g58952(.A (w1[18] ), .B (n_28484), .Y (n_22772));
INVX1 g57159(.A (n_23323), .Y (n_23010));
XOR2X1 g58956(.A (n_17538), .B (n_28483), .Y (n_22770));
XOR2X1 g58957(.A (n_17539), .B (n_22774), .Y (n_22769));
XOR2X1 g58961(.A (n_2795), .B (n_28483), .Y (n_22768));
NAND2X1 g56884(.A (n_22764), .B (n_6400), .Y (n_22767));
NAND2X1 g57185(.A (n_29326), .B (n_9), .Y (n_22766));
NAND2X1 g56886(.A (n_22764), .B (n_14866), .Y (n_22765));
NAND2X1 g57187(.A (n_29327), .B (n_22762), .Y (n_22763));
NAND2X1 g56888(.A (n_27949), .B (n_5151), .Y (n_25790));
INVX2 g57197(.A (n_26987), .Y (n_23276));
NAND2X1 g56891(.A (n_23210), .B (n_2251), .Y (n_22759));
CLKBUFX3 g57200(.A (n_26987), .Y (n_23278));
NAND2X1 g59114(.A (n_26441), .B (n_22755), .Y (n_22757));
NAND2X1 g56894(.A (n_27949), .B (n_9202), .Y (n_22754));
NAND4X1 g59130(.A (n_25776), .B (n_21986), .C (n_25777), .D(n_16217), .Y (n_22956));
INVX2 g59136(.A (n_26327), .Y (n_22954));
INVX1 g59137(.A (n_26327), .Y (n_22752));
NAND2X1 g59140(.A (n_23296), .B (n_22750), .Y (n_22751));
NAND2X1 g59147(.A (n_22748), .B (n_23296), .Y (n_22749));
NAND2X1 g59148(.A (n_22746), .B (n_22745), .Y (n_22747));
INVX1 g59152(.A (n_22744), .Y (n_23967));
INVX1 g59172(.A (n_27364), .Y (n_22743));
INVX1 g59174(.A (n_27364), .Y (n_22941));
NOR4X1 g59177(.A (n_25885), .B (n_25883), .C (n_25882), .D (n_25880),.Y (n_23674));
INVX2 g59183(.A (n_22738), .Y (n_22939));
INVX1 g59184(.A (n_22738), .Y (n_22737));
NAND2X1 g56900(.A (n_27949), .B (n_2870), .Y (n_22736));
NAND4X1 g59190(.A (n_25685), .B (n_21533), .C (n_22252), .D(n_25686), .Y (n_23031));
OR4X1 g59201(.A (n_20750), .B (n_21532), .C (n_22196), .D (n_26937),.Y (n_22735));
INVX1 g59207(.A (n_27574), .Y (n_22734));
INVX1 g59209(.A (n_27574), .Y (n_22934));
INVX1 g59217(.A (n_28324), .Y (n_22931));
INVX2 g59222(.A (n_26949), .Y (n_23006));
NOR2X1 g59225(.A (n_22008), .B (n_22480), .Y (n_22730));
NAND2X1 g57230(.A (n_22727), .B (n_1039), .Y (n_22728));
NAND2X1 g57231(.A (n_22725), .B (w2[1] ), .Y (n_22726));
NAND2X1 g57232(.A (n_22725), .B (w2[3] ), .Y (n_22724));
NAND2X1 g57233(.A (n_22727), .B (n_1235), .Y (n_22723));
NAND2X1 g57235(.A (n_23182), .B (n_1163), .Y (n_22721));
NAND2X1 g57237(.A (n_23182), .B (n_1632), .Y (n_22719));
XOR2X1 g59281(.A (n_22717), .B (n_22715), .Y (n_22718));
XOR2X1 g59282(.A (n_1500), .B (n_22715), .Y (n_22716));
XOR2X1 g59283(.A (w1[23] ), .B (n_22715), .Y (n_22714));
NAND2X1 g57238(.A (n_22725), .B (w2[31] ), .Y (n_22713));
XOR2X1 g59284(.A (n_13952), .B (n_22715), .Y (n_22712));
NAND2X1 g57240(.A (n_23182), .B (n_2174), .Y (n_22711));
NOR4X1 g56917(.A (n_22709), .B (n_22708), .C (n_27248), .D (n_26910),.Y (n_23004));
NAND2X1 g57247(.A (n_23182), .B (n_2009), .Y (n_22710));
OR4X1 g56918(.A (n_22709), .B (n_22708), .C (n_27248), .D (n_26910),.Y (n_23344));
INVX1 g57253(.A (n_23584), .Y (n_22911));
XOR2X1 g59341(.A (n_22704), .B (n_22702), .Y (n_22705));
OR4X1 g57261(.A (n_21375), .B (n_20319), .C (n_21939), .D (n_22388),.Y (n_22909));
XOR2X1 g59346(.A (n_2511), .B (n_22702), .Y (n_22703));
XOR2X1 g59348(.A (w1[1] ), .B (n_22702), .Y (n_22701));
XOR2X1 g59351(.A (n_12115), .B (n_22702), .Y (n_22700));
NAND2X1 g59377(.A (n_29005), .B (w0[10] ), .Y (n_22699));
NAND2X1 g59379(.A (n_22697), .B (n_9203), .Y (n_22698));
NAND2X1 g59380(.A (n_22693), .B (n_22717), .Y (n_22696));
NAND2X1 g59381(.A (n_22697), .B (n_1103), .Y (n_22695));
NAND2X1 g59382(.A (n_22693), .B (w0[31] ), .Y (n_22694));
NAND2X1 g59383(.A (n_22697), .B (n_29005), .Y (n_22692));
NAND2X1 g59384(.A (n_22467), .B (n_29007), .Y (n_22691));
NAND2X1 g59385(.A (n_22697), .B (n_6404), .Y (n_22689));
NAND2X1 g59386(.A (n_22693), .B (n_23580), .Y (n_22688));
NAND2X1 g59388(.A (n_22748), .B (w0[1] ), .Y (n_25727));
NAND2X1 g59389(.A (n_22697), .B (n_16938), .Y (n_22686));
NAND2X1 g59390(.A (n_22467), .B (w0[3] ), .Y (n_22685));
NAND2X1 g59392(.A (n_22748), .B (w0[4] ), .Y (n_25714));
INVX1 g59403(.A (n_29200), .Y (n_22906));
INVX2 g59407(.A (n_29201), .Y (n_23231));
INVX4 g59415(.A (n_27323), .Y (n_23560));
INVX1 g59417(.A (n_22807), .Y (n_24032));
INVX1 g59419(.A (n_24031), .Y (n_22681));
INVX2 g59422(.A (n_29133), .Y (n_23326));
INVX2 g59426(.A (n_29134), .Y (n_23887));
CLKBUFX3 g59427(.A (n_29134), .Y (n_23714));
INVX1 g59430(.A (n_26944), .Y (n_24028));
INVX2 g59432(.A (n_26944), .Y (n_23025));
INVX1 g59437(.A (n_24275), .Y (n_22678));
INVX2 g59440(.A (n_27005), .Y (n_23232));
INVX2 g59444(.A (n_27005), .Y (n_23888));
CLKBUFX3 g59445(.A (n_27005), .Y (n_23348));
INVX1 g59456(.A (n_22810), .Y (n_24038));
INVX1 g59458(.A (n_24037), .Y (n_22676));
NAND4X1 g59463(.A (n_18888), .B (n_22431), .C (n_20861), .D(n_13530), .Y (n_29210));
NAND2X1 g59476(.A (n_22674), .B (n_27666), .Y (n_23496));
INVX1 g59487(.A (n_22979), .Y (n_22671));
INVX2 g59503(.A (n_22949), .Y (n_24236));
INVX1 g59517(.A (n_23023), .Y (n_22668));
INVX2 g59518(.A (n_23023), .Y (n_23954));
INVX2 g57294(.A (n_27856), .Y (n_23869));
CLKBUFX3 g57296(.A (n_27856), .Y (n_23181));
INVX2 g59530(.A (n_22536), .Y (n_22892));
NAND4X1 g59533(.A (n_29365), .B (n_21974), .C (n_29366), .D(n_22275), .Y (n_23570));
NAND4X1 g59535(.A (n_15464), .B (n_22414), .C (n_19884), .D(n_21784), .Y (n_22891));
AOI21X1 g59536(.A0 (n_18219), .A1 (n_196), .B0 (n_22462), .Y(n_22666));
NAND3X1 g59538(.A (n_13764), .B (n_22417), .C (n_21859), .Y(n_23594));
NAND3X1 g59540(.A (n_15461), .B (n_22413), .C (n_22024), .Y(n_22890));
INVX1 g59544(.A (n_22535), .Y (n_22665));
NAND4X1 g59546(.A (n_18362), .B (n_22149), .C (n_22362), .D(n_22109), .Y (n_23596));
INVX2 g59556(.A (n_22662), .Y (n_22663));
INVX2 g59562(.A (n_22660), .Y (n_23235));
INVX1 g59564(.A (n_22660), .Y (n_23556));
INVX2 g59565(.A (n_22660), .Y (n_23896));
INVX1 g56942(.A (n_22994), .Y (n_22886));
NOR3X1 g59589(.A (n_21220), .B (n_21526), .C (n_22412), .Y (n_22657));
CLKBUFX1 g59594(.A (n_22655), .Y (n_23576));
XOR2X1 g59600(.A (n_22653), .B (n_22649), .Y (n_22654));
XOR2X1 g59601(.A (n_23551), .B (n_22651), .Y (n_22652));
XOR2X1 g59604(.A (w1[20] ), .B (n_22649), .Y (n_22650));
XOR2X1 g59606(.A (n_15855), .B (n_22649), .Y (n_22648));
XOR2X1 g59608(.A (n_1308), .B (n_22651), .Y (n_22647));
XOR2X1 g59609(.A (n_2201), .B (n_22649), .Y (n_22646));
INVX2 g56952(.A (n_26680), .Y (n_22876));
INVX1 g59650(.A (n_22899), .Y (n_22643));
INVX1 g59651(.A (n_22899), .Y (n_22642));
INVX1 g59667(.A (n_22798), .Y (n_22868));
INVX1 g59668(.A (n_22798), .Y (n_22641));
INVX1 g59670(.A (n_22639), .Y (n_22640));
INVX1 g59674(.A (n_28211), .Y (n_22638));
INVX2 g59677(.A (n_28211), .Y (n_23139));
INVX2 g59679(.A (n_27018), .Y (n_23499));
CLKBUFX3 g59682(.A (n_27018), .Y (n_23498));
INVX1 g59683(.A (n_27018), .Y (n_22636));
INVX2 g59684(.A (n_27018), .Y (n_23881));
INVX1 g59695(.A (n_23138), .Y (n_22632));
INVX1 g59696(.A (n_23138), .Y (n_22631));
INVX1 g59700(.A (n_25866), .Y (n_22628));
INVX2 g59703(.A (n_25866), .Y (n_24512));
INVX1 g59710(.A (n_26252), .Y (n_22863));
INVX1 g59711(.A (n_26252), .Y (n_22625));
INVX2 g59719(.A (n_26055), .Y (n_23093));
INVX1 g59721(.A (n_23013), .Y (n_22622));
INVX2 g59724(.A (n_23013), .Y (n_23455));
INVX2 g59741(.A (n_23503), .Y (n_24496));
INVX1 g59746(.A (n_26218), .Y (n_22620));
INVX2 g59753(.A (n_23193), .Y (n_24289));
INVX1 g59766(.A (n_22618), .Y (n_23473));
INVX2 g59774(.A (n_26135), .Y (n_23155));
INVX1 g59789(.A (n_27521), .Y (n_22855));
NAND2X2 g59794(.A (n_25816), .B (n_25817), .Y (n_23693));
INVX1 g59801(.A (n_23486), .Y (n_22852));
INVX1 g59810(.A (n_26303), .Y (n_22851));
INVX2 g59828(.A (n_27918), .Y (n_22849));
OAI21X1 g59834(.A0 (n_22405), .A1 (n_22423), .B0 (n_22042), .Y(n_22609));
INVX2 g59865(.A (n_23720), .Y (n_22608));
INVX2 g59875(.A (n_23445), .Y (n_22847));
INVX2 g59880(.A (n_23350), .Y (n_22605));
INVX1 g59887(.A (n_23883), .Y (n_22603));
INVX2 g59909(.A (n_23305), .Y (n_22844));
INVX2 g59921(.A (n_23303), .Y (n_22842));
INVX1 g59928(.A (n_23956), .Y (n_22600));
INVX2 g59940(.A (n_22597), .Y (n_23955));
INVX1 g59941(.A (n_22597), .Y (n_22598));
INVX1 g59999(.A (n_22596), .Y (n_22840));
INVX1 g60000(.A (n_22596), .Y (n_22595));
INVX4 g60021(.A (n_23446), .Y (n_23811));
INVX1 g57503(.A (n_23402), .Y (n_23091));
NAND2X1 g57521(.A (n_23378), .B (n_22591), .Y (n_22592));
INVX2 g57533(.A (n_26404), .Y (n_23083));
CLKBUFX1 g57536(.A (n_26404), .Y (n_23081));
INVX2 g56809(.A (n_27034), .Y (n_22821));
NAND2X1 g57561(.A (n_23044), .B (w1[31] ), .Y (n_22588));
NAND2X1 g57562(.A (n_22586), .B (n_338), .Y (n_22587));
NAND2X1 g57565(.A (n_23044), .B (n_982), .Y (n_22585));
NAND2X1 g57571(.A (n_23044), .B (n_255), .Y (n_22584));
NAND2X1 g57573(.A (n_22582), .B (n_1040), .Y (n_22583));
NAND2X1 g57574(.A (n_22586), .B (w1[1] ), .Y (n_22581));
NAND2X1 g57575(.A (n_22582), .B (n_1236), .Y (n_22580));
NAND2X1 g57576(.A (n_22586), .B (w1[3] ), .Y (n_22579));
NAND2X1 g57577(.A (n_23044), .B (n_1164), .Y (n_22578));
OR4X1 g57591(.A (n_21372), .B (n_20313), .C (n_21758), .D (n_22334),.Y (n_22815));
INVX2 g57604(.A (n_27353), .Y (n_23726));
CLKBUFX3 g57606(.A (n_27353), .Y (n_23043));
NAND2X1 g56833(.A (n_28345), .B (n_21552), .Y (n_22573));
NAND2X1 g58720(.A (n_25826), .B (n_26522), .Y (n_22572));
NAND2X1 g58763(.A (n_26775), .B (n_22437), .Y (n_22571));
CLKBUFX3 g57160(.A (n_28226), .Y (n_23323));
NAND2X1 g59036(.A (n_28287), .B (n_22569), .Y (n_22570));
NAND2X1 g59040(.A (n_28288), .B (n_22567), .Y (n_22568));
NAND2X1 g56885(.A (n_27948), .B (w3[1] ), .Y (n_22566));
NAND2X1 g59044(.A (n_28288), .B (n_22564), .Y (n_22565));
NAND2X1 g56887(.A (n_27948), .B (n_14878), .Y (n_22563));
NAND2X1 g59120(.A (n_22482), .B (n_27015), .Y (n_22560));
NAND2X1 g59146(.A (n_28511), .B (n_22557), .Y (n_22559));
INVX2 g59153(.A (n_22556), .Y (n_22744));
INVX1 g59154(.A (n_22556), .Y (n_22555));
INVX1 g59185(.A (n_26521), .Y (n_22738));
NOR2X1 g59226(.A (n_22000), .B (n_28200), .Y (n_22554));
XOR2X1 g59229(.A (u0_rcon_1054), .B (n_22550), .Y (n_23068));
CLKBUFX3 g57254(.A (n_29327), .Y (n_23584));
XOR2X1 g59342(.A (w0[25] ), .B (n_22550), .Y (n_22551));
XOR2X1 g59358(.A (n_153), .B (n_22550), .Y (n_22549));
NAND2X1 g59376(.A (n_29007), .B (n_16921), .Y (n_22548));
NAND2X1 g59378(.A (n_29007), .B (n_22546), .Y (n_22547));
NAND2X1 g59387(.A (n_22745), .B (n_6401), .Y (n_25728));
NAND2X1 g59391(.A (n_22745), .B (n_9624), .Y (n_25715));
INVX2 g59418(.A (n_26316), .Y (n_22807));
INVX1 g59420(.A (n_26316), .Y (n_24031));
CLKBUFX1 g59436(.A (n_26061), .Y (n_24276));
INVX2 g59438(.A (n_26061), .Y (n_24275));
INVX2 g59457(.A (n_29136), .Y (n_22810));
INVX1 g59459(.A (n_29136), .Y (n_24037));
INVX2 g57281(.A (n_22727), .Y (n_22917));
INVX2 g57286(.A (n_23182), .Y (n_23543));
INVX2 g59490(.A (n_26691), .Y (n_22979));
INVX2 g59493(.A (n_22746), .Y (n_23297));
NAND3X1 g59497(.A (n_21293), .B (n_21754), .C (n_22363), .Y(n_23284));
INVX1 g59499(.A (n_22755), .Y (n_22539));
INVX2 g59504(.A (n_22755), .Y (n_22949));
INVX2 g59519(.A (n_26822), .Y (n_23023));
OR4X1 g59531(.A (n_16297), .B (n_21361), .C (n_21538), .D (n_26367),.Y (n_22536));
NAND2X1 g59537(.A (n_22435), .B (n_19031), .Y (n_23288));
NAND3X1 g59542(.A (n_18344), .B (n_22378), .C (n_22015), .Y(n_23251));
NAND4X1 g59543(.A (n_29412), .B (n_21875), .C (n_29413), .D(n_22150), .Y (n_23270));
NAND3X1 g59545(.A (n_17523), .B (n_22389), .C (n_22041), .Y(n_22535));
AOI21X1 g59547(.A0 (n_15549), .A1 (n_2826), .B0 (n_22432), .Y(n_22534));
NAND3X1 g59548(.A (n_29304), .B (n_29305), .C (n_22146), .Y(n_23253));
INVX2 g59558(.A (n_22984), .Y (n_22662));
INVX2 g59567(.A (n_26029), .Y (n_22660));
INVX2 g56939(.A (n_22764), .Y (n_22962));
INVX1 g56943(.A (n_27949), .Y (n_22994));
INVX1 g56945(.A (n_27949), .Y (n_22529));
NOR3X1 g59593(.A (n_21195), .B (n_21517), .C (n_22371), .Y (n_22528));
NAND4X1 g59595(.A (n_22422), .B (n_11378), .C (n_21659), .D(n_13531), .Y (n_22655));
INVX1 g59634(.A (n_22674), .Y (n_22644));
INVX1 g59635(.A (n_22674), .Y (n_22527));
INVX1 g59637(.A (n_22525), .Y (n_22526));
INVX1 g59649(.A (n_27666), .Y (n_22524));
INVX2 g59652(.A (n_27666), .Y (n_22899));
NAND3X1 g59654(.A (n_22424), .B (n_18394), .C (n_21603), .Y(n_23171));
INVX2 g59669(.A (n_26169), .Y (n_22798));
INVX1 g59671(.A (n_26169), .Y (n_22639));
NAND2X2 g59673(.A (n_22419), .B (n_21996), .Y (n_23166));
INVX1 g59694(.A (n_27043), .Y (n_22522));
INVX2 g59697(.A (n_27043), .Y (n_23138));
INVX2 g59725(.A (n_26943), .Y (n_23013));
INVX1 g59733(.A (n_27946), .Y (n_22621));
INVX2 g59739(.A (n_22521), .Y (n_23373));
CLKBUFX3 g59742(.A (n_22521), .Y (n_23503));
INVX1 g59754(.A (n_22519), .Y (n_23193));
INVX2 g59756(.A (n_23623), .Y (n_23663));
NAND2X1 g59764(.A (n_22651), .B (u0_rcon_1057), .Y (n_22517));
INVX2 g59767(.A (n_26481), .Y (n_22618));
INVX1 g59770(.A (n_26306), .Y (n_23176));
INVX2 g59802(.A (n_22697), .Y (n_23486));
INVX1 g59867(.A (n_25997), .Y (n_23720));
NAND2X2 g59876(.A (n_22409), .B (n_22246), .Y (n_23445));
INVX1 g59882(.A (n_22875), .Y (n_23350));
INVX1 g59888(.A (n_28119), .Y (n_23883));
INVX2 g59911(.A (n_27459), .Y (n_23305));
INVX1 g59912(.A (n_27459), .Y (n_22511));
INVX2 g59923(.A (n_22508), .Y (n_23303));
INVX1 g59924(.A (n_22508), .Y (n_22509));
INVX1 g59930(.A (n_22507), .Y (n_23956));
INVX2 g59932(.A (n_22507), .Y (n_22505));
OAI21X1 g59942(.A0 (n_22160), .A1 (sa00[0] ), .B0 (n_22403), .Y(n_22597));
INVX1 g60001(.A (n_22504), .Y (n_22596));
INVX1 g60002(.A (n_22504), .Y (n_22503));
NAND2X2 g60022(.A (n_29381), .B (n_29382), .Y (n_23446));
INVX1 g60025(.A (n_22502), .Y (n_22594));
INVX1 g60026(.A (n_22502), .Y (n_22501));
INVX1 g60033(.A (n_22500), .Y (n_22593));
CLKBUFX3 g57504(.A (n_26180), .Y (n_23402));
NAND2X1 g57520(.A (n_26977), .B (w1[25] ), .Y (n_22498));
NAND2X1 g57522(.A (n_26977), .B (n_22496), .Y (n_22497));
INVX1 g57583(.A (n_23378), .Y (n_22576));
INVX2 g57595(.A (n_22582), .Y (n_22819));
INVX2 g57600(.A (n_23044), .Y (n_23374));
NAND2X1 g58719(.A (n_26145), .B (n_22448), .Y (n_22493));
INVX1 g59155(.A (n_26144), .Y (n_22556));
NAND4X1 g59465(.A (n_19628), .B (n_21738), .C (n_22090), .D(n_22154), .Y (n_22986));
CLKBUFX3 g57280(.A (n_22490), .Y (n_22725));
INVX2 g57283(.A (n_22490), .Y (n_22727));
INVX2 g57287(.A (n_22490), .Y (n_23182));
INVX2 g59494(.A (n_28511), .Y (n_22746));
INVX2 g59505(.A (n_27015), .Y (n_22755));
INVX1 g59507(.A (n_22487), .Y (n_22488));
INVX2 g59508(.A (n_22487), .Y (n_23304));
INVX2 g59521(.A (n_22482), .Y (n_22483));
NAND4X1 g59549(.A (n_25652), .B (n_14900), .C (n_25653), .D(n_21620), .Y (n_22480));
CLKBUFX3 g59560(.A (n_28288), .Y (n_22984));
INVX1 g56938(.A (n_27948), .Y (n_23210));
INVX2 g56940(.A (n_27948), .Y (n_22764));
INVX2 g59636(.A (n_27468), .Y (n_22674));
INVX1 g59638(.A (n_27468), .Y (n_22525));
INVX2 g59743(.A (n_26212), .Y (n_22521));
INVX1 g59751(.A (n_22471), .Y (n_24062));
INVX1 g59755(.A (n_22471), .Y (n_22519));
CLKBUFX3 g59758(.A (n_22471), .Y (n_23623));
INVX2 g59795(.A (n_22745), .Y (n_22693));
INVX2 g59796(.A (n_22745), .Y (n_22467));
CLKBUFX3 g59799(.A (n_22465), .Y (n_22748));
INVX2 g59803(.A (n_22465), .Y (n_22697));
OAI21X1 g59831(.A0 (n_22093), .A1 (n_22377), .B0 (n_22356), .Y(n_22463));
OAI21X1 g59841(.A0 (n_22288), .A1 (n_22372), .B0 (n_21686), .Y(n_22462));
NAND2X2 g59883(.A (n_29114), .B (n_22128), .Y (n_22875));
INVX1 g59891(.A (n_22425), .Y (n_25816));
NAND4X1 g59899(.A (n_17277), .B (n_21970), .C (n_22119), .D(n_21675), .Y (n_29217));
OAI21X1 g59925(.A0 (n_22259), .A1 (n_1593), .B0 (n_22339), .Y(n_22508));
NAND2X2 g59933(.A (n_27273), .B (n_22361), .Y (n_22507));
NAND2X2 g60003(.A (n_22343), .B (n_22053), .Y (n_22504));
INVX1 g60027(.A (n_22456), .Y (n_22502));
INVX1 g60028(.A (n_22456), .Y (n_22455));
INVX1 g60035(.A (n_28118), .Y (n_22500));
CLKBUFX3 g57584(.A (n_26977), .Y (n_23378));
CLKBUFX3 g57594(.A (n_22451), .Y (n_22586));
INVX2 g57597(.A (n_22451), .Y (n_22582));
INVX2 g57601(.A (n_22451), .Y (n_23044));
NAND4X1 g59464(.A (n_20218), .B (n_21739), .C (n_22091), .D(n_22030), .Y (n_28484));
NAND4X1 g59466(.A (n_18886), .B (n_21737), .C (n_22089), .D(n_22028), .Y (n_22774));
INVX2 g57288(.A (n_22396), .Y (n_22490));
NAND3X1 g59498(.A (n_21295), .B (n_21553), .C (n_22224), .Y(n_22783));
INVX2 g59509(.A (n_27537), .Y (n_22487));
INVX1 g59510(.A (n_27537), .Y (n_22448));
INVX2 g59523(.A (n_26441), .Y (n_22482));
INVX2 g59642(.A (n_26640), .Y (n_23500));
INVX2 g59643(.A (n_26640), .Y (n_22442));
INVX1 g59644(.A (n_26640), .Y (n_22441));
NAND4X1 g59655(.A (n_22302), .B (n_22035), .C (n_21601), .D(n_18387), .Y (n_22702));
NAND3X1 g59656(.A (n_22317), .B (n_21755), .C (n_21495), .Y(n_22715));
INVX2 g59727(.A (n_27944), .Y (n_23416));
INVX1 g59730(.A (n_27944), .Y (n_22437));
NAND2X2 g59759(.A (n_27211), .B (n_21769), .Y (n_22471));
CLKBUFX3 g59798(.A (n_27421), .Y (n_22745));
INVX2 g59804(.A (n_27421), .Y (n_22465));
AOI21X1 g59818(.A0 (n_21605), .A1 (n_22418), .B0 (n_22327), .Y(n_22435));
NAND2X1 g59832(.A (n_22229), .B (n_22299), .Y (n_22434));
OAI21X1 g59833(.A0 (n_22092), .A1 (n_1138), .B0 (n_22298), .Y(n_22433));
OAI21X1 g59835(.A0 (n_22200), .A1 (n_22223), .B0 (n_21899), .Y(n_22432));
AOI21X1 g59859(.A0 (n_20639), .A1 (n_196), .B0 (n_22287), .Y(n_22431));
AOI21X1 g59861(.A0 (n_22163), .A1 (n_18480), .B0 (n_27526), .Y(n_22429));
AOI21X1 g59884(.A0 (n_22161), .A1 (n_18470), .B0 (n_825), .Y(n_22427));
NAND4X1 g59892(.A (n_25770), .B (n_25771), .C (n_21992), .D(n_20275), .Y (n_22425));
AOI21X1 g59893(.A0 (n_22187), .A1 (n_22423), .B0 (n_22036), .Y(n_22424));
AOI21X1 g59895(.A0 (n_22067), .A1 (n_21687), .B0 (n_22289), .Y(n_22422));
NAND4X1 g59896(.A (n_18382), .B (n_22113), .C (n_21984), .D(n_22017), .Y (n_22649));
NAND4X1 g59898(.A (n_17289), .B (n_21797), .C (n_21983), .D(n_22013), .Y (n_22651));
NAND2X1 g56971(.A (n_25702), .B (n_25703), .Y (n_22420));
AOI21X1 g59902(.A0 (n_21353), .A1 (n_22418), .B0 (n_22297), .Y(n_22419));
AOI21X1 g59914(.A0 (n_21802), .A1 (n_22353), .B0 (n_22313), .Y(n_22417));
AOI22X1 g59945(.A0 (n_22168), .A1 (n_1138), .B0 (n_21093), .B1(n_22301), .Y (n_22414));
AOI22X1 g59947(.A0 (n_22167), .A1 (w3[8] ), .B0 (n_21811), .B1(n_22423), .Y (n_22413));
OAI21X1 g59948(.A0 (n_22178), .A1 (n_26619), .B0 (n_22152), .Y(n_22412));
INVX1 g59979(.A (n_22359), .Y (n_22409));
NAND2X2 g60029(.A (n_22277), .B (n_22164), .Y (n_22456));
INVX1 g60060(.A (n_22348), .Y (n_22405));
AOI21X1 g60104(.A0 (n_27504), .A1 (n_26833), .B0 (n_22117), .Y(n_29382));
AOI21X1 g60197(.A0 (n_21806), .A1 (sa00[0] ), .B0 (n_25942), .Y(n_22403));
INVX2 g57602(.A (n_28071), .Y (n_22451));
NAND3X1 g57289(.A (n_21781), .B (n_21718), .C (n_22101), .Y(n_22396));
NAND4X1 g59657(.A (n_22215), .B (n_22033), .C (n_21364), .D(n_13754), .Y (n_22550));
OAI21X1 g59853(.A0 (n_22056), .A1 (n_19020), .B0 (w3[16] ), .Y(n_22389));
AOI21X1 g57344(.A0 (n_22076), .A1 (n_18478), .B0 (n_21717), .Y(n_22388));
OAI21X1 g59870(.A0 (n_22054), .A1 (n_19072), .B0 (sa00[0] ), .Y(n_25685));
NAND2X1 g59900(.A (n_21381), .B (n_22218), .Y (n_22381));
AOI21X1 g59915(.A0 (n_21509), .A1 (n_22377), .B0 (n_22222), .Y(n_22378));
AOI21X1 g59917(.A0 (n_21505), .A1 (n_1138), .B0 (n_22221), .Y(n_29304));
OAI21X1 g59952(.A0 (n_22057), .A1 (n_21843), .B0 (n_21844), .Y(n_22371));
AOI21X1 g59962(.A0 (n_22082), .A1 (n_28179), .B0 (n_21930), .Y(n_25776));
AOI22X1 g59964(.A0 (n_22062), .A1 (w3[16] ), .B0 (n_21374), .B1(n_22214), .Y (n_22363));
NOR2X1 g59969(.A (n_20282), .B (n_22176), .Y (n_22362));
NAND2X1 g59972(.A (n_27237), .B (n_26553), .Y (n_22361));
NAND4X1 g59980(.A (n_22027), .B (n_20243), .C (n_21821), .D(n_21492), .Y (n_22359));
INVX1 g59983(.A (n_26792), .Y (n_22357));
NAND2X1 g59993(.A (n_22190), .B (w3[8] ), .Y (n_22356));
NAND2X1 g60006(.A (n_22175), .B (n_22353), .Y (n_29365));
NAND2X1 g60010(.A (n_22174), .B (sa10[0] ), .Y (n_25503));
AOI22X1 g60056(.A0 (n_27817), .A1 (n_29147), .B0 (n_21271), .B1(n_3538), .Y (n_22349));
NAND2X1 g60061(.A (n_22169), .B (n_19028), .Y (n_22348));
NOR2X1 g60103(.A (n_21822), .B (n_22118), .Y (n_22343));
INVX1 g60155(.A (n_22270), .Y (n_22341));
AOI21X1 g60195(.A0 (n_21808), .A1 (n_28207), .B0 (n_22111), .Y(n_22339));
AOI21X1 g57626(.A0 (n_22074), .A1 (n_18474), .B0 (n_344), .Y(n_22334));
NAND2X1 g59852(.A (n_22094), .B (n_21405), .Y (n_22327));
OAI21X1 g59860(.A0 (n_27342), .A1 (n_19079), .B0 (n_26012), .Y(n_22325));
OAI21X1 g59885(.A0 (n_27561), .A1 (n_19065), .B0 (sa21[0] ), .Y(n_25775));
OAI21X1 g59886(.A0 (n_21917), .A1 (n_18469), .B0 (sa03[0] ), .Y(n_22320));
OAI21X1 g57349(.A0 (n_27109), .A1 (n_20926), .B0 (n_21938), .Y(n_25812));
AOI21X1 g59916(.A0 (n_21699), .A1 (n_22377), .B0 (n_22014), .Y(n_22317));
OAI21X1 g59967(.A0 (n_17381), .A1 (n_17069), .B0 (n_22064), .Y(n_22313));
OAI21X1 g59974(.A0 (n_21870), .A1 (n_14472), .B0 (n_26920), .Y(n_22311));
OAI21X1 g59985(.A0 (n_21855), .A1 (n_18126), .B0 (n_21843), .Y(n_25477));
OAI21X1 g59992(.A0 (n_21832), .A1 (n_17307), .B0 (n_22301), .Y(n_22302));
NAND2X1 g59994(.A (n_22055), .B (n_880), .Y (n_29412));
NAND2X1 g59996(.A (n_22079), .B (w3[16] ), .Y (n_22299));
NAND2X1 g60004(.A (n_22078), .B (n_341), .Y (n_22298));
AOI21X1 g60007(.A0 (n_21831), .A1 (n_18348), .B0 (n_22418), .Y(n_22297));
NAND2X1 g60015(.A (n_22060), .B (sa03[0] ), .Y (n_22295));
NAND2X1 g60043(.A (n_22070), .B (n_22251), .Y (n_22292));
OAI21X1 g60058(.A0 (n_21860), .A1 (n_22274), .B0 (n_21630), .Y(n_22289));
AOI21X1 g60059(.A0 (n_13526), .A1 (n_20406), .B0 (n_22069), .Y(n_22288));
NAND2X1 g60065(.A (n_22077), .B (n_21688), .Y (n_22287));
NAND2X1 g60084(.A (n_21993), .B (n_27817), .Y (n_25774));
NOR2X1 g60105(.A (n_21976), .B (n_21978), .Y (n_22277));
OAI21X1 g60125(.A0 (n_21770), .A1 (n_18684), .B0 (n_22274), .Y(n_22275));
NAND4X1 g60156(.A (n_21981), .B (n_13087), .C (n_13753), .D(n_16890), .Y (n_22270));
NAND4X1 g60161(.A (n_29195), .B (n_17342), .C (n_20547), .D(n_29196), .Y (n_22269));
NOR2X1 g60174(.A (n_15182), .B (n_21979), .Y (n_22268));
NAND4X1 g60184(.A (n_25666), .B (n_17167), .C (n_21187), .D(n_25667), .Y (n_22267));
NAND4X1 g60186(.A (n_25598), .B (n_17150), .C (n_21186), .D(n_25599), .Y (n_22266));
AOI21X1 g60208(.A0 (n_20935), .A1 (n_21314), .B0 (n_22020), .Y(n_22261));
NOR2X1 g60222(.A (n_21504), .B (n_22007), .Y (n_22259));
OAI21X1 g57006(.A0 (n_26273), .A1 (n_14371), .B0 (n_27239), .Y(n_25702));
NAND2X1 g60346(.A (n_21955), .B (n_22251), .Y (n_22252));
AOI21X1 g60426(.A0 (n_21747), .A1 (sa11[0] ), .B0 (n_18759), .Y(n_22246));
OAI21X1 g57630(.A0 (n_26669), .A1 (n_20910), .B0 (n_21757), .Y(n_22240));
NAND2X1 g59854(.A (n_21937), .B (n_22214), .Y (n_22229));
AOI22X1 g59965(.A0 (n_21697), .A1 (n_341), .B0 (n_21081), .B1(n_22223), .Y (n_22224));
OAI21X1 g59968(.A0 (n_18381), .A1 (n_2718), .B0 (n_21924), .Y(n_22222));
OAI21X1 g59970(.A0 (n_17287), .A1 (n_19797), .B0 (n_21923), .Y(n_22221));
OAI21X1 g59975(.A0 (n_21683), .A1 (n_10051), .B0 (n_27786), .Y(n_22219));
OAI21X1 g59976(.A0 (n_21682), .A1 (n_17283), .B0 (n_22231), .Y(n_22218));
OAI21X1 g59995(.A0 (n_21662), .A1 (n_17296), .B0 (n_22214), .Y(n_22215));
NAND2X1 g60008(.A (n_21929), .B (n_26535), .Y (n_25652));
NAND2X2 g60009(.A (n_21910), .B (sa20[0] ), .Y (n_25476));
NAND2X1 g60041(.A (n_21928), .B (n_26405), .Y (n_25481));
NAND2X1 g60048(.A (n_27429), .B (n_22203), .Y (n_28252));
AOI21X1 g60062(.A0 (n_15205), .A1 (n_1132), .B0 (n_21920), .Y(n_22200));
AOI21X1 g60077(.A0 (n_21563), .A1 (n_20933), .B0 (n_22203), .Y(n_22197));
AOI21X1 g60082(.A0 (n_27726), .A1 (n_20916), .B0 (n_22195), .Y(n_22196));
NAND4X1 g60108(.A (n_20889), .B (n_16583), .C (n_21478), .D(n_15617), .Y (n_22190));
NAND2X1 g60114(.A (n_21839), .B (sa20[0] ), .Y (n_22189));
OR4X1 g60119(.A (n_18396), .B (n_17308), .C (n_17314), .D (n_21463),.Y (n_22187));
NOR2X1 g60162(.A (n_13563), .B (n_21826), .Y (n_22179));
NOR2X1 g60166(.A (n_13485), .B (n_21825), .Y (n_22178));
OAI21X1 g60170(.A0 (n_21632), .A1 (w3[16] ), .B0 (n_17170), .Y(n_22176));
NAND4X1 g60175(.A (n_16548), .B (n_18419), .C (n_20410), .D(n_21304), .Y (n_22175));
NAND4X1 g60176(.A (n_25706), .B (n_17257), .C (n_20882), .D(n_25707), .Y (n_22174));
NAND4X1 g60178(.A (n_16773), .B (n_17247), .C (n_20543), .D(n_21300), .Y (n_22173));
AOI21X1 g60188(.A0 (n_19569), .A1 (n_933), .B0 (n_21869), .Y(n_22169));
NAND4X1 g60191(.A (n_13543), .B (n_13758), .C (n_21343), .D(n_21240), .Y (n_22168));
NAND4X1 g60192(.A (n_16818), .B (n_15697), .C (n_21340), .D(n_21239), .Y (n_22167));
AOI21X1 g60203(.A0 (n_21609), .A1 (sa00[0] ), .B0 (n_20227), .Y(n_29381));
AOI21X1 g60204(.A0 (n_21608), .A1 (sa01[0] ), .B0 (n_20699), .Y(n_22164));
AOI21X1 g60206(.A0 (n_20936), .A1 (n_20457), .B0 (n_21857), .Y(n_22163));
AOI21X1 g60212(.A0 (n_26618), .A1 (n_21108), .B0 (n_21850), .Y(n_22161));
NOR2X1 g60214(.A (n_21513), .B (n_21863), .Y (n_22160));
NAND4X1 g60226(.A (n_25717), .B (n_19279), .C (n_20286), .D(n_25718), .Y (n_22156));
INVX1 g60275(.A (n_22029), .Y (n_22154));
NAND2X1 g60332(.A (n_21810), .B (n_26619), .Y (n_22152));
OAI21X1 g60338(.A0 (n_21730), .A1 (n_19344), .B0 (n_22214), .Y(n_22150));
AND2X1 g60342(.A (n_21765), .B (n_10805), .Y (n_22149));
NAND2X1 g60343(.A (n_21809), .B (n_26833), .Y (n_22148));
AND2X1 g60349(.A (n_21764), .B (n_11086), .Y (n_22146));
NAND2X1 g60351(.A (n_21762), .B (n_16512), .Y (n_22145));
NAND2X2 g60370(.A (n_21767), .B (n_26553), .Y (n_22143));
NAND2X1 g60387(.A (n_27261), .B (n_29324), .Y (n_25770));
AOI21X1 g60427(.A0 (n_21519), .A1 (sa12[0] ), .B0 (n_19579), .Y(n_22128));
AOI21X1 g60428(.A0 (n_21518), .A1 (sa10[0] ), .B0 (n_16310), .Y(n_22126));
AOI21X1 g60446(.A0 (n_20971), .A1 (n_1558), .B0 (n_21798), .Y(n_22119));
NAND2X1 g60462(.A (n_21800), .B (n_21647), .Y (n_22118));
NAND2X1 g60463(.A (n_21792), .B (n_21642), .Y (n_22117));
NAND2X1 g60553(.A (n_21743), .B (w3[8] ), .Y (n_22113));
NAND3X1 g60569(.A (n_28279), .B (n_28280), .C (n_20367), .Y(n_22111));
NAND2X1 g60637(.A (n_21742), .B (w3[16] ), .Y (n_22109));
NAND2X1 g57342(.A (n_26702), .B (sa31[0] ), .Y (n_22101));
NAND2X1 g59991(.A (n_21694), .B (n_22195), .Y (n_22099));
AOI21X1 g60051(.A0 (n_21406), .A1 (n_21687), .B0 (n_21626), .Y(n_22094));
NOR2X1 g60052(.A (n_21712), .B (n_18112), .Y (n_22093));
NOR2X1 g60054(.A (n_21711), .B (n_18108), .Y (n_22092));
AOI21X1 g60066(.A0 (n_21078), .A1 (n_21708), .B0 (n_21709), .Y(n_22091));
AOI21X1 g60067(.A0 (n_21363), .A1 (n_250), .B0 (n_21707), .Y(n_22090));
AOI21X1 g60068(.A0 (n_21362), .A1 (n_22223), .B0 (n_21705), .Y(n_22089));
NOR2X1 g60087(.A (n_20716), .B (n_21657), .Y (n_25515));
NAND4X1 g60092(.A (n_25612), .B (n_25613), .C (n_25596), .D(n_19928), .Y (n_22086));
NAND4X1 g60096(.A (n_28258), .B (n_18993), .C (n_28259), .D(n_19389), .Y (n_22082));
NAND4X1 g60109(.A (n_20546), .B (n_15149), .C (n_21263), .D(n_17284), .Y (n_22079));
NAND4X1 g60110(.A (n_20884), .B (n_15189), .C (n_21261), .D(n_15658), .Y (n_22078));
OAI21X1 g60115(.A0 (n_21393), .A1 (n_20098), .B0 (w3[0] ), .Y(n_22077));
AOI21X1 g60118(.A0 (n_20995), .A1 (n_20397), .B0 (n_21677), .Y(n_22076));
NAND4X1 g60127(.A (n_21635), .B (n_20573), .C (n_17725), .D(n_19646), .Y (n_22075));
AOI21X1 g60129(.A0 (n_20994), .A1 (n_20386), .B0 (n_21671), .Y(n_22074));
NAND4X1 g60150(.A (n_20274), .B (n_18820), .C (n_18285), .D(n_21002), .Y (n_22070));
NAND4X1 g60151(.A (n_21061), .B (n_21660), .C (n_17382), .D(n_21029), .Y (n_22069));
NAND4X1 g60154(.A (n_21656), .B (n_20093), .C (n_18115), .D(n_14868), .Y (n_22067));
INVX1 g60157(.A (n_21926), .Y (n_22066));
NOR2X1 g60163(.A (n_16862), .B (n_21655), .Y (n_22065));
AOI22X1 g60164(.A0 (n_21392), .A1 (n_22274), .B0 (n_15294), .B1(n_20162), .Y (n_22064));
NAND4X1 g60165(.A (n_18634), .B (n_14556), .C (n_21092), .D(n_17453), .Y (n_22063));
NAND4X1 g60171(.A (n_19292), .B (n_14157), .C (n_21087), .D(n_19145), .Y (n_22062));
NAND4X1 g60179(.A (n_16752), .B (n_19006), .C (n_20544), .D(n_21014), .Y (n_22060));
NOR2X1 g60185(.A (n_18810), .B (n_21651), .Y (n_22057));
NAND4X1 g60189(.A (n_20214), .B (n_6970), .C (n_18374), .D (n_21020),.Y (n_22056));
NAND4X1 g60193(.A (n_16845), .B (n_17335), .C (n_21060), .D(n_21238), .Y (n_22055));
NAND4X1 g60199(.A (n_20970), .B (n_21120), .C (n_18662), .D(n_21016), .Y (n_22054));
AOI21X1 g60202(.A0 (sa02[0] ), .A1 (n_28284), .B0 (n_19015), .Y(n_22053));
AOI21X1 g60211(.A0 (n_20914), .A1 (n_21133), .B0 (n_21680), .Y(n_22047));
NAND4X1 g60223(.A (n_28592), .B (n_28593), .C (n_21041), .D(n_16226), .Y (n_22046));
OAI21X1 g60249(.A0 (n_21460), .A1 (n_20594), .B0 (n_27617), .Y(n_22044));
NAND2X1 g60251(.A (n_21607), .B (n_22423), .Y (n_22042));
NAND2X1 g60253(.A (n_21606), .B (n_250), .Y (n_22041));
AOI21X1 g60267(.A0 (n_21476), .A1 (n_19360), .B0 (n_22423), .Y(n_22036));
OAI21X1 g60268(.A0 (n_21475), .A1 (n_19358), .B0 (n_1138), .Y(n_22035));
OAI21X1 g60269(.A0 (n_21474), .A1 (n_19909), .B0 (w3[16] ), .Y(n_22033));
INVX1 g60273(.A (n_21891), .Y (n_22030));
AOI21X1 g60276(.A0 (n_21477), .A1 (n_13468), .B0 (w3[17] ), .Y(n_22029));
INVX1 g60277(.A (n_21889), .Y (n_22028));
OAI21X1 g60288(.A0 (n_21493), .A1 (n_21820), .B0 (n_27192), .Y(n_22027));
AND2X1 g60297(.A (n_21604), .B (n_19882), .Y (n_22024));
NAND3X1 g60308(.A (n_25809), .B (n_20955), .C (n_19902), .Y(n_22020));
NAND2X1 g60334(.A (n_21567), .B (n_22423), .Y (n_22017));
OAI21X1 g60335(.A0 (n_17755), .A1 (n_933), .B0 (n_21599), .Y(n_22016));
AND2X1 g60336(.A (n_21585), .B (n_11139), .Y (n_22015));
AOI21X1 g60337(.A0 (n_21288), .A1 (n_20590), .B0 (w3[8] ), .Y(n_22014));
NAND2X1 g60341(.A (n_21566), .B (n_22214), .Y (n_22013));
AOI21X1 g60352(.A0 (n_21485), .A1 (n_21214), .B0 (n_27456), .Y(n_22008));
NAND4X1 g60358(.A (n_21210), .B (n_15354), .C (n_19676), .D(n_21175), .Y (n_22007));
NAND4X1 g60365(.A (n_21454), .B (n_19003), .C (n_21233), .D(n_19841), .Y (n_22005));
NAND4X1 g60373(.A (n_20428), .B (n_17203), .C (n_21200), .D(n_17594), .Y (n_29147));
NAND2X1 g60379(.A (n_21574), .B (n_16644), .Y (n_25709));
AOI21X1 g60382(.A0 (n_21484), .A1 (n_21197), .B0 (n_26553), .Y(n_22000));
NAND2X1 g60385(.A (n_21571), .B (n_16715), .Y (n_21999));
AND2X1 g60389(.A (n_21570), .B (n_15860), .Y (n_25771));
INVX1 g60403(.A (n_21837), .Y (n_21996));
NAND2X1 g60412(.A (n_18355), .B (n_21597), .Y (n_21995));
NAND2X1 g60416(.A (n_21558), .B (n_21202), .Y (n_21993));
AOI21X1 g60422(.A0 (n_21317), .A1 (n_25911), .B0 (n_18979), .Y(n_21992));
OAI21X1 g60423(.A0 (n_21316), .A1 (sa01[0] ), .B0 (n_19662), .Y(n_21991));
INVX1 g60440(.A (n_21827), .Y (n_21986));
AOI21X1 g60444(.A0 (n_21462), .A1 (n_1699), .B0 (n_21624), .Y(n_21984));
AOI21X1 g60445(.A0 (n_21461), .A1 (n_19532), .B0 (n_21622), .Y(n_21983));
AOI22X1 g60448(.A0 (n_21470), .A1 (n_20153), .B0 (n_19576), .B1(n_15516), .Y (n_21982));
AOI22X1 g60449(.A0 (n_21467), .A1 (w3[17] ), .B0 (n_3739), .B1(n_14048), .Y (n_21981));
NAND4X1 g60456(.A (n_25456), .B (n_21303), .C (n_25457), .D(n_14772), .Y (n_21979));
NAND2X1 g60464(.A (n_21615), .B (n_21638), .Y (n_21978));
NAND2X1 g60465(.A (n_21614), .B (n_21637), .Y (n_21977));
INVX1 g60492(.A (n_26360), .Y (n_21976));
INVX1 g60495(.A (n_21816), .Y (n_21975));
AND2X1 g60503(.A (n_21494), .B (n_19295), .Y (n_21974));
NAND2X1 g60562(.A (n_21506), .B (n_1138), .Y (n_21970));
NAND4X1 g60618(.A (n_21723), .B (n_19243), .C (n_20761), .D(n_17856), .Y (n_21963));
OAI21X1 g60657(.A0 (n_21431), .A1 (n_20370), .B0 (sa12[0] ), .Y(n_21960));
AOI21X1 g60664(.A0 (n_21430), .A1 (n_19974), .B0 (n_22231), .Y(n_21959));
NAND2X1 g60676(.A (n_21254), .B (n_21511), .Y (n_21956));
OAI21X1 g60677(.A0 (n_21148), .A1 (n_20862), .B0 (n_21728), .Y(n_21955));
NAND2X1 g60678(.A (n_21252), .B (n_21501), .Y (n_21954));
NAND3X1 g61016(.A (n_28552), .B (n_21113), .C (n_28553), .Y(n_21945));
AOI21X1 g57338(.A0 (n_21066), .A1 (n_21225), .B0 (n_21938), .Y(n_21939));
NAND4X1 g60053(.A (n_18887), .B (n_19930), .C (n_20688), .D(n_19311), .Y (n_21937));
NAND4X1 g60131(.A (n_21399), .B (n_20565), .C (n_12113), .D(n_18918), .Y (n_21933));
AOI21X1 g60146(.A0 (n_20874), .A1 (n_21071), .B0 (n_825), .Y(n_21930));
NAND4X1 g60147(.A (n_29424), .B (n_17974), .C (n_18283), .D(n_29425), .Y (n_21929));
NAND4X1 g60149(.A (n_29125), .B (n_19602), .C (n_18292), .D(n_29126), .Y (n_21928));
INVX1 g60152(.A (n_21701), .Y (n_21927));
NAND4X1 g60158(.A (n_21404), .B (n_13066), .C (n_18386), .D(n_16903), .Y (n_21926));
AOI22X1 g60167(.A0 (n_21095), .A1 (n_21708), .B0 (n_16524), .B1(w3[9] ), .Y (n_21924));
AOI22X1 g60172(.A0 (n_21094), .A1 (n_22223), .B0 (n_15217), .B1(n_20577), .Y (n_21923));
AND2X1 g56999(.A (n_21384), .B (sa32[0] ), .Y (n_21922));
NAND4X1 g60190(.A (n_19614), .B (n_5798), .C (n_17279), .D (n_20657),.Y (n_21920));
NAND4X1 g60201(.A (n_21243), .B (n_20948), .C (n_18658), .D(n_20644), .Y (n_21917));
NAND4X1 g60215(.A (n_19549), .B (n_19148), .C (n_20682), .D(n_16263), .Y (n_21911));
NAND4X1 g60220(.A (n_21124), .B (n_20261), .C (n_20679), .D(n_16267), .Y (n_21910));
NAND4X1 g60224(.A (n_20444), .B (n_18529), .C (n_20678), .D(n_16223), .Y (n_21909));
NAND4X1 g60235(.A (n_29383), .B (n_19742), .C (n_29384), .D(n_16164), .Y (n_21905));
NAND2X1 g60246(.A (n_21369), .B (n_26140), .Y (n_21901));
NAND2X1 g60254(.A (n_21373), .B (n_22223), .Y (n_21899));
NAND2X1 g60258(.A (n_21358), .B (n_825), .Y (n_21897));
AOI21X1 g60274(.A0 (n_21267), .A1 (n_13505), .B0 (n_1699), .Y(n_21891));
AOI21X1 g60278(.A0 (n_21262), .A1 (n_9577), .B0 (n_1558), .Y(n_21889));
AND2X1 g60298(.A (n_21366), .B (n_19872), .Y (n_21875));
NAND4X1 g60305(.A (n_19944), .B (n_15591), .C (n_20931), .D(n_17634), .Y (n_21870));
NAND3X1 g60309(.A (n_7073), .B (n_21025), .C (n_17309), .Y (n_21869));
NAND2X1 g60315(.A (n_21391), .B (n_27456), .Y (n_21867));
NAND2X1 g60316(.A (n_21390), .B (n_22231), .Y (n_21865));
NAND4X1 g60317(.A (n_21215), .B (n_16859), .C (n_19687), .D(n_20863), .Y (n_21863));
NAND3X1 g60322(.A (n_18640), .B (n_21054), .C (n_19805), .Y(n_21861));
NOR2X1 g60325(.A (n_21192), .B (n_21368), .Y (n_21860));
AND2X1 g60326(.A (n_21352), .B (n_17139), .Y (n_21859));
NAND4X1 g60327(.A (n_15702), .B (n_20595), .C (n_20859), .D(n_19693), .Y (n_21858));
NAND3X1 g60329(.A (n_28255), .B (n_15931), .C (n_28256), .Y(n_21857));
NAND4X1 g60354(.A (n_25511), .B (n_17317), .C (n_25512), .D(n_18145), .Y (n_21855));
NAND3X1 g60357(.A (n_18615), .B (n_21050), .C (n_19784), .Y(n_21853));
NAND2X1 g60361(.A (n_21389), .B (n_28194), .Y (n_21852));
NAND3X1 g60369(.A (n_12271), .B (n_21010), .C (n_19340), .Y(n_21850));
NAND3X1 g60380(.A (n_8324), .B (n_21047), .C (n_20277), .Y (n_21848));
NAND2X1 g60383(.A (n_21348), .B (n_16665), .Y (n_21847));
NAND4X1 g60390(.A (n_28322), .B (n_18281), .C (n_28323), .D(n_18148), .Y (n_21846));
NAND4X1 g60394(.A (n_25582), .B (n_19247), .C (n_25583), .D(n_17029), .Y (n_21845));
NAND2X1 g60395(.A (n_21388), .B (n_21843), .Y (n_21844));
OAI21X1 g60399(.A0 (n_21273), .A1 (n_19895), .B0 (n_825), .Y(n_21842));
NAND3X1 g60401(.A (n_20792), .B (n_21056), .C (n_20348), .Y(n_21839));
NAND4X1 g60404(.A (n_21700), .B (n_20013), .C (n_20954), .D(n_20656), .Y (n_21837));
NAND3X1 g60406(.A (n_21125), .B (n_21052), .C (n_20733), .Y(n_21835));
NAND3X1 g60407(.A (n_20762), .B (n_21046), .C (n_19927), .Y(n_21834));
NAND4X1 g60410(.A (n_29395), .B (n_29396), .C (n_21290), .D(n_14758), .Y (n_21832));
INVX1 g60413(.A (n_21661), .Y (n_21831));
AOI21X1 g60421(.A0 (n_21274), .A1 (n_20742), .B0 (n_27817), .Y(n_25708));
NAND4X1 g60441(.A (n_19084), .B (n_16651), .C (n_20856), .D(n_19153), .Y (n_21827));
NAND4X1 g60451(.A (n_17343), .B (n_21031), .C (n_18722), .D(n_14428), .Y (n_21826));
NAND4X1 g60453(.A (n_25483), .B (n_21023), .C (n_25484), .D(n_14863), .Y (n_21825));
INVX1 g60477(.A (n_21648), .Y (n_21822));
OAI21X1 g60482(.A0 (n_21209), .A1 (n_21820), .B0 (n_20729), .Y(n_21821));
OAI21X1 g60496(.A0 (n_26957), .A1 (n_18908), .B0 (n_26553), .Y(n_21816));
INVX1 g60511(.A (n_21631), .Y (n_21815));
NAND3X1 g60518(.A (n_21286), .B (n_14870), .C (n_19702), .Y(n_21814));
NAND3X1 g60519(.A (n_21284), .B (n_13139), .C (n_17419), .Y(n_21813));
NAND3X1 g60523(.A (n_28853), .B (n_17638), .C (n_28854), .Y(n_21812));
NAND4X1 g60524(.A (n_20327), .B (n_18715), .C (n_20739), .D(n_15472), .Y (n_21811));
NAND4X1 g60525(.A (n_25623), .B (n_19538), .C (n_17992), .D(n_25624), .Y (n_21810));
NAND4X1 g60527(.A (n_19898), .B (n_19524), .C (n_18847), .D(n_20783), .Y (n_21809));
NAND3X1 g60531(.A (n_20134), .B (n_17618), .C (n_21191), .Y(n_21808));
NAND3X1 g60534(.A (n_20814), .B (n_15900), .C (n_21185), .Y(n_21806));
NAND3X1 g60544(.A (n_16829), .B (n_21162), .C (n_20369), .Y(n_21803));
NAND2X1 g60546(.A (n_21469), .B (n_20375), .Y (n_21802));
NAND2X1 g60559(.A (n_21481), .B (n_16362), .Y (n_21800));
AOI21X1 g60563(.A0 (n_21149), .A1 (n_16776), .B0 (n_21552), .Y(n_21798));
NAND2X1 g60570(.A (n_21307), .B (n_880), .Y (n_21797));
NAND2X1 g60585(.A (n_27157), .B (n_21520), .Y (n_21792));
OAI21X1 g60598(.A0 (n_21194), .A1 (n_20109), .B0 (n_27192), .Y(n_28251));
NAND4X1 g60615(.A (n_21435), .B (n_20023), .C (n_20422), .D(n_15126), .Y (n_29324));
NAND4X1 g60616(.A (n_21434), .B (n_19811), .C (n_20766), .D(n_16592), .Y (n_21786));
NAND4X1 g60617(.A (n_21437), .B (n_19814), .C (n_20795), .D(n_15163), .Y (n_21785));
AOI21X1 g60622(.A0 (n_19960), .A1 (n_21552), .B0 (n_21291), .Y(n_21784));
AOI21X1 g60640(.A0 (n_21153), .A1 (n_19985), .B0 (n_26920), .Y(n_21782));
NOR2X1 g60643(.A (n_21168), .B (n_21339), .Y (n_21781));
AND2X1 g60648(.A (n_21294), .B (sa23[0] ), .Y (n_21779));
AOI21X1 g60665(.A0 (n_21154), .A1 (n_19971), .B0 (n_27786), .Y(n_21772));
NAND4X1 g60672(.A (n_19520), .B (n_10690), .C (n_20745), .D (n_7256),.Y (n_21770));
AOI21X1 g60674(.A0 (n_21169), .A1 (n_487), .B0 (n_21333), .Y(n_21769));
OAI21X1 g60679(.A0 (n_19172), .A1 (n_21396), .B0 (n_21329), .Y(n_25643));
OAI21X1 g60680(.A0 (n_21139), .A1 (n_21569), .B0 (n_21472), .Y(n_21767));
AOI22X1 g60693(.A0 (n_21163), .A1 (n_3264), .B0 (n_13475), .B1(n_1667), .Y (n_21765));
AOI22X1 g60696(.A0 (n_21165), .A1 (n_2826), .B0 (n_14698), .B1(n_1132), .Y (n_21764));
AOI22X1 g60697(.A0 (n_21146), .A1 (n_21055), .B0 (n_11389), .B1(n_638), .Y (n_21762));
AOI21X1 g57619(.A0 (n_21065), .A1 (n_21208), .B0 (n_21757), .Y(n_21758));
AOI22X1 g60716(.A0 (n_21138), .A1 (n_5131), .B0 (n_20315), .B1(n_3886), .Y (n_21756));
OAI21X1 g60740(.A0 (n_21112), .A1 (n_20808), .B0 (n_20153), .Y(n_21755));
OAI21X1 g60743(.A0 (n_21116), .A1 (n_20499), .B0 (n_19532), .Y(n_21754));
NAND2X1 g60811(.A (n_21429), .B (n_13481), .Y (n_21751));
AOI21X1 g60816(.A0 (n_13964), .A1 (n_15074), .B0 (n_21427), .Y(n_21750));
NAND3X1 g60834(.A (n_21426), .B (n_19968), .C (n_17954), .Y(n_21747));
NAND4X1 g60874(.A (n_20462), .B (n_21126), .C (n_20853), .D(n_17691), .Y (n_21743));
NAND2X1 g60892(.A (n_21433), .B (n_19989), .Y (n_21742));
AOI21X1 g60959(.A0 (n_14205), .A1 (n_21598), .B0 (n_21450), .Y(n_21739));
AOI21X1 g60962(.A0 (n_16086), .A1 (n_2702), .B0 (n_21452), .Y(n_21738));
NOR2X1 g60963(.A (n_15216), .B (n_21451), .Y (n_21737));
NAND3X1 g61052(.A (n_19533), .B (n_13680), .C (n_20747), .Y(n_21730));
NAND4X1 g61063(.A (n_19187), .B (n_14644), .C (n_20341), .D(n_13914), .Y (n_21729));
INVX1 g61074(.A (n_21473), .Y (n_21728));
OAI21X1 g61106(.A0 (n_20725), .A1 (n_869), .B0 (n_19205), .Y(n_21727));
OAI21X1 g61367(.A0 (n_20724), .A1 (n_17222), .B0 (n_21398), .Y(n_21725));
OAI21X1 g61386(.A0 (n_20720), .A1 (n_17147), .B0 (n_21447), .Y(n_21724));
NOR3X1 g61419(.A (n_18267), .B (n_7865), .C (n_20711), .Y (n_21723));
NOR2X1 g61422(.A (n_19630), .B (n_21128), .Y (n_28279));
NAND4X1 g61977(.A (n_14942), .B (n_16390), .C (n_19423), .D(n_20216), .Y (n_29323));
OAI21X1 g57341(.A0 (n_20946), .A1 (n_20780), .B0 (n_21717), .Y(n_21718));
NAND2X1 g60078(.A (n_19931), .B (n_21101), .Y (n_21712));
NAND3X1 g60079(.A (n_19401), .B (n_15836), .C (n_20686), .Y(n_21711));
AOI21X1 g60120(.A0 (n_20698), .A1 (n_19539), .B0 (n_21708), .Y(n_21709));
AOI21X1 g60121(.A0 (n_20695), .A1 (n_20080), .B0 (n_250), .Y(n_21707));
NAND4X1 g60122(.A (n_25781), .B (n_25782), .C (n_16366), .D(n_17076), .Y (n_21706));
AOI21X1 g60123(.A0 (n_20694), .A1 (n_19525), .B0 (n_22301), .Y(n_21705));
NAND4X1 g60139(.A (n_21098), .B (n_20600), .C (n_12779), .D(n_17091), .Y (n_21704));
NAND4X1 g60153(.A (n_21100), .B (n_21700), .C (n_12925), .D(n_15433), .Y (n_21701));
NAND4X1 g60168(.A (n_17528), .B (n_16477), .C (n_19640), .D(n_20267), .Y (n_21699));
NAND4X1 g60173(.A (n_19300), .B (n_16488), .C (n_20221), .D(n_19144), .Y (n_21697));
NAND4X1 g60216(.A (n_20470), .B (n_19142), .C (n_20212), .D(n_16175), .Y (n_21694));
OAI21X1 g57005(.A0 (n_20818), .A1 (n_20180), .B0 (sa32[0] ), .Y(n_21693));
NAND2X1 g60247(.A (n_21079), .B (n_21687), .Y (n_21688));
NAND2X1 g60248(.A (n_21073), .B (n_22372), .Y (n_21686));
OAI21X1 g60296(.A0 (n_20978), .A1 (n_12322), .B0 (n_19414), .Y(n_21684));
NAND4X1 g60306(.A (n_20351), .B (n_15652), .C (n_20575), .D(n_18703), .Y (n_21683));
NAND4X1 g60307(.A (n_19937), .B (n_17219), .C (n_20562), .D(n_17601), .Y (n_21682));
NAND3X1 g60310(.A (n_20952), .B (n_20660), .C (n_19339), .Y(n_21681));
NAND3X1 g60311(.A (n_20743), .B (n_20651), .C (n_19897), .Y(n_21680));
NOR3X1 g60318(.A (n_16112), .B (n_20615), .C (n_20982), .Y (n_21678));
NAND3X1 g60328(.A (n_11182), .B (n_20664), .C (n_18665), .Y(n_21677));
NAND4X1 g60339(.A (n_25584), .B (n_15232), .C (n_25585), .D(n_13603), .Y (n_21676));
NAND2X1 g60344(.A (n_21067), .B (n_22301), .Y (n_21675));
NAND4X1 g60353(.A (n_19476), .B (n_15321), .C (n_20548), .D(n_11575), .Y (n_29197));
NAND3X1 g60359(.A (n_11092), .B (n_20654), .C (n_18660), .Y(n_21671));
NAND4X1 g60367(.A (n_25640), .B (n_16695), .C (n_25641), .D(n_15397), .Y (n_21668));
NAND4X1 g60371(.A (n_19487), .B (n_18835), .C (n_20555), .D(n_15396), .Y (n_21666));
NAND4X1 g60372(.A (n_18866), .B (n_19062), .C (n_20552), .D(n_19914), .Y (n_21665));
AND2X1 g60378(.A (n_21068), .B (n_15014), .Y (n_21663));
NAND4X1 g60411(.A (n_16905), .B (n_20972), .C (n_20634), .D(n_14754), .Y (n_21662));
NAND4X1 g60414(.A (n_21660), .B (n_20974), .C (n_21659), .D(n_11419), .Y (n_21661));
AOI21X1 g60418(.A0 (n_20981), .A1 (n_20182), .B0 (sa33[0] ), .Y(n_21658));
NAND2X1 g60420(.A (n_18300), .B (n_21075), .Y (n_21657));
AOI22X1 g60429(.A0 (n_20638), .A1 (w3[1] ), .B0 (n_18113), .B1(n_19433), .Y (n_21656));
NAND4X1 g60452(.A (n_18406), .B (n_20668), .C (n_20476), .D(n_13435), .Y (n_21655));
NAND4X1 g60461(.A (n_28315), .B (n_28316), .C (n_20027), .D(n_14778), .Y (n_21651));
OAI21X1 g60478(.A0 (n_20925), .A1 (n_18900), .B0 (n_26535), .Y(n_21648));
OAI21X1 g60479(.A0 (n_20924), .A1 (n_15811), .B0 (n_1196), .Y(n_21647));
OAI21X1 g60490(.A0 (n_20905), .A1 (n_18164), .B0 (n_1008), .Y(n_21642));
OAI21X1 g60494(.A0 (n_20900), .A1 (n_26704), .B0 (n_21174), .Y(n_21638));
OAI21X1 g60497(.A0 (n_20898), .A1 (n_15670), .B0 (n_2909), .Y(n_21637));
NAND2X1 g60501(.A (n_20989), .B (n_19414), .Y (n_21635));
NAND2X1 g60502(.A (n_21005), .B (n_27910), .Y (n_21634));
NOR2X1 g60509(.A (n_21037), .B (n_19704), .Y (n_21632));
NAND3X1 g60512(.A (n_15496), .B (n_20858), .C (n_20448), .Y(n_21631));
NOR2X1 g60517(.A (n_20993), .B (n_18538), .Y (n_21630));
NAND4X1 g60529(.A (n_20326), .B (n_20781), .C (n_13572), .D(n_20066), .Y (n_21629));
OAI21X1 g60543(.A0 (n_20939), .A1 (n_20095), .B0 (n_26844), .Y(n_21627));
AND2X1 g60545(.A (n_21249), .B (n_17444), .Y (n_21626));
NOR3X1 g60550(.A (n_17908), .B (n_12771), .C (n_20890), .Y (n_21625));
AOI21X1 g60554(.A0 (n_20838), .A1 (n_15244), .B0 (n_1699), .Y(n_21624));
AOI21X1 g60557(.A0 (n_20927), .A1 (n_18836), .B0 (n_21581), .Y(n_21623));
AOI21X1 g60558(.A0 (n_20837), .A1 (n_15329), .B0 (n_20632), .Y(n_21622));
OAI21X1 g60567(.A0 (n_20852), .A1 (n_19058), .B0 (n_1196), .Y(n_21620));
NAND2X1 g60568(.A (n_21272), .B (sa22[1] ), .Y (n_21618));
AOI21X1 g60582(.A0 (n_20911), .A1 (n_16701), .B0 (n_15766), .Y(n_21616));
NAND2X1 g60589(.A (n_21270), .B (n_903), .Y (n_21615));
NAND2X1 g60591(.A (n_21269), .B (n_20610), .Y (n_21614));
OAI21X1 g60593(.A0 (n_20850), .A1 (n_19689), .B0 (n_21174), .Y(n_21613));
OAI21X1 g60597(.A0 (n_20849), .A1 (n_19055), .B0 (n_1008), .Y(n_21611));
NAND3X1 g60603(.A (n_19707), .B (n_20809), .C (n_20902), .Y(n_21609));
NAND3X1 g60604(.A (n_20247), .B (n_20508), .C (n_20899), .Y(n_21608));
NAND4X1 g60607(.A (n_20637), .B (n_19232), .C (n_20515), .D (n_9426),.Y (n_21607));
NAND4X1 g60608(.A (n_20633), .B (n_19819), .C (n_20513), .D (n_9466),.Y (n_21606));
NAND4X1 g60624(.A (n_20467), .B (n_20860), .C (n_20360), .D(n_13732), .Y (n_21605));
AOI21X1 g60627(.A0 (n_20363), .A1 (w3[9] ), .B0 (n_20991), .Y(n_21604));
AOI21X1 g60628(.A0 (n_19429), .A1 (w3[9] ), .B0 (n_21027), .Y(n_21603));
AOI21X1 g60630(.A0 (n_19956), .A1 (n_1558), .B0 (n_21024), .Y(n_21601));
AOI21X1 g60632(.A0 (n_7031), .A1 (n_21598), .B0 (n_20990), .Y(n_21599));
OAI21X1 g60639(.A0 (n_27218), .A1 (n_20189), .B0 (n_27526), .Y(n_21597));
NAND4X1 g60654(.A (n_19669), .B (n_16703), .C (n_20482), .D(n_15399), .Y (n_21594));
OAI21X1 g60659(.A0 (n_20819), .A1 (n_20187), .B0 (n_28179), .Y(n_21593));
NAND2X1 g60684(.A (n_21040), .B (n_20202), .Y (n_21587));
NAND2X1 g60688(.A (n_21053), .B (n_20346), .Y (n_21586));
AOI22X1 g60690(.A0 (n_20854), .A1 (n_933), .B0 (n_9457), .B1(n_20010), .Y (n_21585));
NOR3X1 g60691(.A (n_17285), .B (n_19870), .C (n_20957), .Y (n_29123));
NOR3X1 g60692(.A (n_18363), .B (n_20317), .C (n_20956), .Y (n_21583));
NOR3X1 g60701(.A (n_18999), .B (n_19838), .C (n_20953), .Y (n_21579));
NOR3X1 g60702(.A (n_17208), .B (n_19835), .C (n_20719), .Y (n_25833));
NOR3X1 g60703(.A (n_18994), .B (n_20312), .C (n_20744), .Y (n_21577));
AOI22X1 g60705(.A0 (n_20834), .A1 (n_15766), .B0 (n_11346), .B1(n_18456), .Y (n_21576));
AOI22X1 g60709(.A0 (n_20833), .A1 (n_2681), .B0 (n_17669), .B1(n_29039), .Y (n_21574));
AOI22X1 g60710(.A0 (n_20831), .A1 (n_26903), .B0 (n_11281), .B1(n_290), .Y (n_21573));
AOI22X1 g60712(.A0 (n_20830), .A1 (n_21275), .B0 (n_11305), .B1(n_1295), .Y (n_21571));
AOI22X1 g60713(.A0 (n_26730), .A1 (n_21569), .B0 (n_13830), .B1(n_28631), .Y (n_21570));
AOI22X1 g60714(.A0 (n_20828), .A1 (n_21174), .B0 (n_19844), .B1(n_1310), .Y (n_21568));
NAND4X1 g60718(.A (n_21222), .B (n_17113), .C (n_15691), .D(n_18702), .Y (n_21567));
NAND4X1 g60719(.A (n_21217), .B (n_15583), .C (n_15677), .D(n_19436), .Y (n_21566));
AOI22X1 g60724(.A0 (n_27143), .A1 (n_20564), .B0 (n_18066), .B1(n_20332), .Y (n_21563));
AOI22X1 g60729(.A0 (n_20851), .A1 (n_3538), .B0 (n_18054), .B1(n_21396), .Y (n_21558));
INVX1 g60737(.A (n_21341), .Y (n_25453));
OAI21X1 g60745(.A0 (n_20005), .A1 (n_20806), .B0 (n_21552), .Y(n_21553));
NAND3X1 g60749(.A (n_28501), .B (n_18535), .C (n_28502), .Y(n_21550));
AOI21X1 g60750(.A0 (n_14210), .A1 (n_20771), .B0 (n_20157), .Y(n_21549));
NAND2X1 g60763(.A (n_21181), .B (n_2978), .Y (n_21540));
INVX1 g60788(.A (n_21328), .Y (n_21538));
NAND2X1 g60809(.A (n_21152), .B (n_15053), .Y (n_21535));
AOI21X1 g60812(.A0 (n_17547), .A1 (n_13575), .B0 (n_21147), .Y(n_21533));
NAND2X1 g60813(.A (n_28061), .B (n_15114), .Y (n_21532));
NAND2X1 g60815(.A (n_21140), .B (n_15027), .Y (n_21530));
AND2X1 g60826(.A (n_21211), .B (n_21174), .Y (n_21526));
NAND3X1 g60827(.A (n_21132), .B (n_19969), .C (n_18002), .Y(n_21524));
NAND3X1 g60838(.A (n_21131), .B (n_19438), .C (n_18842), .Y(n_21519));
NAND3X1 g60839(.A (n_21130), .B (n_17584), .C (n_18834), .Y(n_21518));
INVX1 g60845(.A (n_21315), .Y (n_21517));
NOR2X1 g60848(.A (n_29429), .B (n_29428), .Y (n_21516));
NAND3X1 g60853(.A (n_28269), .B (n_14762), .C (n_28270), .Y(n_21513));
NOR2X1 g60855(.A (n_16140), .B (n_21241), .Y (n_29195));
NAND2X1 g60875(.A (n_21150), .B (n_16362), .Y (n_21511));
NAND2X1 g60877(.A (n_21159), .B (n_19446), .Y (n_21509));
NAND4X1 g60896(.A (n_20071), .B (n_20784), .C (n_21164), .D(n_14739), .Y (n_21506));
NAND2X1 g60898(.A (n_21158), .B (n_19987), .Y (n_21505));
NAND3X1 g60905(.A (n_19825), .B (n_14763), .C (n_20798), .Y(n_21504));
NAND2X1 g60924(.A (n_21142), .B (n_903), .Y (n_21501));
OAI21X1 g60926(.A0 (n_20805), .A1 (sa11[1] ), .B0 (n_19158), .Y(n_21499));
NAND2X1 g60946(.A (n_19751), .B (n_21172), .Y (n_21498));
NOR2X1 g60952(.A (n_14527), .B (n_21236), .Y (n_25666));
NOR2X1 g60957(.A (n_14235), .B (n_21235), .Y (n_25598));
AOI21X1 g60961(.A0 (n_11508), .A1 (n_16466), .B0 (n_21247), .Y(n_21495));
AOI21X1 g60992(.A0 (n_20361), .A1 (n_869), .B0 (n_21180), .Y(n_21494));
NAND3X1 g60996(.A (n_20919), .B (n_19982), .C (n_18340), .Y(n_21493));
OAI21X1 g60997(.A0 (n_20494), .A1 (n_11206), .B0 (n_20767), .Y(n_21492));
AOI21X1 g61018(.A0 (n_20353), .A1 (n_20102), .B0 (n_19850), .Y(n_21486));
AOI21X1 g61019(.A0 (n_20365), .A1 (n_1196), .B0 (n_20951), .Y(n_21485));
AOI21X1 g61020(.A0 (n_20364), .A1 (n_21569), .B0 (n_20949), .Y(n_21484));
NAND4X1 g61031(.A (n_28253), .B (n_12873), .C (n_28254), .D(n_14475), .Y (n_21481));
AOI22X1 g61037(.A0 (n_20431), .A1 (n_3538), .B0 (n_11764), .B1(n_19750), .Y (n_21479));
NOR2X1 g61051(.A (n_15337), .B (n_20932), .Y (n_21478));
AOI21X1 g61053(.A0 (n_16420), .A1 (n_19310), .B0 (n_20958), .Y(n_21477));
AOI21X1 g61066(.A0 (n_18920), .A1 (n_20010), .B0 (n_20867), .Y(n_21476));
NAND4X1 g61067(.A (n_12741), .B (n_18675), .C (n_8465), .D (n_19731),.Y (n_21475));
NAND4X1 g61068(.A (n_12714), .B (n_19920), .C (n_12673), .D(n_19730), .Y (n_21474));
NAND4X1 g61075(.A (n_20734), .B (n_12668), .C (n_18580), .D (n_8192),.Y (n_21473));
AOI21X1 g61079(.A0 (n_18053), .A1 (n_14627), .B0 (n_20903), .Y(n_21472));
NAND4X1 g61080(.A (n_25719), .B (n_19735), .C (n_25720), .D(n_10193), .Y (n_21471));
NAND4X1 g61082(.A (n_11827), .B (n_16810), .C (n_18849), .D(n_19719), .Y (n_21470));
AOI22X1 g61083(.A0 (n_20408), .A1 (n_17444), .B0 (n_19165), .B1(n_196), .Y (n_21469));
NAND4X1 g61084(.A (n_8610), .B (n_13058), .C (n_18010), .D (n_19718),.Y (n_21467));
NAND4X1 g61089(.A (n_25467), .B (n_25468), .C (n_19376), .D (n_9802),.Y (n_21465));
NOR2X1 g61090(.A (n_17593), .B (n_20879), .Y (n_21464));
OAI21X1 g61091(.A0 (n_20405), .A1 (n_19319), .B0 (n_20550), .Y(n_21463));
NAND4X1 g61096(.A (n_17991), .B (n_16817), .C (n_19747), .D(n_11156), .Y (n_21462));
NAND4X1 g61097(.A (n_16596), .B (n_16092), .C (n_19746), .D(n_12485), .Y (n_21461));
OAI21X1 g61099(.A0 (n_27784), .A1 (n_20041), .B0 (n_19945), .Y(n_21460));
NAND4X1 g61244(.A (n_27238), .B (n_16411), .C (n_19638), .D(n_19671), .Y (n_21458));
OAI21X1 g61305(.A0 (n_20302), .A1 (n_21055), .B0 (n_19886), .Y(n_21455));
INVX1 g61327(.A (n_21189), .Y (n_21454));
OAI21X1 g61370(.A0 (n_20294), .A1 (n_19908), .B0 (n_14859), .Y(n_21452));
OAI21X1 g61372(.A0 (n_20292), .A1 (n_124), .B0 (n_13212), .Y(n_21451));
OAI21X1 g61375(.A0 (n_20297), .A1 (n_933), .B0 (n_17768), .Y(n_21450));
OAI21X1 g61380(.A0 (n_20259), .A1 (n_10323), .B0 (n_21447), .Y(n_25591));
OAI21X1 g61385(.A0 (n_20306), .A1 (n_17337), .B0 (n_27449), .Y(n_21446));
OAI21X1 g61388(.A0 (n_20301), .A1 (n_487), .B0 (n_18103), .Y(n_21445));
OAI21X1 g61396(.A0 (n_20288), .A1 (n_28170), .B0 (n_18088), .Y(n_21439));
OAI21X1 g61397(.A0 (n_20287), .A1 (sa21[1] ), .B0 (n_19626), .Y(n_21438));
NOR3X1 g61409(.A (n_17261), .B (n_8109), .C (n_20266), .Y (n_21437));
NAND3X1 g61413(.A (n_6167), .B (n_20334), .C (n_19842), .Y (n_21436));
NOR3X1 g61415(.A (n_17179), .B (n_9698), .C (n_20265), .Y (n_21435));
NOR3X1 g61418(.A (n_17172), .B (n_8104), .C (n_20263), .Y (n_21434));
AOI21X1 g61437(.A0 (n_19793), .A1 (n_663), .B0 (n_20785), .Y(n_21433));
OAI21X1 g61439(.A0 (n_18522), .A1 (n_487), .B0 (n_27448), .Y(n_21432));
OAI21X1 g61443(.A0 (n_19126), .A1 (n_20758), .B0 (n_20811), .Y(n_21431));
AOI22X1 g61446(.A0 (n_20279), .A1 (sa23[1] ), .B0 (n_18521), .B1(n_164), .Y (n_21430));
AOI22X1 g61456(.A0 (n_27311), .A1 (n_20564), .B0 (n_8638), .B1(n_19157), .Y (n_21429));
NAND2X1 g61477(.A (n_16104), .B (n_20803), .Y (n_21427));
AOI21X1 g61495(.A0 (n_20303), .A1 (n_21188), .B0 (n_20337), .Y(n_21426));
OAI21X1 g61601(.A0 (n_25580), .A1 (n_25581), .B0 (n_20579), .Y(n_21423));
OAI21X1 g61655(.A0 (n_16578), .A1 (n_20236), .B0 (n_20564), .Y(n_21422));
AND2X1 g61901(.A (n_20229), .B (n_20723), .Y (n_21420));
NOR2X1 g62434(.A (n_20685), .B (n_18853), .Y (n_21419));
NAND4X1 g60130(.A (n_28850), .B (n_28851), .C (n_28161), .D(n_18182), .Y (n_21417));
NAND4X1 g60140(.A (n_25710), .B (n_25711), .C (n_20628), .D(n_17088), .Y (n_21416));
NAND3X1 g60252(.A (n_20344), .B (n_20205), .C (n_19312), .Y(n_21413));
NAND3X1 g60257(.A (n_19941), .B (n_20200), .C (n_19282), .Y(n_21412));
NAND3X1 g60261(.A (n_20340), .B (n_20199), .C (n_19275), .Y(n_21411));
NAND3X1 g60262(.A (n_19391), .B (n_20197), .C (n_17511), .Y(n_21410));
OAI21X1 g60282(.A0 (n_20623), .A1 (n_8849), .B0 (n_20397), .Y(n_21409));
OAI21X1 g60287(.A0 (n_20622), .A1 (n_8085), .B0 (n_20386), .Y(n_25690));
NAND3X1 g60312(.A (n_17442), .B (n_20191), .C (n_17578), .Y(n_21406));
OAI21X1 g60323(.A0 (n_20625), .A1 (n_16719), .B0 (n_196), .Y(n_21405));
AOI22X1 g60450(.A0 (n_20619), .A1 (n_1558), .B0 (n_4048), .B1(n_14017), .Y (n_21404));
OAI21X1 g60480(.A0 (n_20583), .A1 (n_16078), .B0 (n_21447), .Y(n_21400));
OAI21X1 g60485(.A0 (n_20568), .A1 (n_16017), .B0 (n_21398), .Y(n_21399));
OAI21X1 g60486(.A0 (n_20566), .A1 (n_14327), .B0 (n_21396), .Y(n_28882));
AND2X1 g60487(.A (n_20988), .B (n_21442), .Y (n_21395));
NAND2X1 g60504(.A (n_20684), .B (n_17445), .Y (n_21393));
NAND4X1 g60507(.A (n_17424), .B (n_19411), .C (n_20118), .D(n_16481), .Y (n_21392));
NAND4X1 g60520(.A (n_29414), .B (n_29415), .C (n_18009), .D(n_20107), .Y (n_21391));
NAND4X1 g60521(.A (n_18668), .B (n_19551), .C (n_16863), .D(n_20103), .Y (n_21390));
NAND4X1 g60530(.A (n_19342), .B (n_20443), .C (n_17951), .D(n_20054), .Y (n_21389));
NAND4X1 g60533(.A (n_19893), .B (n_19473), .C (n_16549), .D(n_20029), .Y (n_21388));
NAND2X1 g60555(.A (n_20980), .B (n_804), .Y (n_21386));
NAND4X1 g60574(.A (n_20289), .B (n_12231), .C (n_19367), .D(n_20056), .Y (n_21384));
NAND2X1 g60576(.A (n_20985), .B (n_21382), .Y (n_21383));
NAND2X1 g60578(.A (n_20979), .B (n_788), .Y (n_21381));
NAND4X1 g60586(.A (n_25734), .B (n_15781), .C (n_20045), .D(n_25735), .Y (n_21379));
NAND3X1 g60602(.A (n_20250), .B (n_20132), .C (n_20581), .Y(n_28284));
NAND3X1 g60605(.A (n_20246), .B (n_20128), .C (n_20549), .Y(n_21376));
NAND3X1 g60606(.A (n_19686), .B (n_16002), .C (n_20593), .Y(n_21375));
NAND4X1 g60609(.A (n_20921), .B (n_19868), .C (n_18686), .D(n_19309), .Y (n_21374));
NAND4X1 g60610(.A (n_19607), .B (n_19230), .C (n_20143), .D(n_11384), .Y (n_21373));
NAND3X1 g60612(.A (n_19673), .B (n_14366), .C (n_20572), .Y(n_21372));
NAND3X1 g60613(.A (n_18319), .B (n_14262), .C (n_20557), .Y(n_22709));
NAND4X1 g60619(.A (n_18402), .B (n_9569), .C (n_20121), .D (n_11587),.Y (n_21371));
NAND4X1 g60620(.A (n_20237), .B (n_9586), .C (n_20120), .D (n_13594),.Y (n_21370));
NAND4X1 g60621(.A (n_18399), .B (n_15301), .C (n_20119), .D(n_13616), .Y (n_21369));
NAND4X1 g60625(.A (n_15277), .B (n_17306), .C (n_20016), .D(n_15300), .Y (n_21368));
NAND4X1 g60626(.A (n_19664), .B (n_11519), .C (n_20117), .D(n_15431), .Y (n_28283));
AOI21X1 g60633(.A0 (n_20362), .A1 (n_20632), .B0 (n_20635), .Y(n_21366));
AOI21X1 g60634(.A0 (n_19954), .A1 (w3[17] ), .B0 (n_20659), .Y(n_21364));
NAND4X1 g60635(.A (n_18365), .B (n_20078), .C (n_13465), .D(n_20152), .Y (n_21363));
NAND3X1 g60636(.A (n_17162), .B (n_20523), .C (n_9572), .Y (n_21362));
AOI21X1 g60641(.A0 (n_20519), .A1 (n_19722), .B0 (n_21), .Y(n_21361));
NAND4X1 g60644(.A (n_18969), .B (n_17846), .C (n_20110), .D(n_13582), .Y (n_21360));
NAND4X1 g60650(.A (n_17215), .B (n_17934), .C (n_20113), .D(n_11581), .Y (n_21358));
NAND4X1 g60651(.A (n_28893), .B (n_11460), .C (n_28894), .D(n_15400), .Y (n_21357));
OAI21X1 g60656(.A0 (n_20516), .A1 (n_20188), .B0 (n_0), .Y (n_21356));
NAND4X1 g60668(.A (n_17175), .B (n_13290), .C (n_20112), .D(n_11578), .Y (n_21355));
NAND4X1 g60670(.A (n_18277), .B (n_17865), .C (n_20111), .D(n_15389), .Y (n_21354));
NAND4X1 g60685(.A (n_19354), .B (n_11083), .C (n_19727), .D(n_19517), .Y (n_21353));
AOI22X1 g60689(.A0 (n_20527), .A1 (n_196), .B0 (n_14621), .B1(n_19433), .Y (n_21352));
AOI22X1 g60698(.A0 (n_20522), .A1 (n_1196), .B0 (n_19862), .B1(n_19651), .Y (n_21350));
AOI22X1 g60706(.A0 (n_20521), .A1 (n_20729), .B0 (n_20567), .B1(n_624), .Y (n_21349));
AOI22X1 g60711(.A0 (n_20520), .A1 (n_20102), .B0 (n_11227), .B1(n_3910), .Y (n_21348));
NAND2X1 g60715(.A (n_20683), .B (n_19925), .Y (n_21346));
NOR2X1 g60731(.A (n_18231), .B (n_20941), .Y (n_21345));
NOR2X1 g60734(.A (n_13113), .B (n_20893), .Y (n_21343));
NOR2X1 g60736(.A (n_18215), .B (n_20938), .Y (n_21342));
NAND3X1 g60738(.A (n_18953), .B (n_20272), .C (n_20022), .Y(n_21341));
AOI21X1 g60739(.A0 (n_11699), .A1 (n_16466), .B0 (n_20891), .Y(n_21340));
NAND3X1 g60746(.A (n_17798), .B (n_18890), .C (n_20398), .Y(n_21339));
NAND3X1 g60762(.A (n_29367), .B (n_19150), .C (n_29368), .Y(n_21333));
NAND2X1 g60769(.A (n_20865), .B (n_20018), .Y (n_21332));
NAND2X1 g60772(.A (n_20864), .B (n_14630), .Y (n_21331));
OAI21X1 g60773(.A0 (n_20439), .A1 (n_12516), .B0 (n_27242), .Y(n_25717));
OAI21X1 g60775(.A0 (n_20437), .A1 (n_15999), .B0 (n_21396), .Y(n_21329));
NAND2X1 g60789(.A (n_20894), .B (n_21382), .Y (n_21328));
OAI21X1 g60801(.A0 (n_20352), .A1 (n_12330), .B0 (n_21275), .Y(n_21327));
OAI21X1 g60823(.A0 (n_20478), .A1 (n_19559), .B0 (n_20767), .Y(n_21326));
OAI21X1 g60825(.A0 (n_20466), .A1 (n_19558), .B0 (n_20068), .Y(n_21323));
NOR2X1 g60832(.A (n_20821), .B (n_20609), .Y (n_21320));
NAND3X1 g60841(.A (n_20608), .B (n_19996), .C (n_20511), .Y(n_21317));
NOR2X1 g60843(.A (n_20816), .B (n_20607), .Y (n_21316));
OAI21X1 g60846(.A0 (n_20383), .A1 (n_15387), .B0 (n_21314), .Y(n_21315));
NAND4X1 g60858(.A (n_20794), .B (n_19885), .C (n_16864), .D(n_17814), .Y (n_21312));
OAI21X1 g60868(.A0 (n_20463), .A1 (n_14434), .B0 (sa20[1] ), .Y(n_25809));
NOR3X1 g60881(.A (n_17421), .B (n_19921), .C (n_20456), .Y (n_21308));
NAND4X1 g60890(.A (n_20077), .B (n_20455), .C (n_16084), .D(n_14743), .Y (n_21307));
OAI21X1 g60893(.A0 (n_20500), .A1 (n_804), .B0 (n_19159), .Y(n_21306));
AOI22X1 g60899(.A0 (n_20452), .A1 (n_196), .B0 (n_7822), .B1(n_14142), .Y (n_21304));
AOI22X1 g60901(.A0 (n_20450), .A1 (n_5131), .B0 (n_11672), .B1(n_18266), .Y (n_21303));
NOR2X1 g60904(.A (n_14420), .B (n_20964), .Y (n_25706));
NOR2X1 g60908(.A (n_12586), .B (n_20962), .Y (n_21300));
NOR3X1 g60930(.A (n_17418), .B (n_19375), .C (n_20432), .Y (n_21298));
NAND4X1 g60956(.A (n_14928), .B (n_19173), .C (n_11887), .D(n_19759), .Y (n_21297));
AOI21X1 g60964(.A0 (n_13420), .A1 (n_4582), .B0 (n_20968), .Y(n_21295));
NAND3X1 g60965(.A (n_20248), .B (n_19918), .C (n_20441), .Y(n_21294));
AOI21X1 g60966(.A0 (n_14901), .A1 (n_13466), .B0 (n_20969), .Y(n_21293));
NAND4X1 g60973(.A (n_20735), .B (n_20335), .C (n_13324), .D(n_19100), .Y (n_21292));
AOI21X1 g60978(.A0 (n_20471), .A1 (n_21290), .B0 (n_1558), .Y(n_21291));
NAND4X1 g60984(.A (n_15667), .B (n_20003), .C (n_19877), .D(n_17530), .Y (n_21289));
NOR2X1 g60985(.A (n_20866), .B (n_19315), .Y (n_21288));
AOI21X1 g60989(.A0 (n_20403), .A1 (n_3264), .B0 (n_19198), .Y(n_21286));
AOI21X1 g60991(.A0 (n_20401), .A1 (n_124), .B0 (n_19790), .Y(n_21284));
NAND4X1 g60995(.A (n_14007), .B (n_19450), .C (n_19284), .D(n_19285), .Y (n_21283));
NAND3X1 g61007(.A (n_20591), .B (n_19990), .C (n_18377), .Y(n_21279));
AOI21X1 g61015(.A0 (n_19959), .A1 (n_21055), .B0 (n_19321), .Y(n_21278));
AOI21X1 g61017(.A0 (n_19958), .A1 (n_21275), .B0 (n_19287), .Y(n_21276));
AOI22X1 g61025(.A0 (n_19998), .A1 (sa21[1] ), .B0 (n_19151), .B1(n_27910), .Y (n_21274));
NAND4X1 g61032(.A (n_20061), .B (n_15161), .C (n_19368), .D(n_15891), .Y (n_21273));
NAND4X1 g61033(.A (n_17970), .B (n_16772), .C (n_19196), .D(n_15916), .Y (n_21272));
NAND4X1 g61039(.A (n_28275), .B (n_14635), .C (n_19181), .D(n_28276), .Y (n_21271));
NAND4X1 g61040(.A (n_25589), .B (n_12678), .C (n_25590), .D(n_14217), .Y (n_21270));
NAND4X1 g61041(.A (n_25810), .B (n_14354), .C (n_25811), .D(n_14473), .Y (n_21269));
NAND4X1 g61045(.A (n_19212), .B (n_16265), .C (n_19410), .D(n_15822), .Y (n_21268));
AOI21X1 g61046(.A0 (n_16496), .A1 (n_19445), .B0 (n_20606), .Y(n_21267));
NAND4X1 g61047(.A (n_28581), .B (n_11040), .C (n_28582), .D (n_8844),.Y (n_21266));
NAND4X1 g61048(.A (n_17489), .B (n_16076), .C (n_19407), .D(n_12079), .Y (n_21265));
NAND4X1 g61050(.A (n_19208), .B (n_14708), .C (n_19406), .D(n_15833), .Y (n_21264));
NOR2X1 g61054(.A (n_17875), .B (n_20584), .Y (n_21263));
AOI21X1 g61055(.A0 (n_16491), .A1 (n_1132), .B0 (n_20605), .Y(n_21262));
NOR2X1 g61056(.A (n_16777), .B (n_20576), .Y (n_21261));
NAND4X1 g61057(.A (n_28320), .B (n_10870), .C (n_28321), .D (n_7407),.Y (n_21260));
NAND4X1 g61058(.A (n_17485), .B (n_12404), .C (n_19384), .D(n_13896), .Y (n_21259));
NAND4X1 g61060(.A (n_19192), .B (n_14672), .C (n_19397), .D(n_15824), .Y (n_21258));
NAND4X1 g61062(.A (n_25617), .B (n_10873), .C (n_25618), .D(n_10294), .Y (n_21257));
NAND4X1 g61064(.A (n_25487), .B (n_12429), .C (n_19386), .D(n_25488), .Y (n_21256));
NOR2X1 g61071(.A (n_19416), .B (n_20596), .Y (n_21254));
NOR2X1 g61078(.A (n_19938), .B (n_20563), .Y (n_21252));
AOI22X1 g61092(.A0 (n_20012), .A1 (n_4357), .B0 (n_20084), .B1(n_21552), .Y (n_29395));
NAND4X1 g61095(.A (n_15209), .B (n_11204), .C (n_19147), .D(n_10833), .Y (n_21249));
OAI21X1 g61107(.A0 (n_19815), .A1 (n_14435), .B0 (n_1196), .Y(n_21248));
OAI21X1 g61108(.A0 (n_19873), .A1 (n_20153), .B0 (n_20295), .Y(n_21247));
OAI21X1 g61112(.A0 (n_19812), .A1 (n_17604), .B0 (n_21174), .Y(n_21246));
OAI21X1 g61114(.A0 (n_19808), .A1 (n_14477), .B0 (n_21242), .Y(n_21243));
AOI21X1 g61115(.A0 (n_14893), .A1 (n_19721), .B0 (n_21188), .Y(n_21241));
INVX1 g61116(.A (n_20967), .Y (n_21240));
INVX1 g61119(.A (n_20966), .Y (n_21239));
INVX1 g61121(.A (n_20965), .Y (n_21238));
AOI21X1 g61128(.A0 (n_13939), .A1 (n_19716), .B0 (n_20412), .Y(n_21236));
AOI21X1 g61129(.A0 (n_13250), .A1 (n_19715), .B0 (n_20068), .Y(n_21235));
NOR3X1 g61148(.A (n_20535), .B (n_13362), .C (n_19839), .Y (n_21233));
AOI22X1 g61163(.A0 (n_19829), .A1 (n_11277), .B0 (n_15960), .B1(n_673), .Y (n_21230));
AOI22X1 g61164(.A0 (n_19828), .A1 (n_20325), .B0 (n_17591), .B1(n_477), .Y (n_21229));
NAND4X1 g61171(.A (n_21227), .B (n_15830), .C (n_18941), .D(n_19038), .Y (n_21228));
INVX1 g61192(.A (n_20937), .Y (n_21225));
NAND2X1 g61201(.A (n_20461), .B (w3[9] ), .Y (n_21222));
AOI21X1 g61205(.A0 (n_19878), .A1 (n_17906), .B0 (n_21174), .Y(n_21220));
NAND3X1 g61213(.A (n_25837), .B (n_17525), .C (n_25838), .Y(n_21219));
NAND2X1 g61214(.A (n_20454), .B (sa22[1] ), .Y (n_21218));
NAND2X1 g61215(.A (n_20451), .B (n_19532), .Y (n_21217));
NAND4X1 g61216(.A (n_21215), .B (n_16435), .C (n_18948), .D(n_19018), .Y (n_21216));
NOR3X1 g61228(.A (n_20239), .B (n_17704), .C (n_19864), .Y (n_21214));
NAND4X1 g61234(.A (n_21210), .B (n_16432), .C (n_18926), .D(n_19027), .Y (n_21211));
NAND3X1 g61237(.A (n_29310), .B (n_17217), .C (n_19860), .Y(n_21209));
INVX1 g61238(.A (n_20918), .Y (n_21208));
NAND2X1 g61251(.A (n_20442), .B (n_788), .Y (n_21207));
NAND3X1 g61264(.A (n_15035), .B (n_17516), .C (n_19836), .Y(n_21205));
INVX1 g61272(.A (n_20906), .Y (n_21202));
NAND3X1 g61279(.A (n_16671), .B (n_17514), .C (n_19833), .Y(n_21201));
NAND2X1 g61283(.A (n_20426), .B (n_3538), .Y (n_21200));
NOR3X1 g61293(.A (n_28138), .B (n_16329), .C (n_19827), .Y (n_21197));
NAND2X1 g61300(.A (n_20268), .B (n_20382), .Y (n_21196));
AOI21X1 g61301(.A0 (n_19823), .A1 (n_27801), .B0 (n_21314), .Y(n_21195));
NAND2X1 g61304(.A (n_20378), .B (n_19234), .Y (n_21194));
NOR2X1 g61308(.A (n_20505), .B (n_19732), .Y (n_28853));
OAI21X1 g61309(.A0 (n_19741), .A1 (n_17444), .B0 (n_18217), .Y(n_21192));
NOR2X1 g61320(.A (n_20496), .B (n_19726), .Y (n_21191));
AOI22X1 g61322(.A0 (n_19780), .A1 (sa22[1] ), .B0 (n_18184), .B1(n_6244), .Y (n_21190));
OAI21X1 g61328(.A0 (n_19740), .A1 (n_21188), .B0 (n_17580), .Y(n_21189));
AOI21X1 g61334(.A0 (n_10849), .A1 (n_19408), .B0 (n_20416), .Y(n_21187));
AOI21X1 g61335(.A0 (n_12721), .A1 (n_19398), .B0 (n_20411), .Y(n_21186));
NOR2X1 g61337(.A (n_20485), .B (n_20257), .Y (n_21185));
NAND4X1 g61339(.A (n_20339), .B (n_10801), .C (n_19092), .D(n_16020), .Y (n_21184));
NAND4X1 g61341(.A (n_20338), .B (n_28901), .C (n_19090), .D(n_16054), .Y (n_21183));
OR4X1 g61346(.A (n_16093), .B (n_10171), .C (n_17643), .D (n_18891),.Y (n_21181));
AOI21X1 g61354(.A0 (n_19866), .A1 (n_21659), .B0 (w3[1] ), .Y(n_21180));
NAND2X1 g61366(.A (n_20465), .B (n_1196), .Y (n_21179));
OAI21X1 g61371(.A0 (n_19738), .A1 (n_10605), .B0 (n_27449), .Y(n_21177));
NAND2X1 g61374(.A (n_20447), .B (n_21174), .Y (n_21175));
OAI21X1 g61378(.A0 (n_19737), .A1 (n_9041), .B0 (n_21275), .Y(n_21173));
OAI21X1 g61384(.A0 (n_19736), .A1 (n_8907), .B0 (n_2681), .Y(n_21172));
OAI21X1 g61403(.A0 (n_19760), .A1 (n_877), .B0 (n_20487), .Y(n_21169));
NAND2X1 g61404(.A (n_20049), .B (n_20400), .Y (n_21168));
NAND4X1 g61410(.A (n_18739), .B (n_21164), .C (n_15659), .D(n_19102), .Y (n_21165));
NAND4X1 g61417(.A (n_17842), .B (n_19019), .C (n_18964), .D (n_9505),.Y (n_21163));
NOR2X1 g61421(.A (n_19654), .B (n_20504), .Y (n_21162));
MX2X1 g61436(.A (n_19210), .B (n_19794), .S0 (n_933), .Y (n_21159));
MX2X1 g61440(.A (n_19788), .B (n_19764), .S0 (n_124), .Y (n_21158));
OAI21X1 g61441(.A0 (n_19127), .A1 (n_20767), .B0 (n_20509), .Y(n_21157));
AOI22X1 g61444(.A0 (n_19773), .A1 (n_778), .B0 (n_17443), .B1(n_177), .Y (n_21156));
AOI22X1 g61445(.A0 (n_19771), .A1 (sa32[1] ), .B0 (n_17457), .B1(n_1397), .Y (n_21155));
AOI22X1 g61447(.A0 (n_19767), .A1 (n_20574), .B0 (n_19125), .B1(n_21275), .Y (n_21154));
AOI22X1 g61448(.A0 (n_19787), .A1 (sa20[1] ), .B0 (n_19739), .B1(n_21055), .Y (n_21153));
AOI22X1 g61451(.A0 (n_19710), .A1 (n_21151), .B0 (n_10209), .B1(n_19160), .Y (n_21152));
NAND4X1 g61453(.A (n_15248), .B (n_14709), .C (n_19026), .D(n_11342), .Y (n_21150));
INVX1 g61461(.A (n_20836), .Y (n_21149));
NOR2X1 g61465(.A (n_15185), .B (n_20453), .Y (n_21148));
NAND2X1 g61467(.A (n_16073), .B (n_20498), .Y (n_21147));
NAND4X1 g61468(.A (n_29321), .B (n_13946), .C (n_29322), .D(n_12955), .Y (n_21146));
NAND2X1 g61471(.A (n_16098), .B (n_20502), .Y (n_21145));
NAND4X1 g61473(.A (n_15079), .B (n_14679), .C (n_19004), .D(n_12966), .Y (n_21142));
NAND2X1 g61474(.A (n_16008), .B (n_20493), .Y (n_21141));
AOI22X1 g61475(.A0 (n_19712), .A1 (n_778), .B0 (n_10217), .B1(n_19152), .Y (n_21140));
NOR2X1 g61476(.A (n_16682), .B (n_20430), .Y (n_21139));
NAND4X1 g61488(.A (n_14919), .B (n_19071), .C (n_17406), .D(n_19557), .Y (n_21138));
AOI21X1 g61489(.A0 (n_19650), .A1 (n_21314), .B0 (n_20004), .Y(n_21137));
AOI21X1 g61490(.A0 (n_18907), .A1 (n_21396), .B0 (n_20394), .Y(n_21135));
AOI21X1 g61492(.A0 (n_19635), .A1 (n_21133), .B0 (n_20393), .Y(n_21134));
NOR2X1 g61493(.A (n_19922), .B (n_20458), .Y (n_21132));
NOR2X1 g61496(.A (n_19917), .B (n_20435), .Y (n_21131));
NOR2X1 g61498(.A (n_19915), .B (n_20429), .Y (n_21130));
OAI21X1 g61508(.A0 (n_19754), .A1 (n_19934), .B0 (n_19992), .Y(n_29428));
NAND3X1 g61559(.A (n_28505), .B (n_28506), .C (n_19010), .Y(n_21128));
NOR2X1 g61617(.A (n_15690), .B (n_20318), .Y (n_21127));
NAND2X1 g61662(.A (n_20304), .B (n_20153), .Y (n_21126));
INVX1 g61711(.A (n_20778), .Y (n_21125));
NOR2X1 g61714(.A (n_20260), .B (n_6672), .Y (n_21124));
OAI21X1 g61716(.A0 (n_19684), .A1 (n_21122), .B0 (n_27493), .Y(n_25456));
NAND4X1 g61156(.A (n_28586), .B (n_16606), .C (n_21120), .D(n_14544), .Y (n_21121));
OAI21X1 g61818(.A0 (n_16560), .A1 (n_19661), .B0 (n_21151), .Y(n_21119));
NOR2X1 g61819(.A (n_20258), .B (n_6449), .Y (n_21118));
AOI21X1 g61872(.A0 (n_19629), .A1 (n_17250), .B0 (n_19310), .Y(n_21116));
AND2X1 g61879(.A (n_19022), .B (n_20316), .Y (n_25686));
NAND3X1 g61885(.A (n_25546), .B (n_25547), .C (n_17046), .Y(n_21114));
AOI21X1 g61887(.A0 (n_14379), .A1 (n_20677), .B0 (n_20314), .Y(n_21113));
AOI21X1 g61926(.A0 (n_19632), .A1 (n_17303), .B0 (n_19445), .Y(n_21112));
NAND4X1 g61976(.A (n_16612), .B (n_19430), .C (n_19585), .D(n_12390), .Y (n_21110));
NOR2X1 g62432(.A (n_20219), .B (n_17961), .Y (n_21106));
INVX1 g62575(.A (n_20717), .Y (n_21104));
AOI22X1 g60430(.A0 (n_19610), .A1 (w3[9] ), .B0 (n_13682), .B1(n_20010), .Y (n_21101));
AOI22X1 g60447(.A0 (n_20190), .A1 (n_869), .B0 (n_19692), .B1(n_10139), .Y (n_21100));
NAND2X1 g60469(.A (n_20206), .B (n_171), .Y (n_21098));
OAI21X1 g60470(.A0 (n_20179), .A1 (n_16132), .B0 (n_27449), .Y(n_29405));
NAND2X1 g60499(.A (n_20193), .B (n_21133), .Y (n_25781));
NAND4X1 g60508(.A (n_17422), .B (n_19933), .C (n_17647), .D(n_16445), .Y (n_21095));
NAND4X1 g60510(.A (n_18511), .B (n_19932), .C (n_19554), .D(n_13140), .Y (n_21094));
NAND4X1 g60522(.A (n_19347), .B (n_18719), .C (n_19447), .D(n_15474), .Y (n_21093));
AOI22X1 g60549(.A0 (n_20177), .A1 (n_196), .B0 (n_9230), .B1(n_14142), .Y (n_21092));
AOI21X1 g60560(.A0 (n_9299), .A1 (n_13606), .B0 (n_20211), .Y(n_21087));
NAND2X1 g60590(.A (n_20627), .B (n_1397), .Y (n_21085));
AND2X1 g63776(.A (n_20618), .B (n_16835), .Y (n_21083));
NAND4X1 g60601(.A (n_20273), .B (n_12264), .C (n_19371), .D(n_19467), .Y (n_21082));
NAND3X1 g60611(.A (n_20616), .B (n_19301), .C (n_19400), .Y(n_21081));
NOR3X1 g60614(.A (n_19667), .B (n_19264), .C (n_20171), .Y (n_25700));
NAND3X1 g60623(.A (n_15706), .B (n_20156), .C (n_15293), .Y(n_21079));
NAND3X1 g60629(.A (n_17154), .B (n_20154), .C (n_11542), .Y(n_21078));
NAND4X1 g60642(.A (n_18263), .B (n_13344), .C (n_19553), .D(n_11577), .Y (n_21077));
NAND4X1 g60649(.A (n_17221), .B (n_11464), .C (n_19561), .D(n_15403), .Y (n_21076));
OAI21X1 g60660(.A0 (n_20148), .A1 (n_20186), .B0 (n_26844), .Y(n_21075));
NAND4X1 g60687(.A (n_20469), .B (n_20175), .C (n_18734), .D(n_11375), .Y (n_21073));
AOI22X1 g60695(.A0 (n_378), .A1 (n_28606), .B0 (n_20178), .B1(n_2981), .Y (n_21072));
NOR3X1 g60704(.A (n_17199), .B (n_19266), .C (n_20185), .Y (n_21071));
AOI21X1 g60707(.A0 (n_20150), .A1 (n_28169), .B0 (n_14204), .Y(n_21070));
AOI22X1 g60708(.A0 (n_20149), .A1 (n_20018), .B0 (n_20582), .B1(n_27128), .Y (n_21068));
NAND4X1 g60720(.A (n_20578), .B (n_16775), .C (n_15656), .D(n_18700), .Y (n_21067));
AOI22X1 g60722(.A0 (n_20161), .A1 (n_20841), .B0 (n_18069), .B1(n_20144), .Y (n_21066));
AOI22X1 g60725(.A0 (sa30[1] ), .A1 (n_28605), .B0 (n_18058), .B1(n_129), .Y (n_21065));
NAND2X1 g60735(.A (n_20528), .B (n_12788), .Y (n_21061));
NOR3X1 g60741(.A (n_14727), .B (n_17801), .C (n_20081), .Y (n_21060));
NAND2X1 g60764(.A (n_20541), .B (n_27449), .Y (n_21057));
NAND2X1 g60765(.A (n_20540), .B (n_21055), .Y (n_21056));
OAI21X1 g60767(.A0 (n_20097), .A1 (n_12804), .B0 (n_20397), .Y(n_21054));
NAND2X1 g60768(.A (n_20539), .B (n_1196), .Y (n_21053));
NAND2X1 g60770(.A (n_20534), .B (n_164), .Y (n_21052));
OAI21X1 g60771(.A0 (n_20063), .A1 (n_12348), .B0 (n_20386), .Y(n_21050));
NAND2X1 g60774(.A (n_20538), .B (n_20677), .Y (n_21049));
NAND2X1 g60776(.A (n_20537), .B (n_21242), .Y (n_21048));
NAND2X1 g60777(.A (n_20536), .B (n_21398), .Y (n_21047));
NAND2X1 g60778(.A (n_20533), .B (n_21275), .Y (n_21046));
NAND2X1 g60784(.A (n_20592), .B (n_20386), .Y (n_21043));
OAI21X1 g60790(.A0 (n_19950), .A1 (n_14394), .B0 (n_21242), .Y(n_21041));
NAND2X1 g60792(.A (n_20571), .B (n_1397), .Y (n_21040));
OAI21X1 g60799(.A0 (n_19948), .A1 (n_14154), .B0 (n_20102), .Y(n_21038));
OAI21X1 g60807(.A0 (n_18196), .A1 (w3[17] ), .B0 (n_20603), .Y(n_21037));
NAND3X1 g60817(.A (n_15296), .B (n_16894), .C (n_20133), .Y(n_21036));
NAND3X1 g60818(.A (n_16581), .B (n_11589), .C (n_20130), .Y(n_21035));
OAI21X1 g60831(.A0 (n_19508), .A1 (n_20126), .B0 (n_804), .Y(n_21034));
AOI22X1 g60850(.A0 (n_20104), .A1 (n_1196), .B0 (n_11668), .B1(n_19791), .Y (n_21031));
NAND2X1 g60862(.A (n_20532), .B (n_869), .Y (n_21029));
OAI21X1 g60866(.A0 (n_20089), .A1 (n_12767), .B0 (n_20412), .Y(n_28256));
OR2X1 g60867(.A (n_19800), .B (n_20530), .Y (n_21027));
OAI21X1 g60870(.A0 (n_20087), .A1 (n_9331), .B0 (n_19319), .Y(n_21025));
OR2X1 g60872(.A (n_19798), .B (n_20529), .Y (n_21024));
AOI22X1 g60876(.A0 (n_20083), .A1 (n_21174), .B0 (n_11661), .B1(n_16279), .Y (n_21023));
OAI21X1 g60884(.A0 (n_20002), .A1 (n_13640), .B0 (n_20198), .Y(n_21022));
OAI21X1 g60888(.A0 (n_20079), .A1 (n_11066), .B0 (w3[17] ), .Y(n_21020));
NAND2X1 g60889(.A (n_20525), .B (sa22[1] ), .Y (n_21018));
OAI21X1 g60891(.A0 (n_20074), .A1 (n_18197), .B0 (sa20[1] ), .Y(n_25672));
OAI21X1 g60897(.A0 (n_20072), .A1 (n_12692), .B0 (n_19934), .Y(n_21016));
OAI21X1 g60903(.A0 (n_20064), .A1 (n_17072), .B0 (n_487), .Y(n_21015));
NOR2X1 g60915(.A (n_14350), .B (n_20611), .Y (n_21014));
OAI21X1 g60923(.A0 (n_20053), .A1 (n_17049), .B0 (sa11[1] ), .Y(n_25613));
OAI21X1 g60928(.A0 (n_20050), .A1 (n_15540), .B0 (n_20574), .Y(n_21012));
OAI21X1 g60932(.A0 (n_27413), .A1 (n_14258), .B0 (sa10[1] ), .Y(n_21010));
OAI21X1 g60937(.A0 (n_20046), .A1 (n_13708), .B0 (n_20810), .Y(n_25696));
NAND4X1 g60938(.A (n_20044), .B (n_19832), .C (n_16867), .D(n_18776), .Y (n_21008));
OAI21X1 g60939(.A0 (n_20043), .A1 (n_17042), .B0 (sa23[1] ), .Y(n_21007));
OAI21X1 g60940(.A0 (n_20123), .A1 (n_20585), .B0 (n_19154), .Y(n_21006));
NAND3X1 g60941(.A (n_18831), .B (n_19270), .C (n_20040), .Y(n_21005));
NAND4X1 g60943(.A (n_25496), .B (n_20438), .C (n_25497), .D(n_13170), .Y (n_21004));
OAI21X1 g60944(.A0 (n_20039), .A1 (n_17039), .B0 (sa10[1] ), .Y(n_28258));
OAI21X1 g60949(.A0 (n_20033), .A1 (n_17032), .B0 (n_19934), .Y(n_21002));
OAI21X1 g60951(.A0 (n_20088), .A1 (n_18552), .B0 (n_20198), .Y(n_21000));
AOI21X1 g60955(.A0 (n_19991), .A1 (n_14907), .B0 (n_26368), .Y(n_20997));
OR4X1 g60969(.A (n_12780), .B (n_13858), .C (n_10175), .D (n_19098),.Y (n_20995));
OR4X1 g60971(.A (n_12580), .B (n_28803), .C (n_9935), .D (n_19096),.Y (n_20994));
AOI21X1 g60980(.A0 (n_18449), .A1 (n_20015), .B0 (n_869), .Y(n_20993));
AOI21X1 g60981(.A0 (n_20091), .A1 (n_19314), .B0 (n_1699), .Y(n_20991));
AOI21X1 g60983(.A0 (n_18422), .A1 (n_20011), .B0 (n_20153), .Y(n_20990));
NAND4X1 g60994(.A (n_20417), .B (n_14674), .C (n_19353), .D(n_16238), .Y (n_20989));
NAND4X1 g61000(.A (n_13745), .B (n_20392), .C (n_18604), .D(n_18605), .Y (n_20988));
NAND2X1 g61006(.A (n_20168), .B (n_20986), .Y (n_20987));
NAND4X1 g61009(.A (n_18459), .B (n_7136), .C (n_9108), .D (n_18672),.Y (n_20985));
NAND3X1 g61013(.A (n_20141), .B (n_19456), .C (n_27341), .Y(n_20984));
NAND4X1 g61014(.A (n_25578), .B (n_17791), .C (n_25579), .D(n_14874), .Y (n_20982));
AOI21X1 g61026(.A0 (n_18706), .A1 (n_26368), .B0 (n_20000), .Y(n_20981));
NAND4X1 g61029(.A (n_17981), .B (n_18809), .C (n_18563), .D(n_17635), .Y (n_20980));
NAND4X1 g61035(.A (n_19605), .B (n_16861), .C (n_18556), .D(n_17602), .Y (n_20979));
NAND4X1 g61065(.A (n_19174), .B (n_14181), .C (n_18681), .D(n_10273), .Y (n_20978));
INVX1 g61072(.A (n_20620), .Y (n_20976));
AOI22X1 g61093(.A0 (n_19459), .A1 (n_196), .B0 (n_19518), .B1(n_17444), .Y (n_20974));
AOI22X1 g61094(.A0 (n_19462), .A1 (n_3264), .B0 (n_19528), .B1(w3[17] ), .Y (n_20972));
NAND4X1 g61098(.A (n_15197), .B (n_13542), .C (n_18530), .D(n_12288), .Y (n_20971));
OAI21X1 g61109(.A0 (n_19220), .A1 (n_18712), .B0 (n_5131), .Y(n_20970));
OAI21X1 g61110(.A0 (n_19236), .A1 (w3[17] ), .B0 (n_19200), .Y(n_20969));
OAI21X1 g61111(.A0 (n_19296), .A1 (n_1558), .B0 (n_19199), .Y(n_20968));
AOI21X1 g61117(.A0 (n_19116), .A1 (n_16497), .B0 (n_1558), .Y(n_20967));
AOI21X1 g61120(.A0 (n_19115), .A1 (n_16506), .B0 (w3[9] ), .Y(n_20966));
AOI21X1 g61122(.A0 (n_19112), .A1 (n_14890), .B0 (n_15482), .Y(n_20965));
AOI21X1 g61123(.A0 (n_16500), .A1 (n_19106), .B0 (sa10[1] ), .Y(n_20964));
AOI21X1 g61126(.A0 (n_14887), .A1 (n_19105), .B0 (n_17246), .Y(n_20962));
OAI21X1 g61139(.A0 (n_19245), .A1 (n_3886), .B0 (n_17359), .Y(n_29429));
NAND2X1 g61142(.A (n_20009), .B (n_19953), .Y (n_20958));
NAND4X1 g61143(.A (n_25806), .B (n_12279), .C (n_15931), .D(n_18368), .Y (n_20957));
NAND4X1 g61145(.A (n_29303), .B (n_14912), .C (n_20955), .D(n_12818), .Y (n_20956));
NAND2X1 g61146(.A (n_19952), .B (n_869), .Y (n_20954));
NAND4X1 g61149(.A (n_29380), .B (n_15040), .C (n_20952), .D(n_12358), .Y (n_20953));
NAND4X1 g61150(.A (n_11077), .B (n_16597), .C (n_20950), .D(n_18257), .Y (n_20951));
NAND4X1 g61154(.A (n_10930), .B (n_17893), .C (n_20948), .D(n_18296), .Y (n_20949));
AOI22X1 g61159(.A0 (n_19298), .A1 (n_11261), .B0 (n_16069), .B1(n_1000), .Y (n_20947));
NAND3X1 g61166(.A (n_19294), .B (n_19348), .C (n_15372), .Y(n_20946));
NAND3X1 g61167(.A (n_18591), .B (n_19351), .C (n_15374), .Y(n_20945));
NAND3X1 g61169(.A (n_19253), .B (n_19349), .C (n_15378), .Y(n_20943));
NAND2X1 g61174(.A (n_19164), .B (n_20021), .Y (n_20941));
NAND2X1 g61180(.A (n_18106), .B (n_19967), .Y (n_20940));
NAND2X1 g61186(.A (n_20019), .B (n_19327), .Y (n_20939));
NAND2X1 g61189(.A (n_19162), .B (n_20017), .Y (n_20938));
NAND4X1 g61193(.A (n_12775), .B (n_7255), .C (n_18212), .D (n_13072),.Y (n_20937));
NAND3X1 g61195(.A (n_10976), .B (n_19223), .C (n_18000), .Y(n_20936));
NAND3X1 g61198(.A (n_29306), .B (n_29307), .C (n_15435), .Y(n_20935));
NAND2X1 g61200(.A (n_20085), .B (n_804), .Y (n_20934));
NOR3X1 g61202(.A (n_13307), .B (n_6848), .C (n_19231), .Y (n_20933));
NAND3X1 g61203(.A (n_10192), .B (n_19320), .C (n_10667), .Y(n_20932));
NAND2X1 g61204(.A (n_20082), .B (sa20[1] ), .Y (n_20931));
NAND3X1 g61209(.A (n_25677), .B (n_17526), .C (n_18619), .Y(n_20929));
NAND3X1 g61210(.A (n_12368), .B (n_19221), .C (n_17972), .Y(n_20928));
NOR3X1 g61211(.A (n_20926), .B (n_14488), .C (n_19203), .Y (n_20927));
NAND4X1 g61219(.A (n_17461), .B (n_18134), .C (n_18357), .D(n_15416), .Y (n_20925));
NAND3X1 g61220(.A (n_18648), .B (n_19308), .C (n_19307), .Y(n_20924));
NAND2X1 g61226(.A (n_18105), .B (n_19965), .Y (n_20923));
OAI21X1 g61229(.A0 (n_19293), .A1 (n_11898), .B0 (n_804), .Y(n_25511));
NAND2X1 g61231(.A (n_20073), .B (n_20632), .Y (n_20921));
NAND2X1 g61235(.A (n_20058), .B (n_20564), .Y (n_20919));
NAND4X1 g61239(.A (n_28263), .B (n_7042), .C (n_28264), .D (n_13002),.Y (n_20918));
NOR3X1 g61245(.A (n_13303), .B (n_5872), .C (n_27289), .Y (n_20916));
NAND3X1 g61247(.A (n_29407), .B (n_29408), .C (n_16793), .Y(n_20914));
NAND2X1 g61253(.A (n_18104), .B (n_19963), .Y (n_20913));
NAND3X1 g61260(.A (n_25627), .B (n_17517), .C (n_16637), .Y(n_20912));
NOR3X1 g61261(.A (n_20910), .B (n_14271), .C (n_19184), .Y (n_20911));
NAND4X1 g61273(.A (n_20832), .B (n_11727), .C (n_18163), .D(n_12944), .Y (n_20906));
NAND3X1 g61274(.A (n_18582), .B (n_19274), .C (n_19273), .Y(n_20905));
NAND2X1 g61275(.A (n_20047), .B (n_20661), .Y (n_20904));
NAND4X1 g61276(.A (n_26721), .B (n_11853), .C (n_18160), .D(n_12943), .Y (n_20903));
OAI21X1 g61277(.A0 (n_19272), .A1 (n_13871), .B0 (n_1991), .Y(n_20902));
NAND3X1 g61281(.A (n_17197), .B (n_17512), .C (n_19271), .Y(n_20901));
NAND3X1 g61285(.A (n_18587), .B (n_19268), .C (n_18596), .Y(n_20900));
OAI21X1 g61286(.A0 (n_19267), .A1 (n_17427), .B0 (sa01[1] ), .Y(n_20899));
NAND3X1 g61291(.A (n_14673), .B (n_19260), .C (n_19259), .Y(n_20898));
OAI21X1 g61297(.A0 (n_19251), .A1 (n_12191), .B0 (n_788), .Y(n_28322));
NAND2X1 g61298(.A (n_19749), .B (n_19993), .Y (n_20896));
OAI21X1 g61299(.A0 (n_19249), .A1 (n_14761), .B0 (n_20574), .Y(n_25582));
NAND3X1 g61302(.A (n_28557), .B (n_19286), .C (n_28558), .Y(n_20894));
OR2X1 g61306(.A (n_16489), .B (n_20099), .Y (n_20893));
OR2X1 g61311(.A (n_16478), .B (n_20092), .Y (n_20891));
AOI21X1 g61312(.A0 (n_19362), .A1 (n_15554), .B0 (n_26368), .Y(n_20890));
AOI21X1 g61313(.A0 (n_19137), .A1 (n_933), .B0 (n_18630), .Y(n_20889));
NAND2X1 g61314(.A (n_20145), .B (n_18937), .Y (n_20888));
AOI21X1 g61315(.A0 (n_19136), .A1 (n_27449), .B0 (n_19880), .Y(n_29124));
OAI21X1 g61317(.A0 (n_19202), .A1 (n_20102), .B0 (n_19869), .Y(n_20886));
AOI21X1 g61318(.A0 (n_19134), .A1 (n_124), .B0 (n_12641), .Y(n_20884));
AOI22X1 g61319(.A0 (n_19257), .A1 (n_17474), .B0 (n_10831), .B1(n_19857), .Y (n_20882));
OAI21X1 g61325(.A0 (n_19189), .A1 (n_21396), .B0 (n_19846), .Y(n_20880));
NAND4X1 g61326(.A (n_19280), .B (n_26952), .C (n_18494), .D(n_12526), .Y (n_20879));
NAND2X1 g61329(.A (n_20140), .B (n_18922), .Y (n_20878));
AOI21X1 g61330(.A0 (n_19133), .A1 (n_20018), .B0 (n_19854), .Y(n_25834));
OAI21X1 g61331(.A0 (n_19132), .A1 (sa32[1] ), .B0 (n_19276), .Y(n_20875));
AOI21X1 g61332(.A0 (n_19131), .A1 (n_20677), .B0 (n_18602), .Y(n_20874));
AOI21X1 g61333(.A0 (n_19129), .A1 (n_21396), .B0 (n_17633), .Y(n_25701));
NAND4X1 g61338(.A (n_19383), .B (n_18645), .C (n_18510), .D(n_12860), .Y (n_20870));
NAND4X1 g61340(.A (n_19379), .B (n_13443), .C (n_18503), .D(n_12709), .Y (n_20869));
NAND4X1 g61342(.A (n_19377), .B (n_18333), .C (n_18497), .D(n_12542), .Y (n_20868));
NAND3X1 g61345(.A (n_19923), .B (n_19118), .C (n_19799), .Y(n_20867));
NAND4X1 g61351(.A (n_15518), .B (n_12657), .C (n_18421), .D(n_18379), .Y (n_20866));
OR4X1 g61353(.A (n_10821), .B (n_28053), .C (n_16119), .D (n_18118),.Y (n_20865));
OR4X1 g61356(.A (n_14398), .B (n_10049), .C (n_27694), .D (n_18123),.Y (n_20864));
NAND2X1 g61362(.A (n_20101), .B (n_20862), .Y (n_20863));
AOI22X1 g61363(.A0 (n_19211), .A1 (n_869), .B0 (n_4470), .B1(n_13076), .Y (n_20861));
AOI22X1 g61365(.A0 (n_19225), .A1 (n_17444), .B0 (n_13237), .B1(n_16480), .Y (n_20860));
AOI21X1 g61368(.A0 (n_12137), .A1 (n_196), .B0 (n_20014), .Y(n_20859));
OAI21X1 g61373(.A0 (n_19331), .A1 (n_15644), .B0 (n_20677), .Y(n_20858));
AOI21X1 g61377(.A0 (n_19352), .A1 (n_11819), .B0 (n_16358), .Y(n_20857));
OAI21X1 g61382(.A0 (n_19123), .A1 (n_12009), .B0 (n_21108), .Y(n_20856));
OAI21X1 g61402(.A0 (n_19190), .A1 (n_2001), .B0 (n_18725), .Y(n_20855));
NAND4X1 g61407(.A (n_19568), .B (n_20853), .C (n_16801), .D(n_18513), .Y (n_20854));
NAND3X1 g61408(.A (n_5896), .B (n_19369), .C (n_14009), .Y (n_20852));
NAND4X1 g61411(.A (n_28267), .B (n_16645), .C (n_28268), .D(n_12946), .Y (n_20851));
NAND3X1 g61414(.A (n_6059), .B (n_19365), .C (n_17563), .Y (n_20850));
NAND3X1 g61416(.A (n_7091), .B (n_19363), .C (n_18682), .Y (n_20849));
NAND4X1 g61426(.A (n_15112), .B (n_16853), .C (n_18447), .D(n_14701), .Y (n_20847));
NAND4X1 g61431(.A (n_13390), .B (n_14588), .C (n_18434), .D(n_11279), .Y (n_20844));
OAI21X1 g61438(.A0 (n_18536), .A1 (n_20841), .B0 (n_20138), .Y(n_20842));
OAI21X1 g61442(.A0 (n_18533), .A1 (sa30[1] ), .B0 (n_20135), .Y(n_20840));
INVX1 g61454(.A (n_20524), .Y (n_20838));
NOR2X1 g61458(.A (n_20075), .B (n_18670), .Y (n_20837));
NAND3X1 g61462(.A (n_19356), .B (n_19109), .C (n_18220), .Y(n_20836));
NAND4X1 g61464(.A (n_14933), .B (n_12072), .C (n_18481), .D(n_14593), .Y (n_20835));
NAND4X1 g61478(.A (n_13440), .B (n_12058), .C (n_18487), .D(n_14625), .Y (n_20834));
NAND4X1 g61482(.A (n_25621), .B (n_20832), .C (n_25622), .D(n_14690), .Y (n_20833));
NAND4X1 g61483(.A (n_14975), .B (n_12012), .C (n_18485), .D(n_11237), .Y (n_20831));
NAND4X1 g61485(.A (n_17887), .B (n_12025), .C (n_18483), .D(n_12902), .Y (n_20830));
NAND4X1 g61487(.A (n_17866), .B (n_19690), .C (n_17410), .D(n_18729), .Y (n_20828));
AOI21X1 g61491(.A0 (n_18906), .A1 (n_21275), .B0 (n_19451), .Y(n_20827));
AOI21X1 g61499(.A0 (n_19169), .A1 (n_191), .B0 (n_19458), .Y(n_20823));
OAI21X1 g61501(.A0 (n_18541), .A1 (n_19942), .B0 (n_20020), .Y(n_20821));
AOI21X1 g61502(.A0 (n_19168), .A1 (n_15766), .B0 (n_19453), .Y(n_20820));
OAI21X1 g61504(.A0 (n_18539), .A1 (n_778), .B0 (n_19999), .Y(n_20819));
OAI21X1 g61506(.A0 (n_19167), .A1 (sa32[1] ), .B0 (n_19448), .Y(n_20818));
OAI21X1 g61507(.A0 (n_19166), .A1 (n_903), .B0 (n_19994), .Y(n_20816));
NAND2X1 g61518(.A (n_19779), .B (n_20648), .Y (n_20815));
OAI21X1 g61522(.A0 (n_27753), .A1 (n_17652), .B0 (n_5131), .Y(n_20814));
OAI21X1 g61531(.A0 (n_18884), .A1 (n_17192), .B0 (n_20810), .Y(n_20811));
OAI21X1 g61538(.A0 (n_18915), .A1 (n_14604), .B0 (n_5131), .Y(n_20809));
AOI21X1 g61551(.A0 (n_14236), .A1 (n_19042), .B0 (n_16466), .Y(n_20808));
AOI21X1 g61557(.A0 (n_17620), .A1 (n_19041), .B0 (n_15166), .Y(n_20806));
NOR3X1 g61565(.A (n_12112), .B (n_7043), .C (n_19057), .Y (n_20805));
AOI21X1 g61568(.A0 (n_14360), .A1 (n_19040), .B0 (n_16835), .Y(n_20804));
OAI21X1 g61569(.A0 (n_18314), .A1 (n_18913), .B0 (n_844), .Y(n_20803));
OAI21X1 g61575(.A0 (n_18865), .A1 (n_13926), .B0 (sa22[1] ), .Y(n_20802));
NAND2X1 g61580(.A (n_19817), .B (n_1991), .Y (n_28269));
NAND2X1 g61590(.A (n_19813), .B (n_903), .Y (n_20798));
AOI21X1 g61595(.A0 (n_4904), .A1 (n_19361), .B0 (n_19776), .Y(n_20796));
AOI21X1 g61602(.A0 (n_9044), .A1 (n_20105), .B0 (n_19943), .Y(n_20795));
INVX1 g61618(.A (n_20473), .Y (n_20794));
INVX1 g61624(.A (n_20472), .Y (n_20792));
NAND2X1 g61629(.A (n_19761), .B (n_1991), .Y (n_20791));
AOI22X1 g61661(.A0 (n_18936), .A1 (n_21174), .B0 (n_8605), .B1(n_20765), .Y (n_25623));
OAI21X1 g61668(.A0 (n_19023), .A1 (n_20786), .B0 (n_1310), .Y(n_25483));
NOR2X1 g61688(.A (n_19762), .B (w3[17] ), .Y (n_20785));
NAND2X1 g61693(.A (n_19807), .B (n_19143), .Y (n_20784));
AOI22X1 g61694(.A0 (n_18930), .A1 (n_5131), .B0 (n_8500), .B1(n_20760), .Y (n_20783));
OAI21X1 g61699(.A0 (n_18971), .A1 (n_7117), .B0 (n_17246), .Y(n_20781));
AOI21X1 g61708(.A0 (n_18804), .A1 (n_18963), .B0 (n_20144), .Y(n_20780));
NAND3X1 g61712(.A (n_17623), .B (n_20192), .C (n_19013), .Y(n_20778));
OAI21X1 g61720(.A0 (n_17973), .A1 (n_19068), .B0 (n_19414), .Y(n_20777));
NAND2X1 g61735(.A (n_19782), .B (n_903), .Y (n_20775));
NAND2X1 g61746(.A (n_19847), .B (n_3538), .Y (n_28881));
NAND2X1 g61762(.A (n_19778), .B (n_19995), .Y (n_20772));
NOR3X1 g61788(.A (n_12776), .B (n_9395), .C (n_19085), .Y (n_20771));
AOI21X1 g61799(.A0 (n_15192), .A1 (n_18957), .B0 (n_129), .Y(n_20770));
OAI21X1 g61802(.A0 (n_19045), .A1 (n_9775), .B0 (n_20767), .Y(n_20768));
AOI21X1 g61808(.A0 (n_11978), .A1 (n_20765), .B0 (n_19936), .Y(n_20766));
OAI21X1 g61812(.A0 (n_19044), .A1 (n_8306), .B0 (n_487), .Y(n_20764));
INVX1 g61814(.A (n_20418), .Y (n_20762));
AOI21X1 g61824(.A0 (n_9135), .A1 (n_20760), .B0 (n_19935), .Y(n_20761));
OAI21X1 g61831(.A0 (n_19043), .A1 (n_9541), .B0 (n_20758), .Y(n_20759));
NAND3X1 g61841(.A (n_17470), .B (n_19037), .C (n_19648), .Y(n_20757));
NAND3X1 g61842(.A (n_16139), .B (n_19082), .C (n_15509), .Y(n_20756));
INVX1 g61853(.A (n_20407), .Y (n_20755));
NAND3X1 g61858(.A (n_19881), .B (n_18097), .C (n_11641), .Y(n_20754));
NAND3X1 g61862(.A (n_19875), .B (n_18880), .C (n_13751), .Y(n_20753));
NAND3X1 g61863(.A (n_28804), .B (n_19075), .C (n_15513), .Y(n_20752));
NAND2X1 g61888(.A (n_19856), .B (n_20677), .Y (n_28501));
NAND3X1 g61889(.A (n_19855), .B (n_18090), .C (n_13810), .Y(n_20750));
OAI21X1 g61922(.A0 (n_18973), .A1 (n_13976), .B0 (n_19940), .Y(n_20748));
AOI22X1 g61937(.A0 (n_18934), .A1 (n_282), .B0 (n_3266), .B1(n_19226), .Y (n_20747));
NAND2X1 g61940(.A (n_16788), .B (n_19867), .Y (n_20746));
AOI22X1 g61943(.A0 (n_18929), .A1 (n_196), .B0 (n_6567), .B1(n_5887), .Y (n_20745));
NAND4X1 g61152(.A (n_12669), .B (n_15000), .C (n_20743), .D(n_18308), .Y (n_20744));
AOI22X1 g61959(.A0 (n_18883), .A1 (n_29039), .B0 (n_14403), .B1(n_29074), .Y (n_20742));
AOI22X1 g61965(.A0 (n_18940), .A1 (n_933), .B0 (n_4264), .B1(n_4965), .Y (n_20739));
NAND2X1 g61989(.A (n_14569), .B (n_19911), .Y (n_20738));
NAND2X1 g61993(.A (n_12636), .B (n_19910), .Y (n_20737));
AOI21X1 g62002(.A0 (n_18871), .A1 (sa33[1] ), .B0 (n_12457), .Y(n_20735));
NAND2X1 g62037(.A (n_19620), .B (n_1008), .Y (n_20734));
NAND2X1 g62071(.A (n_19649), .B (n_20585), .Y (n_20733));
NAND2X1 g62079(.A (n_19639), .B (n_16358), .Y (n_20732));
OAI21X1 g62110(.A0 (n_19580), .A1 (n_17936), .B0 (n_20729), .Y(n_20730));
NAND2X1 g62134(.A (n_19631), .B (n_27216), .Y (n_20728));
AND2X1 g62230(.A (n_19681), .B (n_7847), .Y (n_20725));
NAND2X1 g62295(.A (n_19682), .B (n_19046), .Y (n_20724));
AND2X1 g62343(.A (n_19637), .B (n_11819), .Y (n_20723));
NOR2X1 g62384(.A (n_19619), .B (n_21174), .Y (n_20722));
OAI21X1 g62389(.A0 (n_16605), .A1 (n_18846), .B0 (sa00[1] ), .Y(n_20721));
NAND2X1 g62420(.A (n_19658), .B (n_18437), .Y (n_20720));
NAND4X1 g61151(.A (n_12816), .B (n_15007), .C (n_27131), .D(n_18313), .Y (n_20719));
AOI21X1 g62576(.A0 (n_19588), .A1 (n_9435), .B0 (n_16649), .Y(n_20717));
AOI21X1 g62577(.A0 (n_19586), .A1 (n_13031), .B0 (n_18617), .Y(n_20716));
AOI21X1 g62601(.A0 (n_19595), .A1 (n_12892), .B0 (n_18643), .Y(n_20715));
AND2X1 g62604(.A (n_19663), .B (n_13423), .Y (n_20713));
NAND2X1 g62692(.A (n_19660), .B (n_18970), .Y (n_20711));
INVX1 g62787(.A (n_20251), .Y (n_20710));
INVX1 g63288(.A (n_20232), .Y (n_25612));
OAI21X1 g63295(.A0 (n_19564), .A1 (n_20705), .B0 (n_21174), .Y(n_20706));
INVX1 g63336(.A (n_20230), .Y (n_20701));
AND2X1 g63371(.A (n_20172), .B (n_26874), .Y (n_20699));
AOI21X1 g60471(.A0 (n_19577), .A1 (n_933), .B0 (n_18656), .Y(n_20698));
NAND2X1 g60474(.A (n_19612), .B (n_187), .Y (n_25711));
AOI21X1 g60475(.A0 (n_19575), .A1 (n_20213), .B0 (n_19332), .Y(n_20695));
AOI21X1 g60476(.A0 (n_19574), .A1 (n_124), .B0 (n_18653), .Y(n_20694));
NAND2X1 g60483(.A (n_19611), .B (n_27242), .Y (n_20693));
OAI21X1 g60484(.A0 (n_19591), .A1 (n_16023), .B0 (n_20677), .Y(n_28850));
OAI21X1 g60489(.A0 (n_19587), .A1 (n_14244), .B0 (n_20680), .Y(n_20690));
NAND2X1 g60498(.A (n_19609), .B (n_21314), .Y (n_25455));
OAI21X1 g60526(.A0 (n_19566), .A1 (n_15551), .B0 (n_15482), .Y(n_20688));
OAI21X1 g60528(.A0 (n_19565), .A1 (n_15547), .B0 (n_16944), .Y(n_20686));
OAI21X1 g63770(.A0 (n_12681), .A1 (n_3886), .B0 (n_21215), .Y(n_20685));
OAI21X1 g60766(.A0 (n_19548), .A1 (n_14536), .B0 (n_196), .Y(n_20684));
OAI21X1 g60779(.A0 (n_19471), .A1 (n_12314), .B0 (n_20517), .Y(n_20683));
OAI21X1 g60781(.A0 (n_19431), .A1 (n_14468), .B0 (n_21174), .Y(n_20682));
OAI21X1 g60787(.A0 (n_19418), .A1 (n_16115), .B0 (n_21055), .Y(n_20679));
OAI21X1 g60791(.A0 (n_19427), .A1 (n_14382), .B0 (n_20677), .Y(n_20678));
OAI21X1 g60798(.A0 (n_19424), .A1 (n_17585), .B0 (n_1008), .Y(n_20675));
OAI21X1 g60804(.A0 (n_19421), .A1 (n_14095), .B0 (n_1196), .Y(n_29383));
AOI22X1 g60854(.A0 (n_19550), .A1 (n_19372), .B0 (n_9719), .B1(n_19896), .Y (n_20668));
OAI21X1 g60861(.A0 (n_19464), .A1 (n_15447), .B0 (n_20204), .Y(n_20667));
OAI21X1 g60865(.A0 (n_19544), .A1 (n_14514), .B0 (n_20587), .Y(n_20664));
OAI21X1 g60873(.A0 (n_19536), .A1 (n_12736), .B0 (n_20116), .Y(n_20663));
OAI21X1 g60879(.A0 (n_19531), .A1 (n_9968), .B0 (n_20661), .Y(n_20662));
OAI21X1 g60882(.A0 (n_19530), .A1 (n_14253), .B0 (sa22[1] ), .Y(n_20660));
OR2X1 g60883(.A (n_19796), .B (n_20164), .Y (n_20659));
NAND4X1 g60887(.A (n_19983), .B (n_20096), .C (n_18624), .D(n_14856), .Y (n_20658));
OAI21X1 g60895(.A0 (n_19522), .A1 (n_7673), .B0 (n_20577), .Y(n_20657));
NOR2X1 g60900(.A (n_17070), .B (n_20163), .Y (n_20656));
OAI21X1 g60902(.A0 (n_19516), .A1 (n_15545), .B0 (n_20116), .Y(n_29424));
OAI21X1 g60909(.A0 (n_19504), .A1 (n_14376), .B0 (n_20558), .Y(n_20654));
OAI21X1 g60918(.A0 (n_19500), .A1 (n_14345), .B0 (n_20585), .Y(n_20651));
OAI21X1 g60922(.A0 (n_19498), .A1 (n_14326), .B0 (sa01[1] ), .Y(n_20650));
OAI21X1 g60931(.A0 (n_19491), .A1 (n_14269), .B0 (n_20648), .Y(n_20647));
NAND4X1 g60935(.A (n_19980), .B (n_20062), .C (n_18601), .D(n_13178), .Y (n_20645));
OAI21X1 g60936(.A0 (n_26468), .A1 (n_12719), .B0 (n_20610), .Y(n_20644));
NAND2X1 g60945(.A (n_20165), .B (sa21[1] ), .Y (n_20643));
OAI21X1 g60948(.A0 (n_19481), .A1 (n_15532), .B0 (n_903), .Y(n_29125));
AOI22X1 g60953(.A0 (n_19472), .A1 (n_21055), .B0 (n_8079), .B1(n_11261), .Y (n_28315));
NAND4X1 g60958(.A (n_11559), .B (n_17402), .C (n_19951), .D(n_18568), .Y (n_20639));
OR2X1 g60968(.A (n_20155), .B (n_13522), .Y (n_20638));
AOI21X1 g60982(.A0 (n_19439), .A1 (w3[9] ), .B0 (n_15941), .Y(n_20637));
AOI21X1 g60987(.A0 (n_19515), .A1 (n_20634), .B0 (w3[17] ), .Y(n_20635));
AOI21X1 g60988(.A0 (n_19432), .A1 (n_20632), .B0 (n_17630), .Y(n_20633));
NAND4X1 g61008(.A (n_18462), .B (n_5818), .C (n_12779), .D (n_17554),.Y (n_20631));
NAND4X1 g61010(.A (n_18457), .B (n_6278), .C (n_20628), .D (n_17551),.Y (n_20629));
NAND4X1 g61011(.A (n_18455), .B (n_8292), .C (n_20626), .D (n_17549),.Y (n_20627));
NAND4X1 g61027(.A (n_19434), .B (n_17062), .C (n_15240), .D(n_13129), .Y (n_20625));
NAND4X1 g61038(.A (n_16675), .B (n_14370), .C (n_17473), .D(n_14237), .Y (n_20624));
NAND4X1 g61049(.A (n_17487), .B (n_8482), .C (n_17572), .D (n_10580),.Y (n_20623));
NAND4X1 g61059(.A (n_17479), .B (n_8744), .C (n_17568), .D (n_10441),.Y (n_20622));
NAND4X1 g61061(.A (n_25550), .B (n_8655), .C (n_25551), .D (n_13917),.Y (n_20621));
NAND4X1 g61073(.A (n_19415), .B (n_15935), .C (n_17499), .D (n_5907),.Y (n_20620));
NAND4X1 g61086(.A (n_8535), .B (n_13495), .C (n_16790), .D (n_17437),.Y (n_20619));
NAND2X1 g65178(.A (n_17031), .B (n_20617), .Y (n_20618));
AOI21X1 g61087(.A0 (n_17629), .A1 (n_19143), .B0 (n_19302), .Y(n_20616));
AOI21X1 g61105(.A0 (n_18519), .A1 (n_13614), .B0 (sa33[1] ), .Y(n_20615));
AOI21X1 g61127(.A0 (n_13253), .A1 (n_18514), .B0 (n_20610), .Y(n_20611));
OAI21X1 g61133(.A0 (n_18616), .A1 (n_19651), .B0 (n_17386), .Y(n_20609));
AOI21X1 g61137(.A0 (n_18590), .A1 (n_28692), .B0 (n_18423), .Y(n_20608));
OAI21X1 g61138(.A0 (n_18586), .A1 (sa01[2] ), .B0 (n_17361), .Y(n_20607));
NAND2X1 g61141(.A (n_19463), .B (n_19428), .Y (n_20606));
NAND2X1 g61144(.A (n_19461), .B (n_19955), .Y (n_20605));
NAND3X1 g61147(.A (n_25780), .B (n_14742), .C (n_15555), .Y(n_20604));
AOI21X1 g61157(.A0 (n_18651), .A1 (n_18369), .B0 (n_12674), .Y(n_20603));
AOI22X1 g61162(.A0 (n_18593), .A1 (n_29062), .B0 (n_14202), .B1(n_29039), .Y (n_20602));
NAND3X1 g61170(.A (n_17346), .B (n_18236), .C (n_18680), .Y(n_20601));
OAI21X1 g61173(.A0 (n_11566), .A1 (n_18578), .B0 (n_20204), .Y(n_20600));
OAI21X1 g61176(.A0 (n_25732), .A1 (n_25733), .B0 (n_804), .Y(n_25454));
OAI21X1 g61178(.A0 (n_18003), .A1 (n_18577), .B0 (n_21151), .Y(n_20598));
NAND4X1 g61181(.A (n_16127), .B (n_8140), .C (n_17080), .D (n_14714),.Y (n_20596));
NAND2X1 g61190(.A (n_19545), .B (n_869), .Y (n_20595));
NAND4X1 g61191(.A (n_12777), .B (n_9928), .C (n_17067), .D (n_11856),.Y (n_20594));
NAND2X1 g61194(.A (n_19543), .B (n_20841), .Y (n_20593));
NAND3X1 g61197(.A (n_17312), .B (n_18797), .C (n_18678), .Y(n_20592));
NAND2X1 g61206(.A (n_19535), .B (n_21151), .Y (n_20591));
NAND2X1 g61208(.A (n_19534), .B (n_20153), .Y (n_20590));
NAND2X1 g61212(.A (n_19526), .B (n_20587), .Y (n_25584));
OAI21X1 g61217(.A0 (n_17986), .A1 (n_18575), .B0 (n_20585), .Y(n_25782));
NAND3X1 g61218(.A (n_6969), .B (n_18622), .C (n_9525), .Y (n_20584));
OR4X1 g61221(.A (n_20582), .B (n_11333), .C (n_7653), .D (n_17074),.Y (n_20583));
OAI21X1 g61222(.A0 (n_18585), .A1 (n_15792), .B0 (n_2204), .Y(n_20581));
OAI21X1 g61223(.A0 (n_17978), .A1 (n_18574), .B0 (n_20579), .Y(n_20580));
NAND2X1 g61224(.A (n_19521), .B (n_20577), .Y (n_20578));
NAND3X1 g61225(.A (n_6511), .B (n_18621), .C (n_7609), .Y (n_20576));
NAND2X1 g61232(.A (n_19511), .B (n_20574), .Y (n_20575));
OAI21X1 g61236(.A0 (n_17963), .A1 (n_18573), .B0 (n_20574), .Y(n_20573));
NAND2X1 g61240(.A (n_19503), .B (sa30[1] ), .Y (n_20572));
NAND3X1 g61241(.A (n_17238), .B (n_17770), .C (n_18676), .Y(n_20571));
OAI21X1 g61243(.A0 (n_11534), .A1 (n_18576), .B0 (n_20198), .Y(n_25710));
OAI21X1 g61250(.A0 (n_28239), .A1 (n_28240), .B0 (n_778), .Y(n_28851));
OR4X1 g61252(.A (n_7656), .B (n_11275), .C (n_20567), .D (n_17053),.Y (n_20568));
NAND4X1 g61255(.A (n_18996), .B (n_14660), .C (n_28607), .D(n_17129), .Y (n_20566));
OAI21X1 g61256(.A0 (n_17944), .A1 (n_18571), .B0 (n_20564), .Y(n_20565));
NAND4X1 g61257(.A (n_16010), .B (n_8247), .C (n_17050), .D (n_16215),.Y (n_20563));
NAND2X1 g61258(.A (n_19497), .B (sa23[1] ), .Y (n_20562));
NAND2X1 g61259(.A (n_19496), .B (n_20579), .Y (n_20560));
NAND2X1 g61263(.A (n_19492), .B (n_20558), .Y (n_25640));
NAND2X1 g61267(.A (n_19490), .B (n_2249), .Y (n_20557));
NAND2X1 g61278(.A (n_19485), .B (n_20055), .Y (n_20555));
NAND2X1 g61280(.A (n_19482), .B (n_778), .Y (n_20554));
OAI21X1 g61282(.A0 (n_18599), .A1 (n_20551), .B0 (sa21[1] ), .Y(n_20552));
NAND2X1 g61289(.A (n_19541), .B (n_20153), .Y (n_20550));
OAI21X1 g61292(.A0 (n_18594), .A1 (n_15743), .B0 (n_16358), .Y(n_20549));
NAND2X1 g61303(.A (n_19552), .B (n_20157), .Y (n_20548));
AOI21X1 g61307(.A0 (n_12810), .A1 (n_19385), .B0 (n_19547), .Y(n_20547));
AOI21X1 g61316(.A0 (n_18523), .A1 (n_282), .B0 (n_17522), .Y(n_20546));
AOI22X1 g61323(.A0 (n_18611), .A1 (n_28689), .B0 (n_14279), .B1(n_28692), .Y (n_20544));
AOI22X1 g61324(.A0 (n_18610), .A1 (n_477), .B0 (n_10969), .B1(n_9106), .Y (n_20543));
OR4X1 g61347(.A (n_12831), .B (n_10209), .C (n_15906), .D (n_17015),.Y (n_20541));
OR4X1 g61348(.A (n_11134), .B (n_12246), .C (n_16121), .D (n_17013),.Y (n_20540));
OR4X1 g61349(.A (n_14570), .B (n_9913), .C (n_14503), .D (n_17010),.Y (n_20539));
OR4X1 g61357(.A (n_14294), .B (n_10217), .C (n_12510), .D (n_17009),.Y (n_20538));
OR4X1 g61358(.A (n_14153), .B (n_9787), .C (n_14277), .D (n_17007),.Y (n_20537));
OR4X1 g61359(.A (n_10866), .B (n_8638), .C (n_20535), .D (n_17006),.Y (n_20536));
OR4X1 g61360(.A (n_12360), .B (n_14037), .C (n_16059), .D (n_17001),.Y (n_20534));
OR4X1 g61361(.A (n_12355), .B (n_12664), .C (n_15937), .D (n_17002),.Y (n_20533));
NAND4X1 g61364(.A (n_11063), .B (n_18635), .C (n_7847), .D (n_17174),.Y (n_20532));
OAI21X1 g61389(.A0 (n_18567), .A1 (w3[9] ), .B0 (n_18101), .Y(n_20530));
OAI21X1 g61390(.A0 (n_18565), .A1 (n_20577), .B0 (n_18093), .Y(n_20529));
NAND4X1 g61398(.A (n_11557), .B (n_20526), .C (n_11378), .D(n_16935), .Y (n_20528));
NAND4X1 g61412(.A (n_20526), .B (n_13536), .C (n_20468), .D(n_17429), .Y (n_20527));
NAND4X1 g61428(.A (n_15228), .B (n_15116), .C (n_17376), .D(n_13050), .Y (n_20525));
NAND4X1 g61455(.A (n_19113), .B (n_18210), .C (n_16210), .D(n_16994), .Y (n_20524));
AOI22X1 g61460(.A0 (n_18559), .A1 (n_20577), .B0 (n_12906), .B1(n_16978), .Y (n_20523));
NAND4X1 g61470(.A (n_17850), .B (n_10469), .C (n_17408), .D(n_16182), .Y (n_20522));
NAND4X1 g61480(.A (n_13308), .B (n_17935), .C (n_17415), .D(n_12932), .Y (n_20521));
NAND4X1 g61484(.A (n_14974), .B (n_11956), .C (n_17413), .D(n_14623), .Y (n_20520));
AOI22X1 g61497(.A0 (n_18570), .A1 (n_20518), .B0 (n_20517), .B1(n_29180), .Y (n_20519));
OAI21X1 g61503(.A0 (n_18540), .A1 (sa11[1] ), .B0 (n_19452), .Y(n_20516));
NAND2X1 g61512(.A (n_19107), .B (n_933), .Y (n_20515));
OAI21X1 g61515(.A0 (n_18410), .A1 (n_10796), .B0 (n_3264), .Y(n_20513));
NAND2X1 g61520(.A (n_19177), .B (n_20157), .Y (n_20512));
OAI21X1 g61521(.A0 (n_18821), .A1 (n_17176), .B0 (n_21242), .Y(n_20511));
OAI21X1 g61529(.A0 (n_13696), .A1 (n_18302), .B0 (n_20767), .Y(n_20509));
OAI21X1 g61539(.A0 (n_18154), .A1 (n_14656), .B0 (n_14630), .Y(n_20508));
AOI21X1 g61543(.A0 (n_14522), .A1 (n_18418), .B0 (n_19364), .Y(n_20506));
NAND3X1 g61546(.A (n_12312), .B (n_18150), .C (n_16554), .Y(n_20505));
NAND3X1 g61547(.A (n_18099), .B (n_15561), .C (n_18398), .Y(n_20504));
OAI21X1 g61549(.A0 (n_12763), .A1 (n_18479), .B0 (n_19433), .Y(n_20503));
OAI21X1 g61550(.A0 (n_17305), .A1 (n_18207), .B0 (n_2204), .Y(n_20502));
OAI21X1 g61552(.A0 (n_18442), .A1 (n_3612), .B0 (n_12341), .Y(n_20501));
NOR3X1 g61553(.A (n_10548), .B (n_9537), .C (n_18460), .Y (n_20500));
AOI21X1 g61554(.A0 (n_15924), .A1 (n_18415), .B0 (n_18369), .Y(n_20499));
OAI21X1 g61555(.A0 (n_17271), .A1 (n_18192), .B0 (sa00[1] ), .Y(n_20498));
NAND3X1 g61558(.A (n_11154), .B (n_18234), .C (n_13424), .Y(n_20496));
AOI21X1 g61560(.A0 (n_14408), .A1 (n_18413), .B0 (n_28642), .Y(n_20495));
OAI21X1 g61561(.A0 (n_18436), .A1 (n_20477), .B0 (n_14582), .Y(n_20494));
OAI21X1 g61563(.A0 (n_17224), .A1 (n_18177), .B0 (sa01[1] ), .Y(n_20493));
AOI21X1 g61567(.A0 (n_18027), .A1 (n_17130), .B0 (n_2681), .Y(n_20491));
OAI21X1 g61570(.A0 (n_18425), .A1 (n_27407), .B0 (n_12393), .Y(n_20489));
AOI21X1 g61576(.A0 (n_14438), .A1 (n_18411), .B0 (n_14474), .Y(n_20488));
NAND2X1 g61578(.A (n_19237), .B (n_2981), .Y (n_20487));
NAND3X1 g61579(.A (n_27496), .B (n_18129), .C (n_13576), .Y(n_20485));
NAND2X1 g61584(.A (n_19224), .B (n_16362), .Y (n_20484));
NAND2X1 g61592(.A (n_19213), .B (n_844), .Y (n_20483));
OAI21X1 g61594(.A0 (n_18429), .A1 (n_14816), .B0 (n_844), .Y(n_20482));
OAI21X1 g61600(.A0 (n_18420), .A1 (n_11423), .B0 (sa33[1] ), .Y(n_20480));
NAND2X1 g61606(.A (n_19149), .B (n_20116), .Y (n_29414));
AOI21X1 g61610(.A0 (n_18232), .A1 (n_7478), .B0 (n_20477), .Y(n_20478));
OAI21X1 g61614(.A0 (n_18405), .A1 (n_12266), .B0 (n_18326), .Y(n_20476));
AOI21X1 g61616(.A0 (n_18229), .A1 (n_15835), .B0 (n_1310), .Y(n_20475));
AOI21X1 g61619(.A0 (n_13553), .A1 (n_18073), .B0 (n_21174), .Y(n_20473));
NAND3X1 g61625(.A (n_15912), .B (n_19608), .C (n_18401), .Y(n_20472));
AOI21X1 g61627(.A0 (n_18255), .A1 (n_4582), .B0 (n_11424), .Y(n_20471));
NOR2X1 g61628(.A (n_12720), .B (n_28242), .Y (n_20470));
AND2X1 g61634(.A (n_19328), .B (n_20468), .Y (n_20469));
NOR2X1 g61636(.A (n_19334), .B (n_15939), .Y (n_20467));
AOI21X1 g61637(.A0 (n_18216), .A1 (n_10574), .B0 (n_1756), .Y(n_20466));
NAND3X1 g61639(.A (n_9870), .B (n_18214), .C (n_16543), .Y (n_20465));
NAND3X1 g61640(.A (n_17592), .B (n_11730), .C (n_18397), .Y(n_20464));
NAND4X1 g61653(.A (n_25508), .B (n_19297), .C (n_14930), .D(n_17328), .Y (n_20463));
AOI21X1 g61663(.A0 (n_15693), .A1 (n_16466), .B0 (n_19333), .Y(n_20462));
NAND3X1 g61664(.A (n_19228), .B (n_13700), .C (n_17083), .Y(n_20461));
OAI21X1 g61665(.A0 (n_15306), .A1 (n_18443), .B0 (n_804), .Y(n_20460));
AOI21X1 g61672(.A0 (n_17987), .A1 (n_18441), .B0 (n_20457), .Y(n_20458));
AOI21X1 g61675(.A0 (n_15234), .A1 (n_18439), .B0 (n_171), .Y(n_20456));
NAND2X1 g61682(.A (n_19217), .B (n_663), .Y (n_20455));
NAND3X1 g61684(.A (n_15223), .B (n_18233), .C (n_16879), .Y(n_20454));
NAND2X1 g61697(.A (n_19103), .B (n_16510), .Y (n_20453));
NAND2X1 g61701(.A (n_14885), .B (n_19108), .Y (n_20452));
NAND3X1 g61702(.A (n_19227), .B (n_13697), .C (n_18199), .Y(n_20451));
NAND3X1 g61707(.A (n_14783), .B (n_9352), .C (n_18350), .Y (n_20450));
OAI21X1 g61721(.A0 (n_13422), .A1 (n_18345), .B0 (n_778), .Y(n_20448));
NAND3X1 g61725(.A (n_13843), .B (n_18189), .C (n_16426), .Y(n_20447));
INVX1 g61733(.A (n_20057), .Y (n_20444));
OAI21X1 g61742(.A0 (n_18337), .A1 (n_8405), .B0 (n_908), .Y(n_20443));
NAND3X1 g61745(.A (n_15095), .B (n_18183), .C (n_16878), .Y(n_20442));
OAI21X1 g61749(.A0 (n_16731), .A1 (n_18433), .B0 (n_788), .Y(n_20441));
NAND4X1 g61750(.A (n_20438), .B (n_17744), .C (n_17937), .D(n_12963), .Y (n_20439));
NAND4X1 g61755(.A (n_13795), .B (n_20169), .C (n_17932), .D(n_11266), .Y (n_20437));
NAND4X1 g61756(.A (n_19001), .B (n_18801), .C (n_14328), .D(n_13329), .Y (n_25642));
AOI21X1 g61758(.A0 (n_18843), .A1 (n_18431), .B0 (n_26931), .Y(n_20435));
AOI21X1 g61760(.A0 (n_16707), .A1 (n_18430), .B0 (n_187), .Y(n_20432));
NAND3X1 g61769(.A (n_18838), .B (n_18162), .C (n_18013), .Y(n_20431));
NAND2X1 g61773(.A (n_19101), .B (n_15076), .Y (n_20430));
AOI21X1 g61782(.A0 (n_16660), .A1 (n_18424), .B0 (n_21108), .Y(n_20429));
AOI21X1 g61784(.A0 (n_18156), .A1 (n_27910), .B0 (n_13023), .Y(n_20428));
NAND3X1 g61785(.A (n_14226), .B (n_6966), .C (n_18412), .Y (n_20426));
AOI21X1 g61798(.A0 (n_18109), .A1 (n_14627), .B0 (n_14052), .Y(n_20422));
NOR2X1 g61806(.A (n_19121), .B (n_9556), .Y (n_20419));
NAND3X1 g61815(.A (n_12345), .B (n_20417), .C (n_18279), .Y(n_20418));
AOI21X1 g61817(.A0 (n_18273), .A1 (n_27900), .B0 (n_27604), .Y(n_20416));
NAND2X1 g61833(.A (n_19240), .B (n_20412), .Y (n_29315));
AOI21X1 g61834(.A0 (n_18258), .A1 (n_12042), .B0 (n_15574), .Y(n_20411));
AOI21X1 g61836(.A0 (n_18270), .A1 (n_19433), .B0 (n_17787), .Y(n_20410));
NAND2X1 g61852(.A (n_16989), .B (n_19325), .Y (n_20408));
AOI21X1 g61854(.A0 (n_18213), .A1 (n_17321), .B0 (n_20406), .Y(n_20407));
NOR2X1 g61856(.A (n_16811), .B (n_19204), .Y (n_20405));
NAND3X1 g61864(.A (n_17797), .B (n_18367), .C (n_18142), .Y(n_20404));
INVX1 g61867(.A (n_20008), .Y (n_20403));
INVX1 g61874(.A (n_20007), .Y (n_20401));
NAND2X1 g61881(.A (n_19313), .B (n_20399), .Y (n_20400));
OAI21X1 g61882(.A0 (n_18280), .A1 (n_12154), .B0 (n_20397), .Y(n_20398));
NAND3X1 g61898(.A (n_18603), .B (n_18084), .C (n_9904), .Y (n_20396));
AOI21X1 g61900(.A0 (n_18161), .A1 (n_27910), .B0 (n_18997), .Y(n_25506));
AOI21X1 g61908(.A0 (n_18033), .A1 (n_17734), .B0 (n_21396), .Y(n_20394));
AOI21X1 g61911(.A0 (n_18032), .A1 (n_20392), .B0 (n_21133), .Y(n_20393));
NAND2X1 g61917(.A (n_19252), .B (n_20388), .Y (n_20389));
OAI21X1 g61918(.A0 (n_18288), .A1 (n_12161), .B0 (n_20386), .Y(n_20387));
OAI21X1 g61919(.A0 (n_18282), .A1 (n_10129), .B0 (n_21133), .Y(n_20385));
NAND2X1 g61921(.A (n_19250), .B (n_19830), .Y (n_20384));
NAND3X1 g61924(.A (n_18767), .B (n_18271), .C (n_18946), .Y(n_20383));
NAND2X1 g61925(.A (n_19248), .B (n_21275), .Y (n_20382));
OAI21X1 g61928(.A0 (n_18261), .A1 (n_19207), .B0 (n_1196), .Y(n_20380));
AOI21X1 g61930(.A0 (n_10804), .A1 (n_378), .B0 (n_19242), .Y(n_29314));
AOI21X1 g61931(.A0 (n_10788), .A1 (n_27481), .B0 (n_26839), .Y(n_20378));
OAI21X1 g61932(.A0 (n_18260), .A1 (n_17491), .B0 (n_27216), .Y(n_29367));
AOI22X1 g61934(.A0 (n_18117), .A1 (n_19433), .B0 (n_11108), .B1(n_12827), .Y (n_20375));
NAND2X1 g61939(.A (n_16576), .B (n_19304), .Y (n_20374));
NOR2X1 g61947(.A (n_15402), .B (n_19413), .Y (n_20373));
NAND2X1 g61955(.A (n_16636), .B (n_19263), .Y (n_20372));
NAND2X1 g61956(.A (n_17896), .B (n_19261), .Y (n_20371));
NAND2X1 g61958(.A (n_16624), .B (n_19258), .Y (n_20370));
AOI22X1 g61964(.A0 (n_18039), .A1 (n_16553), .B0 (n_13827), .B1(n_14548), .Y (n_20369));
AOI22X1 g61966(.A0 (n_18044), .A1 (n_13423), .B0 (n_15774), .B1(n_16895), .Y (n_20367));
NAND4X1 g61974(.A (n_15178), .B (n_19420), .C (n_17721), .D(n_12317), .Y (n_20365));
NAND3X1 g61975(.A (n_17890), .B (n_18082), .C (n_19949), .Y(n_20364));
NAND4X1 g61986(.A (n_12834), .B (n_18343), .C (n_13962), .D(n_16933), .Y (n_20363));
NAND4X1 g61987(.A (n_19216), .B (n_18361), .C (n_13676), .D(n_16929), .Y (n_20362));
NAND4X1 g61988(.A (n_16564), .B (n_11056), .C (n_20360), .D(n_16928), .Y (n_20361));
OAI21X1 g61990(.A0 (n_18041), .A1 (n_20457), .B0 (n_14553), .Y(n_20359));
OAI21X1 g61996(.A0 (n_18037), .A1 (n_26931), .B0 (n_14458), .Y(n_20358));
OAI21X1 g61997(.A0 (n_18036), .A1 (n_26903), .B0 (n_14342), .Y(n_20357));
NAND3X1 g62003(.A (n_15003), .B (n_18071), .C (n_19947), .Y(n_20353));
NAND4X1 g62021(.A (n_14123), .B (n_14252), .C (n_19957), .D(n_16926), .Y (n_20352));
OAI21X1 g62028(.A0 (n_12290), .A1 (n_18746), .B0 (n_21275), .Y(n_20351));
NAND2X1 g62050(.A (n_18949), .B (n_19934), .Y (n_20349));
NAND2X1 g62052(.A (n_18947), .B (n_804), .Y (n_20348));
NAND2X1 g62056(.A (n_18942), .B (n_2204), .Y (n_20346));
OAI21X1 g62059(.A0 (n_11527), .A1 (n_18748), .B0 (n_171), .Y(n_20344));
NAND2X1 g62073(.A (n_18927), .B (sa01[1] ), .Y (n_20343));
OAI21X1 g62078(.A0 (n_18841), .A1 (n_26728), .B0 (n_28692), .Y(n_20341));
OAI21X1 g62080(.A0 (n_13348), .A1 (n_18747), .B0 (n_129), .Y(n_20340));
OAI21X1 g62096(.A0 (n_18764), .A1 (n_15327), .B0 (n_27216), .Y(n_20339));
OAI21X1 g62104(.A0 (n_18763), .A1 (n_15194), .B0 (n_27718), .Y(n_20338));
AOI21X1 g62105(.A0 (n_18783), .A1 (n_27313), .B0 (n_20564), .Y(n_20337));
OAI21X1 g62107(.A0 (n_18762), .A1 (n_15089), .B0 (n_17933), .Y(n_20336));
OAI21X1 g62116(.A0 (n_18761), .A1 (n_14223), .B0 (n_20680), .Y(n_20335));
OAI21X1 g62131(.A0 (n_18795), .A1 (n_11003), .B0 (n_28642), .Y(n_20334));
NAND2X1 g62135(.A (n_18899), .B (n_20332), .Y (n_20333));
NAND2X1 g62136(.A (n_18898), .B (n_27718), .Y (n_20331));
AOI21X1 g62141(.A0 (n_16854), .A1 (n_18004), .B0 (n_21055), .Y(n_20329));
AOI21X1 g62155(.A0 (n_13374), .A1 (n_17943), .B0 (n_2681), .Y(n_20328));
INVX1 g62167(.A (n_19904), .Y (n_20327));
NAND2X1 g62177(.A (n_19011), .B (n_20325), .Y (n_20326));
NAND2X1 g62185(.A (n_18998), .B (n_8708), .Y (n_20324));
XOR2X1 g59836(.A (u0_rcon_1057), .B (n_1429), .Y (n_20322));
AOI21X1 g62211(.A0 (n_15349), .A1 (n_16835), .B0 (n_18627), .Y(n_28270));
NOR2X1 g62233(.A (n_18938), .B (n_20204), .Y (n_20319));
NAND2X1 g62241(.A (n_19024), .B (n_16452), .Y (n_20318));
AOI21X1 g62265(.A0 (n_17985), .A1 (n_16792), .B0 (n_21055), .Y(n_20317));
NOR2X1 g62288(.A (n_18928), .B (n_20315), .Y (n_20316));
NAND3X1 g62306(.A (n_18856), .B (n_14836), .C (n_12853), .Y(n_20314));
NOR2X1 g62311(.A (n_18923), .B (n_20198), .Y (n_20313));
AOI21X1 g62351(.A0 (n_16658), .A1 (n_18833), .B0 (n_164), .Y(n_20312));
NOR3X1 g62387(.A (n_8803), .B (n_8128), .C (n_18822), .Y (n_20311));
XOR2X1 g59953(.A (u0_rcon_1055), .B (n_1158), .Y (n_20310));
XOR2X1 g59954(.A (u0_rcon_1056), .B (n_1271), .Y (n_20309));
INVX1 g59955(.A (n_20307), .Y (n_20308));
NAND2X1 g62402(.A (n_18972), .B (n_19052), .Y (n_20306));
NOR2X1 g62431(.A (n_18905), .B (n_18840), .Y (n_20305));
NAND4X1 g62460(.A (n_29208), .B (n_12834), .C (n_13701), .D(n_17805), .Y (n_20304));
NAND3X1 g62468(.A (n_19051), .B (n_17939), .C (n_16577), .Y(n_20303));
AOI22X1 g62478(.A0 (n_17942), .A1 (n_15894), .B0 (n_4427), .B1(n_6748), .Y (n_20302));
NOR2X1 g62480(.A (n_18001), .B (n_19081), .Y (n_20301));
NAND2X1 g62481(.A (n_19053), .B (n_21151), .Y (n_20300));
INVX1 g62494(.A (n_19802), .Y (n_20299));
INVX1 g62496(.A (n_19801), .Y (n_20298));
AOI21X1 g62502(.A0 (n_13067), .A1 (n_16466), .B0 (n_18921), .Y(n_20297));
AOI21X1 g62508(.A0 (n_6294), .A1 (n_7579), .B0 (n_18896), .Y(n_20295));
AOI21X1 g62515(.A0 (n_11208), .A1 (n_18369), .B0 (n_18932), .Y(n_20294));
NOR2X1 g62516(.A (n_17983), .B (n_19070), .Y (n_20293));
AOI21X1 g62519(.A0 (n_15156), .A1 (n_4582), .B0 (n_18931), .Y(n_20292));
OAI21X1 g62534(.A0 (n_18796), .A1 (n_3910), .B0 (n_16794), .Y(n_20290));
NOR2X1 g62544(.A (n_19007), .B (n_11488), .Y (n_20289));
AOI21X1 g62548(.A0 (n_18781), .A1 (n_15039), .B0 (n_16744), .Y(n_20288));
AOI21X1 g62549(.A0 (n_18780), .A1 (n_29102), .B0 (n_15081), .Y(n_20287));
NAND2X1 g62552(.A (n_19050), .B (n_20648), .Y (n_20286));
NAND2X1 g62554(.A (n_19049), .B (n_28170), .Y (n_20285));
AOI21X1 g62580(.A0 (n_18793), .A1 (n_10794), .B0 (n_19795), .Y(n_20282));
INVX1 g62582(.A (n_19770), .Y (n_20281));
NAND2X1 g62588(.A (n_18881), .B (n_18295), .Y (n_20279));
NOR2X1 g62589(.A (n_18870), .B (n_17122), .Y (n_20278));
NAND2X1 g62591(.A (n_19047), .B (n_20564), .Y (n_20277));
NOR2X1 g62592(.A (n_18869), .B (n_17119), .Y (n_29126));
INVX1 g62595(.A (n_19766), .Y (n_20275));
NOR2X1 g62598(.A (n_18868), .B (n_18239), .Y (n_20274));
INVX1 g62614(.A (n_19757), .Y (n_20273));
OAI21X1 g62640(.A0 (n_17975), .A1 (n_10197), .B0 (n_20271), .Y(n_20272));
OAI21X1 g62653(.A0 (n_18819), .A1 (n_10149), .B0 (n_20269), .Y(n_20270));
OAI21X1 g62655(.A0 (n_18812), .A1 (n_8590), .B0 (n_20065), .Y(n_20268));
AOI22X1 g62666(.A0 (n_18766), .A1 (n_20153), .B0 (n_10837), .B1(n_21598), .Y (n_20267));
NAND2X1 g62676(.A (n_13719), .B (n_19039), .Y (n_20266));
NAND2X1 g62684(.A (n_18289), .B (n_18980), .Y (n_20265));
NOR2X1 g62686(.A (n_29401), .B (n_29400), .Y (n_20264));
NAND2X1 g62687(.A (n_18975), .B (n_18974), .Y (n_20263));
NOR2X1 g62690(.A (n_17860), .B (n_19059), .Y (n_20262));
NOR2X1 g62694(.A (n_16778), .B (n_19083), .Y (n_20261));
NAND2X1 g62719(.A (n_7165), .B (n_18955), .Y (n_20260));
OAI21X1 g62721(.A0 (n_18760), .A1 (n_15574), .B0 (n_7688), .Y(n_20259));
NAND2X1 g62727(.A (n_8322), .B (n_18954), .Y (n_20258));
NAND2X1 g62730(.A (n_17636), .B (n_19094), .Y (n_20257));
AOI22X1 g62737(.A0 (n_18750), .A1 (n_17411), .B0 (n_12085), .B1(n_11731), .Y (n_20256));
AOI22X1 g62742(.A0 (n_18751), .A1 (n_29048), .B0 (n_12303), .B1(n_4689), .Y (n_25467));
NAND2X1 g62788(.A (n_19025), .B (n_18506), .Y (n_20251));
AOI21X1 g62789(.A0 (n_16789), .A1 (n_12986), .B0 (n_19016), .Y(n_20250));
INVX1 g62792(.A (n_19708), .Y (n_20248));
AOI21X1 g62795(.A0 (n_17907), .A1 (n_27688), .B0 (n_18992), .Y(n_20247));
AOI21X1 g62796(.A0 (n_16629), .A1 (n_28642), .B0 (n_18988), .Y(n_20246));
OR2X1 g62833(.A (n_19590), .B (n_21275), .Y (n_20245));
OR2X1 g62886(.A (n_19593), .B (n_20729), .Y (n_20243));
NAND3X1 g63051(.A (n_17235), .B (n_9508), .C (n_18745), .Y (n_25580));
OAI21X1 g63064(.A0 (n_20239), .A1 (n_28274), .B0 (n_1196), .Y(n_20240));
INVX1 g63088(.A (n_19683), .Y (n_20237));
NAND3X1 g63129(.A (n_18391), .B (n_9397), .C (n_18741), .Y (n_20236));
NAND2X1 g73100(.A (n_18864), .B (n_19755), .Y (n_20234));
INVX1 g63237(.A (n_19678), .Y (n_20233));
AOI21X1 g63289(.A0 (n_10962), .A1 (n_18688), .B0 (n_17414), .Y(n_20232));
AOI21X1 g63337(.A0 (n_10911), .A1 (n_18690), .B0 (n_15574), .Y(n_20230));
OAI21X1 g63340(.A0 (n_18732), .A1 (n_28138), .B0 (n_2909), .Y(n_20229));
AOI21X1 g63344(.A0 (n_18731), .A1 (n_17752), .B0 (n_9084), .Y(n_20227));
NAND2X1 g63470(.A (n_19582), .B (n_13801), .Y (n_20226));
NAND2X1 g63471(.A (n_18853), .B (n_19934), .Y (n_20225));
NAND2X1 g63582(.A (n_18855), .B (n_5131), .Y (n_20222));
AOI22X1 g60564(.A0 (n_18782), .A1 (n_124), .B0 (n_18254), .B1(n_4582), .Y (n_20221));
OAI21X1 g63763(.A0 (n_19781), .A1 (n_1310), .B0 (n_21210), .Y(n_20219));
AOI21X1 g63839(.A0 (n_10700), .A1 (n_3301), .B0 (n_18850), .Y(n_20218));
OAI21X1 g63870(.A0 (n_18683), .A1 (n_12872), .B0 (n_20760), .Y(n_20217));
AOI21X1 g63908(.A0 (n_12468), .A1 (n_16835), .B0 (n_19583), .Y(n_20216));
NAND2X1 g64028(.A (n_16841), .B (n_18848), .Y (n_20215));
NAND2X1 g60742(.A (n_19567), .B (n_20213), .Y (n_20214));
OAI21X1 g60782(.A0 (n_18698), .A1 (n_14518), .B0 (n_20018), .Y(n_20212));
AOI21X1 g60786(.A0 (n_18696), .A1 (n_11064), .B0 (n_663), .Y(n_20211));
OAI21X1 g60800(.A0 (n_18692), .A1 (n_12350), .B0 (n_19475), .Y(n_20208));
NAND4X1 g60852(.A (n_7252), .B (n_14722), .C (n_17544), .D (n_13094),.Y (n_20206));
NAND2X1 g60885(.A (n_19573), .B (n_20204), .Y (n_20205));
NOR2X1 g60906(.A (n_11407), .B (n_19599), .Y (n_20203));
OAI21X1 g60910(.A0 (n_18713), .A1 (n_17472), .B0 (n_20055), .Y(n_20202));
NAND2X1 g60914(.A (n_19572), .B (n_20518), .Y (n_20200));
NAND2X1 g60933(.A (n_19571), .B (n_20198), .Y (n_20199));
NAND2X1 g60942(.A (n_19570), .B (n_20648), .Y (n_20197));
OAI21X1 g60947(.A0 (n_18709), .A1 (n_17034), .B0 (n_19995), .Y(n_20195));
NAND4X1 g60976(.A (n_20192), .B (n_14619), .C (n_17545), .D(n_16183), .Y (n_20193));
NOR2X1 g60979(.A (n_19596), .B (n_18641), .Y (n_20191));
NAND4X1 g61081(.A (n_8411), .B (n_11371), .C (n_16832), .D (n_15798),.Y (n_20190));
OAI21X1 g61132(.A0 (n_17519), .A1 (n_3612), .B0 (n_15731), .Y(n_20189));
OAI21X1 g61134(.A0 (n_17506), .A1 (n_624), .B0 (n_15734), .Y(n_20188));
OAI21X1 g61135(.A0 (n_17505), .A1 (n_2001), .B0 (n_15733), .Y(n_20187));
OAI21X1 g61136(.A0 (n_17504), .A1 (n_1756), .B0 (n_15732), .Y(n_20186));
NAND4X1 g61153(.A (n_9261), .B (n_14985), .C (n_12271), .D (n_15611),.Y (n_20185));
AOI21X1 g61158(.A0 (n_17532), .A1 (n_18679), .B0 (n_18194), .Y(n_20184));
NAND2X1 g65408(.A (n_18718), .B (n_19966), .Y (n_20183));
AOI21X1 g61160(.A0 (n_17510), .A1 (n_17912), .B0 (n_11643), .Y(n_20182));
AOI21X1 g61161(.A0 (n_17509), .A1 (n_16754), .B0 (n_15533), .Y(n_20181));
OAI21X1 g61165(.A0 (n_17894), .A1 (n_14807), .B0 (n_18723), .Y(n_20180));
OR4X1 g61177(.A (n_20178), .B (n_11230), .C (n_7629), .D (n_15559),.Y (n_20179));
NAND4X1 g61179(.A (n_12796), .B (n_12829), .C (n_7552), .D (n_15699),.Y (n_20177));
AND2X1 g65468(.A (n_18714), .B (n_13291), .Y (n_20176));
NAND2X1 g61187(.A (n_18699), .B (n_869), .Y (n_20175));
OAI21X1 g61248(.A0 (n_15110), .A1 (n_17495), .B0 (sa32[1] ), .Y(n_20173));
NAND2X1 g65704(.A (n_18738), .B (n_14800), .Y (n_20172));
NAND4X1 g61287(.A (n_27560), .B (n_16640), .C (n_20169), .D(n_15608), .Y (n_20171));
NAND3X1 g61288(.A (n_10087), .B (n_17562), .C (n_15689), .Y(n_20168));
NAND2X1 g65800(.A (n_18711), .B (n_19964), .Y (n_29423));
INVX1 g65803(.A (n_19581), .Y (n_20166));
NAND4X1 g61383(.A (n_17901), .B (n_17902), .C (n_13803), .D(n_14796), .Y (n_20165));
OAI21X1 g61391(.A0 (n_17484), .A1 (w3[17] ), .B0 (n_18096), .Y(n_20164));
OAI21X1 g61394(.A0 (n_17480), .A1 (n_20162), .B0 (n_18081), .Y(n_20163));
NAND4X1 g61424(.A (n_29420), .B (n_13093), .C (n_29421), .D(n_13074), .Y (n_20161));
NAND4X1 g61429(.A (n_29312), .B (n_13043), .C (n_29313), .D(n_13004), .Y (n_28605));
AOI21X1 g61435(.A0 (n_17448), .A1 (n_20157), .B0 (n_18674), .Y(n_20158));
AOI21X1 g61449(.A0 (n_17462), .A1 (n_17423), .B0 (n_11580), .Y(n_20156));
NAND4X1 g61450(.A (n_11551), .B (n_18633), .C (n_15761), .D (n_6457),.Y (n_20155));
AOI22X1 g61452(.A0 (n_17486), .A1 (n_20153), .B0 (n_16176), .B1(n_20010), .Y (n_20154));
AOI22X1 g61457(.A0 (n_17482), .A1 (w3[17] ), .B0 (n_13022), .B1(n_19310), .Y (n_20152));
NAND4X1 g61466(.A (n_15006), .B (n_15326), .C (n_15786), .D(n_12920), .Y (n_28606));
NAND4X1 g61479(.A (n_13309), .B (n_15087), .C (n_15780), .D(n_11242), .Y (n_20150));
NAND4X1 g61481(.A (n_29390), .B (n_27135), .C (n_29391), .D(n_16228), .Y (n_20149));
OAI21X1 g61505(.A0 (n_17458), .A1 (n_20068), .B0 (n_18704), .Y(n_20148));
OAI21X1 g61514(.A0 (n_16561), .A1 (n_17116), .B0 (n_20144), .Y(n_20145));
NAND2X1 g61516(.A (n_18516), .B (n_124), .Y (n_20143));
OAI21X1 g61517(.A0 (n_25785), .A1 (n_25786), .B0 (n_310), .Y(n_20141));
OAI21X1 g61519(.A0 (n_16686), .A1 (n_17133), .B0 (n_129), .Y(n_20140));
OAI21X1 g61526(.A0 (n_29432), .A1 (n_29433), .B0 (sa31[1] ), .Y(n_20138));
OAI21X1 g61528(.A0 (n_17106), .A1 (n_14261), .B0 (n_14627), .Y(n_20137));
OAI21X1 g61530(.A0 (n_15514), .A1 (n_17196), .B0 (n_20198), .Y(n_20135));
OAI21X1 g61532(.A0 (n_17108), .A1 (n_17617), .B0 (n_21174), .Y(n_20134));
OAI21X1 g61533(.A0 (n_17326), .A1 (n_13242), .B0 (n_20587), .Y(n_20133));
OAI21X1 g61534(.A0 (n_17065), .A1 (n_14678), .B0 (n_1196), .Y(n_20132));
OAI21X1 g61535(.A0 (n_17259), .A1 (n_11569), .B0 (n_20558), .Y(n_20130));
OAI21X1 g61537(.A0 (n_17213), .A1 (n_13182), .B0 (n_3538), .Y(n_28893));
OAI21X1 g61540(.A0 (n_17036), .A1 (n_14638), .B0 (n_21242), .Y(n_20128));
AND2X1 g61544(.A (n_18632), .B (n_16301), .Y (n_20127));
AOI21X1 g61556(.A0 (n_17622), .A1 (n_15727), .B0 (n_15894), .Y(n_20126));
OAI21X1 g61566(.A0 (n_17366), .A1 (n_1756), .B0 (n_12282), .Y(n_20124));
NOR3X1 g61571(.A (n_12518), .B (n_5859), .C (n_17395), .Y (n_20123));
AOI21X1 g61573(.A0 (n_17641), .A1 (n_17349), .B0 (n_14155), .Y(n_20122));
OAI21X1 g61581(.A0 (n_17385), .A1 (n_14881), .B0 (sa13[1] ), .Y(n_20121));
OAI21X1 g61582(.A0 (n_17384), .A1 (n_17724), .B0 (n_1991), .Y(n_20120));
OAI21X1 g61583(.A0 (n_17383), .A1 (n_16486), .B0 (sa20[1] ), .Y(n_20119));
NAND2X1 g61585(.A (n_18636), .B (n_16480), .Y (n_20118));
OAI21X1 g61586(.A0 (n_17380), .A1 (n_14865), .B0 (n_20116), .Y(n_20117));
OAI21X1 g61591(.A0 (n_17373), .A1 (n_17777), .B0 (n_903), .Y(n_20115));
OAI21X1 g61593(.A0 (n_17367), .A1 (n_13184), .B0 (sa10[1] ), .Y(n_20113));
OAI21X1 g61597(.A0 (n_17362), .A1 (n_16352), .B0 (n_20767), .Y(n_20112));
OAI21X1 g61598(.A0 (n_17360), .A1 (n_13151), .B0 (n_20574), .Y(n_20111));
OAI21X1 g61599(.A0 (n_17374), .A1 (n_16347), .B0 (sa23[1] ), .Y(n_20110));
AOI21X1 g61604(.A0 (n_15357), .A1 (n_17142), .B0 (n_123), .Y(n_20109));
NAND4X1 g61605(.A (n_11179), .B (n_19097), .C (n_15359), .D(n_13098), .Y (n_20108));
AOI22X1 g61607(.A0 (n_17093), .A1 (n_1196), .B0 (n_8755), .B1(n_20105), .Y (n_20107));
NAND3X1 g61609(.A (n_14895), .B (n_12440), .C (n_17341), .Y(n_20104));
AOI22X1 g61611(.A0 (n_17092), .A1 (n_20102), .B0 (n_8348), .B1(n_20269), .Y (n_20103));
NAND3X1 g61615(.A (n_10137), .B (n_17090), .C (n_16334), .Y(n_20101));
NAND2X1 g61622(.A (n_18569), .B (n_20412), .Y (n_20100));
AOI21X1 g61626(.A0 (n_17327), .A1 (n_11516), .B0 (n_4582), .Y(n_20099));
NAND3X1 g61631(.A (n_18642), .B (n_13524), .C (n_14922), .Y(n_20098));
NAND4X1 g61632(.A (n_20096), .B (n_28580), .C (n_15073), .D(n_12959), .Y (n_20097));
AOI21X1 g61635(.A0 (n_15181), .A1 (n_17138), .B0 (n_20018), .Y(n_20095));
AOI21X1 g61638(.A0 (n_17141), .A1 (n_196), .B0 (n_17096), .Y(n_20093));
AOI21X1 g61645(.A0 (n_17255), .A1 (n_14512), .B0 (n_13083), .Y(n_20092));
AOI21X1 g61646(.A0 (n_17114), .A1 (n_16466), .B0 (n_11439), .Y(n_20091));
NAND4X1 g61650(.A (n_25460), .B (n_17297), .C (n_12209), .D(n_11228), .Y (n_20089));
NAND4X1 g61652(.A (n_11060), .B (n_19095), .C (n_15171), .D(n_13032), .Y (n_20088));
NAND4X1 g61654(.A (n_18046), .B (n_15692), .C (n_9309), .D (n_16689),.Y (n_20087));
NAND3X1 g61657(.A (n_16732), .B (n_17082), .C (n_16880), .Y(n_20085));
NAND4X1 g61658(.A (n_11151), .B (n_17021), .C (n_15694), .D(n_14786), .Y (n_20084));
NAND3X1 g61666(.A (n_25803), .B (n_12676), .C (n_25804), .Y(n_20083));
NAND3X1 g61667(.A (n_14131), .B (n_6945), .C (n_17354), .Y (n_20082));
AOI21X1 g61674(.A0 (n_17173), .A1 (n_14493), .B0 (n_13606), .Y(n_20081));
AND2X1 g61680(.A (n_18626), .B (n_15231), .Y (n_20080));
NAND4X1 g61681(.A (n_20078), .B (n_8293), .C (n_9340), .D (n_15229),.Y (n_20079));
AOI21X1 g61683(.A0 (n_13750), .A1 (n_18369), .B0 (n_18654), .Y(n_20077));
NAND2X1 g61685(.A (n_18517), .B (n_18203), .Y (n_20075));
NAND3X1 g61686(.A (n_12625), .B (n_17789), .C (n_17388), .Y(n_20074));
NAND3X1 g61689(.A (n_12673), .B (n_17118), .C (n_17687), .Y(n_20073));
NAND4X1 g61692(.A (n_28594), .B (n_16271), .C (n_16812), .D(n_12907), .Y (n_20072));
AOI21X1 g61695(.A0 (n_13742), .A1 (n_4582), .B0 (n_18652), .Y(n_20071));
NAND2X1 g61704(.A (n_18558), .B (n_20068), .Y (n_29422));
AOI22X1 g61713(.A0 (n_17094), .A1 (n_19414), .B0 (n_6835), .B1(n_20065), .Y (n_20066));
NAND3X1 g61715(.A (n_11030), .B (n_17794), .C (n_13814), .Y(n_20064));
NAND4X1 g61718(.A (n_20062), .B (n_12224), .C (n_15356), .D(n_12911), .Y (n_20063));
OAI21X1 g61719(.A0 (n_17358), .A1 (n_8423), .B0 (n_21487), .Y(n_20061));
OAI21X1 g61723(.A0 (n_17363), .A1 (n_12871), .B0 (n_3538), .Y(n_20060));
NOR2X1 g61724(.A (n_10733), .B (n_18673), .Y (n_20059));
NAND3X1 g61730(.A (n_16046), .B (n_11865), .C (n_17399), .Y(n_20058));
NAND3X1 g61734(.A (n_10830), .B (n_9940), .C (n_17107), .Y (n_20057));
OAI21X1 g61739(.A0 (n_17369), .A1 (n_8469), .B0 (n_20055), .Y(n_20056));
AOI22X1 g61743(.A0 (n_17057), .A1 (n_21242), .B0 (n_9922), .B1(n_19752), .Y (n_20054));
NAND3X1 g61748(.A (n_25768), .B (n_17765), .C (n_25769), .Y(n_20053));
NAND2X1 g61753(.A (n_18554), .B (n_28170), .Y (n_20052));
NAND3X1 g61757(.A (n_14285), .B (n_16400), .C (n_17387), .Y(n_20050));
NAND2X1 g61767(.A (n_18557), .B (n_14854), .Y (n_20049));
NAND3X1 g61770(.A (n_13342), .B (n_17746), .C (n_13731), .Y(n_20047));
NAND3X1 g61772(.A (n_10910), .B (n_17747), .C (n_15759), .Y(n_20046));
OAI21X1 g61774(.A0 (n_15010), .A1 (n_17364), .B0 (n_20055), .Y(n_20045));
INVX1 g61778(.A (n_19484), .Y (n_20044));
NAND3X1 g61781(.A (n_14228), .B (n_17741), .C (n_15758), .Y(n_20043));
NAND2X1 g61783(.A (n_18551), .B (n_20041), .Y (n_20042));
OAI21X1 g61786(.A0 (n_13330), .A1 (n_17201), .B0 (n_29039), .Y(n_20040));
NAND3X1 g61787(.A (n_12439), .B (n_17737), .C (n_13805), .Y(n_20039));
NOR3X1 g61789(.A (n_5160), .B (n_9931), .C (n_17105), .Y (n_20038));
NAND2X1 g61796(.A (n_18546), .B (n_20767), .Y (n_20036));
NAND2X1 g61803(.A (n_18545), .B (n_13176), .Y (n_20034));
NAND3X1 g61804(.A (n_12797), .B (n_17719), .C (n_15752), .Y(n_20033));
NAND2X1 g61807(.A (n_18579), .B (n_19924), .Y (n_25542));
INVX1 g61809(.A (n_19477), .Y (n_20031));
NAND2X1 g61813(.A (n_18512), .B (n_14741), .Y (n_20030));
AOI22X1 g61822(.A0 (n_17026), .A1 (n_21055), .B0 (n_8449), .B1(n_20271), .Y (n_20029));
OAI21X1 g61825(.A0 (n_17159), .A1 (n_14537), .B0 (n_638), .Y(n_20027));
INVX1 g61828(.A (n_19469), .Y (n_28509));
NOR2X1 g61837(.A (n_14839), .B (n_18613), .Y (n_25635));
NAND4X1 g61839(.A (n_11883), .B (n_16031), .C (n_20023), .D(n_16282), .Y (n_20024));
OAI21X1 g61843(.A0 (n_17318), .A1 (n_8163), .B0 (n_21314), .Y(n_20022));
OAI21X1 g61844(.A0 (n_17339), .A1 (n_17467), .B0 (n_19981), .Y(n_20021));
NAND2X1 g61845(.A (n_18649), .B (n_20116), .Y (n_20020));
AOI21X1 g61848(.A0 (n_11073), .A1 (n_20018), .B0 (n_27655), .Y(n_20019));
OAI21X1 g61849(.A0 (n_17323), .A1 (n_17465), .B0 (n_19834), .Y(n_20017));
AOI21X1 g61850(.A0 (n_16964), .A1 (w3[1] ), .B0 (n_13234), .Y(n_20016));
AOI21X1 g61851(.A0 (n_17322), .A1 (n_19433), .B0 (n_18347), .Y(n_20015));
NAND4X1 g61855(.A (n_12789), .B (n_20013), .C (n_21659), .D(n_15430), .Y (n_20014));
NAND4X1 g61859(.A (n_13496), .B (n_14935), .C (n_12746), .D(n_15386), .Y (n_20012));
AOI21X1 g61861(.A0 (n_17304), .A1 (n_20010), .B0 (n_11233), .Y(n_20011));
AOI22X1 g61866(.A0 (n_17291), .A1 (n_13466), .B0 (n_5025), .B1(n_18792), .Y (n_20009));
AOI21X1 g61868(.A0 (n_17251), .A1 (n_1667), .B0 (n_10724), .Y(n_20008));
AOI21X1 g61875(.A0 (n_17275), .A1 (n_15655), .B0 (n_9459), .Y(n_20007));
AOI21X1 g61877(.A0 (n_17073), .A1 (n_17274), .B0 (n_16978), .Y(n_20005));
AOI21X1 g61878(.A0 (n_16943), .A1 (n_20003), .B0 (n_21314), .Y(n_20004));
NAND4X1 g61884(.A (n_15413), .B (n_7470), .C (n_16526), .D (n_13425),.Y (n_20002));
OAI21X1 g61886(.A0 (n_17244), .A1 (n_19186), .B0 (n_21242), .Y(n_20001));
AOI21X1 g61902(.A0 (n_16940), .A1 (n_14949), .B0 (n_20517), .Y(n_20000));
OAI21X1 g61906(.A0 (n_16937), .A1 (n_13008), .B0 (n_778), .Y(n_19999));
NAND2X1 g61909(.A (n_18110), .B (n_18592), .Y (n_19998));
OAI21X1 g61914(.A0 (n_17182), .A1 (n_17477), .B0 (n_1397), .Y(n_19997));
OAI21X1 g61916(.A0 (n_16936), .A1 (n_11303), .B0 (n_19995), .Y(n_19996));
NAND2X1 g61920(.A (n_18588), .B (sa01[1] ), .Y (n_19994));
NAND2X1 g61923(.A (n_18584), .B (n_20862), .Y (n_19993));
NAND2X1 g61927(.A (n_18583), .B (n_19934), .Y (n_19992));
NOR2X1 g61929(.A (n_11195), .B (n_18581), .Y (n_19991));
NOR2X1 g61936(.A (n_13596), .B (n_18689), .Y (n_19990));
AOI22X1 g61938(.A0 (n_16960), .A1 (n_1667), .B0 (n_12520), .B1(n_15674), .Y (n_19989));
AOI22X1 g61941(.A0 (n_16958), .A1 (n_1132), .B0 (n_12658), .B1(n_4582), .Y (n_19987));
AOI22X1 g61942(.A0 (n_16965), .A1 (n_638), .B0 (n_16067), .B1(n_15894), .Y (n_19985));
INVX1 g61944(.A (n_19444), .Y (n_19983));
AOI22X1 g61946(.A0 (n_17060), .A1 (n_19981), .B0 (n_17211), .B1(n_9819), .Y (n_19982));
INVX1 g61948(.A (n_19443), .Y (n_19980));
NOR2X1 g61950(.A (n_13587), .B (n_18687), .Y (n_19979));
INVX1 g61952(.A (n_19442), .Y (n_25497));
AOI21X1 g61960(.A0 (n_16950), .A1 (n_26271), .B0 (n_16616), .Y(n_19976));
AOI22X1 g61961(.A0 (n_16949), .A1 (n_3910), .B0 (n_12869), .B1(n_17411), .Y (n_19974));
AOI22X1 g61962(.A0 (n_16948), .A1 (n_1295), .B0 (n_15955), .B1(n_263), .Y (n_19971));
AOI21X1 g61968(.A0 (n_17298), .A1 (n_1547), .B0 (n_13672), .Y(n_19969));
AOI21X1 g61970(.A0 (n_17242), .A1 (n_5329), .B0 (n_13666), .Y(n_19968));
AOI21X1 g61978(.A0 (n_19966), .A1 (n_10348), .B0 (n_18644), .Y(n_19967));
AOI21X1 g61982(.A0 (n_19964), .A1 (n_10249), .B0 (n_18618), .Y(n_19965));
AOI22X1 g61983(.A0 (n_17226), .A1 (n_3168), .B0 (n_17760), .B1(n_10515), .Y (n_19963));
NAND4X1 g61985(.A (n_12814), .B (n_17266), .C (n_11615), .D(n_15466), .Y (n_19960));
NAND3X1 g61995(.A (n_13455), .B (n_16972), .C (n_19417), .Y(n_19959));
NAND3X1 g62001(.A (n_15044), .B (n_16968), .C (n_19957), .Y(n_19958));
NAND3X1 g62008(.A (n_9304), .B (n_17081), .C (n_19955), .Y (n_19956));
NAND3X1 g62009(.A (n_9341), .B (n_17077), .C (n_19953), .Y (n_19954));
NAND3X1 g62011(.A (n_11142), .B (n_17068), .C (n_19951), .Y(n_19952));
NAND4X1 g62013(.A (n_14396), .B (n_12718), .C (n_19949), .D(n_15457), .Y (n_19950));
NAND4X1 g62018(.A (n_15945), .B (n_14344), .C (n_19947), .D(n_15453), .Y (n_19948));
NAND2X1 g62029(.A (n_18070), .B (n_21055), .Y (n_19946));
NAND2X1 g62031(.A (n_18067), .B (n_20041), .Y (n_19945));
OAI21X1 g62033(.A0 (n_14416), .A1 (n_17678), .B0 (n_21314), .Y(n_19944));
AOI21X1 g62035(.A0 (n_16529), .A1 (n_16850), .B0 (n_19942), .Y(n_19943));
NAND2X1 g62038(.A (n_18253), .B (n_19940), .Y (n_19941));
NAND2X1 g62039(.A (n_18057), .B (n_20102), .Y (n_19939));
AOI21X1 g62040(.A0 (n_12528), .A1 (n_16896), .B0 (n_903), .Y(n_19938));
OAI21X1 g62041(.A0 (n_14298), .A1 (n_17677), .B0 (n_21133), .Y(n_19937));
AOI21X1 g62044(.A0 (n_29387), .A1 (n_29388), .B0 (sa01[1] ), .Y(n_19936));
AOI21X1 g62045(.A0 (n_16840), .A1 (n_17854), .B0 (n_19934), .Y(n_19935));
NAND2X1 g62047(.A (n_18130), .B (n_933), .Y (n_19933));
NAND2X1 g62048(.A (n_18193), .B (n_124), .Y (n_19932));
INVX1 g62057(.A (n_19405), .Y (n_19931));
INVX1 g62061(.A (n_19402), .Y (n_19930));
OAI21X1 g62063(.A0 (n_16513), .A1 (n_17680), .B0 (n_21055), .Y(n_19929));
OAI21X1 g62074(.A0 (n_13373), .A1 (n_17679), .B0 (n_27045), .Y(n_19928));
NAND2X1 g62088(.A (n_18143), .B (sa22[1] ), .Y (n_19927));
NAND2X1 g62090(.A (n_18138), .B (n_19924), .Y (n_19925));
OAI21X1 g62097(.A0 (n_17701), .A1 (n_13510), .B0 (n_933), .Y(n_19923));
AOI21X1 g62100(.A0 (n_17715), .A1 (n_19709), .B0 (n_21151), .Y(n_19922));
AOI21X1 g62101(.A0 (n_17799), .A1 (n_13071), .B0 (n_20587), .Y(n_19921));
OAI21X1 g62102(.A0 (n_17700), .A1 (n_11531), .B0 (n_3264), .Y(n_19920));
OAI21X1 g62109(.A0 (n_17764), .A1 (n_14662), .B0 (n_20102), .Y(n_19918));
AOI21X1 g62111(.A0 (n_17759), .A1 (n_28064), .B0 (sa12[1] ), .Y(n_19917));
OAI21X1 g62113(.A0 (n_17745), .A1 (n_16207), .B0 (n_19486), .Y(n_25734));
AOI21X1 g62114(.A0 (n_17740), .A1 (n_19711), .B0 (n_28170), .Y(n_19915));
NAND2X1 g62115(.A (n_18311), .B (n_21396), .Y (n_19914));
OAI21X1 g62117(.A0 (n_17552), .A1 (n_17702), .B0 (n_21055), .Y(n_25719));
NAND2X1 g62139(.A (n_18042), .B (sa31[1] ), .Y (n_19911));
NAND2X1 g62146(.A (n_18040), .B (n_20198), .Y (n_19910));
AOI21X1 g62147(.A0 (n_17858), .A1 (n_14914), .B0 (n_19908), .Y(n_19909));
NAND2X1 g62162(.A (n_18409), .B (n_12986), .Y (n_29415));
XOR2X1 g68817(.A (n_1237), .B (n_16939), .Y (n_19905));
AOI21X1 g62168(.A0 (n_16820), .A1 (n_12752), .B0 (n_20010), .Y(n_19904));
NAND2X1 g62170(.A (n_18390), .B (n_15894), .Y (n_19902));
OAI21X1 g62171(.A0 (n_16800), .A1 (n_19889), .B0 (n_12298), .Y(n_19901));
XOR2X1 g68829(.A (n_1127), .B (n_16922), .Y (n_19900));
NAND2X1 g62173(.A (n_18287), .B (n_19364), .Y (n_25624));
NAND2X1 g62176(.A (n_18354), .B (n_16434), .Y (n_19898));
NAND2X1 g62181(.A (n_18336), .B (n_19896), .Y (n_19897));
INVX1 g62183(.A (n_19341), .Y (n_19895));
NAND2X1 g62191(.A (n_18269), .B (n_11261), .Y (n_19893));
INVX1 g62213(.A (n_19329), .Y (n_19887));
OR2X1 g62215(.A (n_18228), .B (n_27160), .Y (n_19886));
NOR2X1 g62216(.A (n_18225), .B (n_16849), .Y (n_19885));
NAND2X1 g62221(.A (n_18221), .B (n_2826), .Y (n_19884));
NAND2X1 g62234(.A (n_18211), .B (n_933), .Y (n_19882));
OAI21X1 g62235(.A0 (n_16807), .A1 (n_19880), .B0 (n_378), .Y(n_19881));
INVX1 g62243(.A (n_19318), .Y (n_19878));
OAI21X1 g62246(.A0 (n_15239), .A1 (n_17763), .B0 (n_1000), .Y(n_19877));
OAI21X1 g62248(.A0 (n_25725), .A1 (n_25726), .B0 (n_123), .Y(n_19875));
NOR2X1 g62250(.A (n_18376), .B (n_16931), .Y (n_19873));
OR2X1 g62253(.A (n_18204), .B (n_20632), .Y (n_19872));
NAND2X1 g62255(.A (n_18202), .B (n_27100), .Y (n_25837));
AOI21X1 g62261(.A0 (n_28559), .A1 (n_28560), .B0 (n_27216), .Y(n_19870));
OR2X1 g62266(.A (n_18195), .B (n_27028), .Y (n_19869));
AND2X1 g62267(.A (n_18141), .B (n_13752), .Y (n_19868));
NAND2X1 g62276(.A (n_18045), .B (n_2981), .Y (n_19867));
AOI21X1 g62286(.A0 (n_17820), .A1 (n_12827), .B0 (n_11125), .Y(n_19866));
NOR2X1 g62289(.A (n_18059), .B (n_1196), .Y (n_19864));
NOR2X1 g62299(.A (n_18206), .B (n_19862), .Y (n_19863));
OAI21X1 g62305(.A0 (n_16759), .A1 (n_16422), .B0 (n_624), .Y(n_19860));
AOI21X1 g62307(.A0 (n_15125), .A1 (n_19857), .B0 (n_17956), .Y(n_28552));
NAND3X1 g62309(.A (n_13310), .B (n_17607), .C (n_17955), .Y(n_19856));
OAI21X1 g62313(.A0 (n_16748), .A1 (n_19854), .B0 (n_20018), .Y(n_19855));
NAND2X1 g62315(.A (n_18334), .B (n_19852), .Y (n_19853));
OAI21X1 g62318(.A0 (n_16746), .A1 (n_19850), .B0 (n_20102), .Y(n_19851));
INVX1 g62319(.A (n_19281), .Y (n_19848));
NAND3X1 g62321(.A (n_13381), .B (n_14826), .C (n_16742), .Y(n_19847));
NAND2X1 g62323(.A (n_18179), .B (n_27914), .Y (n_19846));
NOR2X1 g62325(.A (n_18176), .B (n_19844), .Y (n_19845));
OAI21X1 g62327(.A0 (n_17940), .A1 (n_13363), .B0 (sa11[1] ), .Y(n_19841));
NAND2X1 g62328(.A (n_18325), .B (n_25758), .Y (n_19839));
AOI21X1 g62334(.A0 (n_17927), .A1 (n_17926), .B0 (n_21275), .Y(n_19838));
NAND2X1 g62336(.A (n_18170), .B (n_18456), .Y (n_19836));
AOI21X1 g62345(.A0 (n_28313), .A1 (n_28314), .B0 (n_19834), .Y(n_19835));
NAND2X1 g62347(.A (n_18157), .B (n_26271), .Y (n_19833));
NOR2X1 g62356(.A (n_18155), .B (n_16648), .Y (n_19832));
NAND2X1 g62362(.A (n_18303), .B (n_19830), .Y (n_19831));
NAND4X1 g62378(.A (n_25526), .B (n_9715), .C (n_14194), .D (n_19499),.Y (n_19829));
NAND4X1 g62380(.A (n_29411), .B (n_7985), .C (n_19529), .D (n_11784),.Y (n_19828));
AND2X1 g62381(.A (n_18052), .B (n_16358), .Y (n_19827));
AOI21X1 g62394(.A0 (n_14950), .A1 (n_15688), .B0 (n_18818), .Y(n_25543));
XOR2X1 g59956(.A (u0_rcon_1058), .B (n_1020), .Y (n_20307));
AOI21X1 g62399(.A0 (n_15145), .A1 (n_19364), .B0 (n_13882), .Y(n_19825));
INVX1 g62404(.A (n_19246), .Y (n_19823));
NOR2X1 g62408(.A (n_18137), .B (n_17849), .Y (n_19822));
INVX1 g62409(.A (n_19244), .Y (n_19821));
AOI21X1 g62425(.A0 (n_14858), .A1 (n_11312), .B0 (n_18201), .Y(n_19819));
NOR2X1 g62428(.A (n_18152), .B (n_17996), .Y (n_19818));
NAND3X1 g62451(.A (n_17340), .B (n_17646), .C (n_18275), .Y(n_19817));
NOR2X1 g62456(.A (n_16384), .B (n_18392), .Y (n_19816));
NAND4X1 g62458(.A (n_28852), .B (n_19814), .C (n_11554), .D(n_12238), .Y (n_19815));
NAND3X1 g62466(.A (n_17249), .B (n_17616), .C (n_15531), .Y(n_19813));
NAND4X1 g62471(.A (n_25535), .B (n_18827), .C (n_19811), .D(n_10738), .Y (n_19812));
NAND4X1 g62475(.A (n_15070), .B (n_17748), .C (n_20023), .D(n_12248), .Y (n_19808));
NAND4X1 g62476(.A (n_9305), .B (n_12814), .C (n_13704), .D (n_16444),.Y (n_19807));
OAI21X1 g62477(.A0 (n_16808), .A1 (n_638), .B0 (n_15344), .Y(n_19806));
NAND2X1 g62486(.A (n_18450), .B (sa31[1] ), .Y (n_19805));
NAND3X1 g62491(.A (n_16822), .B (n_16823), .C (n_18151), .Y(n_19803));
NAND3X1 g62495(.A (n_17993), .B (n_17786), .C (n_15427), .Y(n_19802));
NAND3X1 g62497(.A (n_15265), .B (n_17811), .C (n_14150), .Y(n_19801));
AOI21X1 g62499(.A0 (n_17611), .A1 (n_19799), .B0 (n_2718), .Y(n_19800));
AOI21X1 g62503(.A0 (n_17806), .A1 (n_8465), .B0 (n_19797), .Y(n_19798));
AOI21X1 g62505(.A0 (n_17795), .A1 (n_12673), .B0 (n_19795), .Y(n_19796));
AOI21X1 g62507(.A0 (n_7441), .A1 (n_19445), .B0 (n_18049), .Y(n_19794));
NAND2X1 g62520(.A (n_16996), .B (n_18359), .Y (n_19793));
OAI21X1 g62522(.A0 (n_17749), .A1 (n_11917), .B0 (n_19791), .Y(n_28253));
AOI21X1 g62524(.A0 (n_16442), .A1 (n_16782), .B0 (n_21552), .Y(n_19790));
AOI21X1 g62525(.A0 (n_17710), .A1 (n_1132), .B0 (n_16986), .Y(n_19788));
NAND2X1 g62529(.A (n_18107), .B (n_18352), .Y (n_19787));
NAND2X1 g62530(.A (n_18438), .B (n_20579), .Y (n_19786));
NAND2X1 g62537(.A (n_18432), .B (n_20198), .Y (n_19784));
NAND3X1 g62542(.A (n_16763), .B (n_16764), .C (n_19781), .Y(n_19782));
NAND2X1 g62546(.A (n_9909), .B (n_18453), .Y (n_19780));
NAND2X1 g62547(.A (n_9915), .B (n_18451), .Y (n_19779));
NAND3X1 g62561(.A (n_17924), .B (n_17925), .C (n_18904), .Y(n_19778));
NAND2X1 g62566(.A (n_18309), .B (n_15275), .Y (n_19776));
AOI21X1 g62568(.A0 (n_17738), .A1 (n_9108), .B0 (n_16579), .Y(n_19775));
NAND3X1 g62574(.A (n_18301), .B (n_7326), .C (n_15325), .Y (n_19773));
NAND3X1 g62581(.A (n_18297), .B (n_9008), .C (n_15119), .Y (n_19771));
AOI21X1 g62583(.A0 (n_17727), .A1 (n_8069), .B0 (n_2663), .Y(n_19770));
NAND3X1 g62590(.A (n_18293), .B (n_10608), .C (n_16745), .Y(n_19767));
AOI21X1 g62596(.A0 (n_17722), .A1 (n_15132), .B0 (n_2800), .Y(n_19766));
AOI21X1 g62602(.A0 (n_7513), .A1 (n_1132), .B0 (n_18062), .Y(n_19764));
AOI21X1 g62605(.A0 (n_9069), .A1 (n_19111), .B0 (n_18065), .Y(n_19762));
NAND3X1 g62609(.A (n_16836), .B (n_16837), .C (n_12681), .Y(n_19761));
AOI21X1 g62611(.A0 (n_17834), .A1 (n_2022), .B0 (n_8795), .Y(n_19760));
NOR2X1 g62612(.A (n_10248), .B (n_18463), .Y (n_19759));
NOR2X1 g62613(.A (n_18028), .B (n_17136), .Y (n_29425));
NAND3X1 g62615(.A (n_16509), .B (n_17705), .C (n_14489), .Y(n_19757));
NAND2X1 g70759(.A (n_18024), .B (n_19755), .Y (n_19756));
NOR2X1 g62631(.A (n_18808), .B (n_15597), .Y (n_19754));
OAI21X1 g62641(.A0 (n_16766), .A1 (n_9943), .B0 (n_19752), .Y(n_19753));
OAI21X1 g62649(.A0 (n_17735), .A1 (n_10939), .B0 (n_19750), .Y(n_19751));
NAND2X1 g62654(.A (n_18276), .B (n_20760), .Y (n_19749));
OAI21X1 g62656(.A0 (n_17845), .A1 (n_8203), .B0 (n_20105), .Y(n_19748));
AOI21X1 g62665(.A0 (n_8113), .A1 (n_7194), .B0 (n_18383), .Y(n_19747));
AOI21X1 g62668(.A0 (n_6829), .A1 (n_7101), .B0 (n_18370), .Y(n_19746));
NOR2X1 g62677(.A (n_17962), .B (n_18475), .Y (n_28592));
NOR2X1 g62683(.A (n_18839), .B (n_18466), .Y (n_19743));
NOR2X1 g62695(.A (n_17847), .B (n_18464), .Y (n_19742));
INVX1 g62699(.A (n_19138), .Y (n_19741));
NOR2X1 g62705(.A (n_13364), .B (n_18252), .Y (n_19740));
NAND4X1 g62711(.A (n_12245), .B (n_17628), .C (n_18965), .D(n_18966), .Y (n_19739));
OAI21X1 g62717(.A0 (n_17698), .A1 (n_15708), .B0 (n_7040), .Y(n_19738));
OAI21X1 g62720(.A0 (n_17694), .A1 (n_18320), .B0 (n_8318), .Y(n_19737));
OAI21X1 g62724(.A0 (n_17693), .A1 (n_29048), .B0 (n_5753), .Y(n_19736));
AOI22X1 g62731(.A0 (n_17690), .A1 (n_15894), .B0 (n_10324), .B1(n_6534), .Y (n_19735));
NAND2X1 g62733(.A (n_15964), .B (n_18508), .Y (n_19732));
AOI22X1 g62735(.A0 (n_17684), .A1 (n_9527), .B0 (n_7556), .B1(n_8679), .Y (n_19731));
AOI22X1 g62736(.A0 (n_17688), .A1 (n_13606), .B0 (n_4511), .B1(n_11312), .Y (n_19730));
AOI22X1 g62739(.A0 (n_17686), .A1 (n_16480), .B0 (n_4613), .B1(n_14866), .Y (n_19727));
NAND2X1 g62740(.A (n_16065), .B (n_18500), .Y (n_19726));
AOI22X1 g62741(.A0 (n_17682), .A1 (n_18320), .B0 (n_10424), .B1(n_14484), .Y (n_19725));
OR2X1 g62744(.A (n_18823), .B (n_17183), .Y (n_19723));
AND2X1 g62746(.A (n_18351), .B (n_15777), .Y (n_19722));
AND2X1 g62748(.A (n_14545), .B (n_18404), .Y (n_19721));
NAND2X1 g71341(.A (n_18023), .B (n_8520), .Y (n_19720));
AOI21X1 g62756(.A0 (n_17819), .A1 (n_19114), .B0 (n_13097), .Y(n_19719));
AOI21X1 g62759(.A0 (n_17793), .A1 (n_19110), .B0 (n_12916), .Y(n_19718));
NAND2X1 g62769(.A (n_14374), .B (n_18339), .Y (n_19717));
AND2X1 g62774(.A (n_12339), .B (n_18274), .Y (n_19716));
AND2X1 g62775(.A (n_12274), .B (n_18259), .Y (n_19715));
NAND3X1 g62782(.A (n_28585), .B (n_16720), .C (n_19711), .Y(n_19712));
NAND3X1 g62785(.A (n_18208), .B (n_15308), .C (n_19709), .Y(n_19710));
NAND2X1 g62793(.A (n_29416), .B (n_29417), .Y (n_19708));
AOI22X1 g62794(.A0 (n_17916), .A1 (n_16835), .B0 (n_15451), .B1(n_3886), .Y (n_19707));
AOI21X1 g62804(.A0 (n_17792), .A1 (n_11417), .B0 (n_20213), .Y(n_19704));
OR2X1 g62815(.A (n_18789), .B (n_20457), .Y (n_19703));
OR2X1 g62816(.A (n_18794), .B (n_3264), .Y (n_19702));
AOI21X1 g62817(.A0 (n_16063), .A1 (n_18967), .B0 (n_21314), .Y(n_19701));
OAI21X1 g62830(.A0 (n_14288), .A1 (n_17600), .B0 (n_17414), .Y(n_19700));
OR2X1 g62852(.A (n_18754), .B (n_21174), .Y (n_25482));
OR2X1 g62854(.A (n_18753), .B (n_20862), .Y (n_19696));
OR2X1 g62855(.A (n_18752), .B (n_1196), .Y (n_25653));
AOI21X1 g62871(.A0 (n_19692), .A1 (n_4838), .B0 (n_19679), .Y(n_19693));
AOI21X1 g62924(.A0 (n_17589), .A1 (n_13370), .B0 (n_19364), .Y(n_19689));
NAND2X1 g72317(.A (n_18026), .B (n_19755), .Y (n_19688));
OR2X1 g63073(.A (n_18407), .B (n_19934), .Y (n_19687));
NOR2X1 g63075(.A (n_18758), .B (n_11391), .Y (n_19686));
NAND3X1 g63078(.A (n_18859), .B (n_18353), .C (n_15352), .Y(n_19684));
NAND2X1 g63089(.A (n_18852), .B (n_12907), .Y (n_19683));
OAI21X1 g63113(.A0 (n_17561), .A1 (n_16169), .B0 (n_12298), .Y(n_19682));
AOI21X1 g63192(.A0 (n_8903), .A1 (n_16480), .B0 (n_19679), .Y(n_19681));
AOI21X1 g63238(.A0 (n_11005), .A1 (n_17577), .B0 (n_15708), .Y(n_19678));
NAND2X1 g63239(.A (n_18802), .B (n_29062), .Y (n_25546));
OR2X1 g63247(.A (n_18784), .B (sa01[1] ), .Y (n_19676));
INVX1 g63253(.A (n_19009), .Y (n_19674));
NOR2X1 g63264(.A (n_11346), .B (n_29386), .Y (n_19673));
OAI21X1 g63268(.A0 (n_17560), .A1 (n_16225), .B0 (n_28642), .Y(n_19671));
INVX1 g63318(.A (n_19000), .Y (n_19669));
AND2X1 g63377(.A (n_18777), .B (n_29102), .Y (n_19667));
AND2X1 g63383(.A (n_18774), .B (n_1241), .Y (n_19666));
OR2X1 g63407(.A (n_18772), .B (n_2204), .Y (n_19665));
INVX1 g63411(.A (n_18983), .Y (n_19664));
NAND2X1 g63440(.A (n_18768), .B (n_15340), .Y (n_19663));
NAND2X1 g63441(.A (n_17961), .B (sa01[1] ), .Y (n_19662));
NAND3X1 g63456(.A (n_17315), .B (n_9382), .C (n_17658), .Y (n_19661));
NAND2X1 g63465(.A (n_18816), .B (n_19934), .Y (n_19660));
NAND2X1 g63494(.A (n_17996), .B (n_2204), .Y (n_19659));
OAI21X1 g63498(.A0 (n_17559), .A1 (n_16174), .B0 (n_12896), .Y(n_19658));
INVX1 g63506(.A (n_18968), .Y (n_25673));
INVX1 g63532(.A (n_18959), .Y (n_19656));
INVX1 g63607(.A (n_18943), .Y (n_19654));
NAND2X1 g63626(.A (n_17977), .B (n_15688), .Y (n_19653));
NAND3X1 g63667(.A (n_18790), .B (n_17980), .C (n_11885), .Y(n_19650));
NAND3X1 g63670(.A (n_6841), .B (n_17569), .C (n_19648), .Y (n_19649));
NAND2X1 g63675(.A (n_18828), .B (n_21174), .Y (n_28505));
NAND2X1 g63682(.A (n_17958), .B (n_9106), .Y (n_19646));
AOI21X1 g63683(.A0 (n_17555), .A1 (n_1310), .B0 (n_15128), .Y(n_19645));
OR2X1 g63684(.A (n_11493), .B (n_19643), .Y (n_19644));
NAND2X1 g63699(.A (n_15218), .B (n_18862), .Y (n_19641));
AOI22X1 g60556(.A0 (n_17788), .A1 (n_933), .B0 (n_10023), .B1(n_16466), .Y (n_19640));
NAND3X1 g63717(.A (n_29418), .B (n_29419), .C (n_19638), .Y(n_19639));
INVX1 g63734(.A (n_18912), .Y (n_19637));
NAND3X1 g63759(.A (n_17728), .B (n_19604), .C (n_13767), .Y(n_19635));
AND2X1 g63774(.A (n_18019), .B (n_7467), .Y (n_19632));
NAND2X1 g63778(.A (n_18815), .B (n_12723), .Y (n_19631));
INVX1 g63783(.A (n_18901), .Y (n_19630));
AOI21X1 g63791(.A0 (n_17625), .A1 (n_18792), .B0 (n_8828), .Y(n_19629));
AOI21X1 g63843(.A0 (n_9173), .A1 (n_13679), .B0 (n_18011), .Y(n_19628));
OAI21X1 g63871(.A0 (n_17564), .A1 (n_12617), .B0 (n_20765), .Y(n_28506));
NAND2X1 g63897(.A (n_18799), .B (n_1289), .Y (n_19626));
NAND2X1 g63917(.A (n_11871), .B (n_18845), .Y (n_19623));
MX2X1 g63940(.A (n_16172), .B (n_17446), .S0 (n_11261), .Y (n_19621));
NAND3X1 g63954(.A (n_17595), .B (n_17576), .C (n_16545), .Y(n_19620));
NOR2X1 g63974(.A (n_17889), .B (n_18825), .Y (n_19619));
NOR2X1 g63992(.A (n_15094), .B (n_17948), .Y (n_19618));
NAND3X1 g63993(.A (n_8917), .B (n_18911), .C (n_26952), .Y (n_19617));
NAND2X1 g60744(.A (n_18740), .B (n_4357), .Y (n_19614));
INVX1 g64170(.A (n_18860), .Y (n_21215));
NAND4X1 g60880(.A (n_7723), .B (n_14695), .C (n_15862), .D (n_11349),.Y (n_19612));
NAND4X1 g60917(.A (n_16000), .B (n_14663), .C (n_15857), .D(n_12985), .Y (n_19611));
NAND4X1 g60970(.A (n_13712), .B (n_12333), .C (n_17527), .D(n_15796), .Y (n_19610));
NAND4X1 g60974(.A (n_19608), .B (n_14719), .C (n_15865), .D(n_16275), .Y (n_19609));
AOI21X1 g60993(.A0 (n_17579), .A1 (n_21552), .B0 (n_12696), .Y(n_19607));
AND2X1 g64850(.A (n_19604), .B (n_19060), .Y (n_19605));
NOR2X1 g65057(.A (n_14626), .B (n_13012), .Y (n_25811));
NAND2X1 g65110(.A (n_17541), .B (n_14630), .Y (n_19602));
INVX1 g65201(.A (n_18814), .Y (n_25636));
NAND2X1 g65219(.A (n_17582), .B (n_6244), .Y (n_19600));
AOI21X1 g61124(.A0 (n_14888), .A1 (n_15791), .B0 (sa21[1] ), .Y(n_19599));
INVX1 g65298(.A (n_18806), .Y (n_19598));
NAND3X1 g65453(.A (n_9371), .B (n_13912), .C (sa00[1] ), .Y(n_19597));
AOI21X1 g61188(.A0 (n_12452), .A1 (n_15821), .B0 (n_196), .Y(n_19596));
INVX1 g65558(.A (n_18786), .Y (n_19595));
NAND3X1 g65573(.A (n_12624), .B (n_16005), .C (sa01[1] ), .Y(n_19594));
AND2X1 g65577(.A (n_17609), .B (n_11452), .Y (n_19593));
AND2X1 g65633(.A (n_17626), .B (n_13305), .Y (n_19592));
OR4X1 g61249(.A (n_9903), .B (n_11280), .C (n_7843), .D (n_13710), .Y(n_19591));
AOI21X1 g65648(.A0 (n_14128), .A1 (n_523), .B0 (n_17599), .Y(n_19590));
NAND2X1 g65670(.A (n_17587), .B (n_14266), .Y (n_19589));
INVX1 g65672(.A (n_18779), .Y (n_19588));
OR4X1 g61271(.A (n_16300), .B (n_9405), .C (n_11050), .D (n_13709),.Y (n_19587));
INVX1 g65718(.A (n_18773), .Y (n_19586));
INVX1 g65736(.A (n_18771), .Y (n_19585));
AOI21X1 g65745(.A0 (n_15848), .A1 (n_9930), .B0 (n_16835), .Y(n_19583));
NOR2X1 g65798(.A (n_14313), .B (n_18627), .Y (n_19582));
OAI21X1 g65804(.A0 (n_17048), .A1 (n_9264), .B0 (n_12113), .Y(n_19581));
NAND2X1 g65852(.A (n_17667), .B (n_11927), .Y (n_19580));
OAI22X1 g65874(.A0 (n_8089), .A1 (n_4188), .B0 (n_3471), .B1(n_27290), .Y (n_19579));
OAI22X1 g65882(.A0 (n_7700), .A1 (n_4521), .B0 (n_3102), .B1(n_18716), .Y (n_19578));
OR4X1 g61350(.A (n_14505), .B (n_19576), .C (n_16582), .D (n_13702),.Y (n_19577));
NAND4X1 g61352(.A (n_17483), .B (n_11798), .C (n_10937), .D (n_6126),.Y (n_19575));
NAND4X1 g61355(.A (n_17481), .B (n_11820), .C (n_10915), .D (n_7876),.Y (n_19574));
NAND4X1 g61369(.A (n_16456), .B (n_14409), .C (n_13816), .D(n_13204), .Y (n_19573));
NAND4X1 g61376(.A (n_13397), .B (n_12556), .C (n_13811), .D(n_13197), .Y (n_19572));
NAND4X1 g61379(.A (n_16393), .B (n_14254), .C (n_13809), .D(n_13179), .Y (n_19571));
NAND4X1 g61381(.A (n_14798), .B (n_10892), .C (n_13806), .D(n_13205), .Y (n_19570));
NAND4X1 g61399(.A (n_17494), .B (n_19568), .C (n_6064), .D (n_16551),.Y (n_19569));
NAND4X1 g61401(.A (n_17493), .B (n_17841), .C (n_5941), .D (n_15675),.Y (n_19567));
NAND4X1 g61459(.A (n_12325), .B (n_19291), .C (n_13813), .D (n_3677),.Y (n_19566));
NAND3X1 g61463(.A (n_12328), .B (n_15797), .C (n_19299), .Y(n_19565));
NOR2X1 g66486(.A (n_17888), .B (n_27688), .Y (n_19564));
OAI21X1 g61525(.A0 (n_15573), .A1 (n_14529), .B0 (n_1196), .Y(n_28854));
OAI21X1 g61536(.A0 (n_15633), .A1 (n_13188), .B0 (sa32[1] ), .Y(n_19561));
AOI21X1 g61542(.A0 (n_16141), .A1 (n_15730), .B0 (n_5329), .Y(n_19559));
INVX1 g66695(.A (n_18728), .Y (n_20617));
AOI21X1 g61548(.A0 (n_15982), .A1 (n_15729), .B0 (n_15574), .Y(n_19558));
INVX1 g66761(.A (n_18724), .Y (n_19557));
AOI21X1 g61572(.A0 (n_14320), .A1 (n_15768), .B0 (n_29065), .Y(n_19556));
AOI21X1 g61574(.A0 (n_14132), .A1 (n_15717), .B0 (n_14589), .Y(n_19555));
NAND2X1 g61588(.A (n_17521), .B (n_4582), .Y (n_19554));
OAI21X1 g61589(.A0 (n_15750), .A1 (n_16423), .B0 (sa12[1] ), .Y(n_19553));
NAND3X1 g61603(.A (n_25820), .B (n_8683), .C (n_25821), .Y (n_19552));
NAND2X1 g61608(.A (n_17454), .B (n_20585), .Y (n_19551));
NAND3X1 g61613(.A (n_14894), .B (n_12859), .C (n_15711), .Y(n_19550));
NOR3X1 g61621(.A (n_6435), .B (n_10172), .C (n_15578), .Y (n_19549));
NAND4X1 g61630(.A (n_12256), .B (n_12807), .C (n_13535), .D (n_9399),.Y (n_19548));
AOI21X1 g61633(.A0 (n_15704), .A1 (n_12885), .B0 (n_12298), .Y(n_19547));
NAND3X1 g61642(.A (n_5779), .B (n_15492), .C (n_17685), .Y (n_19545));
NAND4X1 g61644(.A (n_11362), .B (n_17531), .C (n_12203), .D(n_13515), .Y (n_19544));
NAND3X1 g61647(.A (n_17438), .B (n_19542), .C (n_13071), .Y(n_19543));
NAND3X1 g61648(.A (n_17496), .B (n_11094), .C (n_18895), .Y(n_19541));
OAI21X1 g61649(.A0 (n_15745), .A1 (n_10154), .B0 (n_20558), .Y(n_19540));
AND2X1 g61651(.A (n_17533), .B (n_16806), .Y (n_19539));
NAND2X1 g61659(.A (n_17451), .B (n_903), .Y (n_19538));
NAND4X1 g61660(.A (n_18982), .B (n_28815), .C (n_13561), .D(n_13489), .Y (n_19536));
NAND3X1 g61669(.A (n_17586), .B (n_11716), .C (n_15775), .Y(n_19535));
NAND3X1 g61670(.A (n_19799), .B (n_15589), .C (n_8990), .Y (n_19534));
NAND2X1 g61671(.A (n_17450), .B (n_19532), .Y (n_19533));
NAND4X1 g61673(.A (n_10894), .B (n_28450), .C (n_13367), .D(n_14694), .Y (n_19531));
NAND4X1 g61676(.A (n_25763), .B (n_19529), .C (n_12234), .D (n_9143),.Y (n_19530));
NAND4X1 g61677(.A (n_12846), .B (n_17024), .C (n_13756), .D(n_14862), .Y (n_19528));
AOI21X1 g61678(.A0 (n_15553), .A1 (n_20144), .B0 (n_28988), .Y(n_25585));
NAND3X1 g61679(.A (n_12716), .B (n_7874), .C (n_15726), .Y (n_19526));
AND2X1 g61687(.A (n_15845), .B (n_17837), .Y (n_19525));
NAND2X1 g61690(.A (n_17449), .B (n_1991), .Y (n_19524));
NAND4X1 g61691(.A (n_11517), .B (n_9365), .C (n_9303), .D (n_14918),.Y (n_19522));
NAND3X1 g61696(.A (n_17498), .B (n_13703), .C (n_16956), .Y(n_19521));
NAND2X1 g61700(.A (n_17435), .B (n_869), .Y (n_19520));
NAND4X1 g61703(.A (n_17018), .B (n_12772), .C (n_13739), .D(n_14773), .Y (n_19518));
AOI21X1 g61705(.A0 (n_15585), .A1 (n_196), .B0 (n_9286), .Y(n_19517));
NAND3X1 g61706(.A (n_14079), .B (n_16482), .C (n_13812), .Y(n_19516));
AOI21X1 g61717(.A0 (n_15584), .A1 (n_15674), .B0 (n_13156), .Y(n_19515));
NAND3X1 g61722(.A (n_16050), .B (n_7232), .C (n_15725), .Y (n_19511));
AOI21X1 g61726(.A0 (n_15542), .A1 (n_10438), .B0 (n_28631), .Y(n_19510));
AOI21X1 g61727(.A0 (n_15524), .A1 (n_10467), .B0 (n_638), .Y(n_19508));
NOR3X1 g61731(.A (n_5177), .B (n_8439), .C (n_15571), .Y (n_28593));
OAI21X1 g61736(.A0 (n_11491), .A1 (n_15582), .B0 (sa10[1] ), .Y(n_28553));
NAND4X1 g61737(.A (n_10465), .B (n_17508), .C (n_12251), .D(n_13410), .Y (n_19504));
NAND3X1 g61738(.A (n_17431), .B (n_19502), .C (n_12993), .Y(n_19503));
NAND4X1 g61744(.A (n_18264), .B (n_19499), .C (n_15350), .D(n_13395), .Y (n_19500));
NAND4X1 g61747(.A (n_19008), .B (n_16236), .C (n_16599), .D(n_13379), .Y (n_19498));
NAND3X1 g61751(.A (n_14299), .B (n_8370), .C (n_15724), .Y (n_19497));
NAND3X1 g61752(.A (n_28837), .B (n_9952), .C (n_28838), .Y (n_19496));
AOI21X1 g61754(.A0 (n_15541), .A1 (n_13910), .B0 (n_3886), .Y(n_19495));
AOI21X1 g61763(.A0 (n_15537), .A1 (n_129), .B0 (n_18614), .Y(n_25641));
NAND3X1 g61764(.A (n_12497), .B (n_8344), .C (n_15723), .Y (n_19492));
NAND4X1 g61765(.A (n_17455), .B (n_15825), .C (n_14044), .D(n_15038), .Y (n_19491));
NAND3X1 g61766(.A (n_17430), .B (n_26673), .C (n_16208), .Y(n_19490));
AOI21X1 g61775(.A0 (n_15536), .A1 (n_19486), .B0 (n_16670), .Y(n_19487));
NAND3X1 g61777(.A (n_12463), .B (n_7259), .C (n_15722), .Y (n_19485));
AOI21X1 g61779(.A0 (n_16668), .A1 (n_15491), .B0 (n_1008), .Y(n_19484));
NAND3X1 g61780(.A (n_15977), .B (n_15721), .C (n_15770), .Y(n_19482));
NAND3X1 g61795(.A (n_14177), .B (n_16382), .C (n_15754), .Y(n_19481));
AOI21X1 g61797(.A0 (n_15530), .A1 (n_9146), .B0 (n_29039), .Y(n_19480));
AOI21X1 g61805(.A0 (n_15529), .A1 (n_12061), .B0 (n_3910), .Y(n_19479));
NAND3X1 g61810(.A (n_28260), .B (n_7616), .C (n_11112), .Y (n_19477));
AOI21X1 g61811(.A0 (n_15523), .A1 (n_19475), .B0 (n_13025), .Y(n_19476));
AOI21X1 g61816(.A0 (n_15527), .A1 (n_10493), .B0 (n_1295), .Y(n_19474));
NAND2X1 g61821(.A (n_17447), .B (n_804), .Y (n_19473));
NAND3X1 g61823(.A (n_14292), .B (n_14114), .C (n_15598), .Y(n_19472));
NAND4X1 g61826(.A (n_25628), .B (n_18707), .C (n_27708), .D (n_6207),.Y (n_19471));
AOI21X1 g61827(.A0 (n_15522), .A1 (n_7305), .B0 (n_19651), .Y(n_19470));
AOI21X1 g61829(.A0 (n_16530), .A1 (n_15486), .B0 (n_1196), .Y(n_19469));
NOR3X1 g61830(.A (n_6440), .B (n_9745), .C (n_15563), .Y (n_29384));
OAI21X1 g61835(.A0 (n_15751), .A1 (n_9763), .B0 (n_20587), .Y(n_19467));
NAND4X1 g61838(.A (n_28507), .B (n_15642), .C (n_9108), .D (n_7076),.Y (n_19466));
NAND4X1 g61840(.A (n_17156), .B (n_14245), .C (n_17824), .D(n_10074), .Y (n_19465));
NAND4X1 g61847(.A (n_15434), .B (n_9040), .C (n_14925), .D (n_13528),.Y (n_19464));
AOI22X1 g61857(.A0 (n_15599), .A1 (n_16466), .B0 (n_6135), .B1(n_583), .Y (n_19463));
NAND4X1 g61865(.A (n_16722), .B (n_13477), .C (n_12706), .D(n_13605), .Y (n_19462));
AOI22X1 g61869(.A0 (n_15660), .A1 (n_4582), .B0 (n_3287), .B1(n_1626), .Y (n_19461));
NAND4X1 g61871(.A (n_25507), .B (n_18691), .C (n_17356), .D (n_8867),.Y (n_19460));
NAND4X1 g61880(.A (n_14923), .B (n_13438), .C (n_12925), .D(n_13581), .Y (n_19459));
AOI21X1 g61883(.A0 (n_15481), .A1 (n_14909), .B0 (n_191), .Y(n_19458));
NAND3X1 g61890(.A (n_12541), .B (n_15773), .C (n_14991), .Y(n_19457));
INVX1 g61891(.A (n_18708), .Y (n_19456));
NAND4X1 g61896(.A (n_13590), .B (n_8784), .C (n_15059), .D (n_15061),.Y (n_19455));
NAND4X1 g61899(.A (n_25823), .B (n_16621), .C (n_26913), .D (n_9200),.Y (n_19454));
AOI21X1 g61904(.A0 (n_15479), .A1 (n_15034), .B0 (n_129), .Y(n_19453));
NAND2X1 g61905(.A (n_17507), .B (sa11[1] ), .Y (n_19452));
AOI21X1 g61910(.A0 (n_15478), .A1 (n_19450), .B0 (n_21275), .Y(n_19451));
OAI21X1 g61912(.A0 (n_15475), .A1 (n_7718), .B0 (n_875), .Y(n_19448));
AOI22X1 g61933(.A0 (n_15558), .A1 (n_4357), .B0 (n_4358), .B1(n_14757), .Y (n_19447));
AOI22X1 g61935(.A0 (n_15485), .A1 (n_19445), .B0 (n_9235), .B1(n_13083), .Y (n_19446));
NAND3X1 g61945(.A (n_13281), .B (n_15604), .C (n_11182), .Y(n_19444));
NAND3X1 g61949(.A (n_13345), .B (n_15623), .C (n_11092), .Y(n_19443));
NAND3X1 g61953(.A (n_14993), .B (n_15614), .C (n_9539), .Y (n_19442));
AOI22X1 g61957(.A0 (n_15484), .A1 (n_27407), .B0 (n_10869), .B1(n_19395), .Y (n_19441));
NAND4X1 g61969(.A (n_15257), .B (n_15313), .C (n_11584), .D(n_14611), .Y (n_19439));
AOI21X1 g61971(.A0 (n_15629), .A1 (n_15574), .B0 (n_13665), .Y(n_19438));
AOI21X1 g61980(.A0 (n_15552), .A1 (n_3264), .B0 (n_12662), .Y(n_19436));
AOI22X1 g61991(.A0 (n_15641), .A1 (n_19433), .B0 (n_14534), .B1(n_20406), .Y (n_19434));
NAND4X1 g61994(.A (n_16587), .B (n_16574), .C (n_13626), .D(n_14691), .Y (n_19432));
NAND4X1 g62005(.A (n_12738), .B (n_14325), .C (n_19430), .D(n_13671), .Y (n_19431));
NAND3X1 g62007(.A (n_9310), .B (n_15519), .C (n_19428), .Y (n_19429));
NAND4X1 g62014(.A (n_14385), .B (n_14257), .C (n_19130), .D(n_13667), .Y (n_19427));
NAND4X1 g62019(.A (n_12365), .B (n_12691), .C (n_19423), .D(n_13661), .Y (n_19424));
NAND4X1 g62022(.A (n_14097), .B (n_14506), .C (n_18251), .D(n_13659), .Y (n_19422));
NAND4X1 g62023(.A (n_15917), .B (n_12735), .C (n_19420), .D(n_13660), .Y (n_19421));
NAND4X1 g62025(.A (n_14498), .B (n_14433), .C (n_19417), .D(n_13674), .Y (n_19418));
AOI21X1 g62032(.A0 (n_16106), .A1 (n_13608), .B0 (n_20116), .Y(n_19416));
NAND2X1 g62036(.A (n_16947), .B (n_19414), .Y (n_19415));
AOI21X1 g62042(.A0 (n_16125), .A1 (n_14730), .B0 (sa12[1] ), .Y(n_19413));
NAND2X1 g62046(.A (n_17086), .B (n_196), .Y (n_19411));
OAI21X1 g62049(.A0 (n_15318), .A1 (n_10640), .B0 (n_16835), .Y(n_19410));
OAI21X1 g62051(.A0 (n_15307), .A1 (n_7895), .B0 (n_19408), .Y(n_28581));
OAI21X1 g62053(.A0 (n_15298), .A1 (n_12098), .B0 (n_15894), .Y(n_19407));
OAI21X1 g62055(.A0 (n_15179), .A1 (n_14528), .B0 (n_19791), .Y(n_19406));
AOI21X1 g62058(.A0 (n_15242), .A1 (n_16291), .B0 (w3[9] ), .Y(n_19405));
OAI21X1 g62060(.A0 (n_11523), .A1 (n_16293), .B0 (n_27216), .Y(n_19404));
AOI21X1 g62062(.A0 (n_16575), .A1 (n_11414), .B0 (n_15482), .Y(n_19402));
INVX1 g62065(.A (n_18685), .Y (n_19401));
AOI21X1 g62067(.A0 (n_4951), .A1 (n_3668), .B0 (n_16945), .Y(n_19400));
OAI21X1 g62069(.A0 (n_15168), .A1 (n_11988), .B0 (n_19398), .Y(n_28320));
OAI21X1 g62072(.A0 (n_15129), .A1 (n_10448), .B0 (n_19364), .Y(n_19397));
OAI21X1 g62076(.A0 (n_16718), .A1 (n_8912), .B0 (n_19395), .Y(n_25617));
OAI21X1 g62077(.A0 (n_16716), .A1 (n_16289), .B0 (n_21275), .Y(n_19394));
OAI21X1 g62081(.A0 (n_15015), .A1 (n_16288), .B0 (n_19834), .Y(n_19393));
OAI21X1 g62082(.A0 (n_16666), .A1 (n_16287), .B0 (n_20102), .Y(n_19392));
OAI21X1 g62083(.A0 (n_14998), .A1 (n_16286), .B0 (n_26903), .Y(n_19391));
OAI21X1 g62084(.A0 (n_14989), .A1 (n_16292), .B0 (n_28172), .Y(n_19389));
OAI21X1 g62085(.A0 (n_16646), .A1 (n_16285), .B0 (n_21396), .Y(n_19388));
OAI21X1 g62087(.A0 (n_16603), .A1 (n_10370), .B0 (n_19385), .Y(n_19386));
OAI21X1 g62091(.A0 (n_15172), .A1 (n_10264), .B0 (n_17411), .Y(n_19384));
OAI21X1 g62095(.A0 (n_16319), .A1 (n_15347), .B0 (n_171), .Y(n_19383));
OAI21X1 g62099(.A0 (n_16465), .A1 (n_11296), .B0 (n_21055), .Y(n_19381));
OAI21X1 g62103(.A0 (n_16318), .A1 (n_16567), .B0 (n_129), .Y(n_19379));
OAI21X1 g62106(.A0 (n_16315), .A1 (n_15107), .B0 (n_27242), .Y(n_19377));
OAI21X1 g62108(.A0 (n_13378), .A1 (n_16314), .B0 (n_2681), .Y(n_19376));
AOI21X1 g62112(.A0 (n_16397), .A1 (n_12993), .B0 (sa30[1] ), .Y(n_19375));
OAI21X1 g62118(.A0 (n_16417), .A1 (n_16316), .B0 (n_21275), .Y(n_19374));
OAI21X1 g62119(.A0 (n_16333), .A1 (n_14764), .B0 (n_19372), .Y(n_19373));
NAND2X1 g62120(.A (n_17095), .B (n_15371), .Y (n_19371));
NAND2X1 g62121(.A (n_17085), .B (n_129), .Y (n_19370));
OAI21X1 g62123(.A0 (n_16433), .A1 (n_11076), .B0 (n_19791), .Y(n_19369));
NAND2X1 g62125(.A (n_17061), .B (n_28172), .Y (n_19368));
NAND2X1 g62127(.A (n_17059), .B (n_1397), .Y (n_19367));
OAI21X1 g62132(.A0 (n_16361), .A1 (n_12599), .B0 (n_19364), .Y(n_19365));
OAI21X1 g62133(.A0 (n_16357), .A1 (n_5006), .B0 (n_18266), .Y(n_19363));
AOI21X1 g62142(.A0 (n_15311), .A1 (n_19361), .B0 (n_16074), .Y(n_19362));
NAND2X1 g62143(.A (n_16946), .B (n_20153), .Y (n_19360));
AOI21X1 g62144(.A0 (n_15157), .A1 (n_9580), .B0 (n_124), .Y(n_19358));
NOR2X1 g62150(.A (n_16993), .B (n_19355), .Y (n_19356));
NAND2X1 g62151(.A (n_16942), .B (n_869), .Y (n_19354));
AOI21X1 g62152(.A0 (n_15136), .A1 (n_14589), .B0 (n_12605), .Y(n_19353));
AOI21X1 g62156(.A0 (n_15065), .A1 (n_28645), .B0 (n_10949), .Y(n_19352));
NOR2X1 g62158(.A (n_11596), .B (n_17184), .Y (n_19351));
NOR2X1 g62159(.A (n_11594), .B (n_17181), .Y (n_19350));
NOR2X1 g62160(.A (n_13622), .B (n_17178), .Y (n_19349));
NOR2X1 g62161(.A (n_13618), .B (n_17263), .Y (n_19348));
INVX1 g62164(.A (n_18666), .Y (n_19347));
NAND2X1 g62169(.A (n_17313), .B (n_27604), .Y (n_28255));
XOR2X1 g68827(.A (n_1386), .B (n_15458), .Y (n_19345));
AOI21X1 g62174(.A0 (n_15235), .A1 (n_12626), .B0 (n_19310), .Y(n_19344));
NAND2X1 g62180(.A (n_17233), .B (n_28645), .Y (n_19342));
OAI21X1 g62184(.A0 (n_15160), .A1 (n_10288), .B0 (n_15039), .Y(n_19341));
NAND2X1 g62186(.A (n_17210), .B (n_15039), .Y (n_19340));
NAND2X1 g62188(.A (n_17294), .B (n_14589), .Y (n_19339));
OAI21X1 g62196(.A0 (n_12257), .A1 (n_869), .B0 (n_16984), .Y(n_19334));
OAI21X1 g62199(.A0 (n_10770), .A1 (n_20153), .B0 (n_16980), .Y(n_19333));
INVX1 g62200(.A (n_18655), .Y (n_19332));
NAND2X1 g62208(.A (n_17344), .B (n_19048), .Y (n_19331));
INVX1 g62209(.A (n_18647), .Y (n_19330));
NAND3X1 g62214(.A (n_14565), .B (n_16284), .C (n_17228), .Y(n_19329));
AOI21X1 g62225(.A0 (n_15286), .A1 (n_12827), .B0 (n_16572), .Y(n_19328));
AOI21X1 g62226(.A0 (n_16638), .A1 (n_12896), .B0 (n_15284), .Y(n_19327));
NAND2X1 g62227(.A (n_17320), .B (n_20406), .Y (n_19325));
OAI21X1 g62237(.A0 (n_15252), .A1 (n_19321), .B0 (n_21055), .Y(n_19322));
NAND2X1 g62240(.A (n_16962), .B (n_19319), .Y (n_19320));
NAND3X1 g62244(.A (n_15930), .B (n_16281), .C (n_19811), .Y(n_19318));
NAND3X1 g62249(.A (n_18393), .B (n_15426), .C (n_19314), .Y(n_19315));
NAND2X1 g62252(.A (n_11036), .B (n_17348), .Y (n_19313));
NAND2X1 g62257(.A (n_17290), .B (n_828), .Y (n_19312));
NAND2X1 g62262(.A (n_16955), .B (n_19310), .Y (n_19311));
NOR2X1 g62268(.A (n_17186), .B (n_15175), .Y (n_19309));
OAI21X1 g62269(.A0 (n_15206), .A1 (n_13921), .B0 (n_14474), .Y(n_19308));
NAND2X1 g62270(.A (n_17030), .B (n_503), .Y (n_19307));
OAI21X1 g62272(.A0 (n_15237), .A1 (n_16462), .B0 (n_2981), .Y(n_25677));
OAI21X1 g62273(.A0 (n_15200), .A1 (n_14081), .B0 (n_27100), .Y(n_19304));
NAND3X1 g62281(.A (n_18385), .B (n_13598), .C (n_21290), .Y(n_19302));
NOR2X1 g62282(.A (n_17272), .B (n_16781), .Y (n_19301));
AND2X1 g62283(.A (n_16979), .B (n_19299), .Y (n_19300));
NAND4X1 g62284(.A (n_25502), .B (n_8121), .C (n_14448), .D (n_19297),.Y (n_19298));
NOR2X1 g62285(.A (n_17270), .B (n_15465), .Y (n_19296));
OR2X1 g62287(.A (n_17063), .B (n_869), .Y (n_19295));
AOI21X1 g62290(.A0 (n_13332), .A1 (n_15712), .B0 (n_17869), .Y(n_19294));
NAND2X1 g62291(.A (n_16969), .B (n_17689), .Y (n_19293));
AND2X1 g62292(.A (n_16977), .B (n_19291), .Y (n_19292));
AOI21X1 g62293(.A0 (n_16544), .A1 (n_14474), .B0 (n_13942), .Y(n_19290));
OAI21X1 g62294(.A0 (n_15219), .A1 (n_19287), .B0 (n_21275), .Y(n_19288));
OAI21X1 g62296(.A0 (n_15320), .A1 (n_8857), .B0 (n_17912), .Y(n_19286));
OAI21X1 g62301(.A0 (n_15139), .A1 (n_13926), .B0 (n_20325), .Y(n_19285));
OAI21X1 g62302(.A0 (n_15138), .A1 (n_16428), .B0 (n_485), .Y(n_19284));
NAND2X1 g62314(.A (n_17230), .B (n_27336), .Y (n_19282));
NAND4X1 g62320(.A (n_19218), .B (n_15681), .C (n_14658), .D(n_12971), .Y (n_19281));
AOI21X1 g62324(.A0 (n_15077), .A1 (n_16358), .B0 (n_16740), .Y(n_19280));
AND2X1 g62329(.A (n_17220), .B (n_14668), .Y (n_19279));
OAI21X1 g62333(.A0 (n_16712), .A1 (n_16401), .B0 (n_27128), .Y(n_25627));
AOI21X1 g62337(.A0 (n_13350), .A1 (n_19276), .B0 (n_20055), .Y(n_22708));
NAND2X1 g62339(.A (n_17209), .B (n_18456), .Y (n_19275));
OAI21X1 g62341(.A0 (n_16685), .A1 (n_11940), .B0 (n_18266), .Y(n_19274));
OAI21X1 g62342(.A0 (n_14239), .A1 (n_16392), .B0 (n_3886), .Y(n_19273));
NAND3X1 g62344(.A (n_17650), .B (n_14809), .C (n_6986), .Y (n_19272));
OAI21X1 g62349(.A0 (n_16664), .A1 (n_14806), .B0 (n_2001), .Y(n_19271));
NAND2X1 g62353(.A (n_17131), .B (n_29102), .Y (n_19270));
OAI21X1 g62355(.A0 (n_16656), .A1 (n_14992), .B0 (n_875), .Y(n_25496));
OAI21X1 g62358(.A0 (n_15078), .A1 (n_13927), .B0 (n_19364), .Y(n_19268));
NAND3X1 g62360(.A (n_15930), .B (n_16373), .C (n_7222), .Y (n_19267));
AOI21X1 g62361(.A0 (n_28878), .A1 (n_28879), .B0 (n_28172), .Y(n_19266));
AOI21X1 g62363(.A0 (n_14984), .A1 (n_16641), .B0 (n_27910), .Y(n_19264));
OAI21X1 g62364(.A0 (n_16633), .A1 (n_14127), .B0 (n_18456), .Y(n_19263));
NAND2X1 g62365(.A (n_16952), .B (n_624), .Y (n_19261));
OAI21X1 g62366(.A0 (n_16630), .A1 (n_13907), .B0 (n_28692), .Y(n_19260));
NAND2X1 g62368(.A (n_17038), .B (n_28631), .Y (n_19259));
NAND2X1 g62372(.A (n_16951), .B (n_2983), .Y (n_19258));
NAND2X1 g62382(.A (n_17227), .B (n_10900), .Y (n_19257));
NAND2X1 g62385(.A (n_12765), .B (n_17351), .Y (n_19256));
AOI21X1 g62386(.A0 (n_14965), .A1 (n_29062), .B0 (n_17921), .Y(n_19255));
AOI21X1 g62390(.A0 (n_13294), .A1 (n_17567), .B0 (n_17883), .Y(n_19253));
NAND2X1 g62392(.A (n_10853), .B (n_17350), .Y (n_19252));
NAND2X1 g62393(.A (n_16967), .B (n_18749), .Y (n_19251));
NAND2X1 g62397(.A (n_14135), .B (n_17397), .Y (n_19250));
NAND2X1 g62401(.A (n_16966), .B (n_17681), .Y (n_19249));
NAND3X1 g62403(.A (n_13301), .B (n_15923), .C (n_19247), .Y(n_19248));
NAND3X1 g62405(.A (n_12320), .B (n_16278), .C (n_17310), .Y(n_19246));
NOR3X1 g62407(.A (n_11900), .B (n_9710), .C (n_16298), .Y (n_19245));
NAND3X1 g62410(.A (n_17650), .B (n_13120), .C (n_19243), .Y(n_19244));
NAND3X1 g62412(.A (n_16882), .B (n_14777), .C (n_19033), .Y(n_19242));
AOI21X1 g62413(.A0 (n_16522), .A1 (n_17864), .B0 (n_17836), .Y(n_19241));
NAND2X1 g62414(.A (n_14905), .B (n_17112), .Y (n_19240));
NAND2X1 g62416(.A (n_14086), .B (n_17347), .Y (n_19237));
NOR2X1 g62417(.A (n_17152), .B (n_7245), .Y (n_19236));
AOI21X1 g62419(.A0 (n_16508), .A1 (n_9819), .B0 (n_15363), .Y(n_19234));
AOI21X1 g62423(.A0 (n_13082), .A1 (n_7410), .B0 (n_17084), .Y(n_19232));
NAND2X1 g62424(.A (n_16224), .B (n_17078), .Y (n_19231));
AOI22X1 g62426(.A0 (n_15204), .A1 (n_15166), .B0 (n_13211), .B1(n_5817), .Y (n_19230));
AOI22X1 g62437(.A0 (n_15247), .A1 (n_13083), .B0 (n_15588), .B1(n_5400), .Y (n_19228));
AOI22X1 g62438(.A0 (n_15212), .A1 (n_11603), .B0 (n_19226), .B1(n_3552), .Y (n_19227));
NAND4X1 g62452(.A (n_11056), .B (n_9214), .C (n_8544), .D (n_14875),.Y (n_19225));
NAND3X1 g62453(.A (n_17324), .B (n_15927), .C (n_15544), .Y(n_19224));
NOR2X1 g62454(.A (n_16476), .B (n_17316), .Y (n_19223));
NOR2X1 g62455(.A (n_16340), .B (n_17311), .Y (n_29306));
NOR2X1 g62459(.A (n_17802), .B (n_15683), .Y (n_19221));
NAND4X1 g62462(.A (n_18854), .B (n_16446), .C (n_19243), .D(n_12220), .Y (n_19220));
NAND4X1 g62465(.A (n_17757), .B (n_19218), .C (n_7168), .D (n_14843),.Y (n_19219));
NAND4X1 g62467(.A (n_13482), .B (n_19216), .C (n_13698), .D(n_14853), .Y (n_19217));
NOR2X1 g62469(.A (n_16415), .B (n_17237), .Y (n_25678));
NOR2X1 g62470(.A (n_16409), .B (n_17229), .Y (n_29407));
NAND3X1 g62472(.A (n_15635), .B (n_16004), .C (n_17033), .Y(n_19213));
OAI21X1 g62479(.A0 (n_16336), .A1 (n_9585), .B0 (n_3886), .Y(n_19212));
NAND3X1 g62487(.A (n_16834), .B (n_15292), .C (n_13521), .Y(n_19211));
AOI21X1 g62489(.A0 (n_16429), .A1 (n_19445), .B0 (n_16998), .Y(n_19210));
OAI21X1 g62490(.A0 (n_16484), .A1 (n_19207), .B0 (n_19651), .Y(n_19208));
AOI21X1 g62493(.A0 (n_7864), .A1 (n_19030), .B0 (n_17019), .Y(n_19205));
NAND3X1 g62498(.A (n_13430), .B (n_15419), .C (n_12466), .Y(n_19204));
INVX1 g62510(.A (n_18561), .Y (n_19203));
AOI22X1 g62521(.A0 (n_15208), .A1 (n_14155), .B0 (n_2701), .B1(n_11901), .Y (n_19202));
AOI21X1 g62523(.A0 (n_6216), .A1 (n_17288), .B0 (n_17025), .Y(n_19200));
AOI21X1 g62528(.A0 (n_5017), .A1 (n_7507), .B0 (n_17022), .Y(n_19199));
AOI21X1 g62533(.A0 (n_16470), .A1 (n_15176), .B0 (w3[17] ), .Y(n_19198));
OAI21X1 g62538(.A0 (n_15887), .A1 (n_26253), .B0 (n_20325), .Y(n_19196));
OAI21X1 g62539(.A0 (n_19182), .A1 (n_14201), .B0 (n_29048), .Y(n_19195));
NAND3X1 g62540(.A (n_25861), .B (n_16283), .C (n_13016), .Y(n_19194));
OAI21X1 g62541(.A0 (n_16427), .A1 (n_19191), .B0 (n_1310), .Y(n_19192));
AOI21X1 g62543(.A0 (n_15123), .A1 (n_975), .B0 (n_4706), .Y(n_19190));
AOI22X1 g62550(.A0 (n_15080), .A1 (n_29062), .B0 (n_5936), .B1(n_15997), .Y (n_19189));
OAI21X1 g62557(.A0 (n_16709), .A1 (n_29018), .B0 (n_7393), .Y(n_19188));
OAI21X1 g62558(.A0 (n_16399), .A1 (n_19186), .B0 (n_28689), .Y(n_19187));
INVX1 g62559(.A (n_18553), .Y (n_19184));
OAI21X1 g62567(.A0 (n_16381), .A1 (n_25860), .B0 (n_29048), .Y(n_19181));
OAI21X1 g62569(.A0 (n_16377), .A1 (n_13835), .B0 (n_19364), .Y(n_25589));
OAI21X1 g62572(.A0 (n_16369), .A1 (n_11882), .B0 (n_28692), .Y(n_25810));
NAND2X1 g62573(.A (n_8275), .B (n_17390), .Y (n_19177));
AOI21X1 g62593(.A0 (n_16608), .A1 (n_1830), .B0 (n_4605), .Y(n_19175));
OAI21X1 g62606(.A0 (n_16407), .A1 (n_12970), .B0 (n_1295), .Y(n_19174));
NAND2X1 g62610(.A (n_17357), .B (n_27336), .Y (n_19173));
NOR2X1 g62618(.A (n_7272), .B (n_17047), .Y (n_19172));
NAND3X1 g62622(.A (n_13447), .B (n_15153), .C (n_15879), .Y(n_19169));
NAND3X1 g62625(.A (n_14980), .B (n_13313), .C (n_15873), .Y(n_19168));
NOR2X1 g62629(.A (n_13299), .B (n_17187), .Y (n_19167));
NOR2X1 g62630(.A (n_17867), .B (n_13721), .Y (n_19166));
NAND3X1 g62632(.A (n_17097), .B (n_15705), .C (n_19951), .Y(n_19165));
OAI21X1 g62633(.A0 (n_15343), .A1 (n_7260), .B0 (n_18876), .Y(n_19164));
OAI21X1 g62635(.A0 (n_15268), .A1 (n_6888), .B0 (n_18094), .Y(n_19162));
OAI21X1 g62637(.A0 (n_16453), .A1 (n_12278), .B0 (n_19160), .Y(n_19161));
OAI21X1 g62638(.A0 (n_16450), .A1 (n_9759), .B0 (n_9326), .Y(n_19159));
NAND2X1 g62643(.A (n_17218), .B (n_19157), .Y (n_19158));
OAI21X1 g62645(.A0 (n_16386), .A1 (n_12815), .B0 (n_28054), .Y(n_19156));
OAI21X1 g62646(.A0 (n_16380), .A1 (n_5913), .B0 (n_9272), .Y(n_19154));
NAND2X1 g62647(.A (n_17198), .B (n_19152), .Y (n_19153));
NAND4X1 g62650(.A (n_25522), .B (n_25523), .C (n_18958), .D (n_9720),.Y (n_19151));
OAI21X1 g62657(.A0 (n_16518), .A1 (n_7823), .B0 (n_18102), .Y(n_19150));
NAND4X1 g62658(.A (n_8757), .B (n_13690), .C (n_6528), .D (n_14723),.Y (n_19149));
NOR2X1 g62660(.A (n_16843), .B (n_17404), .Y (n_19148));
AOI22X1 g62662(.A0 (n_16565), .A1 (n_16480), .B0 (n_15497), .B1(n_16934), .Y (n_19147));
AOI22X1 g62670(.A0 (n_16330), .A1 (n_15482), .B0 (n_11039), .B1(n_2702), .Y (n_19145));
AOI21X1 g62674(.A0 (n_16320), .A1 (n_19143), .B0 (n_13293), .Y(n_19144));
NOR2X1 g62680(.A (n_15297), .B (n_17400), .Y (n_19142));
NAND4X1 g62700(.A (n_15640), .B (n_18114), .C (n_7219), .D (n_14749),.Y (n_19138));
NAND4X1 g62701(.A (n_17302), .B (n_15245), .C (n_6983), .D (n_14751),.Y (n_19137));
NAND3X1 g62702(.A (n_15046), .B (n_16306), .C (n_26040), .Y(n_19136));
NAND4X1 g62703(.A (n_16501), .B (n_17619), .C (n_7228), .D (n_14748),.Y (n_19134));
NAND3X1 g62706(.A (n_15013), .B (n_16304), .C (n_18697), .Y(n_19133));
NOR2X1 g62707(.A (n_13323), .B (n_17128), .Y (n_19132));
NAND3X1 g62708(.A (n_13321), .B (n_16302), .C (n_19130), .Y(n_19131));
NAND3X1 g62709(.A (n_17899), .B (n_14746), .C (n_26912), .Y(n_19129));
NOR2X1 g62712(.A (n_17575), .B (n_16987), .Y (n_19127));
NOR2X1 g62713(.A (n_17573), .B (n_15512), .Y (n_19126));
NAND4X1 g62716(.A (n_12239), .B (n_15954), .C (n_18248), .D(n_18249), .Y (n_19125));
NAND2X1 g62718(.A (n_10131), .B (n_17110), .Y (n_28242));
OAI21X1 g62722(.A0 (n_16309), .A1 (n_15039), .B0 (n_6957), .Y(n_19123));
NAND2X1 g62726(.A (n_9074), .B (n_17100), .Y (n_19121));
AOI22X1 g62734(.A0 (n_16296), .A1 (n_16466), .B0 (n_4634), .B1(n_7410), .Y (n_19118));
AOI22X1 g62752(.A0 (n_16490), .A1 (n_16978), .B0 (n_9755), .B1(n_5417), .Y (n_19116));
AOI22X1 g62755(.A0 (n_16479), .A1 (n_20010), .B0 (n_19114), .B1(n_16290), .Y (n_19115));
AOI21X1 g62757(.A0 (n_15246), .A1 (n_19445), .B0 (n_12327), .Y(n_19113));
AOI22X1 g62758(.A0 (n_16461), .A1 (n_19111), .B0 (n_19110), .B1(n_11412), .Y (n_19112));
AOI21X1 g62763(.A0 (n_15146), .A1 (n_15655), .B0 (n_12671), .Y(n_19109));
AND2X1 g62765(.A (n_11178), .B (n_17268), .Y (n_19108));
NAND4X1 g62766(.A (n_11409), .B (n_18342), .C (n_7206), .D (n_12751),.Y (n_19107));
NOR2X1 g62767(.A (n_10907), .B (n_17164), .Y (n_19106));
NOR2X1 g62771(.A (n_10978), .B (n_17231), .Y (n_19105));
NAND2X1 g62776(.A (n_16053), .B (n_17146), .Y (n_19104));
AOI21X1 g62777(.A0 (n_16430), .A1 (n_3886), .B0 (n_13060), .Y(n_19103));
NOR2X1 g62780(.A (n_7711), .B (n_17137), .Y (n_19102));
AOI21X1 g62783(.A0 (n_16388), .A1 (n_28689), .B0 (n_12941), .Y(n_19101));
AOI21X1 g62784(.A0 (n_16294), .A1 (n_17912), .B0 (n_11120), .Y(n_19100));
NAND4X1 g62797(.A (n_19097), .B (n_7065), .C (n_25736), .D (n_10098),.Y (n_19098));
NAND4X1 g62798(.A (n_19095), .B (n_6732), .C (n_25639), .D (n_9937),.Y (n_19096));
OAI21X1 g62806(.A0 (n_14501), .A1 (n_16154), .B0 (n_16835), .Y(n_19094));
OAI21X1 g62808(.A0 (n_14551), .A1 (n_16129), .B0 (n_27604), .Y(n_19092));
OAI21X1 g62818(.A0 (n_14470), .A1 (n_16094), .B0 (n_15574), .Y(n_19090));
OAI21X1 g62820(.A0 (n_15976), .A1 (n_18400), .B0 (n_11261), .Y(n_29321));
OR2X1 g62836(.A (n_17743), .B (n_26931), .Y (n_25592));
AOI21X1 g62837(.A0 (n_15970), .A1 (n_18245), .B0 (n_21442), .Y(n_19086));
INVX1 g62839(.A (n_18488), .Y (n_19085));
OR2X1 g62841(.A (n_17736), .B (n_28169), .Y (n_19084));
AOI21X1 g62861(.A0 (n_11773), .A1 (n_17979), .B0 (n_21055), .Y(n_19083));
NAND2X1 g62862(.A (n_17919), .B (n_17571), .Y (n_19082));
AND2X1 g62864(.A (n_16761), .B (n_27604), .Y (n_19081));
AOI21X1 g62869(.A0 (n_16257), .A1 (n_14222), .B0 (n_15776), .Y(n_19079));
OR2X1 g62873(.A (n_17804), .B (n_11261), .Y (n_19078));
NAND2X1 g62877(.A (n_17803), .B (n_14624), .Y (n_19075));
AOI21X1 g62880(.A0 (n_16250), .A1 (n_19071), .B0 (n_16835), .Y(n_19072));
AND2X1 g62881(.A (n_17783), .B (n_15574), .Y (n_19070));
AND2X1 g62883(.A (n_17758), .B (n_18320), .Y (n_19068));
AOI21X1 g62897(.A0 (n_16246), .A1 (n_13376), .B0 (n_29102), .Y(n_19065));
NAND2X1 g62901(.A (n_17739), .B (n_29102), .Y (n_19062));
AOI21X1 g62906(.A0 (n_9792), .A1 (n_19060), .B0 (n_19372), .Y(n_29401));
AOI21X1 g62909(.A0 (n_9767), .A1 (n_18811), .B0 (n_21275), .Y(n_19059));
AOI21X1 g62917(.A0 (n_16041), .A1 (n_14978), .B0 (n_14474), .Y(n_19058));
AOI21X1 g62919(.A0 (n_16131), .A1 (n_17821), .B0 (n_12298), .Y(n_19057));
AOI21X1 g62925(.A0 (n_16083), .A1 (n_14942), .B0 (n_16835), .Y(n_19055));
NAND2X1 g62952(.A (n_16313), .B (n_19052), .Y (n_19053));
AOI21X1 g62980(.A0 (n_16039), .A1 (n_5329), .B0 (n_9918), .Y(n_19051));
NAND2X1 g62988(.A (n_17697), .B (n_11486), .Y (n_19050));
NAND2X1 g62989(.A (n_17695), .B (n_19048), .Y (n_19049));
NAND2X1 g63008(.A (n_14752), .B (n_19046), .Y (n_19047));
NAND3X1 g63010(.A (n_6354), .B (n_16186), .C (n_5226), .Y (n_19045));
NAND3X1 g63013(.A (n_25614), .B (n_7927), .C (n_7939), .Y (n_19044));
NAND3X1 g63018(.A (n_6392), .B (n_16162), .C (n_4516), .Y (n_19043));
INVX1 g63029(.A (n_18417), .Y (n_19042));
INVX1 g63034(.A (n_18414), .Y (n_19041));
OAI21X1 g63040(.A0 (n_16081), .A1 (n_9370), .B0 (n_27746), .Y(n_19040));
NAND2X1 g63053(.A (n_17782), .B (n_16553), .Y (n_19039));
OAI21X1 g63055(.A0 (n_15882), .A1 (n_16163), .B0 (n_18205), .Y(n_19038));
OAI21X1 g63056(.A0 (n_15881), .A1 (n_16184), .B0 (n_17411), .Y(n_19037));
NAND2X1 g72539(.A (n_16924), .B (n_5114), .Y (n_19036));
NAND2X1 g63074(.A (n_16911), .B (n_14560), .Y (n_19035));
OAI21X1 g63087(.A0 (n_16124), .A1 (n_17405), .B0 (n_9371), .Y(n_19032));
OAI21X1 g63099(.A0 (n_16168), .A1 (n_19030), .B0 (n_14878), .Y(n_19031));
NAND2X1 g63127(.A (n_16802), .B (n_19445), .Y (n_19028));
OAI21X1 g63131(.A0 (n_15880), .A1 (n_11718), .B0 (n_27688), .Y(n_19027));
INVX1 g63138(.A (n_18384), .Y (n_19026));
OAI21X1 g63143(.A0 (n_15943), .A1 (n_10760), .B0 (n_638), .Y(n_19025));
NAND2X1 g63149(.A (n_17825), .B (n_27344), .Y (n_19024));
NAND3X1 g63150(.A (n_18286), .B (n_18826), .C (n_17897), .Y(n_19023));
OAI21X1 g63164(.A0 (n_16188), .A1 (n_19021), .B0 (n_1008), .Y(n_19022));
AOI21X1 g63166(.A0 (n_15908), .A1 (n_19019), .B0 (n_13466), .Y(n_19020));
OAI21X1 g63184(.A0 (n_15871), .A1 (n_27152), .B0 (n_16835), .Y(n_19018));
AOI21X1 g63193(.A0 (n_12660), .A1 (n_15883), .B0 (n_12986), .Y(n_19016));
AND2X1 g63194(.A (n_17812), .B (n_29262), .Y (n_19015));
NAND2X1 g63215(.A (n_16813), .B (n_1991), .Y (n_25457));
OAI21X1 g63222(.A0 (n_15940), .A1 (n_17412), .B0 (n_1497), .Y(n_19013));
OR2X1 g63226(.A (n_17818), .B (n_11261), .Y (n_19012));
NAND3X1 g63235(.A (n_17293), .B (n_17292), .C (n_17590), .Y(n_19011));
NAND2X1 g63241(.A (n_17898), .B (n_16007), .Y (n_19010));
NAND2X1 g63254(.A (n_17960), .B (n_19008), .Y (n_19009));
NAND2X1 g63263(.A (n_17771), .B (n_14367), .Y (n_19007));
NAND2X1 g63272(.A (n_16751), .B (n_908), .Y (n_19006));
INVX1 g63292(.A (n_18329), .Y (n_19004));
OR2X1 g63303(.A (n_17938), .B (n_20332), .Y (n_19003));
NAND2X1 g63309(.A (n_17817), .B (n_1295), .Y (n_19002));
NAND2X1 g63314(.A (n_17931), .B (n_18074), .Y (n_19001));
NAND2X1 g63319(.A (n_18978), .B (n_11945), .Y (n_19000));
INVX1 g63322(.A (n_18321), .Y (n_18999));
NAND3X1 g63324(.A (n_10417), .B (n_14372), .C (n_10328), .Y(n_18998));
NAND3X1 g63333(.A (n_18330), .B (n_14247), .C (n_18996), .Y(n_18997));
OR2X1 g63347(.A (n_17816), .B (n_14155), .Y (n_18995));
INVX1 g63355(.A (n_18307), .Y (n_18994));
INVX1 g63365(.A (n_18304), .Y (n_18993));
AOI21X1 g63367(.A0 (n_15884), .A1 (n_12435), .B0 (n_19364), .Y(n_18992));
OR2X1 g63374(.A (n_17815), .B (n_29102), .Y (n_18991));
AOI21X1 g63382(.A0 (n_15892), .A1 (n_12688), .B0 (n_28692), .Y(n_18988));
OR2X1 g63405(.A (n_16925), .B (n_14589), .Y (n_18986));
NAND2X1 g63412(.A (n_17995), .B (n_18982), .Y (n_18983));
OAI21X1 g63414(.A0 (n_17645), .A1 (n_4853), .B0 (n_16434), .Y(n_28586));
NAND2X1 g63418(.A (n_17772), .B (n_15074), .Y (n_18980));
NOR2X1 g63421(.A (n_18978), .B (n_21569), .Y (n_18979));
NOR2X1 g63429(.A (n_17718), .B (n_14561), .Y (n_28323));
NAND2X1 g63436(.A (n_16749), .B (n_903), .Y (n_18975));
NAND2X1 g63437(.A (n_17716), .B (n_13423), .Y (n_18974));
NAND2X1 g63445(.A (n_18817), .B (n_28245), .Y (n_18973));
OAI21X1 g63454(.A0 (n_17653), .A1 (n_29404), .B0 (n_18440), .Y(n_18972));
NAND3X1 g63458(.A (n_13684), .B (n_16161), .C (n_5856), .Y (n_18971));
NAND2X1 g63466(.A (n_17708), .B (n_13575), .Y (n_18970));
INVX1 g63473(.A (n_18265), .Y (n_18969));
NAND4X1 g63507(.A (n_18967), .B (n_18966), .C (n_10609), .D(n_18965), .Y (n_18968));
NOR2X1 g63508(.A (n_17785), .B (n_13476), .Y (n_18964));
NOR2X1 g63512(.A (n_6892), .B (n_16917), .Y (n_18963));
NOR2X1 g63518(.A (n_16739), .B (n_14310), .Y (n_25596));
INVX1 g63520(.A (n_18250), .Y (n_18961));
INVX1 g63525(.A (n_18246), .Y (n_18960));
NAND4X1 g63533(.A (n_17416), .B (n_18958), .C (n_18882), .D(n_13741), .Y (n_18959));
NOR2X1 g63537(.A (n_7119), .B (n_16918), .Y (n_18957));
INVX1 g63545(.A (n_18238), .Y (n_18955));
INVX1 g63567(.A (n_18235), .Y (n_18954));
OAI21X1 g63575(.A0 (n_17655), .A1 (n_15590), .B0 (n_15894), .Y(n_18953));
NAND2X1 g63587(.A (n_16860), .B (n_25895), .Y (n_18952));
NAND2X1 g63590(.A (n_16856), .B (n_15894), .Y (n_18951));
NAND3X1 g63598(.A (n_13852), .B (n_15896), .C (n_18948), .Y(n_18949));
NAND3X1 g63601(.A (n_6287), .B (n_15895), .C (n_18946), .Y (n_18947));
AOI21X1 g63605(.A0 (n_15868), .A1 (n_3886), .B0 (n_15289), .Y(n_18945));
NAND2X1 g63608(.A (n_16826), .B (n_17703), .Y (n_18943));
NAND3X1 g63614(.A (n_8390), .B (n_15893), .C (n_18941), .Y (n_18942));
OAI21X1 g63616(.A0 (n_18018), .A1 (n_583), .B0 (n_12192), .Y(n_18940));
AND2X1 g63619(.A (n_16816), .B (n_18937), .Y (n_18938));
NAND2X1 g63629(.A (n_16798), .B (n_18153), .Y (n_18936));
OAI21X1 g63637(.A0 (n_17624), .A1 (n_751), .B0 (n_10720), .Y(n_18934));
NAND2X1 g63640(.A (n_16852), .B (n_26872), .Y (n_18933));
NAND2X1 g63644(.A (n_16784), .B (n_12713), .Y (n_18932));
NAND2X1 g63650(.A (n_16851), .B (n_12740), .Y (n_18931));
NAND2X1 g63658(.A (n_13446), .B (n_18914), .Y (n_18930));
NAND2X1 g63662(.A (n_16786), .B (n_12198), .Y (n_18929));
OAI21X1 g63664(.A0 (n_16146), .A1 (n_18266), .B0 (n_16868), .Y(n_18928));
NAND3X1 g63680(.A (n_11791), .B (n_15890), .C (n_18926), .Y(n_18927));
NAND2X1 g63681(.A (n_16769), .B (n_28692), .Y (n_18925));
AND2X1 g63687(.A (n_16756), .B (n_18922), .Y (n_18923));
OR2X1 g63689(.A (n_16805), .B (n_18920), .Y (n_18921));
NAND2X1 g63709(.A (n_16733), .B (n_5329), .Y (n_18918));
AOI21X1 g63718(.A0 (n_15866), .A1 (n_28689), .B0 (n_17923), .Y(n_18916));
NAND4X1 g63731(.A (n_18914), .B (n_5659), .C (n_11889), .D (n_7524),.Y (n_18915));
AOI21X1 g63732(.A0 (n_16113), .A1 (n_3122), .B0 (n_9999), .Y(n_18913));
OAI21X1 g63735(.A0 (n_18911), .A1 (n_28645), .B0 (n_27266), .Y(n_18912));
NOR2X1 g63737(.A (n_17914), .B (n_15428), .Y (n_18910));
NAND2X1 g63753(.A (n_17596), .B (n_16874), .Y (n_18908));
NAND3X1 g63757(.A (n_17731), .B (n_14635), .C (n_13771), .Y(n_18907));
NAND3X1 g63758(.A (n_17729), .B (n_17969), .C (n_11732), .Y(n_18906));
OAI21X1 g63761(.A0 (n_18904), .A1 (n_28689), .B0 (n_27238), .Y(n_18905));
AOI21X1 g63766(.A0 (n_9175), .A1 (n_624), .B0 (n_17877), .Y(n_18903));
NAND2X1 g63771(.A (n_17872), .B (n_14155), .Y (n_18902));
NAND2X1 g63784(.A (n_16774), .B (n_17459), .Y (n_18901));
NAND2X1 g63785(.A (n_13879), .B (n_16873), .Y (n_18900));
NAND2X1 g63792(.A (n_17852), .B (n_17773), .Y (n_18899));
NAND2X1 g63799(.A (n_17840), .B (n_12506), .Y (n_18898));
AOI21X1 g63808(.A0 (n_18765), .A1 (n_18895), .B0 (n_18100), .Y(n_18896));
OR2X1 g63814(.A (n_13624), .B (n_16884), .Y (n_18893));
NAND4X1 g63819(.A (n_17665), .B (n_6986), .C (n_13960), .D (n_8166),.Y (n_18891));
NAND2X1 g63823(.A (n_16757), .B (n_18889), .Y (n_18890));
AOI21X1 g63837(.A0 (n_12158), .A1 (n_5151), .B0 (n_16833), .Y(n_18888));
INVX1 g63844(.A (n_18111), .Y (n_18887));
AOI21X1 g63846(.A0 (n_10694), .A1 (n_15473), .B0 (n_16791), .Y(n_18886));
NAND3X1 g63858(.A (n_14587), .B (n_25626), .C (n_12648), .Y(n_18884));
NAND3X1 g63860(.A (n_14391), .B (n_16639), .C (n_18882), .Y(n_18883));
NOR2X1 g63861(.A (n_12056), .B (n_16858), .Y (n_18881));
NOR2X1 g63881(.A (n_12612), .B (n_18016), .Y (n_18880));
AND2X1 g63882(.A (n_16796), .B (n_15233), .Y (n_18879));
NAND2X1 g63898(.A (n_17111), .B (n_19752), .Y (n_18878));
AND2X1 g63901(.A (n_17928), .B (n_16706), .Y (n_18875));
AND2X1 g63904(.A (n_17918), .B (n_15008), .Y (n_25735));
NAND3X1 g63979(.A (n_7590), .B (n_16146), .C (n_27496), .Y (n_18873));
NAND3X1 g63995(.A (n_17910), .B (n_7795), .C (n_15272), .Y (n_18871));
NAND2X1 g64024(.A (n_14852), .B (n_16919), .Y (n_18870));
NAND2X1 g64025(.A (n_17713), .B (n_15441), .Y (n_18869));
NAND2X1 g64026(.A (n_17720), .B (n_15440), .Y (n_18868));
NAND2X1 g64029(.A (n_16871), .B (n_16780), .Y (n_18867));
AND2X1 g64031(.A (n_28885), .B (n_28886), .Y (n_18866));
NAND2X1 g64032(.A (n_17863), .B (n_17862), .Y (n_18865));
XOR2X1 g76256(.A (text_in_r[19] ), .B (n_18792), .Y (n_18864));
INVX1 g64149(.A (n_18021), .Y (n_21210));
INVX1 g64163(.A (n_19643), .Y (n_18861));
NOR2X1 g64171(.A (n_18859), .B (n_16835), .Y (n_18860));
NAND2X1 g64234(.A (n_17548), .B (n_28169), .Y (n_18856));
NAND2X1 g64287(.A (n_18854), .B (n_18859), .Y (n_18855));
INVX1 g64363(.A (n_18852), .Y (n_18853));
INVX1 g64479(.A (n_18849), .Y (n_18850));
NAND2X1 g64566(.A (n_17557), .B (n_15894), .Y (n_18848));
OR2X1 g64614(.A (n_17556), .B (n_16835), .Y (n_18847));
NAND2X1 g64663(.A (n_13171), .B (n_18859), .Y (n_18846));
NAND2X1 g64865(.A (n_27022), .B (n_17411), .Y (n_18845));
NAND2X1 g64866(.A (n_16024), .B (n_16663), .Y (n_18844));
NOR2X1 g64889(.A (n_14161), .B (n_13431), .Y (n_18843));
OR2X1 g64892(.A (n_15996), .B (n_12896), .Y (n_18842));
NAND2X1 g64895(.A (n_14673), .B (n_14405), .Y (n_18841));
INVX1 g64901(.A (n_18978), .Y (n_18840));
AOI21X1 g64928(.A0 (n_13759), .A1 (n_8092), .B0 (n_2470), .Y(n_18839));
AND2X1 g64953(.A (n_18085), .B (n_16253), .Y (n_18838));
NOR2X1 g64965(.A (n_11256), .B (n_16262), .Y (n_18836));
INVX1 g64980(.A (n_17911), .Y (n_18835));
OR2X1 g64995(.A (n_16048), .B (n_19395), .Y (n_18834));
NOR2X1 g65000(.A (n_6994), .B (n_13095), .Y (n_18833));
AND2X1 g65001(.A (n_14961), .B (n_15914), .Y (n_28276));
NOR2X1 g65005(.A (n_14647), .B (n_13023), .Y (n_18831));
NOR2X1 g65019(.A (n_16197), .B (n_11260), .Y (n_25590));
NAND2X1 g65091(.A (n_15861), .B (n_2909), .Y (n_18829));
NAND2X1 g65094(.A (n_18827), .B (n_18826), .Y (n_18828));
NAND2X1 g65098(.A (n_13256), .B (n_18826), .Y (n_18825));
NAND2X1 g65105(.A (n_16018), .B (n_16758), .Y (n_18823));
INVX1 g65112(.A (n_17886), .Y (n_18822));
NAND2X1 g65124(.A (n_17660), .B (n_11921), .Y (n_18821));
NAND2X1 g65138(.A (n_15859), .B (n_20862), .Y (n_18820));
NAND2X1 g65148(.A (n_10105), .B (n_19060), .Y (n_18819));
INVX1 g65157(.A (n_18817), .Y (n_18818));
NAND2X1 g65176(.A (n_17672), .B (n_15352), .Y (n_18816));
NAND2X1 g65180(.A (n_15967), .B (n_18785), .Y (n_18815));
NAND2X1 g65202(.A (n_15914), .B (n_12416), .Y (n_18814));
NAND2X1 g65215(.A (n_13743), .B (n_18811), .Y (n_18812));
NAND2X1 g65224(.A (n_18809), .B (n_8648), .Y (n_18810));
NAND2X1 g65244(.A (n_18807), .B (n_9785), .Y (n_18808));
AOI21X1 g65299(.A0 (n_13864), .A1 (n_9552), .B0 (n_17411), .Y(n_18806));
INVX1 g65315(.A (n_17828), .Y (n_18804));
NAND3X1 g65327(.A (n_28877), .B (n_12059), .C (n_12779), .Y(n_18803));
NAND2X1 g65332(.A (n_15875), .B (n_18801), .Y (n_18802));
NAND3X1 g65344(.A (n_28809), .B (n_12057), .C (n_20628), .Y(n_18800));
NAND3X1 g65353(.A (n_16639), .B (n_10354), .C (n_10384), .Y(n_18799));
INVX1 g65445(.A (n_17809), .Y (n_18797));
NOR2X1 g65495(.A (n_14421), .B (n_14437), .Y (n_18796));
NAND2X1 g65500(.A (n_9032), .B (n_14673), .Y (n_18795));
AOI21X1 g65504(.A0 (n_9322), .A1 (n_751), .B0 (n_14076), .Y(n_18794));
AOI21X1 g65512(.A0 (n_11854), .A1 (n_18792), .B0 (n_10724), .Y(n_18793));
NOR2X1 g65532(.A (n_16071), .B (n_12183), .Y (n_18790));
AND2X1 g65536(.A (n_16064), .B (n_15226), .Y (n_18789));
AND2X1 g65551(.A (n_16143), .B (n_9048), .Y (n_18788));
OAI21X1 g65559(.A0 (n_16492), .A1 (n_18785), .B0 (n_14014), .Y(n_18786));
NOR2X1 g65564(.A (n_11848), .B (n_16237), .Y (n_18784));
INVX1 g65579(.A (n_17774), .Y (n_18783));
NAND4X1 g61227(.A (n_12848), .B (n_10851), .C (n_7672), .D (n_11690),.Y (n_18782));
NAND2X1 g65608(.A (n_16019), .B (n_7645), .Y (n_18781));
NAND2X1 g65616(.A (n_15936), .B (n_18598), .Y (n_18780));
OAI21X1 g65673(.A0 (n_16394), .A1 (n_6185), .B0 (n_28161), .Y(n_18779));
AND2X1 g65692(.A (n_14219), .B (n_18241), .Y (n_18778));
AOI21X1 g65710(.A0 (n_13735), .A1 (n_4938), .B0 (n_21396), .Y(n_18777));
NAND2X1 g65715(.A (n_15963), .B (n_9371), .Y (n_18776));
NAND2X1 g65717(.A (n_16195), .B (n_16359), .Y (n_18774));
OAI21X1 g65719(.A0 (n_29202), .A1 (n_28373), .B0 (n_14362), .Y(n_18773));
NOR2X1 g65728(.A (n_11729), .B (n_16259), .Y (n_18772));
AOI21X1 g65737(.A0 (n_13899), .A1 (n_8022), .B0 (n_19364), .Y(n_18771));
NOR2X1 g65767(.A (n_14145), .B (n_13882), .Y (n_18768));
INVX1 g65783(.A (n_17712), .Y (n_18767));
NAND2X1 g65832(.A (n_10696), .B (n_18765), .Y (n_18766));
NAND2X1 g65839(.A (n_16268), .B (n_10180), .Y (n_18764));
NAND2X1 g65846(.A (n_16249), .B (n_10008), .Y (n_18763));
NAND2X1 g65850(.A (n_16221), .B (n_10026), .Y (n_18762));
NAND2X1 g65853(.A (n_9843), .B (n_16200), .Y (n_18761));
NOR2X1 g65856(.A (n_15979), .B (n_11010), .Y (n_18760));
OAI21X1 g65870(.A0 (n_2617), .A1 (n_13885), .B0 (n_9701), .Y(n_18759));
NAND2X1 g65892(.A (n_12336), .B (n_18007), .Y (n_18758));
NAND2X1 g65897(.A (n_12569), .B (n_18756), .Y (n_29386));
AOI21X1 g65903(.A0 (n_10429), .A1 (n_2112), .B0 (n_15956), .Y(n_18755));
AOI21X1 g65904(.A0 (n_10531), .A1 (n_16006), .B0 (n_15987), .Y(n_18754));
AOI21X1 g65905(.A0 (n_10618), .A1 (n_10147), .B0 (n_16101), .Y(n_18753));
AOI21X1 g65910(.A0 (n_10556), .A1 (n_14107), .B0 (n_15901), .Y(n_18752));
NAND2X1 g65921(.A (n_16016), .B (n_12305), .Y (n_18751));
NAND4X1 g65924(.A (n_8062), .B (n_18749), .C (n_9127), .D (n_17717),.Y (n_18750));
NAND2X1 g65928(.A (n_16055), .B (n_8573), .Y (n_18748));
NAND2X1 g65937(.A (n_16027), .B (n_8277), .Y (n_18747));
NAND2X1 g65954(.A (n_11985), .B (n_16240), .Y (n_18746));
INVX1 g65986(.A (n_17676), .Y (n_18745));
NAND2X1 g66025(.A (n_27152), .B (n_18266), .Y (n_18744));
INVX1 g66054(.A (n_17675), .Y (n_18741));
NAND4X1 g61400(.A (n_15819), .B (n_18739), .C (n_4593), .D (n_15414),.Y (n_18740));
NAND2X1 g66405(.A (n_19364), .B (n_16005), .Y (n_18738));
NAND2X1 g61511(.A (n_15794), .B (n_12788), .Y (n_18734));
NOR2X1 g66573(.A (n_15068), .B (n_28692), .Y (n_18732));
NAND2X1 g66581(.A (n_16835), .B (n_13912), .Y (n_18731));
INVX1 g66678(.A (n_17659), .Y (n_18729));
NOR2X1 g66696(.A (n_13801), .B (n_13593), .Y (n_18728));
NOR2X1 g66730(.A (n_27077), .B (n_12986), .Y (n_28274));
OR2X1 g61562(.A (n_15834), .B (n_15039), .Y (n_18725));
NOR2X1 g66762(.A (n_15764), .B (n_16434), .Y (n_18724));
NAND2X1 g61596(.A (n_15826), .B (n_15986), .Y (n_18723));
OAI21X1 g61612(.A0 (n_13777), .A1 (n_18721), .B0 (n_503), .Y(n_18722));
NAND2X1 g61623(.A (n_15802), .B (n_20577), .Y (n_18719));
NOR2X1 g67009(.A (n_15708), .B (n_18716), .Y (n_18718));
NAND2X1 g61643(.A (n_15795), .B (n_1699), .Y (n_18715));
OR2X1 g67220(.A (n_13744), .B (n_27604), .Y (n_18714));
NAND4X1 g61740(.A (n_10983), .B (n_17425), .C (n_11485), .D (n_9431),.Y (n_18713));
NAND2X1 g67441(.A (n_18682), .B (n_4276), .Y (n_18712));
NOR2X1 g67599(.A (n_15574), .B (n_27290), .Y (n_18711));
NAND3X1 g61790(.A (n_14191), .B (n_14795), .C (n_13802), .Y(n_18709));
NAND3X1 g61892(.A (n_11478), .B (n_13733), .C (n_18707), .Y(n_18708));
OR4X1 g61903(.A (n_26362), .B (n_12342), .C (n_10711), .D (n_13325),.Y (n_18706));
NAND2X1 g61907(.A (n_15829), .B (sa12[1] ), .Y (n_18704));
NAND2X1 g68276(.A (n_14761), .B (n_20325), .Y (n_18703));
AOI21X1 g61979(.A0 (n_13713), .A1 (n_933), .B0 (n_12838), .Y(n_18702));
AOI21X1 g61981(.A0 (n_13711), .A1 (n_124), .B0 (n_12378), .Y(n_18700));
NAND4X1 g61992(.A (n_18116), .B (n_16941), .C (n_17140), .D(n_11621), .Y (n_18699));
NAND4X1 g62006(.A (n_12805), .B (n_14358), .C (n_18697), .D(n_11614), .Y (n_18698));
AOI21X1 g62010(.A0 (n_19226), .A1 (n_7567), .B0 (n_15838), .Y(n_18696));
NAND4X1 g62012(.A (n_28887), .B (n_14513), .C (n_17115), .D(n_28888), .Y (n_18695));
NAND4X1 g62015(.A (n_8246), .B (n_14268), .C (n_17127), .D (n_11612),.Y (n_18694));
NAND4X1 g62020(.A (n_9782), .B (n_18691), .C (n_17134), .D (n_11628),.Y (n_18692));
NOR2X1 g68479(.A (n_5538), .B (n_15813), .Y (n_18690));
AOI21X1 g62034(.A0 (n_14427), .A1 (n_14729), .B0 (n_20412), .Y(n_18689));
NOR2X1 g68528(.A (n_7015), .B (n_15801), .Y (n_18688));
AOI21X1 g62043(.A0 (n_12459), .A1 (n_14731), .B0 (sa10[1] ), .Y(n_18687));
AOI21X1 g62064(.A0 (n_5128), .A1 (n_5064), .B0 (n_15483), .Y(n_18686));
AOI21X1 g62066(.A0 (n_11513), .A1 (n_14735), .B0 (n_20577), .Y(n_18685));
AOI21X1 g62068(.A0 (n_14904), .A1 (n_12655), .B0 (n_20406), .Y(n_18684));
NAND2X1 g68597(.A (n_10630), .B (n_18682), .Y (n_18683));
OAI21X1 g62089(.A0 (n_14938), .A1 (n_10414), .B0 (n_9106), .Y(n_18681));
OAI21X1 g62092(.A0 (n_13517), .A1 (n_10537), .B0 (n_18679), .Y(n_18680));
OAI21X1 g62093(.A0 (n_13503), .A1 (n_10277), .B0 (n_17567), .Y(n_18678));
OAI21X1 g62094(.A0 (n_13405), .A1 (n_10410), .B0 (n_14807), .Y(n_18676));
OAI21X1 g62098(.A0 (n_13132), .A1 (n_13493), .B0 (n_4357), .Y(n_18675));
AOI21X1 g62124(.A0 (n_13492), .A1 (n_6862), .B0 (sa33[1] ), .Y(n_18674));
AOI21X1 g62126(.A0 (n_13369), .A1 (n_18310), .B0 (n_3538), .Y(n_18673));
OAI21X1 g62128(.A0 (n_14828), .A1 (n_10815), .B0 (n_15776), .Y(n_18672));
OAI21X1 g68764(.A0 (n_3281), .A1 (n_9654), .B0 (n_15764), .Y(n_18671));
NAND3X1 g62148(.A (n_14692), .B (n_4540), .C (n_17295), .Y (n_18670));
XOR2X1 g68816(.A (n_1073), .B (n_13654), .Y (n_18669));
NAND2X1 g62163(.A (n_15715), .B (n_11277), .Y (n_18668));
AOI21X1 g62165(.A0 (n_13544), .A1 (n_12632), .B0 (n_1132), .Y(n_18666));
NAND2X1 g62166(.A (n_15698), .B (n_9410), .Y (n_18665));
OAI21X1 g62172(.A0 (n_13433), .A1 (n_10522), .B0 (n_11300), .Y(n_18664));
XOR2X1 g68830(.A (n_1006), .B (n_13670), .Y (n_18663));
OAI21X1 g62175(.A0 (n_14944), .A1 (n_10480), .B0 (n_16835), .Y(n_18662));
XOR2X1 g68836(.A (n_1217), .B (n_13675), .Y (n_18661));
NAND2X1 g62178(.A (n_15647), .B (n_15568), .Y (n_18660));
OAI21X1 g62182(.A0 (n_13375), .A1 (n_10585), .B0 (n_19364), .Y(n_18659));
OAI21X1 g62187(.A0 (n_15016), .A1 (n_10397), .B0 (n_28692), .Y(n_18658));
INVX1 g62197(.A (n_17537), .Y (n_18656));
AOI21X1 g62201(.A0 (n_14789), .A1 (w3[17] ), .B0 (n_10771), .Y(n_18655));
OAI21X1 g62202(.A0 (n_14049), .A1 (n_20632), .B0 (n_15506), .Y(n_18654));
INVX1 g62203(.A (n_17535), .Y (n_18653));
OAI21X1 g62205(.A0 (n_14019), .A1 (n_20577), .B0 (n_15502), .Y(n_18652));
NAND4X1 g62206(.A (n_8293), .B (n_6830), .C (n_12761), .D (n_7274),.Y (n_18651));
NAND3X1 g62207(.A (n_18648), .B (n_9479), .C (n_13388), .Y (n_18649));
NAND3X1 g62210(.A (n_16151), .B (n_13117), .C (n_19814), .Y(n_18647));
AOI21X1 g62217(.A0 (n_14883), .A1 (n_10801), .B0 (n_18643), .Y(n_18644));
AOI21X1 g62222(.A0 (n_13534), .A1 (n_15507), .B0 (n_18641), .Y(n_18642));
AOI21X1 g62223(.A0 (n_13396), .A1 (n_12335), .B0 (n_28988), .Y(n_18640));
NAND2X1 g62228(.A (n_15498), .B (n_18635), .Y (n_18636));
AND2X1 g62229(.A (n_15508), .B (n_18633), .Y (n_18634));
NAND2X1 g62232(.A (n_15557), .B (n_20986), .Y (n_18632));
OAI21X1 g62236(.A0 (n_13499), .A1 (n_18630), .B0 (n_933), .Y(n_18631));
NAND2X1 g62239(.A (n_27715), .B (n_3724), .Y (n_28557));
AOI21X1 g62256(.A0 (n_13467), .A1 (n_16976), .B0 (n_11023), .Y(n_18626));
OAI21X1 g62259(.A0 (n_13568), .A1 (n_13462), .B0 (n_20587), .Y(n_18624));
OAI21X1 g62263(.A0 (n_13457), .A1 (n_13483), .B0 (n_15482), .Y(n_18622));
OAI21X1 g62275(.A0 (n_11521), .A1 (n_13442), .B0 (w3[25] ), .Y(n_18621));
NAND3X1 g62277(.A (n_18619), .B (n_11315), .C (n_13441), .Y(n_18620));
AOI21X1 g62278(.A0 (n_14782), .A1 (n_28901), .B0 (n_18617), .Y(n_18618));
NOR3X1 g62297(.A (n_28816), .B (n_9705), .C (n_14744), .Y (n_18616));
AOI21X1 g62298(.A0 (n_13573), .A1 (n_12568), .B0 (n_18614), .Y(n_18615));
AOI21X1 g62300(.A0 (n_13417), .A1 (n_15142), .B0 (n_29048), .Y(n_18613));
NAND4X1 g62312(.A (n_18050), .B (n_18051), .C (n_15067), .D(n_14981), .Y (n_18611));
NAND4X1 g62316(.A (n_9227), .B (n_17292), .C (n_15090), .D (n_15091),.Y (n_18610));
OAI21X1 g62317(.A0 (n_13389), .A1 (n_11469), .B0 (sa33[1] ), .Y(n_25780));
OAI21X1 g62322(.A0 (n_14929), .A1 (n_15274), .B0 (n_27336), .Y(n_25578));
OAI21X1 g62330(.A0 (n_15057), .A1 (n_28998), .B0 (n_17411), .Y(n_18605));
OAI21X1 g62331(.A0 (n_15056), .A1 (n_14822), .B0 (n_3910), .Y(n_18604));
OAI21X1 g62338(.A0 (n_15026), .A1 (n_18602), .B0 (n_20677), .Y(n_18603));
OAI21X1 g62340(.A0 (n_15020), .A1 (n_15018), .B0 (sa30[1] ), .Y(n_18601));
NAND3X1 g62350(.A (n_18598), .B (n_14802), .C (n_16713), .Y(n_18599));
OAI21X1 g62352(.A0 (n_14999), .A1 (n_14225), .B0 (n_3724), .Y(n_18597));
NAND2X1 g62359(.A (n_15535), .B (n_1310), .Y (n_18596));
NAND3X1 g62369(.A (n_16031), .B (n_13200), .C (n_6911), .Y (n_18594));
OR4X1 g62375(.A (n_7018), .B (n_9700), .C (n_5891), .D (n_12417), .Y(n_18593));
OAI21X1 g62377(.A0 (n_14976), .A1 (n_28609), .B0 (n_29070), .Y(n_18592));
AOI21X1 g62383(.A0 (n_13296), .A1 (n_26270), .B0 (n_16611), .Y(n_18591));
NAND4X1 g62391(.A (n_29143), .B (n_8112), .C (n_12382), .D (n_26469),.Y (n_18590));
NAND3X1 g62395(.A (n_18587), .B (n_12914), .C (n_14948), .Y(n_18588));
NOR3X1 g62396(.A (n_11795), .B (n_9713), .C (n_14740), .Y (n_18586));
NAND3X1 g62398(.A (n_16149), .B (n_13935), .C (n_7608), .Y (n_18585));
NAND3X1 g62400(.A (n_13118), .B (n_14098), .C (n_16647), .Y(n_18584));
NAND3X1 g62406(.A (n_18582), .B (n_14596), .C (n_14921), .Y(n_18583));
NAND3X1 g62411(.A (n_7347), .B (n_14908), .C (n_13267), .Y (n_18581));
DFFX1 u0_r0_out_reg[28] (.CK (clk), .D (n_15814), .Q (), .QN(u0_rcon_1057));
AOI22X1 g62427(.A0 (n_14943), .A1 (n_18266), .B0 (n_10357), .B1(n_9084), .Y (n_18580));
NAND2X1 g62435(.A (n_16542), .B (n_15490), .Y (n_18579));
NAND2X1 g62440(.A (n_14884), .B (n_15713), .Y (n_18578));
OAI21X1 g62442(.A0 (n_12843), .A1 (n_16787), .B0 (n_15709), .Y(n_18577));
NAND2X1 g62444(.A (n_14886), .B (n_15680), .Y (n_18576));
NAND2X1 g62445(.A (n_14791), .B (n_15669), .Y (n_18575));
OAI21X1 g62446(.A0 (n_12695), .A1 (n_12896), .B0 (n_15595), .Y(n_18574));
NAND2X1 g62447(.A (n_14837), .B (n_15650), .Y (n_18573));
NAND2X1 g62449(.A (n_29319), .B (n_29320), .Y (n_28239));
OAI21X1 g62450(.A0 (n_12527), .A1 (n_17414), .B0 (n_15637), .Y(n_18571));
NAND4X1 g62464(.A (n_10894), .B (n_15556), .C (n_7014), .D (n_13246),.Y (n_18570));
NAND3X1 g62482(.A (n_13546), .B (n_13547), .C (n_11029), .Y(n_18569));
AOI22X1 g62485(.A0 (n_13538), .A1 (n_14142), .B0 (n_3518), .B1(n_14878), .Y (n_18568));
AOI21X1 g62500(.A0 (n_13143), .A1 (n_16466), .B0 (n_16552), .Y(n_18567));
AOI21X1 g62504(.A0 (n_13203), .A1 (n_4582), .B0 (n_15174), .Y(n_18565));
OAI21X1 g62506(.A0 (n_13206), .A1 (n_27807), .B0 (n_11261), .Y(n_18563));
OAI21X1 g62511(.A0 (n_14787), .A1 (n_28220), .B0 (n_9410), .Y(n_18561));
NAND3X1 g62518(.A (n_11438), .B (n_13645), .C (n_17683), .Y(n_18559));
NAND3X1 g62531(.A (n_13436), .B (n_13437), .C (n_10909), .Y(n_18558));
OAI21X1 g62535(.A0 (n_13498), .A1 (n_11052), .B0 (n_5978), .Y(n_18557));
OAI21X1 g62551(.A0 (n_14824), .A1 (n_26048), .B0 (n_11277), .Y(n_18556));
XOR2X1 g60063(.A (u0_rcon_1054), .B (n_1227), .Y (n_18555));
NAND3X1 g62555(.A (n_15051), .B (n_15052), .C (n_10921), .Y(n_18554));
OAI21X1 g62560(.A0 (n_14814), .A1 (n_18552), .B0 (n_16754), .Y(n_18553));
NAND4X1 g62565(.A (n_14043), .B (n_14499), .C (n_12549), .D(n_16990), .Y (n_18551));
DFFX1 u0_r0_out_reg[26] (.CK (clk), .D (n_15686), .Q (u0_rcon_1055),.QN ());
DFFX1 u0_r0_out_reg[27] (.CK (clk), .D (n_15685), .Q (u0_rcon_1056),.QN ());
INVX1 g60074(.A (u0_rcon_1058), .Y (n_18549));
NAND3X1 g62594(.A (n_14960), .B (n_14963), .C (n_10957), .Y(n_18546));
OAI21X1 g62599(.A0 (n_14959), .A1 (n_7201), .B0 (n_5960), .Y(n_18545));
OR2X1 g70711(.A (n_15444), .B (n_13846), .Y (n_18544));
NOR2X1 g62624(.A (n_13566), .B (n_15601), .Y (n_18541));
NOR2X1 g62626(.A (n_11453), .B (n_15606), .Y (n_18540));
NOR2X1 g62627(.A (n_16623), .B (n_13726), .Y (n_18539));
OAI21X1 g62636(.A0 (n_14869), .A1 (n_196), .B0 (n_10749), .Y(n_18538));
NOR2X1 g62639(.A (n_14039), .B (n_15505), .Y (n_18536));
NAND2X1 g62642(.A (n_15649), .B (n_18087), .Y (n_18535));
OAI21X1 g62644(.A0 (n_14813), .A1 (n_10223), .B0 (n_12663), .Y(n_18534));
NOR2X1 g62648(.A (n_14020), .B (n_15501), .Y (n_18533));
AOI21X1 g62672(.A0 (n_6822), .A1 (n_6510), .B0 (n_15663), .Y(n_18530));
AOI22X1 g62678(.A0 (n_14771), .A1 (n_778), .B0 (n_14387), .B1(n_3168), .Y (n_18529));
NOR2X1 g62688(.A (n_16580), .B (n_15765), .Y (n_18524));
NAND4X1 g62704(.A (n_16503), .B (n_11338), .C (n_15837), .D(n_13128), .Y (n_18523));
NOR2X1 g62710(.A (n_15898), .B (n_15515), .Y (n_18522));
NAND4X1 g62715(.A (n_12216), .B (n_14192), .C (n_18243), .D(n_18244), .Y (n_18521));
OAI21X1 g62723(.A0 (n_14766), .A1 (n_10613), .B0 (n_18119), .Y(n_18520));
INVX1 g62749(.A (n_17439), .Y (n_18519));
NAND2X1 g62754(.A (n_16091), .B (n_15703), .Y (n_18518));
NOR2X1 g62761(.A (n_12677), .B (n_15676), .Y (n_18517));
NAND4X1 g62762(.A (n_13107), .B (n_17265), .C (n_17286), .D(n_12631), .Y (n_18516));
NAND2X1 g71387(.A (n_15450), .B (n_5114), .Y (n_18515));
AOI21X1 g62772(.A0 (n_14834), .A1 (n_28631), .B0 (n_9284), .Y(n_18514));
AOI21X1 g62786(.A0 (n_5760), .A1 (n_20010), .B0 (n_15579), .Y(n_18513));
NAND2X1 g62800(.A (n_15528), .B (n_10289), .Y (n_18512));
AOI21X1 g62805(.A0 (n_14846), .A1 (n_16944), .B0 (n_9938), .Y(n_18511));
OAI21X1 g62807(.A0 (n_14568), .A1 (n_11167), .B0 (n_15712), .Y(n_18510));
OAI21X1 g62809(.A0 (n_12582), .A1 (n_14221), .B0 (n_11300), .Y(n_18508));
NAND2X1 g62810(.A (n_16584), .B (n_15894), .Y (n_18506));
OAI21X1 g62814(.A0 (n_14479), .A1 (n_10807), .B0 (n_26670), .Y(n_18503));
NAND2X1 g62821(.A (n_15154), .B (n_20325), .Y (n_18502));
OAI21X1 g62822(.A0 (n_12630), .A1 (n_14443), .B0 (n_19364), .Y(n_18500));
OAI21X1 g62825(.A0 (n_14533), .A1 (n_14341), .B0 (n_18168), .Y(n_18497));
OAI21X1 g62826(.A0 (n_14331), .A1 (n_14170), .B0 (n_15039), .Y(n_18496));
OAI21X1 g62827(.A0 (n_14315), .A1 (n_10954), .B0 (n_28632), .Y(n_18494));
NAND2X1 g62828(.A (n_16728), .B (n_17411), .Y (n_29416));
AOI21X1 g62829(.A0 (n_14295), .A1 (n_16738), .B0 (n_19981), .Y(n_18491));
NAND2X1 g62840(.A (n_16653), .B (n_17912), .Y (n_18488));
OAI21X1 g62843(.A0 (n_14206), .A1 (n_9828), .B0 (n_17567), .Y(n_18487));
OAI21X1 g62847(.A0 (n_14198), .A1 (n_17253), .B0 (n_29062), .Y(n_25621));
OAI21X1 g62848(.A0 (n_14469), .A1 (n_9765), .B0 (n_15986), .Y(n_18485));
OAI21X1 g62851(.A0 (n_14180), .A1 (n_18278), .B0 (n_18320), .Y(n_18483));
OAI21X1 g62860(.A0 (n_14422), .A1 (n_9995), .B0 (n_14592), .Y(n_18481));
OR2X1 g62863(.A (n_16474), .B (n_18440), .Y (n_18480));
AOI21X1 g62870(.A0 (n_14520), .A1 (n_5327), .B0 (n_14878), .Y(n_18479));
OR2X1 g62872(.A (n_16473), .B (n_27099), .Y (n_18478));
AOI21X1 g62885(.A0 (n_9947), .A1 (n_16765), .B0 (n_14627), .Y(n_18475));
OR2X1 g62887(.A (n_16419), .B (n_16754), .Y (n_18474));
OR2X1 g62890(.A (n_16408), .B (n_11277), .Y (n_18473));
AND2X1 g62894(.A (n_16396), .B (n_19385), .Y (n_18472));
OR2X1 g62896(.A (n_16405), .B (n_19395), .Y (n_18470));
AOI21X1 g62898(.A0 (n_14640), .A1 (n_26731), .B0 (n_28645), .Y(n_18469));
AOI21X1 g62905(.A0 (n_10188), .A1 (n_18465), .B0 (n_1008), .Y(n_18466));
AOI21X1 g62911(.A0 (n_8142), .A1 (n_17844), .B0 (n_1196), .Y(n_18464));
AND2X1 g62912(.A (n_16517), .B (n_15776), .Y (n_18463));
OAI21X1 g62914(.A0 (n_14483), .A1 (n_28875), .B0 (n_828), .Y(n_18462));
AOI21X1 g62915(.A0 (n_14291), .A1 (n_11539), .B0 (n_18237), .Y(n_18460));
OAI21X1 g62918(.A0 (n_14329), .A1 (n_12427), .B0 (n_27336), .Y(n_18459));
OAI21X1 g62920(.A0 (n_14243), .A1 (n_28807), .B0 (n_18456), .Y(n_18457));
OAI21X1 g62922(.A0 (n_14214), .A1 (n_12553), .B0 (n_290), .Y(n_18455));
AOI21X1 g62923(.A0 (n_14187), .A1 (n_16683), .B0 (n_28645), .Y(n_18454));
NAND2X1 g62928(.A (n_15106), .B (n_18320), .Y (n_18453));
OAI21X1 g62929(.A0 (n_14338), .A1 (n_12178), .B0 (n_14807), .Y(n_18451));
NAND2X1 g62956(.A (n_16312), .B (n_13569), .Y (n_18450));
AND2X1 g62958(.A (n_16487), .B (n_15701), .Y (n_18449));
NAND2X1 g62967(.A (n_15255), .B (n_638), .Y (n_18447));
NAND2X1 g72208(.A (n_15477), .B (n_8520), .Y (n_18445));
NAND2X1 g62970(.A (n_16464), .B (n_17012), .Y (n_18443));
NOR2X1 g62971(.A (n_16437), .B (n_14605), .Y (n_18442));
AOI21X1 g62972(.A0 (n_14495), .A1 (n_18440), .B0 (n_8375), .Y(n_18441));
AOI21X1 g62973(.A0 (n_14429), .A1 (n_9410), .B0 (n_15072), .Y(n_18439));
NAND2X1 g62974(.A (n_14756), .B (n_18437), .Y (n_18438));
NOR2X1 g62979(.A (n_16424), .B (n_14680), .Y (n_18436));
NAND2X1 g62985(.A (n_15099), .B (n_510), .Y (n_18434));
NAND2X1 g62986(.A (n_16402), .B (n_17000), .Y (n_18433));
NAND2X1 g62987(.A (n_16308), .B (n_13506), .Y (n_18432));
AOI21X1 g62992(.A0 (n_14283), .A1 (n_12896), .B0 (n_8763), .Y(n_18431));
AOI21X1 g62993(.A0 (n_14148), .A1 (n_15568), .B0 (n_15355), .Y(n_18430));
NAND2X1 g62994(.A (n_15443), .B (n_14314), .Y (n_18429));
INVX1 g62998(.A (n_17365), .Y (n_28267));
NOR2X1 g63001(.A (n_16385), .B (n_9445), .Y (n_18425));
AOI21X1 g63002(.A0 (n_14276), .A1 (n_19857), .B0 (n_5906), .Y(n_18424));
AOI21X1 g63009(.A0 (n_17232), .A1 (n_26952), .B0 (n_28632), .Y(n_18423));
AND2X1 g63015(.A (n_16463), .B (n_18421), .Y (n_18422));
NAND2X1 g63019(.A (n_15439), .B (n_16652), .Y (n_18420));
OAI21X1 g63023(.A0 (n_14164), .A1 (n_11141), .B0 (n_17423), .Y(n_18419));
OAI21X1 g63025(.A0 (n_14167), .A1 (n_6202), .B0 (n_11253), .Y(n_18418));
AND2X1 g63030(.A (n_15183), .B (n_7410), .Y (n_18417));
INVX1 g63032(.A (n_17353), .Y (n_18415));
AND2X1 g63035(.A (n_15184), .B (n_5817), .Y (n_18414));
OAI21X1 g63037(.A0 (n_14406), .A1 (n_10950), .B0 (n_12019), .Y(n_18413));
OAI21X1 g63042(.A0 (n_14051), .A1 (n_7390), .B0 (n_29062), .Y(n_18412));
OAI21X1 g63049(.A0 (n_14511), .A1 (n_6197), .B0 (n_29286), .Y(n_18411));
NAND2X1 g63054(.A (n_13102), .B (n_18360), .Y (n_18410));
NAND3X1 g63058(.A (n_10523), .B (n_16704), .C (n_9592), .Y (n_18409));
NAND2X1 g63063(.A (n_15353), .B (n_16072), .Y (n_18408));
NOR2X1 g65390(.A (n_11876), .B (n_16272), .Y (n_18407));
NAND2X1 g63066(.A (n_15351), .B (n_20585), .Y (n_18406));
NAND3X1 g63070(.A (n_18335), .B (n_16912), .C (n_16857), .Y(n_18405));
INVX1 g63082(.A (n_17333), .Y (n_18404));
AND2X1 g63084(.A (n_15312), .B (n_11810), .Y (n_18403));
INVX1 g63085(.A (n_17332), .Y (n_18402));
OAI21X1 g63090(.A0 (n_14106), .A1 (n_18400), .B0 (n_1361), .Y(n_18401));
INVX1 g63091(.A (n_17330), .Y (n_18399));
NAND2X1 g63098(.A (n_15165), .B (n_16097), .Y (n_18398));
OAI21X1 g63105(.A0 (n_14077), .A1 (n_28832), .B0 (n_17706), .Y(n_18397));
NAND2X1 g63118(.A (n_15263), .B (n_6064), .Y (n_18396));
AND2X1 g63120(.A (n_18388), .B (n_18393), .Y (n_18394));
NAND3X1 g63123(.A (n_18391), .B (n_10003), .C (n_17005), .Y(n_18392));
NAND3X1 g63124(.A (n_10359), .B (n_18268), .C (n_10549), .Y(n_18390));
AND2X1 g63125(.A (n_18388), .B (n_13040), .Y (n_28890));
AND2X1 g63135(.A (n_18386), .B (n_18385), .Y (n_18387));
AOI21X1 g63139(.A0 (n_14558), .A1 (n_8379), .B0 (n_17260), .Y(n_18384));
AND2X1 g63141(.A (n_15314), .B (n_13083), .Y (n_18383));
NAND2X1 g63142(.A (n_16468), .B (n_3943), .Y (n_18382));
AND2X1 g63148(.A (n_16061), .B (n_7206), .Y (n_18381));
AOI21X1 g63152(.A0 (n_6084), .A1 (n_13083), .B0 (n_18375), .Y(n_18379));
INVX1 g63153(.A (n_17299), .Y (n_18377));
OR2X1 g63161(.A (n_11074), .B (n_18375), .Y (n_18376));
AOI21X1 g63165(.A0 (n_12627), .A1 (n_13466), .B0 (n_16904), .Y(n_18374));
NAND2X1 g63168(.A (n_15421), .B (n_14562), .Y (n_18372));
AND2X1 g63173(.A (n_15224), .B (n_18369), .Y (n_18370));
OAI21X1 g63176(.A0 (n_15992), .A1 (n_8820), .B0 (n_16787), .Y(n_18368));
OAI21X1 g63179(.A0 (n_14008), .A1 (n_14600), .B0 (n_14589), .Y(n_18367));
NAND2X1 g63183(.A (n_18365), .B (n_20634), .Y (n_18366));
OAI21X1 g63185(.A0 (n_16137), .A1 (n_6217), .B0 (n_18237), .Y(n_29303));
INVX1 g63186(.A (n_17281), .Y (n_18363));
AND2X1 g63188(.A (n_18361), .B (n_18360), .Y (n_18362));
NAND2X1 g63189(.A (n_16449), .B (n_1667), .Y (n_18359));
NAND2X1 g63190(.A (n_14502), .B (n_16848), .Y (n_18358));
NAND2X1 g63191(.A (n_15903), .B (n_503), .Y (n_18357));
NAND2X1 g63203(.A (n_17161), .B (n_21290), .Y (n_18356));
NAND2X1 g63204(.A (n_16717), .B (n_21151), .Y (n_18355));
NAND3X1 g63206(.A (n_10481), .B (n_18353), .C (n_10512), .Y(n_18354));
NAND2X1 g63212(.A (n_16443), .B (n_638), .Y (n_18352));
OR2X1 g63220(.A (n_16349), .B (n_17912), .Y (n_18351));
NAND2X1 g63224(.A (n_16436), .B (n_27493), .Y (n_18350));
NOR2X1 g63225(.A (n_16339), .B (n_14559), .Y (n_25512));
NOR2X1 g63229(.A (n_15241), .B (n_18347), .Y (n_18348));
NAND2X1 g73157(.A (n_15480), .B (n_19755), .Y (n_18346));
NAND3X1 g63234(.A (n_18316), .B (n_13028), .C (n_14669), .Y(n_18345));
AND2X1 g63240(.A (n_18343), .B (n_18342), .Y (n_18344));
OAI21X1 g63250(.A0 (n_14395), .A1 (n_17409), .B0 (n_17813), .Y(n_18341));
INVX1 g63251(.A (n_17245), .Y (n_18340));
INVX1 g63258(.A (n_17243), .Y (n_18339));
NAND3X1 g63269(.A (n_13686), .B (n_14666), .C (n_6347), .Y (n_18337));
NAND3X1 g63277(.A (n_10622), .B (n_18335), .C (n_12067), .Y(n_18336));
NAND2X1 g63279(.A (n_14832), .B (n_18333), .Y (n_18334));
AOI21X1 g63293(.A0 (n_14318), .A1 (n_8686), .B0 (n_27688), .Y(n_18329));
NAND2X1 g63296(.A (n_15069), .B (n_16103), .Y (n_18328));
OAI21X1 g63298(.A0 (n_14303), .A1 (n_10746), .B0 (n_18326), .Y(n_29417));
OAI21X1 g63301(.A0 (n_16013), .A1 (n_7824), .B0 (n_17414), .Y(n_18325));
INVX1 g63312(.A (n_17214), .Y (n_18324));
AND2X1 g63320(.A (n_15124), .B (n_11850), .Y (n_18323));
OAI21X1 g63321(.A0 (n_16044), .A1 (n_7969), .B0 (n_18320), .Y(n_29380));
NAND3X1 g63323(.A (sa22[1] ), .B (n_14069), .C (n_18320), .Y(n_18321));
NOR2X1 g63326(.A (n_16299), .B (n_11281), .Y (n_18319));
NAND2X1 g63339(.A (n_17922), .B (n_14639), .Y (n_18314));
OAI21X1 g63341(.A0 (n_16057), .A1 (n_7288), .B0 (n_16414), .Y(n_18313));
INVX1 g63348(.A (n_17207), .Y (n_18312));
NAND4X1 g63351(.A (n_16253), .B (n_14031), .C (n_18310), .D(n_13166), .Y (n_18311));
INVX1 g63352(.A (n_17205), .Y (n_18309));
OAI21X1 g63354(.A0 (n_15947), .A1 (n_7397), .B0 (n_17500), .Y(n_18308));
NAND3X1 g63356(.A (n_20585), .B (n_14070), .C (n_14155), .Y(n_18307));
AOI21X1 g63366(.A0 (n_14417), .A1 (n_14050), .B0 (n_15039), .Y(n_18304));
NAND2X1 g63373(.A (n_16372), .B (n_13324), .Y (n_18303));
AOI21X1 g63378(.A0 (n_14220), .A1 (n_13385), .B0 (n_9819), .Y(n_18302));
INVX1 g63384(.A (n_17193), .Y (n_18301));
NAND2X1 g63390(.A (n_15173), .B (sa12[1] ), .Y (n_18300));
INVX1 g63395(.A (n_17188), .Y (n_18297));
OAI21X1 g63399(.A0 (n_16003), .A1 (n_5487), .B0 (n_28692), .Y(n_18296));
NAND2X1 g63400(.A (n_16364), .B (n_18326), .Y (n_18295));
NAND2X1 g63402(.A (n_16327), .B (n_21242), .Y (n_18294));
INVX1 g63403(.A (n_17185), .Y (n_18293));
NAND2X1 g63413(.A (n_16326), .B (n_21174), .Y (n_18292));
NAND2X1 g63416(.A (n_15951), .B (n_17920), .Y (n_18290));
NAND2X1 g63417(.A (n_15115), .B (n_908), .Y (n_18289));
NAND2X1 g63423(.A (n_14160), .B (n_17882), .Y (n_18288));
NAND3X1 g63424(.A (n_10586), .B (n_18286), .C (n_10456), .Y(n_18287));
NAND2X1 g63427(.A (n_16332), .B (n_20862), .Y (n_18285));
NAND2X1 g63430(.A (n_16600), .B (n_903), .Y (n_25484));
NAND2X1 g63431(.A (n_16324), .B (n_1196), .Y (n_18283));
NAND2X1 g63434(.A (n_15944), .B (n_18281), .Y (n_18282));
NAND2X1 g63435(.A (n_14175), .B (n_17868), .Y (n_18280));
OAI21X1 g63443(.A0 (n_14134), .A1 (n_18278), .B0 (n_2895), .Y(n_18279));
INVX1 g63446(.A (n_17169), .Y (n_18277));
NAND3X1 g63449(.A (n_18275), .B (n_8554), .C (n_18465), .Y (n_18276));
INVX1 g63451(.A (n_17165), .Y (n_18274));
NOR2X1 g63453(.A (n_15147), .B (n_16563), .Y (n_18273));
NOR2X1 g63455(.A (n_16343), .B (n_17605), .Y (n_25583));
OAI21X1 g63457(.A0 (n_14001), .A1 (n_16266), .B0 (n_18237), .Y(n_18271));
NAND3X1 g63459(.A (n_15211), .B (n_12801), .C (n_16963), .Y(n_18270));
NAND3X1 g63461(.A (n_10359), .B (n_18268), .C (n_16068), .Y(n_18269));
AOI21X1 g63467(.A0 (n_14111), .A1 (n_14942), .B0 (n_18266), .Y(n_18267));
NAND2X1 g63474(.A (n_18298), .B (n_18264), .Y (n_18265));
INVX1 g63475(.A (n_17158), .Y (n_18263));
NAND2X1 g63479(.A (n_16337), .B (n_16527), .Y (n_18262));
NAND2X1 g63483(.A (n_14125), .B (n_17848), .Y (n_18261));
NAND2X1 g63487(.A (n_14270), .B (n_17835), .Y (n_18260));
INVX1 g63490(.A (n_17145), .Y (n_18259));
NOR2X1 g63495(.A (n_16676), .B (n_16515), .Y (n_18258));
OAI21X1 g63497(.A0 (n_15926), .A1 (n_9077), .B0 (n_18205), .Y(n_18257));
NOR2X1 g63504(.A (n_15227), .B (n_14455), .Y (n_18256));
OR2X1 g63514(.A (n_16317), .B (n_18254), .Y (n_18255));
NAND3X1 g63516(.A (n_16032), .B (n_10980), .C (n_9436), .Y (n_18253));
NAND3X1 g63519(.A (n_18251), .B (n_14304), .C (n_12576), .Y(n_18252));
NAND4X1 g63521(.A (n_17598), .B (n_18249), .C (n_15105), .D(n_18248), .Y (n_18250));
NOR2X1 g63524(.A (n_16681), .B (n_12769), .Y (n_25697));
NAND4X1 g63526(.A (n_18245), .B (n_18244), .C (n_15969), .D(n_18243), .Y (n_18246));
NAND4X1 g63528(.A (n_18241), .B (n_8642), .C (n_14336), .D (n_17456),.Y (n_18242));
INVX1 g63530(.A (n_17126), .Y (n_28259));
NAND3X1 g63538(.A (n_15950), .B (n_17879), .C (n_16537), .Y(n_18239));
AOI21X1 g63546(.A0 (n_14013), .A1 (n_16439), .B0 (n_18237), .Y(n_18238));
INVX1 g65372(.A (n_17345), .Y (n_18236));
AOI21X1 g63568(.A0 (n_13996), .A1 (n_8925), .B0 (n_18320), .Y(n_18235));
NAND2X1 g63580(.A (n_16696), .B (n_1368), .Y (n_18234));
NAND2X1 g63581(.A (n_16454), .B (n_1085), .Y (n_18233));
OAI21X1 g63584(.A0 (n_17851), .A1 (n_28843), .B0 (n_819), .Y(n_18232));
AND2X1 g63588(.A (n_15346), .B (n_5329), .Y (n_18231));
OAI21X1 g63592(.A0 (n_6058), .A1 (n_16797), .B0 (n_26874), .Y(n_18229));
NOR2X1 g63593(.A (n_15965), .B (n_11898), .Y (n_18228));
NAND2X1 g63596(.A (n_15333), .B (n_1547), .Y (n_18227));
AND2X1 g63597(.A (n_15341), .B (n_27688), .Y (n_18225));
AOI21X1 g63599(.A0 (n_12166), .A1 (n_877), .B0 (n_15309), .Y(n_18224));
OAI21X1 g63603(.A0 (n_18739), .A1 (n_4582), .B0 (n_18220), .Y(n_18221));
OAI21X1 g63606(.A0 (n_9214), .A1 (n_16480), .B0 (n_18217), .Y(n_18219));
OAI21X1 g63610(.A0 (n_6011), .A1 (n_17839), .B0 (n_28380), .Y(n_18216));
AND2X1 g63611(.A (n_15282), .B (n_15574), .Y (n_18215));
NAND2X1 g63612(.A (n_15279), .B (n_12986), .Y (n_18214));
AOI21X1 g63615(.A0 (n_16785), .A1 (n_430), .B0 (n_4845), .Y(n_18213));
OAI21X1 g63617(.A0 (n_28875), .A1 (n_12715), .B0 (n_27099), .Y(n_18212));
OAI21X1 g63620(.A0 (n_19568), .A1 (n_16466), .B0 (n_18210), .Y(n_18211));
NAND2X1 g63623(.A (n_15261), .B (n_18440), .Y (n_18209));
NAND2X1 g63624(.A (n_16493), .B (n_6941), .Y (n_18208));
AOI21X1 g63632(.A0 (n_14519), .A1 (n_11067), .B0 (n_6527), .Y(n_18207));
OAI21X1 g63633(.A0 (n_18038), .A1 (n_18205), .B0 (n_16828), .Y(n_18206));
AND2X1 g63638(.A (n_10099), .B (n_18203), .Y (n_18204));
NAND3X1 g63641(.A (n_16095), .B (n_14487), .C (n_12803), .Y(n_18202));
AOI21X1 g63645(.A0 (n_16503), .A1 (n_18199), .B0 (n_1667), .Y(n_18201));
NAND3X1 g63649(.A (n_16142), .B (n_18005), .C (n_16172), .Y(n_18197));
NOR2X1 g63651(.A (n_13415), .B (n_16448), .Y (n_18196));
NOR2X1 g63652(.A (n_16431), .B (n_12191), .Y (n_18195));
AOI21X1 g63656(.A0 (n_14074), .A1 (n_18645), .B0 (n_18679), .Y(n_18194));
NAND4X1 g63659(.A (n_15196), .B (n_9232), .C (n_12181), .D (n_11047),.Y (n_18193));
AOI21X1 g63661(.A0 (n_14159), .A1 (n_11110), .B0 (n_3281), .Y(n_18192));
NAND2X1 g63676(.A (n_15141), .B (n_17775), .Y (n_18189));
AND2X1 g63678(.A (n_15133), .B (n_28632), .Y (n_18188));
NAND2X1 g63685(.A (n_15122), .B (n_19395), .Y (n_28502));
OAI21X1 g63686(.A0 (n_28807), .A1 (n_12496), .B0 (n_17567), .Y(n_28263));
OAI21X1 g63693(.A0 (n_14346), .A1 (n_14484), .B0 (n_11843), .Y(n_18184));
OAI21X1 g63697(.A0 (n_14334), .A1 (n_10333), .B0 (n_12858), .Y(n_18183));
NAND2X1 g63698(.A (n_15096), .B (n_19857), .Y (n_18182));
NAND2X1 g63702(.A (n_15082), .B (n_29048), .Y (n_18181));
NAND2X1 g63704(.A (n_16404), .B (n_9802), .Y (n_18179));
AOI21X1 g63705(.A0 (n_14316), .A1 (n_12436), .B0 (n_4208), .Y(n_18177));
OAI21X1 g63707(.A0 (n_18043), .A1 (n_27688), .B0 (n_16865), .Y(n_18176));
NAND2X1 g63710(.A (n_15071), .B (n_21242), .Y (n_18174));
NAND2X1 g63711(.A (n_15066), .B (n_28642), .Y (n_18173));
AOI21X1 g63712(.A0 (n_12146), .A1 (n_2001), .B0 (n_16721), .Y(n_18172));
NAND3X1 g63720(.A (n_15991), .B (n_14263), .C (n_12347), .Y(n_18170));
NAND2X1 g63721(.A (n_16694), .B (n_18168), .Y (n_18169));
NAND2X1 g63724(.A (n_16395), .B (n_1928), .Y (n_28585));
NAND2X1 g63727(.A (n_16687), .B (n_29062), .Y (n_18163));
OAI21X1 g63728(.A0 (n_14461), .A1 (n_27431), .B0 (n_8846), .Y(n_18162));
OAI21X1 g63729(.A0 (n_18598), .A1 (n_29048), .B0 (n_17632), .Y(n_18161));
NAND2X1 g63730(.A (n_16684), .B (n_28645), .Y (n_18160));
NAND3X1 g63739(.A (n_12461), .B (n_14581), .C (n_12177), .Y(n_18157));
NAND3X1 g63741(.A (n_29369), .B (n_12095), .C (n_29370), .Y(n_18156));
AND2X1 g63744(.A (n_16655), .B (n_16835), .Y (n_18155));
NAND4X1 g63747(.A (n_18153), .B (n_5652), .C (n_11792), .D (n_7359),.Y (n_18154));
OAI21X1 g63750(.A0 (n_18151), .A1 (n_688), .B0 (n_21227), .Y(n_18152));
NAND2X1 g63751(.A (n_15287), .B (n_20116), .Y (n_18150));
NAND2X1 g63769(.A (n_16602), .B (n_19896), .Y (n_18148));
NAND2X1 g63772(.A (n_16594), .B (n_11576), .Y (n_18147));
NAND2X1 g63773(.A (n_16535), .B (n_15894), .Y (n_18145));
NAND3X1 g63775(.A (n_5717), .B (n_14066), .C (n_18142), .Y (n_18143));
NOR2X1 g63780(.A (n_15393), .B (n_15424), .Y (n_18141));
AOI21X1 g63794(.A0 (n_12149), .A1 (n_1756), .B0 (n_15214), .Y(n_18140));
NAND3X1 g63795(.A (n_29301), .B (n_29302), .C (n_15687), .Y(n_18138));
AND2X1 g63796(.A (n_16528), .B (n_18205), .Y (n_18137));
NAND2X1 g63798(.A (n_16525), .B (n_14474), .Y (n_18136));
AOI21X1 g63800(.A0 (n_13959), .A1 (n_1196), .B0 (n_14842), .Y(n_18134));
NAND2X1 g63801(.A (n_16520), .B (n_18440), .Y (n_29368));
NAND4X1 g63803(.A (n_17990), .B (n_7807), .C (n_12170), .D (n_12445),.Y (n_18130));
NAND2X1 g63805(.A (n_16511), .B (n_19934), .Y (n_18129));
NAND2X1 g63811(.A (n_13628), .B (n_15384), .Y (n_18127));
OR2X1 g63812(.A (n_13625), .B (n_15381), .Y (n_18126));
OR2X1 g63815(.A (n_15437), .B (n_15376), .Y (n_18125));
NAND4X1 g63825(.A (n_16229), .B (n_7222), .C (n_13965), .D (n_9948),.Y (n_18123));
NAND2X1 g63830(.A (n_16607), .B (n_18121), .Y (n_18122));
NAND2X1 g63834(.A (n_16571), .B (n_18119), .Y (n_18120));
NAND4X1 g63836(.A (n_17236), .B (n_11925), .C (n_25463), .D(n_10170), .Y (n_18118));
NAND4X1 g63838(.A (n_15285), .B (n_18116), .C (n_18115), .D(n_18114), .Y (n_18117));
NAND4X1 g63840(.A (n_11374), .B (n_11550), .C (n_5645), .D (n_16927),.Y (n_18113));
NAND4X1 g63841(.A (n_17754), .B (n_18048), .C (n_11543), .D(n_18047), .Y (n_18112));
NAND4X1 g63845(.A (n_10785), .B (n_18064), .C (n_16959), .D(n_18063), .Y (n_18111));
NOR2X1 g63859(.A (n_8847), .B (n_15143), .Y (n_18110));
NAND3X1 g63862(.A (n_15207), .B (n_17121), .C (n_9896), .Y (n_18109));
NAND4X1 g63863(.A (n_11011), .B (n_18061), .C (n_13487), .D(n_18060), .Y (n_18108));
NOR2X1 g63865(.A (n_10457), .B (n_16541), .Y (n_18107));
NAND3X1 g63867(.A (n_15317), .B (n_15708), .C (n_487), .Y (n_18106));
NAND3X1 g63868(.A (n_15188), .B (n_19398), .C (n_20810), .Y(n_18105));
NAND3X1 g63869(.A (n_15086), .B (n_15039), .C (n_778), .Y (n_18104));
OAI21X1 g63872(.A0 (n_14015), .A1 (n_11150), .B0 (n_18102), .Y(n_18103));
OR2X1 g63873(.A (n_16505), .B (n_18100), .Y (n_18101));
OAI21X1 g63875(.A0 (n_14010), .A1 (n_12792), .B0 (n_20105), .Y(n_18099));
NOR2X1 g63879(.A (n_16102), .B (n_16910), .Y (n_18098));
NOR2X1 g63883(.A (n_12759), .B (n_16908), .Y (n_18097));
OR2X1 g63884(.A (n_16504), .B (n_17023), .Y (n_18096));
OAI21X1 g63888(.A0 (n_13994), .A1 (n_11010), .B0 (n_18094), .Y(n_18095));
OR2X1 g63889(.A (n_16502), .B (n_17020), .Y (n_18093));
OAI21X1 g63892(.A0 (n_13999), .A1 (n_12694), .B0 (n_20065), .Y(n_18092));
NOR2X1 g63893(.A (n_14466), .B (n_16897), .Y (n_18091));
NOR2X1 g63894(.A (n_14349), .B (n_16891), .Y (n_18090));
NOR2X1 g63895(.A (n_16022), .B (n_15420), .Y (n_18089));
NAND2X1 g63896(.A (n_16499), .B (n_18087), .Y (n_18088));
OAI21X1 g63899(.A0 (n_10682), .A1 (n_4755), .B0 (n_18085), .Y(n_18086));
NOR2X1 g63902(.A (n_12488), .B (n_18083), .Y (n_18084));
NOR2X1 g63906(.A (n_12403), .B (n_16365), .Y (n_18082));
OR2X1 g63909(.A (n_17017), .B (n_16495), .Y (n_18081));
NAND2X1 g63912(.A (n_16514), .B (n_18094), .Y (n_18080));
AOI22X1 g63923(.A0 (n_14064), .A1 (n_19364), .B0 (n_16006), .B1(n_8524), .Y (n_18073));
AOI22X1 g63930(.A0 (n_14060), .A1 (n_28642), .B0 (n_2112), .B1(n_6368), .Y (n_25637));
NOR2X1 g63935(.A (n_12733), .B (n_15456), .Y (n_18071));
NAND3X1 g63944(.A (n_14543), .B (n_12254), .C (n_27802), .Y(n_18070));
NAND3X1 g63946(.A (n_15994), .B (n_13110), .C (n_28221), .Y(n_18069));
NAND3X1 g63947(.A (n_15190), .B (n_13109), .C (n_28257), .Y(n_18068));
NAND3X1 g63948(.A (n_28247), .B (n_28248), .C (n_16661), .Y(n_18067));
NAND3X1 g63949(.A (n_14400), .B (n_14728), .C (n_17904), .Y(n_18066));
NAND4X1 g63952(.A (n_19953), .B (n_18064), .C (n_18063), .D(n_20078), .Y (n_18065));
NAND4X1 g63956(.A (n_19955), .B (n_18061), .C (n_18060), .D(n_11517), .Y (n_18062));
NOR2X1 g63959(.A (n_16705), .B (n_13317), .Y (n_18059));
NAND3X1 g63960(.A (n_16038), .B (n_13105), .C (n_16642), .Y(n_18058));
NAND3X1 g63962(.A (n_15972), .B (n_14041), .C (n_26050), .Y(n_18057));
NAND3X1 g63965(.A (n_15983), .B (n_11404), .C (n_25858), .Y(n_18054));
NAND3X1 g63966(.A (n_12475), .B (n_14033), .C (n_12474), .Y(n_18053));
NAND4X1 g63971(.A (n_15068), .B (n_18051), .C (n_18050), .D(n_11461), .Y (n_18052));
NAND4X1 g63976(.A (n_19428), .B (n_18048), .C (n_18047), .D(n_18046), .Y (n_18049));
NAND4X1 g63977(.A (n_15260), .B (n_11714), .C (n_6363), .D (n_15259),.Y (n_18045));
NAND3X1 g63978(.A (n_9136), .B (n_18043), .C (n_11154), .Y (n_18044));
NAND3X1 g63980(.A (n_15348), .B (n_13093), .C (n_11473), .Y(n_18042));
NOR2X1 g63981(.A (n_15332), .B (n_15330), .Y (n_18041));
NAND3X1 g63984(.A (n_16555), .B (n_13043), .C (n_13217), .Y(n_18040));
NAND3X1 g63986(.A (n_8932), .B (n_18038), .C (n_12312), .Y (n_18039));
NOR2X1 g63987(.A (n_15199), .B (n_13448), .Y (n_18037));
NOR2X1 g63991(.A (n_15108), .B (n_13393), .Y (n_18036));
NAND3X1 g63994(.A (n_16726), .B (n_27144), .C (n_10691), .Y(n_18035));
NOR2X1 g63999(.A (n_11240), .B (n_16622), .Y (n_18033));
AOI21X1 g64001(.A0 (n_14188), .A1 (n_1057), .B0 (n_16617), .Y(n_18032));
AND2X1 g64021(.A (n_15152), .B (n_10342), .Y (n_25504));
NAND2X1 g64027(.A (n_14779), .B (n_15445), .Y (n_18028));
AOI21X1 g64030(.A0 (n_15021), .A1 (n_29102), .B0 (n_16708), .Y(n_18027));
XOR2X1 g76192(.A (text_in_r[27] ), .B (n_1626), .Y (n_18026));
XOR2X1 g76235(.A (text_in_r[10] ), .B (n_19445), .Y (n_18024));
XOR2X1 g76279(.A (text_in_r[3] ), .B (n_14878), .Y (n_18023));
INVX1 g64120(.A (n_16913), .Y (n_18862));
NOR2X1 g64150(.A (n_18826), .B (n_27688), .Y (n_18021));
OR2X1 g64153(.A (n_18018), .B (n_7410), .Y (n_18019));
NOR2X1 g64164(.A (n_15091), .B (n_20325), .Y (n_19643));
INVX1 g64198(.A (n_18016), .Y (n_18017));
INVX1 g64256(.A (n_16877), .Y (n_18013));
NAND4X1 g64279(.A (n_16100), .B (n_15596), .C (n_16391), .D(n_10632), .Y (n_18012));
INVX1 g64280(.A (n_18010), .Y (n_18011));
OR2X1 g64283(.A (n_15870), .B (n_18205), .Y (n_18009));
NAND2X1 g64310(.A (n_16138), .B (n_18005), .Y (n_25733));
INVX1 g64313(.A (n_16855), .Y (n_18004));
NAND2X1 g64321(.A (n_15993), .B (n_17071), .Y (n_18003));
OR2X1 g64328(.A (n_16134), .B (n_16787), .Y (n_18002));
NAND2X1 g64343(.A (n_18000), .B (n_27446), .Y (n_18001));
NAND2X1 g64348(.A (n_16079), .B (n_16711), .Y (n_17999));
NAND2X1 g64349(.A (n_16133), .B (n_15236), .Y (n_17998));
NAND2X1 g64365(.A (n_17649), .B (n_17104), .Y (n_18852));
NAND2X1 g64390(.A (n_16116), .B (n_13575), .Y (n_17997));
INVX1 g64428(.A (n_17995), .Y (n_17996));
AND2X1 g64431(.A (n_16096), .B (n_16480), .Y (n_19679));
INVX1 g64465(.A (n_16809), .Y (n_17993));
NAND2X1 g64480(.A (n_16110), .B (n_16466), .Y (n_18849));
OR2X1 g64504(.A (n_15869), .B (n_27688), .Y (n_17992));
AND2X1 g64509(.A (n_17990), .B (n_18765), .Y (n_17991));
NAND2X1 g64519(.A (n_16118), .B (n_11261), .Y (n_17989));
NOR2X1 g64523(.A (n_14227), .B (n_15048), .Y (n_17987));
NAND2X1 g64557(.A (n_15948), .B (n_17041), .Y (n_17986));
NOR2X1 g64573(.A (n_12855), .B (n_15922), .Y (n_17985));
NOR2X1 g64577(.A (n_11191), .B (n_10489), .Y (n_17984));
NAND2X1 g64615(.A (n_17982), .B (n_14587), .Y (n_17983));
AND2X1 g64627(.A (n_17980), .B (n_17979), .Y (n_17981));
NAND2X1 g64628(.A (n_16058), .B (n_10947), .Y (n_17978));
NAND3X1 g64653(.A (n_29179), .B (n_27779), .C (n_13277), .Y(n_17977));
NAND2X1 g64659(.A (n_8186), .B (n_17979), .Y (n_17975));
NAND2X1 g64680(.A (n_15864), .B (n_1196), .Y (n_17974));
NAND2X1 g64681(.A (n_17972), .B (n_15091), .Y (n_17973));
AND2X1 g64683(.A (n_17969), .B (n_18811), .Y (n_17970));
OR2X1 g64698(.A (n_27969), .B (n_29062), .Y (n_17968));
NAND2X1 g64702(.A (n_15985), .B (n_14589), .Y (n_17966));
NOR2X1 g64703(.A (n_12996), .B (n_12894), .Y (n_28254));
NAND2X1 g64711(.A (n_16045), .B (n_15539), .Y (n_17963));
AOI21X1 g64712(.A0 (n_13857), .A1 (n_8094), .B0 (n_2800), .Y(n_17962));
INVX1 g64713(.A (n_17960), .Y (n_17961));
NAND2X1 g64725(.A (n_16406), .B (n_17292), .Y (n_17958));
INVX1 g64732(.A (n_17955), .Y (n_17956));
NAND2X1 g64744(.A (n_16037), .B (n_624), .Y (n_17954));
AOI21X1 g64757(.A0 (n_13800), .A1 (n_9685), .B0 (n_27028), .Y(n_29400));
OR2X1 g64760(.A (n_15867), .B (n_28642), .Y (n_17951));
OR2X1 g64776(.A (n_15878), .B (n_8708), .Y (n_17950));
AOI21X1 g64795(.A0 (n_13853), .A1 (n_6087), .B0 (n_15039), .Y(n_17948));
NAND2X1 g64816(.A (n_16014), .B (n_10202), .Y (n_17944));
OR2X1 g64818(.A (n_15920), .B (n_29062), .Y (n_17943));
NAND4X1 g64833(.A (n_10609), .B (n_16070), .C (n_17762), .D(n_12093), .Y (n_17942));
NAND2X1 g64845(.A (n_17939), .B (n_17832), .Y (n_17940));
OAI21X1 g64852(.A0 (n_11760), .A1 (n_15636), .B0 (n_9819), .Y(n_17938));
NOR2X1 g64854(.A (n_14053), .B (n_10078), .Y (n_17937));
NAND3X1 g64872(.A (n_13885), .B (n_5105), .C (n_17935), .Y (n_17936));
NAND2X1 g64878(.A (n_13982), .B (n_17933), .Y (n_17934));
INVX1 g64882(.A (n_16714), .Y (n_17932));
NAND3X1 g64886(.A (n_13838), .B (n_9406), .C (n_4767), .Y (n_17931));
NAND2X1 g64896(.A (n_17929), .B (n_13695), .Y (n_17930));
OR2X1 g64899(.A (n_14273), .B (n_15568), .Y (n_17928));
NAND2X1 g64902(.A (n_16030), .B (n_28645), .Y (n_18978));
NOR2X1 g64904(.A (n_12614), .B (n_16128), .Y (n_17927));
NOR2X1 g64906(.A (n_6944), .B (n_11325), .Y (n_17926));
NAND2X1 g64907(.A (n_13980), .B (n_28632), .Y (n_17925));
NAND2X1 g64909(.A (n_11273), .B (n_28642), .Y (n_17924));
INVX1 g64914(.A (n_17922), .Y (n_17923));
INVX1 g64933(.A (n_17920), .Y (n_17921));
NAND2X1 g65382(.A (n_14575), .B (n_12865), .Y (n_17919));
INVX1 g64968(.A (n_16679), .Y (n_17918));
NOR2X1 g64973(.A (n_7083), .B (n_16159), .Y (n_28313));
NAND3X1 g64977(.A (n_17915), .B (n_17723), .C (n_16271), .Y(n_17916));
AND2X1 g64978(.A (n_11050), .B (n_17912), .Y (n_17914));
AOI21X1 g64981(.A0 (n_15952), .A1 (n_7372), .B0 (n_14807), .Y(n_17911));
INVX1 g64993(.A (n_16659), .Y (n_17910));
NAND3X1 g65029(.A (n_17906), .B (n_17776), .C (n_16236), .Y(n_17907));
NOR2X1 g65036(.A (n_7352), .B (n_27970), .Y (n_17902));
NOR2X1 g65038(.A (n_14209), .B (n_17900), .Y (n_17901));
NOR2X1 g65039(.A (n_14319), .B (n_17692), .Y (n_17899));
NAND3X1 g65048(.A (n_17888), .B (n_14138), .C (n_17897), .Y(n_17898));
NAND2X1 g65049(.A (n_14508), .B (n_17414), .Y (n_17896));
NOR2X1 g65084(.A (n_5522), .B (n_26802), .Y (n_17894));
OR2X1 g65086(.A (n_16683), .B (n_28642), .Y (n_17893));
AND2X1 g65087(.A (n_16683), .B (n_17037), .Y (n_17890));
NAND2X1 g65099(.A (n_17888), .B (n_18286), .Y (n_17889));
NOR2X1 g65103(.A (n_12366), .B (n_15934), .Y (n_17887));
NAND2X1 g65113(.A (n_14029), .B (n_29014), .Y (n_17886));
AOI22X1 g65116(.A0 (n_11946), .A1 (n_17884), .B0 (n_1365), .B1(n_11831), .Y (n_25817));
INVX1 g65118(.A (n_17882), .Y (n_17883));
NAND2X1 g65120(.A (n_14169), .B (n_3483), .Y (n_17881));
OR2X1 g65123(.A (n_17879), .B (n_1008), .Y (n_17880));
INVX1 g65126(.A (n_27312), .Y (n_17877));
NOR2X1 g65131(.A (n_16503), .B (n_13606), .Y (n_17875));
NOR2X1 g65140(.A (n_6897), .B (n_27450), .Y (n_28559));
NAND2X1 g65147(.A (n_17040), .B (n_14650), .Y (n_17872));
INVX1 g65155(.A (n_16589), .Y (n_29387));
NAND2X1 g65158(.A (n_14147), .B (n_17912), .Y (n_18817));
INVX1 g65161(.A (n_17868), .Y (n_17869));
NAND2X1 g65165(.A (n_16196), .B (n_10037), .Y (n_17867));
NOR2X1 g65172(.A (n_12747), .B (n_16009), .Y (n_17866));
NAND2X1 g65197(.A (n_13979), .B (n_21275), .Y (n_17865));
NAND2X1 g65198(.A (n_15932), .B (n_17864), .Y (n_19052));
NAND2X1 g65203(.A (n_11291), .B (n_18320), .Y (n_17863));
NAND2X1 g65205(.A (n_13990), .B (n_18320), .Y (n_17862));
OR2X1 g65208(.A (n_15984), .B (n_4851), .Y (n_17861));
AOI21X1 g65209(.A0 (n_11753), .A1 (n_9694), .B0 (n_4851), .Y(n_17860));
NOR2X1 g65212(.A (n_11208), .B (n_10603), .Y (n_17858));
NAND2X1 g65229(.A (n_14108), .B (n_16835), .Y (n_17856));
INVX1 g65233(.A (n_16538), .Y (n_17854));
NAND2X1 g65246(.A (n_17851), .B (n_5558), .Y (n_17852));
NOR2X1 g65251(.A (n_5762), .B (n_16126), .Y (n_17850));
INVX1 g65254(.A (n_17848), .Y (n_17849));
AOI21X1 g65263(.A0 (n_11746), .A1 (n_8091), .B0 (n_1610), .Y(n_17847));
NAND2X1 g65267(.A (n_13984), .B (n_21442), .Y (n_17846));
NAND2X1 g65273(.A (n_10052), .B (n_17844), .Y (n_17845));
OR2X1 g65276(.A (n_13977), .B (n_20157), .Y (n_17843));
AND2X1 g65279(.A (n_17841), .B (n_16084), .Y (n_17842));
NAND2X1 g65281(.A (n_17839), .B (n_28444), .Y (n_17840));
OR2X1 g65283(.A (n_13975), .B (n_15574), .Y (n_17838));
NOR2X1 g65284(.A (n_15299), .B (n_14687), .Y (n_17837));
INVX1 g65290(.A (n_17835), .Y (n_17836));
NAND3X1 g65295(.A (n_7039), .B (n_8824), .C (n_15966), .Y (n_17834));
NAND2X1 g65301(.A (n_17832), .B (n_8852), .Y (n_17833));
NAND2X1 g65305(.A (n_14115), .B (n_15113), .Y (n_17831));
OR2X1 g65307(.A (n_13973), .B (n_15776), .Y (n_17830));
NAND2X1 g65316(.A (n_18645), .B (n_17325), .Y (n_17828));
NAND3X1 g65329(.A (n_11539), .B (n_12102), .C (n_9048), .Y (n_17827));
NAND2X1 g65338(.A (n_13997), .B (n_17824), .Y (n_17825));
NAND3X1 g65351(.A (n_13322), .B (n_12015), .C (n_20626), .Y(n_17823));
NAND3X1 g65356(.A (n_17821), .B (n_11999), .C (n_12113), .Y(n_17822));
OR2X1 g65357(.A (n_14004), .B (n_18641), .Y (n_17820));
OR2X1 g65397(.A (n_14580), .B (n_12731), .Y (n_17819));
NOR2X1 g65367(.A (n_12703), .B (n_14063), .Y (n_17818));
NAND4X1 g65368(.A (n_10311), .B (n_5716), .C (n_14657), .D (n_6137),.Y (n_17817));
NOR2X1 g65369(.A (n_14583), .B (n_14056), .Y (n_17816));
NOR2X1 g65370(.A (n_14414), .B (n_14027), .Y (n_17815));
NAND2X1 g65403(.A (n_14419), .B (n_17813), .Y (n_17814));
DFFX1 dcnt_reg[3] (.CK (clk), .D (n_15041), .Q (dcnt[3] ), .QN ());
NAND2X1 g65424(.A (n_14682), .B (n_14841), .Y (n_17812));
NAND2X1 g65440(.A (n_14232), .B (n_26670), .Y (n_17811));
AOI21X1 g65446(.A0 (n_13825), .A1 (n_12578), .B0 (n_17567), .Y(n_17809));
INVX1 g65449(.A (n_16471), .Y (n_17808));
AOI21X1 g65452(.A0 (n_16130), .A1 (n_28728), .B0 (n_13915), .Y(n_17807));
AND2X1 g65454(.A (n_4626), .B (n_16902), .Y (n_17806));
INVX1 g65457(.A (n_16467), .Y (n_17805));
AOI21X1 g65465(.A0 (n_14290), .A1 (n_3503), .B0 (n_12098), .Y(n_17804));
NAND2X1 g65467(.A (n_14121), .B (n_12329), .Y (n_17803));
AND2X1 g65470(.A (n_14554), .B (n_14589), .Y (n_17802));
AND2X1 g65472(.A (n_14158), .B (n_11603), .Y (n_17801));
NOR2X1 g65473(.A (n_10858), .B (n_14058), .Y (n_17799));
INVX1 g65474(.A (n_16460), .Y (n_17798));
INVX1 g65478(.A (n_16459), .Y (n_17797));
AOI21X1 g65480(.A0 (n_11683), .A1 (n_1198), .B0 (n_10414), .Y(n_17796));
AND2X1 g65481(.A (n_5796), .B (n_16889), .Y (n_17795));
INVX1 g65496(.A (n_16455), .Y (n_17794));
NAND3X1 g65499(.A (n_4145), .B (n_10091), .C (n_4017), .Y (n_17793));
AOI21X1 g65502(.A0 (n_9322), .A1 (n_18369), .B0 (n_12922), .Y(n_17792));
AND2X1 g65506(.A (n_14532), .B (n_7173), .Y (n_17791));
INVX1 g65514(.A (n_16447), .Y (n_17790));
INVX1 g65533(.A (n_16440), .Y (n_17789));
NAND4X1 g61207(.A (n_10994), .B (n_10843), .C (n_9330), .D (n_9789),.Y (n_17788));
AND2X1 g65535(.A (n_14557), .B (n_14142), .Y (n_17787));
NAND2X1 g65541(.A (n_14430), .B (n_17912), .Y (n_17786));
NAND2X1 g65542(.A (n_14351), .B (n_10785), .Y (n_17785));
NAND2X1 g65544(.A (n_12650), .B (n_9821), .Y (n_17783));
NAND2X1 g65550(.A (n_14137), .B (n_15278), .Y (n_17782));
OR2X1 g65554(.A (n_15741), .B (n_14653), .Y (n_17781));
NAND2X1 g65555(.A (n_14426), .B (n_18205), .Y (n_28852));
AOI21X1 g65571(.A0 (n_17776), .A1 (n_11743), .B0 (n_17775), .Y(n_17777));
NAND4X1 g65580(.A (n_17773), .B (n_5682), .C (n_11725), .D (n_7427),.Y (n_17774));
NAND2X1 g65581(.A (n_14171), .B (n_15064), .Y (n_17772));
NAND2X1 g65585(.A (n_14369), .B (n_18168), .Y (n_17771));
OR2X1 g65587(.A (n_14365), .B (n_8708), .Y (n_17770));
NAND2X1 g65598(.A (n_14317), .B (n_21598), .Y (n_17768));
NAND2X1 g65612(.A (n_14140), .B (n_27688), .Y (n_25535));
INVX1 g65619(.A (n_16403), .Y (n_17765));
NAND2X1 g65621(.A (n_14307), .B (n_14038), .Y (n_17764));
NAND3X1 g65626(.A (n_17762), .B (n_11931), .C (n_17621), .Y(n_17763));
NAND2X1 g65628(.A (n_14579), .B (n_17760), .Y (n_17761));
NOR2X1 g65637(.A (n_12507), .B (n_14059), .Y (n_17759));
NAND2X1 g65638(.A (n_14412), .B (n_17757), .Y (n_17758));
NAND3X1 g65643(.A (n_11816), .B (n_28136), .C (n_908), .Y (n_17756));
AND2X1 g65649(.A (n_14555), .B (n_17754), .Y (n_17755));
AOI21X1 g65651(.A0 (n_17752), .A1 (n_16883), .B0 (n_19934), .Y(n_17753));
NAND2X1 g65656(.A (n_14439), .B (n_29074), .Y (n_25796));
NAND2X1 g65658(.A (n_13781), .B (n_16331), .Y (n_17750));
NAND2X1 g65660(.A (n_13820), .B (n_16323), .Y (n_17749));
NAND2X1 g65661(.A (n_14241), .B (n_28632), .Y (n_17748));
INVX1 g65663(.A (n_16389), .Y (n_17747));
INVX1 g65666(.A (n_16387), .Y (n_17746));
NAND4X1 g65669(.A (n_17058), .B (n_5664), .C (n_17744), .D (n_7545),.Y (n_17745));
AND2X1 g65676(.A (n_14233), .B (n_16680), .Y (n_17743));
AND2X1 g65679(.A (n_14230), .B (n_11251), .Y (n_17742));
INVX1 g65681(.A (n_16383), .Y (n_17741));
NOR2X1 g65683(.A (n_10906), .B (n_14032), .Y (n_17740));
NAND3X1 g65687(.A (n_25861), .B (n_12973), .C (n_13181), .Y(n_17739));
INVX1 g65690(.A (n_16379), .Y (n_17738));
INVX1 g65701(.A (n_16374), .Y (n_17737));
AND2X1 g65707(.A (n_12280), .B (n_17125), .Y (n_17736));
NAND2X1 g65711(.A (n_7330), .B (n_17734), .Y (n_17735));
INVX1 g65712(.A (n_16371), .Y (n_17733));
NAND2X1 g65714(.A (n_10318), .B (n_16767), .Y (n_17732));
NOR2X1 g65720(.A (n_14203), .B (n_13998), .Y (n_17731));
AND2X1 g65721(.A (n_14200), .B (n_14964), .Y (n_17730));
NOR2X1 g65722(.A (n_14196), .B (n_10707), .Y (n_17729));
NOR2X1 g65723(.A (n_12413), .B (n_14006), .Y (n_17728));
AND2X1 g65724(.A (n_14195), .B (n_20626), .Y (n_17727));
AND2X1 g65730(.A (n_14486), .B (n_17725), .Y (n_17726));
AOI21X1 g65739(.A0 (n_17723), .A1 (n_13773), .B0 (n_17089), .Y(n_17724));
AND2X1 g65747(.A (n_14424), .B (n_19842), .Y (n_17722));
INVX1 g65749(.A (n_16356), .Y (n_17721));
INVX1 g65751(.A (n_16355), .Y (n_17720));
INVX1 g65754(.A (n_16354), .Y (n_17719));
AOI21X1 g65756(.A0 (n_17717), .A1 (n_11190), .B0 (n_12850), .Y(n_17718));
NAND2X1 g65764(.A (n_14149), .B (n_15140), .Y (n_17716));
NOR2X1 g65772(.A (n_12724), .B (n_14034), .Y (n_17715));
INVX1 g65773(.A (n_16345), .Y (n_17714));
INVX1 g65780(.A (n_16341), .Y (n_17713));
AOI21X1 g65784(.A0 (n_15238), .A1 (n_5313), .B0 (n_18237), .Y(n_17712));
NAND3X1 g65785(.A (n_14697), .B (n_29336), .C (n_6344), .Y (n_17710));
NAND2X1 g65793(.A (n_14112), .B (n_13556), .Y (n_17708));
NAND2X1 g65801(.A (n_14101), .B (n_17706), .Y (n_17707));
NAND2X1 g65821(.A (n_14075), .B (n_17571), .Y (n_17705));
AND2X1 g65831(.A (n_14068), .B (n_17703), .Y (n_17704));
NAND2X1 g65838(.A (n_14718), .B (n_11738), .Y (n_17702));
NAND2X1 g65840(.A (n_14705), .B (n_8538), .Y (n_17701));
OAI21X1 g65843(.A0 (n_10091), .A1 (n_18792), .B0 (n_7180), .Y(n_17700));
NOR2X1 g65869(.A (n_14275), .B (n_11150), .Y (n_17698));
MX2X1 g65872(.A (n_11078), .B (n_11670), .S0 (n_26276), .Y (n_17697));
NOR2X1 g65873(.A (n_6779), .B (n_14293), .Y (n_17695));
NOR2X1 g65875(.A (n_14259), .B (n_12694), .Y (n_17694));
AOI21X1 g65878(.A0 (n_16245), .A1 (n_9959), .B0 (n_17692), .Y(n_17693));
AOI21X1 g65894(.A0 (n_4233), .A1 (n_15588), .B0 (n_13963), .Y(n_17691));
NAND4X1 g65912(.A (n_8648), .B (n_17689), .C (n_8814), .D (n_16338),.Y (n_17690));
NAND3X1 g65916(.A (n_12387), .B (n_17687), .C (n_8934), .Y (n_17688));
NAND4X1 g65918(.A (n_17685), .B (n_9350), .C (n_13532), .D (n_9208),.Y (n_17686));
NAND4X1 g65919(.A (n_9211), .B (n_9573), .C (n_10943), .D (n_17683),.Y (n_17684));
NAND4X1 g65920(.A (n_9951), .B (n_17681), .C (n_16416), .D (n_16342),.Y (n_17682));
NAND2X1 g65933(.A (n_14105), .B (n_9910), .Y (n_17680));
NAND2X1 g65935(.A (n_14322), .B (n_8233), .Y (n_17679));
NAND2X1 g65945(.A (n_7320), .B (n_14652), .Y (n_17678));
NAND2X1 g65950(.A (n_9514), .B (n_14648), .Y (n_17677));
NOR3X1 g65987(.A (n_12896), .B (n_15812), .C (n_11728), .Y (n_17676));
NOR3X1 g66055(.A (n_12298), .B (n_15800), .C (n_15799), .Y (n_17675));
CLKBUFX2 g66217(.A (n_17672), .Y (n_18859));
INVX1 g66463(.A (n_18996), .Y (n_17669));
NAND2X1 g66469(.A (n_17588), .B (n_26879), .Y (n_17668));
INVX1 g66495(.A (n_16213), .Y (n_19604));
NAND2X1 g66511(.A (n_12635), .B (n_9264), .Y (n_17667));
NAND2X1 g66555(.A (n_15846), .B (n_16434), .Y (n_17665));
NOR2X1 g66679(.A (n_13849), .B (n_27688), .Y (n_17659));
INVX1 g66713(.A (n_16177), .Y (n_17658));
NAND2X1 g66739(.A (n_15816), .B (n_13247), .Y (n_17657));
NAND2X1 g66840(.A (n_19071), .B (n_15817), .Y (n_17652));
OR2X1 g66842(.A (n_7724), .B (n_13826), .Y (n_17651));
INVX1 g66844(.A (n_17649), .Y (n_17650));
NAND2X1 g61587(.A (n_13949), .B (n_13083), .Y (n_17647));
INVX1 g66902(.A (n_17645), .Y (n_17646));
NOR2X1 g67016(.A (n_12823), .B (n_18164), .Y (n_17642));
AND2X1 g67031(.A (n_15002), .B (n_12052), .Y (n_17641));
OR2X1 g67051(.A (n_7253), .B (n_13881), .Y (n_17640));
OR2X1 g67066(.A (n_11710), .B (n_29065), .Y (n_28275));
OR2X1 g67069(.A (n_18151), .B (n_12986), .Y (n_17638));
NAND2X1 g67094(.A (n_10316), .B (n_9084), .Y (n_17636));
OR2X1 g67112(.A (n_11701), .B (n_11261), .Y (n_17635));
NAND2X1 g67208(.A (n_11898), .B (n_11261), .Y (n_17634));
INVX1 g67212(.A (n_17632), .Y (n_17633));
NAND4X1 g61698(.A (n_8465), .B (n_17683), .C (n_11437), .D (n_3758),.Y (n_17629));
NAND2X1 g67293(.A (n_14082), .B (n_15894), .Y (n_18967));
INVX1 g67329(.A (n_16077), .Y (n_17628));
NAND2X1 g67340(.A (n_15847), .B (n_16835), .Y (n_18914));
OR2X1 g67392(.A (n_11821), .B (n_19398), .Y (n_17626));
INVX1 g67410(.A (n_17624), .Y (n_17625));
NOR2X1 g67412(.A (n_10229), .B (n_17283), .Y (n_17623));
AND2X1 g67448(.A (n_17621), .B (n_11989), .Y (n_17622));
AND2X1 g67466(.A (n_17619), .B (n_7309), .Y (n_17620));
OR2X1 g67486(.A (n_19781), .B (n_19364), .Y (n_17618));
NAND2X1 g67493(.A (n_19690), .B (n_14442), .Y (n_17617));
INVX1 g67524(.A (n_27684), .Y (n_17616));
AND2X1 g65395(.A (n_4640), .B (n_16906), .Y (n_17611));
NOR2X1 g67562(.A (n_12748), .B (n_26704), .Y (n_17610));
OR2X1 g67582(.A (n_11893), .B (n_12298), .Y (n_17609));
OR2X1 g67593(.A (n_14284), .B (n_14589), .Y (n_17608));
NAND2X1 g67594(.A (n_13819), .B (n_19857), .Y (n_17607));
INVX1 g67659(.A (n_17605), .Y (n_17606));
NAND2X1 g67738(.A (n_17563), .B (n_6493), .Y (n_17604));
NOR2X1 g67782(.A (n_8921), .B (n_10292), .Y (n_28838));
OR2X1 g67801(.A (n_11923), .B (n_11277), .Y (n_17602));
NAND2X1 g67803(.A (n_12191), .B (n_11277), .Y (n_17601));
NAND2X1 g67833(.A (n_7548), .B (n_13886), .Y (n_17600));
INVX1 g67842(.A (n_17598), .Y (n_17599));
AND2X1 g67863(.A (n_9182), .B (n_17596), .Y (n_17597));
NOR2X1 g67866(.A (n_10297), .B (n_10616), .Y (n_17595));
NAND2X1 g67991(.A (n_11975), .B (n_29102), .Y (n_17594));
NOR2X1 g68010(.A (n_18904), .B (n_28645), .Y (n_17593));
NOR2X1 g68061(.A (n_12881), .B (n_15811), .Y (n_17592));
NAND2X1 g68090(.A (n_11843), .B (n_17590), .Y (n_17591));
NAND2X1 g68121(.A (n_17588), .B (n_13837), .Y (n_17589));
NOR2X1 g68132(.A (n_5329), .B (n_13884), .Y (n_17587));
NOR2X1 g68189(.A (n_9094), .B (n_10600), .Y (n_17586));
NAND2X1 g68218(.A (n_9817), .B (n_27151), .Y (n_17585));
AOI21X1 g61972(.A0 (n_11656), .A1 (n_15039), .B0 (n_13663), .Y(n_17584));
NAND2X1 g68301(.A (n_5414), .B (n_8009), .Y (n_17582));
INVX1 g68348(.A (n_17580), .Y (n_25725));
NAND3X1 g62004(.A (n_14947), .B (n_11617), .C (n_11512), .Y(n_17579));
NAND2X1 g62030(.A (n_13714), .B (n_12788), .Y (n_17578));
NOR2X1 g68514(.A (n_8559), .B (n_13778), .Y (n_17577));
INVX1 g68540(.A (n_15888), .Y (n_17576));
AOI21X1 g68553(.A0 (n_4370), .A1 (n_15799), .B0 (n_5329), .Y(n_17575));
AOI21X1 g68555(.A0 (n_5261), .A1 (n_11728), .B0 (n_11576), .Y(n_17573));
OAI21X1 g62054(.A0 (n_11499), .A1 (n_16472), .B0 (n_17571), .Y(n_17572));
NAND2X1 g68568(.A (n_13734), .B (n_28632), .Y (n_29418));
NAND2X1 g68571(.A (n_13736), .B (n_17411), .Y (n_17569));
OAI21X1 g62070(.A0 (n_11505), .A1 (n_9017), .B0 (n_17567), .Y(n_17568));
OAI21X1 g62075(.A0 (n_13361), .A1 (n_16375), .B0 (n_18168), .Y(n_25550));
NAND3X1 g65360(.A (n_11470), .B (n_10286), .C (n_16366), .Y(n_17565));
NAND2X1 g68634(.A (n_10516), .B (n_17563), .Y (n_17564));
OAI21X1 g62086(.A0 (n_11411), .A1 (n_8464), .B0 (n_15776), .Y(n_17562));
NAND2X1 g68638(.A (n_13931), .B (n_7796), .Y (n_17561));
NAND2X1 g68640(.A (n_10407), .B (n_13749), .Y (n_17560));
NAND2X1 g68646(.A (n_13920), .B (n_26842), .Y (n_17559));
AOI21X1 g68693(.A0 (n_9704), .A1 (n_29139), .B0 (n_11924), .Y(n_17558));
NAND2X1 g68698(.A (n_6437), .B (n_11989), .Y (n_17557));
NAND2X1 g68706(.A (n_13828), .B (n_13875), .Y (n_17556));
AOI21X1 g68711(.A0 (n_9712), .A1 (n_9668), .B0 (n_12494), .Y(n_17555));
OAI21X1 g62122(.A0 (n_13168), .A1 (n_13602), .B0 (n_27099), .Y(n_17554));
NAND3X1 g65393(.A (n_14542), .B (n_5169), .C (n_13946), .Y (n_17552));
OAI21X1 g62129(.A0 (n_13175), .A1 (n_11015), .B0 (n_16754), .Y(n_17551));
OAI21X1 g62130(.A0 (n_13169), .A1 (n_15395), .B0 (n_15986), .Y(n_17549));
NAND2X1 g68746(.A (n_13873), .B (n_8421), .Y (n_17548));
OR2X1 g68755(.A (n_6565), .B (n_11900), .Y (n_17547));
OR2X1 g68760(.A (n_7929), .B (n_28816), .Y (n_17546));
AOI21X1 g62137(.A0 (n_11561), .A1 (n_14155), .B0 (n_8700), .Y(n_17545));
AOI21X1 g62138(.A0 (n_11568), .A1 (n_15712), .B0 (n_9366), .Y(n_17544));
NAND2X1 g68766(.A (n_10077), .B (n_13849), .Y (n_17543));
OR2X1 g68781(.A (n_7923), .B (n_11795), .Y (n_17542));
NAND2X1 g68784(.A (n_10085), .B (n_17540), .Y (n_17541));
XOR2X1 g68810(.A (n_974), .B (n_11636), .Y (n_17539));
XOR2X1 g68821(.A (n_1224), .B (n_11623), .Y (n_17538));
AOI21X1 g62198(.A0 (n_13232), .A1 (n_20153), .B0 (n_10756), .Y(n_17537));
AOI21X1 g62204(.A0 (n_13146), .A1 (w3[25] ), .B0 (n_10754), .Y(n_17535));
AOI21X1 g62218(.A0 (n_11502), .A1 (n_7832), .B0 (n_11035), .Y(n_17533));
NAND4X1 g62238(.A (n_25695), .B (n_9605), .C (n_17531), .D (n_8772),.Y (n_17532));
OAI21X1 g62245(.A0 (n_11535), .A1 (n_11994), .B0 (n_18237), .Y(n_17530));
INVX1 g69039(.A (n_18682), .Y (n_18627));
AND2X1 g62247(.A (n_13694), .B (n_17527), .Y (n_17528));
OAI21X1 g62251(.A0 (n_13283), .A1 (n_10604), .B0 (n_19408), .Y(n_17526));
OAI21X1 g62254(.A0 (n_11529), .A1 (n_10539), .B0 (n_9410), .Y(n_17525));
OAI21X1 g62260(.A0 (n_11445), .A1 (n_17522), .B0 (n_3264), .Y(n_17523));
NAND4X1 g62279(.A (n_9365), .B (n_6823), .C (n_11059), .D (n_4536),.Y (n_17521));
NOR3X1 g62280(.A (n_7554), .B (n_8107), .C (n_13123), .Y (n_17519));
OAI21X1 g62304(.A0 (n_11494), .A1 (n_10374), .B0 (n_12298), .Y(n_29310));
OAI21X1 g62332(.A0 (n_13358), .A1 (n_10444), .B0 (n_19398), .Y(n_17517));
OAI21X1 g62335(.A0 (n_13352), .A1 (n_8992), .B0 (n_15568), .Y(n_17516));
OAI21X1 g62346(.A0 (n_13335), .A1 (n_10498), .B0 (n_8708), .Y(n_17514));
OAI21X1 g62348(.A0 (n_13334), .A1 (n_10391), .B0 (n_19395), .Y(n_17512));
NAND2X1 g62354(.A (n_13727), .B (sa32[2] ), .Y (n_17511));
NAND4X1 g62357(.A (n_14523), .B (n_9644), .C (n_10881), .D (n_8715),.Y (n_17510));
NAND4X1 g62367(.A (n_25478), .B (n_9702), .C (n_17508), .D (n_8219),.Y (n_17509));
NAND3X1 g62370(.A (n_17217), .B (n_11361), .C (n_13312), .Y(n_17507));
NOR3X1 g62371(.A (n_27471), .B (n_8108), .C (n_13126), .Y (n_17506));
NOR3X1 g62373(.A (n_27409), .B (n_8008), .C (n_13125), .Y (n_17505));
NOR3X1 g62376(.A (n_7146), .B (n_6821), .C (n_13124), .Y (n_17504));
AOI22X1 g62422(.A0 (n_11540), .A1 (n_15894), .B0 (n_8813), .B1(n_6534), .Y (n_17503));
AOI22X1 g62430(.A0 (n_11471), .A1 (n_17500), .B0 (n_9126), .B1(n_9118), .Y (n_17501));
AOI22X1 g62433(.A0 (n_11525), .A1 (n_18320), .B0 (n_10460), .B1(n_14484), .Y (n_17499));
AOI22X1 g62439(.A0 (n_11518), .A1 (n_11354), .B0 (n_14757), .B1(n_12133), .Y (n_17498));
NAND2X1 g62441(.A (n_13900), .B (n_13772), .Y (n_25732));
AOI21X1 g62443(.A0 (n_11504), .A1 (n_16466), .B0 (n_13202), .Y(n_17496));
NAND2X1 g62448(.A (n_14833), .B (n_11663), .Y (n_17495));
NOR2X1 g62457(.A (n_13678), .B (n_14646), .Y (n_17494));
NOR2X1 g62461(.A (n_13677), .B (n_13054), .Y (n_17493));
OAI21X1 g62483(.A0 (n_13164), .A1 (n_17491), .B0 (n_3612), .Y(n_28582));
OAI21X1 g62484(.A0 (n_13149), .A1 (n_8163), .B0 (n_638), .Y(n_17489));
NAND2X1 g62488(.A (n_13798), .B (n_27100), .Y (n_17487));
OAI21X1 g62501(.A0 (n_9226), .A1 (n_13083), .B0 (n_13797), .Y(n_17486));
OAI21X1 g62509(.A0 (n_13141), .A1 (n_10129), .B0 (n_510), .Y(n_17485));
AOI21X1 g62512(.A0 (n_13223), .A1 (n_13466), .B0 (n_13555), .Y(n_17484));
NOR2X1 g62513(.A (n_13699), .B (n_16469), .Y (n_17483));
NAND3X1 g62514(.A (n_14860), .B (n_11604), .C (n_17687), .Y(n_17482));
NOR2X1 g62517(.A (n_13705), .B (n_16441), .Y (n_17481));
AOI21X1 g62532(.A0 (n_13227), .A1 (n_12827), .B0 (n_13548), .Y(n_17480));
NAND2X1 g62545(.A (n_13791), .B (n_18456), .Y (n_17479));
OAI21X1 g62553(.A0 (n_13187), .A1 (n_17477), .B0 (n_290), .Y(n_25551));
OAI21X1 g62556(.A0 (n_13185), .A1 (n_10005), .B0 (n_17474), .Y(n_25618));
OAI21X1 g62564(.A0 (n_13174), .A1 (n_17472), .B0 (n_26270), .Y(n_17473));
DFFX1 u0_r0_out_reg[29] (.CK (clk), .D (n_13729), .Q (u0_rcon_1058),.QN ());
INVX1 g65374(.A (n_15818), .Y (n_17470));
OAI21X1 g62597(.A0 (n_13160), .A1 (n_17467), .B0 (n_20477), .Y(n_25488));
OAI21X1 g62608(.A0 (n_13136), .A1 (n_17465), .B0 (n_1756), .Y(n_28321));
NAND3X1 g62616(.A (n_14877), .B (n_11599), .C (n_17685), .Y(n_17462));
AOI21X1 g62617(.A0 (n_13263), .A1 (n_17703), .B0 (n_14597), .Y(n_17461));
NOR2X1 g62628(.A (n_13306), .B (n_13723), .Y (n_17458));
NAND4X1 g62651(.A (n_12217), .B (n_11072), .C (n_17456), .D(n_17455), .Y (n_17457));
NAND4X1 g62659(.A (n_6358), .B (n_15493), .C (n_6637), .D (n_11397),.Y (n_17454));
AOI21X1 g62663(.A0 (n_13133), .A1 (w3[1] ), .B0 (n_13551), .Y(n_17453));
NAND4X1 g62664(.A (n_11744), .B (n_15487), .C (n_4209), .D (n_11324),.Y (n_17451));
NAND4X1 g62667(.A (n_14738), .B (n_15468), .C (n_13219), .D(n_16954), .Y (n_17450));
NAND4X1 g62669(.A (n_13774), .B (n_16970), .C (n_6551), .D (n_9462),.Y (n_17449));
NAND4X1 g62689(.A (n_5708), .B (n_5162), .C (n_11358), .D (n_6657),.Y (n_17448));
NAND4X1 g62691(.A (n_8181), .B (n_17446), .C (n_5317), .D (n_11288),.Y (n_17447));
AOI21X1 g62698(.A0 (n_13241), .A1 (n_17444), .B0 (n_11127), .Y(n_17445));
NAND4X1 g62714(.A (n_17124), .B (n_12425), .C (n_17123), .D(n_28840), .Y (n_17443));
AOI22X1 g62745(.A0 (n_13115), .A1 (n_19433), .B0 (n_9286), .B1(n_14142), .Y (n_17442));
OAI21X1 g62750(.A0 (n_13165), .A1 (n_1424), .B0 (n_11143), .Y(n_17439));
AOI21X1 g62751(.A0 (n_13233), .A1 (n_16052), .B0 (n_11574), .Y(n_17438));
AOI21X1 g62760(.A0 (n_13209), .A1 (n_9755), .B0 (n_13046), .Y(n_17437));
NAND4X1 g62764(.A (n_14737), .B (n_13239), .C (n_5645), .D (n_13688),.Y (n_17435));
AOI21X1 g62770(.A0 (n_13199), .A1 (n_16090), .B0 (n_9596), .Y(n_17431));
AOI21X1 g62773(.A0 (n_13180), .A1 (n_6406), .B0 (n_11572), .Y(n_17430));
NOR2X1 g62778(.A (n_11328), .B (n_13717), .Y (n_17429));
NAND4X1 g62799(.A (n_8282), .B (n_8588), .C (n_17425), .D (n_8276),.Y (n_17426));
AOI21X1 g62802(.A0 (n_13130), .A1 (n_17423), .B0 (n_13762), .Y(n_17424));
AOI21X1 g62803(.A0 (n_13230), .A1 (w3[9] ), .B0 (n_13822), .Y(n_17422));
INVX1 g62811(.A (n_15788), .Y (n_17421));
OR2X1 g62819(.A (n_14781), .B (n_124), .Y (n_17419));
INVX1 g62831(.A (n_15784), .Y (n_17418));
AOI21X1 g62842(.A0 (n_12426), .A1 (n_17416), .B0 (n_2681), .Y(n_17417));
OAI21X1 g62845(.A0 (n_12432), .A1 (n_10215), .B0 (n_17414), .Y(n_17415));
OAI21X1 g62849(.A0 (n_12396), .A1 (n_17412), .B0 (n_17411), .Y(n_17413));
OAI21X1 g62856(.A0 (n_12356), .A1 (n_17409), .B0 (n_27688), .Y(n_17410));
OAI21X1 g62857(.A0 (n_12310), .A1 (n_28832), .B0 (n_17260), .Y(n_17408));
OAI21X1 g62858(.A0 (n_12307), .A1 (n_17405), .B0 (n_18266), .Y(n_17406));
AOI21X1 g62865(.A0 (n_8347), .A1 (n_15302), .B0 (n_21174), .Y(n_17404));
OR2X1 g62866(.A (n_14879), .B (n_16480), .Y (n_17402));
AOI21X1 g62867(.A0 (n_15267), .A1 (n_28584), .B0 (n_26931), .Y(n_17400));
OAI21X1 g62884(.A0 (n_12603), .A1 (n_8442), .B0 (n_9819), .Y(n_17399));
OAI21X1 g62908(.A0 (n_12346), .A1 (n_7077), .B0 (n_16198), .Y(n_17397));
AOI21X1 g62910(.A0 (n_11689), .A1 (n_15342), .B0 (n_27045), .Y(n_17396));
AOI21X1 g62921(.A0 (n_12447), .A1 (n_11470), .B0 (n_17411), .Y(n_17395));
OAI21X1 g62926(.A0 (n_12857), .A1 (n_12200), .B0 (n_9410), .Y(n_17393));
OAI21X1 g62927(.A0 (n_12670), .A1 (n_12182), .B0 (n_15568), .Y(n_17392));
OAI21X1 g62930(.A0 (n_25827), .A1 (n_25828), .B0 (n_1424), .Y(n_17390));
OR2X1 g72069(.A (n_13657), .B (n_25926), .Y (n_17389));
OAI21X1 g62936(.A0 (n_12702), .A1 (n_10514), .B0 (n_15894), .Y(n_17388));
OAI21X1 g62939(.A0 (n_12504), .A1 (n_7454), .B0 (n_263), .Y(n_17387));
OAI21X1 g62950(.A0 (n_13947), .A1 (n_15415), .B0 (n_688), .Y(n_17386));
NAND2X1 g62953(.A (n_13652), .B (n_9085), .Y (n_17385));
NAND2X1 g62954(.A (n_13651), .B (n_12306), .Y (n_17384));
NAND2X1 g62955(.A (n_13649), .B (n_17689), .Y (n_17383));
AOI21X1 g62959(.A0 (n_12798), .A1 (n_16480), .B0 (n_15276), .Y(n_17382));
NOR2X1 g62960(.A (n_14867), .B (n_18347), .Y (n_17381));
NAND2X1 g62961(.A (n_13642), .B (n_12309), .Y (n_17380));
NAND2X1 g62975(.A (n_13461), .B (n_1295), .Y (n_17376));
XOR2X1 g60241(.A (u0_rcon_1059), .B (n_1226), .Y (n_17375));
NAND2X1 g62977(.A (n_13632), .B (n_18749), .Y (n_17374));
NAND2X1 g62978(.A (n_13638), .B (n_12628), .Y (n_17373));
XOR2X1 g60242(.A (u0_rcon_1060), .B (n_1104), .Y (n_17372));
NAND3X1 g62982(.A (n_6733), .B (n_12994), .C (n_6407), .Y (n_17369));
NAND2X1 g62990(.A (n_13637), .B (n_14330), .Y (n_17367));
NOR2X1 g62991(.A (n_28311), .B (n_28310), .Y (n_17366));
AOI21X1 g62999(.A0 (n_16634), .A1 (n_7650), .B0 (n_29102), .Y(n_17365));
NAND2X1 g63000(.A (n_14808), .B (n_10079), .Y (n_17364));
NAND3X1 g63007(.A (n_27435), .B (n_12909), .C (n_6669), .Y (n_17363));
NAND2X1 g63011(.A (n_13633), .B (n_14286), .Y (n_17362));
OAI21X1 g63012(.A0 (n_13932), .A1 (n_13585), .B0 (n_1310), .Y(n_17361));
NAND2X1 g63014(.A (n_13630), .B (n_17681), .Y (n_17360));
OAI21X1 g63016(.A0 (n_13936), .A1 (n_27505), .B0 (n_3886), .Y(n_17359));
NAND3X1 g63017(.A (n_6529), .B (n_13030), .C (n_9638), .Y (n_17358));
NAND3X1 g63021(.A (n_17356), .B (n_5182), .C (n_15319), .Y (n_17357));
OAI21X1 g63022(.A0 (n_12800), .A1 (n_8868), .B0 (n_20157), .Y(n_25579));
OAI21X1 g63028(.A0 (n_12213), .A1 (n_14082), .B0 (n_15894), .Y(n_17354));
AND2X1 g63033(.A (n_13525), .B (n_11312), .Y (n_17353));
NAND2X1 g63043(.A (n_14967), .B (n_4898), .Y (n_17351));
OAI21X1 g63044(.A0 (n_9329), .A1 (n_16089), .B0 (n_28037), .Y(n_17350));
OAI21X1 g63045(.A0 (n_12372), .A1 (n_8088), .B0 (n_15968), .Y(n_17349));
OAI21X1 g63046(.A0 (n_9300), .A1 (n_16051), .B0 (n_11052), .Y(n_17348));
NAND2X1 g63050(.A (n_14903), .B (n_13247), .Y (n_17347));
NOR2X1 g63052(.A (n_13570), .B (n_25894), .Y (n_17346));
AOI21X1 g65373(.A0 (n_13880), .A1 (n_12778), .B0 (n_15712), .Y(n_17345));
NAND2X1 g63057(.A (n_14892), .B (n_19395), .Y (n_17344));
NAND2X1 g63059(.A (n_13562), .B (n_20116), .Y (n_17343));
OAI21X1 g63060(.A0 (n_12263), .A1 (n_28618), .B0 (n_20767), .Y(n_17342));
NAND2X1 g63061(.A (n_14116), .B (n_19651), .Y (n_17341));
OAI21X1 g63068(.A0 (n_12120), .A1 (n_10777), .B0 (n_16434), .Y(n_17340));
NAND2X1 g63071(.A (n_12851), .B (n_15362), .Y (n_17339));
OAI21X1 g63081(.A0 (n_9205), .A1 (n_10204), .B0 (n_663), .Y(n_17335));
NOR2X1 g63083(.A (n_14882), .B (n_9819), .Y (n_17333));
NAND2X1 g63086(.A (n_17331), .B (n_10322), .Y (n_17332));
NAND2X1 g63092(.A (n_17329), .B (n_17328), .Y (n_17330));
NOR2X1 g63093(.A (n_13584), .B (n_16985), .Y (n_17327));
NAND2X1 g63095(.A (n_13647), .B (n_17325), .Y (n_17326));
OAI21X1 g63100(.A0 (n_12119), .A1 (n_14067), .B0 (n_19791), .Y(n_17324));
NAND2X1 g63101(.A (n_11001), .B (n_15283), .Y (n_17323));
NAND3X1 g63102(.A (n_17321), .B (n_12126), .C (n_18114), .Y(n_17322));
NAND3X1 g63104(.A (n_11104), .B (n_13065), .C (n_11620), .Y(n_17320));
NOR2X1 g63112(.A (n_11098), .B (n_13514), .Y (n_17319));
NAND2X1 g63115(.A (n_14516), .B (n_17317), .Y (n_17318));
NAND3X1 g63116(.A (n_17014), .B (n_11777), .C (n_17315), .Y(n_17316));
NAND2X1 g63117(.A (n_14759), .B (n_19314), .Y (n_17314));
NAND3X1 g63119(.A (n_10382), .B (n_16568), .C (n_26042), .Y(n_17313));
NOR2X1 g63121(.A (n_13507), .B (n_26867), .Y (n_17312));
NAND3X1 g63122(.A (n_17011), .B (n_9790), .C (n_17310), .Y (n_17311));
AOI21X1 g63126(.A0 (n_12753), .A1 (n_16466), .B0 (n_17308), .Y(n_17309));
NAND2X1 g63132(.A (n_16992), .B (n_4593), .Y (n_17307));
OAI21X1 g63133(.A0 (n_6692), .A1 (n_12773), .B0 (n_12827), .Y(n_17306));
NAND2X1 g63140(.A (n_15269), .B (n_14677), .Y (n_17305));
NAND3X1 g63145(.A (n_17303), .B (n_12124), .C (n_17302), .Y(n_17304));
NAND2X1 g63146(.A (n_17153), .B (n_19314), .Y (n_17301));
NAND2X1 g63147(.A (n_14785), .B (n_1310), .Y (n_25803));
AOI21X1 g63154(.A0 (n_11957), .A1 (n_16519), .B0 (n_15708), .Y(n_17299));
NAND3X1 g63155(.A (n_14880), .B (n_17297), .C (n_16559), .Y(n_17298));
NAND2X1 g63158(.A (n_17295), .B (n_5941), .Y (n_17296));
NAND3X1 g63159(.A (n_17293), .B (n_17292), .C (n_12082), .Y(n_17294));
NAND3X1 g63162(.A (n_19019), .B (n_15328), .C (n_6723), .Y (n_17291));
NAND3X1 g63163(.A (n_14436), .B (n_7115), .C (n_15358), .Y (n_17290));
OAI21X1 g63174(.A0 (n_13034), .A1 (n_17288), .B0 (n_18792), .Y(n_17289));
AND2X1 g63175(.A (n_14848), .B (n_17286), .Y (n_17287));
INVX1 g63177(.A (n_15673), .Y (n_17285));
OAI21X1 g63181(.A0 (n_12847), .A1 (n_6023), .B0 (n_15674), .Y(n_17284));
INVX2 g72983(.A (n_13745), .Y (n_17283));
NAND3X1 g63187(.A (sa20[1] ), .B (n_12265), .C (n_11261), .Y(n_17281));
AOI21X1 g63195(.A0 (n_12633), .A1 (n_4582), .B0 (n_15390), .Y(n_17279));
AOI21X1 g63196(.A0 (n_12819), .A1 (n_11567), .B0 (n_15712), .Y(n_29432));
NAND2X1 g63200(.A (n_14849), .B (n_1626), .Y (n_17277));
NAND3X1 g63202(.A (n_17274), .B (n_12122), .C (n_16501), .Y(n_17275));
OR2X1 g63208(.A (n_7666), .B (n_17269), .Y (n_17272));
NAND2X1 g63209(.A (n_15288), .B (n_14603), .Y (n_17271));
OR2X1 g63211(.A (n_9233), .B (n_17269), .Y (n_17270));
INVX1 g63213(.A (n_15661), .Y (n_17268));
AND2X1 g63217(.A (n_17266), .B (n_17265), .Y (n_29305));
NAND3X1 g63218(.A (n_12923), .B (n_10840), .C (n_12261), .Y(n_29180));
NAND2X1 g63219(.A (n_14776), .B (n_17262), .Y (n_17263));
AOI21X1 g63227(.A0 (n_12530), .A1 (n_14978), .B0 (n_17260), .Y(n_17261));
NAND2X1 g63231(.A (n_13656), .B (n_14478), .Y (n_17259));
NAND3X1 g63232(.A (n_15222), .B (n_12353), .C (n_12205), .Y(n_17258));
OAI21X1 g63233(.A0 (n_12237), .A1 (n_7075), .B0 (sa10[1] ), .Y(n_17257));
NOR2X1 g63243(.A (n_12725), .B (n_16997), .Y (n_17255));
OAI21X1 g63244(.A0 (n_9201), .A1 (n_17253), .B0 (n_3538), .Y(n_17254));
NAND3X1 g63245(.A (n_17250), .B (n_9164), .C (n_16503), .Y (n_17251));
OAI21X1 g63246(.A0 (n_12118), .A1 (n_10775), .B0 (n_19364), .Y(n_17249));
OAI21X1 g63248(.A0 (n_12235), .A1 (n_18278), .B0 (n_17246), .Y(n_17247));
AOI21X1 g63252(.A0 (n_10425), .A1 (n_15345), .B0 (n_17414), .Y(n_17245));
NAND2X1 g63255(.A (n_14388), .B (n_15130), .Y (n_17244));
AOI21X1 g63259(.A0 (n_12026), .A1 (n_28880), .B0 (n_26276), .Y(n_17243));
NAND3X1 g63261(.A (n_16351), .B (n_27472), .C (n_17240), .Y(n_17242));
NOR2X1 g63262(.A (n_16034), .B (n_15118), .Y (n_17239));
NOR2X1 g63265(.A (n_11487), .B (n_25945), .Y (n_17238));
NAND3X1 g63266(.A (n_17236), .B (n_9827), .C (n_17235), .Y (n_17237));
NAND3X1 g63267(.A (n_10251), .B (n_16593), .C (n_11122), .Y(n_17234));
NAND3X1 g63270(.A (n_10398), .B (n_18051), .C (n_17232), .Y(n_17233));
NOR2X1 g63271(.A (n_14835), .B (n_9106), .Y (n_17231));
NAND3X1 g63273(.A (n_14042), .B (n_13366), .C (n_3829), .Y (n_17230));
NAND3X1 g63274(.A (n_16999), .B (n_11875), .C (n_17228), .Y(n_17229));
NOR2X1 g63276(.A (n_14986), .B (n_15324), .Y (n_17227));
NAND2X1 g63283(.A (n_14827), .B (n_13725), .Y (n_17226));
NAND2X1 g63294(.A (n_15127), .B (n_14655), .Y (n_17224));
OR2X1 g63297(.A (n_13365), .B (n_17222), .Y (n_17223));
AND2X1 g63300(.A (n_15612), .B (n_17455), .Y (n_17221));
NAND2X1 g63304(.A (n_15063), .B (n_16973), .Y (n_17220));
OAI21X1 g63305(.A0 (n_10372), .A1 (n_14649), .B0 (n_3910), .Y(n_17219));
NAND3X1 g63306(.A (n_8691), .B (n_7404), .C (n_17217), .Y (n_17218));
AND2X1 g63308(.A (n_15054), .B (n_2606), .Y (n_17216));
INVX1 g63310(.A (n_15631), .Y (n_17215));
AOI21X1 g63313(.A0 (n_12001), .A1 (n_15281), .B0 (n_15574), .Y(n_17214));
NAND2X1 g63315(.A (n_11600), .B (n_11949), .Y (n_17213));
NOR2X1 g63325(.A (n_14812), .B (n_17211), .Y (n_17212));
NAND3X1 g63329(.A (n_10287), .B (n_15159), .C (n_14384), .Y(n_17210));
NAND3X1 g63331(.A (n_14251), .B (n_7816), .C (n_15170), .Y (n_17209));
INVX1 g63342(.A (n_15620), .Y (n_17208));
AOI21X1 g63349(.A0 (n_12055), .A1 (n_15121), .B0 (n_15039), .Y(n_17207));
AOI21X1 g63353(.A0 (n_12450), .A1 (n_11456), .B0 (n_17912), .Y(n_17205));
OAI21X1 g63357(.A0 (n_10629), .A1 (n_12937), .B0 (n_29106), .Y(n_17203));
NAND3X1 g63358(.A (n_10964), .B (n_15404), .C (n_15998), .Y(n_17201));
AND2X1 g63364(.A (n_14133), .B (n_15630), .Y (n_25777));
INVX1 g63369(.A (n_15609), .Y (n_17199));
NAND3X1 g63372(.A (n_7726), .B (n_10285), .C (n_17197), .Y (n_17198));
AOI21X1 g63375(.A0 (n_12428), .A1 (n_11447), .B0 (n_26670), .Y(n_17196));
NAND2X1 g63381(.A (n_14955), .B (sa11[1] ), .Y (n_17195));
AOI21X1 g63385(.A0 (n_12406), .A1 (n_9559), .B0 (n_15039), .Y(n_17193));
AOI21X1 g63387(.A0 (n_12418), .A1 (n_13469), .B0 (n_11576), .Y(n_17192));
NAND3X1 g63388(.A (n_21487), .B (n_13359), .C (n_19395), .Y(n_17191));
AOI21X1 g63396(.A0 (n_12708), .A1 (n_9561), .B0 (n_15986), .Y(n_17188));
NAND3X1 g63398(.A (n_10726), .B (n_14337), .C (n_26796), .Y(n_17187));
OR2X1 g63401(.A (n_7644), .B (n_17151), .Y (n_17186));
AOI21X1 g63404(.A0 (n_12270), .A1 (n_15135), .B0 (n_9106), .Y(n_17185));
NAND2X1 g63408(.A (n_14794), .B (n_15100), .Y (n_17184));
AND2X1 g63409(.A (n_14966), .B (n_3967), .Y (n_17183));
NAND2X1 g63410(.A (n_12423), .B (n_16610), .Y (n_17182));
NAND2X1 g63415(.A (n_14793), .B (n_17180), .Y (n_17181));
AOI21X1 g63419(.A0 (n_12592), .A1 (n_16683), .B0 (n_28692), .Y(n_17179));
NAND2X1 g63420(.A (n_14792), .B (n_17177), .Y (n_17178));
NAND3X1 g63422(.A (n_14005), .B (n_26952), .C (n_12587), .Y(n_17176));
INVX1 g63425(.A (n_15602), .Y (n_17175));
NOR2X1 g63432(.A (n_14932), .B (n_7551), .Y (n_17174));
NOR2X1 g63433(.A (n_15423), .B (n_16995), .Y (n_17173));
AOI21X1 g63438(.A0 (n_12363), .A1 (n_13370), .B0 (n_27688), .Y(n_17172));
OR2X1 g63439(.A (n_18365), .B (n_3264), .Y (n_17170));
NAND2X1 g63447(.A (n_17189), .B (n_9143), .Y (n_17169));
OAI21X1 g63448(.A0 (n_12210), .A1 (n_8514), .B0 (sa13[1] ), .Y(n_17167));
NOR2X1 g63452(.A (n_14784), .B (n_9982), .Y (n_17165));
NOR2X1 g63460(.A (n_14861), .B (n_15039), .Y (n_17164));
NAND2X1 g63463(.A (n_14931), .B (n_804), .Y (n_28316));
AND2X1 g63464(.A (n_17161), .B (n_11517), .Y (n_17162));
NAND3X1 g63469(.A (n_18268), .B (n_16540), .C (n_16539), .Y(n_17159));
NAND2X1 g63476(.A (n_17157), .B (n_11287), .Y (n_17158));
NAND2X1 g63478(.A (n_14915), .B (n_7649), .Y (n_17156));
INVX1 g63480(.A (n_15593), .Y (n_17155));
AND2X1 g63482(.A (n_17153), .B (n_18046), .Y (n_17154));
OR2X1 g63484(.A (n_9213), .B (n_17151), .Y (n_17152));
OAI21X1 g63485(.A0 (n_12215), .A1 (n_9872), .B0 (sa12[1] ), .Y(n_17150));
INVX1 g63488(.A (n_15592), .Y (n_17146));
NOR2X1 g63491(.A (n_14774), .B (n_11576), .Y (n_17145));
NOR2X1 g63496(.A (n_11159), .B (n_14898), .Y (n_17143));
AOI22X1 g63499(.A0 (n_12877), .A1 (n_5329), .B0 (n_15919), .B1(n_8425), .Y (n_17142));
NAND3X1 g63500(.A (n_14736), .B (n_17140), .C (n_17139), .Y(n_17141));
AOI22X1 g63505(.A0 (n_12794), .A1 (n_27133), .B0 (n_8317), .B1(n_8491), .Y (n_17138));
NAND3X1 g63509(.A (n_14934), .B (n_12620), .C (n_11011), .Y(n_17137));
NAND3X1 g63511(.A (n_14452), .B (n_14899), .C (n_15322), .Y(n_17136));
NAND3X1 g63517(.A (n_17134), .B (n_12538), .C (n_10967), .Y(n_25785));
NAND3X1 g63523(.A (n_28029), .B (n_12483), .C (n_9313), .Y (n_17133));
NAND3X1 g63527(.A (n_17130), .B (n_9842), .C (n_17129), .Y (n_17131));
NAND3X1 g63529(.A (n_17127), .B (n_12443), .C (n_12441), .Y(n_17128));
NAND4X1 g63531(.A (n_17125), .B (n_17124), .C (n_15085), .D(n_17123), .Y (n_17126));
NAND3X1 g63534(.A (n_14185), .B (n_16614), .C (n_17121), .Y(n_17122));
NAND3X1 g63536(.A (n_14179), .B (n_14969), .C (n_16588), .Y(n_17119));
AOI21X1 g63539(.A0 (n_19226), .A1 (n_7568), .B0 (n_14851), .Y(n_17118));
NAND3X1 g63541(.A (n_17115), .B (n_12281), .C (n_9318), .Y (n_17116));
NAND3X1 g63542(.A (n_10992), .B (n_5935), .C (n_17113), .Y (n_17114));
AOI22X1 g63543(.A0 (n_12782), .A1 (n_27604), .B0 (n_6422), .B1(n_10163), .Y (n_17112));
NAND2X1 g65354(.A (n_12176), .B (n_16683), .Y (n_17111));
INVX1 g63548(.A (n_15576), .Y (n_17110));
NAND3X1 g63553(.A (n_6619), .B (n_13027), .C (n_9793), .Y (n_17108));
OR2X1 g63555(.A (n_13412), .B (n_15610), .Y (n_17107));
NAND3X1 g63556(.A (n_6235), .B (n_12965), .C (n_9871), .Y (n_17106));
AOI21X1 g63557(.A0 (n_12167), .A1 (n_9115), .B0 (n_17104), .Y(n_17105));
INVX1 g63558(.A (n_15570), .Y (n_17103));
OAI21X1 g63560(.A0 (n_12173), .A1 (n_9024), .B0 (n_29018), .Y(n_17102));
INVX1 g63561(.A (n_15569), .Y (n_17101));
INVX1 g63563(.A (n_15567), .Y (n_17100));
INVX1 g63569(.A (n_15564), .Y (n_17099));
OR2X1 g63572(.A (n_14911), .B (n_27604), .Y (n_17098));
NOR2X1 g63573(.A (n_10861), .B (n_17096), .Y (n_17097));
NAND2X1 g63574(.A (n_13574), .B (n_10857), .Y (n_17095));
NAND2X1 g63576(.A (n_9991), .B (n_13427), .Y (n_17094));
NAND2X1 g63579(.A (n_13565), .B (n_17064), .Y (n_17093));
NAND2X1 g63583(.A (n_11800), .B (n_13560), .Y (n_17092));
AOI21X1 g63586(.A0 (n_9366), .A1 (n_17571), .B0 (n_14490), .Y(n_17091));
NAND2X1 g63589(.A (n_13557), .B (n_17089), .Y (n_17090));
AOI21X1 g63595(.A0 (n_9346), .A1 (n_14624), .B0 (n_14151), .Y(n_17088));
NAND4X1 g63613(.A (n_11204), .B (n_8902), .C (n_10710), .D (n_10912),.Y (n_17086));
NAND2X1 g63622(.A (n_15001), .B (n_10932), .Y (n_17085));
AOI21X1 g63625(.A0 (n_17302), .A1 (n_17083), .B0 (n_20010), .Y(n_17084));
OAI21X1 g63627(.A0 (n_12374), .A1 (n_10513), .B0 (n_14113), .Y(n_17082));
AOI21X1 g63628(.A0 (n_4191), .A1 (n_9755), .B0 (n_13488), .Y(n_17081));
NAND2X1 g63631(.A (n_14979), .B (n_12986), .Y (n_17080));
NAND2X1 g63635(.A (n_14952), .B (n_12298), .Y (n_17078));
AOI21X1 g63642(.A0 (n_5444), .A1 (n_19110), .B0 (n_13473), .Y(n_17077));
NAND2X1 g63648(.A (n_14946), .B (n_17411), .Y (n_17076));
AND2X1 g63653(.A (n_13471), .B (n_15574), .Y (n_17074));
AOI21X1 g63660(.A0 (n_12513), .A1 (n_1626), .B0 (n_5973), .Y(n_17073));
NAND3X1 g63663(.A (n_16492), .B (n_17071), .C (n_16557), .Y(n_17072));
AOI21X1 g63665(.A0 (n_12255), .A1 (n_15432), .B0 (n_17069), .Y(n_17070));
AOI21X1 g63666(.A0 (n_16988), .A1 (n_6713), .B0 (n_13434), .Y(n_17068));
NAND2X1 g63669(.A (n_13513), .B (n_1424), .Y (n_17067));
NAND4X1 g63672(.A (n_17064), .B (n_5607), .C (n_11774), .D (n_7472),.Y (n_17065));
AND2X1 g63673(.A (n_8529), .B (n_17062), .Y (n_17063));
NAND2X1 g63674(.A (n_14917), .B (n_10905), .Y (n_17061));
NAND3X1 g63679(.A (n_14397), .B (n_8942), .C (n_13013), .Y (n_17060));
NAND2X1 g63688(.A (n_13407), .B (n_17058), .Y (n_17059));
NAND2X1 g63690(.A (n_13403), .B (n_17035), .Y (n_17057));
AOI21X1 g63694(.A0 (n_9279), .A1 (n_26270), .B0 (n_14368), .Y(n_17054));
AND2X1 g63700(.A (n_13387), .B (n_9819), .Y (n_17053));
NAND2X1 g63701(.A (n_13384), .B (n_29014), .Y (n_28607));
NAND2X1 g63703(.A (n_13371), .B (n_17775), .Y (n_17050));
NAND3X1 g63706(.A (n_17048), .B (n_10202), .C (n_16532), .Y(n_17049));
NAND2X1 g63713(.A (n_11051), .B (n_17046), .Y (n_17047));
AOI21X1 g63715(.A0 (n_9198), .A1 (n_17129), .B0 (n_29062), .Y(n_17045));
NAND2X1 g63722(.A (n_15029), .B (n_19395), .Y (n_17043));
NAND3X1 g63740(.A (n_12399), .B (n_17041), .C (n_17040), .Y(n_17042));
NAND3X1 g63748(.A (n_16394), .B (n_15648), .C (n_15151), .Y(n_17039));
NAND4X1 g63755(.A (n_10876), .B (n_14152), .C (n_17037), .D(n_14393), .Y (n_17038));
NAND4X1 g63756(.A (n_17035), .B (n_6762), .C (n_11707), .D (n_8856),.Y (n_17036));
NAND3X1 g63760(.A (n_12383), .B (n_17033), .C (n_16768), .Y(n_17034));
NAND3X1 g63768(.A (n_27744), .B (n_18275), .C (n_17031), .Y(n_17032));
NAND4X1 g63781(.A (n_15177), .B (n_16825), .C (n_28556), .D(n_14094), .Y (n_17030));
NAND2X1 g63782(.A (n_14941), .B (n_14589), .Y (n_17029));
AOI21X1 g63786(.A0 (n_15538), .A1 (n_13019), .B0 (n_1295), .Y(n_17028));
NAND2X1 g63787(.A (n_9883), .B (n_14937), .Y (n_17026));
AOI21X1 g63806(.A0 (n_16595), .A1 (n_17024), .B0 (n_17023), .Y(n_17025));
AOI21X1 g63809(.A0 (n_15195), .A1 (n_17021), .B0 (n_17020), .Y(n_17022));
AOI21X1 g63810(.A0 (n_11579), .A1 (n_17018), .B0 (n_17017), .Y(n_17019));
OR2X1 g63817(.A (n_13621), .B (n_13578), .Y (n_17016));
NAND4X1 g63820(.A (n_11380), .B (n_12414), .C (n_17014), .D (n_8188),.Y (n_17015));
NAND4X1 g63821(.A (n_28590), .B (n_17012), .C (n_17011), .D(n_28591), .Y (n_17013));
NAND4X1 g63826(.A (n_12987), .B (n_7608), .C (n_13955), .D (n_8302),.Y (n_17010));
NAND4X1 g63827(.A (n_11267), .B (n_8726), .C (n_28164), .D (n_10203),.Y (n_17009));
NAND4X1 g63828(.A (n_12953), .B (n_6911), .C (n_10361), .D (n_8235),.Y (n_17007));
NAND4X1 g63829(.A (n_12930), .B (n_13807), .C (n_17005), .D (n_9818),.Y (n_17006));
NAND2X1 g63831(.A (n_14957), .B (n_17003), .Y (n_17004));
NAND4X1 g63832(.A (n_11220), .B (n_7168), .C (n_15682), .D (n_9807),.Y (n_17002));
NAND4X1 g63835(.A (n_13039), .B (n_17000), .C (n_16999), .D(n_10165), .Y (n_17001));
OR2X1 g63842(.A (n_8980), .B (n_16997), .Y (n_16998));
AOI21X1 g63847(.A0 (n_6432), .A1 (n_19110), .B0 (n_16995), .Y(n_16996));
NOR2X1 g63849(.A (n_5736), .B (n_15262), .Y (n_16994));
NAND2X1 g63851(.A (n_3407), .B (n_16992), .Y (n_16993));
NAND3X1 g63852(.A (n_12550), .B (n_16412), .C (n_16990), .Y(n_16991));
AOI21X1 g63853(.A0 (n_5152), .A1 (n_16988), .B0 (n_15210), .Y(n_16989));
NAND3X1 g63854(.A (n_14207), .B (n_16737), .C (n_14309), .Y(n_16987));
OR2X1 g63864(.A (n_7412), .B (n_16985), .Y (n_16986));
AOI21X1 g63874(.A0 (n_12199), .A1 (n_196), .B0 (n_12795), .Y(n_16984));
NAND2X1 g63876(.A (n_13520), .B (n_18876), .Y (n_16982));
OAI21X1 g63878(.A0 (n_15700), .A1 (n_14866), .B0 (n_13617), .Y(n_16981));
AOI21X1 g63880(.A0 (n_12193), .A1 (n_933), .B0 (n_12502), .Y(n_16980));
AOI22X1 g63890(.A0 (n_12190), .A1 (n_16978), .B0 (n_5997), .B1(n_12134), .Y (n_16979));
AOI22X1 g63891(.A0 (n_12188), .A1 (n_1667), .B0 (n_7084), .B1(n_16976), .Y (n_16977));
NOR2X1 g63925(.A (n_14471), .B (n_13668), .Y (n_16972));
NOR2X1 g63929(.A (n_7098), .B (n_13428), .Y (n_16969));
NOR2X1 g63933(.A (n_10928), .B (n_13664), .Y (n_16968));
NOR2X1 g63936(.A (n_8584), .B (n_14953), .Y (n_16967));
NOR2X1 g63938(.A (n_8130), .B (n_14939), .Y (n_16966));
NAND3X1 g63942(.A (n_14547), .B (n_11539), .C (n_15942), .Y(n_16965));
NAND4X1 g63945(.A (n_10854), .B (n_16963), .C (n_9214), .D (n_13588),.Y (n_16964));
NAND4X1 g63951(.A (n_12786), .B (n_9323), .C (n_16550), .D (n_29208),.Y (n_16962));
NAND4X1 g63953(.A (n_16503), .B (n_16586), .C (n_16959), .D(n_18199), .Y (n_16960));
NAND4X1 g63957(.A (n_16501), .B (n_10231), .C (n_13487), .D(n_16956), .Y (n_16958));
NAND4X1 g63958(.A (n_14451), .B (n_9465), .C (n_16954), .D (n_12324),.Y (n_16955));
NAND4X1 g63967(.A (n_17821), .B (n_27141), .C (n_5731), .D (n_14951),.Y (n_16952));
NAND4X1 g63969(.A (n_15012), .B (n_8251), .C (n_15187), .D (n_13398),.Y (n_16951));
NAND3X1 g63970(.A (n_12411), .B (n_13322), .C (n_16678), .Y(n_16950));
NAND3X1 g63972(.A (n_14189), .B (n_11470), .C (n_8730), .Y (n_16949));
NAND3X1 g63973(.A (n_14129), .B (n_11524), .C (n_7354), .Y (n_16948));
NAND3X1 g63975(.A (n_14444), .B (n_12208), .C (n_26247), .Y(n_16947));
NAND3X1 g63982(.A (n_9581), .B (n_15425), .C (n_14510), .Y (n_16946));
AOI21X1 g63983(.A0 (n_12135), .A1 (n_13539), .B0 (n_16944), .Y(n_16945));
AOI21X1 g63989(.A0 (n_14546), .A1 (n_11261), .B0 (n_13419), .Y(n_16943));
NAND3X1 g63990(.A (n_13349), .B (n_16941), .C (n_12762), .Y(n_16942));
NOR2X1 g63996(.A (n_11246), .B (n_14995), .Y (n_16940));
XOR2X1 g76112(.A (n_16938), .B (n_14866), .Y (n_16939));
NAND2X1 g63998(.A (n_11198), .B (n_14977), .Y (n_16937));
OAI21X1 g64003(.A0 (n_12168), .A1 (n_28692), .B0 (n_13033), .Y(n_16936));
AOI21X1 g64009(.A0 (n_16934), .A1 (n_5215), .B0 (n_13527), .Y(n_16935));
AOI22X1 g64017(.A0 (n_12880), .A1 (n_20010), .B0 (n_16931), .B1(n_13083), .Y (n_16933));
AOI22X1 g64019(.A0 (n_14450), .A1 (n_267), .B0 (n_7245), .B1(n_15674), .Y (n_16929));
MX2X1 g64020(.A (n_16927), .B (n_7847), .S0 (n_14142), .Y (n_16928));
OAI21X1 g64057(.A0 (n_11709), .A1 (n_5318), .B0 (n_20325), .Y(n_16926));
INVX1 g64061(.A (n_15452), .Y (n_16925));
XOR2X1 g76274(.A (text_in_r[18] ), .B (n_19310), .Y (n_16924));
XOR2X1 g76278(.A (n_16921), .B (n_13083), .Y (n_16922));
NOR2X1 g64080(.A (n_14036), .B (n_15986), .Y (n_16920));
INVX1 g64085(.A (n_15442), .Y (n_16919));
AND2X1 g64106(.A (n_14165), .B (n_14624), .Y (n_16918));
AND2X1 g64108(.A (n_14525), .B (n_9410), .Y (n_16917));
AND2X1 g64109(.A (n_14143), .B (n_19475), .Y (n_16916));
NOR2X1 g64121(.A (n_16912), .B (n_17411), .Y (n_16913));
INVX1 g64122(.A (n_16910), .Y (n_16911));
INVX1 g64126(.A (n_16908), .Y (n_16909));
NOR2X1 g64146(.A (n_16906), .B (n_13083), .Y (n_16907));
INVX1 g64158(.A (n_16904), .Y (n_16905));
OR2X1 g64174(.A (n_16902), .B (n_15166), .Y (n_16903));
INVX1 g64184(.A (n_16897), .Y (n_16898));
AOI21X1 g64189(.A0 (n_16590), .A1 (n_16895), .B0 (n_14040), .Y(n_16896));
NOR2X1 g64199(.A (n_17929), .B (n_17414), .Y (n_18016));
OR2X1 g64208(.A (n_16893), .B (n_18679), .Y (n_16894));
INVX1 g64211(.A (n_16891), .Y (n_16892));
INVX1 g64221(.A (n_15387), .Y (n_18014));
OR2X1 g64224(.A (n_16889), .B (n_18369), .Y (n_16890));
AOI21X1 g64235(.A0 (n_9729), .A1 (n_16883), .B0 (sa00[1] ), .Y(n_16884));
NAND2X1 g64244(.A (n_13967), .B (n_62), .Y (n_16882));
INVX1 g64248(.A (n_15368), .Y (n_16880));
INVX1 g64250(.A (n_15367), .Y (n_16879));
INVX1 g64253(.A (n_15365), .Y (n_16878));
AOI21X1 g64257(.A0 (n_5219), .A1 (n_12973), .B0 (n_29048), .Y(n_16877));
NAND2X1 g64258(.A (n_13966), .B (n_1368), .Y (n_16875));
NAND2X1 g64259(.A (n_13958), .B (n_19995), .Y (n_16874));
NAND2X1 g64260(.A (n_13956), .B (n_20116), .Y (n_16873));
NAND2X1 g64274(.A (n_11191), .B (n_17411), .Y (n_16871));
NAND2X1 g64281(.A (n_16844), .B (n_13466), .Y (n_18010));
AND2X1 g64286(.A (n_16865), .B (n_16864), .Y (n_28280));
OR2X1 g64292(.A (n_13992), .B (n_14155), .Y (n_16863));
NAND2X1 g64294(.A (n_16861), .B (n_8062), .Y (n_16862));
OR2X1 g64298(.A (n_14012), .B (n_18679), .Y (n_16860));
OR2X1 g64303(.A (n_14011), .B (n_16835), .Y (n_16859));
NAND2X1 g64304(.A (n_16912), .B (n_16857), .Y (n_16858));
NAND2X1 g64311(.A (n_13148), .B (n_18268), .Y (n_16856));
AOI21X1 g64314(.A0 (n_11895), .A1 (n_8817), .B0 (n_18237), .Y(n_16855));
AND2X1 g64315(.A (n_16853), .B (n_11989), .Y (n_16854));
OR2X1 g64317(.A (n_13995), .B (n_17567), .Y (n_16852));
OAI21X1 g64331(.A0 (n_6353), .A1 (n_12895), .B0 (n_9527), .Y(n_16851));
INVX1 g64334(.A (n_15323), .Y (n_16850));
INVX1 g64339(.A (n_16848), .Y (n_16849));
NOR2X1 g64346(.A (n_16844), .B (n_13052), .Y (n_16845));
AOI21X1 g64352(.A0 (n_11685), .A1 (n_9690), .B0 (n_2290), .Y(n_16843));
NAND2X1 g64354(.A (n_14296), .B (n_4930), .Y (n_16842));
NAND2X1 g64372(.A (n_11388), .B (n_15894), .Y (n_16841));
NOR2X1 g64374(.A (n_11020), .B (n_16264), .Y (n_16840));
NAND2X1 g64383(.A (n_13989), .B (n_17089), .Y (n_16837));
NAND2X1 g64386(.A (n_11188), .B (n_16835), .Y (n_16836));
NAND2X1 g64394(.A (n_13077), .B (n_16480), .Y (n_16834));
INVX1 g64395(.A (n_16832), .Y (n_16833));
AND2X1 g64412(.A (n_16828), .B (n_16827), .Y (n_16829));
NAND4X1 g64413(.A (n_11951), .B (n_15600), .C (n_16825), .D (n_9082),.Y (n_16826));
NAND2X1 g64430(.A (n_28326), .B (n_12986), .Y (n_17995));
NAND2X1 g64435(.A (n_13986), .B (n_12986), .Y (n_16823));
NAND2X1 g64439(.A (n_11373), .B (n_19791), .Y (n_16822));
NOR2X1 g64446(.A (n_12725), .B (n_12637), .Y (n_16820));
AND2X1 g64447(.A (n_16817), .B (n_7603), .Y (n_16818));
OR2X1 g64451(.A (n_12865), .B (n_27099), .Y (n_16816));
NAND3X1 g64452(.A (n_10241), .B (n_5205), .C (n_16812), .Y (n_16813));
NAND2X1 g64453(.A (n_16108), .B (n_9819), .Y (n_19046));
NAND2X1 g64457(.A (n_11034), .B (n_16810), .Y (n_16811));
NOR2X1 g64466(.A (n_13988), .B (n_17912), .Y (n_16809));
NOR2X1 g65389(.A (n_12856), .B (n_12855), .Y (n_16808));
NOR2X1 g64472(.A (n_10896), .B (n_27604), .Y (n_16807));
NOR2X1 g64474(.A (n_15266), .B (n_14706), .Y (n_16806));
AND2X1 g64476(.A (n_13987), .B (n_13083), .Y (n_16805));
INVX1 g64477(.A (n_15258), .Y (n_25508));
NAND3X1 g64481(.A (n_16801), .B (n_11501), .C (n_9523), .Y (n_16802));
NAND2X1 g64493(.A (n_17832), .B (n_12299), .Y (n_16800));
INVX1 g64501(.A (n_15250), .Y (n_28886));
NAND2X1 g64503(.A (n_16797), .B (n_9783), .Y (n_16798));
OR2X1 g64528(.A (n_14492), .B (n_9410), .Y (n_16796));
AND2X1 g64552(.A (n_16793), .B (n_16912), .Y (n_16794));
NOR2X1 g64574(.A (n_8171), .B (n_11213), .Y (n_16792));
INVX1 g64575(.A (n_16790), .Y (n_16791));
NAND3X1 g64591(.A (n_16830), .B (n_14864), .C (n_28815), .Y(n_16789));
NAND2X1 g64616(.A (n_14102), .B (n_16787), .Y (n_16788));
NAND2X1 g64626(.A (n_16785), .B (n_14866), .Y (n_16786));
OAI21X1 g64646(.A0 (n_4051), .A1 (n_10603), .B0 (n_13606), .Y(n_16784));
INVX1 g64651(.A (n_16781), .Y (n_16782));
OAI21X1 g64657(.A0 (n_5137), .A1 (n_10489), .B0 (n_14155), .Y(n_16780));
AOI21X1 g64658(.A0 (n_11862), .A1 (n_9692), .B0 (n_27160), .Y(n_16778));
NOR2X1 g64664(.A (n_16501), .B (n_11354), .Y (n_16777));
AND2X1 g64672(.A (n_16775), .B (n_14845), .Y (n_16776));
NAND4X1 g64685(.A (n_7596), .B (n_13720), .C (n_15534), .D (n_8875),.Y (n_16774));
AND2X1 g64695(.A (n_16772), .B (n_9951), .Y (n_16773));
NAND2X1 g64715(.A (n_26882), .B (n_27688), .Y (n_17960));
NAND2X1 g64716(.A (n_16768), .B (n_16767), .Y (n_16769));
NAND2X1 g64717(.A (n_9944), .B (n_16765), .Y (n_16766));
NAND2X1 g64721(.A (n_13985), .B (n_19364), .Y (n_16764));
NAND2X1 g64722(.A (n_11309), .B (n_19364), .Y (n_16763));
NAND2X1 g64724(.A (n_14383), .B (n_13423), .Y (n_16762));
NAND2X1 g65402(.A (n_12840), .B (n_10896), .Y (n_16761));
NAND2X1 g64729(.A (n_14642), .B (n_16758), .Y (n_16759));
NAND2X1 g64733(.A (n_14378), .B (n_15039), .Y (n_17955));
NAND3X1 g64741(.A (n_16893), .B (n_7155), .C (n_12644), .Y (n_16757));
OR2X1 g64747(.A (n_12329), .B (n_16754), .Y (n_16756));
OR2X1 g64758(.A (n_14356), .B (n_18320), .Y (n_16753));
AND2X1 g64762(.A (n_14354), .B (n_7662), .Y (n_16752));
NAND3X1 g64763(.A (n_8633), .B (n_5371), .C (n_26467), .Y (n_16751));
NAND2X1 g64767(.A (n_18826), .B (n_17897), .Y (n_16749));
NOR2X1 g64769(.A (n_9821), .B (n_15574), .Y (n_16748));
NOR2X1 g64796(.A (n_16730), .B (n_14155), .Y (n_16746));
INVX1 g64797(.A (n_15092), .Y (n_16745));
NAND2X1 g64803(.A (n_26614), .B (n_14637), .Y (n_16744));
NAND2X1 g64809(.A (n_13970), .B (n_29014), .Y (n_16742));
INVX1 g64827(.A (n_15075), .Y (n_16740));
NAND2X1 g64829(.A (n_16738), .B (n_16737), .Y (n_16739));
NAND2X1 g64834(.A (n_13159), .B (n_17832), .Y (n_16733));
AND2X1 g64839(.A (n_14538), .B (n_11295), .Y (n_16732));
NAND2X1 g64840(.A (n_16730), .B (n_14565), .Y (n_16731));
NAND3X1 g64844(.A (n_26047), .B (n_16346), .C (n_19499), .Y(n_16728));
NOR2X1 g64849(.A (n_15254), .B (n_27160), .Y (n_16727));
INVX1 g64855(.A (n_15062), .Y (n_16726));
NOR2X1 g64857(.A (n_16724), .B (n_19961), .Y (n_16725));
AND2X1 g64863(.A (n_14431), .B (n_13058), .Y (n_16722));
INVX1 g64873(.A (n_16720), .Y (n_16721));
OR2X1 g64875(.A (n_9489), .B (n_18641), .Y (n_16719));
NAND2X1 g64876(.A (n_17197), .B (n_9564), .Y (n_16718));
INVX1 g64879(.A (n_17331), .Y (n_16717));
NAND2X1 g64881(.A (n_15886), .B (n_16715), .Y (n_16716));
NAND3X1 g64883(.A (n_16713), .B (n_9992), .C (n_7394), .Y (n_16714));
NAND2X1 g64885(.A (n_17982), .B (n_16711), .Y (n_16712));
NOR2X1 g64887(.A (n_13051), .B (n_15961), .Y (n_28894));
NOR2X1 g64890(.A (n_12503), .B (n_14647), .Y (n_16709));
AND2X1 g64893(.A (n_12207), .B (n_29074), .Y (n_16708));
NOR2X1 g64898(.A (n_14122), .B (n_13272), .Y (n_16707));
OR2X1 g64900(.A (n_12223), .B (n_15568), .Y (n_16706));
NAND2X1 g64903(.A (n_27077), .B (n_16704), .Y (n_16705));
OAI21X1 g64905(.A0 (n_6154), .A1 (n_19186), .B0 (n_21242), .Y(n_16703));
NOR2X1 g64908(.A (n_11258), .B (n_12912), .Y (n_16701));
NAND2X1 g64910(.A (n_12499), .B (n_15074), .Y (n_16700));
NAND2X1 g64915(.A (n_14353), .B (n_28692), .Y (n_17922));
NAND2X1 g64916(.A (n_14679), .B (n_14521), .Y (n_16696));
INVX1 g64921(.A (n_15036), .Y (n_16695));
NAND2X1 g64926(.A (n_13322), .B (n_10344), .Y (n_16694));
NAND2X1 g64929(.A (n_12302), .B (n_16754), .Y (n_16693));
NAND2X1 g64934(.A (n_12386), .B (n_29085), .Y (n_17920));
NAND2X1 g64937(.A (n_16650), .B (n_8719), .Y (n_16690));
INVX1 g64941(.A (n_15024), .Y (n_16689));
NAND2X1 g64943(.A (n_12221), .B (n_12907), .Y (n_16688));
NAND2X1 g64951(.A (n_14390), .B (n_16639), .Y (n_16687));
NAND2X1 g64952(.A (n_28809), .B (n_9472), .Y (n_16686));
NAND2X1 g64957(.A (n_9464), .B (n_16334), .Y (n_16685));
NAND2X1 g64962(.A (n_16683), .B (n_10543), .Y (n_16684));
NAND2X1 g64963(.A (n_16368), .B (n_9921), .Y (n_16682));
NAND2X1 g64964(.A (n_16680), .B (n_15511), .Y (n_16681));
AOI21X1 g64969(.A0 (n_3676), .A1 (n_16678), .B0 (n_15986), .Y(n_16679));
NOR2X1 g64972(.A (n_14161), .B (n_16676), .Y (n_28314));
AND2X1 g64976(.A (n_13298), .B (n_16674), .Y (n_16675));
OR2X1 g64979(.A (n_16672), .B (n_18617), .Y (n_16673));
NOR2X1 g64982(.A (n_16670), .B (n_7718), .Y (n_16671));
OR2X1 g64984(.A (n_12174), .B (n_17912), .Y (n_16669));
NOR2X1 g64987(.A (n_27505), .B (n_6036), .Y (n_16668));
NAND2X1 g64988(.A (n_14823), .B (n_16665), .Y (n_16666));
NAND2X1 g64990(.A (n_26614), .B (n_16663), .Y (n_16664));
NOR2X1 g64992(.A (n_10878), .B (n_13359), .Y (n_16660));
AOI21X1 g64994(.A0 (n_10082), .A1 (n_6991), .B0 (n_15776), .Y(n_16659));
NOR2X1 g64999(.A (n_14437), .B (n_12864), .Y (n_16658));
NOR2X1 g65004(.A (n_15098), .B (n_27028), .Y (n_16657));
NAND2X1 g65015(.A (n_15009), .B (n_14372), .Y (n_16656));
NAND2X1 g65020(.A (n_12935), .B (n_13801), .Y (n_16655));
NOR2X1 g65024(.A (n_7208), .B (n_14636), .Y (n_28878));
NAND2X1 g65028(.A (n_12433), .B (n_16652), .Y (n_16653));
OR2X1 g65030(.A (n_16650), .B (n_16649), .Y (n_16651));
INVX1 g65031(.A (n_16647), .Y (n_16648));
NAND2X1 g65035(.A (n_16645), .B (n_16644), .Y (n_16646));
NOR2X1 g65041(.A (n_9407), .B (n_10961), .Y (n_16641));
OR2X1 g65042(.A (n_16639), .B (n_29014), .Y (n_16640));
NAND2X1 g65043(.A (n_16637), .B (n_13031), .Y (n_16638));
OAI21X1 g65044(.A0 (n_9099), .A1 (n_6938), .B0 (n_15568), .Y(n_16636));
NOR2X1 g65045(.A (n_16634), .B (n_27919), .Y (n_16635));
NAND2X1 g65046(.A (n_28809), .B (n_14272), .Y (n_16633));
NAND2X1 g65058(.A (n_9743), .B (n_16398), .Y (n_16630));
NAND3X1 g65061(.A (n_11883), .B (n_14815), .C (n_26469), .Y(n_16629));
AND2X1 g65062(.A (n_15626), .B (n_27724), .Y (n_25516));
NAND2X1 g65065(.A (n_12508), .B (n_12896), .Y (n_16624));
NAND2X1 g65068(.A (n_11251), .B (n_13818), .Y (n_16623));
AOI21X1 g65073(.A0 (n_10547), .A1 (n_16621), .B0 (n_29102), .Y(n_16622));
AOI21X1 g65079(.A0 (n_10518), .A1 (n_14343), .B0 (n_17500), .Y(n_16617));
AND2X1 g65080(.A (n_12412), .B (n_14807), .Y (n_16616));
AND2X1 g65093(.A (n_13370), .B (n_16049), .Y (n_16612));
INVX1 g65096(.A (n_16610), .Y (n_16611));
NAND2X1 g65104(.A (n_5099), .B (n_12567), .Y (n_16608));
NAND3X1 g65107(.A (n_16674), .B (n_6948), .C (n_15109), .Y (n_16607));
OR2X1 g65109(.A (n_14942), .B (n_18266), .Y (n_16606));
NAND2X1 g65119(.A (n_12596), .B (n_11489), .Y (n_17882));
NAND2X1 g65122(.A (n_16187), .B (n_18353), .Y (n_16605));
AOI21X1 g65128(.A0 (n_9801), .A1 (n_9686), .B0 (n_2682), .Y(n_16604));
NAND2X1 g65133(.A (n_17217), .B (n_9363), .Y (n_16603));
NAND2X1 g65135(.A (n_20392), .B (n_16601), .Y (n_16602));
NAND3X1 g65141(.A (n_10048), .B (n_6291), .C (n_16599), .Y (n_16600));
NAND2X1 g65142(.A (n_12371), .B (n_14155), .Y (n_18281));
OR2X1 g65144(.A (n_14978), .B (n_18205), .Y (n_16597));
AND2X1 g65145(.A (n_13414), .B (n_16595), .Y (n_16596));
NAND2X1 g65150(.A (n_13357), .B (n_16593), .Y (n_16594));
NAND2X1 g65152(.A (n_12361), .B (n_27688), .Y (n_16592));
NOR2X1 g65153(.A (n_16590), .B (n_14671), .Y (n_29388));
NAND2X1 g65156(.A (n_16588), .B (n_7877), .Y (n_16589));
AND2X1 g65159(.A (n_16586), .B (n_15392), .Y (n_16587));
NAND2X1 g65162(.A (n_12315), .B (n_9410), .Y (n_17868));
NAND3X1 g65167(.A (n_27801), .B (n_16485), .C (n_19297), .Y(n_16584));
NOR2X1 g65168(.A (n_5819), .B (n_16582), .Y (n_16583));
OR2X1 g65170(.A (n_12163), .B (n_20558), .Y (n_16581));
AOI21X1 g65171(.A0 (n_9845), .A1 (n_6806), .B0 (n_16579), .Y(n_16580));
NAND2X1 g65174(.A (n_16577), .B (n_17240), .Y (n_16578));
OAI21X1 g65179(.A0 (n_9144), .A1 (n_7125), .B0 (n_9410), .Y(n_16576));
AND2X1 g65182(.A (n_16574), .B (n_10805), .Y (n_16575));
OR2X1 g65183(.A (n_12143), .B (n_27604), .Y (n_16573));
NAND2X1 g65184(.A (n_16572), .B (n_19433), .Y (n_18217));
NAND2X1 g65185(.A (n_12344), .B (n_16570), .Y (n_16571));
NAND2X1 g65186(.A (n_16568), .B (n_10320), .Y (n_16569));
NAND3X1 g65187(.A (n_10835), .B (n_3990), .C (n_12058), .Y (n_16567));
NOR2X1 g65188(.A (n_27899), .B (n_10012), .Y (n_25667));
NAND2X1 g65191(.A (n_17140), .B (n_16564), .Y (n_16565));
NAND2X1 g65193(.A (n_27446), .B (n_27445), .Y (n_16563));
NAND2X1 g65196(.A (n_12338), .B (n_9106), .Y (n_19247));
NAND2X1 g65199(.A (n_28877), .B (n_9509), .Y (n_16561));
NAND2X1 g65200(.A (n_12334), .B (n_16559), .Y (n_16560));
OR2X1 g65204(.A (n_16557), .B (n_16787), .Y (n_16558));
OR2X1 g65206(.A (n_12707), .B (n_16754), .Y (n_16555));
OAI21X1 g65207(.A0 (n_11436), .A1 (n_4436), .B0 (n_16553), .Y(n_16554));
NAND2X1 g65211(.A (n_16551), .B (n_16550), .Y (n_16552));
OR2X1 g65217(.A (n_12153), .B (n_15894), .Y (n_16549));
NOR2X1 g65220(.A (n_15291), .B (n_8701), .Y (n_16548));
NAND2X1 g65225(.A (n_16543), .B (n_16704), .Y (n_16544));
INVX1 g65230(.A (n_14926), .Y (n_16542));
NAND2X1 g65232(.A (n_16540), .B (n_16539), .Y (n_16541));
NAND2X1 g65234(.A (n_16537), .B (n_15949), .Y (n_16538));
AOI21X1 g65235(.A0 (n_8173), .A1 (n_9681), .B0 (n_19961), .Y(n_16536));
NAND2X1 g65237(.A (n_20003), .B (n_16534), .Y (n_16535));
OR2X1 g65243(.A (n_16532), .B (n_12298), .Y (n_16533));
NOR2X1 g65250(.A (n_15415), .B (n_7302), .Y (n_16530));
NOR2X1 g65252(.A (n_13607), .B (n_14707), .Y (n_16529));
NAND2X1 g65253(.A (n_18648), .B (n_16527), .Y (n_16528));
NAND2X1 g65255(.A (n_12811), .B (n_18205), .Y (n_17848));
NAND2X1 g65257(.A (n_12150), .B (n_17567), .Y (n_16526));
NAND2X1 g65270(.A (n_15543), .B (n_15902), .Y (n_16525));
INVX1 g65274(.A (n_17153), .Y (n_16524));
NAND2X1 g65286(.A (n_16593), .B (n_10254), .Y (n_16523));
NAND2X1 g65289(.A (n_18619), .B (n_12892), .Y (n_16522));
NAND2X1 g65291(.A (n_12286), .B (n_16787), .Y (n_17835));
NOR2X1 g65293(.A (n_13454), .B (n_9727), .Y (n_25599));
NAND2X1 g65297(.A (n_16557), .B (n_16519), .Y (n_16520));
NAND2X1 g65300(.A (n_9726), .B (n_16321), .Y (n_16518));
NAND2X1 g65302(.A (n_12277), .B (n_11319), .Y (n_16517));
NAND2X1 g65309(.A (n_14587), .B (n_12648), .Y (n_16515));
NAND2X1 g65313(.A (n_16711), .B (n_14361), .Y (n_16514));
NAND2X1 g65318(.A (n_15111), .B (n_16512), .Y (n_16513));
NAND2X1 g65319(.A (n_16510), .B (n_14571), .Y (n_16511));
INVX1 g65320(.A (n_14897), .Y (n_16509));
NAND2X1 g65322(.A (n_27130), .B (n_11576), .Y (n_18437));
NAND2X1 g65323(.A (n_17217), .B (n_10242), .Y (n_16508));
NAND2X1 g65324(.A (n_14564), .B (n_17411), .Y (n_18298));
NAND3X1 g65335(.A (n_29198), .B (n_4909), .C (n_10121), .Y (n_16507));
NOR2X1 g65336(.A (n_12787), .B (n_10562), .Y (n_16506));
AND2X1 g65337(.A (n_12195), .B (n_17302), .Y (n_16505));
AND2X1 g65340(.A (n_10725), .B (n_16503), .Y (n_16504));
AND2X1 g65341(.A (n_12185), .B (n_16501), .Y (n_16502));
INVX1 g65342(.A (n_14889), .Y (n_16500));
NAND3X1 g65352(.A (n_12532), .B (n_10390), .C (n_28161), .Y(n_16499));
NOR2X1 g65355(.A (n_12728), .B (n_8962), .Y (n_16497));
OAI21X1 g65398(.A0 (n_2109), .A1 (n_7410), .B0 (n_12466), .Y(n_16496));
AND2X1 g65358(.A (n_10717), .B (n_18114), .Y (n_16495));
NAND3X1 g65364(.A (n_12802), .B (n_6314), .C (n_10065), .Y (n_16494));
NAND3X1 g65404(.A (n_5525), .B (n_16492), .C (n_12292), .Y (n_16493));
OAI21X1 g65412(.A0 (n_7411), .A1 (n_5817), .B0 (n_12746), .Y(n_16491));
NAND3X1 g65413(.A (n_9328), .B (n_9450), .C (n_8643), .Y (n_16490));
AOI21X1 g65414(.A0 (n_16488), .A1 (n_9093), .B0 (n_1132), .Y(n_16489));
AOI21X1 g65415(.A0 (n_6269), .A1 (n_16988), .B0 (n_12806), .Y(n_16487));
AOI21X1 g65417(.A0 (n_16485), .A1 (n_11861), .B0 (n_15894), .Y(n_16486));
OAI21X1 g65422(.A0 (n_4026), .A1 (n_29297), .B0 (n_16543), .Y(n_16484));
INVX1 g65429(.A (n_14873), .Y (n_16482));
OR2X1 g65436(.A (n_12656), .B (n_16480), .Y (n_16481));
NAND3X1 g65438(.A (n_9348), .B (n_7733), .C (n_14598), .Y (n_16479));
AOI21X1 g65439(.A0 (n_16477), .A1 (n_8995), .B0 (n_20010), .Y(n_16478));
AND2X1 g65442(.A (n_12675), .B (n_16787), .Y (n_16476));
AOI21X1 g65443(.A0 (n_14274), .A1 (n_26386), .B0 (n_12100), .Y(n_16474));
AOI21X1 g65444(.A0 (n_14482), .A1 (n_2720), .B0 (n_16472), .Y(n_16473));
AND2X1 g65450(.A (n_12377), .B (n_16754), .Y (n_16471));
AOI21X1 g65451(.A0 (n_19110), .A1 (n_2479), .B0 (n_16469), .Y(n_16470));
NAND2X1 g65456(.A (n_13084), .B (n_6066), .Y (n_16468));
AND2X1 g65458(.A (n_12732), .B (n_16466), .Y (n_16467));
NAND2X1 g65459(.A (n_12661), .B (n_12247), .Y (n_16465));
NAND2X1 g65460(.A (n_12276), .B (n_15894), .Y (n_16464));
AOI21X1 g65461(.A0 (n_19114), .A1 (n_5462), .B0 (n_16582), .Y(n_16463));
NAND3X1 g65466(.A (n_15315), .B (n_15909), .C (n_15045), .Y(n_16462));
NAND3X1 g65471(.A (n_9209), .B (n_11321), .C (n_8486), .Y (n_16461));
AND2X1 g65475(.A (n_12845), .B (n_27099), .Y (n_16460));
AOI21X1 g65479(.A0 (n_15137), .A1 (n_9647), .B0 (n_14589), .Y(n_16459));
AND2X1 g65485(.A (n_12710), .B (n_15586), .Y (n_16457));
NOR2X1 g65486(.A (n_12645), .B (n_13073), .Y (n_16456));
AOI21X1 g65497(.A0 (n_12722), .A1 (n_11193), .B0 (n_15708), .Y(n_16455));
NAND3X1 g65501(.A (n_4784), .B (n_8884), .C (n_10272), .Y (n_16454));
NAND2X1 g65503(.A (n_7458), .B (n_18619), .Y (n_16453));
OR2X1 g65505(.A (n_12727), .B (n_15776), .Y (n_16452));
NAND2X1 g65510(.A (n_9047), .B (n_20003), .Y (n_16450));
OR2X1 g65511(.A (n_12379), .B (n_13604), .Y (n_16449));
NAND4X1 g65513(.A (n_12673), .B (n_13472), .C (n_6918), .D (n_9005),.Y (n_16448));
OAI21X1 g65515(.A0 (n_9167), .A1 (n_10495), .B0 (n_12779), .Y(n_16447));
NAND2X1 g65519(.A (n_12682), .B (n_18266), .Y (n_16446));
OR2X1 g65521(.A (n_12639), .B (n_13083), .Y (n_16445));
INVX1 g65522(.A (n_14850), .Y (n_16444));
NAND2X1 g65524(.A (n_12750), .B (n_9593), .Y (n_16443));
AOI21X1 g65527(.A0 (n_9755), .A1 (n_3317), .B0 (n_16441), .Y(n_16442));
AOI21X1 g65534(.A0 (n_7679), .A1 (n_16439), .B0 (n_15894), .Y(n_16440));
NAND2X1 g65545(.A (n_11836), .B (n_13508), .Y (n_16437));
NAND3X1 g65546(.A (n_10266), .B (n_9115), .C (n_12918), .Y (n_16436));
OR2X1 g65547(.A (n_12824), .B (n_16434), .Y (n_16435));
NAND2X1 g65548(.A (n_7318), .B (n_18648), .Y (n_16433));
OR2X1 g65549(.A (n_12749), .B (n_27688), .Y (n_16432));
AOI21X1 g65552(.A0 (n_9513), .A1 (n_12052), .B0 (n_14055), .Y(n_16431));
NAND2X1 g65557(.A (n_12640), .B (n_9236), .Y (n_16430));
OR2X1 g65561(.A (n_12326), .B (n_15418), .Y (n_16429));
OAI21X1 g65562(.A0 (n_4767), .A1 (n_4689), .B0 (n_9369), .Y(n_19182));
NAND3X1 g65565(.A (n_15103), .B (n_8447), .C (n_15042), .Y (n_16428));
OAI21X1 g65566(.A0 (n_3087), .A1 (n_8452), .B0 (n_16426), .Y(n_16427));
AND2X1 g65568(.A (n_12529), .B (n_15580), .Y (n_16425));
NAND2X1 g65572(.A (n_11888), .B (n_27140), .Y (n_16424));
AOI21X1 g65575(.A0 (n_15628), .A1 (n_6989), .B0 (n_12896), .Y(n_16423));
NAND3X1 g65576(.A (n_16421), .B (n_14087), .C (n_14616), .Y(n_16422));
OAI21X1 g65578(.A0 (n_3421), .A1 (n_11307), .B0 (n_12706), .Y(n_16420));
AOI21X1 g65582(.A0 (n_14242), .A1 (n_1340), .B0 (n_9017), .Y(n_16419));
NAND3X1 g65584(.A (n_16416), .B (n_6451), .C (n_12025), .Y (n_16417));
AND2X1 g65588(.A (n_12562), .B (n_16414), .Y (n_16415));
AND2X1 g65589(.A (n_12561), .B (n_16412), .Y (n_16413));
OR2X1 g65590(.A (n_12558), .B (n_28692), .Y (n_16411));
NAND3X1 g65597(.A (n_29204), .B (n_6556), .C (n_7406), .Y (n_16410));
AND2X1 g65600(.A (n_12548), .B (n_14155), .Y (n_16409));
AOI21X1 g65603(.A0 (n_12446), .A1 (n_1238), .B0 (n_10264), .Y(n_16408));
OAI21X1 g65607(.A0 (n_5014), .A1 (n_15388), .B0 (n_16406), .Y(n_16407));
AOI21X1 g65615(.A0 (n_12478), .A1 (n_3394), .B0 (n_12006), .Y(n_16405));
INVX1 g65617(.A (n_14825), .Y (n_16404));
AOI21X1 g65620(.A0 (n_5682), .A1 (n_8922), .B0 (n_13571), .Y(n_16403));
NAND2X1 g65622(.A (n_12521), .B (n_11277), .Y (n_16402));
NAND3X1 g65632(.A (n_15186), .B (n_14517), .C (n_15011), .Y(n_16401));
INVX1 g65634(.A (n_14818), .Y (n_16400));
OAI21X1 g65639(.A0 (n_5324), .A1 (n_12019), .B0 (n_16398), .Y(n_16399));
NOR2X1 g65640(.A (n_10933), .B (n_12225), .Y (n_16397));
NAND2X1 g65641(.A (n_12501), .B (n_17939), .Y (n_16396));
NAND3X1 g65654(.A (n_4243), .B (n_16394), .C (n_14386), .Y (n_16395));
NOR2X1 g65655(.A (n_12487), .B (n_13003), .Y (n_16393));
NAND3X1 g65662(.A (n_16391), .B (n_9817), .C (n_16390), .Y (n_16392));
AOI21X1 g65664(.A0 (n_12505), .A1 (n_15575), .B0 (n_11400), .Y(n_16389));
NAND2X1 g65665(.A (n_12471), .B (n_9803), .Y (n_16388));
AOI21X1 g65667(.A0 (n_14146), .A1 (n_5589), .B0 (n_17912), .Y(n_16387));
NAND2X1 g65675(.A (n_7371), .B (n_16637), .Y (n_16386));
NAND2X1 g65677(.A (n_11686), .B (n_26375), .Y (n_16385));
AND2X1 g65680(.A (n_12755), .B (n_9819), .Y (n_16384));
AOI21X1 g65682(.A0 (n_8037), .A1 (n_15566), .B0 (n_17500), .Y(n_16383));
INVX1 g65684(.A (n_14804), .Y (n_16382));
NAND2X1 g65688(.A (n_9846), .B (n_16645), .Y (n_16381));
NAND2X1 g65689(.A (n_10356), .B (n_20392), .Y (n_16380));
OAI21X1 g65691(.A0 (n_15310), .A1 (n_12559), .B0 (n_6819), .Y(n_16379));
NAND2X1 g65693(.A (n_12049), .B (n_15304), .Y (n_16378));
NAND2X1 g65697(.A (n_11742), .B (n_16325), .Y (n_16377));
AOI21X1 g65699(.A0 (n_14213), .A1 (n_1347), .B0 (n_16375), .Y(n_16376));
AOI21X1 g65702(.A0 (n_10904), .A1 (n_11495), .B0 (n_15039), .Y(n_16374));
NAND2X1 g65703(.A (n_12437), .B (n_15411), .Y (n_16373));
INVX1 g65705(.A (n_14797), .Y (n_16372));
OAI21X1 g65713(.A0 (n_8289), .A1 (n_28037), .B0 (n_8805), .Y(n_16371));
NAND2X1 g65716(.A (n_11857), .B (n_16368), .Y (n_16369));
AND2X1 g65725(.A (n_12408), .B (n_16366), .Y (n_16367));
AOI21X1 g65729(.A0 (n_10510), .A1 (n_8438), .B0 (n_28642), .Y(n_16365));
NAND2X1 g65731(.A (n_12400), .B (n_11560), .Y (n_16364));
NAND2X1 g65740(.A (n_7384), .B (n_18587), .Y (n_16361));
AOI21X1 g65743(.A0 (n_16359), .A1 (n_13971), .B0 (n_16358), .Y(n_16360));
NAND2X1 g65748(.A (n_7488), .B (n_18582), .Y (n_16357));
AOI21X1 g65750(.A0 (n_10634), .A1 (n_27991), .B0 (n_19791), .Y(n_16356));
AOI21X1 g65752(.A0 (n_13119), .A1 (n_13851), .B0 (n_16434), .Y(n_16355));
AOI21X1 g65755(.A0 (n_5659), .A1 (n_9115), .B0 (n_16835), .Y(n_16354));
AOI21X1 g65759(.A0 (n_16351), .A1 (n_8172), .B0 (n_9819), .Y(n_16352));
INVX1 g65760(.A (n_14790), .Y (n_16349));
INVX1 g65765(.A (n_14788), .Y (n_16348));
AOI21X1 g65768(.A0 (n_16346), .A1 (n_13799), .B0 (n_17500), .Y(n_16347));
AND2X1 g65774(.A (n_12244), .B (n_17912), .Y (n_16345));
AOI21X1 g65779(.A0 (n_16342), .A1 (n_11290), .B0 (n_6889), .Y(n_16343));
AOI21X1 g65781(.A0 (n_16280), .A1 (n_11864), .B0 (n_27688), .Y(n_16341));
AND2X1 g65789(.A (n_12565), .B (n_18237), .Y (n_16340));
AOI21X1 g65802(.A0 (n_16338), .A1 (n_11387), .B0 (n_12849), .Y(n_16339));
NOR2X1 g65806(.A (n_12352), .B (n_13942), .Y (n_16337));
OAI21X1 g65808(.A0 (n_4143), .A1 (n_27746), .B0 (n_16334), .Y(n_16336));
NAND3X1 g65811(.A (n_9127), .B (n_5175), .C (n_11956), .Y (n_16333));
NAND2X1 g65822(.A (n_10115), .B (n_16331), .Y (n_16332));
NAND2X1 g65824(.A (n_6929), .B (n_16595), .Y (n_16330));
AOI21X1 g65826(.A0 (n_8634), .A1 (n_6755), .B0 (n_16328), .Y(n_16329));
NAND2X1 g65827(.A (n_8397), .B (n_16368), .Y (n_16327));
NAND2X1 g65829(.A (n_10213), .B (n_16325), .Y (n_16326));
NAND2X1 g65833(.A (n_9850), .B (n_16323), .Y (n_16324));
NAND2X1 g65834(.A (n_9736), .B (n_16321), .Y (n_16322));
NAND2X1 g65835(.A (n_9756), .B (n_15195), .Y (n_16320));
NAND2X1 g65837(.A (n_13090), .B (n_10134), .Y (n_16319));
NAND2X1 g65844(.A (n_13055), .B (n_10220), .Y (n_16318));
NAND2X1 g65847(.A (n_6189), .B (n_16775), .Y (n_16317));
NAND2X1 g65848(.A (n_12998), .B (n_9929), .Y (n_16316));
NAND2X1 g65849(.A (n_12981), .B (n_9916), .Y (n_16315));
NAND2X1 g65851(.A (n_9987), .B (n_12972), .Y (n_16314));
NOR2X1 g65859(.A (n_8704), .B (n_12830), .Y (n_16313));
AOI21X1 g65860(.A0 (n_9706), .A1 (n_9410), .B0 (n_8667), .Y(n_16312));
OAI22X1 g65876(.A0 (n_6797), .A1 (n_6620), .B0 (n_2327), .B1(n_9142), .Y (n_16310));
NOR2X1 g65877(.A (n_12479), .B (n_12531), .Y (n_16309));
AOI21X1 g65881(.A0 (n_9627), .A1 (n_14624), .B0 (n_8291), .Y(n_16308));
AOI21X1 g65885(.A0 (n_10345), .A1 (n_27604), .B0 (n_12593), .Y(n_16306));
AOI21X1 g65888(.A0 (n_9814), .A1 (n_11400), .B0 (n_12785), .Y(n_16304));
AOI21X1 g65889(.A0 (n_26381), .A1 (n_13804), .B0 (n_12422), .Y(n_16302));
AOI21X1 g65893(.A0 (n_8883), .A1 (n_7649), .B0 (n_16300), .Y(n_16301));
NAND2X1 g65899(.A (n_12481), .B (n_15101), .Y (n_16299));
OAI21X1 g65909(.A0 (n_14500), .A1 (n_8945), .B0 (n_9753), .Y(n_16298));
NAND2X1 g65911(.A (n_12647), .B (n_10238), .Y (n_16297));
NAND4X1 g65915(.A (n_7603), .B (n_11500), .C (n_7531), .D (n_8990),.Y (n_16296));
NAND3X1 g65923(.A (n_10890), .B (n_7296), .C (n_16652), .Y (n_16294));
NAND2X1 g65929(.A (n_12654), .B (n_11811), .Y (n_16293));
NAND2X1 g65931(.A (n_12699), .B (n_11839), .Y (n_16292));
AOI22X1 g65934(.A0 (n_4408), .A1 (n_7832), .B0 (n_16290), .B1(n_7410), .Y (n_16291));
NAND2X1 g65936(.A (n_12509), .B (n_11758), .Y (n_16289));
NAND2X1 g65938(.A (n_12473), .B (n_11851), .Y (n_16288));
NAND2X1 g65939(.A (n_12369), .B (n_11750), .Y (n_16287));
NAND2X1 g65940(.A (n_12444), .B (n_8294), .Y (n_16286));
NAND2X1 g65941(.A (n_12701), .B (n_11740), .Y (n_16285));
MX2X1 g65944(.A (n_14054), .B (n_14343), .S0 (n_19896), .Y (n_16284));
MX2X1 g65948(.A (n_14413), .B (n_16621), .S0 (n_29048), .Y (n_16283));
AOI21X1 g65949(.A0 (n_19186), .A1 (n_28632), .B0 (n_11286), .Y(n_16282));
MX2X1 g65953(.A (n_16280), .B (n_14324), .S0 (n_16279), .Y (n_16281));
MX2X1 g65955(.A (n_14061), .B (n_13418), .S0 (n_15894), .Y (n_16278));
INVX1 g66023(.A (n_14721), .Y (n_16275));
NOR2X1 g66034(.A (n_16271), .B (n_16434), .Y (n_16272));
NAND2X1 g66052(.A (n_9905), .B (n_18785), .Y (n_16268));
NAND2X1 g66056(.A (n_16266), .B (n_15894), .Y (n_16267));
INVX1 g66058(.A (n_16264), .Y (n_16265));
NAND2X1 g66067(.A (n_11718), .B (n_19364), .Y (n_16263));
INVX1 g66070(.A (n_14712), .Y (n_17979));
INVX1 g66086(.A (n_16893), .Y (n_16262));
NOR2X1 g66114(.A (n_28815), .B (n_19791), .Y (n_16259));
NAND2X1 g66116(.A (n_11834), .B (n_101), .Y (n_16257));
INVX1 g66147(.A (n_14702), .Y (n_19060));
NAND2X1 g66210(.A (n_16040), .B (n_1268), .Y (n_16254));
OR4X1 g66218(.A (n_4709), .B (n_8945), .C (n_16204), .D (n_7858), .Y(n_17672));
INVX1 g66228(.A (n_16251), .Y (n_16253));
NAND2X1 g66233(.A (n_16082), .B (n_3932), .Y (n_16250));
INVX1 g66240(.A (n_14689), .Y (n_17969));
NAND2X2 g66249(.A (n_29203), .B (n_28444), .Y (n_16249));
NAND2X1 g66275(.A (n_16245), .B (n_4755), .Y (n_16246));
NAND2X1 g66336(.A (n_15958), .B (n_18320), .Y (n_16240));
INVX1 g66350(.A (n_14676), .Y (n_16238));
NOR2X1 g66352(.A (n_16236), .B (n_19364), .Y (n_16237));
INVX1 g66354(.A (n_14675), .Y (n_17980));
NAND2X1 g66368(.A (n_13882), .B (n_27688), .Y (n_16229));
INVX1 g66369(.A (n_14670), .Y (n_16228));
NAND2X1 g66375(.A (n_16225), .B (n_28692), .Y (n_16226));
NAND2X1 g66379(.A (n_15918), .B (n_9264), .Y (n_16224));
NAND2X1 g66382(.A (n_11878), .B (n_19395), .Y (n_16223));
NAND2X1 g66454(.A (n_10182), .B (n_6185), .Y (n_16221));
INVX2 g66464(.A (n_14659), .Y (n_18996));
NAND2X1 g66472(.A (n_10391), .B (n_15039), .Y (n_16217));
NAND2X1 g66476(.A (n_16005), .B (n_9783), .Y (n_16215));
NOR2X1 g66496(.A (n_17411), .B (n_12061), .Y (n_16213));
NAND2X1 g66544(.A (n_15990), .B (n_4898), .Y (n_16209));
INVX1 g66547(.A (n_16207), .Y (n_16208));
OR4X1 g66564(.A (n_18266), .B (n_27757), .C (n_16204), .D (n_9482),.Y (n_18807));
NAND2X1 g66598(.A (n_16199), .B (n_16198), .Y (n_16200));
INVX1 g66602(.A (n_16196), .Y (n_16197));
INVX1 g66616(.A (n_14626), .Y (n_17660));
NAND2X1 g66619(.A (n_28692), .B (n_28136), .Y (n_16195));
NOR2X1 g66667(.A (n_16187), .B (n_16434), .Y (n_16188));
INVX1 g66668(.A (n_14617), .Y (n_16186));
NAND2X1 g66671(.A (n_16184), .B (n_14155), .Y (n_16185));
INVX1 g66680(.A (n_14615), .Y (n_16183));
INVX1 g66687(.A (n_14610), .Y (n_16182));
INVX1 g66689(.A (n_14608), .Y (n_25614));
INVX1 g66701(.A (n_14607), .Y (n_18811));
NOR3X1 g66714(.A (n_16787), .B (n_8116), .C (n_9838), .Y (n_16177));
INVX1 g66728(.A (n_16176), .Y (n_18765));
NAND2X1 g66737(.A (n_16174), .B (n_12896), .Y (n_16175));
INVX1 g66742(.A (n_16172), .Y (n_17655));
AND2X1 g66771(.A (n_13076), .B (n_16480), .Y (n_16168));
NAND2X1 g66777(.A (n_16163), .B (n_11300), .Y (n_16164));
INVX1 g66778(.A (n_14594), .Y (n_16162));
INVX1 g66798(.A (n_14590), .Y (n_16161));
INVX1 g66816(.A (n_17147), .Y (n_16157));
NAND2X1 g66830(.A (n_16123), .B (n_8892), .Y (n_16154));
NOR2X1 g66833(.A (n_12023), .B (n_9038), .Y (n_16153));
NOR2X1 g66846(.A (n_9084), .B (n_16080), .Y (n_17649));
INVX1 g66868(.A (n_28326), .Y (n_16151));
INVX1 g66869(.A (n_28327), .Y (n_16149));
INVX1 g66888(.A (n_16144), .Y (n_16146));
OR2X1 g66892(.A (n_16142), .B (n_6534), .Y (n_16143));
NOR2X1 g66893(.A (n_10302), .B (n_9418), .Y (n_16141));
NAND2X1 g66903(.A (n_17723), .B (n_16390), .Y (n_17645));
AND2X1 g66911(.A (n_11677), .B (n_5329), .Y (n_16140));
OR2X1 g66912(.A (n_16139), .B (n_17571), .Y (n_18007));
INVX1 g66931(.A (n_16137), .Y (n_16138));
OR2X1 g66934(.A (n_12564), .B (n_11261), .Y (n_25720));
AND2X1 g66952(.A (n_12113), .B (n_13519), .Y (n_16135));
AOI21X1 g66954(.A0 (n_1744), .A1 (n_1353), .B0 (n_11715), .Y(n_16134));
INVX1 g66957(.A (n_16132), .Y (n_16133));
NAND2X1 g66969(.A (n_16130), .B (n_8105), .Y (n_16131));
NAND2X1 g66974(.A (n_10782), .B (n_8824), .Y (n_16129));
INVX1 g66994(.A (n_16126), .Y (n_16127));
INVX1 g67002(.A (n_14544), .Y (n_17643));
NOR2X1 g67010(.A (n_8261), .B (n_7212), .Y (n_16125));
NAND2X1 g67015(.A (n_16123), .B (n_4881), .Y (n_16124));
INVX1 g67032(.A (n_27161), .Y (n_16118));
NAND2X1 g67052(.A (n_5537), .B (n_12918), .Y (n_16116));
NAND2X1 g67061(.A (n_11931), .B (n_11701), .Y (n_16115));
NOR2X1 g67102(.A (n_5686), .B (n_12023), .Y (n_28248));
NOR2X1 g67111(.A (n_12964), .B (n_5319), .Y (n_16113));
INVX1 g67116(.A (n_16111), .Y (n_16112));
INVX1 g67119(.A (n_16817), .Y (n_16110));
INVX1 g67145(.A (n_16108), .Y (n_25758));
NOR2X1 g67151(.A (n_11948), .B (n_6056), .Y (n_16106));
NOR2X1 g67160(.A (n_2409), .B (n_8824), .Y (n_19880));
NAND2X1 g67166(.A (n_16103), .B (n_9787), .Y (n_16104));
AND2X1 g67174(.A (n_1361), .B (n_10332), .Y (n_16102));
NOR2X1 g67191(.A (n_16100), .B (n_9084), .Y (n_16101));
NAND2X1 g67193(.A (n_16097), .B (n_9913), .Y (n_16098));
NAND2X1 g67196(.A (n_12077), .B (n_13134), .Y (n_16096));
NAND2X1 g67213(.A (n_10680), .B (n_29173), .Y (n_17632));
INVX1 g67215(.A (n_14497), .Y (n_16095));
NAND2X1 g67218(.A (n_14585), .B (n_27290), .Y (n_16094));
NAND2X1 g67226(.A (n_16391), .B (n_13172), .Y (n_16093));
INVX1 g67230(.A (n_16844), .Y (n_16092));
NAND2X1 g67232(.A (n_16090), .B (n_16089), .Y (n_16091));
OR2X1 g67264(.A (n_28804), .B (n_17567), .Y (n_18756));
OR2X1 g67265(.A (n_29000), .B (n_11277), .Y (n_16087));
NAND2X1 g67266(.A (n_11647), .B (n_8486), .Y (n_16086));
INVX1 g67273(.A (n_16084), .Y (n_17630));
NAND2X1 g67282(.A (n_16082), .B (n_11916), .Y (n_16083));
NAND2X1 g67300(.A (n_16080), .B (n_3080), .Y (n_16081));
INVX1 g67309(.A (n_16078), .Y (n_16079));
NAND2X1 g67330(.A (n_16076), .B (n_10269), .Y (n_16077));
INVX1 g67352(.A (n_16074), .Y (n_16075));
NAND2X1 g67354(.A (n_16072), .B (n_10171), .Y (n_16073));
NAND2X1 g67355(.A (n_10193), .B (n_16070), .Y (n_16071));
NAND2X1 g67356(.A (n_10193), .B (n_16068), .Y (n_16069));
NOR2X1 g67357(.A (n_13082), .B (n_10136), .Y (n_18018));
NAND2X1 g67369(.A (n_10693), .B (n_16070), .Y (n_16067));
NOR2X1 g67375(.A (n_12032), .B (n_8427), .Y (n_28257));
NAND2X1 g67377(.A (n_8927), .B (n_9783), .Y (n_16065));
INVX1 g67380(.A (n_14440), .Y (n_16064));
OR2X1 g67387(.A (n_10609), .B (n_6534), .Y (n_16063));
AOI21X1 g65396(.A0 (n_14704), .A1 (n_3943), .B0 (n_11233), .Y(n_16061));
NOR2X1 g67411(.A (n_11530), .B (n_10046), .Y (n_17624));
INVX1 g67419(.A (n_16057), .Y (n_16058));
NAND2X1 g67446(.A (n_8473), .B (n_8968), .Y (n_16055));
NAND2X1 g67456(.A (n_10575), .B (n_28444), .Y (n_16054));
NAND2X1 g67489(.A (n_16052), .B (n_16051), .Y (n_16053));
NOR2X1 g67503(.A (n_8830), .B (n_10484), .Y (n_16050));
AOI21X1 g67530(.A0 (n_1883), .A1 (n_3566), .B0 (n_26381), .Y(n_16048));
NOR2X1 g67544(.A (n_8842), .B (n_9265), .Y (n_16046));
INVX1 g67552(.A (n_16044), .Y (n_16045));
NAND2X1 g67579(.A (n_16040), .B (n_27070), .Y (n_16041));
NAND2X1 g67592(.A (n_13898), .B (n_27688), .Y (n_18153));
NAND2X1 g67598(.A (n_7767), .B (n_10174), .Y (n_16039));
NOR2X1 g67602(.A (n_12029), .B (n_11845), .Y (n_16038));
OAI21X1 g67608(.A0 (n_4712), .A1 (n_2254), .B0 (n_27141), .Y(n_16037));
AND2X1 g67631(.A (n_10147), .B (n_13912), .Y (n_19021));
INVX1 g67643(.A (n_14357), .Y (n_16032));
NOR2X1 g67660(.A (n_15105), .B (n_6889), .Y (n_17605));
INVX1 g67663(.A (n_16030), .Y (n_16031));
NOR2X1 g67667(.A (n_3467), .B (n_27290), .Y (n_19854));
NAND2X1 g67694(.A (n_8213), .B (n_6005), .Y (n_16027));
INVX1 g67696(.A (n_26802), .Y (n_18333));
INVX1 g67714(.A (n_16023), .Y (n_16024));
AND2X1 g67723(.A (n_1497), .B (n_10489), .Y (n_16022));
NAND2X1 g67725(.A (n_10279), .B (n_11835), .Y (n_16020));
NOR2X1 g67730(.A (n_7282), .B (n_11815), .Y (n_16019));
INVX1 g67742(.A (n_16017), .Y (n_16018));
NOR2X1 g67747(.A (n_8803), .B (n_11778), .Y (n_16016));
INVX1 g67748(.A (n_16013), .Y (n_16014));
INVX1 g67761(.A (n_16009), .Y (n_16010));
NAND2X1 g67768(.A (n_16007), .B (n_10049), .Y (n_16008));
AND2X1 g67779(.A (n_16006), .B (n_16005), .Y (n_20705));
INVX1 g67788(.A (n_14306), .Y (n_18911));
INVX1 g67794(.A (n_16003), .Y (n_16004));
NAND3X1 g67798(.A (n_28578), .B (n_27099), .C (n_15371), .Y(n_16002));
AND2X1 g67802(.A (n_16000), .B (n_12014), .Y (n_25718));
NAND2X1 g67829(.A (n_10295), .B (n_15998), .Y (n_15999));
NAND2X1 g67840(.A (n_10598), .B (n_15997), .Y (n_18085));
AOI21X1 g67841(.A0 (n_13974), .A1 (n_1989), .B0 (n_9814), .Y(n_15996));
NAND2X1 g67843(.A (n_12613), .B (n_9106), .Y (n_17598));
NOR2X1 g67850(.A (n_12071), .B (n_11914), .Y (n_15994));
INVX1 g67871(.A (n_15992), .Y (n_15993));
INVX1 g67883(.A (n_14264), .Y (n_15991));
NAND2X1 g67887(.A (n_14725), .B (n_15990), .Y (n_19276));
NOR2X1 g67899(.A (n_12091), .B (n_5689), .Y (n_15988));
NOR2X1 g67900(.A (n_7596), .B (n_9783), .Y (n_15987));
NAND2X1 g67910(.A (n_12495), .B (n_15986), .Y (n_18241));
INVX1 g67916(.A (n_15984), .Y (n_15985));
NOR2X1 g67918(.A (n_11993), .B (n_6128), .Y (n_15983));
NOR2X1 g67927(.A (n_11981), .B (n_9404), .Y (n_15982));
AND2X1 g67957(.A (n_27122), .B (n_5620), .Y (n_15979));
NOR2X1 g67962(.A (n_12099), .B (n_12420), .Y (n_15977));
NAND2X1 g67964(.A (n_17328), .B (n_17689), .Y (n_15976));
NOR2X1 g67980(.A (n_13940), .B (n_11027), .Y (n_15972));
OR2X1 g67997(.A (n_15969), .B (n_15968), .Y (n_15970));
NAND2X1 g68022(.A (n_8824), .B (n_15966), .Y (n_15967));
AOI21X1 g65394(.A0 (n_7319), .A1 (n_11989), .B0 (n_6534), .Y(n_15965));
NAND2X1 g68056(.A (n_9429), .B (n_29256), .Y (n_15964));
NAND2X1 g68057(.A (n_16123), .B (n_7344), .Y (n_15963));
NOR2X1 g68081(.A (n_13740), .B (n_15961), .Y (n_25522));
NAND2X1 g68088(.A (n_9906), .B (n_15714), .Y (n_15960));
NAND2X1 g68094(.A (n_15958), .B (n_1198), .Y (n_29411));
NOR2X1 g68109(.A (n_12073), .B (n_8928), .Y (n_15956));
NAND2X1 g68115(.A (n_11102), .B (n_15104), .Y (n_15955));
INVX1 g68123(.A (n_14182), .Y (n_15954));
NAND2X1 g68126(.A (n_15952), .B (n_11084), .Y (n_15953));
NAND2X1 g68135(.A (n_13770), .B (n_29102), .Y (n_15951));
AND2X1 g68158(.A (n_15949), .B (n_16100), .Y (n_15950));
INVX1 g68159(.A (n_15947), .Y (n_15948));
INVX1 g68180(.A (n_14156), .Y (n_15945));
NAND2X1 g68187(.A (n_13766), .B (n_19896), .Y (n_15944));
NAND2X1 g68192(.A (n_4386), .B (n_15942), .Y (n_15943));
INVX1 g68202(.A (n_20853), .Y (n_15941));
NAND2X1 g68208(.A (n_9635), .B (n_4486), .Y (n_15940));
INVX1 g68211(.A (n_20468), .Y (n_15939));
NOR2X1 g68224(.A (n_11768), .B (n_3398), .Y (n_15936));
INVX1 g68230(.A (n_15934), .Y (n_15935));
INVX1 g68233(.A (n_15932), .Y (n_15931));
INVX1 g68235(.A (n_26882), .Y (n_15930));
INVX1 g68261(.A (n_15926), .Y (n_15927));
NOR2X1 g68273(.A (n_7315), .B (n_10603), .Y (n_15924));
NAND2X1 g68297(.A (n_11733), .B (n_9106), .Y (n_15923));
INVX1 g68299(.A (n_18268), .Y (n_15922));
OR2X1 g68303(.A (n_10268), .B (n_6534), .Y (n_18809));
NOR2X1 g68332(.A (n_12890), .B (n_9841), .Y (n_15920));
NAND2X1 g68349(.A (n_15919), .B (n_15918), .Y (n_17580));
INVX1 g68362(.A (n_14096), .Y (n_15917));
OR2X1 g68365(.A (n_9988), .B (n_20325), .Y (n_15916));
INVX1 g68376(.A (n_15913), .Y (n_15914));
NOR2X1 g68379(.A (n_11700), .B (n_14472), .Y (n_15912));
NAND2X1 g68383(.A (n_15909), .B (n_13744), .Y (n_15910));
NOR2X1 g68384(.A (n_10204), .B (n_11412), .Y (n_15908));
NAND2X1 g65377(.A (n_11980), .B (n_15902), .Y (n_15903));
NOR2X1 g68429(.A (n_11951), .B (n_29269), .Y (n_15901));
OR2X1 g68433(.A (n_12681), .B (n_16835), .Y (n_15900));
AOI21X1 g68454(.A0 (n_6170), .A1 (n_9838), .B0 (n_1547), .Y(n_15898));
NAND2X1 g68459(.A (n_11802), .B (n_18119), .Y (n_15897));
NAND2X1 g68463(.A (n_11676), .B (n_16434), .Y (n_15896));
NAND2X1 g68464(.A (n_11664), .B (n_15894), .Y (n_15895));
NAND2X1 g68473(.A (n_11666), .B (n_17260), .Y (n_15893));
NOR2X1 g68506(.A (n_9636), .B (n_9781), .Y (n_15892));
NAND2X1 g68512(.A (n_11860), .B (n_18087), .Y (n_15891));
NAND2X1 g68519(.A (n_11674), .B (n_27688), .Y (n_15890));
OAI21X1 g68541(.A0 (n_9588), .A1 (n_18266), .B0 (n_6815), .Y(n_15888));
NAND2X1 g65378(.A (n_8187), .B (n_15886), .Y (n_15887));
INVX1 g68559(.A (n_14025), .Y (n_25523));
NOR2X1 g68561(.A (n_5688), .B (n_11897), .Y (n_15884));
NOR2X1 g68582(.A (n_7875), .B (n_9754), .Y (n_15883));
NAND2X1 g68595(.A (n_9138), .B (n_13879), .Y (n_15882));
NAND2X1 g68596(.A (n_10278), .B (n_13745), .Y (n_15881));
NAND2X1 g68611(.A (n_11977), .B (n_26713), .Y (n_15880));
INVX1 g68628(.A (n_14003), .Y (n_15879));
AOI21X1 g68641(.A0 (n_4327), .A1 (n_3445), .B0 (n_12027), .Y(n_15878));
AOI21X1 g68645(.A0 (n_5273), .A1 (n_12019), .B0 (n_10882), .Y(n_15877));
NOR2X1 g68651(.A (n_10405), .B (n_15874), .Y (n_15875));
INVX1 g68655(.A (n_14000), .Y (n_15873));
NAND2X1 g68669(.A (n_11965), .B (n_8301), .Y (n_29404));
NAND2X1 g68674(.A (n_9051), .B (n_13765), .Y (n_15871));
OAI21X1 g68677(.A0 (n_7096), .A1 (n_29137), .B0 (n_4676), .Y(n_15870));
OAI21X1 g68680(.A0 (n_6730), .A1 (n_11996), .B0 (n_13037), .Y(n_15869));
AOI21X1 g68688(.A0 (n_4334), .A1 (n_13909), .B0 (n_3900), .Y(n_15868));
OAI21X1 g68699(.A0 (n_4893), .A1 (n_9646), .B0 (n_14667), .Y(n_15867));
AND2X1 g68722(.A (n_11735), .B (n_1365), .Y (n_15866));
AOI21X1 g62140(.A0 (n_9594), .A1 (n_15894), .B0 (n_9354), .Y(n_15865));
NAND2X1 g68774(.A (n_9820), .B (n_15863), .Y (n_15864));
AOI21X1 g62145(.A0 (n_11448), .A1 (n_11489), .B0 (n_9346), .Y(n_15862));
NAND2X1 g68783(.A (n_11817), .B (n_15860), .Y (n_15861));
NAND2X1 g68786(.A (n_10218), .B (n_15858), .Y (n_15859));
AOI21X1 g62154(.A0 (n_9562), .A1 (n_26270), .B0 (n_9279), .Y(n_15857));
XOR2X1 g68808(.A (n_1614), .B (n_11302), .Y (n_15856));
XOR2X1 g68809(.A (n_1409), .B (n_9602), .Y (n_15855));
XOR2X1 g68814(.A (n_1309), .B (n_9621), .Y (n_15854));
XOR2X1 g68815(.A (n_1165), .B (n_9625), .Y (n_15853));
XOR2X1 g68820(.A (n_993), .B (n_9617), .Y (n_15852));
INVX1 g68831(.A (n_15850), .Y (n_15851));
XOR2X1 g68835(.A (n_1109), .B (n_9612), .Y (n_15849));
INVX1 g68969(.A (n_15847), .Y (n_15848));
INVX1 g69040(.A (n_15846), .Y (n_18682));
AOI21X1 g62264(.A0 (n_9575), .A1 (n_12134), .B0 (n_10826), .Y(n_15845));
NAND3X1 g62271(.A (n_11065), .B (n_9615), .C (n_15837), .Y (n_15838));
NAND2X1 g62274(.A (n_11627), .B (n_1132), .Y (n_15836));
OR2X1 g69182(.A (n_9668), .B (n_26883), .Y (n_15835));
AOI21X1 g62308(.A0 (n_9566), .A1 (n_6185), .B0 (n_10995), .Y(n_15834));
OR2X1 g69328(.A (n_7840), .B (n_29256), .Y (n_15833));
OR2X1 g65376(.A (n_12882), .B (n_12986), .Y (n_15830));
NAND3X1 g62374(.A (n_16637), .B (n_11241), .C (n_11451), .Y(n_15829));
NAND4X1 g62379(.A (n_15825), .B (n_6756), .C (n_8064), .D (n_8703),.Y (n_15826));
OR2X1 g69863(.A (n_6563), .B (n_9783), .Y (n_15824));
OR2X1 g69882(.A (n_6952), .B (n_9084), .Y (n_15822));
AOI22X1 g62436(.A0 (n_9582), .A1 (n_12827), .B0 (n_8556), .B1(n_5887), .Y (n_15821));
NOR2X1 g62463(.A (n_11616), .B (n_19355), .Y (n_15819));
AOI21X1 g65375(.A0 (n_15055), .A1 (n_5513), .B0 (n_17411), .Y(n_15818));
INVX1 g70422(.A (n_15816), .Y (n_18716));
AOI21X1 g60090(.A0 (n_9648), .A1 (n_13728), .B0 (n_25052), .Y(n_15814));
NOR2X1 g70667(.A (n_15812), .B (n_11728), .Y (n_15813));
NAND4X1 g62661(.A (n_13122), .B (n_15462), .C (n_9528), .D (n_11626),.Y (n_15802));
NOR2X1 g70942(.A (n_15800), .B (n_15799), .Y (n_15801));
AOI21X1 g62671(.A0 (n_9584), .A1 (n_16988), .B0 (n_13006), .Y(n_15798));
AOI22X1 g62673(.A0 (n_11420), .A1 (n_9527), .B0 (n_12134), .B1(n_2716), .Y (n_15797));
AOI22X1 g62679(.A0 (n_11421), .A1 (n_16466), .B0 (n_7832), .B1(n_4965), .Y (n_15796));
NAND4X1 g62696(.A (n_13121), .B (n_15460), .C (n_10836), .D(n_13681), .Y (n_15795));
NAND4X1 g62753(.A (n_10769), .B (n_13763), .C (n_13114), .D(n_12828), .Y (n_15794));
AOI21X1 g62768(.A0 (n_9568), .A1 (n_29070), .B0 (n_11007), .Y(n_15791));
INVX1 g71495(.A (n_17888), .Y (n_17427));
NAND2X1 g71506(.A (n_11618), .B (n_5114), .Y (n_15789));
OAI21X1 g62812(.A0 (n_11146), .A1 (n_28220), .B0 (n_9410), .Y(n_15788));
OAI21X1 g62823(.A0 (n_11021), .A1 (n_8514), .B0 (n_15708), .Y(n_15786));
OAI21X1 g62832(.A0 (n_10927), .A1 (n_18552), .B0 (n_11489), .Y(n_15784));
NAND2X1 g71656(.A (n_9651), .B (n_11731), .Y (n_25526));
OAI21X1 g62835(.A0 (n_11115), .A1 (n_17472), .B0 (n_8708), .Y(n_15781));
OAI21X1 g62844(.A0 (n_10863), .A1 (n_7075), .B0 (n_13804), .Y(n_15780));
OAI21X1 g62846(.A0 (n_10998), .A1 (n_9872), .B0 (n_11400), .Y(n_29390));
NAND2X1 g62859(.A (n_13278), .B (n_15776), .Y (n_15777));
OAI21X1 g62876(.A0 (n_11019), .A1 (n_7177), .B0 (n_16787), .Y(n_15775));
NOR2X1 g71863(.A (n_29331), .B (n_21174), .Y (n_15774));
NAND2X1 g62889(.A (n_13196), .B (n_15986), .Y (n_15773));
OAI21X1 g62892(.A0 (n_10860), .A1 (n_6903), .B0 (n_16414), .Y(n_28837));
OAI21X1 g62899(.A0 (n_10901), .A1 (n_7242), .B0 (n_15039), .Y(n_15770));
OAI21X1 g62903(.A0 (n_10960), .A1 (n_6919), .B0 (n_9368), .Y(n_15768));
AOI21X1 g62904(.A0 (n_9901), .A1 (n_14956), .B0 (n_15766), .Y(n_15767));
AOI21X1 g62907(.A0 (n_8419), .A1 (n_16570), .B0 (n_310), .Y(n_15765));
INVX1 g71962(.A (n_15762), .Y (n_15764));
OAI21X1 g62931(.A0 (n_11132), .A1 (n_7369), .B0 (n_16480), .Y(n_15761));
OAI21X1 g62938(.A0 (n_10955), .A1 (n_10326), .B0 (n_9917), .Y(n_25768));
OAI21X1 g62941(.A0 (n_9254), .A1 (n_10550), .B0 (n_11400), .Y(n_15759));
OAI21X1 g62942(.A0 (n_9251), .A1 (n_10334), .B0 (n_17500), .Y(n_15758));
OAI21X1 g62947(.A0 (n_9245), .A1 (n_10331), .B0 (n_27688), .Y(n_15754));
OAI21X1 g62948(.A0 (n_11137), .A1 (n_9105), .B0 (n_16835), .Y(n_15752));
NAND3X1 g62949(.A (n_25791), .B (n_6623), .C (n_7702), .Y (n_15751));
NAND2X1 g62951(.A (n_11601), .B (n_9034), .Y (n_15750));
OAI21X1 g62962(.A0 (n_13646), .A1 (n_15748), .B0 (n_27111), .Y(n_29420));
NAND3X1 g62963(.A (n_5303), .B (n_11351), .C (n_6655), .Y (n_15745));
INVX1 g72246(.A (n_15741), .Y (n_15742));
OAI21X1 g62981(.A0 (n_13655), .A1 (n_15738), .B0 (n_2888), .Y(n_29312));
INVX1 g62995(.A (n_13786), .Y (n_15735));
OAI21X1 g63003(.A0 (n_8851), .A1 (n_17211), .B0 (n_624), .Y(n_15734));
INVX1 g63004(.A (n_13783), .Y (n_15733));
OAI21X1 g63006(.A0 (n_10253), .A1 (n_15180), .B0 (n_27128), .Y(n_15732));
OAI21X1 g63020(.A0 (n_10319), .A1 (n_13595), .B0 (n_2981), .Y(n_15731));
OAI21X1 g63024(.A0 (n_9364), .A1 (n_14321), .B0 (n_9264), .Y(n_15730));
OAI21X1 g63026(.A0 (n_11173), .A1 (n_12472), .B0 (n_28433), .Y(n_15729));
OAI21X1 g63027(.A0 (n_11145), .A1 (n_11088), .B0 (n_6534), .Y(n_15727));
OAI21X1 g63031(.A0 (n_10731), .A1 (n_9353), .B0 (n_13815), .Y(n_15726));
OAI21X1 g63036(.A0 (n_11071), .A1 (n_12613), .B0 (n_263), .Y(n_15725));
OAI21X1 g63038(.A0 (n_10761), .A1 (n_10968), .B0 (n_17500), .Y(n_15724));
OAI21X1 g63039(.A0 (n_10745), .A1 (n_27671), .B0 (n_17567), .Y(n_15723));
OAI21X1 g63041(.A0 (n_10744), .A1 (n_12495), .B0 (n_8708), .Y(n_15722));
OR2X1 g72477(.A (n_2289), .B (n_11650), .Y (n_15721));
NAND2X1 g72480(.A (n_11592), .B (n_5114), .Y (n_15720));
OAI21X1 g63047(.A0 (n_13609), .A1 (n_29129), .B0 (n_1424), .Y(n_25820));
OAI21X1 g63048(.A0 (n_10126), .A1 (n_5991), .B0 (n_14484), .Y(n_15717));
NAND3X1 g63065(.A (n_10622), .B (n_18335), .C (n_15714), .Y(n_15715));
OAI21X1 g63067(.A0 (n_10665), .A1 (n_14855), .B0 (n_15712), .Y(n_15713));
NAND2X1 g63069(.A (n_13249), .B (n_673), .Y (n_15711));
NAND2X1 g72583(.A (n_11606), .B (n_8520), .Y (n_15710));
OAI21X1 g63076(.A0 (n_10664), .A1 (n_7812), .B0 (n_15708), .Y(n_15709));
NAND2X1 g63094(.A (n_15678), .B (n_11362), .Y (n_15707));
AND2X1 g63096(.A (n_13531), .B (n_15705), .Y (n_15706));
NOR2X1 g63097(.A (n_14084), .B (n_11556), .Y (n_15704));
INVX1 g63107(.A (n_13761), .Y (n_15703));
AND2X1 g63109(.A (n_15701), .B (n_15700), .Y (n_15702));
AOI21X1 g63110(.A0 (n_11105), .A1 (n_12827), .B0 (n_7218), .Y(n_15699));
NAND3X1 g63111(.A (n_10245), .B (n_13567), .C (n_12070), .Y(n_15698));
OAI21X1 g63114(.A0 (n_9225), .A1 (n_11042), .B0 (n_20153), .Y(n_15697));
OAI21X1 g63130(.A0 (n_10656), .A1 (n_14734), .B0 (n_9527), .Y(n_15694));
NAND3X1 g63136(.A (n_9332), .B (n_15692), .C (n_18343), .Y (n_15693));
NAND2X1 g63137(.A (n_13231), .B (n_20010), .Y (n_15691));
OAI21X1 g63144(.A0 (n_15689), .A1 (n_15688), .B0 (n_15687), .Y(n_15690));
NOR2X1 g60320(.A (n_11609), .B (n_24548), .Y (n_15686));
NOR2X1 g60321(.A (n_11624), .B (n_24548), .Y (n_15685));
NAND3X1 g63156(.A (n_15682), .B (n_10069), .C (n_15681), .Y(n_15683));
OAI21X1 g63157(.A0 (n_10660), .A1 (n_13177), .B0 (n_14624), .Y(n_15680));
NAND2X1 g63171(.A (n_13214), .B (n_19310), .Y (n_15677));
AOI21X1 g63172(.A0 (n_11062), .A1 (n_15675), .B0 (n_15674), .Y(n_15676));
NAND3X1 g63178(.A (sa13[1] ), .B (n_10781), .C (n_16787), .Y(n_15673));
INVX1 g72950(.A (n_17596), .Y (n_15670));
OAI21X1 g63180(.A0 (n_10662), .A1 (n_11749), .B0 (n_17500), .Y(n_15669));
AND2X1 g63199(.A (n_11509), .B (n_15166), .Y (n_15663));
AOI21X1 g63214(.A0 (n_11075), .A1 (n_11365), .B0 (n_16480), .Y(n_15661));
NAND3X1 g63221(.A (n_15659), .B (n_14845), .C (n_9456), .Y (n_15660));
OAI21X1 g63223(.A0 (n_11152), .A1 (n_4397), .B0 (n_4582), .Y(n_15658));
NAND2X1 g63228(.A (n_15621), .B (n_11298), .Y (n_15657));
NAND2X1 g63230(.A (n_13208), .B (n_15655), .Y (n_15656));
NAND2X1 g63236(.A (n_11503), .B (n_29039), .Y (n_25547));
OAI21X1 g63242(.A0 (n_10443), .A1 (n_13018), .B0 (n_485), .Y(n_15652));
OAI21X1 g63249(.A0 (n_10659), .A1 (n_12106), .B0 (n_263), .Y(n_15650));
NAND3X1 g63256(.A (n_15648), .B (n_10222), .C (n_14770), .Y(n_15649));
NAND3X1 g63257(.A (n_10474), .B (n_15019), .C (n_12028), .Y(n_15647));
OAI21X1 g63280(.A0 (n_10658), .A1 (n_7820), .B0 (n_13804), .Y(n_29319));
OR2X1 g63281(.A (n_9558), .B (n_15644), .Y (n_15645));
NAND3X1 g63285(.A (n_10207), .B (n_15640), .C (n_13610), .Y(n_15641));
OAI21X1 g63290(.A0 (n_10657), .A1 (n_15636), .B0 (n_17377), .Y(n_15637));
OAI21X1 g63299(.A0 (n_10661), .A1 (n_12020), .B0 (n_28692), .Y(n_15635));
NAND2X1 g63302(.A (n_11476), .B (n_26798), .Y (n_15633));
NAND2X1 g63311(.A (n_15630), .B (n_27412), .Y (n_15631));
NAND3X1 g63316(.A (n_15628), .B (n_15627), .C (n_15626), .Y(n_15629));
OAI21X1 g63317(.A0 (n_10926), .A1 (n_5881), .B0 (n_11816), .Y(n_15625));
OAI21X1 g63332(.A0 (n_11184), .A1 (n_9101), .B0 (n_17567), .Y(n_15623));
NAND3X1 g63343(.A (n_20068), .B (n_10780), .C (n_11400), .Y(n_15620));
OAI21X1 g63346(.A0 (n_11095), .A1 (n_9058), .B0 (n_16466), .Y(n_15617));
NOR2X1 g63359(.A (n_15615), .B (n_20986), .Y (n_15616));
OAI21X1 g63362(.A0 (n_12544), .A1 (n_7357), .B0 (n_14807), .Y(n_15614));
OAI21X1 g63368(.A0 (n_12533), .A1 (n_10453), .B0 (n_15610), .Y(n_15611));
NAND3X1 g63370(.A (n_778), .B (n_10779), .C (n_13804), .Y (n_15609));
OAI21X1 g63376(.A0 (n_8001), .A1 (n_13380), .B0 (n_29065), .Y(n_15608));
NAND3X1 g63386(.A (n_10708), .B (n_11045), .C (n_15605), .Y(n_15606));
OAI21X1 g63394(.A0 (n_11168), .A1 (n_8788), .B0 (n_9410), .Y(n_15604));
OR2X1 g63397(.A (n_15612), .B (n_26903), .Y (n_15603));
NAND2X1 g63426(.A (n_14954), .B (n_27483), .Y (n_15602));
NAND3X1 g63444(.A (n_12202), .B (n_12312), .C (n_15600), .Y(n_15601));
NAND3X1 g63462(.A (n_16801), .B (n_15243), .C (n_8714), .Y (n_15599));
NAND2X1 g63468(.A (n_13145), .B (n_638), .Y (n_15598));
NAND3X1 g63472(.A (n_9186), .B (n_27496), .C (n_15596), .Y (n_15597));
OAI21X1 g63477(.A0 (n_10663), .A1 (n_6744), .B0 (n_27133), .Y(n_15595));
NAND2X1 g63481(.A (n_15615), .B (n_9000), .Y (n_15593));
AOI21X1 g63489(.A0 (n_10792), .A1 (n_10519), .B0 (n_9410), .Y(n_15592));
OAI21X1 g63492(.A0 (n_8797), .A1 (n_15590), .B0 (n_638), .Y(n_15591));
AOI21X1 g63502(.A0 (n_15588), .A1 (n_4124), .B0 (n_13229), .Y(n_15589));
NAND4X1 g63503(.A (n_15586), .B (n_7931), .C (n_14080), .D (n_15503),.Y (n_15587));
NAND3X1 g63510(.A (n_13265), .B (n_7143), .C (n_11329), .Y (n_15585));
NAND3X1 g63513(.A (n_12484), .B (n_7446), .C (n_15583), .Y (n_15584));
NAND2X1 g63515(.A (n_7263), .B (n_11597), .Y (n_15582));
NAND4X1 g63522(.A (n_15580), .B (n_8331), .C (n_14126), .D (n_15499),.Y (n_15581));
NAND3X1 g63540(.A (n_13429), .B (n_10839), .C (n_17754), .Y(n_15579));
AOI21X1 g63547(.A0 (n_10718), .A1 (n_14803), .B0 (n_19364), .Y(n_15578));
AOI21X1 g63549(.A0 (n_10727), .A1 (n_15575), .B0 (n_15574), .Y(n_15576));
NAND3X1 g63550(.A (n_6639), .B (n_11368), .C (n_9996), .Y (n_15573));
AOI21X1 g63552(.A0 (n_10712), .A1 (n_7732), .B0 (n_9410), .Y(n_15572));
AOI21X1 g63554(.A0 (n_10714), .A1 (n_13162), .B0 (n_28642), .Y(n_15571));
AOI21X1 g63559(.A0 (n_10706), .A1 (n_7717), .B0 (n_13326), .Y(n_15570));
AOI21X1 g63562(.A0 (n_11331), .A1 (n_28996), .B0 (n_15568), .Y(n_15569));
AOI21X1 g63564(.A0 (n_10713), .A1 (n_15566), .B0 (n_17500), .Y(n_15567));
INVX1 g63565(.A (n_13716), .Y (n_28260));
AOI21X1 g63570(.A0 (n_10719), .A1 (n_8922), .B0 (n_9819), .Y(n_15564));
AOI21X1 g63571(.A0 (n_10705), .A1 (n_14872), .B0 (n_12986), .Y(n_15563));
NAND2X1 g63585(.A (n_11555), .B (n_1196), .Y (n_15561));
AND2X1 g63594(.A (n_11564), .B (n_27604), .Y (n_15559));
OAI21X1 g63600(.A0 (n_12512), .A1 (n_1626), .B0 (n_9183), .Y(n_15558));
OAI21X1 g63618(.A0 (n_15556), .A1 (n_17912), .B0 (n_15555), .Y(n_15557));
NOR2X1 g63621(.A (n_11573), .B (n_12924), .Y (n_15554));
NAND3X1 g63639(.A (n_12717), .B (n_7519), .C (n_7741), .Y (n_15553));
NAND4X1 g63646(.A (n_13053), .B (n_9504), .C (n_7464), .D (n_8329),.Y (n_15552));
NAND3X1 g63647(.A (n_10091), .B (n_17024), .C (n_15469), .Y(n_15551));
OAI21X1 g63654(.A0 (n_9305), .A1 (n_15166), .B0 (n_12642), .Y(n_15549));
NAND3X1 g63657(.A (n_29336), .B (n_17021), .C (n_15463), .Y(n_15547));
NAND3X1 g63668(.A (n_7709), .B (n_15544), .C (n_15543), .Y (n_15545));
OAI21X1 g63677(.A0 (n_6166), .A1 (n_13402), .B0 (n_294), .Y(n_15542));
OAI21X1 g63714(.A0 (n_7486), .A1 (n_13445), .B0 (n_27747), .Y(n_15541));
NAND3X1 g63716(.A (n_8884), .B (n_15539), .C (n_15538), .Y (n_15540));
NAND3X1 g63719(.A (n_12498), .B (n_7385), .C (n_6928), .Y (n_15537));
NAND3X1 g63736(.A (n_12467), .B (n_7597), .C (n_7714), .Y (n_15536));
NAND4X1 g63746(.A (n_10883), .B (n_15534), .C (n_16049), .D(n_14467), .Y (n_15535));
AOI21X1 g63754(.A0 (n_14231), .A1 (n_13443), .B0 (n_16754), .Y(n_15533));
NAND3X1 g63762(.A (n_10018), .B (n_15531), .C (n_15488), .Y(n_15532));
OAI21X1 g63764(.A0 (n_5807), .A1 (n_13368), .B0 (n_2102), .Y(n_15530));
OAI21X1 g63767(.A0 (n_5857), .A1 (n_13559), .B0 (n_2805), .Y(n_15529));
OAI21X1 g63777(.A0 (n_26993), .A1 (n_13491), .B0 (n_399), .Y(n_15528));
OAI21X1 g63779(.A0 (n_9336), .A1 (n_13426), .B0 (n_523), .Y(n_15527));
OAI21X1 g63789(.A0 (n_28991), .A1 (n_14936), .B0 (n_826), .Y(n_15524));
NAND3X1 g63790(.A (n_11033), .B (n_11207), .C (n_8972), .Y (n_15523));
OAI21X1 g63793(.A0 (n_5895), .A1 (n_13564), .B0 (n_29266), .Y(n_15522));
AOI21X1 g63802(.A0 (n_6213), .A1 (n_19114), .B0 (n_11544), .Y(n_15519));
AOI22X1 g63807(.A0 (n_10677), .A1 (n_933), .B0 (n_5079), .B1(n_15516), .Y (n_15518));
NAND3X1 g63848(.A (n_12672), .B (n_15225), .C (n_14454), .Y(n_15515));
NAND3X1 g63855(.A (n_8872), .B (n_15513), .C (n_14120), .Y (n_15514));
NAND3X1 g63857(.A (n_12424), .B (n_15511), .C (n_12768), .Y(n_15512));
NAND3X1 g63866(.A (n_10377), .B (n_15509), .C (n_14574), .Y(n_29433));
AOI21X1 g63877(.A0 (n_9078), .A1 (n_15507), .B0 (n_11546), .Y(n_15508));
AOI21X1 g63885(.A0 (n_10721), .A1 (n_282), .B0 (n_12646), .Y(n_15506));
NAND3X1 g63886(.A (n_11049), .B (n_11362), .C (n_15503), .Y(n_15505));
AOI21X1 g63887(.A0 (n_9184), .A1 (n_124), .B0 (n_12737), .Y(n_15502));
NAND3X1 g63905(.A (n_10891), .B (n_11298), .C (n_15499), .Y(n_15501));
AOI21X1 g63907(.A0 (n_4194), .A1 (n_15497), .B0 (n_13127), .Y(n_15498));
NAND2X1 g63911(.A (n_13268), .B (n_18087), .Y (n_15496));
NAND2X1 g63913(.A (n_13280), .B (n_18102), .Y (n_15495));
AOI21X1 g63924(.A0 (n_5887), .A1 (n_4786), .B0 (n_11547), .Y(n_15492));
AOI22X1 g63934(.A0 (n_10743), .A1 (n_18266), .B0 (n_10147), .B1(n_9463), .Y (n_15491));
NOR2X1 g63937(.A (n_6992), .B (n_13288), .Y (n_15490));
MX2X1 g63939(.A (n_15488), .B (n_15487), .S0 (n_19364), .Y (n_15489));
AOI22X1 g63941(.A0 (n_10751), .A1 (n_19791), .B0 (n_14107), .B1(n_11435), .Y (n_15486));
NAND4X1 g63943(.A (n_17302), .B (n_15256), .C (n_11543), .D(n_17083), .Y (n_15485));
NAND3X1 g63968(.A (n_12421), .B (n_15028), .C (n_26372), .Y(n_15484));
AOI21X1 g63985(.A0 (n_10678), .A1 (n_13479), .B0 (n_15482), .Y(n_15483));
NOR2X1 g63988(.A (n_11332), .B (n_11515), .Y (n_15481));
XOR2X1 g76106(.A (text_in_r[12] ), .B (n_5306), .Y (n_15480));
NOR2X1 g63997(.A (n_11244), .B (n_13315), .Y (n_15479));
AOI21X1 g64000(.A0 (n_14128), .A1 (n_18320), .B0 (n_13302), .Y(n_15478));
XOR2X1 g76118(.A (text_in_r[26] ), .B (n_16978), .Y (n_15477));
NAND2X1 g64002(.A (n_12931), .B (n_13300), .Y (n_15475));
AOI21X1 g64004(.A0 (n_10728), .A1 (n_15473), .B0 (n_8389), .Y(n_15474));
AOI21X1 g64005(.A0 (n_10729), .A1 (n_3301), .B0 (n_10108), .Y(n_15472));
MX2X1 g64014(.A (n_15469), .B (n_15468), .S0 (n_13466), .Y (n_29413));
AOI22X1 g64015(.A0 (n_10935), .A1 (n_15655), .B0 (n_15465), .B1(n_9527), .Y (n_15466));
MX2X1 g64016(.A (n_15463), .B (n_15462), .S0 (n_4582), .Y (n_15464));
MX2X1 g64018(.A (n_11507), .B (n_15460), .S0 (n_13083), .Y (n_15461));
XOR2X1 g76188(.A (n_22750), .B (n_11312), .Y (n_15458));
OAI21X1 g64042(.A0 (n_10142), .A1 (n_9946), .B0 (n_28645), .Y(n_15457));
AOI21X1 g64048(.A0 (n_10552), .A1 (n_9073), .B0 (n_1057), .Y(n_15456));
OR2X1 g64049(.A (n_12219), .B (n_29102), .Y (n_28885));
OAI21X1 g64054(.A0 (n_10645), .A1 (n_4136), .B0 (n_17411), .Y(n_15453));
NAND4X1 g64062(.A (n_4743), .B (n_10812), .C (n_8349), .D (n_7783),.Y (n_15452));
NAND2X1 g64063(.A (n_12260), .B (n_12470), .Y (n_15451));
XOR2X1 g76259(.A (text_in_r[11] ), .B (n_3943), .Y (n_15450));
XOR2X1 g60721(.A (u0_rcon_1053), .B (n_1319), .Y (n_15448));
NOR2X1 g64069(.A (n_12242), .B (n_17571), .Y (n_15447));
INVX1 g64073(.A (n_13644), .Y (n_15445));
XOR2X1 g76284(.A (text_in_r[2] ), .B (n_16480), .Y (n_15444));
OAI21X1 g64083(.A0 (n_9805), .A1 (n_9716), .B0 (n_28645), .Y(n_15443));
AOI21X1 g64086(.A0 (n_9847), .A1 (n_9028), .B0 (n_28645), .Y(n_15442));
INVX1 g64087(.A (n_13636), .Y (n_15441));
INVX1 g64089(.A (n_13635), .Y (n_15440));
OAI21X1 g64094(.A0 (n_9739), .A1 (n_14531), .B0 (n_1424), .Y(n_15439));
AOI21X1 g64107(.A0 (n_7982), .A1 (n_16857), .B0 (n_20585), .Y(n_15437));
NOR2X1 g64123(.A (n_15435), .B (n_15894), .Y (n_16910));
NOR2X1 g64127(.A (n_18000), .B (n_27604), .Y (n_16908));
INVX1 g64133(.A (n_13613), .Y (n_21290));
INVX1 g64135(.A (n_13611), .Y (n_15434));
OR2X1 g64138(.A (n_16480), .B (n_15432), .Y (n_15433));
OR4X1 g64140(.A (n_17260), .B (n_29286), .C (n_8090), .D (n_6461), .Y(n_15431));
OR2X1 g64141(.A (n_16941), .B (n_12827), .Y (n_15430));
OR2X1 g64143(.A (n_16551), .B (n_13083), .Y (n_18388));
INVX1 g64144(.A (n_15427), .Y (n_15428));
OR2X1 g64152(.A (n_15425), .B (n_16466), .Y (n_15426));
INVX1 g64154(.A (n_15424), .Y (n_20634));
AND2X1 g64159(.A (n_15423), .B (n_11603), .Y (n_16904));
INVX1 g64165(.A (n_15420), .Y (n_15421));
NAND2X1 g64168(.A (n_15418), .B (n_16466), .Y (n_15419));
NAND2X1 g64172(.A (n_15415), .B (n_19791), .Y (n_15416));
OR2X1 g64175(.A (n_15414), .B (n_4582), .Y (n_18386));
INVX1 g64176(.A (n_13592), .Y (n_15413));
OR4X1 g64178(.A (n_15411), .B (n_11253), .C (n_26880), .D (n_7975),.Y (n_15412));
NOR2X1 g64185(.A (n_17972), .B (n_263), .Y (n_16897));
NOR2X1 g64188(.A (n_26614), .B (n_15039), .Y (n_18083));
OR2X1 g64190(.A (n_15404), .B (n_29048), .Y (n_18330));
OR2X1 g64191(.A (n_16674), .B (n_8708), .Y (n_15403));
AND2X1 g64193(.A (n_15180), .B (n_11576), .Y (n_15402));
NAND2X1 g64195(.A (n_12958), .B (n_29039), .Y (n_15400));
OR4X1 g64196(.A (n_28645), .B (n_8928), .C (n_28134), .D (n_8025), .Y(n_15399));
NAND2X1 g64197(.A (n_10824), .B (n_17567), .Y (n_15397));
INVX1 g64200(.A (n_13589), .Y (n_21659));
NAND3X1 g64203(.A (n_14807), .B (n_15395), .C (n_4898), .Y (n_15396));
NOR2X1 g64209(.A (n_15392), .B (n_11603), .Y (n_15393));
NOR2X1 g64212(.A (n_17982), .B (n_15574), .Y (n_16891));
INVX1 g64214(.A (n_15390), .Y (n_29396));
OR4X1 g64218(.A (n_263), .B (n_15388), .C (n_3834), .D (n_7937), .Y(n_15389));
NOR2X1 g64222(.A (n_16540), .B (n_15894), .Y (n_15387));
NAND2X1 g64223(.A (n_14696), .B (n_9527), .Y (n_15386));
NAND2X1 g64230(.A (n_12139), .B (n_21174), .Y (n_15384));
AOI21X1 g64232(.A0 (n_7293), .A1 (n_14415), .B0 (sa20[1] ), .Y(n_15381));
NAND2X1 g64236(.A (n_12132), .B (n_2681), .Y (n_15379));
NAND2X1 g64237(.A (n_12128), .B (n_129), .Y (n_15378));
AOI21X1 g64238(.A0 (n_8636), .A1 (n_14297), .B0 (sa23[1] ), .Y(n_15376));
NAND2X1 g64240(.A (n_12130), .B (n_27242), .Y (n_15374));
NAND2X1 g64242(.A (n_12141), .B (n_15371), .Y (n_15372));
AOI21X1 g64243(.A0 (n_9734), .A1 (n_14840), .B0 (n_20116), .Y(n_15370));
AOI21X1 g64249(.A0 (n_6246), .A1 (n_19297), .B0 (n_15894), .Y(n_15368));
AOI21X1 g64251(.A0 (n_7919), .A1 (n_19529), .B0 (n_9106), .Y(n_15367));
AOI21X1 g64254(.A0 (n_4270), .A1 (n_19499), .B0 (n_17411), .Y(n_15365));
NAND2X1 g64261(.A (n_12887), .B (n_15626), .Y (n_25581));
INVX1 g64266(.A (n_15362), .Y (n_15363));
NOR2X1 g64271(.A (n_15360), .B (n_9977), .Y (n_29196));
OR2X1 g64273(.A (n_15358), .B (n_27099), .Y (n_15359));
NOR2X1 g64275(.A (n_17211), .B (n_9140), .Y (n_15357));
NOR2X1 g64276(.A (n_12211), .B (n_15355), .Y (n_15356));
OR2X1 g64289(.A (n_12180), .B (n_19364), .Y (n_15354));
NAND3X1 g64290(.A (n_16187), .B (n_12680), .C (n_15352), .Y(n_15353));
NAND3X1 g64296(.A (n_8745), .B (n_5467), .C (n_15350), .Y (n_15351));
NAND2X1 g64297(.A (n_16334), .B (n_18353), .Y (n_15349));
OR2X1 g64299(.A (n_12861), .B (n_13815), .Y (n_15348));
NAND3X1 g64300(.A (n_11165), .B (n_5297), .C (n_12072), .Y (n_15347));
NAND2X1 g64301(.A (n_16532), .B (n_15345), .Y (n_15346));
AND2X1 g64305(.A (n_15435), .B (n_16540), .Y (n_15344));
NAND2X1 g64306(.A (n_10124), .B (n_15342), .Y (n_15343));
NAND2X1 g64307(.A (n_18587), .B (n_15340), .Y (n_15341));
OR2X1 g64312(.A (n_12197), .B (n_11261), .Y (n_15339));
NOR2X1 g64316(.A (n_17302), .B (n_13083), .Y (n_15337));
NAND2X1 g64322(.A (n_13282), .B (n_16568), .Y (n_15333));
NAND2X1 g64325(.A (n_27609), .B (n_14085), .Y (n_15332));
AOI21X1 g64326(.A0 (n_10164), .A1 (n_8487), .B0 (n_1547), .Y(n_15330));
AND2X1 g64327(.A (n_15583), .B (n_15328), .Y (n_15329));
NAND3X1 g64330(.A (n_8824), .B (n_6612), .C (n_15326), .Y (n_15327));
INVX1 g64332(.A (n_15324), .Y (n_15325));
NAND2X1 g64335(.A (n_15322), .B (n_8164), .Y (n_15323));
INVX1 g64336(.A (n_13549), .Y (n_15321));
NAND2X1 g64338(.A (n_15319), .B (n_29300), .Y (n_15320));
NAND2X1 g64340(.A (n_12886), .B (n_27688), .Y (n_16848));
NAND2X1 g64342(.A (n_18582), .B (n_16080), .Y (n_15318));
NAND4X1 g64344(.A (n_6363), .B (n_15316), .C (n_15315), .D (n_8933),.Y (n_15317));
NAND2X1 g64347(.A (n_15313), .B (n_18343), .Y (n_15314));
NAND3X1 g64350(.A (n_11563), .B (n_14130), .C (n_5586), .Y (n_15312));
NAND3X1 g64355(.A (n_6681), .B (n_4185), .C (n_15310), .Y (n_15311));
INVX1 g64357(.A (n_15308), .Y (n_15309));
NAND2X1 g64359(.A (n_18619), .B (n_14902), .Y (n_15307));
NAND2X1 g64361(.A (n_9356), .B (n_12320), .Y (n_15306));
NAND2X1 g64367(.A (n_15488), .B (n_15304), .Y (n_15305));
NAND2X1 g64369(.A (n_10043), .B (n_15302), .Y (n_15303));
NAND2X1 g64371(.A (n_12165), .B (n_21314), .Y (n_15301));
OR2X1 g64373(.A (n_18114), .B (n_12827), .Y (n_15300));
NAND2X1 g64377(.A (n_15299), .B (n_16978), .Y (n_18220));
NAND2X1 g64378(.A (n_13081), .B (n_11144), .Y (n_15298));
AOI21X1 g64381(.A0 (n_6990), .A1 (n_9688), .B0 (n_18617), .Y(n_15297));
OR2X1 g64384(.A (n_12156), .B (n_20587), .Y (n_15296));
NAND2X1 g64391(.A (n_12160), .B (n_196), .Y (n_15293));
NAND2X1 g64393(.A (n_12148), .B (n_16480), .Y (n_15292));
NAND2X1 g64396(.A (n_15291), .B (n_16480), .Y (n_16832));
INVX1 g64397(.A (n_15288), .Y (n_15289));
NAND2X1 g64406(.A (n_14709), .B (n_14526), .Y (n_15287));
NAND2X1 g64407(.A (n_15285), .B (n_18114), .Y (n_15286));
INVX1 g64408(.A (n_15283), .Y (n_15284));
NAND2X1 g64419(.A (n_13706), .B (n_15281), .Y (n_15282));
OR2X1 g64420(.A (n_12194), .B (n_14474), .Y (n_15280));
NAND2X1 g64421(.A (n_28829), .B (n_15278), .Y (n_15279));
NOR2X1 g64424(.A (n_12806), .B (n_15276), .Y (n_15277));
INVX1 g64432(.A (n_15274), .Y (n_15275));
NAND2X1 g64443(.A (n_8592), .B (n_15267), .Y (n_15268));
NAND2X1 g64454(.A (n_15266), .B (n_19445), .Y (n_18210));
INVX1 g64455(.A (n_13512), .Y (n_15265));
INVX1 g64458(.A (n_13511), .Y (n_25460));
INVX1 g64460(.A (n_15262), .Y (n_15263));
NAND2X1 g64468(.A (n_15260), .B (n_15259), .Y (n_15261));
AOI21X1 g64478(.A0 (n_9950), .A1 (n_7292), .B0 (n_18237), .Y(n_15258));
AND2X1 g64482(.A (n_15256), .B (n_13068), .Y (n_15257));
INVX1 g64484(.A (n_13502), .Y (n_18342));
NAND2X1 g64486(.A (n_15254), .B (n_5884), .Y (n_15255));
NOR2X1 g64491(.A (n_9356), .B (n_15894), .Y (n_15252));
AOI21X1 g64502(.A0 (n_6558), .A1 (n_8454), .B0 (n_29062), .Y(n_15250));
AND2X1 g64505(.A (n_16323), .B (n_11394), .Y (n_15248));
NAND3X1 g64506(.A (n_18046), .B (n_9361), .C (n_14512), .Y (n_15247));
NAND3X1 g64507(.A (n_16551), .B (n_10993), .C (n_15245), .Y(n_15246));
AND2X1 g64508(.A (n_17113), .B (n_15243), .Y (n_15244));
AND2X1 g64511(.A (n_15313), .B (n_11139), .Y (n_15242));
INVX1 g64513(.A (n_15240), .Y (n_15241));
NAND2X1 g64518(.A (n_15238), .B (n_15435), .Y (n_15239));
AND2X1 g64520(.A (n_12653), .B (n_16466), .Y (n_18375));
NAND2X1 g64522(.A (n_13036), .B (n_15236), .Y (n_15237));
NOR2X1 g64524(.A (n_15423), .B (n_8823), .Y (n_15235));
NOR2X1 g64526(.A (n_14573), .B (n_27373), .Y (n_15234));
OR2X1 g64529(.A (n_12250), .B (n_9410), .Y (n_15233));
OR2X1 g64530(.A (n_15230), .B (n_11603), .Y (n_18203));
INVX1 g64535(.A (n_13474), .Y (n_15232));
AND2X1 g64543(.A (n_15230), .B (n_15583), .Y (n_15231));
INVX1 g64546(.A (n_13463), .Y (n_15229));
AND2X1 g64550(.A (n_15886), .B (n_7354), .Y (n_15228));
NAND2X1 g64551(.A (n_14076), .B (n_18792), .Y (n_18360));
NAND2X1 g64555(.A (n_15226), .B (n_15225), .Y (n_15227));
NAND2X1 g64556(.A (n_16574), .B (n_18361), .Y (n_15224));
AND2X1 g64558(.A (n_12323), .B (n_15222), .Y (n_15223));
OR2X1 g64559(.A (n_27601), .B (n_18643), .Y (n_15221));
NOR2X1 g64563(.A (n_17757), .B (n_263), .Y (n_15219));
OR2X1 g64564(.A (n_12977), .B (n_17411), .Y (n_15218));
INVX1 g64568(.A (n_17161), .Y (n_15217));
AOI21X1 g64572(.A0 (n_9650), .A1 (n_8643), .B0 (n_19797), .Y(n_15216));
NAND2X1 g64576(.A (n_12817), .B (n_9527), .Y (n_16790));
INVX1 g64578(.A (n_28063), .Y (n_15214));
NAND3X1 g64580(.A (n_20078), .B (n_8607), .C (n_14493), .Y (n_15212));
INVX1 g64582(.A (n_15210), .Y (n_15211));
NOR2X1 g64584(.A (n_12960), .B (n_15291), .Y (n_15209));
NAND4X1 g64585(.A (n_15969), .B (n_12868), .C (n_14821), .D (n_8958),.Y (n_15208));
NOR2X1 g64587(.A (n_26470), .B (n_14643), .Y (n_15207));
NAND2X1 g64588(.A (n_8216), .B (n_16543), .Y (n_15206));
NAND3X1 g64592(.A (n_15659), .B (n_9574), .C (n_10827), .Y (n_15205));
NAND2X1 g64593(.A (n_16501), .B (n_16956), .Y (n_15204));
INVX1 g64594(.A (n_13451), .Y (n_28594));
NAND2X1 g64598(.A (n_28877), .B (n_14491), .Y (n_15200));
NAND2X1 g64599(.A (n_27645), .B (n_10687), .Y (n_15199));
AND2X1 g64605(.A (n_15196), .B (n_15195), .Y (n_15197));
NAND3X1 g64606(.A (n_27135), .B (n_4189), .C (n_27290), .Y (n_15194));
INVX1 g64609(.A (n_13444), .Y (n_15192));
NOR2X1 g64612(.A (n_7759), .B (n_16441), .Y (n_15189));
NAND4X1 g64617(.A (n_15187), .B (n_13722), .C (n_15186), .D (n_8976),.Y (n_15188));
NAND2X1 g64620(.A (n_16331), .B (n_8354), .Y (n_15185));
NAND3X1 g64622(.A (n_10827), .B (n_9456), .C (n_6578), .Y (n_15184));
NAND3X1 g64624(.A (n_9523), .B (n_8714), .C (n_4903), .Y (n_15183));
OR2X1 g64625(.A (n_27153), .B (n_11678), .Y (n_15182));
NOR2X1 g64629(.A (n_15180), .B (n_5755), .Y (n_15181));
NAND2X1 g64630(.A (n_18648), .B (n_14577), .Y (n_15179));
AND2X1 g64632(.A (n_14978), .B (n_15177), .Y (n_15178));
INVX1 g64638(.A (n_15175), .Y (n_15176));
NAND2X1 g64640(.A (n_15414), .B (n_13612), .Y (n_15174));
INVX1 g64641(.A (n_17157), .Y (n_15173));
NAND2X1 g64644(.A (n_20392), .B (n_12852), .Y (n_15172));
OR2X1 g64647(.A (n_15170), .B (n_14624), .Y (n_15171));
NAND2X1 g64649(.A (n_16637), .B (n_11186), .Y (n_15168));
AND2X1 g64652(.A (n_9451), .B (n_15166), .Y (n_16781));
NAND3X1 g64660(.A (n_27077), .B (n_14425), .C (n_13776), .Y(n_15165));
NAND2X1 g64661(.A (n_12308), .B (n_18205), .Y (n_15163));
OR2X1 g64665(.A (n_12152), .B (n_15039), .Y (n_15161));
NAND2X1 g64666(.A (n_15159), .B (n_13782), .Y (n_15160));
AND2X1 g64668(.A (n_12393), .B (n_8768), .Y (n_25707));
NOR2X1 g64669(.A (n_15156), .B (n_12895), .Y (n_15157));
NAND3X1 g64671(.A (n_26246), .B (n_14399), .C (n_19529), .Y(n_15154));
NOR2X1 g64675(.A (n_9144), .B (n_14567), .Y (n_15153));
OR2X1 g64676(.A (n_15151), .B (n_19857), .Y (n_15152));
NOR2X1 g64678(.A (n_9469), .B (n_16469), .Y (n_15149));
NOR2X1 g64682(.A (n_14227), .B (n_15147), .Y (n_28560));
NAND3X1 g64684(.A (n_15414), .B (n_7066), .C (n_17619), .Y (n_15146));
NAND2X1 g64688(.A (n_16426), .B (n_18286), .Y (n_15145));
INVX1 g64692(.A (n_15142), .Y (n_15143));
NAND2X1 g64696(.A (n_10048), .B (n_15140), .Y (n_15141));
NAND2X1 g64697(.A (n_9957), .B (n_16406), .Y (n_15139));
NAND2X1 g64700(.A (n_15137), .B (n_17972), .Y (n_15138));
NAND2X1 g64701(.A (n_11304), .B (n_15135), .Y (n_15136));
NOR2X1 g64706(.A (n_26958), .B (n_13928), .Y (n_25638));
NAND2X1 g64707(.A (n_14673), .B (n_15132), .Y (n_15133));
INVX1 g64708(.A (n_15130), .Y (n_15131));
NAND2X1 g64710(.A (n_18587), .B (n_26881), .Y (n_15129));
INVX1 g64726(.A (n_15127), .Y (n_15128));
NAND2X1 g64728(.A (n_12588), .B (n_28645), .Y (n_15126));
NAND2X1 g64731(.A (n_17197), .B (n_9435), .Y (n_15125));
NAND3X1 g64734(.A (n_13470), .B (n_14585), .C (n_26192), .Y(n_15124));
NAND3X1 g64736(.A (n_6956), .B (n_9142), .C (n_8268), .Y (n_15123));
NAND2X1 g64738(.A (n_15151), .B (n_15121), .Y (n_15122));
INVX1 g64745(.A (n_15118), .Y (n_15119));
AND2X1 g64756(.A (n_15116), .B (n_14464), .Y (n_15117));
NAND2X1 g64765(.A (n_12989), .B (n_15067), .Y (n_15115));
NAND2X1 g64766(.A (n_12125), .B (n_15113), .Y (n_15114));
AND2X1 g64770(.A (n_15111), .B (n_15942), .Y (n_15112));
NAND2X1 g64773(.A (n_12545), .B (n_15109), .Y (n_15110));
NAND2X1 g64777(.A (n_12984), .B (n_10701), .Y (n_15108));
NAND3X1 g64780(.A (n_12012), .B (n_4250), .C (n_12024), .Y (n_15107));
NAND4X1 g64781(.A (n_15105), .B (n_15104), .C (n_15103), .D (n_8914),.Y (n_15106));
AND2X1 g64783(.A (n_15101), .B (n_15100), .Y (n_15102));
NAND2X1 g64787(.A (n_15098), .B (n_8048), .Y (n_15099));
NAND2X1 g64788(.A (n_12534), .B (n_15648), .Y (n_28240));
NAND2X1 g64790(.A (n_13333), .B (n_15159), .Y (n_15096));
AND2X1 g64793(.A (n_12267), .B (n_14661), .Y (n_15095));
NAND2X1 g64794(.A (n_26380), .B (n_13190), .Y (n_15094));
NAND2X1 g64798(.A (n_15091), .B (n_15090), .Y (n_15092));
NAND3X1 g64799(.A (n_9142), .B (n_6621), .C (n_15087), .Y (n_15089));
NAND4X1 g64804(.A (n_15085), .B (n_13724), .C (n_14805), .D (n_8909),.Y (n_15086));
NAND2X1 g64805(.A (n_12698), .B (n_27099), .Y (n_15084));
NAND2X1 g64810(.A (n_9369), .B (n_17129), .Y (n_15082));
NAND2X1 g64820(.A (n_13416), .B (n_15404), .Y (n_15081));
NAND4X1 g64822(.A (n_14402), .B (n_18882), .C (n_15998), .D (n_5955),.Y (n_15080));
AND2X1 g64823(.A (n_16325), .B (n_11221), .Y (n_15079));
NAND2X1 g64824(.A (n_8525), .B (n_12610), .Y (n_15078));
NAND2X1 g64826(.A (n_15076), .B (n_14407), .Y (n_15077));
NAND2X1 g64828(.A (n_12462), .B (n_15074), .Y (n_15075));
NOR2X1 g64831(.A (n_12258), .B (n_15072), .Y (n_15073));
NAND2X1 g64835(.A (n_15070), .B (n_18050), .Y (n_15071));
NAND3X1 g64836(.A (n_15068), .B (n_14240), .C (n_15067), .Y(n_15069));
NAND2X1 g64841(.A (n_16398), .B (n_18051), .Y (n_15066));
NAND2X1 g64843(.A (n_8633), .B (n_15064), .Y (n_15065));
NAND3X1 g64853(.A (n_11696), .B (n_14340), .C (n_5591), .Y (n_15063));
AOI21X1 g64856(.A0 (n_8368), .A1 (n_5619), .B0 (n_9819), .Y(n_15062));
NAND2X1 g64858(.A (n_12983), .B (n_18168), .Y (n_15061));
NAND2X1 g64859(.A (n_10702), .B (n_18168), .Y (n_15059));
NAND2X1 g64861(.A (n_10158), .B (n_14945), .Y (n_15057));
NAND2X1 g64864(.A (n_15055), .B (n_16793), .Y (n_15056));
NAND3X1 g64867(.A (n_8462), .B (n_12340), .C (n_5685), .Y (n_15054));
NAND2X1 g64868(.A (n_10674), .B (n_4930), .Y (n_15053));
NAND2X1 g64869(.A (n_10697), .B (n_19857), .Y (n_15052));
NAND2X1 g64870(.A (n_26379), .B (n_19857), .Y (n_15051));
NAND2X1 g64871(.A (n_10940), .B (n_3168), .Y (n_15050));
NAND2X1 g64874(.A (n_12392), .B (n_19857), .Y (n_16720));
NAND2X1 g64880(.A (n_15048), .B (n_16787), .Y (n_17331));
AOI21X1 g64891(.A0 (n_6329), .A1 (n_9414), .B0 (n_27919), .Y(n_15047));
AND2X1 g64894(.A (n_15260), .B (n_15045), .Y (n_15046));
AND2X1 g64897(.A (n_11524), .B (n_15042), .Y (n_15044));
OAI21X1 g61012(.A0 (n_9228), .A1 (n_10999), .B0 (n_9249), .Y(n_15041));
INVX1 g64911(.A (n_13356), .Y (n_15040));
NAND2X1 g64917(.A (n_12272), .B (n_15039), .Y (n_19048));
INVX1 g64918(.A (n_13355), .Y (n_15038));
OR2X1 g64920(.A (n_13460), .B (n_4851), .Y (n_15037));
AOI21X1 g64922(.A0 (n_12376), .A1 (n_7383), .B0 (n_17567), .Y(n_15036));
AND2X1 g64923(.A (n_9550), .B (n_15034), .Y (n_15035));
AND2X1 g64924(.A (n_14996), .B (n_16678), .Y (n_15033));
NAND2X1 g64938(.A (n_15028), .B (n_10353), .Y (n_15029));
NAND2X1 g64939(.A (n_10668), .B (n_3168), .Y (n_15027));
NOR2X1 g64940(.A (n_7645), .B (n_15039), .Y (n_15026));
AOI21X1 g64942(.A0 (n_8587), .A1 (n_10676), .B0 (n_12760), .Y(n_15024));
INVX1 g64944(.A (n_13346), .Y (n_25823));
NOR2X1 g64947(.A (n_14745), .B (n_15021), .Y (n_28268));
NAND2X1 g64948(.A (n_12329), .B (n_15019), .Y (n_15020));
NAND2X1 g64949(.A (n_10121), .B (n_15513), .Y (n_15018));
NAND2X1 g64960(.A (n_18051), .B (n_12597), .Y (n_15016));
NAND2X1 g64961(.A (n_14819), .B (n_15014), .Y (n_15015));
AND2X1 g64966(.A (n_15012), .B (n_15011), .Y (n_15013));
NAND2X1 g64967(.A (n_15009), .B (n_10983), .Y (n_15010));
INVX1 g64970(.A (n_13337), .Y (n_15008));
INVX1 g64974(.A (n_13336), .Y (n_15007));
NOR2X1 g64985(.A (n_5198), .B (n_28123), .Y (n_15006));
NOR2X1 g64986(.A (n_12756), .B (n_12380), .Y (n_29322));
AND2X1 g64996(.A (n_11470), .B (n_15002), .Y (n_15003));
NAND2X1 g64998(.A (n_14958), .B (n_7201), .Y (n_15001));
INVX1 g65002(.A (n_13331), .Y (n_15000));
NAND2X1 g65008(.A (n_12560), .B (n_14765), .Y (n_14999));
NAND2X1 g65009(.A (n_14997), .B (n_14996), .Y (n_14998));
AOI21X1 g65010(.A0 (n_8866), .A1 (n_17356), .B0 (n_1424), .Y(n_14995));
INVX1 g65012(.A (n_13327), .Y (n_14993));
NAND2X1 g65016(.A (n_7046), .B (n_14991), .Y (n_14992));
NAND2X1 g65018(.A (n_10924), .B (n_19852), .Y (n_14990));
NAND2X1 g65021(.A (n_26375), .B (n_14988), .Y (n_14989));
NOR2X1 g65025(.A (n_10878), .B (n_14986), .Y (n_28879));
INVX1 g65026(.A (n_13319), .Y (n_14985));
NAND2X1 g65032(.A (n_10879), .B (n_16835), .Y (n_16647));
AOI21X1 g65040(.A0 (n_15961), .A1 (n_4689), .B0 (n_6885), .Y(n_14984));
NAND3X1 g65051(.A (n_26464), .B (n_6978), .C (n_14981), .Y (n_14983));
INVX1 g65053(.A (n_13314), .Y (n_14980));
NAND2X1 g65055(.A (n_14978), .B (n_10502), .Y (n_14979));
INVX1 g65066(.A (n_13311), .Y (n_14977));
NAND2X1 g65076(.A (n_13382), .B (n_14460), .Y (n_14976));
NOR2X1 g65085(.A (n_14364), .B (n_12476), .Y (n_14975));
NOR2X1 g65089(.A (n_12517), .B (n_12535), .Y (n_14974));
NAND2X1 g65097(.A (n_10818), .B (n_26276), .Y (n_16610));
OR2X1 g65101(.A (n_14969), .B (n_21174), .Y (n_14970));
NAND3X1 g65106(.A (n_13360), .B (n_8815), .C (n_3571), .Y (n_14967));
NAND3X1 g65108(.A (n_28619), .B (n_7548), .C (n_4407), .Y (n_14966));
NAND2X1 g65111(.A (n_12957), .B (n_14964), .Y (n_14965));
NAND2X1 g65114(.A (n_10692), .B (n_9819), .Y (n_14963));
NAND2X1 g65115(.A (n_9866), .B (n_14961), .Y (n_14962));
NAND2X1 g65121(.A (n_27137), .B (n_17414), .Y (n_14960));
NOR2X1 g65130(.A (n_6277), .B (n_14958), .Y (n_14959));
NAND3X1 g65132(.A (n_14956), .B (n_6926), .C (n_12486), .Y (n_14957));
INVX1 g65136(.A (n_14954), .Y (n_14955));
AND2X1 g65139(.A (n_10759), .B (n_17500), .Y (n_14953));
NAND2X1 g65143(.A (n_17821), .B (n_14951), .Y (n_14952));
NAND2X1 g65154(.A (n_14949), .B (n_6819), .Y (n_14950));
INVX1 g65163(.A (n_13285), .Y (n_14948));
NOR2X1 g65166(.A (n_14747), .B (n_15156), .Y (n_14947));
NAND2X1 g65169(.A (n_14945), .B (n_18335), .Y (n_14946));
NAND2X1 g65173(.A (n_18353), .B (n_8833), .Y (n_14944));
NAND2X1 g65175(.A (n_14942), .B (n_12075), .Y (n_14943));
NAND2X1 g65189(.A (n_12524), .B (n_9106), .Y (n_17189));
NAND2X1 g65192(.A (n_19450), .B (n_14940), .Y (n_14941));
AND2X1 g65195(.A (n_10735), .B (n_18320), .Y (n_14939));
NAND2X1 g65214(.A (n_19450), .B (n_10952), .Y (n_14938));
NAND2X1 g65216(.A (n_14936), .B (n_6534), .Y (n_14937));
AND2X1 g65218(.A (n_14934), .B (n_13066), .Y (n_14935));
NOR2X1 g65223(.A (n_6618), .B (n_12774), .Y (n_14933));
AOI21X1 g65226(.A0 (n_8557), .A1 (n_2480), .B0 (n_12827), .Y(n_14932));
NAND3X1 g65227(.A (n_8176), .B (n_4310), .C (n_14930), .Y (n_14931));
NAND2X1 g65228(.A (n_14928), .B (n_14927), .Y (n_14929));
NAND2X1 g65231(.A (n_13324), .B (n_16652), .Y (n_14926));
NAND2X1 g65236(.A (n_10703), .B (n_15712), .Y (n_14925));
NOR2X1 g65239(.A (n_10730), .B (n_13458), .Y (n_25628));
AND2X1 g65240(.A (n_14922), .B (n_11371), .Y (n_14923));
INVX1 g65241(.A (n_13276), .Y (n_14921));
NAND2X1 g65247(.A (n_12705), .B (n_18369), .Y (n_17295));
INVX1 g65248(.A (n_13275), .Y (n_25806));
NOR2X1 g65256(.A (n_12822), .B (n_12667), .Y (n_14919));
INVX1 g65258(.A (n_13274), .Y (n_14918));
NAND2X1 g65260(.A (n_11185), .B (n_6185), .Y (n_14917));
AND2X1 g65261(.A (n_14949), .B (n_17824), .Y (n_28558));
NAND3X1 g65262(.A (n_7489), .B (n_7786), .C (n_9037), .Y (n_14915));
NAND2X1 g65264(.A (n_10809), .B (n_19310), .Y (n_14914));
NAND2X1 g65268(.A (n_20910), .B (n_17567), .Y (n_19502));
OR2X1 g65269(.A (n_10683), .B (n_12298), .Y (n_14913));
INVX1 g65271(.A (n_13271), .Y (n_14912));
NAND2X1 g65275(.A (n_12833), .B (n_16466), .Y (n_17153));
INVX1 g65277(.A (n_13270), .Y (n_14911));
AND2X1 g65282(.A (n_28986), .B (n_14909), .Y (n_25838));
NAND2X1 g65285(.A (n_12938), .B (n_17912), .Y (n_14908));
OR2X1 g65288(.A (n_10802), .B (n_15688), .Y (n_14907));
NOR2X1 g65292(.A (n_13595), .B (n_6053), .Y (n_14905));
NOR2X1 g65294(.A (n_10486), .B (n_9278), .Y (n_14904));
NAND3X1 g65296(.A (n_29343), .B (n_14902), .C (n_3652), .Y (n_14903));
NAND2X1 g65303(.A (n_15469), .B (n_13213), .Y (n_14901));
OR2X1 g65310(.A (n_14899), .B (n_1196), .Y (n_14900));
NAND2X1 g65312(.A (n_27559), .B (n_29062), .Y (n_17046));
NAND2X1 g65314(.A (n_15509), .B (n_14574), .Y (n_14898));
NOR2X1 g65321(.A (n_10679), .B (n_10495), .Y (n_14897));
INVX1 g65325(.A (n_13261), .Y (n_14895));
NOR2X1 g65328(.A (n_9362), .B (n_10392), .Y (n_14894));
NOR2X1 g65330(.A (n_11162), .B (n_8848), .Y (n_14893));
NAND3X1 g65331(.A (n_14380), .B (n_8845), .C (n_26783), .Y (n_14892));
INVX1 g65333(.A (n_13258), .Y (n_25804));
NOR2X1 g65339(.A (n_10798), .B (n_7506), .Y (n_14890));
NAND3X1 g65343(.A (n_14377), .B (n_4224), .C (n_7207), .Y (n_14889));
NOR2X1 g65345(.A (n_9337), .B (n_11972), .Y (n_14888));
INVX1 g65346(.A (n_13255), .Y (n_14887));
INVX1 g65400(.A (n_13252), .Y (n_14886));
NOR2X1 g65361(.A (n_10855), .B (n_14535), .Y (n_14885));
INVX1 g65383(.A (n_11583), .Y (n_14884));
INVX1 g65405(.A (n_13248), .Y (n_14883));
INVX1 g65409(.A (n_13244), .Y (n_14882));
AOI21X1 g65411(.A0 (n_14880), .A1 (n_12291), .B0 (n_18440), .Y(n_14881));
AOI21X1 g65416(.A0 (n_1839), .A1 (n_14878), .B0 (n_13484), .Y(n_14879));
INVX1 g65420(.A (n_13240), .Y (n_14877));
INVX1 g65426(.A (n_13235), .Y (n_14875));
NAND2X1 g65428(.A (n_11113), .B (n_1424), .Y (n_14874));
AOI21X1 g65430(.A0 (n_5607), .A1 (n_14872), .B0 (n_19791), .Y(n_14873));
NAND3X1 g65432(.A (n_19226), .B (n_6024), .C (w3[17] ), .Y(n_14870));
AND2X1 g65434(.A (n_11012), .B (n_14868), .Y (n_14869));
OAI21X1 g65435(.A0 (n_11620), .A1 (n_14866), .B0 (n_13114), .Y(n_14867));
AOI21X1 g65437(.A0 (n_14864), .A1 (n_11745), .B0 (n_12986), .Y(n_14865));
NAND2X1 g65462(.A (n_11119), .B (n_27688), .Y (n_14863));
INVX1 g65476(.A (n_13225), .Y (n_14862));
INVX1 g65483(.A (n_13222), .Y (n_14861));
INVX1 g65487(.A (n_13221), .Y (n_14860));
NAND3X1 g65489(.A (n_16976), .B (n_14858), .C (n_663), .Y (n_14859));
INVX1 g65490(.A (n_13218), .Y (n_14857));
OAI21X1 g65492(.A0 (n_8115), .A1 (n_14855), .B0 (n_14854), .Y(n_14856));
INVX1 g65493(.A (n_13216), .Y (n_14853));
INVX1 g65516(.A (n_13210), .Y (n_14852));
AND2X1 g65518(.A (n_10737), .B (n_13466), .Y (n_14851));
AND2X1 g65523(.A (n_10828), .B (n_8217), .Y (n_14850));
NAND2X1 g65526(.A (n_11326), .B (n_5751), .Y (n_14849));
AOI21X1 g65529(.A0 (n_29337), .A1 (n_1626), .B0 (n_9459), .Y(n_14848));
NAND2X1 g65530(.A (n_9409), .B (n_14845), .Y (n_14846));
NAND2X1 g65556(.A (n_11014), .B (n_9106), .Y (n_14843));
AOI21X1 g65560(.A0 (n_14841), .A1 (n_14840), .B0 (n_2204), .Y(n_14842));
AND2X1 g65563(.A (n_10845), .B (n_29102), .Y (n_14839));
INVX1 g65569(.A (n_13201), .Y (n_14837));
NAND2X1 g65574(.A (n_10997), .B (n_13872), .Y (n_14836));
INVX1 g65592(.A (n_13198), .Y (n_14835));
NAND3X1 g65596(.A (n_10454), .B (n_13162), .C (n_9179), .Y (n_14834));
INVX1 g65601(.A (n_13194), .Y (n_14833));
OAI21X1 g65604(.A0 (n_14831), .A1 (n_12480), .B0 (n_1830), .Y(n_14832));
INVX1 g65605(.A (n_13193), .Y (n_29320));
NAND2X1 g65609(.A (n_10313), .B (n_14949), .Y (n_14828));
INVX1 g65610(.A (n_13191), .Y (n_14827));
INVX1 g65613(.A (n_13189), .Y (n_14826));
AOI21X1 g65618(.A0 (n_12206), .A1 (n_6753), .B0 (n_14026), .Y(n_14825));
NAND2X1 g65623(.A (n_9893), .B (n_14823), .Y (n_14824));
NAND3X1 g65627(.A (n_14821), .B (n_8267), .C (n_15002), .Y (n_14822));
NAND2X1 g65631(.A (n_9885), .B (n_14819), .Y (n_28310));
AOI21X1 g65635(.A0 (n_6773), .A1 (n_8925), .B0 (n_18320), .Y(n_14818));
AOI21X1 g65642(.A0 (n_14815), .A1 (n_13855), .B0 (n_28642), .Y(n_14816));
NAND2X1 g65644(.A (n_9810), .B (n_13408), .Y (n_14814));
NAND2X1 g65645(.A (n_8890), .B (n_19450), .Y (n_14813));
AOI21X1 g65646(.A0 (n_29190), .A1 (n_10691), .B0 (n_11998), .Y(n_14812));
NAND2X1 g65668(.A (n_11111), .B (n_16434), .Y (n_14809));
NAND2X1 g65671(.A (n_11109), .B (n_14807), .Y (n_14808));
NAND3X1 g65678(.A (n_14805), .B (n_14381), .C (n_13320), .Y(n_14806));
AOI21X1 g65685(.A0 (n_5652), .A1 (n_14803), .B0 (n_19364), .Y(n_14804));
NAND2X1 g65686(.A (n_10897), .B (n_29102), .Y (n_14802));
AOI21X1 g65694(.A0 (n_14800), .A1 (n_12138), .B0 (sa01[1] ), .Y(n_14801));
NOR2X1 g65695(.A (n_11085), .B (n_12980), .Y (n_14798));
AOI21X1 g65706(.A0 (n_8971), .A1 (n_7795), .B0 (n_12559), .Y(n_14797));
INVX1 g65708(.A (n_13167), .Y (n_14796));
INVX1 g65733(.A (n_13163), .Y (n_14795));
NAND2X1 g65738(.A (n_10842), .B (n_9276), .Y (n_14794));
NAND2X1 g65744(.A (n_10920), .B (n_11739), .Y (n_14793));
NAND2X1 g65746(.A (n_11032), .B (n_12568), .Y (n_14792));
INVX1 g65757(.A (n_13158), .Y (n_14791));
NAND4X1 g65761(.A (n_3212), .B (n_8523), .C (n_11097), .D (n_5288),.Y (n_14790));
INVX1 g65762(.A (n_13157), .Y (n_14789));
AOI21X1 g65766(.A0 (n_7489), .A1 (n_11249), .B0 (n_7614), .Y(n_14788));
NAND2X1 g65769(.A (n_10053), .B (n_13452), .Y (n_14787));
INVX1 g65770(.A (n_13154), .Y (n_14786));
NAND3X1 g65775(.A (n_9095), .B (n_14803), .C (n_11259), .Y (n_14785));
INVX1 g65776(.A (n_13153), .Y (n_14784));
INVX1 g65365(.A (n_13173), .Y (n_14783));
INVX1 g65786(.A (n_13147), .Y (n_14782));
AOI21X1 g65790(.A0 (n_9281), .A1 (n_1626), .B0 (n_13450), .Y(n_14781));
INVX1 g65795(.A (n_13144), .Y (n_14779));
NAND2X1 g65797(.A (n_10822), .B (n_15894), .Y (n_14778));
NAND2X1 g65810(.A (n_10783), .B (n_11810), .Y (n_14777));
NAND2X1 g65813(.A (n_10847), .B (n_12335), .Y (n_14776));
INVX1 g65815(.A (n_13138), .Y (n_14774));
INVX1 g65818(.A (n_13135), .Y (n_14773));
NAND2X1 g65820(.A (n_11155), .B (n_16434), .Y (n_14772));
NAND2X1 g65825(.A (n_10179), .B (n_14770), .Y (n_14771));
NAND2X1 g65828(.A (n_8472), .B (n_14961), .Y (n_14769));
AND2X1 g65830(.A (n_10778), .B (n_19170), .Y (n_14768));
AND2X1 g65836(.A (n_10776), .B (n_17459), .Y (n_14767));
NAND2X1 g65854(.A (n_10350), .B (n_14765), .Y (n_14766));
NAND2X1 g65855(.A (n_11337), .B (n_10133), .Y (n_14764));
OAI21X1 g65857(.A0 (n_3911), .A1 (n_8336), .B0 (n_13423), .Y(n_14763));
OAI21X1 g65858(.A0 (n_3350), .A1 (n_8286), .B0 (n_13575), .Y(n_14762));
OAI21X1 g65861(.A0 (n_3463), .A1 (n_8274), .B0 (n_16553), .Y(n_14760));
AOI21X1 g65863(.A0 (n_3489), .A1 (n_15588), .B0 (n_12825), .Y(n_14759));
AOI21X1 g65864(.A0 (n_2988), .A1 (n_14757), .B0 (n_12742), .Y(n_14758));
NOR2X1 g65865(.A (n_8177), .B (n_11103), .Y (n_14756));
NAND2X1 g65871(.A (n_10985), .B (n_15074), .Y (n_14755));
AOI21X1 g65879(.A0 (n_3945), .A1 (n_19226), .B0 (n_12296), .Y(n_14754));
MX2X1 g65880(.A (n_6276), .B (n_8106), .S0 (n_9819), .Y (n_14752));
MX2X1 g65883(.A (n_6935), .B (n_15256), .S0 (n_16466), .Y (n_14751));
MX2X1 g65884(.A (n_8576), .B (n_18116), .S0 (n_12827), .Y (n_14749));
AOI21X1 g65887(.A0 (n_14747), .A1 (n_4582), .B0 (n_9307), .Y(n_14748));
AOI21X1 g65890(.A0 (n_14745), .A1 (n_29074), .B0 (n_10903), .Y(n_14746));
OAI21X1 g65895(.A0 (n_12581), .A1 (n_8090), .B0 (n_9960), .Y(n_14744));
AOI21X1 g65896(.A0 (n_4106), .A1 (n_19226), .B0 (n_10670), .Y(n_14743));
OAI21X1 g65898(.A0 (n_8111), .A1 (n_13730), .B0 (n_14741), .Y(n_14742));
OAI21X1 g65906(.A0 (n_12629), .A1 (n_26880), .B0 (n_9784), .Y(n_14740));
AOI21X1 g65908(.A0 (n_3310), .A1 (n_14757), .B0 (n_10672), .Y(n_14739));
AOI21X1 g65914(.A0 (n_19110), .A1 (n_2400), .B0 (n_11339), .Y(n_14738));
AOI21X1 g65917(.A0 (n_29215), .A1 (n_16988), .B0 (n_11330), .Y(n_14737));
NAND2X1 g65925(.A (n_11336), .B (n_7831), .Y (n_17096));
AOI21X1 g65927(.A0 (n_13738), .A1 (n_15507), .B0 (n_11116), .Y(n_14736));
AOI22X1 g65932(.A0 (n_14734), .A1 (n_12134), .B0 (n_5417), .B1(n_8679), .Y (n_14735));
AOI21X1 g65947(.A0 (n_10232), .A1 (n_15610), .B0 (n_9054), .Y(n_14731));
AOI21X1 g65951(.A0 (n_9727), .A1 (n_11400), .B0 (n_7291), .Y(n_14730));
AOI21X1 g65952(.A0 (n_10012), .A1 (n_15708), .B0 (n_8812), .Y(n_14729));
AND2X1 g65964(.A (n_6844), .B (n_10088), .Y (n_14728));
AND2X1 g65965(.A (n_9863), .B (n_15674), .Y (n_14727));
AOI21X1 g65974(.A0 (n_6644), .A1 (n_14725), .B0 (n_9873), .Y(n_14726));
AND2X1 g65975(.A (n_9695), .B (n_6222), .Y (n_14724));
OR2X1 g65996(.A (n_15712), .B (n_14491), .Y (n_19097));
OR2X1 g66002(.A (n_15177), .B (n_17260), .Y (n_14723));
INVX2 g66005(.A (n_13095), .Y (n_16912));
NOR2X1 g66024(.A (n_19297), .B (n_15894), .Y (n_14721));
NAND2X1 g66035(.A (n_14700), .B (n_6534), .Y (n_14718));
AND2X1 g66059(.A (n_11842), .B (n_18266), .Y (n_16264));
NAND2X1 g66064(.A (n_14681), .B (n_29256), .Y (n_14714));
NOR2X1 g66071(.A (n_8167), .B (n_7598), .Y (n_14712));
INVX2 g66087(.A (n_13079), .Y (n_16893));
INVX1 g66117(.A (n_14707), .Y (n_14708));
INVX1 g66125(.A (n_17113), .Y (n_14706));
OR2X1 g66135(.A (n_15692), .B (n_13083), .Y (n_16810));
NAND2X1 g66137(.A (n_14704), .B (n_7410), .Y (n_14705));
NOR2X1 g66148(.A (n_8737), .B (n_11731), .Y (n_14702));
NAND2X1 g66152(.A (n_14700), .B (n_18237), .Y (n_14701));
INVX1 g66160(.A (n_14696), .Y (n_14697));
INVX1 g66173(.A (n_13062), .Y (n_18391));
NAND2X1 g66190(.A (n_13976), .B (n_15776), .Y (n_14694));
NAND2X1 g66202(.A (n_11854), .B (n_13466), .Y (n_14691));
NOR2X1 g66230(.A (n_29065), .B (n_8897), .Y (n_16251));
INVX1 g66238(.A (n_13044), .Y (n_14690));
NOR2X1 g66241(.A (n_263), .B (n_10493), .Y (n_14689));
INVX1 g66242(.A (n_16775), .Y (n_14687));
OR2X1 g66265(.A (n_9868), .B (n_12910), .Y (n_19095));
NAND2X1 g66295(.A (n_12986), .B (n_14681), .Y (n_14682));
INVX1 g66296(.A (n_17240), .Y (n_14680));
OR4X1 g66306(.A (n_9783), .B (n_5413), .C (n_28459), .D (n_6096), .Y(n_18826));
INVX1 g66330(.A (n_14677), .Y (n_14678));
NOR2X1 g66351(.A (n_19529), .B (n_20325), .Y (n_14676));
NOR2X1 g66355(.A (n_15894), .B (n_10467), .Y (n_14675));
INVX1 g66366(.A (n_14671), .Y (n_14672));
NOR2X1 g66370(.A (n_11805), .B (n_11400), .Y (n_14670));
INVX1 g66373(.A (n_13012), .Y (n_16765));
INVX1 g66377(.A (n_13010), .Y (n_16767));
INVX1 g66389(.A (n_13005), .Y (n_14669));
INVX1 g66408(.A (n_16670), .Y (n_14668));
NAND3X1 g66415(.A (n_28642), .B (n_14667), .C (n_8015), .Y (n_19638));
OR2X1 g66419(.A (n_17037), .B (n_28692), .Y (n_14666));
INVX1 g66450(.A (n_14661), .Y (n_14662));
INVX1 g66460(.A (n_12974), .Y (n_14660));
NOR2X1 g66465(.A (n_13383), .B (n_4689), .Y (n_14659));
OR2X1 g66477(.A (n_14657), .B (n_9106), .Y (n_14658));
INVX1 g66481(.A (n_14655), .Y (n_14656));
NOR2X1 g66490(.A (n_26469), .B (n_28680), .Y (n_14653));
NAND2X1 g66491(.A (n_14447), .B (n_11261), .Y (n_14652));
INVX1 g66503(.A (n_14649), .Y (n_14650));
NAND2X1 g66505(.A (n_14193), .B (n_1057), .Y (n_14648));
INVX1 g66521(.A (n_14647), .Y (n_17734));
INVX1 g66528(.A (n_14646), .Y (n_16210));
INVX1 g66533(.A (n_14643), .Y (n_14644));
INVX1 g66535(.A (n_14641), .Y (n_17929));
INVX1 g66536(.A (n_14641), .Y (n_14642));
NOR2X1 g66548(.A (n_8937), .B (n_8708), .Y (n_16207));
NAND2X1 g66567(.A (n_14186), .B (n_28133), .Y (n_14640));
INVX1 g66571(.A (n_14638), .Y (n_14639));
INVX1 g66576(.A (n_14636), .Y (n_14637));
INVX1 g66591(.A (n_14633), .Y (n_14635));
NAND2X1 g66594(.A (n_11778), .B (n_29048), .Y (n_29369));
OR4X1 g66603(.A (n_27688), .B (n_8452), .C (n_28459), .D (n_6096), .Y(n_16196));
NOR2X1 g66614(.A (n_10543), .B (n_14627), .Y (n_14628));
NOR2X1 g66617(.A (n_28680), .B (n_10438), .Y (n_14626));
OR2X1 g66618(.A (n_9875), .B (n_14624), .Y (n_14625));
INVX1 g66629(.A (n_12929), .Y (n_14623));
INVX1 g66662(.A (n_12919), .Y (n_18465));
NOR2X1 g66669(.A (n_14616), .B (n_17414), .Y (n_14617));
NOR2X1 g66681(.A (n_19499), .B (n_17500), .Y (n_14615));
NAND2X1 g66685(.A (n_9626), .B (n_27344), .Y (n_14613));
NAND2X1 g66686(.A (n_14704), .B (n_16466), .Y (n_14611));
NOR2X1 g66688(.A (n_10195), .B (n_17260), .Y (n_14610));
NOR2X1 g66690(.A (n_15045), .B (n_16787), .Y (n_14608));
NOR2X1 g66702(.A (n_8009), .B (n_14484), .Y (n_14607));
INVX1 g66710(.A (n_16559), .Y (n_14605));
INVX1 g66718(.A (n_14603), .Y (n_14604));
NAND3X1 g66723(.A (n_18237), .B (n_5104), .C (n_28611), .Y (n_18946));
NAND2X1 g66724(.A (n_14600), .B (n_263), .Y (n_14601));
NOR2X1 g66729(.A (n_14598), .B (n_7410), .Y (n_16176));
NAND2X1 g66743(.A (n_11762), .B (n_6219), .Y (n_16172));
NOR2X1 g66748(.A (n_10502), .B (n_1196), .Y (n_14597));
NAND2X1 g66749(.A (n_14141), .B (n_16434), .Y (n_14596));
INVX1 g66775(.A (n_12894), .Y (n_17844));
NOR2X1 g66779(.A (n_15011), .B (n_16414), .Y (n_14594));
OR2X1 g66783(.A (n_9956), .B (n_14592), .Y (n_14593));
NOR2X1 g66799(.A (n_15042), .B (n_14589), .Y (n_14590));
INVX1 g66806(.A (n_14587), .Y (n_16159));
NOR2X1 g66817(.A (n_14348), .B (n_14585), .Y (n_17147));
NAND2X1 g66829(.A (n_10339), .B (n_7203), .Y (n_14583));
INVX1 g66831(.A (n_15360), .Y (n_14582));
INVX1 g66837(.A (n_12884), .Y (n_14581));
OR2X1 g66841(.A (n_14704), .B (n_6135), .Y (n_14580));
NOR2X1 g66851(.A (n_15039), .B (n_9142), .Y (n_14579));
AND2X1 g66878(.A (n_10104), .B (n_14574), .Y (n_14575));
OR2X1 g66887(.A (n_9116), .B (n_15968), .Y (n_16861));
NOR2X1 g66890(.A (n_14571), .B (n_13834), .Y (n_16144));
NAND2X1 g66897(.A (n_16825), .B (n_13260), .Y (n_14570));
OR2X1 g66898(.A (n_9040), .B (n_9410), .Y (n_14569));
NAND2X1 g66906(.A (n_5527), .B (n_17325), .Y (n_14568));
NOR2X1 g66919(.A (n_2654), .B (n_16416), .Y (n_19287));
INVX1 g66928(.A (n_14564), .Y (n_14565));
NAND2X1 g66932(.A (n_16485), .B (n_17621), .Y (n_16137));
INVX1 g66935(.A (n_14561), .Y (n_14562));
NAND2X1 g66937(.A (n_14442), .B (n_11008), .Y (n_16797));
INVX1 g66938(.A (n_14559), .Y (n_14560));
NAND2X1 g66941(.A (n_10556), .B (n_29228), .Y (n_14558));
NAND2X1 g66949(.A (n_14556), .B (n_9056), .Y (n_14557));
OR2X1 g66951(.A (n_11543), .B (n_7410), .Y (n_14555));
NOR2X1 g66958(.A (n_8515), .B (n_15708), .Y (n_16132));
NAND2X1 g66959(.A (n_14284), .B (n_10734), .Y (n_14554));
OR2X1 g66971(.A (n_11029), .B (n_16787), .Y (n_14553));
NAND2X1 g66973(.A (n_8515), .B (n_9085), .Y (n_14551));
NAND2X1 g66978(.A (n_10631), .B (n_14548), .Y (n_14549));
NOR2X1 g66985(.A (n_10337), .B (n_14546), .Y (n_14547));
NAND2X1 g66986(.A (n_12362), .B (n_17813), .Y (n_16864));
NAND2X1 g66987(.A (n_27309), .B (n_7063), .Y (n_14545));
INVX1 g66990(.A (n_17292), .Y (n_16128));
NOR2X1 g66995(.A (n_17260), .B (n_10850), .Y (n_16126));
NAND2X1 g67003(.A (n_5006), .B (n_16434), .Y (n_14544));
NOR2X1 g67008(.A (n_12068), .B (n_9355), .Y (n_14543));
INVX1 g67019(.A (n_12818), .Y (n_16121));
INVX1 g67026(.A (n_12816), .Y (n_16119));
NAND2X1 g67038(.A (n_6523), .B (n_8167), .Y (n_14540));
NAND2X1 g67040(.A (n_14537), .B (n_4427), .Y (n_14538));
OR2X1 g67047(.A (n_14535), .B (n_14534), .Y (n_14536));
NAND2X1 g67056(.A (n_4619), .B (n_26798), .Y (n_14533));
OAI21X1 g67073(.A0 (n_8021), .A1 (n_14531), .B0 (n_15776), .Y(n_14532));
OR2X1 g67074(.A (n_14528), .B (n_14681), .Y (n_14529));
AND2X1 g67083(.A (n_9697), .B (n_17864), .Y (n_14527));
OR2X1 g67084(.A (n_14526), .B (n_29228), .Y (n_18038));
NAND2X1 g67085(.A (n_5058), .B (n_10104), .Y (n_14525));
NAND2X1 g67091(.A (n_9000), .B (n_14523), .Y (n_14524));
AND2X1 g67100(.A (n_16049), .B (n_14521), .Y (n_14522));
NOR2X1 g67101(.A (n_7849), .B (n_11177), .Y (n_14520));
NOR2X1 g67104(.A (n_11367), .B (n_4969), .Y (n_14519));
NAND2X1 g67106(.A (n_14517), .B (n_11821), .Y (n_14518));
NAND2X1 g67107(.A (n_11884), .B (n_11261), .Y (n_14516));
NAND2X1 g67115(.A (n_14513), .B (n_11932), .Y (n_14514));
OR2X1 g67117(.A (n_14928), .B (n_13490), .Y (n_16111));
OR2X1 g67120(.A (n_14512), .B (n_7410), .Y (n_16817));
NAND2X1 g67138(.A (n_14577), .B (n_3699), .Y (n_14511));
NOR2X1 g67147(.A (n_7220), .B (n_5558), .Y (n_16108));
OR2X1 g67148(.A (n_14510), .B (n_7410), .Y (n_16906));
NAND2X1 g67167(.A (n_6874), .B (n_15605), .Y (n_14508));
NOR2X1 g67172(.A (n_3198), .B (n_14542), .Y (n_19321));
OR2X1 g67195(.A (n_11386), .B (n_10562), .Y (n_14505));
NAND2X1 g67202(.A (n_10038), .B (n_27688), .Y (n_14502));
NAND2X1 g67206(.A (n_14500), .B (n_12306), .Y (n_14501));
NOR2X1 g67207(.A (n_11886), .B (n_13609), .Y (n_14499));
INVX1 g67209(.A (n_12730), .Y (n_14498));
AOI21X1 g67216(.A0 (n_6250), .A1 (n_3827), .B0 (n_9878), .Y(n_14497));
NAND2X1 g67229(.A (n_5525), .B (n_29343), .Y (n_14495));
NOR2X1 g67231(.A (n_14493), .B (n_11312), .Y (n_16844));
AND2X1 g67235(.A (n_5264), .B (n_14491), .Y (n_14492));
INVX1 g67236(.A (n_14489), .Y (n_14490));
NOR2X1 g67238(.A (n_26492), .B (n_14592), .Y (n_14488));
INVX1 g67244(.A (n_12712), .Y (n_14487));
OR2X1 g67246(.A (n_7574), .B (n_11307), .Y (n_16889));
NAND2X1 g67253(.A (n_27596), .B (n_9170), .Y (n_17904));
OR2X1 g67254(.A (n_8884), .B (n_14484), .Y (n_14486));
AND2X1 g67256(.A (n_14482), .B (n_12249), .Y (n_14483));
OR2X1 g67257(.A (n_10921), .B (n_15039), .Y (n_14481));
NAND2X1 g67260(.A (n_6042), .B (n_14478), .Y (n_14479));
NAND2X1 g67261(.A (n_19842), .B (n_26726), .Y (n_14477));
OR2X1 g67274(.A (n_13466), .B (n_9524), .Y (n_16084));
OR2X1 g67283(.A (n_14093), .B (n_14474), .Y (n_14475));
OR2X1 g67287(.A (n_14392), .B (n_28680), .Y (n_14473));
INVX1 g72980(.A (n_14472), .Y (n_15667));
AND2X1 g67294(.A (n_7632), .B (n_15894), .Y (n_14471));
NAND2X1 g67301(.A (n_14463), .B (n_9034), .Y (n_14470));
NAND2X1 g67302(.A (n_8937), .B (n_10488), .Y (n_14469));
NAND2X1 g67303(.A (n_14467), .B (n_14216), .Y (n_14468));
NOR2X1 g67307(.A (n_6889), .B (n_14464), .Y (n_14466));
NOR2X1 g67310(.A (n_14463), .B (n_11576), .Y (n_16078));
NAND2X1 g67314(.A (n_26464), .B (n_14314), .Y (n_14462));
NAND2X1 g67322(.A (n_4225), .B (n_14460), .Y (n_14461));
INVX1 g67331(.A (n_15638), .Y (n_14459));
OR2X1 g67339(.A (n_10909), .B (n_12896), .Y (n_14458));
NAND2X1 g67341(.A (n_14454), .B (n_6363), .Y (n_14455));
NOR2X1 g67344(.A (n_8165), .B (n_14099), .Y (n_14452));
INVX1 g67346(.A (n_14450), .Y (n_14451));
NOR2X1 g67353(.A (n_14928), .B (n_3630), .Y (n_16074));
NAND2X1 g67358(.A (n_14447), .B (n_1358), .Y (n_14448));
NOR2X1 g67371(.A (n_12081), .B (n_9291), .Y (n_14444));
NAND2X1 g67372(.A (n_14418), .B (n_14442), .Y (n_14443));
NAND2X1 g67374(.A (n_12036), .B (n_16434), .Y (n_17879));
NAND2X1 g67378(.A (n_8675), .B (n_9208), .Y (n_16785));
NOR2X1 g67381(.A (n_6363), .B (n_11835), .Y (n_14440));
INVX1 g67400(.A (n_12669), .Y (n_16059));
NAND2X1 g67407(.A (n_14028), .B (n_14208), .Y (n_14439));
AND2X1 g67414(.A (n_15177), .B (n_14526), .Y (n_14438));
NAND2X1 g67420(.A (n_15628), .B (n_15011), .Y (n_16057));
INVX1 g67423(.A (n_14437), .Y (n_16730));
OR2X1 g67426(.A (n_7309), .B (n_5817), .Y (n_16902));
AND2X1 g67427(.A (n_10638), .B (n_8666), .Y (n_14436));
NAND2X1 g67428(.A (n_14009), .B (n_5761), .Y (n_14435));
NAND2X1 g67431(.A (n_14433), .B (n_13418), .Y (n_14434));
NAND2X1 g67437(.A (n_11642), .B (n_12063), .Y (n_14430));
NAND2X1 g67439(.A (n_4260), .B (n_11808), .Y (n_14429));
NAND2X1 g65380(.A (n_11171), .B (n_12986), .Y (n_14428));
NOR2X1 g67458(.A (n_6028), .B (n_6846), .Y (n_14427));
NAND2X1 g67464(.A (n_14078), .B (n_14425), .Y (n_14426));
OR2X1 g67465(.A (n_12383), .B (n_8928), .Y (n_14424));
NAND2X1 g67467(.A (n_11362), .B (n_17325), .Y (n_14422));
NAND2X1 g67471(.A (n_12546), .B (n_16857), .Y (n_14421));
AND2X1 g67480(.A (n_9711), .B (n_13318), .Y (n_14420));
NAND2X1 g67481(.A (n_14418), .B (n_7573), .Y (n_14419));
NOR2X1 g67482(.A (n_10507), .B (n_4539), .Y (n_14417));
NAND2X1 g67484(.A (n_7110), .B (n_14415), .Y (n_14416));
NAND2X1 g67488(.A (n_14413), .B (n_12870), .Y (n_14414));
NOR2X1 g67502(.A (n_5709), .B (n_9911), .Y (n_14412));
OR2X1 g67518(.A (n_14521), .B (n_11253), .Y (n_18043));
AND2X1 g67528(.A (n_10638), .B (n_9040), .Y (n_14409));
OR2X1 g67531(.A (n_10434), .B (n_15388), .Y (n_16772));
AND2X1 g67533(.A (n_17037), .B (n_14407), .Y (n_14408));
NAND2X1 g67534(.A (n_14405), .B (n_3206), .Y (n_14406));
NAND2X1 g67541(.A (n_12172), .B (n_14402), .Y (n_14403));
NAND2X1 g67546(.A (n_11292), .B (n_8944), .Y (n_14401));
NOR2X1 g67549(.A (n_10436), .B (n_11936), .Y (n_14400));
NAND2X1 g67553(.A (n_14399), .B (n_15042), .Y (n_16044));
NAND2X1 g67557(.A (n_15534), .B (n_13257), .Y (n_14398));
NOR2X1 g67558(.A (n_5808), .B (n_6843), .Y (n_14397));
INVX1 g67559(.A (n_12598), .Y (n_14396));
NAND2X1 g67561(.A (n_14418), .B (n_5953), .Y (n_14395));
NAND2X1 g67563(.A (n_14393), .B (n_14392), .Y (n_14394));
AND2X1 g67565(.A (n_14390), .B (n_8454), .Y (n_14391));
NAND2X1 g67566(.A (n_11920), .B (n_28642), .Y (n_14388));
NAND4X1 g67572(.A (n_14386), .B (n_13183), .C (n_6579), .D (n_3557),.Y (n_14387));
OR2X1 g67575(.A (n_14384), .B (n_13318), .Y (n_14385));
NAND2X1 g67576(.A (n_7971), .B (n_11259), .Y (n_14383));
NAND2X1 g67578(.A (n_14381), .B (n_14380), .Y (n_14382));
NAND2X1 g67581(.A (n_6496), .B (n_13550), .Y (n_14379));
NAND2X1 g67583(.A (n_14377), .B (n_13192), .Y (n_14378));
NAND2X1 g67595(.A (n_28042), .B (n_8371), .Y (n_14376));
OR2X1 g67597(.A (n_7418), .B (n_8815), .Y (n_14374));
INVX1 g67610(.A (n_14372), .Y (n_16034));
INVX1 g67614(.A (n_14370), .Y (n_14371));
NAND2X1 g67618(.A (n_5521), .B (n_10417), .Y (n_14369));
INVX1 g67620(.A (n_14367), .Y (n_14368));
NAND3X1 g67622(.A (n_7089), .B (n_16754), .C (n_129), .Y (n_14366));
NOR2X1 g67630(.A (n_12013), .B (n_14364), .Y (n_14365));
AND2X1 g67634(.A (n_14362), .B (n_14361), .Y (n_25679));
AND2X1 g67638(.A (n_16390), .B (n_14571), .Y (n_14360));
NAND2X1 g67644(.A (n_9894), .B (n_27779), .Y (n_14357));
NOR2X1 g67645(.A (n_10156), .B (n_4460), .Y (n_14356));
INVX1 g67650(.A (n_14353), .Y (n_14354));
NAND2X1 g67655(.A (n_11967), .B (n_13606), .Y (n_14351));
AND2X1 g67657(.A (n_9717), .B (n_28692), .Y (n_14350));
NOR2X1 g67665(.A (n_7498), .B (n_14405), .Y (n_16030));
NOR2X1 g67669(.A (n_14348), .B (n_10687), .Y (n_14349));
AND2X1 g67677(.A (n_11984), .B (n_7437), .Y (n_14346));
NAND2X1 g67690(.A (n_14344), .B (n_14343), .Y (n_14345));
OR2X1 g67691(.A (n_8784), .B (n_8708), .Y (n_14342));
NAND2X1 g67695(.A (n_14340), .B (n_12024), .Y (n_14341));
NAND2X1 g67707(.A (n_14337), .B (n_14336), .Y (n_14338));
NOR2X1 g67715(.A (n_19857), .B (n_8768), .Y (n_16023));
NAND2X1 g67719(.A (n_12399), .B (n_13895), .Y (n_14334));
NAND2X1 g67721(.A (n_10110), .B (n_19830), .Y (n_14333));
NOR2X1 g67722(.A (n_3021), .B (n_9127), .Y (n_19850));
NAND2X1 g67724(.A (n_8959), .B (n_10389), .Y (n_14332));
NAND2X1 g67726(.A (n_8768), .B (n_14330), .Y (n_14331));
NOR2X1 g67732(.A (n_1746), .B (n_11833), .Y (n_14329));
INVX1 g67735(.A (n_14327), .Y (n_14328));
NOR2X1 g67743(.A (n_8466), .B (n_17414), .Y (n_16017));
NAND2X1 g67746(.A (n_14325), .B (n_14324), .Y (n_14326));
NAND2X1 g67749(.A (n_16351), .B (n_14616), .Y (n_16013));
NAND2X1 g67751(.A (n_10341), .B (n_16895), .Y (n_14323));
INVX1 g67754(.A (n_16639), .Y (n_17692));
NAND2X1 g67756(.A (n_14321), .B (n_5558), .Y (n_14322));
NOR2X1 g67762(.A (n_15411), .B (n_11008), .Y (n_16009));
NOR2X1 g67764(.A (n_14319), .B (n_14246), .Y (n_14320));
NAND2X1 g67766(.A (n_10531), .B (n_8452), .Y (n_14318));
NOR2X1 g67770(.A (n_7531), .B (n_7410), .Y (n_14317));
NOR2X1 g67771(.A (n_13026), .B (n_7925), .Y (n_14316));
NAND2X1 g67773(.A (n_7662), .B (n_14314), .Y (n_14315));
NAND2X1 g67775(.A (n_27596), .B (n_17377), .Y (n_16738));
NOR2X1 g67778(.A (n_27744), .B (n_9084), .Y (n_14313));
NAND2X1 g67780(.A (n_14309), .B (n_14308), .Y (n_14310));
NOR2X1 g67787(.A (n_11799), .B (n_8038), .Y (n_14307));
NOR2X1 g67789(.A (n_14407), .B (n_8928), .Y (n_14306));
NAND2X1 g67795(.A (n_14815), .B (n_17037), .Y (n_16003));
NAND2X1 g67796(.A (n_27145), .B (n_17414), .Y (n_14304));
NAND2X1 g67797(.A (n_4220), .B (n_8730), .Y (n_14303));
NOR2X1 g67800(.A (n_10957), .B (n_12298), .Y (n_14301));
NOR2X1 g67804(.A (n_7550), .B (n_10395), .Y (n_14299));
NAND2X1 g67806(.A (n_15395), .B (n_26276), .Y (n_20438));
NAND2X1 g67810(.A (n_8621), .B (n_14297), .Y (n_14298));
NAND2X1 g67813(.A (n_6645), .B (n_8298), .Y (n_14296));
OR2X1 g67814(.A (n_14308), .B (n_8637), .Y (n_14295));
NAND2X1 g67818(.A (n_14805), .B (n_14377), .Y (n_14294));
AND2X1 g67819(.A (n_9709), .B (n_15610), .Y (n_14293));
NOR2X1 g65362(.A (n_10823), .B (n_9045), .Y (n_14292));
NAND2X1 g67822(.A (n_14290), .B (n_10127), .Y (n_14291));
NAND2X1 g67823(.A (n_8003), .B (n_11998), .Y (n_14289));
NAND2X1 g67831(.A (n_8466), .B (n_14286), .Y (n_14288));
AND2X1 g67832(.A (n_10311), .B (n_14284), .Y (n_14285));
NAND2X1 g67837(.A (n_6556), .B (n_8511), .Y (n_14283));
NOR2X1 g67839(.A (n_12591), .B (n_9835), .Y (n_14281));
NAND2X1 g67852(.A (n_5178), .B (n_8944), .Y (n_14279));
NAND2X1 g67856(.A (n_4243), .B (n_9565), .Y (n_14276));
AND2X1 g67859(.A (n_14274), .B (n_6446), .Y (n_14275));
AND2X1 g67860(.A (n_3261), .B (n_14272), .Y (n_14273));
NOR2X1 g67865(.A (n_28041), .B (n_14624), .Y (n_14271));
NAND2X1 g67869(.A (n_9981), .B (n_15708), .Y (n_14270));
NAND2X1 g67872(.A (n_14880), .B (n_15045), .Y (n_15992));
NAND2X1 g67874(.A (n_14268), .B (n_11449), .Y (n_14269));
NAND2X1 g67878(.A (n_14266), .B (n_10569), .Y (n_14267));
NOR2X1 g67880(.A (n_10329), .B (n_7081), .Y (n_14265));
AOI21X1 g67884(.A0 (n_1513), .A1 (n_2259), .B0 (n_9673), .Y(n_14264));
INVX1 g67885(.A (n_12493), .Y (n_14263));
OR2X1 g67888(.A (n_1582), .B (n_17744), .Y (n_14262));
NAND2X1 g67889(.A (n_26731), .B (n_28137), .Y (n_14261));
AOI21X1 g67890(.A0 (n_11682), .A1 (n_7769), .B0 (n_3459), .Y(n_14259));
NAND2X1 g67894(.A (n_14257), .B (n_13310), .Y (n_14258));
AND2X1 g67903(.A (n_10402), .B (n_7470), .Y (n_14254));
NAND2X1 g67904(.A (n_14252), .B (n_13301), .Y (n_14253));
NOR2X1 g67906(.A (n_2289), .B (n_9142), .Y (n_18602));
AND2X1 g67909(.A (n_10402), .B (n_8290), .Y (n_14251));
NAND2X1 g67913(.A (n_12973), .B (n_8897), .Y (n_14250));
OR2X1 g67917(.A (n_16416), .B (n_14484), .Y (n_15984));
NAND2X1 g67922(.A (n_18074), .B (n_14246), .Y (n_14247));
INVX1 g67923(.A (n_14244), .Y (n_14245));
AND2X1 g67926(.A (n_14242), .B (n_12222), .Y (n_14243));
NAND2X1 g67928(.A (n_14190), .B (n_14240), .Y (n_14241));
NAND2X1 g67932(.A (n_9976), .B (n_18854), .Y (n_14239));
OR2X1 g67947(.A (n_14183), .B (n_26270), .Y (n_14237));
AND2X1 g67958(.A (n_15245), .B (n_14510), .Y (n_14236));
AND2X1 g67959(.A (n_9696), .B (n_11576), .Y (n_14235));
INVX1 g67960(.A (n_12460), .Y (n_14233));
NAND2X1 g67971(.A (n_14231), .B (n_10474), .Y (n_14232));
OR2X1 g67972(.A (n_14380), .B (n_15039), .Y (n_14230));
NAND2X1 g67981(.A (n_10968), .B (n_19896), .Y (n_18245));
AND2X1 g67983(.A (n_10339), .B (n_29000), .Y (n_14228));
NOR2X1 g67993(.A (n_14046), .B (n_10347), .Y (n_14226));
NAND2X1 g67994(.A (n_9061), .B (n_8523), .Y (n_14225));
NAND2X1 g67998(.A (n_8098), .B (n_14222), .Y (n_14223));
NAND2X1 g67999(.A (n_14100), .B (n_8801), .Y (n_14221));
NOR2X1 g68000(.A (n_12635), .B (n_10181), .Y (n_14220));
OR2X1 g68001(.A (n_14336), .B (n_4898), .Y (n_14219));
OR2X1 g68012(.A (n_14216), .B (n_19364), .Y (n_14217));
AND2X1 g68016(.A (n_14213), .B (n_11669), .Y (n_14214));
NAND2X1 g68031(.A (n_27411), .B (n_19857), .Y (n_17125));
AND2X1 g68032(.A (n_5282), .B (n_14222), .Y (n_14210));
NOR2X1 g68034(.A (n_10087), .B (n_15688), .Y (n_17908));
NAND2X1 g68047(.A (n_7088), .B (n_14208), .Y (n_14209));
INVX1 g68049(.A (n_12430), .Y (n_14207));
NAND2X1 g68062(.A (n_11298), .B (n_14478), .Y (n_14206));
NAND2X1 g68063(.A (n_9672), .B (n_14598), .Y (n_14205));
NOR2X1 g68076(.A (n_9904), .B (n_15039), .Y (n_14204));
NAND2X1 g68077(.A (n_9802), .B (n_14402), .Y (n_14203));
OR2X1 g68078(.A (n_11975), .B (n_14201), .Y (n_14202));
OR2X1 g68080(.A (n_14460), .B (n_14026), .Y (n_14200));
NAND2X1 g68082(.A (n_8897), .B (n_11949), .Y (n_14198));
NAND2X1 g68084(.A (n_11843), .B (n_15104), .Y (n_14196));
OR2X1 g68087(.A (n_10135), .B (n_12979), .Y (n_14195));
NAND2X1 g68089(.A (n_14193), .B (n_1238), .Y (n_14194));
INVX1 g68095(.A (n_12405), .Y (n_14192));
AND2X1 g68097(.A (n_9028), .B (n_14190), .Y (n_14191));
NOR2X1 g68102(.A (n_10395), .B (n_14188), .Y (n_14189));
NAND2X1 g68103(.A (n_14186), .B (n_12268), .Y (n_14187));
NOR2X1 g68104(.A (n_9897), .B (n_12591), .Y (n_14185));
INVX1 g68107(.A (n_12395), .Y (n_20535));
NAND2X1 g68122(.A (n_8546), .B (n_14183), .Y (n_14184));
NAND2X1 g68124(.A (n_14181), .B (n_9143), .Y (n_14182));
NAND2X1 g68125(.A (n_9143), .B (n_17681), .Y (n_14180));
NOR2X1 g68127(.A (n_7878), .B (n_12362), .Y (n_14179));
AND2X1 g68128(.A (n_7339), .B (n_14139), .Y (n_14177));
NAND2X1 g68130(.A (n_5745), .B (n_11710), .Y (n_14176));
NAND2X1 g68133(.A (n_10062), .B (n_13815), .Y (n_14175));
NAND2X1 g68134(.A (n_8020), .B (n_8737), .Y (n_14173));
INVX1 g68136(.A (n_12384), .Y (n_14171));
NAND2X1 g68138(.A (n_9402), .B (n_9142), .Y (n_14170));
NAND2X1 g68139(.A (n_7912), .B (n_8691), .Y (n_14169));
NAND2X1 g68141(.A (n_26881), .B (n_3582), .Y (n_14167));
NAND2X1 g68142(.A (n_3634), .B (n_9748), .Y (n_14165));
NAND2X1 g68145(.A (n_5448), .B (n_9526), .Y (n_14164));
NAND2X1 g68160(.A (n_16346), .B (n_9133), .Y (n_15947));
NAND2X1 g68165(.A (n_9832), .B (n_16754), .Y (n_14160));
NOR2X1 g68167(.A (n_27745), .B (n_7911), .Y (n_14159));
NAND2X1 g68178(.A (n_14157), .B (n_9075), .Y (n_14158));
NOR2X1 g68181(.A (n_14155), .B (n_12067), .Y (n_14156));
NAND2X1 g68186(.A (n_8267), .B (n_11923), .Y (n_14154));
NAND2X1 g68193(.A (n_14152), .B (n_11462), .Y (n_14153));
INVX1 g68195(.A (n_14150), .Y (n_14151));
INVX1 g68197(.A (n_12364), .Y (n_14149));
NAND2X1 g68200(.A (n_4344), .B (n_11712), .Y (n_14148));
OR2X1 g68203(.A (n_16466), .B (n_8671), .Y (n_20853));
NAND2X1 g68204(.A (n_14146), .B (n_12313), .Y (n_14147));
NOR2X1 g68205(.A (n_10018), .B (n_8452), .Y (n_14145));
NAND2X1 g68209(.A (n_6480), .B (n_13518), .Y (n_14143));
OR2X1 g68212(.A (n_8675), .B (n_14142), .Y (n_20468));
NAND2X1 g68213(.A (n_14141), .B (n_9371), .Y (n_16867));
INVX1 g68215(.A (n_12358), .Y (n_15937));
NAND2X1 g68222(.A (n_14139), .B (n_14138), .Y (n_14140));
INVX1 g68227(.A (n_12351), .Y (n_14137));
NOR2X1 g68231(.A (n_263), .B (n_10812), .Y (n_15934));
NOR2X1 g68234(.A (n_7635), .B (n_11322), .Y (n_15932));
NOR2X1 g68239(.A (n_7386), .B (n_8883), .Y (n_14135));
NAND2X1 g68241(.A (n_16342), .B (n_9020), .Y (n_14134));
INVX1 g68255(.A (n_15644), .Y (n_14133));
AND2X1 g68257(.A (n_15042), .B (n_14464), .Y (n_14132));
NAND2X1 g68262(.A (n_14864), .B (n_15177), .Y (n_15926));
NOR2X1 g68263(.A (n_6542), .B (n_10337), .Y (n_14131));
NOR2X1 g68268(.A (n_1063), .B (n_14130), .Y (n_17337));
NOR2X1 g68269(.A (n_10484), .B (n_14128), .Y (n_14129));
NAND2X1 g68274(.A (n_10418), .B (n_14126), .Y (n_14127));
NAND2X1 g68275(.A (n_9738), .B (n_12986), .Y (n_14125));
INVX1 g68284(.A (n_12331), .Y (n_14123));
AND2X1 g68296(.A (n_9748), .B (n_14120), .Y (n_14121));
NAND2X2 g68300(.A (n_11958), .B (n_9357), .Y (n_18268));
NAND3X1 g65379(.A (n_9129), .B (n_14872), .C (n_8152), .Y (n_14116));
NAND2X1 g68315(.A (n_5366), .B (n_8552), .Y (n_14115));
NAND2X1 g68316(.A (n_14113), .B (n_11088), .Y (n_14114));
INVX1 g68317(.A (n_12321), .Y (n_14112));
NOR2X1 g68319(.A (n_10581), .B (n_14141), .Y (n_14111));
NAND2X1 g68320(.A (n_8650), .B (n_26492), .Y (n_14110));
NAND2X1 g68322(.A (n_9006), .B (n_15596), .Y (n_14108));
AND2X1 g68329(.A (n_14107), .B (n_14681), .Y (n_20239));
NAND2X1 g68331(.A (n_16338), .B (n_9522), .Y (n_14106));
NAND2X1 g68335(.A (n_11088), .B (n_6534), .Y (n_14105));
NAND2X1 g68338(.A (n_11953), .B (n_5700), .Y (n_17851));
NAND2X1 g68347(.A (n_13269), .B (n_15316), .Y (n_14102));
NAND2X1 g68350(.A (n_14100), .B (n_7414), .Y (n_14101));
NAND2X1 g68352(.A (n_14099), .B (n_17706), .Y (n_16827));
NAND2X1 g68353(.A (n_9786), .B (n_17104), .Y (n_14098));
INVX1 g68360(.A (n_12300), .Y (n_14097));
NOR2X1 g68363(.A (n_13432), .B (n_19791), .Y (n_14096));
NAND2X1 g68364(.A (n_14094), .B (n_14093), .Y (n_14095));
NOR2X1 g68377(.A (n_4689), .B (n_6463), .Y (n_15913));
NAND2X1 g68378(.A (n_27287), .B (n_9285), .Y (n_17839));
NAND2X1 g68385(.A (n_14087), .B (n_11893), .Y (n_14088));
AND2X1 g68400(.A (n_15045), .B (n_14085), .Y (n_14086));
INVX1 g68408(.A (n_12279), .Y (n_15906));
NAND2X1 g68416(.A (n_10462), .B (n_14080), .Y (n_14081));
AND2X1 g68419(.A (n_7511), .B (n_14078), .Y (n_14079));
NAND2X1 g68428(.A (n_14100), .B (n_4444), .Y (n_14077));
NAND2X1 g68439(.A (n_14074), .B (n_10245), .Y (n_14075));
NAND3X1 g68448(.A (n_7637), .B (n_5037), .C (n_7996), .Y (n_14070));
INVX1 g72211(.A (n_15068), .Y (n_15743));
NAND3X1 g68449(.A (n_6784), .B (n_5263), .C (n_5542), .Y (n_14069));
OR2X1 g68451(.A (n_10025), .B (n_14067), .Y (n_14068));
NAND2X1 g68458(.A (n_9707), .B (n_18320), .Y (n_14066));
NAND2X1 g68471(.A (n_8013), .B (n_14138), .Y (n_14064));
OAI21X1 g68475(.A0 (n_5884), .A1 (n_6534), .B0 (n_14061), .Y(n_14063));
NAND2X1 g68476(.A (n_9660), .B (n_14240), .Y (n_14060));
NAND2X1 g68483(.A (n_7391), .B (n_28062), .Y (n_14059));
NAND2X1 g68486(.A (n_8963), .B (n_28580), .Y (n_14058));
OAI21X1 g68488(.A0 (n_8048), .A1 (n_14055), .B0 (n_14054), .Y(n_14056));
NAND2X1 g68490(.A (n_9891), .B (n_8588), .Y (n_14053));
AND2X1 g68491(.A (n_10306), .B (n_19752), .Y (n_14052));
NAND2X1 g68501(.A (n_9912), .B (n_6463), .Y (n_14051));
NOR2X1 g68504(.A (n_8325), .B (n_10036), .Y (n_14050));
NOR2X1 g68509(.A (n_5603), .B (n_14048), .Y (n_14049));
NOR2X1 g68517(.A (n_14046), .B (n_25801), .Y (n_14047));
NAND2X1 g68520(.A (n_4646), .B (n_14044), .Y (n_14045));
INVX1 g68521(.A (n_12233), .Y (n_14043));
NOR2X1 g68525(.A (n_9769), .B (n_12555), .Y (n_14042));
INVX1 g68526(.A (n_12227), .Y (n_14041));
OAI21X1 g68529(.A0 (n_8036), .A1 (n_27688), .B0 (n_6813), .Y(n_14040));
AOI21X1 g68530(.A0 (n_5957), .A1 (n_6601), .B0 (n_27099), .Y(n_14039));
NOR2X1 g68531(.A (n_10396), .B (n_14037), .Y (n_14038));
AOI21X1 g68533(.A0 (n_4327), .A1 (n_2592), .B0 (n_15395), .Y(n_14036));
NAND2X1 g68542(.A (n_7351), .B (n_11909), .Y (n_14034));
AOI21X1 g68545(.A0 (n_7917), .A1 (n_2112), .B0 (n_9039), .Y(n_14033));
NAND2X1 g68547(.A (n_10346), .B (n_11918), .Y (n_14032));
AOI21X1 g68548(.A0 (n_7329), .A1 (n_29102), .B0 (n_11764), .Y(n_14031));
NAND2X1 g68551(.A (n_14028), .B (n_29426), .Y (n_14029));
OAI21X1 g68552(.A0 (n_7650), .A1 (n_14026), .B0 (n_7353), .Y(n_14027));
AOI21X1 g68560(.A0 (n_6742), .A1 (n_7902), .B0 (n_29065), .Y(n_14025));
NAND2X1 g68579(.A (n_9966), .B (n_18876), .Y (n_14021));
AOI21X1 g68580(.A0 (n_4912), .A1 (n_6390), .B0 (n_16754), .Y(n_14020));
AOI21X1 g68583(.A0 (n_2716), .A1 (n_1626), .B0 (n_14017), .Y(n_14019));
NAND2X1 g68584(.A (n_9703), .B (n_15776), .Y (n_29301));
NAND2X1 g68598(.A (n_10250), .B (n_14014), .Y (n_14015));
NOR2X1 g68599(.A (n_7599), .B (n_11705), .Y (n_14013));
AOI21X1 g68600(.A0 (n_5410), .A1 (n_28575), .B0 (n_10520), .Y(n_14012));
AOI21X1 g68602(.A0 (n_4429), .A1 (n_9084), .B0 (n_10267), .Y(n_14011));
NAND2X1 g68607(.A (n_10296), .B (n_14009), .Y (n_14010));
NAND2X1 g68609(.A (n_10263), .B (n_14007), .Y (n_14008));
NAND2X1 g68615(.A (n_7520), .B (n_10089), .Y (n_14006));
INVX1 g68624(.A (n_12186), .Y (n_14005));
NAND2X1 g68626(.A (n_10290), .B (n_10832), .Y (n_14004));
NAND2X1 g68629(.A (n_7102), .B (n_10496), .Y (n_14003));
AOI21X1 g68637(.A0 (n_5019), .A1 (n_12019), .B0 (n_10455), .Y(n_14002));
NAND2X1 g68648(.A (n_10373), .B (n_11698), .Y (n_14001));
NAND2X1 g68656(.A (n_5634), .B (n_10535), .Y (n_14000));
NAND2X1 g68660(.A (n_10449), .B (n_17725), .Y (n_13999));
NAND2X1 g68661(.A (n_7345), .B (n_9825), .Y (n_13998));
NOR2X1 g68668(.A (n_6027), .B (n_9626), .Y (n_13997));
NOR2X1 g68670(.A (n_7310), .B (n_11756), .Y (n_13996));
AOI21X1 g68672(.A0 (n_3160), .A1 (n_2674), .B0 (n_10367), .Y(n_13995));
NAND2X1 g68675(.A (n_10400), .B (n_14362), .Y (n_13994));
OAI21X1 g68676(.A0 (n_6636), .A1 (n_13991), .B0 (n_11902), .Y(n_13993));
OAI21X1 g68678(.A0 (n_6444), .A1 (n_13991), .B0 (n_4093), .Y(n_13992));
OAI21X1 g68683(.A0 (n_3459), .A1 (n_3144), .B0 (n_14464), .Y(n_13990));
NAND2X1 g68685(.A (n_5130), .B (n_14571), .Y (n_13989));
NAND2X1 g68695(.A (n_10183), .B (n_11350), .Y (n_13988));
OAI21X1 g68702(.A0 (n_1777), .A1 (n_3119), .B0 (n_14510), .Y(n_13987));
NAND2X1 g68709(.A (n_5176), .B (n_14526), .Y (n_13986));
NAND2X1 g68710(.A (n_5168), .B (n_14521), .Y (n_13985));
OAI21X1 g68718(.A0 (n_2052), .A1 (n_4165), .B0 (n_14343), .Y(n_13984));
OAI21X1 g68721(.A0 (n_2327), .A1 (n_4187), .B0 (n_13310), .Y(n_13982));
NAND2X1 g68723(.A (n_5159), .B (n_14407), .Y (n_13980));
OAI21X1 g68730(.A0 (n_1807), .A1 (n_1825), .B0 (n_13301), .Y(n_13979));
AOI21X1 g68733(.A0 (n_8097), .A1 (n_12784), .B0 (n_13976), .Y(n_13977));
NAND2X1 g68734(.A (n_9949), .B (n_13974), .Y (n_13975));
OAI21X1 g68737(.A0 (n_4301), .A1 (n_4770), .B0 (n_4367), .Y(n_13973));
NAND2X1 g68741(.A (n_9852), .B (n_13971), .Y (n_13972));
NAND3X1 g68747(.A (n_10385), .B (n_4938), .C (n_8137), .Y (n_13970));
NAND2X1 g68753(.A (n_9732), .B (n_9730), .Y (n_13967));
NAND2X1 g68757(.A (n_9884), .B (n_13965), .Y (n_13966));
NAND2X1 g68761(.A (n_5471), .B (n_26469), .Y (n_13964));
OAI21X1 g68763(.A0 (n_9385), .A1 (n_2215), .B0 (n_13962), .Y(n_13963));
NAND2X1 g68770(.A (n_9864), .B (n_13960), .Y (n_13961));
NAND2X1 g68771(.A (n_10084), .B (n_10195), .Y (n_13959));
NAND2X1 g68777(.A (n_9834), .B (n_10361), .Y (n_13958));
NAND2X1 g68782(.A (n_10000), .B (n_9809), .Y (n_13957));
NAND2X1 g68785(.A (n_10028), .B (n_13955), .Y (n_13956));
XOR2X1 g68807(.A (n_1088), .B (n_7893), .Y (n_13954));
XOR2X1 g68813(.A (n_1281), .B (n_7888), .Y (n_13953));
XOR2X1 g68825(.A (n_983), .B (n_9204), .Y (n_13952));
XOR2X1 g68832(.A (n_1038), .B (n_8915), .Y (n_15850));
XOR2X1 g68834(.A (n_1074), .B (n_7882), .Y (n_13951));
XOR2X1 g68837(.A (n_977), .B (n_7883), .Y (n_13950));
NOR2X1 g68970(.A (n_9588), .B (n_12917), .Y (n_15847));
NAND4X1 g62242(.A (n_15692), .B (n_8114), .C (n_7674), .D (n_6136),.Y (n_13949));
INVX1 g69041(.A (n_12108), .Y (n_15846));
NOR2X1 g65359(.A (n_10829), .B (n_10283), .Y (n_13939));
NAND2X1 g65399(.A (n_11068), .B (n_17260), .Y (n_13935));
NAND2X1 g69795(.A (n_11632), .B (n_5558), .Y (n_13931));
INVX1 g69902(.A (n_13927), .Y (n_19781));
INVX1 g69966(.A (n_13921), .Y (n_18151));
NAND2X1 g69996(.A (n_8068), .B (n_28433), .Y (n_13920));
OR2X1 g70098(.A (n_9796), .B (n_9257), .Y (n_13917));
INVX1 g70109(.A (n_17935), .Y (n_13915));
OR2X1 g70129(.A (n_9424), .B (n_8928), .Y (n_13914));
INVX1 g70138(.A (n_13912), .Y (n_15817));
OR2X1 g70195(.A (n_13909), .B (n_9084), .Y (n_13910));
INVX1 g70238(.A (n_13907), .Y (n_18904));
INVX1 g65391(.A (n_11990), .Y (n_13900));
INVX1 g70303(.A (n_13898), .Y (n_13899));
OR2X1 g70315(.A (n_13895), .B (n_14055), .Y (n_13896));
INVX1 g70423(.A (n_8824), .Y (n_15816));
INVX1 g70525(.A (n_15918), .Y (n_13886));
INVX2 g70526(.A (n_15918), .Y (n_13885));
INVX1 g70527(.A (n_15918), .Y (n_13884));
INVX1 g70561(.A (n_13882), .Y (n_17563));
INVX1 g70665(.A (n_13880), .Y (n_13881));
INVX1 g70703(.A (n_13879), .Y (n_15811));
NAND2X1 g70739(.A (n_13875), .B (n_10146), .Y (n_21120));
NAND2X1 g72002(.A (n_11649), .B (n_13872), .Y (n_13873));
INVX1 g70760(.A (n_16187), .Y (n_13871));
NOR2X1 g70883(.A (n_10157), .B (n_9641), .Y (n_13864));
INVX1 g70994(.A (n_16139), .Y (n_13858));
AND2X1 g71088(.A (n_9424), .B (n_13855), .Y (n_13857));
NAND2X1 g71094(.A (n_9614), .B (n_13768), .Y (n_25565));
NOR2X1 g71102(.A (n_7262), .B (n_8030), .Y (n_13853));
OR2X1 g71165(.A (n_13851), .B (n_16434), .Y (n_13852));
INVX1 g71175(.A (n_13848), .Y (n_13849));
NAND2X1 g71199(.A (n_16006), .B (n_29333), .Y (n_17540));
OR2X1 g71249(.A (n_9601), .B (n_13846), .Y (n_13847));
NOR2X1 g71964(.A (n_13851), .B (n_13834), .Y (n_15762));
NAND2X1 g71276(.A (n_9610), .B (n_13787), .Y (n_25660));
INVX1 g71291(.A (n_13843), .Y (n_19844));
NOR2X1 g71317(.A (n_9962), .B (n_5131), .Y (n_13842));
INVX1 g71352(.A (n_27077), .Y (n_15792));
NAND2X1 g71438(.A (n_10376), .B (n_8520), .Y (n_13839));
INVX1 g71467(.A (n_17253), .Y (n_13838));
NAND2X1 g71496(.A (n_29333), .B (n_13837), .Y (n_17888));
INVX1 g71555(.A (n_13835), .Y (n_17906));
NAND2X1 g71653(.A (n_7997), .B (n_6534), .Y (n_25502));
INVX1 g71710(.A (n_11818), .Y (n_29179));
NAND2X1 g71716(.A (n_7610), .B (n_13909), .Y (n_13828));
NOR2X1 g71850(.A (n_9674), .B (n_1196), .Y (n_13827));
INVX1 g71872(.A (n_13825), .Y (n_13826));
AOI21X1 g62913(.A0 (n_6766), .A1 (n_13504), .B0 (n_933), .Y(n_13822));
INVX1 g72006(.A (n_11787), .Y (n_13820));
INVX1 g72017(.A (n_13818), .Y (n_13819));
OR2X1 g72054(.A (n_9607), .B (n_10226), .Y (n_13817));
OAI21X1 g62932(.A0 (n_9290), .A1 (n_7443), .B0 (n_13815), .Y(n_13816));
OAI21X1 g62933(.A0 (n_9306), .A1 (n_8986), .B0 (n_27604), .Y(n_13814));
OAI21X1 g62934(.A0 (n_9215), .A1 (n_7490), .B0 (n_13466), .Y(n_13813));
OAI21X1 g62935(.A0 (n_9308), .A1 (n_7365), .B0 (n_12986), .Y(n_13812));
OAI21X1 g62937(.A0 (n_9282), .A1 (n_5979), .B0 (n_15776), .Y(n_13811));
INVX1 g72094(.A (n_20582), .Y (n_13810));
OAI21X1 g62940(.A0 (n_9255), .A1 (n_7594), .B0 (n_26670), .Y(n_13809));
OAI21X1 g62943(.A0 (n_9247), .A1 (n_7495), .B0 (n_26276), .Y(n_13806));
OAI21X1 g62944(.A0 (n_9343), .A1 (n_7542), .B0 (n_13804), .Y(n_13805));
OAI21X1 g62945(.A0 (n_9241), .A1 (n_7348), .B0 (n_29065), .Y(n_13803));
OAI21X1 g62946(.A0 (n_9238), .A1 (n_7528), .B0 (n_28642), .Y(n_13802));
AND2X1 g72162(.A (n_13895), .B (n_13799), .Y (n_13800));
NAND3X1 g62957(.A (n_8769), .B (n_5354), .C (n_11528), .Y (n_13798));
AOI21X1 g62966(.A0 (n_9222), .A1 (n_16466), .B0 (n_10838), .Y(n_13797));
NAND3X1 g62976(.A (n_9961), .B (n_5194), .C (n_13351), .Y (n_13791));
NOR2X1 g72247(.A (n_28130), .B (n_9543), .Y (n_15741));
DFFX1 u0_r0_out_reg[25] (.CK (clk), .D (n_9649), .Q (u0_rcon_1054),.QN ());
NAND2X1 g72290(.A (n_9609), .B (n_13787), .Y (n_25669));
AOI21X1 g62996(.A0 (n_4997), .A1 (n_10923), .B0 (n_8708), .Y(n_13786));
NOR2X1 g72316(.A (n_11658), .B (n_21242), .Y (n_13784));
AOI21X1 g63005(.A0 (n_13782), .A1 (n_13725), .B0 (n_13804), .Y(n_13783));
OR2X1 g72416(.A (n_9629), .B (n_13593), .Y (n_13781));
NOR2X1 g72463(.A (n_8116), .B (n_9838), .Y (n_13778));
NAND3X1 g63062(.A (n_16704), .B (n_13316), .C (n_13776), .Y(n_13777));
INVX1 g72556(.A (n_17915), .Y (n_13775));
AND2X1 g72558(.A (n_13851), .B (n_13773), .Y (n_13774));
OAI21X1 g63072(.A0 (n_9162), .A1 (n_10305), .B0 (n_15894), .Y(n_13772));
INVX1 g72584(.A (n_13770), .Y (n_13771));
NAND2X1 g72605(.A (n_9619), .B (n_13768), .Y (n_13769));
INVX1 g72658(.A (n_13766), .Y (n_13767));
INVX1 g72665(.A (n_13765), .Y (n_18164));
AND2X1 g63103(.A (n_13763), .B (n_16564), .Y (n_13764));
AOI21X1 g63106(.A0 (n_9387), .A1 (n_13537), .B0 (n_12788), .Y(n_13762));
AOI21X1 g63108(.A0 (n_9219), .A1 (n_10366), .B0 (n_16754), .Y(n_13761));
INVX1 g72709(.A (n_11880), .Y (n_13760));
AND2X1 g72744(.A (n_6952), .B (n_13773), .Y (n_13759));
OAI21X1 g63128(.A0 (n_9192), .A1 (n_8353), .B0 (n_19143), .Y(n_13758));
OAI21X1 g63134(.A0 (n_9161), .A1 (n_11413), .B0 (n_18369), .Y(n_13756));
AND2X1 g63160(.A (n_13753), .B (n_13752), .Y (n_13754));
INVX1 g72916(.A (n_20567), .Y (n_13751));
NAND3X1 g63170(.A (n_13220), .B (n_8293), .C (n_18361), .Y (n_13750));
INVX1 g72951(.A (n_13748), .Y (n_17596));
INVX1 g72952(.A (n_13748), .Y (n_13749));
NAND2X1 g72960(.A (n_9604), .B (n_13768), .Y (n_29379));
INVX1 g72997(.A (n_13744), .Y (n_17653));
NAND2X1 g73012(.A (n_9676), .B (n_14484), .Y (n_13743));
NAND3X1 g63197(.A (n_9529), .B (n_9365), .C (n_17266), .Y (n_13742));
INVX1 g73039(.A (n_13740), .Y (n_13741));
OAI21X1 g63216(.A0 (n_9159), .A1 (n_13738), .B0 (n_12827), .Y(n_13739));
NAND2X1 g73183(.A (n_8346), .B (n_9656), .Y (n_17588));
NAND2X1 g73257(.A (n_7964), .B (n_8197), .Y (n_13736));
NOR2X1 g73258(.A (n_3082), .B (n_7753), .Y (n_13735));
NAND2X1 g73264(.A (n_7868), .B (n_9424), .Y (n_13734));
OAI21X1 g63278(.A0 (n_13340), .A1 (n_8879), .B0 (n_1424), .Y(n_13733));
AOI21X1 g73302(.A0 (n_10768), .A1 (n_11418), .B0 (n_9628), .Y(n_13732));
OAI21X1 g63338(.A0 (n_9158), .A1 (n_13730), .B0 (n_17912), .Y(n_13731));
AOI21X1 g60409(.A0 (n_7862), .A1 (n_13728), .B0 (n_2711), .Y(n_13729));
NAND3X1 g63361(.A (n_11079), .B (n_8615), .C (n_11484), .Y (n_13727));
NAND4X1 g63389(.A (n_13725), .B (n_13724), .C (n_6878), .D (n_7298),.Y (n_13726));
NAND3X1 g63391(.A (n_10723), .B (n_28902), .C (n_13722), .Y(n_13723));
NAND3X1 g63442(.A (n_9188), .B (n_11154), .C (n_13720), .Y (n_13721));
NAND2X1 g63450(.A (n_9595), .B (n_20116), .Y (n_13719));
NAND3X1 g63501(.A (n_11025), .B (n_7727), .C (n_14868), .Y (n_13717));
AOI21X1 g63566(.A0 (n_9180), .A1 (n_11431), .B0 (n_17912), .Y(n_13716));
NAND4X1 g63609(.A (n_11366), .B (n_11327), .C (n_7546), .D (n_12136),.Y (n_13714));
NAND4X1 g63630(.A (n_11353), .B (n_5759), .C (n_6066), .D (n_10675),.Y (n_13713));
NOR2X1 g63634(.A (n_9579), .B (n_14704), .Y (n_13712));
NAND4X1 g63655(.A (n_11316), .B (n_7710), .C (n_5751), .D (n_8613),.Y (n_13711));
AND2X1 g63696(.A (n_9560), .B (n_15039), .Y (n_13710));
AND2X1 g63726(.A (n_11457), .B (n_1424), .Y (n_13709));
NAND3X1 g63733(.A (n_29202), .B (n_10947), .C (n_13706), .Y(n_13708));
NAND4X1 g63822(.A (n_9460), .B (n_13704), .C (n_13703), .D (n_5402),.Y (n_13705));
NAND4X1 g63824(.A (n_11234), .B (n_13701), .C (n_13700), .D (n_7099),.Y (n_13702));
NAND4X1 g63833(.A (n_11192), .B (n_13698), .C (n_13697), .D (n_6906),.Y (n_13699));
NAND3X1 g63856(.A (n_9023), .B (n_13695), .C (n_12500), .Y (n_13696));
AOI22X1 g63910(.A0 (n_9187), .A1 (n_20010), .B0 (n_7576), .B1(n_7832), .Y (n_13694));
MX2X1 g63926(.A (n_11549), .B (n_13688), .S0 (n_16480), .Y (n_29366));
MX2X1 g63932(.A (n_15538), .B (n_13684), .S0 (n_20325), .Y (n_13685));
NAND4X1 g63950(.A (n_12879), .B (n_9425), .C (n_13681), .D (n_8859),.Y (n_13682));
AOI21X1 g64007(.A0 (n_9189), .A1 (n_13679), .B0 (n_10029), .Y(n_13680));
NAND4X1 g64010(.A (n_6233), .B (n_13962), .C (n_13700), .D (n_7056),.Y (n_13678));
NAND4X1 g64011(.A (n_7605), .B (n_13676), .C (n_13697), .D (n_4487),.Y (n_13677));
XOR2X1 g76146(.A (n_22964), .B (n_5817), .Y (n_13675));
OAI21X1 g64035(.A0 (n_8189), .A1 (n_4046), .B0 (n_18237), .Y(n_13674));
AOI21X1 g64036(.A0 (n_8034), .A1 (n_15966), .B0 (n_18440), .Y(n_13672));
OAI21X1 g64037(.A0 (n_8632), .A1 (n_4783), .B0 (n_27688), .Y(n_13671));
XOR2X1 g76195(.A (n_23545), .B (n_3301), .Y (n_13670));
AOI21X1 g64039(.A0 (n_8979), .A1 (n_7164), .B0 (n_11261), .Y(n_13668));
OAI21X1 g64043(.A0 (n_8424), .A1 (n_5494), .B0 (n_28167), .Y(n_13667));
AOI21X1 g64044(.A0 (n_8014), .A1 (n_5700), .B0 (n_12298), .Y(n_13666));
AOI21X1 g64045(.A0 (n_5193), .A1 (n_9285), .B0 (n_11576), .Y(n_13665));
AOI21X1 g64046(.A0 (n_8835), .A1 (n_8321), .B0 (n_18320), .Y(n_13664));
AOI21X1 g64047(.A0 (n_7948), .A1 (n_8268), .B0 (n_19857), .Y(n_13663));
OAI21X1 g64055(.A0 (n_8206), .A1 (n_7867), .B0 (n_18266), .Y(n_13661));
OAI21X1 g64058(.A0 (n_8364), .A1 (n_9823), .B0 (n_17260), .Y(n_13660));
OAI21X1 g64059(.A0 (n_8132), .A1 (n_10181), .B0 (n_9917), .Y(n_13659));
XOR2X1 g76247(.A (text_in_r[25] ), .B (n_124), .Y (n_13657));
OAI21X1 g64064(.A0 (n_8391), .A1 (n_13655), .B0 (n_12910), .Y(n_13656));
XOR2X1 g76254(.A (n_22557), .B (n_7410), .Y (n_13654));
OAI21X1 g64065(.A0 (n_8488), .A1 (n_6588), .B0 (n_16787), .Y(n_13652));
OAI21X1 g64066(.A0 (n_8612), .A1 (n_11671), .B0 (n_16835), .Y(n_13651));
OAI21X1 g64067(.A0 (n_8366), .A1 (n_8078), .B0 (n_15894), .Y(n_13649));
OAI21X1 g64068(.A0 (n_9338), .A1 (n_13646), .B0 (n_15712), .Y(n_13647));
INVX1 g64071(.A (n_11602), .Y (n_13645));
AOI21X1 g64074(.A0 (n_7900), .A1 (n_7511), .B0 (n_17260), .Y(n_13644));
OAI21X1 g64076(.A0 (n_8381), .A1 (n_11667), .B0 (n_17260), .Y(n_13642));
NOR2X1 g64077(.A (n_10774), .B (n_14624), .Y (n_13640));
OAI21X1 g64078(.A0 (n_8688), .A1 (n_11660), .B0 (n_27688), .Y(n_13638));
OAI21X1 g64081(.A0 (n_8720), .A1 (n_7755), .B0 (n_13804), .Y(n_13637));
AOI21X1 g64088(.A0 (n_8595), .A1 (n_7339), .B0 (n_27688), .Y(n_13636));
AOI21X1 g64090(.A0 (n_9237), .A1 (n_7324), .B0 (n_16434), .Y(n_13635));
OAI21X1 g64091(.A0 (n_8210), .A1 (n_7953), .B0 (n_9819), .Y(n_13633));
OAI21X1 g64092(.A0 (n_9553), .A1 (n_9718), .B0 (n_14155), .Y(n_13632));
OAI21X1 g64093(.A0 (n_8297), .A1 (n_8118), .B0 (n_263), .Y (n_13630));
NAND2X1 g64095(.A (n_11106), .B (n_21174), .Y (n_13628));
INVX1 g64096(.A (n_11598), .Y (n_13626));
AOI21X1 g64098(.A0 (n_6569), .A1 (n_16539), .B0 (sa20[1] ), .Y(n_13625));
AND2X1 g64101(.A (n_10867), .B (n_5131), .Y (n_13624));
AND2X1 g64103(.A (n_10864), .B (n_13326), .Y (n_13623));
AOI21X1 g64105(.A0 (n_6555), .A1 (n_14120), .B0 (sa30[1] ), .Y(n_13622));
AOI21X1 g64110(.A0 (n_5345), .A1 (n_15090), .B0 (n_20574), .Y(n_13621));
AND2X1 g64111(.A (n_10810), .B (n_1196), .Y (n_13619));
AOI21X1 g64112(.A0 (n_7952), .A1 (n_14574), .B0 (sa31[1] ), .Y(n_13618));
INVX1 g64116(.A (n_11590), .Y (n_21227));
NAND2X1 g64124(.A (n_11223), .B (n_16480), .Y (n_13617));
OR2X1 g64125(.A (n_16550), .B (n_13083), .Y (n_19314));
OR4X1 g64130(.A (n_18237), .B (n_6534), .C (n_8816), .D (n_6715), .Y(n_13616));
INVX1 g64131(.A (n_11586), .Y (n_13614));
NOR2X1 g64134(.A (n_13612), .B (n_4582), .Y (n_13613));
NOR2X1 g64136(.A (n_12697), .B (n_18679), .Y (n_13611));
OR2X1 g64139(.A (n_13610), .B (n_16480), .Y (n_21700));
AND2X1 g64142(.A (n_12725), .B (n_16466), .Y (n_17308));
NAND3X1 g64145(.A (n_17912), .B (n_13609), .C (n_16198), .Y(n_15427));
AOI21X1 g64151(.A0 (n_13607), .A1 (n_14548), .B0 (n_10763), .Y(n_13608));
NOR2X1 g64155(.A (n_13554), .B (n_13606), .Y (n_15424));
NAND2X1 g64156(.A (n_13604), .B (n_15674), .Y (n_13605));
NAND3X1 g64157(.A (n_27099), .B (n_13602), .C (n_11052), .Y(n_13603));
NOR2X1 g64166(.A (n_14155), .B (n_16793), .Y (n_15420));
NAND2X1 g64167(.A (n_15156), .B (n_16978), .Y (n_13598));
AND2X1 g64169(.A (n_13595), .B (n_15708), .Y (n_13596));
OR4X1 g64173(.A (n_18266), .B (n_13593), .C (n_12469), .D (n_6616),.Y (n_13594));
NOR2X1 g64177(.A (n_12301), .B (n_17567), .Y (n_13592));
OR2X1 g64192(.A (n_12514), .B (n_18168), .Y (n_13590));
NOR2X1 g64201(.A (n_13588), .B (n_14142), .Y (n_13589));
AND2X1 g64204(.A (n_12584), .B (n_19857), .Y (n_13587));
AND2X1 g64215(.A (n_13584), .B (n_11354), .Y (n_15390));
OR4X1 g64216(.A (n_14155), .B (n_14055), .C (n_4113), .D (n_6482), .Y(n_13582));
NAND2X1 g64217(.A (n_13064), .B (n_14142), .Y (n_13581));
AOI21X1 g64239(.A0 (n_8249), .A1 (n_8497), .B0 (sa33[1] ), .Y(n_13579));
AOI21X1 g64241(.A0 (n_6890), .A1 (n_12289), .B0 (n_20574), .Y(n_13578));
OAI21X1 g64262(.A0 (n_8627), .A1 (n_4451), .B0 (n_13575), .Y(n_13576));
NAND2X1 g64263(.A (n_13497), .B (n_26491), .Y (n_13574));
NAND3X1 g64264(.A (n_11345), .B (n_11031), .C (n_3991), .Y (n_13573));
OR2X1 g64265(.A (n_10698), .B (n_20325), .Y (n_13572));
NAND2X1 g64267(.A (n_11183), .B (n_13571), .Y (n_15362));
INVX1 g64268(.A (n_13569), .Y (n_13570));
NAND2X1 g64270(.A (n_12865), .B (n_13567), .Y (n_13568));
NAND2X1 g64278(.A (n_12995), .B (n_9737), .Y (n_13566));
NAND2X1 g64282(.A (n_13564), .B (n_29228), .Y (n_13565));
OR2X1 g64284(.A (n_13516), .B (n_10221), .Y (n_13563));
NAND3X1 g64285(.A (n_28829), .B (n_5415), .C (n_13561), .Y (n_13562));
NAND2X1 g64291(.A (n_13559), .B (n_14055), .Y (n_13560));
NAND2X1 g64308(.A (n_10241), .B (n_13556), .Y (n_13557));
NAND2X1 g64319(.A (n_15675), .B (n_13554), .Y (n_13555));
NOR2X1 g64323(.A (n_13585), .B (n_6001), .Y (n_13553));
AOI21X1 g64324(.A0 (n_8075), .A1 (n_13152), .B0 (n_16787), .Y(n_13552));
AOI21X1 g64329(.A0 (n_8444), .A1 (n_8096), .B0 (n_17069), .Y(n_13551));
NAND2X1 g64333(.A (n_12939), .B (n_13550), .Y (n_15324));
AOI21X1 g64337(.A0 (n_12243), .A1 (n_8973), .B0 (n_15688), .Y(n_13549));
NAND2X1 g64345(.A (n_13588), .B (n_13610), .Y (n_13548));
NAND2X1 g64351(.A (n_10704), .B (n_18440), .Y (n_13547));
NAND2X1 g64353(.A (n_27611), .B (n_18440), .Y (n_13546));
NAND2X1 g64358(.A (n_27899), .B (n_17864), .Y (n_15308));
NOR2X1 g64362(.A (n_13584), .B (n_9314), .Y (n_13544));
AND2X1 g64366(.A (n_13542), .B (n_9211), .Y (n_13543));
NAND2X1 g64368(.A (n_12319), .B (n_11261), .Y (n_17329));
NAND2X1 g64370(.A (n_13612), .B (n_13539), .Y (n_16985));
NAND3X1 g64379(.A (n_13537), .B (n_6971), .C (n_13536), .Y (n_13538));
NOR2X1 g64382(.A (n_10748), .B (n_8543), .Y (n_13535));
NAND3X1 g64385(.A (n_9526), .B (n_13532), .C (n_3999), .Y (n_13534));
INVX1 g64388(.A (n_13531), .Y (n_15294));
OR2X1 g64392(.A (n_10757), .B (n_17069), .Y (n_13530));
NAND2X1 g64398(.A (n_27153), .B (n_17089), .Y (n_15288));
NAND2X1 g64399(.A (n_13092), .B (n_17571), .Y (n_13528));
NAND3X1 g64400(.A (n_20360), .B (n_8668), .C (n_12451), .Y (n_13527));
NAND3X1 g64403(.A (n_9526), .B (n_13536), .C (n_9319), .Y (n_13526));
NAND2X1 g64409(.A (n_11117), .B (n_16414), .Y (n_15283));
NAND3X1 g64410(.A (n_7708), .B (n_6723), .C (n_6607), .Y (n_13525));
OR2X1 g64416(.A (n_13524), .B (n_16480), .Y (n_17062));
INVX1 g64417(.A (n_11553), .Y (n_25507));
NAND3X1 g64423(.A (n_17018), .B (n_11620), .C (n_13521), .Y(n_13522));
NAND2X1 g64426(.A (n_16758), .B (n_13519), .Y (n_13520));
NAND2X1 g64433(.A (n_15689), .B (n_13518), .Y (n_15274));
NAND2X1 g64434(.A (n_28986), .B (n_26492), .Y (n_13517));
NAND2X1 g64442(.A (n_13516), .B (n_17260), .Y (n_15269));
INVX1 g64444(.A (n_11545), .Y (n_13515));
NAND2X1 g64448(.A (n_15513), .B (n_14120), .Y (n_13514));
NAND2X1 g64449(.A (n_14765), .B (n_9061), .Y (n_13513));
NAND2X1 g64450(.A (n_16550), .B (n_13142), .Y (n_16997));
NOR2X1 g64456(.A (n_10686), .B (n_28037), .Y (n_13512));
AOI21X1 g64459(.A0 (n_7195), .A1 (n_7887), .B0 (n_1547), .Y(n_13511));
AND2X1 g64461(.A (n_12465), .B (n_16466), .Y (n_15262));
OR2X1 g64462(.A (n_10669), .B (n_13082), .Y (n_13510));
INVX1 g64469(.A (n_13506), .Y (n_13507));
AND2X1 g64471(.A (n_14512), .B (n_13504), .Y (n_13505));
NAND2X1 g64473(.A (n_9550), .B (n_28041), .Y (n_13503));
NOR2X1 g64485(.A (n_17754), .B (n_7410), .Y (n_13502));
NOR2X1 g64489(.A (n_29208), .B (n_13083), .Y (n_13499));
NOR2X1 g64490(.A (n_5839), .B (n_13497), .Y (n_13498));
AND2X1 g64492(.A (n_10825), .B (n_13495), .Y (n_13496));
NAND2X1 g64494(.A (n_12745), .B (n_9527), .Y (n_16992));
OR2X1 g64495(.A (n_10673), .B (n_13211), .Y (n_13493));
NAND2X1 g64496(.A (n_13491), .B (n_13490), .Y (n_13492));
INVX1 g64498(.A (n_11538), .Y (n_13489));
AOI21X1 g64500(.A0 (n_13487), .A1 (n_5514), .B0 (n_1132), .Y(n_13488));
OR2X1 g64510(.A (n_13411), .B (n_9892), .Y (n_13485));
NAND2X1 g64514(.A (n_13484), .B (n_12827), .Y (n_15240));
NAND2X1 g64515(.A (n_13482), .B (n_11348), .Y (n_13483));
NAND2X1 g64516(.A (n_10671), .B (n_3483), .Y (n_13481));
NOR2X1 g64521(.A (n_17939), .B (n_17414), .Y (n_25726));
NAND2X1 g64525(.A (n_13554), .B (n_13479), .Y (n_16995));
INVX1 g64531(.A (n_11532), .Y (n_25763));
NOR2X1 g64533(.A (n_13476), .B (n_13475), .Y (n_13477));
AOI21X1 g64536(.A0 (n_12844), .A1 (n_7459), .B0 (n_18679), .Y(n_13474));
AOI21X1 g64538(.A0 (n_16959), .A1 (n_13472), .B0 (n_1667), .Y(n_13473));
NAND2X1 g64539(.A (n_13470), .B (n_13469), .Y (n_13471));
AND2X1 g64540(.A (n_14493), .B (n_11416), .Y (n_13468));
NAND3X1 g64542(.A (n_8736), .B (n_7505), .C (n_4471), .Y (n_13467));
NAND2X1 g64544(.A (n_11138), .B (n_13466), .Y (n_18365));
OAI21X1 g64545(.A0 (n_4098), .A1 (n_7245), .B0 (n_3264), .Y(n_13465));
AOI21X1 g64547(.A0 (n_8145), .A1 (n_3551), .B0 (n_18369), .Y(n_13463));
NAND2X1 g64548(.A (n_10065), .B (n_15509), .Y (n_13462));
NAND2X1 g64553(.A (n_13460), .B (n_8295), .Y (n_13461));
NAND2X2 g64560(.A (n_20926), .B (n_14592), .Y (n_19542));
NOR2X1 g64561(.A (n_10767), .B (n_13458), .Y (n_28507));
NAND2X1 g64562(.A (n_10797), .B (n_12739), .Y (n_13457));
NAND2X1 g64569(.A (n_12813), .B (n_4582), .Y (n_17161));
AND2X1 g64570(.A (n_11539), .B (n_17621), .Y (n_13455));
AND2X1 g64581(.A (n_13452), .B (n_14491), .Y (n_29421));
NAND2X1 g64583(.A (n_13588), .B (n_13226), .Y (n_15210));
AND2X1 g64586(.A (n_10938), .B (n_18369), .Y (n_17151));
AOI21X1 g64595(.A0 (n_8489), .A1 (n_6654), .B0 (n_18266), .Y(n_13451));
NAND2X1 g64596(.A (n_13450), .B (n_1626), .Y (n_17265));
INVX1 g65386(.A (n_11474), .Y (n_13449));
AOI21X1 g64600(.A0 (n_8492), .A1 (n_7170), .B0 (n_15574), .Y(n_13448));
INVX1 g64603(.A (n_11514), .Y (n_13447));
NAND2X1 g64608(.A (n_13445), .B (n_13593), .Y (n_13446));
NAND2X1 g64610(.A (n_13443), .B (n_14478), .Y (n_13444));
NAND2X1 g64613(.A (n_9305), .B (n_13612), .Y (n_13442));
INVX1 g64618(.A (n_11511), .Y (n_13441));
NOR2X1 g64621(.A (n_4259), .B (n_12573), .Y (n_13440));
AND2X1 g64623(.A (n_10916), .B (n_8217), .Y (n_17269));
NOR2X1 g64633(.A (n_11024), .B (n_13484), .Y (n_13438));
NAND2X1 g64634(.A (n_10688), .B (n_12896), .Y (n_13437));
NAND2X1 g64635(.A (n_27646), .B (n_12896), .Y (n_13436));
NAND2X1 g65388(.A (n_11163), .B (n_17411), .Y (n_13435));
AND2X1 g64636(.A (n_10941), .B (n_16480), .Y (n_13434));
NAND2X1 g64637(.A (n_16704), .B (n_13432), .Y (n_13433));
AND2X1 g64639(.A (n_12922), .B (n_15674), .Y (n_15175));
NAND2X1 g64642(.A (n_13431), .B (n_27133), .Y (n_17157));
AND2X1 g64648(.A (n_13429), .B (n_13040), .Y (n_13430));
AND2X1 g64654(.A (n_10750), .B (n_18237), .Y (n_13428));
NAND2X1 g64656(.A (n_11158), .B (n_11261), .Y (n_17317));
NAND2X1 g64662(.A (n_13426), .B (n_12105), .Y (n_13427));
DFFX1 dcnt_reg[2] (.CK (clk), .D (n_11000), .Q (dcnt[2] ), .QN ());
NAND2X1 g64667(.A (n_13042), .B (n_26670), .Y (n_13425));
OAI21X1 g64673(.A0 (n_8412), .A1 (n_4570), .B0 (n_13423), .Y(n_13424));
NAND2X1 g64674(.A (n_12294), .B (n_13421), .Y (n_13422));
NAND2X1 g64686(.A (n_15463), .B (n_13207), .Y (n_13420));
AOI21X1 g64687(.A0 (n_8969), .A1 (n_13418), .B0 (n_18237), .Y(n_13419));
NOR2X1 g64691(.A (n_10598), .B (n_12875), .Y (n_13417));
AND2X1 g64693(.A (n_13416), .B (n_11593), .Y (n_15142));
NAND2X1 g64694(.A (n_13414), .B (n_9212), .Y (n_13415));
NAND2X1 g64709(.A (n_11002), .B (n_28692), .Y (n_15130));
INVX1 g64719(.A (n_11496), .Y (n_13412));
NAND2X1 g64727(.A (n_13411), .B (n_27688), .Y (n_15127));
INVX1 g64739(.A (n_11490), .Y (n_13410));
AND2X1 g64742(.A (n_13408), .B (n_14272), .Y (n_29313));
NAND2X1 g64746(.A (n_14991), .B (n_13195), .Y (n_15118));
NAND2X1 g64749(.A (n_12566), .B (n_9257), .Y (n_13407));
NAND2X1 g64752(.A (n_12990), .B (n_14183), .Y (n_13405));
INVX1 g64754(.A (n_11483), .Y (n_13404));
NAND2X1 g64759(.A (n_13402), .B (n_8928), .Y (n_13403));
NAND2X1 g64764(.A (n_15012), .B (n_13398), .Y (n_13399));
NOR2X1 g64768(.A (n_10977), .B (n_13341), .Y (n_13397));
NAND3X1 g64771(.A (n_11390), .B (n_29363), .C (n_4441), .Y (n_13396));
INVX1 g64774(.A (n_11480), .Y (n_13395));
AOI21X1 g64778(.A0 (n_8549), .A1 (n_7137), .B0 (n_18168), .Y(n_13393));
NAND2X1 g64782(.A (n_27710), .B (n_14765), .Y (n_25786));
AND2X1 g64785(.A (n_14823), .B (n_8730), .Y (n_13390));
NAND2X1 g64789(.A (n_11585), .B (n_15689), .Y (n_13389));
INVX1 g64801(.A (n_11468), .Y (n_13388));
NAND2X1 g64806(.A (n_28620), .B (n_13385), .Y (n_13387));
NAND2X1 g64807(.A (n_13383), .B (n_13382), .Y (n_13384));
NOR2X1 g64808(.A (n_17900), .B (n_13380), .Y (n_13381));
INVX1 g64812(.A (n_11465), .Y (n_13379));
NAND3X1 g64814(.A (n_29171), .B (n_4368), .C (n_13376), .Y (n_13378));
NAND2X1 g64815(.A (n_18286), .B (n_11080), .Y (n_13375));
NOR2X1 g64817(.A (n_15021), .B (n_14246), .Y (n_13374));
NAND2X1 g64819(.A (n_27140), .B (n_13372), .Y (n_13373));
NAND2X1 g64821(.A (n_13370), .B (n_10381), .Y (n_13371));
NAND2X1 g64825(.A (n_13368), .B (n_6008), .Y (n_13369));
OR2X1 g64832(.A (n_13366), .B (n_17912), .Y (n_13367));
AOI21X1 g64837(.A0 (n_8073), .A1 (n_13243), .B0 (n_12298), .Y(n_13365));
NAND2X1 g64838(.A (n_17821), .B (n_14616), .Y (n_13364));
NAND2X1 g64846(.A (n_11161), .B (n_13695), .Y (n_13363));
NAND2X1 g64847(.A (n_10982), .B (n_26276), .Y (n_15612));
NOR2X1 g64848(.A (n_17821), .B (n_9819), .Y (n_13362));
NAND2X1 g64860(.A (n_13295), .B (n_13360), .Y (n_13361));
NAND2X1 g64877(.A (n_13359), .B (n_19857), .Y (n_15630));
NAND2X1 g64884(.A (n_8215), .B (n_13357), .Y (n_13358));
NOR2X1 g64912(.A (n_11524), .B (n_9106), .Y (n_13356));
AOI21X1 g64919(.A0 (n_6709), .A1 (n_7258), .B0 (n_26276), .Y(n_13355));
NAND2X1 g64925(.A (n_6996), .B (n_13351), .Y (n_13352));
OR2X1 g64927(.A (n_15009), .B (n_15986), .Y (n_13350));
NAND2X1 g64930(.A (n_9210), .B (n_19433), .Y (n_13349));
NAND2X1 g64935(.A (n_13347), .B (n_13408), .Y (n_13348));
AOI21X1 g64945(.A0 (n_7132), .A1 (n_10732), .B0 (n_29048), .Y(n_13346));
OR2X1 g64946(.A (n_28809), .B (n_14624), .Y (n_13345));
OAI21X1 g64955(.A0 (n_7834), .A1 (n_17465), .B0 (n_27718), .Y(n_13344));
NOR2X1 g64956(.A (n_13341), .B (n_13340), .Y (n_13342));
AOI21X1 g64971(.A0 (n_7712), .A1 (n_10913), .B0 (n_15986), .Y(n_13337));
NOR2X1 g64975(.A (n_15012), .B (n_11576), .Y (n_13336));
NAND2X1 g64983(.A (n_4548), .B (n_13186), .Y (n_13335));
NAND2X1 g64989(.A (n_6922), .B (n_13333), .Y (n_13334));
NAND2X1 g64997(.A (n_14909), .B (n_10216), .Y (n_13332));
NOR2X1 g65003(.A (n_11470), .B (n_19896), .Y (n_13331));
NAND2X1 g65007(.A (n_5745), .B (n_13329), .Y (n_13330));
NAND3X1 g65011(.A (n_19008), .B (n_6964), .C (n_11043), .Y (n_13328));
NOR2X1 g65013(.A (n_13322), .B (n_13326), .Y (n_13327));
NAND2X1 g65014(.A (n_13324), .B (n_12448), .Y (n_13325));
NAND2X1 g65017(.A (n_13322), .B (n_12883), .Y (n_13323));
AND2X1 g65023(.A (n_15028), .B (n_13320), .Y (n_13321));
NOR2X1 g65027(.A (n_15028), .B (n_13318), .Y (n_13319));
NAND2X1 g65047(.A (n_13259), .B (n_13316), .Y (n_13317));
AOI21X1 g65050(.A0 (n_7455), .A1 (n_8371), .B0 (n_11489), .Y(n_13315));
NAND2X1 g65054(.A (n_11257), .B (n_9831), .Y (n_13314));
NOR2X1 g65056(.A (n_9099), .B (n_10824), .Y (n_13313));
INVX1 g65059(.A (n_11454), .Y (n_13312));
AOI21X1 g65067(.A0 (n_7286), .A1 (n_13310), .B0 (n_13804), .Y(n_13311));
NOR2X1 g65069(.A (n_28159), .B (n_10917), .Y (n_13309));
NOR2X1 g65070(.A (n_5932), .B (n_13307), .Y (n_13308));
NAND2X1 g65074(.A (n_13305), .B (n_7204), .Y (n_13306));
NOR2X1 g65075(.A (n_5393), .B (n_13303), .Y (n_29391));
AOI21X1 g65077(.A0 (n_7471), .A1 (n_13301), .B0 (n_263), .Y(n_13302));
INVX1 g65081(.A (n_11450), .Y (n_13300));
NAND2X1 g65083(.A (n_13298), .B (n_8258), .Y (n_13299));
NAND2X1 g65095(.A (n_13295), .B (n_8069), .Y (n_13296));
NAND2X1 g65117(.A (n_15034), .B (n_10072), .Y (n_13294));
AOI21X1 g65129(.A0 (n_6371), .A1 (n_5687), .B0 (n_19797), .Y(n_13293));
NAND2X1 g65137(.A (n_11096), .B (n_5329), .Y (n_14954));
OR2X1 g65146(.A (n_9171), .B (n_20767), .Y (n_13290));
AND2X1 g65151(.A (n_9199), .B (n_15776), .Y (n_13288));
NAND2X1 g65160(.A (n_27373), .B (n_15712), .Y (n_15678));
AOI21X1 g65164(.A0 (n_7316), .A1 (n_14324), .B0 (n_27688), .Y(n_13285));
NAND2X1 g65177(.A (n_8581), .B (n_13282), .Y (n_13283));
OR2X1 g65190(.A (n_28877), .B (n_9410), .Y (n_13281));
NAND2X1 g65194(.A (n_15236), .B (n_10975), .Y (n_13280));
NOR2X1 g70304(.A (n_8036), .B (n_8452), .Y (n_13898));
INVX1 g61100(.A (u0_rcon_1053), .Y (n_13279));
NAND3X1 g65238(.A (n_13277), .B (n_11422), .C (n_14523), .Y(n_13278));
AOI21X1 g65242(.A0 (n_7306), .A1 (n_13118), .B0 (n_18266), .Y(n_13276));
NOR2X1 g65249(.A (n_15260), .B (n_15708), .Y (n_13275));
AOI21X1 g65259(.A0 (n_7250), .A1 (n_5216), .B0 (n_9527), .Y(n_13274));
NAND2X1 g65265(.A (n_10893), .B (n_15776), .Y (n_15615));
NAND2X1 g65266(.A (n_13272), .B (n_17567), .Y (n_15621));
NOR2X1 g65272(.A (n_11539), .B (n_11261), .Y (n_13271));
NAND3X1 g65278(.A (n_11193), .B (n_7297), .C (n_13269), .Y (n_13270));
NAND2X1 g65280(.A (n_16663), .B (n_28160), .Y (n_13268));
NAND2X1 g65287(.A (n_9169), .B (n_17912), .Y (n_13267));
NOR2X1 g65306(.A (n_9165), .B (n_13076), .Y (n_13265));
NAND3X1 g65311(.A (n_18982), .B (n_5992), .C (n_11175), .Y (n_13263));
AOI21X1 g65317(.A0 (n_6780), .A1 (n_13137), .B0 (n_12896), .Y(n_13262));
NAND3X1 g65326(.A (n_13260), .B (n_5424), .C (n_13259), .Y (n_13261));
NAND3X1 g65334(.A (n_13257), .B (n_6283), .C (n_13256), .Y (n_13258));
NAND3X1 g65347(.A (n_12354), .B (n_4782), .C (n_6943), .Y (n_13255));
NAND3X1 g65348(.A (n_10817), .B (n_4814), .C (n_7046), .Y (n_13254));
INVX1 g65349(.A (n_11463), .Y (n_13253));
AOI21X1 g65401(.A0 (n_5575), .A1 (n_12594), .B0 (n_12910), .Y(n_13252));
NOR2X1 g65363(.A (n_9269), .B (n_8791), .Y (n_13250));
NAND3X1 g65385(.A (n_9111), .B (n_11200), .C (n_8737), .Y (n_13249));
AOI21X1 g65406(.A0 (n_8811), .A1 (n_14085), .B0 (n_13247), .Y(n_13248));
NAND2X1 g65407(.A (n_9301), .B (n_17912), .Y (n_13246));
NAND3X1 g65410(.A (n_13243), .B (n_8922), .C (n_8691), .Y (n_13244));
AOI21X1 g65418(.A0 (n_11565), .A1 (n_9907), .B0 (n_13815), .Y(n_13242));
OAI21X1 g65419(.A0 (n_5645), .A1 (n_14142), .B0 (n_11124), .Y(n_13241));
AOI21X1 g65421(.A0 (n_13239), .A1 (n_13236), .B0 (n_16480), .Y(n_13240));
NAND3X1 g65425(.A (n_16564), .B (n_13236), .C (n_18635), .Y(n_13237));
AND2X1 g65427(.A (n_9320), .B (n_14142), .Y (n_13235));
AOI21X1 g65433(.A0 (n_7153), .A1 (n_4195), .B0 (n_11126), .Y(n_13234));
NAND3X1 g65441(.A (n_4260), .B (n_9167), .C (n_5147), .Y (n_13233));
INVX1 g65447(.A (n_11440), .Y (n_13232));
NAND2X1 g65455(.A (n_7577), .B (n_11506), .Y (n_13231));
NAND2X1 g65463(.A (n_9449), .B (n_15243), .Y (n_13230));
AND2X1 g65464(.A (n_9191), .B (n_13083), .Y (n_13229));
NAND3X1 g65469(.A (n_9214), .B (n_13226), .C (n_9193), .Y (n_13227));
AOI21X1 g65477(.A0 (n_3438), .A1 (n_10936), .B0 (n_18369), .Y(n_13225));
NAND3X1 g65482(.A (n_13482), .B (n_7595), .C (n_13479), .Y (n_13223));
NAND3X1 g65484(.A (n_9557), .B (n_11495), .C (n_7726), .Y (n_13222));
AOI21X1 g65488(.A0 (n_13220), .A1 (n_13219), .B0 (n_13466), .Y(n_13221));
AOI21X1 g65491(.A0 (n_6247), .A1 (n_13217), .B0 (n_28037), .Y(n_13218));
AND2X1 g65494(.A (n_9297), .B (n_15674), .Y (n_13216));
NAND2X1 g65498(.A (n_6000), .B (n_13213), .Y (n_13214));
NAND3X1 g65509(.A (n_8534), .B (n_13211), .C (n_20577), .Y (n_13212));
AOI21X1 g65517(.A0 (n_11285), .A1 (n_8404), .B0 (n_28645), .Y(n_13210));
NAND3X1 g65520(.A (n_3237), .B (n_29336), .C (n_2923), .Y (n_13209));
NAND2X1 g65525(.A (n_5998), .B (n_13207), .Y (n_13208));
NAND2X1 g65528(.A (n_9428), .B (n_15111), .Y (n_13206));
INVX1 g65537(.A (n_11434), .Y (n_13205));
INVX1 g65539(.A (n_11433), .Y (n_13204));
NAND3X1 g65543(.A (n_9305), .B (n_7625), .C (n_13539), .Y (n_13203));
AOI21X1 g65553(.A0 (n_4461), .A1 (n_12652), .B0 (n_16466), .Y(n_13202));
AOI21X1 g65570(.A0 (n_5568), .A1 (n_12337), .B0 (n_20325), .Y(n_13201));
NAND2X1 g65583(.A (n_9312), .B (n_28692), .Y (n_13200));
NAND3X1 g65586(.A (n_10440), .B (n_8289), .C (n_4344), .Y (n_13199));
NAND3X1 g65593(.A (n_11492), .B (n_9380), .C (n_8009), .Y (n_13198));
INVX1 g65594(.A (n_11432), .Y (n_13197));
NAND3X1 g65599(.A (n_15009), .B (n_7002), .C (n_13195), .Y (n_13196));
AOI21X1 g65602(.A0 (n_3349), .A1 (n_10816), .B0 (n_13326), .Y(n_13194));
AOI21X1 g65606(.A0 (n_9004), .A1 (n_13192), .B0 (n_13318), .Y(n_13193));
AOI21X1 g65611(.A0 (n_9053), .A1 (n_13190), .B0 (n_10389), .Y(n_13191));
AOI21X1 g65614(.A0 (n_12385), .A1 (n_3456), .B0 (n_29102), .Y(n_13189));
AOI21X1 g65624(.A0 (n_11114), .A1 (n_9795), .B0 (n_26270), .Y(n_13188));
NAND2X1 g65625(.A (n_5490), .B (n_13186), .Y (n_13187));
NAND2X1 g65629(.A (n_5641), .B (n_13333), .Y (n_13185));
AOI21X1 g65630(.A0 (n_11655), .A1 (n_13183), .B0 (n_13804), .Y(n_13184));
AOI21X1 g65636(.A0 (n_27435), .A1 (n_13181), .B0 (n_29062), .Y(n_13182));
NAND3X1 g65647(.A (n_4269), .B (n_8670), .C (n_9796), .Y (n_13180));
INVX1 g65652(.A (n_11428), .Y (n_13179));
OAI21X1 g65657(.A0 (n_6828), .A1 (n_13177), .B0 (n_13176), .Y(n_13178));
NAND2X1 g65659(.A (n_9013), .B (n_15034), .Y (n_13175));
NAND2X1 g65674(.A (n_8309), .B (n_14996), .Y (n_13174));
NAND3X1 g65366(.A (n_13172), .B (n_5385), .C (n_13171), .Y (n_13173));
OAI21X1 g65696(.A0 (n_6818), .A1 (n_11662), .B0 (n_2362), .Y(n_13170));
NAND2X1 g65698(.A (n_7536), .B (n_13295), .Y (n_13169));
NAND2X1 g65700(.A (n_8779), .B (n_14909), .Y (n_13168));
AOI21X1 g65709(.A0 (n_13166), .A1 (n_11263), .B0 (n_29102), .Y(n_13167));
INVX1 g65726(.A (n_11426), .Y (n_13165));
NAND2X1 g65732(.A (n_5442), .B (n_13282), .Y (n_13164));
AOI21X1 g65734(.A0 (n_6762), .A1 (n_13162), .B0 (n_28692), .Y(n_13163));
NAND2X1 g65753(.A (n_4981), .B (n_13159), .Y (n_13160));
AOI21X1 g65758(.A0 (n_5668), .A1 (n_12370), .B0 (n_17500), .Y(n_13158));
NOR2X1 g65763(.A (n_5784), .B (n_13156), .Y (n_13157));
AOI21X1 g65771(.A0 (n_2665), .A1 (n_10914), .B0 (n_9527), .Y(n_13154));
NAND3X1 g65777(.A (n_13152), .B (n_11193), .C (n_8298), .Y (n_13153));
AOI21X1 g65778(.A0 (n_14399), .A1 (n_4554), .B0 (n_9106), .Y(n_13151));
OAI21X1 g65782(.A0 (n_6426), .A1 (n_6534), .B0 (n_13148), .Y(n_13149));
AOI21X1 g65787(.A0 (n_7290), .A1 (n_10687), .B0 (n_28375), .Y(n_13147));
INVX1 g65791(.A (n_11425), .Y (n_13146));
NAND3X1 g65794(.A (n_7870), .B (n_11381), .C (n_8167), .Y (n_13145));
AOI21X1 g65796(.A0 (n_13116), .A1 (n_8756), .B0 (n_17260), .Y(n_13144));
NAND3X1 g65799(.A (n_29208), .B (n_9190), .C (n_13142), .Y (n_13143));
OAI21X1 g65805(.A0 (n_8101), .A1 (n_14055), .B0 (n_14945), .Y(n_13141));
OR2X1 g65809(.A (n_9316), .B (n_15166), .Y (n_13140));
NAND2X1 g65812(.A (n_9375), .B (n_14757), .Y (n_13139));
NAND3X1 g65816(.A (n_13137), .B (n_11235), .C (n_5855), .Y (n_13138));
NAND2X1 g65817(.A (n_5387), .B (n_13357), .Y (n_13136));
AOI21X1 g65819(.A0 (n_13134), .A1 (n_4599), .B0 (n_12827), .Y(n_13135));
NAND2X1 g65823(.A (n_6141), .B (n_11579), .Y (n_13133));
OAI21X1 g65841(.A0 (n_29336), .A1 (n_1626), .B0 (n_8583), .Y(n_13132));
NAND2X1 g65862(.A (n_5888), .B (n_11558), .Y (n_13130));
AOI21X1 g65866(.A0 (n_4786), .A1 (n_16988), .B0 (n_11377), .Y(n_13129));
MX2X1 g65886(.A (n_7086), .B (n_16586), .S0 (n_11603), .Y (n_13128));
OAI21X1 g65891(.A0 (n_9350), .A1 (n_5151), .B0 (n_8360), .Y(n_13127));
OAI21X1 g65900(.A0 (n_8466), .A1 (n_28757), .B0 (n_5781), .Y(n_13126));
OAI21X1 g65901(.A0 (n_8768), .A1 (n_8910), .B0 (n_8264), .Y(n_13125));
OAI21X1 g65902(.A0 (n_9534), .A1 (n_10255), .B0 (n_5712), .Y(n_13124));
OAI21X1 g65907(.A0 (n_8515), .A1 (n_9500), .B0 (n_6108), .Y(n_13123));
AOI21X1 g65913(.A0 (n_9755), .A1 (n_2827), .B0 (n_9495), .Y(n_13122));
AOI21X1 g65922(.A0 (n_19114), .A1 (n_2929), .B0 (n_9394), .Y(n_13121));
MX2X1 g65942(.A (n_13119), .B (n_13118), .S0 (n_18266), .Y (n_13120));
MX2X1 g65943(.A (n_13116), .B (n_12734), .S0 (n_19791), .Y (n_13117));
OAI21X1 g65946(.A0 (n_13114), .A1 (n_9388), .B0 (n_9079), .Y(n_13115));
AND2X1 g65960(.A (n_8663), .B (n_11354), .Y (n_13113));
AOI21X1 g65961(.A0 (n_3669), .A1 (n_28340), .B0 (n_8100), .Y(n_28247));
AOI21X1 g65962(.A0 (n_6557), .A1 (n_12836), .B0 (n_8680), .Y(n_13110));
AND2X1 g65963(.A (n_6423), .B (n_8539), .Y (n_13109));
NAND2X1 g65966(.A (n_8480), .B (n_17567), .Y (n_13108));
AOI21X1 g65967(.A0 (n_6553), .A1 (n_14757), .B0 (n_7142), .Y(n_13107));
AOI21X1 g65970(.A0 (n_5224), .A1 (n_12571), .B0 (n_8420), .Y(n_13105));
INVX1 g65971(.A (n_11406), .Y (n_13104));
AOI21X1 g65977(.A0 (n_7642), .A1 (n_19226), .B0 (n_9321), .Y(n_13102));
NAND2X1 g65978(.A (n_7851), .B (n_14592), .Y (n_13101));
INVX1 g65983(.A (n_15626), .Y (n_28311));
INVX1 g65988(.A (n_11401), .Y (n_17235));
NAND2X1 g65995(.A (n_12154), .B (n_14592), .Y (n_13098));
NOR2X1 g65997(.A (n_18046), .B (n_13083), .Y (n_13097));
NAND4X1 g66003(.A (n_17500), .B (n_4093), .C (n_2231), .D (n_4681),.Y (n_19648));
NOR2X1 g66006(.A (n_9635), .B (n_14055), .Y (n_13095));
INVX1 g66009(.A (n_11395), .Y (n_19814));
INVX1 g66011(.A (n_11393), .Y (n_13094));
INVX1 g66015(.A (n_11391), .Y (n_14722));
INVX1 g66017(.A (n_13092), .Y (n_13093));
NAND2X1 g66020(.A (n_13073), .B (n_26491), .Y (n_13090));
OR2X1 g66021(.A (n_8774), .B (n_8637), .Y (n_15345));
OR2X1 g66022(.A (n_12275), .B (n_7598), .Y (n_15435));
INVX1 g66030(.A (n_11389), .Y (n_14719));
INVX1 g66037(.A (n_11388), .Y (n_16853));
INVX1 g66041(.A (n_13475), .Y (n_13087));
NAND2X1 g66045(.A (n_10603), .B (n_13466), .Y (n_18063));
AND2X1 g66048(.A (n_13063), .B (n_12169), .Y (n_15418));
NAND2X1 g66057(.A (n_10565), .B (n_11312), .Y (n_15230));
NAND2X1 g66063(.A (n_13083), .B (n_13082), .Y (n_13084));
INVX1 g66077(.A (n_13080), .Y (n_20003));
INVX1 g66078(.A (n_13080), .Y (n_13081));
NOR2X1 g66088(.A (n_11052), .B (n_25654), .Y (n_13079));
INVX1 g66090(.A (n_11379), .Y (n_15267));
INVX1 g66094(.A (n_13077), .Y (n_16941));
NAND2X1 g66100(.A (n_10144), .B (n_14866), .Y (n_17140));
INVX1 g66104(.A (n_11373), .Y (n_14709));
AND2X1 g66106(.A (n_13076), .B (n_14866), .Y (n_16572));
AND2X1 g66118(.A (n_10027), .B (n_17260), .Y (n_14707));
NAND2X1 g66123(.A (n_13073), .B (n_17571), .Y (n_13074));
NAND2X1 g66124(.A (n_12835), .B (n_11052), .Y (n_13072));
NAND2X1 g66126(.A (n_10185), .B (n_12169), .Y (n_17113));
INVX1 g66128(.A (n_13069), .Y (n_13071));
INVX1 g66139(.A (n_13067), .Y (n_15425));
INVX1 g66140(.A (n_13067), .Y (n_13068));
INVX1 g66142(.A (n_11359), .Y (n_16551));
NAND2X1 g66151(.A (n_10136), .B (n_12169), .Y (n_15313));
INVX1 g66157(.A (n_13066), .Y (n_14698));
AND2X1 g66161(.A (n_12895), .B (n_2779), .Y (n_14696));
INVX1 g66162(.A (n_11356), .Y (n_15414));
INVX1 g66165(.A (n_13064), .Y (n_13065));
NAND2X1 g66168(.A (n_9754), .B (n_29256), .Y (n_16323));
NAND2X1 g66169(.A (n_13063), .B (n_13083), .Y (n_18047));
NOR2X1 g66174(.A (n_27141), .B (n_5329), .Y (n_13062));
AND2X1 g66177(.A (n_27745), .B (n_16835), .Y (n_13060));
INVX1 g66185(.A (n_11346), .Y (n_14695));
INVX1 g66192(.A (n_13056), .Y (n_13058));
NAND2X1 g66198(.A (n_13003), .B (n_7201), .Y (n_13055));
INVX1 g66200(.A (n_13054), .Y (n_14692));
NAND2X1 g66203(.A (n_10046), .B (n_11312), .Y (n_16574));
NAND2X1 g66208(.A (n_13052), .B (n_13606), .Y (n_13053));
NAND2X1 g66212(.A (n_10332), .B (n_15894), .Y (n_18966));
INVX1 g66214(.A (n_14972), .Y (n_13051));
NAND2X1 g66221(.A (n_12997), .B (n_20325), .Y (n_13050));
INVX2 g66222(.A (n_13047), .Y (n_18587));
NOR2X1 g66231(.A (n_11517), .B (n_4582), .Y (n_13046));
NAND3X1 g66237(.A (n_4689), .B (n_5617), .C (n_9442), .Y (n_16645));
NOR2X1 g66239(.A (n_8288), .B (n_29102), .Y (n_13044));
NAND2X1 g66243(.A (n_9750), .B (n_7325), .Y (n_16775));
NAND2X1 g66248(.A (n_12893), .B (n_11300), .Y (n_15322));
INVX2 g66254(.A (n_11325), .Y (n_15091));
INVX1 g66256(.A (n_13042), .Y (n_13043));
NAND2X1 g66264(.A (n_12518), .B (n_17411), .Y (n_13039));
NAND3X1 g66266(.A (n_15411), .B (n_13037), .C (n_10094), .Y(n_18926));
INVX1 g66268(.A (n_13035), .Y (n_18000));
INVX1 g66269(.A (n_13035), .Y (n_13036));
AND2X1 g66273(.A (n_18369), .B (n_14858), .Y (n_13034));
NAND2X1 g66280(.A (n_12591), .B (n_28642), .Y (n_13033));
NAND2X1 g66282(.A (n_12161), .B (n_17567), .Y (n_13032));
OR2X1 g66285(.A (n_13031), .B (n_28375), .Y (n_15281));
INVX1 g66292(.A (n_11313), .Y (n_13030));
NAND2X1 g66297(.A (n_10747), .B (n_5558), .Y (n_17240));
INVX1 g66311(.A (n_11309), .Y (n_14679));
NAND3X1 g66315(.A (n_13804), .B (n_5602), .C (n_6185), .Y (n_13028));
NAND4X1 g66316(.A (n_10452), .B (n_8910), .C (n_2007), .D (n_5053),.Y (n_15151));
NAND2X1 g66318(.A (n_13026), .B (n_8452), .Y (n_13027));
INVX1 g66319(.A (n_17824), .Y (n_13025));
INVX1 g66323(.A (n_18801), .Y (n_13023));
INVX1 g66325(.A (n_13022), .Y (n_16595));
INVX1 g66327(.A (n_13020), .Y (n_17972));
OR2X1 g66331(.A (n_9134), .B (n_11300), .Y (n_14677));
INVX1 g66332(.A (n_13018), .Y (n_13019));
INVX1 g66341(.A (n_13015), .Y (n_13016));
NAND2X1 g66346(.A (n_12928), .B (n_9783), .Y (n_15140));
NAND3X1 g66353(.A (n_14484), .B (n_5349), .C (n_10031), .Y (n_15135));
INVX1 g66358(.A (n_11305), .Y (n_14674));
INVX1 g66364(.A (n_11303), .Y (n_14673));
AND2X1 g66367(.A (n_9764), .B (n_27688), .Y (n_14671));
NAND2X1 g66371(.A (n_9977), .B (n_13571), .Y (n_13013));
NOR2X1 g66374(.A (n_9179), .B (n_12019), .Y (n_13012));
NAND2X1 g72360(.A (n_6750), .B (n_16973), .Y (n_13011));
NOR2X1 g66378(.A (n_15132), .B (n_12019), .Y (n_13010));
INVX1 g66383(.A (n_13008), .Y (n_17197));
NOR2X1 g66388(.A (n_15705), .B (n_14142), .Y (n_13006));
NOR3X1 g66390(.A (n_13804), .B (n_9708), .C (n_6583), .Y (n_13005));
NAND2X1 g66392(.A (n_13003), .B (n_17567), .Y (n_13004));
NAND2X1 g66393(.A (n_12570), .B (n_7201), .Y (n_13002));
NOR4X1 g66396(.A (n_26270), .B (n_2548), .C (n_2592), .D (n_1707), .Y(n_13000));
NAND2X1 g66397(.A (n_12997), .B (n_15388), .Y (n_12998));
INVX1 g66398(.A (n_12995), .Y (n_12996));
INVX1 g66400(.A (n_11299), .Y (n_12994));
INVX1 g66402(.A (n_12991), .Y (n_12993));
INVX1 g66409(.A (n_12990), .Y (n_16670));
INVX1 g66416(.A (n_12988), .Y (n_18050));
INVX1 g66417(.A (n_12988), .Y (n_12989));
INVX1 g66421(.A (n_11291), .Y (n_15116));
INVX1 g66430(.A (n_11284), .Y (n_20023));
NAND2X1 g66432(.A (n_13942), .B (n_12986), .Y (n_12987));
INVX1 g66433(.A (n_11282), .Y (n_12985));
INVX1 g66438(.A (n_11281), .Y (n_14663));
INVX1 g66441(.A (n_12983), .Y (n_12984));
NAND2X1 g66444(.A (n_12980), .B (n_12979), .Y (n_12981));
OR2X1 g66451(.A (n_18264), .B (n_17500), .Y (n_14661));
AOI21X1 g68649(.A0 (n_5008), .A1 (n_14055), .B0 (n_9112), .Y(n_12977));
NAND2X1 g66459(.A (n_10152), .B (n_9264), .Y (n_16532));
NOR2X1 g66461(.A (n_12973), .B (n_29074), .Y (n_12974));
NAND2X1 g66468(.A (n_12945), .B (n_4689), .Y (n_12972));
NAND2X1 g66470(.A (n_12970), .B (n_9106), .Y (n_12971));
INVX1 g66473(.A (n_12968), .Y (n_15404));
INVX1 g66474(.A (n_12968), .Y (n_12969));
NAND2X1 g66478(.A (n_11897), .B (n_26877), .Y (n_16325));
NAND2X1 g66479(.A (n_13026), .B (n_15411), .Y (n_12966));
OR2X1 g66482(.A (n_8874), .B (n_15411), .Y (n_14655));
INVX1 g66484(.A (n_11273), .Y (n_15076));
NAND2X1 g66487(.A (n_12964), .B (n_12019), .Y (n_12965));
NAND3X1 g66489(.A (n_11272), .B (n_8024), .C (n_8093), .Y (n_15064));
INVX1 g66492(.A (n_11271), .Y (n_16674));
NAND2X1 g66497(.A (n_10314), .B (n_13326), .Y (n_12963));
NOR2X1 g66504(.A (n_14055), .B (n_16601), .Y (n_14649));
NAND2X1 g66513(.A (n_9125), .B (n_27099), .Y (n_12959));
INVX1 g66516(.A (n_14961), .Y (n_12958));
INVX1 g66522(.A (n_12957), .Y (n_14647));
NAND2X1 g66524(.A (n_10862), .B (n_14589), .Y (n_18249));
INVX1 g66525(.A (n_11262), .Y (n_12955));
AND2X1 g66529(.A (n_18920), .B (n_11385), .Y (n_14646));
INVX1 g66531(.A (n_11260), .Y (n_15302));
AND2X1 g66534(.A (n_10882), .B (n_28642), .Y (n_14643));
NOR2X1 g66537(.A (n_10174), .B (n_5558), .Y (n_14641));
NAND2X1 g66538(.A (n_12175), .B (n_28642), .Y (n_12953));
NAND2X1 g66543(.A (n_12980), .B (n_15986), .Y (n_12952));
NAND2X1 g66551(.A (n_10644), .B (n_10389), .Y (n_12950));
OR2X1 g66552(.A (n_27412), .B (n_15039), .Y (n_19711));
INVX1 g66553(.A (n_11254), .Y (n_15304));
NAND2X1 g66560(.A (n_12945), .B (n_29074), .Y (n_12946));
NAND3X1 g66561(.A (n_18266), .B (n_13875), .C (n_10146), .Y(n_18948));
NAND2X1 g66562(.A (n_29173), .B (n_14026), .Y (n_12944));
NAND2X1 g66568(.A (n_28136), .B (n_8928), .Y (n_12943));
NAND2X1 g66569(.A (n_9781), .B (n_7498), .Y (n_16368));
AND2X1 g66570(.A (n_12964), .B (n_28692), .Y (n_12941));
NOR2X1 g66572(.A (n_26464), .B (n_28642), .Y (n_14638));
INVX1 g66577(.A (n_12939), .Y (n_14636));
NAND2X1 g66586(.A (n_10489), .B (n_14155), .Y (n_18244));
INVX1 g66587(.A (n_12938), .Y (n_15272));
NOR2X1 g66593(.A (n_9146), .B (n_29065), .Y (n_14633));
INVX1 g66595(.A (n_27964), .Y (n_12937));
INVX1 g66605(.A (n_12934), .Y (n_18582));
INVX1 g66606(.A (n_12934), .Y (n_12935));
INVX1 g66624(.A (n_11238), .Y (n_12932));
NAND2X1 g66626(.A (n_12409), .B (n_9486), .Y (n_12931));
NAND2X1 g66628(.A (n_10463), .B (n_9819), .Y (n_12930));
NOR2X1 g66630(.A (n_8621), .B (n_14155), .Y (n_12929));
NAND2X1 g66632(.A (n_12928), .B (n_27688), .Y (n_16588));
INVX1 g66633(.A (n_12926), .Y (n_16637));
INVX1 g66638(.A (n_12925), .Y (n_14621));
INVX1 g66640(.A (n_11231), .Y (n_18641));
INVX1 g66646(.A (n_12923), .Y (n_12924));
INVX1 g66654(.A (n_11227), .Y (n_14619));
INVX1 g66657(.A (n_12922), .Y (n_15328));
NAND2X1 g66659(.A (n_10471), .B (n_18266), .Y (n_16537));
INVX1 g66660(.A (n_11224), .Y (n_12920));
NOR2X1 g66663(.A (n_12918), .B (n_12917), .Y (n_12919));
NOR2X1 g66672(.A (n_20078), .B (n_13466), .Y (n_12916));
NAND2X1 g66673(.A (n_28834), .B (n_13593), .Y (n_16331));
INVX1 g66674(.A (n_11222), .Y (n_19811));
NAND2X1 g66676(.A (n_12362), .B (n_27688), .Y (n_12914));
AND2X1 g66682(.A (n_9068), .B (n_8679), .Y (n_15299));
INVX1 g66683(.A (n_11219), .Y (n_19243));
INVX1 g66691(.A (n_14956), .Y (n_12912));
NAND2X1 g66694(.A (n_8806), .B (n_12910), .Y (n_12911));
NAND2X1 g66697(.A (n_10819), .B (n_13593), .Y (n_17031));
INVX1 g66698(.A (n_11217), .Y (n_12909));
NAND2X1 g66703(.A (n_10014), .B (n_14484), .Y (n_15886));
NAND2X2 g66711(.A (n_8818), .B (n_18785), .Y (n_16559));
INVX1 g66715(.A (n_11214), .Y (n_17315));
NAND2X1 g66717(.A (n_10841), .B (n_10599), .Y (n_16557));
OR2X1 g66719(.A (n_12907), .B (n_16434), .Y (n_14603));
INVX1 g66720(.A (n_12906), .Y (n_15195));
INVX2 g66726(.A (n_11213), .Y (n_16540));
INVX1 g66734(.A (n_12903), .Y (n_17982));
AND2X1 g66738(.A (n_10260), .B (n_7410), .Y (n_15266));
OR2X1 g66740(.A (n_10096), .B (n_15894), .Y (n_17310));
INVX1 g66745(.A (n_11209), .Y (n_12902));
NAND2X1 g66747(.A (n_10431), .B (n_28692), .Y (n_17121));
INVX1 g66752(.A (n_11208), .Y (n_15392));
INVX2 g66755(.A (n_12900), .Y (n_18648));
INVX1 g66759(.A (n_11206), .Y (n_15342));
INVX2 g66768(.A (n_12898), .Y (n_20392));
NAND2X1 g66772(.A (n_10323), .B (n_12896), .Y (n_25463));
NAND2X1 g66773(.A (n_12895), .B (n_11354), .Y (n_18060));
NOR2X1 g66776(.A (n_8152), .B (n_29269), .Y (n_12894));
INVX1 g66785(.A (n_11199), .Y (n_15902));
NAND2X1 g66787(.A (n_12893), .B (n_29256), .Y (n_15278));
INVX1 g66790(.A (n_11196), .Y (n_16321));
INVX1 g66794(.A (n_11194), .Y (n_18619));
OR2X1 g66797(.A (n_12892), .B (n_18785), .Y (n_16519));
INVX1 g66802(.A (n_11191), .Y (n_14588));
NAND2X1 g73070(.A (n_7376), .B (n_5140), .Y (n_12890));
INVX1 g66807(.A (n_11189), .Y (n_14587));
NAND2X2 g66811(.A (n_10447), .B (n_28433), .Y (n_16711));
INVX1 g66814(.A (n_11188), .Y (n_16510));
INVX1 g66818(.A (n_13431), .Y (n_12887));
NAND2X1 g66828(.A (n_13257), .B (n_8335), .Y (n_12886));
NOR2X1 g66832(.A (n_12885), .B (n_8637), .Y (n_15360));
NAND2X1 g66834(.A (n_5418), .B (n_7266), .Y (n_15358));
NAND2X1 g66838(.A (n_8546), .B (n_12883), .Y (n_12884));
NOR2X1 g66843(.A (n_12881), .B (n_5762), .Y (n_12882));
INVX1 g66848(.A (n_12879), .Y (n_12880));
NAND2X1 g66850(.A (n_10633), .B (n_18205), .Y (n_17064));
NAND2X1 g66852(.A (n_4172), .B (n_12754), .Y (n_12877));
INVX1 g66858(.A (n_13516), .Y (n_12873));
NAND2X1 g66865(.A (n_8877), .B (n_12870), .Y (n_12871));
NAND2X1 g66867(.A (n_6900), .B (n_12868), .Y (n_12869));
INVX1 g66880(.A (n_12865), .Y (n_14573));
INVX1 g66882(.A (n_18335), .Y (n_12864));
INVX1 g66894(.A (n_12862), .Y (n_16334));
NOR2X1 g66900(.A (n_8077), .B (n_5678), .Y (n_12861));
NAND2X1 g66904(.A (n_4588), .B (n_11052), .Y (n_12860));
NAND2X1 g66905(.A (n_12858), .B (n_8088), .Y (n_12859));
INVX1 g66909(.A (n_18645), .Y (n_14567));
NAND2X1 g66914(.A (n_7600), .B (n_14080), .Y (n_12857));
NAND2X1 g66918(.A (n_12563), .B (n_16539), .Y (n_12856));
INVX1 g66924(.A (n_12853), .Y (n_12854));
NOR2X1 g66930(.A (n_12852), .B (n_9118), .Y (n_14564));
NAND2X1 g66933(.A (n_8725), .B (n_17377), .Y (n_12851));
NOR2X1 g66936(.A (n_10475), .B (n_12850), .Y (n_14561));
NOR2X1 g66939(.A (n_10609), .B (n_12849), .Y (n_14559));
NOR2X1 g66942(.A (n_7067), .B (n_18254), .Y (n_12848));
INVX1 g66955(.A (n_12846), .Y (n_12847));
NAND2X1 g66960(.A (n_12844), .B (n_12643), .Y (n_12845));
NOR2X1 g66961(.A (n_3040), .B (n_8567), .Y (n_12843));
AND2X1 g66979(.A (n_12781), .B (n_27445), .Y (n_12840));
AND2X1 g66980(.A (n_12638), .B (n_13083), .Y (n_12838));
NAND2X1 g66981(.A (n_12836), .B (n_12835), .Y (n_18937));
INVX1 g66982(.A (n_12833), .Y (n_12834));
NAND2X1 g66991(.A (n_6078), .B (n_8997), .Y (n_17292));
NAND2X1 g66999(.A (n_15315), .B (n_12285), .Y (n_12831));
AND2X1 g67000(.A (n_8117), .B (n_27604), .Y (n_12830));
OR2X1 g67004(.A (n_12828), .B (n_12827), .Y (n_12829));
NOR2X1 g67011(.A (n_12823), .B (n_12822), .Y (n_12824));
NOR2X1 g67017(.A (n_13073), .B (n_26489), .Y (n_12819));
NAND2X1 g67020(.A (n_9759), .B (n_18237), .Y (n_12818));
INVX1 g67022(.A (n_13542), .Y (n_12817));
NAND2X1 g67027(.A (n_12815), .B (n_11576), .Y (n_12816));
INVX1 g67028(.A (n_12813), .Y (n_12814));
NAND2X1 g67034(.A (n_13260), .B (n_8273), .Y (n_12811));
OR2X1 g67039(.A (n_27424), .B (n_7547), .Y (n_12810));
INVX1 g67045(.A (n_12807), .Y (n_12806));
INVX1 g67053(.A (n_11123), .Y (n_12805));
NAND2X1 g67055(.A (n_13602), .B (n_9410), .Y (n_20096));
NAND2X1 g67057(.A (n_12803), .B (n_12802), .Y (n_12804));
NOR2X1 g67060(.A (n_9388), .B (n_12801), .Y (n_15291));
NAND2X1 g67062(.A (n_5656), .B (n_7786), .Y (n_12800));
NAND2X1 g67064(.A (n_12828), .B (n_10485), .Y (n_12798));
AND2X1 g67071(.A (n_7324), .B (n_12681), .Y (n_12797));
NOR2X1 g67075(.A (n_10206), .B (n_9230), .Y (n_12796));
NOR2X1 g67076(.A (n_17017), .B (n_15705), .Y (n_12795));
NAND2X1 g67077(.A (n_6341), .B (n_12649), .Y (n_12794));
NAND2X1 g67086(.A (n_8157), .B (n_12788), .Y (n_12789));
OAI21X1 g67092(.A0 (n_3060), .A1 (n_2239), .B0 (n_12786), .Y(n_12787));
AOI21X1 g67095(.A0 (n_5196), .A1 (n_10130), .B0 (n_15574), .Y(n_12785));
NAND2X1 g67098(.A (n_12784), .B (n_13609), .Y (n_16661));
NAND2X1 g67103(.A (n_7257), .B (n_8152), .Y (n_12783));
NAND2X1 g67105(.A (n_4761), .B (n_12781), .Y (n_12782));
NAND2X1 g67113(.A (n_12779), .B (n_12778), .Y (n_12780));
NAND2X1 g67114(.A (n_10321), .B (n_17864), .Y (n_15226));
INVX1 g67124(.A (n_12776), .Y (n_12777));
INVX1 g67128(.A (n_12774), .Y (n_12775));
INVX1 g67130(.A (n_12772), .Y (n_12773));
NOR2X1 g67132(.A (n_5033), .B (n_8155), .Y (n_12771));
NAND2X1 g67139(.A (n_12768), .B (n_15187), .Y (n_12769));
NAND2X1 g67140(.A (n_10351), .B (n_11576), .Y (n_16680));
NAND2X1 g67141(.A (n_26034), .B (n_11510), .Y (n_12767));
NOR2X1 g67142(.A (n_8498), .B (n_12480), .Y (n_12765));
NAND2X1 g67149(.A (n_6003), .B (n_12169), .Y (n_17302));
NAND2X1 g67153(.A (n_15640), .B (n_12762), .Y (n_12763));
INVX1 g67157(.A (n_11089), .Y (n_12761));
AND2X1 g67159(.A (n_10035), .B (n_12760), .Y (n_16582));
AND2X1 g67161(.A (n_11810), .B (n_7444), .Y (n_12759));
NOR2X1 g67162(.A (n_10548), .B (n_12756), .Y (n_29307));
NAND2X1 g67163(.A (n_10957), .B (n_12754), .Y (n_12755));
NAND2X1 g67165(.A (n_12752), .B (n_12751), .Y (n_12753));
NAND2X1 g67168(.A (n_10566), .B (n_6534), .Y (n_15254));
AND2X1 g67169(.A (n_15588), .B (n_13082), .Y (n_18630));
AND2X1 g67170(.A (n_12373), .B (n_6408), .Y (n_12750));
NOR2X1 g67173(.A (n_12748), .B (n_12747), .Y (n_12749));
INVX1 g67176(.A (n_12745), .Y (n_12746));
OR2X1 g67182(.A (n_12740), .B (n_4582), .Y (n_12741));
INVX1 g67183(.A (n_12739), .Y (n_15423));
INVX1 g67186(.A (n_11081), .Y (n_12738));
NOR2X1 g67188(.A (n_11517), .B (n_17020), .Y (n_12737));
NAND2X1 g67189(.A (n_12735), .B (n_12734), .Y (n_12736));
INVX1 g67198(.A (n_11077), .Y (n_14503));
AND2X1 g67204(.A (n_10198), .B (n_17500), .Y (n_12733));
OR2X1 g67205(.A (n_12731), .B (n_16290), .Y (n_12732));
NOR2X1 g67210(.A (n_10549), .B (n_15894), .Y (n_12730));
OAI21X1 g67211(.A0 (n_2843), .A1 (n_2959), .B0 (n_11520), .Y(n_12728));
AOI21X1 g67219(.A0 (n_4367), .A1 (n_10030), .B0 (n_12228), .Y(n_12727));
NAND2X1 g67225(.A (n_12723), .B (n_12722), .Y (n_12724));
OR2X1 g67227(.A (n_12720), .B (n_27643), .Y (n_12721));
NAND2X1 g67233(.A (n_12718), .B (n_5806), .Y (n_12719));
NAND2X1 g67237(.A (n_12634), .B (n_16052), .Y (n_14489));
NOR2X1 g67239(.A (n_9955), .B (n_12140), .Y (n_12717));
NOR2X1 g67241(.A (n_8456), .B (n_12715), .Y (n_12716));
OR2X1 g67242(.A (n_12713), .B (n_18369), .Y (n_12714));
NAND2X1 g67245(.A (n_8650), .B (n_9509), .Y (n_12712));
NAND2X1 g67248(.A (n_6047), .B (n_3318), .Y (n_16503));
AND2X1 g67250(.A (n_19226), .B (n_14858), .Y (n_17522));
OR2X1 g67255(.A (n_14080), .B (n_11052), .Y (n_12710));
NAND2X1 g67258(.A (n_4133), .B (n_7201), .Y (n_12709));
AND2X1 g67259(.A (n_5436), .B (n_13466), .Y (n_16469));
NOR2X1 g67263(.A (n_8669), .B (n_28812), .Y (n_12708));
NOR2X1 g67275(.A (n_8323), .B (n_4860), .Y (n_12707));
INVX1 g67284(.A (n_12705), .Y (n_12706));
NAND2X1 g67288(.A (n_8984), .B (n_5832), .Y (n_12703));
NAND2X1 g67292(.A (n_10610), .B (n_10693), .Y (n_12702));
NAND2X1 g67295(.A (n_5861), .B (n_9368), .Y (n_12701));
NAND2X1 g67296(.A (n_10044), .B (n_11276), .Y (n_12699));
NAND2X1 g67304(.A (n_6020), .B (n_27434), .Y (n_16634));
INVX1 g67305(.A (n_12697), .Y (n_12698));
INVX1 g67312(.A (n_21164), .Y (n_12696));
NOR2X1 g67316(.A (n_4466), .B (n_8661), .Y (n_12695));
INVX1 g67320(.A (n_11050), .Y (n_15319));
INVX1 g67324(.A (n_11524), .Y (n_12694));
NAND2X1 g67328(.A (n_12691), .B (n_13118), .Y (n_12692));
NOR2X1 g67332(.A (n_9406), .B (n_3386), .Y (n_15638));
NAND2X1 g67333(.A (n_17706), .B (n_6197), .Y (n_16828));
NAND2X1 g67336(.A (n_8858), .B (n_5600), .Y (n_15190));
AOI21X1 g67337(.A0 (n_4392), .A1 (n_28134), .B0 (n_12402), .Y(n_12688));
NOR2X1 g67342(.A (n_9905), .B (n_12604), .Y (n_12686));
AND2X1 g67347(.A (n_10204), .B (n_11312), .Y (n_14450));
NAND2X1 g67364(.A (n_12681), .B (n_12680), .Y (n_12682));
NAND2X1 g67366(.A (n_6057), .B (n_8679), .Y (n_16501));
INVX1 g67367(.A (n_13411), .Y (n_12678));
NAND2X1 g67373(.A (n_10478), .B (n_6790), .Y (n_16724));
NOR2X1 g67376(.A (n_6126), .B (n_15674), .Y (n_12677));
NAND2X1 g67379(.A (n_3626), .B (n_6202), .Y (n_12676));
NAND2X1 g67389(.A (n_11029), .B (n_12781), .Y (n_12675));
AOI21X1 g65381(.A0 (n_12673), .A1 (n_8822), .B0 (n_15674), .Y(n_12674));
INVX1 g67393(.A (n_11041), .Y (n_12672));
NOR2X1 g67395(.A (n_7876), .B (n_15166), .Y (n_12671));
NAND2X1 g67396(.A (n_7566), .B (n_14126), .Y (n_12670));
NAND2X1 g67401(.A (n_5913), .B (n_17411), .Y (n_12669));
INVX1 g67402(.A (n_12667), .Y (n_12668));
OR2X1 g67404(.A (n_12349), .B (n_15776), .Y (n_12666));
NAND2X1 g67413(.A (n_12664), .B (n_12663), .Y (n_12665));
AND2X1 g67418(.A (n_11135), .B (n_18369), .Y (n_12662));
NOR2X1 g67421(.A (n_9882), .B (n_7680), .Y (n_12661));
INVX1 g67424(.A (n_11028), .Y (n_14437));
INVX1 g67433(.A (n_11023), .Y (n_14431));
AOI21X1 g67435(.A0 (n_3494), .A1 (n_8090), .B0 (n_12316), .Y(n_12660));
NAND2X1 g67436(.A (n_5743), .B (n_28037), .Y (n_15170));
NAND2X1 g67440(.A (n_12189), .B (n_5514), .Y (n_12658));
NAND2X1 g67442(.A (n_8555), .B (n_933), .Y (n_12657));
AND2X1 g67444(.A (n_5779), .B (n_12655), .Y (n_12656));
NAND2X1 g67450(.A (n_6117), .B (n_11835), .Y (n_12654));
NAND2X1 g67451(.A (n_10561), .B (n_12652), .Y (n_12653));
AND2X1 g67453(.A (n_12649), .B (n_12648), .Y (n_12650));
NAND2X1 g67455(.A (n_8800), .B (n_15776), .Y (n_12647));
NOR2X1 g67457(.A (n_20078), .B (n_17023), .Y (n_12646));
NAND2X1 g67460(.A (n_12644), .B (n_12643), .Y (n_12645));
INVX1 g67461(.A (n_12641), .Y (n_12642));
NAND2X1 g67469(.A (n_10618), .B (n_13593), .Y (n_12640));
NOR2X1 g67472(.A (n_12638), .B (n_12637), .Y (n_12639));
OR2X1 g67473(.A (n_7470), .B (n_15568), .Y (n_12636));
INVX1 g72284(.A (n_12635), .Y (n_17048));
NAND2X1 g67477(.A (n_12634), .B (n_14592), .Y (n_15586));
NAND2X1 g67483(.A (n_7504), .B (n_7832), .Y (n_18393));
NAND2X1 g67485(.A (n_12632), .B (n_12631), .Y (n_12633));
NAND2X1 g67490(.A (n_12629), .B (n_12628), .Y (n_12630));
NAND2X1 g67491(.A (n_12626), .B (n_10795), .Y (n_12627));
AND2X1 g67494(.A (n_8984), .B (n_12564), .Y (n_12625));
NAND2X1 g67495(.A (n_12624), .B (n_6202), .Y (n_16865));
NAND2X1 g67501(.A (n_10451), .B (n_4582), .Y (n_12620));
AND2X1 g67519(.A (n_3967), .B (n_9418), .Y (n_12612));
INVX1 g67520(.A (n_12609), .Y (n_16426));
INVX1 g67521(.A (n_12609), .Y (n_12610));
AND2X1 g67523(.A (n_12607), .B (n_13376), .Y (n_25622));
INVX1 g67542(.A (n_12605), .Y (n_16406));
NAND2X1 g72998(.A (n_12604), .B (n_11322), .Y (n_13744));
NAND2X1 g67547(.A (n_12885), .B (n_27483), .Y (n_12603));
NAND2X1 g67550(.A (n_7956), .B (n_15067), .Y (n_12601));
NOR2X1 g67560(.A (n_12597), .B (n_28692), .Y (n_12598));
NAND2X1 g67564(.A (n_29198), .B (n_12594), .Y (n_12596));
AOI21X1 g67567(.A0 (n_5251), .A1 (n_10140), .B0 (n_16787), .Y(n_12593));
NOR2X1 g67568(.A (n_10542), .B (n_12591), .Y (n_12592));
INVX1 g67569(.A (n_12589), .Y (n_16543));
NAND2X1 g67573(.A (n_7226), .B (n_12587), .Y (n_12588));
AND2X1 g67577(.A (n_8119), .B (n_18320), .Y (n_12586));
NAND2X1 g67588(.A (n_12581), .B (n_12309), .Y (n_12582));
NAND2X1 g67590(.A (n_8805), .B (n_12578), .Y (n_12580));
NOR2X1 g67600(.A (n_9258), .B (n_9933), .Y (n_28880));
NAND2X1 g67601(.A (n_12162), .B (n_27671), .Y (n_16642));
INVX1 g67603(.A (n_10991), .Y (n_12576));
NAND2X2 g67611(.A (n_12495), .B (n_2260), .Y (n_14372));
INVX1 g67612(.A (n_12573), .Y (n_28264));
INVX1 g67615(.A (n_12572), .Y (n_14370));
NAND2X1 g67617(.A (n_12571), .B (n_12570), .Y (n_18922));
NAND2X1 g67619(.A (n_12568), .B (n_9113), .Y (n_12569));
NAND2X1 g67621(.A (n_12495), .B (n_6406), .Y (n_14367));
NAND2X2 g72986(.A (n_11902), .B (n_13991), .Y (n_13745));
INVX1 g67623(.A (n_12566), .Y (n_12567));
NAND2X1 g67625(.A (n_12564), .B (n_12563), .Y (n_12565));
NAND2X1 g67632(.A (n_10909), .B (n_12649), .Y (n_12562));
OR2X1 g67639(.A (n_12560), .B (n_12559), .Y (n_12561));
AND2X1 g67641(.A (n_9182), .B (n_26726), .Y (n_12558));
NAND2X1 g67642(.A (n_13609), .B (n_15776), .Y (n_16412));
NAND2X1 g67647(.A (n_10509), .B (n_28686), .Y (n_17035));
NOR2X1 g67652(.A (n_7498), .B (n_14981), .Y (n_14353));
NAND2X1 g67654(.A (n_10524), .B (n_28381), .Y (n_16672));
NOR2X1 g67656(.A (n_12555), .B (n_8223), .Y (n_12556));
AND2X1 g67678(.A (n_12549), .B (n_12560), .Y (n_12550));
NAND2X1 g67679(.A (n_29000), .B (n_12546), .Y (n_12548));
INVX1 g67687(.A (n_12544), .Y (n_12545));
NAND2X1 g67689(.A (n_5994), .B (n_10452), .Y (n_16650));
NAND2X1 g67693(.A (n_8936), .B (n_4898), .Y (n_12542));
OR2X1 g67700(.A (n_12541), .B (n_18168), .Y (n_15101));
NAND2X1 g67704(.A (n_5024), .B (n_15776), .Y (n_12538));
INVX1 g67708(.A (n_12535), .Y (n_12536));
NAND2X1 g67710(.A (n_10413), .B (n_14055), .Y (n_15098));
INVX1 g67717(.A (n_12533), .Y (n_12534));
INVX1 g67727(.A (n_12531), .Y (n_12532));
NOR2X1 g67731(.A (n_10501), .B (n_14099), .Y (n_12530));
OR2X1 g67734(.A (n_14126), .B (n_28037), .Y (n_12529));
NOR2X1 g67736(.A (n_12416), .B (n_29102), .Y (n_14327));
NOR2X1 g67750(.A (n_8996), .B (n_5783), .Y (n_12528));
NAND2X1 g67755(.A (n_4983), .B (n_9368), .Y (n_16639));
NOR2X1 g67767(.A (n_3922), .B (n_8459), .Y (n_12527));
NAND2X1 g67772(.A (n_5066), .B (n_12019), .Y (n_12526));
INVX1 g67776(.A (n_12524), .Y (n_19218));
NAND2X2 g67786(.A (n_6119), .B (n_9942), .Y (n_16683));
INVX2 g67791(.A (n_10949), .Y (n_16398));
NAND2X1 g67793(.A (n_7722), .B (n_11311), .Y (n_12521));
NAND2X1 g67799(.A (n_12187), .B (n_13472), .Y (n_12520));
NOR2X1 g67805(.A (n_12518), .B (n_12517), .Y (n_29408));
OR2X1 g67807(.A (n_9172), .B (n_8861), .Y (n_12516));
INVX1 g67808(.A (n_12514), .Y (n_12515));
INVX1 g67811(.A (n_12512), .Y (n_12513));
NAND2X1 g67828(.A (n_5991), .B (n_15388), .Y (n_12509));
NAND2X1 g67830(.A (n_7036), .B (n_13722), .Y (n_12508));
NAND2X1 g67834(.A (n_12506), .B (n_12505), .Y (n_12507));
NAND2X1 g67836(.A (n_8935), .B (n_11102), .Y (n_12504));
NAND2X1 g67838(.A (n_10959), .B (n_13376), .Y (n_12503));
NOR2X1 g67851(.A (n_18046), .B (n_18100), .Y (n_12502));
INVX1 g67854(.A (n_10930), .Y (n_14277));
AND2X1 g67862(.A (n_12754), .B (n_12500), .Y (n_12501));
NAND2X1 g67867(.A (n_8049), .B (n_9179), .Y (n_12499));
NOR2X1 g67868(.A (n_12127), .B (n_9874), .Y (n_12498));
NOR2X1 g67873(.A (n_4402), .B (n_12496), .Y (n_12497));
NAND2X1 g67879(.A (n_9914), .B (n_12495), .Y (n_16618));
NAND2X1 g67886(.A (n_8314), .B (n_9472), .Y (n_12493));
NAND2X1 g67895(.A (n_27671), .B (n_14624), .Y (n_15580));
NAND2X1 g67898(.A (n_27411), .B (n_7126), .Y (n_16625));
AND2X1 g67907(.A (n_2606), .B (n_7592), .Y (n_12488));
NAND2X1 g67908(.A (n_12486), .B (n_12375), .Y (n_12487));
OR2X1 g67912(.A (n_12484), .B (n_13606), .Y (n_12485));
NAND2X1 g67920(.A (n_9869), .B (n_26670), .Y (n_12483));
NAND2X1 g67921(.A (n_16973), .B (n_12480), .Y (n_12481));
NOR2X1 g67924(.A (n_7173), .B (n_17912), .Y (n_14244));
AND2X1 g67925(.A (n_12478), .B (n_5155), .Y (n_12479));
INVX1 g67929(.A (n_12476), .Y (n_12477));
NOR2X1 g72953(.A (n_10160), .B (n_11734), .Y (n_13748));
AND2X1 g67934(.A (n_12597), .B (n_15132), .Y (n_12475));
NAND2X1 g67935(.A (n_12397), .B (n_17884), .Y (n_12474));
NAND2X1 g67936(.A (n_12472), .B (n_28427), .Y (n_12473));
NAND2X1 g67940(.A (n_10429), .B (n_12019), .Y (n_12471));
AOI21X1 g67944(.A0 (n_3331), .A1 (n_12469), .B0 (n_12468), .Y(n_12470));
NOR2X1 g67948(.A (n_7243), .B (n_12129), .Y (n_12467));
INVX1 g67949(.A (n_12465), .Y (n_12466));
NOR2X1 g67952(.A (n_5864), .B (n_12410), .Y (n_12463));
NAND3X1 g67953(.A (n_9804), .B (n_6673), .C (n_4393), .Y (n_12462));
INVX1 g67955(.A (n_10902), .Y (n_12461));
NOR2X1 g67961(.A (n_15187), .B (n_28375), .Y (n_12460));
NOR2X1 g67965(.A (n_4687), .B (n_8422), .Y (n_12459));
NOR2X1 g67970(.A (n_7347), .B (n_17912), .Y (n_12457));
AND2X1 g67984(.A (n_12451), .B (n_15285), .Y (n_12452));
INVX1 g67987(.A (n_10896), .Y (n_14227));
NOR2X1 g67989(.A (n_9632), .B (n_4196), .Y (n_12450));
AND2X1 g67992(.A (n_5312), .B (n_12448), .Y (n_12449));
NAND2X1 g67995(.A (n_12446), .B (n_10199), .Y (n_12447));
NOR2X1 g67996(.A (n_12638), .B (n_7744), .Y (n_12445));
NAND2X1 g68005(.A (n_5048), .B (n_4898), .Y (n_12444));
NAND2X1 g68013(.A (n_10150), .B (n_9486), .Y (n_12443));
INVX1 g68014(.A (n_10887), .Y (n_12441));
NAND2X1 g68017(.A (n_1378), .B (n_6197), .Y (n_12440));
AND2X1 g68029(.A (n_10506), .B (n_10921), .Y (n_12439));
NOR3X1 g68030(.A (n_17912), .B (n_27225), .C (n_5503), .Y (n_12438));
NAND2X1 g68033(.A (n_12436), .B (n_9487), .Y (n_12437));
AOI21X1 g68035(.A0 (n_3173), .A1 (n_26880), .B0 (n_12389), .Y(n_12435));
NOR2X1 g68036(.A (n_4517), .B (n_13609), .Y (n_12433));
NAND2X1 g68037(.A (n_27483), .B (n_14286), .Y (n_12432));
NAND2X1 g68048(.A (n_15961), .B (n_29062), .Y (n_17416));
NAND2X1 g68050(.A (n_12429), .B (n_27483), .Y (n_12430));
NOR2X1 g68051(.A (n_13003), .B (n_28045), .Y (n_12428));
INVX1 g68052(.A (n_14765), .Y (n_12427));
OR2X1 g68055(.A (n_18882), .B (n_14026), .Y (n_12426));
INVX1 g68064(.A (n_10874), .Y (n_12425));
INVX1 g68066(.A (n_10871), .Y (n_12424));
NAND2X1 g68068(.A (n_8259), .B (n_8708), .Y (n_12423));
AOI21X1 g68070(.A0 (n_4321), .A1 (n_9939), .B0 (n_15039), .Y(n_12422));
NOR2X1 g68071(.A (n_12420), .B (n_11197), .Y (n_12421));
NAND2X1 g68072(.A (n_27708), .B (n_12448), .Y (n_25827));
NOR2X1 g68073(.A (n_29205), .B (n_28156), .Y (n_12418));
NOR2X1 g68079(.A (n_12416), .B (n_9442), .Y (n_12417));
NAND2X1 g68083(.A (n_9906), .B (n_12868), .Y (n_12413));
NAND2X1 g68085(.A (n_14337), .B (n_7160), .Y (n_12412));
NOR2X1 g68086(.A (n_12410), .B (n_12409), .Y (n_12411));
OR2X1 g68091(.A (n_12399), .B (n_15968), .Y (n_12408));
NOR2X1 g68093(.A (n_10182), .B (n_7745), .Y (n_12406));
NAND2X1 g68096(.A (n_12404), .B (n_18264), .Y (n_12405));
AND2X1 g68098(.A (n_12402), .B (n_28642), .Y (n_12403));
AND2X1 g68099(.A (n_12399), .B (n_6409), .Y (n_12400));
NOR2X1 g68100(.A (n_6847), .B (n_7548), .Y (n_17222));
NAND2X1 g68101(.A (n_12397), .B (n_28692), .Y (n_16614));
NAND2X1 g68105(.A (n_18264), .B (n_8840), .Y (n_12396));
NAND2X1 g68108(.A (n_7241), .B (n_5329), .Y (n_12395));
INVX1 g68110(.A (n_12392), .Y (n_12393));
NAND2X1 g68113(.A (n_12389), .B (n_19364), .Y (n_12390));
OR2X1 g68118(.A (n_12762), .B (n_9388), .Y (n_15432));
NOR2X1 g68129(.A (n_13052), .B (n_4511), .Y (n_12387));
NAND2X1 g68131(.A (n_10295), .B (n_12385), .Y (n_12386));
NAND2X1 g68137(.A (n_12383), .B (n_6491), .Y (n_12384));
NAND2X1 g68143(.A (n_9889), .B (n_2570), .Y (n_12382));
AND2X1 g68146(.A (n_6041), .B (n_9527), .Y (n_16441));
INVX1 g68148(.A (n_12380), .Y (n_12381));
NAND2X1 g68151(.A (n_10091), .B (n_5322), .Y (n_12379));
AND2X1 g68154(.A (n_9315), .B (n_15166), .Y (n_12378));
NAND2X1 g68157(.A (n_12376), .B (n_12375), .Y (n_12377));
INVX1 g68163(.A (n_9821), .Y (n_14161));
NAND2X1 g68166(.A (n_12373), .B (n_12078), .Y (n_12374));
NAND2X1 g68168(.A (n_12852), .B (n_5820), .Y (n_12372));
NAND2X1 g68172(.A (n_12359), .B (n_12370), .Y (n_12371));
NAND2X1 g68177(.A (n_8088), .B (n_14055), .Y (n_12369));
NOR2X1 g68179(.A (n_9041), .B (n_12366), .Y (n_12368));
INVX1 g68184(.A (n_10844), .Y (n_12365));
NAND2X1 g68196(.A (n_27671), .B (n_16090), .Y (n_14150));
NAND2X1 g68198(.A (n_8527), .B (n_6611), .Y (n_12364));
NOR2X1 g68199(.A (n_10380), .B (n_12362), .Y (n_12363));
NAND2X1 g68201(.A (n_7719), .B (n_13720), .Y (n_12361));
INVX1 g68206(.A (n_9924), .Y (n_17129));
NAND2X1 g68210(.A (n_14821), .B (n_12359), .Y (n_12360));
NAND2X1 g68216(.A (n_10223), .B (n_20325), .Y (n_12358));
NAND2X1 g68217(.A (n_8874), .B (n_12628), .Y (n_12356));
NAND2X1 g68219(.A (n_15103), .B (n_12354), .Y (n_12355));
NOR2X1 g68221(.A (n_9990), .B (n_6774), .Y (n_12353));
NOR2X1 g68225(.A (n_7709), .B (n_29269), .Y (n_12352));
NAND2X1 g68228(.A (n_7709), .B (n_6670), .Y (n_12351));
NAND2X1 g68229(.A (n_7428), .B (n_12349), .Y (n_12350));
NAND2X1 g68238(.A (n_12347), .B (n_29199), .Y (n_12348));
NAND2X1 g68240(.A (n_2595), .B (n_8262), .Y (n_12346));
AND2X1 g68242(.A (n_15137), .B (n_14007), .Y (n_12345));
AOI21X1 g68243(.A0 (n_10237), .A1 (n_16198), .B0 (n_13341), .Y(n_12344));
NAND2X1 g68248(.A (n_12342), .B (n_17912), .Y (n_28245));
INVX1 g68249(.A (n_27899), .Y (n_12341));
NOR2X1 g68256(.A (n_8227), .B (n_12340), .Y (n_15644));
NAND2X1 g68258(.A (n_6941), .B (n_6117), .Y (n_12339));
NAND2X1 g68264(.A (n_12354), .B (n_12337), .Y (n_12338));
NAND2X1 g68270(.A (n_12335), .B (n_9029), .Y (n_12336));
INVX1 g68271(.A (n_15048), .Y (n_12334));
NOR2X1 g72917(.A (n_2912), .B (n_11823), .Y (n_20567));
NOR2X1 g68277(.A (n_8860), .B (n_18920), .Y (n_12333));
NOR2X1 g68285(.A (n_10589), .B (n_14589), .Y (n_12331));
NAND2X1 g68286(.A (n_7161), .B (n_8878), .Y (n_16927));
NAND2X1 g68287(.A (n_8447), .B (n_9988), .Y (n_12330));
INVX1 g68290(.A (n_12329), .Y (n_14122));
AND2X1 g68298(.A (n_11625), .B (n_12740), .Y (n_12328));
NOR2X1 g68302(.A (n_8568), .B (n_13083), .Y (n_12327));
NAND2X1 g68304(.A (n_9856), .B (n_6144), .Y (n_12326));
AND2X1 g68305(.A (n_12324), .B (n_12713), .Y (n_12325));
NAND2X1 g68314(.A (n_12322), .B (n_6870), .Y (n_12323));
NAND2X1 g68318(.A (n_27744), .B (n_6475), .Y (n_12321));
INVX1 g68324(.A (n_12319), .Y (n_12320));
NAND2X1 g68327(.A (n_12316), .B (n_19791), .Y (n_12317));
NAND2X1 g68334(.A (n_12802), .B (n_11582), .Y (n_12315));
NAND2X1 g68336(.A (n_12313), .B (n_8155), .Y (n_12314));
INVX1 g68341(.A (n_12312), .Y (n_15415));
NAND2X1 g68344(.A (n_9134), .B (n_12309), .Y (n_12310));
NAND2X1 g68346(.A (n_7035), .B (n_15600), .Y (n_12308));
NAND2X1 g68351(.A (n_12907), .B (n_12306), .Y (n_12307));
NOR2X1 g68356(.A (n_29173), .B (n_12303), .Y (n_12305));
INVX1 g68358(.A (n_12301), .Y (n_12302));
NOR2X1 g68361(.A (n_12299), .B (n_12298), .Y (n_12300));
NAND4X1 g68374(.A (n_12292), .B (n_12291), .C (n_6298), .D (n_4060),.Y (n_12293));
NAND2X1 g68382(.A (n_6980), .B (n_12289), .Y (n_12290));
NAND2X1 g68387(.A (n_18254), .B (n_16978), .Y (n_12288));
NAND2X1 g68390(.A (n_12285), .B (n_8566), .Y (n_12286));
INVX1 g68396(.A (n_13454), .Y (n_12282));
NAND2X1 g68399(.A (n_10071), .B (n_14592), .Y (n_12281));
OR2X1 g68401(.A (n_15085), .B (n_10389), .Y (n_12280));
INVX1 g68405(.A (n_17832), .Y (n_14084));
NAND2X1 g68409(.A (n_12278), .B (n_9982), .Y (n_12279));
NOR2X1 g68410(.A (n_7077), .B (n_10265), .Y (n_12277));
NAND2X1 g68415(.A (n_6714), .B (n_12275), .Y (n_12276));
NAND2X1 g68417(.A (n_7023), .B (n_5136), .Y (n_12274));
INVX1 g68421(.A (n_12272), .Y (n_12271));
NOR2X1 g68424(.A (n_8885), .B (n_5318), .Y (n_12270));
INVX1 g68430(.A (n_16676), .Y (n_16593));
NAND2X2 g72212(.A (n_12268), .B (n_11831), .Y (n_15068));
NAND2X1 g68434(.A (n_12266), .B (n_2701), .Y (n_12267));
INVX1 g68437(.A (n_10785), .Y (n_14076));
NAND3X1 g68446(.A (n_4993), .B (n_5874), .C (n_6660), .Y (n_12265));
NAND2X1 g68453(.A (n_8255), .B (n_18889), .Y (n_12264));
NAND2X1 g68456(.A (n_5330), .B (n_27475), .Y (n_12263));
AOI21X1 g68461(.A0 (n_10312), .A1 (n_1424), .B0 (n_6238), .Y(n_12261));
NOR2X1 g68465(.A (n_5929), .B (n_28834), .Y (n_12260));
NAND2X1 g68467(.A (n_8672), .B (n_7065), .Y (n_12258));
AND2X1 g68470(.A (n_8059), .B (n_12256), .Y (n_12257));
NOR2X1 g68474(.A (n_6063), .B (n_9286), .Y (n_12255));
INVX1 g68477(.A (n_10765), .Y (n_12254));
NAND2X1 g68480(.A (n_8695), .B (n_17003), .Y (n_12253));
NAND2X1 g68482(.A (n_3533), .B (n_12251), .Y (n_12252));
AOI21X1 g68489(.A0 (n_12249), .A1 (n_28575), .B0 (n_7278), .Y(n_12250));
NOR2X1 g68492(.A (n_9515), .B (n_10362), .Y (n_12248));
NOR2X1 g68493(.A (n_9123), .B (n_12246), .Y (n_12247));
INVX1 g68494(.A (n_10758), .Y (n_12245));
NAND2X1 g68499(.A (n_12243), .B (n_8224), .Y (n_12244));
AOI21X1 g68500(.A0 (n_5410), .A1 (n_28574), .B0 (n_13602), .Y(n_12242));
INVX1 g68502(.A (n_10752), .Y (n_12239));
NOR2X1 g68510(.A (n_6999), .B (n_10521), .Y (n_12238));
NAND2X1 g68513(.A (n_5763), .B (n_27403), .Y (n_12237));
NAND2X1 g68518(.A (n_8017), .B (n_12234), .Y (n_12235));
AOI21X1 g68522(.A0 (n_4459), .A1 (n_5503), .B0 (n_17912), .Y(n_12233));
NAND2X1 g68523(.A (n_8415), .B (n_18121), .Y (n_12231));
OR2X1 g68524(.A (n_27716), .B (n_12228), .Y (n_12230));
OAI21X1 g68527(.A0 (n_10551), .A1 (n_17500), .B0 (n_6812), .Y(n_12227));
NAND2X1 g68536(.A (n_8388), .B (n_18094), .Y (n_12226));
NAND2X1 g68537(.A (n_8895), .B (n_12224), .Y (n_12225));
AOI21X1 g68538(.A0 (n_12222), .A1 (n_2674), .B0 (n_7064), .Y(n_12223));
AOI21X1 g68543(.A0 (n_8499), .A1 (n_13593), .B0 (n_21122), .Y(n_12221));
NOR2X1 g68544(.A (n_6955), .B (n_10476), .Y (n_12220));
AND2X1 g68549(.A (n_7983), .B (n_11172), .Y (n_12219));
INVX1 g68556(.A (n_10742), .Y (n_28840));
INVX1 g68562(.A (n_10741), .Y (n_12217));
INVX1 g68564(.A (n_10740), .Y (n_12216));
NAND2X1 g68567(.A (n_5229), .B (n_12214), .Y (n_12215));
NAND2X1 g68572(.A (n_8565), .B (n_10268), .Y (n_12213));
NAND2X1 g68574(.A (n_8129), .B (n_18102), .Y (n_12212));
NAND2X1 g68575(.A (n_8402), .B (n_6732), .Y (n_12211));
NAND2X1 g68576(.A (n_5563), .B (n_12209), .Y (n_12210));
AOI21X1 g68581(.A0 (n_4374), .A1 (n_3791), .B0 (n_8940), .Y(n_12208));
NAND2X1 g68585(.A (n_8138), .B (n_12206), .Y (n_12207));
NOR2X1 g68586(.A (n_9107), .B (n_12664), .Y (n_12205));
NAND2X1 g68590(.A (n_3577), .B (n_12203), .Y (n_12204));
AOI21X1 g68594(.A0 (n_4309), .A1 (n_29269), .B0 (n_8356), .Y(n_12202));
NAND2X1 g68601(.A (n_9091), .B (n_12803), .Y (n_12200));
NAND2X1 g68603(.A (n_9081), .B (n_12198), .Y (n_12199));
AOI21X1 g68604(.A0 (n_4754), .A1 (n_6534), .B0 (n_7871), .Y(n_12197));
AOI21X1 g68605(.A0 (n_12123), .A1 (n_7410), .B0 (n_11233), .Y(n_12195));
AOI21X1 g68610(.A0 (n_6365), .A1 (n_29297), .B0 (n_9130), .Y(n_12194));
NAND2X1 g68612(.A (n_8905), .B (n_12192), .Y (n_12193));
NAND2X1 g68621(.A (n_8793), .B (n_12189), .Y (n_12190));
NAND2X1 g68622(.A (n_8956), .B (n_12187), .Y (n_12188));
NAND2X1 g68625(.A (n_7835), .B (n_8513), .Y (n_12186));
AOI21X1 g68630(.A0 (n_12121), .A1 (n_7325), .B0 (n_9459), .Y(n_12185));
NAND2X1 g68631(.A (n_8977), .B (n_8519), .Y (n_12183));
NAND2X1 g68632(.A (n_9015), .B (n_12347), .Y (n_12182));
AOI21X1 g68633(.A0 (n_6634), .A1 (n_2779), .B0 (n_5697), .Y(n_12181));
AOI21X1 g68635(.A0 (n_3514), .A1 (n_9783), .B0 (n_9096), .Y(n_12180));
NAND2X1 g68642(.A (n_8913), .B (n_12177), .Y (n_12178));
NOR2X1 g68643(.A (n_8900), .B (n_12175), .Y (n_12176));
AOI21X1 g68650(.A0 (n_7846), .A1 (n_16198), .B0 (n_7558), .Y(n_12174));
NAND2X1 g68654(.A (n_9103), .B (n_12172), .Y (n_12173));
NAND2X1 g68657(.A (n_7340), .B (n_12560), .Y (n_25828));
AOI21X1 g68658(.A0 (n_6697), .A1 (n_12169), .B0 (n_7249), .Y(n_12170));
NOR2X1 g68664(.A (n_8428), .B (n_28583), .Y (n_12168));
NOR2X1 g68667(.A (n_7327), .B (n_10122), .Y (n_12167));
AOI21X1 g68682(.A0 (n_5073), .A1 (n_8794), .B0 (n_4159), .Y(n_12166));
OAI21X1 g68684(.A0 (n_3818), .A1 (n_3391), .B0 (n_13418), .Y(n_12165));
AOI21X1 g68686(.A0 (n_12162), .A1 (n_4144), .B0 (n_12161), .Y(n_12163));
NAND2X1 g68687(.A (n_7905), .B (n_7847), .Y (n_12160));
OR2X1 g68689(.A (n_8019), .B (n_6375), .Y (n_12159));
AND2X1 g68690(.A (n_8572), .B (n_5887), .Y (n_12158));
AOI21X1 g68697(.A0 (n_12155), .A1 (n_6439), .B0 (n_12154), .Y(n_12156));
OAI21X1 g68701(.A0 (n_5167), .A1 (n_12144), .B0 (n_5104), .Y(n_12153));
NAND2X1 g68704(.A (n_8443), .B (n_1883), .Y (n_12152));
NAND2X1 g68707(.A (n_8095), .B (n_13217), .Y (n_12150));
AOI21X1 g68708(.A0 (n_28870), .A1 (n_10573), .B0 (n_4832), .Y(n_12149));
NAND2X1 g68713(.A (n_4147), .B (n_12762), .Y (n_12148));
AOI21X1 g68717(.A0 (n_6386), .A1 (n_4181), .B0 (n_2466), .Y(n_12146));
OAI21X1 g68720(.A0 (n_5316), .A1 (n_12144), .B0 (n_11694), .Y(n_12145));
NAND2X1 g68728(.A (n_8222), .B (n_1744), .Y (n_12143));
OR2X1 g68739(.A (n_8504), .B (n_12140), .Y (n_12141));
NAND2X1 g68740(.A (n_8542), .B (n_12138), .Y (n_12139));
NAND2X1 g68743(.A (n_8460), .B (n_12136), .Y (n_12137));
AOI21X1 g68744(.A0 (n_12134), .A1 (n_12133), .B0 (n_8614), .Y(n_12135));
NAND2X1 g68748(.A (n_7694), .B (n_8320), .Y (n_12132));
OR2X1 g68751(.A (n_6882), .B (n_12129), .Y (n_12130));
OR2X1 g68752(.A (n_8234), .B (n_12127), .Y (n_12128));
OAI21X1 g68758(.A0 (n_5215), .A1 (n_10716), .B0 (n_5778), .Y(n_12126));
NAND2X1 g68759(.A (n_8006), .B (n_15627), .Y (n_12125));
OAI21X1 g68765(.A0 (n_12123), .A1 (n_6232), .B0 (n_2357), .Y(n_12124));
OAI21X1 g68767(.A0 (n_12121), .A1 (n_6188), .B0 (n_7803), .Y(n_12122));
AND2X1 g68789(.A (n_4354), .B (n_8585), .Y (n_12120));
AND2X1 g68792(.A (n_4177), .B (n_8221), .Y (n_12119));
AND2X1 g68793(.A (n_5346), .B (n_8333), .Y (n_12118));
XOR2X1 g68826(.A (n_972), .B (n_7775), .Y (n_12117));
XOR2X1 g68828(.A (n_1012), .B (n_6398), .Y (n_12116));
XOR2X1 g68838(.A (n_1041), .B (n_6402), .Y (n_12115));
XOR2X1 g68840(.A (n_1140), .B (n_6405), .Y (n_12114));
INVX1 g69728(.A (n_12112), .Y (n_12113));
INVX1 g69024(.A (n_9592), .Y (n_13947));
NAND2X1 g69042(.A (n_9675), .B (n_27757), .Y (n_12108));
NAND2X1 g69053(.A (n_12106), .B (n_12105), .Y (n_17590));
INVX2 g72127(.A (n_10616), .Y (n_13801));
NAND2X1 g69108(.A (n_11772), .B (n_6534), .Y (n_12102));
INVX1 g69110(.A (n_15326), .Y (n_12100));
INVX1 g69113(.A (n_28164), .Y (n_12099));
INVX1 g69125(.A (n_12098), .Y (n_13946));
INVX1 g69130(.A (n_14442), .Y (n_16005));
INVX1 g69132(.A (n_12096), .Y (n_17689));
OR2X1 g69138(.A (n_29062), .B (n_6753), .Y (n_12095));
NAND2X1 g69143(.A (n_7967), .B (n_6534), .Y (n_12093));
INVX1 g69163(.A (n_14384), .Y (n_12091));
INVX1 g69176(.A (n_10600), .Y (n_15259));
INVX1 g69200(.A (n_12085), .Y (n_17717));
INVX1 g69205(.A (n_12518), .Y (n_16366));
INVX1 g69222(.A (n_12081), .Y (n_12082));
OR2X1 g69245(.A (n_12078), .B (n_6534), .Y (n_12079));
INVX1 g69253(.A (n_14535), .Y (n_12077));
INVX1 g69317(.A (n_12591), .Y (n_12073));
INVX1 g69352(.A (n_12072), .Y (n_16472));
INVX1 g69357(.A (n_12070), .Y (n_12071));
INVX2 g69378(.A (n_14009), .Y (n_13942));
INVX1 g69413(.A (n_12067), .Y (n_13940));
INVX1 g69469(.A (n_12060), .Y (n_12061));
NAND2X1 g69527(.A (n_25597), .B (n_11052), .Y (n_12059));
NAND2X1 g69542(.A (n_11801), .B (n_7201), .Y (n_12057));
INVX1 g69579(.A (n_10512), .Y (n_13936));
AND2X1 g69584(.A (n_8103), .B (n_12858), .Y (n_12056));
NAND2X1 g69592(.A (n_7910), .B (n_6185), .Y (n_12055));
NAND2X1 g69613(.A (n_8007), .B (n_9084), .Y (n_12054));
NAND2X2 g69629(.A (n_9311), .B (n_18266), .Y (n_16812));
INVX2 g69659(.A (n_14188), .Y (n_15969));
NAND2X1 g69691(.A (n_9665), .B (n_9783), .Y (n_12049));
INVX1 g69764(.A (n_10456), .Y (n_13932));
INVX1 g69803(.A (n_12042), .Y (n_12043));
INVX1 g69854(.A (n_14314), .Y (n_13928));
INVX1 g69865(.A (n_14141), .Y (n_16100));
INVX1 g69879(.A (n_26042), .Y (n_12032));
INVX1 g69903(.A (n_14139), .Y (n_13927));
INVX1 g69909(.A (n_14284), .Y (n_13926));
INVX1 g69912(.A (n_12028), .Y (n_12029));
INVX1 g69916(.A (n_12026), .Y (n_12027));
NAND2X1 g68323(.A (n_6038), .B (n_8878), .Y (n_18114));
INVX1 g69951(.A (n_12024), .Y (n_15990));
INVX1 g69967(.A (n_14078), .Y (n_13921));
INVX1 g69970(.A (n_12021), .Y (n_12023));
NAND2X1 g69980(.A (n_12020), .B (n_12019), .Y (n_17232));
NAND2X1 g70003(.A (n_7946), .B (n_4898), .Y (n_12015));
INVX1 g72055(.A (n_12013), .Y (n_12014));
INVX1 g70018(.A (n_12012), .Y (n_16375));
INVX1 g70043(.A (n_15087), .Y (n_12006));
NAND2X1 g70107(.A (n_7943), .B (n_28404), .Y (n_12001));
INVX1 g70110(.A (n_10370), .Y (n_17935));
NAND2X1 g70121(.A (n_11687), .B (n_11998), .Y (n_11999));
INVX1 g70139(.A (n_8892), .Y (n_13912));
INVX1 g70174(.A (n_26916), .Y (n_11993));
AOI21X1 g65392(.A0 (n_4592), .A1 (n_11157), .B0 (n_15894), .Y(n_11990));
INVX1 g70239(.A (n_14190), .Y (n_13907));
INVX1 g70254(.A (n_27135), .Y (n_11988));
INVX1 g70313(.A (n_10316), .Y (n_16123));
OR2X1 g70332(.A (n_11984), .B (n_20325), .Y (n_11985));
INVX1 g70344(.A (n_15011), .Y (n_11981));
NAND2X1 g70352(.A (n_7965), .B (n_29297), .Y (n_11980));
OR2X1 g70363(.A (n_5892), .B (n_11976), .Y (n_11978));
NAND2X1 g70368(.A (n_11976), .B (n_9783), .Y (n_11977));
INVX1 g70407(.A (n_10292), .Y (n_17236));
INVX1 g70429(.A (n_11967), .Y (n_17687));
NAND2X1 g70451(.A (n_7705), .B (n_11322), .Y (n_11965));
NAND2X1 g70462(.A (n_7928), .B (n_15708), .Y (n_11963));
INVX1 g70487(.A (n_14082), .Y (n_17328));
NAND2X1 g70497(.A (n_8010), .B (n_18785), .Y (n_11957));
INVX2 g70528(.A (n_11953), .Y (n_15918));
INVX1 g70536(.A (n_14099), .Y (n_11951));
INVX1 g70554(.A (n_13432), .Y (n_11948));
INVX1 g70562(.A (n_10258), .Y (n_13882));
INVX1 g70585(.A (n_11945), .Y (n_11946));
NAND2X1 g70666(.A (n_5410), .B (n_25597), .Y (n_13880));
INVX1 g70669(.A (n_26492), .Y (n_11934));
INVX1 g70684(.A (n_11929), .Y (n_11931));
NAND2X1 g70695(.A (n_5211), .B (n_5329), .Y (n_11927));
OR2X1 g70704(.A (n_11924), .B (n_29139), .Y (n_13879));
INVX1 g70708(.A (n_11923), .Y (n_16184));
INVX1 g70728(.A (n_11920), .Y (n_11921));
INVX1 g70757(.A (n_11917), .Y (n_16830));
NAND2X1 g70761(.A (n_11916), .B (n_11812), .Y (n_16187));
OR2X1 g70791(.A (n_2839), .B (n_8709), .Y (n_15952));
INVX2 g70800(.A (n_10208), .Y (n_17723));
INVX1 g70853(.A (n_10197), .Y (n_18005));
NAND2X2 g70862(.A (n_28246), .B (n_8342), .Y (n_28804));
INVX1 g70870(.A (n_11900), .Y (n_16271));
INVX1 g70885(.A (n_11008), .Y (n_11897));
NOR2X1 g70889(.A (n_4166), .B (n_6711), .Y (n_11895));
INVX1 g70917(.A (n_11893), .Y (n_16169));
OR2X1 g70973(.A (n_7906), .B (n_9264), .Y (n_11888));
INVX1 g70974(.A (n_11886), .Y (n_11887));
INVX1 g70981(.A (n_10060), .Y (n_16883));
INVX1 g70988(.A (n_11884), .Y (n_11885));
INVX1 g70991(.A (n_11882), .Y (n_11883));
NAND2X2 g70995(.A (n_25597), .B (n_8363), .Y (n_16139));
NOR2X1 g72710(.A (n_7979), .B (n_15039), .Y (n_11880));
INVX1 g71011(.A (n_14380), .Y (n_11878));
INVX1 g71038(.A (n_11876), .Y (n_11877));
INVX1 g71049(.A (n_10138), .Y (n_11875));
NAND2X1 g71058(.A (n_2757), .B (n_28614), .Y (n_19608));
OR2X1 g71069(.A (n_12850), .B (n_9513), .Y (n_11871));
OR2X1 g71116(.A (n_7112), .B (n_6601), .Y (n_25736));
OR2X1 g71145(.A (n_3228), .B (n_7027), .Y (n_11865));
NOR2X1 g71176(.A (n_8452), .B (n_11864), .Y (n_13848));
AND2X1 g71187(.A (n_12078), .B (n_11861), .Y (n_11862));
NAND2X1 g71195(.A (n_8198), .B (n_27199), .Y (n_11860));
INVX1 g71243(.A (n_7632), .Y (n_15942));
OR2X1 g71250(.A (n_6889), .B (n_11984), .Y (n_11858));
INVX1 g71252(.A (n_10095), .Y (n_11857));
NAND2X1 g71256(.A (n_6397), .B (n_12559), .Y (n_11856));
NAND2X1 g71281(.A (n_8052), .B (n_11816), .Y (n_11853));
NAND2X1 g71287(.A (n_6744), .B (n_11850), .Y (n_11851));
INVX1 g71288(.A (n_11848), .Y (n_11849));
NAND2X1 g71292(.A (n_9965), .B (n_11976), .Y (n_13843));
NAND2X1 g71369(.A (n_6397), .B (n_2043), .Y (n_15555));
INVX1 g71412(.A (n_11843), .Y (n_14761));
OR2X1 g71430(.A (n_12436), .B (n_11323), .Y (n_17776));
INVX1 g71468(.A (n_13383), .Y (n_17253));
NAND2X1 g71497(.A (n_7820), .B (n_13872), .Y (n_11839));
OR2X1 g71507(.A (n_8966), .B (n_13846), .Y (n_11837));
OR2X1 g71511(.A (n_8029), .B (n_11835), .Y (n_11836));
NAND2X1 g71512(.A (n_8141), .B (n_6548), .Y (n_16040));
INVX1 g71518(.A (n_11833), .Y (n_11834));
NAND2X1 g71529(.A (n_2112), .B (n_11831), .Y (n_15860));
NOR2X1 g71556(.A (n_12494), .B (n_29329), .Y (n_13835));
NAND2X1 g71936(.A (n_7898), .B (n_13768), .Y (n_25676));
INVX1 g71565(.A (n_14700), .Y (n_16142));
NAND2X1 g71568(.A (n_2757), .B (n_6748), .Y (n_16512));
NAND3X1 g71586(.A (n_7832), .B (n_6587), .C (n_3301), .Y (n_11827));
NAND2X1 g71608(.A (n_5319), .B (n_9942), .Y (n_29143));
NAND2X1 g71636(.A (n_7961), .B (n_11823), .Y (n_16130));
INVX1 g71673(.A (n_11821), .Y (n_16174));
INVX1 g71682(.A (n_14017), .Y (n_11820));
INVX1 g71707(.A (n_11819), .Y (n_13830));
NOR2X1 g71711(.A (n_9420), .B (n_13490), .Y (n_11818));
NAND2X1 g71712(.A (n_12020), .B (n_11816), .Y (n_11817));
INVX1 g71719(.A (n_13550), .Y (n_11815));
NAND2X1 g71731(.A (n_10147), .B (n_11812), .Y (n_15858));
NAND2X1 g71732(.A (n_7812), .B (n_11810), .Y (n_11811));
INVX1 g71786(.A (n_11808), .Y (n_16051));
NAND2X1 g71794(.A (n_7006), .B (n_6476), .Y (n_16082));
INVX1 g72642(.A (n_14093), .Y (n_16163));
NAND2X1 g71849(.A (n_7936), .B (n_5389), .Y (n_11802));
NAND2X1 g71853(.A (n_28611), .B (n_11261), .Y (n_19417));
INVX1 g71866(.A (n_9963), .Y (n_18275));
NAND2X1 g71873(.A (n_3160), .B (n_11801), .Y (n_13825));
INVX1 g71879(.A (n_11799), .Y (n_11800));
INVX1 g71881(.A (n_14048), .Y (n_11798));
INVX1 g71904(.A (n_11795), .Y (n_16236));
INVX1 g71925(.A (n_9951), .Y (n_15958));
OR2X1 g71948(.A (n_11864), .B (n_27688), .Y (n_11791));
INVX1 g71956(.A (n_14392), .Y (n_16225));
INVX1 g71972(.A (n_9943), .Y (n_17033));
INVX1 g71981(.A (n_10149), .Y (n_17041));
NOR2X1 g72007(.A (n_7881), .B (n_29228), .Y (n_11787));
OR2X1 g72011(.A (n_7789), .B (n_6390), .Y (n_25639));
OR2X1 g72018(.A (n_9669), .B (n_9003), .Y (n_13818));
NAND2X1 g72051(.A (n_11752), .B (n_15388), .Y (n_11784));
INVX1 g72060(.A (n_14183), .Y (n_11782));
NOR2X1 g72095(.A (n_4188), .B (n_11728), .Y (n_20582));
INVX1 g72103(.A (n_9920), .Y (n_11777));
INVX1 g72108(.A (n_9918), .Y (n_13807));
OR2X1 g72129(.A (n_6746), .B (n_12850), .Y (n_11776));
NAND2X1 g72164(.A (n_14113), .B (n_11772), .Y (n_11773));
INVX1 g72200(.A (n_14028), .Y (n_11768));
NAND2X1 g72213(.A (n_7902), .B (n_8470), .Y (n_16245));
INVX1 g72215(.A (n_11764), .Y (n_13795));
NAND2X1 g72258(.A (n_8023), .B (n_4223), .Y (n_11760));
NAND2X1 g72300(.A (n_12106), .B (n_2895), .Y (n_11758));
NAND2X1 g72402(.A (n_5104), .B (n_28614), .Y (n_20955));
NOR2X1 g72419(.A (n_11752), .B (n_7116), .Y (n_11753));
NAND2X1 g72421(.A (n_7945), .B (n_8945), .Y (n_16080));
NAND2X1 g72481(.A (n_11749), .B (n_1497), .Y (n_11750));
AND2X1 g72505(.A (n_7840), .B (n_11745), .Y (n_11746));
AND2X1 g72516(.A (n_11864), .B (n_11743), .Y (n_11744));
INVX1 g72549(.A (n_9837), .Y (n_11742));
OR2X1 g72552(.A (n_7892), .B (n_13846), .Y (n_11741));
NAND2X1 g72577(.A (n_6764), .B (n_11739), .Y (n_11740));
NAND2X1 g72578(.A (n_7940), .B (n_15894), .Y (n_11738));
NOR2X1 g72585(.A (n_9368), .B (n_5140), .Y (n_13770));
NAND2X1 g72655(.A (n_6346), .B (n_11734), .Y (n_11735));
INVX1 g72656(.A (n_11732), .Y (n_11733));
NOR2X1 g72659(.A (n_9640), .B (n_11731), .Y (n_13766));
INVX1 g72661(.A (n_11729), .Y (n_11730));
NAND2X1 g72666(.A (n_11648), .B (n_9639), .Y (n_13765));
OR2X1 g72683(.A (n_8080), .B (n_3386), .Y (n_11727));
NAND2X1 g72739(.A (n_14667), .B (n_8015), .Y (n_20948));
INVX1 g72741(.A (n_14216), .Y (n_11718));
OR2X1 g72764(.A (n_2409), .B (n_7887), .Y (n_11716));
INVX1 g72766(.A (n_11714), .Y (n_11715));
NAND2X1 g72808(.A (n_7885), .B (n_19755), .Y (n_11713));
INVX1 g72828(.A (n_11712), .Y (n_16089));
INVX1 g72844(.A (n_11710), .Y (n_15874));
NAND2X1 g72850(.A (n_7784), .B (n_9444), .Y (n_11709));
INVX1 g72963(.A (n_11701), .Y (n_16266));
INVX1 g72965(.A (n_11700), .Y (n_15238));
NAND2X1 g72977(.A (n_7957), .B (n_9221), .Y (n_11699));
NAND2X1 g72978(.A (n_2281), .B (n_11901), .Y (n_16665));
INVX1 g72981(.A (n_11698), .Y (n_14472));
NOR2X1 g73040(.A (n_1768), .B (n_9661), .Y (n_13740));
AOI21X1 g63210(.A0 (n_7640), .A1 (n_11354), .B0 (n_7227), .Y(n_11690));
NAND2X1 g73102(.A (n_27309), .B (n_11687), .Y (n_11689));
OR2X1 g73120(.A (n_7904), .B (n_10389), .Y (n_11686));
AND2X1 g73132(.A (n_6563), .B (n_11743), .Y (n_11685));
NAND2X1 g73163(.A (n_11682), .B (n_7769), .Y (n_11683));
OR2X1 g73173(.A (n_7889), .B (n_13846), .Y (n_11681));
INVX1 g73191(.A (n_14500), .Y (n_11678));
OAI21X1 g73218(.A0 (n_4018), .A1 (n_9264), .B0 (n_7954), .Y(n_11677));
NAND2X1 g73222(.A (n_5228), .B (n_6952), .Y (n_11676));
NAND2X1 g73224(.A (n_5894), .B (n_6563), .Y (n_11674));
OR2X1 g73225(.A (n_5276), .B (n_11671), .Y (n_11672));
AOI21X1 g73229(.A0 (n_11669), .A1 (n_9682), .B0 (n_7830), .Y(n_11670));
OR2X1 g73243(.A (n_7978), .B (n_11667), .Y (n_11668));
NAND2X1 g73245(.A (n_6275), .B (n_7840), .Y (n_11666));
NAND2X1 g73248(.A (n_5875), .B (n_6809), .Y (n_11664));
OAI21X1 g63275(.A0 (n_7811), .A1 (n_11662), .B0 (n_9486), .Y(n_11663));
OR2X1 g73269(.A (n_4726), .B (n_11660), .Y (n_11661));
NAND3X1 g63350(.A (n_11655), .B (n_27410), .C (n_13421), .Y(n_11656));
INVX1 g74104(.A (n_11649), .Y (n_11650));
DFFX1 u0_r0_out_reg[30] (.CK (clk), .D (n_7854), .Q (u0_rcon_1059),.QN ());
DFFX1 u0_r0_out_reg[31] (.CK (clk), .D (n_7859), .Q (u0_rcon_1060),.QN ());
NAND2X1 g72557(.A (n_11648), .B (n_11812), .Y (n_17915));
NAND3X1 g75083(.A (n_13679), .B (n_3868), .C (n_11312), .Y (n_11647));
AOI21X1 g63745(.A0 (n_11642), .A1 (n_13324), .B0 (n_17912), .Y(n_11643));
INVX1 g72540(.A (n_20178), .Y (n_11641));
XOR2X1 g76345(.A (n_2434), .B (n_16480), .Y (n_11636));
INVX2 g75774(.A (n_11632), .Y (n_15799));
INVX1 g72525(.A (n_15310), .Y (n_16199));
OAI21X1 g64056(.A0 (n_6904), .A1 (n_5004), .B0 (n_17912), .Y(n_11628));
NAND4X1 g63955(.A (n_10934), .B (n_11383), .C (n_11626), .D(n_11625), .Y (n_11627));
MX2X1 g60675(.A (n_11608), .B (n_13728), .S0 (u0_r0_rcnt[0] ), .Y(n_11624));
XOR2X1 g76111(.A (n_2769), .B (n_13466), .Y (n_11623));
MX2X1 g64006(.A (n_7618), .B (n_11620), .S0 (n_14142), .Y (n_11621));
XOR2X1 g76129(.A (text_in_r[28] ), .B (n_2838), .Y (n_11618));
MX2X1 g64008(.A (n_7804), .B (n_29336), .S0 (n_4582), .Y (n_11617));
NAND4X1 g64012(.A (n_5374), .B (n_11615), .C (n_13703), .D (n_6127),.Y (n_11616));
OAI21X1 g64038(.A0 (n_6924), .A1 (n_28156), .B0 (n_27133), .Y(n_11614));
NAND3X1 g64041(.A (n_9442), .B (n_6933), .C (n_11739), .Y (n_11613));
OAI21X1 g64050(.A0 (n_7233), .A1 (n_28812), .B0 (n_13326), .Y(n_11612));
OAI21X1 g64052(.A0 (n_7140), .A1 (n_28045), .B0 (n_14624), .Y(n_11611));
OAI21X1 g64053(.A0 (n_7187), .A1 (n_26489), .B0 (n_9410), .Y(n_28887));
MX2X1 g60717(.A (n_13728), .B (n_11608), .S0 (u0_r0_rcnt[0] ), .Y(n_11609));
XOR2X1 g76236(.A (text_in_r[4] ), .B (n_3955), .Y (n_11606));
NAND2X1 g64070(.A (n_9296), .B (n_11603), .Y (n_11604));
AND2X1 g64072(.A (n_9229), .B (n_9527), .Y (n_11602));
OAI21X1 g64075(.A0 (n_7171), .A1 (n_6574), .B0 (n_11400), .Y(n_11601));
OAI21X1 g64082(.A0 (n_7004), .A1 (n_10546), .B0 (n_29048), .Y(n_11600));
OAI21X1 g64084(.A0 (n_7217), .A1 (n_7617), .B0 (n_16480), .Y(n_11599));
AOI21X1 g64097(.A0 (n_6872), .A1 (n_9293), .B0 (n_15674), .Y(n_11598));
NAND2X1 g64100(.A (n_9532), .B (n_15039), .Y (n_11597));
AOI21X1 g64102(.A0 (n_6627), .A1 (n_13195), .B0 (n_875), .Y(n_11596));
AOI21X1 g64104(.A0 (n_6705), .A1 (n_11593), .B0 (n_3538), .Y(n_11594));
XOR2X1 g76334(.A (text_in_r[20] ), .B (n_530), .Y (n_11592));
NOR2X1 g64117(.A (n_13316), .B (n_18205), .Y (n_11590));
OR4X1 g64128(.A (n_15568), .B (n_7201), .C (n_4721), .D (n_5333), .Y(n_11589));
OR4X1 g64129(.A (n_17864), .B (n_13247), .C (n_9500), .D (n_4163), .Y(n_11587));
NAND3X1 g64132(.A (n_12313), .B (n_5477), .C (n_11585), .Y (n_11586));
NAND2X1 g64137(.A (n_9278), .B (n_12827), .Y (n_21660));
INVX1 g64147(.A (n_9599), .Y (n_11584));
AOI21X1 g65384(.A0 (n_5626), .A1 (n_11582), .B0 (n_27099), .Y(n_11583));
OR4X1 g64194(.A (n_15039), .B (n_6185), .C (n_7947), .D (n_5750), .Y(n_11581));
NOR2X1 g64205(.A (n_11579), .B (n_16480), .Y (n_11580));
OR4X1 g64210(.A (n_17377), .B (n_9264), .C (n_28744), .D (n_5259), .Y(n_11578));
OR4X1 g64213(.A (n_11576), .B (n_28433), .C (n_27124), .D (n_5428),.Y (n_11577));
NAND2X1 g64225(.A (n_10885), .B (n_17912), .Y (n_11575));
AOI21X1 g64246(.A0 (n_5547), .A1 (n_17531), .B0 (n_17571), .Y(n_11574));
AOI21X1 g64247(.A0 (n_6181), .A1 (n_14523), .B0 (n_15776), .Y(n_11573));
AOI21X1 g64255(.A0 (n_4340), .A1 (n_15825), .B0 (n_18168), .Y(n_11572));
NAND2X1 g64269(.A (n_11181), .B (n_9410), .Y (n_13569));
OR2X1 g64272(.A (n_13706), .B (n_12896), .Y (n_11570));
AOI21X1 g65371(.A0 (n_11533), .A1 (n_9800), .B0 (n_16754), .Y(n_11569));
NAND2X1 g64293(.A (n_11390), .B (n_11567), .Y (n_11568));
NAND3X1 g64295(.A (n_12644), .B (n_11565), .C (n_9509), .Y (n_11566));
NAND2X1 g64320(.A (n_11563), .B (n_11562), .Y (n_11564));
NAND2X1 g64356(.A (n_8745), .B (n_11560), .Y (n_11561));
AND2X1 g64380(.A (n_11558), .B (n_12801), .Y (n_11559));
NAND2X1 g64389(.A (n_11057), .B (n_14142), .Y (n_13531));
NOR2X1 g64401(.A (n_18347), .B (n_11317), .Y (n_11557));
NAND2X1 g64402(.A (n_13695), .B (n_12500), .Y (n_11556));
NAND2X1 g64414(.A (n_11554), .B (n_13316), .Y (n_11555));
AOI21X1 g64418(.A0 (n_6908), .A1 (n_8682), .B0 (n_1424), .Y(n_11553));
AND2X1 g64422(.A (n_11550), .B (n_11549), .Y (n_11551));
NAND2X1 g64425(.A (n_9489), .B (n_12827), .Y (n_15701));
AND2X1 g64438(.A (n_9196), .B (n_16480), .Y (n_11547));
AOI21X1 g64440(.A0 (n_7534), .A1 (n_11131), .B0 (n_16480), .Y(n_11546));
AOI21X1 g64445(.A0 (n_7211), .A1 (n_8503), .B0 (n_15712), .Y(n_11545));
AOI21X1 g64467(.A0 (n_11543), .A1 (n_3366), .B0 (n_20010), .Y(n_11544));
NAND2X1 g64470(.A (n_11091), .B (n_15568), .Y (n_13506));
OAI21X1 g64475(.A0 (n_5144), .A1 (n_16931), .B0 (n_933), .Y(n_11542));
NAND2X1 g64483(.A (n_11539), .B (n_10336), .Y (n_11540));
AOI21X1 g64499(.A0 (n_6425), .A1 (n_6512), .B0 (n_17260), .Y(n_11538));
NAND2X1 g64517(.A (n_8510), .B (n_13148), .Y (n_11535));
NAND3X1 g64527(.A (n_12486), .B (n_11533), .C (n_9472), .Y (n_11534));
AOI21X1 g64532(.A0 (n_7166), .A1 (n_7230), .B0 (n_14589), .Y(n_11532));
OR2X1 g64534(.A (n_9166), .B (n_11530), .Y (n_11531));
NAND2X1 g64537(.A (n_6927), .B (n_11528), .Y (n_11529));
NAND2X1 g64541(.A (n_28217), .B (n_13452), .Y (n_11527));
NAND2X1 g64549(.A (n_11524), .B (n_10483), .Y (n_11525));
NAND2X1 g64554(.A (n_13508), .B (n_11522), .Y (n_11523));
NAND2X1 g64589(.A (n_11520), .B (n_10880), .Y (n_11521));
OAI21X1 g64590(.A0 (n_6413), .A1 (n_19207), .B0 (n_1196), .Y(n_11519));
NAND3X1 g64601(.A (n_11517), .B (n_7051), .C (n_11516), .Y (n_11518));
AOI21X1 g64602(.A0 (n_7456), .A1 (n_8769), .B0 (n_15712), .Y(n_11515));
NAND2X1 g64604(.A (n_11255), .B (n_10061), .Y (n_11514));
AND2X1 g64607(.A (n_11512), .B (n_11086), .Y (n_11513));
AOI21X1 g64619(.A0 (n_7461), .A1 (n_11510), .B0 (n_16787), .Y(n_11511));
NAND2X1 g64643(.A (n_11512), .B (n_17266), .Y (n_11509));
DFFX1 dcnt_reg[1] (.CK (clk), .D (n_9250), .Q (dcnt[1] ), .QN ());
NAND2X1 g64645(.A (n_9501), .B (n_13083), .Y (n_18421));
NAND2X1 g64655(.A (n_11507), .B (n_11506), .Y (n_11508));
NAND2X1 g64670(.A (n_15034), .B (n_9345), .Y (n_11505));
NAND2X1 g64677(.A (n_9160), .B (n_5559), .Y (n_11504));
NAND2X1 g64679(.A (n_12607), .B (n_13329), .Y (n_11503));
NAND3X1 g64699(.A (n_11501), .B (n_11500), .C (n_4727), .Y (n_11502));
NAND2X1 g64705(.A (n_14909), .B (n_27372), .Y (n_11499));
OAI21X1 g64718(.A0 (n_6434), .A1 (n_19191), .B0 (n_21174), .Y(n_11498));
NAND3X1 g64720(.A (n_11495), .B (n_7433), .C (n_10868), .Y (n_11496));
NAND2X1 g64723(.A (n_8426), .B (n_13159), .Y (n_11494));
AOI21X1 g64730(.A0 (n_6804), .A1 (n_11492), .B0 (n_9106), .Y(n_11493));
NAND2X1 g64735(.A (n_13725), .B (n_14330), .Y (n_11491));
AOI21X1 g64740(.A0 (n_7276), .A1 (n_8343), .B0 (n_11489), .Y(n_11490));
NOR2X1 g64748(.A (n_9174), .B (n_4898), .Y (n_11488));
INVX1 g64750(.A (n_11486), .Y (n_11487));
OR2X1 g64753(.A (n_11484), .B (n_26276), .Y (n_11485));
AOI21X1 g64755(.A0 (n_7038), .A1 (n_6333), .B0 (n_11576), .Y(n_11483));
NAND2X1 g72478(.A (n_14107), .B (n_27076), .Y (n_15863));
AOI21X1 g64775(.A0 (n_7033), .A1 (n_8635), .B0 (n_17411), .Y(n_11480));
OR2X1 g64779(.A (n_14765), .B (n_15776), .Y (n_11478));
OAI21X1 g64079(.A0 (n_7138), .A1 (n_6750), .B0 (n_13326), .Y(n_11476));
AOI21X1 g65387(.A0 (n_6034), .A1 (n_11473), .B0 (n_11052), .Y(n_11474));
NAND2X1 g64784(.A (n_11470), .B (n_11247), .Y (n_11471));
NAND2X1 g64791(.A (n_15556), .B (n_14927), .Y (n_11469));
AOI21X1 g64802(.A0 (n_7529), .A1 (n_12734), .B0 (n_17260), .Y(n_11468));
AOI21X1 g64811(.A0 (n_6801), .A1 (n_9567), .B0 (n_29074), .Y(n_11466));
AOI21X1 g64813(.A0 (n_6905), .A1 (n_8541), .B0 (n_27688), .Y(n_11465));
OAI21X1 g64851(.A0 (n_5170), .A1 (n_17477), .B0 (n_1397), .Y(n_11464));
NAND3X1 g65350(.A (n_11462), .B (n_3797), .C (n_11461), .Y (n_11463));
OAI21X1 g64888(.A0 (n_4151), .A1 (n_5813), .B0 (n_27910), .Y(n_11460));
NAND2X1 g64950(.A (n_11456), .B (n_7786), .Y (n_11457));
INVX1 g71566(.A (n_12373), .Y (n_14700));
AOI21X1 g65060(.A0 (n_5961), .A1 (n_5853), .B0 (n_9819), .Y(n_11454));
NAND2X1 g65063(.A (n_11452), .B (n_8724), .Y (n_11453));
INVX1 g65071(.A (n_9548), .Y (n_11451));
AOI21X1 g65082(.A0 (n_6045), .A1 (n_11449), .B0 (n_15986), .Y(n_11450));
NAND2X1 g73192(.A (n_5077), .B (n_4709), .Y (n_14500));
NAND2X1 g65181(.A (n_11345), .B (n_11447), .Y (n_11448));
DFFX1 u0_r0_out_reg[24] (.CK (clk), .D (n_7713), .Q (u0_rcon_1053),.QN ());
NAND2X1 g73186(.A (n_1784), .B (n_25440), .Y (n_25825));
NOR2X1 g65304(.A (n_13482), .B (n_18369), .Y (n_11445));
NOR2X1 g65448(.A (n_3959), .B (n_11439), .Y (n_11440));
NAND2X1 g70240(.A (n_8024), .B (n_8974), .Y (n_14190));
INVX1 g65507(.A (n_9530), .Y (n_11438));
NAND2X1 g65531(.A (n_7626), .B (n_4582), .Y (n_11437));
OR2X1 g72420(.A (n_11435), .B (n_6724), .Y (n_11436));
AOI21X1 g65538(.A0 (n_5664), .A1 (n_7717), .B0 (n_8708), .Y(n_11434));
AOI21X1 g65540(.A0 (n_10856), .A1 (n_7732), .B0 (n_15712), .Y(n_11433));
AOI21X1 g65595(.A0 (n_6237), .A1 (n_11431), .B0 (n_1424), .Y(n_11432));
AOI21X1 g65653(.A0 (n_10931), .A1 (n_28996), .B0 (n_11489), .Y(n_11428));
NAND3X1 g65727(.A (n_7557), .B (n_6942), .C (n_11431), .Y (n_11426));
NOR2X1 g65792(.A (n_4758), .B (n_11424), .Y (n_11425));
AOI21X1 g65807(.A0 (n_11422), .A1 (n_9844), .B0 (n_17912), .Y(n_11423));
NAND3X1 g65842(.A (n_7463), .B (n_7417), .C (n_9234), .Y (n_11421));
NAND3X1 g65845(.A (n_5996), .B (n_7452), .C (n_12189), .Y (n_11420));
AOI21X1 g65867(.A0 (n_11418), .A1 (n_6372), .B0 (n_7630), .Y(n_11419));
AND2X1 g65868(.A (n_7175), .B (n_11416), .Y (n_11417));
NAND2X2 g71413(.A (n_3460), .B (n_5349), .Y (n_11843));
AOI22X1 g65930(.A0 (n_11413), .A1 (n_16976), .B0 (n_11412), .B1(n_11307), .Y (n_11414));
NAND2X1 g65052(.A (n_5776), .B (n_15556), .Y (n_11411));
AOI21X1 g65968(.A0 (n_5217), .A1 (n_15588), .B0 (n_7090), .Y(n_11409));
AND2X1 g65969(.A (n_7184), .B (n_29102), .Y (n_11407));
AND2X1 g65972(.A (n_6914), .B (n_26276), .Y (n_11406));
AND2X1 g65976(.A (n_6831), .B (n_5531), .Y (n_11404));
INVX1 g65979(.A (n_9510), .Y (n_25791));
OR4X1 g65982(.A (n_276), .B (n_28757), .C (n_6546), .D (n_7725), .Y(n_17217));
NAND4X1 g65984(.A (n_28433), .B (n_27124), .C (n_28781), .D (n_4414),.Y (n_15626));
NOR2X1 g65989(.A (n_8251), .B (n_11400), .Y (n_11401));
NAND4X1 g65999(.A (n_17260), .B (n_4676), .C (n_29163), .D (n_4073),.Y (n_18941));
AND2X1 g66007(.A (n_8970), .B (n_9527), .Y (n_19355));
OR4X1 g66008(.A (n_17500), .B (n_11731), .C (n_3069), .D (n_7675), .Y(n_11397));
NOR2X1 g66010(.A (n_11394), .B (n_17260), .Y (n_11395));
NOR2X1 g66012(.A (n_17531), .B (n_27099), .Y (n_11393));
NOR2X1 g66016(.A (n_11390), .B (n_10495), .Y (n_11391));
NOR2X1 g66019(.A (n_10846), .B (n_27365), .Y (n_13092));
OR2X1 g66026(.A (n_8730), .B (n_17411), .Y (n_17228));
NOR2X1 g66031(.A (n_8176), .B (n_6534), .Y (n_11389));
NAND3X1 g66032(.A (n_4709), .B (n_6183), .C (n_10315), .Y (n_13556));
NAND3X1 g66033(.A (n_15968), .B (n_8729), .C (n_4113), .Y (n_17040));
NOR2X1 g66038(.A (n_11387), .B (n_6534), .Y (n_11388));
NOR2X1 g66042(.A (n_8736), .B (n_11312), .Y (n_13475));
NAND2X1 g66046(.A (n_11386), .B (n_11385), .Y (n_19428));
INVX1 g66060(.A (n_9497), .Y (n_13604));
OR2X1 g66066(.A (n_11383), .B (n_9527), .Y (n_11384));
NAND2X1 g69904(.A (n_7974), .B (n_7559), .Y (n_14139));
INVX1 g66072(.A (n_9491), .Y (n_13612));
NAND2X1 g66076(.A (n_11046), .B (n_7325), .Y (n_15463));
NOR2X1 g66079(.A (n_11381), .B (n_2318), .Y (n_13080));
NAND4X1 g66085(.A (n_9500), .B (n_11835), .C (n_27604), .D (n_4438),.Y (n_11380));
NOR2X1 g66091(.A (n_8552), .B (n_28381), .Y (n_11379));
NAND2X1 g66092(.A (n_9088), .B (n_14866), .Y (n_13524));
NOR2X1 g66096(.A (n_9056), .B (n_9388), .Y (n_13077));
INVX1 g66097(.A (n_11377), .Y (n_11378));
OR2X1 g66101(.A (n_11374), .B (n_12827), .Y (n_11375));
NOR2X1 g66105(.A (n_7414), .B (n_29286), .Y (n_11373));
INVX1 g66107(.A (n_11369), .Y (n_11371));
NAND2X1 g66110(.A (n_11367), .B (n_29228), .Y (n_11368));
NAND2X1 g66113(.A (n_8701), .B (n_14142), .Y (n_11366));
OR2X1 g66115(.A (n_11365), .B (n_16480), .Y (n_18633));
INVX2 g66121(.A (n_11363), .Y (n_15689));
NOR2X1 g66130(.A (n_11362), .B (n_9410), .Y (n_13069));
INVX1 g66132(.A (n_9483), .Y (n_16550));
NAND4X1 g66134(.A (n_5558), .B (n_28757), .C (n_7725), .D (n_6452),.Y (n_16758));
NAND2X1 g66136(.A (n_10747), .B (n_9819), .Y (n_11361));
NOR2X1 g66141(.A (n_8995), .B (n_12169), .Y (n_13067));
NOR2X1 g66143(.A (n_9523), .B (n_12169), .Y (n_11359));
INVX1 g66144(.A (n_9480), .Y (n_13588));
INVX1 g66149(.A (n_9477), .Y (n_11358));
INVX1 g66158(.A (n_9475), .Y (n_13066));
NOR2X1 g66163(.A (n_10827), .B (n_2779), .Y (n_11356));
NAND2X1 g66164(.A (n_8516), .B (n_11354), .Y (n_19955));
AND2X1 g66166(.A (n_11334), .B (n_9388), .Y (n_13064));
NAND2X1 g66167(.A (n_6093), .B (n_16466), .Y (n_11353));
INVX1 g66170(.A (n_9473), .Y (n_11351));
NAND3X1 g66172(.A (n_1424), .B (n_11350), .C (n_4695), .Y (n_15687));
NOR2X1 g66175(.A (n_16534), .B (n_6534), .Y (n_15590));
INVX1 g66179(.A (n_9471), .Y (n_11349));
INVX1 g66181(.A (n_29186), .Y (n_13554));
INVX1 g66182(.A (n_29185), .Y (n_11348));
NOR2X1 g66186(.A (n_11345), .B (n_6005), .Y (n_11346));
NAND2X1 g66191(.A (n_8713), .B (n_11307), .Y (n_15469));
NOR2X1 g66194(.A (n_8293), .B (n_18369), .Y (n_13056));
NAND2X1 g66196(.A (n_11367), .B (n_17260), .Y (n_11342));
NAND2X1 g66197(.A (n_8600), .B (n_13466), .Y (n_19953));
AND2X1 g66201(.A (n_8939), .B (n_18369), .Y (n_13054));
AOI21X1 g68671(.A0 (n_5450), .A1 (n_11215), .B0 (n_7191), .Y(n_11340));
NOR2X1 g66206(.A (n_11338), .B (n_18369), .Y (n_11339));
NAND2X1 g66213(.A (n_11278), .B (n_11731), .Y (n_11337));
NAND3X1 g66215(.A (n_29074), .B (n_2456), .C (n_10681), .Y (n_14972));
NAND2X1 g66219(.A (n_12827), .B (n_11334), .Y (n_11336));
NOR2X1 g66220(.A (n_15627), .B (n_11400), .Y (n_11333));
NOR2X1 g66224(.A (n_9033), .B (n_26883), .Y (n_13047));
AND2X1 g66236(.A (n_9114), .B (n_13815), .Y (n_11332));
NOR2X1 g68665(.A (n_6006), .B (n_6938), .Y (n_11331));
NOR2X1 g66245(.A (n_15640), .B (n_14142), .Y (n_11330));
NAND2X1 g66246(.A (n_8760), .B (n_9388), .Y (n_11329));
NOR2X1 g66247(.A (n_11327), .B (n_16480), .Y (n_11328));
NAND2X1 g66250(.A (n_15166), .B (n_13211), .Y (n_11326));
NOR2X1 g66255(.A (n_8997), .B (n_8941), .Y (n_11325));
NOR2X1 g66258(.A (n_11099), .B (n_6005), .Y (n_13042));
INVX1 g66261(.A (n_9457), .Y (n_13040));
OR4X1 g66263(.A (n_8435), .B (n_11323), .C (n_28459), .D (n_4573), .Y(n_11324));
NOR2X1 g66270(.A (n_29343), .B (n_11322), .Y (n_13035));
OR2X1 g66271(.A (n_11321), .B (n_13606), .Y (n_19291));
OR2X1 g66272(.A (n_12760), .B (n_7467), .Y (n_17990));
INVX1 g66276(.A (n_11318), .Y (n_14949));
INVX1 g66277(.A (n_11318), .Y (n_11319));
INVX1 g66283(.A (n_11317), .Y (n_13610));
NAND2X1 g66286(.A (n_8685), .B (n_9527), .Y (n_11316));
NAND2X1 g66287(.A (n_8818), .B (n_15708), .Y (n_11315));
INVX1 g66290(.A (n_9451), .Y (n_14845));
NOR2X1 g66293(.A (n_13320), .B (n_15610), .Y (n_11313));
NOR2X1 g66299(.A (n_9093), .B (n_9474), .Y (n_15156));
OR2X1 g66301(.A (n_9527), .B (n_8898), .Y (n_15196));
NAND2X1 g66307(.A (n_8478), .B (n_11312), .Y (n_15583));
OR2X1 g66308(.A (n_11731), .B (n_11311), .Y (n_16793));
NOR2X1 g66312(.A (n_7573), .B (n_8452), .Y (n_11309));
NAND2X1 g66320(.A (n_7077), .B (n_8865), .Y (n_17824));
NAND2X1 g66324(.A (n_7147), .B (n_9368), .Y (n_18801));
NOR2X1 g66326(.A (n_8486), .B (n_11307), .Y (n_13022));
NOR2X1 g66329(.A (n_11013), .B (n_12105), .Y (n_13020));
NOR2X1 g66333(.A (n_14940), .B (n_12105), .Y (n_13018));
NAND3X1 g66335(.A (n_11253), .B (n_10094), .C (n_8560), .Y (n_15488));
NOR2X1 g66342(.A (n_8454), .B (n_29062), .Y (n_13015));
NOR2X1 g66359(.A (n_11304), .B (n_15388), .Y (n_11305));
NOR2X1 g66365(.A (n_7436), .B (n_8974), .Y (n_11303));
NOR2X1 g66385(.A (n_11495), .B (n_10452), .Y (n_13008));
XOR2X1 g76328(.A (n_22569), .B (n_124), .Y (n_11302));
INVX1 g66394(.A (n_9433), .Y (n_14991));
OR2X1 g66399(.A (n_11300), .B (n_7305), .Y (n_12995));
NOR2X1 g66401(.A (n_12883), .B (n_14807), .Y (n_11299));
NOR2X1 g66404(.A (n_11298), .B (n_16754), .Y (n_12991));
INVX1 g66406(.A (n_11295), .Y (n_11296));
NAND2X1 g66410(.A (n_8414), .B (n_4898), .Y (n_12990));
OR2X1 g66412(.A (n_8708), .B (n_8681), .Y (n_17425));
INVX2 g66413(.A (n_9430), .Y (n_15513));
NOR2X1 g66418(.A (n_11292), .B (n_9942), .Y (n_12988));
NOR2X1 g66422(.A (n_11290), .B (n_12105), .Y (n_11291));
NAND2X1 g66424(.A (n_8431), .B (n_28418), .Y (n_14819));
OR4X1 g66427(.A (n_18237), .B (n_6219), .C (n_488), .D (n_4777), .Y(n_11288));
NOR2X1 g66429(.A (n_11285), .B (n_28642), .Y (n_11286));
NOR2X1 g66431(.A (n_8398), .B (n_28692), .Y (n_11284));
NOR2X1 g66434(.A (n_15825), .B (n_14807), .Y (n_11282));
NAND2X1 g66435(.A (n_8883), .B (n_15776), .Y (n_16990));
NOR2X1 g66439(.A (n_8184), .B (n_12979), .Y (n_11281));
INVX2 g70044(.A (n_8912), .Y (n_15087));
NOR2X1 g66443(.A (n_10987), .B (n_2260), .Y (n_12983));
NOR2X1 g66447(.A (n_7028), .B (n_15610), .Y (n_11280));
NAND2X1 g66448(.A (n_11278), .B (n_11277), .Y (n_11279));
NOR2X1 g66455(.A (n_27472), .B (n_9819), .Y (n_11275));
NOR2X1 g66471(.A (n_10919), .B (n_5799), .Y (n_15021));
NOR2X1 g66475(.A (n_11006), .B (n_9368), .Y (n_12968));
NOR2X1 g66485(.A (n_8944), .B (n_11272), .Y (n_11273));
NOR2X1 g66493(.A (n_8417), .B (n_5854), .Y (n_11271));
INVX1 g66501(.A (n_11579), .Y (n_12960));
NAND2X1 g66510(.A (n_28166), .B (n_13804), .Y (n_11267));
NAND2X1 g66514(.A (n_8907), .B (n_29062), .Y (n_11266));
INVX1 g66517(.A (n_11264), .Y (n_14961));
OR2X1 g66523(.A (n_11263), .B (n_5799), .Y (n_12957));
NOR2X1 g66526(.A (n_7110), .B (n_11261), .Y (n_11262));
NOR2X1 g66532(.A (n_11253), .B (n_11259), .Y (n_11260));
INVX1 g66539(.A (n_11257), .Y (n_11258));
INVX1 g66545(.A (n_11255), .Y (n_11256));
NOR2X1 g66554(.A (n_15340), .B (n_11253), .Y (n_11254));
INVX1 g66557(.A (n_9407), .Y (n_13416));
INVX1 g66578(.A (n_9403), .Y (n_12939));
INVX1 g66584(.A (n_11250), .Y (n_11251));
NOR2X1 g66588(.A (n_11249), .B (n_12559), .Y (n_12938));
AND2X1 g66600(.A (n_8870), .B (n_15776), .Y (n_11246));
NOR2X1 g66607(.A (n_9115), .B (n_9084), .Y (n_12934));
AND2X1 g66613(.A (n_11017), .B (n_17567), .Y (n_11244));
INVX1 g66620(.A (n_9390), .Y (n_11242));
NAND2X1 g66622(.A (n_11118), .B (n_11400), .Y (n_11241));
AND2X1 g66623(.A (n_10956), .B (n_29074), .Y (n_11240));
NOR2X1 g66625(.A (n_8433), .B (n_9819), .Y (n_11238));
OR2X1 g66627(.A (n_7244), .B (n_15986), .Y (n_11237));
NOR2X1 g66635(.A (n_11235), .B (n_28410), .Y (n_12926));
NAND2X1 g66636(.A (n_11233), .B (n_13083), .Y (n_11234));
OR2X1 g66639(.A (n_9526), .B (n_14866), .Y (n_12925));
NAND2X1 g66641(.A (n_7849), .B (n_9388), .Y (n_11231));
NOR2X1 g66644(.A (n_17297), .B (n_27604), .Y (n_11230));
OR2X1 g66647(.A (n_1424), .B (n_9000), .Y (n_12923));
OR2X1 g66648(.A (n_11228), .B (n_16787), .Y (n_19709));
NOR2X1 g66655(.A (n_8745), .B (n_9118), .Y (n_11227));
NOR2X1 g66658(.A (n_11321), .B (n_3318), .Y (n_12922));
NOR2X1 g66661(.A (n_9035), .B (n_27604), .Y (n_11224));
INVX1 g66664(.A (n_11549), .Y (n_11223));
INVX2 g70019(.A (n_9386), .Y (n_12012));
OR2X1 g66670(.A (n_18369), .B (n_8827), .Y (n_13414));
NOR2X1 g66675(.A (n_11221), .B (n_27688), .Y (n_11222));
NAND2X1 g66677(.A (n_9041), .B (n_20325), .Y (n_11220));
NOR2X1 g66684(.A (n_8354), .B (n_16434), .Y (n_11219));
INVX2 g66692(.A (n_9384), .Y (n_14956));
NOR2X1 g66699(.A (n_10964), .B (n_29065), .Y (n_11217));
NOR2X1 g66716(.A (n_8880), .B (n_17864), .Y (n_11214));
NOR2X1 g66722(.A (n_8643), .B (n_8679), .Y (n_12906));
NOR2X1 g66727(.A (n_8862), .B (n_6534), .Y (n_11213));
INVX1 g66731(.A (n_11211), .Y (n_19450));
NOR2X1 g66736(.A (n_8511), .B (n_28410), .Y (n_12903));
OR2X1 g66744(.A (n_9365), .B (n_11354), .Y (n_13495));
NOR2X1 g66746(.A (n_6980), .B (n_18320), .Y (n_11209));
NOR2X1 g66753(.A (n_9075), .B (n_11312), .Y (n_11208));
NAND2X1 g66754(.A (n_10889), .B (n_1424), .Y (n_11207));
NOR2X1 g66757(.A (n_14872), .B (n_29275), .Y (n_12900));
NOR2X1 g66760(.A (n_8691), .B (n_5558), .Y (n_11206));
INVX1 g66764(.A (n_11203), .Y (n_11204));
NOR2X1 g66770(.A (n_11200), .B (n_14055), .Y (n_12898));
OR2X1 g66780(.A (n_26372), .B (n_13318), .Y (n_18316));
INVX1 g66781(.A (n_9377), .Y (n_16570));
NOR2X1 g66786(.A (n_16527), .B (n_29256), .Y (n_11199));
NAND2X1 g66788(.A (n_11197), .B (n_13804), .Y (n_11198));
NOR2X1 g66791(.A (n_8298), .B (n_11322), .Y (n_11196));
NOR2X1 g66793(.A (n_8799), .B (n_1424), .Y (n_11195));
NOR2X1 g66795(.A (n_11193), .B (n_11322), .Y (n_11194));
NAND2X1 g66796(.A (n_10724), .B (n_13466), .Y (n_11192));
NOR2X1 g66803(.A (n_11190), .B (n_11731), .Y (n_11191));
NOR2X1 g66808(.A (n_10971), .B (n_28402), .Y (n_11189));
INVX2 g66809(.A (n_9374), .Y (n_15509));
NOR2X1 g66815(.A (n_7344), .B (n_4709), .Y (n_11188));
NOR2X1 g66819(.A (n_28410), .B (n_11186), .Y (n_13431));
NAND2X1 g66820(.A (n_9142), .B (n_5742), .Y (n_11185));
NAND2X1 g66821(.A (n_11533), .B (n_9472), .Y (n_11184));
NAND2X1 g66824(.A (n_10865), .B (n_8458), .Y (n_11183));
INVX1 g66825(.A (n_11181), .Y (n_11182));
INVX1 g66835(.A (n_27373), .Y (n_11179));
NAND2X1 g66839(.A (n_11177), .B (n_16988), .Y (n_11178));
NAND2X1 g66849(.A (n_11042), .B (n_7410), .Y (n_12879));
INVX1 g66855(.A (n_9369), .Y (n_12875));
NAND2X2 g66857(.A (n_13607), .B (n_29225), .Y (n_16704));
NOR2X1 g66859(.A (n_11175), .B (n_29244), .Y (n_13516));
NAND2X1 g66860(.A (n_11186), .B (n_3199), .Y (n_11173));
NAND2X1 g66861(.A (n_29176), .B (n_11172), .Y (n_13368));
INVX1 g66863(.A (n_14942), .Y (n_12872));
NAND2X1 g66866(.A (n_6441), .B (n_7414), .Y (n_11171));
NAND2X1 g66871(.A (n_9127), .B (n_7634), .Y (n_13559));
NAND2X1 g66881(.A (n_8746), .B (n_10495), .Y (n_12865));
NAND2X2 g66883(.A (n_10968), .B (n_11731), .Y (n_18335));
NAND2X1 g66891(.A (n_11565), .B (n_9509), .Y (n_11168));
OR2X1 g67313(.A (n_9527), .B (n_11087), .Y (n_21164));
NOR2X1 g66896(.A (n_28836), .B (n_12917), .Y (n_12862));
NAND2X1 g66907(.A (n_29363), .B (n_11165), .Y (n_11167));
NAND2X2 g66910(.A (n_10791), .B (n_26491), .Y (n_18645));
NAND2X1 g66915(.A (n_9555), .B (n_11190), .Y (n_11163));
INVX1 g66922(.A (n_9356), .Y (n_12855));
NAND2X1 g66925(.A (n_11197), .B (n_13872), .Y (n_12853));
NAND2X1 g66940(.A (n_6478), .B (n_11161), .Y (n_11162));
INVX1 g66946(.A (n_13567), .Y (n_11159));
NAND2X1 g66948(.A (n_11133), .B (n_11157), .Y (n_11158));
OR2X1 g66950(.A (n_10992), .B (n_13083), .Y (n_11156));
NAND2X1 g66953(.A (n_5161), .B (n_7344), .Y (n_11155));
AND2X1 g66956(.A (n_13220), .B (n_11338), .Y (n_12846));
INVX1 g66964(.A (n_11154), .Y (n_13585));
INVX1 g66967(.A (n_11151), .Y (n_11152));
INVX1 g66975(.A (n_15260), .Y (n_11150));
NOR2X1 g66984(.A (n_8714), .B (n_7410), .Y (n_12833));
NAND2X1 g66988(.A (n_11565), .B (n_17531), .Y (n_11146));
NAND2X1 g66992(.A (n_11144), .B (n_5867), .Y (n_11145));
NAND2X1 g66993(.A (n_19361), .B (n_10979), .Y (n_11143));
NAND2X1 g66996(.A (n_11141), .B (n_14878), .Y (n_11142));
INVX1 g67006(.A (n_11139), .Y (n_12825));
INVX1 g67012(.A (n_19216), .Y (n_11138));
NAND2X1 g67014(.A (n_9139), .B (n_9006), .Y (n_11137));
NAND2X1 g67021(.A (n_17762), .B (n_11133), .Y (n_11134));
OR2X1 g67023(.A (n_11516), .B (n_7325), .Y (n_13542));
NAND2X1 g67024(.A (n_11131), .B (n_5974), .Y (n_11132));
NOR2X1 g67030(.A (n_9456), .B (n_8679), .Y (n_12813));
NOR2X1 g67041(.A (n_8675), .B (n_8878), .Y (n_13484));
NAND2X1 g67046(.A (n_16480), .B (n_5850), .Y (n_12807));
AOI21X1 g67048(.A0 (n_4323), .A1 (n_5532), .B0 (n_11126), .Y(n_11127));
INVX1 g67049(.A (n_11124), .Y (n_11125));
NOR2X1 g67054(.A (n_11576), .B (n_11122), .Y (n_11123));
AND2X1 g67058(.A (n_10888), .B (n_12559), .Y (n_11120));
NAND2X1 g67063(.A (n_6436), .B (n_7573), .Y (n_11119));
NOR2X1 g67065(.A (n_11107), .B (n_9388), .Y (n_15276));
NAND2X1 g67072(.A (n_10820), .B (n_8660), .Y (n_11117));
INVX1 g67081(.A (n_14978), .Y (n_12792));
AND2X1 g67088(.A (n_11177), .B (n_14866), .Y (n_11116));
NAND2X1 g67089(.A (n_11114), .B (n_15825), .Y (n_11115));
NAND2X1 g67090(.A (n_11112), .B (n_11249), .Y (n_11113));
NAND2X1 g67093(.A (n_11110), .B (n_7181), .Y (n_11111));
NAND2X1 g67096(.A (n_4269), .B (n_8815), .Y (n_11109));
NAND2X1 g67097(.A (n_11131), .B (n_11107), .Y (n_11108));
NAND2X1 g67108(.A (n_5213), .B (n_17897), .Y (n_11106));
NAND3X1 g67109(.A (n_5532), .B (n_11104), .C (n_6062), .Y (n_11105));
AND2X1 g67110(.A (n_6824), .B (n_15574), .Y (n_11103));
INVX1 g72312(.A (n_11102), .Y (n_11756));
INVX1 g67122(.A (n_15019), .Y (n_11098));
NOR2X1 g67125(.A (n_11097), .B (n_17912), .Y (n_12776));
INVX1 g67126(.A (n_9334), .Y (n_15748));
NOR2X1 g67129(.A (n_9410), .B (n_5928), .Y (n_12774));
AND2X1 g67131(.A (n_15640), .B (n_13236), .Y (n_12772));
INVX1 g67134(.A (n_11096), .Y (n_16577));
INVX1 g67136(.A (n_11094), .Y (n_11095));
INVX1 g67154(.A (n_11091), .Y (n_11092));
NOR2X1 g67158(.A (n_11022), .B (n_13679), .Y (n_11089));
INVX2 g73036(.A (n_12275), .Y (n_11088));
NOR2X1 g67178(.A (n_11087), .B (n_7325), .Y (n_12745));
INVX1 g67180(.A (n_11086), .Y (n_12742));
NAND2X1 g67251(.A (n_15109), .B (n_11084), .Y (n_11085));
NAND2X1 g67184(.A (n_10784), .B (n_11307), .Y (n_12739));
OR2X1 g67185(.A (n_13521), .B (n_16480), .Y (n_11083));
NOR2X1 g67187(.A (n_11080), .B (n_19364), .Y (n_11081));
NAND2X1 g69968(.A (n_7913), .B (n_29221), .Y (n_14078));
AND2X1 g67194(.A (n_7483), .B (n_11078), .Y (n_11079));
NAND2X1 g67199(.A (n_11076), .B (n_12986), .Y (n_11077));
INVX1 g67200(.A (n_9325), .Y (n_11075));
AND2X1 g67217(.A (n_7808), .B (n_13083), .Y (n_11074));
INVX1 g67223(.A (n_9323), .Y (n_12725));
NAND2X1 g67243(.A (n_6065), .B (n_12648), .Y (n_11073));
NOR2X1 g67234(.A (n_8654), .B (n_8641), .Y (n_11072));
NAND2X1 g68587(.A (n_7059), .B (n_9227), .Y (n_11071));
NAND2X1 g67240(.A (n_4517), .B (n_8865), .Y (n_13366));
NAND2X1 g67249(.A (n_11165), .B (n_5928), .Y (n_13497));
NAND2X1 g67267(.A (n_11067), .B (n_9176), .Y (n_11068));
NAND2X1 g67268(.A (n_11065), .B (n_5805), .Y (n_11066));
NOR2X1 g67269(.A (n_11061), .B (n_9299), .Y (n_11064));
NAND2X1 g67277(.A (n_8924), .B (n_2810), .Y (n_13460));
NOR2X1 g67278(.A (n_8887), .B (n_11141), .Y (n_11063));
NOR2X1 g67279(.A (n_11061), .B (n_7315), .Y (n_11062));
INVX1 g67280(.A (n_13272), .Y (n_11060));
NOR2X1 g67286(.A (n_9524), .B (n_11312), .Y (n_12705));
INVX1 g67289(.A (n_9317), .Y (n_11059));
INVX1 g67298(.A (n_11057), .Y (n_11056));
OR2X1 g67306(.A (n_11165), .B (n_27365), .Y (n_12697));
NOR2X1 g67308(.A (n_11053), .B (n_11052), .Y (n_20926));
NAND2X1 g67315(.A (n_6414), .B (n_29074), .Y (n_11051));
NOR2X1 g67321(.A (n_10100), .B (n_11097), .Y (n_11050));
NOR2X1 g67323(.A (n_8481), .B (n_7930), .Y (n_11049));
NAND2X1 g67334(.A (n_6104), .B (n_14142), .Y (n_15700));
NAND2X1 g67335(.A (n_9071), .B (n_2720), .Y (n_25695));
NOR2X1 g67345(.A (n_9315), .B (n_11046), .Y (n_11047));
INVX1 g67350(.A (n_11045), .Y (n_17211));
INVX1 g67362(.A (n_28901), .Y (n_15180));
NOR2X1 g67368(.A (n_11043), .B (n_26877), .Y (n_13411));
NAND2X1 g67391(.A (n_11042), .B (n_12760), .Y (n_13429));
NAND2X1 g67394(.A (n_11040), .B (n_11228), .Y (n_11041));
NAND3X1 g67398(.A (n_6808), .B (n_4017), .C (n_13219), .Y (n_11039));
NOR2X1 g67403(.A (n_18266), .B (n_28836), .Y (n_12667));
AND2X1 g67405(.A (n_9509), .B (n_11473), .Y (n_11036));
INVX1 g67408(.A (n_11034), .Y (n_11035));
NOR2X1 g67415(.A (n_5723), .B (n_8496), .Y (n_11033));
NAND2X1 g67416(.A (n_11031), .B (n_11099), .Y (n_11032));
AND2X1 g67417(.A (n_7448), .B (n_11029), .Y (n_11030));
NAND2X1 g67425(.A (n_11027), .B (n_11731), .Y (n_11028));
INVX1 g67429(.A (n_11024), .Y (n_11025));
NOR2X1 g67434(.A (n_11022), .B (n_1512), .Y (n_11023));
NAND2X1 g67438(.A (n_11228), .B (n_9085), .Y (n_11021));
NAND2X1 g67443(.A (n_7296), .B (n_11097), .Y (n_13491));
NAND2X1 g67445(.A (n_11020), .B (n_12917), .Y (n_18353));
NAND2X1 g67447(.A (n_27900), .B (n_11228), .Y (n_11019));
NAND2X1 g67449(.A (n_11017), .B (n_12568), .Y (n_17177));
AND2X1 g67462(.A (n_14757), .B (n_13211), .Y (n_12641));
NAND2X1 g67463(.A (n_11015), .B (n_16754), .Y (n_20062));
NAND2X1 g67470(.A (n_7494), .B (n_11385), .Y (n_17754));
INVX1 g67475(.A (n_15159), .Y (n_14986));
NAND2X1 g67479(.A (n_4784), .B (n_11013), .Y (n_11014));
OR2X1 g67487(.A (n_18115), .B (n_9388), .Y (n_11012));
INVX1 g67499(.A (n_11011), .Y (n_13450));
INVX1 g67507(.A (n_13370), .Y (n_12617));
INVX1 g67510(.A (n_17757), .Y (n_12614));
INVX1 g67512(.A (n_15012), .Y (n_11010));
NOR2X1 g67522(.A (n_11008), .B (n_11323), .Y (n_12609));
NOR2X1 g67526(.A (n_8471), .B (n_11006), .Y (n_11007));
AND2X1 g67527(.A (n_7448), .B (n_4600), .Y (n_11005));
NAND2X1 g67529(.A (n_8876), .B (n_29074), .Y (n_11004));
NAND2X1 g67532(.A (n_28135), .B (n_10948), .Y (n_13402));
NOR2X1 g67543(.A (n_15388), .B (n_10812), .Y (n_12605));
NAND2X1 g67545(.A (n_11462), .B (n_10984), .Y (n_11002));
NAND2X1 g67551(.A (n_7205), .B (n_15574), .Y (n_11001));
NOR2X1 g67571(.A (n_10850), .B (n_29275), .Y (n_12589));
NAND2X1 g72982(.A (n_11694), .B (n_12144), .Y (n_11698));
NOR3X1 g61776(.A (n_7192), .B (n_10999), .C (n_25052), .Y (n_11000));
NAND2X1 g67574(.A (n_11287), .B (n_9034), .Y (n_10998));
NAND2X1 g67580(.A (n_9402), .B (n_10996), .Y (n_10997));
INVX1 g67586(.A (n_13725), .Y (n_12584));
NAND2X1 g67591(.A (n_13320), .B (n_13190), .Y (n_10995));
AND2X1 g67596(.A (n_10993), .B (n_10992), .Y (n_10994));
AOI21X1 g67604(.A0 (n_4109), .A1 (n_8951), .B0 (n_9819), .Y(n_10991));
INVX1 g67605(.A (n_9288), .Y (n_15738));
NOR2X1 g67613(.A (n_16754), .B (n_10834), .Y (n_12573));
NOR2X1 g67616(.A (n_10986), .B (n_4898), .Y (n_12572));
NAND2X1 g67624(.A (n_10945), .B (n_6082), .Y (n_12566));
NAND2X1 g67629(.A (n_4476), .B (n_10984), .Y (n_10985));
INVX1 g67635(.A (n_10982), .Y (n_10983));
NAND2X1 g67649(.A (n_10979), .B (n_13490), .Y (n_10980));
NOR2X1 g67653(.A (n_10607), .B (n_11013), .Y (n_10978));
NAND2X1 g67668(.A (n_8300), .B (n_7347), .Y (n_10977));
AND2X1 g67670(.A (n_14014), .B (n_10975), .Y (n_10976));
NAND2X1 g72903(.A (n_2227), .B (n_5114), .Y (n_10974));
INVX1 g67674(.A (n_13322), .Y (n_12553));
NAND2X1 g67683(.A (n_27642), .B (n_10971), .Y (n_10972));
NAND2X1 g67688(.A (n_11114), .B (n_12883), .Y (n_12544));
NAND2X1 g67692(.A (n_6448), .B (n_11290), .Y (n_10969));
INVX1 g67705(.A (n_9274), .Y (n_10967));
NOR2X1 g67709(.A (n_17411), .B (n_7634), .Y (n_12535));
NAND2X1 g67718(.A (n_11655), .B (n_13320), .Y (n_12533));
NAND2X1 g67720(.A (n_13607), .B (n_11300), .Y (n_14899));
INVX1 g67728(.A (n_15028), .Y (n_12531));
NAND2X1 g67737(.A (n_10964), .B (n_13181), .Y (n_13380));
NOR2X1 g67745(.A (n_7409), .B (n_9774), .Y (n_10962));
NAND2X1 g67760(.A (n_10959), .B (n_11006), .Y (n_10960));
AND2X1 g67763(.A (n_7408), .B (n_10957), .Y (n_25769));
NAND2X1 g67765(.A (n_11739), .B (n_10956), .Y (n_17180));
NAND2X1 g67769(.A (n_10369), .B (n_6874), .Y (n_10955));
NAND2X1 g67774(.A (n_11292), .B (n_28135), .Y (n_10954));
NOR2X1 g67777(.A (n_10952), .B (n_14484), .Y (n_12524));
NOR2X1 g67792(.A (n_10948), .B (n_11272), .Y (n_10949));
NAND2X1 g72964(.A (n_4046), .B (n_7598), .Y (n_11701));
OR2X1 g67809(.A (n_10945), .B (n_2260), .Y (n_12514));
AND2X1 g67812(.A (n_10943), .B (n_11087), .Y (n_12512));
INVX1 g67816(.A (n_9261), .Y (n_12510));
NAND2X1 g67820(.A (n_11107), .B (n_18115), .Y (n_10941));
NAND2X1 g67821(.A (n_6580), .B (n_7726), .Y (n_10940));
NAND2X1 g67827(.A (n_29065), .B (n_10939), .Y (n_20169));
NAND2X1 g67845(.A (n_10937), .B (n_10936), .Y (n_10938));
INVX1 g67846(.A (n_10934), .Y (n_10935));
NAND2X1 g67848(.A (n_8892), .B (n_28836), .Y (n_13445));
NAND2X1 g67849(.A (n_10932), .B (n_10931), .Y (n_10933));
NAND2X1 g67855(.A (n_11003), .B (n_28692), .Y (n_10930));
AND2X1 g67857(.A (n_8351), .B (n_263), .Y (n_10928));
NAND2X1 g67858(.A (n_11533), .B (n_17508), .Y (n_10927));
NAND2X1 g67861(.A (n_11292), .B (n_4435), .Y (n_10926));
NAND2X1 g67864(.A (n_8775), .B (n_5558), .Y (n_17939));
INVX1 g67881(.A (n_10923), .Y (n_10924));
NAND2X1 g67891(.A (n_10921), .B (n_9531), .Y (n_10922));
NAND2X1 g67892(.A (n_9406), .B (n_10919), .Y (n_10920));
INVX1 g67901(.A (n_10917), .Y (n_10918));
NAND2X1 g67911(.A (n_10915), .B (n_10914), .Y (n_10916));
OR2X1 g67919(.A (n_11172), .B (n_29048), .Y (n_20832));
NOR2X1 g67930(.A (n_15986), .B (n_10913), .Y (n_12476));
NOR2X1 g67931(.A (n_9286), .B (n_9389), .Y (n_10912));
AND2X1 g67933(.A (n_7378), .B (n_3449), .Y (n_10911));
AND2X1 g67939(.A (n_7378), .B (n_10909), .Y (n_10910));
INVX1 g67942(.A (n_9253), .Y (n_28556));
NOR2X1 g67945(.A (n_9637), .B (n_9565), .Y (n_10907));
NAND2X1 g67946(.A (n_10905), .B (n_10904), .Y (n_10906));
NOR2X1 g67951(.A (n_8671), .B (n_12169), .Y (n_12465));
AOI21X1 g67954(.A0 (n_3411), .A1 (n_8243), .B0 (n_29102), .Y(n_10903));
AOI21X1 g67956(.A0 (n_2548), .A1 (n_2839), .B0 (n_10393), .Y(n_10902));
NAND2X1 g67963(.A (n_10900), .B (n_27412), .Y (n_10901));
NAND2X1 g67982(.A (n_4225), .B (n_11006), .Y (n_10897));
NAND2X1 g67988(.A (n_8427), .B (n_4173), .Y (n_10896));
NOR2X1 g67990(.A (n_8287), .B (n_8319), .Y (n_29370));
INVX1 g68002(.A (n_10893), .Y (n_10894));
AND2X1 g68006(.A (n_7483), .B (n_8784), .Y (n_10892));
NOR2X1 g68009(.A (n_8743), .B (n_8330), .Y (n_10891));
NOR2X1 g68011(.A (n_10889), .B (n_10888), .Y (n_10890));
AOI21X1 g68015(.A0 (n_6489), .A1 (n_4403), .B0 (n_8708), .Y(n_10887));
INVX1 g68023(.A (n_9244), .Y (n_10883));
INVX1 g72241(.A (n_10882), .Y (n_14152));
NAND2X1 g68026(.A (n_10889), .B (n_1603), .Y (n_10881));
INVX1 g68038(.A (n_10880), .Y (n_13584));
NAND2X1 g68040(.A (n_8818), .B (n_11810), .Y (n_19033));
NAND2X1 g68041(.A (n_13172), .B (n_8285), .Y (n_10879));
NOR2X1 g68058(.A (n_9181), .B (n_8377), .Y (n_10876));
NAND2X1 g68059(.A (n_9064), .B (n_1340), .Y (n_25478));
NAND2X1 g68065(.A (n_10873), .B (n_27412), .Y (n_10874));
NAND2X1 g68067(.A (n_10870), .B (n_11287), .Y (n_10871));
NAND2X1 g68069(.A (n_10868), .B (n_13724), .Y (n_10869));
NAND2X1 g68075(.A (n_3964), .B (n_15352), .Y (n_10867));
INVX1 g72236(.A (n_8375), .Y (n_12414));
NOR2X1 g68112(.A (n_10900), .B (n_10389), .Y (n_12392));
NAND2X1 g68114(.A (n_16421), .B (n_10865), .Y (n_10866));
NAND2X1 g68116(.A (n_4205), .B (n_7002), .Y (n_10864));
NAND2X1 g68117(.A (n_16590), .B (n_15411), .Y (n_14969));
NAND2X1 g68119(.A (n_27412), .B (n_14330), .Y (n_10863));
INVX1 g69849(.A (n_10862), .Y (n_14464));
AOI21X1 g68472(.A0 (n_4434), .A1 (n_5803), .B0 (n_12827), .Y(n_10861));
NAND2X1 g68140(.A (n_10799), .B (n_11287), .Y (n_10860));
NAND2X1 g68144(.A (n_11020), .B (n_10859), .Y (n_16545));
NAND2X1 g68147(.A (n_10857), .B (n_10856), .Y (n_10858));
NOR2X1 g68149(.A (n_15894), .B (n_6879), .Y (n_12380));
NAND2X1 g68152(.A (n_3498), .B (n_10854), .Y (n_10855));
AND2X1 g68155(.A (n_9472), .B (n_13217), .Y (n_10853));
NOR2X1 g68169(.A (n_9060), .B (n_13458), .Y (n_25821));
OR2X1 g68170(.A (n_12631), .B (n_8217), .Y (n_10851));
NAND2X1 g68171(.A (n_8801), .B (n_10850), .Y (n_13564));
OR2X1 g68174(.A (n_26096), .B (n_9349), .Y (n_10849));
NAND2X1 g68182(.A (n_29363), .B (n_10846), .Y (n_10847));
NAND2X1 g68183(.A (n_28023), .B (n_10919), .Y (n_10845));
NOR2X1 g68185(.A (n_8833), .B (n_16434), .Y (n_10844));
OR2X1 g68188(.A (n_12751), .B (n_16466), .Y (n_10843));
NAND2X1 g68194(.A (n_14340), .B (n_10987), .Y (n_10842));
INVX1 g72922(.A (n_10841), .Y (n_15316));
NOR2X1 g68220(.A (n_6861), .B (n_8154), .Y (n_10840));
NAND2X1 g68223(.A (n_10838), .B (n_11385), .Y (n_10839));
NAND3X1 g68226(.A (n_6810), .B (n_3728), .C (n_10836), .Y (n_10837));
INVX1 g68245(.A (n_16568), .Y (n_15147));
NAND2X1 g68247(.A (n_10835), .B (n_10834), .Y (n_14958));
OR2X1 g68251(.A (n_10832), .B (n_12827), .Y (n_10833));
NAND2X1 g68252(.A (n_10830), .B (n_10996), .Y (n_10831));
NAND2X1 g68253(.A (n_6652), .B (n_6896), .Y (n_10829));
NOR2X1 g68272(.A (n_14902), .B (n_11322), .Y (n_15048));
NAND2X1 g68288(.A (n_3237), .B (n_10827), .Y (n_10828));
NAND2X2 g68291(.A (n_8586), .B (n_6005), .Y (n_12329));
NAND2X1 g68292(.A (n_8814), .B (n_7624), .Y (n_14936));
INVX1 g68294(.A (n_10825), .Y (n_10826));
INVX2 g68309(.A (n_10824), .Y (n_13443));
NAND2X1 g68312(.A (n_4232), .B (n_8170), .Y (n_10823));
NAND2X1 g68321(.A (n_6671), .B (n_11387), .Y (n_10822));
NOR2X1 g68326(.A (n_11144), .B (n_7598), .Y (n_12319));
NAND2X1 g68328(.A (n_15186), .B (n_10820), .Y (n_10821));
INVX1 g72904(.A (n_10819), .Y (n_15596));
NAND2X1 g68333(.A (n_10817), .B (n_10816), .Y (n_10818));
NAND2X2 g68337(.A (n_10815), .B (n_1424), .Y (n_18707));
NAND2X2 g68343(.A (n_11076), .B (n_29279), .Y (n_12312));
NAND2X1 g68345(.A (n_16416), .B (n_10812), .Y (n_13426));
NAND2X2 g68354(.A (n_16590), .B (n_8452), .Y (n_18286));
NAND2X1 g68355(.A (n_6540), .B (n_13776), .Y (n_10810));
NAND2X1 g68357(.A (n_7569), .B (n_9294), .Y (n_10809));
OR2X1 g68359(.A (n_10835), .B (n_7201), .Y (n_12301));
NAND2X1 g68366(.A (n_11031), .B (n_10835), .Y (n_10807));
NOR2X1 g68367(.A (n_10806), .B (n_7201), .Y (n_20910));
INVX1 g68369(.A (n_10805), .Y (n_12296));
INVX1 g68372(.A (n_13359), .Y (n_12294));
NAND2X1 g68386(.A (n_6604), .B (n_27445), .Y (n_10804));
NAND2X2 g68388(.A (n_26470), .B (n_5085), .Y (n_18051));
AOI21X1 g68389(.A0 (n_6479), .A1 (n_16198), .B0 (n_10815), .Y(n_10802));
INVX1 g68393(.A (n_10801), .Y (n_13595));
NOR2X1 g68397(.A (n_28427), .B (n_10799), .Y (n_13454));
OAI21X1 g68398(.A0 (n_1930), .A1 (n_6431), .B0 (n_10797), .Y(n_10798));
NAND2X1 g68402(.A (n_10795), .B (n_10794), .Y (n_10796));
NAND2X2 g68406(.A (n_27596), .B (n_7496), .Y (n_17832));
NOR2X1 g68418(.A (n_9333), .B (n_10791), .Y (n_10792));
NOR2X1 g72216(.A (n_3979), .B (n_9368), .Y (n_11764));
NOR2X1 g68422(.A (n_13724), .B (n_11276), .Y (n_12272));
NAND2X1 g68423(.A (n_7548), .B (n_10789), .Y (n_10790));
NAND2X1 g68426(.A (n_5512), .B (n_12500), .Y (n_10788));
INVX2 g68431(.A (n_9207), .Y (n_16676));
NAND2X1 g68438(.A (n_10784), .B (n_7158), .Y (n_10785));
NAND2X1 g68440(.A (n_10782), .B (n_7399), .Y (n_10783));
NAND3X1 g68444(.A (n_4417), .B (n_4295), .C (n_5421), .Y (n_10781));
NAND3X1 g68445(.A (n_4102), .B (n_3339), .C (n_3605), .Y (n_10780));
NAND3X1 g68447(.A (n_4499), .B (n_4140), .C (n_5456), .Y (n_10779));
OR2X1 g68450(.A (n_6940), .B (n_10777), .Y (n_10778));
OR2X1 g68452(.A (n_7667), .B (n_10775), .Y (n_10776));
AOI21X1 g68455(.A0 (n_3160), .A1 (n_6554), .B0 (n_11015), .Y(n_10774));
AOI21X1 g68460(.A0 (n_5232), .A1 (n_4017), .B0 (n_1530), .Y(n_10771));
AOI21X1 g68462(.A0 (n_4965), .A1 (n_3943), .B0 (n_19576), .Y(n_10770));
AOI21X1 g68468(.A0 (n_10768), .A1 (n_2583), .B0 (n_6816), .Y(n_10769));
NAND2X1 g68469(.A (n_7663), .B (n_28450), .Y (n_10767));
OAI21X1 g68478(.A0 (n_8978), .A1 (n_18237), .B0 (n_6772), .Y(n_10765));
OAI21X1 g68481(.A0 (n_5545), .A1 (n_17260), .B0 (n_7022), .Y(n_10763));
NAND2X1 g68484(.A (n_5780), .B (n_9116), .Y (n_10761));
NAND2X1 g68485(.A (n_5540), .B (n_7624), .Y (n_10760));
NAND2X1 g68487(.A (n_7818), .B (n_12546), .Y (n_10759));
AOI21X1 g68495(.A0 (n_5452), .A1 (n_9970), .B0 (n_15894), .Y(n_10758));
AOI21X1 g68496(.A0 (n_5369), .A1 (n_4837), .B0 (n_5850), .Y(n_10757));
AOI21X1 g68497(.A0 (n_5307), .A1 (n_3728), .B0 (n_2384), .Y(n_10756));
AOI21X1 g68498(.A0 (n_5237), .A1 (n_2923), .B0 (n_2385), .Y(n_10754));
AOI21X1 g68503(.A0 (n_4678), .A1 (n_7769), .B0 (n_263), .Y (n_10752));
NAND2X1 g68505(.A (n_6592), .B (n_14425), .Y (n_10751));
NAND2X1 g68508(.A (n_5398), .B (n_12563), .Y (n_10750));
OR2X1 g68511(.A (n_5009), .B (n_11365), .Y (n_10749));
NAND2X1 g68515(.A (n_7047), .B (n_12451), .Y (n_10748));
NAND2X1 g68532(.A (n_6537), .B (n_7634), .Y (n_10746));
NAND2X1 g68539(.A (n_6962), .B (n_10806), .Y (n_10745));
NAND2X1 g68546(.A (n_7239), .B (n_10986), .Y (n_10744));
NAND2X1 g68550(.A (n_6370), .B (n_12680), .Y (n_10743));
AOI21X1 g68557(.A0 (n_5011), .A1 (n_9511), .B0 (n_13804), .Y(n_10742));
AOI21X1 g68563(.A0 (n_5938), .A1 (n_9645), .B0 (n_13326), .Y(n_10741));
AOI21X1 g68565(.A0 (n_6376), .A1 (n_8392), .B0 (n_17411), .Y(n_10740));
NOR2X1 g68566(.A (n_7016), .B (n_8943), .Y (n_10738));
NAND2X1 g68570(.A (n_4265), .B (n_7595), .Y (n_10737));
NAND2X1 g68573(.A (n_8908), .B (n_29144), .Y (n_29129));
NAND2X1 g68577(.A (n_6531), .B (n_10734), .Y (n_10735));
AOI21X1 g68578(.A0 (n_3279), .A1 (n_10732), .B0 (n_2342), .Y(n_10733));
NAND2X1 g68588(.A (n_7026), .B (n_11053), .Y (n_10731));
NAND2X1 g68589(.A (n_7139), .B (n_7014), .Y (n_10730));
AOI21X1 g68591(.A0 (n_3816), .A1 (n_3306), .B0 (n_2215), .Y(n_10729));
AOI21X1 g68593(.A0 (n_1609), .A1 (n_3269), .B0 (n_4006), .Y(n_10728));
NOR2X1 g68606(.A (n_7382), .B (n_8406), .Y (n_10727));
AOI21X1 g68608(.A0 (n_5937), .A1 (n_8708), .B0 (n_7541), .Y(n_10726));
AOI21X1 g68616(.A0 (n_9163), .A1 (n_11312), .B0 (n_10724), .Y(n_10725));
AOI21X1 g68617(.A0 (n_5463), .A1 (n_28373), .B0 (n_6965), .Y(n_10723));
NAND2X1 g68618(.A (n_4625), .B (n_10720), .Y (n_10721));
NOR2X1 g68620(.A (n_7497), .B (n_8174), .Y (n_10719));
NOR2X1 g68623(.A (n_7492), .B (n_8658), .Y (n_10718));
AOI21X1 g68627(.A0 (n_10716), .A1 (n_14866), .B0 (n_18347), .Y(n_10717));
NOR2X1 g68636(.A (n_7434), .B (n_8652), .Y (n_10714));
NOR2X1 g68644(.A (n_7380), .B (n_8195), .Y (n_10713));
INVX1 g72884(.A (n_8203), .Y (n_15544));
NOR2X1 g68647(.A (n_7349), .B (n_7125), .Y (n_10712));
NAND2X1 g68652(.A (n_7346), .B (n_5871), .Y (n_10711));
AOI21X1 g68653(.A0 (n_5388), .A1 (n_14866), .B0 (n_5885), .Y(n_10710));
AOI21X1 g68659(.A0 (n_6689), .A1 (n_7496), .B0 (n_5812), .Y(n_10708));
NAND2X1 g68662(.A (n_7336), .B (n_7197), .Y (n_10707));
NOR2X1 g68663(.A (n_7332), .B (n_8550), .Y (n_10706));
NOR2X1 g68673(.A (n_7540), .B (n_8399), .Y (n_10705));
NAND2X1 g68681(.A (n_6447), .B (n_14085), .Y (n_10704));
NAND2X1 g68691(.A (n_6613), .B (n_11473), .Y (n_10703));
NAND2X1 g68694(.A (n_5164), .B (n_10701), .Y (n_10702));
AND2X1 g68696(.A (n_7130), .B (n_15588), .Y (n_10700));
OR2X1 g68703(.A (n_6282), .B (n_6857), .Y (n_10699));
OAI21X1 g68705(.A0 (n_5383), .A1 (n_7121), .B0 (n_2811), .Y(n_10698));
NAND2X1 g68716(.A (n_5156), .B (n_13190), .Y (n_10697));
NAND2X1 g72836(.A (n_19114), .B (n_12123), .Y (n_10696));
AND2X1 g68719(.A (n_6840), .B (n_14757), .Y (n_10694));
INVX1 g72868(.A (n_10693), .Y (n_11705));
NAND2X1 g68724(.A (n_6453), .B (n_10691), .Y (n_10692));
NAND3X1 g68725(.A (n_6987), .B (n_15507), .C (n_5151), .Y (n_10690));
NAND2X1 g68727(.A (n_5621), .B (n_10687), .Y (n_10688));
NAND2X1 g68729(.A (n_6837), .B (n_6281), .Y (n_10686));
OAI21X1 g68731(.A0 (n_3849), .A1 (n_7121), .B0 (n_9899), .Y(n_10685));
NAND2X1 g68732(.A (n_6850), .B (n_1988), .Y (n_10683));
OAI21X1 g68736(.A0 (n_6749), .A1 (n_10681), .B0 (n_10680), .Y(n_10682));
NAND2X1 g68738(.A (n_6834), .B (n_8018), .Y (n_10679));
AOI21X1 g68742(.A0 (n_16976), .A1 (n_3552), .B0 (n_8328), .Y(n_10678));
OAI21X1 g68745(.A0 (n_2215), .A1 (n_10676), .B0 (n_10675), .Y(n_10677));
NAND2X1 g68754(.A (n_6571), .B (n_17297), .Y (n_10674));
OAI21X1 g68762(.A0 (n_6694), .A1 (n_1333), .B0 (n_15659), .Y(n_10673));
OAI21X1 g68769(.A0 (n_5013), .A1 (n_4006), .B0 (n_11615), .Y(n_10672));
OAI21X1 g68773(.A0 (n_4712), .A1 (n_6767), .B0 (n_27472), .Y(n_10671));
OAI21X1 g68775(.A0 (n_6319), .A1 (n_2291), .B0 (n_13676), .Y(n_10670));
NAND2X1 g68779(.A (n_4376), .B (n_8929), .Y (n_10669));
NAND2X1 g68780(.A (n_6573), .B (n_27410), .Y (n_10668));
OAI21X1 g68787(.A0 (n_4408), .A1 (n_7193), .B0 (n_10191), .Y(n_10667));
AND2X1 g68788(.A (n_6721), .B (n_4512), .Y (n_10665));
AND2X1 g68791(.A (n_4381), .B (n_7108), .Y (n_10664));
AND2X1 g68795(.A (n_4246), .B (n_6976), .Y (n_10663));
AND2X1 g68797(.A (n_4714), .B (n_7190), .Y (n_10662));
AND2X1 g68799(.A (n_3966), .B (n_6369), .Y (n_10661));
AND2X1 g68800(.A (n_6610), .B (n_4135), .Y (n_10660));
AND2X1 g68801(.A (n_5269), .B (n_7061), .Y (n_10659));
AND2X1 g68803(.A (n_4281), .B (n_7025), .Y (n_10658));
AND2X1 g68804(.A (n_5172), .B (n_7828), .Y (n_10657));
AND2X1 g68805(.A (n_6464), .B (n_3601), .Y (n_10656));
XOR2X1 g68818(.A (n_1633), .B (n_5117), .Y (n_10655));
XOR2X1 g68819(.A (n_1253), .B (n_6121), .Y (n_10654));
XOR2X1 g68824(.A (n_1135), .B (n_5129), .Y (n_10653));
NAND2X1 g68988(.A (n_6393), .B (n_19398), .Y (n_10646));
NAND2X1 g72837(.A (n_8197), .B (n_6231), .Y (n_10645));
INVX1 g68999(.A (n_10640), .Y (n_19071));
INVX1 g69002(.A (n_10637), .Y (n_10638));
INVX2 g69006(.A (n_10635), .Y (n_15042));
INVX1 g69012(.A (n_10633), .Y (n_10634));
NAND2X1 g69014(.A (n_6459), .B (n_9084), .Y (n_10632));
INVX1 g69019(.A (n_18982), .Y (n_10631));
NAND2X1 g69036(.A (n_5202), .B (n_13593), .Y (n_10630));
AND2X1 g69043(.A (n_7794), .B (n_4689), .Y (n_10629));
NAND4X1 g69076(.A (n_14055), .B (n_4113), .C (n_3069), .D (n_10619),.Y (n_15714));
INVX1 g69078(.A (n_10621), .Y (n_10622));
NAND4X1 g69090(.A (n_1057), .B (n_3069), .C (n_7586), .D (n_10619),.Y (n_15350));
NOR2X1 g72128(.A (n_7664), .B (n_6997), .Y (n_10616));
INVX2 g69111(.A (n_7895), .Y (n_15326));
NAND2X1 g69116(.A (n_6688), .B (n_13318), .Y (n_14257));
NAND2X1 g69122(.A (n_6545), .B (n_19398), .Y (n_14358));
NOR2X1 g69126(.A (n_9691), .B (n_10610), .Y (n_12098));
NAND2X1 g69131(.A (n_9779), .B (n_8560), .Y (n_14442));
INVX1 g69136(.A (n_10609), .Y (n_14546));
OR2X1 g69139(.A (n_6429), .B (n_10607), .Y (n_10608));
NAND2X2 g69164(.A (n_8030), .B (n_1147), .Y (n_14384));
NOR2X1 g69177(.A (n_7942), .B (n_10599), .Y (n_10600));
INVX1 g69192(.A (n_10595), .Y (n_17325));
INVX2 g69219(.A (n_10590), .Y (n_15045));
INVX1 g69223(.A (n_10589), .Y (n_12081));
INVX1 g69229(.A (n_9094), .Y (n_17014));
INVX1 g69247(.A (n_10585), .Y (n_10586));
AND2X1 g69254(.A (n_6692), .B (n_9388), .Y (n_14535));
INVX1 g69267(.A (n_10581), .Y (n_12075));
OR2X1 g69271(.A (n_5147), .B (n_11052), .Y (n_10580));
INVX1 g69293(.A (n_10575), .Y (n_14585));
OR2X1 g69298(.A (n_10573), .B (n_28375), .Y (n_10574));
INVX1 g69310(.A (n_27475), .Y (n_10569));
INVX1 g69332(.A (n_10566), .Y (n_16439));
INVX1 g69353(.A (n_8071), .Y (n_12072));
NAND2X1 g69358(.A (n_9997), .B (n_11052), .Y (n_12070));
INVX1 g69370(.A (n_10561), .Y (n_10562));
NAND2X1 g69382(.A (n_7620), .B (n_15712), .Y (n_14513));
INVX1 g69389(.A (n_12409), .Y (n_14336));
INVX1 g69392(.A (n_14872), .Y (n_10556));
OR2X1 g69403(.A (n_10551), .B (n_11731), .Y (n_10552));
AND2X1 g69405(.A (n_7963), .B (n_28381), .Y (n_10550));
INVX1 g69410(.A (n_10549), .Y (n_12068));
NAND2X2 g69414(.A (n_9502), .B (n_14055), .Y (n_12067));
NAND2X1 g69428(.A (n_10546), .B (n_9368), .Y (n_10547));
INVX1 g69439(.A (n_10747), .Y (n_14308));
INVX1 g69447(.A (n_10542), .Y (n_10543));
INVX1 g69462(.A (n_9038), .Y (n_12063));
AND2X1 g69464(.A (n_6243), .B (n_8968), .Y (n_10537));
NAND2X1 g69466(.A (n_6717), .B (n_6005), .Y (n_10535));
NOR2X1 g69470(.A (n_7999), .B (n_11731), .Y (n_12060));
INVX2 g69479(.A (n_14803), .Y (n_10531));
INVX1 g69503(.A (n_10524), .Y (n_15575));
INVX1 g69528(.A (n_9021), .Y (n_17293));
INVX1 g69537(.A (n_9017), .Y (n_12058));
INVX1 g69539(.A (n_10522), .Y (n_10523));
NAND2X1 g69541(.A (n_7758), .B (n_20325), .Y (n_14252));
INVX1 g69544(.A (n_10521), .Y (n_13955));
INVX1 g69553(.A (n_10519), .Y (n_10520));
NAND2X1 g69556(.A (n_8047), .B (n_9118), .Y (n_10518));
NAND2X1 g69557(.A (n_10212), .B (n_9783), .Y (n_10516));
INVX1 g69559(.A (n_27403), .Y (n_10515));
AND2X1 g69567(.A (n_10513), .B (n_2318), .Y (n_10514));
NAND2X1 g69569(.A (n_6641), .B (n_27688), .Y (n_14325));
NAND2X1 g69580(.A (n_10777), .B (n_13593), .Y (n_10512));
INVX1 g69585(.A (n_10509), .Y (n_10510));
NAND2X1 g69588(.A (n_6355), .B (n_5329), .Y (n_10508));
INVX1 g69589(.A (n_10506), .Y (n_10507));
INVX1 g69610(.A (n_10501), .Y (n_10502));
NAND2X1 g69618(.A (n_6488), .B (n_10495), .Y (n_10496));
INVX1 g69620(.A (n_10492), .Y (n_10493));
INVX1 g69637(.A (n_10489), .Y (n_12052));
INVX1 g69641(.A (n_26797), .Y (n_10488));
INVX1 g69643(.A (n_10485), .Y (n_10486));
INVX1 g69645(.A (n_10483), .Y (n_10484));
INVX1 g69648(.A (n_10480), .Y (n_10481));
INVX1 g69656(.A (n_10476), .Y (n_13960));
INVX2 g69660(.A (n_10475), .Y (n_14188));
INVX1 g69662(.A (n_10472), .Y (n_10474));
INVX1 g69670(.A (n_10471), .Y (n_14571));
INVX1 g69683(.A (n_14528), .Y (n_10469));
INVX1 g69698(.A (n_10466), .Y (n_10467));
INVX1 g69705(.A (n_27671), .Y (n_10465));
NAND2X1 g69717(.A (n_29333), .B (n_8435), .Y (n_16599));
CLKBUFX1 g69729(.A (n_10463), .Y (n_12112));
NAND2X1 g69734(.A (n_6685), .B (n_15894), .Y (n_14433));
INVX1 g69748(.A (n_12715), .Y (n_10462));
AND2X1 g69762(.A (n_6427), .B (n_14113), .Y (n_10457));
NAND2X1 g69765(.A (n_10775), .B (n_8452), .Y (n_10456));
NAND2X1 g69766(.A (n_6594), .B (n_17414), .Y (n_14506));
INVX1 g69767(.A (n_10454), .Y (n_10455));
NAND2X2 g69773(.A (n_10453), .B (n_10452), .Y (n_14377));
INVX1 g69774(.A (n_10451), .Y (n_17683));
NAND2X1 g69787(.A (n_7141), .B (n_14484), .Y (n_10449));
INVX1 g69796(.A (n_10448), .Y (n_19690));
INVX1 g69804(.A (n_10447), .Y (n_12042));
INVX2 g69808(.A (n_10445), .Y (n_15177));
INVX1 g72072(.A (n_12416), .Y (n_11778));
AND2X1 g69819(.A (n_7799), .B (n_12105), .Y (n_10443));
INVX1 g69822(.A (n_12907), .Y (n_12036));
OR2X1 g69827(.A (n_10440), .B (n_28037), .Y (n_10441));
INVX1 g69833(.A (n_10437), .Y (n_10438));
INVX1 g69835(.A (n_12299), .Y (n_10436));
INVX1 g69838(.A (n_12322), .Y (n_10434));
INVX1 g69842(.A (n_10432), .Y (n_17037));
INVX2 g69855(.A (n_8948), .Y (n_14314));
INVX1 g69866(.A (n_8946), .Y (n_14141));
NAND2X1 g69878(.A (n_6356), .B (n_9264), .Y (n_10425));
INVX1 g69885(.A (n_10424), .Y (n_16342));
INVX1 g69891(.A (n_9265), .Y (n_14951));
NAND2X1 g69910(.A (n_5349), .B (n_9335), .Y (n_14284));
NAND2X1 g69911(.A (n_6734), .B (n_16974), .Y (n_25703));
NAND2X1 g69913(.A (n_9798), .B (n_7201), .Y (n_12028));
INVX1 g69914(.A (n_12885), .Y (n_10421));
NAND2X2 g69917(.A (n_10034), .B (n_9257), .Y (n_12026));
INVX1 g69927(.A (n_12495), .Y (n_17455));
INVX1 g69933(.A (n_12496), .Y (n_10418));
INVX1 g69939(.A (n_10415), .Y (n_10417));
INVX1 g69944(.A (n_10414), .Y (n_12025));
INVX1 g69946(.A (n_10413), .Y (n_15566));
INVX1 g69952(.A (n_10411), .Y (n_12024));
AND2X1 g69956(.A (n_6468), .B (n_12979), .Y (n_10410));
INVX1 g69957(.A (n_10408), .Y (n_17681));
NAND2X1 g69964(.A (n_28132), .B (n_7498), .Y (n_10407));
AND2X1 g69969(.A (n_9958), .B (n_5799), .Y (n_10405));
NAND2X1 g69972(.A (n_10081), .B (n_13490), .Y (n_12021));
INVX1 g69977(.A (n_10401), .Y (n_10402));
NAND2X1 g69979(.A (n_10020), .B (n_28445), .Y (n_10400));
INVX1 g69981(.A (n_10397), .Y (n_10398));
INVX1 g69987(.A (n_8927), .Y (n_14418));
INVX1 g69994(.A (n_8921), .Y (n_13398));
INVX1 g70000(.A (n_15105), .Y (n_14128));
AND2X1 g70015(.A (n_10355), .B (n_17500), .Y (n_10396));
NAND2X1 g70016(.A (n_6648), .B (n_1057), .Y (n_14344));
INVX1 g70023(.A (n_9429), .Y (n_14100));
INVX1 g70027(.A (n_11247), .Y (n_10395));
NOR2X1 g72056(.A (n_2548), .B (n_10393), .Y (n_12013));
INVX1 g70031(.A (n_28161), .Y (n_12009));
INVX1 g70035(.A (n_12359), .Y (n_10392));
NAND2X1 g70047(.A (n_10177), .B (n_10389), .Y (n_10390));
INVX1 g70049(.A (n_10387), .Y (n_14928));
NAND2X1 g70053(.A (n_6624), .B (n_27099), .Y (n_25813));
INVX1 g70054(.A (n_12206), .Y (n_14246));
INVX1 g70056(.A (n_9439), .Y (n_10385));
INVX1 g70065(.A (n_10382), .Y (n_10383));
INVX1 g70071(.A (n_10380), .Y (n_10381));
INVX1 g70076(.A (n_12175), .Y (n_19842));
NAND2X1 g70081(.A (n_6863), .B (n_16052), .Y (n_10377));
XOR2X1 g76107(.A (text_in_r[21] ), .B (n_6431), .Y (n_10376));
NAND2X1 g70091(.A (n_7810), .B (n_6534), .Y (n_10373));
AND2X1 g70095(.A (n_6600), .B (n_11731), .Y (n_10372));
NOR2X1 g70111(.A (n_28733), .B (n_10369), .Y (n_10370));
INVX1 g70117(.A (n_10366), .Y (n_10367));
INVX1 g70132(.A (n_10362), .Y (n_10361));
INVX1 g70135(.A (n_10358), .Y (n_10359));
INVX1 g70147(.A (n_12564), .Y (n_11994));
NAND2X1 g70156(.A (n_6533), .B (n_8708), .Y (n_14268));
NAND2X1 g70160(.A (n_10355), .B (n_15968), .Y (n_10356));
NAND2X1 g70162(.A (n_5408), .B (n_4689), .Y (n_10354));
INVX1 g70164(.A (n_12420), .Y (n_10353));
INVX1 g70166(.A (n_8888), .Y (n_16390));
INVX1 g73367(.A (n_11831), .Y (n_11658));
NAND2X1 g70182(.A (n_10030), .B (n_12559), .Y (n_10350));
INVX1 g70183(.A (n_12209), .Y (n_10348));
INVX1 g70185(.A (n_14390), .Y (n_10347));
NAND2X1 g70196(.A (n_10284), .B (n_15039), .Y (n_10346));
INVX2 g72767(.A (n_10345), .Y (n_11714));
INVX1 g70202(.A (n_12410), .Y (n_10344));
NAND2X1 g70206(.A (n_6530), .B (n_15039), .Y (n_10342));
INVX1 g70220(.A (n_19008), .Y (n_10341));
INVX1 g70227(.A (n_10338), .Y (n_10339));
INVX1 g70230(.A (n_10336), .Y (n_10337));
AND2X1 g70236(.A (n_10333), .B (n_9118), .Y (n_10334));
INVX1 g70245(.A (n_10332), .Y (n_11989));
AND2X1 g70251(.A (n_8035), .B (n_8452), .Y (n_10331));
INVX1 g70252(.A (n_10328), .Y (n_10329));
INVX1 g70259(.A (n_10327), .Y (n_16652));
AND2X1 g70262(.A (n_7934), .B (n_7496), .Y (n_10326));
INVX1 g70265(.A (n_10324), .Y (n_16338));
INVX1 g70272(.A (n_10323), .Y (n_14362));
INVX1 g70281(.A (n_10321), .Y (n_10322));
INVX1 g70289(.A (n_10319), .Y (n_10320));
NAND2X1 g70298(.A (n_6595), .B (n_7498), .Y (n_10318));
OR2X1 g72763(.A (n_7418), .B (n_10393), .Y (n_10317));
NOR2X1 g70314(.A (n_7944), .B (n_10315), .Y (n_10316));
INVX1 g70316(.A (n_10314), .Y (n_20626));
NAND2X1 g70329(.A (n_10312), .B (n_16198), .Y (n_10313));
INVX1 g70335(.A (n_10309), .Y (n_10311));
INVX1 g70342(.A (n_8842), .Y (n_17005));
INVX2 g70345(.A (n_10307), .Y (n_15011));
NAND2X1 g70357(.A (n_6599), .B (n_9860), .Y (n_10306));
NAND2X1 g69622(.A (n_10305), .B (n_6534), .Y (n_16068));
INVX1 g70369(.A (n_14981), .Y (n_10304));
INVX2 g70372(.A (n_10302), .Y (n_14616));
INVX1 g70380(.A (n_10299), .Y (n_14478));
NAND2X1 g70392(.A (n_9849), .B (n_29256), .Y (n_10296));
INVX1 g70394(.A (n_10295), .Y (n_11972));
OR2X1 g70396(.A (n_14386), .B (n_10389), .Y (n_10294));
INVX1 g70404(.A (n_8830), .Y (n_15682));
NOR2X1 g70408(.A (n_11400), .B (n_25665), .Y (n_10292));
NAND2X1 g70415(.A (n_5215), .B (n_8878), .Y (n_10290));
OR2X1 g70416(.A (n_5804), .B (n_12559), .Y (n_10289));
INVX1 g70417(.A (n_10287), .Y (n_10288));
NAND2X1 g70419(.A (n_9791), .B (n_15968), .Y (n_10286));
NOR2X1 g70430(.A (n_5289), .B (n_11312), .Y (n_11967));
NAND2X1 g70431(.A (n_10284), .B (n_10389), .Y (n_10285));
INVX1 g70434(.A (n_12285), .Y (n_10283));
INVX1 g70443(.A (n_10279), .Y (n_14130));
NAND2X1 g70448(.A (n_6586), .B (n_11731), .Y (n_10278));
AND2X1 g70449(.A (n_7921), .B (n_6005), .Y (n_10277));
OR2X1 g70450(.A (n_6344), .B (n_7325), .Y (n_16956));
NAND2X2 g70459(.A (n_10034), .B (n_8708), .Y (n_14044));
OR2X1 g70475(.A (n_10272), .B (n_12105), .Y (n_10273));
INVX1 g70477(.A (n_8813), .Y (n_14542));
INVX1 g70485(.A (n_10269), .Y (n_11958));
INVX1 g70488(.A (n_10269), .Y (n_14082));
INVX1 g70493(.A (n_10268), .Y (n_14537));
INVX1 g70502(.A (n_10266), .Y (n_10267));
INVX1 g70505(.A (n_10265), .Y (n_14222));
INVX1 g70514(.A (n_10264), .Y (n_11956));
INVX1 g70516(.A (n_12893), .Y (n_14526));
NAND2X1 g70529(.A (n_8240), .B (n_28744), .Y (n_11953));
CLKBUFX1 g70531(.A (n_8805), .Y (n_20628));
NAND2X1 g70534(.A (n_7950), .B (n_14484), .Y (n_10263));
INVX1 g70552(.A (n_8803), .Y (n_11949));
NAND2X2 g70555(.A (n_6724), .B (n_29297), .Y (n_13432));
NAND2X1 g70563(.A (n_8083), .B (n_8452), .Y (n_10258));
INVX1 g70567(.A (n_8801), .Y (n_14681));
INVX1 g70579(.A (n_10253), .Y (n_10254));
INVX1 g70581(.A (n_10251), .Y (n_10252));
NAND2X1 g70584(.A (n_9735), .B (n_11835), .Y (n_10250));
INVX1 g70586(.A (n_12397), .Y (n_11945));
INVX1 g70593(.A (n_12214), .Y (n_10249));
NOR2X1 g70597(.A (n_6681), .B (n_12559), .Y (n_10248));
INVX1 g70634(.A (n_12681), .Y (n_11940));
INVX1 g70636(.A (n_10243), .Y (n_10245));
INVX1 g70647(.A (n_10242), .Y (n_11936));
INVX1 g70656(.A (n_17405), .Y (n_10241));
INVX1 g70659(.A (n_17472), .Y (n_10239));
NAND2X1 g70663(.A (n_10237), .B (n_7649), .Y (n_10238));
NAND2X1 g70664(.A (n_2220), .B (n_5114), .Y (n_10235));
INVX1 g70673(.A (n_12154), .Y (n_11932));
INVX1 g70680(.A (n_14747), .Y (n_10231));
NOR2X1 g70686(.A (n_7966), .B (n_7598), .Y (n_11929));
INVX1 g70687(.A (n_10229), .Y (n_15055));
NAND2X1 g70696(.A (n_8674), .B (n_5202), .Y (n_18854));
INVX1 g70699(.A (n_8763), .Y (n_11925));
OR2X1 g70706(.A (n_7214), .B (n_10226), .Y (n_10227));
NAND2X1 g70709(.A (n_4136), .B (n_9118), .Y (n_11923));
NAND2X1 g70723(.A (n_7334), .B (n_10389), .Y (n_10222));
INVX1 g70725(.A (n_12581), .Y (n_10221));
NAND2X1 g70727(.A (n_4241), .B (n_16754), .Y (n_10220));
NOR2X1 g70729(.A (n_4393), .B (n_12019), .Y (n_11920));
NAND2X1 g70737(.A (n_10777), .B (n_9371), .Y (n_10218));
INVX1 g70750(.A (n_10217), .Y (n_11918));
NOR2X1 g70758(.A (n_11924), .B (n_27075), .Y (n_11917));
INVX1 g70768(.A (n_10216), .Y (n_11914));
INVX1 g70777(.A (n_8062), .Y (n_14193));
NAND2X1 g70795(.A (n_13837), .B (n_10212), .Y (n_10213));
INVX1 g70798(.A (n_10209), .Y (n_11909));
NOR2X1 g70801(.A (n_11110), .B (n_13593), .Y (n_10208));
INVX1 g70807(.A (n_10206), .Y (n_10207));
INVX1 g70820(.A (n_8735), .Y (n_10203));
NAND2X1 g70841(.A (n_3244), .B (n_5114), .Y (n_10201));
NAND2X1 g70842(.A (n_10199), .B (n_6586), .Y (n_14054));
NOR2X1 g70854(.A (n_6747), .B (n_6534), .Y (n_10197));
INVX1 g70864(.A (n_8723), .Y (n_16485));
INVX1 g70867(.A (n_10194), .Y (n_10195));
INVX1 g70879(.A (n_10193), .Y (n_11898));
NAND3X1 g70881(.A (n_6158), .B (n_10191), .C (n_3301), .Y (n_10192));
NAND2X1 g70891(.A (n_9351), .B (n_5202), .Y (n_10188));
NAND2X1 g70900(.A (n_7721), .B (n_5804), .Y (n_10183));
NAND2X1 g70918(.A (n_10181), .B (n_8637), .Y (n_11893));
NAND2X1 g70927(.A (n_4319), .B (n_17864), .Y (n_10180));
INVX1 g70928(.A (n_8712), .Y (n_14138));
NAND2X1 g70930(.A (n_9878), .B (n_6601), .Y (n_14482));
NAND2X1 g70943(.A (n_1928), .B (n_10177), .Y (n_10179));
INVX1 g70955(.A (n_10174), .Y (n_14321));
NOR2X1 g70959(.A (n_8022), .B (n_8540), .Y (n_10172));
INVX1 g70961(.A (n_10171), .Y (n_11889));
INVX1 g70967(.A (n_8702), .Y (n_10170));
NOR2X1 g70975(.A (n_5804), .B (n_8418), .Y (n_11886));
INVX1 g70976(.A (n_12541), .Y (n_10166));
INVX1 g70978(.A (n_8699), .Y (n_10165));
NOR2X1 g70983(.A (n_10163), .B (n_10162), .Y (n_10164));
NOR2X1 g70989(.A (n_8026), .B (n_6534), .Y (n_11884));
NOR2X1 g70993(.A (n_10160), .B (n_10125), .Y (n_11882));
NAND2X1 g71004(.A (n_10157), .B (n_14055), .Y (n_10158));
OR2X1 g71005(.A (n_6739), .B (n_9098), .Y (n_10156));
INVX1 g71006(.A (n_8690), .Y (n_28590));
NAND2X2 g71012(.A (n_7745), .B (n_10452), .Y (n_14380));
OR2X1 g71018(.A (n_6102), .B (n_4468), .Y (n_10154));
INVX1 g71019(.A (n_10152), .Y (n_15605));
INVX1 g71023(.A (n_10150), .Y (n_16678));
NOR2X1 g71982(.A (n_8086), .B (n_15968), .Y (n_10149));
AND2X1 g71039(.A (n_10147), .B (n_10146), .Y (n_11876));
NAND2X1 g71045(.A (n_9424), .B (n_8916), .Y (n_10142));
OR2X1 g71046(.A (n_10140), .B (n_1063), .Y (n_10141));
INVX1 g71047(.A (n_12256), .Y (n_10139));
NOR2X1 g71050(.A (n_4572), .B (n_1057), .Y (n_10138));
INVX1 g71051(.A (n_10137), .Y (n_20315));
INVX1 g71065(.A (n_12980), .Y (n_10135));
NAND2X1 g71071(.A (n_4112), .B (n_9410), .Y (n_10134));
NAND2X1 g71073(.A (n_4170), .B (n_17411), .Y (n_10133));
OR2X1 g71076(.A (n_10130), .B (n_14348), .Y (n_10131));
NAND2X1 g71085(.A (n_10127), .B (n_7810), .Y (n_14061));
NAND2X1 g68259(.A (n_10952), .B (n_3289), .Y (n_10126));
OR2X1 g71110(.A (n_10125), .B (n_28692), .Y (n_13971));
NAND2X1 g71117(.A (n_29191), .B (n_9264), .Y (n_10124));
INVX1 g71121(.A (n_8648), .Y (n_14447));
INVX1 g71133(.A (n_10119), .Y (n_10121));
NAND2X1 g71147(.A (n_11916), .B (n_5202), .Y (n_10115));
NAND2X1 g71162(.A (n_2811), .B (n_28862), .Y (n_20952));
INVX1 g71166(.A (n_10109), .Y (n_10110));
NOR2X1 g71169(.A (n_4778), .B (n_18100), .Y (n_10108));
NAND2X1 g71196(.A (n_4676), .B (n_10083), .Y (n_20950));
NAND2X1 g71201(.A (n_5951), .B (n_11731), .Y (n_10105));
OR2X1 g71214(.A (n_8086), .B (n_14155), .Y (n_14297));
INVX1 g71223(.A (n_10102), .Y (n_10104));
NAND2X2 g71226(.A (n_10101), .B (n_10100), .Y (n_14146));
OR2X1 g71228(.A (n_17841), .B (n_13606), .Y (n_10099));
NAND2X2 g71236(.A (n_7973), .B (n_7728), .Y (n_14405));
OR2X1 g71239(.A (n_4601), .B (n_15712), .Y (n_10098));
NOR2X1 g71253(.A (n_6516), .B (n_12019), .Y (n_10095));
NAND2X1 g71267(.A (n_3743), .B (n_5114), .Y (n_10093));
INVX1 g71274(.A (n_10091), .Y (n_11854));
NAND2X1 g71279(.A (n_2415), .B (n_5114), .Y (n_10090));
NAND2X1 g71280(.A (n_6377), .B (n_14155), .Y (n_10089));
AND2X1 g71289(.A (n_16006), .B (n_10094), .Y (n_11848));
INVX1 g71293(.A (n_8597), .Y (n_10088));
INVX1 g71295(.A (n_27716), .Y (n_10087));
NAND2X1 g71299(.A (n_10775), .B (n_17813), .Y (n_10085));
NAND2X1 g71304(.A (n_1378), .B (n_10083), .Y (n_10084));
NOR2X1 g71313(.A (n_4463), .B (n_10081), .Y (n_10082));
INVX1 g71328(.A (n_10078), .Y (n_10079));
NAND2X1 g71330(.A (n_3626), .B (n_10094), .Y (n_10077));
INVX1 g71339(.A (n_27707), .Y (n_10074));
INVX1 g71343(.A (n_10072), .Y (n_11845));
INVX1 g71346(.A (n_10071), .Y (n_14491));
OR2X1 g71363(.A (n_7968), .B (n_9106), .Y (n_10069));
INVX1 g71375(.A (n_10063), .Y (n_10065));
INVX1 g71378(.A (n_10061), .Y (n_10062));
NOR2X1 g70982(.A (n_9962), .B (n_16434), .Y (n_10060));
OR2X1 g71390(.A (n_12849), .B (n_7319), .Y (n_10058));
NAND2X1 g71400(.A (n_2420), .B (n_5114), .Y (n_10057));
INVX1 g71414(.A (n_8571), .Y (n_10053));
NAND2X1 g71418(.A (n_5571), .B (n_29256), .Y (n_10052));
INVX1 g71426(.A (n_14007), .Y (n_10051));
NAND2X1 g71431(.A (n_3896), .B (n_5114), .Y (n_10050));
INVX1 g71436(.A (n_16391), .Y (n_11842));
INVX1 g71944(.A (n_10049), .Y (n_11792));
INVX1 g71442(.A (n_17409), .Y (n_10048));
NAND2X1 g71461(.A (n_5671), .B (n_11253), .Y (n_10043));
INVX2 g71469(.A (n_8553), .Y (n_13383));
NAND2X1 g71471(.A (n_2732), .B (n_5114), .Y (n_10041));
INVX1 g71485(.A (n_10037), .Y (n_10038));
NOR2X1 g71487(.A (n_9708), .B (n_6583), .Y (n_10036));
INVX1 g71490(.A (n_10035), .Y (n_14598));
NAND2X1 g71493(.A (n_14725), .B (n_10034), .Y (n_14997));
NAND2X1 g71513(.A (n_28862), .B (n_10031), .Y (n_15104));
NOR2X1 g71519(.A (n_4771), .B (n_10030), .Y (n_11833));
AND2X1 g72662(.A (n_14107), .B (n_10083), .Y (n_11729));
NOR2X1 g71548(.A (n_5289), .B (n_17023), .Y (n_10029));
NAND2X1 g71550(.A (n_14107), .B (n_4963), .Y (n_10028));
INVX1 g71558(.A (n_8532), .Y (n_15628));
NAND2X1 g71572(.A (n_4380), .B (n_15039), .Y (n_10026));
NAND2X1 g71575(.A (n_6680), .B (n_5311), .Y (n_10025));
NAND2X1 g71584(.A (n_7023), .B (n_10020), .Y (n_28584));
INVX1 g71588(.A (n_13026), .Y (n_10018));
NAND2X1 g71591(.A (n_1565), .B (n_5114), .Y (n_10017));
NAND2X1 g71650(.A (n_4519), .B (n_11576), .Y (n_10008));
NAND2X1 g71663(.A (n_6490), .B (n_9486), .Y (n_17058));
INVX1 g71664(.A (n_8505), .Y (n_10003));
NAND2X1 g71674(.A (n_28156), .B (n_28410), .Y (n_11821));
OR2X1 g71677(.A (n_9999), .B (n_9543), .Y (n_10000));
NOR2X1 g71683(.A (n_6578), .B (n_8679), .Y (n_14017));
NAND2X1 g71684(.A (n_12836), .B (n_9997), .Y (n_28888));
NAND2X1 g71713(.A (n_4691), .B (n_12986), .Y (n_9996));
NAND2X1 g71715(.A (n_6492), .B (n_9838), .Y (n_14274));
INVX1 g71720(.A (n_8495), .Y (n_13550));
INVX1 g71737(.A (n_9993), .Y (n_15692));
INVX1 g71744(.A (n_7992), .Y (n_9992));
INVX1 g71746(.A (n_9990), .Y (n_9991));
INVX1 g71757(.A (n_9988), .Y (n_14600));
NAND2X1 g71778(.A (n_4484), .B (n_29102), .Y (n_9987));
INVX1 g71788(.A (n_8473), .Y (n_11808));
INVX1 g71790(.A (n_12945), .Y (n_14460));
INVX1 g72648(.A (n_8261), .Y (n_11805));
INVX1 g71810(.A (n_9980), .Y (n_9981));
NAND2X1 g71812(.A (n_4389), .B (n_9978), .Y (n_9979));
INVX1 g71817(.A (n_12823), .Y (n_9976));
INVX1 g71825(.A (n_8464), .Y (n_13518));
NAND2X1 g71827(.A (n_9772), .B (n_9970), .Y (n_14290));
INVX1 g71839(.A (n_17356), .Y (n_13976));
NAND2X1 g71852(.A (n_5508), .B (n_6653), .Y (n_9966));
NAND2X1 g71854(.A (n_9965), .B (n_10212), .Y (n_18827));
NOR2X1 g71862(.A (n_8000), .B (n_29065), .Y (n_25801));
INVX2 g71912(.A (n_9953), .Y (n_19529));
NOR2X1 g71867(.A (n_9962), .B (n_13593), .Y (n_9963));
NOR2X1 g71880(.A (n_10551), .B (n_2052), .Y (n_11799));
NOR2X1 g71882(.A (n_6607), .B (n_11307), .Y (n_14048));
INVX1 g71885(.A (n_12161), .Y (n_9961));
NAND2X1 g71888(.A (n_4969), .B (n_29256), .Y (n_9960));
NAND2X1 g71896(.A (n_9959), .B (n_9958), .Y (n_14413));
NAND2X1 g71902(.A (n_5554), .B (n_15388), .Y (n_9957));
INVX1 g71909(.A (n_9955), .Y (n_9956));
OR2X1 g71919(.A (n_3467), .B (n_6333), .Y (n_9952));
NAND2X1 g71926(.A (n_28862), .B (n_8997), .Y (n_9951));
NOR2X1 g71930(.A (n_7739), .B (n_8564), .Y (n_9950));
NAND2X1 g71939(.A (n_5368), .B (n_10573), .Y (n_9949));
INVX1 g71941(.A (n_8436), .Y (n_9948));
INVX1 g71953(.A (n_8590), .Y (n_15539));
OR2X1 g71955(.A (n_9999), .B (n_7821), .Y (n_9947));
NAND2X1 g71957(.A (n_9946), .B (n_9942), .Y (n_14392));
NAND2X1 g71970(.A (n_5614), .B (n_8928), .Y (n_9944));
NOR2X1 g71973(.A (n_5674), .B (n_9942), .Y (n_9943));
INVX1 g71976(.A (n_5806), .Y (n_19186));
OR2X1 g71983(.A (n_9939), .B (n_8227), .Y (n_9940));
AOI21X1 g62916(.A0 (n_5829), .A1 (n_9576), .B0 (n_4357), .Y (n_9938));
OR2X1 g72014(.A (n_4036), .B (n_12910), .Y (n_9937));
INVX1 g72015(.A (n_9935), .Y (n_9936));
CLKBUFX3 g72029(.A (n_9933), .Y (n_15395));
NOR2X1 g72049(.A (n_9930), .B (n_8191), .Y (n_9931));
NAND2X1 g72050(.A (n_4103), .B (n_18320), .Y (n_9929));
OR2X1 g72053(.A (n_7614), .B (n_9927), .Y (n_9928));
NAND2X1 g72061(.A (n_28812), .B (n_5854), .Y (n_14183));
NAND2X1 g72080(.A (n_9900), .B (n_6390), .Y (n_14242));
NOR2X1 g68207(.A (n_11172), .B (n_9923), .Y (n_9924));
OR2X1 g72086(.A (n_6521), .B (n_7185), .Y (n_9922));
INVX1 g72099(.A (n_12402), .Y (n_9921));
NOR2X1 g72104(.A (n_4171), .B (n_27604), .Y (n_9920));
NOR2X1 g72109(.A (n_6171), .B (n_9917), .Y (n_9918));
NAND2X1 g72123(.A (n_4127), .B (n_13326), .Y (n_9916));
NAND2X1 g72130(.A (n_9914), .B (n_10034), .Y (n_9915));
INVX1 g72133(.A (n_9913), .Y (n_11774));
NAND2X1 g72139(.A (n_6149), .B (n_5799), .Y (n_9912));
NAND2X1 g72152(.A (n_3791), .B (n_28862), .Y (n_20417));
INVX1 g72153(.A (n_15090), .Y (n_9911));
NAND2X1 g72156(.A (n_10305), .B (n_1361), .Y (n_9910));
NAND2X1 g72160(.A (n_6870), .B (n_5670), .Y (n_9909));
AND2X1 g72161(.A (n_5147), .B (n_9907), .Y (n_9908));
INVX1 g72189(.A (n_9906), .Y (n_12191));
INVX2 g72201(.A (n_8382), .Y (n_14028));
INVX1 g72221(.A (n_9903), .Y (n_9904));
OR2X1 g72225(.A (n_7899), .B (n_9900), .Y (n_9901));
INVX1 g72231(.A (n_16070), .Y (n_11762));
INVX1 g72233(.A (n_9896), .Y (n_9897));
OR2X1 g72254(.A (n_9714), .B (n_11731), .Y (n_9893));
INVX1 g72256(.A (n_12629), .Y (n_9892));
INVX1 g72259(.A (n_9262), .Y (n_9891));
INVX1 g72262(.A (n_9268), .Y (n_17744));
INVX1 g72285(.A (n_9298), .Y (n_12635));
OR2X1 g72295(.A (n_6450), .B (n_28427), .Y (n_9885));
NAND2X1 g72297(.A (n_3791), .B (n_5670), .Y (n_16715));
NAND2X1 g72299(.A (n_16006), .B (n_4945), .Y (n_9884));
INVX1 g72306(.A (n_9882), .Y (n_9883));
NAND2X1 g72315(.A (n_10146), .B (n_18266), .Y (n_19423));
OR2X1 g72328(.A (n_8706), .B (n_9878), .Y (n_9879));
INVX1 g72329(.A (n_9876), .Y (n_19297));
INVX1 g72350(.A (n_9874), .Y (n_9875));
INVX1 g72357(.A (n_8341), .Y (n_9873));
INVX1 g72363(.A (n_9872), .Y (n_13470));
INVX1 g72376(.A (n_12638), .Y (n_19799));
NAND2X1 g72381(.A (n_4827), .B (n_28645), .Y (n_9871));
INVX1 g72385(.A (n_9870), .Y (n_19862));
INVX1 g72388(.A (n_9869), .Y (n_14272));
INVX1 g72389(.A (n_9869), .Y (n_9868));
NAND2X1 g72397(.A (n_4614), .B (n_4689), .Y (n_9866));
NAND2X1 g72407(.A (n_10147), .B (n_4335), .Y (n_9864));
NAND2X1 g72412(.A (n_6505), .B (n_9295), .Y (n_9863));
NAND2X1 g72432(.A (n_7821), .B (n_9860), .Y (n_14186));
NAND2X1 g72449(.A (n_3460), .B (n_7950), .Y (n_14657));
NAND2X1 g72466(.A (n_2423), .B (n_5114), .Y (n_9858));
INVX1 g72469(.A (n_9856), .Y (n_14704));
OR2X1 g72491(.A (n_26457), .B (n_8437), .Y (n_9852));
NAND2X1 g72492(.A (n_27070), .B (n_9849), .Y (n_9850));
NAND2X1 g72495(.A (n_2701), .B (n_7995), .Y (n_18243));
OR2X1 g72498(.A (n_5884), .B (n_12849), .Y (n_9848));
OR2X1 g72506(.A (n_4962), .B (n_11272), .Y (n_9847));
OR2X1 g72507(.A (n_9699), .B (n_4689), .Y (n_9846));
AND2X1 g72513(.A (n_29115), .B (n_9844), .Y (n_9845));
NAND2X1 g72517(.A (n_4891), .B (n_15776), .Y (n_9843));
NAND2X1 g72518(.A (n_9841), .B (n_4689), .Y (n_9842));
NOR2X1 g72541(.A (n_4521), .B (n_9838), .Y (n_20178));
NOR2X1 g72550(.A (n_6731), .B (n_8452), .Y (n_9837));
OR2X1 g72555(.A (n_6747), .B (n_18237), .Y (n_14415));
INVX1 g72573(.A (n_12587), .Y (n_9835));
OR2X1 g72587(.A (n_28130), .B (n_26457), .Y (n_9834));
INVX1 g72588(.A (n_9831), .Y (n_9832));
INVX1 g72597(.A (n_9829), .Y (n_9830));
INVX1 g74638(.A (n_9651), .Y (n_13895));
INVX1 g72619(.A (n_8272), .Y (n_9827));
NAND2X1 g72635(.A (n_6743), .B (n_29102), .Y (n_9825));
NAND2X1 g72643(.A (n_9823), .B (n_29269), .Y (n_14093));
NAND2X1 g68164(.A (n_8477), .B (n_28402), .Y (n_9821));
OR2X1 g72657(.A (n_4256), .B (n_9417), .Y (n_11732));
NAND2X1 g72668(.A (n_14067), .B (n_17706), .Y (n_9820));
NAND2X1 g72677(.A (n_6791), .B (n_9819), .Y (n_18251));
INVX1 g72678(.A (n_8598), .Y (n_9818));
INVX1 g72680(.A (n_9815), .Y (n_9817));
INVX1 g72687(.A (n_8638), .Y (n_11725));
INVX1 g72702(.A (n_9811), .Y (n_19499));
INVX1 g72712(.A (n_8245), .Y (n_9810));
INVX2 g75776(.A (n_11823), .Y (n_11632));
INVX1 g72725(.A (n_9808), .Y (n_9809));
INVX1 g72736(.A (n_8239), .Y (n_9807));
NAND2X1 g72743(.A (n_4783), .B (n_11323), .Y (n_14216));
NAND2X1 g72753(.A (n_9804), .B (n_9803), .Y (n_9805));
INVX1 g72757(.A (n_9802), .Y (n_11975));
INVX1 g72773(.A (n_8231), .Y (n_16346));
AND2X1 g72778(.A (n_6245), .B (n_9800), .Y (n_9801));
NAND2X1 g72784(.A (n_2872), .B (n_9798), .Y (n_9799));
AND2X1 g72801(.A (n_9796), .B (n_9795), .Y (n_9797));
NAND2X1 g72802(.A (n_28862), .B (n_9106), .Y (n_19957));
NAND2X1 g72804(.A (n_1858), .B (n_5114), .Y (n_9794));
NAND2X1 g72819(.A (n_4700), .B (n_17775), .Y (n_9793));
INVX1 g72830(.A (n_8213), .Y (n_11712));
NAND2X1 g72835(.A (n_12858), .B (n_9791), .Y (n_9792));
INVX1 g72841(.A (n_9149), .Y (n_9790));
NAND2X2 g72845(.A (n_28609), .B (n_9368), .Y (n_11710));
AOI21X1 g63151(.A0 (n_6145), .A1 (n_11385), .B0 (n_6982), .Y(n_9789));
INVX1 g72860(.A (n_9787), .Y (n_11707));
INVX1 g72862(.A (n_9785), .Y (n_9786));
NAND2X1 g72882(.A (n_7925), .B (n_9783), .Y (n_9784));
INVX1 g72890(.A (n_8201), .Y (n_16351));
NAND2X1 g72900(.A (n_2043), .B (n_10081), .Y (n_9782));
NAND2X1 g72926(.A (n_13837), .B (n_9779), .Y (n_16280));
OR2X1 g72945(.A (n_9774), .B (n_6745), .Y (n_9775));
INVX1 g72955(.A (n_9773), .Y (n_14402));
NOR2X1 g72966(.A (n_4974), .B (n_9772), .Y (n_11700));
NOR2X1 g72987(.A (n_9927), .B (n_12559), .Y (n_9769));
NAND2X1 g72988(.A (n_1085), .B (n_7141), .Y (n_9767));
INVX1 g72990(.A (n_9765), .Y (n_11696));
OR2X1 g73008(.A (n_5975), .B (n_6759), .Y (n_9763));
NAND2X1 g73011(.A (n_2616), .B (n_5114), .Y (n_9762));
INVX1 g73060(.A (n_8161), .Y (n_15531));
NAND2X1 g73066(.A (n_9755), .B (n_12121), .Y (n_9756));
INVX1 g73067(.A (n_9372), .Y (n_16857));
NAND2X1 g73087(.A (n_29142), .B (n_27990), .Y (n_14577));
NAND2X1 g73099(.A (n_7911), .B (n_13593), .Y (n_9753));
INVX1 g73116(.A (n_9746), .Y (n_9748));
NOR2X1 g73130(.A (n_27991), .B (n_8139), .Y (n_9745));
NAND2X1 g73133(.A (n_6674), .B (n_7498), .Y (n_9743));
NAND2X1 g73134(.A (n_1706), .B (n_25440), .Y (n_9742));
NAND2X1 g73142(.A (n_6396), .B (n_13787), .Y (n_29178));
NAND2X1 g73143(.A (n_10083), .B (n_17260), .Y (n_19420));
NAND2X1 g73152(.A (n_4464), .B (n_9927), .Y (n_9739));
INVX1 g73153(.A (n_9737), .Y (n_9738));
NAND2X1 g73161(.A (n_6941), .B (n_9735), .Y (n_9736));
NAND2X1 g73162(.A (n_4963), .B (n_17706), .Y (n_9734));
NAND2X1 g73169(.A (n_26388), .B (n_11810), .Y (n_9732));
NAND2X1 g73176(.A (n_4335), .B (n_9371), .Y (n_9729));
INVX1 g73179(.A (n_9727), .Y (n_14463));
NAND2X1 g73187(.A (n_5638), .B (n_13247), .Y (n_9726));
INVX1 g73200(.A (n_9720), .Y (n_9721));
OR2X1 g73217(.A (n_6720), .B (n_9718), .Y (n_9719));
OR2X1 g73220(.A (n_6564), .B (n_9716), .Y (n_9717));
OR2X1 g73223(.A (n_3364), .B (n_9714), .Y (n_9715));
AOI21X1 g73226(.A0 (n_4736), .A1 (n_9712), .B0 (n_4079), .Y (n_9713));
NAND2X1 g73227(.A (n_6394), .B (n_7756), .Y (n_9711));
AOI21X1 g73228(.A0 (n_7610), .A1 (n_4334), .B0 (n_3003), .Y (n_9710));
OAI21X1 g73232(.A0 (n_9708), .A1 (n_3566), .B0 (n_14386), .Y(n_9709));
NAND2X1 g73233(.A (n_6635), .B (n_10272), .Y (n_9707));
NAND2X1 g73234(.A (n_6498), .B (n_6418), .Y (n_9706));
AOI21X1 g73241(.A0 (n_7095), .A1 (n_9704), .B0 (n_3502), .Y (n_9705));
NAND2X1 g73247(.A (n_3142), .B (n_29115), .Y (n_9703));
NAND2X1 g73253(.A (n_976), .B (n_6438), .Y (n_9702));
OR2X1 g73254(.A (n_6768), .B (n_2912), .Y (n_9701));
NOR2X1 g73259(.A (n_2216), .B (n_9699), .Y (n_9700));
AOI21X1 g73262(.A0 (n_2356), .A1 (n_5324), .B0 (n_2452), .Y (n_9698));
OAI21X1 g73266(.A0 (n_5946), .A1 (n_11835), .B0 (n_6589), .Y(n_9697));
OAI21X1 g73271(.A0 (n_4003), .A1 (n_28418), .B0 (n_6575), .Y(n_9696));
NAND2X1 g73273(.A (n_6678), .B (n_8759), .Y (n_9695));
AOI21X1 g73285(.A0 (n_9416), .A1 (n_3824), .B0 (n_6590), .Y (n_9694));
AOI21X1 g73286(.A0 (n_4261), .A1 (n_6497), .B0 (n_6803), .Y (n_9693));
AOI21X1 g73291(.A0 (n_9691), .A1 (n_2972), .B0 (n_6535), .Y (n_9692));
AOI21X1 g73292(.A0 (n_26880), .A1 (n_28542), .B0 (n_6361), .Y(n_9690));
AOI21X1 g73294(.A0 (n_27124), .A1 (n_1850), .B0 (n_7776), .Y(n_9688));
AOI21X1 g73297(.A0 (n_4721), .A1 (n_1065), .B0 (n_6802), .Y (n_9686));
AOI21X1 g73298(.A0 (n_4113), .A1 (n_4926), .B0 (n_7676), .Y (n_9685));
AOI21X1 g73299(.A0 (n_3807), .A1 (n_9682), .B0 (n_6469), .Y (n_9683));
AOI21X1 g73301(.A0 (n_28744), .A1 (n_2254), .B0 (n_6547), .Y(n_9681));
NAND2X1 g73623(.A (n_9481), .B (n_7485), .Y (n_13773));
INVX1 g73696(.A (n_11984), .Y (n_9676));
INVX1 g73709(.A (n_9675), .Y (n_13851));
INVX1 g73843(.A (n_27076), .Y (n_9674));
INVX1 g74026(.A (n_11801), .Y (n_9673));
NAND3X1 g74024(.A (n_3301), .B (n_6335), .C (n_7410), .Y (n_9672));
INVX1 g74099(.A (n_9668), .Y (n_11996));
INVX1 g74105(.A (n_28858), .Y (n_11649));
INVX1 g74378(.A (n_8012), .Y (n_9660));
INVX1 g74484(.A (n_11976), .Y (n_9656));
NAND3X1 g74721(.A (n_15473), .B (n_3667), .C (n_5817), .Y (n_9650));
AOI21X1 g60539(.A0 (n_6079), .A1 (n_13728), .B0 (n_25052), .Y(n_9649));
NAND3X1 g60540(.A (n_2848), .B (n_7860), .C (u0_r0_rcnt[0] ), .Y(n_9648));
INVX1 g74887(.A (n_12366), .Y (n_9647));
INVX1 g74906(.A (n_11734), .Y (n_9646));
NAND2X1 g72553(.A (n_5047), .B (n_9645), .Y (n_14213));
NAND2X1 g73255(.A (n_9419), .B (n_11350), .Y (n_9644));
NAND2X1 g71708(.A (n_6234), .B (n_28132), .Y (n_11819));
INVX1 g75199(.A (n_9640), .Y (n_9641));
INVX1 g75283(.A (n_9639), .Y (n_13909));
OR2X1 g75336(.A (n_9637), .B (n_6386), .Y (n_9638));
NOR2X1 g75460(.A (n_7792), .B (n_28134), .Y (n_9636));
INVX1 g69202(.A (n_9635), .Y (n_12085));
INVX2 g72526(.A (n_9632), .Y (n_15310));
NOR2X1 g75868(.A (n_6285), .B (n_2266), .Y (n_9629));
NOR2X1 g75891(.A (n_9195), .B (n_6373), .Y (n_9628));
NAND2X1 g73244(.A (n_4238), .B (n_10440), .Y (n_9627));
INVX1 g71638(.A (n_12349), .Y (n_9626));
XOR2X1 g76096(.A (n_9624), .B (n_5151), .Y (n_9625));
NOR2X1 g69134(.A (n_6754), .B (n_6534), .Y (n_12096));
XOR2X1 g76142(.A (n_23551), .B (n_15473), .Y (n_9621));
XOR2X1 g76160(.A (text_in_r[30] ), .B (n_5236), .Y (n_9619));
XOR2X1 g76182(.A (n_22546), .B (n_4582), .Y (n_9617));
OAI21X1 g64040(.A0 (n_5752), .A1 (n_7008), .B0 (n_15674), .Y(n_9615));
XOR2X1 g76216(.A (text_in_r[23] ), .B (n_3868), .Y (n_9614));
XOR2X1 g76229(.A (n_23087), .B (n_3038), .Y (n_9612));
XOR2X1 g76252(.A (text_in_r[7] ), .B (n_4837), .Y (n_9610));
XOR2X1 g76273(.A (text_in_r[14] ), .B (n_5305), .Y (n_9609));
XOR2X1 g76280(.A (text_in_r[5] ), .B (n_4750), .Y (n_9607));
NAND2X1 g73236(.A (n_6313), .B (n_6785), .Y (n_9605));
XOR2X1 g76333(.A (text_in_r[22] ), .B (n_5231), .Y (n_9604));
XOR2X1 g76346(.A (n_23547), .B (n_13679), .Y (n_9602));
XOR2X1 g76347(.A (text_in_r[13] ), .B (n_3038), .Y (n_9601));
AOI21X1 g64148(.A0 (n_7030), .A1 (n_9220), .B0 (n_16466), .Y(n_9599));
OR2X1 g64160(.A (n_15675), .B (n_13466), .Y (n_13753));
OR4X1 g64226(.A (n_17912), .B (n_16198), .C (n_5924), .D (n_4752), .Y(n_9597));
AOI21X1 g64252(.A0 (n_4219), .A1 (n_17508), .B0 (n_26670), .Y(n_9596));
NAND2X1 g64288(.A (n_13316), .B (n_13776), .Y (n_9595));
NAND2X1 g64309(.A (n_8176), .B (n_9593), .Y (n_9594));
NAND2X1 g69025(.A (n_14067), .B (n_29244), .Y (n_9592));
NAND2X1 g67870(.A (n_8850), .B (n_5454), .Y (n_9590));
INVX1 g75313(.A (n_9587), .Y (n_9588));
OAI21X1 g64376(.A0 (n_5012), .A1 (n_9585), .B0 (n_5131), .Y (n_9586));
OR2X1 g64405(.A (n_14868), .B (n_14866), .Y (n_13763));
NAND3X1 g64411(.A (n_5532), .B (n_4343), .C (n_11620), .Y (n_9584));
NAND3X1 g64415(.A (n_7381), .B (n_5765), .C (n_7555), .Y (n_9582));
NAND2X1 g64463(.A (n_7687), .B (n_20010), .Y (n_9581));
NAND2X1 g64497(.A (n_7771), .B (n_15655), .Y (n_9580));
NAND2X1 g64512(.A (n_18895), .B (n_11507), .Y (n_9579));
AND2X1 g64565(.A (n_11516), .B (n_9576), .Y (n_9577));
NAND3X1 g64567(.A (n_9574), .B (n_9573), .C (n_4412), .Y (n_9575));
OAI21X1 g64571(.A0 (n_5174), .A1 (n_15465), .B0 (n_124), .Y (n_9572));
DFFX1 dcnt_reg[0] (.CK (clk), .D (n_6421), .Q (dcnt[0] ), .QN ());
OAI21X1 g64631(.A0 (n_5601), .A1 (n_17491), .B0 (n_27216), .Y(n_9569));
NAND3X1 g64690(.A (n_11263), .B (n_9567), .C (n_9414), .Y (n_9568));
NAND3X1 g64737(.A (n_9565), .B (n_9564), .C (n_3248), .Y (n_9566));
DFFX1 u0_r0_rcnt_reg[3] (.CK (clk), .D (n_7806), .Q (u0_r0_rcnt[3]), .QN ());
NAND2X1 g64751(.A (n_9538), .B (n_15986), .Y (n_11486));
NAND2X1 g64772(.A (n_8184), .B (n_9561), .Y (n_9562));
NAND2X1 g64786(.A (n_8462), .B (n_9559), .Y (n_9560));
AOI21X1 g64792(.A0 (n_5680), .A1 (n_9557), .B0 (n_15039), .Y(n_9558));
INVX1 g75884(.A (n_9555), .Y (n_9556));
NAND2X1 g73202(.A (n_9552), .B (n_6746), .Y (n_9553));
INVX1 g66154(.A (n_9550), .Y (n_18614));
NOR2X1 g70374(.A (n_7496), .B (n_6337), .Y (n_10302));
NAND2X1 g73193(.A (n_2954), .B (n_8520), .Y (n_9549));
AOI21X1 g65072(.A0 (n_4597), .A1 (n_9547), .B0 (n_27133), .Y(n_9548));
NAND2X1 g72456(.A (n_3419), .B (n_8520), .Y (n_9545));
AND2X1 g74888(.A (n_9899), .B (n_8016), .Y (n_12366));
OR2X1 g71530(.A (n_7813), .B (n_5569), .Y (n_9541));
NAND2X1 g67633(.A (n_7797), .B (n_7331), .Y (n_11484));
INVX1 g67627(.A (n_9538), .Y (n_9539));
AND2X1 g73184(.A (n_1361), .B (n_28991), .Y (n_9537));
INVX1 g73180(.A (n_9534), .Y (n_9727));
NAND2X2 g67587(.A (n_9260), .B (n_10452), .Y (n_13725));
NAND2X1 g67589(.A (n_3567), .B (n_9531), .Y (n_9532));
NAND2X2 g70148(.A (n_8250), .B (n_6534), .Y (n_12564));
INVX1 g73166(.A (n_6849), .Y (n_14087));
AOI21X1 g65508(.A0 (n_9529), .A1 (n_9528), .B0 (n_9527), .Y (n_9530));
NAND2X1 g73164(.A (n_5197), .B (n_16414), .Y (n_12506));
OAI21X1 g68768(.A0 (n_11413), .A1 (n_7100), .B0 (n_1531), .Y(n_9525));
OR2X1 g73154(.A (n_6725), .B (n_29256), .Y (n_9737));
INVX1 g71448(.A (n_9524), .Y (n_10046));
INVX1 g73148(.A (n_9523), .Y (n_16290));
NOR2X1 g70136(.A (n_9522), .B (n_6219), .Y (n_10358));
INVX1 g72041(.A (n_8884), .Y (n_12997));
NAND2X1 g67476(.A (n_27411), .B (n_8263), .Y (n_15159));
NOR2X1 g71405(.A (n_3329), .B (n_28692), .Y (n_9515));
OR2X1 g70096(.A (n_9513), .B (n_1057), .Y (n_9514));
NAND2X1 g72386(.A (n_6931), .B (n_6420), .Y (n_9870));
NAND2X1 g72379(.A (n_7429), .B (n_9511), .Y (n_12478));
NOR2X1 g65980(.A (n_9509), .B (n_15712), .Y (n_9510));
NAND3X1 g65985(.A (n_11576), .B (n_4466), .C (n_28373), .Y (n_9508));
NAND4X1 g65993(.A (n_28433), .B (n_27124), .C (n_28780), .D (n_5612),.Y (n_13706));
OR2X1 g65994(.A (n_9504), .B (n_18369), .Y (n_9505));
INVX1 g75200(.A (n_9502), .Y (n_9640));
NAND4X1 g66013(.A (n_7266), .B (n_7601), .C (n_28476), .D (n_2447),.Y (n_11567));
INVX1 g66039(.A (n_15243), .Y (n_9501));
NAND4X1 g66044(.A (n_9500), .B (n_27604), .C (n_2124), .D (n_6486),.Y (n_15225));
OR2X1 g66047(.A (n_7206), .B (n_7410), .Y (n_11506));
NAND3X1 g66051(.A (n_9118), .B (n_7367), .C (n_7636), .Y (n_11560));
NAND4X1 g66053(.A (n_11276), .B (n_8910), .C (n_7734), .D (n_5154),.Y (n_16663));
NAND4X1 g66061(.A (n_11312), .B (n_3307), .C (n_9467), .D (n_4764),.Y (n_9497));
NAND2X1 g66062(.A (n_7473), .B (n_11322), .Y (n_13508));
NOR2X1 g66068(.A (n_17619), .B (n_11354), .Y (n_9495));
NAND4X1 g66069(.A (n_15894), .B (n_6534), .C (n_6303), .D (n_3718),.Y (n_28591));
NOR2X1 g66073(.A (n_9573), .B (n_8679), .Y (n_9491));
INVX1 g66081(.A (n_13537), .Y (n_9489));
NAND2X1 g66083(.A (n_14534), .B (n_12827), .Y (n_19951));
AND2X1 g66099(.A (n_7355), .B (n_12827), .Y (n_11377));
NOR2X1 g66109(.A (n_18635), .B (n_12827), .Y (n_11369));
NAND4X1 g66119(.A (n_9486), .B (n_3807), .C (n_3464), .D (n_5148), .Y(n_17456));
NOR2X1 g66122(.A (n_10100), .B (n_7489), .Y (n_11363));
NOR2X1 g66133(.A (n_11500), .B (n_12169), .Y (n_9483));
INVX1 g72368(.A (n_11022), .Y (n_13052));
INVX1 g77729(.A (n_9481), .Y (n_9482));
NOR2X1 g66145(.A (n_13532), .B (n_8878), .Y (n_9480));
NAND4X1 g66146(.A (n_12986), .B (n_8090), .C (n_29166), .D (n_27072),.Y (n_9479));
NOR2X1 g66150(.A (n_27710), .B (n_15776), .Y (n_9477));
NOR2X1 g66159(.A (n_9574), .B (n_9474), .Y (n_9475));
INVX1 g73710(.A (n_6775), .Y (n_9675));
NOR2X1 g66171(.A (n_9472), .B (n_12910), .Y (n_9473));
OR4X1 g66178(.A (n_26041), .B (n_11322), .C (n_2124), .D (n_4030), .Y(n_13291));
NOR2X1 g66180(.A (n_17508), .B (n_17567), .Y (n_9471));
NAND2X1 g66187(.A (n_7278), .B (n_27365), .Y (n_13452));
AND2X1 g66188(.A (n_9469), .B (n_9342), .Y (n_13156));
NAND4X1 g66189(.A (n_11312), .B (n_3307), .C (n_9467), .D (n_3053),.Y (n_18361));
OR2X1 g66204(.A (n_9465), .B (n_13606), .Y (n_9466));
OR2X1 g66205(.A (n_6051), .B (n_7496), .Y (n_13695));
OR2X1 g66209(.A (n_10794), .B (n_11312), .Y (n_13213));
NAND4X1 g66216(.A (n_9410), .B (n_4261), .C (n_28472), .D (n_6142),.Y (n_15503));
NAND2X1 g71388(.A (n_9463), .B (n_13593), .Y (n_9464));
NAND2X1 g66225(.A (n_9404), .B (n_28398), .Y (n_13469));
OR4X1 g66226(.A (n_18266), .B (n_4709), .C (n_16204), .D (n_3106), .Y(n_9462));
NAND3X1 g66227(.A (n_8679), .B (n_7182), .C (n_2632), .Y (n_11512));
NAND4X1 g66232(.A (n_263), .B (n_2811), .C (n_2368), .D (n_9415), .Y(n_18142));
NAND2X1 g66251(.A (n_9459), .B (n_11354), .Y (n_9460));
NOR2X1 g66262(.A (n_7157), .B (n_12169), .Y (n_9457));
INVX1 g73114(.A (n_9456), .Y (n_9750));
NAND2X1 g66267(.A (n_7668), .B (n_6534), .Y (n_15111));
NOR2X1 g66278(.A (n_11431), .B (n_10100), .Y (n_11318));
OR2X1 g66279(.A (n_17286), .B (n_8679), .Y (n_13207));
OR4X1 g66281(.A (n_263), .B (n_10031), .C (n_9089), .D (n_3144), .Y(n_15222));
NOR2X1 g66284(.A (n_9319), .B (n_14866), .Y (n_11317));
NOR2X1 g66291(.A (n_9450), .B (n_9474), .Y (n_9451));
OR2X1 g66294(.A (n_9450), .B (n_9527), .Y (n_19299));
NAND2X1 g66300(.A (n_7504), .B (n_13083), .Y (n_9449));
INVX1 g66302(.A (n_9446), .Y (n_15034));
INVX1 g66313(.A (n_13421), .Y (n_9445));
INVX1 g73698(.A (n_8063), .Y (n_9444));
NAND4X1 g66321(.A (n_4689), .B (n_9442), .C (n_9392), .D (n_3664), .Y(n_13329));
INVX1 g66337(.A (n_9440), .Y (n_14909));
NAND2X1 g70055(.A (n_4215), .B (n_6462), .Y (n_12206));
NOR2X1 g70057(.A (n_8127), .B (n_5799), .Y (n_9439));
INVX1 g66380(.A (n_14770), .Y (n_9437));
NAND2X1 g72361(.A (n_13730), .B (n_7649), .Y (n_9436));
OR2X1 g66387(.A (n_9435), .B (n_11276), .Y (n_15121));
NAND2X1 g66391(.A (n_7064), .B (n_6005), .Y (n_13408));
NOR2X1 g66395(.A (n_7421), .B (n_2260), .Y (n_9433));
OR4X1 g66407(.A (n_11261), .B (n_1584), .C (n_488), .D (n_5457), .Y(n_11295));
NAND2X1 g66411(.A (n_17477), .B (n_18168), .Y (n_9431));
NOR2X1 g66414(.A (n_11031), .B (n_352), .Y (n_9430));
NOR2X1 g70024(.A (n_29140), .B (n_27990), .Y (n_9429));
OR2X1 g72332(.A (n_8120), .B (n_6534), .Y (n_9428));
OR2X1 g66445(.A (n_9425), .B (n_13083), .Y (n_9426));
NAND2X1 g66446(.A (n_7269), .B (n_9118), .Y (n_14823));
NAND4X1 g66462(.A (n_6008), .B (n_6462), .C (n_3081), .D (n_3702), .Y(n_13382));
NAND2X1 g66466(.A (n_9418), .B (n_7496), .Y (n_13385));
INVX1 g75875(.A (n_9419), .Y (n_9420));
OR2X1 g66480(.A (n_7354), .B (n_18320), .Y (n_15681));
NAND2X1 g66488(.A (n_9418), .B (n_17414), .Y (n_16737));
NAND4X1 g66494(.A (n_9417), .B (n_9416), .C (n_2368), .D (n_9415), .Y(n_15538));
OR2X1 g66502(.A (n_5851), .B (n_8878), .Y (n_11579));
INVX1 g66508(.A (n_7718), .Y (n_13295));
OR4X1 g66515(.A (n_11400), .B (n_28418), .C (n_28781), .D (n_4015),.Y (n_13305));
NOR2X1 g66519(.A (n_4689), .B (n_9414), .Y (n_11264));
OR2X1 g70029(.A (n_6409), .B (n_9118), .Y (n_11247));
OR2X1 g66540(.A (n_14624), .B (n_5960), .Y (n_11257));
NAND2X1 g66542(.A (n_7602), .B (n_5854), .Y (n_14996));
OR2X1 g66546(.A (n_9410), .B (n_5978), .Y (n_11255));
NAND2X1 g66549(.A (n_9281), .B (n_4582), .Y (n_9409));
NOR2X1 g66558(.A (n_9406), .B (n_9368), .Y (n_9407));
NOR2X1 g66559(.A (n_14523), .B (n_1424), .Y (n_9405));
NAND2X1 g66574(.A (n_9404), .B (n_11576), .Y (n_15511));
OR2X1 g66575(.A (n_8708), .B (n_7373), .Y (n_13298));
NOR2X1 g66579(.A (n_9402), .B (n_10389), .Y (n_9403));
NOR2X1 g66585(.A (n_13804), .B (n_7430), .Y (n_11250));
NAND2X1 g66599(.A (n_18347), .B (n_16480), .Y (n_9399));
NAND2X1 g66604(.A (n_17467), .B (n_17377), .Y (n_9397));
NAND2X1 g66608(.A (n_7592), .B (n_6877), .Y (n_17124));
NOR2X1 g66609(.A (n_5724), .B (n_15688), .Y (n_9395));
NOR2X1 g66610(.A (n_15245), .B (n_16466), .Y (n_9394));
NAND4X1 g66612(.A (n_29065), .B (n_9442), .C (n_9392), .D (n_3702),.Y (n_18958));
NOR2X1 g66621(.A (n_7188), .B (n_15610), .Y (n_9390));
NAND2X2 g66642(.A (n_7444), .B (n_4173), .Y (n_11562));
NAND2X1 g66665(.A (n_9389), .B (n_9388), .Y (n_11549));
NAND2X1 g66666(.A (n_9344), .B (n_14142), .Y (n_9387));
NOR2X1 g70020(.A (n_9246), .B (n_7419), .Y (n_9386));
NAND2X1 g77704(.A (n_3301), .B (n_23418), .Y (n_9385));
NOR2X1 g66693(.A (n_7068), .B (n_7201), .Y (n_9384));
NAND4X1 g66709(.A (n_9500), .B (n_11835), .C (n_2124), .D (n_6445),.Y (n_15236));
NAND2X1 g66712(.A (n_17491), .B (n_16787), .Y (n_9382));
NOR2X1 g66733(.A (n_9380), .B (n_15388), .Y (n_11211));
NOR2X1 g66765(.A (n_7395), .B (n_12827), .Y (n_11203));
NOR2X1 g66782(.A (n_6942), .B (n_12559), .Y (n_9377));
NAND2X1 g67327(.A (n_7333), .B (n_2810), .Y (n_11524));
NOR2X1 g66800(.A (n_9450), .B (n_124), .Y (n_9375));
NOR2X1 g66810(.A (n_27365), .B (n_29363), .Y (n_9374));
NOR2X1 g66827(.A (n_7600), .B (n_11052), .Y (n_11181));
NOR2X1 g73068(.A (n_6716), .B (n_11731), .Y (n_9372));
NAND2X1 g66847(.A (n_9371), .B (n_9370), .Y (n_16868));
NAND2X1 g66856(.A (n_7390), .B (n_9368), .Y (n_9369));
NAND2X1 g66864(.A (n_7343), .B (n_1647), .Y (n_14942));
NAND2X1 g66877(.A (n_26491), .B (n_7283), .Y (n_28877));
INVX1 g66885(.A (n_9366), .Y (n_11528));
NAND2X1 g66899(.A (n_9363), .B (n_3193), .Y (n_9364));
NAND2X1 g66901(.A (n_4555), .B (n_6993), .Y (n_9362));
NAND2X1 g71350(.A (n_8308), .B (n_12169), .Y (n_9361));
NAND4X1 g66913(.A (n_12335), .B (n_4261), .C (n_28472), .D (n_3559),.Y (n_17262));
NAND2X1 g66917(.A (n_7307), .B (n_9357), .Y (n_11539));
NAND2X1 g66923(.A (n_9355), .B (n_7598), .Y (n_9356));
INVX1 g66926(.A (n_9354), .Y (n_13148));
INVX1 g66944(.A (n_7629), .Y (n_13282));
NAND2X1 g66947(.A (n_9353), .B (n_10495), .Y (n_13567));
NAND2X2 g66966(.A (n_6915), .B (n_11323), .Y (n_11154));
AND2X1 g66968(.A (n_9529), .B (n_17619), .Y (n_11151));
NAND2X1 g66970(.A (n_9351), .B (n_9370), .Y (n_9352));
OR2X1 g66972(.A (n_9350), .B (n_12827), .Y (n_14922));
NAND2X1 g66977(.A (n_9349), .B (n_10599), .Y (n_15260));
OR2X1 g67007(.A (n_9348), .B (n_13083), .Y (n_11139));
NOR2X1 g71348(.A (n_27365), .B (n_3918), .Y (n_10071));
OR2X1 g67013(.A (n_6723), .B (n_11307), .Y (n_19216));
INVX1 g67036(.A (n_9346), .Y (n_13351));
NOR2X1 g67281(.A (n_6005), .B (n_9345), .Y (n_13272));
NAND2X1 g67042(.A (n_15507), .B (n_9344), .Y (n_20013));
OR2X1 g67043(.A (n_7847), .B (n_12827), .Y (n_11558));
NAND2X1 g67050(.A (n_16934), .B (n_9389), .Y (n_11124));
NAND2X1 g67059(.A (n_8911), .B (n_10868), .Y (n_9343));
AND2X1 g67067(.A (n_6811), .B (n_9342), .Y (n_13476));
NAND2X1 g67082(.A (n_7703), .B (n_29256), .Y (n_14978));
OR2X1 g67087(.A (n_9340), .B (n_11307), .Y (n_9341));
NAND2X1 g71337(.A (n_5507), .B (n_5677), .Y (n_9338));
NAND2X1 g67099(.A (n_7481), .B (n_4861), .Y (n_14927));
NAND2X1 g67262(.A (n_2457), .B (n_6884), .Y (n_9337));
NAND2X2 g72313(.A (n_9336), .B (n_9335), .Y (n_11102));
NAND2X1 g67127(.A (n_9333), .B (n_8968), .Y (n_9334));
NOR2X1 g67135(.A (n_9363), .B (n_8637), .Y (n_11096));
AND2X1 g67137(.A (n_9332), .B (n_15245), .Y (n_11094));
NOR2X1 g67156(.A (n_7566), .B (n_7201), .Y (n_11091));
NAND2X1 g67164(.A (n_9330), .B (n_9217), .Y (n_9331));
NAND2X1 g67175(.A (n_9345), .B (n_2733), .Y (n_9329));
OR2X1 g67181(.A (n_9328), .B (n_9527), .Y (n_11086));
NAND2X1 g67190(.A (n_12246), .B (n_9326), .Y (n_9327));
NAND2X1 g67192(.A (n_27710), .B (n_11422), .Y (n_13340));
NAND2X1 g67201(.A (n_6107), .B (n_5851), .Y (n_9325));
NOR2X1 g67203(.A (n_12298), .B (n_5700), .Y (n_13307));
NAND2X1 g67224(.A (n_7494), .B (n_9057), .Y (n_9323));
NAND2X1 g67228(.A (n_9322), .B (n_16976), .Y (n_13752));
INVX1 g73028(.A (n_6873), .Y (n_9321));
NAND2X1 g67252(.A (n_4343), .B (n_9319), .Y (n_9320));
INVX1 g73583(.A (n_9962), .Y (n_11812));
INVX1 g67270(.A (n_7690), .Y (n_9318));
NOR2X1 g67290(.A (n_9211), .B (n_7182), .Y (n_9317));
NOR2X1 g67291(.A (n_9315), .B (n_9314), .Y (n_9316));
NOR2X1 g67299(.A (n_6971), .B (n_14866), .Y (n_11057));
INVX1 g67317(.A (n_7671), .Y (n_9313));
NAND2X1 g67338(.A (n_3122), .B (n_9283), .Y (n_9312));
NAND2X1 g67351(.A (n_7241), .B (n_7496), .Y (n_11045));
INVX1 g73584(.A (n_9962), .Y (n_9311));
OR2X1 g67370(.A (n_9309), .B (n_7410), .Y (n_9310));
NAND2X1 g67382(.A (n_8039), .B (n_7035), .Y (n_9308));
AOI21X1 g67383(.A0 (n_4286), .A1 (n_3334), .B0 (n_4582), .Y (n_9307));
NAND2X1 g67384(.A (n_7894), .B (n_13269), .Y (n_9306));
OR2X1 g67388(.A (n_9303), .B (n_5817), .Y (n_9304));
NAND2X1 g67390(.A (n_4185), .B (n_6950), .Y (n_9301));
NAND2X1 g67406(.A (n_27372), .B (n_3214), .Y (n_9300));
INVX1 g72288(.A (n_9299), .Y (n_12484));
OR2X1 g67409(.A (n_7603), .B (n_16466), .Y (n_11034));
AND2X1 g67430(.A (n_7161), .B (n_12827), .Y (n_11024));
INVX1 g73003(.A (n_15534), .Y (n_9764));
INVX4 g69930(.A (n_8937), .Y (n_12495));
NAND2X1 g72286(.A (n_8441), .B (n_28734), .Y (n_9298));
NAND2X1 g67478(.A (n_4145), .B (n_7708), .Y (n_9297));
NAND3X1 g67492(.A (n_9295), .B (n_9294), .C (n_9293), .Y (n_9296));
NAND2X1 g67500(.A (n_7976), .B (n_8217), .Y (n_11011));
NAND2X1 g67508(.A (n_7572), .B (n_9783), .Y (n_13370));
NAND2X1 g67511(.A (n_9291), .B (n_2810), .Y (n_17757));
NAND2X2 g67514(.A (n_27643), .B (n_28418), .Y (n_15012));
NAND2X1 g67517(.A (n_8070), .B (n_7124), .Y (n_9290));
NAND2X1 g71305(.A (n_5126), .B (n_8520), .Y (n_9289));
NAND2X1 g67606(.A (n_28993), .B (n_6005), .Y (n_9288));
NOR2X1 g67637(.A (n_7416), .B (n_4898), .Y (n_10982));
NOR2X1 g67658(.A (n_12896), .B (n_9285), .Y (n_13303));
NOR2X1 g67661(.A (n_9999), .B (n_9283), .Y (n_9284));
NAND2X1 g67662(.A (n_5312), .B (n_7879), .Y (n_9282));
NAND2X1 g67666(.A (n_9281), .B (n_12134), .Y (n_18385));
NAND2X1 g67675(.A (n_7422), .B (n_12979), .Y (n_13322));
NAND2X1 g67676(.A (n_7081), .B (n_2260), .Y (n_15009));
INVX1 g67681(.A (n_9279), .Y (n_13186));
INVX1 g67684(.A (n_16963), .Y (n_9278));
NAND4X1 g67701(.A (n_9276), .B (n_3807), .C (n_3464), .D (n_3925), .Y(n_15100));
AOI21X1 g67706(.A0 (n_7615), .A1 (n_3253), .B0 (n_15776), .Y(n_9274));
INVX1 g67712(.A (n_7843), .Y (n_13333));
NAND2X1 g67716(.A (n_14037), .B (n_9272), .Y (n_9273));
NAND2X1 g67123(.A (n_27671), .B (n_6005), .Y (n_15019));
NAND2X1 g67729(.A (n_7450), .B (n_6185), .Y (n_15028));
NAND2X1 g67733(.A (n_4390), .B (n_7082), .Y (n_9269));
NOR2X1 g72263(.A (n_3571), .B (n_5854), .Y (n_9268));
INVX1 g67740(.A (n_7656), .Y (n_13159));
OR2X1 g67744(.A (n_14208), .B (n_29102), .Y (n_25468));
INVX1 g67758(.A (n_18598), .Y (n_10961));
NOR2X1 g69892(.A (n_6597), .B (n_9264), .Y (n_9265));
NAND2X2 g67784(.A (n_7585), .B (n_11731), .Y (n_11470));
NOR2X1 g72260(.A (n_6532), .B (n_26276), .Y (n_9262));
NAND2X1 g67817(.A (n_9260), .B (n_13318), .Y (n_9261));
NAND2X2 g67844(.A (n_7547), .B (n_8637), .Y (n_17821));
NAND2X1 g67847(.A (n_5772), .B (n_8679), .Y (n_10934));
INVX1 g67876(.A (n_7653), .Y (n_13357));
NAND2X1 g67882(.A (n_9258), .B (n_9257), .Y (n_10923));
NOR2X1 g67902(.A (n_13804), .B (n_5742), .Y (n_10917));
NAND2X1 g67905(.A (n_9016), .B (n_6937), .Y (n_9255));
NAND2X1 g67941(.A (n_8863), .B (n_7036), .Y (n_9254));
AOI21X1 g67943(.A0 (n_11924), .A1 (n_3085), .B0 (n_8141), .Y(n_9253));
NAND2X1 g72245(.A (n_2043), .B (n_4757), .Y (n_9894));
NAND2X1 g67978(.A (n_7532), .B (n_352), .Y (n_28809));
NAND2X1 g67979(.A (n_8809), .B (n_6900), .Y (n_9251));
OAI21X1 g61897(.A0 (n_4421), .A1 (n_10999), .B0 (n_9249), .Y(n_9250));
NOR2X1 g68004(.A (n_7079), .B (n_13490), .Y (n_10893));
NAND2X1 g68007(.A (n_9246), .B (n_7160), .Y (n_9247));
NAND2X1 g68008(.A (n_8954), .B (n_7719), .Y (n_9245));
INVX1 g72242(.A (n_7011), .Y (n_10882));
INVX1 g68020(.A (n_13324), .Y (n_10885));
AOI21X1 g68024(.A0 (n_12494), .A1 (n_2295), .B0 (n_8346), .Y(n_9244));
INVX1 g68027(.A (n_9242), .Y (n_9243));
NAND2X1 g68042(.A (n_12172), .B (n_8780), .Y (n_9241));
INVX1 g68045(.A (n_7645), .Y (n_10878));
NAND2X2 g68054(.A (n_7521), .B (n_4861), .Y (n_14765));
NAND2X1 g68106(.A (n_8904), .B (n_7226), .Y (n_9238));
INVX1 g69850(.A (n_7437), .Y (n_10862));
OR2X1 g72795(.A (n_9236), .B (n_12917), .Y (n_9237));
NAND2X1 g68150(.A (n_9234), .B (n_3366), .Y (n_9235));
NOR2X1 g68156(.A (n_9232), .B (n_16978), .Y (n_9233));
NAND2X2 g72232(.A (n_28614), .B (n_6092), .Y (n_16070));
INVX1 g71260(.A (n_10832), .Y (n_9230));
NAND3X1 g68175(.A (n_8662), .B (n_7770), .C (n_3931), .Y (n_9229));
NOR2X1 g69834(.A (n_12019), .B (n_7844), .Y (n_10437));
AOI21X1 g61954(.A0 (n_6301), .A1 (dcnt[3] ), .B0 (n_6302), .Y(n_9228));
INVX1 g69840(.A (n_9227), .Y (n_12322));
AND2X1 g68191(.A (n_9332), .B (n_10836), .Y (n_9226));
NAND2X1 g68466(.A (n_4283), .B (n_9309), .Y (n_9225));
NAND2X1 g68246(.A (n_7815), .B (n_4173), .Y (n_16568));
INVX1 g72920(.A (n_10948), .Y (n_9781));
NAND3X1 g68254(.A (n_9221), .B (n_7686), .C (n_9220), .Y (n_9222));
NOR2X1 g68260(.A (n_28993), .B (n_7388), .Y (n_9219));
OR2X1 g66997(.A (n_9217), .B (n_11385), .Y (n_13504));
NAND2X1 g68278(.A (n_6018), .B (n_12187), .Y (n_9215));
NOR2X1 g68293(.A (n_9212), .B (n_1667), .Y (n_9213));
OR2X1 g68295(.A (n_9211), .B (n_9527), .Y (n_10825));
INVX1 g68310(.A (n_7389), .Y (n_10824));
NAND3X1 g68313(.A (n_3982), .B (n_7215), .C (n_7415), .Y (n_9210));
INVX1 g69813(.A (n_10909), .Y (n_10444));
OR2X1 g68370(.A (n_9209), .B (n_18369), .Y (n_10805));
NOR2X1 g68373(.A (n_9564), .B (n_11276), .Y (n_13359));
NOR2X1 g69810(.A (n_7641), .B (n_29221), .Y (n_10445));
INVX1 g69800(.A (n_9208), .Y (n_13076));
NAND2X1 g68432(.A (n_26550), .B (n_28423), .Y (n_9207));
NAND2X1 g68457(.A (n_4328), .B (n_9340), .Y (n_9205));
XOR2X1 g76296(.A (n_9203), .B (n_9202), .Y (n_9204));
NAND2X1 g68516(.A (n_5201), .B (n_9200), .Y (n_9201));
INVX1 g72895(.A (n_7623), .Y (n_14094));
NAND2X1 g68534(.A (n_5181), .B (n_5776), .Y (n_9199));
NOR2X1 g68535(.A (n_5397), .B (n_5813), .Y (n_9198));
NOR2X1 g72894(.A (n_3289), .B (n_8997), .Y (n_12664));
INVX1 g69782(.A (n_8959), .Y (n_12340));
OR2X1 g72893(.A (n_1811), .B (n_25926), .Y (n_9197));
OAI21X1 g68554(.A0 (n_9195), .A1 (n_5151), .B0 (n_9193), .Y (n_9196));
NAND2X1 g68558(.A (n_4257), .B (n_9303), .Y (n_9192));
NAND2X1 g68569(.A (n_5380), .B (n_9190), .Y (n_9191));
AOI21X1 g68592(.A0 (n_2444), .A1 (n_3372), .B0 (n_2291), .Y (n_9189));
AOI21X1 g68613(.A0 (n_4130), .A1 (n_11323), .B0 (n_5893), .Y(n_9188));
NAND2X1 g68614(.A (n_6046), .B (n_9234), .Y (n_9187));
AOI21X1 g68619(.A0 (n_4071), .A1 (n_1647), .B0 (n_5789), .Y (n_9186));
NAND2X1 g68639(.A (n_5939), .B (n_9183), .Y (n_9184));
NAND2X1 g72190(.A (n_2527), .B (n_7367), .Y (n_9906));
INVX1 g72078(.A (n_9181), .Y (n_9182));
NOR2X1 g68666(.A (n_5949), .B (n_7104), .Y (n_9180));
INVX1 g71209(.A (n_11003), .Y (n_9179));
NAND2X1 g68395(.A (n_3305), .B (n_11322), .Y (n_10801));
AOI21X1 g68700(.A0 (n_4388), .A1 (n_7477), .B0 (n_4382), .Y (n_9175));
OAI21X1 g68712(.A0 (n_3247), .A1 (n_7583), .B0 (n_7932), .Y (n_9174));
AND2X1 g68714(.A (n_5837), .B (n_19226), .Y (n_9173));
INVX1 g72864(.A (n_12177), .Y (n_9172));
AOI21X1 g68726(.A0 (n_9170), .A1 (n_3654), .B0 (n_17467), .Y(n_9171));
NAND2X1 g68735(.A (n_5180), .B (n_7795), .Y (n_9169));
OAI21X1 g68756(.A0 (n_6609), .A1 (n_473), .B0 (n_19019), .Y (n_9166));
OAI21X1 g68772(.A0 (n_3640), .A1 (n_2934), .B0 (n_13536), .Y(n_9165));
OAI21X1 g68776(.A0 (n_9163), .A1 (n_7678), .B0 (n_6871), .Y (n_9164));
AND2X1 g68790(.A (n_5458), .B (n_5917), .Y (n_9162));
AND2X1 g68794(.A (n_5187), .B (n_4558), .Y (n_9161));
MX2X1 g68796(.A (n_7685), .B (n_3119), .S0 (n_7777), .Y (n_9160));
NOR2X1 g68798(.A (n_5134), .B (n_4787), .Y (n_9159));
AND2X1 g68806(.A (n_4356), .B (n_5886), .Y (n_9158));
INVX1 g68811(.A (n_9156), .Y (n_9157));
XOR2X1 g68822(.A (n_1087), .B (n_4111), .Y (n_9155));
OR2X1 g71186(.A (n_8603), .B (n_12169), .Y (n_12786));
NAND2X1 g72848(.A (n_2418), .B (n_8520), .Y (n_9152));
INVX1 g69730(.A (n_7457), .Y (n_10463));
NOR2X1 g72842(.A (n_3858), .B (n_15894), .Y (n_9149));
INVX1 g68971(.A (n_11165), .Y (n_12835));
INVX1 g68974(.A (n_9145), .Y (n_9146));
INVX1 g68985(.A (n_9143), .Y (n_12613));
INVX1 g68993(.A (n_9142), .Y (n_10644));
INVX1 g68996(.A (n_9140), .Y (n_14286));
NOR2X1 g72134(.A (n_3699), .B (n_29244), .Y (n_9913));
NOR2X1 g69000(.A (n_9139), .B (n_12469), .Y (n_10640));
NOR2X1 g69003(.A (n_5626), .B (n_26491), .Y (n_10637));
NAND2X1 g69004(.A (n_6420), .B (n_29269), .Y (n_9138));
OR2X1 g69008(.A (n_8380), .B (n_8090), .Y (n_13690));
OR2X1 g69011(.A (n_9018), .B (n_9783), .Y (n_9136));
NOR2X1 g69013(.A (n_5545), .B (n_29244), .Y (n_10633));
OR2X1 g69015(.A (n_5788), .B (n_9050), .Y (n_9135));
OR2X1 g69016(.A (n_5322), .B (n_11312), .Y (n_18199));
INVX1 g69017(.A (n_13607), .Y (n_9134));
INVX1 g69020(.A (n_13607), .Y (n_18982));
INVX1 g69029(.A (n_7596), .Y (n_12362));
NAND2X1 g69032(.A (n_27076), .B (n_17260), .Y (n_13561));
INVX1 g69033(.A (n_9132), .Y (n_15002));
INVX1 g69034(.A (n_9132), .Y (n_9133));
INVX1 g69047(.A (n_9129), .Y (n_9130));
INVX1 g69061(.A (n_9127), .Y (n_9126));
INVX1 g69063(.A (n_9124), .Y (n_9125));
CLKBUFX3 g69065(.A (n_9124), .Y (n_12779));
AND2X1 g69067(.A (n_9046), .B (n_15894), .Y (n_9123));
INVX2 g69069(.A (n_10968), .Y (n_18264));
NOR2X1 g69079(.A (n_4486), .B (n_9118), .Y (n_10621));
NAND2X1 g72834(.A (n_2074), .B (n_13768), .Y (n_25616));
INVX1 g69088(.A (n_9116), .Y (n_12266));
INVX1 g69096(.A (n_9115), .Y (n_10618));
INVX1 g69099(.A (n_9114), .Y (n_14080));
INVX1 g69102(.A (n_13217), .Y (n_9113));
INVX1 g69104(.A (n_9111), .Y (n_9112));
INVX1 g69120(.A (n_9108), .Y (n_10613));
NAND2X2 g69137(.A (n_6748), .B (n_9691), .Y (n_10609));
AND2X1 g69140(.A (n_8889), .B (n_9106), .Y (n_9107));
INVX1 g69141(.A (n_6416), .Y (n_16049));
INVX1 g69145(.A (n_14521), .Y (n_12928));
NAND2X1 g69150(.A (n_8664), .B (n_12910), .Y (n_12251));
AND2X1 g69151(.A (n_6679), .B (n_9084), .Y (n_9105));
INVX1 g69153(.A (n_14014), .Y (n_10605));
INVX1 g69155(.A (n_10701), .Y (n_12480));
INVX1 g69160(.A (n_11029), .Y (n_10604));
INVX1 g69167(.A (n_7574), .Y (n_10603));
INVX1 g69187(.A (n_6463), .Y (n_10598));
NAND2X1 g69189(.A (n_6919), .B (n_9368), .Y (n_9103));
NOR2X1 g69194(.A (n_8254), .B (n_27365), .Y (n_10595));
INVX1 g69203(.A (n_7565), .Y (n_9635));
INVX1 g69208(.A (n_7564), .Y (n_12518));
NAND2X2 g69210(.A (n_6417), .B (n_14484), .Y (n_12354));
OR2X1 g69211(.A (n_11104), .B (n_14866), .Y (n_15285));
INVX1 g69213(.A (n_6542), .Y (n_17011));
NOR2X1 g69221(.A (n_11322), .B (n_6614), .Y (n_10590));
NAND2X2 g69224(.A (n_9098), .B (n_8997), .Y (n_10589));
OR2X1 g69225(.A (n_4412), .B (n_7325), .Y (n_12632));
INVX1 g69226(.A (n_9095), .Y (n_9096));
NOR2X1 g69230(.A (n_6614), .B (n_15708), .Y (n_9094));
INVX1 g69242(.A (n_17130), .Y (n_9092));
NAND2X1 g69246(.A (n_5496), .B (n_26491), .Y (n_9091));
NOR2X1 g69248(.A (n_5953), .B (n_9783), .Y (n_10585));
NAND4X1 g69249(.A (n_20325), .B (n_9089), .C (n_8918), .D (n_2910),.Y (n_12234));
INVX1 g69250(.A (n_9088), .Y (n_12801));
NAND2X1 g69255(.A (n_6728), .B (n_12019), .Y (n_12597));
INVX1 g69258(.A (n_11334), .Y (n_12762));
NOR2X1 g69268(.A (n_6475), .B (n_9084), .Y (n_10581));
NAND2X1 g69272(.A (n_5233), .B (n_11323), .Y (n_13257));
NAND2X1 g69281(.A (n_5358), .B (n_29256), .Y (n_9082));
NAND2X1 g69282(.A (n_6269), .B (n_14142), .Y (n_9081));
NAND2X1 g69291(.A (n_9078), .B (n_9388), .Y (n_9079));
INVX1 g69295(.A (n_10971), .Y (n_10575));
NAND2X1 g69299(.A (n_9077), .B (n_29221), .Y (n_13260));
OR2X1 g72821(.A (n_9073), .B (n_12850), .Y (n_9074));
INVX2 g69319(.A (n_7544), .Y (n_12591));
NAND2X1 g69329(.A (n_4178), .B (n_5912), .Y (n_9069));
INVX1 g69333(.A (n_11381), .Y (n_10566));
INVX1 g69342(.A (n_11516), .Y (n_9068));
INVX1 g69344(.A (n_9066), .Y (n_17621));
INVX1 g69366(.A (n_9060), .Y (n_9061));
NAND2X1 g69372(.A (n_9058), .B (n_9057), .Y (n_10561));
INVX1 g72817(.A (n_7527), .Y (n_17012));
INVX2 g69390(.A (n_7522), .Y (n_12409));
NOR2X1 g69408(.A (n_9053), .B (n_13804), .Y (n_9054));
NAND2X1 g69411(.A (n_6711), .B (n_2318), .Y (n_10549));
NAND2X1 g69418(.A (n_9050), .B (n_13593), .Y (n_9051));
INVX1 g69420(.A (n_9048), .Y (n_10548));
NAND2X1 g69423(.A (n_9046), .B (n_6534), .Y (n_9047));
INVX1 g69424(.A (n_11133), .Y (n_9045));
INVX1 g69426(.A (n_7518), .Y (n_18920));
OR2X1 g69434(.A (n_8355), .B (n_6420), .Y (n_9044));
INVX1 g69435(.A (n_9043), .Y (n_21122));
NOR2X1 g69449(.A (n_6491), .B (n_8974), .Y (n_10542));
INVX1 g69452(.A (n_9040), .Y (n_10539));
NOR2X1 g69460(.A (n_5243), .B (n_28692), .Y (n_9039));
NOR2X1 g69463(.A (n_9037), .B (n_8865), .Y (n_9038));
CLKBUFX3 g69481(.A (n_9033), .Y (n_14803));
NAND2X1 g69484(.A (n_8855), .B (n_7498), .Y (n_9032));
INVX1 g69504(.A (n_11235), .Y (n_10524));
INVX1 g69507(.A (n_11473), .Y (n_9029));
INVX1 g69509(.A (n_9026), .Y (n_9028));
INVX1 g69513(.A (n_14510), .Y (n_13063));
INVX1 g69516(.A (n_11263), .Y (n_9024));
AND2X1 g69519(.A (n_6764), .B (n_6008), .Y (n_14201));
NAND2X1 g69524(.A (n_5714), .B (n_27309), .Y (n_9023));
OR2X1 g69526(.A (n_8916), .B (n_28686), .Y (n_16359));
NOR2X1 g69529(.A (n_9020), .B (n_8997), .Y (n_9021));
OR2X1 g69532(.A (n_9018), .B (n_27688), .Y (n_14800));
INVX1 g69533(.A (n_10784), .Y (n_20078));
NOR2X1 g69538(.A (n_9016), .B (n_7607), .Y (n_9017));
NOR2X1 g69540(.A (n_4444), .B (n_29256), .Y (n_10522));
NAND2X1 g69543(.A (n_6106), .B (n_7201), .Y (n_9015));
NOR2X1 g69545(.A (n_5629), .B (n_11300), .Y (n_10521));
INVX1 g69546(.A (n_7494), .Y (n_18046));
NAND2X1 g69554(.A (n_4703), .B (n_10495), .Y (n_10519));
NAND2X1 g69558(.A (n_8894), .B (n_7201), .Y (n_9013));
OR2X1 g69570(.A (n_5153), .B (n_7418), .Y (n_9008));
INVX1 g71124(.A (n_9006), .Y (n_10122));
NAND2X1 g69574(.A (n_5253), .B (n_3318), .Y (n_9005));
NOR2X1 g69586(.A (n_5243), .B (n_11272), .Y (n_10509));
OR2X1 g69590(.A (n_9004), .B (n_9003), .Y (n_10506));
NAND2X1 g69591(.A (n_5728), .B (n_7023), .Y (n_25626));
INVX1 g69596(.A (n_10964), .Y (n_14319));
INVX4 g69606(.A (n_9000), .Y (n_13609));
OR2X1 g69609(.A (n_8611), .B (n_12469), .Y (n_16970));
NOR2X1 g69612(.A (n_6670), .B (n_29256), .Y (n_10501));
NOR2X1 g69621(.A (n_5221), .B (n_8997), .Y (n_10492));
INVX1 g69624(.A (n_11080), .Y (n_8996));
OR2X1 g69628(.A (n_5440), .B (n_14866), .Y (n_17321));
INVX1 g69638(.A (n_7368), .Y (n_10489));
OR2X1 g69644(.A (n_3999), .B (n_14866), .Y (n_10485));
OR2X1 g69647(.A (n_6200), .B (n_14484), .Y (n_10483));
NOR2X1 g69649(.A (n_4881), .B (n_13593), .Y (n_10480));
NOR2X1 g69657(.A (n_6384), .B (n_18266), .Y (n_10476));
NAND2X1 g69661(.A (n_7294), .B (n_383), .Y (n_10475));
NOR2X1 g69664(.A (n_3991), .B (n_28037), .Y (n_10472));
OR2X1 g69665(.A (n_8931), .B (n_17260), .Y (n_14841));
INVX1 g69674(.A (n_10838), .Y (n_8990));
INVX1 g69671(.A (n_7469), .Y (n_10471));
OR2X1 g69692(.A (n_8687), .B (n_26880), .Y (n_15487));
AND2X1 g69693(.A (n_6703), .B (n_11322), .Y (n_8986));
INVX1 g69695(.A (n_8983), .Y (n_8984));
NOR2X1 g69699(.A (n_6851), .B (n_7598), .Y (n_10466));
INVX1 g69710(.A (n_7550), .Y (n_16999));
AOI21X1 g69713(.A0 (n_4901), .A1 (n_2109), .B0 (n_5735), .Y (n_8980));
OR2X1 g69714(.A (n_8978), .B (n_7598), .Y (n_8979));
NAND2X1 g69715(.A (n_5309), .B (n_6534), .Y (n_8977));
INVX1 g69718(.A (n_11043), .Y (n_20786));
NAND2X1 g69720(.A (n_5341), .B (n_28427), .Y (n_8976));
AND2X1 g69721(.A (n_6758), .B (n_8974), .Y (n_28583));
INVX1 g69736(.A (n_10835), .Y (n_12570));
NAND2X1 g69738(.A (n_5510), .B (n_13490), .Y (n_8973));
OR2X1 g69743(.A (n_8971), .B (n_1424), .Y (n_8972));
INVX1 g69745(.A (n_8970), .Y (n_12740));
NAND2X1 g69747(.A (n_6794), .B (n_7598), .Y (n_8969));
NOR2X1 g69749(.A (n_26488), .B (n_8968), .Y (n_12715));
INVX1 g69752(.A (n_16416), .Y (n_10460));
XOR2X1 g76243(.A (text_in_r[9] ), .B (n_933), .Y (n_8966));
NAND2X1 g69757(.A (n_7367), .B (n_14055), .Y (n_29000));
NAND2X1 g69768(.A (n_7800), .B (n_8974), .Y (n_10454));
NAND2X1 g69769(.A (n_8778), .B (n_13815), .Y (n_8963));
INVX1 g69771(.A (n_10915), .Y (n_8962));
NOR2X1 g69775(.A (n_4203), .B (n_9474), .Y (n_10451));
NAND2X1 g72074(.A (n_6304), .B (n_4689), .Y (n_12416));
NAND2X1 g69788(.A (n_5296), .B (n_14055), .Y (n_8958));
NAND2X1 g69794(.A (n_6606), .B (n_11307), .Y (n_8956));
NOR2X1 g69797(.A (n_8954), .B (n_26880), .Y (n_10448));
INVX1 g69805(.A (n_10799), .Y (n_10447));
OR2X1 g72070(.A (n_8951), .B (n_6847), .Y (n_8952));
INVX2 g69823(.A (n_11020), .Y (n_12907));
INVX1 g69829(.A (n_10956), .Y (n_18882));
NAND2X2 g69836(.A (n_8367), .B (n_7496), .Y (n_12299));
NOR2X1 g69844(.A (n_4950), .B (n_8974), .Y (n_10432));
INVX1 g69846(.A (n_14407), .Y (n_10431));
NOR2X1 g69856(.A (n_5474), .B (n_8974), .Y (n_8948));
INVX1 g69859(.A (n_13162), .Y (n_10429));
NAND2X1 g69867(.A (n_8810), .B (n_8945), .Y (n_8946));
INVX1 g69873(.A (n_8943), .Y (n_13965));
OR2X1 g69877(.A (n_29192), .B (n_17414), .Y (n_8942));
INVX1 g69887(.A (n_8941), .Y (n_10424));
NOR2X1 g69899(.A (n_8834), .B (n_20325), .Y (n_8940));
INVX1 g69900(.A (n_8939), .Y (n_12713));
NAND2X2 g69915(.A (n_7052), .B (n_28757), .Y (n_12885));
NOR2X1 g69934(.A (n_28035), .B (n_6005), .Y (n_12496));
INVX1 g69935(.A (n_14340), .Y (n_8936));
NOR2X1 g69941(.A (n_7331), .B (n_5591), .Y (n_10415));
NOR2X1 g69945(.A (n_8935), .B (n_9416), .Y (n_10414));
INVX1 g69947(.A (n_11200), .Y (n_10413));
INVX1 g69954(.A (n_10945), .Y (n_10411));
NOR2X1 g69959(.A (n_4636), .B (n_14484), .Y (n_10408));
INVX1 g69960(.A (n_11530), .Y (n_8934));
CLKBUFX1 g69961(.A (n_11530), .Y (n_14858));
NAND2X1 g69963(.A (n_5166), .B (n_13247), .Y (n_8933));
OR2X1 g69965(.A (n_8931), .B (n_29256), .Y (n_8932));
OR2X1 g69973(.A (n_9804), .B (n_28134), .Y (n_13686));
CLKBUFX1 g69974(.A (n_8929), .Y (n_16801));
NOR2X1 g69978(.A (n_5575), .B (n_6005), .Y (n_10401));
NOR2X1 g69982(.A (n_4435), .B (n_8928), .Y (n_10397));
NOR2X1 g69985(.A (n_5589), .B (n_13490), .Y (n_12555));
NOR2X1 g69988(.A (n_9668), .B (n_8560), .Y (n_8927));
INVX1 g69989(.A (n_8924), .Y (n_8925));
INVX1 g69652(.A (n_8922), .Y (n_10478));
NOR2X1 g69995(.A (n_7837), .B (n_28375), .Y (n_8921));
NAND4X1 g70001(.A (n_2910), .B (n_9089), .C (n_8918), .D (n_10031),.Y (n_15105));
OR2X1 g70021(.A (n_8916), .B (n_12019), .Y (n_8917));
XOR2X1 g76108(.A (n_1019), .B (n_3888), .Y (n_8915));
NAND2X1 g70025(.A (n_6228), .B (n_14484), .Y (n_8914));
NAND2X1 g70026(.A (n_5146), .B (n_2260), .Y (n_8913));
NAND2X1 g70036(.A (n_7397), .B (n_9118), .Y (n_12359));
INVX1 g70040(.A (n_10921), .Y (n_10391));
NOR2X1 g70045(.A (n_8911), .B (n_8910), .Y (n_8912));
NAND2X1 g70048(.A (n_5529), .B (n_10389), .Y (n_8909));
INVX1 g70051(.A (n_8908), .Y (n_10387));
INVX1 g70061(.A (n_8907), .Y (n_10384));
OR2X1 g70066(.A (n_5586), .B (n_11322), .Y (n_10382));
NAND2X1 g70067(.A (n_5462), .B (n_16466), .Y (n_8905));
NOR2X1 g70073(.A (n_6611), .B (n_8452), .Y (n_10380));
INVX1 g72779(.A (n_8902), .Y (n_8903));
INVX1 g70077(.A (n_7748), .Y (n_12175));
INVX1 g70079(.A (n_10900), .Y (n_8901));
AND2X1 g70083(.A (n_8396), .B (n_12019), .Y (n_8900));
INVX1 g70089(.A (n_10957), .Y (n_10374));
NAND2X1 g70118(.A (n_4741), .B (n_6005), .Y (n_10366));
INVX1 g70122(.A (n_8897), .Y (n_15961));
INVX1 g70126(.A (n_8897), .Y (n_8896));
NAND2X1 g70130(.A (n_8894), .B (n_11489), .Y (n_8895));
NOR2X1 g70133(.A (n_4950), .B (n_28680), .Y (n_10362));
INVX1 g70141(.A (n_8892), .Y (n_10357));
OR2X1 g70143(.A (n_8296), .B (n_3834), .Y (n_13684));
OR2X1 g70144(.A (n_9552), .B (n_4113), .Y (n_15493));
OR2X1 g70152(.A (n_4727), .B (n_12169), .Y (n_12752));
NAND2X1 g70155(.A (n_5544), .B (n_9264), .Y (n_8891));
NAND2X1 g70159(.A (n_8889), .B (n_14484), .Y (n_8890));
NOR2X1 g70165(.A (n_10452), .B (n_7746), .Y (n_12420));
NOR2X1 g70167(.A (n_6384), .B (n_4709), .Y (n_8888));
INVX1 g70169(.A (n_8887), .Y (n_15705));
INVX1 g70178(.A (n_11287), .Y (n_10351));
INVX1 g72042(.A (n_8884), .Y (n_8885));
NAND2X1 g70184(.A (n_5015), .B (n_9982), .Y (n_12209));
OR2X1 g70186(.A (n_28610), .B (n_9368), .Y (n_14390));
INVX1 g70193(.A (n_10986), .Y (n_8881));
INVX2 g73368(.A (n_10125), .Y (n_11831));
INVX1 g72769(.A (n_8880), .Y (n_10345));
NOR2X1 g70203(.A (n_28810), .B (n_9257), .Y (n_12410));
NAND2X2 g70205(.A (n_8879), .B (n_10100), .Y (n_12313));
INVX1 g70207(.A (n_11175), .Y (n_18721));
NAND2X1 g70209(.A (n_6306), .B (n_8878), .Y (n_12828));
INVX1 g70210(.A (n_8876), .Y (n_8877));
NAND2X1 g70215(.A (n_5299), .B (n_26877), .Y (n_8875));
INVX1 g70218(.A (n_16590), .Y (n_8874));
INVX1 g70221(.A (n_16590), .Y (n_19008));
NAND2X1 g70225(.A (n_5738), .B (n_16090), .Y (n_8872));
NOR2X1 g70228(.A (n_5668), .B (n_9118), .Y (n_10338));
NAND2X1 g70229(.A (n_5304), .B (n_16754), .Y (n_8871));
OR2X1 g70232(.A (n_6408), .B (n_2318), .Y (n_10336));
NAND2X2 g72758(.A (n_9959), .B (n_4215), .Y (n_9802));
INVX1 g70246(.A (n_7363), .Y (n_10332));
INVX1 g70248(.A (n_8867), .Y (n_8868));
NAND2X1 g70250(.A (n_7235), .B (n_8865), .Y (n_8866));
NAND2X1 g70253(.A (n_8548), .B (n_9257), .Y (n_10328));
NOR2X1 g70261(.A (n_5389), .B (n_10100), .Y (n_10327));
INVX1 g70267(.A (n_8862), .Y (n_10324));
INVX1 g70273(.A (n_7814), .Y (n_10323));
INVX1 g70275(.A (n_10817), .Y (n_8861));
INVX1 g70277(.A (n_8859), .Y (n_8860));
INVX1 g70282(.A (n_11228), .Y (n_10321));
INVX1 g70283(.A (n_11228), .Y (n_8858));
AND2X1 g70290(.A (n_7812), .B (n_1946), .Y (n_10319));
NAND2X1 g70305(.A (n_8855), .B (n_28642), .Y (n_8856));
INVX2 g74100(.A (n_26878), .Y (n_9668));
INVX1 g70309(.A (n_8851), .Y (n_8852));
INVX1 g70317(.A (n_8850), .Y (n_10314));
INVX1 g70320(.A (n_11053), .Y (n_8849));
INVX1 g70322(.A (n_10865), .Y (n_8848));
AND2X1 g70328(.A (n_5150), .B (n_8846), .Y (n_8847));
NAND2X1 g70331(.A (n_6584), .B (n_10389), .Y (n_8845));
OR2X1 g70334(.A (n_12292), .B (n_11835), .Y (n_8844));
NOR2X1 g70337(.A (n_5568), .B (n_9417), .Y (n_10309));
NOR2X1 g70343(.A (n_6337), .B (n_9819), .Y (n_8842));
NOR2X1 g70347(.A (n_28427), .B (n_25665), .Y (n_10307));
INVX1 g70354(.A (n_8839), .Y (n_18749));
INVX1 g70355(.A (n_8839), .Y (n_8840));
OR2X1 g70367(.A (n_8837), .B (n_11998), .Y (n_25487));
NAND2X1 g70370(.A (n_8396), .B (n_28134), .Y (n_14981));
NOR2X1 g70382(.A (n_27669), .B (n_6005), .Y (n_10299));
OR2X1 g70383(.A (n_8834), .B (n_8997), .Y (n_8835));
INVX1 g70388(.A (n_8833), .Y (n_10297));
NAND2X1 g70395(.A (n_6477), .B (n_6008), .Y (n_10295));
NOR2X1 g70405(.A (n_28865), .B (n_14589), .Y (n_8830));
NAND2X1 g70409(.A (n_6132), .B (n_16434), .Y (n_12691));
INVX1 g70410(.A (n_8827), .Y (n_8828));
OR2X1 g70418(.A (n_5685), .B (n_10389), .Y (n_10287));
NAND2X2 g70426(.A (n_7705), .B (n_9500), .Y (n_8824));
INVX1 g70427(.A (n_8822), .Y (n_8823));
INVX1 g70432(.A (n_27900), .Y (n_8821));
NAND2X2 g70435(.A (n_8820), .B (n_8467), .Y (n_12285));
INVX1 g70445(.A (n_10782), .Y (n_10279));
OR2X1 g70474(.A (n_8817), .B (n_8816), .Y (n_17446));
INVX1 g70480(.A (n_8814), .Y (n_8813));
NOR2X1 g70483(.A (n_8811), .B (n_27604), .Y (n_8812));
INVX1 g70489(.A (n_7308), .Y (n_10269));
NAND2X1 g70503(.A (n_8810), .B (n_9084), .Y (n_10266));
NOR2X1 g70515(.A (n_8809), .B (n_383), .Y (n_10264));
INVX1 g70517(.A (n_6399), .Y (n_12893));
OR2X1 g70519(.A (n_4471), .B (n_11307), .Y (n_12626));
NAND2X1 g72019(.A (n_2555), .B (n_8520), .Y (n_8808));
INVX1 g70530(.A (n_8805), .Y (n_8806));
INVX1 g70538(.A (n_7301), .Y (n_14099));
NAND2X1 g70540(.A (n_7820), .B (n_9003), .Y (n_13782));
INVX1 g70547(.A (n_14512), .Y (n_10260));
NOR2X1 g70553(.A (n_27434), .B (n_28892), .Y (n_8803));
NAND2X1 g70556(.A (n_5119), .B (n_12986), .Y (n_12735));
INVX1 g70564(.A (n_11118), .Y (n_15187));
INVX1 g70576(.A (n_8799), .Y (n_8800));
AND2X1 g70580(.A (n_6744), .B (n_28381), .Y (n_10253));
OR2X1 g70582(.A (n_26192), .B (n_28404), .Y (n_10251));
AND2X1 g70583(.A (n_5517), .B (n_6534), .Y (n_8797));
CLKBUFX3 g70587(.A (n_26470), .Y (n_12397));
NOR2X1 g70591(.A (n_8794), .B (n_13247), .Y (n_8795));
NAND2X1 g70594(.A (n_5930), .B (n_11400), .Y (n_12214));
NAND2X1 g70595(.A (n_6577), .B (n_5817), .Y (n_8793));
INVX1 g70604(.A (n_10820), .Y (n_8791));
NAND2X2 g70612(.A (n_8788), .B (n_10495), .Y (n_12802));
NAND2X1 g70614(.A (n_8362), .B (n_27099), .Y (n_12203));
INVX2 g70623(.A (n_11362), .Y (n_12634));
NOR2X1 g70626(.A (n_5034), .B (n_9264), .Y (n_19889));
INVX1 g69616(.A (n_8784), .Y (n_10498));
NAND2X1 g68283(.A (n_5772), .B (n_11354), .Y (n_14934));
NAND2X1 g70635(.A (n_6183), .B (n_9084), .Y (n_12681));
NOR2X1 g70638(.A (n_5631), .B (n_8968), .Y (n_10243));
OR2X1 g70639(.A (n_6462), .B (n_8780), .Y (n_13376));
NAND2X1 g70640(.A (n_8778), .B (n_11052), .Y (n_8779));
NAND2X1 g70641(.A (n_5355), .B (n_8339), .Y (n_13722));
OR2X1 g70645(.A (n_1965), .B (n_25926), .Y (n_8777));
INVX1 g70648(.A (n_8775), .Y (n_10242));
INVX1 g70649(.A (n_8775), .Y (n_8774));
NOR2X1 g70658(.A (n_10315), .B (n_28319), .Y (n_17405));
NOR2X1 g70660(.A (n_2548), .B (n_8709), .Y (n_17472));
NAND2X1 g70668(.A (n_6738), .B (n_7266), .Y (n_8772));
NAND2X1 g70671(.A (n_2013), .B (n_19755), .Y (n_8770));
INVX1 g70675(.A (n_8769), .Y (n_12154));
INVX1 g70678(.A (n_8768), .Y (n_10232));
NOR2X1 g70681(.A (n_6494), .B (n_7325), .Y (n_14747));
NOR2X1 g70688(.A (n_4928), .B (n_8393), .Y (n_10229));
OR2X1 g70693(.A (n_1283), .B (n_8696), .Y (n_28318));
NOR2X1 g70697(.A (n_11924), .B (n_8141), .Y (n_12881));
NOR2X1 g70700(.A (n_4978), .B (n_19398), .Y (n_8763));
NAND2X1 g70705(.A (n_8759), .B (n_4413), .Y (n_14988));
AND2X1 g70710(.A (n_8756), .B (n_11745), .Y (n_8757));
OR2X1 g70713(.A (n_5425), .B (n_28724), .Y (n_8755));
INVX1 g70721(.A (n_7275), .Y (n_15648));
NAND2X1 g70726(.A (n_5628), .B (n_29269), .Y (n_12581));
NAND2X1 g70748(.A (n_2683), .B (n_19755), .Y (n_8749));
NOR2X1 g70751(.A (n_3248), .B (n_9003), .Y (n_10217));
NAND2X1 g70752(.A (n_1907), .B (n_13768), .Y (n_8748));
INVX1 g70754(.A (n_11394), .Y (n_12316));
NAND2X1 g70766(.A (n_1758), .B (n_8520), .Y (n_8747));
INVX1 g70769(.A (n_8746), .Y (n_10216));
NOR2X1 g70771(.A (n_8644), .B (n_11489), .Y (n_15355));
NOR2X1 g70774(.A (n_8569), .B (n_28742), .Y (n_10215));
INVX1 g70782(.A (n_7267), .Y (n_12644));
INVX1 g70787(.A (n_8745), .Y (n_17412));
INVX1 g70793(.A (n_8743), .Y (n_8744));
NOR2X1 g70799(.A (n_3652), .B (n_8742), .Y (n_10209));
NOR2X1 g70808(.A (n_6712), .B (n_14866), .Y (n_10206));
INVX1 g70817(.A (n_8736), .Y (n_10204));
NOR2X1 g70821(.A (n_6687), .B (n_6877), .Y (n_8735));
OR2X1 g70822(.A (n_2433), .B (n_25926), .Y (n_8734));
INVX1 g70834(.A (n_7260), .Y (n_10202));
INVX1 g70844(.A (n_8730), .Y (n_10198));
NAND2X1 g70847(.A (n_8490), .B (n_7366), .Y (n_12852));
NAND2X1 g70855(.A (n_8729), .B (n_383), .Y (n_12868));
INVX1 g70859(.A (n_8724), .Y (n_8725));
NOR2X1 g70865(.A (n_6714), .B (n_2318), .Y (n_8723));
NOR2X1 g70873(.A (n_6616), .B (n_9084), .Y (n_11900));
NAND2X1 g70874(.A (n_8110), .B (n_12784), .Y (n_12549));
NAND2X1 g70882(.A (n_2431), .B (n_8520), .Y (n_8721));
NAND2X1 g70884(.A (n_6087), .B (n_8719), .Y (n_8720));
NAND2X1 g70895(.A (n_7763), .B (n_8865), .Y (n_8715));
INVX1 g70898(.A (n_8714), .Y (n_10185));
INVX1 g70904(.A (n_8713), .Y (n_13472));
INVX1 g70910(.A (n_16394), .Y (n_10182));
INVX1 g70912(.A (n_11027), .Y (n_16601));
INVX1 g70925(.A (n_16492), .Y (n_9905));
NOR2X1 g70929(.A (n_8561), .B (n_8452), .Y (n_8712));
NAND2X1 g70931(.A (n_1608), .B (n_8520), .Y (n_8711));
NOR2X1 g70937(.A (n_8709), .B (n_8708), .Y (n_12129));
NOR2X1 g70940(.A (n_3214), .B (n_26491), .Y (n_8707));
NOR2X1 g70946(.A (n_8706), .B (n_28859), .Y (n_10175));
INVX1 g70957(.A (n_7063), .Y (n_10174));
NOR2X1 g70963(.A (n_4600), .B (n_1547), .Y (n_8704));
NAND2X1 g70964(.A (n_7830), .B (n_7331), .Y (n_8703));
NOR2X1 g70968(.A (n_6544), .B (n_19398), .Y (n_8702));
INVX1 g68265(.A (n_8700), .Y (n_14945));
NAND2X1 g70977(.A (n_5149), .B (n_6342), .Y (n_12541));
NOR2X1 g70979(.A (n_6647), .B (n_17500), .Y (n_8699));
OR2X1 g70980(.A (n_2700), .B (n_8696), .Y (n_25601));
NAND2X1 g70990(.A (n_27367), .B (n_27365), .Y (n_12803));
NAND2X1 g70997(.A (n_4694), .B (n_27669), .Y (n_8695));
NOR2X1 g71007(.A (n_6684), .B (n_11261), .Y (n_8690));
NAND2X1 g71009(.A (n_8687), .B (n_8686), .Y (n_8688));
NAND2X1 g71016(.A (n_28610), .B (n_6753), .Y (n_8684));
OR2X1 g71017(.A (n_8099), .B (n_8682), .Y (n_8683));
INVX1 g71021(.A (n_7220), .Y (n_10152));
INVX1 g71024(.A (n_8681), .Y (n_10150));
INVX1 g71027(.A (n_7240), .Y (n_8680));
AND2X1 g71030(.A (n_3887), .B (n_8679), .Y (n_18254));
INVX1 g71032(.A (n_7237), .Y (n_16539));
NAND2X1 g71034(.A (n_1809), .B (n_8520), .Y (n_8678));
NAND2X1 g71035(.A (n_2281), .B (n_8729), .Y (n_20192));
NAND2X1 g71036(.A (n_5252), .B (n_16787), .Y (n_12723));
INVX1 g71043(.A (n_8675), .Y (n_10144));
OR2X1 g71048(.A (n_5327), .B (n_14866), .Y (n_12256));
NAND2X1 g71052(.A (n_8674), .B (n_9050), .Y (n_10137));
OR2X1 g71059(.A (n_2543), .B (n_13846), .Y (n_8673));
OR2X1 g71060(.A (n_7619), .B (n_27099), .Y (n_8672));
INVX1 g71063(.A (n_8671), .Y (n_10136));
INVX1 g71066(.A (n_8670), .Y (n_12980));
INVX1 g71067(.A (n_8670), .Y (n_8669));
OR2X1 g71070(.A (n_7683), .B (n_14142), .Y (n_8668));
NOR2X1 g71072(.A (n_8666), .B (n_9410), .Y (n_8667));
OR2X1 g71075(.A (n_995), .B (n_13846), .Y (n_8665));
NAND2X1 g71077(.A (n_2872), .B (n_8664), .Y (n_13347));
INVX1 g71081(.A (n_14343), .Y (n_10129));
NAND2X1 g71087(.A (n_5191), .B (n_8662), .Y (n_8663));
INVX1 g71089(.A (n_8660), .Y (n_8661));
NAND2X1 g71096(.A (n_1845), .B (n_8520), .Y (n_8657));
INVX1 g71097(.A (n_8654), .Y (n_8655));
INVX1 g71114(.A (n_8649), .Y (n_8650));
NAND2X1 g71122(.A (n_28611), .B (n_2318), .Y (n_8648));
INVX1 g71126(.A (n_8645), .Y (n_15067));
NOR2X1 g71135(.A (n_8644), .B (n_6005), .Y (n_10119));
INVX1 g71143(.A (n_8641), .Y (n_8642));
NAND2X1 g72674(.A (n_2173), .B (n_8520), .Y (n_8640));
NOR2X1 g72688(.A (n_3193), .B (n_8637), .Y (n_8638));
OR2X1 g71152(.A (n_8635), .B (n_12850), .Y (n_8636));
AOI21X1 g71153(.A0 (n_2973), .A1 (n_28134), .B0 (n_8169), .Y(n_8634));
NAND2X1 g71158(.A (n_10680), .B (n_5936), .Y (n_16644));
INVX1 g71160(.A (n_7212), .Y (n_10112));
NAND2X1 g71163(.A (n_6563), .B (n_9018), .Y (n_8632));
NAND2X1 g71167(.A (n_5179), .B (n_4695), .Y (n_10109));
INVX1 g71170(.A (n_7209), .Y (n_15132));
OR2X1 g71189(.A (n_3401), .B (n_10226), .Y (n_8629));
NAND2X1 g71190(.A (n_2494), .B (n_8520), .Y (n_8628));
INVX2 g71192(.A (n_9167), .Y (n_13073));
OR2X1 g71200(.A (n_9463), .B (n_7321), .Y (n_8627));
NAND2X1 g71216(.A (n_2547), .B (n_13768), .Y (n_28562));
INVX1 g71218(.A (n_8620), .Y (n_8621));
NOR2X1 g71225(.A (n_10495), .B (n_4852), .Y (n_10102));
NAND2X1 g71227(.A (n_29182), .B (n_11850), .Y (n_8619));
NAND2X1 g71235(.A (n_4730), .B (n_16198), .Y (n_29300));
INVX1 g71237(.A (n_7202), .Y (n_8615));
INVX1 g71240(.A (n_8613), .Y (n_8614));
INVX1 g71245(.A (n_7632), .Y (n_10096));
NAND2X1 g71247(.A (n_8611), .B (n_9236), .Y (n_8612));
NAND3X1 g71251(.A (n_16976), .B (n_6696), .C (n_13679), .Y (n_8610));
NAND2X1 g71254(.A (n_2918), .B (n_8520), .Y (n_8608));
NAND2X1 g71255(.A (n_8604), .B (n_3318), .Y (n_8607));
OR2X1 g71268(.A (n_5262), .B (n_6963), .Y (n_8605));
NAND2X2 g71275(.A (n_8604), .B (n_3736), .Y (n_10091));
OR2X1 g71277(.A (n_8603), .B (n_12760), .Y (n_13701));
NOR2X1 g72679(.A (n_6593), .B (n_9917), .Y (n_8598));
NOR2X1 g72682(.A (n_6458), .B (n_13593), .Y (n_9815));
NOR3X1 g71294(.A (n_9819), .B (n_3805), .C (n_28757), .Y (n_8597));
OR2X1 g71302(.A (n_8686), .B (n_11323), .Y (n_8595));
AND2X1 g71303(.A (n_2456), .B (n_10681), .Y (n_20551));
NAND2X1 g71306(.A (n_3183), .B (n_8520), .Y (n_8593));
NAND2X1 g71307(.A (n_5653), .B (n_28433), .Y (n_8592));
NOR2X1 g71954(.A (n_4642), .B (n_9417), .Y (n_8590));
NOR2X1 g71329(.A (n_4164), .B (n_26270), .Y (n_10078));
AOI21X1 g71335(.A0 (n_2990), .A1 (n_12169), .B0 (n_8308), .Y(n_8587));
INVX1 g71344(.A (n_8586), .Y (n_10072));
OR2X1 g71349(.A (n_9463), .B (n_4709), .Y (n_8585));
NOR2X1 g71356(.A (n_3021), .B (n_6366), .Y (n_8584));
NAND2X1 g71357(.A (n_5378), .B (n_15166), .Y (n_8583));
NAND2X1 g71360(.A (n_10163), .B (n_18785), .Y (n_8581));
OR2X1 g71370(.A (n_2590), .B (n_25926), .Y (n_8580));
NAND2X1 g71371(.A (n_2408), .B (n_13787), .Y (n_25722));
OR2X1 g71372(.A (n_4642), .B (n_263), .Y (n_12289));
NOR2X1 g71373(.A (n_6148), .B (n_9078), .Y (n_8576));
NOR2X1 g71377(.A (n_8493), .B (n_27365), .Y (n_10063));
OR2X1 g71379(.A (n_8076), .B (n_10495), .Y (n_10061));
NOR2X1 g71403(.A (n_8090), .B (n_4979), .Y (n_28832));
NAND2X1 g71404(.A (n_14855), .B (n_12335), .Y (n_8573));
NAND2X1 g71407(.A (n_29214), .B (n_4612), .Y (n_8572));
AOI21X1 g71415(.A0 (n_7701), .A1 (n_6833), .B0 (n_26491), .Y(n_8571));
NAND2X1 g71417(.A (n_2868), .B (n_13787), .Y (n_8570));
OR2X1 g71419(.A (n_8569), .B (n_7496), .Y (n_12754));
INVX1 g71424(.A (n_11386), .Y (n_8568));
NAND2X1 g71427(.A (n_7121), .B (n_9899), .Y (n_14007));
INVX1 g71428(.A (n_8566), .Y (n_8567));
NAND2X1 g71432(.A (n_8564), .B (n_6219), .Y (n_8565));
NAND2X1 g71437(.A (n_6350), .B (n_1647), .Y (n_16391));
NOR2X1 g71444(.A (n_8561), .B (n_8560), .Y (n_17409));
NOR2X1 g71445(.A (n_27603), .B (n_18785), .Y (n_8559));
AOI21X1 g71453(.A0 (n_5923), .A1 (n_6226), .B0 (n_8556), .Y (n_8557));
INVX1 g71454(.A (n_13142), .Y (n_8555));
INVX1 g71457(.A (n_9565), .Y (n_10044));
NAND2X1 g71462(.A (n_4418), .B (n_27746), .Y (n_8554));
NOR2X1 g71470(.A (n_6462), .B (n_6470), .Y (n_8553));
INVX1 g71473(.A (n_8552), .Y (n_12815));
NOR2X1 g71481(.A (n_4547), .B (n_8548), .Y (n_8549));
INVX1 g71483(.A (n_8545), .Y (n_8546));
OR2X1 g71486(.A (n_3806), .B (n_9783), .Y (n_10037));
NOR2X1 g71491(.A (n_3039), .B (n_3920), .Y (n_10035));
INVX1 g71499(.A (n_11042), .Y (n_11501));
INVX1 g71534(.A (n_8543), .Y (n_8544));
OR2X1 g71537(.A (n_8541), .B (n_8540), .Y (n_8542));
INVX1 g71539(.A (n_7826), .Y (n_8539));
NAND2X1 g71542(.A (n_5334), .B (n_16466), .Y (n_8538));
OR2X1 g71543(.A (n_1542), .B (n_25926), .Y (n_8537));
OR2X1 g71547(.A (n_3541), .B (n_10226), .Y (n_8536));
NAND3X1 g71549(.A (n_8534), .B (n_5271), .C (n_15473), .Y (n_8535));
NAND2X1 g71551(.A (n_1727), .B (n_13768), .Y (n_25731));
NOR2X1 g71559(.A (n_6556), .B (n_28375), .Y (n_8532));
INVX1 g71561(.A (n_16825), .Y (n_10027));
NAND2X1 g71567(.A (n_8564), .B (n_6043), .Y (n_12373));
OR2X1 g71574(.A (n_20526), .B (n_14142), .Y (n_8529));
INVX1 g71578(.A (n_10992), .Y (n_10023));
INVX1 g71589(.A (n_8527), .Y (n_13026));
OR2X1 g71597(.A (n_1961), .B (n_25926), .Y (n_8526));
NAND2X1 g71598(.A (n_8524), .B (n_9783), .Y (n_8525));
OR2X1 g71605(.A (n_1749), .B (n_13846), .Y (n_8522));
NAND2X1 g71609(.A (n_6113), .B (n_8520), .Y (n_8521));
NAND2X1 g71610(.A (n_5453), .B (n_15894), .Y (n_8519));
NAND2X1 g71611(.A (n_2550), .B (n_8520), .Y (n_8518));
INVX1 g71615(.A (n_10812), .Y (n_10014));
OR2X1 g71618(.A (n_29329), .B (n_27688), .Y (n_12138));
INVX1 g71628(.A (n_8515), .Y (n_10012));
INVX1 g71632(.A (n_8514), .Y (n_11563));
NAND2X1 g71634(.A (n_6598), .B (n_28642), .Y (n_8513));
NAND2X1 g71639(.A (n_4196), .B (n_8865), .Y (n_12349));
INVX1 g71641(.A (n_8511), .Y (n_12472));
NAND2X1 g71645(.A (n_4166), .B (n_6534), .Y (n_8510));
NAND2X1 g71649(.A (n_2436), .B (n_19755), .Y (n_8508));
NAND2X1 g71658(.A (n_3201), .B (n_8520), .Y (n_8507));
INVX1 g71661(.A (n_13310), .Y (n_10005));
NOR2X1 g71665(.A (n_3871), .B (n_12298), .Y (n_8505));
NOR2X1 g71669(.A (n_8503), .B (n_5691), .Y (n_8504));
INVX1 g71680(.A (n_18552), .Y (n_8502));
OR2X1 g71694(.A (n_5250), .B (n_8499), .Y (n_8500));
INVX1 g71696(.A (n_12883), .Y (n_8498));
INVX1 g71704(.A (n_8496), .Y (n_8497));
NOR2X1 g71721(.A (n_6536), .B (n_10389), .Y (n_8495));
NOR2X1 g71722(.A (n_8493), .B (n_13815), .Y (n_15072));
NOR2X1 g71724(.A (n_8491), .B (n_7553), .Y (n_8492));
INVX1 g71727(.A (n_11390), .Y (n_9995));
NAND2X1 g71735(.A (n_12858), .B (n_8490), .Y (n_12404));
NOR2X1 g71739(.A (n_3039), .B (n_7777), .Y (n_9993));
NOR2X1 g71743(.A (n_4989), .B (n_8499), .Y (n_8489));
NOR2X1 g71747(.A (n_8834), .B (n_1807), .Y (n_9990));
NAND2X1 g71750(.A (n_8487), .B (n_27603), .Y (n_8488));
CLKBUFX3 g71759(.A (n_10791), .Y (n_13602));
INVX1 g71760(.A (n_10791), .Y (n_25654));
OR2X1 g71763(.A (n_2532), .B (n_13846), .Y (n_8484));
OR2X1 g71764(.A (n_2524), .B (n_25926), .Y (n_8483));
INVX1 g71765(.A (n_8481), .Y (n_8482));
OAI21X1 g71771(.A0 (n_6827), .A1 (n_6554), .B0 (n_6258), .Y (n_8480));
INVX1 g72652(.A (n_8477), .Y (n_13031));
NOR2X1 g71789(.A (n_6972), .B (n_3017), .Y (n_8473));
OR2X1 g71796(.A (n_8471), .B (n_8470), .Y (n_8472));
NAND2X1 g71803(.A (n_11078), .B (n_9795), .Y (n_8469));
OR2X1 g71809(.A (n_2676), .B (n_8696), .Y (n_25760));
OR2X1 g71811(.A (n_6581), .B (n_8467), .Y (n_9980));
INVX1 g71815(.A (n_8466), .Y (n_9977));
NOR2X1 g71818(.A (n_3900), .B (n_7006), .Y (n_12823));
NOR2X1 g71826(.A (n_6701), .B (n_10100), .Y (n_8464));
INVX1 g71833(.A (n_13277), .Y (n_9968));
NAND2X1 g71843(.A (n_8556), .B (n_15507), .Y (n_8460));
INVX1 g71847(.A (n_7072), .Y (n_12781));
INVX1 g71857(.A (n_8458), .Y (n_8459));
NAND2X1 g71878(.A (n_4427), .B (n_6659), .Y (n_18965));
INVX1 g71898(.A (n_8454), .Y (n_14745));
NOR2X1 g70962(.A (n_3080), .B (n_13593), .Y (n_10171));
NOR2X1 g71907(.A (n_7841), .B (n_8452), .Y (n_11795));
NAND2X1 g71908(.A (n_2413), .B (n_19755), .Y (n_8451));
NOR2X1 g71910(.A (n_26491), .B (n_3705), .Y (n_9955));
NOR2X1 g71913(.A (n_7937), .B (n_9335), .Y (n_9953));
OR2X1 g71914(.A (n_4908), .B (n_8564), .Y (n_8449));
NAND2X1 g71915(.A (n_1589), .B (n_19755), .Y (n_8448));
INVX1 g71916(.A (n_8445), .Y (n_8447));
AND2X1 g71921(.A (n_5532), .B (n_13239), .Y (n_8444));
NAND2X1 g71927(.A (n_5502), .B (n_4181), .Y (n_8443));
OR2X1 g71929(.A (n_8218), .B (n_7325), .Y (n_11520));
AND2X1 g71935(.A (n_8441), .B (n_8637), .Y (n_8442));
INVX1 g71937(.A (n_7144), .Y (n_15909));
NOR2X1 g71940(.A (n_8438), .B (n_8437), .Y (n_8439));
NOR2X1 g71942(.A (n_6640), .B (n_8435), .Y (n_8436));
NOR2X1 g71945(.A (n_3582), .B (n_11253), .Y (n_10049));
INVX1 g71965(.A (n_7199), .Y (n_14393));
NAND2X1 g71968(.A (n_6422), .B (n_5015), .Y (n_11522));
OR2X1 g71975(.A (n_2416), .B (n_10226), .Y (n_8429));
INVX1 g71987(.A (n_8427), .Y (n_12892));
NAND2X1 g71991(.A (n_8425), .B (n_5558), .Y (n_8426));
NAND2X1 g71992(.A (n_14386), .B (n_6312), .Y (n_8424));
INVX1 g71998(.A (n_7053), .Y (n_14381));
OR2X1 g72000(.A (n_4539), .B (n_3480), .Y (n_8423));
INVX1 g72003(.A (n_8421), .Y (n_8422));
INVX1 g72008(.A (n_7050), .Y (n_8420));
OR2X1 g72020(.A (n_8418), .B (n_7787), .Y (n_8419));
INVX2 g72030(.A (n_8417), .Y (n_9933));
OR2X1 g72034(.A (n_3122), .B (n_8974), .Y (n_14815));
NAND2X1 g72052(.A (n_3616), .B (n_5255), .Y (n_8415));
INVX1 g72057(.A (n_8414), .Y (n_13360));
OR2X1 g72067(.A (n_8524), .B (n_7479), .Y (n_8412));
NAND3X1 g72068(.A (n_15507), .B (n_5447), .C (n_5151), .Y (n_8411));
NAND2X1 g72076(.A (n_8490), .B (n_9118), .Y (n_14821));
NAND2X1 g72081(.A (n_2051), .B (n_8520), .Y (n_8408));
NAND2X1 g72085(.A (n_8404), .B (n_13855), .Y (n_8405));
INVX1 g72087(.A (n_7476), .Y (n_8403));
OR2X1 g72090(.A (n_6699), .B (n_14624), .Y (n_8402));
INVX1 g72100(.A (n_8398), .Y (n_12402));
NAND2X1 g72106(.A (n_12268), .B (n_8396), .Y (n_8397));
NAND2X1 g72111(.A (n_3192), .B (n_8520), .Y (n_8395));
NAND2X1 g72121(.A (n_8393), .B (n_8392), .Y (n_12446));
NAND2X1 g72122(.A (n_6258), .B (n_4859), .Y (n_8391));
OR2X1 g72138(.A (n_8756), .B (n_17260), .Y (n_8390));
NOR2X1 g72140(.A (n_4203), .B (n_17020), .Y (n_8389));
INVX2 g72154(.A (n_7606), .Y (n_15090));
NAND2X1 g72163(.A (n_5042), .B (n_5247), .Y (n_8388));
INVX1 g72177(.A (n_7018), .Y (n_12973));
NAND2X1 g72184(.A (n_1854), .B (n_19755), .Y (n_8386));
NAND2X1 g72191(.A (n_2588), .B (n_13768), .Y (n_25611));
NAND2X1 g72192(.A (n_2516), .B (n_8520), .Y (n_8384));
NAND2X1 g72196(.A (n_1658), .B (n_8520), .Y (n_8383));
NOR2X1 g72202(.A (n_27434), .B (n_25664), .Y (n_8382));
NAND2X1 g72206(.A (n_4855), .B (n_4689), .Y (n_15998));
NAND2X1 g72207(.A (n_8380), .B (n_8379), .Y (n_8381));
NAND2X1 g72217(.A (n_15919), .B (n_8378), .Y (n_13372));
INVX1 g72219(.A (n_8377), .Y (n_15070));
NOR2X1 g72223(.A (n_6620), .B (n_9511), .Y (n_9903));
NAND2X1 g72224(.A (n_2591), .B (n_13768), .Y (n_25788));
NOR2X1 g72237(.A (n_3992), .B (n_17864), .Y (n_8375));
INVX1 g71886(.A (n_8371), .Y (n_12161));
NAND2X1 g72257(.A (n_10094), .B (n_11323), .Y (n_12629));
OR2X1 g72261(.A (n_3021), .B (n_8635), .Y (n_8370));
INVX1 g72267(.A (n_7662), .Y (n_9889));
NOR2X1 g72274(.A (n_8425), .B (n_8367), .Y (n_8368));
NAND2X1 g72275(.A (n_8817), .B (n_5884), .Y (n_8366));
NAND2X1 g72277(.A (n_2455), .B (n_13768), .Y (n_25603));
NAND2X1 g72278(.A (n_7840), .B (n_8931), .Y (n_8364));
NAND2X1 g72279(.A (n_8363), .B (n_8362), .Y (n_12844));
OR2X1 g72293(.A (n_1968), .B (n_25926), .Y (n_8361));
NAND2X1 g72296(.A (n_3518), .B (n_9388), .Y (n_8360));
NOR2X1 g72307(.A (n_8978), .B (n_3818), .Y (n_9882));
INVX1 g72321(.A (n_12673), .Y (n_11135));
OR2X1 g70919(.A (n_2660), .B (n_10226), .Y (n_8358));
NAND2X1 g72323(.A (n_2148), .B (n_13787), .Y (n_8357));
AND2X1 g72325(.A (n_8355), .B (n_18205), .Y (n_8356));
NOR2X1 g72331(.A (n_2318), .B (n_4385), .Y (n_9876));
INVX1 g72624(.A (n_8354), .Y (n_12468));
INVX1 g72334(.A (n_9574), .Y (n_8353));
INVX1 g72343(.A (n_8351), .Y (n_8349));
OR2X1 g72349(.A (n_5315), .B (n_7032), .Y (n_8348));
NOR2X1 g72351(.A (n_28037), .B (n_3644), .Y (n_9874));
OR2X1 g72352(.A (n_4208), .B (n_8346), .Y (n_8347));
OR2X1 g72353(.A (n_2846), .B (n_13846), .Y (n_8345));
OR2X1 g72354(.A (n_2900), .B (n_8343), .Y (n_8344));
NAND2X1 g72355(.A (n_8342), .B (n_8664), .Y (n_12376));
OR2X1 g72358(.A (n_5491), .B (n_8708), .Y (n_8341));
NOR2X1 g72364(.A (n_8339), .B (n_8253), .Y (n_9872));
INVX1 g72365(.A (n_8338), .Y (n_14574));
NAND2X1 g72371(.A (n_12162), .B (n_8664), .Y (n_8337));
INVX1 g72374(.A (n_8335), .Y (n_8336));
INVX1 g72377(.A (n_7802), .Y (n_12638));
NAND2X1 g72387(.A (n_2429), .B (n_8520), .Y (n_8334));
NOR2X1 g72390(.A (n_7593), .B (n_29385), .Y (n_9869));
INVX1 g72393(.A (n_12383), .Y (n_12964));
OR2X1 g72396(.A (n_8524), .B (n_11253), .Y (n_8333));
INVX1 g72398(.A (n_8330), .Y (n_8331));
INVX1 g72400(.A (n_8328), .Y (n_8329));
INVX1 g72404(.A (n_8326), .Y (n_14120));
NOR2X1 g72411(.A (n_8719), .B (n_6185), .Y (n_8325));
INVX1 g72413(.A (n_21820), .Y (n_8324));
NAND2X1 g72424(.A (n_4094), .B (n_8284), .Y (n_8323));
OR2X1 g72425(.A (n_8321), .B (n_6889), .Y (n_8322));
INVX1 g72430(.A (n_8319), .Y (n_8320));
NAND2X1 g72433(.A (n_2895), .B (n_9336), .Y (n_8318));
NAND2X1 g72434(.A (n_8317), .B (n_5930), .Y (n_15014));
INVX1 g72436(.A (n_28038), .Y (n_8314));
NAND2X1 g72457(.A (n_8015), .B (n_28642), .Y (n_19949));
INVX1 g72460(.A (n_7833), .Y (n_8309));
NAND2X1 g72471(.A (n_8308), .B (n_3301), .Y (n_9856));
NAND2X1 g72472(.A (n_4695), .B (n_15776), .Y (n_17134));
OR2X1 g72479(.A (n_7578), .B (n_5630), .Y (n_8306));
INVX1 g72485(.A (n_5006), .Y (n_12918));
NAND2X1 g72499(.A (n_8729), .B (n_1057), .Y (n_19947));
INVX1 g72502(.A (n_11221), .Y (n_12389));
INVX4 g75789(.A (n_9878), .Y (n_25597));
INVX1 g72511(.A (n_6967), .Y (n_8302));
INVX1 g72523(.A (n_8301), .Y (n_21649));
INVX2 g72527(.A (n_8300), .Y (n_9632));
OR2X1 g72529(.A (n_2585), .B (n_13846), .Y (n_8299));
INVX1 g72531(.A (n_8298), .Y (n_12278));
NAND2X1 g72536(.A (n_8296), .B (n_8295), .Y (n_8297));
NAND2X1 g72538(.A (n_11662), .B (n_9276), .Y (n_8294));
NAND2X1 g72551(.A (n_16973), .B (n_4258), .Y (n_8292));
NOR2X1 g72559(.A (n_8290), .B (n_16754), .Y (n_8291));
INVX2 g72563(.A (n_8289), .Y (n_13003));
INVX1 g72566(.A (n_8287), .Y (n_8288));
INVX1 g72570(.A (n_11304), .Y (n_18278));
INVX1 g72581(.A (n_8285), .Y (n_8286));
OR2X1 g72589(.A (n_8284), .B (n_6005), .Y (n_9831));
NAND2X1 g72590(.A (n_1473), .B (n_8520), .Y (n_8283));
OR2X1 g72591(.A (n_7213), .B (n_9645), .Y (n_8282));
NAND2X1 g72599(.A (n_13177), .B (n_12568), .Y (n_8277));
OR2X1 g72600(.A (n_3162), .B (n_9486), .Y (n_8276));
NAND2X1 g72601(.A (n_12784), .B (n_4757), .Y (n_8275));
INVX1 g72603(.A (n_8273), .Y (n_8274));
NOR2X1 g72620(.A (n_3646), .B (n_11400), .Y (n_8272));
INVX1 g72608(.A (n_11345), .Y (n_9828));
INVX1 g72613(.A (n_8269), .Y (n_8268));
INVX1 g70892(.A (n_8266), .Y (n_8267));
NAND2X1 g72628(.A (n_2505), .B (n_8520), .Y (n_8265));
NAND2X1 g72629(.A (n_6698), .B (n_8263), .Y (n_8264));
INVX1 g72630(.A (n_10979), .Y (n_8262));
INVX1 g72644(.A (n_6947), .Y (n_14517));
NOR2X1 g72649(.A (n_5921), .B (n_28423), .Y (n_8261));
NAND2X1 g72660(.A (n_1477), .B (n_8520), .Y (n_8260));
INVX1 g72663(.A (n_8258), .Y (n_8259));
NAND2X1 g72667(.A (n_5355), .B (n_11400), .Y (n_18697));
NAND2X1 g72675(.A (n_2055), .B (n_8520), .Y (n_8256));
NAND2X1 g72690(.A (n_4162), .B (n_8254), .Y (n_8255));
OR2X1 g72693(.A (n_8253), .B (n_28373), .Y (n_12649));
INVX1 g72697(.A (n_8251), .Y (n_9814));
NAND2X2 g70880(.A (n_10127), .B (n_8250), .Y (n_10193));
OR2X1 g72701(.A (n_7614), .B (n_8682), .Y (n_8249));
NOR2X1 g72704(.A (n_4788), .B (n_14055), .Y (n_9811));
OR2X1 g72705(.A (n_8686), .B (n_8540), .Y (n_8247));
NAND2X1 g72706(.A (n_14725), .B (n_8548), .Y (n_8246));
AOI21X1 g72713(.A0 (n_6836), .A1 (n_6856), .B0 (n_7593), .Y (n_8245));
OR2X1 g72717(.A (n_8243), .B (n_3386), .Y (n_8244));
NOR2X1 g72718(.A (n_6633), .B (n_13490), .Y (n_12342));
NOR2X1 g72727(.A (n_8404), .B (n_9942), .Y (n_9808));
INVX2 g75777(.A (n_8240), .Y (n_11823));
NOR2X1 g72737(.A (n_7757), .B (n_18320), .Y (n_8239));
NOR2X1 g72751(.A (n_6461), .B (n_29244), .Y (n_28816));
NAND2X1 g72752(.A (n_10094), .B (n_8560), .Y (n_13720));
INVX1 g72759(.A (n_7328), .Y (n_8235));
NOR2X1 g72761(.A (n_8343), .B (n_5704), .Y (n_8234));
NAND2X1 g72765(.A (n_15636), .B (n_9978), .Y (n_8233));
NAND2X1 g72772(.A (n_2441), .B (n_13768), .Y (n_25773));
NOR2X1 g72774(.A (n_7722), .B (n_14055), .Y (n_8231));
OR2X1 g72783(.A (n_2198), .B (n_25926), .Y (n_8229));
OR2X1 g72786(.A (n_8719), .B (n_8227), .Y (n_8228));
INVX1 g72797(.A (n_8223), .Y (n_8224));
NAND2X1 g72805(.A (n_6327), .B (n_8794), .Y (n_8222));
OR2X1 g72809(.A (n_11435), .B (n_29228), .Y (n_8221));
INVX1 g72810(.A (n_6923), .Y (n_14880));
INVX1 g72813(.A (n_7523), .Y (n_14467));
NAND2X1 g72815(.A (n_7778), .B (n_28037), .Y (n_8219));
OR2X1 g72816(.A (n_8218), .B (n_8217), .Y (n_13704));
NAND2X1 g72820(.A (n_11435), .B (n_29269), .Y (n_8216));
NAND2X1 g72826(.A (n_8491), .B (n_28375), .Y (n_8215));
NOR2X1 g72831(.A (n_6727), .B (n_4721), .Y (n_8213));
OR2X1 g72832(.A (n_2185), .B (n_25926), .Y (n_8212));
NAND2X1 g72833(.A (n_5619), .B (n_8209), .Y (n_8210));
NAND2X1 g72846(.A (n_10094), .B (n_8435), .Y (n_19430));
OR2X1 g72847(.A (n_8404), .B (n_28692), .Y (n_29419));
INVX1 g72853(.A (n_11259), .Y (n_12599));
NAND2X1 g72857(.A (n_6952), .B (n_7420), .Y (n_8206));
NAND2X1 g72858(.A (n_3811), .B (n_8520), .Y (n_8205));
NOR2X1 g70868(.A (n_8756), .B (n_29228), .Y (n_10194));
NOR2X1 g72861(.A (n_3206), .B (n_5085), .Y (n_9787));
OR2X1 g72863(.A (n_3260), .B (n_1647), .Y (n_9785));
NAND2X1 g72869(.A (n_28991), .B (n_7598), .Y (n_10693));
NOR2X1 g72885(.A (n_29275), .B (n_9674), .Y (n_8203));
OR2X1 g72886(.A (n_1321), .B (n_25926), .Y (n_8202));
OR2X1 g72889(.A (n_6661), .B (n_7410), .Y (n_15256));
NOR2X1 g72891(.A (n_7767), .B (n_7496), .Y (n_8201));
OR2X1 g72892(.A (n_5122), .B (n_13846), .Y (n_8199));
NAND2X1 g74047(.A (n_6338), .B (n_11276), .Y (n_8198));
INVX1 g74640(.A (n_8197), .Y (n_9651));
INVX1 g72905(.A (n_6901), .Y (n_10819));
NAND2X1 g72910(.A (n_3186), .B (n_19755), .Y (n_8194));
INVX1 g72924(.A (n_7635), .Y (n_10841));
OR2X1 g72927(.A (n_4684), .B (n_25926), .Y (n_8193));
OR2X1 g72928(.A (n_9236), .B (n_8191), .Y (n_8192));
NOR2X1 g72931(.A (n_12494), .B (n_8346), .Y (n_12748));
NAND2X1 g72939(.A (n_6809), .B (n_7319), .Y (n_8189));
INVX1 g72940(.A (n_6895), .Y (n_8188));
OR2X1 g72943(.A (n_7984), .B (n_12105), .Y (n_8187));
NAND2X1 g72944(.A (n_4457), .B (n_6534), .Y (n_8186));
INVX1 g72956(.A (n_8185), .Y (n_9773));
INVX1 g72969(.A (n_6888), .Y (n_10947));
INVX1 g72975(.A (n_13301), .Y (n_12970));
INVX1 g72991(.A (n_8184), .Y (n_9765));
NAND2X1 g72995(.A (n_2024), .B (n_19755), .Y (n_8183));
AND2X1 g73006(.A (n_5832), .B (n_11861), .Y (n_8181));
NOR2X1 g73018(.A (n_5921), .B (n_11576), .Y (n_8177));
INVX1 g73021(.A (n_8176), .Y (n_18400));
AND2X1 g73030(.A (n_8837), .B (n_8172), .Y (n_8173));
INVX1 g73031(.A (n_8170), .Y (n_8171));
NAND2X1 g72234(.A (n_17884), .B (n_8169), .Y (n_9896));
INVX1 g73037(.A (n_7682), .Y (n_12275));
NAND2X1 g73041(.A (n_4093), .B (n_8729), .Y (n_20743));
INVX2 g73044(.A (n_8167), .Y (n_9759));
INVX1 g73047(.A (n_7696), .Y (n_8166));
INVX1 g73051(.A (n_8164), .Y (n_8165));
NOR2X1 g73061(.A (n_29329), .B (n_11253), .Y (n_8161));
OR2X1 g73069(.A (n_2403), .B (n_25926), .Y (n_8159));
INVX1 g73073(.A (n_10850), .Y (n_9754));
NAND2X1 g73075(.A (n_2552), .B (n_13787), .Y (n_25705));
INVX1 g73076(.A (n_13226), .Y (n_8157));
INVX1 g73088(.A (n_6865), .Y (n_12486));
INVX1 g73090(.A (n_8154), .Y (n_8155));
INVX1 g73093(.A (n_11076), .Y (n_8152));
OR2X1 g73098(.A (n_1656), .B (n_13846), .Y (n_8149));
NOR2X1 g73110(.A (n_8441), .B (n_29427), .Y (n_8148));
NOR2X1 g73118(.A (n_5103), .B (n_6005), .Y (n_9746));
AOI21X1 g73128(.A0 (n_2373), .A1 (n_7658), .B0 (n_8604), .Y (n_8145));
OR2X1 g73129(.A (n_27075), .B (n_17260), .Y (n_14840));
OR2X1 g73131(.A (n_1760), .B (n_25926), .Y (n_8144));
NAND2X1 g73137(.A (n_2234), .B (n_13787), .Y (n_8143));
OR2X1 g73138(.A (n_6527), .B (n_8141), .Y (n_8142));
OR2X1 g73139(.A (n_8379), .B (n_8139), .Y (n_8140));
OR2X1 g73140(.A (n_8137), .B (n_9442), .Y (n_8138));
NAND2X1 g73141(.A (n_2556), .B (n_8520), .Y (n_8135));
NAND2X1 g73144(.A (n_5628), .B (n_27990), .Y (n_15600));
NAND2X1 g73155(.A (n_4289), .B (n_29189), .Y (n_8132));
NAND2X1 g73165(.A (n_12292), .B (n_8811), .Y (n_25571));
INVX1 g73171(.A (n_6846), .Y (n_9730));
NOR2X1 g73177(.A (n_2654), .B (n_6740), .Y (n_8130));
OR2X1 g73182(.A (n_11067), .B (n_29269), .Y (n_14864));
NAND2X1 g73185(.A (n_5981), .B (n_4819), .Y (n_8129));
INVX1 g73189(.A (n_7823), .Y (n_17071));
NOR2X1 g73195(.A (n_1233), .B (n_8127), .Y (n_8128));
INVX1 g73197(.A (n_6843), .Y (n_9722));
OR2X1 g73199(.A (n_2935), .B (n_13846), .Y (n_8126));
NAND2X1 g73201(.A (n_8846), .B (n_4855), .Y (n_9720));
NAND2X1 g73205(.A (n_5163), .B (n_15776), .Y (n_8125));
NAND2X1 g73208(.A (n_12155), .B (n_8362), .Y (n_8124));
OR2X1 g73210(.A (n_1712), .B (n_13846), .Y (n_8123));
NAND2X1 g73212(.A (n_4695), .B (n_6805), .Y (n_12448));
OR2X1 g73216(.A (n_4732), .B (n_8120), .Y (n_8121));
OR2X1 g73219(.A (n_5492), .B (n_8118), .Y (n_8119));
OAI21X1 g73230(.A0 (n_8116), .A1 (n_1353), .B0 (n_12292), .Y(n_8117));
OAI21X1 g73231(.A0 (n_4828), .A1 (n_28472), .B0 (n_7113), .Y(n_8115));
NAND2X1 g73235(.A (n_2090), .B (n_8113), .Y (n_8114));
NAND2X1 g73238(.A (n_14667), .B (n_6515), .Y (n_8112));
OR2X1 g73240(.A (n_5472), .B (n_8110), .Y (n_8111));
AOI21X1 g73246(.A0 (n_3774), .A1 (n_4026), .B0 (n_1939), .Y (n_8109));
AOI21X1 g73251(.A0 (n_7730), .A1 (n_4388), .B0 (n_3749), .Y (n_8108));
AOI21X1 g73256(.A0 (n_6327), .A1 (n_5073), .B0 (n_3443), .Y (n_8107));
AOI21X1 g73261(.A0 (n_8105), .A1 (n_2254), .B0 (n_6211), .Y (n_8106));
AOI21X1 g73263(.A0 (n_3170), .A1 (n_3087), .B0 (n_3258), .Y (n_8104));
OAI21X1 g75953(.A0 (n_383), .A1 (n_2231), .B0 (n_8101), .Y (n_8103));
AOI21X1 g73283(.A0 (n_29119), .A1 (n_4581), .B0 (n_8099), .Y(n_8100));
AOI21X1 g73284(.A0 (n_7196), .A1 (n_8097), .B0 (n_6397), .Y (n_8098));
AOI21X1 g73287(.A0 (n_1142), .A1 (n_5151), .B0 (n_5405), .Y (n_8096));
NAND2X1 g75952(.A (n_12222), .B (n_4100), .Y (n_8095));
AOI21X1 g73290(.A0 (n_8093), .A1 (n_3936), .B0 (n_5504), .Y (n_8094));
AOI21X1 g73293(.A0 (n_8945), .A1 (n_3512), .B0 (n_5210), .Y (n_8092));
AOI21X1 g73295(.A0 (n_8090), .A1 (n_3493), .B0 (n_5550), .Y (n_8091));
OR2X1 g73324(.A (n_3422), .B (n_11576), .Y (n_8089));
INVX1 g70804(.A (n_11311), .Y (n_8088));
INVX2 g73340(.A (n_8086), .Y (n_11901));
INVX1 g69373(.A (n_10806), .Y (n_8085));
NOR2X1 g72598(.A (n_7418), .B (n_5294), .Y (n_9829));
INVX1 g73457(.A (n_8083), .Y (n_11864));
INVX1 g73495(.A (n_7637), .Y (n_11749));
INVX1 g73520(.A (n_6784), .Y (n_12106));
INVX1 g73523(.A (n_10546), .Y (n_8080));
OR2X1 g73267(.A (n_6220), .B (n_8078), .Y (n_8079));
NAND2X1 g70792(.A (n_4342), .B (n_8076), .Y (n_8077));
NAND2X1 g73588(.A (n_5947), .B (n_11835), .Y (n_8075));
NAND2X1 g73607(.A (n_4019), .B (n_11998), .Y (n_8073));
NOR2X1 g69354(.A (n_27371), .B (n_8070), .Y (n_8071));
INVX2 g75440(.A (n_8068), .Y (n_11728));
NAND2X1 g68092(.A (n_7424), .B (n_1347), .Y (n_8064));
INVX1 g73697(.A (n_8063), .Y (n_11984));
NAND2X1 g70778(.A (n_8729), .B (n_9118), .Y (n_8062));
OR2X1 g73753(.A (n_2864), .B (n_9388), .Y (n_8059));
INVX1 g71784(.A (n_7089), .Y (n_12224));
INVX1 g69338(.A (n_14493), .Y (n_10565));
INVX1 g73857(.A (n_9803), .Y (n_8052));
INVX1 g71792(.A (n_7088), .Y (n_12945));
NAND2X1 g75535(.A (n_7955), .B (n_8928), .Y (n_8049));
NAND2X1 g73911(.A (n_7698), .B (n_8452), .Y (n_11743));
INVX1 g73924(.A (n_8047), .Y (n_8048));
NOR2X1 g69684(.A (n_8039), .B (n_8090), .Y (n_14528));
INVX1 g73955(.A (n_8037), .Y (n_8038));
INVX1 g73967(.A (n_7890), .Y (n_8036));
OR2X1 g73994(.A (n_3809), .B (n_9500), .Y (n_8034));
NOR2X1 g74002(.A (n_8452), .B (n_4736), .Y (n_11660));
NOR2X1 g74013(.A (n_7095), .B (n_29286), .Y (n_11667));
INVX1 g74027(.A (n_9900), .Y (n_11801));
INVX2 g74028(.A (n_9900), .Y (n_28246));
INVX1 g74055(.A (n_8030), .Y (n_9669));
NOR2X1 g75929(.A (n_4084), .B (n_7938), .Y (n_8029));
INVX1 g74126(.A (n_8024), .Y (n_8025));
NAND2X1 g74143(.A (n_6255), .B (n_28733), .Y (n_8023));
INVX1 g74183(.A (n_8022), .Y (n_9665));
NOR2X1 g74206(.A (n_7845), .B (n_13490), .Y (n_8021));
NAND2X1 g74227(.A (n_7981), .B (n_15968), .Y (n_8020));
NAND2X1 g74231(.A (n_8018), .B (n_11052), .Y (n_8019));
NAND2X1 g74273(.A (n_8016), .B (n_20325), .Y (n_8017));
INVX1 g74291(.A (n_7753), .Y (n_9661));
NAND2X2 g72574(.A (n_8015), .B (n_8093), .Y (n_12587));
OR2X1 g74329(.A (n_5030), .B (n_28733), .Y (n_8014));
INVX1 g74338(.A (n_6676), .Y (n_8013));
NOR2X1 g74379(.A (n_6735), .B (n_7728), .Y (n_8012));
INVX1 g74417(.A (n_10140), .Y (n_8010));
INVX1 g70718(.A (n_8009), .Y (n_10223));
AOI21X1 g73265(.A0 (n_5502), .A1 (n_6706), .B0 (n_3938), .Y (n_8008));
CLKBUFX1 g74485(.A (n_9779), .Y (n_11976));
INVX1 g74491(.A (n_9930), .Y (n_8007));
NAND2X1 g71758(.A (n_5318), .B (n_9417), .Y (n_9988));
OR2X1 g74516(.A (n_4772), .B (n_3422), .Y (n_8006));
INVX1 g74531(.A (n_10146), .Y (n_9654));
INVX1 g74583(.A (n_8000), .Y (n_8001));
INVX1 g74624(.A (n_7999), .Y (n_13991));
INVX1 g74632(.A (n_7997), .Y (n_12078));
INVX1 g74645(.A (n_7995), .Y (n_7996));
NOR2X1 g71745(.A (n_5468), .B (n_29065), .Y (n_7992));
OR2X1 g73260(.A (n_4077), .B (n_7984), .Y (n_7985));
INVX1 g74831(.A (n_10272), .Y (n_11752));
OR2X1 g74850(.A (n_5021), .B (n_9442), .Y (n_7983));
NAND2X1 g74869(.A (n_7981), .B (n_17411), .Y (n_7982));
INVX1 g74883(.A (n_10453), .Y (n_7979));
NOR2X1 g74894(.A (n_6364), .B (n_29256), .Y (n_7978));
NAND2X1 g68039(.A (n_7976), .B (n_2779), .Y (n_10880));
INVX1 g74901(.A (n_7974), .Y (n_7975));
INVX1 g74907(.A (n_7973), .Y (n_11734));
NOR2X1 g74933(.A (n_7610), .B (n_13834), .Y (n_11671));
NAND2X1 g74935(.A (n_5212), .B (n_9783), .Y (n_7971));
INVX1 g75001(.A (n_7968), .Y (n_7969));
INVX1 g75018(.A (n_7966), .Y (n_7967));
INVX1 g75041(.A (n_27991), .Y (n_7965));
OR2X1 g75049(.A (n_5068), .B (n_7563), .Y (n_7964));
INVX1 g75109(.A (n_7961), .Y (n_11687));
NAND2X1 g75167(.A (n_6336), .B (n_3301), .Y (n_7957));
NAND2X1 g75180(.A (n_7955), .B (n_28692), .Y (n_7956));
INVX1 g75182(.A (n_7953), .Y (n_7954));
NAND3X1 g75187(.A (n_9410), .B (n_4261), .C (n_28574), .Y (n_7952));
OR2X1 g75259(.A (n_5950), .B (n_7947), .Y (n_7948));
INVX1 g75274(.A (n_10393), .Y (n_7946));
INVX1 g75285(.A (n_7944), .Y (n_7945));
INVX1 g75296(.A (n_10130), .Y (n_7943));
INVX1 g75306(.A (n_7942), .Y (n_12604));
INVX1 g75325(.A (n_10610), .Y (n_7940));
INVX1 g75340(.A (n_9772), .Y (n_11772));
NAND2X1 g75367(.A (n_6941), .B (n_7938), .Y (n_7939));
INVX1 g75043(.A (n_5349), .Y (n_7937));
NAND2X1 g75392(.A (n_3984), .B (n_16198), .Y (n_7936));
INVX1 g75686(.A (n_7934), .Y (n_7935));
NAND2X1 g75491(.A (n_7932), .B (n_4898), .Y (n_7933));
INVX1 g71688(.A (n_7930), .Y (n_7931));
NOR2X1 g75503(.A (n_3502), .B (n_4416), .Y (n_7929));
INVX1 g75510(.A (n_7927), .Y (n_7928));
NOR2X1 g75624(.A (n_4079), .B (n_3030), .Y (n_7923));
NAND2X1 g75683(.A (n_2811), .B (n_8016), .Y (n_7919));
NAND2X1 g75697(.A (n_2594), .B (n_2862), .Y (n_7917));
NAND2X1 g75769(.A (n_5511), .B (n_11998), .Y (n_7912));
INVX1 g75795(.A (n_9939), .Y (n_7910));
NOR2X1 g75918(.A (n_4773), .B (n_5225), .Y (n_7906));
NAND2X1 g75928(.A (n_16934), .B (n_5509), .Y (n_7905));
NOR2X1 g75950(.A (n_5093), .B (n_6853), .Y (n_7904));
OAI21X1 g75958(.A0 (n_9500), .A1 (n_2164), .B0 (n_5441), .Y (n_7903));
INVX1 g75670(.A (n_9958), .Y (n_7902));
OR2X1 g72514(.A (n_8379), .B (n_29244), .Y (n_7900));
NOR2X1 g72016(.A (n_7899), .B (n_5333), .Y (n_9935));
XOR2X1 g76109(.A (text_in_r[15] ), .B (n_6335), .Y (n_7898));
NOR2X1 g69112(.A (n_9500), .B (n_7894), .Y (n_7895));
XOR2X1 g76139(.A (n_23234), .B (n_23418), .Y (n_7893));
XOR2X1 g76168(.A (text_in_r[17] ), .B (n_19908), .Y (n_7892));
INVX1 g70522(.A (n_7302), .Y (n_12309));
XOR2X1 g76214(.A (text_in_r[29] ), .B (n_3888), .Y (n_7889));
XOR2X1 g76220(.A (n_22564), .B (n_933), .Y (n_7888));
INVX1 g75644(.A (n_26388), .Y (n_7887));
XOR2X1 g76249(.A (text_in_r[6] ), .B (n_1142), .Y (n_7885));
XOR2X1 g76258(.A (n_23238), .B (n_23422), .Y (n_7883));
XOR2X1 g76304(.A (n_23241), .B (n_3014), .Y (n_7882));
NOR2X1 g75894(.A (n_27988), .B (n_4939), .Y (n_7881));
NOR2X1 g70506(.A (n_7879), .B (n_5924), .Y (n_10265));
INVX1 g72500(.A (n_7877), .Y (n_7878));
INVX1 g71622(.A (n_8516), .Y (n_7876));
NOR2X1 g74177(.A (n_6081), .B (n_8090), .Y (n_7875));
OR2X1 g72959(.A (n_2931), .B (n_8503), .Y (n_7874));
INVX1 g70498(.A (n_7870), .Y (n_7871));
NAND2X2 g70494(.A (n_6500), .B (n_6043), .Y (n_10268));
OR2X1 g75630(.A (n_5086), .B (n_8093), .Y (n_7868));
NOR2X1 g75315(.A (n_7742), .B (n_4300), .Y (n_9587));
AOI21X1 g73221(.A0 (n_3765), .A1 (n_4143), .B0 (n_3282), .Y (n_7865));
INVX1 g70472(.A (n_7309), .Y (n_12895));
NOR2X1 g69007(.A (n_28865), .B (n_8997), .Y (n_10635));
AND2X1 g77553(.A (n_196), .B (n_14866), .Y (n_7864));
NAND2X1 g60859(.A (n_2848), .B (n_7860), .Y (n_7862));
AND2X1 g60860(.A (n_5044), .B (n_7860), .Y (n_7859));
INVX1 g77730(.A (n_9481), .Y (n_7858));
NOR2X1 g78001(.A (n_11998), .B (n_19981), .Y (n_14266));
INVX1 g73880(.A (n_6755), .Y (n_12020));
AND2X1 g60977(.A (n_3973), .B (n_7860), .Y (n_7854));
NAND2X1 g73209(.A (n_2745), .B (n_13768), .Y (n_7853));
OAI21X1 g73207(.A0 (n_4828), .A1 (n_28574), .B0 (n_5507), .Y(n_7851));
INVX1 g75284(.A (n_7944), .Y (n_9639));
NAND3X1 g66155(.A (n_6005), .B (n_5810), .C (n_4721), .Y (n_9550));
INVX1 g77871(.A (n_7845), .Y (n_7846));
INVX1 g74908(.A (n_7844), .Y (n_7973));
NOR2X1 g67713(.A (n_5742), .B (n_9003), .Y (n_7843));
INVX1 g75275(.A (n_6342), .Y (n_10393));
INVX1 g74902(.A (n_7841), .Y (n_7974));
NAND2X2 g71562(.A (n_29142), .B (n_29225), .Y (n_16825));
NAND2X1 g70358(.A (n_3954), .B (n_8974), .Y (n_7835));
INVX1 g74445(.A (n_8015), .Y (n_9543));
NOR2X1 g75882(.A (n_3471), .B (n_4299), .Y (n_7834));
NAND2X1 g71552(.A (n_5617), .B (n_4689), .Y (n_12385));
AOI21X1 g72461(.A0 (n_3157), .A1 (n_2366), .B0 (n_2260), .Y (n_7833));
NAND2X1 g73194(.A (n_7832), .B (n_7299), .Y (n_13962));
NAND2X1 g71544(.A (n_16934), .B (n_7152), .Y (n_7831));
INVX1 g74436(.A (n_7830), .Y (n_9796));
OR2X1 g72446(.A (n_5419), .B (n_7496), .Y (n_7828));
NOR3X1 g71540(.A (n_2921), .B (n_4030), .C (n_9500), .Y (n_7826));
NAND2X2 g70323(.A (n_7824), .B (n_7496), .Y (n_10865));
NOR2X1 g73190(.A (n_2962), .B (n_11322), .Y (n_7823));
NAND2X1 g71531(.A (n_3753), .B (n_7216), .Y (n_7822));
INVX1 g74424(.A (n_8396), .Y (n_7821));
NAND2X1 g70318(.A (n_5599), .B (n_7331), .Y (n_8850));
INVX2 g74884(.A (n_5382), .Y (n_10453));
AND2X1 g70310(.A (n_5609), .B (n_7496), .Y (n_8851));
INVX1 g74879(.A (n_6310), .Y (n_7818));
INVX1 g71520(.A (n_5852), .Y (n_7816));
INVX2 g70284(.A (n_7815), .Y (n_11228));
NAND2X1 g70274(.A (n_7813), .B (n_28423), .Y (n_7814));
INVX1 g70268(.A (n_5963), .Y (n_8862));
AND2X1 g68802(.A (n_4206), .B (n_4483), .Y (n_7811));
INVX1 g74863(.A (n_9970), .Y (n_7810));
DFFX1 done_reg(.CK (clk), .D (n_4509), .Q (done), .QN ());
INVX1 g73174(.A (n_7807), .Y (n_7808));
NAND3X1 g61183(.A (n_7805), .B (n_6289), .C (n_1827), .Y (n_11608));
INVX1 g76401(.A (n_6391), .Y (n_25440));
NOR2X1 g61185(.A (n_7805), .B (n_24548), .Y (n_7806));
INVX1 g71394(.A (n_7173), .Y (n_10889));
AOI21X1 g68679(.A0 (n_7803), .A1 (n_2071), .B0 (n_5828), .Y (n_7804));
NAND2X1 g72378(.A (n_2357), .B (n_7517), .Y (n_7802));
INVX1 g74854(.A (n_8321), .Y (n_7799));
NOR2X1 g71484(.A (n_5145), .B (n_5854), .Y (n_8545));
INVX1 g71474(.A (n_7798), .Y (n_8552));
INVX1 g72992(.A (n_7797), .Y (n_8184));
INVX1 g72414(.A (n_7796), .Y (n_21820));
INVX1 g70191(.A (n_7795), .Y (n_8883));
INVX1 g74363(.A (n_8243), .Y (n_7794));
INVX2 g70180(.A (n_26550), .Y (n_11287));
NAND2X1 g78309(.A (n_28271), .B (n_8928), .Y (n_7792));
INVX1 g72770(.A (n_5730), .Y (n_8880));
INVX1 g76395(.A (n_7628), .Y (n_25335));
NOR2X1 g72399(.A (n_6825), .B (n_7789), .Y (n_8330));
NAND2X1 g72403(.A (n_12568), .B (n_3656), .Y (n_7785));
INVX1 g74833(.A (n_7782), .Y (n_7784));
NAND2X1 g75373(.A (n_2612), .B (n_9416), .Y (n_7783));
INVX1 g74832(.A (n_7782), .Y (n_10272));
NAND2X1 g70142(.A (n_6582), .B (n_4300), .Y (n_8892));
AND2X1 g71425(.A (n_1929), .B (n_7777), .Y (n_11386));
NOR2X1 g74801(.A (n_4682), .B (n_28381), .Y (n_7776));
XOR2X1 g76297(.A (n_2560), .B (n_6352), .Y (n_7775));
NAND2X2 g73004(.A (n_26878), .B (n_9783), .Y (n_15534));
NAND3X1 g67459(.A (n_7770), .B (n_2886), .C (n_5823), .Y (n_7771));
INVX1 g75206(.A (n_7769), .Y (n_7950));
NAND3X1 g65992(.A (n_8968), .B (n_27367), .C (n_4261), .Y (n_28986));
NAND2X1 g70090(.A (n_5258), .B (n_7496), .Y (n_10957));
INVX1 g75688(.A (n_7767), .Y (n_7934));
OR4X1 g66001(.A (n_29269), .B (n_2487), .C (n_29153), .D (n_3562), .Y(n_13316));
INVX1 g75201(.A (n_6218), .Y (n_9502));
INVX1 g74304(.A (n_7763), .Y (n_29115));
OR4X1 g66040(.A (n_12169), .B (n_3920), .C (n_3038), .D (n_4501), .Y(n_15243));
AND2X1 g66074(.A (n_7759), .B (n_11354), .Y (n_11424));
NAND4X1 g66075(.A (n_2779), .B (n_379), .C (n_827), .D (n_2530), .Y(n_17266));
INVX1 g74730(.A (n_7757), .Y (n_7758));
INVX1 g74268(.A (n_7755), .Y (n_7756));
OR4X1 g66082(.A (n_1376), .B (n_4882), .C (n_2492), .D (n_5404), .Y(n_13537));
NAND4X1 g66084(.A (n_12169), .B (n_3301), .C (n_3038), .D (n_2541),.Y (n_18343));
NOR2X1 g74292(.A (n_4028), .B (n_4568), .Y (n_7753));
NAND4X1 g66111(.A (n_14866), .B (n_5151), .C (n_2492), .D (n_2583),.Y (n_16564));
NAND4X1 g66112(.A (n_17912), .B (n_13490), .C (n_2968), .D (n_29120),.Y (n_15642));
NAND2X1 g72375(.A (n_6958), .B (n_26883), .Y (n_8335));
NAND4X1 g70078(.A (n_7543), .B (n_7438), .C (n_28271), .D (n_4391),.Y (n_7748));
AND2X1 g66127(.A (n_5819), .B (n_12760), .Y (n_11439));
INVX2 g74294(.A (n_7746), .Y (n_7745));
NAND2X1 g66131(.A (n_7744), .B (n_12169), .Y (n_11507));
INVX1 g75568(.A (n_8346), .Y (n_10212));
INVX1 g77731(.A (n_7742), .Y (n_9481));
NAND4X1 g66195(.A (n_27099), .B (n_7266), .C (n_28575), .D (n_5546),.Y (n_7741));
AND2X1 g75560(.A (n_2883), .B (n_2318), .Y (n_7739));
NAND2X1 g73115(.A (n_6838), .B (n_7182), .Y (n_9456));
NAND4X1 g66298(.A (n_14624), .B (n_4721), .C (n_1186), .D (n_4920),.Y (n_15499));
NOR2X1 g66304(.A (n_28996), .B (n_7593), .Y (n_9446));
NAND4X1 g66314(.A (n_10389), .B (n_7947), .C (n_7734), .D (n_2705),.Y (n_13421));
INVX1 g70063(.A (n_6205), .Y (n_8907));
OR2X1 g66317(.A (n_7733), .B (n_16466), .Y (n_17527));
NOR2X1 g66339(.A (n_7732), .B (n_26491), .Y (n_9440));
OR2X1 g73109(.A (n_3931), .B (n_8679), .Y (n_11383));
INVX1 g71382(.A (n_5861), .Y (n_11006));
NOR2X1 g75183(.A (n_7730), .B (n_6790), .Y (n_7953));
NAND2X1 g70052(.A (n_27227), .B (n_636), .Y (n_8908));
NAND4X1 g66376(.A (n_9942), .B (n_7728), .C (n_28362), .D (n_5985),.Y (n_16768));
NAND2X1 g67397(.A (n_5972), .B (n_16480), .Y (n_7727));
OR2X1 g66381(.A (n_7726), .B (n_9003), .Y (n_14770));
OR4X1 g66386(.A (n_9819), .B (n_6790), .C (n_7725), .D (n_3805), .Y(n_11452));
INVX1 g71354(.A (n_7723), .Y (n_7724));
NAND2X1 g66449(.A (n_6074), .B (n_1147), .Y (n_9559));
INVX1 g74266(.A (n_7722), .Y (n_10333));
NOR2X1 g71374(.A (n_4437), .B (n_13490), .Y (n_13341));
NAND2X1 g70041(.A (n_5749), .B (n_8263), .Y (n_10921));
NAND2X1 g75876(.A (n_7721), .B (n_6656), .Y (n_9419));
INVX1 g71092(.A (n_7719), .Y (n_8658));
NOR2X1 g66509(.A (n_7717), .B (n_12979), .Y (n_7718));
INVX1 g75172(.A (n_5319), .Y (n_9424));
NAND3X1 g66563(.A (n_4861), .B (n_6265), .C (n_4825), .Y (n_11456));
NAND4X1 g66580(.A (n_9486), .B (n_5854), .C (n_3445), .D (n_4326), .Y(n_7714));
INVX1 g61523(.A (n_6184), .Y (n_7713));
NAND2X1 g74249(.A (n_11669), .B (n_3445), .Y (n_7712));
NOR2X1 g66645(.A (n_7710), .B (n_15166), .Y (n_7711));
INVX1 g73458(.A (n_5661), .Y (n_8083));
NAND4X1 g66700(.A (n_6005), .B (n_7607), .C (n_1186), .D (n_2329), .Y(n_11447));
INVX1 g73080(.A (n_7709), .Y (n_11367));
OR2X1 g66767(.A (n_7708), .B (n_3318), .Y (n_15675));
NAND4X1 g66784(.A (n_29225), .B (n_27990), .C (n_29163), .D (n_4115),.Y (n_15543));
INVX4 g74236(.A (n_7705), .Y (n_9838));
OR2X1 g74732(.A (n_8706), .B (n_7701), .Y (n_7702));
OR2X1 g73639(.A (n_4158), .B (n_18440), .Y (n_7700));
NOR2X1 g66886(.A (n_5928), .B (n_8968), .Y (n_9366));
INVX1 g73064(.A (n_6162), .Y (n_9365));
NAND2X1 g72193(.A (n_7069), .B (n_28398), .Y (n_15186));
NOR2X1 g73048(.A (n_6131), .B (n_18266), .Y (n_7696));
NAND2X1 g72324(.A (n_7131), .B (n_11739), .Y (n_7694));
NAND2X1 g73052(.A (n_14548), .B (n_5310), .Y (n_8164));
NOR2X1 g67037(.A (n_5767), .B (n_6005), .Y (n_9346));
NAND2X1 g72322(.A (n_6871), .B (n_7659), .Y (n_12673));
NAND2X1 g67070(.A (n_7661), .B (n_14142), .Y (n_14868));
AOI21X1 g67271(.A0 (n_4899), .A1 (n_5692), .B0 (n_14592), .Y(n_7690));
OR2X1 g71338(.A (n_14348), .B (n_4314), .Y (n_7688));
NAND3X1 g67144(.A (n_7686), .B (n_7685), .C (n_5694), .Y (n_7687));
NAND2X2 g67150(.A (n_6084), .B (n_12169), .Y (n_29208));
NOR2X1 g73038(.A (n_7631), .B (n_7362), .Y (n_7682));
OR2X1 g73032(.A (n_7526), .B (n_2318), .Y (n_8170));
INVX1 g73605(.A (n_7679), .Y (n_7680));
AND2X1 g69962(.A (n_7678), .B (n_3736), .Y (n_11530));
INVX2 g69948(.A (n_6140), .Y (n_11200));
NOR2X1 g74722(.A (n_7675), .B (n_11731), .Y (n_7676));
NAND2X1 g67276(.A (n_6093), .B (n_5306), .Y (n_7674));
NAND2X1 g67311(.A (n_7672), .B (n_6134), .Y (n_7673));
AOI21X1 g67318(.A0 (n_4297), .A1 (n_5705), .B0 (n_14624), .Y(n_7671));
NAND2X1 g67386(.A (n_7665), .B (n_5817), .Y (n_9305));
OR2X1 g73010(.A (n_4275), .B (n_6968), .Y (n_7667));
INVX1 g73585(.A (n_8810), .Y (n_9962));
AND2X1 g67454(.A (n_7665), .B (n_8217), .Y (n_7666));
INVX1 g73581(.A (n_8810), .Y (n_7664));
NAND2X1 g72280(.A (n_379), .B (n_2632), .Y (n_11087));
INVX1 g73000(.A (n_5709), .Y (n_10734));
OR2X1 g72276(.A (n_5399), .B (n_17912), .Y (n_7663));
NAND2X1 g72268(.A (n_6332), .B (n_4391), .Y (n_7662));
NOR2X1 g67628(.A (n_14337), .B (n_9257), .Y (n_9538));
INVX1 g74641(.A (n_5722), .Y (n_8197));
NOR2X1 g67682(.A (n_6082), .B (n_2260), .Y (n_9279));
NAND2X1 g67686(.A (n_7661), .B (n_8878), .Y (n_16963));
AND2X1 g69901(.A (n_7659), .B (n_7658), .Y (n_8939));
INVX2 g72698(.A (n_5734), .Y (n_8251));
NAND2X1 g72976(.A (n_5567), .B (n_14484), .Y (n_13301));
NOR2X1 g67741(.A (n_5700), .B (n_8637), .Y (n_7656));
INVX1 g69888(.A (n_5984), .Y (n_8941));
NAND2X1 g67759(.A (n_6128), .B (n_5799), .Y (n_18598));
NAND2X1 g74184(.A (n_6730), .B (n_5660), .Y (n_8022));
NOR2X1 g67877(.A (n_5866), .B (n_28445), .Y (n_7653));
INVX1 g73524(.A (n_7650), .Y (n_10546));
NAND2X1 g68021(.A (n_6249), .B (n_10100), .Y (n_13324));
NAND4X1 g68028(.A (n_7649), .B (n_5924), .C (n_2968), .D (n_28340),.Y (n_9242));
NAND2X1 g68046(.A (n_5689), .B (n_10452), .Y (n_7645));
NAND2X1 g68060(.A (n_5686), .B (n_10100), .Y (n_15556));
AND2X1 g68074(.A (n_7639), .B (n_1512), .Y (n_7644));
NAND2X1 g74168(.A (n_2742), .B (n_3723), .Y (n_7642));
INVX1 g74162(.A (n_7641), .Y (n_10083));
NAND3X1 g68173(.A (n_6344), .B (n_2923), .C (n_4638), .Y (n_7640));
NAND2X1 g68176(.A (n_7639), .B (n_11307), .Y (n_13482));
OR2X1 g68190(.A (n_5805), .B (n_13466), .Y (n_11416));
NAND2X1 g73496(.A (n_5403), .B (n_7636), .Y (n_7637));
NAND2X1 g72925(.A (n_7123), .B (n_9500), .Y (n_7635));
INVX1 g69830(.A (n_5986), .Y (n_10956));
NOR2X1 g68266(.A (n_7634), .B (n_11731), .Y (n_8700));
NOR2X1 g72220(.A (n_2322), .B (n_6031), .Y (n_8377));
NAND2X1 g68280(.A (n_6104), .B (n_14866), .Y (n_9214));
NOR2X1 g71246(.A (n_2318), .B (n_7631), .Y (n_7632));
NAND2X2 g69814(.A (n_5427), .B (n_28402), .Y (n_10909));
INVX1 g68411(.A (n_17139), .Y (n_7630));
INVX1 g76406(.A (n_8696), .Y (n_25353));
NOR2X1 g66945(.A (n_5715), .B (n_11322), .Y (n_7629));
INVX1 g76394(.A (n_7628), .Y (n_25426));
NAND2X1 g68507(.A (n_3927), .B (n_7625), .Y (n_7626));
NOR2X1 g66927(.A (n_7624), .B (n_6219), .Y (n_9354));
INVX1 g69784(.A (n_9402), .Y (n_8959));
NOR2X1 g72896(.A (n_5357), .B (n_29269), .Y (n_7623));
INVX1 g74144(.A (n_7619), .Y (n_7620));
AOI21X1 g68692(.A0 (n_5778), .A1 (n_3726), .B0 (n_7617), .Y (n_7618));
INVX1 g72181(.A (n_6197), .Y (n_9176));
INVX2 g69760(.A (n_5994), .Y (n_11495));
INVX1 g72876(.A (n_5711), .Y (n_11114));
OR2X1 g72872(.A (n_7615), .B (n_7614), .Y (n_7616));
NAND2X1 g72870(.A (n_9899), .B (n_7440), .Y (n_15137));
NAND2X2 g71194(.A (n_7210), .B (n_4261), .Y (n_9167));
OAI21X1 g68778(.A0 (n_14734), .A1 (n_5845), .B0 (n_2386), .Y(n_7609));
INVX1 g72158(.A (n_7020), .Y (n_7608));
NAND2X1 g69737(.A (n_5227), .B (n_7607), .Y (n_10835));
NAND2X1 g71188(.A (n_3167), .B (n_6939), .Y (n_15949));
XOR2X1 g68812(.A (n_3184), .B (n_1221), .Y (n_9156));
NOR2X1 g72155(.A (n_5257), .B (n_2810), .Y (n_7606));
NAND2X1 g72851(.A (n_7101), .B (n_7678), .Y (n_7605));
NAND2X1 g72849(.A (n_6974), .B (n_8742), .Y (n_15315));
INVX1 g72146(.A (n_7602), .Y (n_10913));
INVX1 g72141(.A (n_6080), .Y (n_14425));
NAND2X2 g68972(.A (n_6243), .B (n_7601), .Y (n_11165));
INVX1 g68978(.A (n_7600), .Y (n_9144));
INVX2 g68986(.A (n_6078), .Y (n_9143));
AND2X1 g68989(.A (n_4122), .B (n_7598), .Y (n_7599));
NOR2X1 g68998(.A (n_27594), .B (n_7496), .Y (n_9140));
INVX1 g69009(.A (n_6077), .Y (n_7597));
CLKBUFX3 g69021(.A (n_6076), .Y (n_13607));
NAND2X1 g69030(.A (n_29330), .B (n_5413), .Y (n_7596));
NOR2X1 g69035(.A (n_7549), .B (n_14055), .Y (n_9132));
INVX1 g72838(.A (n_6916), .Y (n_7595));
INVX1 g69045(.A (n_5066), .Y (n_11292));
INVX1 g69050(.A (n_15085), .Y (n_11197));
AND2X1 g69052(.A (n_6256), .B (n_7593), .Y (n_7594));
INVX2 g69055(.A (n_7592), .Y (n_13190));
NAND2X2 g69066(.A (n_5975), .B (n_7512), .Y (n_9124));
INVX2 g69070(.A (n_7591), .Y (n_10968));
INVX2 g73370(.A (n_7800), .Y (n_10125));
OR2X1 g69080(.A (n_7420), .B (n_9084), .Y (n_7590));
INVX1 g69083(.A (n_9418), .Y (n_10691));
NAND2X1 g69089(.A (n_5278), .B (n_7563), .Y (n_9116));
INVX1 g69091(.A (n_9344), .Y (n_18115));
INVX1 g69097(.A (n_6072), .Y (n_9115));
INVX1 g69100(.A (n_6069), .Y (n_9114));
NAND2X1 g69103(.A (n_4567), .B (n_7607), .Y (n_13217));
NAND4X1 g69105(.A (n_9118), .B (n_3069), .C (n_7586), .D (n_2960), .Y(n_9111));
INVX1 g69106(.A (n_7585), .Y (n_11190));
NOR2X1 g71248(.A (n_3138), .B (n_7583), .Y (n_7584));
NAND2X2 g69121(.A (n_5595), .B (n_16198), .Y (n_9108));
NAND2X2 g69146(.A (n_6339), .B (n_4934), .Y (n_14521));
NAND2X1 g69154(.A (n_7578), .B (n_11835), .Y (n_14014));
NAND2X1 g69157(.A (n_7480), .B (n_3807), .Y (n_10701));
NAND2X2 g69161(.A (n_3250), .B (n_4173), .Y (n_11029));
NAND2X1 g69162(.A (n_7576), .B (n_7410), .Y (n_7577));
NAND2X1 g69168(.A (n_7659), .B (n_7537), .Y (n_7574));
INVX1 g69172(.A (n_6064), .Y (n_11233));
INVX1 g69178(.A (n_7572), .Y (n_7573));
NOR2X1 g72120(.A (n_7568), .B (n_7567), .Y (n_7569));
INVX1 g69197(.A (n_7566), .Y (n_9099));
NOR2X1 g69204(.A (n_5576), .B (n_7563), .Y (n_7565));
NAND4X1 g69209(.A (n_367), .B (n_7563), .C (n_3696), .D (n_2960), .Y(n_7564));
INVX1 g69216(.A (n_10943), .Y (n_13211));
NAND2X1 g69227(.A (n_29333), .B (n_7559), .Y (n_9095));
INVX1 g69231(.A (n_7557), .Y (n_7558));
INVX1 g69237(.A (n_6057), .Y (n_9093));
INVX1 g69239(.A (n_9573), .Y (n_7556));
CLKBUFX1 g69243(.A (n_14208), .Y (n_17130));
INVX1 g69251(.A (n_7555), .Y (n_9088));
INVX1 g72822(.A (n_7554), .Y (n_17297));
NAND2X2 g69257(.A (n_7553), .B (n_28445), .Y (n_11122));
INVX1 g69259(.A (n_5423), .Y (n_11334));
INVX1 g69264(.A (n_6053), .Y (n_9085));
INVX1 g69269(.A (n_7551), .Y (n_7552));
NOR2X1 g69711(.A (n_7549), .B (n_14155), .Y (n_7550));
INVX1 g69277(.A (n_7548), .Y (n_8003));
INVX1 g69286(.A (n_7547), .Y (n_10789));
INVX1 g69288(.A (n_19030), .Y (n_7546));
NAND2X1 g69290(.A (n_7535), .B (n_8708), .Y (n_7545));
INVX1 g69296(.A (n_6048), .Y (n_10971));
INVX1 g69302(.A (n_6047), .Y (n_9075));
INVX1 g69306(.A (n_9404), .Y (n_10687));
INVX1 g69315(.A (n_5527), .Y (n_9071));
NAND4X1 g69320(.A (n_7543), .B (n_28364), .C (n_28271), .D (n_6988),.Y (n_7544));
INVX1 g69323(.A (n_9281), .Y (n_13487));
AND2X1 g69326(.A (n_5757), .B (n_10389), .Y (n_7542));
AND2X1 g69327(.A (n_5208), .B (n_6007), .Y (n_7541));
AND2X1 g69330(.A (n_6111), .B (n_29297), .Y (n_7540));
INVX1 g69334(.A (n_6044), .Y (n_11381));
NAND2X1 g69339(.A (n_4868), .B (n_7537), .Y (n_14493));
NAND2X1 g69340(.A (n_7535), .B (n_5854), .Y (n_7536));
NAND2X1 g69341(.A (n_5326), .B (n_14866), .Y (n_7534));
NAND2X1 g69343(.A (n_6960), .B (n_7182), .Y (n_11516));
NOR2X1 g69346(.A (n_28615), .B (n_6534), .Y (n_9066));
INVX1 g69349(.A (n_6042), .Y (n_9064));
INVX1 g69355(.A (n_7532), .Y (n_11099));
INVX1 g69361(.A (n_7531), .Y (n_13082));
NAND2X1 g69365(.A (n_5610), .B (n_29221), .Y (n_7529));
NOR2X1 g69368(.A (n_6151), .B (n_8865), .Y (n_9060));
AND2X1 g69375(.A (n_5363), .B (n_12019), .Y (n_7528));
NOR2X1 g72818(.A (n_7526), .B (n_11261), .Y (n_7527));
NAND2X2 g69381(.A (n_5644), .B (n_29297), .Y (n_14009));
NAND2X1 g69383(.A (n_7487), .B (n_16434), .Y (n_7524));
NOR2X1 g72814(.A (n_5298), .B (n_11323), .Y (n_7523));
NOR2X1 g74646(.A (n_4745), .B (n_7563), .Y (n_7995));
NAND2X1 g69391(.A (n_5613), .B (n_6191), .Y (n_7522));
INVX2 g69395(.A (n_5690), .Y (n_14872));
INVX1 g69397(.A (n_7521), .Y (n_11249));
INVX1 g69401(.A (n_6036), .Y (n_12306));
NAND2X1 g69404(.A (n_4665), .B (n_11731), .Y (n_7520));
INVX1 g69406(.A (n_6035), .Y (n_7519));
INVX1 g69415(.A (n_6880), .Y (n_13320));
NAND2X1 g69422(.A (n_4994), .B (n_6534), .Y (n_9048));
NAND2X1 g69425(.A (n_6217), .B (n_2318), .Y (n_11133));
NAND2X1 g69427(.A (n_7517), .B (n_12169), .Y (n_7518));
NAND2X1 g69436(.A (n_5202), .B (n_8945), .Y (n_9043));
NAND2X1 g69437(.A (n_3706), .B (n_4565), .Y (n_7513));
INVX1 g69441(.A (n_5731), .Y (n_10747));
INVX1 g69445(.A (n_17725), .Y (n_9041));
NAND2X1 g69453(.A (n_7503), .B (n_7512), .Y (n_9040));
OR2X1 g69454(.A (n_4599), .B (n_9388), .Y (n_11550));
INVX1 g69457(.A (n_7509), .Y (n_7511));
INVX1 g69477(.A (n_5755), .Y (n_9034));
INVX1 g69482(.A (n_6026), .Y (n_9033));
INVX1 g69487(.A (n_6024), .Y (n_11321));
INVX1 g69490(.A (n_10937), .Y (n_7506));
INVX1 g69500(.A (n_7504), .Y (n_11543));
INVX1 g69505(.A (n_6022), .Y (n_11235));
NAND2X1 g69508(.A (n_7503), .B (n_27371), .Y (n_11473));
NAND2X1 g69514(.A (n_7517), .B (n_3920), .Y (n_14510));
INVX1 g69517(.A (n_6020), .Y (n_11263));
INVX2 g69520(.A (n_7499), .Y (n_15640));
NOR2X1 g71128(.A (n_5230), .B (n_7498), .Y (n_8645));
AND2X1 g69530(.A (n_5437), .B (n_7496), .Y (n_7497));
AND2X1 g69531(.A (n_5347), .B (n_5854), .Y (n_7495));
AND2X1 g69552(.A (n_5206), .B (n_11323), .Y (n_7492));
AND2X1 g69555(.A (n_5747), .B (n_3318), .Y (n_7490));
INVX1 g69564(.A (n_7489), .Y (n_10888));
NAND2X1 g69568(.A (n_7487), .B (n_13593), .Y (n_7488));
NAND2X2 g71125(.A (n_7486), .B (n_7485), .Y (n_9006));
INVX1 g69576(.A (n_14126), .Y (n_11017));
NOR2X1 g69581(.A (n_5481), .B (n_17912), .Y (n_13458));
NAND2X1 g73074(.A (n_6419), .B (n_2803), .Y (n_10850));
INVX1 g69593(.A (n_5926), .Y (n_12451));
INVX1 g69597(.A (n_6009), .Y (n_10964));
INVX1 g69600(.A (n_7482), .Y (n_7483));
INVX2 g69607(.A (n_7481), .Y (n_9000));
NAND2X1 g69617(.A (n_7480), .B (n_7331), .Y (n_8784));
NAND2X1 g69625(.A (n_7479), .B (n_8452), .Y (n_11080));
OR2X1 g69627(.A (n_7477), .B (n_9264), .Y (n_7478));
NOR3X1 g72088(.A (n_27133), .B (n_4015), .C (n_27124), .Y (n_7476));
INVX2 g69653(.A (n_5982), .Y (n_8922));
NAND2X1 g69655(.A (n_7317), .B (n_11300), .Y (n_7472));
NAND2X1 g69658(.A (n_4480), .B (n_8997), .Y (n_7471));
INVX1 g69668(.A (n_7470), .Y (n_8992));
NAND2X1 g69672(.A (n_6183), .B (n_8945), .Y (n_7469));
NOR2X1 g69675(.A (n_4778), .B (n_7777), .Y (n_10838));
INVX1 g69677(.A (n_6001), .Y (n_12628));
INVX1 g69680(.A (n_7466), .Y (n_7467));
NOR2X1 g69696(.A (n_4592), .B (n_7598), .Y (n_8983));
INVX1 g69701(.A (n_17288), .Y (n_7464));
NAND2X1 g69712(.A (n_12731), .B (n_7410), .Y (n_7463));
NAND2X1 g69716(.A (n_27612), .B (n_11322), .Y (n_7461));
NAND2X1 g69719(.A (n_6209), .B (n_5413), .Y (n_11043));
NAND2X1 g69722(.A (n_4277), .B (n_26491), .Y (n_7459));
NAND2X1 g69724(.A (n_7350), .B (n_11835), .Y (n_7458));
NAND2X1 g69731(.A (n_4420), .B (n_7496), .Y (n_7457));
NAND2X1 g69732(.A (n_4607), .B (n_26491), .Y (n_7456));
NAND2X1 g69740(.A (n_13655), .B (n_7593), .Y (n_7455));
AND2X1 g69741(.A (n_5499), .B (n_8997), .Y (n_7454));
NOR2X1 g72798(.A (n_7453), .B (n_5481), .Y (n_8223));
AND2X1 g69746(.A (n_3997), .B (n_3599), .Y (n_8970));
NAND2X2 g69753(.A (n_6229), .B (n_5483), .Y (n_16416));
OR2X1 g69770(.A (n_7452), .B (n_379), .Y (n_15659));
NAND2X1 g69772(.A (n_4397), .B (n_7325), .Y (n_10915));
INVX1 g69776(.A (n_7450), .Y (n_10996));
INVX1 g69779(.A (n_7447), .Y (n_7448));
NAND2X1 g69789(.A (n_7678), .B (n_11307), .Y (n_7446));
NAND2X1 g69801(.A (n_5215), .B (n_5922), .Y (n_9208));
AND2X1 g69802(.A (n_5360), .B (n_27365), .Y (n_7443));
NAND2X2 g69806(.A (n_5816), .B (n_8339), .Y (n_10799));
NAND2X1 g69818(.A (n_5222), .B (n_6462), .Y (n_29176));
CLKBUFX3 g69825(.A (n_5989), .Y (n_11020));
NAND2X1 g69828(.A (n_4377), .B (n_4248), .Y (n_7441));
NAND2X2 g69841(.A (n_7440), .B (n_10031), .Y (n_9227));
NAND2X1 g69847(.A (n_8024), .B (n_7438), .Y (n_14407));
NAND2X1 g69851(.A (n_5349), .B (n_7127), .Y (n_7437));
INVX1 g69861(.A (n_6443), .Y (n_7436));
NAND2X1 g69864(.A (n_5487), .B (n_8974), .Y (n_11462));
INVX1 g69871(.A (n_6119), .Y (n_8944));
NOR2X1 g69874(.A (n_6415), .B (n_27688), .Y (n_8943));
AND2X1 g69875(.A (n_5552), .B (n_8974), .Y (n_7434));
NAND2X1 g69883(.A (n_5352), .B (n_6185), .Y (n_7433));
INVX1 g71978(.A (n_5806), .Y (n_8428));
INVX1 g69893(.A (n_7432), .Y (n_14330));
INVX1 g74686(.A (n_7429), .Y (n_10177));
INVX1 g71104(.A (n_27712), .Y (n_7428));
NAND2X1 g69906(.A (n_7403), .B (n_9819), .Y (n_7427));
INVX1 g69922(.A (n_7422), .Y (n_10987));
INVX2 g69931(.A (n_6138), .Y (n_8937));
CLKBUFX2 g69936(.A (n_7421), .Y (n_14340));
OR2X1 g69950(.A (n_7420), .B (n_17104), .Y (n_17752));
NAND2X2 g69955(.A (n_6206), .B (n_7419), .Y (n_10945));
NOR2X1 g71098(.A (n_7418), .B (n_4214), .Y (n_8654));
OR2X1 g69975(.A (n_7417), .B (n_3301), .Y (n_8929));
INVX1 g69991(.A (n_9380), .Y (n_8924));
INVX1 g72058(.A (n_7416), .Y (n_8414));
OR2X1 g72780(.A (n_7415), .B (n_9388), .Y (n_8902));
INVX1 g70004(.A (n_7703), .Y (n_7414));
INVX1 g70011(.A (n_6173), .Y (n_11365));
NAND2X2 g70013(.A (n_5670), .B (n_9335), .Y (n_11492));
AOI21X1 g70014(.A0 (n_3783), .A1 (n_7411), .B0 (n_1668), .Y (n_7412));
OR2X1 g70046(.A (n_4292), .B (n_7410), .Y (n_17303));
INVX1 g70068(.A (n_7408), .Y (n_7409));
OR2X1 g70070(.A (n_7406), .B (n_28433), .Y (n_7407));
NAND2X1 g70080(.A (n_5411), .B (n_6977), .Y (n_10900));
INVX1 g70085(.A (n_5973), .Y (n_8898));
NAND2X1 g70092(.A (n_4870), .B (n_15776), .Y (n_18691));
NAND2X1 g70097(.A (n_7403), .B (n_9264), .Y (n_7404));
INVX1 g70104(.A (n_9349), .Y (n_7399));
INVX1 g70115(.A (n_14046), .Y (n_7394));
OR2X1 g70119(.A (n_27432), .B (n_9368), .Y (n_7393));
NAND2X1 g70120(.A (n_7370), .B (n_11400), .Y (n_7391));
INVX1 g70127(.A (n_7390), .Y (n_8897));
NAND2X1 g68311(.A (n_7388), .B (n_6005), .Y (n_7389));
INVX1 g70149(.A (n_27710), .Y (n_7386));
INVX1 g70153(.A (n_6248), .Y (n_7385));
NAND2X1 g70157(.A (n_7358), .B (n_9783), .Y (n_7384));
NAND2X1 g70158(.A (n_4221), .B (n_7201), .Y (n_7383));
AND2X1 g70163(.A (n_5406), .B (n_28375), .Y (n_7382));
INVX1 g70170(.A (n_7381), .Y (n_8887));
NAND2X1 g70194(.A (n_6342), .B (n_6279), .Y (n_10986));
INVX1 g72045(.A (n_6274), .Y (n_13195));
AND2X1 g70198(.A (n_4293), .B (n_9118), .Y (n_7380));
INVX1 g70200(.A (n_7377), .Y (n_7378));
OR2X1 g70204(.A (n_4001), .B (n_11312), .Y (n_17250));
NAND2X1 g70208(.A (n_6930), .B (n_27990), .Y (n_11175));
NOR2X1 g70211(.A (n_7376), .B (n_6462), .Y (n_8876));
NAND2X1 g70216(.A (n_6920), .B (n_12979), .Y (n_7372));
NAND2X1 g70217(.A (n_7370), .B (n_28444), .Y (n_7371));
CLKBUFX3 g70222(.A (n_5967), .Y (n_16590));
AND2X1 g70224(.A (n_6270), .B (n_14866), .Y (n_7369));
NAND2X1 g69639(.A (n_7367), .B (n_7366), .Y (n_7368));
INVX1 g70234(.A (n_12560), .Y (n_8870));
AND2X1 g70237(.A (n_5882), .B (n_29225), .Y (n_7365));
NAND2X1 g70247(.A (n_6223), .B (n_7362), .Y (n_7363));
NAND2X1 g70249(.A (n_4757), .B (n_15776), .Y (n_8867));
NAND2X1 g70258(.A (n_7041), .B (n_13326), .Y (n_17127));
NAND2X1 g70263(.A (n_7358), .B (n_15411), .Y (n_7359));
NAND2X2 g70276(.A (n_7357), .B (n_5854), .Y (n_10817));
OR2X1 g70278(.A (n_4461), .B (n_12169), .Y (n_8859));
INVX1 g70279(.A (n_7355), .Y (n_13521));
INVX1 g72344(.A (n_7354), .Y (n_8351));
INVX1 g69632(.A (n_6003), .Y (n_8995));
INVX1 g70286(.A (n_7352), .Y (n_7353));
NAND2X1 g70288(.A (n_7350), .B (n_16787), .Y (n_7351));
AND2X1 g70291(.A (n_5280), .B (n_7512), .Y (n_7349));
AND2X1 g70292(.A (n_5301), .B (n_27434), .Y (n_7348));
INVX1 g70294(.A (n_7347), .Y (n_8857));
NAND2X1 g70296(.A (n_4371), .B (n_10100), .Y (n_7346));
NAND2X1 g70297(.A (n_4977), .B (n_4689), .Y (n_7345));
INVX1 g70299(.A (n_7343), .Y (n_7344));
INVX1 g70307(.A (n_9322), .Y (n_16959));
NAND2X1 g70319(.A (n_4272), .B (n_16198), .Y (n_7340));
NAND2X1 g70321(.A (n_5038), .B (n_4848), .Y (n_11053));
INVX1 g70325(.A (n_7337), .Y (n_7339));
NAND2X1 g70330(.A (n_4359), .B (n_9417), .Y (n_7336));
NAND2X1 g70333(.A (n_7567), .B (n_11307), .Y (n_10795));
INVX1 g73358(.A (n_9053), .Y (n_7334));
INVX1 g70348(.A (n_7333), .Y (n_11290));
AND2X1 g70350(.A (n_5460), .B (n_7331), .Y (n_7332));
NAND2X1 g70353(.A (n_7329), .B (n_14026), .Y (n_7330));
NOR2X1 g70356(.A (n_4394), .B (n_14055), .Y (n_8839));
NOR2X1 g72760(.A (n_4141), .B (n_28686), .Y (n_7328));
AND2X1 g70360(.A (n_6155), .B (n_4709), .Y (n_7327));
OR2X1 g70361(.A (n_4666), .B (n_9637), .Y (n_7326));
NAND2X1 g70362(.A (n_4279), .B (n_7325), .Y (n_12631));
INVX1 g70364(.A (n_7322), .Y (n_7324));
INVX1 g70385(.A (n_7976), .Y (n_11517));
NAND2X1 g70389(.A (n_7321), .B (n_7485), .Y (n_8833));
OR2X1 g70390(.A (n_7319), .B (n_11261), .Y (n_7320));
NAND2X1 g70391(.A (n_7317), .B (n_29286), .Y (n_7318));
NAND2X1 g70397(.A (n_6010), .B (n_8452), .Y (n_7316));
INVX1 g70400(.A (n_7315), .Y (n_11338));
OR2X1 g70411(.A (n_3372), .B (n_11312), .Y (n_8827));
INVX1 g70413(.A (n_4983), .Y (n_10919));
NAND2X1 g70428(.A (n_11413), .B (n_11307), .Y (n_8822));
INVX2 g70438(.A (n_7312), .Y (n_11193));
INVX2 g70446(.A (n_5945), .Y (n_10782));
NAND2X1 g71068(.A (n_7238), .B (n_2655), .Y (n_8670));
INVX1 g70460(.A (n_5943), .Y (n_13697));
AND2X1 g70463(.A (n_5240), .B (n_8997), .Y (n_7310));
INVX1 g70467(.A (n_5941), .Y (n_10724));
NAND3X1 g70473(.A (n_490), .B (n_2743), .C (n_827), .Y (n_7309));
NAND2X1 g70476(.A (n_4129), .B (n_9057), .Y (n_12751));
NAND2X2 g70481(.A (n_6295), .B (n_6043), .Y (n_8814));
NOR2X1 g70490(.A (n_5214), .B (n_4522), .Y (n_7308));
NAND4X1 g70495(.A (n_15894), .B (n_488), .C (n_2319), .D (n_1750), .Y(n_14930));
NAND2X1 g70499(.A (n_5560), .B (n_6219), .Y (n_7870));
INVX1 g70500(.A (n_7307), .Y (n_11387));
NAND2X1 g70508(.A (n_5648), .B (n_27757), .Y (n_7306));
INVX1 g70509(.A (n_7303), .Y (n_7305));
NOR2X1 g70523(.A (n_28725), .B (n_29297), .Y (n_7302));
NAND2X2 g70533(.A (n_6102), .B (n_7201), .Y (n_8805));
NAND2X1 g70539(.A (n_27076), .B (n_6055), .Y (n_7301));
NAND2X1 g70548(.A (n_7299), .B (n_3920), .Y (n_14512));
NAND2X1 g70549(.A (n_4905), .B (n_10452), .Y (n_7298));
INVX1 g70565(.A (n_5934), .Y (n_11118));
NAND2X1 g70571(.A (n_6308), .B (n_11322), .Y (n_7297));
OR2X1 g70577(.A (n_7296), .B (n_13490), .Y (n_8799));
OR2X1 g72740(.A (n_7292), .B (n_12849), .Y (n_7293));
NOR2X1 g70596(.A (n_7290), .B (n_16414), .Y (n_7291));
NAND2X2 g70605(.A (n_7288), .B (n_28418), .Y (n_10820));
INVX1 g70608(.A (n_9406), .Y (n_12303));
NAND2X1 g70613(.A (n_5580), .B (n_1147), .Y (n_7286));
INVX1 g70618(.A (n_7283), .Y (n_10846));
INVX1 g72012(.A (n_9531), .Y (n_7282));
NOR2X1 g70650(.A (n_4546), .B (n_28733), .Y (n_8775));
NAND2X1 g70651(.A (n_12268), .B (n_28132), .Y (n_11285));
NAND2X2 g70679(.A (n_28163), .B (n_6185), .Y (n_8768));
NOR2X1 g70712(.A (n_5443), .B (n_11312), .Y (n_11061));
NOR2X1 g70714(.A (n_4372), .B (n_6961), .Y (n_7276));
INVX1 g70719(.A (n_5470), .Y (n_8009));
NOR2X1 g70722(.A (n_4984), .B (n_10452), .Y (n_7275));
NAND2X1 g70724(.A (n_5025), .B (n_11312), .Y (n_7274));
NOR2X1 g70730(.A (n_12870), .B (n_29014), .Y (n_7272));
INVX1 g70731(.A (n_5918), .Y (n_13259));
INVX1 g70735(.A (n_5514), .Y (n_11046));
NAND2X1 g70738(.A (n_7106), .B (n_4522), .Y (n_11144));
NAND2X1 g70753(.A (n_27070), .B (n_6420), .Y (n_13116));
INVX1 g70755(.A (n_5594), .Y (n_11394));
INVX1 g72728(.A (n_6751), .Y (n_15352));
NOR2X1 g70770(.A (n_4704), .B (n_3017), .Y (n_8746));
INVX1 g70779(.A (n_6769), .Y (n_11565));
NOR2X1 g70783(.A (n_4704), .B (n_7266), .Y (n_7267));
NAND2X1 g70784(.A (n_6164), .B (n_7512), .Y (n_11582));
INVX1 g70788(.A (n_7264), .Y (n_8745));
NOR2X1 g70794(.A (n_7899), .B (n_6855), .Y (n_8743));
NAND2X1 g70796(.A (n_8759), .B (n_7262), .Y (n_7263));
INVX1 g70805(.A (n_5914), .Y (n_11311));
NAND2X1 g70823(.A (n_5684), .B (n_1147), .Y (n_13192));
INVX1 g70828(.A (n_5911), .Y (n_12563));
INVX1 g70830(.A (n_9355), .Y (n_16534));
NOR2X1 g70835(.A (n_6842), .B (n_8637), .Y (n_7260));
INVX1 g70857(.A (n_5906), .Y (n_8726));
OR2X1 g70860(.A (n_5343), .B (n_7496), .Y (n_8724));
OR2X1 g70863(.A (n_2994), .B (n_7258), .Y (n_7259));
NOR2X1 g70894(.A (n_5295), .B (n_9118), .Y (n_8266));
NAND2X1 g75534(.A (n_6539), .B (n_29244), .Y (n_7257));
NAND2X1 g70899(.A (n_7128), .B (n_3301), .Y (n_8714));
OR2X1 g70901(.A (n_17017), .B (n_2480), .Y (n_7256));
NAND2X1 g70903(.A (n_13646), .B (n_12335), .Y (n_7255));
AND2X1 g70905(.A (n_7159), .B (n_3307), .Y (n_8713));
NAND2X2 g70911(.A (n_7247), .B (n_4598), .Y (n_16394));
NOR2X1 g70913(.A (n_5931), .B (n_7636), .Y (n_11027));
INVX1 g70914(.A (n_7252), .Y (n_7253));
NAND2X1 g70920(.A (n_28163), .B (n_6877), .Y (n_19130));
NOR2X1 g71988(.A (n_3820), .B (n_2962), .Y (n_8427));
AOI21X1 g72700(.A0 (n_1997), .A1 (n_6868), .B0 (n_7183), .Y (n_7250));
INVX1 g70933(.A (n_5783), .Y (n_15340));
AND2X1 g70935(.A (n_4378), .B (n_13083), .Y (n_7249));
NAND2X1 g70941(.A (n_6934), .B (n_11385), .Y (n_12192));
NAND2X1 g70944(.A (n_16976), .B (n_4868), .Y (n_13676));
INVX1 g70947(.A (n_7048), .Y (n_17897));
INVX1 g70965(.A (n_7243), .Y (n_7244));
INVX1 g70971(.A (n_9350), .Y (n_8701));
INVX1 g70985(.A (n_9414), .Y (n_10939));
AND2X1 g70996(.A (n_7247), .B (n_8263), .Y (n_7242));
INVX2 g71000(.A (n_7241), .Y (n_8691));
INVX1 g71014(.A (n_9211), .Y (n_8685));
INVX1 g71025(.A (n_5897), .Y (n_8681));
OR2X1 g71028(.A (n_4262), .B (n_27099), .Y (n_7240));
NAND2X1 g71031(.A (n_7238), .B (n_2260), .Y (n_7239));
NOR2X1 g71033(.A (n_5285), .B (n_7598), .Y (n_7237));
NAND2X1 g72707(.A (n_5469), .B (n_4478), .Y (n_7233));
INVX1 g71055(.A (n_9389), .Y (n_11107));
NAND2X1 g71064(.A (n_3920), .B (n_2794), .Y (n_8671));
OR2X1 g71074(.A (n_2654), .B (n_7230), .Y (n_7232));
NAND2X2 g71082(.A (n_5667), .B (n_14055), .Y (n_14343));
INVX1 g71083(.A (n_7227), .Y (n_7228));
NAND2X1 g71090(.A (n_5555), .B (n_28423), .Y (n_8660));
INVX1 g71100(.A (n_7226), .Y (n_8652));
INVX1 g71107(.A (n_7221), .Y (n_7222));
NOR2X1 g71115(.A (n_5495), .B (n_7266), .Y (n_8649));
NAND2X1 g71022(.A (n_6791), .B (n_28757), .Y (n_7220));
INVX1 g71129(.A (n_7218), .Y (n_7219));
NAND2X1 g71131(.A (n_4900), .B (n_9410), .Y (n_10857));
NAND2X1 g71132(.A (n_7216), .B (n_7215), .Y (n_7217));
OR2X1 g71136(.A (n_7145), .B (n_14866), .Y (n_10854));
INVX1 g71141(.A (n_6041), .Y (n_8643));
XOR2X1 g76094(.A (text_in_r[1] ), .B (n_6400), .Y (n_7214));
NOR2X1 g71144(.A (n_4325), .B (n_7213), .Y (n_8641));
OR2X1 g71146(.A (n_5645), .B (n_8878), .Y (n_11327));
INVX1 g71149(.A (n_6056), .Y (n_16527));
INVX1 g71156(.A (n_5881), .Y (n_8633));
NOR2X1 g71161(.A (n_6887), .B (n_27133), .Y (n_7212));
INVX1 g72544(.A (n_5707), .Y (n_8293));
NOR2X1 g71168(.A (n_4330), .B (n_7210), .Y (n_7211));
NOR2X1 g71171(.A (n_5674), .B (n_4490), .Y (n_7209));
INVX1 g71172(.A (n_7207), .Y (n_7208));
NAND2X1 g71969(.A (n_5646), .B (n_15388), .Y (n_12337));
INVX1 g72691(.A (n_7204), .Y (n_7205));
OR2X1 g71215(.A (n_4820), .B (n_9388), .Y (n_11374));
NOR2X1 g71219(.A (n_7203), .B (n_9118), .Y (n_8620));
INVX1 g71220(.A (n_5870), .Y (n_12680));
OR2X1 g71222(.A (n_3692), .B (n_12169), .Y (n_18895));
INVX1 g71233(.A (n_9283), .Y (n_10950));
NOR2X1 g71238(.A (n_4997), .B (n_4898), .Y (n_7202));
OR2X1 g71241(.A (n_3444), .B (n_9527), .Y (n_8613));
NAND2X1 g71242(.A (n_5564), .B (n_7201), .Y (n_12594));
NOR2X1 g71966(.A (n_5272), .B (n_9942), .Y (n_7199));
NAND2X1 g71258(.A (n_12335), .B (n_3859), .Y (n_7198));
NAND2X1 g71262(.A (n_6334), .B (n_8878), .Y (n_10832));
INVX1 g71263(.A (n_5868), .Y (n_17531));
NAND2X1 g71266(.A (n_4679), .B (n_14589), .Y (n_7197));
NAND2X1 g71278(.A (n_7196), .B (n_4757), .Y (n_12243));
NOR2X1 g71282(.A (n_4174), .B (n_7176), .Y (n_7195));
INVX1 g71285(.A (n_6126), .Y (n_8600));
NAND2X1 g71300(.A (n_7194), .B (n_7193), .Y (n_18048));
NAND2X1 g71301(.A (n_2658), .B (n_6226), .Y (n_13134));
INVX1 g71309(.A (n_9319), .Y (n_11177));
AOI22X1 g62747(.A0 (n_3929), .A1 (dcnt[2] ), .B0 (n_1501), .B1(n_1694), .Y (n_7192));
AND2X1 g71316(.A (n_6169), .B (n_9982), .Y (n_7191));
OR2X1 g71318(.A (n_5367), .B (n_9118), .Y (n_7190));
NAND2X1 g71010(.A (n_5147), .B (n_6034), .Y (n_7187));
INVX1 g71333(.A (n_5864), .Y (n_8588));
NAND2X1 g71336(.A (n_4363), .B (n_7003), .Y (n_7184));
NOR2X1 g71345(.A (n_4721), .B (n_29410), .Y (n_8586));
NAND2X2 g71359(.A (n_7183), .B (n_7182), .Y (n_29336));
INVX1 g71361(.A (n_9370), .Y (n_7181));
INVX1 g71367(.A (n_5417), .Y (n_10827));
NAND2X1 g71380(.A (n_4138), .B (n_18369), .Y (n_7180));
INVX1 g71384(.A (n_7178), .Y (n_12500));
AND2X1 g71389(.A (n_7176), .B (n_4173), .Y (n_7177));
NAND2X1 g71391(.A (n_4447), .B (n_19226), .Y (n_7175));
INVX1 g71397(.A (n_7172), .Y (n_15825));
INVX1 g71950(.A (n_5808), .Y (n_8433));
NAND2X1 g71406(.A (n_7170), .B (n_7169), .Y (n_7171));
INVX1 g71422(.A (n_12399), .Y (n_11278));
NAND2X1 g71429(.A (n_5585), .B (n_6052), .Y (n_8566));
OR2X1 g71433(.A (n_3692), .B (n_12760), .Y (n_10675));
NAND2X1 g71434(.A (n_7085), .B (n_18369), .Y (n_10720));
INVX1 g71439(.A (n_7167), .Y (n_7168));
NAND2X1 g71449(.A (n_3307), .B (n_6060), .Y (n_9524));
NOR2X1 g71451(.A (n_4267), .B (n_7058), .Y (n_7166));
OR2X1 g71452(.A (n_7164), .B (n_12849), .Y (n_7165));
OR2X1 g71455(.A (n_6097), .B (n_7410), .Y (n_13142));
INVX1 g71458(.A (n_7162), .Y (n_9565));
INVX1 g71459(.A (n_7162), .Y (n_7163));
INVX1 g71465(.A (n_7161), .Y (n_9526));
INVX1 g71479(.A (n_7160), .Y (n_8550));
NAND2X1 g71489(.A (n_7159), .B (n_7158), .Y (n_15837));
INVX1 g71931(.A (n_5848), .Y (n_14240));
INVX1 g71500(.A (n_7157), .Y (n_11042));
NAND2X1 g71508(.A (n_3859), .B (n_26491), .Y (n_7155));
OR2X1 g72664(.A (n_6315), .B (n_5854), .Y (n_8258));
OR2X1 g71514(.A (n_3499), .B (n_14142), .Y (n_12136));
NOR2X1 g71517(.A (n_7152), .B (n_13738), .Y (n_7153));
INVX1 g71527(.A (n_10959), .Y (n_7147));
NOR2X1 g72636(.A (n_7114), .B (n_11489), .Y (n_12127));
INVX2 g71532(.A (n_7146), .Y (n_15627));
NOR2X1 g71535(.A (n_7145), .B (n_12827), .Y (n_8543));
NAND2X1 g71538(.A (n_7121), .B (n_10031), .Y (n_10952));
NOR2X1 g71938(.A (n_5165), .B (n_8742), .Y (n_7144));
NAND2X1 g71541(.A (n_4182), .B (n_16480), .Y (n_7143));
INVX1 g71545(.A (n_6330), .Y (n_7142));
INVX1 g74063(.A (n_11682), .Y (n_7141));
OR2X1 g71553(.A (n_6171), .B (n_7496), .Y (n_11161));
OR2X1 g71554(.A (n_3475), .B (n_11312), .Y (n_17024));
NAND2X1 g71557(.A (n_6245), .B (n_6247), .Y (n_7140));
INVX1 g71563(.A (n_5846), .Y (n_7139));
NAND2X1 g71573(.A (n_6913), .B (n_7137), .Y (n_7138));
NAND2X1 g71576(.A (n_26993), .B (n_7649), .Y (n_7136));
NAND2X1 g71579(.A (n_4923), .B (n_12169), .Y (n_10992));
NOR2X1 g71596(.A (n_2503), .B (n_7131), .Y (n_7132));
INVX1 g71599(.A (n_5842), .Y (n_13256));
INVX1 g71603(.A (n_5024), .Y (n_8523));
OR2X1 g71607(.A (n_2929), .B (n_7128), .Y (n_7130));
NAND2X2 g71616(.A (n_7127), .B (n_5646), .Y (n_10812));
NAND2X1 g71617(.A (n_7126), .B (n_5455), .Y (n_17123));
INVX1 g71619(.A (n_7124), .Y (n_7125));
NAND2X1 g71629(.A (n_7123), .B (n_11322), .Y (n_8515));
NOR2X1 g71630(.A (n_4903), .B (n_7410), .Y (n_19576));
NOR2X1 g71633(.A (n_7071), .B (n_9500), .Y (n_8514));
NAND2X1 g71635(.A (n_1085), .B (n_7121), .Y (n_14181));
INVX2 g71643(.A (n_5136), .Y (n_8511));
NOR2X1 g71648(.A (n_7120), .B (n_13815), .Y (n_12140));
INVX1 g71651(.A (n_5838), .Y (n_11655));
AND2X1 g71654(.A (n_12571), .B (n_6995), .Y (n_7119));
NAND2X2 g71662(.A (n_5602), .B (n_6185), .Y (n_13310));
OR2X1 g71671(.A (n_5654), .B (n_7116), .Y (n_7117));
NAND2X1 g71675(.A (n_3610), .B (n_11731), .Y (n_12370));
OR2X1 g71676(.A (n_7005), .B (n_165), .Y (n_13698));
INVX1 g71678(.A (n_5239), .Y (n_7115));
NOR2X1 g71681(.A (n_1513), .B (n_7114), .Y (n_18552));
NOR2X1 g71689(.A (n_7113), .B (n_7112), .Y (n_7930));
INVX1 g71691(.A (n_7109), .Y (n_7110));
OR2X1 g71693(.A (n_5188), .B (n_4173), .Y (n_7108));
NOR2X1 g73092(.A (n_13490), .B (n_2595), .Y (n_8154));
NAND2X1 g71700(.A (n_14113), .B (n_7106), .Y (n_16076));
NOR2X1 g71705(.A (n_4437), .B (n_15776), .Y (n_8496));
NAND2X1 g71709(.A (n_5956), .B (n_9410), .Y (n_7102));
NAND2X1 g71717(.A (n_7101), .B (n_7100), .Y (n_18064));
OR2X1 g71723(.A (n_4346), .B (n_12760), .Y (n_7099));
INVX2 g71729(.A (n_5418), .Y (n_11390));
NOR2X1 g71733(.A (n_3198), .B (n_6068), .Y (n_7098));
NAND2X1 g71736(.A (n_6907), .B (n_4861), .Y (n_29144));
INVX1 g77085(.A (n_7095), .Y (n_7096));
INVX1 g71740(.A (n_7093), .Y (n_11533));
INVX1 g71748(.A (n_5827), .Y (n_12546));
INVX1 g71753(.A (n_5436), .Y (n_8486));
NOR2X1 g71766(.A (n_8706), .B (n_6374), .Y (n_8481));
NAND2X1 g72711(.A (n_9371), .B (n_7486), .Y (n_7091));
INVX1 g71772(.A (n_5822), .Y (n_7090));
NOR2X1 g71785(.A (n_2733), .B (n_7593), .Y (n_7089));
NAND2X1 g71793(.A (n_6149), .B (n_4568), .Y (n_7088));
NOR2X1 g71795(.A (n_7085), .B (n_7084), .Y (n_7086));
INVX1 g71797(.A (n_7082), .Y (n_7083));
INVX1 g71801(.A (n_7081), .Y (n_8069));
INVX1 g71807(.A (n_7079), .Y (n_7077));
OR2X1 g72646(.A (n_3630), .B (n_5503), .Y (n_7076));
INVX1 g71822(.A (n_9315), .Y (n_8465));
INVX1 g71829(.A (n_7075), .Y (n_8462));
NAND2X1 g71834(.A (n_4367), .B (n_4757), .Y (n_13277));
NAND2X1 g71841(.A (n_5588), .B (n_4861), .Y (n_17356));
NAND2X1 g71842(.A (n_2794), .B (n_9057), .Y (n_12652));
NOR2X1 g71848(.A (n_11322), .B (n_7071), .Y (n_7072));
NAND2X1 g71851(.A (n_7069), .B (n_27124), .Y (n_11186));
INVX1 g71855(.A (n_9291), .Y (n_14940));
INVX1 g71859(.A (n_7068), .Y (n_11015));
INVX1 g71864(.A (n_7066), .Y (n_7067));
INVX1 g71869(.A (n_7065), .Y (n_8456));
INVX1 g71875(.A (n_7064), .Y (n_10834));
NAND2X1 g71887(.A (n_5574), .B (n_7201), .Y (n_8371));
INVX1 g71899(.A (n_5801), .Y (n_8454));
NOR2X1 g69534(.A (n_5289), .B (n_3307), .Y (n_10784));
NAND2X2 g71928(.A (n_5617), .B (n_330), .Y (n_11172));
NAND2X1 g71934(.A (n_6898), .B (n_8974), .Y (n_10984));
NOR2X1 g70958(.A (n_7062), .B (n_28749), .Y (n_7063));
INVX1 g71946(.A (n_5809), .Y (n_14399));
INVX2 g71959(.A (n_9285), .Y (n_8431));
NAND2X1 g71967(.A (n_7106), .B (n_7598), .Y (n_17762));
OR2X1 g71984(.A (n_5554), .B (n_8997), .Y (n_7061));
NAND2X1 g71989(.A (n_7058), .B (n_8997), .Y (n_7059));
OR2X1 g71990(.A (n_5548), .B (n_11385), .Y (n_7056));
NOR2X1 g71999(.A (n_5528), .B (n_9003), .Y (n_7053));
OR2X1 g72004(.A (n_4984), .B (n_28167), .Y (n_8421));
INVX1 g75110(.A (n_7052), .Y (n_7961));
NAND2X1 g72005(.A (n_7183), .B (n_9474), .Y (n_7051));
OR2X1 g72009(.A (n_4722), .B (n_17567), .Y (n_7050));
OR2X1 g72010(.A (n_4562), .B (n_12827), .Y (n_7047));
INVX1 g72023(.A (n_5048), .Y (n_8815));
INVX2 g72032(.A (n_5970), .Y (n_8417));
INVX1 g72035(.A (n_7044), .Y (n_7046));
NOR2X1 g72038(.A (n_6847), .B (n_5394), .Y (n_7043));
NAND2X2 g72043(.A (n_7058), .B (n_6783), .Y (n_8884));
NAND2X1 g72044(.A (n_13655), .B (n_12568), .Y (n_7042));
NAND2X1 g72047(.A (n_4327), .B (n_7041), .Y (n_11084));
OR2X1 g72048(.A (n_1063), .B (n_7039), .Y (n_7040));
INVX1 g74056(.A (n_5536), .Y (n_8030));
NOR2X1 g72075(.A (n_4675), .B (n_6902), .Y (n_7038));
NOR2X1 g72079(.A (n_10160), .B (n_6031), .Y (n_9181));
INVX1 g72083(.A (n_7036), .Y (n_8406));
INVX1 g72092(.A (n_7035), .Y (n_8399));
INVX1 g72097(.A (n_6028), .Y (n_9035));
INVX1 g72101(.A (n_6032), .Y (n_8398));
NAND2X2 g72105(.A (n_28163), .B (n_6977), .Y (n_13724));
NAND2X1 g72110(.A (n_14725), .B (n_7041), .Y (n_16000));
INVX1 g72112(.A (n_5792), .Y (n_13220));
INVX1 g72114(.A (n_5791), .Y (n_15109));
NAND2X1 g72116(.A (n_6266), .B (n_2260), .Y (n_10816));
NOR2X1 g72117(.A (n_4664), .B (n_7032), .Y (n_7033));
INVX1 g72118(.A (n_7030), .Y (n_7031));
NAND2X1 g72131(.A (n_7121), .B (n_14484), .Y (n_15103));
INVX1 g72136(.A (n_27409), .Y (n_7028));
NAND2X1 g72144(.A (n_7210), .B (n_7266), .Y (n_7026));
OR2X1 g72145(.A (n_7262), .B (n_1147), .Y (n_7025));
NAND2X1 g72150(.A (n_7023), .B (n_7069), .Y (n_10870));
NAND2X1 g73279(.A (n_4155), .B (n_14107), .Y (n_7022));
NOR2X1 g69511(.A (n_4476), .B (n_7498), .Y (n_9026));
NOR2X1 g72178(.A (n_3241), .B (n_5799), .Y (n_7018));
NOR2X1 g72183(.A (n_27686), .B (n_8435), .Y (n_7016));
NOR2X1 g72194(.A (n_8209), .B (n_8637), .Y (n_7015));
INVX1 g72197(.A (n_7013), .Y (n_7014));
NAND2X1 g72243(.A (n_5375), .B (n_11272), .Y (n_7011));
NAND2X2 g70926(.A (n_7176), .B (n_3820), .Y (n_16492));
INVX1 g72272(.A (n_5779), .Y (n_9286));
AND2X1 g72289(.A (n_7008), .B (n_11312), .Y (n_9299));
OR2X1 g72304(.A (n_7005), .B (n_11312), .Y (n_10797));
NAND2X1 g72305(.A (n_7003), .B (n_7376), .Y (n_7004));
INVX1 g72308(.A (n_7000), .Y (n_7002));
NOR2X1 g72326(.A (n_6280), .B (n_17260), .Y (n_6999));
NAND2X1 g72333(.A (n_4298), .B (n_14624), .Y (n_10932));
INVX1 g72335(.A (n_5772), .Y (n_9574));
NAND2X1 g72340(.A (n_6997), .B (n_6953), .Y (n_28836));
NAND2X1 g72359(.A (n_6995), .B (n_28037), .Y (n_6996));
NOR2X1 g72367(.A (n_5396), .B (n_26491), .Y (n_8338));
NAND2X1 g72369(.A (n_3270), .B (n_7658), .Y (n_11022));
INVX1 g72372(.A (n_6993), .Y (n_6994));
NOR2X1 g72380(.A (n_6991), .B (n_8099), .Y (n_6992));
AND2X1 g72391(.A (n_7406), .B (n_6989), .Y (n_6990));
NAND2X1 g72394(.A (n_7185), .B (n_6988), .Y (n_12383));
NAND2X1 g72395(.A (n_5138), .B (n_4612), .Y (n_6987));
NOR2X1 g72401(.A (n_3475), .B (n_1512), .Y (n_8328));
NOR2X1 g72406(.A (n_6114), .B (n_352), .Y (n_8326));
INVX1 g72409(.A (n_6985), .Y (n_6986));
NOR2X1 g72418(.A (n_27225), .B (n_5503), .Y (n_16300));
INVX1 g72428(.A (n_6982), .Y (n_6983));
NOR2X1 g72431(.A (n_6951), .B (n_29065), .Y (n_8319));
INVX1 g72439(.A (n_6979), .Y (n_6980));
NAND2X1 g72441(.A (n_7185), .B (n_5085), .Y (n_6978));
NAND2X1 g75796(.A (n_5093), .B (n_6977), .Y (n_9939));
OR2X1 g72448(.A (n_5337), .B (n_28410), .Y (n_6976));
NAND2X1 g72462(.A (n_6974), .B (n_27904), .Y (n_14902));
CLKBUFX3 g75790(.A (n_6972), .Y (n_9878));
INVX1 g72625(.A (n_5124), .Y (n_8354));
INVX1 g72475(.A (n_6971), .Y (n_7849));
INVX1 g72488(.A (n_9469), .Y (n_6970));
NAND3X1 g72490(.A (n_3725), .B (n_7101), .C (n_13679), .Y (n_6969));
NAND2X2 g72497(.A (n_5642), .B (n_5924), .Y (n_11097));
NAND2X1 g72501(.A (n_16895), .B (n_6968), .Y (n_7877));
INVX1 g72503(.A (n_5102), .Y (n_11221));
INVX1 g72508(.A (n_5120), .Y (n_13181));
NAND2X1 g72510(.A (n_7649), .B (n_6261), .Y (n_28450));
NOR2X1 g72512(.A (n_5118), .B (n_17260), .Y (n_6967));
NAND2X1 g72515(.A (n_10680), .B (n_7131), .Y (n_6966));
AND2X1 g72537(.A (n_5260), .B (n_27133), .Y (n_6965));
NAND2X1 g72547(.A (n_6963), .B (n_11253), .Y (n_6964));
NAND2X1 g72548(.A (n_6961), .B (n_6005), .Y (n_6962));
NAND2X1 g72560(.A (n_12134), .B (n_6960), .Y (n_11615));
NAND2X2 g70888(.A (n_5660), .B (n_6958), .Y (n_11008));
NAND2X1 g72565(.A (n_6961), .B (n_4721), .Y (n_8289));
NOR2X1 g72567(.A (n_12870), .B (n_4689), .Y (n_8287));
OR2X1 g72568(.A (n_8227), .B (n_6956), .Y (n_6957));
INVX1 g72571(.A (n_5485), .Y (n_11304));
NOR2X1 g72575(.A (n_2426), .B (n_16434), .Y (n_6955));
NAND2X1 g72582(.A (n_6953), .B (n_9084), .Y (n_8285));
INVX1 g75784(.A (n_6952), .Y (n_7911));
NOR2X1 g72617(.A (n_6951), .B (n_4689), .Y (n_17900));
NAND2X1 g72618(.A (n_5600), .B (n_5420), .Y (n_14454));
INVX2 g72631(.A (n_6950), .Y (n_10979));
INVX1 g72633(.A (n_5740), .Y (n_13236));
NAND2X1 g72641(.A (n_14831), .B (n_9257), .Y (n_6948));
NOR2X1 g72645(.A (n_5340), .B (n_28427), .Y (n_6947));
NOR2X1 g72653(.A (n_2699), .B (n_6946), .Y (n_8477));
OR2X1 g72654(.A (n_3198), .B (n_7292), .Y (n_6945));
INVX1 g72621(.A (n_6943), .Y (n_6944));
INVX2 g72669(.A (n_6942), .Y (n_10815));
NAND2X1 g72684(.A (n_6941), .B (n_6974), .Y (n_11040));
INVX1 g75778(.A (n_8569), .Y (n_8240));
OR2X1 g72708(.A (n_4496), .B (n_6939), .Y (n_6940));
NAND2X1 g71858(.A (n_5040), .B (n_7496), .Y (n_8458));
INVX1 g72714(.A (n_6937), .Y (n_6938));
INVX1 g72733(.A (n_11620), .Y (n_8760));
NOR2X1 g72735(.A (n_6934), .B (n_7576), .Y (n_6935));
NAND2X1 g72738(.A (n_5662), .B (n_6534), .Y (n_11157));
INVX1 g72745(.A (n_9217), .Y (n_16931));
NAND2X1 g72762(.A (n_4595), .B (n_6239), .Y (n_6933));
INVX1 g72781(.A (n_5726), .Y (n_17000));
NAND2X1 g72785(.A (n_6931), .B (n_6930), .Y (n_11554));
NAND2X1 g72787(.A (n_19110), .B (n_9163), .Y (n_6929));
NAND4X1 g66541(.A (n_14624), .B (n_7201), .C (n_2674), .D (n_4217),.Y (n_6928));
INVX1 g72791(.A (n_5991), .Y (n_11013));
NAND2X1 g72796(.A (n_6891), .B (n_10495), .Y (n_6927));
NAND2X1 g72799(.A (n_3656), .B (n_7201), .Y (n_6926));
NAND2X1 g72800(.A (n_4274), .B (n_4685), .Y (n_6924));
OR2X1 g72803(.A (n_3444), .B (n_9474), .Y (n_17021));
NOR2X1 g72811(.A (n_5525), .B (n_11322), .Y (n_6923));
NAND2X1 g72812(.A (n_7262), .B (n_11276), .Y (n_6922));
INVX1 g72614(.A (n_5742), .Y (n_8269));
NAND2X1 g72824(.A (n_6920), .B (n_9276), .Y (n_6921));
NAND2X1 g72825(.A (n_4179), .B (n_18369), .Y (n_6918));
INVX2 g72854(.A (n_6915), .Y (n_11259));
NAND2X1 g72865(.A (n_7583), .B (n_5854), .Y (n_12177));
OAI21X1 g72866(.A0 (n_6817), .A1 (n_2592), .B0 (n_6913), .Y (n_6914));
INVX1 g72874(.A (n_6910), .Y (n_6911));
NOR2X1 g72887(.A (n_3024), .B (n_6907), .Y (n_6908));
OR2X1 g72888(.A (n_4915), .B (n_7158), .Y (n_6906));
NOR2X1 g72897(.A (n_4332), .B (n_6963), .Y (n_6905));
OR2X1 g72898(.A (n_6212), .B (n_12169), .Y (n_10993));
NAND2X1 g72901(.A (n_5493), .B (n_6151), .Y (n_6904));
AND2X1 g72902(.A (n_6902), .B (n_28375), .Y (n_6903));
NAND2X1 g72906(.A (n_5077), .B (n_8945), .Y (n_6901));
INVX1 g72908(.A (n_6900), .Y (n_8195));
INVX1 g72911(.A (n_7473), .Y (n_15966));
NAND2X2 g72921(.A (n_4490), .B (n_6898), .Y (n_10948));
INVX1 g72929(.A (n_6896), .Y (n_6897));
NOR2X1 g72941(.A (n_5475), .B (n_17864), .Y (n_6895));
AND2X1 g72949(.A (n_12836), .B (n_6891), .Y (n_6892));
NAND2X1 g72957(.A (n_6304), .B (n_6462), .Y (n_8185));
OR2X1 g72958(.A (n_7230), .B (n_6889), .Y (n_6890));
NOR2X1 g72970(.A (n_6887), .B (n_28375), .Y (n_6888));
INVX1 g72971(.A (n_6884), .Y (n_6885));
INVX1 g72610(.A (n_5743), .Y (n_11345));
NOR2X1 g73005(.A (n_7258), .B (n_967), .Y (n_6882));
INVX1 g73013(.A (n_7668), .Y (n_6879));
NAND2X1 g73019(.A (n_5010), .B (n_6877), .Y (n_6878));
INVX1 g73022(.A (n_6875), .Y (n_8176));
INVX1 g73026(.A (n_6874), .Y (n_8174));
OR2X1 g73029(.A (n_4157), .B (n_1512), .Y (n_6873));
NAND2X1 g73033(.A (n_6871), .B (n_7159), .Y (n_6872));
INVX2 g73045(.A (n_6122), .Y (n_8167));
NAND2X1 g73053(.A (n_6870), .B (n_5541), .Y (n_18248));
INVX1 g73057(.A (n_13418), .Y (n_8163));
NAND2X1 g72932(.A (n_2632), .B (n_6868), .Y (n_10914));
INVX2 g70845(.A (n_5769), .Y (n_8730));
OR2X1 g73077(.A (n_6268), .B (n_1553), .Y (n_13226));
INVX1 g73082(.A (n_6866), .Y (n_12648));
INVX1 g73085(.A (n_6179), .Y (n_13171));
NOR2X1 g73089(.A (n_29410), .B (n_6005), .Y (n_6865));
OAI21X1 g75955(.A0 (n_4261), .A1 (n_28470), .B0 (n_3065), .Y(n_6863));
INVX1 g73105(.A (n_6202), .Y (n_9487));
INVX1 g73107(.A (n_6861), .Y (n_6862));
INVX1 g73121(.A (n_6858), .Y (n_13776));
INVX1 g73125(.A (n_5700), .Y (n_8146));
NAND2X1 g73135(.A (n_4110), .B (n_13571), .Y (n_17773));
AND2X1 g73136(.A (n_6856), .B (n_6855), .Y (n_6857));
INVX1 g73149(.A (n_6254), .Y (n_9523));
NAND2X1 g72604(.A (n_2803), .B (n_29286), .Y (n_8273));
INVX1 g75453(.A (n_6851), .Y (n_12144));
NAND2X1 g73160(.A (n_7730), .B (n_7477), .Y (n_6850));
NOR2X1 g73167(.A (n_5543), .B (n_8637), .Y (n_6849));
NOR2X1 g73168(.A (n_8209), .B (n_6847), .Y (n_6848));
NOR2X1 g73172(.A (n_2962), .B (n_27604), .Y (n_6846));
NAND2X1 g73181(.A (n_5355), .B (n_28427), .Y (n_9534));
NAND2X1 g73276(.A (n_4304), .B (n_15919), .Y (n_6844));
NOR2X1 g73198(.A (n_6842), .B (n_9819), .Y (n_6843));
OR2X1 g73203(.A (n_7203), .B (n_17411), .Y (n_6841));
OR2X1 g73204(.A (n_2827), .B (n_6838), .Y (n_6840));
NAND2X1 g73211(.A (n_6836), .B (n_6855), .Y (n_6837));
OR2X1 g73214(.A (n_4594), .B (n_7058), .Y (n_6835));
NAND2X1 g73215(.A (n_6833), .B (n_6374), .Y (n_6834));
OAI21X1 g73277(.A0 (n_1284), .A1 (n_3702), .B0 (n_10680), .Y(n_6831));
NAND2X1 g73237(.A (n_584), .B (n_6829), .Y (n_6830));
OAI21X1 g73239(.A0 (n_6827), .A1 (n_1186), .B0 (n_6825), .Y (n_6828));
OAI21X1 g73249(.A0 (n_15812), .A1 (n_1989), .B0 (n_7406), .Y(n_6824));
NAND2X1 g73250(.A (n_1173), .B (n_6822), .Y (n_6823));
AOI21X1 g73252(.A0 (n_5368), .A1 (n_28870), .B0 (n_4772), .Y(n_6821));
NAND2X1 g71044(.A (n_2658), .B (n_5422), .Y (n_8675));
OAI21X1 g73268(.A0 (n_6817), .A1 (n_3464), .B0 (n_4325), .Y (n_6818));
INVX1 g69386(.A (n_6038), .Y (n_9056));
AOI21X1 g73275(.A0 (n_2864), .A1 (n_2671), .B0 (n_2873), .Y (n_6816));
NAND2X1 g73278(.A (n_4229), .B (n_10147), .Y (n_6815));
NAND2X1 g73280(.A (n_4406), .B (n_8317), .Y (n_6814));
NAND2X1 g73281(.A (n_4211), .B (n_16006), .Y (n_6813));
NAND2X1 g73282(.A (n_4201), .B (n_2281), .Y (n_6812));
INVX1 g70818(.A (n_6811), .Y (n_8736));
AOI21X1 g73288(.A0 (n_3301), .A1 (n_5305), .B0 (n_4502), .Y (n_6810));
INVX1 g74634(.A (n_6809), .Y (n_7997));
AOI21X1 g73289(.A0 (n_13679), .A1 (n_5231), .B0 (n_4789), .Y(n_6808));
INVX1 g70812(.A (n_5913), .Y (n_8737));
AOI21X1 g73296(.A0 (n_6805), .A1 (n_2181), .B0 (n_4150), .Y (n_6806));
NAND2X1 g73314(.A (n_4830), .B (n_14484), .Y (n_6804));
NOR2X1 g75446(.A (n_26494), .B (n_11052), .Y (n_6803));
INVX2 g73341(.A (n_7294), .Y (n_8086));
NOR2X1 g74630(.A (n_4738), .B (n_7201), .Y (n_6802));
NAND2X1 g69374(.A (n_5590), .B (n_6012), .Y (n_10806));
NAND2X1 g73362(.A (n_5020), .B (n_9442), .Y (n_6801));
OR2X1 g73388(.A (n_4514), .B (n_19857), .Y (n_6797));
INVX1 g73418(.A (n_6094), .Y (n_10777));
NAND2X1 g71816(.A (n_6791), .B (n_6790), .Y (n_8466));
INVX1 g75744(.A (n_5211), .Y (n_10369));
NAND2X1 g75945(.A (n_6833), .B (n_7701), .Y (n_6785));
NAND2X1 g73521(.A (n_6428), .B (n_6783), .Y (n_6784));
INVX1 g73544(.A (n_8971), .Y (n_10237));
INVX2 g73560(.A (n_9037), .Y (n_10101));
NAND2X1 g73589(.A (n_4004), .B (n_28375), .Y (n_6780));
NOR2X1 g70785(.A (n_5578), .B (n_13804), .Y (n_6779));
INVX4 g73682(.A (n_8709), .Y (n_10034));
OR2X1 g73686(.A (n_6677), .B (n_1147), .Y (n_10904));
INVX1 g73691(.A (n_5611), .Y (n_14067));
NOR2X1 g73699(.A (n_6293), .B (n_6252), .Y (n_8063));
INVX1 g73703(.A (n_5608), .Y (n_10775));
NAND2X1 g73711(.A (n_6210), .B (n_5005), .Y (n_6775));
INVX1 g73712(.A (n_6773), .Y (n_6774));
NAND2X1 g73272(.A (n_4453), .B (n_2757), .Y (n_6772));
OR2X1 g73756(.A (n_6767), .B (n_5329), .Y (n_6768));
NAND2X1 g72586(.A (n_4477), .B (n_15588), .Y (n_6766));
INVX1 g73849(.A (n_6760), .Y (n_6762));
INVX1 g73855(.A (n_9907), .Y (n_6759));
INVX1 g73858(.A (n_6758), .Y (n_9803));
NAND2X1 g73270(.A (n_4339), .B (n_4807), .Y (n_6756));
INVX1 g73877(.A (n_4993), .Y (n_10305));
NAND2X1 g73881(.A (n_5323), .B (n_4865), .Y (n_6755));
INVX1 g75734(.A (n_8564), .Y (n_6754));
NOR2X1 g75937(.A (n_6260), .B (n_6749), .Y (n_9699));
INVX1 g73920(.A (n_6748), .Y (n_6747));
INVX1 g73927(.A (n_6746), .Y (n_8047));
INVX1 g73938(.A (n_8172), .Y (n_6745));
NOR2X1 g71918(.A (n_6227), .B (n_9417), .Y (n_8445));
INVX1 g73957(.A (n_6742), .Y (n_6743));
INVX1 g73960(.A (n_6740), .Y (n_6739));
NOR2X1 g73969(.A (n_6096), .B (n_5413), .Y (n_7890));
INVX1 g73979(.A (n_6733), .Y (n_6734));
NOR2X1 g75933(.A (n_6730), .B (n_3016), .Y (n_6731));
CLKBUFX3 g74029(.A (n_6727), .Y (n_9900));
INVX1 g74035(.A (n_6725), .Y (n_6724));
INVX1 g71776(.A (n_6723), .Y (n_8478));
NAND2X1 g74046(.A (n_3594), .B (n_7512), .Y (n_6721));
NOR2X1 g74048(.A (n_5007), .B (n_11731), .Y (n_6720));
INVX1 g74067(.A (n_8644), .Y (n_6717));
INVX1 g74069(.A (n_6716), .Y (n_10355));
INVX1 g74073(.A (n_8250), .Y (n_6715));
INVX1 g74079(.A (n_6714), .Y (n_10513));
INVX1 g74082(.A (n_6712), .Y (n_6713));
INVX1 g74085(.A (n_6711), .Y (n_8026));
NOR2X1 g72576(.A (n_4887), .B (n_7238), .Y (n_6709));
NAND3X1 g74108(.A (n_29062), .B (n_6328), .C (n_9442), .Y (n_6705));
INVX1 g74141(.A (n_6701), .Y (n_10312));
INVX1 g74146(.A (n_6699), .Y (n_6700));
INVX1 g74160(.A (n_8603), .Y (n_6697));
NAND3X1 g74176(.A (n_6696), .B (n_13679), .C (n_11307), .Y (n_17841));
OR2X1 g74185(.A (n_6694), .B (n_3071), .Y (n_15462));
INVX1 g74189(.A (n_6325), .Y (n_29426));
INVX1 g74217(.A (n_7683), .Y (n_6692));
INVX1 g74246(.A (n_6687), .Y (n_6688));
INVX1 g74278(.A (n_6684), .Y (n_6685));
INVX1 g74301(.A (n_7763), .Y (n_6681));
NAND2X1 g74316(.A (n_4976), .B (n_8090), .Y (n_6680));
INVX1 g74323(.A (n_6679), .Y (n_11110));
NAND2X1 g74330(.A (n_6677), .B (n_4663), .Y (n_6678));
NOR2X1 g74339(.A (n_6194), .B (n_5413), .Y (n_6676));
INVX1 g74344(.A (n_6673), .Y (n_6674));
INVX1 g75925(.A (n_6671), .Y (n_6672));
INVX1 g74384(.A (n_6670), .Y (n_9823));
NAND2X1 g74387(.A (n_8846), .B (n_6749), .Y (n_6669));
INVX1 g74402(.A (n_6665), .Y (n_10573));
INVX1 g74411(.A (n_6661), .Y (n_12123));
INVX1 g74415(.A (n_6659), .Y (n_6660));
NAND2X2 g74418(.A (n_4084), .B (n_27904), .Y (n_10140));
OR2X1 g74429(.A (n_8418), .B (n_6656), .Y (n_6657));
OR2X1 g74431(.A (n_7899), .B (n_6856), .Y (n_6655));
NOR2X1 g74457(.A (n_5096), .B (n_11272), .Y (n_9716));
INVX1 g74488(.A (n_8441), .Y (n_6653));
NAND2X1 g74508(.A (n_3147), .B (n_9500), .Y (n_6652));
INVX1 g74517(.A (n_5446), .Y (n_10551));
INVX1 g74521(.A (n_6647), .Y (n_6648));
NAND2X1 g74555(.A (n_6603), .B (n_11835), .Y (n_6645));
NAND2X1 g74579(.A (n_2183), .B (n_3694), .Y (n_6644));
INVX1 g74591(.A (n_8393), .Y (n_9791));
INVX1 g74615(.A (n_6640), .Y (n_6641));
NAND2X1 g74618(.A (n_6931), .B (n_3874), .Y (n_6639));
INVX1 g74625(.A (n_8490), .Y (n_7999));
NAND2X1 g74676(.A (n_12858), .B (n_6636), .Y (n_6637));
OR2X1 g74677(.A (n_4099), .B (n_10031), .Y (n_6635));
INVX1 g74684(.A (n_8218), .Y (n_6634));
INVX1 g74690(.A (n_6633), .Y (n_10081));
NAND3X1 g74723(.A (n_14807), .B (n_3807), .C (n_2592), .Y (n_6627));
INVX1 g74724(.A (n_6623), .Y (n_6624));
OR2X1 g74729(.A (n_6620), .B (n_4187), .Y (n_6621));
NAND2X1 g74733(.A (n_9965), .B (n_3204), .Y (n_6619));
INVX1 g74735(.A (n_12778), .Y (n_6618));
INVX1 g74737(.A (n_6183), .Y (n_6616));
INVX1 g74755(.A (n_6614), .Y (n_6615));
NAND2X1 g75922(.A (n_12249), .B (n_5834), .Y (n_6613));
NAND2X1 g74763(.A (n_4760), .B (n_6442), .Y (n_6612));
NAND2X1 g74771(.A (n_3388), .B (n_7201), .Y (n_6610));
OR2X1 g74778(.A (n_6609), .B (n_3723), .Y (n_15468));
NAND2X2 g70676(.A (n_5625), .B (n_27365), .Y (n_8769));
INVX1 g74788(.A (n_6606), .Y (n_6607));
NAND2X1 g74803(.A (n_6603), .B (n_27604), .Y (n_6604));
INVX1 g74840(.A (n_9073), .Y (n_6600));
INVX1 g74842(.A (n_6598), .Y (n_6599));
INVX1 g74856(.A (n_8438), .Y (n_6595));
INVX1 g74858(.A (n_6593), .Y (n_6594));
OR2X1 g74860(.A (n_5108), .B (n_27990), .Y (n_6592));
NOR2X1 g74882(.A (n_3240), .B (n_14484), .Y (n_6590));
INVX1 g74890(.A (n_6588), .Y (n_6589));
NAND3X1 g74893(.A (n_6587), .B (n_3301), .C (n_7410), .Y (n_19568));
INVX1 g74600(.A (n_8392), .Y (n_6586));
INVX1 g74919(.A (n_6584), .Y (n_6583));
NAND2X1 g72546(.A (n_11916), .B (n_6582), .Y (n_13119));
INVX2 g74928(.A (n_6581), .Y (n_10162));
NAND2X1 g74932(.A (n_6495), .B (n_10389), .Y (n_6580));
OR2X1 g74934(.A (n_5052), .B (n_1147), .Y (n_6579));
INVX1 g74939(.A (n_6577), .Y (n_6578));
INVX1 g74950(.A (n_6574), .Y (n_6575));
OR2X1 g74968(.A (n_3938), .B (n_4514), .Y (n_6573));
OR2X1 g74980(.A (n_3443), .B (n_4158), .Y (n_6571));
NAND2X1 g74988(.A (n_6522), .B (n_15894), .Y (n_6569));
AND2X1 g74996(.A (n_3778), .B (n_6400), .Y (n_6567));
NOR2X1 g75010(.A (n_3003), .B (n_3482), .Y (n_6565));
NAND2X1 g75019(.A (n_2883), .B (n_7362), .Y (n_7966));
NOR2X1 g75029(.A (n_5018), .B (n_11272), .Y (n_6564));
INVX1 g75033(.A (n_6563), .Y (n_7925));
NAND2X1 g75064(.A (n_3225), .B (n_9442), .Y (n_6558));
NAND2X1 g75075(.A (n_25745), .B (n_3755), .Y (n_6557));
INVX1 g75079(.A (n_6556), .Y (n_7963));
NAND3X1 g75081(.A (n_16754), .B (n_4721), .C (n_6554), .Y (n_6555));
NAND2X1 g75091(.A (n_1447), .B (n_3071), .Y (n_6553));
INVX1 g75092(.A (n_8127), .Y (n_9841));
OR2X1 g75698(.A (n_3281), .B (n_4334), .Y (n_6551));
INVX1 g75113(.A (n_6549), .Y (n_10020));
INVX1 g75119(.A (n_6420), .Y (n_6548));
NOR2X1 g75124(.A (n_6546), .B (n_5558), .Y (n_6547));
INVX1 g75129(.A (n_5140), .Y (n_7959));
INVX1 g75132(.A (n_6544), .Y (n_6545));
NOR2X1 g69214(.A (n_28616), .B (n_15894), .Y (n_6542));
NAND2X1 g75155(.A (n_6539), .B (n_19791), .Y (n_6540));
OR2X1 g75160(.A (n_4002), .B (n_4113), .Y (n_6537));
INVX1 g75161(.A (n_6536), .Y (n_10284));
NOR2X1 g75168(.A (n_4777), .B (n_6534), .Y (n_6535));
INVX1 g75175(.A (n_6532), .Y (n_6533));
INVX1 g75184(.A (n_6204), .Y (n_6531));
INVX1 g75189(.A (n_6529), .Y (n_6530));
OR2X1 g75193(.A (n_6527), .B (n_9704), .Y (n_6528));
NAND2X1 g75211(.A (n_6522), .B (n_6534), .Y (n_6523));
AND2X1 g75212(.A (n_3915), .B (n_8928), .Y (n_6521));
INVX1 g75213(.A (n_7778), .Y (n_10440));
INVX1 g75892(.A (n_6515), .Y (n_6516));
NAND3X1 g72542(.A (n_3989), .B (n_6510), .C (n_15473), .Y (n_6511));
NAND2X1 g75297(.A (n_5074), .B (n_27124), .Y (n_10130));
NAND2X1 g75310(.A (n_4864), .B (n_13679), .Y (n_6505));
INVX1 g75341(.A (n_6500), .Y (n_9772));
INVX2 g71697(.A (n_6499), .Y (n_12883));
NAND2X1 g75364(.A (n_12249), .B (n_6497), .Y (n_6498));
NAND2X1 g75372(.A (n_6495), .B (n_15610), .Y (n_6496));
NAND2X1 g71695(.A (n_6060), .B (n_7658), .Y (n_10936));
INVX1 g75399(.A (n_6494), .Y (n_12121));
INVX1 g75403(.A (n_12747), .Y (n_6493));
INVX1 g75413(.A (n_8284), .Y (n_9798));
INVX1 g75432(.A (n_6492), .Y (n_9735));
INVX2 g75441(.A (n_8253), .Y (n_8068));
INVX1 g75469(.A (n_6491), .Y (n_9946));
INVX2 g70624(.A (n_9353), .Y (n_11362));
INVX1 g75505(.A (n_6489), .Y (n_6490));
INVX1 g75507(.A (n_8493), .Y (n_6488));
NAND2X1 g75511(.A (n_4760), .B (n_6486), .Y (n_7927));
INVX1 g75512(.A (n_7787), .Y (n_10030));
INVX1 g75561(.A (n_7367), .Y (n_6482));
NAND2X1 g75578(.A (n_6479), .B (n_1424), .Y (n_6480));
NAND2X1 g75585(.A (n_4083), .B (n_28757), .Y (n_6478));
INVX1 g74584(.A (n_6477), .Y (n_8000));
INVX1 g75602(.A (n_9050), .Y (n_6476));
INVX1 g75627(.A (n_6475), .Y (n_7867));
INVX1 g72532(.A (n_3305), .Y (n_8298));
INVX1 g73992(.A (n_12436), .Y (n_8035));
INVX1 g75671(.A (n_6470), .Y (n_9958));
NOR2X1 g75719(.A (n_3671), .B (n_5854), .Y (n_6469));
INVX1 g75720(.A (n_9645), .Y (n_6468));
NAND2X1 g75750(.A (n_3710), .B (n_7325), .Y (n_6464));
NAND2X1 g69188(.A (n_5408), .B (n_6462), .Y (n_6463));
INVX1 g75765(.A (n_6461), .Y (n_7913));
NAND2X2 g72528(.A (n_6907), .B (n_636), .Y (n_8300));
INVX1 g75681(.A (n_6458), .Y (n_6459));
NAND2X1 g75836(.A (n_3778), .B (n_15507), .Y (n_6457));
INVX1 g75840(.A (n_8076), .Y (n_9997));
NAND2X1 g75866(.A (n_8105), .B (n_6452), .Y (n_6453));
NAND2X1 g75872(.A (n_4824), .B (n_6198), .Y (n_6451));
NOR2X1 g75873(.A (n_5074), .B (n_28869), .Y (n_6450));
INVX1 g75877(.A (n_6448), .Y (n_6449));
NAND2X1 g75883(.A (n_6446), .B (n_6445), .Y (n_6447));
NAND2X1 g75885(.A (n_10199), .B (n_5091), .Y (n_9555));
NAND2X1 g72524(.A (n_3045), .B (n_6974), .Y (n_8301));
NOR2X1 g75890(.A (n_6444), .B (n_6636), .Y (n_9714));
INVX1 g69860(.A (n_6443), .Y (n_13162));
INVX1 g75906(.A (n_6440), .Y (n_6441));
NAND2X1 g75932(.A (n_12249), .B (n_6439), .Y (n_10786));
NAND2X1 g75938(.A (n_6836), .B (n_6856), .Y (n_6438));
NAND2X1 g75941(.A (n_10127), .B (n_4037), .Y (n_6437));
INVX1 g75946(.A (n_6435), .Y (n_6436));
AND2X1 g75949(.A (n_16895), .B (n_3204), .Y (n_6434));
OAI21X1 g75957(.A0 (n_13679), .A1 (n_6431), .B0 (n_2678), .Y(n_6432));
NOR2X1 g75962(.A (n_3835), .B (n_6428), .Y (n_6429));
OAI21X1 g75964(.A0 (n_9691), .A1 (n_3560), .B0 (n_6426), .Y (n_6427));
NOR2X1 g71657(.A (n_4212), .B (n_28724), .Y (n_6425));
OAI21X1 g73274(.A0 (n_2724), .A1 (n_6486), .B0 (n_6422), .Y (n_6423));
OAI21X1 g61895(.A0 (n_3202), .A1 (n_10999), .B0 (n_9249), .Y(n_6421));
NAND2X1 g70570(.A (n_6420), .B (n_6419), .Y (n_8801));
INVX1 g73975(.A (n_6738), .Y (n_6418));
INVX1 g75002(.A (n_6417), .Y (n_7968));
NOR2X1 g69142(.A (n_6415), .B (n_11253), .Y (n_6416));
NAND2X1 g73242(.A (n_4929), .B (n_27432), .Y (n_6414));
AND2X1 g75900(.A (n_14548), .B (n_3874), .Y (n_6413));
NAND2X1 g75000(.A (n_6406), .B (n_3138), .Y (n_6407));
XOR2X1 g76199(.A (n_6404), .B (n_2870), .Y (n_6405));
XOR2X1 g76203(.A (n_6401), .B (n_6400), .Y (n_6402));
NAND2X1 g70518(.A (n_5721), .B (n_27990), .Y (n_6399));
INVX1 g75326(.A (n_5290), .Y (n_10610));
XOR2X1 g76287(.A (n_234), .B (n_4750), .Y (n_6398));
XOR2X1 g76311(.A (text_in_r[31] ), .B (n_3667), .Y (n_6396));
OR2X1 g75647(.A (n_4493), .B (n_10452), .Y (n_6394));
INVX1 g74977(.A (n_6392), .Y (n_6393));
INVX1 g76392(.A (n_7628), .Y (n_25332));
INVX1 g76393(.A (n_7628), .Y (n_25370));
INVX1 g76400(.A (n_6391), .Y (n_25407));
INVX1 g75638(.A (n_6390), .Y (n_7921));
AND2X1 g71624(.A (n_6838), .B (n_6868), .Y (n_8516));
OR2X1 g73956(.A (n_3796), .B (n_11731), .Y (n_8037));
INVX1 g76757(.A (n_6853), .Y (n_6386));
NAND2X2 g69062(.A (n_5430), .B (n_383), .Y (n_9127));
INVX2 g74532(.A (n_6384), .Y (n_10146));
NAND2X1 g69048(.A (n_27076), .B (n_29228), .Y (n_9129));
INVX1 g75631(.A (n_6376), .Y (n_6377));
AND2X1 g72496(.A (n_7701), .B (n_6374), .Y (n_6375));
INVX1 g77040(.A (n_6372), .Y (n_6373));
AND2X1 g72494(.A (n_2923), .B (n_9528), .Y (n_6371));
OR2X1 g75623(.A (n_5061), .B (n_6997), .Y (n_6370));
OR2X1 g71612(.A (n_3499), .B (n_9388), .Y (n_17018));
OR2X1 g72238(.A (n_6368), .B (n_8974), .Y (n_6369));
INVX1 g74952(.A (n_6366), .Y (n_10157));
INVX1 g75308(.A (n_5032), .Y (n_7942));
INVX1 g77657(.A (n_6364), .Y (n_6365));
NAND2X2 g68994(.A (n_5373), .B (n_6977), .Y (n_9142));
INVX1 g75618(.A (n_8141), .Y (n_9849));
INVX2 g70456(.A (n_6363), .Y (n_8818));
NAND2X1 g71606(.A (n_5439), .B (n_1376), .Y (n_11131));
NOR2X1 g68975(.A (n_6239), .B (n_9368), .Y (n_9145));
NOR2X1 g74505(.A (n_4573), .B (n_11253), .Y (n_6361));
NAND2X1 g74492(.A (n_6285), .B (n_8945), .Y (n_9930));
AND2X1 g71592(.A (n_7203), .B (n_13799), .Y (n_6358));
INVX1 g74486(.A (n_8561), .Y (n_9779));
INVX1 g74930(.A (n_8951), .Y (n_6356));
NAND2X1 g71590(.A (n_6963), .B (n_5660), .Y (n_8527));
INVX1 g75607(.A (n_6354), .Y (n_6355));
NOR2X1 g75888(.A (n_1806), .B (n_3710), .Y (n_6353));
INVX1 g80175(.A (n_4837), .Y (n_6352));
INVX1 g75286(.A (n_6350), .Y (n_7944));
NAND2X1 g77872(.A (n_2744), .B (n_5924), .Y (n_7845));
NAND2X1 g73856(.A (n_3010), .B (n_27365), .Y (n_9907));
OR2X1 g74912(.A (n_9999), .B (n_6346), .Y (n_6347));
NOR2X1 g70402(.A (n_5942), .B (n_7658), .Y (n_7315));
DFFX1 text_in_r_reg[116] (.CK (clk), .D (n_3223), .Q(text_in_r[116] ), .QN ());
DFFX1 text_in_r_reg[111] (.CK (clk), .D (n_3870), .Q(text_in_r[111] ), .QN ());
DFFX1 text_in_r_reg[37] (.CK (clk), .D (n_3210), .Q (text_in_r[37]), .QN ());
NOR2X1 g70386(.A (n_4203), .B (n_379), .Y (n_7976));
DFFX1 text_in_r_reg[14] (.CK (clk), .D (n_3565), .Q (text_in_r[14]), .QN ());
DFFX1 text_in_r_reg[67] (.CK (clk), .D (n_3851), .Q (text_in_r[67]), .QN ());
DFFX1 text_in_r_reg[47] (.CK (clk), .D (n_3933), .Q (text_in_r[47]), .QN ());
INVX1 g75599(.A (n_4969), .Y (n_7840));
NAND2X1 g75653(.A (n_2311), .B (n_1989), .Y (n_6341));
INVX1 g74903(.A (n_6339), .Y (n_7841));
INVX1 g77863(.A (n_6677), .Y (n_6338));
INVX1 g74460(.A (n_28156), .Y (n_7837));
INVX1 g75654(.A (n_6791), .Y (n_6337));
DFFX1 text_in_r_reg[18] (.CK (clk), .D (n_3089), .Q (text_in_r[18]), .QN ());
INVX1 g73860(.A (n_4962), .Y (n_6758));
DFFX1 text_in_r_reg[0] (.CK (clk), .D (n_3227), .Q (text_in_r[0] ),.QN ());
INVX1 g75454(.A (n_7106), .Y (n_6851));
NOR2X1 g70366(.A (n_4439), .B (n_4709), .Y (n_7322));
NAND2X1 g75080(.A (n_5612), .B (n_6021), .Y (n_6556));
INVX1 g72464(.A (n_7665), .Y (n_17286));
NOR2X1 g76945(.A (n_6335), .B (n_7410), .Y (n_6336));
INVX1 g74042(.A (n_6334), .Y (n_11104));
CLKBUFX3 g74446(.A (n_6332), .Y (n_8015));
DFFX1 text_in_r_reg[68] (.CK (clk), .D (n_3619), .Q (text_in_r[68]), .QN ());
INVX1 g75587(.A (n_4945), .Y (n_8541));
OR2X1 g71546(.A (n_3304), .B (n_8217), .Y (n_6330));
DFFX1 text_in_r_reg[49] (.CK (clk), .D (n_3216), .Q (text_in_r[49]), .QN ());
NAND2X1 g74889(.A (n_5516), .B (n_6328), .Y (n_6329));
NOR2X1 g74891(.A (n_6327), .B (n_8742), .Y (n_6588));
DFFX1 text_in_r_reg[42] (.CK (clk), .D (n_3328), .Q (text_in_r[42]), .QN ());
NOR2X1 g74190(.A (n_3226), .B (n_6462), .Y (n_6325));
INVX1 g74695(.A (n_4691), .Y (n_8039));
INVX1 g73838(.A (n_4938), .Y (n_6764));
OR2X1 g71536(.A (n_6099), .B (n_13490), .Y (n_11585));
NAND2X1 g77576(.A (n_13679), .B (n_23422), .Y (n_6319));
INVX1 g74432(.A (n_6315), .Y (n_8548));
NAND2X1 g74430(.A (n_6313), .B (n_28472), .Y (n_6314));
AND2X1 g70308(.A (n_6025), .B (n_3307), .Y (n_9322));
INVX1 g73829(.A (n_4499), .Y (n_7820));
NOR2X1 g72440(.A (n_5716), .B (n_15388), .Y (n_6979));
NOR2X1 g75583(.A (n_7721), .B (n_8865), .Y (n_14531));
INVX1 g73360(.A (n_5675), .Y (n_6312));
INVX2 g74425(.A (n_6031), .Y (n_8396));
NOR2X1 g70302(.A (n_5005), .B (n_4881), .Y (n_7343));
NOR2X1 g74880(.A (n_3131), .B (n_383), .Y (n_6310));
NAND2X1 g71528(.A (n_4855), .B (n_6462), .Y (n_10959));
NAND2X1 g73993(.A (n_3831), .B (n_5413), .Y (n_12436));
INVX1 g74875(.A (n_7415), .Y (n_6306));
INVX1 g75111(.A (n_7062), .Y (n_7052));
NOR2X1 g74874(.A (n_3176), .B (n_4042), .Y (n_8110));
INVX1 g73822(.A (n_4927), .Y (n_8817));
NOR2X1 g70285(.A (n_3820), .B (n_25629), .Y (n_7815));
NOR2X1 g74416(.A (n_3837), .B (n_6303), .Y (n_6659));
NOR2X1 g62157(.A (n_6301), .B (n_3286), .Y (n_6302));
DFFX1 text_in_r_reg[127] (.CK (clk), .D (n_3020), .Q(text_in_r[127] ), .QN ());
INVX1 g73820(.A (n_4417), .Y (n_7812));
DFFX1 text_in_r_reg[64] (.CK (clk), .D (n_3224), .Q (text_in_r[64]), .QN ());
DFFX1 text_in_r_reg[54] (.CK (clk), .D (n_3930), .Q (text_in_r[54]), .QN ());
OR2X1 g75813(.A (n_3697), .B (n_10599), .Y (n_6298));
DFFX1 text_in_r_reg[35] (.CK (clk), .D (n_3613), .Q (text_in_r[35]), .QN ());
DFFX1 text_in_r_reg[6] (.CK (clk), .D (n_3292), .Q (text_in_r[6] ),.QN ());
INVX1 g74864(.A (n_6295), .Y (n_9970));
DFFX1 text_in_r_reg[17] (.CK (clk), .D (n_3410), .Q (text_in_r[17]), .QN ());
DFFX1 text_in_r_reg[108] (.CK (clk), .D (n_3703), .Q(text_in_r[108] ), .QN ());
DFFX1 text_in_r_reg[11] (.CK (clk), .D (n_3916), .Q (text_in_r[11]), .QN ());
DFFX1 text_in_r_reg[123] (.CK (clk), .D (n_3804), .Q(text_in_r[123] ), .QN ());
DFFX1 text_in_r_reg[24] (.CK (clk), .D (n_3895), .Q (text_in_r[24]), .QN ());
DFFX1 text_in_r_reg[26] (.CK (clk), .D (n_3362), .Q (text_in_r[26]), .QN ());
DFFX1 text_in_r_reg[29] (.CK (clk), .D (n_3405), .Q (text_in_r[29]), .QN ());
DFFX1 text_in_r_reg[46] (.CK (clk), .D (n_3433), .Q (text_in_r[46]), .QN ());
DFFX1 text_in_r_reg[55] (.CK (clk), .D (n_3466), .Q (text_in_r[55]), .QN ());
DFFX1 text_in_r_reg[61] (.CK (clk), .D (n_3172), .Q (text_in_r[61]), .QN ());
DFFX1 text_in_r_reg[63] (.CK (clk), .D (n_3429), .Q (text_in_r[63]), .QN ());
DFFX1 text_in_r_reg[78] (.CK (clk), .D (n_3642), .Q (text_in_r[78]), .QN ());
DFFX1 text_in_r_reg[81] (.CK (clk), .D (n_3485), .Q (text_in_r[81]), .QN ());
DFFX1 text_in_r_reg[86] (.CK (clk), .D (n_3621), .Q (text_in_r[86]), .QN ());
DFFX1 text_in_r_reg[8] (.CK (clk), .D (n_3367), .Q (text_in_r[8] ),.QN ());
DFFX1 text_in_r_reg[99] (.CK (clk), .D (n_3375), .Q (text_in_r[99]), .QN ());
CLKBUFX1 g74403(.A (n_7069), .Y (n_6665));
AND2X1 g77363(.A (n_7410), .B (n_933), .Y (n_6294));
DFFX1 text_in_r_reg[91] (.CK (clk), .D (n_3406), .Q (text_in_r[91]), .QN ());
DFFX1 text_in_r_reg[39] (.CK (clk), .D (n_3347), .Q (text_in_r[39]), .QN ());
DFFX1 text_in_r_reg[60] (.CK (clk), .D (n_3519), .Q (text_in_r[60]), .QN ());
DFFX1 text_in_r_reg[103] (.CK (clk), .D (n_3926), .Q(text_in_r[103] ), .QN ());
DFFX1 text_in_r_reg[23] (.CK (clk), .D (n_3300), .Q (text_in_r[23]), .QN ());
DFFX1 text_in_r_reg[58] (.CK (clk), .D (n_3295), .Q (text_in_r[58]), .QN ());
DFFX1 text_in_r_reg[3] (.CK (clk), .D (n_3909), .Q (text_in_r[3] ),.QN ());
INVX1 g77519(.A (n_6293), .Y (n_8016));
NAND2X1 g74861(.A (n_6033), .B (n_27688), .Y (n_6291));
NAND3X1 g61182(.A (n_6286), .B (n_6289), .C (n_2848), .Y (n_13728));
OR2X1 g71488(.A (n_5832), .B (n_15894), .Y (n_6287));
NOR2X1 g61184(.A (n_6286), .B (n_6289), .Y (n_7860));
DFFX1 text_in_r_reg[118] (.CK (clk), .D (n_3617), .Q(text_in_r[118] ), .QN ());
INVX1 g76714(.A (n_6285), .Y (n_7610));
DFFX1 text_in_r_reg[59] (.CK (clk), .D (n_3402), .Q (text_in_r[59]), .QN ());
INVX1 g75231(.A (n_4891), .Y (n_7879));
NAND2X1 g74853(.A (n_3177), .B (n_26880), .Y (n_6283));
DFFX1 text_in_r_reg[96] (.CK (clk), .D (n_3948), .Q (text_in_r[96]), .QN ());
NAND2X1 g74382(.A (n_6281), .B (n_7201), .Y (n_6282));
INVX1 g75447(.A (n_6280), .Y (n_9077));
NOR2X1 g72994(.A (n_5774), .B (n_6279), .Y (n_7797));
NAND2X1 g72417(.A (n_12568), .B (n_6277), .Y (n_6278));
INVX1 g73779(.A (n_9774), .Y (n_6276));
DFFX1 text_in_r_reg[70] (.CK (clk), .D (n_3800), .Q (text_in_r[70]), .QN ());
OR2X1 g75229(.A (n_3163), .B (n_8090), .Y (n_6275));
NOR2X1 g72046(.A (n_4216), .B (n_4898), .Y (n_6274));
INVX1 g74368(.A (n_6268), .Y (n_6269));
NOR2X1 g71466(.A (n_5803), .B (n_5422), .Y (n_7161));
INVX1 g74846(.A (n_10181), .Y (n_6597));
NAND2X1 g74354(.A (n_4375), .B (n_2324), .Y (n_15460));
NAND2X2 g70192(.A (n_6265), .B (n_4825), .Y (n_7795));
NAND2X1 g74364(.A (n_6260), .B (n_6462), .Y (n_8243));
NOR2X1 g71460(.A (n_5915), .B (n_4598), .Y (n_7162));
NAND2X1 g73158(.A (n_4137), .B (n_3756), .Y (n_13269));
NAND2X1 g73156(.A (n_26890), .B (n_6185), .Y (n_10868));
NAND2X1 g74841(.A (n_6444), .B (n_7563), .Y (n_9073));
INVX1 g75405(.A (n_5331), .Y (n_6258));
INVX1 g70171(.A (n_7661), .Y (n_7381));
DFFX1 text_in_r_reg[51] (.CK (clk), .D (n_3660), .Q (text_in_r[51]), .QN ());
INVX1 g75514(.A (n_6261), .Y (n_7787));
NOR2X1 g77784(.A (n_7725), .B (n_8637), .Y (n_6255));
NOR2X1 g73150(.A (n_4481), .B (n_3920), .Y (n_6254));
NOR2X1 g74834(.A (n_6252), .B (n_4034), .Y (n_7782));
INVX2 g72670(.A (n_6249), .Y (n_6942));
NOR2X1 g70154(.A (n_6247), .B (n_12910), .Y (n_6248));
INVX1 g74345(.A (n_6368), .Y (n_6673));
AND2X1 g77740(.A (n_14589), .B (n_19414), .Y (n_12663));
OR2X1 g75573(.A (n_4732), .B (n_4973), .Y (n_6246));
INVX1 g75216(.A (n_6245), .Y (n_7778));
INVX1 g74814(.A (n_6243), .Y (n_6601));
INVX1 g76405(.A (ld_r), .Y (n_10226));
INVX1 g74820(.A (n_6239), .Y (n_10681));
INVX1 g73433(.A (n_6237), .Y (n_6238));
NAND2X2 g71423(.A (n_7032), .B (n_383), .Y (n_12399));
AND2X1 g77319(.A (n_8093), .B (n_2777), .Y (n_7955));
NAND2X1 g75328(.A (n_6234), .B (n_6153), .Y (n_6235));
NAND2X1 g71416(.A (n_7194), .B (n_6232), .Y (n_6233));
NOR2X1 g70128(.A (n_9442), .B (n_4650), .Y (n_7390));
INVX1 g74324(.A (n_4350), .Y (n_6679));
INVX1 g73736(.A (n_5951), .Y (n_6231));
INVX1 g74809(.A (n_4847), .Y (n_8978));
INVX1 g74806(.A (n_28132), .Y (n_9860));
NOR2X1 g74802(.A (n_5983), .B (n_28595), .Y (n_9336));
INVX1 g70986(.A (n_4569), .Y (n_9414));
INVX1 g75208(.A (n_6229), .Y (n_7769));
INVX1 g74797(.A (n_6227), .Y (n_6228));
INVX1 g70102(.A (n_4613), .Y (n_13532));
NAND2X1 g71396(.A (n_4695), .B (n_8865), .Y (n_7173));
NOR2X1 g70106(.A (n_27904), .B (n_4419), .Y (n_9349));
AND2X1 g70100(.A (n_4452), .B (n_6226), .Y (n_18347));
INVX1 g72776(.A (n_13118), .Y (n_9585));
CLKBUFX1 g74074(.A (n_6223), .Y (n_8250));
INVX1 g72382(.A (n_4507), .Y (n_6222));
AND2X1 g74790(.A (n_3307), .B (n_4764), .Y (n_6606));
NOR2X1 g75203(.A (n_4753), .B (n_6219), .Y (n_6220));
DFFX1 text_in_r_reg[92] (.CK (clk), .D (n_3495), .Q (text_in_r[92]), .QN ());
NAND4X1 g66027(.A (n_6219), .B (n_4846), .C (n_488), .D (n_3314), .Y(n_9593));
NAND2X1 g75202(.A (n_4038), .B (n_4113), .Y (n_6218));
NAND2X1 g75162(.A (n_4966), .B (n_4804), .Y (n_6536));
AND2X1 g77718(.A (n_11307), .B (n_282), .Y (n_6216));
INVX1 g74783(.A (n_6212), .Y (n_6213));
NAND2X1 g75190(.A (n_755), .B (n_3073), .Y (n_6529));
INVX1 g74779(.A (n_8837), .Y (n_6211));
INVX1 g77732(.A (n_6210), .Y (n_7742));
INVX2 g75569(.A (n_6209), .Y (n_8346));
OR2X1 g70069(.A (n_4957), .B (n_9264), .Y (n_7408));
INVX1 g74756(.A (n_7123), .Y (n_6614));
NAND4X1 g66244(.A (n_1424), .B (n_12559), .C (n_6805), .D (n_28340),.Y (n_6207));
NAND2X1 g74772(.A (n_3664), .B (n_27434), .Y (n_8137));
INVX1 g75721(.A (n_6206), .Y (n_9645));
NAND2X1 g70064(.A (n_4947), .B (n_27434), .Y (n_6205));
NOR2X1 g75185(.A (n_4842), .B (n_5990), .Y (n_6204));
NOR2X1 g71386(.A (n_4268), .B (n_5558), .Y (n_7178));
INVX1 g74767(.A (n_4783), .Y (n_6611));
AND2X1 g73108(.A (n_3254), .B (n_17912), .Y (n_6861));
NOR2X1 g73106(.A (n_5101), .B (n_26880), .Y (n_6202));
INVX1 g75178(.A (n_5318), .Y (n_6200));
NAND2X1 g75878(.A (n_3460), .B (n_6198), .Y (n_6448));
NOR2X1 g72182(.A (n_5593), .B (n_27990), .Y (n_6197));
NAND4X1 g66436(.A (n_2260), .B (n_6191), .C (n_3464), .D (n_3569), .Y(n_9561));
NAND2X2 g73687(.A (n_3925), .B (n_2260), .Y (n_9795));
DFFX1 text_in_r_reg[107] (.CK (clk), .D (n_3603), .Q(text_in_r[107] ), .QN ());
NAND2X1 g70037(.A (n_6188), .B (n_8679), .Y (n_6189));
NAND2X1 g75176(.A (n_4095), .B (n_6007), .Y (n_6532));
NAND2X1 g72356(.A (n_3326), .B (n_15507), .Y (n_20360));
INVX1 g73672(.A (n_5614), .Y (n_8916));
AOI21X1 g61524(.A0 (n_2849), .A1 (n_6289), .B0 (n_25126), .Y(n_6184));
NAND2X1 g74736(.A (n_5410), .B (n_1294), .Y (n_12778));
NAND2X1 g74734(.A (n_11350), .B (n_3823), .Y (n_6181));
NOR2X1 g73086(.A (n_5764), .B (n_7485), .Y (n_6179));
NOR2X1 g73084(.A (n_4379), .B (n_28375), .Y (n_6866));
NOR2X1 g71362(.A (n_5123), .B (n_8945), .Y (n_9370));
NOR2X1 g70012(.A (n_5925), .B (n_5922), .Y (n_6173));
INVX1 g74240(.A (n_6171), .Y (n_6689));
INVX1 g75549(.A (n_6169), .Y (n_6170));
INVX2 g74237(.A (n_7071), .Y (n_7705));
NAND2X1 g72676(.A (n_11816), .B (n_6166), .Y (n_6167));
DFFX1 text_in_r_reg[28] (.CK (clk), .D (n_3907), .Q (text_in_r[28]), .QN ());
NOR2X1 g73065(.A (n_6040), .B (n_3599), .Y (n_6162));
OR2X1 g69992(.A (n_28866), .B (n_3534), .Y (n_9380));
NOR2X1 g77694(.A (n_3038), .B (n_7410), .Y (n_6158));
NAND2X1 g73058(.A (n_4833), .B (n_2318), .Y (n_13418));
AND2X1 g75917(.A (n_17884), .B (n_6153), .Y (n_6154));
DFFX1 text_in_r_reg[77] (.CK (clk), .D (n_3354), .Q (text_in_r[77]), .QN ());
INVX1 g74224(.A (n_6149), .Y (n_28892));
NAND2X1 g73050(.A (n_6148), .B (n_12827), .Y (n_12198));
DFFX1 text_in_r_reg[1] (.CK (clk), .D (n_3732), .Q (text_in_r[1] ),.QN ());
NAND3X1 g67214(.A (n_6144), .B (n_3728), .C (n_4639), .Y (n_6145));
NAND2X1 g74725(.A (n_8363), .B (n_6142), .Y (n_6623));
DFFX1 text_in_r_reg[19] (.CK (clk), .D (n_3650), .Q (text_in_r[19]), .QN ());
NAND2X1 g72298(.A (n_10716), .B (n_16988), .Y (n_6141));
INVX1 g71324(.A (n_4687), .Y (n_7188));
NOR2X1 g69949(.A (n_4872), .B (n_4113), .Y (n_6140));
DFFX1 text_in_r_reg[56] (.CK (clk), .D (n_3543), .Q (text_in_r[56]), .QN ());
NOR2X1 g69932(.A (n_6133), .B (n_4618), .Y (n_6138));
OR2X1 g72294(.A (n_8295), .B (n_12105), .Y (n_6137));
DFFX1 text_in_r_reg[90] (.CK (clk), .D (n_3845), .Q (text_in_r[90]), .QN ());
NAND2X1 g72292(.A (n_6135), .B (n_12169), .Y (n_6136));
INVX1 g73586(.A (n_4835), .Y (n_8810));
OR2X1 g67468(.A (n_6134), .B (n_9527), .Y (n_9576));
INVX1 g73578(.A (n_5638), .Y (n_8811));
NOR2X1 g69923(.A (n_6133), .B (n_4883), .Y (n_7422));
OR2X1 g72632(.A (n_636), .B (n_27223), .Y (n_6950));
NAND2X1 g71298(.A (n_4291), .B (n_7410), .Y (n_9234));
OR2X1 g73606(.A (n_2707), .B (n_6534), .Y (n_7679));
INVX1 g74197(.A (n_6131), .Y (n_6132));
DFFX1 text_in_r_reg[69] (.CK (clk), .D (n_3404), .Q (text_in_r[69]), .QN ());
OR2X1 g72972(.A (n_5786), .B (n_5799), .Y (n_6884));
INVX1 g76372(.A (n_5843), .Y (n_25403));
OR2X1 g71234(.A (n_6031), .B (n_6988), .Y (n_9283));
INVX1 g72204(.A (n_6128), .Y (n_14964));
OR2X1 g72255(.A (n_4396), .B (n_8217), .Y (n_6127));
NAND2X1 g71286(.A (n_5835), .B (n_7658), .Y (n_6126));
NOR2X1 g73046(.A (n_4385), .B (n_6043), .Y (n_6122));
XOR2X1 g76132(.A (n_22567), .B (n_19908), .Y (n_6121));
NOR2X1 g69872(.A (n_596), .B (n_4435), .Y (n_6119));
INVX1 g69792(.A (n_14085), .Y (n_7444));
INVX1 g74635(.A (n_4523), .Y (n_6809));
INVX1 g77086(.A (n_27988), .Y (n_7095));
NOR2X1 g72938(.A (n_27896), .B (n_3820), .Y (n_6117));
DFFX1 text_in_r_reg[12] (.CK (clk), .D (n_3631), .Q (text_in_r[12]), .QN ());
OR2X1 g72930(.A (n_3992), .B (n_4173), .Y (n_6896));
INVX1 g74613(.A (n_6114), .Y (n_8894));
XOR2X1 g76218(.A (text_in_r[125] ), .B (n_497), .Y (n_6113));
INVX1 g76759(.A (n_6706), .Y (n_6853));
DFFX1 text_in_r_reg[85] (.CK (clk), .D (n_3245), .Q (text_in_r[85]), .QN ());
INVX1 g74702(.A (n_4488), .Y (n_9139));
DFFX1 text_in_r_reg[80] (.CK (clk), .D (n_3399), .Q (text_in_r[80]), .QN ());
DFFX1 text_in_r_reg[66] (.CK (clk), .D (n_3942), .Q (text_in_r[66]), .QN ());
NAND2X1 g72218(.A (n_4308), .B (n_11322), .Y (n_6108));
OR2X1 g68412(.A (n_6107), .B (n_12827), .Y (n_17139));
INVX1 g74510(.A (n_6105), .Y (n_6106));
DFFX1 text_in_r_reg[9] (.CK (clk), .D (n_3639), .Q (text_in_r[9] ),.QN ());
INVX1 g71231(.A (n_6104), .Y (n_13114));
NOR2X1 g72199(.A (n_6099), .B (n_1424), .Y (n_7013));
INVX4 g82284(.A (n_27493), .Y (n_16434));
OR2X1 g72692(.A (n_4307), .B (n_28375), .Y (n_7204));
INVX1 g78217(.A (n_6096), .Y (n_7698));
INVX1 g76407(.A (ld_r), .Y (n_8696));
INVX1 g76417(.A (n_6230), .Y (n_8520));
DFFX1 text_in_r_reg[53] (.CK (clk), .D (n_3770), .Q (text_in_r[53]), .QN ());
NAND2X1 g73419(.A (n_4142), .B (n_6997), .Y (n_6094));
NOR2X1 g72840(.A (n_5912), .B (n_7658), .Y (n_6916));
NOR2X1 g73024(.A (n_5910), .B (n_6092), .Y (n_6875));
DFFX1 text_in_r_reg[45] (.CK (clk), .D (n_3504), .Q (text_in_r[45]), .QN ());
OR2X1 g69744(.A (n_3438), .B (n_11307), .Y (n_12324));
DFFX1 text_in_r_reg[52] (.CK (clk), .D (n_3059), .Q (text_in_r[52]), .QN ());
XOR2X1 g68823(.A (n_1417), .B (n_2672), .Y (n_6088));
INVX1 g73438(.A (n_6086), .Y (n_6087));
XOR2X1 g68833(.A (n_980), .B (n_2297), .Y (n_6085));
INVX1 g71184(.A (n_6084), .Y (n_7206));
XOR2X1 g68839(.A (n_1341), .B (n_2540), .Y (n_6083));
INVX1 g72148(.A (n_6082), .Y (n_7602));
INVX1 g76396(.A (n_6067), .Y (n_7628));
NAND2X1 g77975(.A (n_1336), .B (n_29228), .Y (n_6081));
NOR2X1 g72142(.A (n_4979), .B (n_29228), .Y (n_6080));
NAND2X1 g62219(.A (n_3609), .B (n_6289), .Y (n_6079));
NAND2X1 g68979(.A (n_3764), .B (n_7601), .Y (n_7600));
NOR2X1 g68987(.A (n_6252), .B (n_4636), .Y (n_6078));
NOR2X1 g69010(.A (n_4478), .B (n_14807), .Y (n_6077));
NOR2X1 g69022(.A (n_28727), .B (n_2830), .Y (n_6076));
NAND4X1 g69031(.A (n_6008), .B (n_3081), .C (n_1244), .D (n_2323), .Y(n_9567));
NAND4X1 g69051(.A (n_3735), .B (n_3001), .C (n_4627), .D (n_3566), .Y(n_15085));
CLKBUFX2 g69056(.A (n_6074), .Y (n_7592));
AND2X1 g69092(.A (n_6015), .B (n_5922), .Y (n_9344));
NOR2X1 g69098(.A (n_4672), .B (n_5005), .Y (n_6072));
NAND2X1 g69101(.A (n_4703), .B (n_7601), .Y (n_6069));
NOR2X1 g69107(.A (n_383), .B (n_4486), .Y (n_7585));
INVX1 g69148(.A (n_6066), .Y (n_7579));
NAND2X1 g74248(.A (n_5365), .B (n_16414), .Y (n_6065));
NAND4X1 g69173(.A (n_7777), .B (n_3920), .C (n_2870), .D (n_23418),.Y (n_6064));
NOR2X1 g69181(.A (n_3234), .B (n_4550), .Y (n_7572));
NOR2X1 g69190(.A (n_6062), .B (n_9388), .Y (n_6063));
INVX1 g76375(.A (n_5112), .Y (n_25395));
NAND4X1 g69215(.A (n_3597), .B (n_5203), .C (n_7496), .D (n_2140), .Y(n_13243));
NAND2X1 g72827(.A (n_12624), .B (n_6058), .Y (n_6059));
NAND2X1 g69232(.A (n_4757), .B (n_4861), .Y (n_7557));
INVX1 g69233(.A (n_4242), .Y (n_9450));
NOR2X1 g69238(.A (n_5416), .B (n_4412), .Y (n_6057));
INVX1 g69240(.A (n_4647), .Y (n_9573));
NOR2X1 g71150(.A (n_27075), .B (n_6055), .Y (n_6056));
NAND2X1 g69244(.A (n_4215), .B (n_27434), .Y (n_14208));
INVX1 g76382(.A (n_5969), .Y (n_25415));
NAND2X1 g69252(.A (n_3326), .B (n_5922), .Y (n_7555));
NOR2X1 g69265(.A (n_4819), .B (n_6052), .Y (n_6053));
INVX1 g69278(.A (n_6050), .Y (n_7548));
INVX1 g69279(.A (n_6050), .Y (n_6051));
INVX1 g69283(.A (n_4644), .Y (n_11431));
NOR2X1 g69287(.A (n_28749), .B (n_4407), .Y (n_7547));
NOR2X1 g69289(.A (n_12827), .B (n_6062), .Y (n_19030));
NOR2X1 g69297(.A (n_4919), .B (n_4364), .Y (n_6048));
NAND2X1 g74070(.A (n_2875), .B (n_7636), .Y (n_6716));
NOR2X1 g69303(.A (n_4916), .B (n_4471), .Y (n_6047));
INVX2 g69307(.A (n_4365), .Y (n_9404));
NAND2X1 g69312(.A (n_5968), .B (n_11354), .Y (n_9303));
INVX4 g76385(.A (ld_r), .Y (n_25269));
NAND2X1 g69325(.A (n_4902), .B (n_7410), .Y (n_6046));
INVX1 g74114(.A (n_4380), .Y (n_8911));
NAND2X1 g69331(.A (n_3980), .B (n_2260), .Y (n_6045));
NOR2X1 g69335(.A (n_28616), .B (n_6043), .Y (n_6044));
NAND2X1 g69350(.A (n_5944), .B (n_6005), .Y (n_6042));
NAND2X1 g69363(.A (n_6232), .B (n_3301), .Y (n_7531));
NOR2X1 g71142(.A (n_6040), .B (n_7182), .Y (n_6041));
NOR2X1 g69387(.A (n_3999), .B (n_4882), .Y (n_6038));
NAND2X1 g73395(.A (n_3718), .B (n_6534), .Y (n_11861));
NOR2X1 g69398(.A (n_4715), .B (n_5643), .Y (n_7521));
NOR2X1 g69402(.A (n_5988), .B (n_7485), .Y (n_6036));
NOR2X1 g69407(.A (n_6034), .B (n_15712), .Y (n_6035));
NAND2X1 g74147(.A (n_2885), .B (n_352), .Y (n_6699));
NOR2X1 g69417(.A (n_28162), .B (n_6185), .Y (n_6880));
AND2X1 g75404(.A (n_2292), .B (n_6033), .Y (n_12747));
NOR2X1 g72102(.A (n_6031), .B (n_4391), .Y (n_6032));
NAND4X1 g69446(.A (n_8997), .B (n_1206), .C (n_8918), .D (n_2910), .Y(n_17725));
NAND2X1 g69455(.A (n_4853), .B (n_7485), .Y (n_13172));
NOR2X1 g72098(.A (n_4600), .B (n_4173), .Y (n_6028));
NOR2X1 g69459(.A (n_4430), .B (n_29275), .Y (n_7509));
AND2X1 g69467(.A (n_4771), .B (n_8865), .Y (n_6027));
NOR2X1 g69483(.A (n_4658), .B (n_5660), .Y (n_6026));
NAND2X1 g69485(.A (n_6025), .B (n_9342), .Y (n_9340));
NOR2X1 g69488(.A (n_5942), .B (n_3307), .Y (n_6024));
NAND2X1 g69489(.A (n_6025), .B (n_11312), .Y (n_9209));
NAND2X1 g69491(.A (n_6023), .B (n_11312), .Y (n_10937));
INVX1 g69495(.A (n_4511), .Y (n_7505));
AND2X1 g69501(.A (n_6004), .B (n_3301), .Y (n_7504));
NOR2X1 g69506(.A (n_4134), .B (n_6021), .Y (n_6022));
NOR2X1 g69518(.A (n_3277), .B (n_330), .Y (n_6020));
NAND2X1 g69523(.A (n_4914), .B (n_9342), .Y (n_11065));
OR2X1 g69525(.A (n_6018), .B (n_3307), .Y (n_19019));
AND2X1 g71130(.A (n_3726), .B (n_12827), .Y (n_7218));
NOR2X1 g69548(.A (n_4778), .B (n_3301), .Y (n_7494));
INVX1 g69550(.A (n_4634), .Y (n_11500));
AND2X1 g69561(.A (n_6015), .B (n_12827), .Y (n_11141));
INVX2 g69565(.A (n_4537), .Y (n_7489));
INVX1 g69571(.A (n_5862), .Y (n_17619));
NAND2X2 g69577(.A (n_4741), .B (n_6012), .Y (n_14126));
NAND2X1 g72084(.A (n_28402), .B (n_6011), .Y (n_7036));
INVX1 g69582(.A (n_4632), .Y (n_15245));
INVX1 g73381(.A (n_6010), .Y (n_8686));
NOR2X1 g69598(.A (n_5971), .B (n_6008), .Y (n_6009));
NOR2X1 g69601(.A (n_3349), .B (n_6007), .Y (n_7482));
AND2X1 g69623(.A (n_4701), .B (n_6005), .Y (n_6006));
NAND2X1 g69626(.A (n_6004), .B (n_12169), .Y (n_9348));
NOR2X1 g69633(.A (n_3920), .B (n_4727), .Y (n_6003));
DFFX1 text_in_r_reg[97] (.CK (clk), .D (n_3663), .Q (text_in_r[97]), .QN ());
NOR2X1 g69678(.A (n_5966), .B (n_11323), .Y (n_6001));
NOR2X1 g69681(.A (n_3306), .B (n_7777), .Y (n_7466));
DFFX1 text_in_r_reg[10] (.CK (clk), .D (n_3358), .Q (text_in_r[10]), .QN ());
NAND2X1 g69700(.A (n_7084), .B (n_11312), .Y (n_6000));
NOR2X1 g69702(.A (n_5795), .B (n_7158), .Y (n_17288));
NAND2X1 g69669(.A (n_4567), .B (n_7201), .Y (n_7470));
NAND2X1 g69723(.A (n_5997), .B (n_8679), .Y (n_5998));
NAND2X1 g69735(.A (n_4312), .B (n_2779), .Y (n_5996));
DFFX1 text_in_r_reg[34] (.CK (clk), .D (n_3680), .Q (text_in_r[34]), .QN ());
NOR2X1 g69761(.A (n_5381), .B (n_28162), .Y (n_5994));
NOR2X1 g69777(.A (n_4627), .B (n_4543), .Y (n_7450));
NAND2X1 g71109(.A (n_28724), .B (n_29269), .Y (n_5992));
NOR2X1 g69780(.A (n_4410), .B (n_8742), .Y (n_7447));
INVX2 g69785(.A (n_4708), .Y (n_9402));
NOR2X1 g72792(.A (n_5771), .B (n_5990), .Y (n_5991));
NOR2X1 g69826(.A (n_6997), .B (n_5988), .Y (n_5989));
NAND2X1 g69831(.A (n_5936), .B (n_9442), .Y (n_5986));
INVX1 g70764(.A (n_7634), .Y (n_7269));
NOR2X1 g69862(.A (n_4950), .B (n_4961), .Y (n_6443));
DFFX1 text_in_r_reg[110] (.CK (clk), .D (n_3636), .Q(text_in_r[110] ), .QN ());
OR2X1 g69876(.A (n_6144), .B (n_7410), .Y (n_17083));
NAND3X1 g69881(.A (n_28680), .B (n_5985), .C (n_11272), .Y (n_12718));
NOR2X1 g69889(.A (n_4107), .B (n_5983), .Y (n_5984));
NOR2X1 g69895(.A (n_27199), .B (n_6185), .Y (n_7432));
INVX1 g69897(.A (n_4706), .Y (n_7430));
INVX1 g69920(.A (n_4619), .Y (n_7424));
INVX1 g69937(.A (n_4718), .Y (n_7421));
NOR2X1 g69654(.A (n_4123), .B (n_28771), .Y (n_5982));
AND2X1 g69983(.A (n_4408), .B (n_7410), .Y (n_12637));
NAND2X1 g75773(.A (n_2724), .B (n_18785), .Y (n_5981));
AND2X1 g70002(.A (n_4184), .B (n_12559), .Y (n_5979));
NOR2X1 g70007(.A (n_27990), .B (n_4444), .Y (n_7703));
INVX1 g70008(.A (n_5976), .Y (n_5978));
NAND2X1 g71093(.A (n_6058), .B (n_11253), .Y (n_7719));
INVX1 g73374(.A (n_5975), .Y (n_8666));
OR2X1 g70082(.A (n_5974), .B (n_5151), .Y (n_13536));
NOR2X1 g70086(.A (n_3269), .B (n_8679), .Y (n_5973));
INVX1 g70093(.A (n_5972), .Y (n_17685));
INVX1 g70113(.A (n_4845), .Y (n_7395));
NOR2X1 g70116(.A (n_5971), .B (n_29102), .Y (n_14046));
NOR2X1 g72033(.A (n_6133), .B (n_5860), .Y (n_5970));
INVX1 g76380(.A (n_5969), .Y (n_25428));
NAND2X1 g70161(.A (n_6004), .B (n_16466), .Y (n_9309));
NAND2X1 g70168(.A (n_4345), .B (n_12760), .Y (n_9330));
NAND2X1 g70197(.A (n_5968), .B (n_2779), .Y (n_9328));
NOR2X1 g70201(.A (n_4559), .B (n_28398), .Y (n_7377));
INVX1 g70213(.A (n_4605), .Y (n_7373));
NOR2X1 g70223(.A (n_5966), .B (n_26880), .Y (n_5967));
NAND2X1 g70235(.A (n_3716), .B (n_636), .Y (n_12560));
NOR2X1 g70269(.A (n_4202), .B (n_6043), .Y (n_5963));
AND2X1 g70280(.A (n_5777), .B (n_6226), .Y (n_7355));
NOR2X1 g70287(.A (n_3456), .B (n_9368), .Y (n_7352));
NAND2X2 g70295(.A (n_6265), .B (n_12559), .Y (n_7347));
NAND2X1 g70311(.A (n_4462), .B (n_6790), .Y (n_5961));
NOR2X1 g70327(.A (n_4943), .B (n_9783), .Y (n_7337));
INVX1 g70338(.A (n_5958), .Y (n_5960));
INVX1 g73757(.A (n_5956), .Y (n_5957));
NOR2X1 g70349(.A (n_5990), .B (n_4692), .Y (n_7333));
NAND2X1 g70351(.A (n_3862), .B (n_4689), .Y (n_5955));
INVX1 g75852(.A (n_4046), .Y (n_6408));
INVX1 g73354(.A (n_6958), .Y (n_5953));
INVX1 g70378(.A (n_4593), .Y (n_9459));
NAND2X1 g72746(.A (n_4798), .B (n_12169), .Y (n_9217));
INVX1 g73735(.A (n_5951), .Y (n_9513));
NAND2X1 g78080(.A (n_3735), .B (n_11276), .Y (n_5950));
AND2X1 g70398(.A (n_4740), .B (n_8865), .Y (n_5949));
INVX1 g78076(.A (n_5946), .Y (n_5947));
NAND2X1 g70441(.A (n_5015), .B (n_4173), .Y (n_13152));
NOR2X1 g70447(.A (n_3981), .B (n_27904), .Y (n_5945));
NOR2X1 g70461(.A (n_5942), .B (n_9342), .Y (n_5943));
NAND4X1 g70468(.A (n_7658), .B (n_3307), .C (n_9202), .D (n_23422),.Y (n_5941));
NAND2X1 g70482(.A (n_3317), .B (n_9527), .Y (n_5939));
INVX1 g73675(.A (n_5937), .Y (n_5938));
NAND2X1 g70496(.A (n_5766), .B (n_9410), .Y (n_17115));
NOR2X1 g70501(.A (n_6303), .B (n_4465), .Y (n_7307));
NAND2X1 g70507(.A (n_5936), .B (n_29102), .Y (n_9200));
NOR2X1 g70511(.A (n_29140), .B (n_29256), .Y (n_7303));
INVX2 g70543(.A (n_4133), .Y (n_11031));
NAND2X1 g70557(.A (n_6232), .B (n_7410), .Y (n_5935));
NAND2X1 g70566(.A (n_5930), .B (n_27124), .Y (n_5934));
INVX1 g74094(.A (n_5932), .Y (n_13519));
INVX1 g73343(.A (n_5931), .Y (n_7294));
INVX2 g70609(.A (n_4180), .Y (n_9406));
NAND2X2 g70611(.A (n_5930), .B (n_28408), .Y (n_13137));
NOR2X1 g75144(.A (n_3029), .B (n_12469), .Y (n_5929));
INVX1 g75093(.A (n_4596), .Y (n_8127));
NOR2X1 g70619(.A (n_3017), .B (n_4441), .Y (n_7283));
DFFX1 text_in_r_reg[30] (.CK (clk), .D (n_3380), .Q (text_in_r[30]), .QN ());
INVX1 g70654(.A (n_5928), .Y (n_7278));
NOR2X1 g69594(.A (n_5925), .B (n_16480), .Y (n_5926));
NOR2X1 g69608(.A (n_5924), .B (n_4857), .Y (n_7481));
NAND2X1 g74083(.A (n_5923), .B (n_5922), .Y (n_6712));
INVX1 g70661(.A (n_9547), .Y (n_17465));
INVX1 g73332(.A (n_7813), .Y (n_5921));
NOR2X1 g72730(.A (n_4315), .B (n_7485), .Y (n_6751));
NOR2X1 g70732(.A (n_5787), .B (n_29256), .Y (n_5918));
INVX1 g75527(.A (n_4519), .Y (n_8863));
OR2X1 g71040(.A (n_4166), .B (n_9357), .Y (n_5917));
NOR2X1 g70781(.A (n_4260), .B (n_27365), .Y (n_6769));
NOR2X1 g70790(.A (n_5826), .B (n_7636), .Y (n_7264));
NOR2X1 g70806(.A (n_5768), .B (n_7366), .Y (n_5914));
NOR2X1 g70813(.A (n_383), .B (n_4788), .Y (n_5913));
NOR2X1 g70819(.A (n_5912), .B (n_7537), .Y (n_6811));
NOR2X1 g70829(.A (n_5910), .B (n_2318), .Y (n_5911));
NOR2X1 g70831(.A (n_4007), .B (n_7362), .Y (n_9355));
OR2X1 g70840(.A (n_8295), .B (n_6889), .Y (n_5907));
INVX1 g75140(.A (n_4241), .Y (n_9016));
NOR2X1 g70858(.A (n_5878), .B (n_6877), .Y (n_5906));
NAND2X1 g72716(.A (n_6277), .B (n_7593), .Y (n_6937));
OR2X1 g70902(.A (n_4025), .B (n_7410), .Y (n_9332));
INVX1 g73528(.A (n_4454), .Y (n_13177));
NOR2X1 g70949(.A (n_4255), .B (n_11323), .Y (n_7048));
NOR2X1 g70966(.A (n_4424), .B (n_9257), .Y (n_7243));
NAND2X1 g74080(.A (n_4776), .B (n_677), .Y (n_6714));
NAND2X1 g71008(.A (n_4285), .B (n_9527), .Y (n_9183));
NAND2X1 g71015(.A (n_2071), .B (n_6868), .Y (n_9211));
NOR2X1 g71026(.A (n_5047), .B (n_7331), .Y (n_5897));
NAND2X1 g71029(.A (n_17706), .B (n_5895), .Y (n_5896));
INVX1 g71053(.A (n_14324), .Y (n_19191));
INVX1 g71056(.A (n_4563), .Y (n_9389));
OR2X1 g75131(.A (n_3714), .B (n_26880), .Y (n_5894));
OR2X1 g69587(.A (n_7215), .B (n_5151), .Y (n_13688));
AND2X1 g71084(.A (n_2071), .B (n_8217), .Y (n_7227));
AND2X1 g71086(.A (n_5892), .B (n_27688), .Y (n_5893));
AND2X1 g71095(.A (n_27431), .B (n_9368), .Y (n_5891));
NAND2X1 g71101(.A (n_6166), .B (n_12019), .Y (n_7226));
NOR2X1 g71108(.A (n_5841), .B (n_8435), .Y (n_7221));
NAND2X1 g71111(.A (n_7617), .B (n_5887), .Y (n_5888));
OR2X1 g71112(.A (n_4730), .B (n_8865), .Y (n_5886));
NAND2X1 g71118(.A (n_4320), .B (n_15039), .Y (n_10905));
AND2X1 g71137(.A (n_4433), .B (n_12827), .Y (n_5885));
INVX1 g73399(.A (n_5884), .Y (n_6794));
INVX1 g75601(.A (n_6582), .Y (n_28319));
OR2X1 g71151(.A (n_4247), .B (n_11307), .Y (n_9212));
NOR2X1 g71157(.A (n_28131), .B (n_7728), .Y (n_5881));
NAND2X1 g72806(.A (n_27309), .B (n_5770), .Y (n_12429));
OR2X1 g71173(.A (n_5878), .B (n_8263), .Y (n_7207));
NAND2X1 g74068(.A (n_4100), .B (n_4925), .Y (n_8644));
INVX1 g71197(.A (n_4878), .Y (n_11422));
OR2X1 g75280(.A (n_3112), .B (n_6303), .Y (n_5875));
NAND2X1 g74670(.A (n_3101), .B (n_9691), .Y (n_5874));
INVX1 g71205(.A (n_4557), .Y (n_9472));
NOR2X1 g71211(.A (n_4669), .B (n_4490), .Y (n_11003));
NOR2X1 g71212(.A (n_7169), .B (n_14348), .Y (n_5872));
NAND2X1 g71213(.A (n_4458), .B (n_17912), .Y (n_5871));
NOR2X1 g71221(.A (n_3993), .B (n_27757), .Y (n_5870));
AND2X1 g74671(.A (n_3506), .B (n_4882), .Y (n_9078));
NOR2X1 g71264(.A (n_28859), .B (n_7266), .Y (n_5868));
NOR2X1 g71269(.A (n_5867), .B (n_9357), .Y (n_12246));
INVX4 g74038(.A (n_6415), .Y (n_10094));
CLKBUFX3 g71960(.A (n_5866), .Y (n_9285));
INVX1 g71310(.A (n_4731), .Y (n_9319));
NAND2X1 g71312(.A (n_4000), .B (n_7658), .Y (n_12187));
NOR2X1 g71334(.A (n_4739), .B (n_26276), .Y (n_5864));
NAND2X1 g71355(.A (n_12571), .B (n_5944), .Y (n_7723));
NOR2X1 g71383(.A (n_5800), .B (n_6462), .Y (n_5861));
NOR2X1 g71399(.A (n_5860), .B (n_2260), .Y (n_7172));
NOR2X1 g71441(.A (n_5741), .B (n_18320), .Y (n_7167));
AND2X1 g71450(.A (n_1497), .B (n_5857), .Y (n_5859));
OR2X1 g75839(.A (n_10607), .B (n_4884), .Y (n_5856));
NAND2X1 g71480(.A (n_4258), .B (n_5854), .Y (n_7160));
INVX1 g74064(.A (n_7440), .Y (n_11682));
INVX1 g71501(.A (n_4907), .Y (n_7157));
INVX1 g71504(.A (n_5853), .Y (n_17467));
INVX1 g71509(.A (n_7639), .Y (n_10794));
INVX1 g71515(.A (n_4534), .Y (n_18635));
NOR2X1 g71521(.A (n_4841), .B (n_6005), .Y (n_5852));
INVX1 g71525(.A (n_5850), .Y (n_5851));
NOR2X1 g71533(.A (n_28402), .B (n_4366), .Y (n_7146));
NOR2X1 g71932(.A (n_28131), .B (n_4391), .Y (n_5848));
NOR2X1 g71564(.A (n_4869), .B (n_17912), .Y (n_5846));
NAND2X1 g71569(.A (n_3683), .B (n_6868), .Y (n_12189));
NAND2X1 g71570(.A (n_6510), .B (n_5845), .Y (n_18061));
INVX1 g76379(.A (n_5969), .Y (n_25393));
INVX1 g76364(.A (n_5581), .Y (n_25422));
INVX1 g76381(.A (n_5969), .Y (n_25386));
INVX1 g71581(.A (n_7732), .Y (n_9333));
NAND2X1 g71585(.A (n_5833), .B (n_10452), .Y (n_14805));
INVX1 g76371(.A (n_5843), .Y (n_25382));
INVX1 g76370(.A (n_5843), .Y (n_25391));
NOR2X1 g71600(.A (n_5841), .B (n_11323), .Y (n_5842));
NAND2X1 g71621(.A (n_5839), .B (n_26491), .Y (n_7124));
NOR2X1 g71652(.A (n_4243), .B (n_1147), .Y (n_5838));
OR2X1 g71655(.A (n_16954), .B (n_11312), .Y (n_9504));
OR2X1 g71670(.A (n_2400), .B (n_5835), .Y (n_5837));
NAND2X1 g75508(.A (n_5834), .B (n_3017), .Y (n_8493));
NAND2X1 g70972(.A (n_3726), .B (n_6226), .Y (n_9350));
NOR2X1 g71692(.A (n_5832), .B (n_6219), .Y (n_7109));
NOR2X1 g71699(.A (n_3268), .B (n_5854), .Y (n_6499));
NAND2X1 g71714(.A (n_5828), .B (n_14757), .Y (n_5829));
OR2X1 g71718(.A (n_9220), .B (n_7410), .Y (n_9425));
NOR2X1 g71749(.A (n_5826), .B (n_367), .Y (n_5827));
NOR2X1 g71762(.A (n_26486), .B (n_28860), .Y (n_10791));
INVX1 g71768(.A (n_4526), .Y (n_14523));
OR2X1 g71770(.A (n_5823), .B (n_9474), .Y (n_9232));
OR2X1 g71773(.A (n_3302), .B (n_11385), .Y (n_5822));
NAND2X1 g71777(.A (n_5835), .B (n_3307), .Y (n_6723));
NOR2X1 g71920(.A (n_5820), .B (n_11731), .Y (n_14037));
INVX1 g71781(.A (n_4402), .Y (n_6732));
DFFX1 text_in_r_reg[104] (.CK (clk), .D (n_3624), .Q(text_in_r[104] ), .QN ());
NOR2X1 g71823(.A (n_1806), .B (n_6040), .Y (n_9315));
NOR2X1 g71831(.A (n_5802), .B (n_4598), .Y (n_7075));
INVX1 g71836(.A (n_5819), .Y (n_7073));
NAND2X1 g71844(.A (n_1416), .B (n_5944), .Y (n_12375));
NAND2X1 g71846(.A (n_12335), .B (n_5839), .Y (n_5818));
NOR2X1 g71856(.A (n_4642), .B (n_7127), .Y (n_9291));
INVX1 g71860(.A (n_7388), .Y (n_7068));
OR2X1 g71865(.A (n_4190), .B (n_5817), .Y (n_7066));
INVX1 g71870(.A (n_4503), .Y (n_7065));
INVX1 g75114(.A (n_5816), .Y (n_6549));
INVX2 g71893(.A (n_16621), .Y (n_5813));
AND2X1 g71901(.A (n_4369), .B (n_9819), .Y (n_5812));
DFFX1 text_in_r_reg[65] (.CK (clk), .D (n_3044), .Q (text_in_r[65]), .QN ());
INVX1 g71922(.A (n_11510), .Y (n_17491));
NAND2X1 g71933(.A (n_5810), .B (n_7201), .Y (n_12347));
NOR2X1 g71947(.A (n_4784), .B (n_9335), .Y (n_5809));
NOR2X1 g71951(.A (n_4886), .B (n_9264), .Y (n_5808));
NAND2X1 g71974(.A (n_5807), .B (n_5799), .Y (n_12172));
NAND2X1 g71979(.A (n_4475), .B (n_12019), .Y (n_5806));
INVX1 g70952(.A (n_5805), .Y (n_7245));
INVX1 g71995(.A (n_7726), .Y (n_9260));
OR2X1 g72001(.A (n_5803), .B (n_8878), .Y (n_9193));
OR2X1 g72013(.A (n_5802), .B (n_6185), .Y (n_9531));
NOR2X1 g71900(.A (n_5800), .B (n_5799), .Y (n_5801));
INVX1 g72025(.A (n_12734), .Y (n_19207));
INVX1 g72027(.A (n_7759), .Y (n_5798));
NOR2X1 g72037(.A (n_4164), .B (n_5854), .Y (n_7044));
NAND2X1 g72059(.A (n_4213), .B (n_2655), .Y (n_7416));
INVX1 g72065(.A (n_11449), .Y (n_17477));
OR2X1 g72089(.A (n_5719), .B (n_7498), .Y (n_11461));
NAND2X1 g72093(.A (n_5895), .B (n_29228), .Y (n_7035));
OR2X1 g69465(.A (n_5795), .B (n_11312), .Y (n_5796));
NOR2X1 g72113(.A (n_4145), .B (n_11312), .Y (n_5792));
NOR2X1 g72115(.A (n_5616), .B (n_2260), .Y (n_5791));
NAND2X1 g72119(.A (n_2357), .B (n_3365), .Y (n_7030));
NOR2X1 g69522(.A (n_5925), .B (n_8878), .Y (n_7499));
AND2X1 g72151(.A (n_5788), .B (n_16434), .Y (n_5789));
NOR2X1 g72159(.A (n_5787), .B (n_17260), .Y (n_7020));
INVX1 g72170(.A (n_4517), .Y (n_7786));
OR2X1 g72195(.A (n_5786), .B (n_29065), .Y (n_16713));
INVX1 g73498(.A (n_4570), .Y (n_8687));
NOR2X1 g72209(.A (n_16954), .B (n_13466), .Y (n_5784));
NOR2X1 g70934(.A (n_4467), .B (n_5413), .Y (n_5783));
NAND2X1 g73111(.A (n_4801), .B (n_7496), .Y (n_5781));
NAND2X1 g72264(.A (n_7032), .B (n_11731), .Y (n_5780));
NAND2X2 g72273(.A (n_5778), .B (n_5777), .Y (n_5779));
NAND2X1 g72291(.A (n_1928), .B (n_5833), .Y (n_10873));
INVX1 g72301(.A (n_5775), .Y (n_5776));
NOR2X1 g72310(.A (n_5774), .B (n_7331), .Y (n_7000));
NAND2X1 g72327(.A (n_9170), .B (n_4222), .Y (n_14309));
NAND2X1 g73081(.A (n_28724), .B (n_6419), .Y (n_7709));
OR2X1 g72345(.A (n_5771), .B (n_1942), .Y (n_7354));
NAND2X1 g72348(.A (n_5770), .B (n_28757), .Y (n_9363));
NOR2X1 g70846(.A (n_5768), .B (n_14055), .Y (n_5769));
INVX1 g71876(.A (n_5767), .Y (n_7064));
INVX1 g74649(.A (n_4518), .Y (n_8503));
OR2X1 g72373(.A (n_5725), .B (n_9118), .Y (n_6993));
NAND2X1 g70915(.A (n_12836), .B (n_5766), .Y (n_7252));
NAND2X1 g72384(.A (n_5733), .B (n_9388), .Y (n_5765));
NOR2X1 g72410(.A (n_5764), .B (n_18266), .Y (n_6985));
NAND2X1 g75797(.A (n_2042), .B (n_15039), .Y (n_5763));
NAND2X1 g72415(.A (n_2485), .B (n_5770), .Y (n_7796));
INVX1 g74156(.A (n_5761), .Y (n_5762));
INVX1 g72426(.A (n_5759), .Y (n_5760));
AND2X1 g72429(.A (n_3365), .B (n_11385), .Y (n_6982));
NAND2X1 g72445(.A (n_4602), .B (n_9388), .Y (n_7847));
NAND2X1 g72447(.A (n_4875), .B (n_3604), .Y (n_12768));
NOR2X1 g69478(.A (n_4728), .B (n_28381), .Y (n_5755));
INVX1 g72458(.A (n_4505), .Y (n_17508));
NAND2X1 g72467(.A (n_5807), .B (n_18074), .Y (n_5753));
NOR2X1 g72489(.A (n_1930), .B (n_5942), .Y (n_9469));
NAND2X1 g72493(.A (n_4017), .B (n_5795), .Y (n_5752));
INVX1 g69472(.A (n_5751), .Y (n_7507));
INVX1 g75481(.A (n_5749), .Y (n_5750));
INVX1 g72520(.A (n_5744), .Y (n_5745));
NAND2X1 g72561(.A (n_5770), .B (n_6790), .Y (n_16421));
NOR2X1 g72611(.A (n_4553), .B (n_3348), .Y (n_5743));
OR2X1 g72622(.A (n_5741), .B (n_9335), .Y (n_6943));
NOR2X1 g72634(.A (n_4343), .B (n_6226), .Y (n_5740));
OAI21X1 g75963(.A0 (n_4721), .A1 (n_2035), .B0 (n_2461), .Y (n_5738));
NOR2X1 g72689(.A (n_5735), .B (n_7685), .Y (n_5736));
NOR2X1 g72699(.A (n_28408), .B (n_5135), .Y (n_5734));
NAND2X2 g72734(.A (n_5733), .B (n_5151), .Y (n_11620));
NAND2X2 g69442(.A (n_4585), .B (n_28757), .Y (n_5731));
NOR2X1 g72771(.A (n_27893), .B (n_27896), .Y (n_5730));
OAI21X1 g75961(.A0 (n_27124), .A1 (n_28780), .B0 (n_5386), .Y(n_5728));
NOR2X1 g72782(.A (n_5725), .B (n_17500), .Y (n_5726));
OR2X1 g72788(.A (n_4867), .B (n_11312), .Y (n_16586));
INVX1 g72793(.A (n_5723), .Y (n_5724));
NOR2X1 g74642(.A (n_4282), .B (n_7563), .Y (n_5722));
NOR2X1 g72823(.A (n_11322), .B (n_4163), .Y (n_7554));
INVX2 g75766(.A (n_5721), .Y (n_6461));
NOR2X1 g72855(.A (n_3234), .B (n_4967), .Y (n_6915));
AND2X1 g72856(.A (n_4986), .B (n_6226), .Y (n_14534));
NAND2X1 g72871(.A (n_5810), .B (n_7607), .Y (n_9345));
INVX1 g75861(.A (n_4484), .Y (n_8780));
NOR2X1 g72875(.A (n_5719), .B (n_28692), .Y (n_6910));
INVX1 g72879(.A (n_7717), .Y (n_9258));
OR2X1 g72899(.A (n_5716), .B (n_20325), .Y (n_5717));
NAND2X1 g72909(.A (n_5857), .B (n_9118), .Y (n_6900));
INVX1 g72913(.A (n_5715), .Y (n_7473));
OAI21X1 g75956(.A0 (n_28757), .A1 (n_4082), .B0 (n_4980), .Y(n_5714));
NAND2X1 g72954(.A (n_4273), .B (n_28375), .Y (n_5712));
NOR2X1 g72877(.A (n_4269), .B (n_7331), .Y (n_5711));
NOR2X1 g73001(.A (n_5484), .B (n_1942), .Y (n_5709));
AND2X1 g73009(.A (n_9844), .B (n_3829), .Y (n_5708));
INVX1 g73015(.A (n_7624), .Y (n_7668));
NAND2X1 g73027(.A (n_4811), .B (n_7496), .Y (n_6874));
NOR2X1 g72545(.A (n_5435), .B (n_7658), .Y (n_5707));
OR2X1 g73062(.A (n_5705), .B (n_5704), .Y (n_5706));
NOR2X1 g73097(.A (n_4167), .B (n_27990), .Y (n_11076));
OR2X1 g73101(.A (n_3829), .B (n_17912), .Y (n_29302));
NOR2X1 g73123(.A (n_4960), .B (n_29244), .Y (n_6858));
AND2X1 g73151(.A (n_3707), .B (n_9527), .Y (n_5697));
NAND2X1 g73159(.A (n_5833), .B (n_6977), .Y (n_9564));
OR2X1 g73175(.A (n_5694), .B (n_12169), .Y (n_7807));
OR2X1 g73206(.A (n_5692), .B (n_5691), .Y (n_5693));
NAND2X1 g73213(.A (n_2914), .B (n_5766), .Y (n_12643));
NOR2X1 g69396(.A (n_4688), .B (n_27990), .Y (n_5690));
INVX1 g70826(.A (n_5689), .Y (n_9435));
NOR2X1 g75449(.A (n_3203), .B (n_26880), .Y (n_5688));
AOI21X1 g73300(.A0 (n_15473), .A1 (n_5236), .B0 (n_3291), .Y(n_5687));
INVX1 g73311(.A (n_9927), .Y (n_7235));
INVX1 g72595(.A (n_5686), .Y (n_6819));
INVX1 g73319(.A (n_5684), .Y (n_5685));
INVX1 g73325(.A (n_5681), .Y (n_5682));
NAND2X1 g73328(.A (n_5665), .B (n_7438), .Y (n_8404));
NAND2X1 g73329(.A (n_4492), .B (n_10389), .Y (n_5680));
INVX1 g73335(.A (n_6842), .Y (n_8378));
INVX1 g73349(.A (n_5677), .Y (n_5678));
INVX1 g73359(.A (n_5675), .Y (n_9053));
INVX2 g73371(.A (n_5674), .Y (n_7800));
INVX1 g73392(.A (n_5671), .Y (n_9018));
INVX1 g73414(.A (n_5667), .Y (n_5668));
NAND2X1 g73417(.A (n_5665), .B (n_12019), .Y (n_13855));
INVX1 g73441(.A (n_5663), .Y (n_5664));
INVX1 g73448(.A (n_5662), .Y (n_9522));
NAND2X1 g73459(.A (n_4748), .B (n_5660), .Y (n_5661));
INVX1 g73460(.A (n_5657), .Y (n_5659));
INVX1 g73467(.A (n_6102), .Y (n_8290));
INVX1 g73472(.A (n_4460), .Y (n_8296));
NAND2X1 g75685(.A (n_3823), .B (n_1424), .Y (n_5656));
INVX1 g73487(.A (n_7290), .Y (n_5653));
INVX1 g73491(.A (n_5650), .Y (n_5652));
NAND2X1 g74036(.A (n_4939), .B (n_27990), .Y (n_6725));
INVX1 g73509(.A (n_5646), .Y (n_9020));
INVX1 g73514(.A (n_4455), .Y (n_9804));
NAND2X1 g73525(.A (n_4027), .B (n_4568), .Y (n_7650));
INVX1 g73526(.A (n_4697), .Y (n_9552));
INVX1 g73534(.A (n_5644), .Y (n_8756));
INVX1 g73541(.A (n_4451), .Y (n_8611));
NAND2X1 g71808(.A (n_4301), .B (n_5643), .Y (n_7079));
INVX1 g73549(.A (n_7120), .Y (n_8362));
INVX2 g73561(.A (n_5642), .Y (n_9037));
OR2X1 g75082(.A (n_28485), .B (n_11276), .Y (n_5641));
NOR2X1 g69356(.A (n_4721), .B (n_3991), .Y (n_7532));
NAND2X1 g72592(.A (n_4911), .B (n_14624), .Y (n_5634));
INVX2 g73610(.A (n_7114), .Y (n_8664));
INVX1 g73617(.A (n_6164), .Y (n_5631));
INVX1 g75762(.A (n_3979), .Y (n_6919));
INVX1 g73628(.A (n_12291), .Y (n_5630));
INVX1 g74164(.A (n_5628), .Y (n_5629));
INVX1 g73636(.A (n_5625), .Y (n_5626));
INVX1 g73648(.A (n_4436), .Y (n_8380));
NAND2X1 g75942(.A (n_5620), .B (n_3145), .Y (n_5621));
INVX1 g73658(.A (n_5618), .Y (n_5619));
NOR2X1 g71802(.A (n_5616), .B (n_6191), .Y (n_7081));
INVX4 g73683(.A (n_5613), .Y (n_8709));
NAND2X2 g75442(.A (n_5612), .B (n_28792), .Y (n_8253));
NAND2X1 g73692(.A (n_4955), .B (n_3632), .Y (n_5611));
CLKBUFX1 g73701(.A (n_5609), .Y (n_15636));
NAND2X1 g73704(.A (n_4023), .B (n_5413), .Y (n_5608));
OR2X1 g73713(.A (n_3083), .B (n_8997), .Y (n_6773));
INVX1 g73718(.A (n_5605), .Y (n_5607));
NOR2X1 g73721(.A (n_2742), .B (n_11312), .Y (n_5603));
INVX1 g73727(.A (n_4856), .Y (n_11662));
OR2X1 g71798(.A (n_4978), .B (n_28427), .Y (n_7082));
INVX1 g73739(.A (n_5602), .Y (n_9004));
INVX1 g73741(.A (n_4850), .Y (n_14855));
AND2X1 g75940(.A (n_5600), .B (n_6442), .Y (n_5601));
OR2X1 g73743(.A (n_3097), .B (n_7593), .Y (n_10931));
INVX1 g73744(.A (n_5599), .Y (n_11078));
INVX1 g75433(.A (n_27897), .Y (n_6492));
INVX1 g73760(.A (n_4423), .Y (n_13730));
NOR2X1 g70756(.A (n_5593), .B (n_29269), .Y (n_5594));
INVX1 g73771(.A (n_6266), .Y (n_5591));
INVX1 g74030(.A (n_5590), .Y (n_6727));
INVX1 g73790(.A (n_5588), .Y (n_5589));
INVX1 g73793(.A (n_5585), .Y (n_5586));
INVX1 g75732(.A (n_4170), .Y (n_8809));
INVX1 g76366(.A (n_5581), .Y (n_25418));
INVX1 g74626(.A (n_5576), .Y (n_8490));
INVX1 g73824(.A (n_5574), .Y (n_5575));
INVX1 g73832(.A (n_5571), .Y (n_8931));
OR2X1 g73835(.A (n_25746), .B (n_27365), .Y (n_10856));
NAND2X1 g73840(.A (n_27072), .B (n_29244), .Y (n_11745));
NOR2X1 g73851(.A (n_2594), .B (n_12019), .Y (n_6760));
INVX1 g73866(.A (n_6989), .Y (n_5569));
INVX2 g76367(.A (n_5581), .Y (n_25305));
INVX1 g73873(.A (n_5567), .Y (n_5568));
NAND2X1 g75458(.A (n_1985), .B (n_17864), .Y (n_5563));
CLKBUFX3 g73921(.A (n_5560), .Y (n_6748));
NAND2X1 g73939(.A (n_3187), .B (n_5558), .Y (n_8172));
INVX1 g73953(.A (n_4102), .Y (n_6744));
INVX1 g73961(.A (n_5554), .Y (n_6740));
NOR2X1 g73981(.A (n_4072), .B (n_29244), .Y (n_5550));
INVX1 g73982(.A (n_4400), .Y (n_8343));
INVX1 g73987(.A (n_5548), .Y (n_9058));
NAND2X1 g73989(.A (n_6313), .B (n_5546), .Y (n_5547));
NOR2X1 g73990(.A (n_4076), .B (n_6997), .Y (n_9463));
DFFX1 text_in_r_reg[79] (.CK (clk), .D (n_3748), .Q (text_in_r[79]), .QN ());
INVX1 g74003(.A (n_5350), .Y (n_5545));
INVX1 g74008(.A (n_5543), .Y (n_5544));
INVX1 g74014(.A (n_5541), .Y (n_5542));
OR2X1 g74025(.A (n_3454), .B (n_9691), .Y (n_5540));
INVX1 g74031(.A (n_5590), .Y (n_29385));
INVX1 g70746(.A (n_7708), .Y (n_11412));
AND2X1 g69324(.A (n_5968), .B (n_379), .Y (n_9281));
INVX1 g74051(.A (n_4112), .Y (n_8070));
NOR2X1 g72579(.A (n_7169), .B (n_28404), .Y (n_5538));
NAND2X1 g74053(.A (n_3963), .B (n_9084), .Y (n_5537));
NAND2X1 g74057(.A (n_4070), .B (n_26887), .Y (n_5536));
DFFX1 text_in_r_reg[7] (.CK (clk), .D (n_3343), .Q (text_in_r[7] ),.QN ());
NAND2X1 g74096(.A (n_3581), .B (n_5530), .Y (n_5531));
INVX1 g74110(.A (n_5528), .Y (n_5529));
NAND2X1 g69316(.A (n_5766), .B (n_27365), .Y (n_5527));
INVX1 g74117(.A (n_5525), .Y (n_6703));
INVX1 g74135(.A (n_4778), .Y (n_8308));
INVX1 g74139(.A (n_5521), .Y (n_5522));
NAND2X1 g74142(.A (n_3984), .B (n_5643), .Y (n_6701));
NAND2X1 g74145(.A (n_26483), .B (n_27365), .Y (n_7619));
INVX1 g74149(.A (n_14386), .Y (n_6698));
NAND2X1 g74161(.A (n_4762), .B (n_3920), .Y (n_8603));
INVX1 g74163(.A (n_5628), .Y (n_7641));
INVX1 g74173(.A (n_7164), .Y (n_5517));
INVX1 g74179(.A (n_4700), .Y (n_8954));
NAND2X1 g74181(.A (n_5516), .B (n_5218), .Y (n_12607));
NAND2X1 g75930(.A (n_5778), .B (n_5509), .Y (n_14556));
NAND2X1 g70736(.A (n_2071), .B (n_7182), .Y (n_5514));
INVX1 g74195(.A (n_12517), .Y (n_5513));
NAND2X1 g74199(.A (n_5511), .B (n_17414), .Y (n_5512));
INVX1 g74200(.A (n_7615), .Y (n_5510));
NOR2X1 g74202(.A (n_3077), .B (n_7728), .Y (n_8169));
NAND2X1 g74219(.A (n_5509), .B (n_4882), .Y (n_7683));
NAND2X1 g74220(.A (n_2424), .B (n_5558), .Y (n_5508));
INVX1 g74223(.A (n_6149), .Y (n_10732));
INVX1 g74242(.A (n_5505), .Y (n_5507));
NOR2X1 g74245(.A (n_3686), .B (n_5085), .Y (n_5504));
NAND2X1 g74247(.A (n_4021), .B (n_1147), .Y (n_6687));
INVX1 g74256(.A (n_7210), .Y (n_8254));
INVX1 g74259(.A (n_4489), .Y (n_8682));
NAND2X1 g74267(.A (n_3297), .B (n_4113), .Y (n_7722));
NOR2X1 g74269(.A (n_5502), .B (n_6185), .Y (n_7755));
NAND2X1 g74279(.A (n_4776), .B (n_2318), .Y (n_6684));
INVX2 g74281(.A (n_4036), .Y (n_9101));
INVX1 g74287(.A (n_5495), .Y (n_5496));
INVX2 g74295(.A (n_5494), .Y (n_7746));
INVX2 g74305(.A (n_5493), .Y (n_7763));
NOR2X1 g74315(.A (n_4829), .B (n_8997), .Y (n_5492));
INVX1 g74317(.A (n_4844), .Y (n_5491));
OR2X1 g74319(.A (n_29357), .B (n_4898), .Y (n_5490));
INVX4 g74341(.A (n_7549), .Y (n_8729));
NOR2X1 g72572(.A (n_5484), .B (n_5483), .Y (n_5485));
INVX1 g76360(.A (n_4329), .Y (n_13768));
OR2X1 g74377(.A (n_1599), .B (n_12559), .Y (n_5477));
INVX1 g74380(.A (n_5475), .Y (n_5476));
INVX1 g74385(.A (n_4897), .Y (n_6670));
INVX1 g74395(.A (n_7185), .Y (n_5474));
AND2X1 g74406(.A (n_3867), .B (n_6805), .Y (n_5472));
INVX1 g74412(.A (n_7299), .Y (n_6661));
INVX1 g76356(.A (n_5114), .Y (n_13846));
NAND2X1 g74422(.A (n_14667), .B (n_5370), .Y (n_5471));
NOR2X1 g70720(.A (n_4839), .B (n_5983), .Y (n_5470));
INVX1 g74437(.A (n_5469), .Y (n_7830));
NAND2X1 g74440(.A (n_27439), .B (n_5799), .Y (n_5468));
NAND2X1 g74441(.A (n_3197), .B (n_17500), .Y (n_5467));
INVX1 g74454(.A (n_6097), .Y (n_5462));
INVX1 g74469(.A (n_4335), .Y (n_6654));
NAND2X1 g74617(.A (n_5457), .B (n_6534), .Y (n_5458));
INVX1 g74476(.A (n_5455), .Y (n_5456));
INVX1 g74479(.A (n_5454), .Y (n_14364));
NAND2X1 g75926(.A (n_10127), .B (n_2818), .Y (n_6671));
NAND2X2 g74487(.A (n_3831), .B (n_28459), .Y (n_8561));
INVX1 g74489(.A (n_27594), .Y (n_8441));
OR2X1 g71755(.A (n_9293), .B (n_11307), .Y (n_9465));
INVX1 g74493(.A (n_6974), .Y (n_8794));
INVX1 g74499(.A (n_5452), .Y (n_5453));
NAND2X1 g74666(.A (n_12827), .B (n_5447), .Y (n_5448));
NOR2X1 g74518(.A (n_3055), .B (n_383), .Y (n_5446));
INVX1 g74519(.A (n_5443), .Y (n_5444));
INVX1 g74022(.A (n_4393), .Y (n_6728));
OR2X1 g74537(.A (n_5441), .B (n_18785), .Y (n_5442));
INVX1 g74540(.A (n_4316), .Y (n_8834));
INVX1 g74549(.A (n_5439), .Y (n_5440));
INVX1 g75848(.A (n_4601), .Y (n_8788));
NOR2X1 g71754(.A (n_5435), .B (n_7537), .Y (n_5436));
INVX1 g74561(.A (n_4136), .Y (n_6409));
AND2X1 g69270(.A (n_4561), .B (n_12827), .Y (n_7551));
INVX1 g74585(.A (n_4922), .Y (n_6477));
NOR2X1 g74587(.A (n_29214), .B (n_5422), .Y (n_8556));
INVX1 g74601(.A (n_5430), .Y (n_8392));
INVX1 g74619(.A (n_5427), .Y (n_5428));
AND2X1 g74628(.A (n_2719), .B (n_29256), .Y (n_5425));
NAND2X1 g74016(.A (n_3150), .B (n_8090), .Y (n_5424));
NAND2X1 g69260(.A (n_5777), .B (n_5422), .Y (n_5423));
INVX1 g74643(.A (n_5420), .Y (n_5421));
CLKBUFX1 g74647(.A (n_5419), .Y (n_8425));
NOR2X1 g71730(.A (n_4852), .B (n_27371), .Y (n_5418));
INVX1 g74657(.A (n_4389), .Y (n_7027));
NOR2X1 g71368(.A (n_4836), .B (n_5416), .Y (n_5417));
NAND2X1 g74667(.A (n_1791), .B (n_17260), .Y (n_5415));
NAND2X1 g74669(.A (n_5344), .B (n_14484), .Y (n_5414));
NOR2X1 g74604(.A (n_4736), .B (n_5413), .Y (n_8524));
NAND2X1 g75414(.A (n_4671), .B (n_3338), .Y (n_8284));
NAND2X1 g74685(.A (n_4724), .B (n_379), .Y (n_8218));
INVX1 g74687(.A (n_5411), .Y (n_7429));
NAND2X2 g74691(.A (n_4770), .B (n_5924), .Y (n_6633));
NAND2X1 g74697(.A (n_4849), .B (n_5410), .Y (n_14074));
NOR2X1 g71742(.A (n_4344), .B (n_6005), .Y (n_7093));
INVX1 g75708(.A (n_4171), .Y (n_8820));
NAND2X1 g74731(.A (n_9415), .B (n_1942), .Y (n_7757));
INVX1 g75470(.A (n_4491), .Y (n_6491));
INVX1 g74749(.A (n_5408), .Y (n_8470));
NOR2X1 g74762(.A (n_5404), .B (n_14866), .Y (n_5405));
INVX1 g78015(.A (n_5403), .Y (n_8101));
OR2X1 g71734(.A (n_3033), .B (n_9527), .Y (n_5402));
INVX1 g74769(.A (n_10676), .Y (n_5400));
INVX1 g74773(.A (n_5399), .Y (n_8879));
INVX1 g74775(.A (n_4796), .Y (n_5398));
NOR2X1 g74777(.A (n_3034), .B (n_5799), .Y (n_5397));
INVX1 g74785(.A (n_5396), .Y (n_8778));
INVX1 g74791(.A (n_5394), .Y (n_28843));
INVX1 g74799(.A (n_5393), .Y (n_14361));
NAND2X1 g75921(.A (n_7803), .B (n_2401), .Y (n_16488));
INVX1 g74825(.A (n_6907), .Y (n_5389));
INVX1 g74838(.A (n_7145), .Y (n_5388));
NOR3X1 g74843(.A (n_596), .B (n_5085), .C (n_28271), .Y (n_6598));
OR2X1 g74848(.A (n_5386), .B (n_28375), .Y (n_5387));
NAND2X1 g74852(.A (n_3141), .B (n_8945), .Y (n_5385));
NAND2X1 g74855(.A (n_5383), .B (n_10031), .Y (n_8321));
NAND2X1 g74857(.A (n_4893), .B (n_6988), .Y (n_8438));
NAND2X1 g74859(.A (n_5204), .B (n_6790), .Y (n_6593));
NOR2X1 g78018(.A (n_28375), .B (n_27718), .Y (n_19964));
NAND2X2 g74885(.A (n_3257), .B (n_5381), .Y (n_5382));
OR2X1 g74892(.A (n_2785), .B (n_3301), .Y (n_5380));
INVX1 g74895(.A (n_7452), .Y (n_5378));
INVX1 g74909(.A (n_5375), .Y (n_7844));
NAND2X1 g72554(.A (n_6510), .B (n_6188), .Y (n_5374));
INVX1 g74917(.A (n_5373), .Y (n_9511));
NAND2X1 g74931(.A (n_4773), .B (n_28733), .Y (n_8951));
NAND2X1 g74938(.A (n_5370), .B (n_28692), .Y (n_5371));
AND2X1 g74941(.A (n_379), .B (n_2743), .Y (n_6577));
NAND2X1 g74948(.A (n_5369), .B (n_5447), .Y (n_20526));
NOR2X1 g74951(.A (n_5368), .B (n_28375), .Y (n_6574));
INVX1 g74953(.A (n_5367), .Y (n_6366));
NAND2X1 g74956(.A (n_5365), .B (n_28375), .Y (n_5366));
INVX1 g74983(.A (n_7296), .Y (n_6397));
INVX1 g74985(.A (n_5357), .Y (n_5358));
INVX1 g75003(.A (n_4128), .Y (n_6417));
INVX1 g74086(.A (n_4384), .Y (n_6711));
INVX1 g75007(.A (n_5355), .Y (n_25665));
OR2X1 g75013(.A (n_3065), .B (n_8968), .Y (n_5354));
INVX1 g75014(.A (n_4253), .Y (n_8635));
NAND2X1 g75058(.A (n_4699), .B (n_8452), .Y (n_5346));
NAND2X1 g75700(.A (n_5344), .B (n_18320), .Y (n_5345));
INVX2 g75067(.A (n_5343), .Y (n_8367));
INVX1 g75070(.A (n_5340), .Y (n_5341));
INVX1 g74674(.A (n_4572), .Y (n_7397));
NOR2X1 g75077(.A (n_2487), .B (n_27987), .Y (n_11435));
CLKBUFX1 g75089(.A (n_5337), .Y (n_8491));
INVX1 g75125(.A (n_7417), .Y (n_5334));
NAND2X1 g75133(.A (n_5612), .B (n_28375), .Y (n_6544));
INVX1 g75134(.A (n_4567), .Y (n_5333));
NAND2X1 g75145(.A (n_4800), .B (n_5329), .Y (n_5330));
DFFX1 text_in_r_reg[82] (.CK (clk), .D (n_3625), .Q (text_in_r[82]), .QN ());
INVX1 g75152(.A (n_5326), .Y (n_5327));
INVX1 g77960(.A (n_5323), .Y (n_5324));
INVX1 g75156(.A (n_7008), .Y (n_5322));
INVX1 g70643(.A (n_4235), .Y (n_9509));
NOR2X1 g75173(.A (n_4114), .B (n_596), .Y (n_5319));
NAND2X1 g75181(.A (n_14113), .B (n_5316), .Y (n_5317));
AND2X1 g75188(.A (n_2875), .B (n_14055), .Y (n_5315));
INVX1 g75191(.A (n_12756), .Y (n_5313));
INVX1 g71702(.A (n_5312), .Y (n_7104));
INVX1 g75219(.A (n_5310), .Y (n_5311));
INVX1 g75227(.A (n_7526), .Y (n_5309));
NAND3X1 g75236(.A (n_5306), .B (n_5305), .C (n_7410), .Y (n_5307));
INVX1 g75237(.A (n_5303), .Y (n_5304));
INVX1 g75400(.A (n_6960), .Y (n_6494));
INVX1 g75249(.A (n_5298), .Y (n_5299));
NAND2X1 g75251(.A (n_8363), .B (n_6439), .Y (n_5297));
INVX1 g75253(.A (n_5295), .Y (n_5296));
INVX1 g75267(.A (n_4963), .Y (n_6512));
INVX1 g75269(.A (n_7480), .Y (n_5294));
NOR2X1 g77041(.A (n_16480), .B (n_3955), .Y (n_6372));
NOR2X1 g75287(.A (n_4802), .B (n_3511), .Y (n_6350));
NAND2X1 g75689(.A (n_5204), .B (n_28733), .Y (n_7767));
INVX1 g77994(.A (n_18617), .Y (n_15113));
NOR2X1 g75327(.A (n_5457), .B (n_7598), .Y (n_5290));
INVX1 g75331(.A (n_5289), .Y (n_8604));
NAND2X1 g75334(.A (n_2170), .B (n_2744), .Y (n_5288));
NAND2X1 g69218(.A (n_6188), .B (n_379), .Y (n_10943));
INVX1 g75347(.A (n_5285), .Y (n_9046));
INVX1 g75355(.A (n_12228), .Y (n_5282));
INVX1 g74592(.A (n_5278), .Y (n_8393));
NOR2X1 g75383(.A (n_4428), .B (n_13593), .Y (n_5276));
NOR2X1 g75397(.A (n_4894), .B (n_677), .Y (n_28991));
INVX1 g75408(.A (n_5272), .Y (n_5273));
NAND3X1 g75410(.A (n_5271), .B (n_15473), .C (n_7325), .Y (n_18739));
NOR2X1 g70625(.A (n_4668), .B (n_5186), .Y (n_9353));
NAND2X1 g75429(.A (n_3144), .B (n_15388), .Y (n_5269));
NAND2X1 g75395(.A (n_6313), .B (n_1493), .Y (n_5264));
NAND2X1 g75450(.A (n_3940), .B (n_9416), .Y (n_5263));
AND2X1 g75457(.A (n_2265), .B (n_11323), .Y (n_5262));
INVX1 g75461(.A (n_5260), .Y (n_5261));
INVX1 g75463(.A (n_5258), .Y (n_5259));
INVX1 g75475(.A (n_5257), .Y (n_8889));
INVX1 g75493(.A (n_7238), .Y (n_5255));
INVX1 g75498(.A (n_7005), .Y (n_5253));
INVX1 g75500(.A (n_5251), .Y (n_5252));
NAND2X1 g75506(.A (n_5149), .B (n_3925), .Y (n_6489));
AND2X1 g75509(.A (n_2334), .B (n_4709), .Y (n_5250));
INVX1 g75520(.A (n_6902), .Y (n_5247));
INVX1 g75543(.A (n_5242), .Y (n_5243));
NOR2X1 g71679(.A (n_4606), .B (n_10495), .Y (n_5239));
INVX1 g75034(.A (n_4251), .Y (n_6563));
NAND3X1 g75554(.A (n_2838), .B (n_5236), .C (n_5817), .Y (n_5237));
INVX1 g75581(.A (n_27686), .Y (n_5233));
NAND3X1 g75584(.A (n_530), .B (n_5231), .C (n_11307), .Y (n_5232));
INVX1 g75593(.A (n_5230), .Y (n_8855));
CLKBUFX1 g75603(.A (n_6582), .Y (n_9050));
NAND2X1 g75609(.A (n_3079), .B (n_11576), .Y (n_5229));
OR2X1 g75610(.A (n_3149), .B (n_8945), .Y (n_5228));
NAND2X1 g69198(.A (n_5944), .B (n_7607), .Y (n_7566));
INVX1 g75639(.A (n_5227), .Y (n_6390));
NAND2X1 g75652(.A (n_27309), .B (n_5225), .Y (n_5226));
INVX1 g75661(.A (n_4127), .Y (n_9246));
NAND2X1 g75668(.A (n_3097), .B (n_3086), .Y (n_5224));
INVX1 g75673(.A (n_5222), .Y (n_25664));
INVX1 g75692(.A (n_7121), .Y (n_5221));
NAND2X1 g75699(.A (n_2456), .B (n_5218), .Y (n_5219));
NAND2X1 g75704(.A (n_2613), .B (n_1921), .Y (n_5217));
INVX1 g75705(.A (n_12133), .Y (n_5216));
DFFX1 text_in_r_reg[126] (.CK (clk), .D (n_3213), .Q(text_in_r[126] ), .QN ());
INVX1 g75735(.A (n_5214), .Y (n_8564));
NAND2X1 g75680(.A (n_5212), .B (n_27688), .Y (n_5213));
NOR2X1 g75745(.A (n_5171), .B (n_7496), .Y (n_5211));
NOR2X1 g75746(.A (n_3106), .B (n_12917), .Y (n_5210));
NAND2X1 g75756(.A (n_1261), .B (n_16434), .Y (n_5205));
NAND2X2 g75779(.A (n_5203), .B (n_5204), .Y (n_8569));
INVX2 g75785(.A (n_4803), .Y (n_6952));
INVX1 g75801(.A (n_5202), .Y (n_7006));
NAND2X1 g75808(.A (n_29062), .B (n_5218), .Y (n_5201));
NAND2X1 g75682(.A (n_4988), .B (n_4300), .Y (n_6458));
INVX1 g75814(.A (n_5198), .Y (n_10975));
INVX1 g75817(.A (n_5196), .Y (n_5197));
NAND2X1 g70592(.A (n_4413), .B (n_6185), .Y (n_9557));
OR2X1 g75819(.A (n_2461), .B (n_6005), .Y (n_5194));
OR2X1 g75822(.A (n_3883), .B (n_27124), .Y (n_5193));
NAND2X1 g75829(.A (n_3125), .B (n_15473), .Y (n_5191));
CLKBUFX1 g75834(.A (n_5188), .Y (n_10163));
NAND2X1 g75837(.A (n_2741), .B (n_7658), .Y (n_5187));
NAND2X1 g75841(.A (n_4045), .B (n_5186), .Y (n_8076));
OR2X1 g75863(.A (n_3588), .B (n_13490), .Y (n_5182));
INVX1 g75864(.A (n_4152), .Y (n_5181));
NAND2X1 g75867(.A (n_5179), .B (n_3501), .Y (n_5180));
INVX1 g75870(.A (n_5177), .Y (n_5178));
NOR2X1 g75874(.A (n_5383), .B (n_3849), .Y (n_7984));
NAND2X1 g75881(.A (n_27070), .B (n_3171), .Y (n_5176));
OR2X1 g75887(.A (n_3046), .B (n_4165), .Y (n_5175));
NAND2X1 g75889(.A (n_2357), .B (n_5143), .Y (n_16477));
NAND2X1 g75893(.A (n_4866), .B (n_6346), .Y (n_6515));
AND2X1 g75898(.A (n_6510), .B (n_2401), .Y (n_5174));
NAND2X1 g75382(.A (n_5171), .B (n_8637), .Y (n_5172));
AND2X1 g75902(.A (n_9914), .B (n_4249), .Y (n_5170));
NOR2X1 g75907(.A (n_27069), .B (n_4080), .Y (n_6440));
NAND2X1 g75910(.A (n_5155), .B (n_3257), .Y (n_10830));
NAND2X1 g75912(.A (n_3816), .B (n_1177), .Y (n_8113));
OR2X1 g75915(.A (n_3050), .B (n_3391), .Y (n_5169));
NAND2X1 g75916(.A (n_13837), .B (n_3133), .Y (n_5168));
NOR2X1 g75927(.A (n_5167), .B (n_5316), .Y (n_8120));
INVX1 g75820(.A (n_5165), .Y (n_5166));
NAND2X1 g75931(.A (n_11669), .B (n_3105), .Y (n_5164));
INVX1 g75908(.A (n_5162), .Y (n_5163));
INVX1 g75935(.A (n_5160), .Y (n_5161));
NAND2X1 g75939(.A (n_12268), .B (n_3488), .Y (n_5159));
NOR2X1 g75947(.A (n_3777), .B (n_1552), .Y (n_6435));
NAND2X1 g75948(.A (n_5155), .B (n_5154), .Y (n_5156));
NOR2X1 g75954(.A (n_3132), .B (n_29355), .Y (n_5153));
OAI21X1 g75960(.A0 (n_790), .A1 (n_5151), .B0 (n_3517), .Y (n_5152));
OAI21X1 g75965(.A0 (n_2905), .A1 (n_6462), .B0 (n_3034), .Y (n_5150));
NAND2X1 g73980(.A (n_5149), .B (n_5148), .Y (n_6733));
INVX1 g73976(.A (n_5147), .Y (n_6738));
INVX2 g75672(.A (n_5222), .Y (n_6470));
INVX1 g75370(.A (n_5145), .Y (n_5146));
AND2X1 g75904(.A (n_7194), .B (n_5143), .Y (n_5144));
DFFX1 text_in_r_reg[105] (.CK (clk), .D (n_3390), .Q(text_in_r[105] ), .QN ());
DFFX1 text_in_r_reg[13] (.CK (clk), .D (n_3290), .Q (text_in_r[13]), .QN ());
NAND2X2 g75130(.A (n_4039), .B (n_4568), .Y (n_5140));
NAND2X1 g75901(.A (n_29214), .B (n_5138), .Y (n_15497));
AND2X1 g75899(.A (n_10199), .B (n_3689), .Y (n_5137));
NOR2X1 g71644(.A (n_6946), .B (n_5135), .Y (n_5136));
AND2X1 g74558(.A (n_2627), .B (n_1376), .Y (n_5134));
AND2X1 g77953(.A (n_16434), .B (n_5131), .Y (n_16072));
NAND2X1 g75934(.A (n_11916), .B (n_3104), .Y (n_5130));
INVX1 g74994(.A (n_4256), .Y (n_9098));
XOR2X1 g76189(.A (n_23763), .B (n_9467), .Y (n_5129));
INVX1 g80273(.A (n_819), .Y (n_11998));
AND2X1 g77952(.A (n_13606), .B (n_13679), .Y (n_5128));
XOR2X1 g76233(.A (text_in_r[8] ), .B (w3[8] ), .Y (n_5126));
NOR2X1 g72626(.A (n_5123), .B (n_27746), .Y (n_5124));
XOR2X1 g76262(.A (text_in_r[24] ), .B (n_2004), .Y (n_5122));
NOR2X1 g72509(.A (n_4225), .B (n_27434), .Y (n_5120));
INVX1 g74991(.A (n_5118), .Y (n_5119));
XOR2X1 g76293(.A (n_1103), .B (n_2251), .Y (n_5117));
INVX1 g75342(.A (n_7631), .Y (n_6500));
INVX1 g75338(.A (n_4103), .Y (n_8935));
INVX1 g76359(.A (n_4329), .Y (n_19755));
INVX1 g76361(.A (n_4329), .Y (n_13787));
INVX1 g76365(.A (n_5581), .Y (n_25409));
INVX1 g76369(.A (n_5843), .Y (n_25361));
INVX1 g76374(.A (n_5112), .Y (n_25341));
INVX2 g76377(.A (n_5112), .Y (n_25320));
INVX1 g76402(.A (n_5111), .Y (n_6391));
NAND2X1 g73958(.A (n_4544), .B (n_6328), .Y (n_6742));
NAND2X1 g75335(.A (n_4987), .B (n_3654), .Y (n_5105));
NAND2X1 g74978(.A (n_2311), .B (n_2303), .Y (n_6392));
INVX1 g75640(.A (n_5227), .Y (n_5103));
INVX1 g69084(.A (n_4653), .Y (n_9418));
NOR2X1 g72504(.A (n_5101), .B (n_9783), .Y (n_5102));
INVX1 g69074(.A (n_4655), .Y (n_7591));
NAND2X1 g76718(.A (n_3936), .B (n_5085), .Y (n_5086));
NOR2X1 g76767(.A (n_9410), .B (n_2720), .Y (n_8018));
AND2X1 g76809(.A (n_3301), .B (n_6335), .Y (n_5079));
INVX2 g74534(.A (n_5077), .Y (n_6384));
INVX1 g76860(.A (n_5073), .Y (n_7938));
NAND2X1 g76961(.A (n_4926), .B (n_367), .Y (n_5068));
NOR2X1 g69046(.A (n_4970), .B (n_4865), .Y (n_5066));
AND2X1 g77037(.A (n_3868), .B (n_3264), .Y (n_5064));
OR2X1 g75632(.A (n_3532), .B (n_4113), .Y (n_6376));
INVX1 g75628(.A (n_4049), .Y (n_6475));
INVX1 g77069(.A (n_4392), .Y (n_6735));
NAND2X1 g75322(.A (n_8363), .B (n_1493), .Y (n_5058));
INVX1 g77154(.A (n_5052), .Y (n_5053));
INVX1 g74524(.A (n_4319), .Y (n_7894));
NOR2X1 g72024(.A (n_5047), .B (n_2655), .Y (n_5048));
NAND2X1 g74522(.A (n_4681), .B (n_367), .Y (n_6647));
NOR2X1 g64360(.A (n_3785), .B (u0_r0_rcnt[0] ), .Y (n_5044));
INVX1 g76376(.A (n_5112), .Y (n_25432));
AND2X1 g77361(.A (n_383), .B (n_3530), .Y (n_7981));
NOR2X1 g75809(.A (n_2487), .B (n_29371), .Y (n_8355));
INVX2 g75619(.A (n_6930), .Y (n_8141));
NAND2X1 g74955(.A (n_2850), .B (n_28444), .Y (n_5042));
NAND2X1 g75311(.A (n_3070), .B (n_4113), .Y (n_5037));
INVX1 g73934(.A (n_5040), .Y (n_5034));
DFFX1 text_in_r_reg[120] (.CK (clk), .D (n_3219), .Q(text_in_r[120] ), .QN ());
NAND2X1 g77550(.A (n_17912), .B (n_310), .Y (n_5033));
NOR2X1 g75309(.A (n_3697), .B (n_27904), .Y (n_5032));
NAND2X1 g77617(.A (n_3597), .B (n_8637), .Y (n_5030));
DFFX1 text_in_r_reg[84] (.CK (clk), .D (n_3395), .Q (text_in_r[84]), .QN ());
NAND2X1 g73928(.A (n_4744), .B (n_383), .Y (n_6746));
NAND2X1 g77658(.A (n_27990), .B (n_1336), .Y (n_6364));
AND2X1 g77674(.A (n_2681), .B (n_29102), .Y (n_19750));
DFFX1 text_in_r_reg[74] (.CK (clk), .D (n_3418), .Q (text_in_r[74]), .QN ());
NOR2X1 g77726(.A (n_11835), .B (n_27216), .Y (n_19966));
NOR2X1 g71604(.A (n_27223), .B (n_4861), .Y (n_5024));
INVX1 g77810(.A (n_5020), .Y (n_5021));
AND2X1 g77819(.A (n_6352), .B (n_9388), .Y (n_11418));
INVX1 g77825(.A (n_5018), .Y (n_5019));
AND2X1 g77830(.A (n_5817), .B (n_4357), .Y (n_5017));
NAND2X2 g70458(.A (n_5015), .B (n_3820), .Y (n_6363));
INVX1 g77921(.A (n_6428), .Y (n_5014));
NAND2X1 g77968(.A (n_15473), .B (n_3014), .Y (n_5013));
AND2X1 g75886(.A (n_10859), .B (n_2111), .Y (n_5012));
INVX1 g75702(.A (n_5010), .Y (n_5011));
OR2X1 g75300(.A (n_2873), .B (n_196), .Y (n_5009));
INVX1 g78066(.A (n_5007), .Y (n_5008));
INVX2 g75791(.A (n_5038), .Y (n_6972));
NOR2X1 g72487(.A (n_4769), .B (n_5005), .Y (n_5006));
DFFX1 text_in_r_reg[16] (.CK (clk), .D (n_3220), .Q (text_in_r[16]), .QN ());
DFFX1 text_in_r_reg[40] (.CK (clk), .D (n_3587), .Q (text_in_r[40]), .QN ());
INVX1 g73545(.A (n_5004), .Y (n_8971));
DFFX1 text_in_r_reg[15] (.CK (clk), .D (n_3242), .Q (text_in_r[15]), .QN ());
DFFX1 text_in_r_reg[121] (.CK (clk), .D (n_3341), .Q(text_in_r[121] ), .QN ());
NOR2X1 g70440(.A (n_3820), .B (n_4290), .Y (n_7312));
DFFX1 text_in_r_reg[41] (.CK (clk), .D (n_3126), .Q (text_in_r[41]), .QN ());
DFFX1 text_in_r_reg[36] (.CK (clk), .D (n_3231), .Q (text_in_r[36]), .QN ());
NAND2X1 g74616(.A (n_4659), .B (n_26873), .Y (n_6640));
INVX1 g73898(.A (n_4997), .Y (n_6750));
INVX1 g73890(.A (n_4614), .Y (n_6753));
DFFX1 text_in_r_reg[20] (.CK (clk), .D (n_3409), .Q (text_in_r[20]), .QN ());
DFFX1 u0_r0_rcnt_reg[2] (.CK (clk), .D (n_3545), .Q (u0_r0_rcnt[2]), .QN ());
NAND2X1 g73878(.A (n_4009), .B (n_6303), .Y (n_4993));
DFFX1 text_in_r_reg[32] (.CK (clk), .D (n_3754), .Q (text_in_r[32]), .QN ());
DFFX1 text_in_r_reg[75] (.CK (clk), .D (n_3403), .Q (text_in_r[75]), .QN ());
DFFX1 text_in_r_reg[88] (.CK (clk), .D (n_3521), .Q (text_in_r[88]), .QN ());
AND2X1 g75288(.A (n_4988), .B (n_13834), .Y (n_4989));
NAND2X1 g75608(.A (n_4987), .B (n_2748), .Y (n_6354));
INVX1 g75290(.A (n_4827), .Y (n_8904));
NAND2X1 g74929(.A (n_26385), .B (n_9500), .Y (n_6581));
NAND2X1 g72476(.A (n_4986), .B (n_4882), .Y (n_6971));
DFFX1 text_in_r_reg[33] (.CK (clk), .D (n_3236), .Q (text_in_r[33]), .QN ());
NOR2X1 g70414(.A (n_4767), .B (n_6462), .Y (n_4983));
OR2X1 g75606(.A (n_4980), .B (n_9264), .Y (n_4981));
CLKBUFX1 g74920(.A (n_5373), .Y (n_6584));
NOR2X1 g78170(.A (n_10389), .B (n_177), .Y (n_17760));
INVX2 g75121(.A (n_4979), .Y (n_6420));
INVX1 g74452(.A (n_4978), .Y (n_5463));
INVX1 g75591(.A (n_5786), .Y (n_4977));
NOR2X1 g78113(.A (n_29166), .B (n_29228), .Y (n_4976));
NOR2X1 g75192(.A (n_4974), .B (n_4973), .Y (n_12756));
NOR2X1 g75835(.A (n_3890), .B (n_9500), .Y (n_5188));
INVX1 g74910(.A (n_4970), .Y (n_5375));
INVX1 g74464(.A (n_3571), .Y (n_5460));
NOR2X1 g75600(.A (n_3923), .B (n_27990), .Y (n_4969));
INVX2 g74904(.A (n_4967), .Y (n_6339));
INVX1 g77864(.A (n_4966), .Y (n_6677));
INVX2 g74187(.A (n_3646), .Y (n_7288));
NAND2X1 g74456(.A (n_4965), .B (n_3301), .Y (n_6097));
NOR2X1 g75268(.A (n_3903), .B (n_27990), .Y (n_4963));
NAND2X1 g75594(.A (n_3915), .B (n_596), .Y (n_5230));
NAND2X2 g73861(.A (n_3076), .B (n_4961), .Y (n_4962));
INVX1 g75717(.A (n_4960), .Y (n_7317));
INVX1 g75270(.A (n_5860), .Y (n_7480));
NOR2X1 g70340(.A (n_4132), .B (n_7593), .Y (n_5958));
INVX1 g75262(.A (n_29181), .Y (n_6333));
OR2X1 g74896(.A (n_3710), .B (n_2779), .Y (n_7452));
INVX1 g75823(.A (n_5810), .Y (n_6855));
AND2X1 g77383(.A (n_4582), .B (n_15473), .Y (n_4951));
INVX1 g74448(.A (n_4950), .Y (n_6332));
NOR2X1 g75588(.A (n_9712), .B (n_3234), .Y (n_4945));
NAND2X1 g75254(.A (n_1264), .B (n_7366), .Y (n_5295));
INVX1 g76590(.A (n_4941), .Y (n_15588));
INVX4 g82042(.A (n_124), .Y (n_21552));
INVX1 g76937(.A (n_4939), .Y (n_9704));
NAND2X1 g75250(.A (n_4331), .B (n_5413), .Y (n_5298));
NAND2X1 g75501(.A (n_4760), .B (n_4438), .Y (n_5251));
NAND2X1 g73839(.A (n_3041), .B (n_6462), .Y (n_4938));
INVX1 g74438(.A (n_3323), .Y (n_5469));
INVX1 g74393(.A (n_3887), .Y (n_6344));
NOR2X1 g71526(.A (n_4533), .B (n_4882), .Y (n_5850));
INVX1 g78111(.A (n_4930), .Y (n_18643));
NAND2X1 g74881(.A (n_9959), .B (n_719), .Y (n_4929));
NOR2X1 g74196(.A (n_4928), .B (n_4426), .Y (n_12517));
INVX1 g75547(.A (n_3289), .Y (n_5240));
NAND2X1 g74876(.A (n_29215), .B (n_4611), .Y (n_7415));
NOR2X1 g73823(.A (n_2902), .B (n_6219), .Y (n_4927));
INVX1 g78389(.A (n_4926), .Y (n_10619));
NOR2X1 g73826(.A (n_4925), .B (n_25729), .Y (n_5574));
INVX1 g74870(.A (n_6144), .Y (n_4923));
NAND2X1 g74586(.A (n_29150), .B (n_4568), .Y (n_4922));
NAND2X1 g75238(.A (n_8342), .B (n_4920), .Y (n_5303));
INVX1 g74404(.A (n_4919), .Y (n_7069));
NOR2X1 g73792(.A (n_4581), .B (n_4825), .Y (n_5588));
NOR2X1 g71510(.A (n_3475), .B (n_4916), .Y (n_7639));
NOR2X1 g74410(.A (n_3671), .B (n_3807), .Y (n_28812));
INVX1 g74867(.A (n_4914), .Y (n_4915));
INVX1 g73810(.A (n_4911), .Y (n_4912));
NAND2X1 g75529(.A (n_976), .B (n_1186), .Y (n_4909));
INVX1 g73808(.A (n_8719), .Y (n_5580));
AND2X1 g74588(.A (n_4117), .B (n_2318), .Y (n_4908));
NOR2X1 g71502(.A (n_4500), .B (n_3920), .Y (n_4907));
INVX1 g76378(.A (n_4622), .Y (n_5112));
INVX1 g78352(.A (n_3868), .Y (n_9202));
INVX2 g74396(.A (n_4906), .Y (n_7185));
INVX1 g75430(.A (n_5878), .Y (n_4905));
INVX1 g75728(.A (n_5803), .Y (n_5215));
OR2X1 g75496(.A (n_3175), .B (n_4422), .Y (n_4904));
NAND2X1 g74381(.A (n_4635), .B (n_1946), .Y (n_5475));
INVX1 g75240(.A (n_4902), .Y (n_4903));
OR2X1 g76904(.A (n_3301), .B (n_2239), .Y (n_4901));
INVX1 g74388(.A (n_4899), .Y (n_4900));
OR2X1 g75474(.A (n_1911), .B (n_4898), .Y (n_6913));
NOR2X1 g74386(.A (n_2645), .B (n_27990), .Y (n_4897));
INVX1 g76569(.A (n_4893), .Y (n_5096));
NAND2X1 g74140(.A (n_29355), .B (n_4327), .Y (n_5521));
NOR2X1 g75232(.A (n_2345), .B (n_4861), .Y (n_4891));
AND2X1 g75444(.A (n_2890), .B (n_6007), .Y (n_4887));
AND2X1 g77811(.A (n_2323), .B (n_5799), .Y (n_5020));
INVX1 g71476(.A (n_7798), .Y (n_5855));
INVX1 g73780(.A (n_4886), .Y (n_9774));
INVX1 g73773(.A (n_4883), .Y (n_6266));
NAND2X1 g74370(.A (n_3778), .B (n_4882), .Y (n_6268));
INVX1 g73749(.A (n_5936), .Y (n_6951));
INVX1 g73768(.A (n_4881), .Y (n_6953));
INVX1 g74366(.A (n_27669), .Y (n_6961));
NOR2X1 g71198(.A (n_3772), .B (n_8865), .Y (n_4878));
NOR2X1 g73758(.A (n_3827), .B (n_28575), .Y (n_5956));
CLKBUFX3 g74342(.A (n_4872), .Y (n_7549));
NAND2X1 g73755(.A (n_2706), .B (n_8679), .Y (n_9528));
INVX1 g75758(.A (n_4869), .Y (n_4870));
INVX1 g75223(.A (n_4867), .Y (n_4868));
OR2X1 g73754(.A (n_3723), .B (n_7658), .Y (n_9294));
NOR2X1 g74346(.A (n_4866), .B (n_4865), .Y (n_6368));
NOR2X1 g77328(.A (n_3868), .B (n_11312), .Y (n_4864));
INVX1 g75222(.A (n_4867), .Y (n_9163));
INVX1 g73575(.A (n_4859), .Y (n_4860));
INVX2 g74827(.A (n_4857), .Y (n_6907));
INVX1 g74336(.A (n_3329), .Y (n_5487));
INVX1 g74299(.A (n_3799), .Y (n_7230));
NAND2X1 g73728(.A (n_29358), .B (n_6279), .Y (n_4856));
INVX1 g74822(.A (n_4855), .Y (n_6239));
INVX1 g74816(.A (n_4852), .Y (n_6243));
INVX1 g78292(.A (n_4851), .Y (n_6244));
NAND2X1 g73742(.A (n_4849), .B (n_4848), .Y (n_4850));
NOR2X1 g74810(.A (n_3717), .B (n_4846), .Y (n_4847));
NOR2X1 g70114(.A (n_4612), .B (n_6226), .Y (n_4845));
NOR2X1 g74318(.A (n_3924), .B (n_7419), .Y (n_4844));
INVX1 g74321(.A (n_3806), .Y (n_7479));
INVX1 g73729(.A (n_4841), .Y (n_13655));
INVX2 g75047(.A (n_4839), .Y (n_5349));
AND2X1 g77128(.A (n_4837), .B (n_5151), .Y (n_4838));
INVX1 g75401(.A (n_4836), .Y (n_6960));
NAND2X1 g73587(.A (n_3768), .B (n_218), .Y (n_4835));
NOR2X1 g74800(.A (n_4832), .B (n_3422), .Y (n_5393));
NOR2X1 g74043(.A (n_2598), .B (n_4882), .Y (n_6334));
INVX1 g78194(.A (n_4829), .Y (n_4830));
INVX1 g76561(.A (n_6313), .Y (n_4828));
NOR2X1 g75291(.A (n_3965), .B (n_11272), .Y (n_4827));
NAND2X1 g74798(.A (n_4266), .B (n_5483), .Y (n_6227));
NOR2X1 g72672(.A (n_4825), .B (n_4525), .Y (n_6249));
NOR2X1 g78282(.A (n_3834), .B (n_12105), .Y (n_4824));
NOR2X1 g70094(.A (n_2480), .B (n_9388), .Y (n_5972));
INVX1 g73722(.A (n_7617), .Y (n_4820));
INVX2 g74310(.A (n_4819), .Y (n_7176));
INVX2 g74306(.A (n_3330), .Y (n_5493));
NAND2X1 g74794(.A (n_4339), .B (n_3464), .Y (n_4814));
INVX1 g74792(.A (n_4811), .Y (n_5394));
NOR2X1 g73720(.A (n_4154), .B (n_29244), .Y (n_5605));
OR2X1 g75879(.A (n_3247), .B (n_3138), .Y (n_4807));
NAND2X1 g74786(.A (n_25747), .B (n_3017), .Y (n_5396));
INVX1 g74297(.A (n_3769), .Y (n_7258));
NOR2X1 g74296(.A (n_4804), .B (n_3917), .Y (n_5494));
NAND2X1 g74784(.A (n_2990), .B (n_3920), .Y (n_6212));
INVX2 g73376(.A (n_3705), .Y (n_5975));
NOR2X1 g75786(.A (n_5005), .B (n_3235), .Y (n_4803));
INVX1 g77733(.A (n_4802), .Y (n_6210));
INVX1 g74780(.A (n_4801), .Y (n_8837));
NAND2X1 g74774(.A (n_2881), .B (n_4825), .Y (n_5399));
INVX1 g77881(.A (n_4800), .Y (n_6767));
INVX1 g75570(.A (n_5101), .Y (n_6209));
NOR2X1 g74776(.A (n_2397), .B (n_6303), .Y (n_4796));
AND2X1 g76872(.A (n_9500), .B (n_1735), .Y (n_6603));
OR2X1 g74770(.A (n_1177), .B (n_3920), .Y (n_10676));
INVX1 g75482(.A (n_4792), .Y (n_5749));
AND2X1 g73702(.A (n_3622), .B (n_28733), .Y (n_5609));
NOR2X1 g75151(.A (n_2647), .B (n_11307), .Y (n_4789));
INVX2 g75564(.A (n_4788), .Y (n_7367));
NOR2X1 g71315(.A (n_4786), .B (n_6226), .Y (n_4787));
INVX1 g74276(.A (n_4784), .Y (n_5499));
NOR2X1 g74768(.A (n_3830), .B (n_5660), .Y (n_4783));
NAND2X1 g74764(.A (n_2369), .B (n_10031), .Y (n_4782));
INVX1 g76861(.A (n_26385), .Y (n_5073));
INVX1 g76540(.A (n_3173), .Y (n_6194));
OR2X1 g75126(.A (n_3119), .B (n_9057), .Y (n_7417));
INVX1 g74760(.A (n_3199), .Y (n_5406));
INVX2 g73684(.A (n_5616), .Y (n_5613));
INVX1 g76425(.A (n_4776), .Y (n_4777));
INVX1 g76849(.A (n_5368), .Y (n_5074));
AND2X1 g73590(.A (n_3473), .B (n_4916), .Y (n_11413));
NOR2X1 g73676(.A (n_2839), .B (n_2191), .Y (n_5937));
INVX1 g76841(.A (n_4773), .Y (n_7730));
INVX1 g76845(.A (n_4772), .Y (n_13974));
NOR2X1 g73674(.A (n_3651), .B (n_4961), .Y (n_5614));
NAND2X1 g75071(.A (n_2775), .B (n_27124), .Y (n_5340));
INVX2 g74252(.A (n_4771), .Y (n_5503));
INVX1 g77244(.A (n_4770), .Y (n_6656));
INVX1 g74740(.A (n_4769), .Y (n_6183));
INVX1 g75722(.A (n_5774), .Y (n_6206));
INVX1 g75023(.A (n_3248), .Y (n_5352));
NOR2X1 g74244(.A (n_2113), .B (n_27365), .Y (n_5505));
NAND2X1 g74230(.A (n_4760), .B (n_1353), .Y (n_4761));
NAND2X1 g74241(.A (n_4520), .B (n_28744), .Y (n_6171));
NOR2X1 g73017(.A (n_11626), .B (n_4582), .Y (n_4758));
NOR2X1 g70010(.A (n_27366), .B (n_26491), .Y (n_5976));
INVX1 g78230(.A (n_4753), .Y (n_4754));
INVX1 g74997(.A (n_6265), .Y (n_4752));
NOR2X1 g72338(.A (n_4565), .B (n_379), .Y (n_5772));
NOR2X1 g73638(.A (n_4586), .B (n_25746), .Y (n_5625));
INVX1 g73632(.A (n_5930), .Y (n_6887));
OR2X1 g73627(.A (n_3071), .B (n_3599), .Y (n_7770));
INVX2 g78218(.A (n_4748), .Y (n_6096));
INVX1 g77681(.A (n_4744), .Y (n_4745));
OR2X1 g74221(.A (n_2771), .B (n_9416), .Y (n_4743));
INVX2 g74921(.A (n_5802), .Y (n_5373));
NOR2X1 g75742(.A (n_2333), .B (n_5151), .Y (n_7152));
INVX1 g76423(.A (n_3494), .Y (n_5108));
INVX1 g75555(.A (n_4739), .Y (n_7041));
INVX1 g76480(.A (n_2885), .Y (n_4738));
INVX1 g76815(.A (n_4736), .Y (n_6730));
NOR2X1 g71311(.A (n_4552), .B (n_5922), .Y (n_4731));
INVX1 g74209(.A (n_4730), .Y (n_6991));
INVX2 g75521(.A (n_4728), .Y (n_6902));
NOR2X1 g75805(.A (n_3513), .B (n_11253), .Y (n_4726));
OR2X1 g75804(.A (n_2878), .B (n_4721), .Y (n_4722));
NAND2X1 g73016(.A (n_1584), .B (n_3814), .Y (n_7624));
NOR2X1 g69938(.A (n_4604), .B (n_2655), .Y (n_4718));
NOR2X1 g73580(.A (n_4158), .B (n_27904), .Y (n_5638));
INVX2 g75802(.A (n_5123), .Y (n_5202));
INVX2 g73562(.A (n_4715), .Y (n_5642));
NAND2X1 g74787(.A (n_4169), .B (n_14055), .Y (n_4714));
AND2X1 g74829(.A (n_4207), .B (n_4391), .Y (n_4713));
INVX1 g76796(.A (n_1988), .Y (n_4712));
NAND2X1 g74198(.A (n_4349), .B (n_4709), .Y (n_6131));
INVX2 g73612(.A (n_4741), .Y (n_7114));
NOR2X1 g69786(.A (n_5381), .B (n_4705), .Y (n_4708));
NOR2X1 g74714(.A (n_6462), .B (n_27438), .Y (n_5054));
NOR2X1 g69898(.A (n_4705), .B (n_6185), .Y (n_4706));
INVX2 g73548(.A (n_4703), .Y (n_4704));
NOR2X1 g71232(.A (n_3499), .B (n_5922), .Y (n_6104));
NOR2X1 g74180(.A (n_4699), .B (n_8452), .Y (n_4700));
NOR2X1 g73527(.A (n_4200), .B (n_9118), .Y (n_4697));
NAND2X1 g74830(.A (n_4012), .B (n_28037), .Y (n_4694));
NOR2X1 g74696(.A (n_4176), .B (n_29225), .Y (n_4691));
OR2X1 g74942(.A (n_4595), .B (n_4689), .Y (n_7003));
INVX2 g73510(.A (n_4692), .Y (n_5646));
INVX1 g74166(.A (n_4688), .Y (n_5628));
OR2X1 g69852(.A (n_2768), .B (n_13083), .Y (n_13700));
NOR2X1 g71325(.A (n_3417), .B (n_8263), .Y (n_4687));
OR2X1 g74158(.A (n_11924), .B (n_4416), .Y (n_5761));
INVX1 g74597(.A (n_3699), .Y (n_6111));
INVX1 g73489(.A (n_4456), .Y (n_4685));
NAND2X1 g72914(.A (n_27904), .B (n_3865), .Y (n_5715));
XOR2X1 g76303(.A (text_in_r[16] ), .B (n_250), .Y (n_4684));
INVX2 g74150(.A (n_3336), .Y (n_14386));
NOR2X1 g75158(.A (n_2647), .B (n_3307), .Y (n_7008));
INVX1 g76444(.A (n_5612), .Y (n_4682));
INVX1 g74563(.A (n_5966), .Y (n_6963));
INVX1 g76751(.A (n_4681), .Y (n_7675));
INVX1 g74698(.A (n_4678), .Y (n_4679));
INVX1 g74553(.A (n_3193), .Y (n_5437));
AND2X1 g74542(.A (n_2775), .B (n_28375), .Y (n_4675));
INVX1 g74535(.A (n_4672), .Y (n_5077));
INVX1 g77219(.A (n_4671), .Y (n_6856));
NAND2X1 g74520(.A (n_2373), .B (n_3307), .Y (n_5443));
INVX2 g74130(.A (n_4669), .Y (n_8024));
NOR2X1 g73462(.A (n_4228), .B (n_7485), .Y (n_5657));
INVX2 g74257(.A (n_4668), .Y (n_7210));
NOR2X1 g72794(.A (n_3829), .B (n_8865), .Y (n_5723));
NOR2X1 g75959(.A (n_2008), .B (n_28487), .Y (n_4666));
NAND2X1 g75228(.A (n_4108), .B (n_4522), .Y (n_7526));
INVX1 g72880(.A (n_3771), .Y (n_7717));
INVX1 g74371(.A (n_5725), .Y (n_4665));
INVX1 g76403(.A (n_25926), .Y (n_5111));
INVX1 g71180(.A (n_7603), .Y (n_6093));
AND2X1 g74112(.A (n_1264), .B (n_9118), .Y (n_4664));
NOR2X1 g73440(.A (n_4663), .B (n_10389), .Y (n_6086));
CLKBUFX3 g74040(.A (n_4658), .Y (n_6415));
INVX1 g74688(.A (n_5915), .Y (n_5411));
NOR2X1 g75550(.A (n_2694), .B (n_9500), .Y (n_6169));
AND2X1 g69057(.A (n_3273), .B (n_4598), .Y (n_6074));
NOR2X1 g69075(.A (n_3589), .B (n_383), .Y (n_4655));
NAND2X1 g69085(.A (n_3852), .B (n_28742), .Y (n_4653));
NOR2X1 g73416(.A (n_3796), .B (n_383), .Y (n_5667));
OR2X1 g69174(.A (n_3682), .B (n_5817), .Y (n_17274));
INVX1 g74225(.A (n_4650), .Y (n_6149));
NOR2X1 g69241(.A (n_3269), .B (n_7182), .Y (n_4647));
NAND2X1 g74203(.A (n_4326), .B (n_15986), .Y (n_4646));
NOR2X1 g69284(.A (n_4643), .B (n_4825), .Y (n_4644));
INVX2 g73406(.A (n_4642), .Y (n_5670));
AND2X1 g69364(.A (n_14734), .B (n_2779), .Y (n_9314));
OR2X1 g69369(.A (n_2768), .B (n_3301), .Y (n_7733));
OR2X1 g69388(.A (n_4639), .B (n_7410), .Y (n_4640));
INVX1 g75488(.A (n_4196), .Y (n_6151));
NAND2X1 g69456(.A (n_3032), .B (n_9527), .Y (n_7672));
OR2X1 g69473(.A (n_4638), .B (n_9527), .Y (n_5751));
INVX1 g75148(.A (n_4636), .Y (n_7058));
NAND2X1 g74118(.A (n_4635), .B (n_3820), .Y (n_5525));
NAND3X1 g69502(.A (n_6279), .B (n_4326), .C (n_2191), .Y (n_14337));
NOR2X1 g69551(.A (n_3306), .B (n_3920), .Y (n_4634));
BUFX3 g76389(.A (n_25926), .Y (n_25283));
BUFX3 g76388(.A (n_25926), .Y (n_25274));
NOR2X1 g69573(.A (n_4590), .B (n_8679), .Y (n_5862));
NOR2X1 g69583(.A (n_2768), .B (n_7777), .Y (n_4632));
NOR2X1 g73875(.A (n_2750), .B (n_5990), .Y (n_5567));
AND2X1 g74058(.A (n_3135), .B (n_3920), .Y (n_7576));
INVX1 g75856(.A (n_27367), .Y (n_6374));
INVX1 g73382(.A (n_3574), .Y (n_6010));
NAND2X1 g74111(.A (n_2704), .B (n_4627), .Y (n_5528));
OR2X1 g69733(.A (n_4638), .B (n_8679), .Y (n_4626));
INVX2 g75811(.A (n_5988), .Y (n_8499));
OR2X1 g69739(.A (n_2665), .B (n_7325), .Y (n_11625));
NAND2X1 g69742(.A (n_2479), .B (n_13606), .Y (n_4625));
NAND2X2 g69793(.A (n_3250), .B (n_27904), .Y (n_14085));
INVX1 g76383(.A (n_4622), .Y (n_5969));
INVX2 g73977(.A (n_3232), .Y (n_5147));
NAND3X1 g73372(.A (n_2891), .B (n_28358), .C (n_1591), .Y (n_5674));
NOR2X1 g75544(.A (n_3084), .B (n_4490), .Y (n_5242));
INVX1 g73965(.A (n_3206), .Y (n_5552));
NAND2X2 g74238(.A (n_4635), .B (n_3251), .Y (n_7071));
NAND2X1 g72066(.A (n_3469), .B (n_6007), .Y (n_11449));
NAND2X1 g69921(.A (n_3869), .B (n_271), .Y (n_4619));
INVX2 g75494(.A (n_4618), .Y (n_7238));
NOR2X1 g73891(.A (n_3209), .B (n_6462), .Y (n_4614));
INVX1 g76368(.A (n_4622), .Y (n_5581));
NOR2X1 g70103(.A (n_4612), .B (n_4611), .Y (n_4613));
INVX2 g73609(.A (n_4741), .Y (n_29410));
INVX1 g73485(.A (n_4606), .Y (n_4607));
NOR2X1 g70214(.A (n_4604), .B (n_7331), .Y (n_4605));
NAND2X1 g73802(.A (n_2541), .B (n_12169), .Y (n_10836));
NAND2X1 g75849(.A (n_2399), .B (n_3017), .Y (n_4601));
INVX1 g73805(.A (n_4600), .Y (n_7578));
INVX1 g73776(.A (n_4602), .Y (n_4599));
NOR2X1 g73361(.A (n_4514), .B (n_4598), .Y (n_5675));
NAND2X1 g70324(.A (n_3353), .B (n_28410), .Y (n_4597));
NOR2X1 g75094(.A (n_4595), .B (n_6462), .Y (n_4596));
NAND2X1 g70359(.A (n_13738), .B (n_9388), .Y (n_12655));
AND2X1 g74088(.A (n_4373), .B (n_8997), .Y (n_4594));
NOR2X1 g73740(.A (n_3579), .B (n_4598), .Y (n_5602));
NAND4X1 g70379(.A (n_6868), .B (n_490), .C (n_2251), .D (n_3014), .Y(n_4593));
NOR2X1 g74072(.A (n_6609), .B (n_3052), .Y (n_7085));
INVX1 g73724(.A (n_4833), .Y (n_4592));
INVX1 g73694(.A (n_8379), .Y (n_5610));
OR2X1 g70504(.A (n_4590), .B (n_11354), .Y (n_13703));
NOR2X1 g70630(.A (n_27366), .B (n_4586), .Y (n_4588));
NAND2X1 g73344(.A (n_4450), .B (n_3695), .Y (n_5931));
INVX1 g73336(.A (n_4585), .Y (n_6842));
INVX1 g74092(.A (n_3518), .Y (n_5532));
OR2X1 g73434(.A (n_4581), .B (n_12559), .Y (n_6237));
NOR2X1 g73327(.A (n_1581), .B (n_7496), .Y (n_5681));
NAND2X1 g70765(.A (n_383), .B (n_3610), .Y (n_7634));
NOR2X1 g70827(.A (n_3385), .B (n_4627), .Y (n_5689));
INVX1 g70838(.A (n_3366), .Y (n_7744));
INVX1 g73551(.A (n_4703), .Y (n_7120));
AND2X1 g75533(.A (n_2704), .B (n_1147), .Y (n_4575));
NAND2X1 g73312(.A (n_4105), .B (n_2744), .Y (n_9927));
INVX1 g76705(.A (n_4659), .Y (n_4573));
NAND2X1 g74675(.A (n_3159), .B (n_4113), .Y (n_4572));
NAND2X1 g70953(.A (n_3437), .B (n_11312), .Y (n_5805));
NOR2X1 g73499(.A (n_2515), .B (n_11323), .Y (n_4570));
NOR2X1 g70987(.A (n_3241), .B (n_4568), .Y (n_4569));
INVX1 g75531(.A (n_11067), .Y (n_5882));
OR2X1 g71037(.A (n_4565), .B (n_7325), .Y (n_7625));
NOR2X1 g73660(.A (n_4302), .B (n_7496), .Y (n_5618));
INVX1 g73475(.A (n_5716), .Y (n_5654));
NAND2X1 g71054(.A (n_3911), .B (n_26873), .Y (n_14324));
NAND2X1 g71057(.A (n_3726), .B (n_5422), .Y (n_4563));
INVX1 g75747(.A (n_4561), .Y (n_4562));
NOR2X1 g71185(.A (n_3692), .B (n_3920), .Y (n_6084));
OR2X1 g71203(.A (n_7568), .B (n_11307), .Y (n_4558));
NOR2X1 g71206(.A (n_6005), .B (n_4401), .Y (n_4557));
NAND2X1 g74049(.A (n_2625), .B (n_383), .Y (n_4555));
INVX1 g73389(.A (n_4554), .Y (n_7116));
INVX1 g75641(.A (n_4553), .Y (n_5227));
OR2X1 g71265(.A (n_4552), .B (n_14866), .Y (n_18116));
INVX1 g73355(.A (n_4550), .Y (n_6958));
INVX1 g75522(.A (n_4728), .Y (n_4549));
NAND2X1 g71314(.A (n_4547), .B (n_9257), .Y (n_4548));
INVX1 g73337(.A (n_4585), .Y (n_4546));
INVX1 g73333(.A (n_3449), .Y (n_7813));
NAND3X1 g71327(.A (n_29062), .B (n_4544), .C (n_5530), .Y (n_18310));
INVX1 g73321(.A (n_4543), .Y (n_5684));
NAND2X1 g71420(.A (n_19110), .B (n_7568), .Y (n_4540));
INVX1 g73814(.A (n_4539), .Y (n_5578));
INVX1 g75516(.A (n_27223), .Y (n_6261));
INVX1 g75827(.A (n_26890), .Y (n_6956));
NOR2X1 g69566(.A (n_26602), .B (n_4825), .Y (n_4537));
NAND2X1 g71492(.A (n_3287), .B (n_9474), .Y (n_4536));
NAND2X1 g71505(.A (n_3922), .B (n_7496), .Y (n_5853));
NOR2X1 g71516(.A (n_4533), .B (n_9388), .Y (n_4534));
INVX1 g76397(.A (n_25926), .Y (n_6067));
INVX1 g76373(.A (n_4622), .Y (n_5843));
OR2X1 g71647(.A (n_3237), .B (n_8679), .Y (n_9529));
INVX1 g75115(.A (n_5135), .Y (n_5816));
NAND2X2 g71703(.A (n_12559), .B (n_26993), .Y (n_5312));
NOR2X1 g71769(.A (n_4525), .B (n_8865), .Y (n_4526));
OR2X1 g71845(.A (n_11626), .B (n_7325), .Y (n_7710));
NOR2X1 g71861(.A (n_3338), .B (n_4504), .Y (n_7388));
NAND2X1 g71877(.A (n_4721), .B (n_3345), .Y (n_5767));
NAND2X1 g71895(.A (n_3455), .B (n_6008), .Y (n_16621));
NOR2X1 g74636(.A (n_3844), .B (n_4522), .Y (n_4523));
NAND2X1 g71923(.A (n_3040), .B (n_10599), .Y (n_11510));
NAND2X2 g75112(.A (n_4520), .B (n_27599), .Y (n_7062));
NAND2X1 g71961(.A (n_6021), .B (n_27640), .Y (n_5866));
NOR2X1 g75528(.A (n_4245), .B (n_28423), .Y (n_4519));
INVX2 g71996(.A (n_3396), .Y (n_7726));
NOR2X1 g73394(.A (n_3030), .B (n_3234), .Y (n_5671));
INVX1 g71890(.A (n_3398), .Y (n_11593));
NAND2X1 g72149(.A (n_6133), .B (n_3842), .Y (n_6082));
NOR2X1 g74650(.A (n_3698), .B (n_4848), .Y (n_4518));
NOR2X1 g72171(.A (n_4513), .B (n_5643), .Y (n_4517));
INVX1 g72172(.A (n_6134), .Y (n_15465));
NAND2X1 g75806(.A (n_7023), .B (n_28869), .Y (n_4516));
NAND2X1 g73127(.A (n_28744), .B (n_3342), .Y (n_5700));
NOR2X1 g72205(.A (n_3825), .B (n_9442), .Y (n_6128));
NOR2X1 g72303(.A (n_4513), .B (n_12559), .Y (n_5775));
OR2X1 g72314(.A (n_3893), .B (n_26491), .Y (n_4512));
NOR2X1 g69496(.A (n_3372), .B (n_3307), .Y (n_4511));
INVX1 g72346(.A (n_3722), .Y (n_4509));
NOR2X1 g74648(.A (n_3148), .B (n_28757), .Y (n_5419));
NOR3X1 g72383(.A (n_13318), .B (n_3319), .C (n_8910), .Y (n_4507));
OR2X1 g72427(.A (n_13681), .B (n_12169), .Y (n_5759));
NOR2X1 g72459(.A (n_4504), .B (n_6005), .Y (n_4505));
NOR2X1 g72465(.A (n_3444), .B (n_379), .Y (n_7665));
NOR2X1 g71871(.A (n_4234), .B (n_9410), .Y (n_4503));
NOR2X1 g75553(.A (n_4501), .B (n_7410), .Y (n_4502));
OR2X1 g72580(.A (n_4500), .B (n_12169), .Y (n_9190));
NAND2X1 g73830(.A (n_28487), .B (n_4627), .Y (n_4499));
AND2X1 g75780(.A (n_2521), .B (n_8945), .Y (n_4496));
NAND2X1 g72777(.A (n_3350), .B (n_4709), .Y (n_13118));
INVX1 g78078(.A (n_4492), .Y (n_4493));
NOR2X1 g75471(.A (n_2586), .B (n_4490), .Y (n_4491));
NAND2X1 g72616(.A (n_4804), .B (n_3294), .Y (n_5742));
NAND2X1 g74174(.A (n_5167), .B (n_8816), .Y (n_7164));
NOR2X1 g74260(.A (n_3729), .B (n_636), .Y (n_4489));
NOR2X1 g75090(.A (n_5368), .B (n_6946), .Y (n_5337));
OR2X1 g73049(.A (n_3316), .B (n_2779), .Y (n_13539));
NOR2X1 g74703(.A (n_4353), .B (n_9084), .Y (n_4488));
OR2X1 g73119(.A (n_3891), .B (n_165), .Y (n_4487));
NOR2X1 g71837(.A (n_3060), .B (n_2768), .Y (n_5819));
NAND2X2 g73400(.A (n_3836), .B (n_1584), .Y (n_5884));
NOR2X1 g75862(.A (n_3687), .B (n_6008), .Y (n_4484));
OR2X1 g72602(.A (n_4547), .B (n_5854), .Y (n_4483));
INVX1 g74750(.A (n_5800), .Y (n_5408));
XOR2X1 g76105(.A (n_1019), .B (n_23399), .Y (n_4482));
INVX1 g74413(.A (n_4481), .Y (n_7299));
INVX1 g73307(.A (n_8295), .Y (n_4480));
OR2X1 g73313(.A (n_4405), .B (n_28445), .Y (n_12505));
NAND2X1 g75448(.A (n_3874), .B (n_27990), .Y (n_6280));
INVX1 g73345(.A (n_4478), .Y (n_14831));
OR2X1 g73350(.A (n_3755), .B (n_7266), .Y (n_5677));
OR2X1 g73351(.A (n_3049), .B (n_1946), .Y (n_8487));
INVX1 g73363(.A (n_9220), .Y (n_4477));
INVX1 g73379(.A (n_4475), .Y (n_4476));
NOR2X1 g72596(.A (n_3715), .B (n_5643), .Y (n_5686));
NOR2X1 g73423(.A (n_1083), .B (n_196), .Y (n_4470));
INVX1 g73424(.A (n_9800), .Y (n_4468));
NOR2X1 g73443(.A (n_2183), .B (n_2260), .Y (n_5663));
INVX1 g73444(.A (n_4559), .Y (n_4466));
INVX1 g73449(.A (n_4465), .Y (n_5662));
INVX1 g73452(.A (n_4463), .Y (n_4464));
INVX1 g73454(.A (n_4462), .Y (n_8209));
INVX1 g73463(.A (n_4798), .Y (n_4461));
INVX2 g73469(.A (n_3644), .Y (n_6102));
NOR2X1 g73473(.A (n_2017), .B (n_8997), .Y (n_4460));
INVX1 g73477(.A (n_4458), .Y (n_4459));
INVX2 g73481(.A (n_4457), .Y (n_7319));
INVX1 g73484(.A (n_4606), .Y (n_13646));
INVX1 g73488(.A (n_4456), .Y (n_7290));
NOR2X1 g73493(.A (n_4210), .B (n_8452), .Y (n_5650));
INVX1 g73503(.A (n_9236), .Y (n_5648));
INVX1 g75736(.A (n_3013), .Y (n_5214));
NOR2X1 g73515(.A (n_2862), .B (n_8974), .Y (n_4455));
NAND2X1 g73529(.A (n_4168), .B (n_6012), .Y (n_4454));
NAND2X1 g75445(.A (n_2707), .B (n_2145), .Y (n_4453));
INVX1 g73535(.A (n_3633), .Y (n_5644));
NOR2X1 g73542(.A (n_4227), .B (n_7485), .Y (n_4451));
NAND2X1 g73543(.A (n_4450), .B (n_11731), .Y (n_13799));
INVX1 g73554(.A (n_9293), .Y (n_4447));
INVX1 g73602(.A (n_3678), .Y (n_7376));
OR2X1 g73604(.A (n_4404), .B (n_28408), .Y (n_7170));
INVX1 g73618(.A (n_4441), .Y (n_6164));
NAND2X1 g73621(.A (n_4450), .B (n_7563), .Y (n_7203));
NAND2X1 g75818(.A (n_2311), .B (n_4414), .Y (n_5196));
NAND2X1 g73629(.A (n_4438), .B (n_11322), .Y (n_12291));
NOR2X1 g74644(.A (n_2302), .B (n_9500), .Y (n_5420));
INVX1 g73641(.A (n_4757), .Y (n_4437));
NOR2X1 g73649(.A (n_2350), .B (n_29286), .Y (n_4436));
INVX1 g73655(.A (n_4435), .Y (n_6898));
INVX1 g73661(.A (n_4433), .Y (n_4434));
OR2X1 g73663(.A (n_1921), .B (n_7777), .Y (n_7686));
INVX2 g73667(.A (n_4767), .Y (n_5617));
OR2X1 g73700(.A (n_3694), .B (n_6007), .Y (n_7137));
INVX1 g78052(.A (n_4428), .Y (n_4429));
NOR2X1 g73737(.A (n_4426), .B (n_4113), .Y (n_5951));
INVX1 g73745(.A (n_4424), .Y (n_5599));
OR2X1 g73759(.A (n_1503), .B (n_11215), .Y (n_12722));
NAND2X1 g73761(.A (n_4422), .B (n_4825), .Y (n_4423));
INVX1 g73763(.A (n_3829), .Y (n_5595));
AOI21X1 g63903(.A0 (n_6301), .A1 (dcnt[1] ), .B0 (n_2390), .Y(n_4421));
INVX1 g73781(.A (n_4886), .Y (n_4420));
INVX1 g73795(.A (n_4419), .Y (n_5585));
INVX1 g73799(.A (n_4418), .Y (n_7420));
NAND2X1 g73821(.A (n_3425), .B (n_27904), .Y (n_4417));
NOR2X1 g75936(.A (n_3711), .B (n_2376), .Y (n_5160));
NOR2X1 g73834(.A (n_4416), .B (n_27990), .Y (n_5571));
NAND2X1 g73867(.A (n_4414), .B (n_28375), .Y (n_6989));
INVX1 g73869(.A (n_4413), .Y (n_4984));
INVX1 g73930(.A (n_4408), .Y (n_5559));
INVX1 g73935(.A (n_4407), .Y (n_5040));
NAND2X1 g73970(.A (n_4405), .B (n_4404), .Y (n_4406));
INVX1 g73971(.A (n_4403), .Y (n_6920));
NOR2X1 g71782(.A (n_4401), .B (n_14624), .Y (n_4402));
NOR2X1 g73983(.A (n_3701), .B (n_6012), .Y (n_4400));
NOR2X1 g74005(.A (n_3562), .B (n_6055), .Y (n_5350));
NAND2X1 g74009(.A (n_2605), .B (n_28744), .Y (n_5543));
INVX1 g74010(.A (n_4396), .Y (n_4397));
NOR2X1 g74015(.A (n_2609), .B (n_3834), .Y (n_5541));
INVX1 g74017(.A (n_7032), .Y (n_4394));
NAND2X1 g74023(.A (n_3165), .B (n_4490), .Y (n_4393));
INVX2 g74032(.A (n_3505), .Y (n_5590));
NOR2X1 g77070(.A (n_2837), .B (n_4391), .Y (n_4392));
NAND2X1 g74045(.A (n_2819), .B (n_27124), .Y (n_4390));
OR2X1 g70747(.A (n_4867), .B (n_3736), .Y (n_7708));
NOR2X1 g74658(.A (n_28749), .B (n_4388), .Y (n_4389));
INVX1 g74065(.A (n_5771), .Y (n_7440));
NAND2X1 g74071(.A (n_2396), .B (n_8816), .Y (n_4386));
INVX1 g74076(.A (n_4385), .Y (n_6223));
NAND2X1 g74087(.A (n_3134), .B (n_677), .Y (n_4384));
NOR2X1 g74095(.A (n_4382), .B (n_4055), .Y (n_5932));
NAND2X1 g74109(.A (n_4318), .B (n_8742), .Y (n_4381));
NOR2X1 g74115(.A (n_4280), .B (n_6185), .Y (n_4380));
INVX1 g74122(.A (n_4379), .Y (n_7370));
INVX1 g74124(.A (n_4377), .Y (n_4378));
NAND2X1 g74132(.A (n_4375), .B (n_5143), .Y (n_4376));
OR2X1 g75065(.A (n_4373), .B (n_3288), .Y (n_4374));
AND2X1 g74159(.A (n_2393), .B (n_28037), .Y (n_4372));
INVX1 g74169(.A (n_6099), .Y (n_4371));
NAND2X1 g74201(.A (n_3230), .B (n_5643), .Y (n_7615));
INVX1 g74204(.A (n_4369), .Y (n_4370));
NAND2X1 g74207(.A (n_4544), .B (n_29149), .Y (n_4368));
NAND2X1 g74216(.A (n_4422), .B (n_4367), .Y (n_11642));
INVX1 g74620(.A (n_4366), .Y (n_5427));
NAND2X1 g69308(.A (n_3312), .B (n_4364), .Y (n_4365));
NAND2X1 g75502(.A (n_2456), .B (n_2323), .Y (n_4363));
INVX1 g74270(.A (n_5741), .Y (n_4359));
AND2X1 g74272(.A (n_2716), .B (n_4357), .Y (n_4358));
NAND2X1 g74284(.A (n_3500), .B (n_10100), .Y (n_4356));
NAND2X1 g74308(.A (n_4353), .B (n_12917), .Y (n_4354));
NAND2X1 g74325(.A (n_4349), .B (n_5005), .Y (n_4350));
INVX1 g74331(.A (n_5770), .Y (n_7477));
AND2X1 g74347(.A (n_2605), .B (n_276), .Y (n_29427));
INVX1 g74351(.A (n_4695), .Y (n_5481));
INVX1 g74680(.A (n_4345), .Y (n_4346));
INVX1 g74357(.A (n_4344), .Y (n_6256));
INVX1 g74375(.A (n_4343), .Y (n_6270));
INVX2 g74399(.A (n_3871), .Y (n_7824));
NOR2X1 g74401(.A (n_4022), .B (n_9118), .Y (n_9718));
INVX1 g74419(.A (n_4342), .Y (n_6891));
NAND2X1 g74433(.A (n_2367), .B (n_6133), .Y (n_6315));
NAND2X1 g74450(.A (n_4339), .B (n_4326), .Y (n_4340));
NOR2X1 g74470(.A (n_4334), .B (n_8945), .Y (n_4335));
AND2X1 g75069(.A (n_4331), .B (n_26873), .Y (n_4332));
AND2X1 g74474(.A (n_2938), .B (n_26493), .Y (n_4330));
INVX1 g76358(.A (n_4329), .Y (n_5114));
NAND2X1 g74478(.A (n_6696), .B (n_13466), .Y (n_4328));
NAND2X1 g74480(.A (n_4327), .B (n_4326), .Y (n_5454));
INVX1 g74481(.A (n_3975), .Y (n_4325));
NOR2X1 g69280(.A (n_3812), .B (n_28757), .Y (n_6050));
NAND2X1 g74506(.A (n_5778), .B (n_1142), .Y (n_4323));
NOR2X1 g74507(.A (n_4598), .B (n_3218), .Y (n_7262));
INVX1 g74512(.A (n_4320), .Y (n_4321));
NOR2X1 g74525(.A (n_4318), .B (n_11322), .Y (n_4319));
NOR2X1 g74541(.A (n_3000), .B (n_5990), .Y (n_4316));
NAND2X2 g75068(.A (n_2565), .B (n_28757), .Y (n_5343));
INVX1 g75417(.A (n_4315), .Y (n_7487));
INVX1 g74566(.A (n_6011), .Y (n_4314));
NAND2X1 g74572(.A (n_1298), .B (n_15894), .Y (n_4310));
INVX1 g74574(.A (n_5787), .Y (n_4309));
INVX1 g74581(.A (n_4308), .Y (n_12292));
INVX2 g74589(.A (n_4307), .Y (n_7553));
INVX1 g74593(.A (n_5768), .Y (n_5278));
INVX1 g74609(.A (n_3306), .Y (n_7128));
NAND2X1 g74627(.A (n_2460), .B (n_3327), .Y (n_5576));
NOR2X1 g75706(.A (n_1075), .B (n_379), .Y (n_12133));
NAND2X1 g74629(.A (n_1581), .B (n_4302), .Y (n_4304));
INVX1 g74663(.A (n_4301), .Y (n_5804));
NOR2X1 g74678(.A (n_2821), .B (n_4300), .Y (n_6939));
NOR2X1 g75924(.A (n_15812), .B (n_4299), .Y (n_12720));
INVX1 g74704(.A (n_4297), .Y (n_4298));
NAND2X1 g74716(.A (n_2125), .B (n_9500), .Y (n_4295));
INVX1 g74746(.A (n_5820), .Y (n_4293));
INVX1 g74752(.A (n_4291), .Y (n_4292));
INVX1 g74757(.A (n_4290), .Y (n_7123));
INVX1 g74781(.A (n_4801), .Y (n_4289));
INVX1 g74795(.A (n_4285), .Y (n_4286));
INVX1 g77520(.A (n_3841), .Y (n_6293));
NAND2X1 g75411(.A (n_6587), .B (n_16466), .Y (n_4283));
INVX1 g78016(.A (n_4282), .Y (n_5403));
NAND2X1 g74835(.A (n_4280), .B (n_9003), .Y (n_4281));
INVX1 g74836(.A (n_5823), .Y (n_4279));
NAND2X1 g74839(.A (n_4146), .B (n_5422), .Y (n_7145));
NOR2X1 g74847(.A (n_3005), .B (n_28742), .Y (n_10181));
INVX1 g74865(.A (n_5910), .Y (n_6295));
INVX1 g74605(.A (n_5692), .Y (n_4277));
INVX1 g74877(.A (n_12822), .Y (n_4276));
AND2X1 g75504(.A (n_4375), .B (n_2541), .Y (n_6934));
AND2X1 g74897(.A (n_2834), .B (n_8560), .Y (n_4275));
INVX1 g74899(.A (n_4273), .Y (n_4274));
INVX1 g74006(.A (n_4271), .Y (n_4272));
OR2X1 g74913(.A (n_3364), .B (n_4426), .Y (n_4270));
INVX1 g75056(.A (n_4269), .Y (n_5347));
INVX1 g74926(.A (n_4268), .Y (n_7403));
AND2X1 g74945(.A (n_4266), .B (n_1942), .Y (n_4267));
OR2X1 g74947(.A (n_2573), .B (n_3307), .Y (n_4265));
AND2X1 g75701(.A (n_3107), .B (n_7410), .Y (n_4264));
OR2X1 g74962(.A (n_3221), .B (n_4261), .Y (n_4262));
INVX1 g74965(.A (n_4260), .Y (n_5360));
INVX1 g74969(.A (n_12578), .Y (n_4259));
INVX1 g74975(.A (n_4258), .Y (n_5099));
NAND2X1 g74979(.A (n_5271), .B (n_9527), .Y (n_4257));
INVX1 g74602(.A (n_5826), .Y (n_5430));
NAND2X1 g74995(.A (n_2926), .B (n_5983), .Y (n_4256));
INVX1 g75011(.A (n_4255), .Y (n_7358));
NOR2X1 g75015(.A (n_3921), .B (n_4113), .Y (n_4253));
NAND2X1 g70655(.A (n_26486), .B (n_3691), .Y (n_5928));
NOR2X1 g75035(.A (n_3087), .B (n_4934), .Y (n_4251));
INVX1 g75037(.A (n_5942), .Y (n_7159));
NAND2X2 g70662(.A (n_3679), .B (n_28408), .Y (n_9547));
NAND2X1 g75066(.A (n_5149), .B (n_4249), .Y (n_4250));
INVX1 g75072(.A (n_6232), .Y (n_4248));
INVX1 g75084(.A (n_4247), .Y (n_7567));
INVX1 g75087(.A (n_5912), .Y (n_7678));
NAND2X1 g75053(.A (n_4245), .B (n_28381), .Y (n_4246));
INVX1 g75107(.A (n_4243), .Y (n_5757));
NOR2X1 g69234(.A (n_4590), .B (n_490), .Y (n_4242));
NOR2X1 g75141(.A (n_3388), .B (n_28037), .Y (n_4241));
NAND2X1 g75143(.A (n_12222), .B (n_1065), .Y (n_4238));
OR2X1 g75146(.A (n_5138), .B (n_6226), .Y (n_7216));
INVX1 g75165(.A (n_3652), .Y (n_6308));
NOR2X1 g75179(.A (n_3240), .B (n_5983), .Y (n_5318));
NOR2X1 g70644(.A (n_4234), .B (n_27365), .Y (n_4235));
AND2X1 g75186(.A (n_4233), .B (n_3038), .Y (n_7193));
NOR2X1 g75462(.A (n_2519), .B (n_6021), .Y (n_5260));
INVX1 g75197(.A (n_3858), .Y (n_6217));
INVX1 g75209(.A (n_5484), .Y (n_6229));
INVX1 g75217(.A (n_3817), .Y (n_6245));
NOR2X1 g75220(.A (n_2754), .B (n_6419), .Y (n_5310));
NAND2X1 g75226(.A (n_2380), .B (n_8816), .Y (n_4232));
NAND2X1 g75239(.A (n_4228), .B (n_4227), .Y (n_4229));
INVX1 g75246(.A (n_4225), .Y (n_5301));
NAND2X1 g75248(.A (n_2577), .B (n_8910), .Y (n_4224));
INVX1 g75255(.A (n_4222), .Y (n_4223));
INVX1 g75264(.A (n_5705), .Y (n_4221));
INVX1 g73410(.A (n_4471), .Y (n_6060));
NAND2X1 g75272(.A (n_3130), .B (n_4113), .Y (n_4220));
INVX2 g75277(.A (n_5047), .Y (n_6342));
NAND2X1 g75279(.A (n_976), .B (n_4217), .Y (n_4219));
INVX1 g75298(.A (n_5435), .Y (n_7659));
INVX1 g75349(.A (n_4216), .Y (n_7535));
NAND2X1 g75371(.A (n_2890), .B (n_6133), .Y (n_5145));
INVX1 g75378(.A (n_4213), .Y (n_4214));
AND2X1 g75389(.A (n_4104), .B (n_29225), .Y (n_4212));
INVX1 g75390(.A (n_3913), .Y (n_7292));
NAND2X1 g75396(.A (n_4210), .B (n_2515), .Y (n_4211));
OR2X1 g75398(.A (n_4208), .B (n_9712), .Y (n_4209));
NOR2X1 g75407(.A (n_6005), .B (n_6836), .Y (n_5331));
NAND2X1 g75409(.A (n_4207), .B (n_7438), .Y (n_5272));
NAND2X1 g75412(.A (n_4126), .B (n_6007), .Y (n_4206));
NAND2X1 g75419(.A (n_5149), .B (n_1972), .Y (n_4205));
INVX1 g75420(.A (n_4204), .Y (n_7350));
INVX1 g75423(.A (n_5971), .Y (n_6304));
NOR2X1 g75427(.A (n_3776), .B (n_5005), .Y (n_7486));
INVX1 g73998(.A (n_4203), .Y (n_7183));
INVX1 g75455(.A (n_4202), .Y (n_7106));
NAND2X1 g75459(.A (n_3796), .B (n_4200), .Y (n_4201));
INVX1 g75464(.A (n_4199), .Y (n_5258));
NAND2X1 g75497(.A (n_4194), .B (n_790), .Y (n_4195));
NAND2X1 g75499(.A (n_2089), .B (n_3307), .Y (n_7005));
INVX1 g75393(.A (n_4190), .Y (n_4191));
OR2X1 g73995(.A (n_4188), .B (n_4299), .Y (n_4189));
DFFX1 u0_r0_rcnt_reg[1] (.CK (clk), .D (n_3972), .Q (u0_r0_rcnt[1]), .QN ());
INVX1 g77025(.A (n_3257), .Y (n_4187));
INVX1 g75574(.A (n_4184), .Y (n_4185));
INVX1 g75589(.A (n_5974), .Y (n_4182));
INVX1 g75611(.A (n_5833), .Y (n_4181));
NOR2X1 g70610(.A (n_3672), .B (n_4568), .Y (n_4180));
INVX1 g75633(.A (n_4178), .Y (n_4179));
NAND2X1 g75635(.A (n_4176), .B (n_29256), .Y (n_4177));
AND2X1 g75646(.A (n_2641), .B (n_4173), .Y (n_4174));
OR2X1 g75648(.A (n_2352), .B (n_4261), .Y (n_7113));
NAND2X1 g75696(.A (n_2021), .B (n_2140), .Y (n_4172));
NOR2X1 g75703(.A (n_2537), .B (n_4627), .Y (n_5010));
NAND2X1 g75709(.A (n_6442), .B (n_27904), .Y (n_4171));
NOR2X1 g75733(.A (n_4169), .B (n_367), .Y (n_4170));
NAND2X1 g75757(.A (n_4168), .B (n_3160), .Y (n_14231));
INVX1 g75767(.A (n_4167), .Y (n_5721));
INVX1 g75771(.A (n_4166), .Y (n_6068));
INVX1 g76648(.A (n_4165), .Y (n_5091));
NAND2X1 g73988(.A (n_5143), .B (n_3920), .Y (n_5548));
INVX2 g75793(.A (n_3918), .Y (n_5038));
INVX1 g74577(.A (n_4164), .Y (n_5208));
NAND2X1 g75807(.A (n_25744), .B (n_10495), .Y (n_4162));
NOR2X1 g75815(.A (n_4159), .B (n_4158), .Y (n_5198));
NAND2X1 g75821(.A (n_2641), .B (n_3820), .Y (n_5165));
CLKBUFX1 g75379(.A (n_4213), .Y (n_7583));
INVX1 g75832(.A (n_3080), .Y (n_6155));
OR2X1 g75838(.A (n_3052), .B (n_3736), .Y (n_4157));
NAND2X1 g75854(.A (n_4154), .B (n_2350), .Y (n_4155));
NOR2X1 g75865(.A (n_4825), .B (n_29130), .Y (n_4152));
NAND2X1 g75869(.A (n_1609), .B (n_1075), .Y (n_6822));
AND2X1 g75880(.A (n_29149), .B (n_15997), .Y (n_4151));
INVX2 g73985(.A (n_27199), .Y (n_7247));
NOR2X1 g75679(.A (n_4149), .B (n_12559), .Y (n_4150));
AND2X1 g72942(.A (n_14725), .B (n_4547), .Y (n_4148));
NAND2X1 g75903(.A (n_2444), .B (n_1983), .Y (n_6829));
NAND2X1 g75909(.A (n_2709), .B (n_2331), .Y (n_5162));
NAND2X1 g75919(.A (n_5179), .B (n_8097), .Y (n_11112));
NOR2X1 g72521(.A (n_3861), .B (n_5799), .Y (n_5744));
NAND2X1 g75951(.A (n_5778), .B (n_4146), .Y (n_4147));
INVX1 g75479(.A (n_4145), .Y (n_5747));
INVX2 g75674(.A (n_3256), .Y (n_5222));
NAND2X1 g75905(.A (n_12222), .B (n_4144), .Y (n_11100));
INVX1 g77964(.A (n_4142), .Y (n_4143));
NAND2X1 g75369(.A (n_5985), .B (n_12019), .Y (n_4141));
INVX1 g75359(.A (n_3214), .Y (n_5280));
OR2X1 g69149(.A (n_4639), .B (n_12760), .Y (n_6066));
NAND2X1 g75667(.A (n_2306), .B (n_27202), .Y (n_4140));
INVX1 g74538(.A (n_6018), .Y (n_4138));
INVX1 g75362(.A (n_4137), .Y (n_7039));
NOR2X1 g74562(.A (n_3461), .B (n_4113), .Y (n_4136));
OR2X1 g71646(.A (n_3174), .B (n_28037), .Y (n_4135));
INVX1 g75008(.A (n_4134), .Y (n_5355));
NOR2X1 g70544(.A (n_4132), .B (n_4925), .Y (n_4133));
INVX1 g75676(.A (n_5841), .Y (n_4130));
INVX1 g75451(.A (n_5694), .Y (n_4129));
NAND2X1 g75004(.A (n_6198), .B (n_6252), .Y (n_4128));
NOR2X1 g75662(.A (n_4126), .B (n_6007), .Y (n_4127));
INVX1 g75257(.A (n_7685), .Y (n_4124));
NOR2X1 g75356(.A (n_3987), .B (n_7453), .Y (n_12228));
INVX2 g75657(.A (n_4123), .Y (n_6791));
INVX1 g74556(.A (n_5867), .Y (n_4122));
INVX1 g75650(.A (n_3260), .Y (n_7321));
NAND2X1 g75348(.A (n_4117), .B (n_6092), .Y (n_5285));
NAND2X1 g75476(.A (n_4373), .B (n_5990), .Y (n_5257));
INVX1 g75345(.A (n_28859), .Y (n_7503));
NAND2X1 g74992(.A (n_4115), .B (n_29269), .Y (n_5118));
INVX1 g77962(.A (n_4114), .Y (n_5323));
NAND2X1 g78067(.A (n_4113), .B (n_7586), .Y (n_5007));
NOR2X1 g74052(.A (n_3594), .B (n_26493), .Y (n_4112));
NOR2X1 g73962(.A (n_5983), .B (n_4014), .Y (n_5554));
XOR2X1 g76295(.A (n_243), .B (n_2760), .Y (n_4111));
INVX1 g74989(.A (n_4109), .Y (n_4110));
NAND2X1 g75343(.A (n_4108), .B (n_1627), .Y (n_7631));
INVX2 g75694(.A (n_4107), .Y (n_7121));
AND2X1 g74987(.A (n_4106), .B (n_9467), .Y (n_7100));
NAND2X1 g74984(.A (n_4105), .B (n_3802), .Y (n_7296));
NAND2X1 g74986(.A (n_4104), .B (n_2487), .Y (n_5357));
NOR2X1 g75339(.A (n_3144), .B (n_2810), .Y (n_4103));
NOR2X1 g74550(.A (n_3153), .B (n_5422), .Y (n_5439));
INVX1 g75332(.A (n_3180), .Y (n_5289));
NAND2X1 g73954(.A (n_3673), .B (n_6021), .Y (n_4102));
NAND2X1 g76460(.A (n_3824), .B (n_8997), .Y (n_4099));
AND2X1 g75920(.A (n_7101), .B (n_2950), .Y (n_4098));
INVX1 g74546(.A (n_4094), .Y (n_6995));
INVX1 g77009(.A (n_8116), .Y (n_6446));
INVX2 g76633(.A (n_5502), .Y (n_5093));
INVX2 g74972(.A (n_3162), .Y (n_7357));
INVX2 g76669(.A (n_6327), .Y (n_4084));
NOR2X1 g76672(.A (n_4082), .B (n_7496), .Y (n_4083));
INVX1 g76716(.A (n_4076), .Y (n_6285));
INVX1 g76738(.A (n_4072), .Y (n_4073));
INVX1 g74526(.A (n_5764), .Y (n_4071));
NOR2X1 g75871(.A (n_3522), .B (n_3161), .Y (n_5177));
INVX1 g76760(.A (n_4070), .Y (n_6706));
AND2X1 g76880(.A (n_6419), .B (n_1925), .Y (n_6539));
INVX1 g73947(.A (n_26192), .Y (n_5555));
NAND2X1 g76925(.A (n_9500), .B (n_2085), .Y (n_4060));
INVX1 g76971(.A (n_5171), .Y (n_6452));
NOR2X1 g73944(.A (n_4055), .B (n_28733), .Y (n_5072));
INVX1 g62026(.A (n_6286), .Y (n_7805));
AND2X1 g77047(.A (n_9691), .B (n_2999), .Y (n_6522));
INVX1 g77063(.A (n_3331), .Y (n_5061));
AND2X1 g75911(.A (n_6871), .B (n_2089), .Y (n_4051));
NOR2X1 g75629(.A (n_2752), .B (n_5005), .Y (n_4049));
AND2X1 g77924(.A (n_15166), .B (n_4357), .Y (n_4048));
NOR2X1 g75853(.A (n_3575), .B (n_677), .Y (n_4046));
INVX1 g77113(.A (n_4045), .Y (n_7701));
AND2X1 g77116(.A (n_27202), .B (n_3359), .Y (n_6495));
INVX1 g77120(.A (n_4043), .Y (n_12249));
OR2X1 g75312(.A (n_2569), .B (n_4721), .Y (n_6825));
AND2X1 g77143(.A (n_4042), .B (n_5924), .Y (n_6479));
CLKBUFX1 g77195(.A (n_4039), .Y (n_6749));
CLKBUFX1 g77005(.A (n_4038), .Y (n_6636));
INVX1 g74960(.A (n_3122), .Y (n_5363));
INVX1 g77309(.A (n_5457), .Y (n_4037));
NAND2X2 g74282(.A (n_4144), .B (n_4721), .Y (n_4036));
INVX1 g77922(.A (n_4034), .Y (n_6428));
NOR2X1 g77371(.A (n_12827), .B (n_5151), .Y (n_10768));
INVX1 g77381(.A (n_4027), .Y (n_4028));
INVX1 g77384(.A (n_4955), .Y (n_4026));
INVX1 g74943(.A (n_4025), .Y (n_12731));
AND2X1 g77410(.A (n_13318), .B (n_28172), .Y (n_19152));
NOR2X1 g74954(.A (n_4022), .B (n_4113), .Y (n_5367));
INVX1 g77155(.A (n_4021), .Y (n_5052));
INVX2 g75620(.A (n_5593), .Y (n_6930));
INVX1 g77580(.A (n_4018), .Y (n_4019));
NOR2X1 g75551(.A (n_2279), .B (n_5413), .Y (n_6968));
INVX1 g75304(.A (n_4017), .Y (n_5025));
NAND2X1 g74511(.A (n_2393), .B (n_7607), .Y (n_6105));
NOR2X1 g74949(.A (n_4014), .B (n_15388), .Y (n_8118));
NAND2X1 g74614(.A (n_4012), .B (n_4721), .Y (n_6114));
INVX1 g77802(.A (n_4009), .Y (n_6426));
INVX1 g75754(.A (n_3582), .Y (n_5206));
NAND2X1 g77826(.A (n_7728), .B (n_28271), .Y (n_5018));
INVX1 g73922(.A (n_4007), .Y (n_5560));
INVX1 g77833(.A (n_4006), .Y (n_8534));
AND2X1 g75154(.A (n_962), .B (n_5422), .Y (n_5326));
INVX1 g77925(.A (n_4003), .Y (n_4004));
NAND2X1 g77945(.A (n_7586), .B (n_9118), .Y (n_4002));
INVX1 g74682(.A (n_4000), .Y (n_4001));
INVX1 g75281(.A (n_6040), .Y (n_3997));
INVX2 g75604(.A (n_3993), .Y (n_6582));
INVX1 g74502(.A (n_3992), .Y (n_5450));
OR2X1 g74500(.A (n_2320), .B (n_6043), .Y (n_5452));
NAND2X1 g78077(.A (n_9500), .B (n_1569), .Y (n_5946));
INVX1 g73908(.A (n_3991), .Y (n_5564));
NAND2X1 g75443(.A (n_8342), .B (n_4144), .Y (n_3990));
NOR2X1 g78172(.A (n_3888), .B (n_4357), .Y (n_3989));
NOR2X1 g73546(.A (n_5643), .B (n_3987), .Y (n_5004));
INVX1 g74898(.A (n_4273), .Y (n_7406));
INVX1 g75294(.A (n_3039), .Y (n_7517));
INVX1 g74494(.A (n_3981), .Y (n_6974));
NAND2X1 g75913(.A (n_11669), .B (n_4249), .Y (n_10988));
INVX2 g73899(.A (n_3980), .Y (n_4997));
NAND2X1 g75763(.A (n_3702), .B (n_6462), .Y (n_3979));
INVX1 g73894(.A (n_5832), .Y (n_4994));
AND2X1 g64704(.A (n_3972), .B (u0_r0_rcnt[0] ), .Y (n_3973));
NAND2X1 g74288(.A (n_2938), .B (n_4848), .Y (n_5495));
NOR2X1 g72028(.A (n_2843), .B (n_4590), .Y (n_7759));
INVX1 g77887(.A (n_6847), .Y (n_3967));
NAND2X1 g72026(.A (n_3463), .B (n_29269), .Y (n_12734));
NOR2X1 g74477(.A (n_2636), .B (n_6977), .Y (n_5455));
INVX1 g77585(.A (n_5410), .Y (n_6250));
NOR2X1 g75076(.A (n_3666), .B (n_4568), .Y (n_7131));
INVX1 g71582(.A (n_3018), .Y (n_7732));
INVX1 g75538(.A (n_3269), .Y (n_6838));
NAND2X1 g74925(.A (n_3965), .B (n_9942), .Y (n_3966));
NAND2X1 g74475(.A (n_3963), .B (n_16434), .Y (n_3964));
INVX1 g76954(.A (n_5204), .Y (n_6546));
NOR2X1 g71290(.A (n_13681), .B (n_13083), .Y (n_3959));
INVX1 g74472(.A (n_5719), .Y (n_3954));
INVX1 g80008(.A (n_790), .Y (n_4750));
NAND2X1 g73308(.A (n_2608), .B (n_1206), .Y (n_8295));
DFFX1 text_in_r_reg[125] (.CK (clk), .D (n_2047), .Q(text_in_r[125] ), .QN ());
MX2X1 g75989(.A (text_in_r[96] ), .B (text_in[96]), .S0 (n_672), .Y(n_3948));
NAND2X2 g74077(.A (n_2146), .B (n_1627), .Y (n_4385));
NAND2X1 g73555(.A (n_3945), .B (n_9467), .Y (n_9293));
MX2X1 g76038(.A (text_in_r[66] ), .B (text_in[66]), .S0 (n_672), .Y(n_3942));
NOR2X1 g77506(.A (n_9089), .B (n_8997), .Y (n_3940));
INVX1 g80655(.A (n_7543), .Y (n_3936));
NAND2X2 g74905(.A (n_2093), .B (n_28464), .Y (n_4967));
DFFX1 text_in_r_reg[2] (.CK (clk), .D (n_2217), .Q (text_in_r[2] ),.QN ());
NAND2X1 g74453(.A (n_3373), .B (n_4364), .Y (n_4978));
MX2X1 g76007(.A (text_in_r[47] ), .B (text_in[47]), .S0 (n_600), .Y(n_3933));
INVX1 g80778(.A (n_12469), .Y (n_3932));
INVX1 g73863(.A (n_3931), .Y (n_5828));
MX2X1 g76002(.A (text_in_r[54] ), .B (text_in[54]), .S0 (n_600), .Y(n_3930));
NAND2X2 g75122(.A (n_3427), .B (n_29166), .Y (n_4979));
NAND2X2 g75271(.A (n_2026), .B (n_2079), .Y (n_5860));
INVX1 g76688(.A (n_13037), .Y (n_4079));
DFFX1 text_in_r_reg[44] (.CK (clk), .D (n_1578), .Q (text_in_r[44]), .QN ());
NOR2X1 g74900(.A (n_4364), .B (n_2695), .Y (n_4273));
INVX1 g73557(.A (n_3656), .Y (n_6247));
NAND2X1 g73425(.A (n_3643), .B (n_352), .Y (n_9800));
NAND2X1 g65006(.A (n_1501), .B (n_1448), .Y (n_3929));
OR2X1 g75194(.A (n_1779), .B (n_7182), .Y (n_3927));
MX2X1 g76081(.A (text_in_r[103] ), .B (text_in[103]), .S0 (ld), .Y(n_3926));
INVX1 g77375(.A (n_3924), .Y (n_3925));
INVX1 g77386(.A (n_3923), .Y (n_4955));
INVX1 g73853(.A (n_3922), .Y (n_4957));
INVX1 g77006(.A (n_3921), .Y (n_4038));
OR2X1 g75258(.A (n_3816), .B (n_3920), .Y (n_7685));
NAND2X2 g75794(.A (n_1737), .B (n_28476), .Y (n_3918));
OR2X1 g75590(.A (n_2627), .B (n_1701), .Y (n_5974));
DFFX1 text_in_r_reg[72] (.CK (clk), .D (n_1813), .Q (text_in_r[72]), .QN ());
INVX1 g77156(.A (n_3917), .Y (n_4021));
MX2X1 g76051(.A (text_in_r[11] ), .B (text_in[11]), .S0 (n_600), .Y(n_3916));
INVX2 g75613(.A (n_4705), .Y (n_5833));
NAND2X1 g75592(.A (n_3585), .B (n_330), .Y (n_5786));
INVX2 g73552(.A (n_2989), .Y (n_4703));
NOR2X1 g75391(.A (n_2365), .B (n_6043), .Y (n_3913));
INVX1 g73436(.A (n_3911), .Y (n_4943));
DFFX1 text_in_r_reg[101] (.CK (clk), .D (n_1541), .Q(text_in_r[101] ), .QN ());
NAND2X1 g76592(.A (n_19445), .B (n_7777), .Y (n_4941));
MX2X1 g76006(.A (text_in_r[3] ), .B (text_in[3]), .S0 (n_672), .Y(n_3909));
MX2X1 g76074(.A (text_in_r[28] ), .B (text_in[28]), .S0 (n_672), .Y(n_3907));
INVX2 g73338(.A (n_2945), .Y (n_4585));
NOR2X1 g75252(.A (n_3704), .B (n_2937), .Y (n_5839));
INVX1 g76938(.A (n_3903), .Y (n_4939));
INVX2 g77283(.A (n_3760), .Y (n_16934));
NOR2X1 g74878(.A (n_3900), .B (n_3482), .Y (n_12822));
XOR2X1 g76190(.A (text_in_r[71] ), .B (n_22781), .Y (n_3896));
NAND2X1 g75718(.A (n_2719), .B (n_27990), .Y (n_4960));
NAND2X2 g74428(.A (n_1637), .B (n_28358), .Y (n_6031));
NOR2X1 g75243(.A (n_2835), .B (n_4113), .Y (n_5857));
MX2X1 g76087(.A (text_in_r[24] ), .B (text_in[24]), .S0 (n_600), .Y(n_3895));
NAND2X1 g75402(.A (n_2713), .B (n_827), .Y (n_4836));
NAND2X1 g74414(.A (n_2829), .B (n_3038), .Y (n_4481));
AND2X1 g75242(.A (n_3301), .B (n_2324), .Y (n_4902));
INVX1 g78390(.A (n_2960), .Y (n_4926));
INVX1 g74420(.A (n_3893), .Y (n_4342));
INVX1 g76363(.A (ld_r), .Y (n_4329));
DFFX1 text_in_r_reg[106] (.CK (clk), .D (n_1969), .Q(text_in_r[106] ), .QN ());
INVX1 g74872(.A (n_3891), .Y (n_6023));
OR2X1 g74871(.A (n_4501), .B (n_3920), .Y (n_6144));
NAND2X1 g74066(.A (n_3535), .B (n_3840), .Y (n_5771));
CLKBUFX3 g76670(.A (n_3890), .Y (n_6327));
NAND2X1 g73806(.A (n_3322), .B (n_27904), .Y (n_4600));
NOR2X1 g73811(.A (n_2259), .B (n_2674), .Y (n_4911));
INVX2 g75523(.A (n_26547), .Y (n_4728));
NOR2X1 g74394(.A (n_1938), .B (n_379), .Y (n_3887));
DFFX1 text_in_r_reg[4] (.CK (clk), .D (n_1798), .Q (text_in_r[4] ),.QN ());
AND2X1 g74868(.A (n_3536), .B (n_3318), .Y (n_4914));
DFFX1 text_in_r_reg[43] (.CK (clk), .D (n_1816), .Q (text_in_r[43]), .QN ());
NAND2X1 g77827(.A (n_3108), .B (n_28373), .Y (n_3883));
NAND2X1 g74405(.A (n_3448), .B (n_28779), .Y (n_4919));
NAND2X1 g74866(.A (n_3833), .B (n_1627), .Y (n_5910));
DFFX1 text_in_r_reg[112] (.CK (clk), .D (n_2121), .Q(text_in_r[112] ), .QN ());
INVX1 g76680(.A (n_3874), .Y (n_4080));
NAND2X2 g74400(.A (n_2286), .B (n_28757), .Y (n_3871));
MX2X1 g75967(.A (text_in_r[111] ), .B (text_in[111]), .S0 (n_672),.Y (n_3870));
INVX1 g75556(.A (n_3869), .Y (n_4739));
INVX1 g76578(.A (n_3166), .Y (n_10859));
NOR2X1 g78191(.A (n_8865), .B (n_2968), .Y (n_3867));
INVX1 g73796(.A (n_3865), .Y (n_4419));
NAND2X2 g74397(.A (n_3573), .B (n_28351), .Y (n_4906));
NAND2X2 g75495(.A (n_3285), .B (n_1272), .Y (n_4618));
INVX2 g75039(.A (n_3270), .Y (n_5942));
INVX2 g73769(.A (n_2927), .Y (n_4881));
INVX2 g73787(.A (n_3859), .Y (n_6034));
INVX1 g75472(.A (n_3861), .Y (n_3862));
NAND2X1 g75198(.A (n_2818), .B (n_677), .Y (n_3858));
INVX1 g75465(.A (n_3852), .Y (n_4199));
MX2X1 g76044(.A (text_in_r[67] ), .B (text_in[67]), .S0 (n_600), .Y(n_3851));
NAND2X1 g74376(.A (n_3420), .B (n_4611), .Y (n_4343));
INVX1 g77350(.A (n_3849), .Y (n_4884));
DFFX1 text_in_r_reg[93] (.CK (clk), .D (n_1525), .Q (text_in_r[93]), .QN ());
NOR2X1 g73778(.A (n_2864), .B (n_4882), .Y (n_4602));
MX2X1 g75979(.A (text_in_r[90] ), .B (text_in[90]), .S0 (n_672), .Y(n_3845));
INVX1 g75424(.A (n_3276), .Y (n_5971));
INVX1 g77803(.A (n_3844), .Y (n_4009));
INVX1 g77346(.A (n_3102), .Y (n_5600));
NAND2X1 g74372(.A (n_3813), .B (n_383), .Y (n_5725));
INVX1 g73774(.A (n_3842), .Y (n_4883));
INVX1 g76907(.A (n_3471), .Y (n_4875));
INVX2 g73563(.A (n_2884), .Y (n_4715));
NOR2X1 g77521(.A (n_2153), .B (n_3840), .Y (n_3841));
INVX1 g78032(.A (n_3836), .Y (n_3837));
NAND2X1 g75421(.A (n_2724), .B (n_3820), .Y (n_4204));
NOR2X1 g76488(.A (n_3834), .B (n_2368), .Y (n_3835));
NAND2X2 g75716(.A (n_3833), .B (n_3560), .Y (n_28616));
INVX2 g76708(.A (n_3830), .Y (n_3831));
NAND2X1 g77122(.A (n_27370), .B (n_26491), .Y (n_4043));
INVX1 g74360(.A (n_4552), .Y (n_10716));
DFFX1 text_in_r_reg[73] (.CK (clk), .D (n_1653), .Q (text_in_r[73]), .QN ());
NAND2X2 g74358(.A (n_2885), .B (n_4925), .Y (n_4344));
INVX2 g78306(.A (n_3827), .Y (n_8363));
INVX1 g73750(.A (n_3825), .Y (n_5936));
INVX2 g74352(.A (n_4643), .Y (n_4695));
INVX1 g77618(.A (n_3987), .Y (n_3823));
DFFX1 text_in_r_reg[50] (.CK (clk), .D (n_2244), .Q (text_in_r[50]), .QN ());
NAND2X2 g75108(.A (n_3002), .B (n_26887), .Y (n_4243));
NOR2X1 g75363(.A (n_2640), .B (n_3820), .Y (n_4137));
NAND2X2 g74828(.A (n_2344), .B (n_2708), .Y (n_4857));
NAND2X1 g73746(.A (n_3465), .B (n_3807), .Y (n_4424));
NOR2X1 g75218(.A (n_2461), .B (n_4721), .Y (n_3817));
OR2X1 g75366(.A (n_3816), .B (n_7410), .Y (n_9221));
INVX1 g73450(.A (n_3814), .Y (n_4465));
NAND2X1 g74594(.A (n_3813), .B (n_2646), .Y (n_5768));
INVX1 g74332(.A (n_3812), .Y (n_5770));
AND2X1 g78294(.A (n_15894), .B (n_21055), .Y (n_9326));
XOR2X1 g76157(.A (text_in_r[85] ), .B (n_805), .Y (n_3811));
NAND2X1 g77772(.A (n_1569), .B (n_11835), .Y (n_3809));
NAND2X2 g74817(.A (n_26483), .B (n_28478), .Y (n_4852));
NAND2X1 g75350(.A (n_3615), .B (n_3807), .Y (n_4216));
NAND2X1 g74322(.A (n_2958), .B (n_5660), .Y (n_3806));
NAND2X1 g75210(.A (n_3746), .B (n_2383), .Y (n_5484));
AND2X1 g78287(.A (n_27688), .B (n_21174), .Y (n_16007));
MX2X1 g76078(.A (text_in_r[123] ), .B (text_in[123]), .S0 (n_619),.Y (n_3804));
INVX1 g76901(.A (n_2612), .Y (n_4842));
NAND2X1 g75759(.A (n_3802), .B (n_4861), .Y (n_4869));
MX2X1 g76040(.A (text_in_r[70] ), .B (text_in[70]), .S0 (n_672), .Y(n_3800));
NOR2X1 g74300(.A (n_2925), .B (n_5983), .Y (n_3799));
NAND2X1 g75123(.A (n_1688), .B (n_8093), .Y (n_3797));
NOR2X1 g73726(.A (n_2707), .B (n_1584), .Y (n_4833));
DFFX1 text_in_r_reg[100] (.CK (clk), .D (n_1987), .Q(text_in_r[100] ), .QN ());
INVX1 g77304(.A (n_15812), .Y (n_5620));
INVX2 g74312(.A (n_3787), .Y (n_4819));
INVX1 g74313(.A (n_3787), .Y (n_25629));
INVX1 g65957(.A (n_3972), .Y (n_3785));
OR2X1 g77295(.A (n_379), .B (n_2959), .Y (n_3783));
INVX1 g77296(.A (n_3777), .Y (n_13837));
INVX1 g77103(.A (n_3776), .Y (n_4988));
OR2X1 g78276(.A (n_1336), .B (n_29225), .Y (n_29371));
NOR2X1 g74796(.A (n_6694), .B (n_3303), .Y (n_4285));
OR2X1 g76882(.A (n_8090), .B (n_29163), .Y (n_3774));
NAND2X1 g75247(.A (n_27437), .B (n_4568), .Y (n_4225));
INVX1 g75576(.A (n_3772), .Y (n_4184));
NOR2X1 g72881(.A (n_2267), .B (n_3807), .Y (n_3771));
INVX1 g81946(.A (n_2022), .Y (n_13247));
MX2X1 g75984(.A (text_in_r[53] ), .B (text_in[53]), .S0 (ld), .Y(n_3770));
NOR2X1 g74298(.A (n_2366), .B (n_6133), .Y (n_3769));
INVX1 g77734(.A (n_3768), .Y (n_4802));
OR2X1 g77281(.A (n_8945), .B (n_2081), .Y (n_3765));
INVX1 g74717(.A (n_4234), .Y (n_3764));
INVX1 g77134(.A (n_2934), .Y (n_5509));
NAND2X1 g72370(.A (n_14757), .B (n_3600), .Y (n_3758));
DFFX1 text_in_r_reg[114] (.CK (clk), .D (n_1546), .Q(text_in_r[114] ), .QN ());
NOR2X1 g75174(.A (n_1644), .B (n_6997), .Y (n_5788));
NAND2X2 g77011(.A (n_27894), .B (n_3756), .Y (n_8116));
INVX1 g78249(.A (n_3755), .Y (n_6142));
MX2X1 g76013(.A (text_in_r[32] ), .B (text_in[32]), .S0 (n_619), .Y(n_3754));
NAND2X1 g75159(.A (n_4194), .B (n_6352), .Y (n_3753));
DFFX1 text_in_r_reg[25] (.CK (clk), .D (n_2105), .Q (text_in_r[25]), .QN ());
NAND2X2 g75565(.A (n_1902), .B (n_3296), .Y (n_4788));
MX2X1 g76054(.A (text_in_r[79] ), .B (text_in[79]), .S0 (n_672), .Y(n_3748));
NAND2X1 g75695(.A (n_3590), .B (n_1823), .Y (n_4107));
NAND2X1 g74277(.A (n_3746), .B (n_1206), .Y (n_4784));
NAND2X2 g73695(.A (n_2753), .B (n_3632), .Y (n_8379));
XOR2X1 g76159(.A (text_in_r[72] ), .B (n_23567), .Y (n_3743));
NAND2X1 g74758(.A (n_2723), .B (n_2069), .Y (n_4290));
AND2X1 g77719(.A (n_15674), .B (n_282), .Y (n_3739));
OR2X1 g73635(.A (n_2488), .B (n_3736), .Y (n_5795));
AND2X1 g78079(.A (n_27202), .B (n_3735), .Y (n_4492));
NAND2X2 g74258(.A (n_2680), .B (n_28481), .Y (n_4668));
INVX1 g74262(.A (n_2480), .Y (n_5733));
NOR2X1 g74753(.A (n_2991), .B (n_3920), .Y (n_4291));
MX2X1 g75968(.A (text_in_r[1] ), .B (text_in[1]), .S0 (n_600), .Y(n_3732));
NAND2X1 g75085(.A (n_2400), .B (n_7537), .Y (n_4247));
INVX1 g74254(.A (n_4513), .Y (n_4771));
INVX2 g75073(.A (n_4500), .Y (n_6232));
INVX2 g77245(.A (n_3729), .Y (n_4770));
INVX1 g75740(.A (n_3728), .Y (n_6135));
INVX1 g75061(.A (n_4612), .Y (n_4986));
NOR2X1 g78112(.A (n_16787), .B (n_62), .Y (n_4930));
NOR2X1 g78237(.A (n_9467), .B (n_3264), .Y (n_3725));
INVX1 g77662(.A (n_3723), .Y (n_4764));
NAND4X1 g72347(.A (n_1176), .B (dcnt[0] ), .C (n_3721), .D (n_77),.Y (n_3722));
INVX4 g81037(.A (n_27128), .Y (n_11576));
INVX2 g73656(.A (n_2809), .Y (n_4435));
NAND2X1 g78053(.A (n_6997), .B (n_1230), .Y (n_4428));
INVX1 g77310(.A (n_4108), .Y (n_5457));
INVX1 g77699(.A (n_3717), .Y (n_3718));
INVX1 g73640(.A (n_3715), .Y (n_3716));
NAND2X1 g76835(.A (n_28542), .B (n_7559), .Y (n_3714));
NOR2X1 g76516(.A (n_16787), .B (sa13[1] ), .Y (n_18102));
INVX1 g77186(.A (n_3710), .Y (n_4724));
INVX1 g74228(.A (n_3706), .Y (n_3707));
OR2X1 g78293(.A (n_14589), .B (n_21275), .Y (n_4851));
INVX1 g74718(.A (n_4234), .Y (n_5766));
INVX2 g73633(.A (n_2699), .Y (n_5930));
DFFX1 text_in_r_reg[57] (.CK (clk), .D (n_1763), .Q (text_in_r[57]), .QN ());
NAND2X2 g73377(.A (n_3559), .B (n_3704), .Y (n_3705));
NOR2X1 g74976(.A (n_2889), .B (n_386), .Y (n_4258));
MX2X1 g76025(.A (text_in_r[108] ), .B (text_in[108]), .S0 (n_672),.Y (n_3703));
NAND2X1 g74007(.A (n_636), .B (n_3023), .Y (n_4271));
INVX1 g77220(.A (n_3701), .Y (n_4671));
INVX1 g78219(.A (n_3700), .Y (n_4748));
NAND2X1 g74598(.A (n_27990), .B (n_2643), .Y (n_3699));
INVX1 g73600(.A (n_2794), .Y (n_4727));
INVX1 g77114(.A (n_3698), .Y (n_4045));
INVX2 g77210(.A (n_4635), .Y (n_3697));
NOR2X1 g74210(.A (n_2536), .B (n_5924), .Y (n_4730));
AND2X1 g77682(.A (n_3696), .B (n_3695), .Y (n_4744));
INVX1 g78209(.A (n_3694), .Y (n_5148));
INVX1 g73317(.A (n_3692), .Y (n_6004));
INVX1 g73619(.A (n_3691), .Y (n_4441));
INVX1 g77071(.A (n_4169), .Y (n_3689));
NAND2X1 g74927(.A (n_2424), .B (n_28744), .Y (n_4268));
INVX1 g77204(.A (n_5985), .Y (n_3686));
NAND2X1 g75282(.A (n_2743), .B (n_827), .Y (n_6040));
INVX1 g74923(.A (n_3682), .Y (n_3683));
INVX1 g74915(.A (n_2595), .Y (n_4740));
OR2X1 g75634(.A (n_1571), .B (n_3307), .Y (n_4178));
NAND2X2 g74911(.A (n_2684), .B (n_28351), .Y (n_4970));
INVX1 g77677(.A (n_4414), .Y (n_4015));
MX2X1 g76073(.A (text_in_r[34] ), .B (text_in[34]), .S0 (n_672), .Y(n_3680));
DFFX1 text_in_r_reg[95] (.CK (clk), .D (n_1648), .Q (text_in_r[95]), .QN ());
INVX1 g73446(.A (n_3679), .Y (n_4559));
NAND2X1 g74606(.A (n_2596), .B (n_5186), .Y (n_5692));
NOR2X1 g73603(.A (n_2865), .B (n_6008), .Y (n_3678));
NAND2X1 g74849(.A (n_16976), .B (n_1325), .Y (n_3677));
NAND2X1 g74837(.A (n_2827), .B (n_490), .Y (n_5823));
OR2X1 g74851(.A (n_6817), .B (n_9682), .Y (n_3676));
INVX1 g73594(.A (n_2803), .Y (n_4444));
DFFX1 text_in_r_reg[124] (.CK (clk), .D (n_1840), .Q(text_in_r[124] ), .QN ());
INVX1 g77671(.A (n_3673), .Y (n_5386));
NOR2X1 g74205(.A (n_1886), .B (n_28744), .Y (n_4369));
INVX1 g74823(.A (n_3672), .Y (n_4855));
INVX1 g76494(.A (n_3671), .Y (n_4095));
NOR2X1 g77504(.A (n_5924), .B (n_1424), .Y (n_3669));
AND2X1 g76489(.A (n_3667), .B (n_4357), .Y (n_3668));
INVX1 g77196(.A (n_3666), .Y (n_4039));
INVX1 g77172(.A (n_4280), .Y (n_5154));
INVX1 g77198(.A (n_3687), .Y (n_3664));
MX2X1 g76066(.A (text_in_r[97] ), .B (text_in[97]), .S0 (n_672), .Y(n_3663));
NAND2X1 g74012(.A (n_2401), .B (n_7182), .Y (n_4396));
MX2X1 g76003(.A (text_in_r[51] ), .B (text_in[51]), .S0 (n_619), .Y(n_3660));
INVX1 g78082(.A (n_27160), .Y (n_4529));
INVX1 g74497(.A (n_4786), .Y (n_3982));
NAND2X1 g74741(.A (n_883), .B (n_218), .Y (n_4769));
INVX1 g76608(.A (n_3653), .Y (n_3654));
NAND2X1 g75166(.A (n_3820), .B (n_2298), .Y (n_3652));
MX2X1 g75999(.A (text_in_r[19] ), .B (text_in[19]), .S0 (ld), .Y(n_3650));
NAND2X2 g74188(.A (n_2638), .B (n_4364), .Y (n_3646));
NAND2X1 g74131(.A (n_538), .B (n_28357), .Y (n_4669));
NAND2X2 g73470(.A (n_3643), .B (n_3338), .Y (n_3644));
MX2X1 g76092(.A (text_in_r[78] ), .B (text_in[78]), .S0 (n_672), .Y(n_3642));
NOR2X1 g74715(.A (n_3640), .B (n_1430), .Y (n_6148));
MX2X1 g75998(.A (text_in_r[9] ), .B (text_in[9]), .S0 (n_3340), .Y(n_3639));
MX2X1 g76093(.A (text_in_r[110] ), .B (text_in[110]), .S0 (n_600),.Y (n_3636));
NAND2X1 g74705(.A (n_999), .B (n_3643), .Y (n_4297));
DFFX1 text_in_r_reg[115] (.CK (clk), .D (n_2060), .Q(text_in_r[115] ), .QN ());
INVX1 g75415(.A (n_4533), .Y (n_5777));
NAND2X1 g75749(.A (n_8342), .B (n_2236), .Y (n_3634));
NAND2X1 g73536(.A (n_27072), .B (n_3632), .Y (n_3633));
MX2X1 g76070(.A (text_in_r[12] ), .B (text_in[12]), .S0 (n_672), .Y(n_3631));
INVX1 g76771(.A (n_3630), .Y (n_12784));
OR2X1 g73576(.A (n_2611), .B (n_6005), .Y (n_4859));
MX2X1 g76031(.A (text_in_r[82] ), .B (text_in[82]), .S0 (n_600), .Y(n_3625));
INVX1 g74708(.A (n_2733), .Y (n_4701));
MX2X1 g76065(.A (text_in_r[104] ), .B (text_in[104]), .S0 (ld), .Y(n_3624));
INVX1 g78302(.A (n_3622), .Y (n_4980));
MX2X1 g76067(.A (text_in_r[86] ), .B (text_in[86]), .S0 (n_619), .Y(n_3621));
NOR2X1 g74175(.A (n_2349), .B (n_5413), .Y (n_6058));
MX2X1 g76079(.A (text_in_r[68] ), .B (text_in[68]), .S0 (n_600), .Y(n_3619));
DFFX1 text_in_r_reg[98] (.CK (clk), .D (n_1895), .Q (text_in_r[98]), .QN ());
MX2X1 g75981(.A (text_in_r[118] ), .B (text_in[118]), .S0 (n_672),.Y (n_3617));
NAND2X1 g74700(.A (n_3615), .B (n_9257), .Y (n_3616));
INVX1 g76739(.A (n_4115), .Y (n_4072));
MX2X1 g75980(.A (text_in_r[35] ), .B (text_in[35]), .S0 (n_600), .Y(n_3613));
INVX1 g73507(.A (n_3610), .Y (n_4486));
NOR2X1 g68120(.A (n_1827), .B (u0_r0_rcnt[0] ), .Y (n_3609));
INVX1 g74692(.A (n_3604), .Y (n_3605));
MX2X1 g76000(.A (text_in_r[107] ), .B (text_in[107]), .S0 (n_600),.Y (n_3603));
INVX1 g77044(.A (n_4388), .Y (n_5225));
INVX2 g76761(.A (n_2510), .Y (n_4070));
OR2X1 g71257(.A (n_3600), .B (n_3599), .Y (n_3601));
NAND2X1 g77581(.A (n_28757), .B (n_3597), .Y (n_4018));
INVX1 g80435(.A (w3[1] ), .Y (n_6400));
NAND2X1 g78195(.A (n_1206), .B (n_8918), .Y (n_4829));
INVX1 g76674(.A (n_3594), .Y (n_5834));
INVX4 g76445(.A (n_28153), .Y (n_5612));
NOR2X1 g74567(.A (n_4364), .B (n_2774), .Y (n_6011));
INVX1 g76442(.A (n_3467), .Y (n_8317));
NAND2X1 g73476(.A (n_3590), .B (n_6252), .Y (n_5716));
INVX1 g74018(.A (n_3589), .Y (n_7032));
INVX1 g77577(.A (n_4422), .Y (n_3588));
MX2X1 g76057(.A (text_in_r[40] ), .B (text_in[40]), .S0 (n_600), .Y(n_3587));
NAND2X2 g74226(.A (n_3585), .B (n_867), .Y (n_4650));
NAND2X1 g75755(.A (n_3234), .B (n_2514), .Y (n_3582));
NOR2X1 g78201(.A (n_29074), .B (n_6462), .Y (n_3581));
NAND2X1 g74527(.A (n_3246), .B (n_5005), .Y (n_5764));
INVX1 g77865(.A (n_3579), .Y (n_4966));
DFFX1 text_in_r_reg[31] (.CK (clk), .D (n_2212), .Q (text_in_r[31]), .QN ());
NAND2X1 g74504(.A (n_5546), .B (n_9410), .Y (n_3577));
INVX1 g77834(.A (n_12134), .Y (n_4006));
INVX1 g78150(.A (n_4974), .Y (n_11694));
INVX1 g76427(.A (n_3575), .Y (n_4776));
NAND2X1 g73383(.A (n_2278), .B (n_5660), .Y (n_3574));
NAND2X1 g74473(.A (n_3573), .B (n_4490), .Y (n_5719));
NOR2X1 g74471(.A (n_2787), .B (n_4490), .Y (n_6166));
NAND2X1 g74465(.A (n_3807), .B (n_3569), .Y (n_3571));
DFFX1 text_in_r_reg[122] (.CK (clk), .D (n_1588), .Q(text_in_r[122] ), .QN ());
INVX1 g76420(.A (ld_r), .Y (n_6230));
NAND2X1 g74044(.A (n_755), .B (n_3566), .Y (n_3567));
NAND2X1 g74170(.A (n_27220), .B (n_636), .Y (n_6099));
MX2X1 g76015(.A (text_in_r[14] ), .B (text_in[14]), .S0 (n_619), .Y(n_3565));
NAND2X1 g75456(.A (n_3346), .B (n_3560), .Y (n_4202));
NAND2X1 g74389(.A (n_2916), .B (n_3559), .Y (n_4899));
NAND2X1 g76434(.A (n_27202), .B (n_2798), .Y (n_3557));
NAND2X1 g74944(.A (n_2049), .B (n_3920), .Y (n_4025));
DFFX1 text_in_r_reg[119] (.CK (clk), .D (n_1955), .Q(text_in_r[119] ), .QN ());
NOR2X1 g73478(.A (n_2330), .B (n_8865), .Y (n_4458));
AND2X1 g78178(.A (n_196), .B (n_14142), .Y (n_19692));
NOR2X1 g77123(.A (n_9486), .B (n_1347), .Y (n_7932));
INVX1 g74119(.A (n_3551), .Y (n_3552));
NAND2X1 g73432(.A (n_2714), .B (n_28464), .Y (n_4467));
INVX1 g76707(.A (n_3830), .Y (n_4659));
INVX1 g81242(.A (n_21520), .Y (n_3546));
NOR2X1 g62220(.A (n_6289), .B (n_25052), .Y (n_3545));
MX2X1 g76063(.A (text_in_r[56] ), .B (text_in[56]), .S0 (n_600), .Y(n_3543));
XOR2X1 g76121(.A (text_in_r[89] ), .B (w1[25] ), .Y (n_3541));
NAND2X2 g75088(.A (n_3536), .B (n_3283), .Y (n_5912));
NAND2X1 g74271(.A (n_3535), .B (n_3534), .Y (n_5741));
CLKBUFX1 g76384(.A (ld_r), .Y (n_4622));
NAND2X1 g75428(.A (n_4217), .B (n_15568), .Y (n_3533));
OR2X1 g77518(.A (n_3696), .B (n_9118), .Y (n_3532));
INVX1 g76570(.A (n_4866), .Y (n_4893));
DFFX1 text_in_r_reg[102] (.CK (clk), .D (n_1507), .Q(text_in_r[102] ), .QN ());
NAND2X1 g75418(.A (n_2334), .B (n_5005), .Y (n_4315));
INVX1 g81752(.A (n_7586), .Y (n_3530));
INVX1 g77002(.A (n_4014), .Y (n_5383));
NAND2X1 g74167(.A (n_1819), .B (n_29155), .Y (n_4688));
MX2X1 g75993(.A (text_in_r[88] ), .B (text_in[88]), .S0 (n_600), .Y(n_3521));
INVX2 g75149(.A (n_2662), .Y (n_4636));
MX2X1 g75972(.A (text_in_r[60] ), .B (text_in[60]), .S0 (n_600), .Y(n_3519));
OR2X1 g74125(.A (n_2053), .B (n_3920), .Y (n_4377));
NOR2X1 g74093(.A (n_3517), .B (n_5422), .Y (n_3518));
INVX1 g73512(.A (n_2481), .Y (n_4692));
NOR2X1 g77318(.A (n_17912), .B (sa33[1] ), .Y (n_18119));
INVX1 g77927(.A (n_3513), .Y (n_3514));
INVX1 g77065(.A (n_3522), .Y (n_12268));
NAND2X1 g76717(.A (n_3512), .B (n_3511), .Y (n_4076));
NAND2X1 g78231(.A (n_6043), .B (n_2319), .Y (n_4753));
DFFX1 text_in_r_reg[76] (.CK (clk), .D (n_1915), .Q (text_in_r[76]), .QN ());
INVX1 g77277(.A (n_5138), .Y (n_3506));
NAND2X1 g74041(.A (n_2387), .B (n_28463), .Y (n_4658));
NAND2X1 g74033(.A (n_27673), .B (n_27674), .Y (n_3505));
MX2X1 g76058(.A (text_in_r[45] ), .B (text_in[45]), .S0 (n_600), .Y(n_3504));
INVX1 g78915(.A (n_8816), .Y (n_3503));
INVX1 g73999(.A (n_2468), .Y (n_4203));
DFFX1 text_in_r_reg[113] (.CK (clk), .D (n_1528), .Q(text_in_r[113] ), .QN ());
INVX1 g77232(.A (n_3500), .Y (n_3501));
INVX1 g73386(.A (n_3499), .Y (n_6015));
NAND2X1 g75816(.A (n_4194), .B (n_2492), .Y (n_3498));
NAND2X1 g73932(.A (n_3491), .B (n_7658), .Y (n_13219));
NAND2X2 g73486(.A (n_2351), .B (n_27371), .Y (n_4606));
MX2X1 g75991(.A (text_in_r[92] ), .B (text_in[92]), .S0 (n_600), .Y(n_3495));
NOR2X1 g76424(.A (n_3493), .B (n_29297), .Y (n_3494));
NAND2X1 g73905(.A (n_3491), .B (n_3307), .Y (n_16954));
NAND2X1 g73364(.A (n_3489), .B (n_3038), .Y (n_9220));
INVX1 g76846(.A (n_2603), .Y (n_4772));
NAND2X1 g77362(.A (w3[1] ), .B (n_16480), .Y (n_11126));
INVX1 g77055(.A (n_3965), .Y (n_3488));
NOR2X1 g70173(.A (n_2480), .B (n_5422), .Y (n_7661));
NAND2X1 g73809(.A (n_2635), .B (n_5381), .Y (n_8719));
NAND2X1 g73390(.A (n_3590), .B (n_14484), .Y (n_4554));
MX2X1 g76080(.A (text_in_r[81] ), .B (text_in[81]), .S0 (n_672), .Y(n_3485));
INVX1 g78138(.A (n_19961), .Y (n_3483));
NAND2X1 g75321(.A (n_3746), .B (n_1823), .Y (n_28866));
INVX1 g73356(.A (n_2623), .Y (n_4550));
NOR2X1 g73801(.A (n_3482), .B (n_5005), .Y (n_4418));
INVX1 g73784(.A (n_13183), .Y (n_3480));
DFFX1 text_in_r_reg[94] (.CK (clk), .D (n_1752), .Q (text_in_r[94]), .QN ());
AND2X1 g73723(.A (n_2332), .B (n_5422), .Y (n_7617));
INVX1 g73707(.A (n_3475), .Y (n_6025));
MX2X1 g76049(.A (text_in_r[55] ), .B (text_in[55]), .S0 (n_672), .Y(n_3466));
NAND2X2 g73685(.A (n_3465), .B (n_3464), .Y (n_5616));
INVX1 g73678(.A (n_3463), .Y (n_4430));
INVX1 g73346(.A (n_3457), .Y (n_4478));
INVX1 g76856(.A (n_3459), .Y (n_3460));
INVX1 g73650(.A (n_3455), .Y (n_3456));
NOR2X1 g73662(.A (n_3640), .B (n_6352), .Y (n_4433));
NAND2X1 g78236(.A (n_2319), .B (n_2318), .Y (n_3454));
INVX1 g76866(.A (n_2327), .Y (n_7126));
DFFX1 text_in_r_reg[62] (.CK (clk), .D (n_1851), .Q (text_in_r[62]), .QN ());
NAND2X1 g74536(.A (n_1995), .B (n_519), .Y (n_4672));
INVX1 g82279(.A (n_27493), .Y (n_17104));
NAND2X1 g73334(.A (n_3448), .B (n_6021), .Y (n_3449));
DFFX1 text_in_r_reg[48] (.CK (clk), .D (n_1805), .Q (text_in_r[48]), .QN ());
NOR2X1 g75142(.A (n_2446), .B (n_2487), .Y (n_5895));
INVX2 g74153(.A (n_4401), .Y (n_5944));
INVX2 g74664(.A (n_26602), .Y (n_4301));
INVX2 g73573(.A (n_2962), .Y (n_5015));
INVX1 g73567(.A (n_3444), .Y (n_5968));
INVX1 g73516(.A (n_3437), .Y (n_3438));
NOR2X1 g71003(.A (n_2580), .B (n_28771), .Y (n_7241));
MX2X1 g76083(.A (text_in_r[46] ), .B (text_in[46]), .S0 (n_600), .Y(n_3433));
INVX1 g73455(.A (n_2856), .Y (n_4462));
NAND2X1 g71181(.A (n_3365), .B (n_12169), .Y (n_7603));
INVX1 g73412(.A (n_2574), .Y (n_4471));
MX2X1 g76089(.A (text_in_r[63] ), .B (text_in[63]), .S0 (ld), .Y(n_3429));
NAND2X1 g75532(.A (n_3427), .B (n_3632), .Y (n_11067));
INVX1 g77473(.A (n_3425), .Y (n_5441));
NOR2X1 g76520(.A (n_9410), .B (sa31[1] ), .Y (n_18889));
NOR2X1 g73490(.A (n_3422), .B (n_4364), .Y (n_4456));
INVX1 g78068(.A (n_3473), .Y (n_3421));
AND2X1 g75748(.A (n_3420), .B (n_1376), .Y (n_4561));
XOR2X1 g76114(.A (text_in_r[93] ), .B (n_645), .Y (n_3419));
MX2X1 g76039(.A (text_in_r[74] ), .B (text_in[74]), .S0 (n_672), .Y(n_3418));
INVX2 g73815(.A (n_3417), .Y (n_4539));
INVX1 g76466(.A (n_3228), .Y (n_15919));
NOR2X1 g71477(.A (n_4364), .B (n_2823), .Y (n_7798));
INVX1 g80760(.A (n_9442), .Y (n_4755));
DFFX1 text_in_r_reg[27] (.CK (clk), .D (n_2176), .Q (text_in_r[27]), .QN ());
NAND2X1 g74668(.A (n_4544), .B (n_5530), .Y (n_3411));
MX2X1 g76091(.A (text_in_r[17] ), .B (text_in[17]), .S0 (ld), .Y(n_3410));
INVX1 g81117(.A (n_19857), .Y (n_17474));
MX2X1 g76077(.A (text_in_r[20] ), .B (text_in[20]), .S0 (n_672), .Y(n_3409));
NAND2X1 g71625(.A (n_9755), .B (n_3600), .Y (n_3407));
MX2X1 g76032(.A (text_in_r[91] ), .B (text_in[91]), .S0 (n_619), .Y(n_3406));
INVX1 g76698(.A (n_2811), .Y (n_4077));
MX2X1 g75976(.A (text_in_r[29] ), .B (text_in[29]), .S0 (n_600), .Y(n_3405));
DFFX1 text_in_r_reg[109] (.CK (clk), .D (n_1734), .Q(text_in_r[109] ), .QN ());
MX2X1 g76036(.A (text_in_r[69] ), .B (text_in[69]), .S0 (n_600), .Y(n_3404));
MX2X1 g76088(.A (text_in_r[75] ), .B (text_in[75]), .S0 (n_600), .Y(n_3403));
MX2X1 g76035(.A (text_in_r[59] ), .B (text_in[59]), .S0 (n_672), .Y(n_3402));
XOR2X1 g76323(.A (text_in_r[0] ), .B (n_21687), .Y (n_3401));
MX2X1 g76024(.A (text_in_r[80] ), .B (text_in[80]), .S0 (ld), .Y(n_3399));
NOR2X1 g71891(.A (n_2335), .B (n_9368), .Y (n_3398));
INVX1 g78242(.A (n_4760), .Y (n_4521));
NOR2X1 g71997(.A (n_2804), .B (n_4598), .Y (n_3396));
MX2X1 g76033(.A (text_in_r[84] ), .B (text_in[84]), .S0 (n_619), .Y(n_3395));
INVX1 g81725(.A (n_7947), .Y (n_3394));
XOR2X1 g76286(.A (text_in_r[64] ), .B (n_1958), .Y (n_3393));
INVX1 g76451(.A (n_4595), .Y (n_6260));
NAND2X1 g72173(.A (n_2664), .B (n_3599), .Y (n_6134));
NOR2X1 g75490(.A (n_4825), .B (n_25808), .Y (n_4196));
MX2X1 g76034(.A (text_in_r[105] ), .B (text_in[105]), .S0 (ld), .Y(n_3390));
INVX1 g76455(.A (n_3388), .Y (n_4100));
NAND2X1 g75723(.A (n_2755), .B (n_3284), .Y (n_5774));
NAND2X1 g75480(.A (n_3536), .B (n_3307), .Y (n_4145));
INVX1 g78117(.A (n_3386), .Y (n_18074));
INVX1 g73871(.A (n_3385), .Y (n_4413));
OR2X1 g72569(.A (n_2892), .B (n_3318), .Y (n_13479));
INVX2 g77586(.A (n_3384), .Y (n_5410));
DFFX1 text_in_r_reg[117] (.CK (clk), .D (n_1891), .Q(text_in_r[117] ), .QN ());
NOR2X1 g72640(.A (n_2563), .B (n_4721), .Y (n_3381));
MX2X1 g76016(.A (text_in_r[30] ), .B (text_in[30]), .S0 (n_672), .Y(n_3380));
MX2X1 g75985(.A (text_in_r[99] ), .B (text_in[99]), .S0 (n_672), .Y(n_3375));
NAND2X2 g75116(.A (n_3373), .B (n_28792), .Y (n_5135));
INVX1 g75844(.A (n_3372), .Y (n_5835));
NAND2X1 g75768(.A (n_1920), .B (n_29158), .Y (n_4167));
INVX1 g82486(.A (n_2674), .Y (n_6554));
DFFX1 u0_r0_rcnt_reg[0] (.CK (clk), .D (n_2710), .Q (u0_r0_rcnt[0]), .QN ());
MX2X1 g75992(.A (text_in_r[8] ), .B (text_in[8]), .S0 (n_600), .Y(n_3367));
NAND2X1 g70839(.A (n_3365), .B (n_3920), .Y (n_3366));
NOR2X1 g75772(.A (n_3096), .B (n_677), .Y (n_4166));
MX2X1 g75975(.A (text_in_r[26] ), .B (text_in[26]), .S0 (n_600), .Y(n_3362));
MX2X1 g76023(.A (text_in_r[10] ), .B (text_in[10]), .S0 (n_672), .Y(n_3358));
NAND2X2 g75102(.A (n_27072), .B (n_29155), .Y (n_29140));
MX2X1 g76022(.A (text_in_r[77] ), .B (text_in[77]), .S0 (n_3340), .Y(n_3354));
NAND2X2 g73407(.A (n_3590), .B (n_2383), .Y (n_4642));
INVX1 g73420(.A (n_3353), .Y (n_7169));
NOR2X1 g73453(.A (n_8865), .B (n_29119), .Y (n_4463));
NOR2X1 g73465(.A (n_2613), .B (n_3301), .Y (n_4798));
NOR2X1 g73483(.A (n_6043), .B (n_4973), .Y (n_4457));
INVX2 g73613(.A (n_2739), .Y (n_4741));
INVX1 g73625(.A (n_3350), .Y (n_4439));
INVX2 g73645(.A (n_3715), .Y (n_4757));
INVX2 g73669(.A (n_2824), .Y (n_4767));
INVX1 g73688(.A (n_3469), .Y (n_3349));
NOR2X1 g74782(.A (n_2911), .B (n_28733), .Y (n_4801));
OR2X1 g73717(.A (n_2930), .B (n_4882), .Y (n_6062));
NAND2X1 g73731(.A (n_2568), .B (n_3348), .Y (n_4841));
MX2X1 g76019(.A (text_in_r[39] ), .B (text_in[39]), .S0 (n_600), .Y(n_3347));
NAND2X2 g73782(.A (n_3187), .B (n_28733), .Y (n_4886));
OR2X1 g73783(.A (n_2671), .B (n_9388), .Y (n_7215));
NAND2X1 g73865(.A (n_28340), .B (n_8865), .Y (n_9844));
NAND2X1 g73895(.A (n_3346), .B (n_4522), .Y (n_5832));
INVX1 g73909(.A (n_3345), .Y (n_3991));
NAND2X1 g73923(.A (n_3346), .B (n_1627), .Y (n_4007));
MX2X1 g76017(.A (text_in_r[7] ), .B (text_in[7]), .S0 (ld), .Y(n_3343));
INVX2 g73936(.A (n_3342), .Y (n_4407));
NOR2X1 g73380(.A (n_2594), .B (n_4865), .Y (n_4475));
MX2X1 g76021(.A (text_in_r[121] ), .B (text_in[121]), .S0 (n_3340),.Y (n_3341));
NAND2X1 g74001(.A (n_2128), .B (n_10255), .Y (n_3339));
NOR2X1 g74081(.A (n_3338), .B (n_2392), .Y (n_6277));
NAND2X1 g74123(.A (n_2850), .B (n_6021), .Y (n_4379));
INVX1 g74137(.A (n_2796), .Y (n_4778));
NOR2X1 g74151(.A (n_28488), .B (n_5381), .Y (n_3336));
INVX1 g74171(.A (n_3334), .Y (n_5997));
AND2X1 g74283(.A (n_2852), .B (n_3307), .Y (n_7084));
NOR2X1 g77064(.A (n_3512), .B (n_9084), .Y (n_3331));
NOR2X1 g74307(.A (n_6805), .B (n_2772), .Y (n_3330));
NAND2X1 g74337(.A (n_2696), .B (n_4961), .Y (n_3329));
MX2X1 g76011(.A (text_in_r[42] ), .B (text_in[42]), .S0 (ld), .Y(n_3328));
NAND2X2 g74343(.A (n_3297), .B (n_3327), .Y (n_4872));
INVX1 g74359(.A (n_4552), .Y (n_3326));
DFFX1 text_in_r_reg[21] (.CK (clk), .D (n_1698), .Q (text_in_r[21]), .QN ());
NOR2X1 g74439(.A (n_29360), .B (n_3807), .Y (n_3323));
NAND2X2 g74449(.A (n_1923), .B (n_28351), .Y (n_4950));
NAND2X1 g74495(.A (n_3322), .B (n_1568), .Y (n_3981));
NAND2X1 g74503(.A (n_3252), .B (n_9500), .Y (n_3992));
NOR2X1 g74513(.A (n_6620), .B (n_3319), .Y (n_4320));
OR2X1 g74539(.A (n_2741), .B (n_3318), .Y (n_6018));
INVX1 g74543(.A (n_3316), .Y (n_3317));
NAND2X1 g74557(.A (n_6043), .B (n_3314), .Y (n_5867));
NAND2X2 g74565(.A (n_3267), .B (n_28463), .Y (n_5966));
NAND2X1 g74575(.A (n_3091), .B (n_27990), .Y (n_5787));
INVX1 g74621(.A (n_3312), .Y (n_4366));
AND2X1 g74679(.A (n_3310), .B (n_827), .Y (n_5845));
AND2X1 g74681(.A (n_2049), .B (n_9057), .Y (n_4345));
NOR2X1 g74683(.A (n_2372), .B (n_3307), .Y (n_4000));
OR2X1 g74699(.A (n_1943), .B (n_6783), .Y (n_4678));
NOR2X1 g72535(.A (n_2464), .B (n_3820), .Y (n_3305));
NAND2X1 g74747(.A (n_4113), .B (n_2304), .Y (n_5820));
NAND2X2 g74751(.A (n_3585), .B (n_3067), .Y (n_5800));
NOR2X1 g74793(.A (n_28757), .B (n_2604), .Y (n_4811));
NAND2X1 g78017(.A (n_2960), .B (n_3695), .Y (n_4282));
OR2X1 g74886(.A (n_3303), .B (n_7182), .Y (n_3304));
OR2X1 g74946(.A (n_2969), .B (n_3301), .Y (n_3302));
MX2X1 g76059(.A (text_in_r[23] ), .B (text_in[23]), .S0 (n_600), .Y(n_3300));
NAND2X1 g73504(.A (n_2820), .B (n_10315), .Y (n_9236));
NAND2X1 g74603(.A (n_3297), .B (n_3296), .Y (n_5826));
NAND2X1 g75009(.A (n_28779), .B (n_28152), .Y (n_4134));
MX2X1 g75977(.A (text_in_r[58] ), .B (text_in[58]), .S0 (n_600), .Y(n_3295));
INVX1 g73322(.A (n_3294), .Y (n_4543));
INVX1 g75050(.A (n_3726), .Y (n_5925));
NAND2X1 g75057(.A (n_2755), .B (n_386), .Y (n_4269));
MX2X1 g76069(.A (text_in_r[6] ), .B (text_in[6]), .S0 (n_672), .Y(n_3292));
NOR2X1 g75117(.A (n_1938), .B (n_5817), .Y (n_3291));
MX2X1 g76037(.A (text_in_r[13] ), .B (text_in[13]), .S0 (n_672), .Y(n_3290));
INVX1 g75137(.A (n_4504), .Y (n_4567));
NAND2X1 g75548(.A (n_6252), .B (n_3288), .Y (n_3289));
AOI21X1 g63749(.A0 (n_1693), .A1 (dcnt[3] ), .B0 (n_6301), .Y(n_3286));
NAND2X1 g75265(.A (n_2766), .B (n_4721), .Y (n_5705));
NAND2X2 g75278(.A (n_3285), .B (n_3284), .Y (n_5047));
NAND2X1 g75299(.A (n_2628), .B (n_3283), .Y (n_5435));
OR2X1 g75301(.A (n_3281), .B (n_5131), .Y (n_3282));
OR2X1 g75305(.A (n_2678), .B (n_3736), .Y (n_4017));
NAND2X2 g75048(.A (n_671), .B (n_2383), .Y (n_4839));
OR2X1 g77996(.A (n_11400), .B (n_20018), .Y (n_18617));
INVX1 g75353(.A (n_2426), .Y (n_4853));
NAND2X1 g75365(.A (n_1284), .B (n_6008), .Y (n_3279));
INVX1 g75425(.A (n_3276), .Y (n_3277));
NAND2X2 g74590(.A (n_28872), .B (n_6021), .Y (n_4307));
INVX1 g75483(.A (n_3273), .Y (n_4792));
NAND2X1 g75394(.A (n_1997), .B (n_379), .Y (n_4190));
NAND2X2 g74689(.A (n_3128), .B (n_26893), .Y (n_5915));
NOR2X1 g77093(.A (n_11489), .B (sa30[1] ), .Y (n_17003));
INVX1 g75557(.A (n_3869), .Y (n_3268));
NAND2X1 g75571(.A (n_3267), .B (n_28464), .Y (n_5101));
AND2X1 g75579(.A (n_1325), .B (n_3264), .Y (n_3266));
OR2X1 g75684(.A (n_6827), .B (n_1065), .Y (n_3261));
NOR2X1 g74582(.A (n_27904), .B (n_2402), .Y (n_4308));
NAND2X1 g75651(.A (n_2266), .B (n_10315), .Y (n_3260));
OR2X1 g75659(.A (n_4208), .B (n_14630), .Y (n_3258));
INVX2 g77028(.A (n_3195), .Y (n_3257));
NAND2X1 g75675(.A (n_27437), .B (n_2943), .Y (n_3256));
NOR2X1 g75678(.A (n_1491), .B (n_5413), .Y (n_5892));
INVX1 g75690(.A (n_3253), .Y (n_3254));
INVX2 g75386(.A (n_3250), .Y (n_4163));
NAND4X1 g69309(.A (n_9388), .B (n_2492), .C (n_1431), .D (n_2099), .Y(n_6107));
NAND2X1 g75024(.A (n_26887), .B (n_2919), .Y (n_3248));
NAND2X1 g73972(.A (n_3247), .B (n_6133), .Y (n_4403));
NAND2X2 g75812(.A (n_3246), .B (n_2993), .Y (n_5988));
NAND2X2 g75803(.A (n_28312), .B (n_3246), .Y (n_5123));
XOR2X1 g62027(.A (u0_r0_rcnt[3] ), .B (n_1205), .Y (n_6286));
INVX1 g75825(.A (n_4132), .Y (n_5810));
MX2X1 g76090(.A (text_in_r[85] ), .B (text_in[85]), .S0 (n_672), .Y(n_3245));
INVX1 g79717(.A (n_26271), .Y (n_16974));
XOR2X1 g76301(.A (text_in_r[75] ), .B (n_546), .Y (n_3244));
NAND2X1 g75914(.A (n_6871), .B (n_2950), .Y (n_14157));
MX2X1 g75966(.A (text_in_r[15] ), .B (text_in[15]), .S0 (n_600), .Y(n_3242));
INVX1 g75376(.A (n_3241), .Y (n_4215));
INVX1 g76642(.A (n_3240), .Y (n_9415));
NAND2X1 g75677(.A (n_3267), .B (n_5660), .Y (n_5841));
INVX1 g74570(.A (n_3237), .Y (n_4312));
MX2X1 g75983(.A (text_in_r[33] ), .B (text_in[33]), .S0 (n_600), .Y(n_3236));
INVX1 g77966(.A (n_3235), .Y (n_4142));
NAND2X1 g75012(.A (n_2265), .B (n_3234), .Y (n_4255));
NOR2X1 g73978(.A (n_2715), .B (n_3017), .Y (n_3232));
INVX1 g78655(.A (n_3612), .Y (n_19408));
MX2X1 g76012(.A (text_in_r[36] ), .B (text_in[36]), .S0 (n_600), .Y(n_3231));
INVX1 g77117(.A (n_3230), .Y (n_7721));
MX2X1 g76028(.A (text_in_r[0] ), .B (text_in[0]), .S0 (n_672), .Y(n_3227));
INVX1 g76637(.A (n_3225), .Y (n_3226));
MX2X1 g76009(.A (text_in_r[64] ), .B (text_in[64]), .S0 (n_672), .Y(n_3224));
MX2X1 g76043(.A (text_in_r[116] ), .B (text_in[116]), .S0 (n_672),.Y (n_3223));
INVX1 g77016(.A (n_3093), .Y (n_7194));
MX2X1 g76056(.A (text_in_r[16] ), .B (text_in[16]), .S0 (n_3340), .Y(n_3220));
MX2X1 g76062(.A (text_in_r[120] ), .B (text_in[120]), .S0 (ld), .Y(n_3219));
CLKBUFX3 g76635(.A (n_3218), .Y (n_5502));
INVX1 g75665(.A (n_4565), .Y (n_6188));
MX2X1 g76072(.A (text_in_r[49] ), .B (text_in[49]), .S0 (n_672), .Y(n_3216));
NAND2X1 g75360(.A (n_4586), .B (n_2447), .Y (n_3214));
MX2X1 g76086(.A (text_in_r[126] ), .B (text_in[126]), .S0 (n_600),.Y (n_3213));
AND2X1 g76768(.A (n_9416), .B (n_557), .Y (n_5344));
NAND2X1 g75361(.A (n_2360), .B (n_6805), .Y (n_3212));
DFFX1 text_in_r_reg[5] (.CK (clk), .D (n_2247), .Q (text_in_r[5] ),.QN ());
MX2X1 g76010(.A (text_in_r[37] ), .B (text_in[37]), .S0 (n_600), .Y(n_3210));
INVX1 g77481(.A (n_3209), .Y (n_5218));
XOR2X1 g76151(.A (n_22569), .B (w1[25] ), .Y (n_3208));
NAND2X2 g75658(.A (n_2908), .B (n_27593), .Y (n_4123));
NAND2X1 g73966(.A (n_596), .B (n_2861), .Y (n_3206));
NAND2X1 g78075(.A (n_1551), .B (n_8452), .Y (n_3203));
XOR2X1 g64033(.A (dcnt[0] ), .B (n_6301), .Y (n_3202));
XOR2X1 g76187(.A (text_in_r[61] ), .B (n_684), .Y (n_3201));
NAND2X2 g74761(.A (n_6946), .B (n_2303), .Y (n_3199));
INVX1 g77721(.A (n_4426), .Y (n_3197));
INVX1 g74998(.A (n_4525), .Y (n_6265));
NAND2X1 g74554(.A (n_28742), .B (n_2748), .Y (n_3193));
XOR2X1 g76276(.A (text_in_r[44] ), .B (w2[12] ), .Y (n_3192));
NAND2X1 g75729(.A (n_2469), .B (n_2099), .Y (n_5803));
NAND2X1 g74990(.A (n_2021), .B (n_3187), .Y (n_4109));
XOR2X1 g76313(.A (text_in_r[92] ), .B (n_398), .Y (n_3186));
XOR2X1 g76322(.A (n_1318), .B (n_2004), .Y (n_3184));
XOR2X1 g76326(.A (text_in_r[114] ), .B (w0[18] ), .Y (n_3183));
NOR2X1 g75333(.A (n_646), .B (n_3283), .Y (n_3180));
NAND2X1 g75642(.A (n_1747), .B (n_2235), .Y (n_4553));
NOR2X1 g76470(.A (n_11400), .B (sa12[1] ), .Y (n_18094));
NOR2X1 g76471(.A (n_28452), .B (n_11323), .Y (n_3177));
INVX1 g76472(.A (n_7789), .Y (n_12162));
NAND2X1 g75452(.A (n_2929), .B (n_3920), .Y (n_5694));
INVX1 g76506(.A (n_5104), .Y (n_4732));
INVX1 g76514(.A (n_3175), .Y (n_3176));
INVX1 g74547(.A (n_3174), .Y (n_4094));
NOR2X1 g76541(.A (n_28542), .B (n_8452), .Y (n_3173));
MX2X1 g76053(.A (text_in_r[61] ), .B (text_in[61]), .S0 (n_619), .Y(n_3172));
INVX1 g76545(.A (n_4176), .Y (n_3171));
INVX1 g76553(.A (n_2883), .Y (n_4894));
OR2X1 g76559(.A (n_26880), .B (n_28452), .Y (n_3170));
INVX1 g77471(.A (n_3168), .Y (n_16649));
AND2X1 g76573(.A (n_10255), .B (n_1390), .Y (n_5365));
INVX1 g76579(.A (n_3166), .Y (n_3167));
INVX2 g76581(.A (n_3165), .Y (n_6346));
INVX1 g76614(.A (n_2289), .Y (n_8759));
NAND2X1 g76619(.A (n_3493), .B (n_29225), .Y (n_3163));
NAND2X2 g74973(.A (n_4249), .B (n_3807), .Y (n_3162));
INVX1 g76625(.A (n_3161), .Y (n_6153));
NAND2X1 g74970(.A (n_3160), .B (n_4217), .Y (n_12578));
INVX1 g76649(.A (n_3159), .Y (n_4165));
AND2X1 g76655(.A (n_8560), .B (n_575), .Y (n_5212));
INVX1 g73532(.A (n_5645), .Y (n_4452));
INVX1 g76693(.A (n_15800), .Y (n_8105));
INVX1 g76700(.A (n_4318), .Y (n_6445));
INVX1 g76752(.A (n_3461), .Y (n_4681));
NOR2X1 g74289(.A (n_1954), .B (n_6462), .Y (n_5807));
INVX1 g76775(.A (n_4266), .Y (n_28595));
INVX1 g76777(.A (n_3153), .Y (n_5923));
INVX1 g73915(.A (n_2658), .Y (n_3999));
NAND2X1 g76816(.A (n_28540), .B (n_28464), .Y (n_4736));
INVX1 g76817(.A (n_4022), .Y (n_6444));
NOR2X1 g76821(.A (n_29163), .B (n_29228), .Y (n_3150));
INVX1 g76822(.A (n_7112), .Y (n_12155));
INVX1 g79351(.A (n_2102), .Y (n_14026));
INVX1 g76832(.A (n_3711), .Y (n_11916));
NAND2X1 g76839(.A (n_3512), .B (n_9084), .Y (n_3149));
INVX2 g76842(.A (n_3148), .Y (n_4773));
NOR2X1 g76858(.A (n_2164), .B (n_8467), .Y (n_3147));
INVX1 g76868(.A (n_4245), .Y (n_3145));
OR2X1 g75020(.A (n_1509), .B (n_6805), .Y (n_3142));
NOR2X1 g76903(.A (n_2081), .B (n_7485), .Y (n_3141));
NAND2X1 g74966(.A (n_26483), .B (n_27369), .Y (n_4260));
INVX1 g76962(.A (n_7213), .Y (n_9914));
CLKBUFX1 g76982(.A (n_3134), .Y (n_5316));
INVX1 g76989(.A (n_4699), .Y (n_3133));
NOR2X1 g77004(.A (n_7419), .B (n_1213), .Y (n_3132));
INVX1 g77038(.A (n_3130), .Y (n_3131));
NAND2X1 g75431(.A (n_3128), .B (n_5381), .Y (n_5878));
INVX1 g77077(.A (n_3818), .Y (n_4427));
MX2X1 g76075(.A (text_in_r[41] ), .B (text_in[41]), .S0 (n_672), .Y(n_3126));
NOR2X1 g77144(.A (n_3667), .B (n_5817), .Y (n_3125));
NAND2X1 g74961(.A (n_3121), .B (n_28141), .Y (n_3122));
INVX1 g75380(.A (n_4604), .Y (n_4213));
INVX1 g77238(.A (n_3119), .Y (n_4762));
OR2X1 g77490(.A (n_6400), .B (n_16480), .Y (n_17069));
AND2X1 g77253(.A (n_28742), .B (n_1258), .Y (n_5511));
INVX2 g81012(.A (n_1756), .Y (n_19398));
NOR2X1 g76947(.A (n_14624), .B (n_1340), .Y (n_6281));
NAND2X1 g77294(.A (n_2972), .B (n_7598), .Y (n_3112));
NAND2X1 g77926(.A (n_27124), .B (n_3108), .Y (n_4003));
INVX1 g77316(.A (n_3107), .Y (n_18100));
INVX1 g77320(.A (n_4349), .Y (n_3106));
INVX1 g80201(.A (n_2323), .Y (n_6328));
INVX1 g77330(.A (n_4126), .Y (n_3105));
INVX1 g77341(.A (n_4353), .Y (n_3104));
OR2X1 g76935(.A (w3[1] ), .B (n_12827), .Y (n_17017));
INVX2 g77366(.A (n_4438), .Y (n_4030));
NOR2X1 g77370(.A (n_488), .B (n_7598), .Y (n_3101));
INVX1 g77396(.A (n_4012), .Y (n_3097));
NOR2X1 g75622(.A (n_3096), .B (n_2318), .Y (n_8078));
INVX1 g77151(.A (n_9708), .Y (n_5155));
NAND2X2 g75621(.A (n_3091), .B (n_29153), .Y (n_5593));
DFFX1 text_in_r_reg[22] (.CK (clk), .D (n_1457), .Q (text_in_r[22]), .QN ());
MX2X1 g76050(.A (text_in_r[18] ), .B (text_in[18]), .S0 (ld), .Y(n_3089));
INVX1 g77447(.A (n_3087), .Y (n_4023));
DFFX1 text_in_r_reg[83] (.CK (clk), .D (n_1852), .Q (text_in_r[83]), .QN ());
INVX1 g77598(.A (n_4920), .Y (n_3086));
INVX1 g77611(.A (n_3085), .Y (n_6931));
INVX1 g77613(.A (n_3084), .Y (n_5665));
DFFX1 text_in_r_reg[38] (.CK (clk), .D (n_1645), .Q (text_in_r[38]), .QN ());
AND2X1 g73931(.A (n_2859), .B (n_3920), .Y (n_4408));
INVX1 g77654(.A (n_4373), .Y (n_3083));
NOR2X1 g74509(.A (n_2216), .B (n_3081), .Y (n_3082));
NAND2X1 g75833(.A (n_5005), .B (n_2336), .Y (n_3080));
AND2X1 g77720(.A (n_14155), .B (n_20102), .Y (n_9272));
INVX1 g77727(.A (n_3076), .Y (n_3077));
AND2X1 g77783(.A (n_9819), .B (n_123), .Y (n_19157));
INVX1 g77794(.A (n_4663), .Y (n_3073));
NOR2X1 g77813(.A (n_3069), .B (n_11731), .Y (n_3070));
NOR2X1 g75256(.A (n_2210), .B (n_28742), .Y (n_4222));
AND2X1 g77382(.A (n_1502), .B (n_3067), .Y (n_4027));
INVX1 g77901(.A (n_4849), .Y (n_3065));
NAND2X1 g77923(.A (n_1933), .B (n_1739), .Y (n_4034));
NAND2X1 g77963(.A (n_2044), .B (n_28357), .Y (n_4114));
MX2X1 g76008(.A (text_in_r[52] ), .B (text_in[52]), .S0 (n_672), .Y(n_3059));
INVX1 g77997(.A (n_4450), .Y (n_3055));
NOR2X1 g74483(.A (n_2095), .B (n_6191), .Y (n_3975));
INVX1 g78022(.A (n_3052), .Y (n_3053));
OR2X1 g78040(.A (n_6043), .B (n_2318), .Y (n_3050));
NAND2X1 g74578(.A (n_3285), .B (n_3807), .Y (n_4164));
INVX1 g78096(.A (n_3049), .Y (n_6486));
INVX1 g77431(.A (n_4581), .Y (n_3984));
OR2X1 g78171(.A (n_383), .B (n_9118), .Y (n_3046));
INVX1 g78223(.A (n_4159), .Y (n_3045));
MX2X1 g75978(.A (text_in_r[65] ), .B (text_in[65]), .S0 (n_600), .Y(n_3044));
DFFX1 text_in_r_reg[71] (.CK (clk), .D (n_2066), .Q (text_in_r[71]), .QN ());
INVX1 g76972(.A (n_4520), .Y (n_5171));
DFFX1 text_in_r_reg[89] (.CK (clk), .D (n_1731), .Q (text_in_r[89]), .QN ());
INVX2 g73900(.A (n_2751), .Y (n_3980));
INVX1 g73903(.A (n_3040), .Y (n_4410));
NAND2X2 g75295(.A (n_665), .B (n_3038), .Y (n_3039));
INVX1 g77425(.A (n_3041), .Y (n_3034));
INVX1 g74936(.A (n_3032), .Y (n_3033));
INVX1 g77898(.A (n_3030), .Y (n_6033));
NAND2X1 g78132(.A (n_1230), .B (n_13593), .Y (n_3029));
AND2X1 g75751(.A (n_4861), .B (n_3023), .Y (n_3024));
INVX1 g77420(.A (n_4832), .Y (n_3022));
MX2X1 g76001(.A (text_in_r[127] ), .B (text_in[127]), .S0 (n_672),.Y (n_3020));
NOR2X1 g71583(.A (n_2781), .B (n_3017), .Y (n_3018));
INVX1 g76475(.A (n_9712), .Y (n_3016));
INVX1 g73886(.A (n_2632), .Y (n_4412));
INVX1 g73538(.A (n_12870), .Y (n_4947));
INVX2 g78957(.A (n_9527), .Y (n_15655));
DFFX1 text_in_r_reg[87] (.CK (clk), .D (n_1899), .Q (text_in_r[87]), .QN ());
NAND2X1 g75605(.A (n_2901), .B (n_218), .Y (n_3993));
NOR2X1 g75737(.A (n_2792), .B (n_1627), .Y (n_3013));
AND2X1 g78263(.A (n_5922), .B (n_14866), .Y (n_5369));
INVX2 g77888(.A (n_9978), .Y (n_6847));
INVX1 g77934(.A (n_3221), .Y (n_3010));
INVX2 g76955(.A (n_3005), .Y (n_5204));
INVX1 g77882(.A (n_4055), .Y (n_4800));
NAND2X2 g74922(.A (n_3002), .B (n_3001), .Y (n_5802));
INVX8 g78474(.A (n_975), .Y (n_10389));
INVX1 g77607(.A (n_3590), .Y (n_3000));
INVX1 g80099(.A (n_2319), .Y (n_2999));
NOR2X1 g74466(.A (n_2444), .B (n_4916), .Y (n_7568));
INVX1 g77286(.A (n_2994), .Y (n_14725));
NAND2X1 g77104(.A (n_1601), .B (n_2993), .Y (n_3776));
INVX1 g77166(.A (n_2991), .Y (n_2990));
NAND2X1 g73553(.A (n_2382), .B (n_28478), .Y (n_2989));
NAND2X1 g73864(.A (n_2988), .B (n_827), .Y (n_3931));
INVX1 g77866(.A (n_1505), .Y (n_3579));
INVX1 g77395(.A (n_2346), .Y (n_25729));
INVX1 g77274(.A (n_2276), .Y (n_16006));
INVX2 g81933(.A (n_2107), .Y (n_18785));
AND2X1 g77393(.A (n_17864), .B (n_62), .Y (n_19160));
INVX1 g77306(.A (n_2880), .Y (n_8097));
BUFX3 g81118(.A (n_13804), .Y (n_19857));
NOR2X1 g73854(.A (n_1581), .B (n_28744), .Y (n_3922));
NOR2X1 g77853(.A (n_28364), .B (n_7498), .Y (n_2973));
INVX1 g81365(.A (n_16480), .Y (n_19433));
CLKBUFX1 g81753(.A (n_3696), .Y (n_7586));
NAND2X1 g77007(.A (n_1621), .B (n_1315), .Y (n_3921));
NOR2X1 g76940(.A (n_19791), .B (n_2204), .Y (n_20105));
NAND2X2 g76939(.A (n_1925), .B (n_29158), .Y (n_3903));
NAND2X1 g75826(.A (n_2738), .B (n_1947), .Y (n_4132));
NAND3X1 g73574(.A (n_25691), .B (n_2070), .C (n_2096), .Y (n_2962));
INVX1 g80137(.A (n_23422), .Y (n_5231));
AND2X1 g78033(.A (n_2319), .B (n_488), .Y (n_3836));
INVX1 g82110(.A (n_2959), .Y (n_3888));
INVX2 g76476(.A (n_2958), .Y (n_9712));
INVX1 g77639(.A (n_4928), .Y (n_11902));
XOR2X1 g76103(.A (text_in_r[103] ), .B (w0[7] ), .Y (n_2954));
INVX2 g77355(.A (n_2952), .Y (n_19226));
INVX2 g76582(.A (n_2213), .Y (n_3165));
CLKBUFX3 g77367(.A (n_3322), .Y (n_4438));
NAND2X1 g74873(.A (n_2950), .B (n_3307), .Y (n_3891));
NAND2X1 g73816(.A (n_2933), .B (n_27197), .Y (n_3417));
NAND2X1 g73339(.A (n_2691), .B (n_2656), .Y (n_2945));
NOR2X1 g75426(.A (n_2943), .B (n_27436), .Y (n_3276));
NAND2X1 g76580(.A (n_18266), .B (n_27747), .Y (n_3166));
INVX1 g79017(.A (n_3735), .Y (n_3359));
INVX1 g76922(.A (n_2937), .Y (n_2938));
CLKBUFX3 g77655(.A (n_2749), .Y (n_4373));
NOR2X1 g76681(.A (n_400), .B (n_29167), .Y (n_3874));
XOR2X1 g76335(.A (text_in_r[65] ), .B (n_1040), .Y (n_2935));
NOR2X1 g73789(.A (n_2137), .B (n_26486), .Y (n_3859));
NAND2X1 g77135(.A (n_2099), .B (n_1129), .Y (n_2934));
NAND2X1 g73785(.A (n_2933), .B (n_6185), .Y (n_13183));
NAND2X1 g76571(.A (n_2237), .B (n_28357), .Y (n_4866));
INVX1 g77919(.A (n_2930), .Y (n_5447));
NOR2X1 g73770(.A (n_1874), .B (n_218), .Y (n_2927));
INVX1 g77352(.A (n_2925), .Y (n_2926));
XOR2X1 g76179(.A (n_221), .B (w1[16] ), .Y (n_2924));
INVX1 g75027(.A (n_2923), .Y (n_3287));
NAND2X1 g77804(.A (n_1750), .B (n_1627), .Y (n_3844));
INVX1 g77342(.A (n_3246), .Y (n_4353));
NAND2X1 g77348(.A (n_2921), .B (n_2107), .Y (n_3102));
NAND2X1 g73765(.A (n_28340), .B (n_6805), .Y (n_3829));
INVX1 g76429(.A (n_3833), .Y (n_3575));
NAND2X1 g75225(.A (n_2089), .B (n_3283), .Y (n_4867));
INVX1 g77795(.A (n_2919), .Y (n_4663));
XOR2X1 g76104(.A (text_in_r[117] ), .B (n_24366), .Y (n_2918));
INVX1 g77792(.A (n_2917), .Y (n_20399));
INVX1 g77935(.A (n_3559), .Y (n_3221));
INVX1 g77331(.A (n_3285), .Y (n_4126));
INVX1 g78307(.A (n_2916), .Y (n_3827));
INVX2 g78057(.A (n_8191), .Y (n_9371));
INVX1 g77587(.A (n_2914), .Y (n_3384));
XOR2X1 g76338(.A (n_23087), .B (n_23096), .Y (n_2913));
INVX1 g77742(.A (n_2912), .Y (n_4987));
INVX1 g78303(.A (n_2911), .Y (n_3622));
INVX1 g77173(.A (n_3128), .Y (n_4280));
INVX1 g80813(.A (n_2910), .Y (n_3824));
INVX4 g79759(.A (n_2720), .Y (n_4261));
INVX2 g76957(.A (n_2908), .Y (n_3005));
NAND2X1 g76857(.A (n_1941), .B (n_1942), .Y (n_3459));
INVX1 g79240(.A (n_2905), .Y (n_9392));
INVX1 g77775(.A (n_3314), .Y (n_2902));
INVX1 g78297(.A (n_1985), .Y (n_4158));
CLKBUFX1 g77322(.A (n_2901), .Y (n_4349));
INVX1 g76883(.A (n_2900), .Y (n_12571));
NOR2X1 g77317(.A (n_13083), .B (w3[9] ), .Y (n_3107));
XOR2X1 g76219(.A (n_1004), .B (n_23545), .Y (n_2894));
INVX1 g77762(.A (n_3187), .Y (n_3805));
NOR2X1 g73451(.A (n_2145), .B (n_1627), .Y (n_3814));
CLKBUFX3 g80657(.A (n_2891), .Y (n_7543));
INVX1 g77314(.A (n_2889), .Y (n_2890));
INVX1 g75323(.A (n_3600), .Y (n_2886));
INVX1 g76564(.A (n_2394), .Y (n_14548));
NOR2X1 g73564(.A (n_2343), .B (n_29116), .Y (n_2884));
NOR2X1 g76554(.A (n_1396), .B (n_1627), .Y (n_2883));
INVX1 g77307(.A (n_2880), .Y (n_2881));
INVX1 g78283(.A (n_3643), .Y (n_2878));
AND2X1 g77753(.A (n_28686), .B (n_21242), .Y (n_16103));
INVX1 g77756(.A (n_2875), .Y (n_3796));
INVX1 g76885(.A (n_2900), .Y (n_2872));
NAND2X2 g77305(.A (n_1717), .B (n_28423), .Y (n_15812));
INVX1 g79678(.A (n_2870), .Y (n_6335));
NAND2X1 g77298(.A (n_1792), .B (n_11253), .Y (n_3777));
XOR2X1 g76318(.A (text_in_r[126] ), .B (w0[30] ), .Y (n_2868));
INVX2 g78036(.A (n_2865), .Y (n_3702));
INVX1 g78280(.A (n_2864), .Y (n_3778));
NAND2X1 g75577(.A (n_2522), .B (n_5643), .Y (n_3772));
INVX1 g77644(.A (n_4208), .Y (n_3626));
INVX1 g77458(.A (n_2861), .Y (n_2862));
NAND2X1 g73456(.A (n_2209), .B (n_28771), .Y (n_2856));
OR2X1 g74229(.A (n_1441), .B (n_379), .Y (n_3706));
INVX1 g77735(.A (n_2228), .Y (n_3768));
INVX1 g76877(.A (n_3535), .Y (n_3144));
INVX1 g78266(.A (n_2850), .Y (n_4405));
AND2X1 g65959(.A (n_2848), .B (u0_r0_rcnt[0] ), .Y (n_2849));
INVX1 g76546(.A (n_3091), .Y (n_4176));
NOR2X1 g65958(.A (n_2848), .B (ld), .Y (n_3972));
NAND2X2 g73708(.A (n_3491), .B (n_2462), .Y (n_3475));
XOR2X1 g76277(.A (text_in_r[112] ), .B (n_221), .Y (n_2846));
AND2X1 g77728(.A (n_1036), .B (n_28357), .Y (n_3076));
CLKBUFX1 g80779(.A (n_10315), .Y (n_12469));
INVX1 g77271(.A (n_2090), .Y (n_3060));
NOR2X1 g76563(.A (n_2241), .B (n_26493), .Y (n_6313));
NOR2X1 g74314(.A (n_251), .B (n_29409), .Y (n_3787));
OR2X1 g75741(.A (n_2109), .B (n_3920), .Y (n_3728));
NOR2X1 g73447(.A (n_2100), .B (n_6021), .Y (n_3679));
INVX2 g78590(.A (n_2838), .Y (n_15473));
INVX1 g80658(.A (n_2891), .Y (n_2837));
NOR2X1 g78108(.A (n_28459), .B (n_7559), .Y (n_2834));
INVX1 g77257(.A (n_2409), .Y (n_6422));
DFFX1 ld_r_reg(.CK (clk), .D (n_24548), .Q (ld_r), .QN ());
NAND2X2 g78002(.A (n_2830), .B (n_29269), .Y (n_11924));
INVX1 g77239(.A (n_2829), .Y (n_3119));
NOR2X1 g76960(.A (n_15986), .B (sa32[1] ), .Y (n_18121));
NOR2X1 g73670(.A (n_1223), .B (n_2943), .Y (n_2824));
INVX1 g76701(.A (n_3252), .Y (n_4318));
NOR2X1 g78243(.A (n_27904), .B (n_3756), .Y (n_4760));
INVX1 g74622(.A (n_2823), .Y (n_3312));
INVX1 g77625(.A (n_2820), .Y (n_2821));
NOR2X1 g77242(.A (n_28780), .B (n_28375), .Y (n_2819));
INVX1 g76529(.A (n_2818), .Y (n_3391));
INVX2 g78234(.A (n_1791), .Y (n_4416));
NOR2X1 g76699(.A (n_2084), .B (n_2810), .Y (n_2811));
NOR2X1 g73657(.A (n_1522), .B (n_28357), .Y (n_2809));
NOR2X1 g73652(.A (n_1246), .B (n_6462), .Y (n_3455));
INVX1 g76810(.A (n_2807), .Y (n_5143));
INVX2 g79070(.A (n_2805), .Y (n_15968));
INVX1 g75484(.A (n_2804), .Y (n_3273));
NOR2X1 g73595(.A (n_2206), .B (n_29167), .Y (n_2803));
INVX1 g77233(.A (n_27220), .Y (n_3500));
NAND3X1 g73646(.A (n_2211), .B (n_2744), .C (n_27222), .Y (n_3715));
NOR2X1 g74138(.A (n_2062), .B (n_3038), .Y (n_2796));
XOR2X1 g76113(.A (n_23352), .B (n_2769), .Y (n_2795));
NOR2X1 g73601(.A (n_1921), .B (n_3038), .Y (n_2794));
INVX2 g77311(.A (n_2792), .Y (n_4108));
INVX4 g80577(.A (n_2777), .Y (n_28271));
INVX1 g77225(.A (n_3802), .Y (n_4149));
INVX1 g77222(.A (n_2787), .Y (n_4207));
NAND2X2 g77221(.A (n_2218), .B (n_2235), .Y (n_3701));
CLKBUFX1 g77205(.A (n_3121), .Y (n_5985));
OR2X1 g77094(.A (n_5305), .B (n_7777), .Y (n_2785));
INVX1 g77523(.A (n_5370), .Y (n_3651));
INVX1 g76511(.A (n_2398), .Y (n_6439));
NAND2X1 g77080(.A (n_106), .B (n_826), .Y (n_3818));
NAND2X1 g73622(.A (n_2583), .B (n_6226), .Y (n_13239));
CLKBUFX2 g74719(.A (n_2781), .Y (n_4234));
NAND2X1 g76823(.A (n_27099), .B (n_656), .Y (n_7112));
INVX1 g78210(.A (n_3569), .Y (n_3694));
AND2X1 g74937(.A (n_2484), .B (n_2779), .Y (n_3032));
INVX1 g76509(.A (n_2774), .Y (n_2775));
INVX1 g77578(.A (n_2772), .Y (n_4422));
NAND2X1 g77545(.A (n_8918), .B (n_9335), .Y (n_2771));
XOR2X1 g76321(.A (n_23494), .B (n_2769), .Y (n_2770));
INVX1 g74214(.A (n_3365), .Y (n_2768));
NOR2X1 g76507(.A (n_2187), .B (n_9357), .Y (n_5104));
NOR2X1 g74194(.A (n_1480), .B (n_29158), .Y (n_3332));
NAND2X1 g76468(.A (n_624), .B (n_7496), .Y (n_3228));
NOR2X1 g77194(.A (n_14155), .B (sa23[1] ), .Y (n_20269));
INVX1 g77899(.A (n_1488), .Y (n_3030));
INVX1 g76495(.A (n_2755), .Y (n_3671));
INVX1 g75062(.A (n_2160), .Y (n_4612));
NAND2X2 g77197(.A (n_1887), .B (n_2943), .Y (n_3666));
INVX1 g77779(.A (n_2753), .Y (n_2754));
INVX1 g77323(.A (n_2901), .Y (n_2752));
NAND2X1 g73901(.A (n_2094), .B (n_3807), .Y (n_2751));
INVX1 g77653(.A (n_2749), .Y (n_2750));
INVX1 g78203(.A (n_2748), .Y (n_4302));
NAND2X1 g74824(.A (n_2621), .B (n_2150), .Y (n_3672));
INVX1 g76897(.A (n_2873), .Y (n_5887));
NAND2X1 g73568(.A (n_2530), .B (n_827), .Y (n_3444));
XOR2X1 g76230(.A (text_in_r[110] ), .B (n_23599), .Y (n_2745));
INVX1 g79507(.A (n_2744), .Y (n_4042));
INVX1 g78047(.A (n_2743), .Y (n_3071));
NOR2X1 g73518(.A (n_2742), .B (n_3307), .Y (n_3437));
INVX1 g74611(.A (n_1929), .Y (n_3306));
NAND2X1 g73614(.A (n_2738), .B (n_27674), .Y (n_2739));
INVX1 g76781(.A (n_13875), .Y (n_3003));
INVX1 g77157(.A (n_3002), .Y (n_3917));
INVX1 g76980(.A (n_3816), .Y (n_3135));
CLKBUFX1 g77678(.A (n_3448), .Y (n_4414));
NAND2X1 g74709(.A (n_3338), .B (n_2534), .Y (n_2733));
XOR2X1 g76134(.A (text_in_r[124] ), .B (w0[28] ), .Y (n_2732));
NOR2X1 g77329(.A (n_3920), .B (n_1616), .Y (n_4233));
NOR2X1 g75052(.A (n_1771), .B (n_1711), .Y (n_3726));
NAND2X1 g74172(.A (n_1835), .B (n_7182), .Y (n_3334));
NOR2X1 g74693(.A (n_1371), .B (n_27124), .Y (n_3604));
NAND2X2 g77153(.A (n_1745), .B (n_6185), .Y (n_9708));
NOR2X1 g73620(.A (n_1685), .B (n_28480), .Y (n_3691));
INVX1 g79601(.A (n_19385), .Y (n_20477));
CLKBUFX3 g77211(.A (n_2723), .Y (n_4635));
INVX1 g76456(.A (n_27673), .Y (n_3388));
NOR2X1 g76985(.A (n_28642), .B (n_844), .Y (n_19752));
INVX1 g78030(.A (n_3281), .Y (n_9351));
INVX1 g78092(.A (n_2719), .Y (n_4154));
NAND2X2 g76909(.A (n_27133), .B (n_28419), .Y (n_3471));
INVX1 g76584(.A (n_2526), .Y (n_10199));
INVX1 g81498(.A (n_17411), .Y (n_3910));
INVX1 g77894(.A (n_2718), .Y (n_21598));
NAND2X1 g74362(.A (n_1837), .B (n_2492), .Y (n_4552));
INVX2 g77059(.A (n_1570), .Y (n_6442));
NAND2X1 g77967(.A (n_1601), .B (n_218), .Y (n_3235));
INVX1 g78023(.A (n_3491), .Y (n_3052));
NOR2X1 g73626(.A (n_1918), .B (n_10315), .Y (n_3350));
NAND2X1 g74545(.A (n_2716), .B (n_379), .Y (n_3316));
INVX1 g77903(.A (n_2715), .Y (n_4849));
INVX1 g77351(.A (n_2925), .Y (n_3849));
INVX1 g78220(.A (n_2714), .Y (n_3700));
INVX1 g77620(.A (n_1548), .Y (n_3987));
INVX1 g77187(.A (n_2713), .Y (n_3710));
INVX1 g77847(.A (n_2710), .Y (n_2711));
NOR2X1 g77546(.A (n_10100), .B (n_2180), .Y (n_2709));
NOR2X1 g76515(.A (n_636), .B (n_2708), .Y (n_3175));
INVX1 g78062(.A (n_2707), .Y (n_4117));
INVX1 g77786(.A (n_3303), .Y (n_2706));
INVX1 g77689(.A (n_3319), .Y (n_2705));
INVX1 g77141(.A (n_26889), .Y (n_2704));
INVX1 g77800(.A (n_2702), .Y (n_19795));
INVX8 g80997(.A (n_1310), .Y (n_19364));
INVX2 g75540(.A (n_1594), .Y (n_3269));
XOR2X1 g76257(.A (text_in_r[70] ), .B (n_141), .Y (n_2700));
OR2X1 g74121(.A (n_1983), .B (n_7537), .Y (n_3551));
NOR2X1 g74421(.A (n_2113), .B (n_4586), .Y (n_3893));
NAND3X1 g73634(.A (n_28793), .B (n_1989), .C (n_627), .Y (n_2699));
INVX1 g77072(.A (n_3813), .Y (n_4169));
NAND2X1 g78224(.A (n_27904), .B (n_4173), .Y (n_4159));
INVX1 g77494(.A (n_16579), .Y (n_19830));
INVX1 g77708(.A (n_3422), .Y (n_3079));
INVX1 g77217(.A (n_4676), .Y (n_3502));
INVX1 g76626(.A (n_2696), .Y (n_3161));
INVX1 g77672(.A (n_2695), .Y (n_3673));
INVX1 g78176(.A (n_7418), .Y (n_6406));
INVX1 g78192(.A (n_1821), .Y (n_2694));
XOR2X1 g76205(.A (n_2692), .B (n_112), .Y (n_2693));
AND2X1 g76620(.A (n_6997), .B (n_2119), .Y (n_3963));
NAND2X2 g74353(.A (n_1243), .B (n_26601), .Y (n_4643));
OR2X1 g77612(.A (n_2830), .B (n_29244), .Y (n_3085));
NAND2X1 g74333(.A (n_2691), .B (n_27593), .Y (n_3812));
INVX2 g76915(.A (n_2374), .Y (n_4144));
INVX1 g76517(.A (n_2687), .Y (n_10127));
NOR2X1 g73437(.A (n_1817), .B (n_5413), .Y (n_3911));
INVX1 g77614(.A (n_2684), .Y (n_3084));
XOR2X1 g76175(.A (text_in_r[107] ), .B (n_23363), .Y (n_2683));
INVX1 g78155(.A (n_2682), .Y (n_20388));
INVX1 g81243(.A (n_20862), .Y (n_21520));
INVX2 g76675(.A (n_2680), .Y (n_3594));
INVX1 g73421(.A (n_1775), .Y (n_3353));
NAND2X1 g75074(.A (n_2049), .B (n_3038), .Y (n_4500));
INVX1 g78070(.A (n_2678), .Y (n_3473));
XOR2X1 g76196(.A (text_in_r[102] ), .B (n_243), .Y (n_2676));
XOR2X1 g76207(.A (n_221), .B (n_250), .Y (n_2672));
INVX1 g73402(.A (n_2664), .Y (n_2665));
INVX1 g78104(.A (n_2663), .Y (n_19852));
NOR2X1 g75150(.A (n_818), .B (n_1534), .Y (n_2662));
XOR2X1 g76332(.A (text_in_r[81] ), .B (n_22591), .Y (n_2660));
NOR2X1 g73916(.A (n_2671), .B (n_1711), .Y (n_2658));
INVX1 g82295(.A (n_27493), .Y (n_17089));
NOR2X1 g73937(.A (n_1772), .B (n_2656), .Y (n_3342));
NOR2X1 g73348(.A (n_1707), .B (n_2655), .Y (n_3457));
INVX1 g77302(.A (n_2654), .Y (n_3791));
NAND2X2 g77115(.A (n_28566), .B (n_28466), .Y (n_3698));
XOR2X1 g76164(.A (n_221), .B (n_2648), .Y (n_2650));
INVX1 g77200(.A (n_3585), .Y (n_3687));
INVX1 g77535(.A (n_5735), .Y (n_19114));
NAND2X1 g77928(.A (n_26880), .B (n_1551), .Y (n_3513));
INVX1 g77162(.A (n_3536), .Y (n_2647));
NOR2X1 g73508(.A (n_2162), .B (n_2646), .Y (n_3610));
INVX1 g76737(.A (n_3427), .Y (n_2645));
NAND2X2 g76671(.A (n_2085), .B (n_1540), .Y (n_3890));
INVX1 g77091(.A (n_2640), .Y (n_2641));
XOR2X1 g76161(.A (n_22557), .B (n_1072), .Y (n_2639));
NAND2X1 g76443(.A (n_1756), .B (n_28423), .Y (n_3467));
INVX1 g77124(.A (n_2638), .Y (n_4299));
INVX1 g77931(.A (n_2635), .Y (n_2636));
XOR2X1 g76122(.A (n_234), .B (n_194), .Y (n_2633));
NOR2X1 g73887(.A (n_2048), .B (n_2467), .Y (n_2632));
INVX1 g77664(.A (n_2628), .Y (n_3723));
INVX1 g76523(.A (n_2627), .Y (n_4146));
AND2X1 g77030(.A (n_19364), .B (sa01[1] ), .Y (n_17459));
INVX1 g77701(.A (n_3346), .Y (n_3717));
NOR2X1 g76995(.A (n_2231), .B (n_9118), .Y (n_2625));
NOR2X1 g73797(.A (n_26395), .B (n_1789), .Y (n_3865));
NOR2X1 g73357(.A (n_2092), .B (n_28464), .Y (n_2623));
NAND2X1 g76963(.A (n_26276), .B (n_902), .Y (n_7213));
NAND2X1 g73751(.A (n_2621), .B (n_3067), .Y (n_3825));
OR2X1 g73732(.A (n_2214), .B (n_379), .Y (n_4638));
OR2X1 g73352(.A (n_1246), .B (n_27434), .Y (n_13166));
INVX1 g76927(.A (n_2617), .Y (n_9170));
XOR2X1 g76289(.A (text_in_r[108] ), .B (n_23290), .Y (n_2616));
NAND2X2 g76818(.A (n_2483), .B (n_1484), .Y (n_4022));
INVX1 g78130(.A (n_2613), .Y (n_4965));
INVX1 g76869(.A (n_3373), .Y (n_4245));
INVX1 g76754(.A (n_3297), .Y (n_3461));
NOR2X1 g76902(.A (n_2337), .B (n_1942), .Y (n_2612));
INVX1 g77599(.A (n_2611), .Y (n_4920));
INVX1 g77705(.A (n_2608), .Y (n_2609));
INVX1 g77822(.A (n_8227), .Y (n_2606));
INVX1 g76874(.A (n_2604), .Y (n_2605));
NOR2X1 g76847(.A (n_27641), .B (n_28410), .Y (n_2603));
AND2X1 g77400(.A (n_17260), .B (n_1196), .Y (n_16097));
INVX1 g76829(.A (n_3420), .Y (n_2598));
OR2X1 g73615(.A (n_1822), .B (n_3920), .Y (n_4639));
INVX1 g76805(.A (n_2596), .Y (n_6833));
INVX1 g77108(.A (n_2049), .Y (n_4501));
NAND2X1 g74916(.A (n_29121), .B (n_636), .Y (n_2595));
INVX1 g77630(.A (n_2594), .Y (n_3915));
INVX1 g80091(.A (n_2592), .Y (n_3445));
XOR2X1 g76217(.A (text_in_r[119] ), .B (n_22717), .Y (n_2591));
XOR2X1 g76150(.A (text_in_r[121] ), .B (n_22569), .Y (n_2590));
NAND2X1 g73539(.A (n_2621), .B (n_330), .Y (n_12870));
XOR2X1 g76213(.A (text_in_r[94] ), .B (n_2587), .Y (n_2588));
INVX1 g77203(.A (n_3121), .Y (n_2586));
CLKBUFX1 g76740(.A (n_3427), .Y (n_4115));
XOR2X1 g76248(.A (text_in_r[120] ), .B (n_1318), .Y (n_2585));
NAND2X2 g73533(.A (n_2583), .B (n_4611), .Y (n_5645));
NAND2X2 g76695(.A (n_28754), .B (n_6790), .Y (n_15800));
NAND2X1 g73501(.A (n_2541), .B (n_3920), .Y (n_13681));
INVX1 g75466(.A (n_2580), .Y (n_3852));
NOR2X1 g76639(.A (n_13804), .B (sa10[1] ), .Y (n_18087));
NOR2X1 g76640(.A (n_2007), .B (n_8263), .Y (n_2577));
INVX1 g76765(.A (n_1744), .Y (n_3443));
INVX1 g76941(.A (n_2575), .Y (n_7101));
INVX1 g76587(.A (n_3096), .Y (n_5167));
NOR2X1 g73413(.A (n_2040), .B (n_1273), .Y (n_2574));
OR2X1 g76572(.A (n_1641), .B (n_3318), .Y (n_2573));
INVX4 g80943(.A (n_14624), .Y (n_18456));
INVX1 g81657(.A (n_28134), .Y (n_2570));
INVX1 g77828(.A (n_2568), .Y (n_2569));
NOR2X1 g74548(.A (n_1998), .B (n_4925), .Y (n_3174));
NOR2X1 g73323(.A (n_27204), .B (n_1905), .Y (n_3294));
NOR2X1 g77472(.A (n_13804), .B (n_177), .Y (n_3168));
NAND2X2 g76452(.A (n_868), .B (n_719), .Y (n_4595));
INVX1 g77042(.A (n_2496), .Y (n_2565));
CLKBUFX3 g74154(.A (n_2563), .Y (n_4401));
NAND2X2 g76843(.A (n_2254), .B (n_2656), .Y (n_3148));
NAND2X1 g76778(.A (n_997), .B (n_1431), .Y (n_3153));
INVX1 g77590(.A (n_3900), .Y (n_11648));
NOR2X1 g73775(.A (n_3284), .B (n_2025), .Y (n_3842));
XOR2X1 g76337(.A (n_2560), .B (n_97), .Y (n_2561));
XOR2X1 g76210(.A (n_23551), .B (n_1308), .Y (n_2559));
XOR2X1 g76316(.A (text_in_r[99] ), .B (w0[3] ), .Y (n_2556));
INVX2 g78119(.A (n_11739), .Y (n_3386));
XOR2X1 g76306(.A (text_in_r[84] ), .B (w1[20] ), .Y (n_2555));
XOR2X1 g76348(.A (text_in_r[78] ), .B (w1[14] ), .Y (n_2552));
XOR2X1 g76288(.A (text_in_r[122] ), .B (w0[26] ), .Y (n_2550));
NOR2X1 g75730(.A (n_1911), .B (n_3807), .Y (n_4547));
XOR2X1 g76265(.A (text_in_r[118] ), .B (n_23255), .Y (n_2547));
INVX1 g77711(.A (n_8540), .Y (n_17813));
XOR2X1 g76145(.A (text_in_r[73] ), .B (n_22496), .Y (n_2544));
XOR2X1 g76239(.A (text_in_r[56] ), .B (n_1220), .Y (n_2543));
INVX1 g77056(.A (n_3573), .Y (n_3965));
NAND2X1 g73318(.A (n_2541), .B (n_3038), .Y (n_3692));
XOR2X1 g76231(.A (n_2692), .B (n_21708), .Y (n_2540));
OR2X1 g77575(.A (n_2359), .B (n_1147), .Y (n_2537));
INVX1 g77118(.A (n_2536), .Y (n_3230));
NAND2X2 g75138(.A (n_2534), .B (n_2235), .Y (n_4504));
NAND2X1 g75691(.A (n_27224), .B (n_28340), .Y (n_3253));
INVX1 g77998(.A (n_2459), .Y (n_4450));
XOR2X1 g76209(.A (text_in_r[37] ), .B (n_194), .Y (n_2532));
NAND2X1 g73500(.A (n_2530), .B (n_379), .Y (n_11626));
NAND2X1 g75473(.A (n_2502), .B (n_4568), .Y (n_3861));
INVX1 g76585(.A (n_2526), .Y (n_2527));
XOR2X1 g76194(.A (text_in_r[66] ), .B (n_245), .Y (n_2524));
NAND2X1 g74255(.A (n_2522), .B (n_27222), .Y (n_4513));
NOR2X1 g78181(.A (n_16204), .B (n_9084), .Y (n_2521));
INVX1 g78122(.A (n_1671), .Y (n_2519));
INVX1 g81104(.A (n_27407), .Y (n_19395));
XOR2X1 g76169(.A (text_in_r[116] ), .B (n_22653), .Y (n_2516));
INVX1 g77970(.A (n_2514), .Y (n_2515));
INVX2 g77100(.A (n_2513), .Y (n_10147));
XOR2X1 g76162(.A (n_1934), .B (n_1040), .Y (n_2511));
NAND2X2 g76762(.A (n_1037), .B (n_27204), .Y (n_2510));
CLKBUFX1 g81726(.A (n_27202), .Y (n_7947));
XOR2X1 g76152(.A (n_1318), .B (n_23261), .Y (n_2509));
INVX1 g78133(.A (n_8139), .Y (n_17706));
XOR2X1 g76137(.A (text_in_r[76] ), .B (w1[12] ), .Y (n_2505));
AND2X1 g74742(.A (n_2502), .B (n_27434), .Y (n_2503));
CLKBUFX1 g77045(.A (n_2496), .Y (n_4388));
XOR2X1 g76154(.A (text_in_r[115] ), .B (n_24266), .Y (n_2494));
NAND2X1 g73387(.A (n_2583), .B (n_2492), .Y (n_3499));
AND2X1 g77084(.A (n_19791), .B (n_2204), .Y (n_17703));
INVX1 g78179(.A (n_2488), .Y (n_6696));
NOR2X1 g73559(.A (n_2076), .B (n_4721), .Y (n_3656));
NOR2X1 g73679(.A (n_2078), .B (n_2487), .Y (n_3463));
AND2X1 g73917(.A (n_1402), .B (n_490), .Y (n_14734));
INVX1 g77568(.A (n_4382), .Y (n_2485));
NAND2X2 g75666(.A (n_2484), .B (n_2467), .Y (n_4565));
OR2X1 g74019(.A (n_1782), .B (n_2483), .Y (n_3589));
NOR2X1 g73513(.A (n_2017), .B (n_3840), .Y (n_2481));
INVX1 g74326(.A (n_2892), .Y (n_2479));
NAND2X1 g77018(.A (n_13083), .B (n_583), .Y (n_3093));
INVX1 g77138(.A (n_1883), .Y (n_3938));
NAND2X1 g74571(.A (n_2484), .B (n_490), .Y (n_3237));
INVX1 g77377(.A (n_3465), .Y (n_3924));
NAND2X2 g74999(.A (n_29121), .B (n_2343), .Y (n_4525));
INVX1 g78245(.A (n_13575), .Y (n_2470));
INVX1 g77278(.A (n_2469), .Y (n_5138));
NOR2X1 g74000(.A (n_1897), .B (n_2467), .Y (n_2468));
INVX1 g78115(.A (n_2466), .Y (n_3047));
NAND2X1 g75381(.A (n_1516), .B (n_1539), .Y (n_4604));
INVX2 g75387(.A (n_2464), .Y (n_3250));
NOR2X1 g75040(.A (n_2253), .B (n_2462), .Y (n_3270));
INVX1 g78148(.A (n_2461), .Y (n_4168));
INVX1 g78688(.A (n_2981), .Y (n_18440));
INVX1 g77999(.A (n_2459), .Y (n_2460));
INVX1 g75845(.A (n_1781), .Y (n_3372));
NOR2X1 g73690(.A (n_2183), .B (n_386), .Y (n_3469));
NAND2X1 g74573(.A (n_2456), .B (n_3081), .Y (n_2457));
NOR2X1 g77039(.A (n_1484), .B (n_367), .Y (n_3130));
XOR2X1 g76131(.A (text_in_r[95] ), .B (n_338), .Y (n_2455));
NAND2X1 g75416(.A (n_962), .B (n_1711), .Y (n_4533));
OR2X1 g75368(.A (n_9999), .B (n_14627), .Y (n_2452));
XOR2X1 g76310(.A (n_234), .B (w1[5] ), .Y (n_2450));
INVX1 g78250(.A (n_2447), .Y (n_3755));
INVX1 g76432(.A (n_2446), .Y (n_4104));
INVX8 g78786(.A (n_26386), .Y (n_9500));
OR2X1 g75663(.A (n_2444), .B (n_7658), .Y (n_9295));
INVX1 g76643(.A (n_3746), .Y (n_3240));
XOR2X1 g76101(.A (text_in_r[86] ), .B (n_2440), .Y (n_2441));
XOR2X1 g76119(.A (n_243), .B (n_2437), .Y (n_2438));
XOR2X1 g76130(.A (text_in_r[74] ), .B (w1[10] ), .Y (n_2436));
XOR2X1 g76136(.A (n_2434), .B (n_245), .Y (n_2435));
XOR2X1 g76141(.A (text_in_r[101] ), .B (n_234), .Y (n_2433));
XOR2X1 g76174(.A (text_in_r[123] ), .B (n_2430), .Y (n_2431));
XOR2X1 g76177(.A (text_in_r[39] ), .B (w2[7] ), .Y (n_2429));
NAND2X1 g75354(.A (n_2111), .B (n_5005), .Y (n_2426));
XOR2X1 g76206(.A (n_1970), .B (n_22496), .Y (n_2425));
XOR2X1 g76211(.A (text_in_r[100] ), .B (n_22881), .Y (n_2423));
XOR2X1 g76222(.A (n_243), .B (n_141), .Y (n_2422));
XOR2X1 g76225(.A (text_in_r[67] ), .B (w1[3] ), .Y (n_2420));
XOR2X1 g76227(.A (text_in_r[83] ), .B (n_2417), .Y (n_2418));
XOR2X1 g76238(.A (text_in_r[88] ), .B (n_23261), .Y (n_2416));
XOR2X1 g76241(.A (text_in_r[98] ), .B (w0[2] ), .Y (n_2415));
XOR2X1 g76246(.A (text_in_r[90] ), .B (n_2412), .Y (n_2413));
XOR2X1 g76267(.A (text_in_r[111] ), .B (n_23580), .Y (n_2408));
NAND2X1 g75377(.A (n_1102), .B (n_2943), .Y (n_3241));
XOR2X1 g76315(.A (n_22567), .B (n_22591), .Y (n_2406));
XOR2X1 g76329(.A (n_23763), .B (n_23397), .Y (n_2405));
INVX1 g77266(.A (n_2404), .Y (n_9959));
XOR2X1 g76336(.A (text_in_r[77] ), .B (n_23096), .Y (n_2403));
INVX1 g77474(.A (n_2402), .Y (n_3425));
INVX1 g76512(.A (n_2398), .Y (n_2399));
INVX1 g76535(.A (n_4093), .Y (n_3364));
INVX2 g74653(.A (n_2071), .Y (n_4590));
INVX1 g76549(.A (n_2396), .Y (n_2397));
INVX1 g76616(.A (n_2392), .Y (n_2393));
INVX1 g76622(.A (n_2307), .Y (n_14107));
NAND2X2 g76636(.A (n_1229), .B (n_26893), .Y (n_3218));
NOR2X1 g76638(.A (n_719), .B (n_27434), .Y (n_3225));
NOR2X1 g64202(.A (n_6301), .B (n_986), .Y (n_2390));
INVX1 g76664(.A (n_3247), .Y (n_3157));
NOR2X1 g76689(.A (n_932), .B (n_8452), .Y (n_13037));
INVX2 g76709(.A (n_2387), .Y (n_3830));
INVX1 g76729(.A (n_2385), .Y (n_2386));
AND2X1 g76749(.A (n_18266), .B (sa00[1] ), .Y (n_19170));
NAND2X1 g76772(.A (n_399), .B (n_17912), .Y (n_3630));
INVX1 g76773(.A (n_10191), .Y (n_2384));
NOR2X1 g76776(.A (n_2152), .B (n_2383), .Y (n_4266));
INVX1 g76799(.A (n_1988), .Y (n_3749));
NOR2X1 g76820(.A (n_3560), .B (n_7598), .Y (n_2380));
INVX1 g76828(.A (n_3420), .Y (n_5404));
NAND2X1 g76834(.A (n_795), .B (n_27757), .Y (n_3711));
NAND2X2 g76852(.A (n_1850), .B (n_28787), .Y (n_5368));
INVX1 g76918(.A (n_2372), .Y (n_2373));
NOR2X1 g76944(.A (n_2368), .B (n_8997), .Y (n_2369));
INVX1 g76952(.A (n_2366), .Y (n_2367));
INVX2 g76973(.A (n_27598), .Y (n_4520));
INVX1 g76983(.A (n_2365), .Y (n_3134));
INVX2 g76986(.A (n_2364), .Y (n_16895));
INVX1 g77000(.A (n_2362), .Y (n_2363));
INVX2 g77014(.A (n_1552), .Y (n_3204));
INVX1 g77019(.A (n_1695), .Y (n_11669));
INVX1 g77021(.A (n_2360), .Y (n_29130));
INVX1 g77856(.A (n_8706), .Y (n_16052));
NAND2X1 g77029(.A (n_2359), .B (n_27198), .Y (n_3195));
OR2X1 g77061(.A (n_8093), .B (n_28362), .Y (n_2356));
NAND2X1 g77067(.A (n_28133), .B (n_4391), .Y (n_3522));
INVX1 g77081(.A (n_2353), .Y (n_12222));
INVX1 g77929(.A (n_2351), .Y (n_2352));
INVX1 g77464(.A (n_2643), .Y (n_2350));
INVX1 g77106(.A (n_1825), .Y (n_6198));
INVX1 g77126(.A (n_2349), .Y (n_4331));
NAND2X1 g77387(.A (n_27985), .B (n_29167), .Y (n_3923));
INVX1 g77168(.A (n_2931), .Y (n_12836));
INVX2 g77190(.A (n_2766), .Y (n_6836));
CLKBUFX1 g77398(.A (n_2346), .Y (n_4012));
INVX1 g77230(.A (n_2344), .Y (n_2345));
NAND2X1 g77246(.A (n_736), .B (n_2343), .Y (n_3729));
NAND2X1 g77285(.A (n_16480), .B (n_2063), .Y (n_3760));
INVX1 g80988(.A (n_1310), .Y (n_16279));
NAND2X1 g77003(.A (n_2337), .B (n_2383), .Y (n_4014));
INVX1 g77440(.A (n_2336), .Y (n_4227));
INVX1 g77482(.A (n_1748), .Y (n_3209));
INVX1 g74514(.A (n_2335), .Y (n_7329));
INVX1 g77530(.A (n_2334), .Y (n_4228));
INVX1 g77558(.A (n_2332), .Y (n_2333));
INVX1 g77560(.A (n_2330), .Y (n_2331));
INVX1 g77597(.A (n_2611), .Y (n_2329));
NAND2X1 g76867(.A (n_6877), .B (n_897), .Y (n_2327));
NAND2X2 g77448(.A (n_28547), .B (n_28464), .Y (n_3087));
AND2X1 g77693(.A (n_4568), .B (n_9368), .Y (n_5516));
INVX1 g77712(.A (n_8540), .Y (n_12624));
INVX1 g77722(.A (n_2168), .Y (n_4426));
INVX1 g77746(.A (n_2322), .Y (n_6234));
INVX1 g77915(.A (n_27072), .Y (n_3562));
OR2X1 g77766(.A (n_2319), .B (n_2318), .Y (n_2320));
NOR2X1 g76474(.A (n_16434), .B (sa00[1] ), .Y (n_20760));
INVX1 g77869(.A (n_1599), .Y (n_4105));
INVX4 g81170(.A (n_399), .Y (n_12559));
INVX1 g77879(.A (n_2311), .Y (n_4188));
INVX1 g76990(.A (n_3267), .Y (n_4699));
NOR2X1 g77959(.A (n_7734), .B (n_10452), .Y (n_2306));
INVX1 g77565(.A (n_5691), .Y (n_12335));
INVX1 g77427(.A (n_2305), .Y (n_3041));
INVX1 g77981(.A (n_2304), .Y (n_4200));
INVX1 g78009(.A (n_2303), .Y (n_4404));
INVX1 g78013(.A (n_2301), .Y (n_2302));
INVX1 g78097(.A (n_2298), .Y (n_3049));
XOR2X1 g76281(.A (w0[0] ), .B (n_22418), .Y (n_2297));
NOR2X1 g74498(.A (n_1620), .B (n_4611), .Y (n_4786));
INVX1 g77910(.A (n_2295), .Y (n_9965));
INVX2 g77432(.A (n_1494), .Y (n_4581));
INVX1 g78157(.A (n_2292), .Y (n_12494));
NOR2X1 g73910(.A (n_2235), .B (n_29316), .Y (n_3345));
INVX2 g75614(.A (n_1741), .Y (n_4705));
INVX1 g78086(.A (n_13423), .Y (n_2290));
NAND2X1 g76615(.A (n_1576), .B (n_6185), .Y (n_2289));
INVX1 g76610(.A (n_2286), .Y (n_3653));
NOR2X1 g73904(.A (n_1503), .B (n_3820), .Y (n_3040));
NOR2X1 g76650(.A (n_1621), .B (n_2646), .Y (n_3159));
NAND2X1 g77421(.A (n_6021), .B (n_28375), .Y (n_4832));
NAND2X1 g78152(.A (n_4846), .B (n_9357), .Y (n_4974));
AND2X1 g73892(.A (n_1839), .B (n_4611), .Y (n_13738));
INVX1 g79867(.A (n_844), .Y (n_21569));
INVX1 g78238(.A (n_2278), .Y (n_2279));
NAND2X1 g76473(.A (n_14624), .B (n_481), .Y (n_7789));
INVX2 g77417(.A (n_2042), .Y (n_4514));
INVX8 g79074(.A (n_205), .Y (n_9118));
INVX1 g80397(.A (n_7725), .Y (n_4082));
NOR2X1 g76604(.A (n_4916), .B (n_3868), .Y (n_4106));
INVX1 g80342(.A (n_7410), .Y (n_3943));
INVX4 g80761(.A (n_441), .Y (n_9442));
INVX1 g75558(.A (n_2267), .Y (n_3869));
INVX1 g76601(.A (n_2266), .Y (n_4334));
INVX1 g77389(.A (n_2265), .Y (n_4210));
NAND2X1 g73872(.A (n_2933), .B (n_27204), .Y (n_3385));
INVX1 g78470(.A (n_1053), .Y (n_11276));
OR2X1 g74924(.A (n_1996), .B (n_490), .Y (n_3682));
INVX1 g77883(.A (n_1461), .Y (n_4055));
INVX1 g76951(.A (n_2366), .Y (n_3138));
NOR2X1 g76654(.A (n_27688), .B (sa01[1] ), .Y (n_20765));
NAND2X1 g77289(.A (n_494), .B (n_2260), .Y (n_2994));
INVX1 g77402(.A (n_2259), .Y (n_8342));
INVX1 g77163(.A (n_2253), .Y (n_3536));
INVX1 g80246(.A (n_2251), .Y (n_3667));
INVX2 g80376(.A (n_2368), .Y (n_9089));
MX2X1 g76042(.A (text_in_r[5] ), .B (text_in[5]), .S0 (n_24778), .Y(n_2247));
AND2X1 g77588(.A (n_3704), .B (n_27365), .Y (n_2914));
MX2X1 g76004(.A (text_in_r[50] ), .B (text_in[50]), .S0 (n_25123),.Y (n_2244));
NOR2X1 g77399(.A (n_27674), .B (n_926), .Y (n_2346));
NOR2X1 g77892(.A (n_9819), .B (n_276), .Y (n_9978));
NAND2X1 g77646(.A (n_27688), .B (n_8452), .Y (n_4208));
NAND2X1 g76730(.A (n_9527), .B (w3[25] ), .Y (n_2385));
INVX1 g76478(.A (n_1282), .Y (n_2958));
INVX1 g79769(.A (n_2241), .Y (n_7601));
INVX1 g80659(.A (n_2237), .Y (n_2891));
AND2X1 g77451(.A (n_27133), .B (n_28375), .Y (n_7023));
NAND2X2 g78149(.A (n_2236), .B (n_2235), .Y (n_2461));
XOR2X1 g76305(.A (text_in_r[47] ), .B (w2[15] ), .Y (n_2234));
XOR2X1 g76095(.A (n_16938), .B (n_1236), .Y (n_2229));
NAND2X1 g77736(.A (n_630), .B (n_1285), .Y (n_2228));
XOR2X1 g76102(.A (text_in_r[52] ), .B (w2[20] ), .Y (n_2227));
NOR2X1 g77656(.A (n_8918), .B (n_3840), .Y (n_2749));
XOR2X1 g76325(.A (text_in_r[35] ), .B (w2[3] ), .Y (n_2220));
INVX1 g82488(.A (n_2218), .Y (n_2674));
INVX8 g81052(.A (n_1756), .Y (n_11400));
MX2X1 g76014(.A (text_in_r[2] ), .B (text_in[2]), .S0 (n_619), .Y(n_2217));
INVX1 g76933(.A (n_2456), .Y (n_2216));
INVX1 g76710(.A (n_1002), .Y (n_2387));
INVX1 g77372(.A (n_2214), .Y (n_5271));
NAND2X2 g76583(.A (n_2158), .B (n_28357), .Y (n_2213));
MX2X1 g76052(.A (text_in_r[31] ), .B (text_in[31]), .S0 (ld), .Y(n_2212));
NAND2X1 g77579(.A (n_2211), .B (n_2343), .Y (n_2772));
INVX1 g77423(.A (n_2209), .Y (n_2210));
INVX1 g77465(.A (n_2206), .Y (n_2643));
CLKBUFX1 g77226(.A (n_2522), .Y (n_3802));
XOR2X1 g76178(.A (n_23547), .B (n_23079), .Y (n_2201));
XOR2X1 g76155(.A (text_in_r[113] ), .B (n_22567), .Y (n_2198));
NAND2X1 g77167(.A (n_1014), .B (n_2239), .Y (n_2991));
INVX1 g80093(.A (n_2191), .Y (n_2592));
INVX1 g78907(.A (n_2187), .Y (n_7362));
INVX1 g77823(.A (n_13872), .Y (n_8227));
NAND2X1 g77358(.A (n_19310), .B (n_7658), .Y (n_2952));
XOR2X1 g76294(.A (text_in_r[80] ), .B (w1[16] ), .Y (n_2185));
NAND2X1 g76923(.A (n_849), .B (n_28469), .Y (n_2937));
INVX1 g77501(.A (n_7649), .Y (n_7614));
INVX1 g77636(.A (n_2183), .Y (n_3615));
INVX1 g79649(.A (n_2180), .Y (n_2181));
AND2X1 g77812(.A (n_4916), .B (n_437), .Y (n_3945));
INVX1 g79715(.A (n_290), .Y (n_18168));
NAND2X1 g75485(.A (n_1384), .B (n_27204), .Y (n_2804));
MX2X1 g76048(.A (text_in_r[27] ), .B (text_in[27]), .S0 (n_24599),.Y (n_2176));
XOR2X1 g76330(.A (n_2174), .B (n_9203), .Y (n_2175));
XOR2X1 g76204(.A (text_in_r[50] ), .B (w2[18] ), .Y (n_2173));
NAND2X1 g75467(.A (n_1155), .B (n_1079), .Y (n_2580));
INVX4 g81331(.A (n_20406), .Y (n_14142));
INVX8 g81131(.A (n_2001), .Y (n_15039));
NOR2X1 g76550(.A (n_1628), .B (n_2318), .Y (n_2396));
INVX1 g76789(.A (n_1746), .Y (n_2170));
INVX1 g78188(.A (n_27225), .Y (n_7196));
NOR2X1 g77723(.A (n_1118), .B (n_2483), .Y (n_2168));
INVX1 g76913(.A (n_1177), .Y (n_2929));
INVX8 g81967(.A (n_27901), .Y (n_11322));
OR2X1 g77793(.A (n_13815), .B (n_171), .Y (n_2917));
INVX1 g77982(.A (n_2162), .Y (n_2304));
INVX1 g78167(.A (n_6889), .Y (n_2895));
INVX1 g82390(.A (n_27336), .Y (n_15688));
INVX1 g77787(.A (n_2530), .Y (n_3303));
NOR2X1 g75063(.A (n_1430), .B (n_100), .Y (n_2160));
NAND2X1 g78000(.A (n_541), .B (n_1427), .Y (n_2459));
INVX1 g79256(.A (n_1196), .Y (n_16362));
NOR2X1 g76627(.A (n_2158), .B (n_28357), .Y (n_2696));
NOR2X1 g78308(.A (n_3704), .B (n_27365), .Y (n_2916));
INVX1 g80808(.A (n_2152), .Y (n_2153));
NAND2X1 g76487(.A (n_1266), .B (n_2150), .Y (n_2151));
INVX1 g79241(.A (n_3081), .Y (n_2905));
NOR2X1 g77801(.A (n_15674), .B (n_3264), .Y (n_2702));
AND2X1 g77780(.A (n_1336), .B (n_29158), .Y (n_2753));
XOR2X1 g76180(.A (text_in_r[63] ), .B (w2[31] ), .Y (n_2148));
INVX1 g77773(.A (n_2145), .Y (n_2146));
NAND2X1 g76988(.A (n_27688), .B (n_1010), .Y (n_2364));
NAND2X1 g77591(.A (n_4300), .B (n_27746), .Y (n_3900));
INVX1 g79485(.A (n_2254), .Y (n_2140));
INVX1 g77769(.A (n_2137), .Y (n_5546));
XOR2X1 g76208(.A (n_23001), .B (n_23087), .Y (n_2135));
NAND2X1 g77857(.A (n_27098), .B (n_26491), .Y (n_8706));
NOR2X1 g77524(.A (n_28357), .B (n_2044), .Y (n_5370));
CLKBUFX3 g77763(.A (n_2691), .Y (n_3187));
XOR2X1 g76319(.A (n_1674), .B (n_22829), .Y (n_2131));
NOR2X1 g77759(.A (n_28781), .B (n_28445), .Y (n_2128));
INVX4 g81956(.A (n_2022), .Y (n_11835));
NOR2X1 g78271(.A (n_2124), .B (n_4173), .Y (n_2125));
XOR2X1 g65926(.A (u0_r0_rcnt[2] ), .B (n_1204), .Y (n_6289));
MX2X1 g76020(.A (text_in_r[112] ), .B (text_in[112]), .S0 (n_1914),.Y (n_2121));
NOR2X1 g76881(.A (n_1389), .B (n_12559), .Y (n_11350));
OR2X1 g77747(.A (n_28141), .B (n_11272), .Y (n_2322));
NAND2X1 g77303(.A (n_485), .B (n_8997), .Y (n_2654));
INVX1 g77227(.A (n_2522), .Y (n_25808));
INVX1 g76807(.A (n_2113), .Y (n_2596));
INVX1 g76719(.A (n_28130), .Y (n_2112));
INVX1 g76888(.A (n_2111), .Y (n_2376));
INVX1 g77605(.A (n_2109), .Y (n_2859));
INVX1 g78183(.A (n_16976), .Y (n_2291));
INVX4 g80917(.A (n_18456), .Y (n_16754));
MX2X1 g75997(.A (text_in_r[25] ), .B (text_in[25]), .S0 (n_24599),.Y (n_2105));
INVX2 g79355(.A (n_2102), .Y (n_9923));
INVX1 g78267(.A (n_2100), .Y (n_2850));
OR2X1 g78281(.A (n_2099), .B (n_493), .Y (n_2864));
AND2X1 g78014(.A (n_26383), .B (n_2096), .Y (n_2301));
INVX1 g77724(.A (n_2094), .Y (n_2095));
INVX2 g77972(.A (n_2092), .Y (n_2093));
INVX1 g76543(.A (n_2091), .Y (n_16328));
NOR2X1 g77272(.A (n_5306), .B (n_9057), .Y (n_2090));
INVX1 g76658(.A (n_2089), .Y (n_2741));
XOR2X1 g76135(.A (n_22546), .B (n_23053), .Y (n_2086));
NAND2X2 g74720(.A (n_1294), .B (n_28567), .Y (n_2781));
INVX1 g80950(.A (n_15568), .Y (n_2888));
OR2X1 g77911(.A (n_26880), .B (n_8452), .Y (n_2295));
INVX1 g79030(.A (n_16204), .Y (n_2081));
INVX4 g79508(.A (n_736), .Y (n_2744));
NAND2X2 g76953(.A (n_1120), .B (n_2079), .Y (n_2366));
INVX1 g78093(.A (n_2078), .Y (n_2719));
XOR2X1 g76193(.A (text_in_r[127] ), .B (w0[31] ), .Y (n_2074));
NOR2X1 g74654(.A (n_1134), .B (n_827), .Y (n_2071));
NAND2X1 g77092(.A (n_2070), .B (n_2069), .Y (n_2640));
INVX1 g76644(.A (n_1868), .Y (n_3746));
MX2X1 g76005(.A (text_in_r[71] ), .B (text_in[71]), .S0 (n_25123),.Y (n_2066));
CLKBUFX3 g77936(.A (n_2382), .Y (n_3559));
CLKBUFX3 g78284(.A (n_2738), .Y (n_3643));
INVX1 g77240(.A (n_2062), .Y (n_2829));
INVX2 g77709(.A (n_1350), .Y (n_3422));
MX2X1 g75969(.A (text_in_r[115] ), .B (text_in[115]), .S0 (n_1890),.Y (n_2060));
OR2X1 g77713(.A (n_26873), .B (n_27688), .Y (n_8540));
NOR2X1 g78087(.A (n_27688), .B (n_14630), .Y (n_13423));
XOR2X1 g76263(.A (text_in_r[59] ), .B (w2[27] ), .Y (n_2055));
OR2X1 g77832(.A (n_1956), .B (n_9057), .Y (n_2053));
INVX1 g76733(.A (n_2052), .Y (n_2701));
XOR2X1 g76340(.A (text_in_r[42] ), .B (w2[10] ), .Y (n_2051));
NAND2X2 g74155(.A (n_1312), .B (n_926), .Y (n_2563));
INVX1 g77231(.A (n_27228), .Y (n_2344));
INVX1 g78048(.A (n_2048), .Y (n_2743));
MX2X1 g76076(.A (text_in_r[125] ), .B (text_in[125]), .S0 (n_619),.Y (n_2047));
INVX2 g76676(.A (n_1736), .Y (n_2680));
INVX1 g77690(.A (n_2933), .Y (n_3319));
NAND2X1 g77223(.A (n_2044), .B (n_28351), .Y (n_2787));
INVX8 g82397(.A (n_826), .Y (n_6534));
INVX1 g76557(.A (n_8099), .Y (n_2043));
NOR2X1 g77418(.A (n_872), .B (n_27204), .Y (n_2042));
INVX1 g77665(.A (n_2040), .Y (n_2628));
INVX1 g77181(.A (n_1075), .Y (n_2827));
INVX1 g78199(.A (n_15074), .Y (n_2800));
INVX1 g78221(.A (n_988), .Y (n_2714));
INVX2 g76726(.A (n_1585), .Y (n_4249));
NAND2X1 g76566(.A (n_11300), .B (n_29292), .Y (n_2394));
INVX2 g76490(.A (n_1993), .Y (n_17884));
INVX1 g78010(.A (n_26194), .Y (n_2303));
INVX1 g78212(.A (n_2025), .Y (n_2026));
XOR2X1 g76240(.A (text_in_r[106] ), .B (w0[10] ), .Y (n_2024));
INVX2 g81579(.A (n_530), .Y (n_13679));
INVX1 g77744(.A (n_2021), .Y (n_2912));
NAND2X1 g74328(.A (n_1325), .B (n_3307), .Y (n_2892));
INVX1 g76575(.A (n_4339), .Y (n_6817));
INVX1 g79897(.A (n_3566), .Y (n_2798));
INVX1 g76968(.A (n_3021), .Y (n_2281));
XOR2X1 g76339(.A (text_in_r[36] ), .B (w2[4] ), .Y (n_2013));
INVX1 g81879(.A (n_2708), .Y (n_2968));
INVX4 g80483(.A (n_19310), .Y (n_13466));
XOR2X1 g76282(.A (n_2009), .B (n_6404), .Y (n_2010));
NOR2X1 g77177(.A (n_6977), .B (n_2007), .Y (n_2008));
INVX1 g77669(.A (n_1298), .Y (n_4973));
NAND2X1 g76519(.A (n_783), .B (n_2318), .Y (n_2687));
INVX1 g76501(.A (n_1173), .Y (n_2843));
NAND2X1 g77308(.A (n_2744), .B (n_26601), .Y (n_2880));
INVX8 g81342(.A (n_20406), .Y (n_16480));
INVX1 g77192(.A (n_1998), .Y (n_2766));
INVX1 g77129(.A (n_1996), .Y (n_1997));
INVX1 g77325(.A (n_1986), .Y (n_1995));
INVX1 g81248(.A (n_1991), .Y (n_2978));
INVX4 g79765(.A (n_3017), .Y (n_2720));
NAND2X1 g77673(.A (n_1989), .B (n_28786), .Y (n_2695));
NOR2X1 g76800(.A (n_28754), .B (n_8637), .Y (n_1988));
MX2X1 g76085(.A (text_in_r[100] ), .B (text_in[100]), .S0 (ld), .Y(n_1987));
INVX1 g77324(.A (n_1986), .Y (n_2901));
NOR2X1 g78298(.A (n_2070), .B (n_26395), .Y (n_1985));
XOR2X1 g76268(.A (n_1164), .B (n_9624), .Y (n_1984));
INVX1 g76463(.A (n_1983), .Y (n_2400));
XOR2X1 g76317(.A (n_23274), .B (n_23547), .Y (n_1982));
NAND2X1 g77171(.A (n_828), .B (n_27365), .Y (n_2931));
INVX4 g80051(.A (n_18792), .Y (n_11312));
NOR2X1 g76611(.A (n_1258), .B (n_27599), .Y (n_2286));
NAND2X2 g78301(.A (n_1972), .B (n_2079), .Y (n_29360));
XOR2X1 g76271(.A (n_22762), .B (n_1970), .Y (n_1971));
MX2X1 g76026(.A (text_in_r[106] ), .B (text_in[106]), .S0 (n_619),.Y (n_1969));
XOR2X1 g76250(.A (text_in_r[105] ), .B (n_1970), .Y (n_1968));
XOR2X1 g76312(.A (text_in_r[33] ), .B (n_1039), .Y (n_1965));
NAND2X1 g77127(.A (n_28547), .B (n_28463), .Y (n_2349));
INVX1 g76741(.A (n_1818), .Y (n_3427));
INVX1 g77159(.A (n_28329), .Y (n_1963));
AND2X1 g78239(.A (n_1551), .B (n_28464), .Y (n_2278));
XOR2X1 g76228(.A (text_in_r[34] ), .B (n_1960), .Y (n_1961));
XOR2X1 g76291(.A (w0[0] ), .B (n_1958), .Y (n_1959));
INVX1 g76651(.A (n_1572), .Y (n_6871));
AND2X1 g77659(.A (n_3920), .B (n_1956), .Y (n_3489));
INVX1 g79071(.A (n_9118), .Y (n_2805));
MX2X1 g76068(.A (text_in_r[119] ), .B (text_in[119]), .S0 (n_24915),.Y (n_1955));
INVX1 g78211(.A (n_2025), .Y (n_3569));
INVX1 g76537(.A (n_2502), .Y (n_1954));
INVX2 g82520(.A (n_525), .Y (n_13593));
INVX2 g77057(.A (n_1636), .Y (n_3573));
NAND2X1 g78304(.A (n_1483), .B (n_2656), .Y (n_2911));
AND2X1 g78158(.A (n_5660), .B (n_26883), .Y (n_2292));
NAND2X1 g76618(.A (n_464), .B (n_1947), .Y (n_2392));
NAND2X1 g77258(.A (n_877), .B (n_1946), .Y (n_2409));
OR2X1 g77939(.A (n_8918), .B (n_1942), .Y (n_1943));
INVX1 g79438(.A (n_1941), .Y (n_5483));
NOR2X1 g73403(.A (n_1447), .B (n_490), .Y (n_2664));
OR2X1 g75095(.A (n_6527), .B (n_1196), .Y (n_1939));
INVX1 g76824(.A (n_2484), .Y (n_1938));
NAND2X1 g78071(.A (n_1600), .B (n_3283), .Y (n_2678));
XOR2X1 g76158(.A (n_1039), .B (n_1934), .Y (n_1936));
INVX1 g80815(.A (n_2337), .Y (n_1933));
NAND2X1 g76433(.A (n_27985), .B (n_29155), .Y (n_2446));
INVX2 g76755(.A (n_1064), .Y (n_3297));
INVX1 g80814(.A (n_2337), .Y (n_2910));
NOR2X1 g74612(.A (n_1125), .B (n_3038), .Y (n_1929));
INVX1 g78042(.A (n_1928), .Y (n_9637));
NAND2X2 g76513(.A (n_28567), .B (n_28469), .Y (n_2398));
INVX2 g77332(.A (n_1252), .Y (n_3285));
OR2X1 g78051(.A (n_9527), .B (n_4357), .Y (n_19797));
INVX1 g76794(.A (n_1377), .Y (n_5778));
INVX1 g77207(.A (n_1630), .Y (n_1923));
OR2X1 g77561(.A (n_2744), .B (n_636), .Y (n_2330));
INVX1 g77685(.A (n_1921), .Y (n_2324));
NOR2X1 g77125(.A (n_1390), .B (n_28785), .Y (n_2638));
INVX1 g77466(.A (n_2206), .Y (n_1920));
INVX1 g77531(.A (n_1918), .Y (n_2334));
XOR2X1 g76097(.A (n_1678), .B (n_22831), .Y (n_1916));
MX2X1 g76047(.A (text_in_r[76] ), .B (text_in[76]), .S0 (n_1914), .Y(n_1915));
INVX1 g76665(.A (n_1911), .Y (n_3247));
XOR2X1 g76266(.A (text_in_r[54] ), .B (w2[22] ), .Y (n_1907));
INVX1 g77796(.A (n_1905), .Y (n_2919));
INVX2 g77337(.A (n_1904), .Y (n_14757));
INVX2 g77983(.A (n_2162), .Y (n_1902));
CLKBUFX3 g80398(.A (n_5203), .Y (n_7725));
MX2X1 g75994(.A (text_in_r[87] ), .B (text_in[87]), .S0 (ld), .Y(n_1899));
INVX1 g77188(.A (n_1897), .Y (n_2713));
MX2X1 g75986(.A (text_in_r[98] ), .B (text_in[98]), .S0 (ld), .Y(n_1895));
MX2X1 g75970(.A (text_in_r[117] ), .B (text_in[117]), .S0 (n_1890),.Y (n_1891));
NAND2X1 g74515(.A (n_1284), .B (n_4568), .Y (n_2335));
INVX1 g77850(.A (n_1888), .Y (n_12858));
INVX1 g80203(.A (n_1887), .Y (n_2323));
NOR2X1 g77848(.A (u0_r0_rcnt[0] ), .B (ld), .Y (n_2710));
INVX1 g77817(.A (n_1443), .Y (n_1886));
INVX2 g77343(.A (n_1387), .Y (n_3246));
NOR2X1 g76994(.A (n_1339), .B (n_8974), .Y (n_14667));
NOR2X1 g77139(.A (n_674), .B (n_6185), .Y (n_1883));
AND2X1 g77930(.A (n_28576), .B (n_28476), .Y (n_2351));
NOR2X1 g78121(.A (n_29102), .B (n_9368), .Y (n_11739));
NOR2X1 g77752(.A (n_28478), .B (n_28576), .Y (n_2831));
INVX8 g82275(.A (n_3886), .Y (n_16835));
INVX2 g76702(.A (n_29131), .Y (n_3252));
NAND2X1 g77698(.A (n_1228), .B (n_27204), .Y (n_28488));
INVX1 g77437(.A (n_962), .Y (n_2671));
INVX1 g77956(.A (n_2076), .Y (n_4217));
INVX2 g79148(.A (n_713), .Y (n_12105));
XOR2X1 g76156(.A (text_in_r[43] ), .B (w2[11] ), .Y (n_1858));
NAND2X2 g75559(.A (n_1212), .B (n_1292), .Y (n_2267));
INVX2 g78729(.A (n_828), .Y (n_17571));
XOR2X1 g76244(.A (text_in_r[40] ), .B (w2[8] ), .Y (n_1854));
MX2X1 g76064(.A (text_in_r[83] ), .B (text_in[83]), .S0 (n_1914), .Y(n_1852));
MX2X1 g75996(.A (text_in_r[62] ), .B (text_in[62]), .S0 (ld), .Y(n_1851));
OR2X1 g78156(.A (n_11489), .B (n_187), .Y (n_2682));
INVX2 g81244(.A (n_1991), .Y (n_20862));
INVX2 g77615(.A (n_1256), .Y (n_2684));
XOR2X1 g76237(.A (text_in_r[68] ), .B (w1[4] ), .Y (n_1845));
XOR2X1 g76251(.A (n_1842), .B (n_22750), .Y (n_1843));
INVX1 g76998(.A (n_2444), .Y (n_2852));
MX2X1 g76030(.A (text_in_r[124] ), .B (text_in[124]), .S0 (n_619),.Y (n_1840));
INVX1 g77548(.A (n_1839), .Y (n_3517));
NOR2X1 g76924(.A (n_9106), .B (sa22[1] ), .Y (n_20065));
INVX1 g76524(.A (n_1837), .Y (n_2627));
NAND2X2 g77312(.A (n_1395), .B (n_214), .Y (n_2792));
NAND2X1 g76812(.A (n_1956), .B (n_2239), .Y (n_2807));
AND2X1 g76774(.A (n_12760), .B (w3[9] ), .Y (n_10191));
XOR2X1 g76212(.A (w2[10] ), .B (w0[10] ), .Y (n_1833));
NAND2X2 g77046(.A (n_1258), .B (n_1460), .Y (n_2496));
INVX1 g73303(.A (n_2848), .Y (n_1827));
INVX1 g78144(.A (n_5149), .Y (n_2839));
NAND2X2 g77107(.A (n_8918), .B (n_1823), .Y (n_1825));
INVX1 g77551(.A (n_1822), .Y (n_6587));
NOR2X1 g78193(.A (n_1569), .B (n_320), .Y (n_1821));
INVX1 g76742(.A (n_1818), .Y (n_1819));
AND2X1 g77559(.A (n_2099), .B (n_2492), .Y (n_2332));
INVX1 g77390(.A (n_1817), .Y (n_2265));
MX2X1 g76060(.A (text_in_r[43] ), .B (text_in[43]), .S0 (ld), .Y(n_1816));
OR2X1 g76725(.A (n_1142), .B (n_1376), .Y (n_9195));
INVX1 g77359(.A (n_26994), .Y (n_3023));
MX2X1 g76061(.A (text_in_r[72] ), .B (text_in[72]), .S0 (n_24778),.Y (n_1813));
INVX1 g77034(.A (n_1777), .Y (n_2357));
XOR2X1 g76308(.A (text_in_r[49] ), .B (n_22976), .Y (n_1811));
XOR2X1 g76200(.A (text_in_r[58] ), .B (w2[26] ), .Y (n_1809));
INVX1 g76746(.A (n_1807), .Y (n_6870));
INVX1 g76976(.A (n_1806), .Y (n_7803));
MX2X1 g76018(.A (text_in_r[48] ), .B (text_in[48]), .S0 (n_25123),.Y (n_1805));
INVX4 g79176(.A (n_427), .Y (n_15388));
OR2X1 g77567(.A (n_27098), .B (n_26493), .Y (n_5691));
INVX1 g79234(.A (n_27985), .Y (n_3493));
NOR2X1 g77218(.A (n_1110), .B (n_29225), .Y (n_4676));
INVX1 g77212(.A (n_1267), .Y (n_2723));
AND2X1 g77626(.A (n_463), .B (n_218), .Y (n_2820));
NAND2X1 g76984(.A (n_214), .B (n_1627), .Y (n_2365));
AND2X1 g77814(.A (n_1512), .B (n_3318), .Y (n_19110));
MX2X1 g75995(.A (text_in_r[4] ), .B (text_in[4]), .S0 (n_24599), .Y(n_1798));
XOR2X1 g76165(.A (n_22750), .B (n_1385), .Y (n_1797));
NAND2X1 g78177(.A (n_26276), .B (n_7331), .Y (n_7418));
INVX2 g77158(.A (n_28328), .Y (n_3002));
INVX2 g80691(.A (n_1792), .Y (n_8560));
NOR2X1 g78235(.A (n_27985), .B (n_29158), .Y (n_1791));
INVX1 g78098(.A (n_1789), .Y (n_2298));
INVX1 g78063(.A (n_1788), .Y (n_2707));
AND2X1 g76801(.A (n_15776), .B (sa33[1] ), .Y (n_14741));
XOR2X1 g76140(.A (n_23545), .B (n_1005), .Y (n_1786));
XOR2X1 g76221(.A (text_in_r[87] ), .B (w1[23] ), .Y (n_1784));
AND2X1 g76804(.A (n_14592), .B (sa31[1] ), .Y (n_14854));
INVX1 g77073(.A (n_1782), .Y (n_3813));
NOR2X1 g75846(.A (n_1313), .B (n_2462), .Y (n_1781));
OR2X1 g76542(.A (n_1046), .B (n_6868), .Y (n_1779));
NAND2X1 g73422(.A (n_1370), .B (n_6021), .Y (n_1775));
NAND2X1 g76981(.A (n_853), .B (n_3038), .Y (n_3816));
INVX2 g77201(.A (n_1278), .Y (n_3585));
INVX1 g78204(.A (n_1772), .Y (n_2748));
INVX2 g76991(.A (n_1248), .Y (n_3267));
INVX1 g76830(.A (n_1771), .Y (n_3420));
XOR2X1 g76349(.A (n_2560), .B (n_1769), .Y (n_1770));
INVX1 g76836(.A (n_1768), .Y (n_15997));
NAND2X1 g76917(.A (n_1634), .B (n_27668), .Y (n_2374));
MX2X1 g76084(.A (text_in_r[57] ), .B (text_in[57]), .S0 (ld), .Y(n_1763));
OR2X1 g78136(.A (n_11300), .B (n_29244), .Y (n_8139));
XOR2X1 g76242(.A (text_in_r[45] ), .B (n_23001), .Y (n_1760));
XOR2X1 g76327(.A (text_in_r[82] ), .B (w1[18] ), .Y (n_1758));
INVX2 g81020(.A (n_1756), .Y (n_12896));
INVX1 g79453(.A (n_1198), .Y (n_3834));
NOR2X1 g75324(.A (n_1609), .B (n_490), .Y (n_3600));
MX2X1 g75987(.A (text_in_r[94] ), .B (text_in[94]), .S0 (ld), .Y(n_1752));
INVX1 g81601(.A (n_1750), .Y (n_2972));
XOR2X1 g76198(.A (text_in_r[109] ), .B (n_23087), .Y (n_1749));
NOR2X1 g77483(.A (n_2943), .B (n_720), .Y (n_1748));
INVX1 g76484(.A (n_1743), .Y (n_1747));
INVX1 g76791(.A (n_1746), .Y (n_5179));
NOR2X1 g76766(.A (n_791), .B (n_4173), .Y (n_1744));
INVX1 g79442(.A (n_2084), .Y (n_6783));
NAND2X1 g76886(.A (n_18456), .B (n_6005), .Y (n_2900));
OR2X1 g76597(.A (n_9527), .B (w3[25] ), .Y (n_17020));
INVX1 g77510(.A (n_2541), .Y (n_2969));
INVX1 g76483(.A (n_1743), .Y (n_2885));
INVX2 g77608(.A (n_1742), .Y (n_3590));
NOR2X1 g75615(.A (n_1307), .B (n_27204), .Y (n_1741));
INVX1 g78899(.A (n_3014), .Y (n_5236));
AND2X1 g77706(.A (n_8918), .B (n_1739), .Y (n_2608));
NOR2X1 g78246(.A (n_18266), .B (n_5131), .Y (n_13575));
INVX1 g76677(.A (n_1736), .Y (n_1737));
INVX1 g76630(.A (n_976), .Y (n_6827));
MX2X1 g76082(.A (text_in_r[109] ), .B (text_in[109]), .S0 (n_24915),.Y (n_1734));
MX2X1 g75990(.A (text_in_r[89] ), .B (text_in[89]), .S0 (n_24599),.Y (n_1731));
NOR2X1 g77815(.A (n_4300), .B (n_7485), .Y (n_8674));
INVX1 g78378(.A (n_20198), .Y (n_21507));
XOR2X1 g76153(.A (text_in_r[55] ), .B (w2[23] ), .Y (n_1727));
XOR2X1 g76269(.A (n_2434), .B (n_1960), .Y (n_1724));
NAND2X1 g76510(.A (n_1989), .B (n_28779), .Y (n_2774));
INVX4 g82111(.A (n_827), .Y (n_2959));
INVX1 g80618(.A (n_5305), .Y (n_23418));
NOR2X1 g77652(.A (n_9442), .B (n_9368), .Y (n_4544));
OR2X1 g78105(.A (n_8708), .B (n_19486), .Y (n_2663));
INVX2 g80119(.A (n_1717), .Y (n_10255));
XOR2X1 g76100(.A (text_in_r[69] ), .B (w1[5] ), .Y (n_1712));
OR2X1 g74264(.A (n_1324), .B (n_1711), .Y (n_2480));
NAND2X1 g74623(.A (n_26185), .B (n_28786), .Y (n_2823));
INVX1 g77942(.A (n_1707), .Y (n_4326));
INVX1 g81026(.A (n_15574), .Y (n_2983));
NAND2X2 g75388(.A (n_1166), .B (n_2096), .Y (n_2464));
XOR2X1 g76120(.A (text_in_r[46] ), .B (w2[14] ), .Y (n_1706));
AND2X1 g77831(.A (n_12827), .B (n_1701), .Y (n_16988));
INVX1 g76684(.A (n_1233), .Y (n_10680));
INVX2 g77679(.A (n_1306), .Y (n_3448));
INVX2 g76870(.A (n_26546), .Y (n_3373));
INVX1 g81190(.A (sa31[1] ), .Y (n_21581));
MX2X1 g75973(.A (text_in_r[21] ), .B (text_in[21]), .S0 (n_1890), .Y(n_1698));
INVX2 g78918(.A (n_1358), .Y (n_6303));
INVX1 g79881(.A (n_19995), .Y (n_2909));
NAND2X1 g77020(.A (n_1347), .B (n_7331), .Y (n_1695));
INVX1 g66589(.A (n_1693), .Y (n_1694));
OR2X1 g78140(.A (n_9917), .B (n_27045), .Y (n_19961));
XOR2X1 g76148(.A (text_in_r[62] ), .B (w2[30] ), .Y (n_1691));
INVX4 g79317(.A (n_14878), .Y (n_14866));
NOR2X1 g76802(.A (n_28362), .B (n_7498), .Y (n_1688));
INVX1 g77260(.A (n_1289), .Y (n_2342));
INVX1 g78252(.A (n_1685), .Y (n_1686));
INVX1 g81531(.A (n_11277), .Y (n_18326));
XOR2X1 g76226(.A (n_255), .B (n_6404), .Y (n_1683));
INVX1 g77477(.A (n_2017), .Y (n_3288));
INVX1 g82521(.A (n_525), .Y (n_12917));
XOR2X1 g76149(.A (n_22789), .B (n_1678), .Y (n_1679));
INVX1 g82548(.A (n_27747), .Y (n_13834));
INVX1 g77594(.A (n_1261), .Y (n_3482));
NOR2X1 g76530(.A (n_214), .B (n_1627), .Y (n_2818));
XOR2X1 g76184(.A (n_22787), .B (n_1674), .Y (n_1675));
INVX4 g82168(.A (n_26874), .Y (n_9783));
INVX1 g78037(.A (n_1102), .Y (n_2865));
NOR2X1 g78123(.A (n_3108), .B (n_28375), .Y (n_1671));
INVX1 g77492(.A (n_9755), .Y (n_1668));
XOR2X1 g76167(.A (n_1235), .B (n_16938), .Y (n_1666));
NAND2X2 g77149(.A (n_4837), .B (n_493), .Y (n_29214));
INVX1 g76430(.A (n_960), .Y (n_3833));
NOR2X1 g76536(.A (n_393), .B (n_367), .Y (n_4093));
XOR2X1 g76124(.A (text_in_r[79] ), .B (w1[15] ), .Y (n_1658));
NAND2X1 g77536(.A (n_12760), .B (n_12169), .Y (n_5735));
XOR2X1 g76172(.A (text_in_r[41] ), .B (n_22762), .Y (n_1656));
MX2X1 g76055(.A (text_in_r[73] ), .B (text_in[73]), .S0 (n_25123),.Y (n_1653));
NAND2X1 g77569(.A (n_28734), .B (n_7496), .Y (n_4382));
INVX2 g80124(.A (n_1651), .Y (n_8339));
MX2X1 g75982(.A (text_in_r[95] ), .B (text_in[95]), .S0 (n_24915),.Y (n_1648));
NAND2X1 g78031(.A (n_18266), .B (n_1647), .Y (n_3281));
INVX2 g79798(.A (n_26490), .Y (n_11052));
MX2X1 g76046(.A (text_in_r[38] ), .B (text_in[38]), .S0 (ld), .Y(n_1645));
OR2X1 g77846(.A (n_1230), .B (n_27746), .Y (n_1644));
NAND2X1 g77641(.A (n_7636), .B (n_9118), .Y (n_4928));
OR2X1 g77920(.A (n_493), .B (n_1431), .Y (n_2930));
INVX1 g81938(.A (n_1642), .Y (n_8467));
INVX2 g80138(.A (n_1641), .Y (n_23422));
NOR2X1 g77758(.A (n_1427), .B (n_3296), .Y (n_2875));
INVX1 g77054(.A (n_1636), .Y (n_1637));
AND2X1 g77829(.A (n_1634), .B (n_2235), .Y (n_2568));
XOR2X1 g76191(.A (n_1632), .B (w1[31] ), .Y (n_1633));
CLKBUFX1 g78019(.A (n_2621), .Y (n_5530));
INVX1 g76437(.A (n_1333), .Y (n_2401));
INVX2 g77702(.A (n_1051), .Y (n_3346));
INVX1 g77206(.A (n_1630), .Y (n_3121));
NAND2X1 g76588(.A (n_1628), .B (n_1627), .Y (n_3096));
INVX1 g77776(.A (n_2145), .Y (n_3314));
NAND2X1 g76899(.A (n_20406), .B (n_6226), .Y (n_2873));
INVX1 g81754(.A (n_1621), .Y (n_3696));
INVX1 g77279(.A (n_1620), .Y (n_2469));
XOR2X1 g76223(.A (n_16921), .B (n_23047), .Y (n_1618));
INVX1 g79679(.A (n_1616), .Y (n_2870));
INVX1 g76690(.A (n_1615), .Y (n_6510));
OR2X1 g77896(.A (n_12760), .B (n_933), .Y (n_2718));
XOR2X1 g76302(.A (n_9), .B (w1[25] ), .Y (n_1614));
INVX1 g78125(.A (n_16553), .Y (n_1610));
OR2X1 g75572(.A (n_1609), .B (n_3599), .Y (n_8662));
XOR2X1 g76283(.A (text_in_r[60] ), .B (w2[28] ), .Y (n_1608));
XOR2X1 g76186(.A (n_23241), .B (n_22833), .Y (n_1606));
OR2X1 g78180(.A (n_160), .B (n_3283), .Y (n_2488));
OR2X1 g77495(.A (n_17912), .B (n_310), .Y (n_16579));
INVX1 g79635(.A (n_6805), .Y (n_1603));
NAND2X2 g77353(.A (n_2383), .B (n_557), .Y (n_2925));
NAND2X1 g77119(.A (n_931), .B (n_2343), .Y (n_2536));
INVX2 g78882(.A (n_1601), .Y (n_3512));
NAND2X1 g76920(.A (n_1600), .B (n_6431), .Y (n_2372));
NAND2X1 g77870(.A (n_636), .B (n_2343), .Y (n_1599));
CLKBUFX1 g79018(.A (n_2359), .Y (n_3735));
CLKBUFX1 g78744(.A (n_27099), .Y (n_18679));
NOR2X1 g75541(.A (n_1263), .B (n_827), .Y (n_1594));
INVX1 g79556(.A (n_26619), .Y (n_1593));
OR2X1 g78131(.A (n_664), .B (n_3038), .Y (n_2613));
INVX2 g80578(.A (n_1591), .Y (n_2777));
OR2X1 g75028(.A (n_7411), .B (n_379), .Y (n_2923));
XOR2X1 g76138(.A (text_in_r[91] ), .B (n_332), .Y (n_1589));
MX2X1 g75971(.A (text_in_r[122] ), .B (text_in[122]), .S0 (n_24915),.Y (n_1588));
INVX2 g78919(.A (n_1358), .Y (n_1584));
NAND2X1 g77419(.A (n_14807), .B (n_19486), .Y (n_1582));
NOR2X1 g77022(.A (n_4861), .B (n_1508), .Y (n_2360));
INVX1 g77515(.A (n_1581), .Y (n_2424));
NAND2X1 g77428(.A (n_3067), .B (n_1244), .Y (n_2305));
AND2X1 g77001(.A (n_26276), .B (sa32[1] ), .Y (n_2362));
MX2X1 g76041(.A (text_in_r[44] ), .B (text_in[44]), .S0 (n_24778),.Y (n_1578));
INVX1 g78917(.A (n_1358), .Y (n_8816));
NOR2X1 g74215(.A (n_1191), .B (n_3038), .Y (n_3365));
INVX1 g79602(.A (n_624), .Y (n_19385));
OR2X1 g77505(.A (n_9202), .B (n_3318), .Y (n_1571));
NAND2X2 g77060(.A (n_1569), .B (n_1568), .Y (n_1570));
INVX1 g77488(.A (n_4327), .Y (n_2548));
XOR2X1 g76116(.A (text_in_r[104] ), .B (w0[8] ), .Y (n_1565));
XOR2X1 g76123(.A (n_22976), .B (n_22567), .Y (n_1564));
XOR2X1 g76127(.A (n_23309), .B (n_23763), .Y (n_1562));
XOR2X1 g76128(.A (n_22964), .B (w1[27] ), .Y (n_1560));
INVX1 g82068(.A (n_1558), .Y (n_2826));
XOR2X1 g76144(.A (n_1555), .B (n_22557), .Y (n_1556));
INVX1 g79333(.A (n_2063), .Y (n_1553));
NAND2X2 g77015(.A (n_1551), .B (n_28463), .Y (n_1552));
INVX1 g77971(.A (n_2092), .Y (n_2514));
NOR2X1 g77621(.A (n_2211), .B (n_2343), .Y (n_1548));
MX2X1 g76045(.A (text_in_r[114] ), .B (text_in[114]), .S0 (n_24778),.Y (n_1546));
XOR2X1 g76298(.A (n_1163), .B (n_9624), .Y (n_1544));
XOR2X1 g76300(.A (text_in_r[97] ), .B (n_1934), .Y (n_1542));
MX2X1 g76027(.A (text_in_r[101] ), .B (text_in[101]), .S0 (n_1914),.Y (n_1541));
NAND2X2 g77475(.A (n_1540), .B (n_1353), .Y (n_2402));
NAND2X1 g77268(.A (n_274), .B (n_9368), .Y (n_2404));
INVX1 g77631(.A (n_1082), .Y (n_2594));
INVX1 g79664(.A (n_1142), .Y (n_2760));
NAND2X1 g77315(.A (n_896), .B (n_1539), .Y (n_2889));
INVX1 g76496(.A (n_1538), .Y (n_2755));
NOR2X1 g76531(.A (n_12298), .B (sa11[1] ), .Y (n_18876));
INVX1 g76602(.A (n_1335), .Y (n_2266));
INVX1 g77264(.A (n_1264), .Y (n_2835));
NOR2X1 g76803(.A (n_11261), .B (sa20[1] ), .Y (n_20271));
INVX1 g76878(.A (n_1534), .Y (n_3535));
NOR2X1 g76930(.A (n_1423), .B (n_8878), .Y (n_4194));
INVX1 g77023(.A (n_1530), .Y (n_1531));
NAND2X1 g77083(.A (n_706), .B (n_7593), .Y (n_2353));
NAND2X1 g77102(.A (sa00[2] ), .B (n_4709), .Y (n_2513));
MX2X1 g76029(.A (text_in_r[113] ), .B (text_in[113]), .S0 (ld), .Y(n_1528));
XOR2X1 g76272(.A (n_1103), .B (w1[31] ), .Y (n_1526));
INVX1 g78251(.A (n_1685), .Y (n_2447));
MX2X1 g75988(.A (text_in_r[93] ), .B (text_in[93]), .S0 (ld), .Y(n_1525));
INVX2 g77174(.A (n_27203), .Y (n_3128));
INVX1 g77459(.A (n_1522), .Y (n_2861));
OR2X1 g77327(.A (n_9342), .B (w3[17] ), .Y (n_17023));
AND2X1 g77183(.A (n_14624), .B (sa30[1] ), .Y (n_13176));
NAND2X1 g76586(.A (n_1238), .B (n_14055), .Y (n_2526));
NAND2X1 g76929(.A (n_9819), .B (n_1153), .Y (n_2617));
CLKBUFX3 g77378(.A (n_1516), .Y (n_3465));
INVX8 g80941(.A (sa30[2] ), .Y (n_14624));
INVX1 g77542(.A (n_1513), .Y (n_3160));
AND2X1 g77449(.A (n_11385), .B (n_933), .Y (n_15516));
NAND2X1 g76943(.A (n_1512), .B (n_751), .Y (n_2575));
INVX1 g77441(.A (n_1874), .Y (n_2336));
INVX1 g77600(.A (n_2534), .Y (n_2611));
NAND2X1 g76521(.A (n_8865), .B (n_1508), .Y (n_1509));
INVX2 g77368(.A (n_1098), .Y (n_3322));
MX2X1 g76071(.A (text_in_r[102] ), .B (text_in[102]), .S0 (ld), .Y(n_1507));
NAND2X1 g76624(.A (n_688), .B (n_29228), .Y (n_2307));
NOR2X1 g77867(.A (n_1456), .B (n_27204), .Y (n_1505));
INVX1 g77907(.A (n_1503), .Y (n_2724));
INVX1 g80204(.A (n_1887), .Y (n_1502));
INVX1 g67824(.A (n_6301), .Y (n_1501));
XOR2X1 g76201(.A (n_982), .B (n_9203), .Y (n_1500));
INVX1 g77979(.A (n_12850), .Y (n_1497));
INVX1 g77052(.A (n_3198), .Y (n_2757));
OR2X1 g78059(.A (n_18266), .B (n_4709), .Y (n_8191));
NOR2X1 g77433(.A (n_2744), .B (n_26989), .Y (n_1494));
NAND2X2 g77904(.A (n_1493), .B (n_28476), .Y (n_2715));
OR2X1 g78060(.A (n_1551), .B (n_26873), .Y (n_1491));
NOR2X1 g77900(.A (n_28547), .B (n_28464), .Y (n_1488));
NAND2X1 g78116(.A (n_6185), .B (n_4627), .Y (n_2466));
INVX4 g78392(.A (n_1484), .Y (n_2960));
NAND2X1 g76875(.A (n_1483), .B (n_1069), .Y (n_2604));
INVX2 g78432(.A (n_2231), .Y (n_3069));
NAND2X1 g77276(.A (sa01[2] ), .B (n_8452), .Y (n_2276));
INVX4 g78650(.A (n_877), .Y (n_15708));
NOR2X1 g78054(.A (n_3301), .B (n_12169), .Y (n_4375));
INVX1 g76547(.A (n_1480), .Y (n_3091));
INVX1 g80984(.A (n_1310), .Y (n_17775));
INVX1 g81765(.A (n_581), .Y (n_7419));
XOR2X1 g76324(.A (text_in_r[51] ), .B (w2[19] ), .Y (n_1477));
INVX1 g78930(.A (n_2187), .Y (n_9691));
XOR2X1 g76331(.A (text_in_r[53] ), .B (w2[21] ), .Y (n_1473));
INVX1 g79449(.A (n_1198), .Y (n_9416));
NOR2X1 g76946(.A (n_379), .B (n_1251), .Y (n_3310));
NOR2X1 g77884(.A (n_1483), .B (n_1460), .Y (n_1461));
INVX2 g76958(.A (n_1331), .Y (n_2908));
MX2X1 g75974(.A (text_in_r[22] ), .B (text_in[22]), .S0 (n_1890), .Y(n_1457));
AND2X1 g77932(.A (n_1456), .B (n_27204), .Y (n_2635));
INVX1 g79873(.A (n_14627), .Y (n_20610));
NOR2X1 g76782(.A (n_821), .B (n_9084), .Y (n_13875));
NOR2X1 g77880(.A (n_4364), .B (n_28375), .Y (n_2311));
INVX1 g78268(.A (n_749), .Y (n_2100));
INVX2 g81733(.A (n_1124), .Y (n_8910));
NAND2X1 g77852(.A (n_17411), .B (n_9118), .Y (n_1888));
NAND2X1 g66590(.A (n_1448), .B (n_328), .Y (n_1693));
INVX1 g77408(.A (n_1447), .Y (n_2716));
INVX1 g80816(.A (n_1157), .Y (n_2337));
NOR2X1 g77818(.A (n_1080), .B (n_276), .Y (n_1443));
INVX1 g77391(.A (n_435), .Y (n_1817));
INVX1 g80411(.A (n_196), .Y (n_20162));
OR2X1 g77849(.A (n_1332), .B (n_6868), .Y (n_1441));
INVX1 g78433(.A (n_3695), .Y (n_2231));
INVX1 g77555(.A (n_7899), .Y (n_16090));
NOR2X1 g76577(.A (n_264), .B (n_271), .Y (n_4339));
INVX1 g79882(.A (n_21242), .Y (n_19995));
AND2X1 g77549(.A (n_100), .B (n_1431), .Y (n_1839));
INVX2 g77527(.A (n_1430), .Y (n_2583));
XOR2X1 g76290(.A (n_23551), .B (n_1428), .Y (n_1429));
INVX2 g79770(.A (n_26486), .Y (n_2241));
INVX1 g81755(.A (n_1427), .Y (n_1621));
INVX8 g82162(.A (n_26874), .Y (n_8452));
BUFX3 g81030(.A (n_27133), .Y (n_15574));
INVX2 g80503(.A (n_1423), .Y (n_5922));
XOR2X1 g76307(.A (n_2648), .B (w1[16] ), .Y (n_1417));
INVX1 g77543(.A (n_1416), .Y (n_1513));
NAND2X1 g77280(.A (n_100), .B (n_1201), .Y (n_1620));
XOR2X1 g76125(.A (n_23079), .B (n_23274), .Y (n_1409));
INVX1 g81072(.A (n_20661), .Y (n_21382));
NAND2X1 g76999(.A (n_514), .B (n_3283), .Y (n_2444));
AND2X1 g77489(.A (n_386), .B (n_271), .Y (n_4327));
INVX1 g78936(.A (n_783), .Y (n_6092));
INVX2 g78458(.A (n_1053), .Y (n_8263));
INVX1 g77908(.A (n_871), .Y (n_1503));
INVX1 g78106(.A (n_7411), .Y (n_1402));
INVX1 g81854(.A (n_1397), .Y (n_2249));
INVX1 g81605(.A (n_1395), .Y (n_1396));
INVX2 g80288(.A (n_819), .Y (n_5558));
NAND2X1 g76692(.A (n_11354), .B (n_941), .Y (n_1615));
CLKBUFX3 g77601(.A (n_1016), .Y (n_2534));
INVX2 g80120(.A (n_27124), .Y (n_1717));
NAND2X2 g76894(.A (n_1390), .B (n_28793), .Y (n_2067));
NAND2X1 g76792(.A (n_1389), .B (n_4861), .Y (n_1746));
CLKBUFX1 g81031(.A (n_27133), .Y (n_16414));
INVX2 g82489(.A (n_1634), .Y (n_2218));
NAND2X1 g77344(.A (n_1260), .B (n_462), .Y (n_1387));
XOR2X1 g76110(.A (n_1842), .B (n_1385), .Y (n_1386));
NAND2X1 g77340(.A (n_15655), .B (n_7325), .Y (n_1904));
INVX1 g81816(.A (n_4898), .Y (n_1830));
INVX1 g77797(.A (n_1384), .Y (n_1905));
CLKBUFX3 g79019(.A (n_1456), .Y (n_2359));
INVX1 g78274(.A (n_6527), .Y (n_1378));
NAND2X1 g76795(.A (n_3955), .B (n_1376), .Y (n_1377));
INVX4 g82189(.A (n_1373), .Y (n_11323));
NOR2X1 g78065(.A (n_862), .B (n_1627), .Y (n_1788));
INVX1 g77781(.A (n_1370), .Y (n_1371));
INVX1 g79755(.A (n_27370), .Y (n_5186));
INVX1 g79271(.A (n_1196), .Y (n_19942));
NAND2X2 g77058(.A (n_1255), .B (n_167), .Y (n_1636));
INVX2 g77502(.A (n_1363), .Y (n_7649));
INVX1 g78162(.A (n_12849), .Y (n_1361));
INVX1 g77467(.A (n_459), .Y (n_2206));
INVX1 g81643(.A (n_1316), .Y (n_2830));
INVX1 g79650(.A (n_1508), .Y (n_2180));
NAND2X1 g76666(.A (n_454), .B (n_1291), .Y (n_1911));
INVX1 g78316(.A (n_62), .Y (n_21151));
INVX1 g80863(.A (n_688), .Y (n_14474));
INVX2 g80798(.A (n_1353), .Y (n_2085));
INVX2 g81153(.A (n_399), .Y (n_16198));
INVX1 g80661(.A (n_2044), .Y (n_2237));
NOR2X1 g77710(.A (n_1305), .B (n_28793), .Y (n_1350));
INVX1 g80449(.A (n_15674), .Y (n_19111));
INVX1 g79356(.A (n_9368), .Y (n_2102));
NAND2X1 g77053(.A (n_1000), .B (n_2318), .Y (n_3198));
XOR2X1 g76202(.A (n_112), .B (n_1296), .Y (n_1341));
CLKBUFX1 g79435(.A (n_3534), .Y (n_7127));
INVX1 g81183(.A (n_1336), .Y (n_1925));
INVX2 g78020(.A (n_913), .Y (n_2621));
NAND2X1 g76603(.A (n_968), .B (n_218), .Y (n_1335));
INVX1 g78636(.A (n_1569), .Y (n_1735));
INVX4 g79766(.A (n_27370), .Y (n_3017));
NAND2X1 g76438(.A (n_1332), .B (n_348), .Y (n_1333));
NAND2X2 g76959(.A (n_870), .B (n_107), .Y (n_1331));
INVX1 g82319(.A (n_933), .Y (n_1699));
INVX1 g82028(.A (n_3264), .Y (n_20632));
INVX1 g77666(.A (n_917), .Y (n_2040));
INVX2 g77984(.A (n_901), .Y (n_2162));
NAND2X1 g77131(.A (n_607), .B (n_2959), .Y (n_1996));
INVX1 g77413(.A (n_1325), .Y (n_2742));
INVX1 g77228(.A (n_1242), .Y (n_2522));
INVX1 g81936(.A (n_1946), .Y (n_2107));
INVX1 g76525(.A (n_1324), .Y (n_1837));
INVX1 g77097(.A (n_473), .Y (n_2950));
XOR2X1 g76234(.A (text_in_r[48] ), .B (n_2648), .Y (n_1321));
INVX4 g78466(.A (n_1053), .Y (n_10452));
XOR2X1 g76320(.A (n_1318), .B (n_1220), .Y (n_1319));
INVX1 g78439(.A (n_1315), .Y (n_3327));
INVX1 g78026(.A (n_1313), .Y (n_3491));
INVX2 g81791(.A (n_902), .Y (n_9257));
INVX1 g77957(.A (n_1312), .Y (n_2076));
XOR2X1 g76173(.A (n_1428), .B (n_1308), .Y (n_1309));
NAND2X1 g76548(.A (n_1302), .B (n_400), .Y (n_1480));
INVX2 g77516(.A (n_623), .Y (n_1581));
NAND2X1 g77208(.A (n_469), .B (n_537), .Y (n_1630));
INVX2 g77691(.A (n_1307), .Y (n_2933));
NAND2X2 g77680(.A (n_1305), .B (n_748), .Y (n_1306));
NAND2X1 g77074(.A (n_900), .B (n_834), .Y (n_1782));
INVX1 g77379(.A (n_802), .Y (n_1516));
INVX4 g79168(.A (n_523), .Y (n_14484));
CLKBUFX1 g79575(.A (n_9819), .Y (n_17377));
INVX1 g80693(.A (n_3234), .Y (n_1792));
NOR2X1 g77670(.A (n_1050), .B (n_1627), .Y (n_1298));
XOR2X1 g76299(.A (n_1296), .B (n_2692), .Y (n_1297));
NAND2X1 g76646(.A (n_775), .B (n_1043), .Y (n_1868));
INVX1 g77770(.A (n_1294), .Y (n_2137));
INVX2 g78409(.A (n_3038), .Y (n_2239));
AND2X1 g77725(.A (n_1292), .B (n_1291), .Y (n_2094));
NOR2X1 g77261(.A (sa21[1] ), .B (n_29102), .Y (n_1289));
NOR2X1 g76538(.A (n_2943), .B (n_719), .Y (n_2502));
INVX1 g79942(.A (n_360), .Y (n_3340));
INVX2 g77777(.A (n_579), .Y (n_2145));
NAND2X1 g77326(.A (n_629), .B (n_1285), .Y (n_1986));
XOR2X1 g76163(.A (text_in_r[38] ), .B (n_2437), .Y (n_1283));
INVX1 g77292(.A (n_584), .Y (n_1930));
NOR2X1 g77745(.A (n_28749), .B (n_7496), .Y (n_2021));
INVX4 g81156(.A (n_399), .Y (n_13490));
NAND2X1 g76479(.A (n_575), .B (n_28464), .Y (n_1282));
NAND2X1 g76748(.A (n_9106), .B (n_713), .Y (n_1807));
XOR2X1 g76181(.A (n_22496), .B (n_22762), .Y (n_1281));
INVX1 g78253(.A (n_803), .Y (n_1685));
INVX2 g81957(.A (n_6052), .Y (n_2022));
XOR2X1 g76314(.A (u0_r0_rcnt[1] ), .B (n_111), .Y (n_2848));
NAND2X2 g77202(.A (n_479), .B (n_919), .Y (n_1278));
INVX2 g79486(.A (n_1483), .Y (n_2254));
INVX1 g78094(.A (n_632), .Y (n_2078));
INVX1 g77532(.A (n_833), .Y (n_1918));
INVX2 g77937(.A (n_850), .Y (n_2382));
NAND2X1 g76464(.A (n_3868), .B (n_1273), .Y (n_1983));
NAND2X1 g76728(.A (n_1292), .B (n_1272), .Y (n_1585));
XOR2X1 g76270(.A (n_22964), .B (n_1270), .Y (n_1271));
INVX1 g77461(.A (n_538), .Y (n_1522));
OR2X1 g77552(.A (n_1014), .B (n_3038), .Y (n_1822));
NAND2X1 g77213(.A (n_612), .B (n_26382), .Y (n_1267));
INVX2 g80205(.A (n_1266), .Y (n_1887));
AND2X1 g78043(.A (n_28167), .B (n_1147), .Y (n_1928));
NOR2X1 g77265(.A (n_384), .B (n_178), .Y (n_1264));
INVX1 g77788(.A (n_1263), .Y (n_2530));
OR2X1 g78169(.A (n_263), .B (n_2810), .Y (n_6889));
NOR2X1 g77595(.A (n_1260), .B (n_218), .Y (n_1261));
INVX1 g80237(.A (n_1258), .Y (n_3597));
INVX1 g78006(.A (n_11850), .Y (n_14348));
INVX1 g77687(.A (n_665), .Y (n_1921));
NAND2X2 g77616(.A (n_1255), .B (n_1081), .Y (n_1256));
XOR2X1 g76143(.A (n_22591), .B (n_22976), .Y (n_1253));
NAND2X1 g77333(.A (n_896), .B (n_303), .Y (n_1252));
INVX8 g82261(.A (n_18266), .Y (n_3886));
INVX2 g80379(.A (n_1739), .Y (n_2368));
INVX1 g80247(.A (n_1251), .Y (n_2251));
NAND2X1 g76992(.A (n_28549), .B (n_377), .Y (n_1248));
INVX1 g77716(.A (n_1284), .Y (n_1246));
NAND2X1 g76492(.A (n_28692), .B (n_753), .Y (n_1993));
INVX1 g77224(.A (n_1242), .Y (n_1243));
NAND2X2 g76879(.A (n_1044), .B (n_207), .Y (n_1534));
INVX2 g80568(.A (n_1241), .Y (n_8928));
NAND2X1 g77695(.A (key[24]), .B (n_25052), .Y (n_1239));
XOR2X1 g76343(.A (n_1236), .B (n_1235), .Y (n_1237));
INVX2 g78227(.A (n_1083), .Y (n_15507));
NAND2X1 g76685(.A (n_29018), .B (n_5799), .Y (n_1233));
NOR2X1 g78200(.A (n_28686), .B (n_14627), .Y (n_15074));
NAND2X1 g76653(.A (w3[20] ), .B (n_3318), .Y (n_1572));
INVX1 g79471(.A (n_1230), .Y (n_2119));
INVX1 g79899(.A (n_1228), .Y (n_1229));
XOR2X1 g76260(.A (n_22569), .B (n_9), .Y (n_1227));
INVX1 g82018(.A (n_19532), .Y (n_19908));
XOR2X1 g76197(.A (n_23241), .B (n_22794), .Y (n_1226));
AND2X1 g76544(.A (n_28645), .B (n_908), .Y (n_2091));
XOR2X1 g76215(.A (n_23352), .B (n_23494), .Y (n_1224));
INVX1 g78034(.A (n_1102), .Y (n_1223));
INVX2 g78690(.A (n_2981), .Y (n_1547));
INVX1 g81196(.A (n_20397), .Y (n_20841));
XOR2X1 g76341(.A (n_1220), .B (n_23261), .Y (n_1221));
INVX1 g79680(.A (n_1956), .Y (n_1616));
INVX1 g78463(.A (n_1053), .Y (n_9003));
XOR2X1 g76344(.A (n_1270), .B (w1[27] ), .Y (n_1217));
NAND2X2 g76678(.A (n_28577), .B (n_849), .Y (n_1736));
INVX4 g81132(.A (n_28167), .Y (n_2001));
INVX1 g77943(.A (n_1212), .Y (n_1707));
INVX1 g77637(.A (n_571), .Y (n_2183));
INVX1 g80619(.A (n_1014), .Y (n_5305));
INVX4 g79322(.A (n_1701), .Y (n_14878));
INVX1 g78213(.A (n_654), .Y (n_2025));
NAND2X1 g77537(.A (rst), .B (n_698), .Y (n_9249));
INVX1 g79445(.A (n_1206), .Y (n_2084));
NOR2X1 g66065(.A (n_1204), .B (n_63), .Y (n_1205));
CLKBUFX1 g81133(.A (n_28167), .Y (n_15610));
INVX1 g81742(.A (n_1972), .Y (n_9682));
NAND2X1 g76831(.A (n_381), .B (n_1201), .Y (n_1771));
NAND2X1 g77164(.A (n_514), .B (n_916), .Y (n_2253));
INVX1 g79748(.A (n_1989), .Y (n_1850));
INVX1 g78255(.A (n_8471), .Y (n_8846));
INVX4 g79447(.A (n_1198), .Y (n_5990));
INVX1 g80579(.A (n_2158), .Y (n_1591));
NOR2X1 g78126(.A (n_11300), .B (n_1196), .Y (n_16553));
INVX1 g78320(.A (sa13[1] ), .Y (n_20457));
NOR2X1 g78145(.A (n_386), .B (n_271), .Y (n_5149));
INVX1 g78661(.A (n_16787), .Y (n_3612));
NAND2X1 g76838(.A (n_29062), .B (n_829), .Y (n_1768));
INVX1 g82069(.A (n_4357), .Y (n_1558));
INVX2 g77973(.A (n_28018), .Y (n_2092));
INVX1 g77111(.A (n_1191), .Y (n_2049));
INVX2 g81629(.A (n_1268), .Y (n_8090));
BUFX3 g80952(.A (n_14624), .Y (n_15568));
NAND2X1 g77036(.A (n_5306), .B (n_9057), .Y (n_1777));
INVX1 g79439(.A (n_6252), .Y (n_1941));
INVX1 g81532(.A (n_673), .Y (n_11277));
INVX1 g81987(.A (n_1186), .Y (n_2035));
NAND2X1 g76743(.A (n_27984), .B (n_1185), .Y (n_1818));
INVX1 g81274(.A (n_2124), .Y (n_2164));
INVX2 g81880(.A (n_2343), .Y (n_2708));
INVX1 g79887(.A (n_21242), .Y (n_16358));
INVX1 g81728(.A (n_27202), .Y (n_1745));
NAND2X1 g77189(.A (n_731), .B (n_296), .Y (n_1897));
INVX1 g76660(.A (n_646), .Y (n_2089));
INVX1 g77455(.A (n_7453), .Y (n_4367));
INVX1 g82218(.A (n_27718), .Y (n_20579));
INVX1 g77861(.A (n_755), .Y (n_6620));
INVX4 g80706(.A (n_932), .Y (n_5413));
BUFX3 g79436(.A (n_3534), .Y (n_10031));
NAND2X1 g76914(.A (n_964), .B (n_3038), .Y (n_1177));
AND2X1 g67826(.A (n_1448), .B (n_1176), .Y (n_6301));
INVX1 g81837(.A (n_1493), .Y (n_6497));
INVX1 g77649(.A (n_1365), .Y (n_10160));
NOR2X1 g76502(.A (w3[28] ), .B (n_2779), .Y (n_1173));
INVX2 g81113(.A (n_27407), .Y (n_6877));
INVX1 g77573(.A (n_8437), .Y (n_11816));
INVX1 g78099(.A (n_1166), .Y (n_1789));
XOR2X1 g76126(.A (n_1164), .B (n_1163), .Y (n_1165));
INVX4 g78739(.A (n_27100), .Y (n_15712));
XOR2X1 g76342(.A (n_22546), .B (n_23191), .Y (n_1158));
INVX1 g80809(.A (n_1157), .Y (n_2152));
INVX1 g78205(.A (n_1155), .Y (n_1772));
NOR2X1 g77824(.A (n_28167), .B (n_1147), .Y (n_13872));
AND2X1 g78207(.A (n_5983), .B (n_1942), .Y (n_9899));
INVX8 g81021(.A (n_27133), .Y (n_1756));
XOR2X1 g76170(.A (n_2009), .B (n_255), .Y (n_1140));
INVX1 g78500(.A (n_1138), .Y (n_2004));
XOR2X1 g76255(.A (n_23309), .B (n_23397), .Y (n_1135));
INVX1 g76826(.A (n_1134), .Y (n_2484));
INVX4 g80365(.A (n_583), .Y (n_12169));
INVX2 g79002(.A (n_1132), .Y (n_15166));
INVX1 g80014(.A (n_1711), .Y (n_1129));
XOR2X1 g76253(.A (n_23047), .B (n_23184), .Y (n_1127));
NAND2X1 g77024(.A (n_15674), .B (w3[17] ), .Y (n_1530));
INVX2 g81602(.A (n_1628), .Y (n_1750));
INVX1 g77511(.A (n_1125), .Y (n_2541));
AND2X1 g77845(.A (n_379), .B (n_1332), .Y (n_2988));
INVX2 g80299(.A (n_819), .Y (n_9264));
INVX1 g80101(.A (n_214), .Y (n_2319));
INVX1 g80094(.A (n_1120), .Y (n_2191));
INVX4 g78393(.A (n_1118), .Y (n_1484));
INVX1 g80877(.A (n_20677), .Y (n_21487));
INVX2 g82443(.A (n_183), .Y (n_9357));
INVX1 g77843(.A (n_7832), .Y (n_2215));
INVX2 g80958(.A (n_1113), .Y (n_15411));
XOR2X1 g76171(.A (n_23001), .B (n_23096), .Y (n_1109));
NOR2X1 g77838(.A (n_11354), .B (n_6868), .Y (n_12134));
INVX2 g78883(.A (n_1106), .Y (n_1601));
XOR2X1 g76166(.A (n_1103), .B (n_1632), .Y (n_1104));
INVX1 g81638(.A (n_1110), .Y (n_6055));
NAND2X2 g77369(.A (n_1015), .B (n_26382), .Y (n_1098));
INVX2 g78908(.A (n_4522), .Y (n_2187));
CLKBUFX1 g78088(.A (n_9276), .Y (n_16973));
XOR2X1 g76098(.A (n_22829), .B (n_22787), .Y (n_1088));
CLKBUFX1 g78909(.A (n_4522), .Y (n_4846));
XOR2X1 g76117(.A (n_141), .B (n_2437), .Y (n_1087));
INVX1 g78073(.A (n_1085), .Y (n_10607));
NOR2X1 g77632(.A (n_1081), .B (n_28357), .Y (n_1082));
CLKBUFX1 g79898(.A (n_1228), .Y (n_3566));
AND2X1 g77424(.A (n_1080), .B (n_1079), .Y (n_2209));
INVX4 g80849(.A (n_19651), .Y (n_19791));
NAND2X1 g77182(.A (n_370), .B (n_827), .Y (n_1075));
XOR2X1 g76115(.A (n_22794), .B (n_22833), .Y (n_1074));
XOR2X1 g76292(.A (n_1072), .B (n_1555), .Y (n_1073));
INVX2 g80399(.A (n_1069), .Y (n_5203));
NAND2X1 g77193(.A (n_1065), .B (n_27674), .Y (n_1998));
NOR2X1 g76934(.A (n_441), .B (n_27434), .Y (n_2456));
NAND2X2 g76485(.A (n_1065), .B (n_527), .Y (n_1743));
OR2X1 g77373(.A (n_607), .B (n_827), .Y (n_2214));
NAND2X2 g76756(.A (n_540), .B (n_899), .Y (n_1064));
INVX1 g77950(.A (n_1063), .Y (n_11810));
INVX1 g81940(.A (n_10599), .Y (n_1642));
NAND2X1 g76736(.A (n_17411), .B (n_668), .Y (n_2052));
NAND2X2 g77703(.A (n_1050), .B (n_959), .Y (n_1051));
INVX1 g78900(.A (n_1046), .Y (n_3014));
NAND2X2 g77610(.A (n_1044), .B (n_1043), .Y (n_1742));
XOR2X1 g76285(.A (n_1040), .B (n_1039), .Y (n_1041));
XOR2X1 g76183(.A (n_1018), .B (n_23399), .Y (n_1038));
INVX1 g78628(.A (n_2007), .Y (n_7734));
INVX2 g79015(.A (n_1456), .Y (n_1037));
INVX1 g80580(.A (n_2158), .Y (n_1036));
INVX2 g78285(.A (n_529), .Y (n_2738));
NAND2X1 g76808(.A (n_981), .B (n_28480), .Y (n_2113));
INVX1 g81121(.A (n_13804), .Y (n_1576));
XOR2X1 g76264(.A (n_1019), .B (n_1018), .Y (n_1020));
INVX2 g81648(.A (n_1339), .Y (n_7728));
INVX1 g77596(.A (n_1016), .Y (n_29316));
NAND2X1 g77606(.A (n_1014), .B (n_3038), .Y (n_2109));
INVX1 g77737(.A (n_8418), .Y (n_19361));
XOR2X1 g76245(.A (n_194), .B (w1[5] ), .Y (n_1012));
INVX2 g82184(.A (n_1010), .Y (n_7559));
NAND2X1 g76498(.A (n_801), .B (n_454), .Y (n_1538));
INVX2 g81252(.A (n_1008), .Y (n_1991));
INVX1 g80126(.A (n_6946), .Y (n_1651));
XOR2X1 g76261(.A (n_1005), .B (n_1004), .Y (n_1006));
INVX1 g77622(.A (n_1003), .Y (n_14113));
NAND2X1 g76711(.A (n_28548), .B (n_434), .Y (n_1002));
INVX1 g77764(.A (n_773), .Y (n_2691));
INVX1 g77403(.A (n_999), .Y (n_2259));
INVX1 g80012(.A (n_2492), .Y (n_997));
CLKBUFX3 g79771(.A (n_26486), .Y (n_4848));
XOR2X1 g76350(.A (text_in_r[57] ), .B (n_9), .Y (n_995));
XOR2X1 g76133(.A (n_23191), .B (n_23053), .Y (n_993));
INVX2 g80524(.A (n_3955), .Y (n_5151));
NAND2X1 g77854(.A (key[29]), .B (n_25052), .Y (n_989));
INVX1 g79335(.A (n_9388), .Y (n_2063));
INVX2 g77991(.A (n_5704), .Y (n_12568));
AND2X1 g77493(.A (n_9527), .B (n_3599), .Y (n_9755));
NAND2X1 g78222(.A (n_28549), .B (n_434), .Y (n_988));
AOI21X1 g75895(.A0 (dcnt[0] ), .A1 (dcnt[1] ), .B0 (n_1448), .Y(n_986));
OR2X1 g77394(.A (n_379), .B (n_2779), .Y (n_6694));
NAND2X1 g76969(.A (n_673), .B (n_9118), .Y (n_3021));
XOR2X1 g76224(.A (n_2174), .B (n_982), .Y (n_983));
INVX1 g78049(.A (n_732), .Y (n_2048));
XOR2X1 g76176(.A (w2[0] ), .B (n_1958), .Y (n_980));
XOR2X1 g76275(.A (n_22831), .B (n_22789), .Y (n_977));
INVX1 g80139(.A (n_1600), .Y (n_1641));
NOR2X1 g76631(.A (n_706), .B (n_7593), .Y (n_976));
XOR2X1 g76147(.A (n_245), .B (n_1960), .Y (n_974));
XOR2X1 g76099(.A (n_97), .B (n_1769), .Y (n_972));
NAND2X1 g77642(.A (n_28642), .B (n_12019), .Y (n_9999));
INVX1 g77443(.A (n_883), .Y (n_1874));
CLKBUFX3 g79031(.A (n_3511), .Y (n_16204));
INVX1 g79154(.A (n_969), .Y (n_9417));
NOR2X1 g76889(.A (n_968), .B (n_218), .Y (n_2111));
INVX1 g78089(.A (n_9276), .Y (n_967));
INVX1 g76595(.A (n_1609), .Y (n_1835));
OR2X1 g77980(.A (n_17411), .B (n_9118), .Y (n_12850));
NAND2X1 g76977(.A (n_213), .B (n_2779), .Y (n_1806));
NAND2X1 g77241(.A (n_474), .B (n_964), .Y (n_2062));
INVX2 g77479(.A (n_671), .Y (n_2017));
NAND2X1 g76431(.A (n_709), .B (n_959), .Y (n_960));
INVX2 g80182(.A (n_2099), .Y (n_4837));
NAND2X1 g76558(.A (n_4861), .B (n_3724), .Y (n_8099));
INVX1 g81528(.A (n_673), .Y (n_19896));
INVX4 g80068(.A (n_751), .Y (n_11307));
INVX2 g80393(.A (n_735), .Y (n_2656));
INVX1 g81651(.A (n_4865), .Y (n_1339));
INVX8 g79833(.A (n_638), .Y (n_11261));
INVX2 g80639(.A (n_3538), .Y (n_2681));
INVX2 g78481(.A (n_1147), .Y (n_975));
INVX1 g81603(.A (n_1050), .Y (n_1628));
INVX2 g81764(.A (n_581), .Y (n_6133));
INVX1 g78885(.A (n_1260), .Y (n_1106));
INVX4 g80702(.A (n_932), .Y (n_5660));
OR2X1 g77993(.A (n_14624), .B (n_28037), .Y (n_5704));
INVX2 g79653(.A (n_2211), .Y (n_931));
NOR2X1 g77958(.A (n_464), .B (n_68), .Y (n_1312));
INVX2 g82491(.A (n_744), .Y (n_926));
INVX2 g79480(.A (n_870), .Y (n_920));
NOR2X1 g78039(.A (n_919), .B (n_912), .Y (n_1102));
NOR2X1 g77667(.A (n_160), .B (n_916), .Y (n_917));
INVX1 g80504(.A (n_4611), .Y (n_1423));
INVX1 g78440(.A (n_807), .Y (n_1315));
NOR2X1 g78090(.A (n_8708), .B (n_271), .Y (n_9276));
NAND2X1 g78021(.A (n_912), .B (n_919), .Y (n_913));
INVX2 g80694(.A (n_26879), .Y (n_3234));
INVX2 g82087(.A (n_1539), .Y (n_3284));
INVX1 g81760(.A (n_1678), .Y (n_23255));
OR2X1 g77633(.A (n_5422), .B (n_152), .Y (n_3640));
INVX1 g80386(.A (n_631), .Y (n_3840));
INVX1 g79773(.A (n_26485), .Y (n_4586));
INVX8 g81437(.A (n_20010), .Y (n_16466));
INVX1 g81975(.A (n_669), .Y (n_8742));
INVX4 g80856(.A (n_688), .Y (n_18205));
INVX4 g80106(.A (n_27641), .Y (n_6021));
INVX1 g81821(.A (n_902), .Y (n_12979));
INVX1 g81064(.A (n_1674), .Y (n_23599));
NOR2X1 g77985(.A (n_900), .B (n_899), .Y (n_901));
INVX4 g81146(.A (n_399), .Y (n_10100));
INVX8 g82537(.A (n_27747), .Y (n_9084));
INVX8 g78449(.A (n_897), .Y (n_6185));
INVX2 g82514(.A (n_1390), .Y (n_3108));
NOR2X1 g77944(.A (n_896), .B (n_15), .Y (n_1212));
XOR2X1 g76309(.A (text_in_r[32] ), .B (w2[0] ), .Y (n_894));
INVX1 g81958(.A (n_770), .Y (n_6052));
INVX4 g81783(.A (n_902), .Y (n_7331));
NOR2X1 g77439(.A (n_561), .B (n_176), .Y (n_962));
NOR2X1 g77844(.A (n_22), .B (n_9057), .Y (n_7832));
CLKBUFX3 g79455(.A (n_470), .Y (n_1198));
INVX1 g81548(.A (n_21275), .Y (n_20574));
INVX8 g79046(.A (n_563), .Y (n_14055));
XOR2X1 g76232(.A (text_in_r[96] ), .B (w0[0] ), .Y (n_884));
NOR2X1 g77444(.A (n_228), .B (n_2), .Y (n_883));
INVX2 g81738(.A (n_578), .Y (n_6977));
INVX1 g82334(.A (n_933), .Y (n_19319));
INVX1 g79902(.A (n_26891), .Y (n_872));
NOR2X1 g77909(.A (n_26382), .B (n_251), .Y (n_871));
INVX2 g79487(.A (n_870), .Y (n_1483));
NAND2X1 g78275(.A (n_18205), .B (n_29297), .Y (n_6527));
INVX1 g79244(.A (n_867), .Y (n_868));
INVX2 g79687(.A (n_494), .Y (n_9486));
INVX1 g78434(.A (n_509), .Y (n_3695));
NAND2X1 g77624(.A (n_18237), .B (n_2318), .Y (n_1003));
INVX1 g81073(.A (n_19940), .Y (n_20661));
INVX4 g78983(.A (n_16978), .Y (n_4582));
INVX1 g80621(.A (n_1014), .Y (n_853));
INVX4 g80122(.A (n_28154), .Y (n_4364));
NAND2X2 g77938(.A (n_849), .B (n_28568), .Y (n_850));
INVX1 g81197(.A (sa31[1] ), .Y (n_20397));
INVX1 g81076(.A (n_19924), .Y (n_20986));
NOR2X1 g78206(.A (n_772), .B (n_622), .Y (n_1155));
INVX2 g80850(.A (n_18205), .Y (n_19651));
INVX2 g79707(.A (n_290), .Y (n_13326));
CLKBUFX3 g82192(.A (n_26874), .Y (n_1373));
INVX2 g79297(.A (n_718), .Y (n_8878));
INVX1 g81734(.A (n_4598), .Y (n_1124));
INVX2 g81756(.A (n_834), .Y (n_1427));
NOR2X1 g77533(.A (n_1285), .B (n_218), .Y (n_833));
NAND2X1 g77112(.A (w3[14] ), .B (n_664), .Y (n_1191));
CLKBUFX2 g78679(.A (n_2921), .Y (n_17864));
INVX2 g81776(.A (n_3807), .Y (n_1347));
INVX1 g78735(.A (n_828), .Y (n_14592));
OR2X1 g77409(.A (n_730), .B (n_827), .Y (n_1447));
INVX1 g79611(.A (sa10[0] ), .Y (n_825));
INVX4 g79381(.A (n_829), .Y (n_4689));
INVX2 g80789(.A (n_821), .Y (n_4300));
CLKBUFX3 g80380(.A (n_818), .Y (n_1739));
INVX4 g82392(.A (n_27336), .Y (n_15776));
INVX1 g82239(.A (n_27718), .Y (n_20068));
INVX2 g78933(.A (n_783), .Y (n_4522));
INVX4 g81788(.A (n_902), .Y (n_2260));
INVX1 g82447(.A (n_9624), .Y (n_22881));
INVX4 g78792(.A (n_791), .Y (n_3820));
NAND2X1 g77556(.A (n_14624), .B (n_28037), .Y (n_7899));
INVX2 g81110(.A (n_27407), .Y (n_13318));
INVX4 g79864(.A (n_106), .Y (n_1000));
INVX2 g78437(.A (n_807), .Y (n_2483));
INVX1 g79813(.A (sa31[3] ), .Y (n_7512));
INVX4 g81292(.A (n_804), .Y (n_21314));
INVX1 g80359(.A (n_583), .Y (n_7777));
NOR2X1 g78254(.A (n_849), .B (n_28568), .Y (n_803));
CLKBUFX1 g81275(.A (n_3251), .Y (n_2124));
INVX2 g79803(.A (n_547), .Y (n_8968));
INVX2 g81278(.A (n_2069), .Y (n_1540));
NAND2X1 g77380(.A (n_801), .B (n_896), .Y (n_802));
INVX2 g79749(.A (n_28158), .Y (n_1989));
INVX1 g80269(.A (n_6790), .Y (n_1153));
INVX1 g78372(.A (sa30[1] ), .Y (n_20386));
INVX1 g80695(.A (n_26879), .Y (n_4934));
INVX1 g80260(.A (n_1970), .Y (n_23169));
INVX4 g80786(.A (n_795), .Y (n_8945));
INVX4 g81423(.A (n_13083), .Y (n_19445));
NAND2X1 g76526(.A (n_380), .B (n_1431), .Y (n_1324));
INVX1 g79243(.A (n_867), .Y (n_3081));
CLKBUFX1 g81641(.A (n_3632), .Y (n_6419));
INVX1 g78367(.A (n_20198), .Y (n_15766));
INVX4 g79360(.A (n_789), .Y (n_9368));
INVX1 g82141(.A (n_788), .Y (n_21133));
INVX1 g81937(.A (n_408), .Y (n_1946));
INVX2 g79440(.A (n_532), .Y (n_6252));
INVX1 g80889(.A (n_778), .Y (n_17933));
INVX4 g81877(.A (n_569), .Y (n_2343));
INVX1 g80817(.A (n_775), .Y (n_1157));
NAND2X1 g77765(.A (n_772), .B (n_622), .Y (n_773));
NAND2X2 g77692(.A (n_26888), .B (n_767), .Y (n_1307));
INVX4 g80926(.A (n_18456), .Y (n_11489));
NOR2X1 g77798(.A (n_26888), .B (n_767), .Y (n_1384));
INVX1 g81674(.A (n_759), .Y (n_6988));
NOR2X1 g77771(.A (n_849), .B (n_28482), .Y (n_1294));
NOR2X1 g77862(.A (n_4598), .B (n_280), .Y (n_755));
INVX4 g78753(.A (n_27111), .Y (n_9410));
INVX2 g80581(.A (n_1081), .Y (n_2158));
INVX2 g80510(.A (n_3955), .Y (n_4882));
NOR2X1 g78269(.A (n_748), .B (n_28786), .Y (n_749));
INVX8 g82532(.A (n_27747), .Y (n_4709));
INVX2 g82490(.A (n_744), .Y (n_1634));
INVX2 g82333(.A (n_933), .Y (n_20153));
INVX1 g79600(.A (n_624), .Y (n_13571));
INVX4 g79573(.A (n_624), .Y (n_12298));
OR2X1 g77951(.A (n_26041), .B (n_4173), .Y (n_1063));
CLKBUFX3 g80400(.A (n_735), .Y (n_1069));
NOR2X1 g78050(.A (n_731), .B (n_730), .Y (n_732));
AND2X1 g77544(.A (n_3338), .B (n_352), .Y (n_1416));
INVX1 g79937(.A (n_24548), .Y (n_3721));
NAND2X1 g76827(.A (n_440), .B (n_295), .Y (n_1134));
INVX4 g78665(.A (sa13[2] ), .Y (n_16787));
INVX1 g80083(.A (n_719), .Y (n_720));
CLKBUFX3 g80799(.A (n_1015), .Y (n_1353));
INVX8 g79144(.A (n_713), .Y (n_8997));
INVX1 g79156(.A (n_2810), .Y (n_969));
INVX8 g81919(.A (n_481), .Y (n_6005));
INVX2 g81817(.A (n_902), .Y (n_4898));
INVX4 g79020(.A (n_714), .Y (n_1456));
INVX2 g80013(.A (n_790), .Y (n_2492));
INVX8 g79853(.A (n_1000), .Y (n_15894));
INVX2 g81606(.A (n_709), .Y (n_1395));
INVX1 g79681(.A (n_964), .Y (n_1956));
INVX2 g82465(.A (n_706), .Y (n_7607));
INVX2 g78438(.A (n_807), .Y (n_3296));
INVX1 g79900(.A (n_26891), .Y (n_1228));
INVX4 g81123(.A (sa10[2] ), .Y (n_13804));
INVX4 g82196(.A (n_26874), .Y (n_11253));
INVX8 g80749(.A (n_441), .Y (n_6462));
INVX4 g80772(.A (n_795), .Y (n_6997));
INVX8 g81695(.A (n_5306), .Y (n_3301));
INVX1 g80569(.A (n_5085), .Y (n_1241));
INVX2 g78934(.A (n_783), .Y (n_6043));
INVX1 g79249(.A (n_23053), .Y (n_2412));
INVX4 g78822(.A (n_1295), .Y (n_20325));
INVX1 g80963(.A (n_27688), .Y (n_1113));
INVX1 g78929(.A (n_783), .Y (n_677));
INVX1 g82094(.A (n_3464), .Y (n_1213));
CLKBUFX1 g82186(.A (n_26874), .Y (n_1010));
INVX1 g81524(.A (n_673), .Y (n_1057));
NOR2X1 g77480(.A (n_109), .B (n_1043), .Y (n_671));
NAND2X1 g77789(.A (n_18), .B (n_26), .Y (n_1263));
INVX1 g81645(.A (n_2487), .Y (n_1316));
INVX1 g82100(.A (n_1065), .Y (n_2236));
OR2X1 g78229(.A (n_12827), .B (n_1376), .Y (n_1083));
NOR2X1 g77688(.A (n_14), .B (n_664), .Y (n_665));
INVX4 g80525(.A (n_5422), .Y (n_3955));
INVX1 g80464(.A (n_267), .Y (n_13606));
INVX1 g81988(.A (n_27668), .Y (n_1186));
INVX2 g80074(.A (n_508), .Y (n_7658));
INVX1 g78572(.A (n_482), .Y (n_5416));
NOR2X1 g78214(.A (n_896), .B (n_801), .Y (n_654));
INVX1 g81868(.A (n_26903), .Y (n_20648));
INVX1 g81995(.A (n_22833), .Y (n_2587));
INVX1 g81640(.A (n_3632), .Y (n_1110));
INVX2 g79502(.A (n_6431), .Y (n_9467));
INVX1 g81842(.A (n_1385), .Y (n_2417));
NAND2X1 g76661(.A (n_160), .B (w3[23] ), .Y (n_646));
NOR2X1 g78100(.A (n_343), .B (n_26382), .Y (n_1166));
CLKBUFX3 g78921(.A (n_783), .Y (n_1358));
NAND2X2 g77456(.A (n_636), .B (n_4861), .Y (n_7453));
NOR2X1 g78262(.A (n_26597), .B (n_89), .Y (n_29122));
INVX2 g79786(.A (n_656), .Y (n_7266));
NOR2X1 g78095(.A (n_1185), .B (n_29167), .Y (n_632));
INVX4 g80384(.A (n_631), .Y (n_2383));
INVX1 g82227(.A (n_20758), .Y (n_21447));
INVX1 g78887(.A (n_629), .Y (n_630));
AND2X1 g77782(.A (n_627), .B (n_28786), .Y (n_1370));
INVX2 g82458(.A (n_4721), .Y (n_1340));
NOR2X1 g77517(.A (n_622), .B (n_1079), .Y (n_623));
NOR2X1 g77404(.A (n_3348), .B (n_352), .Y (n_999));
INVX4 g79767(.A (n_27369), .Y (n_27370));
INVX1 g80801(.A (n_612), .Y (n_2070));
OR2X1 g78163(.A (n_18237), .B (n_2318), .Y (n_12849));
INVX1 g78901(.A (n_607), .Y (n_1046));
XOR2X1 g76185(.A (w2[0] ), .B (w0[0] ), .Y (n_606));
INVX1 g81655(.A (n_28133), .Y (n_7438));
INVX8 g82365(.A (n_27336), .Y (n_17912));
INVX2 g80381(.A (n_818), .Y (n_1823));
INVX2 g78637(.A (n_26394), .Y (n_1569));
INVX1 g78712(.A (n_14630), .Y (n_1368));
INVX4 g78459(.A (n_1147), .Y (n_1053));
INVX4 g81669(.A (n_881), .Y (n_596));
INVX4 g80282(.A (n_819), .Y (n_8637));
INVX1 g81945(.A (n_770), .Y (n_11215));
INVX1 g81398(.A (n_591), .Y (n_11385));
INVX2 g80965(.A (n_587), .Y (n_8435));
NOR2X1 g77293(.A (w3[20] ), .B (n_3318), .Y (n_584));
INVX8 g80347(.A (n_583), .Y (n_7410));
INVX2 g81855(.A (n_875), .Y (n_1397));
INVX2 g79412(.A (n_1626), .Y (n_9474));
INVX1 g79472(.A (n_968), .Y (n_1230));
INVX1 g80248(.A (n_1332), .Y (n_1251));
INVX1 g80937(.A (sa30[2] ), .Y (n_12910));
INVX2 g81768(.A (n_581), .Y (n_2655));
INVX4 g81253(.A (n_19934), .Y (n_1008));
NOR2X1 g77778(.A (n_199), .B (n_959), .Y (n_579));
INVX2 g82305(.A (n_575), .Y (n_1551));
INVX1 g78593(.A (n_7182), .Y (n_2838));
NOR2X1 g77638(.A (n_801), .B (n_315), .Y (n_571));
INVX1 g80082(.A (n_719), .Y (n_1244));
NAND2X1 g77739(.A (n_4861), .B (n_27344), .Y (n_8418));
INVX4 g79884(.A (n_908), .Y (n_21242));
OR2X1 g77574(.A (n_28686), .B (n_4391), .Y (n_8437));
NAND2X2 g77528(.A (n_561), .B (n_176), .Y (n_1430));
INVX1 g78640(.A (n_26394), .Y (n_25691));
INVX4 g79736(.A (n_557), .Y (n_8918));
INVX1 g78311(.A (w0[18] ), .Y (n_2769));
INVX1 g81822(.A (n_902), .Y (n_6007));
INVX1 g79008(.A (n_11354), .Y (n_1132));
OR2X1 g77503(.A (n_4861), .B (n_27344), .Y (n_1363));
INVX1 g80148(.A (sa11[1] ), .Y (n_19981));
INVX2 g80718(.A (n_4113), .Y (n_1238));
INVX4 g80532(.A (n_544), .Y (n_8974));
INVX2 g80127(.A (n_28154), .Y (n_6946));
INVX1 g78396(.A (n_540), .Y (n_541));
INVX1 g79666(.A (n_1431), .Y (n_1142));
NOR2X1 g77462(.A (n_285), .B (n_537), .Y (n_538));
INVX4 g79299(.A (n_718), .Y (n_6226));
INVX1 g80804(.A (n_1934), .Y (n_22704));
INVX1 g82527(.A (n_525), .Y (n_1647));
INVX1 g79437(.A (n_532), .Y (n_3534));
INVX1 g79323(.A (n_430), .Y (n_1701));
INVX4 g80238(.A (n_1080), .Y (n_1258));
INVX2 g81584(.A (n_530), .Y (n_7537));
NAND2X2 g78286(.A (n_528), .B (n_527), .Y (n_529));
INVX1 g80723(.A (n_393), .Y (n_7366));
INVX1 g82019(.A (n_20213), .Y (n_19532));
INVX4 g81806(.A (n_902), .Y (n_5854));
INVX1 g79032(.A (n_519), .Y (n_3511));
INVX1 g81779(.A (n_264), .Y (n_6279));
AND2X1 g77651(.A (n_4490), .B (n_4391), .Y (n_1365));
INVX1 g78435(.A (n_509), .Y (n_2646));
INVX2 g78395(.A (n_540), .Y (n_1118));
INVX4 g79693(.A (sa32[2] ), .Y (n_8708));
INVX2 g79411(.A (n_1626), .Y (n_5817));
INVX4 g80831(.A (n_503), .Y (n_12986));
INVX2 g80015(.A (n_790), .Y (n_1711));
INVX1 g80459(.A (n_267), .Y (n_11603));
INVX1 g80168(.A (n_20767), .Y (n_21398));
INVX4 g79591(.A (n_624), .Y (n_5329));
INVX2 g80394(.A (n_735), .Y (n_1460));
INVX2 g79774(.A (n_26485), .Y (n_3704));
INVX2 g80018(.A (n_790), .Y (n_493));
INVX1 g81778(.A (n_264), .Y (n_6191));
INVX2 g78576(.A (n_213), .Y (n_490));
INVX4 g80541(.A (n_753), .Y (n_9942));
INVX4 g78841(.A (n_485), .Y (n_14589));
INVX1 g80140(.A (n_514), .Y (n_1600));
INVX4 g81918(.A (n_481), .Y (n_7201));
INVX2 g80206(.A (n_479), .Y (n_1266));
INVX2 g81722(.A (n_674), .Y (n_4627));
INVX1 g81943(.A (n_770), .Y (n_3756));
NAND2X1 g77512(.A (n_474), .B (n_664), .Y (n_1125));
AND2X1 g78074(.A (n_300), .B (n_1942), .Y (n_1085));
NAND2X1 g77098(.A (n_437), .B (w3[21] ), .Y (n_473));
INVX4 g79805(.A (n_547), .Y (n_10495));
INVX1 g79446(.A (n_470), .Y (n_1206));
INVX1 g80095(.A (n_1292), .Y (n_1120));
INVX1 g80662(.A (n_469), .Y (n_2044));
NOR2X1 g78186(.A (n_165), .B (n_3318), .Y (n_16976));
INVX1 g81189(.A (sa31[1] ), .Y (n_15371));
NOR2X1 g77602(.A (n_464), .B (n_527), .Y (n_1016));
INVX1 g79474(.A (n_462), .Y (n_463));
NOR2X1 g77468(.A (n_27983), .B (n_305), .Y (n_459));
INVX2 g80935(.A (sa30[2] ), .Y (n_17567));
NOR2X1 g77717(.A (n_457), .B (n_2943), .Y (n_1284));
NAND2X1 g78027(.A (n_160), .B (n_916), .Y (n_1313));
INVX4 g80645(.A (sa21[1] ), .Y (n_21396));
INVX2 g78692(.A (n_9982), .Y (n_2981));
INVX1 g81743(.A (n_454), .Y (n_1972));
INVX4 g80480(.A (n_1667), .Y (n_18369));
INVX1 g78731(.A (n_828), .Y (n_13815));
NOR2X1 g78007(.A (n_27133), .B (n_28375), .Y (n_11850));
INVX1 g82139(.A (sa23[1] ), .Y (n_19372));
CLKBUFX3 g81002(.A (sa01[2] ), .Y (n_1310));
INVX2 g79592(.A (n_624), .Y (n_9917));
INVX1 g78629(.A (n_3001), .Y (n_2007));
INVX1 g80157(.A (n_20332), .Y (n_20564));
INVX8 g78810(.A (n_1295), .Y (n_18320));
NAND2X1 g76596(.A (n_440), .B (n_827), .Y (n_1609));
INVX4 g82357(.A (n_3724), .Y (n_1424));
NOR2X1 g77414(.A (n_437), .B (n_2462), .Y (n_1325));
INVX1 g81724(.A (sa10[4] ), .Y (n_4804));
NOR2X1 g77392(.A (n_434), .B (n_28464), .Y (n_435));
INVX2 g79336(.A (n_430), .Y (n_9388));
INVX1 g79023(.A (n_2993), .Y (n_28312));
OR2X1 g78264(.A (n_4916), .B (n_3318), .Y (n_6609));
INVX1 g81838(.A (n_981), .Y (n_1493));
INVX4 g81552(.A (sa22[1] ), .Y (n_21275));
NAND2X1 g78257(.A (n_29065), .B (n_27434), .Y (n_8471));
INVX1 g80902(.A (sa10[1] ), .Y (n_21108));
AND2X1 g78102(.A (n_26041), .B (n_4173), .Y (n_6941));
INVX8 g80839(.A (n_503), .Y (n_17260));
INVX1 g82145(.A (n_788), .Y (n_21442));
NAND2X1 g78107(.A (n_731), .B (n_827), .Y (n_7411));
NAND2X1 g77229(.A (n_26597), .B (sa33[6] ), .Y (n_1242));
INVX1 g81941(.A (n_408), .Y (n_10599));
INVX4 g81505(.A (n_510), .Y (n_17500));
INVX2 g81184(.A (n_400), .Y (n_1336));
INVX8 g81149(.A (n_399), .Y (n_8865));
INVX4 g79060(.A (n_668), .Y (n_11731));
INVX4 g80731(.A (n_393), .Y (n_7563));
INVX4 g81285(.A (sa20[1] ), .Y (n_21055));
INVX1 g79651(.A (n_2211), .Y (n_1508));
INVX1 g81828(.A (n_27192), .Y (n_22203));
CLKBUFX3 g80096(.A (n_801), .Y (n_1292));
INVX8 g80555(.A (n_294), .Y (n_12019));
CLKBUFX1 g80159(.A (n_27481), .Y (n_20332));
INVX4 g81263(.A (sa00[1] ), .Y (n_5131));
INVX1 g78387(.A (n_900), .Y (n_384));
INVX4 g80348(.A (n_9057), .Y (n_583));
CLKBUFX1 g81761(.A (n_23238), .Y (n_1678));
INVX4 g82414(.A (n_2318), .Y (n_826));
INVX1 g80186(.A (n_380), .Y (n_381));
INVX1 g79918(.A (n_360), .Y (n_672));
INVX1 g78326(.A (n_378), .Y (n_20412));
INVX1 g81646(.A (sa02[4] ), .Y (n_2487));
INVX1 g82308(.A (n_434), .Y (n_377));
CLKBUFX1 g80261(.A (n_22564), .Y (n_1970));
INVX4 g79009(.A (w3[26] ), .Y (n_11354));
INVX1 g81942(.A (n_320), .Y (n_408));
INVX1 g79392(.A (n_362), .Y (n_7325));
INVX1 g80252(.A (n_730), .Y (n_370));
INVX1 g80792(.A (n_5005), .Y (n_821));
INVX2 g78797(.A (n_26393), .Y (n_791));
INVX4 g79047(.A (n_367), .Y (n_563));
INVX1 g79033(.A (n_218), .Y (n_519));
INVX2 g81758(.A (n_899), .Y (n_834));
INVX1 g81677(.A (n_4490), .Y (n_759));
INVX1 g79425(.A (n_362), .Y (n_3599));
INVX4 g79705(.A (n_290), .Y (n_15986));
INVX4 g80640(.A (n_21396), .Y (n_3538));
INVX1 g81597(.A (w3[20] ), .Y (n_4916));
INVX4 g79652(.A (n_26991), .Y (n_2211));
CLKBUFX3 g81276(.A (n_2096), .Y (n_3251));
INVX1 g80406(.A (n_27817), .Y (n_357));
INVX1 g80258(.A (n_1018), .Y (n_684));
INVX1 g79742(.A (n_1308), .Y (n_398));
INVX2 g82493(.A (n_527), .Y (n_744));
INVX2 g78359(.A (n_437), .Y (n_3868));
INVX1 g82117(.A (n_348), .Y (n_2467));
INVX4 g81883(.A (n_26989), .Y (n_569));
INVX1 g80802(.A (n_343), .Y (n_612));
NOR2X1 g77816(.A (dcnt[0] ), .B (dcnt[1] ), .Y (n_1448));
INVX1 g80077(.A (n_919), .Y (n_342));
INVX1 g78508(.A (n_22223), .Y (n_341));
INVX1 g78902(.A (n_440), .Y (n_607));
INVX1 g81565(.A (n_26844), .Y (n_22195));
INVX1 g79789(.A (n_26493), .Y (n_656));
INVX2 g78381(.A (n_129), .Y (n_20198));
INVX2 g79424(.A (n_362), .Y (n_8679));
INVX2 g81502(.A (n_17411), .Y (n_510));
INVX2 g80084(.A (n_919), .Y (n_719));
INVX1 g79877(.A (n_14627), .Y (n_844));
INVX1 g82020(.A (w3[17] ), .Y (n_20213));
INVX1 g79245(.A (n_2943), .Y (n_867));
INVX1 g82565(.A (n_23397), .Y (n_805));
INVX1 g81074(.A (sa33[1] ), .Y (n_19940));
INVX1 g78693(.A (sa13[2] ), .Y (n_9982));
INVX2 g79737(.A (n_1043), .Y (n_557));
INVX2 g82482(.A (n_527), .Y (n_25783));
INVX2 g82515(.A (n_627), .Y (n_1390));
INVX1 g81959(.A (n_320), .Y (n_770));
INVX2 g82089(.A (n_315), .Y (n_1539));
INVX2 g79376(.A (n_6008), .Y (n_829));
INVX1 g80147(.A (n_20729), .Y (n_21188));
INVX4 g78594(.A (n_213), .Y (n_7182));
INVX1 g81071(.A (sa33[1] ), .Y (n_310));
INVX2 g78714(.A (sa01[1] ), .Y (n_14630));
INVX1 g79972(.A (n_360), .Y (n_24915));
INVX1 g81081(.A (n_19475), .Y (n_20518));
INVX1 g78945(.A (n_21687), .Y (n_22418));
INVX1 g82223(.A (sa12[1] ), .Y (n_19834));
INVX1 g81642(.A (sa02[4] ), .Y (n_3632));
INVX1 g82053(.A (n_124), .Y (n_19143));
INVX2 g81185(.A (n_305), .Y (n_400));
CLKBUFX1 g81065(.A (n_23234), .Y (n_1674));
INVX2 g80086(.A (n_801), .Y (n_303));
INVX2 g78397(.A (n_900), .Y (n_540));
CLKBUFX3 g80383(.A (n_208), .Y (n_818));
INVX1 g78842(.A (n_300), .Y (n_485));
INVX1 g80428(.A (n_12788), .Y (n_17444));
INVX1 g80967(.A (n_27688), .Y (n_587));
INVX1 g80250(.A (n_295), .Y (n_296));
INVX4 g80741(.A (n_274), .Y (n_4568));
CLKBUFX3 g79247(.A (n_2943), .Y (n_3067));
INVX1 g80622(.A (w3[14] ), .Y (n_1014));
INVX4 g80736(.A (n_383), .Y (n_393));
INVX2 g79711(.A (n_290), .Y (n_14807));
INVX2 g79181(.A (n_9335), .Y (n_427));
INVX1 g78631(.A (n_27204), .Y (n_288));
INVX1 g79386(.A (n_2779), .Y (n_941));
INVX2 g82358(.A (n_27344), .Y (n_3724));
INVX4 g80765(.A (n_330), .Y (n_441));
INVX1 g79985(.A (n_360), .Y (n_25052));
CLKBUFX3 g80654(.A (n_285), .Y (n_1255));
INVX1 g80663(.A (n_285), .Y (n_469));
INVX2 g80452(.A (n_267), .Y (n_15674));
CLKBUFX3 g80270(.A (n_276), .Y (n_6790));
INVX2 g82306(.A (n_434), .Y (n_575));
INVX1 g81978(.A (n_4173), .Y (n_669));
INVX1 g79904(.A (n_26888), .Y (n_273));
INVX1 g79964(.A (n_360), .Y (n_25126));
INVX1 g79963(.A (n_360), .Y (n_25123));
INVX2 g81585(.A (n_3307), .Y (n_530));
INVX1 g80453(.A (n_267), .Y (n_7158));
INVX1 g79806(.A (n_27365), .Y (n_547));
INVX1 g82471(.A (sa30[4] ), .Y (n_3348));
INVX8 g81456(.A (n_13083), .Y (n_20010));
INVX1 g79262(.A (n_1196), .Y (n_20116));
INVX4 g81777(.A (n_264), .Y (n_3807));
INVX1 g80534(.A (n_4391), .Y (n_544));
INVX4 g80843(.A (n_688), .Y (n_11300));
INVX1 g78852(.A (n_9106), .Y (n_477));
INVX1 g79969(.A (n_360), .Y (n_24599));
INVX4 g79574(.A (n_9819), .Y (n_624));
CLKBUFX1 g82467(.A (n_3348), .Y (n_6012));
INVX4 g80719(.A (n_277), .Y (n_4113));
INVX1 g79625(.A (n_23096), .Y (n_764));
INVX1 g82528(.A (n_27746), .Y (n_525));
INVX4 g82101(.A (n_464), .Y (n_1065));
INVX4 g78939(.A (n_238), .Y (n_783));
INVX1 g80665(.A (n_21708), .Y (n_22377));
INVX1 g79441(.A (n_162), .Y (n_532));
CLKBUFX1 g80249(.A (n_295), .Y (n_1332));
INVX1 g78573(.A (n_379), .Y (n_482));
INVX2 g81280(.A (n_251), .Y (n_2069));
INVX1 g78948(.A (n_22274), .Y (n_22353));
INVX1 g82507(.A (n_250), .Y (n_880));
INVX2 g78491(.A (n_3560), .Y (n_488));
INVX2 g78455(.A (n_280), .Y (n_897));
CLKBUFX1 g82228(.A (sa12[1] ), .Y (n_20758));
INVX1 g81723(.A (n_27197), .Y (n_674));
INVX1 g79475(.A (n_1285), .Y (n_462));
INVX1 g80545(.A (n_11272), .Y (n_753));
INVX4 g80832(.A (n_11300), .Y (n_503));
INVX1 g82072(.A (n_4357), .Y (n_16944));
INVX2 g79172(.A (n_1942), .Y (n_523));
INVX1 g80072(.A (n_3318), .Y (n_751));
BUFX3 g79413(.A (n_362), .Y (n_1626));
INVX8 g80310(.A (n_319), .Y (n_7496));
INVX1 g79157(.A (sa22[3] ), .Y (n_2810));
CLKBUFX3 g78886(.A (n_228), .Y (n_1260));
INVX4 g81992(.A (n_1947), .Y (n_2235));
INVX4 g79641(.A (n_101), .Y (n_6805));
INVX1 g79931(.A (n_360), .Y (n_619));
INVX1 g79945(.A (n_360), .Y (n_698));
INVX1 g81653(.A (sa03[4] ), .Y (n_4961));
INVX1 g79246(.A (n_2943), .Y (n_2150));
INVX1 g82146(.A (n_164), .Y (n_788));
INVX8 g81699(.A (n_3920), .Y (n_5306));
INVX1 g79024(.A (n_218), .Y (n_2993));
INVX2 g81672(.A (n_28141), .Y (n_881));
INVX1 g80103(.A (n_214), .Y (n_862));
INVX8 g79152(.A (n_1942), .Y (n_713));
CLKBUFX1 g81077(.A (sa33[1] ), .Y (n_19924));
INVX2 g79415(.A (n_362), .Y (n_6868));
CLKBUFX1 g82517(.A (n_27746), .Y (n_7485));
INVX1 g80057(.A (n_3318), .Y (n_508));
INVX1 g80570(.A (sa03[3] ), .Y (n_5085));
INVX2 g80387(.A (n_208), .Y (n_631));
INVX1 g79738(.A (n_1043), .Y (n_207));
INVX2 g81922(.A (n_28032), .Y (n_7593));
INVX8 g81824(.A (n_271), .Y (n_902));
INVX2 g80890(.A (n_28172), .Y (n_778));
INVX1 g81652(.A (sa03[4] ), .Y (n_4865));
INVX2 g79491(.A (w3[21] ), .Y (n_3283));
BUFX3 g79581(.A (n_9819), .Y (n_17414));
CLKBUFX3 g81604(.A (n_199), .Y (n_1050));
INVX1 g80506(.A (w3[4] ), .Y (n_4611));
INVX1 g80414(.A (n_196), .Y (n_17423));
INVX2 g80481(.A (n_1512), .Y (n_1667));
INVX1 g78385(.A (n_187), .Y (n_20558));
INVX2 g81293(.A (n_21055), .Y (n_804));
CLKBUFX3 g79062(.A (n_205), .Y (n_668));
INVX8 g82459(.A (n_230), .Y (n_4721));
INVX1 g82011(.A (n_3264), .Y (n_663));
INVX2 g82441(.A (n_183), .Y (n_6219));
INVX1 g78436(.A (n_178), .Y (n_509));
CLKBUFX3 g80880(.A (n_177), .Y (n_20677));
INVX1 g79669(.A (n_176), .Y (n_1201));
INVX4 g81520(.A (n_673), .Y (n_14155));
INVX1 g79974(.A (n_360), .Y (n_1914));
INVX1 g78503(.A (n_1138), .Y (n_22301));
INVX1 g81210(.A (n_171), .Y (n_20587));
CLKBUFX3 g80730(.A (n_383), .Y (n_7636));
INVX1 g80583(.A (n_537), .Y (n_167));
INVX1 g80454(.A (n_267), .Y (n_165));
INVX1 g81558(.A (n_19414), .Y (n_17246));
INVX1 g79962(.A (n_360), .Y (n_24548));
CLKBUFX3 g79457(.A (n_162), .Y (n_5983));
INVX4 g81920(.A (n_352), .Y (n_481));
INVX2 g80142(.A (n_160), .Y (n_514));
CLKBUFX3 g80538(.A (n_4391), .Y (n_7498));
INVX1 g82092(.A (n_1291), .Y (n_1272));
CLKBUFX3 g82086(.A (n_315), .Y (n_2079));
INVX4 g80401(.A (n_27592), .Y (n_735));
INVX2 g81607(.A (n_199), .Y (n_709));
INVX1 g82233(.A (n_20018), .Y (n_20810));
INVX1 g79683(.A (n_664), .Y (n_964));
INVX4 g80301(.A (n_276), .Y (n_819));
INVX1 g57639(.A (n_344), .Y (n_21757));
INVX2 g79337(.A (n_152), .Y (n_430));
INVX1 g79967(.A (n_360), .Y (n_24778));
INVX2 g82510(.A (n_748), .Y (n_25802));
INVX4 g82435(.A (n_183), .Y (n_7598));
INVX2 g81839(.A (n_849), .Y (n_981));
CLKBUFX3 g79347(.A (n_135), .Y (n_5799));
INVX1 g81740(.A (n_5381), .Y (n_578));
CLKBUFX3 g82095(.A (n_1291), .Y (n_3464));
INVX1 g79975(.A (n_360), .Y (n_1890));
INVX1 g82031(.A (n_3264), .Y (n_15482));
INVX1 g79645(.A (n_4825), .Y (n_1389));
INVX2 g80709(.A (n_26885), .Y (n_932));
INVX1 g81067(.A (sa33[1] ), .Y (n_20517));
CLKBUFX3 g78630(.A (n_27204), .Y (n_3001));
INVX1 g81270(.A (n_2096), .Y (n_1568));
INVX1 g79362(.A (n_135), .Y (n_789));
INVX4 g79488(.A (n_772), .Y (n_870));
INVX4 g79021(.A (n_767), .Y (n_714));
INVX2 g81744(.A (n_896), .Y (n_454));
INVX1 g57365(.A (n_209), .Y (n_21938));
INVX8 g78830(.A (n_263), .Y (n_1295));
INVX4 g79844(.A (n_18237), .Y (n_638));
INVX1 g82466(.A (n_3348), .Y (n_706));
CLKBUFX3 g79233(.A (n_27983), .Y (n_1302));
NOR2X1 g77557(.A (dcnt[2] ), .B (dcnt[3] ), .Y (n_1176));
INVX1 g79968(.A (n_360), .Y (n_24937));
INVX1 g79958(.A (n_360), .Y (n_600));
INVX1 g79456(.A (n_162), .Y (n_470));
INVX8 g81151(.A (n_4861), .Y (n_399));
INVX2 g81769(.A (n_386), .Y (n_581));
INVX1 g79473(.A (n_1285), .Y (n_968));
INVX1 g82061(.A (n_124), .Y (n_20577));
INVX2 g80185(.A (n_380), .Y (n_2099));
INVX1 g81085(.A (n_20157), .Y (n_20041));
CLKBUFX1 g80805(.A (n_6401), .Y (n_1934));
CLKBUFX3 g79744(.A (n_28151), .Y (n_1305));
INVX4 g80498(.A (n_9342), .Y (n_19310));
INVX8 g81372(.A (n_12827), .Y (n_20406));
INVX1 g78342(.A (n_27449), .Y (n_487));
INVX4 g80787(.A (n_10315), .Y (n_795));
INVX1 g79298(.A (n_1376), .Y (n_718));
INVX2 g80169(.A (n_123), .Y (n_20767));
INVX2 g79503(.A (n_1273), .Y (n_6431));
CLKBUFX3 g80582(.A (n_537), .Y (n_1081));
NAND2X1 g77422(.A (u0_r0_rcnt[0] ), .B (u0_r0_rcnt[1] ), .Y(n_1204));
CLKBUFX3 g80800(.A (n_343), .Y (n_1015));
INVX1 g82159(.A (n_20102), .Y (n_20585));
CLKBUFX3 g80807(.A (n_109), .Y (n_1044));
INVX1 g78736(.A (n_27098), .Y (n_828));
INVX4 g80054(.A (n_3318), .Y (n_18792));
INVX1 g78888(.A (n_228), .Y (n_629));
INVX4 g79512(.A (n_26597), .Y (n_736));
INVX1 g81863(.A (n_26903), .Y (n_20055));
CLKBUFX3 g80240(.A (n_107), .Y (n_1080));
INVX2 g78653(.A (n_26041), .Y (n_877));
INVX4 g80019(.A (n_100), .Y (n_790));
INVX1 g81086(.A (n_20157), .Y (n_20680));
INVX1 g80422(.A (n_196), .Y (n_869));
INVX4 g81238(.A (n_5131), .Y (n_19934));
INVX2 g78708(.A (n_21174), .Y (n_903));
INVX1 g79714(.A (n_26276), .Y (n_494));
INVX2 g78984(.A (n_8217), .Y (n_16978));
INVX2 g80207(.A (n_457), .Y (n_479));
INVX2 g78441(.A (n_178), .Y (n_807));
INVX4 g79642(.A (n_101), .Y (n_5924));
INVX1 g81206(.A (n_20144), .Y (n_20204));
INVX1 g81857(.A (n_27242), .Y (n_875));
INVX4 g78482(.A (n_279), .Y (n_1147));
INVX1 g78680(.A (sa13[2] ), .Y (n_2921));
INVX1 g81717(.A (n_26833), .Y (n_98));
INVX1 g80233(.A (n_622), .Y (n_95));
INVX1 g80818(.A (n_109), .Y (n_775));
INVX1 g81399(.A (n_12760), .Y (n_591));
INVX1 g79479(.A (w2[27] ), .Y (n_1270));
CLKBUFX3 g82463(.A (sa30[4] ), .Y (n_230));
INVX1 g80241(.A (sa11[7] ), .Y (n_107));
INVX4 g81457(.A (w3[10] ), .Y (n_13083));
INVX2 g79052(.A (sa23[3] ), .Y (n_367));
INVX1 g80200(.A (w2[5] ), .Y (n_194));
INVX2 g82073(.A (w3[25] ), .Y (n_4357));
INVX1 g82130(.A (w0[8] ), .Y (n_2692));
INVX1 g82478(.A (n_645), .Y (n_23399));
INVX8 g81373(.A (w3[2] ), .Y (n_12827));
INVX2 g80788(.A (sa00[4] ), .Y (n_10315));
INVX4 g80527(.A (w3[4] ), .Y (n_5422));
INVX2 g79657(.A (sa33[6] ), .Y (n_89));
INVX1 g80613(.A (w3[14] ), .Y (n_474));
INVX1 g81681(.A (w1[5] ), .Y (n_23777));
CLKBUFX3 g81535(.A (sa23[2] ), .Y (n_673));
INVX1 g81231(.A (w0[7] ), .Y (n_2560));
INVX4 g82062(.A (w3[25] ), .Y (n_124));
INVX1 g82561(.A (w1[3] ), .Y (n_1236));
INVX1 g82509(.A (w3[16] ), .Y (n_250));
INVX1 g57641(.A (sa30[0] ), .Y (n_344));
INVX1 g78614(.A (n_22717), .Y (n_9203));
INVX2 g81747(.A (sa32[6] ), .Y (n_896));
INVX1 g80429(.A (w3[1] ), .Y (n_12788));
INVX8 g81177(.A (sa33[3] ), .Y (n_4861));
INVX1 g81475(.A (w2[30] ), .Y (n_22794));
INVX1 g79430(.A (w0[31] ), .Y (n_1103));
INVX1 g81886(.A (w2[19] ), .Y (n_1842));
INVX2 g80584(.A (sa03[7] ), .Y (n_537));
INVX4 g79022(.A (sa10[7] ), .Y (n_767));
INVX2 g78442(.A (sa23[5] ), .Y (n_178));
INVX1 g80321(.A (n_23257), .Y (n_141));
INVX1 g78314(.A (dcnt[1] ), .Y (n_77));
INVX2 g82516(.A (sa12[7] ), .Y (n_627));
INVX4 g82344(.A (w3[9] ), .Y (n_933));
INVX1 g79127(.A (w2[3] ), .Y (n_1235));
INVX2 g78398(.A (sa23[6] ), .Y (n_900));
INVX1 g81985(.A (u0_r0_rcnt[0] ), .Y (n_111));
INVX1 g80389(.A (sa11[5] ), .Y (n_1079));
INVX2 g79684(.A (w3[15] ), .Y (n_664));
INVX2 g80208(.A (sa21[7] ), .Y (n_457));
INVX1 g57022(.A (sa32[0] ), .Y (n_21915));
INVX2 g80085(.A (sa21[6] ), .Y (n_919));
INVX4 g78853(.A (sa22[2] ), .Y (n_9106));
INVX1 g78444(.A (w2[26] ), .Y (n_23191));
INVX2 g79387(.A (n_362), .Y (n_2779));
INVX1 g81713(.A (n_22781), .Y (n_97));
INVX1 g80195(.A (w0[2] ), .Y (n_2434));
INVX4 g78831(.A (sa22[2] ), .Y (n_263));
INVX1 g79673(.A (w2[8] ), .Y (n_1296));
INVX2 g82090(.A (sa32[5] ), .Y (n_315));
INVX1 g81460(.A (w2[31] ), .Y (n_1632));
INVX2 g81277(.A (sa13[5] ), .Y (n_2096));
INVX2 g81770(.A (sa32[4] ), .Y (n_386));
INVX1 g82127(.A (n_23567), .Y (n_112));
INVX2 g82234(.A (sa12[1] ), .Y (n_20018));
INVX1 g81871(.A (sa32[1] ), .Y (n_19486));
INVX2 g81608(.A (sa20[6] ), .Y (n_199));
INVX1 g82500(.A (w3[16] ), .Y (n_22214));
INVX4 g78413(.A (w3[13] ), .Y (n_3038));
INVX2 g81759(.A (sa23[7] ), .Y (n_899));
INVX1 g80172(.A (w2[21] ), .Y (n_23309));
INVX1 g81226(.A (n_2440), .Y (n_22831));
INVX2 g80388(.A (sa22[5] ), .Y (n_208));
INVX1 g78361(.A (w3[23] ), .Y (n_916));
INVX1 g80251(.A (w3[31] ), .Y (n_295));
INVX1 g80680(.A (w0[25] ), .Y (n_22569));
CLKBUFX1 g82119(.A (w3[29] ), .Y (n_348));
INVX4 g79845(.A (sa20[2] ), .Y (n_18237));
INVX1 g81991(.A (sa30[5] ), .Y (n_68));
INVX1 g80002(.A (ld), .Y (n_229));
INVX1 g81083(.A (sa33[1] ), .Y (n_19475));
INVX1 g80806(.A (w0[1] ), .Y (n_6401));
INVX2 g80767(.A (sa21[4] ), .Y (n_330));
INVX1 g79461(.A (w2[16] ), .Y (n_2648));
INVX2 g79894(.A (n_908), .Y (n_14627));
INVX1 g78843(.A (sa22[2] ), .Y (n_300));
INVX1 g78456(.A (sa10[3] ), .Y (n_280));
INVX2 g80020(.A (w3[5] ), .Y (n_100));
INVX2 g81562(.A (sa22[1] ), .Y (n_19414));
INVX2 g82464(.A (sa30[4] ), .Y (n_3338));
INVX4 g82264(.A (sa00[2] ), .Y (n_18266));
INVX1 g81097(.A (w0[28] ), .Y (n_23551));
CLKBUFX3 g80315(.A (sa11[3] ), .Y (n_319));
INVX1 g79140(.A (w1[27] ), .Y (n_332));
INVX2 g79739(.A (sa22[7] ), .Y (n_1043));
INVX1 g81480(.A (n_546), .Y (n_1072));
INVX1 g82481(.A (w2[9] ), .Y (n_22762));
INVX1 g82036(.A (w1[4] ), .Y (n_1164));
INVX1 g81094(.A (w2[28] ), .Y (n_1428));
INVX1 g79342(.A (w0[30] ), .Y (n_23241));
INVX1 g81980(.A (u0_r0_rcnt[2] ), .Y (n_63));
INVX2 g78995(.A (w3[26] ), .Y (n_8217));
INVX2 g81736(.A (sa10[4] ), .Y (n_4598));
INVX1 g78325(.A (sa13[1] ), .Y (n_62));
INVX1 g80174(.A (w3[7] ), .Y (n_561));
INVX1 g78334(.A (sa13[1] ), .Y (n_378));
CLKBUFX3 g80187(.A (w3[7] ), .Y (n_380));
INVX1 g81593(.A (w3[20] ), .Y (n_3736));
INVX1 g79458(.A (sa22[4] ), .Y (n_162));
INVX1 g82097(.A (sa30[6] ), .Y (n_528));
CLKBUFX1 g80744(.A (sa21[4] ), .Y (n_274));
INVX1 g81762(.A (w0[22] ), .Y (n_23238));
CLKBUFX3 g78492(.A (sa20[5] ), .Y (n_3560));
INVX2 g81281(.A (sa13[5] ), .Y (n_251));
INVX8 g79981(.A (ld), .Y (n_360));
INVX2 g81960(.A (sa13[3] ), .Y (n_320));
INVX1 g78771(.A (n_925), .Y (n_234));
CLKBUFX3 g78483(.A (sa10[3] ), .Y (n_279));
INVX1 g81201(.A (sa31[1] ), .Y (n_191));
INVX1 g79668(.A (w3[6] ), .Y (n_1431));
INVX4 g78574(.A (w3[28] ), .Y (n_379));
INVX2 g80664(.A (sa03[6] ), .Y (n_285));
INVX1 g78349(.A (w1[1] ), .Y (n_1040));
INVX1 g79660(.A (w0[17] ), .Y (n_22567));
INVX8 g79283(.A (n_2204), .Y (n_1196));
CLKBUFX3 g81994(.A (sa30[5] ), .Y (n_1947));
INVX1 g78950(.A (w3[0] ), .Y (n_22372));
INVX1 g80530(.A (w2[6] ), .Y (n_2437));
INVX4 g81798(.A (sa32[3] ), .Y (n_271));
INVX4 g80539(.A (sa03[3] ), .Y (n_4391));
INVX1 g79303(.A (w3[3] ), .Y (n_1376));
INVX1 g79137(.A (n_23580), .Y (n_6404));
INVX1 g79232(.A (w2[11] ), .Y (n_1555));
INVX4 g80097(.A (sa32[7] ), .Y (n_801));
INVX1 g79494(.A (w3[21] ), .Y (n_2462));
INVX4 g79248(.A (sa21[5] ), .Y (n_2943));
INVX1 g78905(.A (w3[30] ), .Y (n_731));
INVX1 g78510(.A (n_1138), .Y (n_22223));
INVX1 g82449(.A (w0[4] ), .Y (n_9624));
INVX4 g79174(.A (sa22[3] ), .Y (n_1942));
INVX4 g81590(.A (w3[20] ), .Y (n_3307));
INVX8 g81707(.A (w3[12] ), .Y (n_3920));
INVX1 g81007(.A (w2[4] ), .Y (n_1163));
INVX2 g82307(.A (sa01[7] ), .Y (n_434));
INVX2 g81741(.A (sa10[4] ), .Y (n_5381));
CLKBUFX2 g80104(.A (sa20[7] ), .Y (n_214));
INVX2 g80546(.A (sa03[3] ), .Y (n_11272));
INVX1 g79014(.A (w2[14] ), .Y (n_22787));
INVX1 g81178(.A (sa02[7] ), .Y (n_1185));
INVX1 g80030(.A (w0[6] ), .Y (n_243));
INVX4 g82115(.A (w3[29] ), .Y (n_827));
INVX1 g81930(.A (w1[0] ), .Y (n_1958));
INVX8 g79597(.A (sa11[2] ), .Y (n_9819));
INVX2 g79490(.A (sa11[6] ), .Y (n_772));
INVX4 g79630(.A (sa33[4] ), .Y (n_636));
INVX1 g82134(.A (w1[15] ), .Y (n_255));
INVX1 g78949(.A (w3[0] ), .Y (n_22274));
INVX2 g82511(.A (sa12[7] ), .Y (n_748));
INVX1 g80675(.A (w3[8] ), .Y (n_22423));
INVX1 g81211(.A (sa31[1] ), .Y (n_171));
INVX1 g79866(.A (sa20[2] ), .Y (n_106));
INVX1 g80881(.A (sa10[1] ), .Y (n_177));
INVX4 g80076(.A (w3[19] ), .Y (n_3318));
INVX1 g79133(.A (w1[31] ), .Y (n_338));
INVX1 g82085(.A (w1[25] ), .Y (n_153));
INVX1 g78892(.A (w2[10] ), .Y (n_23184));
INVX2 g80105(.A (sa20[7] ), .Y (n_959));
INVX2 g78376(.A (sa30[1] ), .Y (n_129));
INVX2 g80209(.A (sa21[7] ), .Y (n_912));
INVX1 g81390(.A (w2[17] ), .Y (n_22976));
INVX1 g81066(.A (w0[14] ), .Y (n_23234));
INVX2 g80803(.A (sa13[6] ), .Y (n_343));
CLKBUFX1 g82446(.A (sa20[3] ), .Y (n_183));
INVX1 g82557(.A (w1[16] ), .Y (n_23605));
INVX1 g82147(.A (sa23[1] ), .Y (n_164));
INVX1 g80267(.A (w2[24] ), .Y (n_1220));
INVX8 g81511(.A (sa23[2] ), .Y (n_17411));
INVX2 g81840(.A (sa31[6] ), .Y (n_849));
INVX1 g80501(.A (n_267), .Y (n_9342));
INVX1 g81749(.A (w2[18] ), .Y (n_23494));
INVX1 g80254(.A (w3[31] ), .Y (n_26));
INVX1 g78801(.A (w0[13] ), .Y (n_23087));
INVX2 g82032(.A (w3[17] ), .Y (n_3264));
INVX1 g80668(.A (w3[8] ), .Y (n_21708));
INVX1 g79634(.A (sa33[4] ), .Y (n_5643));
INVX1 g78621(.A (n_22653), .Y (n_23547));
INVX1 g79504(.A (w3[21] ), .Y (n_1273));
INVX2 g79670(.A (w3[6] ), .Y (n_176));
INVX1 g81461(.A (rst), .Y (n_10999));
INVX1 g81396(.A (w3[10] ), .Y (n_22));
INVX2 g78940(.A (sa20[4] ), .Y (n_238));
INVX1 g81214(.A (w1[18] ), .Y (n_23352));
INVX4 g78966(.A (w3[26] ), .Y (n_9527));
CLKBUFX3 g79643(.A (sa33[4] ), .Y (n_101));
INVX1 g79182(.A (sa22[3] ), .Y (n_9335));
INVX2 g80234(.A (sa11[7] ), .Y (n_622));
INVX1 g81269(.A (w1[9] ), .Y (n_22496));
INVX1 g80589(.A (w1[12] ), .Y (n_1005));
INVX1 g81380(.A (w1[20] ), .Y (n_23079));
INVX4 g79025(.A (sa00[5] ), .Y (n_218));
INVX1 g82122(.A (w2[1] ), .Y (n_1039));
INVX1 g79289(.A (sa33[0] ), .Y (n_21));
INVX1 g82217(.A (w2[7] ), .Y (n_1769));
INVX4 g80373(.A (w3[11] ), .Y (n_9057));
INVX1 g78598(.A (n_23363), .Y (n_22557));
INVX2 g81207(.A (sa31[1] ), .Y (n_20144));
INVX4 g80776(.A (sa00[4] ), .Y (n_5005));
INVX1 g81403(.A (w3[10] ), .Y (n_12760));
INVX2 g79476(.A (sa00[7] ), .Y (n_1285));
INVX2 g80819(.A (sa22[6] ), .Y (n_109));
INVX2 g80143(.A (w3[22] ), .Y (n_160));
INVX2 g81910(.A (sa30[3] ), .Y (n_352));
INVX1 g80608(.A (n_22778), .Y (n_245));
INVX4 g78709(.A (sa01[1] ), .Y (n_21174));
INVX1 g81382(.A (w2[20] ), .Y (n_23274));
INVX2 g79383(.A (sa21[3] ), .Y (n_6008));
CLKBUFX3 g81088(.A (sa33[1] ), .Y (n_20157));
INVX1 g79363(.A (sa21[3] ), .Y (n_135));
INVX1 g80024(.A (w1[14] ), .Y (n_22829));
INVX4 g82415(.A (sa20[3] ), .Y (n_2318));
INVX1 g78906(.A (w3[30] ), .Y (n_18));
INVX2 g78889(.A (sa00[6] ), .Y (n_228));
CLKBUFX1 g78904(.A (w3[30] ), .Y (n_440));
INVX2 g81979(.A (sa13[3] ), .Y (n_4173));
INVX1 g82244(.A (dcnt[2] ), .Y (n_328));
INVX1 g81376(.A (w2[13] ), .Y (n_23001));
INVX1 g81466(.A (w1[10] ), .Y (n_23047));
CLKBUFX3 g78595(.A (w3[28] ), .Y (n_213));
INVX1 g80262(.A (w0[9] ), .Y (n_22564));
INVX2 g82102(.A (sa30[6] ), .Y (n_464));
INVX1 g78946(.A (w3[0] ), .Y (n_21687));
INVX1 g79621(.A (n_2430), .Y (n_22964));
INVX1 g79338(.A (w3[3] ), .Y (n_152));
INVX1 g80190(.A (w0[3] ), .Y (n_16938));
INVX1 g82091(.A (sa32[5] ), .Y (n_15));
INVX1 g78386(.A (sa30[1] ), .Y (n_187));
INVX1 g78360(.A (w3[23] ), .Y (n_437));
INVX1 g81849(.A (sa20[0] ), .Y (n_21843));
INVX1 g80624(.A (w3[14] ), .Y (n_14));
INVX1 g79467(.A (w1[24] ), .Y (n_23261));
INVX1 g82212(.A (n_497), .Y (n_1019));
INVX1 g80682(.A (w2[15] ), .Y (n_2009));
INVX4 g82494(.A (sa30[7] ), .Y (n_527));
CLKBUFX3 g81782(.A (sa32[4] ), .Y (n_264));
INVX2 g81678(.A (sa03[4] ), .Y (n_4490));
INVX4 g80423(.A (w3[1] ), .Y (n_196));
INVX1 g79036(.A (w2[22] ), .Y (n_22789));
INVX2 g79646(.A (sa33[4] ), .Y (n_4825));
INVX1 g80908(.A (w2[25] ), .Y (n_9));
INVX1 g81892(.A (n_22981), .Y (n_1318));
INVX1 g82450(.A (sa30[4] ), .Y (n_4925));
INVX1 g57370(.A (sa31[0] ), .Y (n_21717));
INVX2 g82160(.A (sa23[1] ), .Y (n_20102));
INVX4 g78495(.A (sa20[5] ), .Y (n_1627));
INVX1 g82096(.A (sa32[5] ), .Y (n_1291));
CLKBUFX3 g80556(.A (sa03[3] ), .Y (n_294));
INVX2 g80302(.A (sa11[3] ), .Y (n_276));
INVX1 g80447(.A (w2[2] ), .Y (n_1960));
INVX1 g78624(.A (n_23290), .Y (n_23545));
CLKBUFX3 g79079(.A (sa23[3] ), .Y (n_205));
INVX1 g57367(.A (sa31[0] ), .Y (n_209));
INVX1 g81395(.A (w1[17] ), .Y (n_22591));
INVX1 g80612(.A (w0[10] ), .Y (n_16921));
CLKBUFX3 g79712(.A (sa32[2] ), .Y (n_290));
INVX1 g79434(.A (n_24366), .Y (n_23763));
INVX1 g80771(.A (w2[12] ), .Y (n_1004));
INVX4 g80737(.A (sa23[4] ), .Y (n_383));
INVX1 g78618(.A (w1[23] ), .Y (n_982));
INVX1 g82003(.A (w3[17] ), .Y (n_282));
CLKBUFX3 g80722(.A (sa23[4] ), .Y (n_277));
INVX1 g81091(.A (n_24266), .Y (n_22750));
INVX1 g79469(.A (sa00[7] ), .Y (n_2));
INVX1 g81716(.A (sa00[0] ), .Y (n_22251));
INVX1 g80253(.A (w3[31] ), .Y (n_730));
INVX2 g81186(.A (sa02[7] ), .Y (n_305));
INVX1 g79287(.A (w0[26] ), .Y (n_22546));
INVX1 g81387(.A (n_424), .Y (n_221));
INVX1 g81826(.A (sa11[0] ), .Y (n_0));
INVX1 g80170(.A (sa11[1] ), .Y (n_123));
INVX1 g82496(.A (w2[23] ), .Y (n_2174));
INVX1 g80482(.A (n_267), .Y (n_1512));
INVX1 g82076(.A (sa23[0] ), .Y (n_22231));
CLKBUFX1 g83097(.A (n_25739), .Y (n_25738));
CLKBUFX3 g83098(.A (n_27834), .Y (n_25739));
INVX1 g83099(.A (n_27834), .Y (n_25741));
INVX1 g83100(.A (n_27834), .Y (n_25826));
INVX1 g83101(.A (n_25745), .Y (n_25744));
CLKBUFX1 g83102(.A (n_25746), .Y (n_25745));
INVX1 g83103(.A (n_25746), .Y (n_25747));
INVX2 g83104(.A (n_2831), .Y (n_25746));
NAND2X1 g46(.A (n_25542), .B (n_25848), .Y (n_28277));
NOR2X1 g50(.A (n_13579), .B (n_16916), .Y (n_25848));
NAND2X1 g45(.A (n_25543), .B (n_25850), .Y (n_28278));
AND2X1 g47(.A (n_16348), .B (n_9242), .Y (n_25850));
NAND3X1 g62(.A (n_25855), .B (n_25857), .C (n_25865), .Y (n_25866));
NOR2X1 g73(.A (n_25709), .B (n_25708), .Y (n_25855));
INVX1 g70(.A (n_25856), .Y (n_25857));
AOI21X1 g71(.A0 (n_21135), .A1 (n_20602), .B0 (sa21[0] ), .Y(n_25856));
NOR2X1 g63(.A (n_25863), .B (n_25864), .Y (n_25865));
OAI21X1 g64(.A0 (n_14972), .A1 (n_27910), .B0 (n_25862), .Y(n_25863));
AND2X1 g65(.A (n_25858), .B (n_25861), .Y (n_25862));
NAND2X1 g72(.A (n_8896), .B (n_15997), .Y (n_25858));
INVX1 g67(.A (n_25861), .Y (n_25860));
NAND4X1 g68(.A (n_9392), .B (n_9442), .C (n_4689), .D (n_5530), .Y(n_25861));
AOI21X1 g69(.A0 (n_17730), .A1 (n_10384), .B0 (n_27919), .Y(n_25864));
NAND2X2 g42(.A (n_25881), .B (n_25888), .Y (n_25889));
INVX1 g83127(.A (n_25880), .Y (n_25881));
AOI21X1 g83128(.A0 (n_25877), .A1 (n_25878), .B0 (n_27786), .Y(n_25880));
NOR2X1 g83129(.A (n_25876), .B (n_21681), .Y (n_25877));
NOR2X1 g52(.A (n_9106), .B (n_17796), .Y (n_25876));
NAND2X1 g83130(.A (n_20928), .B (n_19414), .Y (n_25878));
NOR2X1 g83131(.A (n_25882), .B (n_25887), .Y (n_25888));
AOI21X1 g83132(.A0 (n_20976), .A1 (n_21018), .B0 (sa22[0] ), .Y(n_25882));
NAND2X1 g83133(.A (n_25884), .B (n_25886), .Y (n_25887));
INVX1 g53(.A (n_25883), .Y (n_25884));
NAND2X1 g54(.A (n_21218), .B (n_12665), .Y (n_25883));
INVX1 g83134(.A (n_25885), .Y (n_25886));
NAND3X1 g83135(.A (n_19288), .B (n_18091), .C (n_14674), .Y(n_25885));
NAND3X1 g83136(.A (n_25890), .B (n_25897), .C (n_25898), .Y(n_25899));
OAI21X1 g60(.A0 (n_21413), .A1 (n_15587), .B0 (n_209), .Y (n_25890));
AOI21X1 g57(.A0 (n_20631), .A1 (n_21581), .B0 (n_25896), .Y(n_25897));
NAND4X1 g58(.A (n_25891), .B (n_25893), .C (n_15678), .D (n_25895),.Y (n_25896));
OR2X1 g83137(.A (n_15371), .B (n_16457), .Y (n_25891));
AOI21X1 g61(.A0 (n_15748), .A1 (n_20399), .B0 (n_10175), .Y(n_25893));
INVX1 g83139(.A (n_25894), .Y (n_25895));
NOR2X1 g83140(.A (n_15509), .B (n_13815), .Y (n_25894));
OAI21X1 g59(.A0 (n_20658), .A1 (n_20888), .B0 (sa31[0] ), .Y(n_25898));
AND2X1 g83144(.A (n_18147), .B (n_14362), .Y (n_25901));
NOR2X1 g83145(.A (n_17147), .B (n_13262), .Y (n_25902));
NAND2X1 g83149(.A (n_16892), .B (n_27656), .Y (n_25907));
OAI21X1 g83152(.A0 (n_22046), .A1 (n_25911), .B0 (n_28080), .Y(n_25916));
INVX1 g83153(.A (sa03[0] ), .Y (n_25911));
AOI21X1 g83158(.A0 (n_25917), .A1 (n_20610), .B0 (n_25918), .Y(n_25919));
OR2X1 g83159(.A (n_20495), .B (n_19510), .Y (n_25917));
NAND3X1 g83160(.A (n_19753), .B (n_20001), .C (n_18925), .Y(n_25918));
NAND2X1 g21(.A (n_25923), .B (n_25924), .Y (n_25925));
NAND2X1 g22(.A (n_27491), .B (n_25922), .Y (n_25923));
INVX1 g25(.A (ld_r), .Y (n_25922));
NAND2X1 g24(.A (n_1691), .B (n_13768), .Y (n_25924));
INVX1 g27(.A (ld_r), .Y (n_25926));
NAND4X1 g37(.A (n_25938), .B (n_25940), .C (n_20222), .D (n_25941),.Y (n_25942));
AND2X1 g38(.A (n_18408), .B (n_25937), .Y (n_25938));
AOI21X1 g40(.A0 (n_18012), .A1 (n_19170), .B0 (n_25936), .Y(n_25937));
NAND2X1 g83165(.A (n_16868), .B (n_16867), .Y (n_25936));
AND2X1 g39(.A (n_20217), .B (n_25939), .Y (n_25940));
NAND2X1 g83166(.A (n_13842), .B (n_10859), .Y (n_25939));
NAND2X1 g41(.A (n_18873), .B (n_13575), .Y (n_25941));
NAND4X1 g83167(.A (n_25943), .B (n_25944), .C (n_25949), .D(n_21085), .Y (n_25950));
OAI21X1 g83168(.A0 (n_21410), .A1 (n_18242), .B0 (sa32[0] ), .Y(n_25943));
OAI21X1 g83169(.A0 (n_21004), .A1 (n_20875), .B0 (n_26899), .Y(n_25944));
NOR2X1 g83170(.A (n_25947), .B (n_25948), .Y (n_25949));
NAND4X1 g83171(.A (n_15612), .B (n_14990), .C (n_25946), .D (n_9830),.Y (n_25947));
INVX1 g83172(.A (n_25945), .Y (n_25946));
NOR2X1 g83173(.A (n_14991), .B (n_18168), .Y (n_25945));
NOR2X1 g83174(.A (n_1397), .B (n_18778), .Y (n_25948));
NOR2X1 g83176(.A (n_25951), .B (n_25954), .Y (n_25955));
NAND2X1 g83177(.A (n_17968), .B (n_11004), .Y (n_25951));
NOR2X1 g83178(.A (n_2681), .B (n_25953), .Y (n_25954));
NOR2X1 g83179(.A (n_20551), .B (n_19194), .Y (n_25953));
OAI21X1 g83180(.A0 (n_21114), .A1 (n_15638), .B0 (n_2681), .Y(n_25956));
OAI21X1 g83181(.A0 (n_25957), .A1 (n_25958), .B0 (sa21[0] ), .Y(n_25959));
NAND2X1 g83182(.A (n_25635), .B (n_25636), .Y (n_25957));
NAND2X1 g83183(.A (n_20203), .B (n_17254), .Y (n_25958));
OAI21X1 g83184(.A0 (n_25960), .A1 (n_25961), .B0 (n_27817), .Y(n_25963));
NAND2X1 g83185(.A (n_19195), .B (n_20059), .Y (n_25960));
NAND2X1 g83186(.A (n_20060), .B (n_11613), .Y (n_25961));
CLKBUFX1 g3(.A (n_26775), .Y (n_25965));
NAND4X1 g83210(.A (n_28848), .B (n_28849), .C (n_25995), .D(n_25996), .Y (n_25997));
NAND2X1 g83211(.A (n_21524), .B (sa13[0] ), .Y (n_28849));
AND2X1 g83212(.A (n_25991), .B (n_25992), .Y (n_28848));
OAI21X1 g83213(.A0 (n_20501), .A1 (n_11196), .B0 (n_487), .Y(n_25991));
OAI21X1 g83214(.A0 (n_20929), .A1 (n_21649), .B0 (n_378), .Y(n_25992));
NOR2X1 g83215(.A (n_19578), .B (n_25994), .Y (n_25995));
NOR2X1 g83216(.A (n_378), .B (n_20176), .Y (n_25994));
OAI21X1 g83217(.A0 (n_21279), .A1 (n_21649), .B0 (n_28127), .Y(n_25996));
INVX1 g83219(.A (n_25998), .Y (n_25999));
AOI21X1 g83220(.A0 (n_16672), .A1 (n_7169), .B0 (n_11400), .Y(n_25998));
AOI21X1 g83221(.A0 (n_29205), .A1 (n_11400), .B0 (n_27646), .Y(n_26007));
NAND2X1 g83223(.A (n_4549), .B (n_6946), .Y (n_26000));
NAND3X1 g83231(.A (n_26019), .B (n_26020), .C (n_26028), .Y(n_26029));
NAND2X1 g83232(.A (n_26012), .B (n_26018), .Y (n_26019));
INVX1 g79(.A (n_26011), .Y (n_26012));
INVX1 g80(.A (sa33[0] ), .Y (n_26011));
NAND3X1 g83233(.A (n_20042), .B (n_26015), .C (n_26017), .Y(n_26018));
NAND2X1 g83234(.A (n_26013), .B (n_19924), .Y (n_26015));
INVX1 g81(.A (n_20796), .Y (n_26013));
AND2X1 g83235(.A (n_18597), .B (n_26016), .Y (n_26017));
OR2X1 g83236(.A (n_3724), .B (n_12449), .Y (n_26016));
NOR2X1 g83237(.A (n_21658), .B (n_21549), .Y (n_26020));
AND2X1 g83238(.A (n_26021), .B (n_26027), .Y (n_26028));
INVX1 g83239(.A (n_19775), .Y (n_26021));
NOR2X1 g83240(.A (n_26024), .B (n_26026), .Y (n_26027));
NAND3X1 g83241(.A (n_26022), .B (n_9894), .C (n_16661), .Y (n_26024));
INVX1 g76(.A (n_12438), .Y (n_26022));
NAND2X1 g83242(.A (n_26025), .B (n_13277), .Y (n_26026));
INVX1 g82(.A (n_15616), .Y (n_26025));
NAND2X1 g83243(.A (n_26036), .B (n_26037), .Y (n_26038));
NOR2X1 g83244(.A (n_26030), .B (n_26035), .Y (n_26036));
AND2X1 g49_dup(.A (n_6615), .B (n_9982), .Y (n_26030));
NAND2X1 g83245(.A (n_26033), .B (n_26034), .Y (n_26035));
NAND3X1 g83246(.A (n_10162), .B (n_11215), .C (n_26032), .Y(n_26033));
INVX1 g83247(.A (n_27604), .Y (n_26032));
NAND2X1 g83249(.A (n_5476), .B (n_27604), .Y (n_26034));
OAI21X1 g83250(.A0 (n_25571), .A1 (n_12604), .B0 (n_15708), .Y(n_26037));
INVX1 g83251(.A (n_26039), .Y (n_26040));
AND2X1 g83252(.A (n_9982), .B (n_6615), .Y (n_26039));
INVX2 g83253(.A (sa13[2] ), .Y (n_26041));
NAND2X2 g83254(.A (n_10162), .B (n_11215), .Y (n_26042));
NAND3X1 g83255(.A (n_26043), .B (n_26045), .C (n_26054), .Y(n_26055));
NOR2X1 g83256(.A (n_21847), .B (n_21959), .Y (n_26043));
INVX1 g83257(.A (n_26044), .Y (n_26045));
AOI21X1 g83258(.A0 (n_21134), .A1 (n_21230), .B0 (sa23[0] ), .Y(n_26044));
NOR2X1 g83259(.A (n_26052), .B (n_26053), .Y (n_26054));
OAI21X1 g83260(.A0 (n_18298), .A1 (n_21442), .B0 (n_26051), .Y(n_26052));
AND2X1 g83261(.A (n_26047), .B (n_26050), .Y (n_26051));
INVX1 g83263(.A (n_26047), .Y (n_26048));
NAND2X2 g83264(.A (n_11901), .B (n_11902), .Y (n_26047));
NAND2X1 g83265(.A (n_10968), .B (n_2701), .Y (n_26050));
AOI21X1 g83266(.A0 (n_16367), .A1 (n_16601), .B0 (n_27028), .Y(n_26053));
CLKBUFX1 g83267(.A (n_26061), .Y (n_26062));
NAND4X1 g83268(.A (n_26057), .B (n_26058), .C (n_26059), .D(n_26060), .Y (n_26061));
NAND2X1 g83269(.A (n_26056), .B (sa00[0] ), .Y (n_26057));
NAND4X1 g83270(.A (n_19743), .B (n_20038), .C (n_20675), .D(n_18744), .Y (n_26056));
OAI21X1 g83271(.A0 (n_21008), .A1 (n_18893), .B0 (n_22251), .Y(n_26058));
NOR2X1 g83272(.A (n_20896), .B (n_21083), .Y (n_26059));
OAI21X1 g83273(.A0 (n_20804), .A1 (n_19495), .B0 (n_21520), .Y(n_26060));
NOR2X1 g83275(.A (n_26063), .B (n_26064), .Y (n_26065));
NAND2X1 g83276(.A (n_18017), .B (n_26840), .Y (n_26063));
NOR2X1 g83277(.A (n_19961), .B (n_17212), .Y (n_26064));
NAND2X1 g83278(.A (n_18876), .B (n_17822), .Y (n_26066));
AND2X1 g83279(.A (n_14267), .B (n_26069), .Y (n_26070));
NAND3X1 g83280(.A (n_26068), .B (n_5329), .C (n_20767), .Y (n_26069));
NAND4X1 g83281(.A (n_15605), .B (n_8891), .C (n_14308), .D (n_16421),.Y (n_26068));
OAI21X1 g83283(.A0 (n_18472), .A1 (n_17930), .B0 (n_19981), .Y(n_26071));
NAND4X1 g83285(.A (n_26073), .B (n_26078), .C (n_26080), .D(n_20777), .Y (n_26081));
OAI21X1 g83286(.A0 (n_22075), .A1 (n_19644), .B0 (n_27786), .Y(n_26073));
NAND2X1 g83287(.A (sa22[0] ), .B (n_26077), .Y (n_26078));
NAND4X1 g83288(.A (n_26075), .B (n_26076), .C (n_19725), .D(n_19374), .Y (n_26077));
INVX1 g83289(.A (n_26074), .Y (n_26075));
AOI21X1 g83290(.A0 (n_16753), .A1 (n_15117), .B0 (n_21275), .Y(n_26074));
AND2X1 g83291(.A (n_11843), .B (n_17608), .Y (n_26076));
INVX1 g83292(.A (n_26079), .Y (n_26080));
NAND4X1 g83293(.A (n_21190), .B (n_18092), .C (n_16898), .D(n_17606), .Y (n_26079));
NAND2X2 g83294(.A (n_26086), .B (n_26091), .Y (n_26092));
AOI21X1 g83295(.A0 (n_26083), .A1 (n_28127), .B0 (n_26085), .Y(n_26086));
NAND4X1 g83296(.A (n_20233), .B (n_21015), .C (n_19404), .D(n_18256), .Y (n_26083));
AOI21X1 g83298(.A0 (n_29123), .A1 (n_29124), .B0 (n_27526), .Y(n_26085));
NOR2X1 g83299(.A (n_26089), .B (n_26090), .Y (n_26091));
NAND3X1 g83300(.A (n_21177), .B (n_26088), .C (n_19161), .Y(n_26089));
AOI21X1 g83301(.A0 (n_15708), .A1 (n_10604), .B0 (n_26087), .Y(n_26088));
NAND2X1 g83302(.A (n_27528), .B (n_17331), .Y (n_26087));
NAND2X1 g83303(.A (n_19703), .B (n_15221), .Y (n_26090));
AOI21X1 g83305(.A0 (n_16322), .A1 (n_20412), .B0 (n_26093), .Y(n_26094));
NAND2X1 g83306(.A (n_10141), .B (n_17098), .Y (n_26093));
OAI21X1 g83307(.A0 (n_26038), .A1 (n_15910), .B0 (n_27449), .Y(n_26095));
AOI21X1 g83308(.A0 (n_12293), .A1 (n_4930), .B0 (n_26096), .Y(n_26097));
AND2X1 g83309(.A (n_6446), .B (n_6442), .Y (n_26096));
NAND2X1 g83310(.A (n_17653), .B (n_19408), .Y (n_26098));
NAND2X2 g29(.A (n_26101), .B (n_26103), .Y (n_26104));
AND2X1 g31(.A (n_22349), .B (n_26100), .Y (n_26101));
NAND2X1 g33(.A (n_21665), .B (sa21[0] ), .Y (n_26100));
AND2X1 g30(.A (n_21634), .B (n_26102), .Y (n_26103));
AOI22X1 g32(.A0 (n_4614), .A1 (n_18074), .B0 (n_27913), .B1(n_29062), .Y (n_26102));
NAND4X1 g36(.A (n_26130), .B (n_26134), .C (n_21104), .D (n_21593),.Y (n_26135));
INVX1 g83335(.A (n_26129), .Y (n_26130));
AOI21X1 g83336(.A0 (n_21156), .A1 (n_19441), .B0 (n_825), .Y(n_26129));
NOR2X1 g83337(.A (n_26132), .B (n_26133), .Y (n_26134));
NAND4X1 g83338(.A (n_17191), .B (n_16625), .C (n_13421), .D(n_14988), .Y (n_26132));
INVX1 g83340(.A (n_21070), .Y (n_26133));
CLKBUFX2 g83341(.A (n_26144), .Y (n_26145));
NAND4X1 g83342(.A (n_29308), .B (n_26137), .C (n_29309), .D(n_26143), .Y (n_26144));
NOR2X1 g83343(.A (n_19035), .B (n_21455), .Y (n_29309));
OAI21X1 g83344(.A0 (n_21471), .A1 (n_20329), .B0 (sa20[0] ), .Y(n_26137));
OAI21X1 g83345(.A0 (n_26138), .A1 (n_26139), .B0 (n_26140), .Y(n_29308));
NAND3X1 g83346(.A (n_25454), .B (n_15339), .C (n_18014), .Y(n_26138));
NAND3X1 g83347(.A (n_25455), .B (n_18951), .C (n_9048), .Y (n_26139));
INVX1 g83348(.A (sa20[0] ), .Y (n_26140));
AOI21X1 g83349(.A0 (n_17827), .A1 (n_20271), .B0 (n_26142), .Y(n_26143));
AND2X1 g83350(.A (n_19806), .B (n_21314), .Y (n_26142));
OR2X1 g83364(.A (n_2363), .B (n_19175), .Y (n_26156));
NAND2X1 g83365(.A (n_27847), .B (n_21915), .Y (n_26159));
OAI21X1 g83366(.A0 (n_20945), .A1 (n_26801), .B0 (sa32[0] ), .Y(n_26160));
NAND3X1 g83367(.A (n_26165), .B (n_26167), .C (n_26168), .Y(n_26169));
OAI21X1 g83368(.A0 (n_26162), .A1 (n_26164), .B0 (sa12[0] ), .Y(n_26165));
NAND2X1 g83369(.A (n_21332), .B (n_19786), .Y (n_26162));
NAND2X1 g83370(.A (n_26163), .B (n_26842), .Y (n_26164));
NOR2X1 g83371(.A (n_18323), .B (n_17999), .Y (n_26163));
AOI21X1 g83372(.A0 (n_27624), .A1 (n_21077), .B0 (n_26166), .Y(n_26167));
NAND4X1 g83373(.A (n_29422), .B (n_29423), .C (n_18140), .D(n_17831), .Y (n_26166));
OAI21X1 g83374(.A0 (n_21260), .A1 (n_12043), .B0 (n_27718), .Y(n_26168));
NAND4X1 g83376(.A (n_28249), .B (n_21576), .C (n_26173), .D(n_28250), .Y (n_26180));
OAI21X1 g83377(.A0 (n_20840), .A1 (n_20372), .B0 (n_21757), .Y(n_28250));
INVX1 g83378(.A (n_26172), .Y (n_26173));
AOI21X1 g83379(.A0 (n_20820), .A1 (n_20181), .B0 (sa30[0] ), .Y(n_26172));
AND2X1 g83380(.A (n_26175), .B (n_26178), .Y (n_28249));
INVX1 g83381(.A (n_26174), .Y (n_26175));
AOI21X1 g83382(.A0 (n_17733), .A1 (n_10072), .B0 (n_2682), .Y(n_26174));
NOR2X1 g83383(.A (n_26176), .B (n_26177), .Y (n_26178));
NAND3X1 g83384(.A (n_13347), .B (n_8502), .C (n_16642), .Y (n_26176));
NOR2X1 g83385(.A (n_129), .B (n_15621), .Y (n_26177));
NOR2X1 g83390(.A (n_28151), .B (n_28157), .Y (n_26185));
INVX1 g83393(.A (n_27640), .Y (n_26192));
INVX1 g83395(.A (n_26185), .Y (n_26194));
OAI21X1 g83399(.A0 (n_21704), .A1 (n_18952), .B0 (n_21717), .Y(n_26197));
AOI21X1 g83400(.A0 (n_20756), .A1 (n_20144), .B0 (n_26198), .Y(n_26199));
AOI21X1 g83401(.A0 (n_17393), .A1 (n_8124), .B0 (n_15371), .Y(n_26198));
OAI21X1 g83402(.A0 (n_20738), .A1 (n_20870), .B0 (sa31[0] ), .Y(n_26200));
AOI21X1 g83403(.A0 (n_18803), .A1 (n_18889), .B0 (n_26203), .Y(n_26204));
NAND3X1 g83404(.A (n_26202), .B (n_18007), .C (n_17262), .Y(n_26203));
INVX1 g83405(.A (n_26201), .Y (n_26202));
AOI21X1 g83406(.A0 (n_13449), .A1 (n_18645), .B0 (n_2917), .Y(n_26201));
XOR2X1 g83412(.A (n_26214), .B (n_26215), .Y (n_26216));
CLKBUFX1 g83413(.A (n_26213), .Y (n_26214));
INVX2 g83414(.A (n_26212), .Y (n_26213));
INVX2 g83415(.A (n_26211), .Y (n_26212));
NAND4X1 g83416(.A (n_28251), .B (n_28252), .C (n_21345), .D(n_21326), .Y (n_26211));
NAND2X1 g34_dup(.A (n_27683), .B (n_13685), .Y (n_26215));
NAND2X2 g83417(.A (n_27683), .B (n_13685), .Y (n_26217));
INVX2 g83418(.A (n_26213), .Y (n_26218));
NAND4X1 g83419(.A (n_26219), .B (n_26222), .C (n_21756), .D(n_26224), .Y (n_26225));
NAND2X1 g83420(.A (n_98), .B (n_21963), .Y (n_26219));
NOR2X1 g83421(.A (n_26220), .B (n_26221), .Y (n_26222));
INVX1 g83422(.A (n_20225), .Y (n_26220));
NOR2X1 g83423(.A (sa00[0] ), .B (n_21516), .Y (n_26221));
AOI21X1 g83424(.A0 (n_20226), .A1 (n_13575), .B0 (n_26223), .Y(n_26224));
NAND3X1 g83425(.A (n_15858), .B (n_17915), .C (n_16545), .Y(n_26223));
NAND4X1 g83426(.A (n_26226), .B (n_21383), .C (n_26227), .D(n_26231), .Y (n_26232));
OAI21X1 g83427(.A0 (n_21412), .A1 (n_16991), .B0 (n_26011), .Y(n_26226));
OAI21X1 g83428(.A0 (n_20984), .A1 (n_20604), .B0 (sa33[0] ), .Y(n_26227));
NOR2X1 g83429(.A (n_26229), .B (n_26230), .Y (n_26231));
NAND4X1 g83430(.A (n_26228), .B (n_15615), .C (n_14333), .D(n_15642), .Y (n_26229));
OR2X1 g83431(.A (n_15689), .B (n_17912), .Y (n_26228));
NOR2X1 g83432(.A (n_26368), .B (n_16413), .Y (n_26230));
NAND4X1 g83433(.A (n_26236), .B (n_26237), .C (n_26238), .D(n_26240), .Y (n_26241));
OAI21X1 g83434(.A0 (n_26233), .A1 (n_26234), .B0 (sa22[0] ), .Y(n_26236));
INVX1 g83435(.A (n_21118), .Y (n_26233));
NAND3X1 g83436(.A (n_21327), .B (n_20262), .C (n_14601), .Y(n_26234));
OAI21X1 g83438(.A0 (n_21845), .A1 (n_17016), .B0 (n_27786), .Y(n_26237));
NOR2X1 g83439(.A (n_17028), .B (n_21196), .Y (n_26238));
NAND2X1 g83440(.A (n_26239), .B (sa22[1] ), .Y (n_26240));
OR2X1 g83441(.A (n_19555), .B (n_19474), .Y (n_26239));
CLKBUFX2 g83442(.A (n_26241), .Y (n_26242));
NAND3X1 g83443(.A (n_26243), .B (n_26245), .C (n_26251), .Y(n_26252));
NOR2X1 g83444(.A (n_21772), .B (n_21999), .Y (n_26243));
INVX1 g83445(.A (n_26244), .Y (n_26245));
AOI21X1 g83446(.A0 (n_20827), .A1 (n_21229), .B0 (sa22[0] ), .Y(n_26244));
NOR2X1 g83447(.A (n_26249), .B (n_26250), .Y (n_26251));
OAI21X1 g83448(.A0 (n_21275), .A1 (n_17189), .B0 (n_26248), .Y(n_26249));
AND2X1 g83449(.A (n_26246), .B (n_26247), .Y (n_26248));
NAND2X1 g83450(.A (n_5670), .B (n_9899), .Y (n_26246));
NAND2X1 g83451(.A (n_6870), .B (n_12613), .Y (n_26247));
AOI21X1 g83452(.A0 (n_17726), .A1 (n_14940), .B0 (n_4851), .Y(n_26250));
INVX1 g83453(.A (n_26246), .Y (n_26253));
NAND3X1 g83461(.A (n_26261), .B (n_26268), .C (n_26272), .Y(n_26273));
OAI21X1 g83462(.A0 (n_19717), .A1 (n_13254), .B0 (n_1397), .Y(n_26261));
NOR2X1 g83463(.A (n_26264), .B (n_26267), .Y (n_26268));
NAND3X1 g83464(.A (n_13104), .B (n_26263), .C (n_4619), .Y (n_26264));
INVX1 g83465(.A (n_26262), .Y (n_26263));
AOI21X1 g83466(.A0 (n_10988), .A1 (n_10987), .B0 (sa32[2] ), .Y(n_26262));
NOR2X1 g83467(.A (n_19486), .B (n_26266), .Y (n_26267));
NOR2X1 g83469(.A (n_9765), .B (n_14045), .Y (n_26266));
NAND2X1 g83470(.A (n_26269), .B (n_26271), .Y (n_26272));
NAND2X1 g83471(.A (n_17239), .B (n_10986), .Y (n_26269));
INVX1 g83472(.A (n_26270), .Y (n_26271));
INVX1 g83473(.A (sa32[2] ), .Y (n_26270));
INVX4 g83476(.A (sa32[2] ), .Y (n_26276));
NAND4X1 g83477(.A (n_29145), .B (n_29146), .C (n_26284), .D(n_26286), .Y (n_26287));
OAI21X1 g83478(.A0 (n_26278), .A1 (n_26279), .B0 (sa32[0] ), .Y(n_29146));
NAND3X1 g83479(.A (n_20693), .B (n_20173), .C (n_26277), .Y(n_26278));
AND2X1 g83480(.A (n_17054), .B (n_20626), .Y (n_26277));
NAND2X1 g83481(.A (n_17950), .B (n_25946), .Y (n_26279));
NOR2X1 g83482(.A (n_26281), .B (n_26282), .Y (n_29145));
NAND2X1 g83483(.A (n_19853), .B (n_15102), .Y (n_26281));
INVX1 g83484(.A (n_20815), .Y (n_26282));
OAI21X1 g83485(.A0 (n_20868), .A1 (n_20357), .B0 (n_21915), .Y(n_26284));
AOI21X1 g83486(.A0 (n_19457), .A1 (n_1397), .B0 (n_26285), .Y(n_26286));
AND2X1 g83487(.A (n_17823), .B (n_18121), .Y (n_26285));
NAND4X1 g83498(.A (n_25515), .B (n_21663), .C (n_21960), .D(n_25516), .Y (n_26297));
INVX1 g83499(.A (n_26297), .Y (n_26298));
NAND4X1 g83500(.A (n_26299), .B (n_26300), .C (n_21568), .D(n_26302), .Y (n_26303));
INVX1 g83501(.A (n_21991), .Y (n_26299));
NAND2X1 g83502(.A (n_21786), .B (sa01[0] ), .Y (n_26300));
NOR2X1 g83503(.A (n_26301), .B (n_20713), .Y (n_26302));
NAND3X1 g83504(.A (n_14323), .B (n_17540), .C (n_17906), .Y(n_26301));
INVX1 g83506(.A (n_26297), .Y (n_26306));
CLKBUFX2 g83507(.A (n_26316), .Y (n_26317));
NAND4X1 g83508(.A (n_26307), .B (n_26308), .C (n_26309), .D(n_26315), .Y (n_26316));
NAND2X1 g83509(.A (n_21911), .B (sa01[0] ), .Y (n_26307));
OAI21X1 g83510(.A0 (n_21312), .A1 (n_18127), .B0 (n_28206), .Y(n_26308));
OAI21X1 g83511(.A0 (n_20475), .A1 (n_20506), .B0 (n_903), .Y(n_26309));
AND2X1 g83512(.A (n_26310), .B (n_26314), .Y (n_26315));
OAI21X1 g83513(.A0 (n_18358), .A1 (n_19191), .B0 (n_21174), .Y(n_26310));
AOI21X1 g83514(.A0 (n_15305), .A1 (n_19364), .B0 (n_26313), .Y(n_26314));
NOR2X1 g83515(.A (n_26311), .B (n_26312), .Y (n_26313));
INVX1 g83516(.A (n_20765), .Y (n_26311));
NOR2X1 g83517(.A (n_8161), .B (n_15303), .Y (n_26312));
NAND3X1 g83518(.A (n_26319), .B (n_26322), .C (n_26326), .Y(n_26327));
INVX1 g83519(.A (n_26318), .Y (n_26319));
AOI21X1 g83520(.A0 (n_25700), .A1 (n_25701), .B0 (n_27817), .Y(n_26318));
NAND2X1 g83521(.A (n_27817), .B (n_29325), .Y (n_26322));
NAND4X1 g83522(.A (n_20643), .B (n_18991), .C (n_19388), .D(n_19656), .Y (n_29325));
NOR2X1 g83524(.A (n_26325), .B (n_21498), .Y (n_26326));
NAND4X1 g83525(.A (n_26323), .B (n_26324), .C (n_14459), .D(n_14972), .Y (n_26325));
INVX1 g83526(.A (n_17417), .Y (n_26323));
AOI21X1 g83527(.A0 (n_29102), .A1 (n_9092), .B0 (n_16635), .Y(n_26324));
OAI21X1 g83550(.A0 (n_26710), .A1 (n_26358), .B0 (n_28206), .Y(n_26360));
INVX1 g83553(.A (n_14801), .Y (n_26350));
NAND2X1 g83557(.A (n_26356), .B (n_26357), .Y (n_26358));
NAND2X1 g83558(.A (n_13328), .B (n_17459), .Y (n_26356));
NAND2X1 g83559(.A (n_17543), .B (n_14630), .Y (n_26357));
NAND2X1 g83561(.A (n_26361), .B (n_26366), .Y (n_26367));
NAND2X1 g83562(.A (n_21), .B (n_29197), .Y (n_26361));
NAND2X1 g83563(.A (n_26365), .B (sa33[1] ), .Y (n_26366));
NAND4X1 g83564(.A (n_19653), .B (n_16111), .C (n_26364), .D(n_12666), .Y (n_26365));
NOR2X1 g83565(.A (n_26362), .B (n_26363), .Y (n_26364));
NOR2X1 g83566(.A (n_5804), .B (n_1363), .Y (n_26362));
INVX1 g83567(.A (n_16570), .Y (n_26363));
INVX1 g83568(.A (sa33[1] ), .Y (n_26368));
NAND2X1 g83570(.A (n_16690), .B (n_2001), .Y (n_26369));
NAND2X1 g83571(.A (n_10182), .B (n_13804), .Y (n_26370));
NOR2X1 g83572(.A (n_26374), .B (n_26376), .Y (n_26377));
NAND2X1 g83573(.A (n_26371), .B (n_26372), .Y (n_26374));
OR2X1 g83574(.A (n_11276), .B (n_10996), .Y (n_26371));
OR2X1 g83576(.A (n_6185), .B (n_5915), .Y (n_26372));
INVX1 g83577(.A (n_26375), .Y (n_26376));
NAND2X1 g83578(.A (n_8269), .B (n_10389), .Y (n_26375));
INVX1 g83579(.A (n_26379), .Y (n_26380));
INVX1 g83580(.A (n_26371), .Y (n_26379));
INVX1 g83581(.A (n_26372), .Y (n_26381));
AND2X1 g83582(.A (n_26385), .B (n_26386), .Y (n_26388));
NOR2X1 g83583(.A (n_26383), .B (n_26384), .Y (n_26385));
CLKBUFX1 g83584(.A (n_26382), .Y (n_26383));
INVX2 g83585(.A (sa13[7] ), .Y (n_26382));
CLKBUFX1 g83586(.A (sa13[5] ), .Y (n_26384));
CLKBUFX3 g83588(.A (sa13[4] ), .Y (n_26386));
INVX1 g83593(.A (sa13[4] ), .Y (n_26393));
INVX2 g83594(.A (n_26382), .Y (n_26394));
INVX1 g83595(.A (n_26384), .Y (n_26395));
INVX2 g83596(.A (n_26403), .Y (n_26404));
NAND4X1 g83597(.A (n_26398), .B (n_26399), .C (n_26401), .D(n_26402), .Y (n_26403));
NAND2X1 g83598(.A (n_26396), .B (n_21757), .Y (n_26398));
NAND2X1 g83599(.A (n_21298), .B (n_18875), .Y (n_26396));
NAND2X1 g83601(.A (n_21205), .B (n_21507), .Y (n_26399));
NOR2X1 g83602(.A (n_26400), .B (n_21616), .Y (n_26401));
NAND2X1 g83603(.A (n_16693), .B (n_7785), .Y (n_26400));
NAND2X1 g83604(.A (n_21668), .B (n_344), .Y (n_26402));
INVX1 g83607(.A (sa01[0] ), .Y (n_26405));
NAND4X1 g83608(.A (n_19674), .B (n_20115), .C (n_15412), .D(n_11498), .Y (n_26406));
NAND2X1 g83612(.A (n_16762), .B (n_19594), .Y (n_26410));
NAND2X1 g83613(.A (n_20775), .B (n_19645), .Y (n_26411));
NAND2X2 g83614(.A (n_26417), .B (n_26422), .Y (n_26423));
AOI21X1 g83615(.A0 (n_26414), .A1 (n_26844), .B0 (n_26416), .Y(n_26417));
NAND4X1 g83616(.A (n_25696), .B (n_20701), .C (n_19393), .D(n_25697), .Y (n_26414));
AOI21X1 g83618(.A0 (n_25833), .A1 (n_25834), .B0 (n_27624), .Y(n_26416));
NOR2X1 g83619(.A (n_26420), .B (n_26421), .Y (n_26422));
NAND3X1 g83620(.A (n_25592), .B (n_26419), .C (n_19156), .Y(n_26420));
AOI21X1 g83621(.A0 (n_10444), .A1 (n_19398), .B0 (n_26418), .Y(n_26419));
NAND2X1 g83622(.A (n_16157), .B (n_17157), .Y (n_26418));
NAND2X1 g83623(.A (n_25591), .B (n_16673), .Y (n_26421));
NAND3X1 g83624(.A (n_26424), .B (n_26427), .C (n_26432), .Y(n_26433));
NAND2X1 g83625(.A (n_22195), .B (n_22266), .Y (n_26424));
NOR2X1 g83626(.A (n_26425), .B (n_26426), .Y (n_26427));
NAND3X1 g83627(.A (n_11570), .B (n_10646), .C (n_18080), .Y(n_26425));
NAND2X1 g83628(.A (n_21724), .B (n_21423), .Y (n_26426));
OAI21X1 g83629(.A0 (n_26428), .A1 (n_26430), .B0 (n_27624), .Y(n_26432));
NAND3X1 g83630(.A (n_20759), .B (n_17838), .C (n_12226), .Y(n_26428));
NAND2X1 g83631(.A (n_26429), .B (n_20331), .Y (n_26430));
OAI21X1 g83632(.A0 (n_16523), .A1 (n_10252), .B0 (n_15574), .Y(n_26429));
NAND3X1 g83634(.A (n_26434), .B (n_26437), .C (n_26440), .Y(n_26441));
OAI21X1 g83635(.A0 (n_21417), .A1 (n_15645), .B0 (n_825), .Y(n_26434));
NOR2X1 g83636(.A (n_20913), .B (n_26436), .Y (n_26437));
OR2X1 g83637(.A (n_26435), .B (n_21439), .Y (n_26436));
OR2X1 g83638(.A (n_12854), .B (n_18083), .Y (n_26435));
OAI21X1 g83639(.A0 (n_26438), .A1 (n_26439), .B0 (sa10[0] ), .Y(n_26440));
NAND4X1 g83640(.A (n_20336), .B (n_14481), .C (n_14332), .D(n_13725), .Y (n_26438));
OAI21X1 g83641(.A0 (n_19618), .A1 (n_21108), .B0 (n_18496), .Y(n_26439));
NAND2X1 g83656(.A (n_26466), .B (n_26467), .Y (n_26468));
AOI21X1 g83657(.A0 (n_26458), .A1 (n_28631), .B0 (n_26465), .Y(n_26466));
NAND2X1 g83658(.A (n_26456), .B (n_26457), .Y (n_26458));
NOR2X1 g83659(.A (n_7185), .B (n_4713), .Y (n_26456));
OR2X1 g83660(.A (n_8093), .B (n_6346), .Y (n_26457));
NAND2X1 g83661(.A (n_26461), .B (n_26464), .Y (n_26465));
NAND2X1 g60_dup(.A (n_8024), .B (n_753), .Y (n_26461));
NAND2X2 g83664(.A (n_29389), .B (n_881), .Y (n_26464));
INVX1 g83666(.A (n_4906), .Y (n_29389));
NAND2X1 g83667(.A (n_7800), .B (n_28692), .Y (n_26467));
NAND2X1 g83668(.A (n_8024), .B (n_753), .Y (n_26469));
INVX2 g83669(.A (n_26464), .Y (n_26470));
NAND4X1 g83671(.A (n_26472), .B (n_26473), .C (n_26476), .D(n_26480), .Y (n_26481));
AND2X1 g83672(.A (n_21349), .B (n_21356), .Y (n_26472));
OAI21X1 g83673(.A0 (n_21157), .A1 (n_20371), .B0 (sa11[0] ), .Y(n_26473));
NAND2X1 g83674(.A (n_26474), .B (n_3483), .Y (n_26476));
NAND2X1 g83675(.A (n_20166), .B (n_10242), .Y (n_26474));
INVX1 g83677(.A (n_26479), .Y (n_26480));
NAND2X1 g83678(.A (n_17195), .B (n_26478), .Y (n_26479));
INVX1 g83679(.A (n_26477), .Y (n_26478));
NAND3X1 g83680(.A (n_13372), .B (n_17240), .C (n_17904), .Y(n_26477));
NAND2X2 g83681(.A (n_26489), .B (n_26491), .Y (n_26492));
INVX1 g83682(.A (n_26488), .Y (n_26489));
NAND2X1 g83683(.A (n_26483), .B (n_2241), .Y (n_26488));
INVX2 g83684(.A (n_26482), .Y (n_26483));
NAND2X1 g83685(.A (n_28568), .B (n_981), .Y (n_26482));
INVX2 g83687(.A (n_26485), .Y (n_26486));
INVX1 g83688(.A (n_27368), .Y (n_26485));
INVX4 g83690(.A (n_26490), .Y (n_26491));
CLKBUFX3 g83691(.A (sa31[3] ), .Y (n_26490));
INVX1 g83692(.A (sa31[3] ), .Y (n_26493));
INVX1 g83693(.A (n_26483), .Y (n_26494));
NAND2X1 g83695(.A (n_21785), .B (sa02[0] ), .Y (n_26495));
AND2X1 g83696(.A (n_21350), .B (n_26497), .Y (n_26498));
AOI21X1 g83697(.A0 (n_18262), .A1 (n_16553), .B0 (n_26496), .Y(n_26497));
NAND2X1 g83698(.A (n_16830), .B (n_15863), .Y (n_26496));
NOR2X1 g83699(.A (n_26499), .B (n_26500), .Y (n_26501));
NAND2X1 g83700(.A (n_19659), .B (n_14549), .Y (n_26499));
NOR2X1 g83701(.A (sa02[0] ), .B (n_21320), .Y (n_26500));
NAND4X1 g83702(.A (n_26503), .B (n_26507), .C (n_26508), .D(n_26509), .Y (n_26510));
NAND2X1 g83703(.A (n_22005), .B (sa11[0] ), .Y (n_26503));
NOR2X1 g83704(.A (n_21499), .B (n_26506), .Y (n_26507));
NAND2X1 g83705(.A (n_26504), .B (n_26505), .Y (n_26506));
INVX1 g83706(.A (n_18491), .Y (n_26504));
AOI21X1 g83707(.A0 (n_8003), .A1 (n_3967), .B0 (n_16725), .Y(n_26505));
NAND2X1 g83708(.A (n_27192), .B (n_22086), .Y (n_26508));
AOI22X1 g83709(.A0 (n_11096), .A1 (n_5329), .B0 (n_5329), .B1(n_10374), .Y (n_26509));
CLKBUFX2 g83710(.A (n_26521), .Y (n_26522));
NAND4X1 g83711(.A (n_29317), .B (n_26518), .C (n_26519), .D(n_29318), .Y (n_26521));
AOI21X1 g83712(.A0 (n_20290), .A1 (n_21442), .B0 (n_26512), .Y(n_29318));
INVX1 g83713(.A (n_26511), .Y (n_26512));
AOI21X1 g83714(.A0 (n_17565), .A1 (n_20269), .B0 (n_18372), .Y(n_26511));
NAND2X1 g83715(.A (sa23[0] ), .B (n_26517), .Y (n_26518));
NAND4X1 g83716(.A (n_26515), .B (n_26516), .C (n_20256), .D(n_19373), .Y (n_26517));
INVX1 g83717(.A (n_26514), .Y (n_26515));
AOI21X1 g83718(.A0 (n_17984), .A1 (n_19598), .B0 (n_20102), .Y(n_26514));
AND2X1 g83719(.A (n_16087), .B (n_9906), .Y (n_26516));
INVX1 g83720(.A (n_20886), .Y (n_26519));
OAI21X1 g83721(.A0 (n_21706), .A1 (n_19641), .B0 (n_22231), .Y(n_29317));
NAND2X2 g83722(.A (n_26525), .B (n_26533), .Y (n_26534));
NAND2X1 g83723(.A (n_26523), .B (n_26524), .Y (n_26525));
INVX1 g83724(.A (n_26140), .Y (n_26523));
NAND2X1 g83725(.A (n_22261), .B (n_19078), .Y (n_26524));
NOR2X1 g83726(.A (n_26527), .B (n_26532), .Y (n_26533));
NAND4X1 g83727(.A (n_20934), .B (n_19322), .C (n_18098), .D(n_26526), .Y (n_26527));
AND2X1 g83728(.A (n_14719), .B (n_9327), .Y (n_26526));
AOI21X1 g83729(.A0 (n_26528), .A1 (n_26531), .B0 (sa20[0] ), .Y(n_26532));
NAND2X1 g83730(.A (n_20847), .B (n_804), .Y (n_26528));
NOR2X1 g83731(.A (n_26529), .B (n_26530), .Y (n_26531));
NAND3X1 g83732(.A (n_9848), .B (n_17503), .C (n_12381), .Y (n_26529));
INVX1 g83733(.A (n_19946), .Y (n_26530));
OAI21X1 g83735(.A0 (n_21905), .A1 (n_26535), .B0 (n_26539), .Y(n_26540));
INVX1 g83736(.A (sa02[0] ), .Y (n_26535));
NAND4X1 g83737(.A (n_28508), .B (n_28509), .C (n_19822), .D(n_26535), .Y (n_26539));
NOR2X1 g83738(.A (n_26536), .B (n_26537), .Y (n_28508));
NAND2X1 g83739(.A (n_16827), .B (n_17707), .Y (n_26536));
OR2X1 g83740(.A (n_13619), .B (n_15370), .Y (n_26537));
AOI21X1 g83741(.A0 (n_26541), .A1 (n_2204), .B0 (n_26542), .Y(n_26543));
OR2X1 g83742(.A (n_20488), .B (n_19470), .Y (n_26541));
NAND3X1 g83743(.A (n_20380), .B (n_19748), .C (n_18136), .Y(n_26542));
INVX1 g19(.A (n_26549), .Y (n_26550));
NAND2X1 g20(.A (n_26547), .B (n_28154), .Y (n_26549));
NOR2X1 g83744(.A (n_28786), .B (n_26546), .Y (n_26547));
NAND2X2 g83746(.A (n_25802), .B (n_1305), .Y (n_26546));
INVX1 g83752(.A (sa03[0] ), .Y (n_26553));
NAND2X1 g83755(.A (n_26555), .B (n_28079), .Y (n_26556));
NAND2X1 g83756(.A (n_13784), .B (n_17884), .Y (n_26555));
NAND2X1 g16(.A (n_28341), .B (n_26601), .Y (n_26602));
NOR2X1 g17(.A (sa33[6] ), .B (n_736), .Y (n_28341));
INVX2 g83794(.A (sa33[7] ), .Y (n_26597));
INVX1 g83795(.A (n_26989), .Y (n_26601));
INVX1 g18(.A (sa33[6] ), .Y (n_26603));
NAND3X1 g83805(.A (n_26616), .B (n_13760), .C (n_26617), .Y(n_26618));
NOR2X1 g83806(.A (n_28165), .B (n_26615), .Y (n_26616));
NAND2X1 g83808(.A (n_18316), .B (n_26614), .Y (n_26615));
INVX1 g83809(.A (n_26613), .Y (n_26614));
NOR2X1 g83810(.A (n_10452), .B (n_7163), .Y (n_26613));
NAND2X1 g83811(.A (n_10922), .B (n_15039), .Y (n_26617));
AOI21X1 g83812(.A0 (n_28243), .A1 (n_1593), .B0 (n_26630), .Y(n_26631));
INVX1 g83814(.A (sa01[0] ), .Y (n_26619));
NAND3X1 g83815(.A (n_26621), .B (n_26622), .C (n_26625), .Y(n_28243));
AOI21X1 g83816(.A0 (n_21110), .A1 (n_21174), .B0 (n_20722), .Y(n_26621));
INVX1 g83817(.A (n_27697), .Y (n_26622));
AND2X1 g83818(.A (n_26623), .B (n_26624), .Y (n_26625));
INVX1 g83819(.A (n_14767), .Y (n_26623));
INVX1 g83820(.A (n_20705), .Y (n_26624));
NAND3X1 g83821(.A (n_25481), .B (n_26629), .C (n_21613), .Y(n_26630));
NOR2X1 g83822(.A (n_26627), .B (n_26628), .Y (n_26629));
INVX1 g83823(.A (n_14970), .Y (n_26627));
INVX1 g83824(.A (n_25482), .Y (n_26628));
XOR2X1 g83825(.A (n_28884), .B (n_28883), .Y (n_26637));
INVX2 g83826(.A (n_26634), .Y (n_28883));
CLKBUFX3 g83827(.A (n_26633), .Y (n_26634));
INVX2 g83828(.A (n_26632), .Y (n_26633));
NAND4X1 g83829(.A (n_22099), .B (n_21627), .C (n_21342), .D(n_21323), .Y (n_26632));
NAND2X1 g31_dup(.A (n_22657), .B (n_15489), .Y (n_28884));
NAND2X2 g83830(.A (n_22657), .B (n_15489), .Y (n_26638));
CLKBUFX1 g83831(.A (n_26638), .Y (n_26639));
INVX4 g83832(.A (n_26633), .Y (n_26640));
NAND2X1 g83840(.A (n_20311), .B (n_9802), .Y (n_26646));
XOR2X1 g83843(.A (w0[18] ), .B (n_29003), .Y (n_26654));
NAND4X1 g83849(.A (n_26657), .B (n_26666), .C (n_26667), .D(n_26668), .Y (n_26669));
OAI21X1 g83850(.A0 (n_18518), .A1 (n_16507), .B0 (n_187), .Y(n_26657));
NAND2X1 g83851(.A (n_26662), .B (n_26665), .Y (n_26666));
NAND2X1 g83852(.A (n_17319), .B (n_26661), .Y (n_26662));
AND2X1 g83853(.A (n_10806), .B (n_18456), .Y (n_26661));
NAND2X1 g83857(.A (n_26663), .B (n_14624), .Y (n_26665));
AND2X1 g83858(.A (n_11100), .B (n_11099), .Y (n_26663));
OAI21X1 g83860(.A0 (n_12252), .A1 (n_9828), .B0 (n_20558), .Y(n_26667));
AND2X1 g83861(.A (n_13108), .B (n_6042), .Y (n_26668));
INVX1 g83862(.A (sa30[2] ), .Y (n_26670));
NAND2X2 g83863(.A (n_26676), .B (n_26679), .Y (n_26680));
AOI21X1 g83864(.A0 (n_27239), .A1 (n_22156), .B0 (n_26675), .Y(n_26676));
NAND2X1 g83865(.A (n_26671), .B (n_26674), .Y (n_26675));
NAND2X1 g83866(.A (n_21076), .B (sa32[0] ), .Y (n_26671));
AND2X1 g83867(.A (n_26672), .B (n_26673), .Y (n_26674));
OR2X1 g83868(.A (n_7584), .B (n_7933), .Y (n_26672));
NAND2X1 g83869(.A (n_12572), .B (n_15986), .Y (n_26673));
AND2X1 g83870(.A (n_26677), .B (n_26678), .Y (n_26679));
OAI21X1 g83871(.A0 (n_20621), .A1 (n_8881), .B0 (n_1397), .Y(n_26677));
OAI21X1 g83872(.A0 (n_19455), .A1 (n_16920), .B0 (n_20648), .Y(n_26678));
NAND2X2 g83874(.A (n_26686), .B (n_26690), .Y (n_26691));
NOR2X1 g83875(.A (n_26684), .B (n_26685), .Y (n_26686));
OAI21X1 g83876(.A0 (n_21127), .A1 (n_20157), .B0 (n_26683), .Y(n_26684));
AND2X1 g83877(.A (n_20662), .B (n_26682), .Y (n_26683));
OR4X1 g83878(.A (n_4149), .B (n_2968), .C (n_7453), .D (n_17912), .Y(n_26682));
NOR2X1 g83879(.A (n_21678), .B (n_26011), .Y (n_26685));
AOI21X1 g83880(.A0 (n_26687), .A1 (n_27617), .B0 (n_26689), .Y(n_26690));
NAND3X1 g83881(.A (n_20299), .B (n_20158), .C (n_15897), .Y(n_26687));
INVX1 g83883(.A (n_8125), .Y (n_26689));
NAND3X1 g83884(.A (n_26695), .B (n_26700), .C (n_26701), .Y(n_26702));
AOI21X1 g83885(.A0 (n_26692), .A1 (n_20399), .B0 (n_26694), .Y(n_26695));
NAND2X1 g83886(.A (n_9908), .B (n_9693), .Y (n_26692));
AOI21X1 g83888(.A0 (n_16893), .A1 (n_9879), .B0 (n_191), .Y(n_26694));
NOR2X1 g83889(.A (n_26698), .B (n_15572), .Y (n_26700));
NAND2X1 g83890(.A (n_26696), .B (n_26697), .Y (n_26698));
NAND2X1 g83891(.A (n_11934), .B (n_18679), .Y (n_26696));
AND2X1 g83892(.A (n_5693), .B (n_10786), .Y (n_26697));
OAI21X1 g83894(.A0 (n_18695), .A1 (n_14110), .B0 (n_20144), .Y(n_26701));
NAND3X1 g83895(.A (n_26706), .B (n_26708), .C (n_26709), .Y(n_26710));
AND2X1 g83896(.A (n_26350), .B (n_26705), .Y (n_26706));
NOR2X1 g83897(.A (n_26703), .B (n_26704), .Y (n_26705));
NOR2X1 g83898(.A (n_14630), .B (n_10381), .Y (n_26703));
NOR2X1 g83899(.A (n_12494), .B (n_9668), .Y (n_26704));
AND2X1 g83900(.A (n_16875), .B (n_26707), .Y (n_26708));
NAND2X1 g83901(.A (n_16279), .B (n_13585), .Y (n_26707));
NAND2X1 g83902(.A (n_16378), .B (n_1113), .Y (n_26709));
INVX1 g83905(.A (n_26704), .Y (n_26713));
NAND2X1 g83909(.A (n_20384), .B (n_17714), .Y (n_26715));
NAND3X1 g83910(.A (n_20748), .B (n_20030), .C (n_18120), .Y(n_26716));
NAND4X1 g83912(.A (n_26721), .B (n_26724), .C (n_26725), .D(n_26729), .Y (n_26730));
INVX1 g83913(.A (n_26720), .Y (n_26721));
NOR2X1 g83914(.A (n_28680), .B (n_10948), .Y (n_26720));
NAND2X1 g83915(.A (n_9808), .B (n_28689), .Y (n_26724));
OAI21X1 g48(.A0 (n_14462), .A1 (n_5881), .B0 (n_28645), .Y (n_26725));
NOR2X1 g49(.A (n_26727), .B (n_26728), .Y (n_26729));
INVX1 g83918(.A (n_26726), .Y (n_26727));
NAND2X1 g83919(.A (n_5370), .B (n_1365), .Y (n_26726));
NOR2X1 g83920(.A (n_8904), .B (n_28134), .Y (n_26728));
INVX1 g83921(.A (n_26728), .Y (n_26731));
NAND2X2 g83922(.A (n_26734), .B (n_26742), .Y (n_26743));
NAND2X1 g83923(.A (n_26732), .B (n_26733), .Y (n_26734));
INVX1 g83924(.A (n_22231), .Y (n_26732));
NAND2X1 g83925(.A (n_22047), .B (n_18473), .Y (n_26733));
NOR2X1 g83926(.A (n_26739), .B (n_26741), .Y (n_26742));
AOI21X1 g83927(.A0 (n_26735), .A1 (n_26738), .B0 (sa23[0] ), .Y(n_26739));
NAND2X1 g83928(.A (n_20585), .B (n_20844), .Y (n_26735));
NOR2X1 g83929(.A (n_26736), .B (n_26737), .Y (n_26738));
NAND3X1 g83930(.A (n_11776), .B (n_17501), .C (n_12536), .Y(n_26736));
INVX1 g83931(.A (n_19939), .Y (n_26737));
NAND4X1 g83932(.A (n_21207), .B (n_19851), .C (n_18089), .D(n_26740), .Y (n_26741));
AND2X1 g83933(.A (n_14619), .B (n_9273), .Y (n_26740));
NAND2X2 g83934(.A (n_26746), .B (n_26750), .Y (n_26751));
NOR2X1 g83935(.A (n_26744), .B (n_26745), .Y (n_26746));
INVX1 g83936(.A (n_22148), .Y (n_26744));
NOR2X1 g43(.A (n_26833), .B (n_22268), .Y (n_26745));
AOI21X1 g83937(.A0 (n_21216), .A1 (n_20862), .B0 (n_26749), .Y(n_26750));
OAI21X1 g83938(.A0 (n_26747), .A1 (n_20862), .B0 (n_26748), .Y(n_26749));
AND2X1 g44(.A (n_19821), .B (n_17915), .Y (n_26747));
MX2X1 g83939(.A (n_17031), .B (n_16970), .S0 (n_16835), .Y (n_26748));
NAND2X1 g83963(.A (n_26778), .B (n_26779), .Y (n_26780));
OR2X1 g83964(.A (n_26775), .B (n_26777), .Y (n_26778));
NAND4X1 g83965(.A (n_25955), .B (n_25956), .C (n_25959), .D(n_25963), .Y (n_26775));
INVX1 g83966(.A (n_26776), .Y (n_26777));
NAND4X1 g40_dup(.A (n_25503), .B (n_21815), .C (n_21842), .D(n_25504), .Y (n_26776));
NAND2X1 g83967(.A (n_26777), .B (n_26775), .Y (n_26779));
NAND4X1 g83968(.A (n_21815), .B (n_25503), .C (n_21842), .D(n_25504), .Y (n_26781));
NAND3X1 g83969(.A (n_26786), .B (n_26787), .C (n_26791), .Y(n_26792));
OAI21X1 g83970(.A0 (n_26782), .A1 (n_26784), .B0 (n_28179), .Y(n_26786));
NAND2X1 g83971(.A (n_20554), .B (n_19979), .Y (n_26782));
NAND2X1 g83972(.A (n_18312), .B (n_26783), .Y (n_26784));
NAND2X2 g83973(.A (n_3047), .B (n_5833), .Y (n_26783));
OAI21X1 g83975(.A0 (n_20489), .A1 (n_9437), .B0 (n_21487), .Y(n_26787));
OAI21X1 g83976(.A0 (n_20901), .A1 (n_26788), .B0 (n_26790), .Y(n_26791));
NAND2X1 g83977(.A (n_26783), .B (n_17933), .Y (n_26788));
NAND2X1 g83978(.A (n_17742), .B (n_26789), .Y (n_26790));
INVX1 g83979(.A (n_17933), .Y (n_26789));
NOR2X1 g83981(.A (n_26903), .B (n_26800), .Y (n_26801));
NOR2X1 g83983(.A (n_4148), .B (n_26799), .Y (n_26800));
NAND3X1 g83984(.A (n_26795), .B (n_26796), .C (n_26798), .Y(n_26799));
INVX1 g83985(.A (n_13623), .Y (n_26795));
NAND2X2 g83986(.A (n_9933), .B (n_7331), .Y (n_26796));
INVX1 g83987(.A (n_26797), .Y (n_26798));
NOR2X1 g83988(.A (n_5854), .B (n_5255), .Y (n_26797));
INVX1 g83989(.A (n_26796), .Y (n_26802));
NAND4X1 g84001(.A (n_26814), .B (n_26815), .C (n_26820), .D(n_26821), .Y (n_26822));
OAI21X1 g84002(.A0 (n_21933), .A1 (n_17223), .B0 (n_0), .Y (n_26814));
AND2X1 g84003(.A (n_26065), .B (n_26070), .Y (n_26815));
OAI21X1 g84004(.A0 (n_26817), .A1 (n_26819), .B0 (sa11[0] ), .Y(n_26820));
NAND3X1 g84005(.A (n_20730), .B (n_19700), .C (n_26816), .Y(n_26817));
INVX1 g84006(.A (n_14301), .Y (n_26816));
NAND3X1 g84007(.A (n_26818), .B (n_14289), .C (n_11045), .Y(n_26819));
NAND2X1 g84008(.A (n_18035), .B (n_21188), .Y (n_26818));
AND2X1 g84009(.A (n_26066), .B (n_26071), .Y (n_26821));
AOI21X1 g84011(.A0 (sa00[0] ), .A1 (n_26829), .B0 (n_26831), .Y(n_26832));
NAND4X1 g84013(.A (n_20721), .B (n_26826), .C (n_26827), .D(n_26828), .Y (n_26829));
NAND2X1 g84015(.A (n_1008), .B (n_29323), .Y (n_26826));
INVX1 g84016(.A (n_21121), .Y (n_26827));
NOR2X1 g84017(.A (n_19021), .B (n_14768), .Y (n_26828));
NAND3X1 g84018(.A (n_22292), .B (n_21611), .C (n_26830), .Y(n_26831));
AND2X1 g84019(.A (n_17880), .B (n_19696), .Y (n_26830));
INVX1 g84020(.A (sa00[0] ), .Y (n_26833));
NAND2X1 g84021(.A (n_26836), .B (n_26838), .Y (n_26839));
NAND2X1 g84022(.A (n_26834), .B (n_20729), .Y (n_26836));
NAND2X1 g84023(.A (n_9979), .B (n_9722), .Y (n_26834));
AOI21X1 g84025(.A0 (n_10790), .A1 (n_9978), .B0 (n_26837), .Y(n_26838));
AND2X1 g84026(.A (n_10747), .B (n_9978), .Y (n_26837));
INVX1 g84027(.A (n_26837), .Y (n_26840));
NAND4X1 g84028(.A (n_29372), .B (n_29373), .C (n_26848), .D(n_26850), .Y (n_26851));
OAI21X1 g84029(.A0 (n_26841), .A1 (n_26843), .B0 (n_26844), .Y(n_29373));
NAND2X1 g84030(.A (n_20560), .B (n_20373), .Y (n_26841));
NAND2X1 g84031(.A (n_18324), .B (n_26842), .Y (n_26843));
NAND2X1 g84032(.A (n_6665), .B (n_3022), .Y (n_26842));
INVX1 g84033(.A (sa12[0] ), .Y (n_26844));
OAI21X1 g84034(.A0 (n_20912), .A1 (n_26846), .B0 (n_27718), .Y(n_29372));
INVX1 g84035(.A (n_26842), .Y (n_26846));
OAI21X1 g84036(.A0 (n_20124), .A1 (n_11379), .B0 (n_20810), .Y(n_26848));
INVX1 g84037(.A (n_26849), .Y (n_26850));
NOR2X1 g84038(.A (n_27718), .B (n_19592), .Y (n_26849));
INVX1 g84043(.A (n_18844), .Y (n_26853));
NOR2X1 g84044(.A (n_26854), .B (n_17216), .Y (n_26855));
INVX1 g84045(.A (n_26783), .Y (n_26854));
AND2X1 g84048(.A (n_18172), .B (n_15050), .Y (n_26858));
NAND3X1 g84050(.A (n_26863), .B (n_26864), .C (n_26870), .Y(n_26871));
OAI21X1 g84051(.A0 (n_20645), .A1 (n_20878), .B0 (sa30[0] ), .Y(n_26863));
OAI21X1 g84052(.A0 (n_21411), .A1 (n_15581), .B0 (n_344), .Y(n_26864));
AOI21X1 g84053(.A0 (n_20629), .A1 (n_15766), .B0 (n_26869), .Y(n_26870));
NAND4X1 g84054(.A (n_26866), .B (n_15621), .C (n_26868), .D (n_9936),.Y (n_26869));
INVX1 g84055(.A (n_26865), .Y (n_26866));
NOR2X1 g84056(.A (n_129), .B (n_16425), .Y (n_26865));
AOI21X1 g84057(.A0 (n_15738), .A1 (n_20388), .B0 (n_26867), .Y(n_26868));
NOR2X1 g84058(.A (n_15513), .B (n_16754), .Y (n_26867));
INVX1 g84059(.A (n_26867), .Y (n_26872));
NOR2X1 g84060(.A (n_26877), .B (n_26881), .Y (n_26882));
INVX1 g84061(.A (n_26874), .Y (n_26877));
INVX8 g84064(.A (n_26873), .Y (n_26874));
INVX4 g84065(.A (sa01[3] ), .Y (n_26873));
NAND2X1 g84066(.A (n_26878), .B (n_26880), .Y (n_26881));
NOR2X1 g84067(.A (n_3700), .B (n_28464), .Y (n_26878));
INVX2 g84068(.A (n_26879), .Y (n_26880));
CLKBUFX1 g84069(.A (sa01[4] ), .Y (n_26879));
INVX4 g84070(.A (n_26874), .Y (n_26883));
INVX1 g84072(.A (sa01[4] ), .Y (n_26885));
NOR2X1 g84073(.A (n_26887), .B (n_26889), .Y (n_26890));
INVX1 g84074(.A (sa10[4] ), .Y (n_26887));
NAND2X1 g84076(.A (n_26888), .B (sa10[5] ), .Y (n_26889));
INVX2 g84077(.A (sa10[6] ), .Y (n_26888));
INVX1 g84078(.A (n_26888), .Y (n_26891));
CLKBUFX3 g84079(.A (n_27204), .Y (n_26893));
NOR2X1 g84081(.A (n_26896), .B (n_26897), .Y (n_26898));
NAND2X1 g84082(.A (n_26894), .B (n_26895), .Y (n_26896));
NAND2X1 g84083(.A (n_19256), .B (n_19852), .Y (n_26894));
NAND2X1 g84084(.A (n_15953), .B (n_14807), .Y (n_26895));
NAND3X1 g84085(.A (n_26156), .B (n_19997), .C (n_18122), .Y(n_26897));
INVX2 g84086(.A (n_26909), .Y (n_26910));
NAND2X2 g84087(.A (n_26899), .B (n_26908), .Y (n_26909));
INVX1 g84088(.A (sa32[0] ), .Y (n_26899));
NAND4X1 g84089(.A (n_26904), .B (n_20647), .C (n_26907), .D(n_20324), .Y (n_26908));
NAND2X1 g84090(.A (n_26902), .B (n_26903), .Y (n_26904));
NAND2X1 g84091(.A (n_26900), .B (n_26901), .Y (n_26902));
NOR2X1 g84092(.A (n_10166), .B (n_17426), .Y (n_26900));
NOR2X1 g84093(.A (n_9590), .B (n_9829), .Y (n_26901));
INVX1 g84094(.A (sa32[1] ), .Y (n_26903));
NOR2X1 g84095(.A (n_26905), .B (n_26906), .Y (n_26907));
INVX1 g84096(.A (n_9539), .Y (n_26905));
NOR2X1 g84097(.A (n_16974), .B (n_16376), .Y (n_26906));
NAND4X1 g84098(.A (n_26911), .B (n_26912), .C (n_26913), .D(n_26914), .Y (n_26915));
OAI21X1 g84099(.A0 (n_8684), .A1 (n_27431), .B0 (n_29074), .Y(n_26911));
NAND2X1 g84100(.A (n_6304), .B (n_29102), .Y (n_26912));
NAND3X1 g84101(.A (n_27439), .B (n_5799), .C (n_29065), .Y (n_26913));
NAND3X1 g84102(.A (n_29106), .B (n_6008), .C (n_7959), .Y (n_26914));
NAND2X1 g84103(.A (n_6008), .B (n_7959), .Y (n_26916));
NAND3X1 g84105(.A (n_26922), .B (n_26923), .C (n_26928), .Y(n_26929));
NAND2X1 g84106(.A (n_26918), .B (n_26921), .Y (n_26922));
NAND3X1 g84107(.A (n_21583), .B (n_21278), .C (sa20[0] ), .Y(n_26918));
NAND4X1 g84108(.A (n_26919), .B (n_25672), .C (n_19929), .D(n_26920), .Y (n_26921));
AND2X1 g84109(.A (n_19012), .B (n_25673), .Y (n_26919));
INVX1 g84110(.A (sa20[0] ), .Y (n_26920));
INVX1 g84111(.A (n_21306), .Y (n_26923));
NOR2X1 g84112(.A (n_26927), .B (n_19701), .Y (n_26928));
NAND4X1 g84113(.A (n_18014), .B (n_26924), .C (n_17329), .D(n_26926), .Y (n_26927));
NAND2X1 g84114(.A (n_11994), .B (n_11261), .Y (n_26924));
INVX1 g84116(.A (n_16727), .Y (n_26926));
AOI21X1 g84117(.A0 (n_28588), .A1 (n_28589), .B0 (n_27624), .Y(n_26937));
NAND2X1 g84118(.A (n_26930), .B (n_26931), .Y (n_28589));
NAND3X1 g84119(.A (n_25678), .B (n_25679), .C (n_17982), .Y(n_26930));
INVX1 g84120(.A (sa12[1] ), .Y (n_26931));
NOR2X1 g84121(.A (n_27132), .B (n_27589), .Y (n_28588));
NAND4X1 g84125(.A (n_26938), .B (n_26939), .C (n_26941), .D(n_26942), .Y (n_26943));
OAI21X1 g84126(.A0 (n_21848), .A1 (n_19723), .B0 (sa11[0] ), .Y(n_26938));
OAI21X1 g84127(.A0 (n_21256), .A1 (n_10421), .B0 (n_20729), .Y(n_26939));
AOI21X1 g84128(.A0 (n_21355), .A1 (n_27192), .B0 (n_26940), .Y(n_26941));
NAND2X1 g84129(.A (n_20036), .B (n_18903), .Y (n_26940));
AND2X1 g84130(.A (n_17881), .B (n_19589), .Y (n_26942));
MX2X1 g84131(.A (n_23025), .B (n_26944), .S0 (n_26947), .Y (n_26948));
NAND2X2 g84132(.A (n_25916), .B (n_25919), .Y (n_26944));
NOR2X1 g84133(.A (n_26945), .B (n_26946), .Y (n_26947));
NAND2X1 g84134(.A (n_22320), .B (n_22143), .Y (n_26945));
NAND2X1 g84135(.A (n_21750), .B (n_21420), .Y (n_26946));
NAND4X1 g84136(.A (n_21750), .B (n_21420), .C (n_22320), .D(n_22143), .Y (n_26949));
NAND3X1 g84137(.A (n_26950), .B (n_26951), .C (n_26956), .Y(n_26957));
AOI21X1 g84138(.A0 (n_14983), .A1 (n_2091), .B0 (n_16360), .Y(n_26950));
NAND2X1 g84139(.A (n_17732), .B (n_28631), .Y (n_26951));
AOI21X1 g84140(.A0 (n_13957), .A1 (n_14627), .B0 (n_26955), .Y(n_26956));
OR2X1 g84141(.A (n_14628), .B (n_26954), .Y (n_26955));
NOR2X1 g84142(.A (n_26952), .B (n_28631), .Y (n_26954));
NAND2X2 g84143(.A (n_7498), .B (n_11003), .Y (n_26952));
INVX1 g84145(.A (n_26952), .Y (n_26958));
NAND2X2 g84147(.A (n_26963), .B (n_26966), .Y (n_26967));
NOR2X1 g84148(.A (n_26960), .B (n_26962), .Y (n_26963));
NOR2X1 g84149(.A (n_22231), .B (n_22065), .Y (n_26960));
NAND2X1 g84150(.A (n_21865), .B (n_26961), .Y (n_26962));
MX2X1 g84151(.A (n_17040), .B (n_15493), .S0 (n_17411), .Y (n_26961));
AOI21X1 g84152(.A0 (n_26964), .A1 (n_21442), .B0 (n_26965), .Y(n_26966));
OR2X1 g84153(.A (n_16913), .B (n_20757), .Y (n_26964));
AOI21X1 g84154(.A0 (n_19887), .A1 (n_26047), .B0 (n_21442), .Y(n_26965));
CLKBUFX1 g84156(.A (n_26977), .Y (n_26978));
NAND4X1 g84157(.A (n_26969), .B (n_26970), .C (n_26973), .D(n_26976), .Y (n_26977));
OAI21X1 g84158(.A0 (n_20869), .A1 (n_20737), .B0 (sa30[0] ), .Y(n_26969));
OAI21X1 g84159(.A0 (n_21416), .A1 (n_18933), .B0 (n_344), .Y(n_26970));
AOI21X1 g84160(.A0 (n_20752), .A1 (n_21507), .B0 (n_26972), .Y(n_26973));
NAND3X1 g84161(.A (n_26971), .B (n_18756), .C (n_17177), .Y(n_26972));
NAND2X1 g84162(.A (n_17003), .B (n_18800), .Y (n_26971));
NOR2X1 g84163(.A (n_26974), .B (n_26975), .Y (n_26976));
AOI21X1 g84164(.A0 (n_13443), .A1 (n_14857), .B0 (n_2682), .Y(n_26974));
AOI21X1 g84165(.A0 (n_17392), .A1 (n_8337), .B0 (n_129), .Y(n_26975));
INVX2 g84166(.A (n_26986), .Y (n_26987));
NAND2X2 g84167(.A (n_26983), .B (n_26985), .Y (n_26986));
NOR2X1 g84168(.A (n_26979), .B (n_26982), .Y (n_26983));
NAND2X1 g84169(.A (n_15084), .B (n_7198), .Y (n_26979));
NAND2X1 g84170(.A (n_26980), .B (n_26981), .Y (n_26982));
NAND2X1 g84171(.A (n_21219), .B (n_20144), .Y (n_26980));
NAND2X1 g84172(.A (n_21676), .B (n_209), .Y (n_26981));
NOR2X1 g84173(.A (n_21623), .B (n_26984), .Y (n_26985));
AOI21X1 g84174(.A0 (n_18879), .A1 (n_21308), .B0 (n_21717), .Y(n_26984));
NOR2X1 g14(.A (n_636), .B (n_26992), .Y (n_26993));
OR2X1 g15_dup(.A (n_26990), .B (n_26991), .Y (n_26992));
CLKBUFX1 g84176(.A (n_26989), .Y (n_26990));
INVX4 g84177(.A (sa33[5] ), .Y (n_26989));
CLKBUFX3 g84178(.A (sa33[6] ), .Y (n_26991));
OR2X1 g15(.A (n_26990), .B (n_26991), .Y (n_26994));
OAI21X1 g84179(.A0 (n_26995), .A1 (n_26996), .B0 (n_26997), .Y(n_26998));
XOR2X1 g84180(.A (n_22954), .B (n_23694), .Y (n_26995));
MX2X1 g84181(.A (n_24306), .B (n_24512), .S0 (n_24156), .Y (n_26996));
NAND2X1 g84182(.A (n_26996), .B (n_26995), .Y (n_26997));
NAND4X1 g84183(.A (n_28601), .B (n_28602), .C (n_27003), .D(n_27004), .Y (n_27005));
OAI21X1 g84184(.A0 (n_21846), .A1 (n_18125), .B0 (n_22231), .Y(n_28602));
NAND2X1 g84185(.A (sa23[0] ), .B (n_27000), .Y (n_28601));
NAND4X1 g84186(.A (n_20419), .B (n_21038), .C (n_20264), .D(n_16185), .Y (n_27000));
INVX1 g84187(.A (n_27002), .Y (n_27003));
NAND3X1 g84188(.A (n_20385), .B (n_18902), .C (n_20270), .Y(n_27002));
OAI21X1 g84189(.A0 (n_20122), .A1 (n_19479), .B0 (n_20585), .Y(n_27004));
NAND4X1 g84190(.A (n_27010), .B (n_27011), .C (n_27012), .D(n_27014), .Y (n_27015));
NAND2X2 g84191(.A (n_27817), .B (n_27009), .Y (n_27010));
NAND4X1 g84193(.A (n_28881), .B (n_28882), .C (n_27007), .D(n_27008), .Y (n_27009));
AND2X1 g84194(.A (n_18181), .B (n_10384), .Y (n_27007));
NOR2X1 g84195(.A (n_15638), .B (n_11466), .Y (n_27008));
OAI21X1 g84196(.A0 (n_21465), .A1 (n_20328), .B0 (sa21[0] ), .Y(n_27011));
INVX1 g84197(.A (n_20880), .Y (n_27012));
NOR2X1 g84198(.A (n_27013), .B (n_21438), .Y (n_27014));
NAND2X1 g84199(.A (n_18330), .B (n_17180), .Y (n_27013));
NAND2X2 g84200(.A (n_28261), .B (n_28262), .Y (n_27018));
AOI22X1 g84201(.A0 (sa10[0] ), .A1 (n_21909), .B0 (n_20855), .B1(n_21487), .Y (n_28262));
AOI21X1 g84202(.A0 (n_28179), .A1 (n_21945), .B0 (n_21550), .Y(n_28261));
OAI21X1 g84204(.A0 (n_21259), .A1 (n_12266), .B0 (n_20102), .Y(n_27019));
OAI21X1 g84205(.A0 (n_18867), .A1 (n_28998), .B0 (n_20585), .Y(n_27020));
AND2X1 g84206(.A (n_27021), .B (n_27024), .Y (n_27025));
NAND2X1 g84207(.A (n_14173), .B (n_27023), .Y (n_27021));
NAND2X1 g84208(.A (n_27022), .B (n_27023), .Y (n_27024));
NOR2X1 g84209(.A (n_15968), .B (n_9127), .Y (n_27022));
NOR2X1 g84210(.A (n_19372), .B (n_14155), .Y (n_27023));
INVX1 g84212(.A (n_27023), .Y (n_27028));
NAND4X1 g84213(.A (n_27030), .B (n_27031), .C (n_20281), .D(n_27033), .Y (n_27034));
INVX1 g84214(.A (n_27029), .Y (n_27030));
AOI21X1 g84215(.A0 (n_21155), .A1 (n_19976), .B0 (sa32[0] ), .Y(n_27029));
AND2X1 g84216(.A (n_21693), .B (n_21573), .Y (n_27031));
INVX1 g84217(.A (n_27032), .Y (n_27033));
NAND4X1 g84218(.A (n_15603), .B (n_10239), .C (n_14997), .D(n_16618), .Y (n_27032));
NAND4X1 g84219(.A (n_27037), .B (n_27038), .C (n_27039), .D(n_27042), .Y (n_27043));
NAND2X1 g84220(.A (n_27036), .B (sa03[0] ), .Y (n_27037));
NAND4X1 g84221(.A (n_20732), .B (n_21048), .C (n_27035), .D(n_17597), .Y (n_27036));
AND2X1 g84222(.A (n_15742), .B (n_15625), .Y (n_27035));
NAND2X1 g84223(.A (n_28194), .B (n_21594), .Y (n_27038));
OAI21X1 g84224(.A0 (n_21729), .A1 (n_10304), .B0 (n_2909), .Y(n_27039));
NOR2X1 g84225(.A (n_27040), .B (n_27041), .Y (n_27042));
NAND2X1 g84226(.A (n_20772), .B (n_17756), .Y (n_27040));
NAND2X1 g84227(.A (n_18916), .B (n_16700), .Y (n_27041));
AOI21X1 g84228(.A0 (n_27046), .A1 (n_27049), .B0 (n_0), .Y (n_27051));
NAND2X1 g84229(.A (n_27044), .B (n_27045), .Y (n_27046));
NAND3X1 g84230(.A (n_16135), .B (n_19816), .C (n_17929), .Y(n_27044));
INVX1 g84231(.A (sa11[1] ), .Y (n_27045));
NOR2X1 g84232(.A (n_27047), .B (n_27048), .Y (n_27049));
NOR2X1 g84233(.A (n_12298), .B (n_17807), .Y (n_27047));
NAND3X1 g84234(.A (n_27480), .B (n_19901), .C (n_25758), .Y(n_27048));
INVX1 g84236(.A (sa11[1] ), .Y (n_20729));
NAND2X2 g84237(.A (n_27053), .B (n_27060), .Y (n_27061));
AND2X1 g84238(.A (n_21852), .B (n_22295), .Y (n_27053));
NOR2X1 g84239(.A (n_27056), .B (n_27059), .Y (n_27060));
INVX1 g84240(.A (n_27055), .Y (n_27056));
AOI21X1 g84241(.A0 (n_21458), .A1 (n_2909), .B0 (n_27054), .Y(n_27055));
AND2X1 g84242(.A (n_20024), .B (n_20610), .Y (n_27054));
OAI21X1 g84243(.A0 (n_16768), .A1 (n_28645), .B0 (n_27058), .Y(n_27059));
NAND2X1 g84244(.A (n_28692), .B (n_27057), .Y (n_27058));
INVX1 g84245(.A (n_13686), .Y (n_27057));
NAND4X1 g84247(.A (n_27066), .B (n_21386), .C (n_22311), .D(n_27067), .Y (n_27068));
AOI21X1 g84248(.A0 (n_21289), .A1 (n_21314), .B0 (n_27065), .Y(n_27066));
AOI21X1 g84249(.A0 (n_20710), .A1 (n_27063), .B0 (n_26920), .Y(n_27065));
AND2X1 g84250(.A (n_20460), .B (n_19381), .Y (n_27063));
AND2X1 g84252(.A (n_17989), .B (n_10058), .Y (n_27067));
NAND2X1 g84253(.A (n_27070), .B (n_27076), .Y (n_27077));
INVX1 g84254(.A (n_27069), .Y (n_27070));
NAND2X1 g84255(.A (n_1268), .B (n_29228), .Y (n_27069));
INVX2 g84256(.A (n_27075), .Y (n_27076));
NAND2X2 g84257(.A (n_27072), .B (n_29158), .Y (n_27075));
INVX4 g84258(.A (n_27071), .Y (n_27072));
NAND2X2 g84259(.A (n_1302), .B (n_1185), .Y (n_27071));
NAND2X2 g84264(.A (n_27083), .B (n_27084), .Y (n_27085));
AOI21X1 g84265(.A0 (sa32[0] ), .A1 (n_21666), .B0 (n_27082), .Y(n_27083));
NAND2X1 g84266(.A (n_27080), .B (n_27081), .Y (n_27082));
NAND2X1 g84267(.A (n_20624), .B (n_20055), .Y (n_27080));
AOI22X1 g84268(.A0 (n_14831), .A1 (n_16973), .B0 (n_12515), .B1(n_16974), .Y (n_27081));
AOI22X1 g84269(.A0 (n_21915), .A1 (n_21379), .B0 (n_21201), .B1(n_1397), .Y (n_27084));
NOR2X1 g84277(.A (n_15371), .B (n_15678), .Y (n_27089));
AOI21X1 g84278(.A0 (n_17790), .A1 (n_10216), .B0 (n_2917), .Y(n_27090));
NAND3X1 g84280(.A (n_27096), .B (n_27107), .C (n_27108), .Y(n_27109));
OAI21X1 g84281(.A0 (n_19104), .A1 (n_16494), .B0 (n_171), .Y(n_27096));
AOI21X1 g84282(.A0 (n_27097), .A1 (n_27100), .B0 (n_27106), .Y(n_27107));
NAND2X1 g84283(.A (n_17143), .B (n_11053), .Y (n_27097));
INVX4 g84286(.A (n_27099), .Y (n_27100));
BUFX3 g84287(.A (n_27098), .Y (n_27099));
INVX2 g84288(.A (sa31[2] ), .Y (n_27098));
NAND3X1 g84289(.A (n_27105), .B (n_13101), .C (n_5527), .Y (n_27106));
INVX1 g84290(.A (n_27104), .Y (n_27105));
AOI21X1 g84291(.A0 (n_10786), .A1 (n_10846), .B0 (n_27100), .Y(n_27104));
OAI21X1 g84293(.A0 (n_12204), .A1 (n_9995), .B0 (n_20587), .Y(n_27108));
INVX1 g84295(.A (n_27098), .Y (n_27111));
NAND4X1 g84296(.A (n_27113), .B (n_27116), .C (n_27117), .D(n_27120), .Y (n_27121));
NAND2X1 g84297(.A (n_27112), .B (sa23[0] ), .Y (n_27113));
NAND2X1 g84298(.A (n_21577), .B (n_21486), .Y (n_27112));
NAND2X1 g84299(.A (n_27114), .B (n_22231), .Y (n_27116));
NAND4X1 g84300(.A (n_21007), .B (n_18960), .C (n_18995), .D(n_19392), .Y (n_27114));
NOR2X1 g84302(.A (n_21006), .B (n_19086), .Y (n_27117));
INVX1 g84303(.A (n_27119), .Y (n_27120));
NAND3X1 g84304(.A (n_18862), .B (n_27118), .C (n_18298), .Y(n_27119));
AOI21X1 g84305(.A0 (n_28998), .A1 (n_17411), .B0 (n_16657), .Y(n_27118));
OAI21X1 g84306(.A0 (n_27127), .A1 (n_11576), .B0 (n_27131), .Y(n_27132));
AOI21X1 g84307(.A0 (n_27122), .A1 (n_1717), .B0 (n_27126), .Y(n_27127));
NAND2X1 g84308(.A (n_11728), .B (n_6549), .Y (n_27122));
INVX4 g84310(.A (n_28154), .Y (n_27124));
NOR2X1 g84312(.A (n_27124), .B (n_8863), .Y (n_27126));
CLKBUFX1 g84314(.A (sa12[2] ), .Y (n_27128));
INVX1 g84315(.A (n_27130), .Y (n_27131));
NOR2X1 g84316(.A (n_28398), .B (n_13722), .Y (n_27130));
INVX4 g84317(.A (sa12[2] ), .Y (n_27133));
INVX1 g84319(.A (n_27126), .Y (n_27135));
NAND3X1 g84320(.A (n_27138), .B (n_27139), .C (n_27142), .Y(n_27143));
NOR2X1 g84321(.A (n_27136), .B (n_27137), .Y (n_27138));
AOI21X1 g84322(.A0 (n_16724), .A1 (n_8209), .B0 (n_17377), .Y(n_27136));
NOR2X1 g84323(.A (n_10789), .B (n_8637), .Y (n_27137));
NAND2X1 g84324(.A (n_12635), .B (n_17377), .Y (n_27139));
AND2X1 g84325(.A (n_27140), .B (n_27141), .Y (n_27142));
NAND2X1 g84326(.A (n_8146), .B (n_9264), .Y (n_27140));
OR2X1 g84327(.A (n_7496), .B (n_7062), .Y (n_27141));
INVX1 g84328(.A (n_27137), .Y (n_27144));
INVX1 g84330(.A (n_27141), .Y (n_27145));
OAI21X1 g84331(.A0 (n_27147), .A1 (n_3886), .B0 (n_27156), .Y(n_27157));
NOR2X1 g84332(.A (n_13775), .B (n_17750), .Y (n_27147));
AOI21X1 g84336(.A0 (n_27152), .A1 (n_3886), .B0 (n_27155), .Y(n_27156));
INVX1 g84337(.A (n_27151), .Y (n_27152));
NAND2X1 g84338(.A (n_7867), .B (n_13834), .Y (n_27151));
NAND3X1 g84339(.A (n_27154), .B (n_18807), .C (n_18465), .Y(n_27155));
INVX1 g84340(.A (n_27153), .Y (n_27154));
NOR2X1 g84341(.A (n_9084), .B (n_9043), .Y (n_27153));
NOR2X1 g84346(.A (n_27160), .B (n_27161), .Y (n_27162));
OR2X1 g84347(.A (n_21055), .B (n_11261), .Y (n_27160));
OR2X1 g84348(.A (n_6534), .B (n_14542), .Y (n_27161));
NAND4X1 g84360(.A (n_29430), .B (n_27177), .C (n_29431), .D(n_29399), .Y (n_27185));
AOI21X1 g84361(.A0 (n_28036), .A1 (n_16754), .B0 (n_16604), .Y(n_29399));
INVX1 g84362(.A (n_15767), .Y (n_27177));
INVX1 g84363(.A (n_27179), .Y (n_29430));
NAND2X1 g84364(.A (n_17101), .B (n_27178), .Y (n_27179));
AND2X1 g84365(.A (n_5706), .B (n_11100), .Y (n_27178));
OAI21X1 g84366(.A0 (n_28040), .A1 (n_27182), .B0 (n_129), .Y(n_29431));
NAND2X1 g84368(.A (n_11611), .B (n_9799), .Y (n_27182));
NAND4X1 g84370(.A (n_27186), .B (n_27187), .C (n_27193), .D(n_27195), .Y (n_27196));
NAND2X1 g84371(.A (n_22269), .B (n_22203), .Y (n_27186));
AND2X1 g84372(.A (n_21422), .B (n_21725), .Y (n_27187));
OAI21X1 g84373(.A0 (n_27189), .A1 (n_27191), .B0 (n_27192), .Y(n_27193));
NAND2X1 g84374(.A (n_20768), .B (n_27188), .Y (n_27189));
AND2X1 g84375(.A (n_14021), .B (n_14913), .Y (n_27188));
NAND2X1 g84376(.A (n_20333), .B (n_27190), .Y (n_27191));
OAI21X1 g84377(.A0 (n_17833), .A1 (n_19889), .B0 (n_17414), .Y(n_27190));
INVX1 g84378(.A (sa11[0] ), .Y (n_27192));
INVX1 g84379(.A (n_27194), .Y (n_27195));
NAND3X1 g84380(.A (n_10508), .B (n_16533), .C (n_16982), .Y(n_27194));
INVX2 g84383(.A (sa10[4] ), .Y (n_27197));
NAND3X1 g84384(.A (n_27198), .B (n_714), .C (n_26888), .Y (n_27199));
CLKBUFX1 g84385(.A (sa10[5] ), .Y (n_27198));
CLKBUFX3 g6(.A (n_27197), .Y (n_27202));
NAND2X1 g84386(.A (n_26888), .B (n_714), .Y (n_27203));
INVX4 g84387(.A (sa10[5] ), .Y (n_27204));
NAND2X2 g84388(.A (n_27206), .B (n_27210), .Y (n_27211));
NAND4X1 g84389(.A (n_29314), .B (n_29315), .C (n_19241), .D(n_28127), .Y (n_27206));
NAND3X1 g84391(.A (n_27209), .B (n_26094), .C (n_26095), .Y(n_27210));
NOR2X1 g84392(.A (n_27207), .B (n_27208), .Y (n_27209));
NAND2X1 g84393(.A (n_26097), .B (sa13[0] ), .Y (n_27207));
INVX1 g84394(.A (n_26098), .Y (n_27208));
NAND2X1 g84396(.A (n_27213), .B (n_27217), .Y (n_27218));
NAND2X1 g84397(.A (n_18620), .B (sa13[1] ), .Y (n_27213));
OAI21X1 g84398(.A0 (n_27214), .A1 (n_27215), .B0 (n_27216), .Y(n_27217));
NAND3X1 g84399(.A (n_15316), .B (n_13291), .C (n_10801), .Y(n_27214));
NAND2X1 g84400(.A (n_11340), .B (n_9980), .Y (n_27215));
INVX1 g84401(.A (sa13[1] ), .Y (n_27216));
NAND2X2 g84403(.A (n_27220), .B (n_27222), .Y (n_27223));
INVX2 g84404(.A (n_27219), .Y (n_27220));
NAND2X1 g33_dup(.A (n_736), .B (n_26603), .Y (n_27219));
INVX1 g84405(.A (sa33[5] ), .Y (n_27222));
INVX2 g84407(.A (n_27224), .Y (n_27225));
NOR2X1 g84408(.A (n_4861), .B (n_636), .Y (n_27224));
INVX1 g84409(.A (n_27223), .Y (n_27227));
NAND2X1 g84410(.A (n_736), .B (n_26603), .Y (n_27228));
NAND2X1 g84411(.A (n_27233), .B (n_27236), .Y (n_27237));
AOI21X1 g84412(.A0 (n_17781), .A1 (n_21242), .B0 (n_27232), .Y(n_27233));
NAND2X1 g84413(.A (n_20483), .B (n_27231), .Y (n_27232));
NOR2X1 g84414(.A (n_27229), .B (n_27230), .Y (n_27231));
NOR2X1 g84415(.A (n_28692), .B (n_18050), .Y (n_27229));
NAND2X1 g84416(.A (n_14755), .B (n_19842), .Y (n_27230));
NOR2X1 g84417(.A (n_27235), .B (n_20857), .Y (n_27236));
NAND2X1 g84418(.A (n_18173), .B (n_27234), .Y (n_27235));
OR2X1 g84419(.A (n_28692), .B (n_14002), .Y (n_27234));
INVX1 g84420(.A (n_27229), .Y (n_27238));
NOR2X1 g84421(.A (n_27239), .B (n_27247), .Y (n_27248));
INVX1 g84422(.A (sa32[0] ), .Y (n_27239));
AOI21X1 g84423(.A0 (n_27241), .A1 (n_27244), .B0 (n_27246), .Y(n_27247));
NAND4X1 g84424(.A (n_27240), .B (n_15735), .C (n_12952), .D(n_15033), .Y (n_27241));
AND2X1 g84425(.A (n_12984), .B (sa32[1] ), .Y (n_27240));
NAND3X1 g84426(.A (n_14265), .B (n_14726), .C (n_27243), .Y(n_27244));
AND2X1 g84427(.A (n_16618), .B (n_27242), .Y (n_27243));
INVX1 g84428(.A (sa32[1] ), .Y (n_27242));
NAND3X1 g84429(.A (n_18169), .B (n_16209), .C (n_27245), .Y(n_27246));
AND2X1 g84430(.A (n_13011), .B (n_12477), .Y (n_27245));
AOI21X1 g84442(.A0 (n_27260), .A1 (n_27261), .B0 (n_27272), .Y(n_27273));
NAND2X1 g84443(.A (n_21464), .B (n_20137), .Y (n_27260));
INVX1 g84444(.A (n_26553), .Y (n_27261));
NAND3X1 g84445(.A (n_27265), .B (n_27268), .C (n_27271), .Y(n_27272));
NOR2X1 g84446(.A (n_27262), .B (n_27264), .Y (n_27265));
NAND2X1 g84447(.A (n_18328), .B (n_18174), .Y (n_27262));
NAND2X1 g84448(.A (n_27263), .B (n_18878), .Y (n_27264));
NAND2X1 g84449(.A (n_19617), .B (n_15074), .Y (n_27263));
NOR2X1 g84450(.A (n_27267), .B (n_26556), .Y (n_27268));
INVX1 g84451(.A (n_27266), .Y (n_27267));
NAND2X1 g84452(.A (n_11816), .B (n_10950), .Y (n_27266));
NAND2X1 g84453(.A (n_27269), .B (n_2091), .Y (n_27271));
NAND2X1 g84454(.A (n_14281), .B (n_15877), .Y (n_27269));
NAND2X1 g84464(.A (n_27282), .B (n_27288), .Y (n_27289));
NAND2X1 g84465(.A (n_13399), .B (n_12896), .Y (n_27282));
OR2X1 g84466(.A (n_28419), .B (n_27287), .Y (n_27288));
NAND2X2 g84471(.A (n_8068), .B (n_10255), .Y (n_27287));
CLKBUFX3 g84473(.A (n_27287), .Y (n_27290));
NAND3X1 g84476(.A (n_27301), .B (n_27302), .C (n_27304), .Y(n_27305));
NAND2X1 g84477(.A (n_27297), .B (n_27300), .Y (n_27301));
NAND2X1 g84478(.A (n_27294), .B (n_27296), .Y (n_27297));
INVX1 g84479(.A (n_21346), .Y (n_27294));
NOR2X1 g84480(.A (n_21), .B (n_19465), .Y (n_27296));
NAND4X1 g84482(.A (n_27298), .B (n_20480), .C (n_17843), .D(n_27617), .Y (n_27300));
AND2X1 g84483(.A (n_17155), .B (n_9597), .Y (n_27298));
NAND2X1 g84485(.A (n_21297), .B (n_21382), .Y (n_27302));
NOR2X1 g84486(.A (n_27303), .B (n_20997), .Y (n_27304));
NAND2X1 g84487(.A (n_17830), .B (n_16075), .Y (n_27303));
NAND2X1 g84488(.A (n_27307), .B (n_27310), .Y (n_27311));
AOI21X1 g84489(.A0 (n_15360), .A1 (n_5329), .B0 (n_27306), .Y(n_27307));
NOR2X1 g84490(.A (n_27483), .B (n_17377), .Y (n_27306));
NAND2X1 g84491(.A (n_27308), .B (n_27309), .Y (n_27310));
NAND3X1 g84492(.A (n_17048), .B (n_7935), .C (n_8837), .Y (n_27308));
AND2X1 g84493(.A (n_276), .B (n_9819), .Y (n_27309));
NAND2X1 g84494(.A (n_15360), .B (n_5329), .Y (n_27312));
INVX1 g84495(.A (n_27306), .Y (n_27313));
NOR2X1 g84496(.A (n_27316), .B (n_27322), .Y (n_27323));
NAND2X1 g84497(.A (n_27314), .B (n_27315), .Y (n_27316));
NAND2X1 g84498(.A (n_21834), .B (sa22[0] ), .Y (n_27314));
NAND2X1 g84499(.A (n_21354), .B (n_27786), .Y (n_27315));
NAND3X1 g84500(.A (n_27321), .B (n_21684), .C (n_17861), .Y(n_27322));
INVX1 g84501(.A (n_27320), .Y (n_27321));
NAND3X1 g84502(.A (n_20802), .B (n_27319), .C (n_19600), .Y(n_27320));
NOR2X1 g84503(.A (n_27317), .B (n_27318), .Y (n_27319));
NOR2X1 g84504(.A (n_1807), .B (n_9227), .Y (n_27317));
NOR2X1 g84505(.A (n_14589), .B (n_10685), .Y (n_27318));
NAND4X1 g84516(.A (n_27334), .B (n_27339), .C (n_27340), .D(n_27341), .Y (n_27342));
OAI21X1 g84517(.A0 (n_19466), .A1 (n_12230), .B0 (n_20680), .Y(n_27334));
NAND2X1 g84518(.A (n_27335), .B (n_17912), .Y (n_27339));
NAND2X1 g84519(.A (n_16153), .B (n_14927), .Y (n_27335));
BUFX3 g84522(.A (sa33[2] ), .Y (n_27336));
OAI21X1 g84523(.A0 (n_19460), .A1 (n_14524), .B0 (n_20518), .Y(n_27340));
NAND2X1 g84524(.A (n_4695), .B (n_11350), .Y (n_27341));
INVX1 g84526(.A (sa33[2] ), .Y (n_27344));
NOR2X1 g84527(.A (n_27346), .B (n_27352), .Y (n_27353));
NAND3X1 g84528(.A (n_25690), .B (n_21022), .C (n_27345), .Y(n_27346));
AND2X1 g84529(.A (n_10699), .B (n_19502), .Y (n_27345));
NOR2X1 g84530(.A (n_27348), .B (n_27351), .Y (n_27352));
NOR2X1 g84531(.A (n_21035), .B (n_27347), .Y (n_27348));
OR2X1 g84532(.A (sa30[0] ), .B (n_15657), .Y (n_27347));
NOR2X1 g84533(.A (n_27350), .B (n_21853), .Y (n_27351));
OR2X1 g84534(.A (n_344), .B (n_17651), .Y (n_27350));
NAND3X1 g84537(.A (n_27357), .B (n_27358), .C (n_27363), .Y(n_27364));
NOR2X1 g84538(.A (n_21145), .B (n_27356), .Y (n_27357));
NAND3X1 g84539(.A (n_20240), .B (n_19863), .C (n_27355), .Y(n_27356));
NAND2X1 g84540(.A (n_17546), .B (n_16553), .Y (n_27355));
NAND2X1 g84541(.A (n_21956), .B (n_26535), .Y (n_27358));
NAND2X1 g84542(.A (n_27362), .B (sa02[0] ), .Y (n_27363));
NAND4X1 g84543(.A (n_27361), .B (n_21248), .C (n_20663), .D(n_20950), .Y (n_27362));
NOR2X1 g84544(.A (n_27359), .B (n_27360), .Y (n_27361));
AOI21X1 g84545(.A0 (n_16254), .A1 (n_10469), .B0 (n_14474), .Y(n_27359));
INVX1 g84546(.A (n_18664), .Y (n_27360));
NOR2X1 g84547(.A (n_27365), .B (n_27372), .Y (n_27373));
INVX4 g84548(.A (sa31[3] ), .Y (n_27365));
NAND2X1 g84549(.A (n_27367), .B (n_27371), .Y (n_27372));
INVX2 g84550(.A (n_27366), .Y (n_27367));
NAND2X2 g84551(.A (n_28481), .B (n_2382), .Y (n_27366));
INVX1 g84552(.A (n_27370), .Y (n_27371));
CLKBUFX3 g84554(.A (n_27368), .Y (n_27369));
INVX1 g84555(.A (sa31[4] ), .Y (n_27368));
CLKBUFX1 g84557(.A (n_27384), .Y (n_27385));
NAND2X2 g84558(.A (n_28845), .B (n_28846), .Y (n_27384));
AOI21X1 g84559(.A0 (n_21370), .A1 (n_22251), .B0 (n_27375), .Y(n_28846));
NAND4X1 g84560(.A (n_20791), .B (n_19597), .C (n_18945), .D(n_17997), .Y (n_27375));
AOI21X1 g84561(.A0 (n_27379), .A1 (n_3546), .B0 (n_27382), .Y(n_28845));
NAND2X1 g84562(.A (n_27377), .B (n_9043), .Y (n_27379));
INVX1 g84563(.A (n_21268), .Y (n_27377));
AND2X1 g84565(.A (sa00[0] ), .B (n_27381), .Y (n_27382));
NAND4X1 g84566(.A (n_21540), .B (n_27380), .C (n_20349), .D(n_17642), .Y (n_27381));
AND2X1 g84567(.A (n_19032), .B (n_11877), .Y (n_27380));
NAND3X1 g84568(.A (n_25812), .B (n_27387), .C (n_27390), .Y(n_27391));
AOI22X1 g84569(.A0 (n_21717), .A1 (n_21082), .B0 (n_27386), .B1(n_20204), .Y (n_27387));
OR2X1 g84570(.A (n_28220), .B (n_20108), .Y (n_27386));
AOI21X1 g84571(.A0 (n_20601), .A1 (n_20397), .B0 (n_27389), .Y(n_27390));
NAND2X1 g84572(.A (n_27388), .B (n_25813), .Y (n_27389));
OR4X1 g84573(.A (n_2137), .B (n_17571), .C (n_28574), .D (n_6250), .Y(n_27388));
NAND3X1 g84574(.A (n_29376), .B (n_29377), .C (n_27401), .Y(n_23863));
NOR2X1 g84575(.A (n_27392), .B (n_27393), .Y (n_29377));
NAND3X1 g84576(.A (n_11963), .B (n_15495), .C (n_16558), .Y(n_27392));
NAND2X1 g84577(.A (n_21446), .B (n_21119), .Y (n_27393));
NAND2X1 g84578(.A (n_22267), .B (n_28128), .Y (n_29376));
OAI21X1 g84579(.A0 (n_27397), .A1 (n_27399), .B0 (n_28127), .Y(n_27401));
NAND2X1 g84580(.A (n_27396), .B (n_20764), .Y (n_27397));
AND2X1 g84581(.A (n_16573), .B (n_12212), .Y (n_27396));
NAND2X1 g84582(.A (n_20728), .B (n_27398), .Y (n_27399));
OAI21X1 g84583(.A0 (n_16569), .A1 (n_10383), .B0 (n_15708), .Y(n_27398));
NAND4X1 g84585(.A (n_27403), .B (n_27408), .C (n_27410), .D(n_27412), .Y (n_27413));
NAND2X1 g84586(.A (n_4413), .B (n_13318), .Y (n_27403));
NAND2X1 g84587(.A (n_27406), .B (n_27407), .Y (n_27408));
NAND2X1 g84588(.A (n_28857), .B (n_27405), .Y (n_27406));
NOR2X1 g84590(.A (n_7247), .B (n_4575), .Y (n_27405));
CLKBUFX3 g84591(.A (sa10[2] ), .Y (n_27407));
INVX1 g84592(.A (n_27409), .Y (n_27410));
NOR2X1 g84593(.A (n_6185), .B (n_4792), .Y (n_27409));
INVX1 g84594(.A (n_27411), .Y (n_27412));
NOR2X1 g84595(.A (n_27197), .B (n_27199), .Y (n_27411));
NAND3X1 g84598(.A (n_28598), .B (n_28599), .C (n_27420), .Y(n_27421));
OAI21X1 g84599(.A0 (n_28277), .A1 (n_28278), .B0 (n_21), .Y(n_28599));
NOR2X1 g84600(.A (n_26715), .B (n_26716), .Y (n_28598));
OAI21X1 g84601(.A0 (n_27418), .A1 (n_27419), .B0 (sa33[0] ), .Y(n_27420));
NAND2X1 g84602(.A (n_20031), .B (n_20208), .Y (n_27418));
NAND2X1 g84603(.A (n_18524), .B (n_14613), .Y (n_27419));
NAND3X1 g84604(.A (n_27422), .B (n_27423), .C (n_27428), .Y(n_27429));
OAI21X1 g84605(.A0 (n_19422), .A1 (n_14088), .B0 (n_27481), .Y(n_27422));
NOR2X1 g84606(.A (n_17396), .B (n_16536), .Y (n_27423));
AND2X1 g84607(.A (n_27427), .B (n_17099), .Y (n_27428));
AOI21X1 g84608(.A0 (n_12298), .A1 (n_16169), .B0 (n_27426), .Y(n_27427));
NAND2X1 g84609(.A (n_8952), .B (n_27425), .Y (n_27426));
INVX1 g84610(.A (n_27424), .Y (n_27425));
NOR2X1 g84611(.A (n_15800), .B (n_3653), .Y (n_27424));
NAND4X1 g84612(.A (n_27430), .B (n_27432), .C (n_27435), .D(n_27440), .Y (n_27441));
NAND2X1 g84613(.A (n_719), .B (n_6462), .Y (n_27430));
INVX1 g84614(.A (n_27431), .Y (n_27432));
NOR2X1 g84615(.A (n_6462), .B (n_2305), .Y (n_27431));
NAND2X1 g84616(.A (n_5530), .B (n_27434), .Y (n_27435));
INVX2 g84617(.A (n_27433), .Y (n_27434));
CLKBUFX1 g84618(.A (sa21[3] ), .Y (n_27433));
NAND2X1 g84619(.A (n_27439), .B (n_27433), .Y (n_27440));
INVX1 g84620(.A (n_27438), .Y (n_27439));
INVX1 g84621(.A (n_27437), .Y (n_27438));
INVX1 g84622(.A (n_27436), .Y (n_27437));
NAND2X1 g84623(.A (n_457), .B (n_342), .Y (n_27436));
OAI21X1 g84624(.A0 (n_27442), .A1 (n_27447), .B0 (sa13[1] ), .Y(n_27448));
AOI21X1 g84625(.A0 (n_11562), .A1 (n_12686), .B0 (n_15708), .Y(n_27442));
NAND3X1 g84626(.A (n_27446), .B (n_27445), .C (n_29397), .Y(n_27447));
NAND2X1 g84627(.A (n_7903), .B (n_6941), .Y (n_29397));
INVX1 g84628(.A (n_27444), .Y (n_27445));
NOR2X1 g84629(.A (n_6052), .B (n_4204), .Y (n_27444));
OR2X1 g84630(.A (n_11215), .B (n_10782), .Y (n_27446));
INVX1 g84631(.A (sa13[1] ), .Y (n_27449));
INVX1 g84632(.A (n_27446), .Y (n_27450));
NAND3X1 g84633(.A (n_27451), .B (n_27457), .C (n_27458), .Y(n_27459));
NAND2X1 g84634(.A (n_21812), .B (sa02[0] ), .Y (n_27451));
OAI21X1 g84635(.A0 (n_27453), .A1 (n_27455), .B0 (n_27456), .Y(n_27457));
NAND3X1 g84636(.A (n_21179), .B (n_27452), .C (n_19665), .Y(n_27453));
AND2X1 g84637(.A (n_19290), .B (n_14760), .Y (n_27452));
NAND2X1 g84638(.A (n_20484), .B (n_27454), .Y (n_27455));
AND2X1 g84639(.A (n_15280), .B (n_21227), .Y (n_27454));
INVX1 g84640(.A (sa02[0] ), .Y (n_27456));
INVX1 g84641(.A (n_21803), .Y (n_27458));
NAND4X1 g84642(.A (n_27463), .B (n_27464), .C (n_27465), .D(n_27467), .Y (n_27468));
OAI21X1 g84643(.A0 (n_27460), .A1 (n_27462), .B0 (sa13[0] ), .Y(n_27463));
NAND2X1 g84644(.A (n_21057), .B (n_20300), .Y (n_27460));
NAND2X1 g84645(.A (n_27461), .B (n_8301), .Y (n_27462));
NOR2X1 g84646(.A (n_18403), .B (n_17998), .Y (n_27461));
NAND2X1 g84647(.A (n_21371), .B (n_27526), .Y (n_27464));
OAI21X1 g84648(.A0 (n_21266), .A1 (n_8821), .B0 (n_378), .Y(n_27465));
INVX1 g84649(.A (n_27466), .Y (n_27467));
NAND4X1 g84650(.A (n_20183), .B (n_18224), .C (n_20100), .D(n_16842), .Y (n_27466));
NAND2X1 g84652(.A (n_27479), .B (sa11[1] ), .Y (n_27480));
NAND2X1 g84653(.A (n_27474), .B (n_27478), .Y (n_27479));
NOR2X1 g84654(.A (n_27470), .B (n_27473), .Y (n_27474));
AOI21X1 g84655(.A0 (n_8148), .A1 (n_7027), .B0 (n_9819), .Y(n_27470));
NAND3X1 g84656(.A (n_5853), .B (n_14506), .C (n_27472), .Y (n_27473));
INVX1 g84657(.A (n_27471), .Y (n_27472));
NOR2X1 g84658(.A (n_7496), .B (n_4199), .Y (n_27471));
AND2X1 g84659(.A (n_27475), .B (n_27483), .Y (n_27478));
NAND2X1 g84660(.A (n_8378), .B (n_17414), .Y (n_27475));
INVX1 g84663(.A (sa11[1] ), .Y (n_27481));
INVX2 g84665(.A (n_27596), .Y (n_27483));
XOR2X1 g84666(.A (n_27488), .B (n_27490), .Y (n_27491));
INVX2 g84667(.A (n_27487), .Y (n_27488));
NAND2X2 g84668(.A (n_27485), .B (n_27486), .Y (n_27487));
NAND2X1 g84669(.A (n_26092), .B (n_28900), .Y (n_27485));
OR2X1 g84671(.A (n_26092), .B (n_28900), .Y (n_27486));
MX2X1 g84672(.A (n_25537), .B (n_27489), .S0 (n_25536), .Y (n_27490));
INVX1 g84673(.A (n_25537), .Y (n_27489));
NAND3X1 g84674(.A (n_27494), .B (n_27502), .C (n_27503), .Y(n_27504));
NAND2X1 g84675(.A (n_27492), .B (n_27493), .Y (n_27494));
NAND2X1 g84676(.A (n_20617), .B (n_12054), .Y (n_27492));
CLKBUFX1 g84677(.A (sa00[2] ), .Y (n_27493));
AOI21X1 g84678(.A0 (n_16688), .A1 (n_19170), .B0 (n_27501), .Y(n_27502));
NAND2X1 g84679(.A (n_27495), .B (n_27500), .Y (n_27501));
AOI21X1 g84680(.A0 (n_10581), .A1 (n_19934), .B0 (n_18164), .Y(n_27495));
AOI21X1 g84681(.A0 (n_27505), .A1 (n_16434), .B0 (n_17753), .Y(n_27500));
NAND2X1 g84684(.A (n_5006), .B (n_4709), .Y (n_27496));
AOI22X1 g84686(.A0 (n_1991), .A1 (n_13961), .B0 (n_18671), .B1(n_20862), .Y (n_27503));
INVX1 g84687(.A (n_27496), .Y (n_27505));
NAND2X1 g84692(.A (n_20987), .B (n_19831), .Y (n_27508));
NAND3X1 g84693(.A (n_20512), .B (n_18520), .C (n_27509), .Y(n_27510));
NOR2X1 g84694(.A (n_9243), .B (n_17908), .Y (n_27509));
MX2X1 g84695(.A (n_27519), .B (n_27520), .S0 (n_27521), .Y (n_27522));
NAND4X1 g84696(.A (n_27514), .B (n_27513), .C (n_27517), .D(n_27518), .Y (n_27519));
OAI21X1 g84697(.A0 (n_21432), .A1 (n_20746), .B0 (sa13[0] ), .Y(n_27513));
INVX1 g84698(.A (n_21995), .Y (n_27514));
AND2X1 g84699(.A (n_21072), .B (n_27516), .Y (n_27517));
INVX1 g84700(.A (n_27515), .Y (n_27516));
NAND3X1 g84701(.A (n_11522), .B (n_16559), .C (n_15190), .Y(n_27515));
INVX1 g84702(.A (n_20715), .Y (n_27518));
INVX1 g84703(.A (n_27519), .Y (n_27520));
NAND3X1 g84704(.A (n_26495), .B (n_26498), .C (n_26501), .Y(n_27521));
NOR2X1 g84705(.A (n_27523), .B (n_27524), .Y (n_27525));
INVX1 g84706(.A (n_27513), .Y (n_27523));
NAND3X1 g84707(.A (n_27514), .B (n_27517), .C (n_27518), .Y(n_27524));
NAND4X1 g84708(.A (n_27532), .B (n_27533), .C (n_27534), .D(n_27536), .Y (n_27537));
NAND2X1 g84709(.A (n_27526), .B (n_27531), .Y (n_27532));
INVX1 g84710(.A (sa13[0] ), .Y (n_27526));
NAND3X1 g84711(.A (n_29405), .B (n_29406), .C (n_20598), .Y(n_27531));
INVX1 g84712(.A (n_27529), .Y (n_29406));
NAND4X1 g84713(.A (n_27527), .B (n_18227), .C (n_14014), .D(n_27528), .Y (n_27529));
INVX1 g84714(.A (n_13552), .Y (n_27527));
INVX1 g84715(.A (n_17337), .Y (n_27528));
OAI21X1 g84716(.A0 (n_21184), .A1 (n_20359), .B0 (sa13[0] ), .Y(n_27533));
INVX1 g84717(.A (n_20940), .Y (n_27534));
NOR2X1 g84718(.A (n_27535), .B (n_21445), .Y (n_27536));
NAND2X1 g84719(.A (n_16909), .B (n_19033), .Y (n_27535));
NAND4X1 g84734(.A (n_27556), .B (n_27557), .C (n_27558), .D(n_27560), .Y (n_27561));
OAI21X1 g84735(.A0 (n_27553), .A1 (n_27554), .B0 (n_21396), .Y(n_27556));
NAND3X1 g84736(.A (n_25796), .B (n_27552), .C (n_13016), .Y(n_27553));
AND2X1 g84737(.A (n_12607), .B (n_6205), .Y (n_27552));
NAND2X1 g84738(.A (n_12969), .B (n_14047), .Y (n_27554));
OAI21X1 g84740(.A0 (n_19454), .A1 (n_14250), .B0 (n_3538), .Y(n_27557));
OAI21X1 g84741(.A0 (n_19182), .A1 (n_11993), .B0 (n_29062), .Y(n_27558));
INVX1 g84742(.A (n_27559), .Y (n_27560));
NOR2X1 g84743(.A (n_8185), .B (n_9368), .Y (n_27559));
NAND3X1 g84744(.A (n_27565), .B (n_27566), .C (n_27573), .Y(n_27574));
NOR2X1 g84745(.A (n_21141), .B (n_27564), .Y (n_27565));
NAND2X1 g84746(.A (n_20706), .B (n_27563), .Y (n_27564));
AOI21X1 g84747(.A0 (n_17542), .A1 (n_13423), .B0 (n_27562), .Y(n_27563));
INVX1 g84748(.A (n_19845), .Y (n_27562));
NAND2X1 g84749(.A (n_21954), .B (n_26405), .Y (n_27566));
NAND2X1 g84750(.A (n_28207), .B (n_27572), .Y (n_27573));
NAND4X1 g84753(.A (n_27571), .B (n_21246), .C (n_20650), .D(n_27693), .Y (n_27572));
NOR2X1 g84754(.A (n_27569), .B (n_27570), .Y (n_27571));
INVX1 g84755(.A (n_18659), .Y (n_27569));
AOI21X1 g84756(.A0 (n_17668), .A1 (n_19690), .B0 (n_19364), .Y(n_27570));
NAND2X1 g84767(.A (n_27585), .B (n_27588), .Y (n_27589));
NAND2X1 g84768(.A (n_17234), .B (n_19398), .Y (n_27585));
OAI21X1 g84769(.A0 (n_27586), .A1 (n_27587), .B0 (sa12[1] ), .Y(n_27588));
NAND2X1 g84770(.A (n_13404), .B (n_12214), .Y (n_27586));
NAND4X1 g84771(.A (n_15627), .B (n_14358), .C (n_11287), .D (n_9547),.Y (n_27587));
INVX2 g84773(.A (n_27595), .Y (n_27596));
OR2X1 g84774(.A (n_28744), .B (n_27594), .Y (n_27595));
NAND3X1 g84776(.A (n_27593), .B (n_920), .C (n_95), .Y (n_27594));
INVX2 g84777(.A (n_27592), .Y (n_27593));
INVX2 g84778(.A (sa11[5] ), .Y (n_27592));
NAND2X1 g84780(.A (n_920), .B (n_95), .Y (n_27598));
INVX1 g84781(.A (n_27593), .Y (n_27599));
NAND3X1 g84782(.A (n_27606), .B (n_27607), .C (n_27609), .Y(n_27610));
NOR2X1 g84783(.A (n_27600), .B (n_27605), .Y (n_27606));
NAND2X1 g84784(.A (n_11714), .B (n_13508), .Y (n_27600));
AOI21X1 g84785(.A0 (n_27601), .A1 (n_27603), .B0 (n_27604), .Y(n_27605));
NAND2X1 g84786(.A (n_7312), .B (n_8742), .Y (n_27601));
NAND2X2 g84788(.A (n_2301), .B (n_3820), .Y (n_27603));
INVX2 g84789(.A (sa13[2] ), .Y (n_27604));
NAND2X1 g84790(.A (n_9905), .B (n_16787), .Y (n_27607));
INVX1 g84791(.A (n_27608), .Y (n_27609));
NOR2X1 g52_dup(.A (n_18785), .B (n_7399), .Y (n_27608));
NOR2X1 g84792(.A (n_18785), .B (n_7399), .Y (n_27611));
INVX1 g84793(.A (n_27603), .Y (n_27612));
OAI21X1 g84796(.A0 (n_27615), .A1 (n_27616), .B0 (n_27617), .Y(n_27618));
NAND2X1 g84797(.A (n_27614), .B (n_20690), .Y (n_27615));
AND2X1 g84798(.A (n_18910), .B (n_9108), .Y (n_27614));
NAND3X1 g84799(.A (n_20904), .B (n_16669), .C (n_26228), .Y(n_27616));
INVX1 g84800(.A (sa33[0] ), .Y (n_27617));
NAND2X1 g84801(.A (n_26012), .B (n_21292), .Y (n_27619));
NOR2X1 g84802(.A (n_27508), .B (n_27510), .Y (n_27620));
NAND2X1 g84805(.A (n_21400), .B (n_20580), .Y (n_27622));
NAND2X1 g84806(.A (n_25901), .B (n_25902), .Y (n_27623));
INVX1 g84807(.A (sa12[0] ), .Y (n_27624));
INVX1 g84811(.A (n_20923), .Y (n_27627));
INVX1 g23(.A (n_27645), .Y (n_27646));
NAND2X1 g84820(.A (n_27643), .B (n_28441), .Y (n_27645));
INVX1 g84821(.A (n_27642), .Y (n_27643));
NAND2X1 g84822(.A (n_27640), .B (n_27641), .Y (n_27642));
AND2X1 g84823(.A (n_28779), .B (n_26185), .Y (n_27640));
CLKBUFX3 g84824(.A (sa12[4] ), .Y (n_27641));
NAND2X1 g84829(.A (n_28596), .B (n_28597), .Y (n_27655));
AOI21X1 g84830(.A0 (n_10972), .A1 (n_11850), .B0 (n_27650), .Y(n_28597));
AND2X1 g84831(.A (n_11118), .B (n_11850), .Y (n_27650));
NAND2X1 g84832(.A (n_27652), .B (n_27718), .Y (n_28596));
NAND2X1 g26(.A (n_8619), .B (n_10112), .Y (n_27652));
INVX1 g84834(.A (n_27650), .Y (n_27656));
NAND4X1 g84835(.A (n_27657), .B (n_27658), .C (n_27659), .D(n_27665), .Y (n_27666));
NAND2X1 g84836(.A (n_26535), .B (n_28283), .Y (n_27657));
OAI21X1 g84837(.A0 (n_21586), .A1 (n_20464), .B0 (sa02[0] ), .Y(n_27658));
OAI21X1 g84838(.A0 (n_21264), .A1 (n_18721), .B0 (n_1196), .Y(n_27659));
INVX1 g84839(.A (n_27664), .Y (n_27665));
NAND4X1 g84840(.A (n_27660), .B (n_27661), .C (n_15269), .D(n_27663), .Y (n_27664));
NAND2X1 g84841(.A (n_19803), .B (n_16362), .Y (n_27660));
AOI22X1 g84842(.A0 (n_16553), .A1 (n_12783), .B0 (n_17558), .B1(n_19651), .Y (n_27661));
NAND3X1 g84844(.A (n_16362), .B (n_17706), .C (n_14681), .Y(n_27663));
INVX2 g84845(.A (n_11298), .Y (n_27671));
OR2X1 g84846(.A (n_3338), .B (n_27669), .Y (n_11298));
NAND3X1 g84848(.A (n_528), .B (n_27668), .C (n_25783), .Y (n_27669));
CLKBUFX3 g84849(.A (sa30[5] ), .Y (n_27668));
INVX2 g84850(.A (n_27672), .Y (n_27673));
NAND2X2 g84851(.A (n_25783), .B (n_528), .Y (n_27672));
INVX2 g84852(.A (n_27668), .Y (n_27674));
NOR2X1 g84853(.A (n_27677), .B (n_27682), .Y (n_27683));
NAND2X1 g84854(.A (n_27675), .B (n_27676), .Y (n_27677));
NAND2X1 g84855(.A (n_21629), .B (n_27786), .Y (n_27675));
OAI21X1 g34(.A0 (n_20404), .A1 (n_19643), .B0 (n_19414), .Y(n_27676));
NAND2X1 g84856(.A (n_27678), .B (n_27681), .Y (n_27682));
NAND2X1 g84857(.A (sa22[0] ), .B (n_22173), .Y (n_27678));
NAND2X1 g35(.A (n_27679), .B (n_20574), .Y (n_27681));
NAND2X1 g84858(.A (n_19848), .B (n_26246), .Y (n_27679));
NAND3X1 g84860(.A (n_27691), .B (n_27692), .C (n_27696), .Y(n_27697));
NAND2X1 g84861(.A (n_27687), .B (n_27690), .Y (n_27691));
NAND2X1 g84862(.A (n_17616), .B (n_27686), .Y (n_27687));
NAND2X1 g84864(.A (n_17776), .B (n_16049), .Y (n_27684));
NAND2X2 g84865(.A (n_3204), .B (n_4934), .Y (n_27686));
CLKBUFX1 g55(.A (n_27688), .Y (n_27690));
INVX8 g84867(.A (sa01[2] ), .Y (n_27688));
OR2X1 g84868(.A (n_27690), .B (n_13370), .Y (n_27692));
AND2X1 g84869(.A (n_27693), .B (n_27695), .Y (n_27696));
NAND2X1 g84870(.A (n_10094), .B (n_13037), .Y (n_27693));
INVX1 g84871(.A (n_27694), .Y (n_27695));
AND2X1 g84872(.A (n_12599), .B (n_27688), .Y (n_27694));
NAND2X2 g84874(.A (n_27701), .B (n_27705), .Y (n_27706));
NOR2X1 g84875(.A (n_27699), .B (n_27700), .Y (n_27701));
INVX1 g84876(.A (n_21867), .Y (n_27699));
NOR2X1 g84877(.A (n_27456), .B (n_22179), .Y (n_27700));
AOI21X1 g84878(.A0 (n_21228), .A1 (n_1196), .B0 (n_27704), .Y(n_27705));
OAI21X1 g84879(.A0 (n_27702), .A1 (n_1196), .B0 (n_27703), .Y(n_27704));
AND2X1 g84880(.A (n_19330), .B (n_16830), .Y (n_27702));
MX2X1 g84881(.A (n_15543), .B (n_13690), .S0 (n_14474), .Y (n_27703));
OR2X1 g84882(.A (n_27707), .B (n_27714), .Y (n_27715));
NOR2X1 g84883(.A (n_7453), .B (n_7787), .Y (n_27707));
NAND2X1 g84884(.A (n_27708), .B (n_27713), .Y (n_27714));
NAND2X1 g84885(.A (n_4301), .B (n_8865), .Y (n_27708));
NOR2X1 g84886(.A (n_27711), .B (n_27712), .Y (n_27713));
NAND2X1 g84887(.A (n_27709), .B (n_27710), .Y (n_27711));
OR2X1 g84888(.A (n_27223), .B (n_27225), .Y (n_27709));
OR2X1 g84889(.A (n_4861), .B (n_4643), .Y (n_27710));
NOR2X1 g84890(.A (n_13490), .B (n_4271), .Y (n_27712));
INVX1 g84891(.A (n_27709), .Y (n_27716));
NAND2X1 g84892(.A (n_27720), .B (n_27725), .Y (n_27726));
NAND4X1 g84893(.A (n_27717), .B (n_25999), .C (n_26007), .D(n_20068), .Y (n_27720));
AND2X1 g84894(.A (n_14819), .B (n_8251), .Y (n_27717));
INVX2 g84896(.A (sa12[1] ), .Y (n_27718));
NAND4X1 g84897(.A (n_27723), .B (n_27724), .C (n_8403), .D (n_27718),.Y (n_27725));
NOR2X1 g84898(.A (n_8477), .B (n_27722), .Y (n_27723));
NAND2X1 g84899(.A (n_11122), .B (n_6814), .Y (n_27722));
NAND2X1 g84901(.A (n_10351), .B (n_4875), .Y (n_27724));
NAND4X1 g84902(.A (n_27729), .B (n_27730), .C (n_27732), .D(n_21897), .Y (n_28802));
OAI21X1 g84903(.A0 (n_27727), .A1 (n_27728), .B0 (sa10[0] ), .Y(n_27729));
NAND2X1 g84904(.A (n_21049), .B (n_26853), .Y (n_27727));
NAND2X1 g84905(.A (n_20285), .B (n_26855), .Y (n_27728));
OAI21X1 g84906(.A0 (n_21257), .A1 (n_8901), .B0 (n_17933), .Y(n_27730));
INVX1 g84907(.A (n_27731), .Y (n_27732));
NAND3X1 g84908(.A (n_26858), .B (n_20052), .C (n_17761), .Y(n_27731));
NAND2X2 g84910(.A (n_27736), .B (n_27740), .Y (n_27741));
OAI21X1 g84911(.A0 (n_21858), .A1 (w3[0] ), .B0 (n_27735), .Y(n_27736));
OR2X1 g84913(.A (n_22372), .B (n_22063), .Y (n_27735));
NOR2X1 g84914(.A (n_21727), .B (n_27739), .Y (n_27740));
INVX1 g84915(.A (n_27738), .Y (n_27739));
AOI21X1 g84916(.A0 (n_27737), .A1 (w3[1] ), .B0 (n_16981), .Y(n_27738));
NAND2X1 g84917(.A (n_20503), .B (n_20755), .Y (n_27737));
NAND2X1 g84919(.A (n_27751), .B (n_27752), .Y (n_27753));
AOI22X1 g84920(.A0 (n_16434), .A1 (n_4488), .B0 (n_27745), .B1(n_9084), .Y (n_27751));
INVX1 g84921(.A (n_27744), .Y (n_27745));
NAND2X2 g84922(.A (n_6997), .B (n_8499), .Y (n_27744));
INVX8 g84926(.A (n_27746), .Y (n_27747));
INVX4 g84927(.A (sa00[3] ), .Y (n_27746));
NAND2X1 g84928(.A (n_8674), .B (n_2111), .Y (n_27752));
INVX2 g84932(.A (n_27747), .Y (n_27757));
INVX1 g84953(.A (n_27783), .Y (n_27784));
NAND4X1 g84954(.A (n_27778), .B (n_27780), .C (n_27782), .D(n_15272), .Y (n_27783));
NAND2X1 g84955(.A (n_16199), .B (n_17912), .Y (n_27778));
AND2X1 g84956(.A (n_8523), .B (n_27779), .Y (n_27780));
NAND2X1 g84957(.A (n_10101), .B (n_4367), .Y (n_27779));
INVX1 g84958(.A (n_27781), .Y (n_27782));
AOI21X1 g84959(.A0 (n_10109), .A1 (n_9927), .B0 (n_1424), .Y(n_27781));
CLKBUFX1 g84960(.A (n_27794), .Y (n_27795));
NAND2X1 g84961(.A (n_27788), .B (n_27793), .Y (n_27794));
AOI21X1 g84962(.A0 (n_27785), .A1 (n_27786), .B0 (n_27787), .Y(n_27788));
NAND4X1 g84963(.A (n_21012), .B (n_18961), .C (n_19394), .D(n_19002), .Y (n_27785));
INVX1 g84964(.A (sa22[0] ), .Y (n_27786));
AOI21X1 g84965(.A0 (n_21579), .A1 (n_21276), .B0 (n_27786), .Y(n_27787));
NOR2X1 g84966(.A (n_27789), .B (n_27792), .Y (n_27793));
NAND2X1 g84967(.A (n_20245), .B (n_15037), .Y (n_27789));
NAND4X1 g84968(.A (n_21173), .B (n_18861), .C (n_27791), .D(n_18534), .Y (n_27792));
AOI21X1 g84969(.A0 (n_13926), .A1 (n_20325), .B0 (n_27790), .Y(n_27791));
INVX1 g84970(.A (n_17189), .Y (n_27790));
NAND3X1 g84971(.A (n_27798), .B (n_27800), .C (n_27805), .Y(n_27806));
NOR2X1 g84972(.A (n_27797), .B (n_22145), .Y (n_27798));
AOI21X1 g84973(.A0 (n_18788), .A1 (n_16534), .B0 (n_27160), .Y(n_27797));
INVX1 g84974(.A (n_27799), .Y (n_27800));
AOI21X1 g84975(.A0 (n_21137), .A1 (n_20947), .B0 (sa20[0] ), .Y(n_27799));
NOR2X1 g84976(.A (n_27804), .B (n_21782), .Y (n_27805));
OAI21X1 g84977(.A0 (n_17329), .A1 (n_21314), .B0 (n_27803), .Y(n_27804));
AND2X1 g84978(.A (n_27801), .B (n_27802), .Y (n_27803));
NAND2X1 g84979(.A (n_6748), .B (n_11694), .Y (n_27801));
NAND2X1 g84980(.A (n_4427), .B (n_14082), .Y (n_27802));
INVX1 g84981(.A (n_27801), .Y (n_27807));
NAND4X1 g84982(.A (n_22240), .B (n_27811), .C (n_27814), .D(n_21043), .Y (n_27815));
INVX1 g84983(.A (n_27810), .Y (n_27811));
NAND3X1 g84984(.A (n_21000), .B (n_8871), .C (n_27809), .Y (n_27810));
OR4X1 g84985(.A (n_2076), .B (n_14624), .C (n_6554), .D (n_1513), .Y(n_27809));
NAND2X1 g84987(.A (n_27812), .B (n_344), .Y (n_27814));
NAND4X1 g84988(.A (n_20298), .B (n_19540), .C (n_19370), .D(n_12253), .Y (n_27812));
NAND3X1 g84991(.A (n_19255), .B (n_19350), .C (n_15379), .Y(n_27816));
INVX4 g84992(.A (sa21[0] ), .Y (n_27817));
NAND3X1 g84993(.A (n_27966), .B (n_27819), .C (n_27822), .Y(n_27823));
OAI21X1 g84995(.A0 (n_18290), .A1 (n_5813), .B0 (n_21396), .Y(n_27819));
OR2X1 g84996(.A (n_2342), .B (n_27821), .Y (n_27822));
NOR2X1 g84998(.A (n_17900), .B (n_14962), .Y (n_27821));
NAND4X1 g84999(.A (n_27825), .B (n_27829), .C (n_27830), .D(n_27833), .Y (n_27834));
OAI21X1 g85000(.A0 (n_27622), .A1 (n_27623), .B0 (n_27624), .Y(n_27825));
AND2X1 g85001(.A (n_27627), .B (n_27828), .Y (n_27829));
NAND2X1 g85002(.A (n_27826), .B (n_20018), .Y (n_27828));
INVX1 g85003(.A (n_20293), .Y (n_27826));
OAI21X1 g85005(.A0 (n_21183), .A1 (n_20358), .B0 (sa12[0] ), .Y(n_27830));
NOR2X1 g85006(.A (n_27831), .B (n_25907), .Y (n_27833));
INVX1 g85007(.A (n_18095), .Y (n_27831));
NAND2X1 g85009(.A (n_27841), .B (n_27846), .Y (n_27847));
NOR2X1 g85010(.A (n_27836), .B (n_27840), .Y (n_27841));
NAND2X1 g85011(.A (n_17103), .B (n_27835), .Y (n_27836));
AND2X1 g85012(.A (n_6921), .B (n_10988), .Y (n_27835));
AOI21X1 g85013(.A0 (n_28841), .A1 (n_28842), .B0 (sa32[1] ), .Y(n_27840));
INVX1 g85014(.A (n_14184), .Y (n_28842));
INVX1 g85015(.A (n_18694), .Y (n_28841));
NOR2X1 g85017(.A (n_27842), .B (n_27845), .Y (n_27846));
AOI21X1 g85018(.A0 (n_10317), .A1 (n_16674), .B0 (n_19486), .Y(n_27842));
OAI21X1 g85019(.A0 (n_27843), .A1 (n_2663), .B0 (n_27844), .Y(n_27845));
AND2X1 g85020(.A (n_9797), .B (n_9683), .Y (n_27843));
NAND2X1 g85021(.A (n_11782), .B (n_26270), .Y (n_27844));
NOR2X1 g85022(.A (n_27849), .B (n_27855), .Y (n_27856));
NAND3X1 g85023(.A (n_21409), .B (n_20667), .C (n_27848), .Y(n_27849));
AND2X1 g85024(.A (n_12159), .B (n_19542), .Y (n_27848));
AOI21X1 g85025(.A0 (n_27850), .A1 (n_27851), .B0 (n_27854), .Y(n_27855));
INVX1 g85026(.A (n_21036), .Y (n_27850));
NOR2X1 g85027(.A (sa31[0] ), .B (n_15707), .Y (n_27851));
NOR2X1 g85028(.A (n_27853), .B (n_21861), .Y (n_27854));
OR2X1 g85029(.A (n_21717), .B (n_17640), .Y (n_27853));
XOR2X1 g85045(.A (n_27873), .B (n_27875), .Y (n_27876));
INVX1 g85046(.A (n_27872), .Y (n_27873));
MX2X1 g85047(.A (n_26297), .B (n_26298), .S0 (n_26303), .Y (n_27872));
MX2X1 g28(.A (n_27874), .B (n_23055), .S0 (n_23932), .Y (n_27875));
INVX1 g85048(.A (n_23055), .Y (n_27874));
NAND3X1 g85056(.A (n_27889), .B (n_27890), .C (n_27891), .Y(n_27892));
NAND3X1 g85057(.A (n_27885), .B (n_27887), .C (n_25926), .Y(n_27889));
INVX1 g85058(.A (n_27884), .Y (n_27885));
MX2X1 g85059(.A (n_24899), .B (n_24898), .S0 (n_24860), .Y (n_27884));
INVX1 g85060(.A (n_27886), .Y (n_27887));
NAND2X1 g85061(.A (n_24530), .B (n_24353), .Y (n_27886));
NAND3X1 g85063(.A (n_27884), .B (n_27886), .C (n_25926), .Y(n_27890));
OR2X1 g85064(.A (n_13846), .B (n_2544), .Y (n_27891));
NOR2X1 g85065(.A (n_27893), .B (n_27898), .Y (n_27899));
INVX1 g85066(.A (sa13[3] ), .Y (n_27893));
NAND2X1 g23_dup(.A (n_27904), .B (n_27897), .Y (n_27898));
CLKBUFX3 g85068(.A (sa13[4] ), .Y (n_27894));
INVX1 g85069(.A (n_27896), .Y (n_27897));
NAND2X2 g85070(.A (n_3251), .B (n_3252), .Y (n_27896));
NAND2X1 g85071(.A (n_27904), .B (n_27897), .Y (n_27900));
INVX2 g85073(.A (n_27893), .Y (n_27901));
INVX4 g85075(.A (n_27894), .Y (n_27904));
NAND4X1 g85076(.A (n_27905), .B (n_27906), .C (n_27911), .D(n_27917), .Y (n_27918));
OAI21X1 g85077(.A0 (n_25643), .A1 (n_25642), .B0 (sa21[0] ), .Y(n_27905));
NAND2X1 g85078(.A (n_21357), .B (n_27817), .Y (n_27906));
NAND2X1 g85079(.A (n_27909), .B (n_27910), .Y (n_27911));
NAND2X1 g85080(.A (n_27907), .B (n_27908), .Y (n_27909));
INVX1 g83(.A (n_19188), .Y (n_27907));
NOR3X1 g85081(.A (n_10598), .B (n_9721), .C (n_17045), .Y (n_27908));
INVX1 g87(.A (sa21[1] ), .Y (n_27910));
NOR2X1 g85082(.A (n_27916), .B (n_20491), .Y (n_27917));
NAND2X1 g85083(.A (n_27912), .B (n_27915), .Y (n_27916));
INVX1 g88(.A (n_18086), .Y (n_27912));
AOI21X1 g85084(.A0 (n_27913), .A1 (n_27914), .B0 (n_15047), .Y(n_27915));
NOR2X1 g85085(.A (n_14026), .B (n_29171), .Y (n_27913));
NOR2X1 g85086(.A (n_21396), .B (n_29014), .Y (n_27914));
INVX1 g85087(.A (n_27914), .Y (n_27919));
NAND2X1 g85107(.A (n_27946), .B (n_27949), .Y (n_27950));
INVX4 g85108(.A (n_27945), .Y (n_27946));
CLKBUFX3 g85109(.A (n_27944), .Y (n_27945));
NAND4X1 g85110(.A (n_27939), .B (n_27940), .C (n_27942), .D(n_27943), .Y (n_27944));
AOI21X1 g85111(.A0 (n_27816), .A1 (n_27817), .B0 (n_27823), .Y(n_27939));
NAND2X1 g85112(.A (n_357), .B (n_28028), .Y (n_27940));
NAND2X1 g85113(.A (n_26646), .B (n_27941), .Y (n_27942));
AND2X1 g85114(.A (sa21[1] ), .B (n_27817), .Y (n_27941));
OAI21X1 g85115(.A0 (n_19556), .A1 (n_19480), .B0 (sa21[1] ), .Y(n_27943));
INVX2 g85116(.A (n_27948), .Y (n_27949));
INVX4 g85117(.A (n_27947), .Y (n_27948));
NAND3X1 g85118(.A (n_26898), .B (n_26159), .C (n_26160), .Y(n_27947));
NAND4X1 g85120(.A (n_27019), .B (n_27025), .C (n_27020), .D(n_27953), .Y (n_27954));
NOR2X1 g85121(.A (n_27951), .B (n_27952), .Y (n_27953));
NOR2X1 g85122(.A (n_2052), .B (n_9116), .Y (n_27951));
NOR2X1 g85123(.A (n_11277), .B (n_13993), .Y (n_27952));
NAND2X1 g85124(.A (n_27955), .B (n_27956), .Y (n_27957));
NAND2X1 g85125(.A (n_21360), .B (n_22231), .Y (n_27955));
NAND2X1 g85126(.A (n_21835), .B (sa23[0] ), .Y (n_27956));
OR2X1 g85127(.A (n_29039), .B (n_27965), .Y (n_27966));
AND2X1 g85131(.A (n_27963), .B (n_27964), .Y (n_27965));
NAND2X1 g31_dup85132(.A (n_9923), .B (n_9773), .Y (n_27963));
OR2X1 g85133(.A (n_14964), .B (n_9923), .Y (n_27964));
NAND2X1 g85136(.A (n_9923), .B (n_9773), .Y (n_27969));
INVX1 g85137(.A (n_27969), .Y (n_27970));
NAND2X1 g85148(.A (n_27988), .B (n_27990), .Y (n_27991));
INVX1 g85149(.A (n_27987), .Y (n_27988));
NAND2X2 g85150(.A (n_29153), .B (n_3493), .Y (n_27987));
INVX1 g85155(.A (n_27984), .Y (n_27985));
INVX1 g85156(.A (n_27983), .Y (n_27984));
INVX2 g85157(.A (sa02[6] ), .Y (n_27983));
INVX8 g85158(.A (n_1268), .Y (n_27990));
CLKBUFX3 g85159(.A (sa02[4] ), .Y (n_1268));
NOR2X1 g8(.A (n_28549), .B (n_434), .Y (n_28018));
NAND3X1 g85183(.A (n_28021), .B (n_28022), .C (n_28027), .Y(n_28028));
AND2X1 g85184(.A (n_28019), .B (n_28020), .Y (n_28021));
NAND2X1 g85185(.A (n_14769), .B (sa21[1] ), .Y (n_28019));
NAND2X1 g85186(.A (n_29102), .B (n_15874), .Y (n_28020));
OAI21X1 g85187(.A0 (n_26915), .A1 (n_14176), .B0 (n_21396), .Y(n_28022));
NOR2X1 g85188(.A (n_28024), .B (n_28026), .Y (n_28027));
NAND2X1 g85189(.A (n_17102), .B (n_28023), .Y (n_28024));
NAND2X1 g85190(.A (n_9959), .B (n_29149), .Y (n_28023));
NAND2X1 g85191(.A (n_8244), .B (n_28025), .Y (n_28026));
NAND2X1 g85192(.A (n_27441), .B (n_27914), .Y (n_28025));
NAND2X1 g85193(.A (n_28031), .B (n_28039), .Y (n_28040));
AND2X1 g85194(.A (n_28029), .B (n_28030), .Y (n_28031));
NAND2X1 g85195(.A (n_5944), .B (n_14624), .Y (n_28029));
NAND2X1 g48_dup(.A (n_6700), .B (n_17567), .Y (n_28030));
NOR2X1 g85196(.A (n_28036), .B (n_28038), .Y (n_28039));
NOR2X1 g85197(.A (n_28032), .B (n_28035), .Y (n_28036));
CLKBUFX1 g85198(.A (sa30[3] ), .Y (n_28032));
NAND2X2 g85199(.A (n_2885), .B (n_1340), .Y (n_28035));
NOR2X1 g85202(.A (n_28037), .B (n_6105), .Y (n_28038));
INVX4 g85203(.A (n_28032), .Y (n_28037));
INVX1 g85204(.A (n_28036), .Y (n_28041));
NAND2X1 g85205(.A (n_17567), .B (n_6700), .Y (n_28042));
INVX1 g85208(.A (n_28035), .Y (n_28045));
NAND4X1 g85209(.A (n_28047), .B (n_22219), .C (n_28051), .D(n_21618), .Y (n_28052));
AOI21X1 g85210(.A0 (n_21283), .A1 (n_21275), .B0 (n_28046), .Y(n_28047));
NAND2X1 g85211(.A (n_17966), .B (n_11858), .Y (n_28046));
NAND2X1 g85212(.A (sa22[0] ), .B (n_28050), .Y (n_28051));
NAND4X1 g85213(.A (n_18986), .B (n_28048), .C (n_28049), .D(n_18502), .Y (n_28050));
NAND2X1 g85214(.A (n_19219), .B (n_20574), .Y (n_28048));
NAND2X1 g85215(.A (n_19414), .B (n_17258), .Y (n_28049));
NOR2X1 g85216(.A (n_28055), .B (n_28060), .Y (n_28061));
AND2X1 g85217(.A (n_28053), .B (n_28054), .Y (n_28055));
NOR2X1 g85218(.A (n_28398), .B (n_3199), .Y (n_28053));
AND2X1 g85219(.A (n_11576), .B (n_27718), .Y (n_28054));
AOI21X1 g85220(.A0 (n_29392), .A1 (n_29393), .B0 (n_20018), .Y(n_28060));
NAND2X1 g85221(.A (n_16410), .B (n_7023), .Y (n_29393));
AOI21X1 g85222(.A0 (n_13454), .A1 (n_11576), .B0 (n_28057), .Y(n_29392));
NOR2X1 g85223(.A (n_11287), .B (n_27133), .Y (n_28057));
INVX1 g85225(.A (n_28053), .Y (n_28062));
NAND2X1 g85226(.A (n_13454), .B (n_11576), .Y (n_28063));
INVX1 g85227(.A (n_28057), .Y (n_28064));
NAND3X1 g85228(.A (n_28065), .B (n_28069), .C (n_28070), .Y(n_28071));
OAI21X1 g85229(.A0 (n_20943), .A1 (n_20770), .B0 (n_344), .Y(n_28065));
NOR2X1 g85230(.A (n_28066), .B (n_28068), .Y (n_28069));
NAND2X1 g85231(.A (n_20387), .B (n_20034), .Y (n_28066));
NAND2X1 g85232(.A (n_28067), .B (n_20389), .Y (n_28068));
AND2X1 g85233(.A (n_17808), .B (n_17004), .Y (n_28067));
NAND2X1 g85234(.A (n_27185), .B (sa30[0] ), .Y (n_28070));
NAND4X1 g85235(.A (n_28075), .B (n_28077), .C (n_28078), .D(n_28079), .Y (n_28080));
AOI21X1 g85236(.A0 (n_13972), .A1 (n_21242), .B0 (n_28074), .Y(n_28075));
NAND2X1 g85237(.A (n_28072), .B (n_28073), .Y (n_28074));
NAND2X1 g85238(.A (n_12601), .B (n_21242), .Y (n_28072));
AOI21X1 g85239(.A0 (n_14401), .A1 (n_11816), .B0 (sa03[0] ), .Y(n_28073));
INVX1 g85240(.A (n_28076), .Y (n_28077));
AOI21X1 g85241(.A0 (n_25638), .A1 (n_25637), .B0 (n_14627), .Y(n_28076));
NOR2X1 g85242(.A (n_15131), .B (n_18188), .Y (n_28078));
NAND2X1 g85243(.A (n_11816), .B (n_12591), .Y (n_28079));
MX2X1 g85272(.A (n_28110), .B (n_28109), .S0 (n_28111), .Y (n_28112));
INVX2 g85273(.A (n_28109), .Y (n_28110));
NAND2X2 g85274(.A (n_23033), .B (n_23329), .Y (n_28109));
MX2X1 g85275(.A (n_26218), .B (n_23503), .S0 (n_24265), .Y (n_28111));
XOR2X1 g85276(.A (n_28115), .B (n_28116), .Y (n_28117));
NAND2X1 g85277(.A (n_28113), .B (n_28114), .Y (n_28115));
AOI21X1 g85278(.A0 (n_21376), .A1 (sa03[0] ), .B0 (n_21977), .Y(n_28113));
NOR2X1 g85279(.A (n_19666), .B (n_21975), .Y (n_28114));
NAND2X1 g85280(.A (n_22126), .B (n_22357), .Y (n_28116));
NAND2X1 g85281(.A (n_28113), .B (n_28114), .Y (n_28118));
NAND2X1 g85282(.A (n_22357), .B (n_22126), .Y (n_28119));
AOI21X1 g85283(.A0 (n_28121), .A1 (n_28126), .B0 (n_28128), .Y(n_28129));
AOI21X1 g85284(.A0 (n_27610), .A1 (n_21151), .B0 (n_28120), .Y(n_28121));
AND2X1 g85285(.A (n_27216), .B (n_18068), .Y (n_28120));
NOR2X1 g85286(.A (n_28124), .B (n_28125), .Y (n_28126));
OR2X1 g85287(.A (n_28122), .B (n_28123), .Y (n_28124));
NOR2X1 g85288(.A (n_1063), .B (n_27603), .Y (n_28122));
NOR2X1 g85289(.A (n_27604), .B (n_15966), .Y (n_28123));
NAND2X1 g85290(.A (n_17657), .B (n_18209), .Y (n_28125));
INVX1 g85291(.A (n_28127), .Y (n_28128));
INVX1 g85292(.A (sa13[0] ), .Y (n_28127));
NOR2X1 g85293(.A (n_28130), .B (n_28137), .Y (n_28138));
NAND2X1 g85294(.A (n_4391), .B (n_28631), .Y (n_28130));
INVX1 g85295(.A (n_28136), .Y (n_28137));
INVX1 g85296(.A (n_28135), .Y (n_28136));
NAND2X2 g85297(.A (n_28132), .B (n_28134), .Y (n_28135));
INVX2 g85298(.A (n_28131), .Y (n_28132));
NAND2X1 g85299(.A (n_28365), .B (n_3121), .Y (n_28131));
INVX1 g85300(.A (n_28133), .Y (n_28134));
CLKBUFX1 g85301(.A (sa03[4] ), .Y (n_28133));
INVX1 g85303(.A (n_28133), .Y (n_8093));
INVX1 g85304(.A (sa03[4] ), .Y (n_28141));
NOR2X1 g85314(.A (n_28153), .B (n_4364), .Y (n_28156));
INVX2 g85315(.A (n_28152), .Y (n_28153));
NOR2X1 g85316(.A (sa12[7] ), .B (n_28151), .Y (n_28152));
INVX2 g85317(.A (sa12[6] ), .Y (n_28151));
CLKBUFX3 g85319(.A (sa12[4] ), .Y (n_28154));
INVX1 g85320(.A (sa12[7] ), .Y (n_28157));
INVX1 g85321(.A (n_28151), .Y (n_28158));
NAND3X1 g85322(.A (n_28160), .B (n_28161), .C (n_28164), .Y(n_28165));
INVX1 g85323(.A (n_28159), .Y (n_28160));
NOR2X1 g85324(.A (n_4514), .B (n_2466), .Y (n_28159));
NAND2X2 g85325(.A (n_4539), .B (n_6185), .Y (n_28161));
NAND2X1 g85326(.A (n_28163), .B (sa10[2] ), .Y (n_28164));
INVX1 g85327(.A (n_28162), .Y (n_28163));
NAND2X2 g85328(.A (n_1963), .B (n_288), .Y (n_28162));
INVX2 g85329(.A (n_28161), .Y (n_28166));
INVX1 g85330(.A (sa10[2] ), .Y (n_28167));
NOR2X1 g85331(.A (sa10[0] ), .B (n_28177), .Y (n_28178));
AOI21X1 g85332(.A0 (n_28168), .A1 (n_28170), .B0 (n_28176), .Y(n_28177));
NAND3X1 g85333(.A (n_26377), .B (n_26369), .C (n_26370), .Y(n_28168));
INVX1 g85334(.A (n_28169), .Y (n_28170));
INVX1 g85335(.A (sa10[1] ), .Y (n_28169));
NAND3X1 g85336(.A (n_28173), .B (n_28175), .C (n_17043), .Y(n_28176));
NAND2X1 g85337(.A (n_28171), .B (n_28172), .Y (n_28173));
NAND3X1 g85338(.A (n_14724), .B (n_15988), .C (n_16625), .Y(n_28171));
INVX1 g85339(.A (sa10[1] ), .Y (n_28172));
INVX1 g85340(.A (n_28174), .Y (n_28175));
NAND3X1 g85341(.A (n_12950), .B (n_10918), .C (n_8228), .Y (n_28174));
INVX1 g85342(.A (sa10[0] ), .Y (n_28179));
NOR2X1 g85344(.A (n_28185), .B (n_28189), .Y (n_28825));
NAND2X1 g85345(.A (n_21901), .B (n_28184), .Y (n_28185));
AND2X1 g85346(.A (n_28182), .B (n_28183), .Y (n_28184));
NOR2X1 g85347(.A (n_28181), .B (n_27162), .Y (n_28182));
OAI21X1 g85348(.A0 (n_12145), .A1 (n_11261), .B0 (n_28180), .Y(n_28181));
OR2X1 g85349(.A (n_3818), .B (n_10268), .Y (n_28180));
NAND2X1 g85350(.A (n_14540), .B (n_4529), .Y (n_28183));
NAND2X1 g85351(.A (n_28188), .B (n_22189), .Y (n_28189));
AND2X1 g85352(.A (n_28186), .B (n_28187), .Y (n_28188));
OAI21X1 g85353(.A0 (n_20215), .A1 (n_11994), .B0 (n_804), .Y(n_28186));
OAI21X1 g85354(.A0 (n_21265), .A1 (n_14537), .B0 (n_21055), .Y(n_28187));
NAND3X1 g85355(.A (n_28195), .B (n_28196), .C (n_28199), .Y(n_28200));
NAND2X1 g85356(.A (n_28193), .B (n_28194), .Y (n_28195));
NAND3X1 g85357(.A (n_28192), .B (n_20278), .C (n_20195), .Y(n_28193));
AND2X1 g85358(.A (n_18829), .B (n_18294), .Y (n_28192));
INVX1 g85359(.A (sa03[0] ), .Y (n_28194));
OAI21X1 g85360(.A0 (n_21436), .A1 (n_18454), .B0 (n_2909), .Y(n_28196));
NAND2X1 g85361(.A (n_28197), .B (n_19995), .Y (n_28199));
NAND2X1 g85362(.A (n_18755), .B (n_16614), .Y (n_28197));
NAND4X1 g85364(.A (n_29374), .B (n_29375), .C (n_28209), .D(n_28210), .Y (n_28211));
NAND2X1 g85365(.A (n_26406), .B (n_26405), .Y (n_29375));
NAND2X1 g85366(.A (n_28205), .B (n_28207), .Y (n_29374));
NAND2X1 g85367(.A (n_28204), .B (n_21331), .Y (n_28205));
NOR2X1 g85368(.A (n_28202), .B (n_28203), .Y (n_28204));
NAND3X1 g85369(.A (n_17610), .B (n_18341), .C (n_11849), .Y(n_28202));
INVX1 g85370(.A (n_20343), .Y (n_28203));
INVX1 g85371(.A (n_28206), .Y (n_28207));
INVX1 g85372(.A (sa01[0] ), .Y (n_28206));
OAI21X1 g85373(.A0 (n_21258), .A1 (n_20786), .B0 (n_21174), .Y(n_28209));
NOR2X1 g85374(.A (n_26410), .B (n_26411), .Y (n_28210));
NAND3X1 g85375(.A (n_28212), .B (n_28214), .C (n_28225), .Y(n_28226));
OAI21X1 g85376(.A0 (n_20842), .A1 (n_20374), .B0 (n_21938), .Y(n_28212));
INVX1 g85377(.A (n_28213), .Y (n_28214));
AOI21X1 g85378(.A0 (n_20823), .A1 (n_20184), .B0 (sa31[0] ), .Y(n_28213));
AOI21X1 g85379(.A0 (n_20835), .A1 (n_21581), .B0 (n_28224), .Y(n_28225));
NAND4X1 g85380(.A (n_28897), .B (n_28898), .C (n_28219), .D(n_28223), .Y (n_28224));
INVX1 g85381(.A (n_27089), .Y (n_28898));
INVX1 g85382(.A (n_27090), .Y (n_28897));
AOI21X1 g85383(.A0 (n_11391), .A1 (n_27100), .B0 (n_28218), .Y(n_28219));
INVX1 g85384(.A (n_28217), .Y (n_28218));
NAND2X1 g85385(.A (n_12836), .B (n_8362), .Y (n_28217));
NOR2X1 g85386(.A (n_28220), .B (n_28222), .Y (n_28223));
NOR2X1 g85387(.A (n_3384), .B (n_7120), .Y (n_28220));
INVX1 g85388(.A (n_28221), .Y (n_28222));
NAND2X1 g85389(.A (n_12155), .B (n_12634), .Y (n_28221));
NAND3X1 g85402(.A (n_27618), .B (n_27619), .C (n_27620), .Y(n_28287));
NAND3X1 g84795_dup(.A (n_27618), .B (n_27619), .C (n_27620), .Y(n_28288));
NAND4X1 g85421(.A (n_25774), .B (n_21479), .C (n_25775), .D(n_25506), .Y (n_28324));
NAND4X1 g59219_dup(.A (n_25774), .B (n_21479), .C (n_25775), .D(n_25506), .Y (n_28325));
NOR2X1 g85422(.A (n_29286), .B (n_14577), .Y (n_28326));
NOR2X1 g66870_dup(.A (n_29297), .B (n_14577), .Y (n_28327));
NAND2X1 g85423(.A (n_273), .B (n_767), .Y (n_28328));
NAND2X1 g77160_dup(.A (n_273), .B (n_767), .Y (n_28329));
CLKBUFX2 g85425(.A (n_28332), .Y (n_28331));
INVX2 g85426(.A (n_24104), .Y (n_28332));
INVX1 g85427(.A (n_23994), .Y (n_28333));
INVX1 g85429(.A (n_23994), .Y (n_28336));
CLKBUFX3 g85432(.A (n_28341), .Y (n_28340));
INVX1 g85435(.A (n_28345), .Y (n_28344));
INVX1 g85436(.A (n_28345), .Y (n_28346));
INVX2 g85438(.A (n_28350), .Y (n_28349));
INVX4 g85439(.A (n_28345), .Y (n_28350));
INVX4 g85440(.A (n_26287), .Y (n_28345));
INVX4 g85441(.A (n_28357), .Y (n_28351));
CLKBUFX1 g85444(.A (n_28357), .Y (n_28358));
INVX1 g85447(.A (n_28364), .Y (n_28362));
CLKBUFX1 g85448(.A (n_28365), .Y (n_28364));
INVX2 g85449(.A (n_28351), .Y (n_28365));
INVX4 g85451(.A (sa03[5] ), .Y (n_28357));
CLKBUFX1 g85455(.A (n_28375), .Y (n_28373));
INVX2 g85460(.A (n_28380), .Y (n_28381));
INVX1 g85461(.A (n_28375), .Y (n_28380));
CLKBUFX3 g85472(.A (n_28408), .Y (n_28398));
CLKBUFX1 g85476(.A (n_28402), .Y (n_28404));
INVX4 g85478(.A (n_28407), .Y (n_28402));
INVX4 g85479(.A (n_28407), .Y (n_28408));
INVX4 g85483(.A (n_28407), .Y (n_28410));
INVX4 g85484(.A (n_28375), .Y (n_28407));
INVX2 g85488(.A (n_28418), .Y (n_28419));
CLKBUFX3 g85489(.A (n_28375), .Y (n_28418));
INVX4 g85491(.A (n_28447), .Y (n_28423));
INVX2 g85496(.A (n_28447), .Y (n_28427));
INVX4 g85499(.A (n_28441), .Y (n_28433));
INVX2 g85506(.A (n_28445), .Y (n_28441));
CLKBUFX3 g85507(.A (n_28445), .Y (n_28444));
INVX2 g85508(.A (n_28447), .Y (n_28445));
INVX4 g85509(.A (n_28375), .Y (n_28447));
INVX8 g85510(.A (sa12[3] ), .Y (n_28375));
INVX1 g85513(.A (n_28459), .Y (n_28452));
CLKBUFX3 g85518(.A (n_28464), .Y (n_28459));
INVX4 g85520(.A (n_28464), .Y (n_28463));
INVX4 g85521(.A (sa01[5] ), .Y (n_28464));
INVX2 g85522(.A (n_28469), .Y (n_28466));
INVX1 g85525(.A (n_28472), .Y (n_28470));
CLKBUFX1 g85528(.A (n_28476), .Y (n_28472));
INVX2 g85531(.A (n_28469), .Y (n_28476));
INVX4 g85532(.A (n_28469), .Y (n_28478));
INVX4 g85533(.A (n_28482), .Y (n_28469));
INVX2 g85534(.A (n_28480), .Y (n_28481));
CLKBUFX3 g85535(.A (n_28482), .Y (n_28480));
INVX4 g85536(.A (sa31[5] ), .Y (n_28482));
CLKBUFX1 g85537(.A (n_28484), .Y (n_28483));
INVX1 g85538(.A (n_28487), .Y (n_28485));
INVX1 g85540(.A (n_28488), .Y (n_28487));
NAND4X1 g85552(.A (n_22325), .B (n_22044), .C (n_21625), .D(n_20127), .Y (n_23296));
NAND4X1 g59496_dup(.A (n_22325), .B (n_22044), .C (n_21625), .D(n_20127), .Y (n_28511));
INVX1 g85579(.A (n_28547), .Y (n_28540));
INVX1 g85581(.A (n_28547), .Y (n_28542));
CLKBUFX2 g85586(.A (n_28549), .Y (n_28547));
INVX1 g85587(.A (n_28549), .Y (n_28548));
INVX2 g85589(.A (sa01[6] ), .Y (n_28549));
NAND2X1 g85590(.A (n_27950), .B (n_22928), .Y (n_28563));
NAND2X1 g56859_dup(.A (n_27950), .B (n_22928), .Y (n_28564));
INVX2 g85591(.A (n_28567), .Y (n_28566));
CLKBUFX3 g85592(.A (n_28568), .Y (n_28567));
INVX1 g85597(.A (n_28575), .Y (n_28574));
CLKBUFX1 g85598(.A (n_28576), .Y (n_28575));
INVX1 g85599(.A (n_28577), .Y (n_28576));
INVX2 g85600(.A (n_28568), .Y (n_28577));
INVX4 g85601(.A (sa31[7] ), .Y (n_28568));
INVX1 g85602(.A (n_28580), .Y (n_28578));
INVX1 g85604(.A (n_8707), .Y (n_28580));
INVX2 g85606(.A (n_28610), .Y (n_28609));
INVX1 g85607(.A (n_5054), .Y (n_28610));
INVX1 g85608(.A (n_28616), .Y (n_28611));
INVX2 g85611(.A (n_28615), .Y (n_28614));
CLKBUFX1 g85612(.A (n_28616), .Y (n_28615));
INVX1 g85614(.A (n_28619), .Y (n_28618));
CLKBUFX1 g85615(.A (n_28620), .Y (n_28619));
INVX1 g85616(.A (n_10215), .Y (n_28620));
INVX1 g85625(.A (n_28631), .Y (n_28632));
INVX2 g85634(.A (n_28631), .Y (n_28645));
INVX8 g85654(.A (n_28631), .Y (n_28642));
INVX8 g85655(.A (n_28680), .Y (n_28631));
INVX2 g85672(.A (n_28631), .Y (n_28686));
INVX1 g85673(.A (n_28692), .Y (n_28689));
INVX8 g85701(.A (n_28631), .Y (n_28692));
INVX4 g85703(.A (sa03[2] ), .Y (n_28680));
INVX1 g85705(.A (n_28724), .Y (n_28725));
INVX2 g85706(.A (n_28727), .Y (n_28724));
INVX1 g85707(.A (n_3332), .Y (n_28727));
INVX1 g85708(.A (n_28733), .Y (n_28728));
CLKBUFX1 g85713(.A (n_28733), .Y (n_28734));
CLKBUFX3 g85715(.A (n_28771), .Y (n_28733));
CLKBUFX2 g85719(.A (n_28771), .Y (n_28742));
CLKBUFX1 g85724(.A (n_28744), .Y (n_28749));
INVX2 g85725(.A (sa11[4] ), .Y (n_28744));
INVX4 g85732(.A (n_28771), .Y (n_28754));
INVX8 g85739(.A (n_28754), .Y (n_28757));
INVX4 g85742(.A (sa11[4] ), .Y (n_28771));
CLKBUFX1 g85744(.A (n_28776), .Y (n_28775));
INVX2 g85745(.A (n_27522), .Y (n_28776));
INVX4 g85747(.A (n_28786), .Y (n_28779));
INVX1 g85748(.A (n_28781), .Y (n_28780));
CLKBUFX1 g85751(.A (n_28785), .Y (n_28781));
CLKBUFX1 g85752(.A (n_28786), .Y (n_28785));
CLKBUFX1 g85753(.A (n_28786), .Y (n_28787));
INVX4 g85755(.A (sa12[5] ), .Y (n_28786));
CLKBUFX1 g85756(.A (n_28793), .Y (n_28792));
INVX2 g85757(.A (sa12[5] ), .Y (n_28793));
CLKBUFX2 g85758(.A (n_28802), .Y (n_28796));
INVX2 g85759(.A (n_28797), .Y (n_28798));
INVX1 g85760(.A (n_28800), .Y (n_28799));
CLKBUFX1 g85761(.A (n_28797), .Y (n_28800));
INVX2 g85762(.A (n_28802), .Y (n_28797));
INVX1 g85763(.A (n_28804), .Y (n_28803));
INVX1 g85765(.A (n_28809), .Y (n_28807));
INVX1 g85767(.A (n_28812), .Y (n_28810));
INVX2 g85771(.A (n_28816), .Y (n_28815));
INVX1 g85775(.A (n_28822), .Y (n_28821));
INVX2 g85776(.A (n_28820), .Y (n_28822));
CLKBUFX3 g85778(.A (n_28825), .Y (n_28820));
INVX1 g85779(.A (n_28826), .Y (n_28827));
INVX2 g85780(.A (n_28825), .Y (n_28826));
INVX1 g85781(.A (n_28832), .Y (n_28829));
INVX1 g85785(.A (n_28836), .Y (n_28834));
OR2X1 g85788(.A (n_27202), .B (n_6706), .Y (n_28857));
OR2X1 g84589_dup(.A (n_27202), .B (n_6706), .Y (n_28858));
NAND2X1 g85789(.A (n_1686), .B (n_28466), .Y (n_28859));
NAND2X1 g75346_dup(.A (n_1686), .B (n_28466), .Y (n_28860));
INVX2 g85791(.A (n_28865), .Y (n_28862));
CLKBUFX1 g85794(.A (n_28866), .Y (n_28865));
INVX1 g85797(.A (n_28870), .Y (n_28869));
CLKBUFX1 g85798(.A (n_28871), .Y (n_28870));
INVX2 g85799(.A (n_28872), .Y (n_28871));
INVX2 g85800(.A (n_2067), .Y (n_28872));
INVX1 g85802(.A (n_28877), .Y (n_28875));
NAND2X1 g85805(.A (n_22730), .B (n_19818), .Y (n_28899));
NAND2X1 g58780_dup(.A (n_22730), .B (n_19818), .Y (n_28900));
NAND2X1 g85806(.A (n_7798), .B (n_28418), .Y (n_28901));
NAND2X1 g67363_dup(.A (n_7798), .B (n_28418), .Y (n_28902));
OR4X1 g85807(.A (n_19623), .B (n_21779), .C (n_21395), .D (n_22381),.Y (n_28903));
OR4X1 g59097_dup(.A (n_19623), .B (n_21779), .C (n_21395), .D(n_22381), .Y (n_28904));
CLKBUFX1 g85808(.A (n_28907), .Y (n_28905));
INVX1 g85868(.A (n_28986), .Y (n_28988));
INVX1 g85871(.A (n_28996), .Y (n_28993));
INVX1 g85874(.A (n_3381), .Y (n_28996));
INVX1 g85876(.A (n_29000), .Y (n_28998));
INVX1 g85879(.A (n_29003), .Y (n_29002));
INVX2 g85880(.A (n_29005), .Y (n_29003));
INVX4 g85882(.A (n_29007), .Y (n_29005));
CLKBUFX3 g85883(.A (n_27305), .Y (n_29007));
INVX1 g85890(.A (n_29018), .Y (n_29014));
INVX8 g85918(.A (n_29039), .Y (n_29048));
INVX4 g85924(.A (n_29062), .Y (n_29039));
INVX8 g85928(.A (n_29018), .Y (n_29062));
INVX8 g85929(.A (n_29065), .Y (n_29018));
INVX1 g85937(.A (n_29074), .Y (n_29070));
CLKBUFX3 g85943(.A (n_29065), .Y (n_29074));
INVX4 g85944(.A (sa21[2] ), .Y (n_29065));
INVX1 g85948(.A (n_29106), .Y (n_29085));
INVX1 g85966(.A (n_29102), .Y (n_29106));
INVX4 g85973(.A (sa21[2] ), .Y (n_29102));
INVX2 g85974(.A (n_26851), .Y (n_29114));
INVX1 g85975(.A (n_29122), .Y (n_29116));
INVX1 g85978(.A (n_29120), .Y (n_29119));
CLKBUFX1 g85979(.A (n_29121), .Y (n_29120));
CLKBUFX3 g85980(.A (n_29122), .Y (n_29121));
NAND2X1 g85981(.A (n_26394), .B (n_1015), .Y (n_29131));
NAND2X1 g76703_dup(.A (n_26394), .B (n_1015), .Y (n_29409));
NAND4X1 g85982(.A (n_25476), .B (n_21034), .C (n_25477), .D(n_25453), .Y (n_29133));
NAND4X1 g59428_dup(.A (n_25476), .B (n_21034), .C (n_25477), .D(n_25453), .Y (n_29134));
NAND2X1 g85983(.A (n_26540), .B (n_26543), .Y (n_29135));
NAND2X1 g83734_dup(.A (n_26540), .B (n_26543), .Y (n_29136));
INVX1 g85984(.A (n_29139), .Y (n_29137));
CLKBUFX1 g85986(.A (n_29140), .Y (n_29139));
INVX1 g85988(.A (n_29140), .Y (n_29142));
CLKBUFX1 g85990(.A (n_29150), .Y (n_29149));
INVX1 g85991(.A (n_2151), .Y (n_29150));
INVX2 g85993(.A (n_29155), .Y (n_29153));
INVX4 g85995(.A (n_29158), .Y (n_29155));
INVX4 g85998(.A (sa02[5] ), .Y (n_29158));
INVX1 g86001(.A (n_29166), .Y (n_29163));
CLKBUFX2 g86003(.A (n_29167), .Y (n_29166));
INVX2 g86005(.A (sa02[5] ), .Y (n_29167));
INVX1 g86006(.A (n_29173), .Y (n_29171));
INVX1 g86009(.A (n_29176), .Y (n_29173));
NOR2X1 g86010(.A (n_28871), .B (n_6021), .Y (n_29181));
NOR2X1 g75263_dup(.A (n_28871), .B (n_6021), .Y (n_29182));
NOR2X1 g86012(.A (n_7505), .B (n_3318), .Y (n_29185));
NOR2X1 g66183_dup(.A (n_7505), .B (n_3318), .Y (n_29186));
XOR2X1 g86013(.A (u0_rcon_1059), .B (n_23596), .Y (n_29187));
XOR2X1 g58863_dup(.A (u0_rcon_1059), .B (n_23596), .Y (n_29188));
INVX1 g86014(.A (n_5072), .Y (n_29189));
INVX1 g86015(.A (n_29191), .Y (n_29190));
CLKBUFX1 g86016(.A (n_29193), .Y (n_29191));
INVX1 g86017(.A (n_29193), .Y (n_29192));
CLKBUFX1 g86018(.A (n_5072), .Y (n_29193));
NAND2X2 g86019(.A (n_9101), .B (n_6005), .Y (n_29198));
NAND2X1 g69191_dup(.A (n_9101), .B (n_6005), .Y (n_29199));
NOR2X1 g86020(.A (n_27954), .B (n_27957), .Y (n_29200));
NOR2X1 g85119_dup(.A (n_27954), .B (n_27957), .Y (n_29201));
INVX2 g86021(.A (n_29203), .Y (n_29202));
INVX2 g86022(.A (n_29204), .Y (n_29203));
INVX2 g86023(.A (n_29205), .Y (n_29204));
INVX2 g86024(.A (n_26000), .Y (n_29205));
INVX1 g86032(.A (n_29214), .Y (n_29215));
CLKBUFX1 g86033(.A (n_29217), .Y (n_29216));
CLKBUFX1 g86036(.A (n_29228), .Y (n_29221));
INVX2 g86039(.A (n_29235), .Y (n_29225));
INVX4 g86045(.A (n_29235), .Y (n_29228));
CLKBUFX1 g86050(.A (n_28933), .Y (n_29235));
INVX4 g86055(.A (n_29266), .Y (n_29244));
INVX4 g86064(.A (n_29262), .Y (n_29256));
CLKBUFX1 g86072(.A (n_29266), .Y (n_29262));
INVX2 g86073(.A (n_29298), .Y (n_29266));
CLKBUFX1 g86078(.A (n_29269), .Y (n_29275));
BUFX3 g86079(.A (n_29298), .Y (n_29269));
INVX1 g86081(.A (n_29292), .Y (n_29279));
INVX2 g86087(.A (n_29292), .Y (n_29286));
INVX4 g86093(.A (n_29297), .Y (n_29292));
CLKBUFX3 g86098(.A (n_29298), .Y (n_29297));
INVX2 g86099(.A (n_28933), .Y (n_29298));
NAND4X1 g86100(.A (n_26197), .B (n_26199), .C (n_26200), .D(n_26204), .Y (n_29326));
NAND4X1 g83398_dup(.A (n_26197), .B (n_26199), .C (n_26200), .D(n_26204), .Y (n_29327));
INVX1 g86102(.A (n_29330), .Y (n_29329));
INVX1 g86103(.A (n_29333), .Y (n_29331));
CLKBUFX2 g86106(.A (n_29330), .Y (n_29333));
INVX1 g86107(.A (n_4467), .Y (n_29330));
INVX1 g86108(.A (n_29336), .Y (n_29337));
INVX2 g86114(.A (n_6117), .Y (n_29343));
INVX2 g86116(.A (n_29351), .Y (n_29347));
INVX1 g86117(.A (n_29351), .Y (n_29349));
INVX1 g86118(.A (n_29351), .Y (n_29350));
INVX2 g86119(.A (n_29353), .Y (n_29351));
INVX1 g86121(.A (n_29357), .Y (n_29355));
CLKBUFX1 g86123(.A (n_29360), .Y (n_29357));
INVX1 g86124(.A (n_29360), .Y (n_29358));
INVX2 g86129(.A (n_4588), .Y (n_29363));
endmodule
