module wb_dma_top ( clk_i, rst_i, wb0s_data_i, wb0s_data_o, wb0_addr_i,wb0_sel_i, wb0_we_i, wb0_cyc_i, wb0_stb_i, wb0_ack_o, wb0_err_o,wb0_rty_o, wb0m_data_i, wb0m_data_o, wb0_addr_o, wb0_sel_o, wb0_we_o,wb0_cyc_o, wb0_stb_o, wb0_ack_i, wb0_err_i, wb0_rty_i, wb1s_data_i,wb1s_data_o, wb1_addr_i, wb1_sel_i, wb1_we_i, wb1_cyc_i, wb1_stb_i,wb1_ack_o, wb1_err_o, wb1_rty_o, wb1m_data_i, wb1m_data_o, wb1_addr_o,wb1_sel_o, wb1_we_o, wb1_cyc_o, wb1_stb_o, wb1_ack_i, wb1_err_i,wb1_rty_i, dma_req_i, dma_ack_o, dma_nd_i, dma_rest_i, inta_o, intb_o, _u2_adr1_cnt_next1, _u2_adr0_cnt_next1);
input [31:0] wb0s_data_i;
output [31:0] wb0s_data_o;
input [31:0] wb0_addr_i;
input [3:0] wb0_sel_i;
input [31:0] wb0m_data_i;
output [31:0] wb0m_data_o;
output [31:0] wb0_addr_o;
output [3:0] wb0_sel_o;
input [31:0] wb1s_data_i;
output [31:0] wb1s_data_o;
input [31:0] wb1_addr_i;
input [3:0] wb1_sel_i;
input [31:0] wb1m_data_i;
output [31:0] wb1m_data_o;
output [31:0] wb1_addr_o;
output [3:0] wb1_sel_o;
input [0:0] dma_req_i;
output [0:0] dma_ack_o;
input [0:0] dma_nd_i;
input [0:0] dma_rest_i;
input clk_i, rst_i, wb0_we_i, wb0_cyc_i, wb0_stb_i, wb0_ack_i, wb0_err_i,wb0_rty_i, wb1_we_i, wb1_cyc_i, wb1_stb_i, wb1_ack_i, wb1_err_i,wb1_rty_i;
output wb0_ack_o, wb0_err_o, wb0_rty_o, wb0_we_o, wb0_cyc_o, wb0_stb_o,wb1_ack_o, wb1_err_o, wb1_rty_o, wb1_we_o, wb1_cyc_o, wb1_stb_o,inta_o, intb_o;
wire   pt1_sel_i, pt0_sel_i, slv0_re, slv0_we, pause_req, paused, dma_abort,dma_busy, dma_err, dma_done, dma_done_all, de_csr_we, de_txsz_we,de_adr0_we, de_adr1_we, de_fetch_descr, ptr_set, de_start, ndr,next_ch, de_ack, mast0_go, mast0_we, mast0_err, mast0_drdy,mast0_wait, mast1_go, mast1_we, mast1_err, mast1_drdy, mast1_wait, n5,SYNOPSYS_UNCONNECTED_7863, SYNOPSYS_UNCONNECTED_7864,SYNOPSYS_UNCONNECTED_7865, SYNOPSYS_UNCONNECTED_7866,SYNOPSYS_UNCONNECTED_7867, SYNOPSYS_UNCONNECTED_7868,SYNOPSYS_UNCONNECTED_7869, SYNOPSYS_UNCONNECTED_7870,SYNOPSYS_UNCONNECTED_7871, SYNOPSYS_UNCONNECTED_7872,SYNOPSYS_UNCONNECTED_7873, SYNOPSYS_UNCONNECTED_7874,SYNOPSYS_UNCONNECTED_7875, SYNOPSYS_UNCONNECTED_7876,SYNOPSYS_UNCONNECTED_7877, SYNOPSYS_UNCONNECTED_7878,SYNOPSYS_UNCONNECTED_7879, SYNOPSYS_UNCONNECTED_7880,SYNOPSYS_UNCONNECTED_7881, SYNOPSYS_UNCONNECTED_7882,SYNOPSYS_UNCONNECTED_7883, SYNOPSYS_UNCONNECTED_7884,SYNOPSYS_UNCONNECTED_7885, SYNOPSYS_UNCONNECTED_7886,SYNOPSYS_UNCONNECTED_7887, SYNOPSYS_UNCONNECTED_7888,SYNOPSYS_UNCONNECTED_7889, SYNOPSYS_UNCONNECTED_7890,SYNOPSYS_UNCONNECTED_7891, SYNOPSYS_UNCONNECTED_7892,SYNOPSYS_UNCONNECTED_7893, SYNOPSYS_UNCONNECTED_7894,SYNOPSYS_UNCONNECTED_7895, SYNOPSYS_UNCONNECTED_7896,SYNOPSYS_UNCONNECTED_7897, SYNOPSYS_UNCONNECTED_7898,SYNOPSYS_UNCONNECTED_7899, SYNOPSYS_UNCONNECTED_7900,SYNOPSYS_UNCONNECTED_7901, SYNOPSYS_UNCONNECTED_7902,SYNOPSYS_UNCONNECTED_7903, SYNOPSYS_UNCONNECTED_7904,SYNOPSYS_UNCONNECTED_7905, SYNOPSYS_UNCONNECTED_7906,SYNOPSYS_UNCONNECTED_7907, SYNOPSYS_UNCONNECTED_7908,SYNOPSYS_UNCONNECTED_7909, SYNOPSYS_UNCONNECTED_7910,SYNOPSYS_UNCONNECTED_7911, SYNOPSYS_UNCONNECTED_7912,SYNOPSYS_UNCONNECTED_7913, SYNOPSYS_UNCONNECTED_7914,SYNOPSYS_UNCONNECTED_7915, SYNOPSYS_UNCONNECTED_7916,SYNOPSYS_UNCONNECTED_7917, SYNOPSYS_UNCONNECTED_7918,SYNOPSYS_UNCONNECTED_7919, SYNOPSYS_UNCONNECTED_7920,SYNOPSYS_UNCONNECTED_7921, SYNOPSYS_UNCONNECTED_7922,SYNOPSYS_UNCONNECTED_7923, SYNOPSYS_UNCONNECTED_7924,SYNOPSYS_UNCONNECTED_7925, SYNOPSYS_UNCONNECTED_7926,SYNOPSYS_UNCONNECTED_7927, SYNOPSYS_UNCONNECTED_7928,SYNOPSYS_UNCONNECTED_7929, SYNOPSYS_UNCONNECTED_7930,SYNOPSYS_UNCONNECTED_7931, SYNOPSYS_UNCONNECTED_7932,SYNOPSYS_UNCONNECTED_7933, SYNOPSYS_UNCONNECTED_7934,SYNOPSYS_UNCONNECTED_7935, SYNOPSYS_UNCONNECTED_7936,SYNOPSYS_UNCONNECTED_7937, SYNOPSYS_UNCONNECTED_7938,SYNOPSYS_UNCONNECTED_7939, SYNOPSYS_UNCONNECTED_7940,SYNOPSYS_UNCONNECTED_7941, SYNOPSYS_UNCONNECTED_7942,SYNOPSYS_UNCONNECTED_7943, SYNOPSYS_UNCONNECTED_7944,SYNOPSYS_UNCONNECTED_7945, SYNOPSYS_UNCONNECTED_7946,SYNOPSYS_UNCONNECTED_7947, SYNOPSYS_UNCONNECTED_7948,SYNOPSYS_UNCONNECTED_7949, SYNOPSYS_UNCONNECTED_7950, _u0_n16309 ,_u0_n16308 , _u0_n16307 , _u0_n16306 , _u0_n16305 , _u0_n16304 ,_u0_n16303 , _u0_n16302 , _u0_n16301 , _u0_n16300 , _u0_n16299 ,_u0_n16298 , _u0_n16297 , _u0_n16296 , _u0_n16295 , _u0_n16294 ,_u0_n16293 , _u0_n16292 , _u0_n16291 , _u0_n16290 , _u0_n16289 ,_u0_n16288 , _u0_n16287 , _u0_n16286 , _u0_n16285 , _u0_n16284 ,_u0_n16283 , _u0_n16282 , _u0_n16281 , _u0_n16280 , _u0_n16279 ,_u0_n16278 , _u0_n16277 , _u0_n16276 , _u0_n16275 , _u0_n16274 ,_u0_n16273 , _u0_n16272 , _u0_n16271 , _u0_n16270 , _u0_n16269 ,_u0_n16268 , _u0_n16267 , _u0_n16266 , _u0_n16265 , _u0_n16264 ,_u0_n16263 , _u0_n16262 , _u0_n16261 , _u0_n16260 , _u0_n16259 ,_u0_n16258 , _u0_n16257 , _u0_n16256 , _u0_n16255 , _u0_n16254 ,_u0_n16253 , _u0_n16252 , _u0_n16251 , _u0_n16250 , _u0_n16249 ,_u0_n16248 , _u0_n16247 , _u0_n16246 , _u0_n16245 , _u0_n16244 ,_u0_n16243 , _u0_n16242 , _u0_n16241 , _u0_n16240 , _u0_n16239 ,_u0_n16238 , _u0_n16237 , _u0_n16236 , _u0_n16235 , _u0_n16234 ,_u0_n16233 , _u0_n16232 , _u0_n16231 , _u0_n16230 , _u0_n16229 ,_u0_n16228 , _u0_n16227 , _u0_n16226 , _u0_n16225 , _u0_n16224 ,_u0_n16223 , _u0_n16222 , _u0_n16221 , _u0_n16220 , _u0_n16219 ,_u0_n16218 , _u0_n16217 , _u0_n16216 , _u0_n16215 , _u0_n16214 ,_u0_n16213 , _u0_n16212 , _u0_n16211 , _u0_n16210 , _u0_n16209 ,_u0_n16208 , _u0_n16207 , _u0_n16206 , _u0_n16205 , _u0_n16204 ,_u0_n16203 , _u0_n16202 , _u0_n16201 , _u0_n16200 , _u0_n16199 ,_u0_n16198 , _u0_n16197 , _u0_n16196 , _u0_n16195 , _u0_n16194 ,_u0_n16193 , _u0_n16192 , _u0_n16191 , _u0_n16190 , _u0_n16189 ,_u0_n16188 , _u0_n16187 , _u0_n16186 , _u0_n16185 , _u0_n16184 ,_u0_n16183 , _u0_n16182 , _u0_n16181 , _u0_n16180 , _u0_n16179 ,_u0_n16178 , _u0_n16177 , _u0_n16176 , _u0_n16175 , _u0_n16174 ,_u0_n16173 , _u0_n16172 , _u0_n16171 , _u0_n16170 , _u0_n16169 ,_u0_n16168 , _u0_n16167 , _u0_n16166 , _u0_n16165 , _u0_n16164 ,_u0_n16163 , _u0_n16162 , _u0_n16161 , _u0_n16160 , _u0_n16159 ,_u0_n16158 , _u0_n16157 , _u0_n16156 , _u0_n16155 , _u0_n16154 ,_u0_n16153 , _u0_n16152 , _u0_n16151 , _u0_n16150 , _u0_n16149 ,_u0_n16148 , _u0_n16147 , _u0_n16146 , _u0_n16145 , _u0_n16144 ,_u0_n16143 , _u0_n16142 , _u0_n16141 , _u0_n16140 , _u0_n16139 ,_u0_n16138 , _u0_n16137 , _u0_n16136 , _u0_n16135 , _u0_n16134 ,_u0_n16133 , _u0_n16132 , _u0_n16131 , _u0_n16130 , _u0_n16129 ,_u0_n16128 , _u0_n16127 , _u0_n16126 , _u0_n16125 , _u0_n16124 ,_u0_n16123 , _u0_n16122 , _u0_n16121 , _u0_n16120 , _u0_n16119 ,_u0_n16118 , _u0_n16117 , _u0_n16116 , _u0_n16115 , _u0_n16114 ,_u0_n16113 , _u0_n16112 , _u0_n16111 , _u0_n16110 , _u0_n16109 ,_u0_n16108 , _u0_n16107 , _u0_n16106 , _u0_n16105 , _u0_n16104 ,_u0_n16103 , _u0_n16102 , _u0_n16101 , _u0_n16100 , _u0_n16099 ,_u0_n16098 , _u0_n16097 , _u0_n16096 , _u0_n16095 , _u0_n16094 ,_u0_n16093 , _u0_n16092 , _u0_n16091 , _u0_n16090 , _u0_n16089 ,_u0_n16088 , _u0_n16087 , _u0_n16086 , _u0_n16085 , _u0_n16084 ,_u0_n16083 , _u0_n16082 , _u0_n16081 , _u0_n16080 , _u0_n16079 ,_u0_n16078 , _u0_n16077 , _u0_n16076 , _u0_n16075 , _u0_n16074 ,_u0_n16073 , _u0_n16072 , _u0_n16071 , _u0_n16070 , _u0_n16069 ,_u0_n16068 , _u0_n16067 , _u0_n16066 , _u0_n16065 , _u0_n16064 ,_u0_n16063 , _u0_n16062 , _u0_n16061 , _u0_n16060 , _u0_n16059 ,_u0_n16058 , _u0_n16057 , _u0_n16056 , _u0_n16055 , _u0_n16054 ,_u0_n16053 , _u0_n16052 , _u0_n16051 , _u0_n16050 , _u0_n16049 ,_u0_n16048 , _u0_n16047 , _u0_n16046 , _u0_n16045 , _u0_n16044 ,_u0_n16043 , _u0_n16042 , _u0_n16041 , _u0_n16040 , _u0_n16039 ,_u0_n16038 , _u0_n16037 , _u0_n16036 , _u0_n16035 , _u0_n16034 ,_u0_n16033 , _u0_n16032 , _u0_n16031 , _u0_n16030 , _u0_n16029 ,_u0_n16028 , _u0_n16027 , _u0_n16026 , _u0_n16025 , _u0_n16024 ,_u0_n16023 , _u0_n16022 , _u0_n16021 , _u0_n16020 , _u0_n16019 ,_u0_n16018 , _u0_pointer0[31] , _u0_pointer0[30] , _u0_pointer0[29] ,_u0_pointer0[28] , _u0_pointer0[27] , _u0_pointer0[26] ,_u0_pointer0[25] , _u0_pointer0[24] , _u0_pointer0[23] ,_u0_pointer0[22] , _u0_pointer0[21] , _u0_pointer0[20] ,_u0_pointer0[19] , _u0_pointer0[18] , _u0_pointer0[17] ,_u0_pointer0[16] , _u0_pointer0[15] , _u0_pointer0[14] ,_u0_pointer0[13] , _u0_pointer0[12] , _u0_pointer0[11] ,_u0_pointer0[10] , _u0_pointer0[9] , _u0_pointer0[8] ,_u0_pointer0[7] , _u0_pointer0[6] , _u0_pointer0[5] ,_u0_pointer0[4] , _u0_pointer0[3] , _u0_pointer0[2] ,_u0_pointer0[1] , _u0_pointer0[0] , _u0_pointer0_s[31] ,_u0_pointer0_s[30] , _u0_pointer0_s[29] , _u0_pointer0_s[28] ,_u0_pointer0_s[27] , _u0_pointer0_s[26] , _u0_pointer0_s[25] ,_u0_pointer0_s[24] , _u0_pointer0_s[23] , _u0_pointer0_s[22] ,_u0_pointer0_s[21] , _u0_pointer0_s[20] , _u0_pointer0_s[19] ,_u0_pointer0_s[18] , _u0_pointer0_s[17] , _u0_pointer0_s[16] ,_u0_pointer0_s[15] , _u0_pointer0_s[14] , _u0_pointer0_s[13] ,_u0_pointer0_s[12] , _u0_pointer0_s[11] , _u0_pointer0_s[10] ,_u0_pointer0_s[9] , _u0_pointer0_s[8] , _u0_pointer0_s[7] ,_u0_pointer0_s[6] , _u0_pointer0_s[5] , _u0_pointer0_s[4] ,_u0_pointer0_s[3] , _u0_pointer0_s[2] , _u0_pointer0_s[1] ,_u0_pointer0_s[0] , _u0_ch0_csr[31] , _u0_ch0_csr[30] ,_u0_ch0_csr[29] , _u0_ch0_csr[28] , _u0_ch0_csr[27] ,_u0_ch0_csr[26] , _u0_ch0_csr[25] , _u0_ch0_csr[24] ,_u0_ch0_csr[23] , _u0_ch0_csr[9] , _u0_ch0_txsz[31] ,_u0_ch0_txsz[30] , _u0_ch0_txsz[29] , _u0_ch0_txsz[28] ,_u0_ch0_txsz[27] , _u0_ch0_txsz[14] , _u0_ch0_txsz[13] ,_u0_ch0_txsz[12] , _u0_ch0_adr0[1] , _u0_ch0_adr0[0] ,_u0_ch0_adr1[1] , _u0_ch0_adr1[0] , _u0_ch0_am0[31] ,_u0_ch0_am0[30] , _u0_ch0_am0[29] , _u0_ch0_am0[28] ,_u0_ch0_am0[27] , _u0_ch0_am0[26] , _u0_ch0_am0[25] ,_u0_ch0_am0[24] , _u0_ch0_am0[23] , _u0_ch0_am0[22] ,_u0_ch0_am0[21] , _u0_ch0_am0[20] , _u0_ch0_am0[19] ,_u0_ch0_am0[18] , _u0_ch0_am0[17] , _u0_ch0_am0[16] ,_u0_ch0_am0[15] , _u0_ch0_am0[14] , _u0_ch0_am0[13] ,_u0_ch0_am0[12] , _u0_ch0_am0[11] , _u0_ch0_am0[10] , _u0_ch0_am0[9] ,_u0_ch0_am0[8] , _u0_ch0_am0[7] , _u0_ch0_am0[6] , _u0_ch0_am0[5] ,_u0_ch0_am0[4] , _u0_ch0_am0[3] , _u0_ch0_am0[2] , _u0_ch0_am0[1] ,_u0_ch0_am0[0] , _u0_ch0_am1[31] , _u0_ch0_am1[30] , _u0_ch0_am1[29] ,_u0_ch0_am1[28] , _u0_ch0_am1[27] , _u0_ch0_am1[26] ,_u0_ch0_am1[25] , _u0_ch0_am1[24] , _u0_ch0_am1[23] ,_u0_ch0_am1[22] , _u0_ch0_am1[21] , _u0_ch0_am1[20] ,_u0_ch0_am1[19] , _u0_ch0_am1[18] , _u0_ch0_am1[17] ,_u0_ch0_am1[16] , _u0_ch0_am1[15] , _u0_ch0_am1[14] ,_u0_ch0_am1[13] , _u0_ch0_am1[12] , _u0_ch0_am1[11] ,_u0_ch0_am1[10] , _u0_ch0_am1[9] , _u0_ch0_am1[8] , _u0_ch0_am1[7] ,_u0_ch0_am1[6] , _u0_ch0_am1[5] , _u0_ch0_am1[4] , _u0_ch0_am1[3] ,_u0_ch0_am1[2] , _u0_ch0_am1[1] , _u0_ch0_am1[0] , _u0_pointer1[31] ,_u0_pointer1[30] , _u0_pointer1[29] , _u0_pointer1[28] ,_u0_pointer1[27] , _u0_pointer1[26] , _u0_pointer1[25] ,_u0_pointer1[24] , _u0_pointer1[23] , _u0_pointer1[22] ,_u0_pointer1[21] , _u0_pointer1[20] , _u0_pointer1[19] ,_u0_pointer1[18] , _u0_pointer1[17] , _u0_pointer1[16] ,_u0_pointer1[15] , _u0_pointer1[14] , _u0_pointer1[13] ,_u0_pointer1[12] , _u0_pointer1[11] , _u0_pointer1[10] ,_u0_pointer1[9] , _u0_pointer1[8] , _u0_pointer1[7] ,_u0_pointer1[6] , _u0_pointer1[5] , _u0_pointer1[4] ,_u0_pointer1[3] , _u0_pointer1[2] , _u0_pointer1[1] ,_u0_pointer1[0] , _u0_pointer1_s[31] , _u0_pointer1_s[30] ,_u0_pointer1_s[29] , _u0_pointer1_s[28] , _u0_pointer1_s[27] ,_u0_pointer1_s[26] , _u0_pointer1_s[25] , _u0_pointer1_s[24] ,_u0_pointer1_s[23] , _u0_pointer1_s[22] , _u0_pointer1_s[21] ,_u0_pointer1_s[20] , _u0_pointer1_s[19] , _u0_pointer1_s[18] ,_u0_pointer1_s[17] , _u0_pointer1_s[16] , _u0_pointer1_s[15] ,_u0_pointer1_s[14] , _u0_pointer1_s[13] , _u0_pointer1_s[12] ,_u0_pointer1_s[11] , _u0_pointer1_s[10] , _u0_pointer1_s[9] ,_u0_pointer1_s[8] , _u0_pointer1_s[7] , _u0_pointer1_s[6] ,_u0_pointer1_s[5] , _u0_pointer1_s[4] , _u0_pointer1_s[3] ,_u0_pointer1_s[2] , _u0_pointer1_s[1] , _u0_pointer1_s[0] ,_u0_ch1_csr[31] , _u0_ch1_csr[30] , _u0_ch1_csr[29] ,_u0_ch1_csr[28] , _u0_ch1_csr[27] , _u0_ch1_csr[26] ,_u0_ch1_csr[25] , _u0_ch1_csr[24] , _u0_ch1_csr[23] ,_u0_ch1_csr[22] , _u0_ch1_csr[21] , _u0_ch1_csr[20] ,_u0_ch1_csr[19] , _u0_ch1_csr[18] , _u0_ch1_csr[17] ,_u0_ch1_csr[16] , _u0_ch1_csr[15] , _u0_ch1_csr[14] ,_u0_ch1_csr[13] , _u0_ch1_csr[12] , _u0_ch1_csr[11] ,_u0_ch1_csr[10] , _u0_ch1_csr[9] , _u0_ch1_csr[8] , _u0_ch1_csr[7] ,_u0_ch1_csr[6] , _u0_ch1_csr[5] , _u0_ch1_csr[4] , _u0_ch1_csr[3] ,_u0_ch1_csr[2] , _u0_ch1_csr[1] , _u0_ch1_csr[0] , _u0_ch1_txsz[31] ,_u0_ch1_txsz[30] , _u0_ch1_txsz[29] , _u0_ch1_txsz[28] ,_u0_ch1_txsz[27] , _u0_ch1_txsz[26] , _u0_ch1_txsz[25] ,_u0_ch1_txsz[24] , _u0_ch1_txsz[23] , _u0_ch1_txsz[22] ,_u0_ch1_txsz[21] , _u0_ch1_txsz[20] , _u0_ch1_txsz[19] ,_u0_ch1_txsz[18] , _u0_ch1_txsz[17] , _u0_ch1_txsz[16] ,_u0_ch1_txsz[15] , _u0_ch1_txsz[14] , _u0_ch1_txsz[13] ,_u0_ch1_txsz[12] , _u0_ch1_txsz[11] , _u0_ch1_txsz[10] ,_u0_ch1_txsz[9] , _u0_ch1_txsz[8] , _u0_ch1_txsz[7] ,_u0_ch1_txsz[6] , _u0_ch1_txsz[5] , _u0_ch1_txsz[4] ,_u0_ch1_txsz[3] , _u0_ch1_txsz[2] , _u0_ch1_txsz[1] ,_u0_ch1_txsz[0] , _u0_ch1_adr0[31] , _u0_ch1_adr0[30] ,_u0_ch1_adr0[29] , _u0_ch1_adr0[28] , _u0_ch1_adr0[27] ,_u0_ch1_adr0[26] , _u0_ch1_adr0[25] , _u0_ch1_adr0[24] ,_u0_ch1_adr0[23] , _u0_ch1_adr0[22] , _u0_ch1_adr0[21] ,_u0_ch1_adr0[20] , _u0_ch1_adr0[19] , _u0_ch1_adr0[18] ,_u0_ch1_adr0[17] , _u0_ch1_adr0[16] , _u0_ch1_adr0[15] ,_u0_ch1_adr0[14] , _u0_ch1_adr0[13] , _u0_ch1_adr0[12] ,_u0_ch1_adr0[11] , _u0_ch1_adr0[10] , _u0_ch1_adr0[9] ,_u0_ch1_adr0[8] , _u0_ch1_adr0[7] , _u0_ch1_adr0[6] ,_u0_ch1_adr0[5] , _u0_ch1_adr0[4] , _u0_ch1_adr0[3] ,_u0_ch1_adr0[2] , _u0_ch1_adr0[1] , _u0_ch1_adr0[0] ,_u0_ch1_adr1[31] , _u0_ch1_adr1[30] , _u0_ch1_adr1[29] ,_u0_ch1_adr1[28] , _u0_ch1_adr1[27] , _u0_ch1_adr1[26] ,_u0_ch1_adr1[25] , _u0_ch1_adr1[24] , _u0_ch1_adr1[23] ,_u0_ch1_adr1[22] , _u0_ch1_adr1[21] , _u0_ch1_adr1[20] ,_u0_ch1_adr1[19] , _u0_ch1_adr1[18] , _u0_ch1_adr1[17] ,_u0_ch1_adr1[16] , _u0_ch1_adr1[15] , _u0_ch1_adr1[14] ,_u0_ch1_adr1[13] , _u0_ch1_adr1[12] , _u0_ch1_adr1[11] ,_u0_ch1_adr1[10] , _u0_ch1_adr1[9] , _u0_ch1_adr1[8] ,_u0_ch1_adr1[7] , _u0_ch1_adr1[6] , _u0_ch1_adr1[5] ,_u0_ch1_adr1[4] , _u0_ch1_adr1[3] , _u0_ch1_adr1[2] ,_u0_ch1_adr1[1] , _u0_ch1_adr1[0] , _u0_ch1_am0[31] ,_u0_ch1_am0[30] , _u0_ch1_am0[29] , _u0_ch1_am0[28] ,_u0_ch1_am0[27] , _u0_ch1_am0[26] , _u0_ch1_am0[25] ,_u0_ch1_am0[24] , _u0_ch1_am0[23] , _u0_ch1_am0[22] ,_u0_ch1_am0[21] , _u0_ch1_am0[20] , _u0_ch1_am0[19] ,_u0_ch1_am0[18] , _u0_ch1_am0[17] , _u0_ch1_am0[16] ,_u0_ch1_am0[15] , _u0_ch1_am0[14] , _u0_ch1_am0[13] ,_u0_ch1_am0[12] , _u0_ch1_am0[11] , _u0_ch1_am0[10] , _u0_ch1_am0[9] ,_u0_ch1_am0[8] , _u0_ch1_am0[7] , _u0_ch1_am0[6] , _u0_ch1_am0[5] ,_u0_ch1_am0[4] , _u0_ch1_am0[3] , _u0_ch1_am0[2] , _u0_ch1_am0[1] ,_u0_ch1_am0[0] , _u0_ch1_am1[31] , _u0_ch1_am1[30] , _u0_ch1_am1[29] ,_u0_ch1_am1[28] , _u0_ch1_am1[27] , _u0_ch1_am1[26] ,_u0_ch1_am1[25] , _u0_ch1_am1[24] , _u0_ch1_am1[23] ,_u0_ch1_am1[22] , _u0_ch1_am1[21] , _u0_ch1_am1[20] ,_u0_ch1_am1[19] , _u0_ch1_am1[18] , _u0_ch1_am1[17] ,_u0_ch1_am1[16] , _u0_ch1_am1[15] , _u0_ch1_am1[14] ,_u0_ch1_am1[13] , _u0_ch1_am1[12] , _u0_ch1_am1[11] ,_u0_ch1_am1[10] , _u0_ch1_am1[9] , _u0_ch1_am1[8] , _u0_ch1_am1[7] ,_u0_ch1_am1[6] , _u0_ch1_am1[5] , _u0_ch1_am1[4] , _u0_ch1_am1[3] ,_u0_ch1_am1[2] , _u0_ch1_am1[1] , _u0_ch1_am1[0] , _u0_pointer2[31] ,_u0_pointer2[30] , _u0_pointer2[29] , _u0_pointer2[28] ,_u0_pointer2[27] , _u0_pointer2[26] , _u0_pointer2[25] ,_u0_pointer2[24] , _u0_pointer2[23] , _u0_pointer2[22] ,_u0_pointer2[21] , _u0_pointer2[20] , _u0_pointer2[19] ,_u0_pointer2[18] , _u0_pointer2[17] , _u0_pointer2[16] ,_u0_pointer2[15] , _u0_pointer2[14] , _u0_pointer2[13] ,_u0_pointer2[12] , _u0_pointer2[11] , _u0_pointer2[10] ,_u0_pointer2[9] , _u0_pointer2[8] , _u0_pointer2[7] ,_u0_pointer2[6] , _u0_pointer2[5] , _u0_pointer2[4] ,_u0_pointer2[3] , _u0_pointer2[2] , _u0_pointer2[1] ,_u0_pointer2[0] , _u0_pointer2_s[31] , _u0_pointer2_s[30] ,_u0_pointer2_s[29] , _u0_pointer2_s[28] , _u0_pointer2_s[27] ,_u0_pointer2_s[26] , _u0_pointer2_s[25] , _u0_pointer2_s[24] ,_u0_pointer2_s[23] , _u0_pointer2_s[22] , _u0_pointer2_s[21] ,_u0_pointer2_s[20] , _u0_pointer2_s[19] , _u0_pointer2_s[18] ,_u0_pointer2_s[17] , _u0_pointer2_s[16] , _u0_pointer2_s[15] ,_u0_pointer2_s[14] , _u0_pointer2_s[13] , _u0_pointer2_s[12] ,_u0_pointer2_s[11] , _u0_pointer2_s[10] , _u0_pointer2_s[9] ,_u0_pointer2_s[8] , _u0_pointer2_s[7] , _u0_pointer2_s[6] ,_u0_pointer2_s[5] , _u0_pointer2_s[4] , _u0_pointer2_s[3] ,_u0_pointer2_s[2] , _u0_pointer2_s[1] , _u0_pointer2_s[0] ,_u0_ch2_csr[31] , _u0_ch2_csr[30] , _u0_ch2_csr[29] ,_u0_ch2_csr[28] , _u0_ch2_csr[27] , _u0_ch2_csr[26] ,_u0_ch2_csr[25] , _u0_ch2_csr[24] , _u0_ch2_csr[23] ,_u0_ch2_csr[22] , _u0_ch2_csr[21] , _u0_ch2_csr[20] ,_u0_ch2_csr[19] , _u0_ch2_csr[18] , _u0_ch2_csr[17] ,_u0_ch2_csr[16] , _u0_ch2_csr[15] , _u0_ch2_csr[14] ,_u0_ch2_csr[13] , _u0_ch2_csr[12] , _u0_ch2_csr[11] ,_u0_ch2_csr[10] , _u0_ch2_csr[9] , _u0_ch2_csr[8] , _u0_ch2_csr[7] ,_u0_ch2_csr[6] , _u0_ch2_csr[5] , _u0_ch2_csr[4] , _u0_ch2_csr[3] ,_u0_ch2_csr[2] , _u0_ch2_csr[1] , _u0_ch2_csr[0] , _u0_ch2_txsz[31] ,_u0_ch2_txsz[30] , _u0_ch2_txsz[29] , _u0_ch2_txsz[28] ,_u0_ch2_txsz[27] , _u0_ch2_txsz[26] , _u0_ch2_txsz[25] ,_u0_ch2_txsz[24] , _u0_ch2_txsz[23] , _u0_ch2_txsz[22] ,_u0_ch2_txsz[21] , _u0_ch2_txsz[20] , _u0_ch2_txsz[19] ,_u0_ch2_txsz[18] , _u0_ch2_txsz[17] , _u0_ch2_txsz[16] ,_u0_ch2_txsz[15] , _u0_ch2_txsz[14] , _u0_ch2_txsz[13] ,_u0_ch2_txsz[12] , _u0_ch2_txsz[11] , _u0_ch2_txsz[10] ,_u0_ch2_txsz[9] , _u0_ch2_txsz[8] , _u0_ch2_txsz[7] ,_u0_ch2_txsz[6] , _u0_ch2_txsz[5] , _u0_ch2_txsz[4] ,_u0_ch2_txsz[3] , _u0_ch2_txsz[2] , _u0_ch2_txsz[1] ,_u0_ch2_txsz[0] , _u0_ch2_adr0[31] , _u0_ch2_adr0[30] ,_u0_ch2_adr0[29] , _u0_ch2_adr0[28] , _u0_ch2_adr0[27] ,_u0_ch2_adr0[26] , _u0_ch2_adr0[25] , _u0_ch2_adr0[24] ,_u0_ch2_adr0[23] , _u0_ch2_adr0[22] , _u0_ch2_adr0[21] ,_u0_ch2_adr0[20] , _u0_ch2_adr0[19] , _u0_ch2_adr0[18] ,_u0_ch2_adr0[17] , _u0_ch2_adr0[16] , _u0_ch2_adr0[15] ,_u0_ch2_adr0[14] , _u0_ch2_adr0[13] , _u0_ch2_adr0[12] ,_u0_ch2_adr0[11] , _u0_ch2_adr0[10] , _u0_ch2_adr0[9] ,_u0_ch2_adr0[8] , _u0_ch2_adr0[7] , _u0_ch2_adr0[6] ,_u0_ch2_adr0[5] , _u0_ch2_adr0[4] , _u0_ch2_adr0[3] ,_u0_ch2_adr0[2] , _u0_ch2_adr0[1] , _u0_ch2_adr0[0] ,_u0_ch2_adr1[31] , _u0_ch2_adr1[30] , _u0_ch2_adr1[29] ,_u0_ch2_adr1[28] , _u0_ch2_adr1[27] , _u0_ch2_adr1[26] ,_u0_ch2_adr1[25] , _u0_ch2_adr1[24] , _u0_ch2_adr1[23] ,_u0_ch2_adr1[22] , _u0_ch2_adr1[21] , _u0_ch2_adr1[20] ,_u0_ch2_adr1[19] , _u0_ch2_adr1[18] , _u0_ch2_adr1[17] ,_u0_ch2_adr1[16] , _u0_ch2_adr1[15] , _u0_ch2_adr1[14] ,_u0_ch2_adr1[13] , _u0_ch2_adr1[12] , _u0_ch2_adr1[11] ,_u0_ch2_adr1[10] , _u0_ch2_adr1[9] , _u0_ch2_adr1[8] ,_u0_ch2_adr1[7] , _u0_ch2_adr1[6] , _u0_ch2_adr1[5] ,_u0_ch2_adr1[4] , _u0_ch2_adr1[3] , _u0_ch2_adr1[2] ,_u0_ch2_adr1[1] , _u0_ch2_adr1[0] , _u0_ch2_am0[31] ,_u0_ch2_am0[30] , _u0_ch2_am0[29] , _u0_ch2_am0[28] ,_u0_ch2_am0[27] , _u0_ch2_am0[26] , _u0_ch2_am0[25] ,_u0_ch2_am0[24] , _u0_ch2_am0[23] , _u0_ch2_am0[22] ,_u0_ch2_am0[21] , _u0_ch2_am0[20] , _u0_ch2_am0[19] ,_u0_ch2_am0[18] , _u0_ch2_am0[17] , _u0_ch2_am0[16] ,_u0_ch2_am0[15] , _u0_ch2_am0[14] , _u0_ch2_am0[13] ,_u0_ch2_am0[12] , _u0_ch2_am0[11] , _u0_ch2_am0[10] , _u0_ch2_am0[9] ,_u0_ch2_am0[8] , _u0_ch2_am0[7] , _u0_ch2_am0[6] , _u0_ch2_am0[5] ,_u0_ch2_am0[4] , _u0_ch2_am0[3] , _u0_ch2_am0[2] , _u0_ch2_am0[1] ,_u0_ch2_am0[0] , _u0_ch2_am1[31] , _u0_ch2_am1[30] , _u0_ch2_am1[29] ,_u0_ch2_am1[28] , _u0_ch2_am1[27] , _u0_ch2_am1[26] ,_u0_ch2_am1[25] , _u0_ch2_am1[24] , _u0_ch2_am1[23] ,_u0_ch2_am1[22] , _u0_ch2_am1[21] , _u0_ch2_am1[20] ,_u0_ch2_am1[19] , _u0_ch2_am1[18] , _u0_ch2_am1[17] ,_u0_ch2_am1[16] , _u0_ch2_am1[15] , _u0_ch2_am1[14] ,_u0_ch2_am1[13] , _u0_ch2_am1[12] , _u0_ch2_am1[11] ,_u0_ch2_am1[10] , _u0_ch2_am1[9] , _u0_ch2_am1[8] , _u0_ch2_am1[7] ,_u0_ch2_am1[6] , _u0_ch2_am1[5] , _u0_ch2_am1[4] , _u0_ch2_am1[3] ,_u0_ch2_am1[2] , _u0_ch2_am1[1] , _u0_ch2_am1[0] , _u0_pointer3[31] ,_u0_pointer3[30] , _u0_pointer3[29] , _u0_pointer3[28] ,_u0_pointer3[27] , _u0_pointer3[26] , _u0_pointer3[25] ,_u0_pointer3[24] , _u0_pointer3[23] , _u0_pointer3[22] ,_u0_pointer3[21] , _u0_pointer3[20] , _u0_pointer3[19] ,_u0_pointer3[18] , _u0_pointer3[17] , _u0_pointer3[16] ,_u0_pointer3[15] , _u0_pointer3[14] , _u0_pointer3[13] ,_u0_pointer3[12] , _u0_pointer3[11] , _u0_pointer3[10] ,_u0_pointer3[9] , _u0_pointer3[8] , _u0_pointer3[7] ,_u0_pointer3[6] , _u0_pointer3[5] , _u0_pointer3[4] ,_u0_pointer3[3] , _u0_pointer3[2] , _u0_pointer3[1] ,_u0_pointer3[0] , _u0_pointer3_s[31] , _u0_pointer3_s[30] ,_u0_pointer3_s[29] , _u0_pointer3_s[28] , _u0_pointer3_s[27] ,_u0_pointer3_s[26] , _u0_pointer3_s[25] , _u0_pointer3_s[24] ,_u0_pointer3_s[23] , _u0_pointer3_s[22] , _u0_pointer3_s[21] ,_u0_pointer3_s[20] , _u0_pointer3_s[19] , _u0_pointer3_s[18] ,_u0_pointer3_s[17] , _u0_pointer3_s[16] , _u0_pointer3_s[15] ,_u0_pointer3_s[14] , _u0_pointer3_s[13] , _u0_pointer3_s[12] ,_u0_pointer3_s[11] , _u0_pointer3_s[10] , _u0_pointer3_s[9] ,_u0_pointer3_s[8] , _u0_pointer3_s[7] , _u0_pointer3_s[6] ,_u0_pointer3_s[5] , _u0_pointer3_s[4] , _u0_pointer3_s[3] ,_u0_pointer3_s[2] , _u0_pointer3_s[1] , _u0_pointer3_s[0] ,_u0_ch3_csr[31] , _u0_ch3_csr[30] , _u0_ch3_csr[29] ,_u0_ch3_csr[28] , _u0_ch3_csr[27] , _u0_ch3_csr[26] ,_u0_ch3_csr[25] , _u0_ch3_csr[24] , _u0_ch3_csr[23] ,_u0_ch3_csr[22] , _u0_ch3_csr[21] , _u0_ch3_csr[20] ,_u0_ch3_csr[19] , _u0_ch3_csr[18] , _u0_ch3_csr[17] ,_u0_ch3_csr[16] , _u0_ch3_csr[15] , _u0_ch3_csr[14] ,_u0_ch3_csr[13] , _u0_ch3_csr[12] , _u0_ch3_csr[11] ,_u0_ch3_csr[10] , _u0_ch3_csr[9] , _u0_ch3_csr[8] , _u0_ch3_csr[7] ,_u0_ch3_csr[6] , _u0_ch3_csr[5] , _u0_ch3_csr[4] , _u0_ch3_csr[3] ,_u0_ch3_csr[2] , _u0_ch3_csr[1] , _u0_ch3_csr[0] , _u0_ch3_txsz[31] ,_u0_ch3_txsz[30] , _u0_ch3_txsz[29] , _u0_ch3_txsz[28] ,_u0_ch3_txsz[27] , _u0_ch3_txsz[26] , _u0_ch3_txsz[25] ,_u0_ch3_txsz[24] , _u0_ch3_txsz[23] , _u0_ch3_txsz[22] ,_u0_ch3_txsz[21] , _u0_ch3_txsz[20] , _u0_ch3_txsz[19] ,_u0_ch3_txsz[18] , _u0_ch3_txsz[17] , _u0_ch3_txsz[16] ,_u0_ch3_txsz[15] , _u0_ch3_txsz[14] , _u0_ch3_txsz[13] ,_u0_ch3_txsz[12] , _u0_ch3_txsz[11] , _u0_ch3_txsz[10] ,_u0_ch3_txsz[9] , _u0_ch3_txsz[8] , _u0_ch3_txsz[7] ,_u0_ch3_txsz[6] , _u0_ch3_txsz[5] , _u0_ch3_txsz[4] ,_u0_ch3_txsz[3] , _u0_ch3_txsz[2] , _u0_ch3_txsz[1] ,_u0_ch3_txsz[0] , _u0_ch3_adr0[31] , _u0_ch3_adr0[30] ,_u0_ch3_adr0[29] , _u0_ch3_adr0[28] , _u0_ch3_adr0[27] ,_u0_ch3_adr0[26] , _u0_ch3_adr0[25] , _u0_ch3_adr0[24] ,_u0_ch3_adr0[23] , _u0_ch3_adr0[22] , _u0_ch3_adr0[21] ,_u0_ch3_adr0[20] , _u0_ch3_adr0[19] , _u0_ch3_adr0[18] ,_u0_ch3_adr0[17] , _u0_ch3_adr0[16] , _u0_ch3_adr0[15] ,_u0_ch3_adr0[14] , _u0_ch3_adr0[13] , _u0_ch3_adr0[12] ,_u0_ch3_adr0[11] , _u0_ch3_adr0[10] , _u0_ch3_adr0[9] ,_u0_ch3_adr0[8] , _u0_ch3_adr0[7] , _u0_ch3_adr0[6] ,_u0_ch3_adr0[5] , _u0_ch3_adr0[4] , _u0_ch3_adr0[3] ,_u0_ch3_adr0[2] , _u0_ch3_adr0[1] , _u0_ch3_adr0[0] ,_u0_ch3_adr1[31] , _u0_ch3_adr1[30] , _u0_ch3_adr1[29] ,_u0_ch3_adr1[28] , _u0_ch3_adr1[27] , _u0_ch3_adr1[26] ,_u0_ch3_adr1[25] , _u0_ch3_adr1[24] , _u0_ch3_adr1[23] ,_u0_ch3_adr1[22] , _u0_ch3_adr1[21] , _u0_ch3_adr1[20] ,_u0_ch3_adr1[19] , _u0_ch3_adr1[18] , _u0_ch3_adr1[17] ,_u0_ch3_adr1[16] , _u0_ch3_adr1[15] , _u0_ch3_adr1[14] ,_u0_ch3_adr1[13] , _u0_ch3_adr1[12] , _u0_ch3_adr1[11] ,_u0_ch3_adr1[10] , _u0_ch3_adr1[9] , _u0_ch3_adr1[8] ,_u0_ch3_adr1[7] , _u0_ch3_adr1[6] , _u0_ch3_adr1[5] ,_u0_ch3_adr1[4] , _u0_ch3_adr1[3] , _u0_ch3_adr1[2] ,_u0_ch3_adr1[1] , _u0_ch3_adr1[0] , _u0_ch3_am0[31] ,_u0_ch3_am0[30] , _u0_ch3_am0[29] , _u0_ch3_am0[28] ,_u0_ch3_am0[27] , _u0_ch3_am0[26] , _u0_ch3_am0[25] ,_u0_ch3_am0[24] , _u0_ch3_am0[23] , _u0_ch3_am0[22] ,_u0_ch3_am0[21] , _u0_ch3_am0[20] , _u0_ch3_am0[19] ,_u0_ch3_am0[18] , _u0_ch3_am0[17] , _u0_ch3_am0[16] ,_u0_ch3_am0[15] , _u0_ch3_am0[14] , _u0_ch3_am0[13] ,_u0_ch3_am0[12] , _u0_ch3_am0[11] , _u0_ch3_am0[10] , _u0_ch3_am0[9] ,_u0_ch3_am0[8] , _u0_ch3_am0[7] , _u0_ch3_am0[6] , _u0_ch3_am0[5] ,_u0_ch3_am0[4] , _u0_ch3_am0[3] , _u0_ch3_am0[2] , _u0_ch3_am0[1] ,_u0_ch3_am0[0] , _u0_ch3_am1[31] , _u0_ch3_am1[30] , _u0_ch3_am1[29] ,_u0_ch3_am1[28] , _u0_ch3_am1[27] , _u0_ch3_am1[26] ,_u0_ch3_am1[25] , _u0_ch3_am1[24] , _u0_ch3_am1[23] ,_u0_ch3_am1[22] , _u0_ch3_am1[21] , _u0_ch3_am1[20] ,_u0_ch3_am1[19] , _u0_ch3_am1[18] , _u0_ch3_am1[17] ,_u0_ch3_am1[16] , _u0_ch3_am1[15] , _u0_ch3_am1[14] ,_u0_ch3_am1[13] , _u0_ch3_am1[12] , _u0_ch3_am1[11] ,_u0_ch3_am1[10] , _u0_ch3_am1[9] , _u0_ch3_am1[8] , _u0_ch3_am1[7] ,_u0_ch3_am1[6] , _u0_ch3_am1[5] , _u0_ch3_am1[4] , _u0_ch3_am1[3] ,_u0_ch3_am1[2] , _u0_ch3_am1[1] , _u0_ch3_am1[0] , _u0_pointer4[31] ,_u0_pointer4[30] , _u0_pointer4[29] , _u0_pointer4[28] ,_u0_pointer4[27] , _u0_pointer4[26] , _u0_pointer4[25] ,_u0_pointer4[24] , _u0_pointer4[23] , _u0_pointer4[22] ,_u0_pointer4[21] , _u0_pointer4[20] , _u0_pointer4[19] ,_u0_pointer4[18] , _u0_pointer4[17] , _u0_pointer4[16] ,_u0_pointer4[15] , _u0_pointer4[14] , _u0_pointer4[13] ,_u0_pointer4[12] , _u0_pointer4[11] , _u0_pointer4[10] ,_u0_pointer4[9] , _u0_pointer4[8] , _u0_pointer4[7] ,_u0_pointer4[6] , _u0_pointer4[5] , _u0_pointer4[4] ,_u0_pointer4[3] , _u0_pointer4[2] , _u0_pointer4[1] ,_u0_pointer4[0] , _u0_pointer4_s[31] , _u0_pointer4_s[30] ,_u0_pointer4_s[29] , _u0_pointer4_s[28] , _u0_pointer4_s[27] ,_u0_pointer4_s[26] , _u0_pointer4_s[25] , _u0_pointer4_s[24] ,_u0_pointer4_s[23] , _u0_pointer4_s[22] , _u0_pointer4_s[21] ,_u0_pointer4_s[20] , _u0_pointer4_s[19] , _u0_pointer4_s[18] ,_u0_pointer4_s[17] , _u0_pointer4_s[16] , _u0_pointer4_s[15] ,_u0_pointer4_s[14] , _u0_pointer4_s[13] , _u0_pointer4_s[12] ,_u0_pointer4_s[11] , _u0_pointer4_s[10] , _u0_pointer4_s[9] ,_u0_pointer4_s[8] , _u0_pointer4_s[7] , _u0_pointer4_s[6] ,_u0_pointer4_s[5] , _u0_pointer4_s[4] , _u0_pointer4_s[3] ,_u0_pointer4_s[2] , _u0_pointer4_s[1] , _u0_pointer4_s[0] ,_u0_ch4_csr[31] , _u0_ch4_csr[30] , _u0_ch4_csr[29] ,_u0_ch4_csr[28] , _u0_ch4_csr[27] , _u0_ch4_csr[26] ,_u0_ch4_csr[25] , _u0_ch4_csr[24] , _u0_ch4_csr[23] ,_u0_ch4_csr[22] , _u0_ch4_csr[21] , _u0_ch4_csr[20] ,_u0_ch4_csr[19] , _u0_ch4_csr[18] , _u0_ch4_csr[17] ,_u0_ch4_csr[16] , _u0_ch4_csr[15] , _u0_ch4_csr[14] ,_u0_ch4_csr[13] , _u0_ch4_csr[12] , _u0_ch4_csr[11] ,_u0_ch4_csr[10] , _u0_ch4_csr[9] , _u0_ch4_csr[8] , _u0_ch4_csr[7] ,_u0_ch4_csr[6] , _u0_ch4_csr[5] , _u0_ch4_csr[4] , _u0_ch4_csr[3] ,_u0_ch4_csr[2] , _u0_ch4_csr[1] , _u0_ch4_csr[0] , _u0_ch4_txsz[31] ,_u0_ch4_txsz[30] , _u0_ch4_txsz[29] , _u0_ch4_txsz[28] ,_u0_ch4_txsz[27] , _u0_ch4_txsz[26] , _u0_ch4_txsz[25] ,_u0_ch4_txsz[24] , _u0_ch4_txsz[23] , _u0_ch4_txsz[22] ,_u0_ch4_txsz[21] , _u0_ch4_txsz[20] , _u0_ch4_txsz[19] ,_u0_ch4_txsz[18] , _u0_ch4_txsz[17] , _u0_ch4_txsz[16] ,_u0_ch4_txsz[15] , _u0_ch4_txsz[14] , _u0_ch4_txsz[13] ,_u0_ch4_txsz[12] , _u0_ch4_txsz[11] , _u0_ch4_txsz[10] ,_u0_ch4_txsz[9] , _u0_ch4_txsz[8] , _u0_ch4_txsz[7] ,_u0_ch4_txsz[6] , _u0_ch4_txsz[5] , _u0_ch4_txsz[4] ,_u0_ch4_txsz[3] , _u0_ch4_txsz[2] , _u0_ch4_txsz[1] ,_u0_ch4_txsz[0] , _u0_ch4_adr0[31] , _u0_ch4_adr0[30] ,_u0_ch4_adr0[29] , _u0_ch4_adr0[28] , _u0_ch4_adr0[27] ,_u0_ch4_adr0[26] , _u0_ch4_adr0[25] , _u0_ch4_adr0[24] ,_u0_ch4_adr0[23] , _u0_ch4_adr0[22] , _u0_ch4_adr0[21] ,_u0_ch4_adr0[20] , _u0_ch4_adr0[19] , _u0_ch4_adr0[18] ,_u0_ch4_adr0[17] , _u0_ch4_adr0[16] , _u0_ch4_adr0[15] ,_u0_ch4_adr0[14] , _u0_ch4_adr0[13] , _u0_ch4_adr0[12] ,_u0_ch4_adr0[11] , _u0_ch4_adr0[10] , _u0_ch4_adr0[9] ,_u0_ch4_adr0[8] , _u0_ch4_adr0[7] , _u0_ch4_adr0[6] ,_u0_ch4_adr0[5] , _u0_ch4_adr0[4] , _u0_ch4_adr0[3] ,_u0_ch4_adr0[2] , _u0_ch4_adr0[1] , _u0_ch4_adr0[0] ,_u0_ch4_adr1[31] , _u0_ch4_adr1[30] , _u0_ch4_adr1[29] ,_u0_ch4_adr1[28] , _u0_ch4_adr1[27] , _u0_ch4_adr1[26] ,_u0_ch4_adr1[25] , _u0_ch4_adr1[24] , _u0_ch4_adr1[23] ,_u0_ch4_adr1[22] , _u0_ch4_adr1[21] , _u0_ch4_adr1[20] ,_u0_ch4_adr1[19] , _u0_ch4_adr1[18] , _u0_ch4_adr1[17] ,_u0_ch4_adr1[16] , _u0_ch4_adr1[15] , _u0_ch4_adr1[14] ,_u0_ch4_adr1[13] , _u0_ch4_adr1[12] , _u0_ch4_adr1[11] ,_u0_ch4_adr1[10] , _u0_ch4_adr1[9] , _u0_ch4_adr1[8] ,_u0_ch4_adr1[7] , _u0_ch4_adr1[6] , _u0_ch4_adr1[5] ,_u0_ch4_adr1[4] , _u0_ch4_adr1[3] , _u0_ch4_adr1[2] ,_u0_ch4_adr1[1] , _u0_ch4_adr1[0] , _u0_ch4_am0[31] ,_u0_ch4_am0[30] , _u0_ch4_am0[29] , _u0_ch4_am0[28] ,_u0_ch4_am0[27] , _u0_ch4_am0[26] , _u0_ch4_am0[25] ,_u0_ch4_am0[24] , _u0_ch4_am0[23] , _u0_ch4_am0[22] ,_u0_ch4_am0[21] , _u0_ch4_am0[20] , _u0_ch4_am0[19] ,_u0_ch4_am0[18] , _u0_ch4_am0[17] , _u0_ch4_am0[16] ,_u0_ch4_am0[15] , _u0_ch4_am0[14] , _u0_ch4_am0[13] ,_u0_ch4_am0[12] , _u0_ch4_am0[11] , _u0_ch4_am0[10] , _u0_ch4_am0[9] ,_u0_ch4_am0[8] , _u0_ch4_am0[7] , _u0_ch4_am0[6] , _u0_ch4_am0[5] ,_u0_ch4_am0[4] , _u0_ch4_am0[3] , _u0_ch4_am0[2] , _u0_ch4_am0[1] ,_u0_ch4_am0[0] , _u0_ch4_am1[31] , _u0_ch4_am1[30] , _u0_ch4_am1[29] ,_u0_ch4_am1[28] , _u0_ch4_am1[27] , _u0_ch4_am1[26] ,_u0_ch4_am1[25] , _u0_ch4_am1[24] , _u0_ch4_am1[23] ,_u0_ch4_am1[22] , _u0_ch4_am1[21] , _u0_ch4_am1[20] ,_u0_ch4_am1[19] , _u0_ch4_am1[18] , _u0_ch4_am1[17] ,_u0_ch4_am1[16] , _u0_ch4_am1[15] , _u0_ch4_am1[14] ,_u0_ch4_am1[13] , _u0_ch4_am1[12] , _u0_ch4_am1[11] ,_u0_ch4_am1[10] , _u0_ch4_am1[9] , _u0_ch4_am1[8] , _u0_ch4_am1[7] ,_u0_ch4_am1[6] , _u0_ch4_am1[5] , _u0_ch4_am1[4] , _u0_ch4_am1[3] ,_u0_ch4_am1[2] , _u0_ch4_am1[1] , _u0_ch4_am1[0] , _u0_pointer5[31] ,_u0_pointer5[30] , _u0_pointer5[29] , _u0_pointer5[28] ,_u0_pointer5[27] , _u0_pointer5[26] , _u0_pointer5[25] ,_u0_pointer5[24] , _u0_pointer5[23] , _u0_pointer5[22] ,_u0_pointer5[21] , _u0_pointer5[20] , _u0_pointer5[19] ,_u0_pointer5[18] , _u0_pointer5[17] , _u0_pointer5[16] ,_u0_pointer5[15] , _u0_pointer5[14] , _u0_pointer5[13] ,_u0_pointer5[12] , _u0_pointer5[11] , _u0_pointer5[10] ,_u0_pointer5[9] , _u0_pointer5[8] , _u0_pointer5[7] ,_u0_pointer5[6] , _u0_pointer5[5] , _u0_pointer5[4] ,_u0_pointer5[3] , _u0_pointer5[2] , _u0_pointer5[1] ,_u0_pointer5[0] , _u0_pointer5_s[31] , _u0_pointer5_s[30] ,_u0_pointer5_s[29] , _u0_pointer5_s[28] , _u0_pointer5_s[27] ,_u0_pointer5_s[26] , _u0_pointer5_s[25] , _u0_pointer5_s[24] ,_u0_pointer5_s[23] , _u0_pointer5_s[22] , _u0_pointer5_s[21] ,_u0_pointer5_s[20] , _u0_pointer5_s[19] , _u0_pointer5_s[18] ,_u0_pointer5_s[17] , _u0_pointer5_s[16] , _u0_pointer5_s[15] ,_u0_pointer5_s[14] , _u0_pointer5_s[13] , _u0_pointer5_s[12] ,_u0_pointer5_s[11] , _u0_pointer5_s[10] , _u0_pointer5_s[9] ,_u0_pointer5_s[8] , _u0_pointer5_s[7] , _u0_pointer5_s[6] ,_u0_pointer5_s[5] , _u0_pointer5_s[4] , _u0_pointer5_s[3] ,_u0_pointer5_s[2] , _u0_pointer5_s[1] , _u0_pointer5_s[0] ,_u0_ch5_csr[31] , _u0_ch5_csr[30] , _u0_ch5_csr[29] ,_u0_ch5_csr[28] , _u0_ch5_csr[27] , _u0_ch5_csr[26] ,_u0_ch5_csr[25] , _u0_ch5_csr[24] , _u0_ch5_csr[23] ,_u0_ch5_csr[22] , _u0_ch5_csr[21] , _u0_ch5_csr[20] ,_u0_ch5_csr[19] , _u0_ch5_csr[18] , _u0_ch5_csr[17] ,_u0_ch5_csr[16] , _u0_ch5_csr[15] , _u0_ch5_csr[14] ,_u0_ch5_csr[13] , _u0_ch5_csr[12] , _u0_ch5_csr[11] ,_u0_ch5_csr[10] , _u0_ch5_csr[9] , _u0_ch5_csr[8] , _u0_ch5_csr[7] ,_u0_ch5_csr[6] , _u0_ch5_csr[5] , _u0_ch5_csr[4] , _u0_ch5_csr[3] ,_u0_ch5_csr[2] , _u0_ch5_csr[1] , _u0_ch5_csr[0] , _u0_ch5_txsz[31] ,_u0_ch5_txsz[30] , _u0_ch5_txsz[29] , _u0_ch5_txsz[28] ,_u0_ch5_txsz[27] , _u0_ch5_txsz[26] , _u0_ch5_txsz[25] ,_u0_ch5_txsz[24] , _u0_ch5_txsz[23] , _u0_ch5_txsz[22] ,_u0_ch5_txsz[21] , _u0_ch5_txsz[20] , _u0_ch5_txsz[19] ,_u0_ch5_txsz[18] , _u0_ch5_txsz[17] , _u0_ch5_txsz[16] ,_u0_ch5_txsz[15] , _u0_ch5_txsz[14] , _u0_ch5_txsz[13] ,_u0_ch5_txsz[12] , _u0_ch5_txsz[11] , _u0_ch5_txsz[10] ,_u0_ch5_txsz[9] , _u0_ch5_txsz[8] , _u0_ch5_txsz[7] ,_u0_ch5_txsz[6] , _u0_ch5_txsz[5] , _u0_ch5_txsz[4] ,_u0_ch5_txsz[3] , _u0_ch5_txsz[2] , _u0_ch5_txsz[1] ,_u0_ch5_txsz[0] , _u0_ch5_adr0[31] , _u0_ch5_adr0[30] ,_u0_ch5_adr0[29] , _u0_ch5_adr0[28] , _u0_ch5_adr0[27] ,_u0_ch5_adr0[26] , _u0_ch5_adr0[25] , _u0_ch5_adr0[24] ,_u0_ch5_adr0[23] , _u0_ch5_adr0[22] , _u0_ch5_adr0[21] ,_u0_ch5_adr0[20] , _u0_ch5_adr0[19] , _u0_ch5_adr0[18] ,_u0_ch5_adr0[17] , _u0_ch5_adr0[16] , _u0_ch5_adr0[15] ,_u0_ch5_adr0[14] , _u0_ch5_adr0[13] , _u0_ch5_adr0[12] ,_u0_ch5_adr0[11] , _u0_ch5_adr0[10] , _u0_ch5_adr0[9] ,_u0_ch5_adr0[8] , _u0_ch5_adr0[7] , _u0_ch5_adr0[6] ,_u0_ch5_adr0[5] , _u0_ch5_adr0[4] , _u0_ch5_adr0[3] ,_u0_ch5_adr0[2] , _u0_ch5_adr0[1] , _u0_ch5_adr0[0] ,_u0_ch5_adr1[31] , _u0_ch5_adr1[30] , _u0_ch5_adr1[29] ,_u0_ch5_adr1[28] , _u0_ch5_adr1[27] , _u0_ch5_adr1[26] ,_u0_ch5_adr1[25] , _u0_ch5_adr1[24] , _u0_ch5_adr1[23] ,_u0_ch5_adr1[22] , _u0_ch5_adr1[21] , _u0_ch5_adr1[20] ,_u0_ch5_adr1[19] , _u0_ch5_adr1[18] , _u0_ch5_adr1[17] ,_u0_ch5_adr1[16] , _u0_ch5_adr1[15] , _u0_ch5_adr1[14] ,_u0_ch5_adr1[13] , _u0_ch5_adr1[12] , _u0_ch5_adr1[11] ,_u0_ch5_adr1[10] , _u0_ch5_adr1[9] , _u0_ch5_adr1[8] ,_u0_ch5_adr1[7] , _u0_ch5_adr1[6] , _u0_ch5_adr1[5] ,_u0_ch5_adr1[4] , _u0_ch5_adr1[3] , _u0_ch5_adr1[2] ,_u0_ch5_adr1[1] , _u0_ch5_adr1[0] , _u0_ch5_am0[31] ,_u0_ch5_am0[30] , _u0_ch5_am0[29] , _u0_ch5_am0[28] ,_u0_ch5_am0[27] , _u0_ch5_am0[26] , _u0_ch5_am0[25] ,_u0_ch5_am0[24] , _u0_ch5_am0[23] , _u0_ch5_am0[22] ,_u0_ch5_am0[21] , _u0_ch5_am0[20] , _u0_ch5_am0[19] ,_u0_ch5_am0[18] , _u0_ch5_am0[17] , _u0_ch5_am0[16] ,_u0_ch5_am0[15] , _u0_ch5_am0[14] , _u0_ch5_am0[13] ,_u0_ch5_am0[12] , _u0_ch5_am0[11] , _u0_ch5_am0[10] , _u0_ch5_am0[9] ,_u0_ch5_am0[8] , _u0_ch5_am0[7] , _u0_ch5_am0[6] , _u0_ch5_am0[5] ,_u0_ch5_am0[4] , _u0_ch5_am0[3] , _u0_ch5_am0[2] , _u0_ch5_am0[1] ,_u0_ch5_am0[0] , _u0_ch5_am1[31] , _u0_ch5_am1[30] , _u0_ch5_am1[29] ,_u0_ch5_am1[28] , _u0_ch5_am1[27] , _u0_ch5_am1[26] ,_u0_ch5_am1[25] , _u0_ch5_am1[24] , _u0_ch5_am1[23] ,_u0_ch5_am1[22] , _u0_ch5_am1[21] , _u0_ch5_am1[20] ,_u0_ch5_am1[19] , _u0_ch5_am1[18] , _u0_ch5_am1[17] ,_u0_ch5_am1[16] , _u0_ch5_am1[15] , _u0_ch5_am1[14] ,_u0_ch5_am1[13] , _u0_ch5_am1[12] , _u0_ch5_am1[11] ,_u0_ch5_am1[10] , _u0_ch5_am1[9] , _u0_ch5_am1[8] , _u0_ch5_am1[7] ,_u0_ch5_am1[6] , _u0_ch5_am1[5] , _u0_ch5_am1[4] , _u0_ch5_am1[3] ,_u0_ch5_am1[2] , _u0_ch5_am1[1] , _u0_ch5_am1[0] , _u0_pointer6[31] ,_u0_pointer6[30] , _u0_pointer6[29] , _u0_pointer6[28] ,_u0_pointer6[27] , _u0_pointer6[26] , _u0_pointer6[25] ,_u0_pointer6[24] , _u0_pointer6[23] , _u0_pointer6[22] ,_u0_pointer6[21] , _u0_pointer6[20] , _u0_pointer6[19] ,_u0_pointer6[18] , _u0_pointer6[17] , _u0_pointer6[16] ,_u0_pointer6[15] , _u0_pointer6[14] , _u0_pointer6[13] ,_u0_pointer6[12] , _u0_pointer6[11] , _u0_pointer6[10] ,_u0_pointer6[9] , _u0_pointer6[8] , _u0_pointer6[7] ,_u0_pointer6[6] , _u0_pointer6[5] , _u0_pointer6[4] ,_u0_pointer6[3] , _u0_pointer6[2] , _u0_pointer6[1] ,_u0_pointer6[0] , _u0_pointer6_s[31] , _u0_pointer6_s[30] ,_u0_pointer6_s[29] , _u0_pointer6_s[28] , _u0_pointer6_s[27] ,_u0_pointer6_s[26] , _u0_pointer6_s[25] , _u0_pointer6_s[24] ,_u0_pointer6_s[23] , _u0_pointer6_s[22] , _u0_pointer6_s[21] ,_u0_pointer6_s[20] , _u0_pointer6_s[19] , _u0_pointer6_s[18] ,_u0_pointer6_s[17] , _u0_pointer6_s[16] , _u0_pointer6_s[15] ,_u0_pointer6_s[14] , _u0_pointer6_s[13] , _u0_pointer6_s[12] ,_u0_pointer6_s[11] , _u0_pointer6_s[10] , _u0_pointer6_s[9] ,_u0_pointer6_s[8] , _u0_pointer6_s[7] , _u0_pointer6_s[6] ,_u0_pointer6_s[5] , _u0_pointer6_s[4] , _u0_pointer6_s[3] ,_u0_pointer6_s[2] , _u0_pointer6_s[1] , _u0_pointer6_s[0] ,_u0_ch6_csr[31] , _u0_ch6_csr[30] , _u0_ch6_csr[29] ,_u0_ch6_csr[28] , _u0_ch6_csr[27] , _u0_ch6_csr[26] ,_u0_ch6_csr[25] , _u0_ch6_csr[24] , _u0_ch6_csr[23] ,_u0_ch6_csr[22] , _u0_ch6_csr[21] , _u0_ch6_csr[20] ,_u0_ch6_csr[19] , _u0_ch6_csr[18] , _u0_ch6_csr[17] ,_u0_ch6_csr[16] , _u0_ch6_csr[15] , _u0_ch6_csr[14] ,_u0_ch6_csr[13] , _u0_ch6_csr[12] , _u0_ch6_csr[11] ,_u0_ch6_csr[10] , _u0_ch6_csr[9] , _u0_ch6_csr[8] , _u0_ch6_csr[7] ,_u0_ch6_csr[6] , _u0_ch6_csr[5] , _u0_ch6_csr[4] , _u0_ch6_csr[3] ,_u0_ch6_csr[2] , _u0_ch6_csr[1] , _u0_ch6_csr[0] , _u0_ch6_txsz[31] ,_u0_ch6_txsz[30] , _u0_ch6_txsz[29] , _u0_ch6_txsz[28] ,_u0_ch6_txsz[27] , _u0_ch6_txsz[26] , _u0_ch6_txsz[25] ,_u0_ch6_txsz[24] , _u0_ch6_txsz[23] , _u0_ch6_txsz[22] ,_u0_ch6_txsz[21] , _u0_ch6_txsz[20] , _u0_ch6_txsz[19] ,_u0_ch6_txsz[18] , _u0_ch6_txsz[17] , _u0_ch6_txsz[16] ,_u0_ch6_txsz[15] , _u0_ch6_txsz[14] , _u0_ch6_txsz[13] ,_u0_ch6_txsz[12] , _u0_ch6_txsz[11] , _u0_ch6_txsz[10] ,_u0_ch6_txsz[9] , _u0_ch6_txsz[8] , _u0_ch6_txsz[7] ,_u0_ch6_txsz[6] , _u0_ch6_txsz[5] , _u0_ch6_txsz[4] ,_u0_ch6_txsz[3] , _u0_ch6_txsz[2] , _u0_ch6_txsz[1] ,_u0_ch6_txsz[0] , _u0_ch6_adr0[31] , _u0_ch6_adr0[30] ,_u0_ch6_adr0[29] , _u0_ch6_adr0[28] , _u0_ch6_adr0[27] ,_u0_ch6_adr0[26] , _u0_ch6_adr0[25] , _u0_ch6_adr0[24] ,_u0_ch6_adr0[23] , _u0_ch6_adr0[22] , _u0_ch6_adr0[21] ,_u0_ch6_adr0[20] , _u0_ch6_adr0[19] , _u0_ch6_adr0[18] ,_u0_ch6_adr0[17] , _u0_ch6_adr0[16] , _u0_ch6_adr0[15] ,_u0_ch6_adr0[14] , _u0_ch6_adr0[13] , _u0_ch6_adr0[12] ,_u0_ch6_adr0[11] , _u0_ch6_adr0[10] , _u0_ch6_adr0[9] ,_u0_ch6_adr0[8] , _u0_ch6_adr0[7] , _u0_ch6_adr0[6] ,_u0_ch6_adr0[5] , _u0_ch6_adr0[4] , _u0_ch6_adr0[3] ,_u0_ch6_adr0[2] , _u0_ch6_adr0[1] , _u0_ch6_adr0[0] ,_u0_ch6_adr1[31] , _u0_ch6_adr1[30] , _u0_ch6_adr1[29] ,_u0_ch6_adr1[28] , _u0_ch6_adr1[27] , _u0_ch6_adr1[26] ,_u0_ch6_adr1[25] , _u0_ch6_adr1[24] , _u0_ch6_adr1[23] ,_u0_ch6_adr1[22] , _u0_ch6_adr1[21] , _u0_ch6_adr1[20] ,_u0_ch6_adr1[19] , _u0_ch6_adr1[18] , _u0_ch6_adr1[17] ,_u0_ch6_adr1[16] , _u0_ch6_adr1[15] , _u0_ch6_adr1[14] ,_u0_ch6_adr1[13] , _u0_ch6_adr1[12] , _u0_ch6_adr1[11] ,_u0_ch6_adr1[10] , _u0_ch6_adr1[9] , _u0_ch6_adr1[8] ,_u0_ch6_adr1[7] , _u0_ch6_adr1[6] , _u0_ch6_adr1[5] ,_u0_ch6_adr1[4] , _u0_ch6_adr1[3] , _u0_ch6_adr1[2] ,_u0_ch6_adr1[1] , _u0_ch6_adr1[0] , _u0_ch6_am0[31] ,_u0_ch6_am0[30] , _u0_ch6_am0[29] , _u0_ch6_am0[28] ,_u0_ch6_am0[27] , _u0_ch6_am0[26] , _u0_ch6_am0[25] ,_u0_ch6_am0[24] , _u0_ch6_am0[23] , _u0_ch6_am0[22] ,_u0_ch6_am0[21] , _u0_ch6_am0[20] , _u0_ch6_am0[19] ,_u0_ch6_am0[18] , _u0_ch6_am0[17] , _u0_ch6_am0[16] ,_u0_ch6_am0[15] , _u0_ch6_am0[14] , _u0_ch6_am0[13] ,_u0_ch6_am0[12] , _u0_ch6_am0[11] , _u0_ch6_am0[10] , _u0_ch6_am0[9] ,_u0_ch6_am0[8] , _u0_ch6_am0[7] , _u0_ch6_am0[6] , _u0_ch6_am0[5] ,_u0_ch6_am0[4] , _u0_ch6_am0[3] , _u0_ch6_am0[2] , _u0_ch6_am0[1] ,_u0_ch6_am0[0] , _u0_ch6_am1[31] , _u0_ch6_am1[30] , _u0_ch6_am1[29] ,_u0_ch6_am1[28] , _u0_ch6_am1[27] , _u0_ch6_am1[26] ,_u0_ch6_am1[25] , _u0_ch6_am1[24] , _u0_ch6_am1[23] ,_u0_ch6_am1[22] , _u0_ch6_am1[21] , _u0_ch6_am1[20] ,_u0_ch6_am1[19] , _u0_ch6_am1[18] , _u0_ch6_am1[17] ,_u0_ch6_am1[16] , _u0_ch6_am1[15] , _u0_ch6_am1[14] ,_u0_ch6_am1[13] , _u0_ch6_am1[12] , _u0_ch6_am1[11] ,_u0_ch6_am1[10] , _u0_ch6_am1[9] , _u0_ch6_am1[8] , _u0_ch6_am1[7] ,_u0_ch6_am1[6] , _u0_ch6_am1[5] , _u0_ch6_am1[4] , _u0_ch6_am1[3] ,_u0_ch6_am1[2] , _u0_ch6_am1[1] , _u0_ch6_am1[0] , _u0_pointer7[31] ,_u0_pointer7[30] , _u0_pointer7[29] , _u0_pointer7[28] ,_u0_pointer7[27] , _u0_pointer7[26] , _u0_pointer7[25] ,_u0_pointer7[24] , _u0_pointer7[23] , _u0_pointer7[22] ,_u0_pointer7[21] , _u0_pointer7[20] , _u0_pointer7[19] ,_u0_pointer7[18] , _u0_pointer7[17] , _u0_pointer7[16] ,_u0_pointer7[15] , _u0_pointer7[14] , _u0_pointer7[13] ,_u0_pointer7[12] , _u0_pointer7[11] , _u0_pointer7[10] ,_u0_pointer7[9] , _u0_pointer7[8] , _u0_pointer7[7] ,_u0_pointer7[6] , _u0_pointer7[5] , _u0_pointer7[4] ,_u0_pointer7[3] , _u0_pointer7[2] , _u0_pointer7[1] ,_u0_pointer7[0] , _u0_pointer7_s[31] , _u0_pointer7_s[30] ,_u0_pointer7_s[29] , _u0_pointer7_s[28] , _u0_pointer7_s[27] ,_u0_pointer7_s[26] , _u0_pointer7_s[25] , _u0_pointer7_s[24] ,_u0_pointer7_s[23] , _u0_pointer7_s[22] , _u0_pointer7_s[21] ,_u0_pointer7_s[20] , _u0_pointer7_s[19] , _u0_pointer7_s[18] ,_u0_pointer7_s[17] , _u0_pointer7_s[16] , _u0_pointer7_s[15] ,_u0_pointer7_s[14] , _u0_pointer7_s[13] , _u0_pointer7_s[12] ,_u0_pointer7_s[11] , _u0_pointer7_s[10] , _u0_pointer7_s[9] ,_u0_pointer7_s[8] , _u0_pointer7_s[7] , _u0_pointer7_s[6] ,_u0_pointer7_s[5] , _u0_pointer7_s[4] , _u0_pointer7_s[3] ,_u0_pointer7_s[2] , _u0_pointer7_s[1] , _u0_pointer7_s[0] ,_u0_ch7_csr[31] , _u0_ch7_csr[30] , _u0_ch7_csr[29] ,_u0_ch7_csr[28] , _u0_ch7_csr[27] , _u0_ch7_csr[26] ,_u0_ch7_csr[25] , _u0_ch7_csr[24] , _u0_ch7_csr[23] ,_u0_ch7_csr[22] , _u0_ch7_csr[21] , _u0_ch7_csr[20] ,_u0_ch7_csr[19] , _u0_ch7_csr[18] , _u0_ch7_csr[17] ,_u0_ch7_csr[16] , _u0_ch7_csr[15] , _u0_ch7_csr[14] ,_u0_ch7_csr[13] , _u0_ch7_csr[12] , _u0_ch7_csr[11] ,_u0_ch7_csr[10] , _u0_ch7_csr[9] , _u0_ch7_csr[8] , _u0_ch7_csr[7] ,_u0_ch7_csr[6] , _u0_ch7_csr[5] , _u0_ch7_csr[4] , _u0_ch7_csr[3] ,_u0_ch7_csr[2] , _u0_ch7_csr[1] , _u0_ch7_csr[0] , _u0_ch7_txsz[31] ,_u0_ch7_txsz[30] , _u0_ch7_txsz[29] , _u0_ch7_txsz[28] ,_u0_ch7_txsz[27] , _u0_ch7_txsz[26] , _u0_ch7_txsz[25] ,_u0_ch7_txsz[24] , _u0_ch7_txsz[23] , _u0_ch7_txsz[22] ,_u0_ch7_txsz[21] , _u0_ch7_txsz[20] , _u0_ch7_txsz[19] ,_u0_ch7_txsz[18] , _u0_ch7_txsz[17] , _u0_ch7_txsz[16] ,_u0_ch7_txsz[15] , _u0_ch7_txsz[14] , _u0_ch7_txsz[13] ,_u0_ch7_txsz[12] , _u0_ch7_txsz[11] , _u0_ch7_txsz[10] ,_u0_ch7_txsz[9] , _u0_ch7_txsz[8] , _u0_ch7_txsz[7] ,_u0_ch7_txsz[6] , _u0_ch7_txsz[5] , _u0_ch7_txsz[4] ,_u0_ch7_txsz[3] , _u0_ch7_txsz[2] , _u0_ch7_txsz[1] ,_u0_ch7_txsz[0] , _u0_ch7_adr0[31] , _u0_ch7_adr0[30] ,_u0_ch7_adr0[29] , _u0_ch7_adr0[28] , _u0_ch7_adr0[27] ,_u0_ch7_adr0[26] , _u0_ch7_adr0[25] , _u0_ch7_adr0[24] ,_u0_ch7_adr0[23] , _u0_ch7_adr0[22] , _u0_ch7_adr0[21] ,_u0_ch7_adr0[20] , _u0_ch7_adr0[19] , _u0_ch7_adr0[18] ,_u0_ch7_adr0[17] , _u0_ch7_adr0[16] , _u0_ch7_adr0[15] ,_u0_ch7_adr0[14] , _u0_ch7_adr0[13] , _u0_ch7_adr0[12] ,_u0_ch7_adr0[11] , _u0_ch7_adr0[10] , _u0_ch7_adr0[9] ,_u0_ch7_adr0[8] , _u0_ch7_adr0[7] , _u0_ch7_adr0[6] ,_u0_ch7_adr0[5] , _u0_ch7_adr0[4] , _u0_ch7_adr0[3] ,_u0_ch7_adr0[2] , _u0_ch7_adr0[1] , _u0_ch7_adr0[0] ,_u0_ch7_adr1[31] , _u0_ch7_adr1[30] , _u0_ch7_adr1[29] ,_u0_ch7_adr1[28] , _u0_ch7_adr1[27] , _u0_ch7_adr1[26] ,_u0_ch7_adr1[25] , _u0_ch7_adr1[24] , _u0_ch7_adr1[23] ,_u0_ch7_adr1[22] , _u0_ch7_adr1[21] , _u0_ch7_adr1[20] ,_u0_ch7_adr1[19] , _u0_ch7_adr1[18] , _u0_ch7_adr1[17] ,_u0_ch7_adr1[16] , _u0_ch7_adr1[15] , _u0_ch7_adr1[14] ,_u0_ch7_adr1[13] , _u0_ch7_adr1[12] , _u0_ch7_adr1[11] ,_u0_ch7_adr1[10] , _u0_ch7_adr1[9] , _u0_ch7_adr1[8] ,_u0_ch7_adr1[7] , _u0_ch7_adr1[6] , _u0_ch7_adr1[5] ,_u0_ch7_adr1[4] , _u0_ch7_adr1[3] , _u0_ch7_adr1[2] ,_u0_ch7_adr1[1] , _u0_ch7_adr1[0] , _u0_ch7_am0[31] ,_u0_ch7_am0[30] , _u0_ch7_am0[29] , _u0_ch7_am0[28] ,_u0_ch7_am0[27] , _u0_ch7_am0[26] , _u0_ch7_am0[25] ,_u0_ch7_am0[24] , _u0_ch7_am0[23] , _u0_ch7_am0[22] ,_u0_ch7_am0[21] , _u0_ch7_am0[20] , _u0_ch7_am0[19] ,_u0_ch7_am0[18] , _u0_ch7_am0[17] , _u0_ch7_am0[16] ,_u0_ch7_am0[15] , _u0_ch7_am0[14] , _u0_ch7_am0[13] ,_u0_ch7_am0[12] , _u0_ch7_am0[11] , _u0_ch7_am0[10] , _u0_ch7_am0[9] ,_u0_ch7_am0[8] , _u0_ch7_am0[7] , _u0_ch7_am0[6] , _u0_ch7_am0[5] ,_u0_ch7_am0[4] , _u0_ch7_am0[3] , _u0_ch7_am0[2] , _u0_ch7_am0[1] ,_u0_ch7_am0[0] , _u0_ch7_am1[31] , _u0_ch7_am1[30] , _u0_ch7_am1[29] ,_u0_ch7_am1[28] , _u0_ch7_am1[27] , _u0_ch7_am1[26] ,_u0_ch7_am1[25] , _u0_ch7_am1[24] , _u0_ch7_am1[23] ,_u0_ch7_am1[22] , _u0_ch7_am1[21] , _u0_ch7_am1[20] ,_u0_ch7_am1[19] , _u0_ch7_am1[18] , _u0_ch7_am1[17] ,_u0_ch7_am1[16] , _u0_ch7_am1[15] , _u0_ch7_am1[14] ,_u0_ch7_am1[13] , _u0_ch7_am1[12] , _u0_ch7_am1[11] ,_u0_ch7_am1[10] , _u0_ch7_am1[9] , _u0_ch7_am1[8] , _u0_ch7_am1[7] ,_u0_ch7_am1[6] , _u0_ch7_am1[5] , _u0_ch7_am1[4] , _u0_ch7_am1[3] ,_u0_ch7_am1[2] , _u0_ch7_am1[1] , _u0_ch7_am1[0] , _u0_pointer8[31] ,_u0_pointer8[30] , _u0_pointer8[29] , _u0_pointer8[28] ,_u0_pointer8[27] , _u0_pointer8[26] , _u0_pointer8[25] ,_u0_pointer8[24] , _u0_pointer8[23] , _u0_pointer8[22] ,_u0_pointer8[21] , _u0_pointer8[20] , _u0_pointer8[19] ,_u0_pointer8[18] , _u0_pointer8[17] , _u0_pointer8[16] ,_u0_pointer8[15] , _u0_pointer8[14] , _u0_pointer8[13] ,_u0_pointer8[12] , _u0_pointer8[11] , _u0_pointer8[10] ,_u0_pointer8[9] , _u0_pointer8[8] , _u0_pointer8[7] ,_u0_pointer8[6] , _u0_pointer8[5] , _u0_pointer8[4] ,_u0_pointer8[3] , _u0_pointer8[2] , _u0_pointer8[1] ,_u0_pointer8[0] , _u0_pointer8_s[31] , _u0_pointer8_s[30] ,_u0_pointer8_s[29] , _u0_pointer8_s[28] , _u0_pointer8_s[27] ,_u0_pointer8_s[26] , _u0_pointer8_s[25] , _u0_pointer8_s[24] ,_u0_pointer8_s[23] , _u0_pointer8_s[22] , _u0_pointer8_s[21] ,_u0_pointer8_s[20] , _u0_pointer8_s[19] , _u0_pointer8_s[18] ,_u0_pointer8_s[17] , _u0_pointer8_s[16] , _u0_pointer8_s[15] ,_u0_pointer8_s[14] , _u0_pointer8_s[13] , _u0_pointer8_s[12] ,_u0_pointer8_s[11] , _u0_pointer8_s[10] , _u0_pointer8_s[9] ,_u0_pointer8_s[8] , _u0_pointer8_s[7] , _u0_pointer8_s[6] ,_u0_pointer8_s[5] , _u0_pointer8_s[4] , _u0_pointer8_s[3] ,_u0_pointer8_s[2] , _u0_pointer8_s[1] , _u0_pointer8_s[0] ,_u0_ch8_csr[31] , _u0_ch8_csr[30] , _u0_ch8_csr[29] ,_u0_ch8_csr[28] , _u0_ch8_csr[27] , _u0_ch8_csr[26] ,_u0_ch8_csr[25] , _u0_ch8_csr[24] , _u0_ch8_csr[23] ,_u0_ch8_csr[22] , _u0_ch8_csr[21] , _u0_ch8_csr[20] ,_u0_ch8_csr[19] , _u0_ch8_csr[18] , _u0_ch8_csr[17] ,_u0_ch8_csr[16] , _u0_ch8_csr[15] , _u0_ch8_csr[14] ,_u0_ch8_csr[13] , _u0_ch8_csr[12] , _u0_ch8_csr[11] ,_u0_ch8_csr[10] , _u0_ch8_csr[9] , _u0_ch8_csr[8] , _u0_ch8_csr[7] ,_u0_ch8_csr[6] , _u0_ch8_csr[5] , _u0_ch8_csr[4] , _u0_ch8_csr[3] ,_u0_ch8_csr[2] , _u0_ch8_csr[1] , _u0_ch8_csr[0] , _u0_ch8_txsz[31] ,_u0_ch8_txsz[30] , _u0_ch8_txsz[29] , _u0_ch8_txsz[28] ,_u0_ch8_txsz[27] , _u0_ch8_txsz[26] , _u0_ch8_txsz[25] ,_u0_ch8_txsz[24] , _u0_ch8_txsz[23] , _u0_ch8_txsz[22] ,_u0_ch8_txsz[21] , _u0_ch8_txsz[20] , _u0_ch8_txsz[19] ,_u0_ch8_txsz[18] , _u0_ch8_txsz[17] , _u0_ch8_txsz[16] ,_u0_ch8_txsz[15] , _u0_ch8_txsz[14] , _u0_ch8_txsz[13] ,_u0_ch8_txsz[12] , _u0_ch8_txsz[11] , _u0_ch8_txsz[10] ,_u0_ch8_txsz[9] , _u0_ch8_txsz[8] , _u0_ch8_txsz[7] ,_u0_ch8_txsz[6] , _u0_ch8_txsz[5] , _u0_ch8_txsz[4] ,_u0_ch8_txsz[3] , _u0_ch8_txsz[2] , _u0_ch8_txsz[1] ,_u0_ch8_txsz[0] , _u0_ch8_adr0[31] , _u0_ch8_adr0[30] ,_u0_ch8_adr0[29] , _u0_ch8_adr0[28] , _u0_ch8_adr0[27] ,_u0_ch8_adr0[26] , _u0_ch8_adr0[25] , _u0_ch8_adr0[24] ,_u0_ch8_adr0[23] , _u0_ch8_adr0[22] , _u0_ch8_adr0[21] ,_u0_ch8_adr0[20] , _u0_ch8_adr0[19] , _u0_ch8_adr0[18] ,_u0_ch8_adr0[17] , _u0_ch8_adr0[16] , _u0_ch8_adr0[15] ,_u0_ch8_adr0[14] , _u0_ch8_adr0[13] , _u0_ch8_adr0[12] ,_u0_ch8_adr0[11] , _u0_ch8_adr0[10] , _u0_ch8_adr0[9] ,_u0_ch8_adr0[8] , _u0_ch8_adr0[7] , _u0_ch8_adr0[6] ,_u0_ch8_adr0[5] , _u0_ch8_adr0[4] , _u0_ch8_adr0[3] ,_u0_ch8_adr0[2] , _u0_ch8_adr0[1] , _u0_ch8_adr0[0] ,_u0_ch8_adr1[31] , _u0_ch8_adr1[30] , _u0_ch8_adr1[29] ,_u0_ch8_adr1[28] , _u0_ch8_adr1[27] , _u0_ch8_adr1[26] ,_u0_ch8_adr1[25] , _u0_ch8_adr1[24] , _u0_ch8_adr1[23] ,_u0_ch8_adr1[22] , _u0_ch8_adr1[21] , _u0_ch8_adr1[20] ,_u0_ch8_adr1[19] , _u0_ch8_adr1[18] , _u0_ch8_adr1[17] ,_u0_ch8_adr1[16] , _u0_ch8_adr1[15] , _u0_ch8_adr1[14] ,_u0_ch8_adr1[13] , _u0_ch8_adr1[12] , _u0_ch8_adr1[11] ,_u0_ch8_adr1[10] , _u0_ch8_adr1[9] , _u0_ch8_adr1[8] ,_u0_ch8_adr1[7] , _u0_ch8_adr1[6] , _u0_ch8_adr1[5] ,_u0_ch8_adr1[4] , _u0_ch8_adr1[3] , _u0_ch8_adr1[2] ,_u0_ch8_adr1[1] , _u0_ch8_adr1[0] , _u0_ch8_am0[31] ,_u0_ch8_am0[30] , _u0_ch8_am0[29] , _u0_ch8_am0[28] ,_u0_ch8_am0[27] , _u0_ch8_am0[26] , _u0_ch8_am0[25] ,_u0_ch8_am0[24] , _u0_ch8_am0[23] , _u0_ch8_am0[22] ,_u0_ch8_am0[21] , _u0_ch8_am0[20] , _u0_ch8_am0[19] ,_u0_ch8_am0[18] , _u0_ch8_am0[17] , _u0_ch8_am0[16] ,_u0_ch8_am0[15] , _u0_ch8_am0[14] , _u0_ch8_am0[13] ,_u0_ch8_am0[12] , _u0_ch8_am0[11] , _u0_ch8_am0[10] , _u0_ch8_am0[9] ,_u0_ch8_am0[8] , _u0_ch8_am0[7] , _u0_ch8_am0[6] , _u0_ch8_am0[5] ,_u0_ch8_am0[4] , _u0_ch8_am0[3] , _u0_ch8_am0[2] , _u0_ch8_am0[1] ,_u0_ch8_am0[0] , _u0_ch8_am1[31] , _u0_ch8_am1[30] , _u0_ch8_am1[29] ,_u0_ch8_am1[28] , _u0_ch8_am1[27] , _u0_ch8_am1[26] ,_u0_ch8_am1[25] , _u0_ch8_am1[24] , _u0_ch8_am1[23] ,_u0_ch8_am1[22] , _u0_ch8_am1[21] , _u0_ch8_am1[20] ,_u0_ch8_am1[19] , _u0_ch8_am1[18] , _u0_ch8_am1[17] ,_u0_ch8_am1[16] , _u0_ch8_am1[15] , _u0_ch8_am1[14] ,_u0_ch8_am1[13] , _u0_ch8_am1[12] , _u0_ch8_am1[11] ,_u0_ch8_am1[10] , _u0_ch8_am1[9] , _u0_ch8_am1[8] , _u0_ch8_am1[7] ,_u0_ch8_am1[6] , _u0_ch8_am1[5] , _u0_ch8_am1[4] , _u0_ch8_am1[3] ,_u0_ch8_am1[2] , _u0_ch8_am1[1] , _u0_ch8_am1[0] , _u0_pointer9[31] ,_u0_pointer9[30] , _u0_pointer9[29] , _u0_pointer9[28] ,_u0_pointer9[27] , _u0_pointer9[26] , _u0_pointer9[25] ,_u0_pointer9[24] , _u0_pointer9[23] , _u0_pointer9[22] ,_u0_pointer9[21] , _u0_pointer9[20] , _u0_pointer9[19] ,_u0_pointer9[18] , _u0_pointer9[17] , _u0_pointer9[16] ,_u0_pointer9[15] , _u0_pointer9[14] , _u0_pointer9[13] ,_u0_pointer9[12] , _u0_pointer9[11] , _u0_pointer9[10] ,_u0_pointer9[9] , _u0_pointer9[8] , _u0_pointer9[7] ,_u0_pointer9[6] , _u0_pointer9[5] , _u0_pointer9[4] ,_u0_pointer9[3] , _u0_pointer9[2] , _u0_pointer9[1] ,_u0_pointer9[0] , _u0_pointer9_s[31] , _u0_pointer9_s[30] ,_u0_pointer9_s[29] , _u0_pointer9_s[28] , _u0_pointer9_s[27] ,_u0_pointer9_s[26] , _u0_pointer9_s[25] , _u0_pointer9_s[24] ,_u0_pointer9_s[23] , _u0_pointer9_s[22] , _u0_pointer9_s[21] ,_u0_pointer9_s[20] , _u0_pointer9_s[19] , _u0_pointer9_s[18] ,_u0_pointer9_s[17] , _u0_pointer9_s[16] , _u0_pointer9_s[15] ,_u0_pointer9_s[14] , _u0_pointer9_s[13] , _u0_pointer9_s[12] ,_u0_pointer9_s[11] , _u0_pointer9_s[10] , _u0_pointer9_s[9] ,_u0_pointer9_s[8] , _u0_pointer9_s[7] , _u0_pointer9_s[6] ,_u0_pointer9_s[5] , _u0_pointer9_s[4] , _u0_pointer9_s[3] ,_u0_pointer9_s[2] , _u0_pointer9_s[1] , _u0_pointer9_s[0] ,_u0_ch9_csr[31] , _u0_ch9_csr[30] , _u0_ch9_csr[29] ,_u0_ch9_csr[28] , _u0_ch9_csr[27] , _u0_ch9_csr[26] ,_u0_ch9_csr[25] , _u0_ch9_csr[24] , _u0_ch9_csr[23] ,_u0_ch9_csr[22] , _u0_ch9_csr[21] , _u0_ch9_csr[20] ,_u0_ch9_csr[19] , _u0_ch9_csr[18] , _u0_ch9_csr[17] ,_u0_ch9_csr[16] , _u0_ch9_csr[15] , _u0_ch9_csr[14] ,_u0_ch9_csr[13] , _u0_ch9_csr[12] , _u0_ch9_csr[11] ,_u0_ch9_csr[10] , _u0_ch9_csr[9] , _u0_ch9_csr[8] , _u0_ch9_csr[7] ,_u0_ch9_csr[6] , _u0_ch9_csr[5] , _u0_ch9_csr[4] , _u0_ch9_csr[3] ,_u0_ch9_csr[2] , _u0_ch9_csr[1] , _u0_ch9_csr[0] , _u0_ch9_txsz[31] ,_u0_ch9_txsz[30] , _u0_ch9_txsz[29] , _u0_ch9_txsz[28] ,_u0_ch9_txsz[27] , _u0_ch9_txsz[26] , _u0_ch9_txsz[25] ,_u0_ch9_txsz[24] , _u0_ch9_txsz[23] , _u0_ch9_txsz[22] ,_u0_ch9_txsz[21] , _u0_ch9_txsz[20] , _u0_ch9_txsz[19] ,_u0_ch9_txsz[18] , _u0_ch9_txsz[17] , _u0_ch9_txsz[16] ,_u0_ch9_txsz[15] , _u0_ch9_txsz[14] , _u0_ch9_txsz[13] ,_u0_ch9_txsz[12] , _u0_ch9_txsz[11] , _u0_ch9_txsz[10] ,_u0_ch9_txsz[9] , _u0_ch9_txsz[8] , _u0_ch9_txsz[7] ,_u0_ch9_txsz[6] , _u0_ch9_txsz[5] , _u0_ch9_txsz[4] ,_u0_ch9_txsz[3] , _u0_ch9_txsz[2] , _u0_ch9_txsz[1] ,_u0_ch9_txsz[0] , _u0_ch9_adr0[31] , _u0_ch9_adr0[30] ,_u0_ch9_adr0[29] , _u0_ch9_adr0[28] , _u0_ch9_adr0[27] ,_u0_ch9_adr0[26] , _u0_ch9_adr0[25] , _u0_ch9_adr0[24] ,_u0_ch9_adr0[23] , _u0_ch9_adr0[22] , _u0_ch9_adr0[21] ,_u0_ch9_adr0[20] , _u0_ch9_adr0[19] , _u0_ch9_adr0[18] ,_u0_ch9_adr0[17] , _u0_ch9_adr0[16] , _u0_ch9_adr0[15] ,_u0_ch9_adr0[14] , _u0_ch9_adr0[13] , _u0_ch9_adr0[12] ,_u0_ch9_adr0[11] , _u0_ch9_adr0[10] , _u0_ch9_adr0[9] ,_u0_ch9_adr0[8] , _u0_ch9_adr0[7] , _u0_ch9_adr0[6] ,_u0_ch9_adr0[5] , _u0_ch9_adr0[4] , _u0_ch9_adr0[3] ,_u0_ch9_adr0[2] , _u0_ch9_adr0[1] , _u0_ch9_adr0[0] ,_u0_ch9_adr1[31] , _u0_ch9_adr1[30] , _u0_ch9_adr1[29] ,_u0_ch9_adr1[28] , _u0_ch9_adr1[27] , _u0_ch9_adr1[26] ,_u0_ch9_adr1[25] , _u0_ch9_adr1[24] , _u0_ch9_adr1[23] ,_u0_ch9_adr1[22] , _u0_ch9_adr1[21] , _u0_ch9_adr1[20] ,_u0_ch9_adr1[19] , _u0_ch9_adr1[18] , _u0_ch9_adr1[17] ,_u0_ch9_adr1[16] , _u0_ch9_adr1[15] , _u0_ch9_adr1[14] ,_u0_ch9_adr1[13] , _u0_ch9_adr1[12] , _u0_ch9_adr1[11] ,_u0_ch9_adr1[10] , _u0_ch9_adr1[9] , _u0_ch9_adr1[8] ,_u0_ch9_adr1[7] , _u0_ch9_adr1[6] , _u0_ch9_adr1[5] ,_u0_ch9_adr1[4] , _u0_ch9_adr1[3] , _u0_ch9_adr1[2] ,_u0_ch9_adr1[1] , _u0_ch9_adr1[0] , _u0_ch9_am0[31] ,_u0_ch9_am0[30] , _u0_ch9_am0[29] , _u0_ch9_am0[28] ,_u0_ch9_am0[27] , _u0_ch9_am0[26] , _u0_ch9_am0[25] ,_u0_ch9_am0[24] , _u0_ch9_am0[23] , _u0_ch9_am0[22] ,_u0_ch9_am0[21] , _u0_ch9_am0[20] , _u0_ch9_am0[19] ,_u0_ch9_am0[18] , _u0_ch9_am0[17] , _u0_ch9_am0[16] ,_u0_ch9_am0[15] , _u0_ch9_am0[14] , _u0_ch9_am0[13] ,_u0_ch9_am0[12] , _u0_ch9_am0[11] , _u0_ch9_am0[10] , _u0_ch9_am0[9] ,_u0_ch9_am0[8] , _u0_ch9_am0[7] , _u0_ch9_am0[6] , _u0_ch9_am0[5] ,_u0_ch9_am0[4] , _u0_ch9_am0[3] , _u0_ch9_am0[2] , _u0_ch9_am0[1] ,_u0_ch9_am0[0] , _u0_ch9_am1[31] , _u0_ch9_am1[30] , _u0_ch9_am1[29] ,_u0_ch9_am1[28] , _u0_ch9_am1[27] , _u0_ch9_am1[26] ,_u0_ch9_am1[25] , _u0_ch9_am1[24] , _u0_ch9_am1[23] ,_u0_ch9_am1[22] , _u0_ch9_am1[21] , _u0_ch9_am1[20] ,_u0_ch9_am1[19] , _u0_ch9_am1[18] , _u0_ch9_am1[17] ,_u0_ch9_am1[16] , _u0_ch9_am1[15] , _u0_ch9_am1[14] ,_u0_ch9_am1[13] , _u0_ch9_am1[12] , _u0_ch9_am1[11] ,_u0_ch9_am1[10] , _u0_ch9_am1[9] , _u0_ch9_am1[8] , _u0_ch9_am1[7] ,_u0_ch9_am1[6] , _u0_ch9_am1[5] , _u0_ch9_am1[4] , _u0_ch9_am1[3] ,_u0_ch9_am1[2] , _u0_ch9_am1[1] , _u0_ch9_am1[0] , _u0_pointer10[31] ,_u0_pointer10[30] , _u0_pointer10[29] , _u0_pointer10[28] ,_u0_pointer10[27] , _u0_pointer10[26] , _u0_pointer10[25] ,_u0_pointer10[24] , _u0_pointer10[23] , _u0_pointer10[22] ,_u0_pointer10[21] , _u0_pointer10[20] , _u0_pointer10[19] ,_u0_pointer10[18] , _u0_pointer10[17] , _u0_pointer10[16] ,_u0_pointer10[15] , _u0_pointer10[14] , _u0_pointer10[13] ,_u0_pointer10[12] , _u0_pointer10[11] , _u0_pointer10[10] ,_u0_pointer10[9] , _u0_pointer10[8] , _u0_pointer10[7] ,_u0_pointer10[6] , _u0_pointer10[5] , _u0_pointer10[4] ,_u0_pointer10[3] , _u0_pointer10[2] , _u0_pointer10[1] ,_u0_pointer10[0] , _u0_pointer10_s[31] , _u0_pointer10_s[30] ,_u0_pointer10_s[29] , _u0_pointer10_s[28] , _u0_pointer10_s[27] ,_u0_pointer10_s[26] , _u0_pointer10_s[25] , _u0_pointer10_s[24] ,_u0_pointer10_s[23] , _u0_pointer10_s[22] , _u0_pointer10_s[21] ,_u0_pointer10_s[20] , _u0_pointer10_s[19] , _u0_pointer10_s[18] ,_u0_pointer10_s[17] , _u0_pointer10_s[16] , _u0_pointer10_s[15] ,_u0_pointer10_s[14] , _u0_pointer10_s[13] , _u0_pointer10_s[12] ,_u0_pointer10_s[11] , _u0_pointer10_s[10] , _u0_pointer10_s[9] ,_u0_pointer10_s[8] , _u0_pointer10_s[7] , _u0_pointer10_s[6] ,_u0_pointer10_s[5] , _u0_pointer10_s[4] , _u0_pointer10_s[3] ,_u0_pointer10_s[2] , _u0_pointer10_s[1] , _u0_pointer10_s[0] ,_u0_ch10_csr[31] , _u0_ch10_csr[30] , _u0_ch10_csr[29] ,_u0_ch10_csr[28] , _u0_ch10_csr[27] , _u0_ch10_csr[26] ,_u0_ch10_csr[25] , _u0_ch10_csr[24] , _u0_ch10_csr[23] ,_u0_ch10_csr[22] , _u0_ch10_csr[21] , _u0_ch10_csr[20] ,_u0_ch10_csr[19] , _u0_ch10_csr[18] , _u0_ch10_csr[17] ,_u0_ch10_csr[16] , _u0_ch10_csr[15] , _u0_ch10_csr[14] ,_u0_ch10_csr[13] , _u0_ch10_csr[12] , _u0_ch10_csr[11] ,_u0_ch10_csr[10] , _u0_ch10_csr[9] , _u0_ch10_csr[8] ,_u0_ch10_csr[7] , _u0_ch10_csr[6] , _u0_ch10_csr[5] ,_u0_ch10_csr[4] , _u0_ch10_csr[3] , _u0_ch10_csr[2] ,_u0_ch10_csr[1] , _u0_ch10_csr[0] , _u0_ch10_txsz[31] ,_u0_ch10_txsz[30] , _u0_ch10_txsz[29] , _u0_ch10_txsz[28] ,_u0_ch10_txsz[27] , _u0_ch10_txsz[26] , _u0_ch10_txsz[25] ,_u0_ch10_txsz[24] , _u0_ch10_txsz[23] , _u0_ch10_txsz[22] ,_u0_ch10_txsz[21] , _u0_ch10_txsz[20] , _u0_ch10_txsz[19] ,_u0_ch10_txsz[18] , _u0_ch10_txsz[17] , _u0_ch10_txsz[16] ,_u0_ch10_txsz[15] , _u0_ch10_txsz[14] , _u0_ch10_txsz[13] ,_u0_ch10_txsz[12] , _u0_ch10_txsz[11] , _u0_ch10_txsz[10] ,_u0_ch10_txsz[9] , _u0_ch10_txsz[8] , _u0_ch10_txsz[7] ,_u0_ch10_txsz[6] , _u0_ch10_txsz[5] , _u0_ch10_txsz[4] ,_u0_ch10_txsz[3] , _u0_ch10_txsz[2] , _u0_ch10_txsz[1] ,_u0_ch10_txsz[0] , _u0_ch10_adr0[31] , _u0_ch10_adr0[30] ,_u0_ch10_adr0[29] , _u0_ch10_adr0[28] , _u0_ch10_adr0[27] ,_u0_ch10_adr0[26] , _u0_ch10_adr0[25] , _u0_ch10_adr0[24] ,_u0_ch10_adr0[23] , _u0_ch10_adr0[22] , _u0_ch10_adr0[21] ,_u0_ch10_adr0[20] , _u0_ch10_adr0[19] , _u0_ch10_adr0[18] ,_u0_ch10_adr0[17] , _u0_ch10_adr0[16] , _u0_ch10_adr0[15] ,_u0_ch10_adr0[14] , _u0_ch10_adr0[13] , _u0_ch10_adr0[12] ,_u0_ch10_adr0[11] , _u0_ch10_adr0[10] , _u0_ch10_adr0[9] ,_u0_ch10_adr0[8] , _u0_ch10_adr0[7] , _u0_ch10_adr0[6] ,_u0_ch10_adr0[5] , _u0_ch10_adr0[4] , _u0_ch10_adr0[3] ,_u0_ch10_adr0[2] , _u0_ch10_adr0[1] , _u0_ch10_adr0[0] ,_u0_ch10_adr1[31] , _u0_ch10_adr1[30] , _u0_ch10_adr1[29] ,_u0_ch10_adr1[28] , _u0_ch10_adr1[27] , _u0_ch10_adr1[26] ,_u0_ch10_adr1[25] , _u0_ch10_adr1[24] , _u0_ch10_adr1[23] ,_u0_ch10_adr1[22] , _u0_ch10_adr1[21] , _u0_ch10_adr1[20] ,_u0_ch10_adr1[19] , _u0_ch10_adr1[18] , _u0_ch10_adr1[17] ,_u0_ch10_adr1[16] , _u0_ch10_adr1[15] , _u0_ch10_adr1[14] ,_u0_ch10_adr1[13] , _u0_ch10_adr1[12] , _u0_ch10_adr1[11] ,_u0_ch10_adr1[10] , _u0_ch10_adr1[9] , _u0_ch10_adr1[8] ,_u0_ch10_adr1[7] , _u0_ch10_adr1[6] , _u0_ch10_adr1[5] ,_u0_ch10_adr1[4] , _u0_ch10_adr1[3] , _u0_ch10_adr1[2] ,_u0_ch10_adr1[1] , _u0_ch10_adr1[0] , _u0_ch10_am0[31] ,_u0_ch10_am0[30] , _u0_ch10_am0[29] , _u0_ch10_am0[28] ,_u0_ch10_am0[27] , _u0_ch10_am0[26] , _u0_ch10_am0[25] ,_u0_ch10_am0[24] , _u0_ch10_am0[23] , _u0_ch10_am0[22] ,_u0_ch10_am0[21] , _u0_ch10_am0[20] , _u0_ch10_am0[19] ,_u0_ch10_am0[18] , _u0_ch10_am0[17] , _u0_ch10_am0[16] ,_u0_ch10_am0[15] , _u0_ch10_am0[14] , _u0_ch10_am0[13] ,_u0_ch10_am0[12] , _u0_ch10_am0[11] , _u0_ch10_am0[10] ,_u0_ch10_am0[9] , _u0_ch10_am0[8] , _u0_ch10_am0[7] ,_u0_ch10_am0[6] , _u0_ch10_am0[5] , _u0_ch10_am0[4] ,_u0_ch10_am0[3] , _u0_ch10_am0[2] , _u0_ch10_am0[1] ,_u0_ch10_am0[0] , _u0_ch10_am1[31] , _u0_ch10_am1[30] ,_u0_ch10_am1[29] , _u0_ch10_am1[28] , _u0_ch10_am1[27] ,_u0_ch10_am1[26] , _u0_ch10_am1[25] , _u0_ch10_am1[24] ,_u0_ch10_am1[23] , _u0_ch10_am1[22] , _u0_ch10_am1[21] ,_u0_ch10_am1[20] , _u0_ch10_am1[19] , _u0_ch10_am1[18] ,_u0_ch10_am1[17] , _u0_ch10_am1[16] , _u0_ch10_am1[15] ,_u0_ch10_am1[14] , _u0_ch10_am1[13] , _u0_ch10_am1[12] ,_u0_ch10_am1[11] , _u0_ch10_am1[10] , _u0_ch10_am1[9] ,_u0_ch10_am1[8] , _u0_ch10_am1[7] , _u0_ch10_am1[6] ,_u0_ch10_am1[5] , _u0_ch10_am1[4] , _u0_ch10_am1[3] ,_u0_ch10_am1[2] , _u0_ch10_am1[1] , _u0_ch10_am1[0] ,_u0_pointer11[31] , _u0_pointer11[30] , _u0_pointer11[29] ,_u0_pointer11[28] , _u0_pointer11[27] , _u0_pointer11[26] ,_u0_pointer11[25] , _u0_pointer11[24] , _u0_pointer11[23] ,_u0_pointer11[22] , _u0_pointer11[21] , _u0_pointer11[20] ,_u0_pointer11[19] , _u0_pointer11[18] , _u0_pointer11[17] ,_u0_pointer11[16] , _u0_pointer11[15] , _u0_pointer11[14] ,_u0_pointer11[13] , _u0_pointer11[12] , _u0_pointer11[11] ,_u0_pointer11[10] , _u0_pointer11[9] , _u0_pointer11[8] ,_u0_pointer11[7] , _u0_pointer11[6] , _u0_pointer11[5] ,_u0_pointer11[4] , _u0_pointer11[3] , _u0_pointer11[2] ,_u0_pointer11[1] , _u0_pointer11[0] , _u0_pointer11_s[31] ,_u0_pointer11_s[30] , _u0_pointer11_s[29] , _u0_pointer11_s[28] ,_u0_pointer11_s[27] , _u0_pointer11_s[26] , _u0_pointer11_s[25] ,_u0_pointer11_s[24] , _u0_pointer11_s[23] , _u0_pointer11_s[22] ,_u0_pointer11_s[21] , _u0_pointer11_s[20] , _u0_pointer11_s[19] ,_u0_pointer11_s[18] , _u0_pointer11_s[17] , _u0_pointer11_s[16] ,_u0_pointer11_s[15] , _u0_pointer11_s[14] , _u0_pointer11_s[13] ,_u0_pointer11_s[12] , _u0_pointer11_s[11] , _u0_pointer11_s[10] ,_u0_pointer11_s[9] , _u0_pointer11_s[8] , _u0_pointer11_s[7] ,_u0_pointer11_s[6] , _u0_pointer11_s[5] , _u0_pointer11_s[4] ,_u0_pointer11_s[3] , _u0_pointer11_s[2] , _u0_pointer11_s[1] ,_u0_pointer11_s[0] , _u0_ch11_csr[31] , _u0_ch11_csr[30] ,_u0_ch11_csr[29] , _u0_ch11_csr[28] , _u0_ch11_csr[27] ,_u0_ch11_csr[26] , _u0_ch11_csr[25] , _u0_ch11_csr[24] ,_u0_ch11_csr[23] , _u0_ch11_csr[22] , _u0_ch11_csr[21] ,_u0_ch11_csr[20] , _u0_ch11_csr[19] , _u0_ch11_csr[18] ,_u0_ch11_csr[17] , _u0_ch11_csr[16] , _u0_ch11_csr[15] ,_u0_ch11_csr[14] , _u0_ch11_csr[13] , _u0_ch11_csr[12] ,_u0_ch11_csr[11] , _u0_ch11_csr[10] , _u0_ch11_csr[9] ,_u0_ch11_csr[8] , _u0_ch11_csr[7] , _u0_ch11_csr[6] ,_u0_ch11_csr[5] , _u0_ch11_csr[4] , _u0_ch11_csr[3] ,_u0_ch11_csr[2] , _u0_ch11_csr[1] , _u0_ch11_csr[0] ,_u0_ch11_txsz[31] , _u0_ch11_txsz[30] , _u0_ch11_txsz[29] ,_u0_ch11_txsz[28] , _u0_ch11_txsz[27] , _u0_ch11_txsz[26] ,_u0_ch11_txsz[25] , _u0_ch11_txsz[24] , _u0_ch11_txsz[23] ,_u0_ch11_txsz[22] , _u0_ch11_txsz[21] , _u0_ch11_txsz[20] ,_u0_ch11_txsz[19] , _u0_ch11_txsz[18] , _u0_ch11_txsz[17] ,_u0_ch11_txsz[16] , _u0_ch11_txsz[15] , _u0_ch11_txsz[14] ,_u0_ch11_txsz[13] , _u0_ch11_txsz[12] , _u0_ch11_txsz[11] ,_u0_ch11_txsz[10] , _u0_ch11_txsz[9] , _u0_ch11_txsz[8] ,_u0_ch11_txsz[7] , _u0_ch11_txsz[6] , _u0_ch11_txsz[5] ,_u0_ch11_txsz[4] , _u0_ch11_txsz[3] , _u0_ch11_txsz[2] ,_u0_ch11_txsz[1] , _u0_ch11_txsz[0] , _u0_ch11_adr0[31] ,_u0_ch11_adr0[30] , _u0_ch11_adr0[29] , _u0_ch11_adr0[28] ,_u0_ch11_adr0[27] , _u0_ch11_adr0[26] , _u0_ch11_adr0[25] ,_u0_ch11_adr0[24] , _u0_ch11_adr0[23] , _u0_ch11_adr0[22] ,_u0_ch11_adr0[21] , _u0_ch11_adr0[20] , _u0_ch11_adr0[19] ,_u0_ch11_adr0[18] , _u0_ch11_adr0[17] , _u0_ch11_adr0[16] ,_u0_ch11_adr0[15] , _u0_ch11_adr0[14] , _u0_ch11_adr0[13] ,_u0_ch11_adr0[12] , _u0_ch11_adr0[11] , _u0_ch11_adr0[10] ,_u0_ch11_adr0[9] , _u0_ch11_adr0[8] , _u0_ch11_adr0[7] ,_u0_ch11_adr0[6] , _u0_ch11_adr0[5] , _u0_ch11_adr0[4] ,_u0_ch11_adr0[3] , _u0_ch11_adr0[2] , _u0_ch11_adr0[1] ,_u0_ch11_adr0[0] , _u0_ch11_adr1[31] , _u0_ch11_adr1[30] ,_u0_ch11_adr1[29] , _u0_ch11_adr1[28] , _u0_ch11_adr1[27] ,_u0_ch11_adr1[26] , _u0_ch11_adr1[25] , _u0_ch11_adr1[24] ,_u0_ch11_adr1[23] , _u0_ch11_adr1[22] , _u0_ch11_adr1[21] ,_u0_ch11_adr1[20] , _u0_ch11_adr1[19] , _u0_ch11_adr1[18] ,_u0_ch11_adr1[17] , _u0_ch11_adr1[16] , _u0_ch11_adr1[15] ,_u0_ch11_adr1[14] , _u0_ch11_adr1[13] , _u0_ch11_adr1[12] ,_u0_ch11_adr1[11] , _u0_ch11_adr1[10] , _u0_ch11_adr1[9] ,_u0_ch11_adr1[8] , _u0_ch11_adr1[7] , _u0_ch11_adr1[6] ,_u0_ch11_adr1[5] , _u0_ch11_adr1[4] , _u0_ch11_adr1[3] ,_u0_ch11_adr1[2] , _u0_ch11_adr1[1] , _u0_ch11_adr1[0] ,_u0_ch11_am0[31] , _u0_ch11_am0[30] , _u0_ch11_am0[29] ,_u0_ch11_am0[28] , _u0_ch11_am0[27] , _u0_ch11_am0[26] ,_u0_ch11_am0[25] , _u0_ch11_am0[24] , _u0_ch11_am0[23] ,_u0_ch11_am0[22] , _u0_ch11_am0[21] , _u0_ch11_am0[20] ,_u0_ch11_am0[19] , _u0_ch11_am0[18] , _u0_ch11_am0[17] ,_u0_ch11_am0[16] , _u0_ch11_am0[15] , _u0_ch11_am0[14] ,_u0_ch11_am0[13] , _u0_ch11_am0[12] , _u0_ch11_am0[11] ,_u0_ch11_am0[10] , _u0_ch11_am0[9] , _u0_ch11_am0[8] ,_u0_ch11_am0[7] , _u0_ch11_am0[6] , _u0_ch11_am0[5] ,_u0_ch11_am0[4] , _u0_ch11_am0[3] , _u0_ch11_am0[2] ,_u0_ch11_am0[1] , _u0_ch11_am0[0] , _u0_ch11_am1[31] ,_u0_ch11_am1[30] , _u0_ch11_am1[29] , _u0_ch11_am1[28] ,_u0_ch11_am1[27] , _u0_ch11_am1[26] , _u0_ch11_am1[25] ,_u0_ch11_am1[24] , _u0_ch11_am1[23] , _u0_ch11_am1[22] ,_u0_ch11_am1[21] , _u0_ch11_am1[20] , _u0_ch11_am1[19] ,_u0_ch11_am1[18] , _u0_ch11_am1[17] , _u0_ch11_am1[16] ,_u0_ch11_am1[15] , _u0_ch11_am1[14] , _u0_ch11_am1[13] ,_u0_ch11_am1[12] , _u0_ch11_am1[11] , _u0_ch11_am1[10] ,_u0_ch11_am1[9] , _u0_ch11_am1[8] , _u0_ch11_am1[7] ,_u0_ch11_am1[6] , _u0_ch11_am1[5] , _u0_ch11_am1[4] ,_u0_ch11_am1[3] , _u0_ch11_am1[2] , _u0_ch11_am1[1] ,_u0_ch11_am1[0] , _u0_pointer12[31] , _u0_pointer12[30] ,_u0_pointer12[29] , _u0_pointer12[28] , _u0_pointer12[27] ,_u0_pointer12[26] , _u0_pointer12[25] , _u0_pointer12[24] ,_u0_pointer12[23] , _u0_pointer12[22] , _u0_pointer12[21] ,_u0_pointer12[20] , _u0_pointer12[19] , _u0_pointer12[18] ,_u0_pointer12[17] , _u0_pointer12[16] , _u0_pointer12[15] ,_u0_pointer12[14] , _u0_pointer12[13] , _u0_pointer12[12] ,_u0_pointer12[11] , _u0_pointer12[10] , _u0_pointer12[9] ,_u0_pointer12[8] , _u0_pointer12[7] , _u0_pointer12[6] ,_u0_pointer12[5] , _u0_pointer12[4] , _u0_pointer12[3] ,_u0_pointer12[2] , _u0_pointer12[1] , _u0_pointer12[0] ,_u0_pointer12_s[31] , _u0_pointer12_s[30] , _u0_pointer12_s[29] ,_u0_pointer12_s[28] , _u0_pointer12_s[27] , _u0_pointer12_s[26] ,_u0_pointer12_s[25] , _u0_pointer12_s[24] , _u0_pointer12_s[23] ,_u0_pointer12_s[22] , _u0_pointer12_s[21] , _u0_pointer12_s[20] ,_u0_pointer12_s[19] , _u0_pointer12_s[18] , _u0_pointer12_s[17] ,_u0_pointer12_s[16] , _u0_pointer12_s[15] , _u0_pointer12_s[14] ,_u0_pointer12_s[13] , _u0_pointer12_s[12] , _u0_pointer12_s[11] ,_u0_pointer12_s[10] , _u0_pointer12_s[9] , _u0_pointer12_s[8] ,_u0_pointer12_s[7] , _u0_pointer12_s[6] , _u0_pointer12_s[5] ,_u0_pointer12_s[4] , _u0_pointer12_s[3] , _u0_pointer12_s[2] ,_u0_pointer12_s[1] , _u0_pointer12_s[0] , _u0_ch12_csr[31] ,_u0_ch12_csr[30] , _u0_ch12_csr[29] , _u0_ch12_csr[28] ,_u0_ch12_csr[27] , _u0_ch12_csr[26] , _u0_ch12_csr[25] ,_u0_ch12_csr[24] , _u0_ch12_csr[23] , _u0_ch12_csr[22] ,_u0_ch12_csr[21] , _u0_ch12_csr[20] , _u0_ch12_csr[19] ,_u0_ch12_csr[18] , _u0_ch12_csr[17] , _u0_ch12_csr[16] ,_u0_ch12_csr[15] , _u0_ch12_csr[14] , _u0_ch12_csr[13] ,_u0_ch12_csr[12] , _u0_ch12_csr[11] , _u0_ch12_csr[10] ,_u0_ch12_csr[9] , _u0_ch12_csr[8] , _u0_ch12_csr[7] ,_u0_ch12_csr[6] , _u0_ch12_csr[5] , _u0_ch12_csr[4] ,_u0_ch12_csr[3] , _u0_ch12_csr[2] , _u0_ch12_csr[1] ,_u0_ch12_csr[0] , _u0_ch12_txsz[31] , _u0_ch12_txsz[30] ,_u0_ch12_txsz[29] , _u0_ch12_txsz[28] , _u0_ch12_txsz[27] ,_u0_ch12_txsz[26] , _u0_ch12_txsz[25] , _u0_ch12_txsz[24] ,_u0_ch12_txsz[23] , _u0_ch12_txsz[22] , _u0_ch12_txsz[21] ,_u0_ch12_txsz[20] , _u0_ch12_txsz[19] , _u0_ch12_txsz[18] ,_u0_ch12_txsz[17] , _u0_ch12_txsz[16] , _u0_ch12_txsz[15] ,_u0_ch12_txsz[14] , _u0_ch12_txsz[13] , _u0_ch12_txsz[12] ,_u0_ch12_txsz[11] , _u0_ch12_txsz[10] , _u0_ch12_txsz[9] ,_u0_ch12_txsz[8] , _u0_ch12_txsz[7] , _u0_ch12_txsz[6] ,_u0_ch12_txsz[5] , _u0_ch12_txsz[4] , _u0_ch12_txsz[3] ,_u0_ch12_txsz[2] , _u0_ch12_txsz[1] , _u0_ch12_txsz[0] ,_u0_ch12_adr0[31] , _u0_ch12_adr0[30] , _u0_ch12_adr0[29] ,_u0_ch12_adr0[28] , _u0_ch12_adr0[27] , _u0_ch12_adr0[26] ,_u0_ch12_adr0[25] , _u0_ch12_adr0[24] , _u0_ch12_adr0[23] ,_u0_ch12_adr0[22] , _u0_ch12_adr0[21] , _u0_ch12_adr0[20] ,_u0_ch12_adr0[19] , _u0_ch12_adr0[18] , _u0_ch12_adr0[17] ,_u0_ch12_adr0[16] , _u0_ch12_adr0[15] , _u0_ch12_adr0[14] ,_u0_ch12_adr0[13] , _u0_ch12_adr0[12] , _u0_ch12_adr0[11] ,_u0_ch12_adr0[10] , _u0_ch12_adr0[9] , _u0_ch12_adr0[8] ,_u0_ch12_adr0[7] , _u0_ch12_adr0[6] , _u0_ch12_adr0[5] ,_u0_ch12_adr0[4] , _u0_ch12_adr0[3] , _u0_ch12_adr0[2] ,_u0_ch12_adr0[1] , _u0_ch12_adr0[0] , _u0_ch12_adr1[31] ,_u0_ch12_adr1[30] , _u0_ch12_adr1[29] , _u0_ch12_adr1[28] ,_u0_ch12_adr1[27] , _u0_ch12_adr1[26] , _u0_ch12_adr1[25] ,_u0_ch12_adr1[24] , _u0_ch12_adr1[23] , _u0_ch12_adr1[22] ,_u0_ch12_adr1[21] , _u0_ch12_adr1[20] , _u0_ch12_adr1[19] ,_u0_ch12_adr1[18] , _u0_ch12_adr1[17] , _u0_ch12_adr1[16] ,_u0_ch12_adr1[15] , _u0_ch12_adr1[14] , _u0_ch12_adr1[13] ,_u0_ch12_adr1[12] , _u0_ch12_adr1[11] , _u0_ch12_adr1[10] ,_u0_ch12_adr1[9] , _u0_ch12_adr1[8] , _u0_ch12_adr1[7] ,_u0_ch12_adr1[6] , _u0_ch12_adr1[5] , _u0_ch12_adr1[4] ,_u0_ch12_adr1[3] , _u0_ch12_adr1[2] , _u0_ch12_adr1[1] ,_u0_ch12_adr1[0] , _u0_ch12_am0[31] , _u0_ch12_am0[30] ,_u0_ch12_am0[29] , _u0_ch12_am0[28] , _u0_ch12_am0[27] ,_u0_ch12_am0[26] , _u0_ch12_am0[25] , _u0_ch12_am0[24] ,_u0_ch12_am0[23] , _u0_ch12_am0[22] , _u0_ch12_am0[21] ,_u0_ch12_am0[20] , _u0_ch12_am0[19] , _u0_ch12_am0[18] ,_u0_ch12_am0[17] , _u0_ch12_am0[16] , _u0_ch12_am0[15] ,_u0_ch12_am0[14] , _u0_ch12_am0[13] , _u0_ch12_am0[12] ,_u0_ch12_am0[11] , _u0_ch12_am0[10] , _u0_ch12_am0[9] ,_u0_ch12_am0[8] , _u0_ch12_am0[7] , _u0_ch12_am0[6] ,_u0_ch12_am0[5] , _u0_ch12_am0[4] , _u0_ch12_am0[3] ,_u0_ch12_am0[2] , _u0_ch12_am0[1] , _u0_ch12_am0[0] ,_u0_ch12_am1[31] , _u0_ch12_am1[30] , _u0_ch12_am1[29] ,_u0_ch12_am1[28] , _u0_ch12_am1[27] , _u0_ch12_am1[26] ,_u0_ch12_am1[25] , _u0_ch12_am1[24] , _u0_ch12_am1[23] ,_u0_ch12_am1[22] , _u0_ch12_am1[21] , _u0_ch12_am1[20] ,_u0_ch12_am1[19] , _u0_ch12_am1[18] , _u0_ch12_am1[17] ,_u0_ch12_am1[16] , _u0_ch12_am1[15] , _u0_ch12_am1[14] ,_u0_ch12_am1[13] , _u0_ch12_am1[12] , _u0_ch12_am1[11] ,_u0_ch12_am1[10] , _u0_ch12_am1[9] , _u0_ch12_am1[8] ,_u0_ch12_am1[7] , _u0_ch12_am1[6] , _u0_ch12_am1[5] ,_u0_ch12_am1[4] , _u0_ch12_am1[3] , _u0_ch12_am1[2] ,_u0_ch12_am1[1] , _u0_ch12_am1[0] , _u0_pointer13[31] ,_u0_pointer13[30] , _u0_pointer13[29] , _u0_pointer13[28] ,_u0_pointer13[27] , _u0_pointer13[26] , _u0_pointer13[25] ,_u0_pointer13[24] , _u0_pointer13[23] , _u0_pointer13[22] ,_u0_pointer13[21] , _u0_pointer13[20] , _u0_pointer13[19] ,_u0_pointer13[18] , _u0_pointer13[17] , _u0_pointer13[16] ,_u0_pointer13[15] , _u0_pointer13[14] , _u0_pointer13[13] ,_u0_pointer13[12] , _u0_pointer13[11] , _u0_pointer13[10] ,_u0_pointer13[9] , _u0_pointer13[8] , _u0_pointer13[7] ,_u0_pointer13[6] , _u0_pointer13[5] , _u0_pointer13[4] ,_u0_pointer13[3] , _u0_pointer13[2] , _u0_pointer13[1] ,_u0_pointer13[0] , _u0_pointer13_s[31] , _u0_pointer13_s[30] ,_u0_pointer13_s[29] , _u0_pointer13_s[28] , _u0_pointer13_s[27] ,_u0_pointer13_s[26] , _u0_pointer13_s[25] , _u0_pointer13_s[24] ,_u0_pointer13_s[23] , _u0_pointer13_s[22] , _u0_pointer13_s[21] ,_u0_pointer13_s[20] , _u0_pointer13_s[19] , _u0_pointer13_s[18] ,_u0_pointer13_s[17] , _u0_pointer13_s[16] , _u0_pointer13_s[15] ,_u0_pointer13_s[14] , _u0_pointer13_s[13] , _u0_pointer13_s[12] ,_u0_pointer13_s[11] , _u0_pointer13_s[10] , _u0_pointer13_s[9] ,_u0_pointer13_s[8] , _u0_pointer13_s[7] , _u0_pointer13_s[6] ,_u0_pointer13_s[5] , _u0_pointer13_s[4] , _u0_pointer13_s[3] ,_u0_pointer13_s[2] , _u0_pointer13_s[1] , _u0_pointer13_s[0] ,_u0_ch13_csr[31] , _u0_ch13_csr[30] , _u0_ch13_csr[29] ,_u0_ch13_csr[28] , _u0_ch13_csr[27] , _u0_ch13_csr[26] ,_u0_ch13_csr[25] , _u0_ch13_csr[24] , _u0_ch13_csr[23] ,_u0_ch13_csr[22] , _u0_ch13_csr[21] , _u0_ch13_csr[20] ,_u0_ch13_csr[19] , _u0_ch13_csr[18] , _u0_ch13_csr[17] ,_u0_ch13_csr[16] , _u0_ch13_csr[15] , _u0_ch13_csr[14] ,_u0_ch13_csr[13] , _u0_ch13_csr[12] , _u0_ch13_csr[11] ,_u0_ch13_csr[10] , _u0_ch13_csr[9] , _u0_ch13_csr[8] ,_u0_ch13_csr[7] , _u0_ch13_csr[6] , _u0_ch13_csr[5] ,_u0_ch13_csr[4] , _u0_ch13_csr[3] , _u0_ch13_csr[2] ,_u0_ch13_csr[1] , _u0_ch13_csr[0] , _u0_ch13_txsz[31] ,_u0_ch13_txsz[30] , _u0_ch13_txsz[29] , _u0_ch13_txsz[28] ,_u0_ch13_txsz[27] , _u0_ch13_txsz[26] , _u0_ch13_txsz[25] ,_u0_ch13_txsz[24] , _u0_ch13_txsz[23] , _u0_ch13_txsz[22] ,_u0_ch13_txsz[21] , _u0_ch13_txsz[20] , _u0_ch13_txsz[19] ,_u0_ch13_txsz[18] , _u0_ch13_txsz[17] , _u0_ch13_txsz[16] ,_u0_ch13_txsz[15] , _u0_ch13_txsz[14] , _u0_ch13_txsz[13] ,_u0_ch13_txsz[12] , _u0_ch13_txsz[11] , _u0_ch13_txsz[10] ,_u0_ch13_txsz[9] , _u0_ch13_txsz[8] , _u0_ch13_txsz[7] ,_u0_ch13_txsz[6] , _u0_ch13_txsz[5] , _u0_ch13_txsz[4] ,_u0_ch13_txsz[3] , _u0_ch13_txsz[2] , _u0_ch13_txsz[1] ,_u0_ch13_txsz[0] , _u0_ch13_adr0[31] , _u0_ch13_adr0[30] ,_u0_ch13_adr0[29] , _u0_ch13_adr0[28] , _u0_ch13_adr0[27] ,_u0_ch13_adr0[26] , _u0_ch13_adr0[25] , _u0_ch13_adr0[24] ,_u0_ch13_adr0[23] , _u0_ch13_adr0[22] , _u0_ch13_adr0[21] ,_u0_ch13_adr0[20] , _u0_ch13_adr0[19] , _u0_ch13_adr0[18] ,_u0_ch13_adr0[17] , _u0_ch13_adr0[16] , _u0_ch13_adr0[15] ,_u0_ch13_adr0[14] , _u0_ch13_adr0[13] , _u0_ch13_adr0[12] ,_u0_ch13_adr0[11] , _u0_ch13_adr0[10] , _u0_ch13_adr0[9] ,_u0_ch13_adr0[8] , _u0_ch13_adr0[7] , _u0_ch13_adr0[6] ,_u0_ch13_adr0[5] , _u0_ch13_adr0[4] , _u0_ch13_adr0[3] ,_u0_ch13_adr0[2] , _u0_ch13_adr0[1] , _u0_ch13_adr0[0] ,_u0_ch13_adr1[31] , _u0_ch13_adr1[30] , _u0_ch13_adr1[29] ,_u0_ch13_adr1[28] , _u0_ch13_adr1[27] , _u0_ch13_adr1[26] ,_u0_ch13_adr1[25] , _u0_ch13_adr1[24] , _u0_ch13_adr1[23] ,_u0_ch13_adr1[22] , _u0_ch13_adr1[21] , _u0_ch13_adr1[20] ,_u0_ch13_adr1[19] , _u0_ch13_adr1[18] , _u0_ch13_adr1[17] ,_u0_ch13_adr1[16] , _u0_ch13_adr1[15] , _u0_ch13_adr1[14] ,_u0_ch13_adr1[13] , _u0_ch13_adr1[12] , _u0_ch13_adr1[11] ,_u0_ch13_adr1[10] , _u0_ch13_adr1[9] , _u0_ch13_adr1[8] ,_u0_ch13_adr1[7] , _u0_ch13_adr1[6] , _u0_ch13_adr1[5] ,_u0_ch13_adr1[4] , _u0_ch13_adr1[3] , _u0_ch13_adr1[2] ,_u0_ch13_adr1[1] , _u0_ch13_adr1[0] , _u0_ch13_am0[31] ,_u0_ch13_am0[30] , _u0_ch13_am0[29] , _u0_ch13_am0[28] ,_u0_ch13_am0[27] , _u0_ch13_am0[26] , _u0_ch13_am0[25] ,_u0_ch13_am0[24] , _u0_ch13_am0[23] , _u0_ch13_am0[22] ,_u0_ch13_am0[21] , _u0_ch13_am0[20] , _u0_ch13_am0[19] ,_u0_ch13_am0[18] , _u0_ch13_am0[17] , _u0_ch13_am0[16] ,_u0_ch13_am0[15] , _u0_ch13_am0[14] , _u0_ch13_am0[13] ,_u0_ch13_am0[12] , _u0_ch13_am0[11] , _u0_ch13_am0[10] ,_u0_ch13_am0[9] , _u0_ch13_am0[8] , _u0_ch13_am0[7] ,_u0_ch13_am0[6] , _u0_ch13_am0[5] , _u0_ch13_am0[4] ,_u0_ch13_am0[3] , _u0_ch13_am0[2] , _u0_ch13_am0[1] ,_u0_ch13_am0[0] , _u0_ch13_am1[31] , _u0_ch13_am1[30] ,_u0_ch13_am1[29] , _u0_ch13_am1[28] , _u0_ch13_am1[27] ,_u0_ch13_am1[26] , _u0_ch13_am1[25] , _u0_ch13_am1[24] ,_u0_ch13_am1[23] , _u0_ch13_am1[22] , _u0_ch13_am1[21] ,_u0_ch13_am1[20] , _u0_ch13_am1[19] , _u0_ch13_am1[18] ,_u0_ch13_am1[17] , _u0_ch13_am1[16] , _u0_ch13_am1[15] ,_u0_ch13_am1[14] , _u0_ch13_am1[13] , _u0_ch13_am1[12] ,_u0_ch13_am1[11] , _u0_ch13_am1[10] , _u0_ch13_am1[9] ,_u0_ch13_am1[8] , _u0_ch13_am1[7] , _u0_ch13_am1[6] ,_u0_ch13_am1[5] , _u0_ch13_am1[4] , _u0_ch13_am1[3] ,_u0_ch13_am1[2] , _u0_ch13_am1[1] , _u0_ch13_am1[0] ,_u0_pointer14[31] , _u0_pointer14[30] , _u0_pointer14[29] ,_u0_pointer14[28] , _u0_pointer14[27] , _u0_pointer14[26] ,_u0_pointer14[25] , _u0_pointer14[24] , _u0_pointer14[23] ,_u0_pointer14[22] , _u0_pointer14[21] , _u0_pointer14[20] ,_u0_pointer14[19] , _u0_pointer14[18] , _u0_pointer14[17] ,_u0_pointer14[16] , _u0_pointer14[15] , _u0_pointer14[14] ,_u0_pointer14[13] , _u0_pointer14[12] , _u0_pointer14[11] ,_u0_pointer14[10] , _u0_pointer14[9] , _u0_pointer14[8] ,_u0_pointer14[7] , _u0_pointer14[6] , _u0_pointer14[5] ,_u0_pointer14[4] , _u0_pointer14[3] , _u0_pointer14[2] ,_u0_pointer14[1] , _u0_pointer14[0] , _u0_pointer14_s[31] ,_u0_pointer14_s[30] , _u0_pointer14_s[29] , _u0_pointer14_s[28] ,_u0_pointer14_s[27] , _u0_pointer14_s[26] , _u0_pointer14_s[25] ,_u0_pointer14_s[24] , _u0_pointer14_s[23] , _u0_pointer14_s[22] ,_u0_pointer14_s[21] , _u0_pointer14_s[20] , _u0_pointer14_s[19] ,_u0_pointer14_s[18] , _u0_pointer14_s[17] , _u0_pointer14_s[16] ,_u0_pointer14_s[15] , _u0_pointer14_s[14] , _u0_pointer14_s[13] ,_u0_pointer14_s[12] , _u0_pointer14_s[11] , _u0_pointer14_s[10] ,_u0_pointer14_s[9] , _u0_pointer14_s[8] , _u0_pointer14_s[7] ,_u0_pointer14_s[6] , _u0_pointer14_s[5] , _u0_pointer14_s[4] ,_u0_pointer14_s[3] , _u0_pointer14_s[2] , _u0_pointer14_s[1] ,_u0_pointer14_s[0] , _u0_ch14_csr[31] , _u0_ch14_csr[30] ,_u0_ch14_csr[29] , _u0_ch14_csr[28] , _u0_ch14_csr[27] ,_u0_ch14_csr[26] , _u0_ch14_csr[25] , _u0_ch14_csr[24] ,_u0_ch14_csr[23] , _u0_ch14_csr[22] , _u0_ch14_csr[21] ,_u0_ch14_csr[20] , _u0_ch14_csr[19] , _u0_ch14_csr[18] ,_u0_ch14_csr[17] , _u0_ch14_csr[16] , _u0_ch14_csr[15] ,_u0_ch14_csr[14] , _u0_ch14_csr[13] , _u0_ch14_csr[12] ,_u0_ch14_csr[11] , _u0_ch14_csr[10] , _u0_ch14_csr[9] ,_u0_ch14_csr[8] , _u0_ch14_csr[7] , _u0_ch14_csr[6] ,_u0_ch14_csr[5] , _u0_ch14_csr[4] , _u0_ch14_csr[3] ,_u0_ch14_csr[2] , _u0_ch14_csr[1] , _u0_ch14_csr[0] ,_u0_ch14_txsz[31] , _u0_ch14_txsz[30] , _u0_ch14_txsz[29] ,_u0_ch14_txsz[28] , _u0_ch14_txsz[27] , _u0_ch14_txsz[26] ,_u0_ch14_txsz[25] , _u0_ch14_txsz[24] , _u0_ch14_txsz[23] ,_u0_ch14_txsz[22] , _u0_ch14_txsz[21] , _u0_ch14_txsz[20] ,_u0_ch14_txsz[19] , _u0_ch14_txsz[18] , _u0_ch14_txsz[17] ,_u0_ch14_txsz[16] , _u0_ch14_txsz[15] , _u0_ch14_txsz[14] ,_u0_ch14_txsz[13] , _u0_ch14_txsz[12] , _u0_ch14_txsz[11] ,_u0_ch14_txsz[10] , _u0_ch14_txsz[9] , _u0_ch14_txsz[8] ,_u0_ch14_txsz[7] , _u0_ch14_txsz[6] , _u0_ch14_txsz[5] ,_u0_ch14_txsz[4] , _u0_ch14_txsz[3] , _u0_ch14_txsz[2] ,_u0_ch14_txsz[1] , _u0_ch14_txsz[0] , _u0_ch14_adr0[31] ,_u0_ch14_adr0[30] , _u0_ch14_adr0[29] , _u0_ch14_adr0[28] ,_u0_ch14_adr0[27] , _u0_ch14_adr0[26] , _u0_ch14_adr0[25] ,_u0_ch14_adr0[24] , _u0_ch14_adr0[23] , _u0_ch14_adr0[22] ,_u0_ch14_adr0[21] , _u0_ch14_adr0[20] , _u0_ch14_adr0[19] ,_u0_ch14_adr0[18] , _u0_ch14_adr0[17] , _u0_ch14_adr0[16] ,_u0_ch14_adr0[15] , _u0_ch14_adr0[14] , _u0_ch14_adr0[13] ,_u0_ch14_adr0[12] , _u0_ch14_adr0[11] , _u0_ch14_adr0[10] ,_u0_ch14_adr0[9] , _u0_ch14_adr0[8] , _u0_ch14_adr0[7] ,_u0_ch14_adr0[6] , _u0_ch14_adr0[5] , _u0_ch14_adr0[4] ,_u0_ch14_adr0[3] , _u0_ch14_adr0[2] , _u0_ch14_adr0[1] ,_u0_ch14_adr0[0] , _u0_ch14_adr1[31] , _u0_ch14_adr1[30] ,_u0_ch14_adr1[29] , _u0_ch14_adr1[28] , _u0_ch14_adr1[27] ,_u0_ch14_adr1[26] , _u0_ch14_adr1[25] , _u0_ch14_adr1[24] ,_u0_ch14_adr1[23] , _u0_ch14_adr1[22] , _u0_ch14_adr1[21] ,_u0_ch14_adr1[20] , _u0_ch14_adr1[19] , _u0_ch14_adr1[18] ,_u0_ch14_adr1[17] , _u0_ch14_adr1[16] , _u0_ch14_adr1[15] ,_u0_ch14_adr1[14] , _u0_ch14_adr1[13] , _u0_ch14_adr1[12] ,_u0_ch14_adr1[11] , _u0_ch14_adr1[10] , _u0_ch14_adr1[9] ,_u0_ch14_adr1[8] , _u0_ch14_adr1[7] , _u0_ch14_adr1[6] ,_u0_ch14_adr1[5] , _u0_ch14_adr1[4] , _u0_ch14_adr1[3] ,_u0_ch14_adr1[2] , _u0_ch14_adr1[1] , _u0_ch14_adr1[0] ,_u0_ch14_am0[31] , _u0_ch14_am0[30] , _u0_ch14_am0[29] ,_u0_ch14_am0[28] , _u0_ch14_am0[27] , _u0_ch14_am0[26] ,_u0_ch14_am0[25] , _u0_ch14_am0[24] , _u0_ch14_am0[23] ,_u0_ch14_am0[22] , _u0_ch14_am0[21] , _u0_ch14_am0[20] ,_u0_ch14_am0[19] , _u0_ch14_am0[18] , _u0_ch14_am0[17] ,_u0_ch14_am0[16] , _u0_ch14_am0[15] , _u0_ch14_am0[14] ,_u0_ch14_am0[13] , _u0_ch14_am0[12] , _u0_ch14_am0[11] ,_u0_ch14_am0[10] , _u0_ch14_am0[9] , _u0_ch14_am0[8] ,_u0_ch14_am0[7] , _u0_ch14_am0[6] , _u0_ch14_am0[5] ,_u0_ch14_am0[4] , _u0_ch14_am0[3] , _u0_ch14_am0[2] ,_u0_ch14_am0[1] , _u0_ch14_am0[0] , _u0_ch14_am1[31] ,_u0_ch14_am1[30] , _u0_ch14_am1[29] , _u0_ch14_am1[28] ,_u0_ch14_am1[27] , _u0_ch14_am1[26] , _u0_ch14_am1[25] ,_u0_ch14_am1[24] , _u0_ch14_am1[23] , _u0_ch14_am1[22] ,_u0_ch14_am1[21] , _u0_ch14_am1[20] , _u0_ch14_am1[19] ,_u0_ch14_am1[18] , _u0_ch14_am1[17] , _u0_ch14_am1[16] ,_u0_ch14_am1[15] , _u0_ch14_am1[14] , _u0_ch14_am1[13] ,_u0_ch14_am1[12] , _u0_ch14_am1[11] , _u0_ch14_am1[10] ,_u0_ch14_am1[9] , _u0_ch14_am1[8] , _u0_ch14_am1[7] ,_u0_ch14_am1[6] , _u0_ch14_am1[5] , _u0_ch14_am1[4] ,_u0_ch14_am1[3] , _u0_ch14_am1[2] , _u0_ch14_am1[1] ,_u0_ch14_am1[0] , _u0_pointer15[31] , _u0_pointer15[30] ,_u0_pointer15[29] , _u0_pointer15[28] , _u0_pointer15[27] ,_u0_pointer15[26] , _u0_pointer15[25] , _u0_pointer15[24] ,_u0_pointer15[23] , _u0_pointer15[22] , _u0_pointer15[21] ,_u0_pointer15[20] , _u0_pointer15[19] , _u0_pointer15[18] ,_u0_pointer15[17] , _u0_pointer15[16] , _u0_pointer15[15] ,_u0_pointer15[14] , _u0_pointer15[13] , _u0_pointer15[12] ,_u0_pointer15[11] , _u0_pointer15[10] , _u0_pointer15[9] ,_u0_pointer15[8] , _u0_pointer15[7] , _u0_pointer15[6] ,_u0_pointer15[5] , _u0_pointer15[4] , _u0_pointer15[3] ,_u0_pointer15[2] , _u0_pointer15[1] , _u0_pointer15[0] ,_u0_pointer15_s[31] , _u0_pointer15_s[30] , _u0_pointer15_s[29] ,_u0_pointer15_s[28] , _u0_pointer15_s[27] , _u0_pointer15_s[26] ,_u0_pointer15_s[25] , _u0_pointer15_s[24] , _u0_pointer15_s[23] ,_u0_pointer15_s[22] , _u0_pointer15_s[21] , _u0_pointer15_s[20] ,_u0_pointer15_s[19] , _u0_pointer15_s[18] , _u0_pointer15_s[17] ,_u0_pointer15_s[16] , _u0_pointer15_s[15] , _u0_pointer15_s[14] ,_u0_pointer15_s[13] , _u0_pointer15_s[12] , _u0_pointer15_s[11] ,_u0_pointer15_s[10] , _u0_pointer15_s[9] , _u0_pointer15_s[8] ,_u0_pointer15_s[7] , _u0_pointer15_s[6] , _u0_pointer15_s[5] ,_u0_pointer15_s[4] , _u0_pointer15_s[3] , _u0_pointer15_s[2] ,_u0_pointer15_s[1] , _u0_pointer15_s[0] , _u0_ch15_csr[31] ,_u0_ch15_csr[30] , _u0_ch15_csr[29] , _u0_ch15_csr[28] ,_u0_ch15_csr[27] , _u0_ch15_csr[26] , _u0_ch15_csr[25] ,_u0_ch15_csr[24] , _u0_ch15_csr[23] , _u0_ch15_csr[22] ,_u0_ch15_csr[21] , _u0_ch15_csr[20] , _u0_ch15_csr[19] ,_u0_ch15_csr[18] , _u0_ch15_csr[17] , _u0_ch15_csr[16] ,_u0_ch15_csr[15] , _u0_ch15_csr[14] , _u0_ch15_csr[13] ,_u0_ch15_csr[12] , _u0_ch15_csr[11] , _u0_ch15_csr[10] ,_u0_ch15_csr[9] , _u0_ch15_csr[8] , _u0_ch15_csr[7] ,_u0_ch15_csr[6] , _u0_ch15_csr[5] , _u0_ch15_csr[4] ,_u0_ch15_csr[3] , _u0_ch15_csr[2] , _u0_ch15_csr[1] ,_u0_ch15_csr[0] , _u0_ch15_txsz[31] , _u0_ch15_txsz[30] ,_u0_ch15_txsz[29] , _u0_ch15_txsz[28] , _u0_ch15_txsz[27] ,_u0_ch15_txsz[26] , _u0_ch15_txsz[25] , _u0_ch15_txsz[24] ,_u0_ch15_txsz[23] , _u0_ch15_txsz[22] , _u0_ch15_txsz[21] ,_u0_ch15_txsz[20] , _u0_ch15_txsz[19] , _u0_ch15_txsz[18] ,_u0_ch15_txsz[17] , _u0_ch15_txsz[16] , _u0_ch15_txsz[15] ,_u0_ch15_txsz[14] , _u0_ch15_txsz[13] , _u0_ch15_txsz[12] ,_u0_ch15_txsz[11] , _u0_ch15_txsz[10] , _u0_ch15_txsz[9] ,_u0_ch15_txsz[8] , _u0_ch15_txsz[7] , _u0_ch15_txsz[6] ,_u0_ch15_txsz[5] , _u0_ch15_txsz[4] , _u0_ch15_txsz[3] ,_u0_ch15_txsz[2] , _u0_ch15_txsz[1] , _u0_ch15_txsz[0] ,_u0_ch15_adr0[31] , _u0_ch15_adr0[30] , _u0_ch15_adr0[29] ,_u0_ch15_adr0[28] , _u0_ch15_adr0[27] , _u0_ch15_adr0[26] ,_u0_ch15_adr0[25] , _u0_ch15_adr0[24] , _u0_ch15_adr0[23] ,_u0_ch15_adr0[22] , _u0_ch15_adr0[21] , _u0_ch15_adr0[20] ,_u0_ch15_adr0[19] , _u0_ch15_adr0[18] , _u0_ch15_adr0[17] ,_u0_ch15_adr0[16] , _u0_ch15_adr0[15] , _u0_ch15_adr0[14] ,_u0_ch15_adr0[13] , _u0_ch15_adr0[12] , _u0_ch15_adr0[11] ,_u0_ch15_adr0[10] , _u0_ch15_adr0[9] , _u0_ch15_adr0[8] ,_u0_ch15_adr0[7] , _u0_ch15_adr0[6] , _u0_ch15_adr0[5] ,_u0_ch15_adr0[4] , _u0_ch15_adr0[3] , _u0_ch15_adr0[2] ,_u0_ch15_adr0[1] , _u0_ch15_adr0[0] , _u0_ch15_adr1[31] ,_u0_ch15_adr1[30] , _u0_ch15_adr1[29] , _u0_ch15_adr1[28] ,_u0_ch15_adr1[27] , _u0_ch15_adr1[26] , _u0_ch15_adr1[25] ,_u0_ch15_adr1[24] , _u0_ch15_adr1[23] , _u0_ch15_adr1[22] ,_u0_ch15_adr1[21] , _u0_ch15_adr1[20] , _u0_ch15_adr1[19] ,_u0_ch15_adr1[18] , _u0_ch15_adr1[17] , _u0_ch15_adr1[16] ,_u0_ch15_adr1[15] , _u0_ch15_adr1[14] , _u0_ch15_adr1[13] ,_u0_ch15_adr1[12] , _u0_ch15_adr1[11] , _u0_ch15_adr1[10] ,_u0_ch15_adr1[9] , _u0_ch15_adr1[8] , _u0_ch15_adr1[7] ,_u0_ch15_adr1[6] , _u0_ch15_adr1[5] , _u0_ch15_adr1[4] ,_u0_ch15_adr1[3] , _u0_ch15_adr1[2] , _u0_ch15_adr1[1] ,_u0_ch15_adr1[0] , _u0_ch15_am0[31] , _u0_ch15_am0[30] ,_u0_ch15_am0[29] , _u0_ch15_am0[28] , _u0_ch15_am0[27] ,_u0_ch15_am0[26] , _u0_ch15_am0[25] , _u0_ch15_am0[24] ,_u0_ch15_am0[23] , _u0_ch15_am0[22] , _u0_ch15_am0[21] ,_u0_ch15_am0[20] , _u0_ch15_am0[19] , _u0_ch15_am0[18] ,_u0_ch15_am0[17] , _u0_ch15_am0[16] , _u0_ch15_am0[15] ,_u0_ch15_am0[14] , _u0_ch15_am0[13] , _u0_ch15_am0[12] ,_u0_ch15_am0[11] , _u0_ch15_am0[10] , _u0_ch15_am0[9] ,_u0_ch15_am0[8] , _u0_ch15_am0[7] , _u0_ch15_am0[6] ,_u0_ch15_am0[5] , _u0_ch15_am0[4] , _u0_ch15_am0[3] ,_u0_ch15_am0[2] , _u0_ch15_am0[1] , _u0_ch15_am0[0] ,_u0_ch15_am1[31] , _u0_ch15_am1[30] , _u0_ch15_am1[29] ,_u0_ch15_am1[28] , _u0_ch15_am1[27] , _u0_ch15_am1[26] ,_u0_ch15_am1[25] , _u0_ch15_am1[24] , _u0_ch15_am1[23] ,_u0_ch15_am1[22] , _u0_ch15_am1[21] , _u0_ch15_am1[20] ,_u0_ch15_am1[19] , _u0_ch15_am1[18] , _u0_ch15_am1[17] ,_u0_ch15_am1[16] , _u0_ch15_am1[15] , _u0_ch15_am1[14] ,_u0_ch15_am1[13] , _u0_ch15_am1[12] , _u0_ch15_am1[11] ,_u0_ch15_am1[10] , _u0_ch15_am1[9] , _u0_ch15_am1[8] ,_u0_ch15_am1[7] , _u0_ch15_am1[6] , _u0_ch15_am1[5] ,_u0_ch15_am1[4] , _u0_ch15_am1[3] , _u0_ch15_am1[2] ,_u0_ch15_am1[1] , _u0_ch15_am1[0] , _u0_pointer16[31] ,_u0_pointer16[30] , _u0_pointer16[29] , _u0_pointer16[28] ,_u0_pointer16[27] , _u0_pointer16[26] , _u0_pointer16[25] ,_u0_pointer16[24] , _u0_pointer16[23] , _u0_pointer16[22] ,_u0_pointer16[21] , _u0_pointer16[20] , _u0_pointer16[19] ,_u0_pointer16[18] , _u0_pointer16[17] , _u0_pointer16[16] ,_u0_pointer16[15] , _u0_pointer16[14] , _u0_pointer16[13] ,_u0_pointer16[12] , _u0_pointer16[11] , _u0_pointer16[10] ,_u0_pointer16[9] , _u0_pointer16[8] , _u0_pointer16[7] ,_u0_pointer16[6] , _u0_pointer16[5] , _u0_pointer16[4] ,_u0_pointer16[3] , _u0_pointer16[2] , _u0_pointer16[1] ,_u0_pointer16[0] , _u0_pointer16_s[31] , _u0_pointer16_s[30] ,_u0_pointer16_s[29] , _u0_pointer16_s[28] , _u0_pointer16_s[27] ,_u0_pointer16_s[26] , _u0_pointer16_s[25] , _u0_pointer16_s[24] ,_u0_pointer16_s[23] , _u0_pointer16_s[22] , _u0_pointer16_s[21] ,_u0_pointer16_s[20] , _u0_pointer16_s[19] , _u0_pointer16_s[18] ,_u0_pointer16_s[17] , _u0_pointer16_s[16] , _u0_pointer16_s[15] ,_u0_pointer16_s[14] , _u0_pointer16_s[13] , _u0_pointer16_s[12] ,_u0_pointer16_s[11] , _u0_pointer16_s[10] , _u0_pointer16_s[9] ,_u0_pointer16_s[8] , _u0_pointer16_s[7] , _u0_pointer16_s[6] ,_u0_pointer16_s[5] , _u0_pointer16_s[4] , _u0_pointer16_s[3] ,_u0_pointer16_s[2] , _u0_pointer16_s[1] , _u0_pointer16_s[0] ,_u0_ch16_csr[31] , _u0_ch16_csr[30] , _u0_ch16_csr[29] ,_u0_ch16_csr[28] , _u0_ch16_csr[27] , _u0_ch16_csr[26] ,_u0_ch16_csr[25] , _u0_ch16_csr[24] , _u0_ch16_csr[23] ,_u0_ch16_csr[22] , _u0_ch16_csr[21] , _u0_ch16_csr[20] ,_u0_ch16_csr[19] , _u0_ch16_csr[18] , _u0_ch16_csr[17] ,_u0_ch16_csr[16] , _u0_ch16_csr[15] , _u0_ch16_csr[14] ,_u0_ch16_csr[13] , _u0_ch16_csr[12] , _u0_ch16_csr[11] ,_u0_ch16_csr[10] , _u0_ch16_csr[9] , _u0_ch16_csr[8] ,_u0_ch16_csr[7] , _u0_ch16_csr[6] , _u0_ch16_csr[5] ,_u0_ch16_csr[4] , _u0_ch16_csr[3] , _u0_ch16_csr[2] ,_u0_ch16_csr[1] , _u0_ch16_csr[0] , _u0_ch16_txsz[31] ,_u0_ch16_txsz[30] , _u0_ch16_txsz[29] , _u0_ch16_txsz[28] ,_u0_ch16_txsz[27] , _u0_ch16_txsz[26] , _u0_ch16_txsz[25] ,_u0_ch16_txsz[24] , _u0_ch16_txsz[23] , _u0_ch16_txsz[22] ,_u0_ch16_txsz[21] , _u0_ch16_txsz[20] , _u0_ch16_txsz[19] ,_u0_ch16_txsz[18] , _u0_ch16_txsz[17] , _u0_ch16_txsz[16] ,_u0_ch16_txsz[15] , _u0_ch16_txsz[14] , _u0_ch16_txsz[13] ,_u0_ch16_txsz[12] , _u0_ch16_txsz[11] , _u0_ch16_txsz[10] ,_u0_ch16_txsz[9] , _u0_ch16_txsz[8] , _u0_ch16_txsz[7] ,_u0_ch16_txsz[6] , _u0_ch16_txsz[5] , _u0_ch16_txsz[4] ,_u0_ch16_txsz[3] , _u0_ch16_txsz[2] , _u0_ch16_txsz[1] ,_u0_ch16_txsz[0] , _u0_ch16_adr0[31] , _u0_ch16_adr0[30] ,_u0_ch16_adr0[29] , _u0_ch16_adr0[28] , _u0_ch16_adr0[27] ,_u0_ch16_adr0[26] , _u0_ch16_adr0[25] , _u0_ch16_adr0[24] ,_u0_ch16_adr0[23] , _u0_ch16_adr0[22] , _u0_ch16_adr0[21] ,_u0_ch16_adr0[20] , _u0_ch16_adr0[19] , _u0_ch16_adr0[18] ,_u0_ch16_adr0[17] , _u0_ch16_adr0[16] , _u0_ch16_adr0[15] ,_u0_ch16_adr0[14] , _u0_ch16_adr0[13] , _u0_ch16_adr0[12] ,_u0_ch16_adr0[11] , _u0_ch16_adr0[10] , _u0_ch16_adr0[9] ,_u0_ch16_adr0[8] , _u0_ch16_adr0[7] , _u0_ch16_adr0[6] ,_u0_ch16_adr0[5] , _u0_ch16_adr0[4] , _u0_ch16_adr0[3] ,_u0_ch16_adr0[2] , _u0_ch16_adr0[1] , _u0_ch16_adr0[0] ,_u0_ch16_adr1[31] , _u0_ch16_adr1[30] , _u0_ch16_adr1[29] ,_u0_ch16_adr1[28] , _u0_ch16_adr1[27] , _u0_ch16_adr1[26] ,_u0_ch16_adr1[25] , _u0_ch16_adr1[24] , _u0_ch16_adr1[23] ,_u0_ch16_adr1[22] , _u0_ch16_adr1[21] , _u0_ch16_adr1[20] ,_u0_ch16_adr1[19] , _u0_ch16_adr1[18] , _u0_ch16_adr1[17] ,_u0_ch16_adr1[16] , _u0_ch16_adr1[15] , _u0_ch16_adr1[14] ,_u0_ch16_adr1[13] , _u0_ch16_adr1[12] , _u0_ch16_adr1[11] ,_u0_ch16_adr1[10] , _u0_ch16_adr1[9] , _u0_ch16_adr1[8] ,_u0_ch16_adr1[7] , _u0_ch16_adr1[6] , _u0_ch16_adr1[5] ,_u0_ch16_adr1[4] , _u0_ch16_adr1[3] , _u0_ch16_adr1[2] ,_u0_ch16_adr1[1] , _u0_ch16_adr1[0] , _u0_ch16_am0[31] ,_u0_ch16_am0[30] , _u0_ch16_am0[29] , _u0_ch16_am0[28] ,_u0_ch16_am0[27] , _u0_ch16_am0[26] , _u0_ch16_am0[25] ,_u0_ch16_am0[24] , _u0_ch16_am0[23] , _u0_ch16_am0[22] ,_u0_ch16_am0[21] , _u0_ch16_am0[20] , _u0_ch16_am0[19] ,_u0_ch16_am0[18] , _u0_ch16_am0[17] , _u0_ch16_am0[16] ,_u0_ch16_am0[15] , _u0_ch16_am0[14] , _u0_ch16_am0[13] ,_u0_ch16_am0[12] , _u0_ch16_am0[11] , _u0_ch16_am0[10] ,_u0_ch16_am0[9] , _u0_ch16_am0[8] , _u0_ch16_am0[7] ,_u0_ch16_am0[6] , _u0_ch16_am0[5] , _u0_ch16_am0[4] ,_u0_ch16_am0[3] , _u0_ch16_am0[2] , _u0_ch16_am0[1] ,_u0_ch16_am0[0] , _u0_ch16_am1[31] , _u0_ch16_am1[30] ,_u0_ch16_am1[29] , _u0_ch16_am1[28] , _u0_ch16_am1[27] ,_u0_ch16_am1[26] , _u0_ch16_am1[25] , _u0_ch16_am1[24] ,_u0_ch16_am1[23] , _u0_ch16_am1[22] , _u0_ch16_am1[21] ,_u0_ch16_am1[20] , _u0_ch16_am1[19] , _u0_ch16_am1[18] ,_u0_ch16_am1[17] , _u0_ch16_am1[16] , _u0_ch16_am1[15] ,_u0_ch16_am1[14] , _u0_ch16_am1[13] , _u0_ch16_am1[12] ,_u0_ch16_am1[11] , _u0_ch16_am1[10] , _u0_ch16_am1[9] ,_u0_ch16_am1[8] , _u0_ch16_am1[7] , _u0_ch16_am1[6] ,_u0_ch16_am1[5] , _u0_ch16_am1[4] , _u0_ch16_am1[3] ,_u0_ch16_am1[2] , _u0_ch16_am1[1] , _u0_ch16_am1[0] ,_u0_pointer17[31] , _u0_pointer17[30] , _u0_pointer17[29] ,_u0_pointer17[28] , _u0_pointer17[27] , _u0_pointer17[26] ,_u0_pointer17[25] , _u0_pointer17[24] , _u0_pointer17[23] ,_u0_pointer17[22] , _u0_pointer17[21] , _u0_pointer17[20] ,_u0_pointer17[19] , _u0_pointer17[18] , _u0_pointer17[17] ,_u0_pointer17[16] , _u0_pointer17[15] , _u0_pointer17[14] ,_u0_pointer17[13] , _u0_pointer17[12] , _u0_pointer17[11] ,_u0_pointer17[10] , _u0_pointer17[9] , _u0_pointer17[8] ,_u0_pointer17[7] , _u0_pointer17[6] , _u0_pointer17[5] ,_u0_pointer17[4] , _u0_pointer17[3] , _u0_pointer17[2] ,_u0_pointer17[1] , _u0_pointer17[0] , _u0_pointer17_s[31] ,_u0_pointer17_s[30] , _u0_pointer17_s[29] , _u0_pointer17_s[28] ,_u0_pointer17_s[27] , _u0_pointer17_s[26] , _u0_pointer17_s[25] ,_u0_pointer17_s[24] , _u0_pointer17_s[23] , _u0_pointer17_s[22] ,_u0_pointer17_s[21] , _u0_pointer17_s[20] , _u0_pointer17_s[19] ,_u0_pointer17_s[18] , _u0_pointer17_s[17] , _u0_pointer17_s[16] ,_u0_pointer17_s[15] , _u0_pointer17_s[14] , _u0_pointer17_s[13] ,_u0_pointer17_s[12] , _u0_pointer17_s[11] , _u0_pointer17_s[10] ,_u0_pointer17_s[9] , _u0_pointer17_s[8] , _u0_pointer17_s[7] ,_u0_pointer17_s[6] , _u0_pointer17_s[5] , _u0_pointer17_s[4] ,_u0_pointer17_s[3] , _u0_pointer17_s[2] , _u0_pointer17_s[1] ,_u0_pointer17_s[0] , _u0_ch17_csr[31] , _u0_ch17_csr[30] ,_u0_ch17_csr[29] , _u0_ch17_csr[28] , _u0_ch17_csr[27] ,_u0_ch17_csr[26] , _u0_ch17_csr[25] , _u0_ch17_csr[24] ,_u0_ch17_csr[23] , _u0_ch17_csr[22] , _u0_ch17_csr[21] ,_u0_ch17_csr[20] , _u0_ch17_csr[19] , _u0_ch17_csr[18] ,_u0_ch17_csr[17] , _u0_ch17_csr[16] , _u0_ch17_csr[15] ,_u0_ch17_csr[14] , _u0_ch17_csr[13] , _u0_ch17_csr[12] ,_u0_ch17_csr[11] , _u0_ch17_csr[10] , _u0_ch17_csr[9] ,_u0_ch17_csr[8] , _u0_ch17_csr[7] , _u0_ch17_csr[6] ,_u0_ch17_csr[5] , _u0_ch17_csr[4] , _u0_ch17_csr[3] ,_u0_ch17_csr[2] , _u0_ch17_csr[1] , _u0_ch17_csr[0] ,_u0_ch17_txsz[31] , _u0_ch17_txsz[30] , _u0_ch17_txsz[29] ,_u0_ch17_txsz[28] , _u0_ch17_txsz[27] , _u0_ch17_txsz[26] ,_u0_ch17_txsz[25] , _u0_ch17_txsz[24] , _u0_ch17_txsz[23] ,_u0_ch17_txsz[22] , _u0_ch17_txsz[21] , _u0_ch17_txsz[20] ,_u0_ch17_txsz[19] , _u0_ch17_txsz[18] , _u0_ch17_txsz[17] ,_u0_ch17_txsz[16] , _u0_ch17_txsz[15] , _u0_ch17_txsz[14] ,_u0_ch17_txsz[13] , _u0_ch17_txsz[12] , _u0_ch17_txsz[11] ,_u0_ch17_txsz[10] , _u0_ch17_txsz[9] , _u0_ch17_txsz[8] ,_u0_ch17_txsz[7] , _u0_ch17_txsz[6] , _u0_ch17_txsz[5] ,_u0_ch17_txsz[4] , _u0_ch17_txsz[3] , _u0_ch17_txsz[2] ,_u0_ch17_txsz[1] , _u0_ch17_txsz[0] , _u0_ch17_adr0[31] ,_u0_ch17_adr0[30] , _u0_ch17_adr0[29] , _u0_ch17_adr0[28] ,_u0_ch17_adr0[27] , _u0_ch17_adr0[26] , _u0_ch17_adr0[25] ,_u0_ch17_adr0[24] , _u0_ch17_adr0[23] , _u0_ch17_adr0[22] ,_u0_ch17_adr0[21] , _u0_ch17_adr0[20] , _u0_ch17_adr0[19] ,_u0_ch17_adr0[18] , _u0_ch17_adr0[17] , _u0_ch17_adr0[16] ,_u0_ch17_adr0[15] , _u0_ch17_adr0[14] , _u0_ch17_adr0[13] ,_u0_ch17_adr0[12] , _u0_ch17_adr0[11] , _u0_ch17_adr0[10] ,_u0_ch17_adr0[9] , _u0_ch17_adr0[8] , _u0_ch17_adr0[7] ,_u0_ch17_adr0[6] , _u0_ch17_adr0[5] , _u0_ch17_adr0[4] ,_u0_ch17_adr0[3] , _u0_ch17_adr0[2] , _u0_ch17_adr0[1] ,_u0_ch17_adr0[0] , _u0_ch17_adr1[31] , _u0_ch17_adr1[30] ,_u0_ch17_adr1[29] , _u0_ch17_adr1[28] , _u0_ch17_adr1[27] ,_u0_ch17_adr1[26] , _u0_ch17_adr1[25] , _u0_ch17_adr1[24] ,_u0_ch17_adr1[23] , _u0_ch17_adr1[22] , _u0_ch17_adr1[21] ,_u0_ch17_adr1[20] , _u0_ch17_adr1[19] , _u0_ch17_adr1[18] ,_u0_ch17_adr1[17] , _u0_ch17_adr1[16] , _u0_ch17_adr1[15] ,_u0_ch17_adr1[14] , _u0_ch17_adr1[13] , _u0_ch17_adr1[12] ,_u0_ch17_adr1[11] , _u0_ch17_adr1[10] , _u0_ch17_adr1[9] ,_u0_ch17_adr1[8] , _u0_ch17_adr1[7] , _u0_ch17_adr1[6] ,_u0_ch17_adr1[5] , _u0_ch17_adr1[4] , _u0_ch17_adr1[3] ,_u0_ch17_adr1[2] , _u0_ch17_adr1[1] , _u0_ch17_adr1[0] ,_u0_ch17_am0[31] , _u0_ch17_am0[30] , _u0_ch17_am0[29] ,_u0_ch17_am0[28] , _u0_ch17_am0[27] , _u0_ch17_am0[26] ,_u0_ch17_am0[25] , _u0_ch17_am0[24] , _u0_ch17_am0[23] ,_u0_ch17_am0[22] , _u0_ch17_am0[21] , _u0_ch17_am0[20] ,_u0_ch17_am0[19] , _u0_ch17_am0[18] , _u0_ch17_am0[17] ,_u0_ch17_am0[16] , _u0_ch17_am0[15] , _u0_ch17_am0[14] ,_u0_ch17_am0[13] , _u0_ch17_am0[12] , _u0_ch17_am0[11] ,_u0_ch17_am0[10] , _u0_ch17_am0[9] , _u0_ch17_am0[8] ,_u0_ch17_am0[7] , _u0_ch17_am0[6] , _u0_ch17_am0[5] ,_u0_ch17_am0[4] , _u0_ch17_am0[3] , _u0_ch17_am0[2] ,_u0_ch17_am0[1] , _u0_ch17_am0[0] , _u0_ch17_am1[31] ,_u0_ch17_am1[30] , _u0_ch17_am1[29] , _u0_ch17_am1[28] ,_u0_ch17_am1[27] , _u0_ch17_am1[26] , _u0_ch17_am1[25] ,_u0_ch17_am1[24] , _u0_ch17_am1[23] , _u0_ch17_am1[22] ,_u0_ch17_am1[21] , _u0_ch17_am1[20] , _u0_ch17_am1[19] ,_u0_ch17_am1[18] , _u0_ch17_am1[17] , _u0_ch17_am1[16] ,_u0_ch17_am1[15] , _u0_ch17_am1[14] , _u0_ch17_am1[13] ,_u0_ch17_am1[12] , _u0_ch17_am1[11] , _u0_ch17_am1[10] ,_u0_ch17_am1[9] , _u0_ch17_am1[8] , _u0_ch17_am1[7] ,_u0_ch17_am1[6] , _u0_ch17_am1[5] , _u0_ch17_am1[4] ,_u0_ch17_am1[3] , _u0_ch17_am1[2] , _u0_ch17_am1[1] ,_u0_ch17_am1[0] , _u0_pointer18[31] , _u0_pointer18[30] ,_u0_pointer18[29] , _u0_pointer18[28] , _u0_pointer18[27] ,_u0_pointer18[26] , _u0_pointer18[25] , _u0_pointer18[24] ,_u0_pointer18[23] , _u0_pointer18[22] , _u0_pointer18[21] ,_u0_pointer18[20] , _u0_pointer18[19] , _u0_pointer18[18] ,_u0_pointer18[17] , _u0_pointer18[16] , _u0_pointer18[15] ,_u0_pointer18[14] , _u0_pointer18[13] , _u0_pointer18[12] ,_u0_pointer18[11] , _u0_pointer18[10] , _u0_pointer18[9] ,_u0_pointer18[8] , _u0_pointer18[7] , _u0_pointer18[6] ,_u0_pointer18[5] , _u0_pointer18[4] , _u0_pointer18[3] ,_u0_pointer18[2] , _u0_pointer18[1] , _u0_pointer18[0] ,_u0_pointer18_s[31] , _u0_pointer18_s[30] , _u0_pointer18_s[29] ,_u0_pointer18_s[28] , _u0_pointer18_s[27] , _u0_pointer18_s[26] ,_u0_pointer18_s[25] , _u0_pointer18_s[24] , _u0_pointer18_s[23] ,_u0_pointer18_s[22] , _u0_pointer18_s[21] , _u0_pointer18_s[20] ,_u0_pointer18_s[19] , _u0_pointer18_s[18] , _u0_pointer18_s[17] ,_u0_pointer18_s[16] , _u0_pointer18_s[15] , _u0_pointer18_s[14] ,_u0_pointer18_s[13] , _u0_pointer18_s[12] , _u0_pointer18_s[11] ,_u0_pointer18_s[10] , _u0_pointer18_s[9] , _u0_pointer18_s[8] ,_u0_pointer18_s[7] , _u0_pointer18_s[6] , _u0_pointer18_s[5] ,_u0_pointer18_s[4] , _u0_pointer18_s[3] , _u0_pointer18_s[2] ,_u0_pointer18_s[1] , _u0_pointer18_s[0] , _u0_ch18_csr[31] ,_u0_ch18_csr[30] , _u0_ch18_csr[29] , _u0_ch18_csr[28] ,_u0_ch18_csr[27] , _u0_ch18_csr[26] , _u0_ch18_csr[25] ,_u0_ch18_csr[24] , _u0_ch18_csr[23] , _u0_ch18_csr[22] ,_u0_ch18_csr[21] , _u0_ch18_csr[20] , _u0_ch18_csr[19] ,_u0_ch18_csr[18] , _u0_ch18_csr[17] , _u0_ch18_csr[16] ,_u0_ch18_csr[15] , _u0_ch18_csr[14] , _u0_ch18_csr[13] ,_u0_ch18_csr[12] , _u0_ch18_csr[11] , _u0_ch18_csr[10] ,_u0_ch18_csr[9] , _u0_ch18_csr[8] , _u0_ch18_csr[7] ,_u0_ch18_csr[6] , _u0_ch18_csr[5] , _u0_ch18_csr[4] ,_u0_ch18_csr[3] , _u0_ch18_csr[2] , _u0_ch18_csr[1] ,_u0_ch18_csr[0] , _u0_ch18_txsz[31] , _u0_ch18_txsz[30] ,_u0_ch18_txsz[29] , _u0_ch18_txsz[28] , _u0_ch18_txsz[27] ,_u0_ch18_txsz[26] , _u0_ch18_txsz[25] , _u0_ch18_txsz[24] ,_u0_ch18_txsz[23] , _u0_ch18_txsz[22] , _u0_ch18_txsz[21] ,_u0_ch18_txsz[20] , _u0_ch18_txsz[19] , _u0_ch18_txsz[18] ,_u0_ch18_txsz[17] , _u0_ch18_txsz[16] , _u0_ch18_txsz[15] ,_u0_ch18_txsz[14] , _u0_ch18_txsz[13] , _u0_ch18_txsz[12] ,_u0_ch18_txsz[11] , _u0_ch18_txsz[10] , _u0_ch18_txsz[9] ,_u0_ch18_txsz[8] , _u0_ch18_txsz[7] , _u0_ch18_txsz[6] ,_u0_ch18_txsz[5] , _u0_ch18_txsz[4] , _u0_ch18_txsz[3] ,_u0_ch18_txsz[2] , _u0_ch18_txsz[1] , _u0_ch18_txsz[0] ,_u0_ch18_adr0[31] , _u0_ch18_adr0[30] , _u0_ch18_adr0[29] ,_u0_ch18_adr0[28] , _u0_ch18_adr0[27] , _u0_ch18_adr0[26] ,_u0_ch18_adr0[25] , _u0_ch18_adr0[24] , _u0_ch18_adr0[23] ,_u0_ch18_adr0[22] , _u0_ch18_adr0[21] , _u0_ch18_adr0[20] ,_u0_ch18_adr0[19] , _u0_ch18_adr0[18] , _u0_ch18_adr0[17] ,_u0_ch18_adr0[16] , _u0_ch18_adr0[15] , _u0_ch18_adr0[14] ,_u0_ch18_adr0[13] , _u0_ch18_adr0[12] , _u0_ch18_adr0[11] ,_u0_ch18_adr0[10] , _u0_ch18_adr0[9] , _u0_ch18_adr0[8] ,_u0_ch18_adr0[7] , _u0_ch18_adr0[6] , _u0_ch18_adr0[5] ,_u0_ch18_adr0[4] , _u0_ch18_adr0[3] , _u0_ch18_adr0[2] ,_u0_ch18_adr0[1] , _u0_ch18_adr0[0] , _u0_ch18_adr1[31] ,_u0_ch18_adr1[30] , _u0_ch18_adr1[29] , _u0_ch18_adr1[28] ,_u0_ch18_adr1[27] , _u0_ch18_adr1[26] , _u0_ch18_adr1[25] ,_u0_ch18_adr1[24] , _u0_ch18_adr1[23] , _u0_ch18_adr1[22] ,_u0_ch18_adr1[21] , _u0_ch18_adr1[20] , _u0_ch18_adr1[19] ,_u0_ch18_adr1[18] , _u0_ch18_adr1[17] , _u0_ch18_adr1[16] ,_u0_ch18_adr1[15] , _u0_ch18_adr1[14] , _u0_ch18_adr1[13] ,_u0_ch18_adr1[12] , _u0_ch18_adr1[11] , _u0_ch18_adr1[10] ,_u0_ch18_adr1[9] , _u0_ch18_adr1[8] , _u0_ch18_adr1[7] ,_u0_ch18_adr1[6] , _u0_ch18_adr1[5] , _u0_ch18_adr1[4] ,_u0_ch18_adr1[3] , _u0_ch18_adr1[2] , _u0_ch18_adr1[1] ,_u0_ch18_adr1[0] , _u0_ch18_am0[31] , _u0_ch18_am0[30] ,_u0_ch18_am0[29] , _u0_ch18_am0[28] , _u0_ch18_am0[27] ,_u0_ch18_am0[26] , _u0_ch18_am0[25] , _u0_ch18_am0[24] ,_u0_ch18_am0[23] , _u0_ch18_am0[22] , _u0_ch18_am0[21] ,_u0_ch18_am0[20] , _u0_ch18_am0[19] , _u0_ch18_am0[18] ,_u0_ch18_am0[17] , _u0_ch18_am0[16] , _u0_ch18_am0[15] ,_u0_ch18_am0[14] , _u0_ch18_am0[13] , _u0_ch18_am0[12] ,_u0_ch18_am0[11] , _u0_ch18_am0[10] , _u0_ch18_am0[9] ,_u0_ch18_am0[8] , _u0_ch18_am0[7] , _u0_ch18_am0[6] ,_u0_ch18_am0[5] , _u0_ch18_am0[4] , _u0_ch18_am0[3] ,_u0_ch18_am0[2] , _u0_ch18_am0[1] , _u0_ch18_am0[0] ,_u0_ch18_am1[31] , _u0_ch18_am1[30] , _u0_ch18_am1[29] ,_u0_ch18_am1[28] , _u0_ch18_am1[27] , _u0_ch18_am1[26] ,_u0_ch18_am1[25] , _u0_ch18_am1[24] , _u0_ch18_am1[23] ,_u0_ch18_am1[22] , _u0_ch18_am1[21] , _u0_ch18_am1[20] ,_u0_ch18_am1[19] , _u0_ch18_am1[18] , _u0_ch18_am1[17] ,_u0_ch18_am1[16] , _u0_ch18_am1[15] , _u0_ch18_am1[14] ,_u0_ch18_am1[13] , _u0_ch18_am1[12] , _u0_ch18_am1[11] ,_u0_ch18_am1[10] , _u0_ch18_am1[9] , _u0_ch18_am1[8] ,_u0_ch18_am1[7] , _u0_ch18_am1[6] , _u0_ch18_am1[5] ,_u0_ch18_am1[4] , _u0_ch18_am1[3] , _u0_ch18_am1[2] ,_u0_ch18_am1[1] , _u0_ch18_am1[0] , _u0_pointer19[31] ,_u0_pointer19[30] , _u0_pointer19[29] , _u0_pointer19[28] ,_u0_pointer19[27] , _u0_pointer19[26] , _u0_pointer19[25] ,_u0_pointer19[24] , _u0_pointer19[23] , _u0_pointer19[22] ,_u0_pointer19[21] , _u0_pointer19[20] , _u0_pointer19[19] ,_u0_pointer19[18] , _u0_pointer19[17] , _u0_pointer19[16] ,_u0_pointer19[15] , _u0_pointer19[14] , _u0_pointer19[13] ,_u0_pointer19[12] , _u0_pointer19[11] , _u0_pointer19[10] ,_u0_pointer19[9] , _u0_pointer19[8] , _u0_pointer19[7] ,_u0_pointer19[6] , _u0_pointer19[5] , _u0_pointer19[4] ,_u0_pointer19[3] , _u0_pointer19[2] , _u0_pointer19[1] ,_u0_pointer19[0] , _u0_pointer19_s[31] , _u0_pointer19_s[30] ,_u0_pointer19_s[29] , _u0_pointer19_s[28] , _u0_pointer19_s[27] ,_u0_pointer19_s[26] , _u0_pointer19_s[25] , _u0_pointer19_s[24] ,_u0_pointer19_s[23] , _u0_pointer19_s[22] , _u0_pointer19_s[21] ,_u0_pointer19_s[20] , _u0_pointer19_s[19] , _u0_pointer19_s[18] ,_u0_pointer19_s[17] , _u0_pointer19_s[16] , _u0_pointer19_s[15] ,_u0_pointer19_s[14] , _u0_pointer19_s[13] , _u0_pointer19_s[12] ,_u0_pointer19_s[11] , _u0_pointer19_s[10] , _u0_pointer19_s[9] ,_u0_pointer19_s[8] , _u0_pointer19_s[7] , _u0_pointer19_s[6] ,_u0_pointer19_s[5] , _u0_pointer19_s[4] , _u0_pointer19_s[3] ,_u0_pointer19_s[2] , _u0_pointer19_s[1] , _u0_pointer19_s[0] ,_u0_ch19_csr[31] , _u0_ch19_csr[30] , _u0_ch19_csr[29] ,_u0_ch19_csr[28] , _u0_ch19_csr[27] , _u0_ch19_csr[26] ,_u0_ch19_csr[25] , _u0_ch19_csr[24] , _u0_ch19_csr[23] ,_u0_ch19_csr[22] , _u0_ch19_csr[21] , _u0_ch19_csr[20] ,_u0_ch19_csr[19] , _u0_ch19_csr[18] , _u0_ch19_csr[17] ,_u0_ch19_csr[16] , _u0_ch19_csr[15] , _u0_ch19_csr[14] ,_u0_ch19_csr[13] , _u0_ch19_csr[12] , _u0_ch19_csr[11] ,_u0_ch19_csr[10] , _u0_ch19_csr[9] , _u0_ch19_csr[8] ,_u0_ch19_csr[7] , _u0_ch19_csr[6] , _u0_ch19_csr[5] ,_u0_ch19_csr[4] , _u0_ch19_csr[3] , _u0_ch19_csr[2] ,_u0_ch19_csr[1] , _u0_ch19_csr[0] , _u0_ch19_txsz[31] ,_u0_ch19_txsz[30] , _u0_ch19_txsz[29] , _u0_ch19_txsz[28] ,_u0_ch19_txsz[27] , _u0_ch19_txsz[26] , _u0_ch19_txsz[25] ,_u0_ch19_txsz[24] , _u0_ch19_txsz[23] , _u0_ch19_txsz[22] ,_u0_ch19_txsz[21] , _u0_ch19_txsz[20] , _u0_ch19_txsz[19] ,_u0_ch19_txsz[18] , _u0_ch19_txsz[17] , _u0_ch19_txsz[16] ,_u0_ch19_txsz[15] , _u0_ch19_txsz[14] , _u0_ch19_txsz[13] ,_u0_ch19_txsz[12] , _u0_ch19_txsz[11] , _u0_ch19_txsz[10] ,_u0_ch19_txsz[9] , _u0_ch19_txsz[8] , _u0_ch19_txsz[7] ,_u0_ch19_txsz[6] , _u0_ch19_txsz[5] , _u0_ch19_txsz[4] ,_u0_ch19_txsz[3] , _u0_ch19_txsz[2] , _u0_ch19_txsz[1] ,_u0_ch19_txsz[0] , _u0_ch19_adr0[31] , _u0_ch19_adr0[30] ,_u0_ch19_adr0[29] , _u0_ch19_adr0[28] , _u0_ch19_adr0[27] ,_u0_ch19_adr0[26] , _u0_ch19_adr0[25] , _u0_ch19_adr0[24] ,_u0_ch19_adr0[23] , _u0_ch19_adr0[22] , _u0_ch19_adr0[21] ,_u0_ch19_adr0[20] , _u0_ch19_adr0[19] , _u0_ch19_adr0[18] ,_u0_ch19_adr0[17] , _u0_ch19_adr0[16] , _u0_ch19_adr0[15] ,_u0_ch19_adr0[14] , _u0_ch19_adr0[13] , _u0_ch19_adr0[12] ,_u0_ch19_adr0[11] , _u0_ch19_adr0[10] , _u0_ch19_adr0[9] ,_u0_ch19_adr0[8] , _u0_ch19_adr0[7] , _u0_ch19_adr0[6] ,_u0_ch19_adr0[5] , _u0_ch19_adr0[4] , _u0_ch19_adr0[3] ,_u0_ch19_adr0[2] , _u0_ch19_adr0[1] , _u0_ch19_adr0[0] ,_u0_ch19_adr1[31] , _u0_ch19_adr1[30] , _u0_ch19_adr1[29] ,_u0_ch19_adr1[28] , _u0_ch19_adr1[27] , _u0_ch19_adr1[26] ,_u0_ch19_adr1[25] , _u0_ch19_adr1[24] , _u0_ch19_adr1[23] ,_u0_ch19_adr1[22] , _u0_ch19_adr1[21] , _u0_ch19_adr1[20] ,_u0_ch19_adr1[19] , _u0_ch19_adr1[18] , _u0_ch19_adr1[17] ,_u0_ch19_adr1[16] , _u0_ch19_adr1[15] , _u0_ch19_adr1[14] ,_u0_ch19_adr1[13] , _u0_ch19_adr1[12] , _u0_ch19_adr1[11] ,_u0_ch19_adr1[10] , _u0_ch19_adr1[9] , _u0_ch19_adr1[8] ,_u0_ch19_adr1[7] , _u0_ch19_adr1[6] , _u0_ch19_adr1[5] ,_u0_ch19_adr1[4] , _u0_ch19_adr1[3] , _u0_ch19_adr1[2] ,_u0_ch19_adr1[1] , _u0_ch19_adr1[0] , _u0_ch19_am0[31] ,_u0_ch19_am0[30] , _u0_ch19_am0[29] , _u0_ch19_am0[28] ,_u0_ch19_am0[27] , _u0_ch19_am0[26] , _u0_ch19_am0[25] ,_u0_ch19_am0[24] , _u0_ch19_am0[23] , _u0_ch19_am0[22] ,_u0_ch19_am0[21] , _u0_ch19_am0[20] , _u0_ch19_am0[19] ,_u0_ch19_am0[18] , _u0_ch19_am0[17] , _u0_ch19_am0[16] ,_u0_ch19_am0[15] , _u0_ch19_am0[14] , _u0_ch19_am0[13] ,_u0_ch19_am0[12] , _u0_ch19_am0[11] , _u0_ch19_am0[10] ,_u0_ch19_am0[9] , _u0_ch19_am0[8] , _u0_ch19_am0[7] ,_u0_ch19_am0[6] , _u0_ch19_am0[5] , _u0_ch19_am0[4] ,_u0_ch19_am0[3] , _u0_ch19_am0[2] , _u0_ch19_am0[1] ,_u0_ch19_am0[0] , _u0_ch19_am1[31] , _u0_ch19_am1[30] ,_u0_ch19_am1[29] , _u0_ch19_am1[28] , _u0_ch19_am1[27] ,_u0_ch19_am1[26] , _u0_ch19_am1[25] , _u0_ch19_am1[24] ,_u0_ch19_am1[23] , _u0_ch19_am1[22] , _u0_ch19_am1[21] ,_u0_ch19_am1[20] , _u0_ch19_am1[19] , _u0_ch19_am1[18] ,_u0_ch19_am1[17] , _u0_ch19_am1[16] , _u0_ch19_am1[15] ,_u0_ch19_am1[14] , _u0_ch19_am1[13] , _u0_ch19_am1[12] ,_u0_ch19_am1[11] , _u0_ch19_am1[10] , _u0_ch19_am1[9] ,_u0_ch19_am1[8] , _u0_ch19_am1[7] , _u0_ch19_am1[6] ,_u0_ch19_am1[5] , _u0_ch19_am1[4] , _u0_ch19_am1[3] ,_u0_ch19_am1[2] , _u0_ch19_am1[1] , _u0_ch19_am1[0] ,_u0_pointer20[31] , _u0_pointer20[30] , _u0_pointer20[29] ,_u0_pointer20[28] , _u0_pointer20[27] , _u0_pointer20[26] ,_u0_pointer20[25] , _u0_pointer20[24] , _u0_pointer20[23] ,_u0_pointer20[22] , _u0_pointer20[21] , _u0_pointer20[20] ,_u0_pointer20[19] , _u0_pointer20[18] , _u0_pointer20[17] ,_u0_pointer20[16] , _u0_pointer20[15] , _u0_pointer20[14] ,_u0_pointer20[13] , _u0_pointer20[12] , _u0_pointer20[11] ,_u0_pointer20[10] , _u0_pointer20[9] , _u0_pointer20[8] ,_u0_pointer20[7] , _u0_pointer20[6] , _u0_pointer20[5] ,_u0_pointer20[4] , _u0_pointer20[3] , _u0_pointer20[2] ,_u0_pointer20[1] , _u0_pointer20[0] , _u0_pointer20_s[31] ,_u0_pointer20_s[30] , _u0_pointer20_s[29] , _u0_pointer20_s[28] ,_u0_pointer20_s[27] , _u0_pointer20_s[26] , _u0_pointer20_s[25] ,_u0_pointer20_s[24] , _u0_pointer20_s[23] , _u0_pointer20_s[22] ,_u0_pointer20_s[21] , _u0_pointer20_s[20] , _u0_pointer20_s[19] ,_u0_pointer20_s[18] , _u0_pointer20_s[17] , _u0_pointer20_s[16] ,_u0_pointer20_s[15] , _u0_pointer20_s[14] , _u0_pointer20_s[13] ,_u0_pointer20_s[12] , _u0_pointer20_s[11] , _u0_pointer20_s[10] ,_u0_pointer20_s[9] , _u0_pointer20_s[8] , _u0_pointer20_s[7] ,_u0_pointer20_s[6] , _u0_pointer20_s[5] , _u0_pointer20_s[4] ,_u0_pointer20_s[3] , _u0_pointer20_s[2] , _u0_pointer20_s[1] ,_u0_pointer20_s[0] , _u0_ch20_csr[31] , _u0_ch20_csr[30] ,_u0_ch20_csr[29] , _u0_ch20_csr[28] , _u0_ch20_csr[27] ,_u0_ch20_csr[26] , _u0_ch20_csr[25] , _u0_ch20_csr[24] ,_u0_ch20_csr[23] , _u0_ch20_csr[22] , _u0_ch20_csr[21] ,_u0_ch20_csr[20] , _u0_ch20_csr[19] , _u0_ch20_csr[18] ,_u0_ch20_csr[17] , _u0_ch20_csr[16] , _u0_ch20_csr[15] ,_u0_ch20_csr[14] , _u0_ch20_csr[13] , _u0_ch20_csr[12] ,_u0_ch20_csr[11] , _u0_ch20_csr[10] , _u0_ch20_csr[9] ,_u0_ch20_csr[8] , _u0_ch20_csr[7] , _u0_ch20_csr[6] ,_u0_ch20_csr[5] , _u0_ch20_csr[4] , _u0_ch20_csr[3] ,_u0_ch20_csr[2] , _u0_ch20_csr[1] , _u0_ch20_csr[0] ,_u0_ch20_txsz[31] , _u0_ch20_txsz[30] , _u0_ch20_txsz[29] ,_u0_ch20_txsz[28] , _u0_ch20_txsz[27] , _u0_ch20_txsz[26] ,_u0_ch20_txsz[25] , _u0_ch20_txsz[24] , _u0_ch20_txsz[23] ,_u0_ch20_txsz[22] , _u0_ch20_txsz[21] , _u0_ch20_txsz[20] ,_u0_ch20_txsz[19] , _u0_ch20_txsz[18] , _u0_ch20_txsz[17] ,_u0_ch20_txsz[16] , _u0_ch20_txsz[15] , _u0_ch20_txsz[14] ,_u0_ch20_txsz[13] , _u0_ch20_txsz[12] , _u0_ch20_txsz[11] ,_u0_ch20_txsz[10] , _u0_ch20_txsz[9] , _u0_ch20_txsz[8] ,_u0_ch20_txsz[7] , _u0_ch20_txsz[6] , _u0_ch20_txsz[5] ,_u0_ch20_txsz[4] , _u0_ch20_txsz[3] , _u0_ch20_txsz[2] ,_u0_ch20_txsz[1] , _u0_ch20_txsz[0] , _u0_ch20_adr0[31] ,_u0_ch20_adr0[30] , _u0_ch20_adr0[29] , _u0_ch20_adr0[28] ,_u0_ch20_adr0[27] , _u0_ch20_adr0[26] , _u0_ch20_adr0[25] ,_u0_ch20_adr0[24] , _u0_ch20_adr0[23] , _u0_ch20_adr0[22] ,_u0_ch20_adr0[21] , _u0_ch20_adr0[20] , _u0_ch20_adr0[19] ,_u0_ch20_adr0[18] , _u0_ch20_adr0[17] , _u0_ch20_adr0[16] ,_u0_ch20_adr0[15] , _u0_ch20_adr0[14] , _u0_ch20_adr0[13] ,_u0_ch20_adr0[12] , _u0_ch20_adr0[11] , _u0_ch20_adr0[10] ,_u0_ch20_adr0[9] , _u0_ch20_adr0[8] , _u0_ch20_adr0[7] ,_u0_ch20_adr0[6] , _u0_ch20_adr0[5] , _u0_ch20_adr0[4] ,_u0_ch20_adr0[3] , _u0_ch20_adr0[2] , _u0_ch20_adr0[1] ,_u0_ch20_adr0[0] , _u0_ch20_adr1[31] , _u0_ch20_adr1[30] ,_u0_ch20_adr1[29] , _u0_ch20_adr1[28] , _u0_ch20_adr1[27] ,_u0_ch20_adr1[26] , _u0_ch20_adr1[25] , _u0_ch20_adr1[24] ,_u0_ch20_adr1[23] , _u0_ch20_adr1[22] , _u0_ch20_adr1[21] ,_u0_ch20_adr1[20] , _u0_ch20_adr1[19] , _u0_ch20_adr1[18] ,_u0_ch20_adr1[17] , _u0_ch20_adr1[16] , _u0_ch20_adr1[15] ,_u0_ch20_adr1[14] , _u0_ch20_adr1[13] , _u0_ch20_adr1[12] ,_u0_ch20_adr1[11] , _u0_ch20_adr1[10] , _u0_ch20_adr1[9] ,_u0_ch20_adr1[8] , _u0_ch20_adr1[7] , _u0_ch20_adr1[6] ,_u0_ch20_adr1[5] , _u0_ch20_adr1[4] , _u0_ch20_adr1[3] ,_u0_ch20_adr1[2] , _u0_ch20_adr1[1] , _u0_ch20_adr1[0] ,_u0_ch20_am0[31] , _u0_ch20_am0[30] , _u0_ch20_am0[29] ,_u0_ch20_am0[28] , _u0_ch20_am0[27] , _u0_ch20_am0[26] ,_u0_ch20_am0[25] , _u0_ch20_am0[24] , _u0_ch20_am0[23] ,_u0_ch20_am0[22] , _u0_ch20_am0[21] , _u0_ch20_am0[20] ,_u0_ch20_am0[19] , _u0_ch20_am0[18] , _u0_ch20_am0[17] ,_u0_ch20_am0[16] , _u0_ch20_am0[15] , _u0_ch20_am0[14] ,_u0_ch20_am0[13] , _u0_ch20_am0[12] , _u0_ch20_am0[11] ,_u0_ch20_am0[10] , _u0_ch20_am0[9] , _u0_ch20_am0[8] ,_u0_ch20_am0[7] , _u0_ch20_am0[6] , _u0_ch20_am0[5] ,_u0_ch20_am0[4] , _u0_ch20_am0[3] , _u0_ch20_am0[2] ,_u0_ch20_am0[1] , _u0_ch20_am0[0] , _u0_ch20_am1[31] ,_u0_ch20_am1[30] , _u0_ch20_am1[29] , _u0_ch20_am1[28] ,_u0_ch20_am1[27] , _u0_ch20_am1[26] , _u0_ch20_am1[25] ,_u0_ch20_am1[24] , _u0_ch20_am1[23] , _u0_ch20_am1[22] ,_u0_ch20_am1[21] , _u0_ch20_am1[20] , _u0_ch20_am1[19] ,_u0_ch20_am1[18] , _u0_ch20_am1[17] , _u0_ch20_am1[16] ,_u0_ch20_am1[15] , _u0_ch20_am1[14] , _u0_ch20_am1[13] ,_u0_ch20_am1[12] , _u0_ch20_am1[11] , _u0_ch20_am1[10] ,_u0_ch20_am1[9] , _u0_ch20_am1[8] , _u0_ch20_am1[7] ,_u0_ch20_am1[6] , _u0_ch20_am1[5] , _u0_ch20_am1[4] ,_u0_ch20_am1[3] , _u0_ch20_am1[2] , _u0_ch20_am1[1] ,_u0_ch20_am1[0] , _u0_pointer21[31] , _u0_pointer21[30] ,_u0_pointer21[29] , _u0_pointer21[28] , _u0_pointer21[27] ,_u0_pointer21[26] , _u0_pointer21[25] , _u0_pointer21[24] ,_u0_pointer21[23] , _u0_pointer21[22] , _u0_pointer21[21] ,_u0_pointer21[20] , _u0_pointer21[19] , _u0_pointer21[18] ,_u0_pointer21[17] , _u0_pointer21[16] , _u0_pointer21[15] ,_u0_pointer21[14] , _u0_pointer21[13] , _u0_pointer21[12] ,_u0_pointer21[11] , _u0_pointer21[10] , _u0_pointer21[9] ,_u0_pointer21[8] , _u0_pointer21[7] , _u0_pointer21[6] ,_u0_pointer21[5] , _u0_pointer21[4] , _u0_pointer21[3] ,_u0_pointer21[2] , _u0_pointer21[1] , _u0_pointer21[0] ,_u0_pointer21_s[31] , _u0_pointer21_s[30] , _u0_pointer21_s[29] ,_u0_pointer21_s[28] , _u0_pointer21_s[27] , _u0_pointer21_s[26] ,_u0_pointer21_s[25] , _u0_pointer21_s[24] , _u0_pointer21_s[23] ,_u0_pointer21_s[22] , _u0_pointer21_s[21] , _u0_pointer21_s[20] ,_u0_pointer21_s[19] , _u0_pointer21_s[18] , _u0_pointer21_s[17] ,_u0_pointer21_s[16] , _u0_pointer21_s[15] , _u0_pointer21_s[14] ,_u0_pointer21_s[13] , _u0_pointer21_s[12] , _u0_pointer21_s[11] ,_u0_pointer21_s[10] , _u0_pointer21_s[9] , _u0_pointer21_s[8] ,_u0_pointer21_s[7] , _u0_pointer21_s[6] , _u0_pointer21_s[5] ,_u0_pointer21_s[4] , _u0_pointer21_s[3] , _u0_pointer21_s[2] ,_u0_pointer21_s[1] , _u0_pointer21_s[0] , _u0_ch21_csr[31] ,_u0_ch21_csr[30] , _u0_ch21_csr[29] , _u0_ch21_csr[28] ,_u0_ch21_csr[27] , _u0_ch21_csr[26] , _u0_ch21_csr[25] ,_u0_ch21_csr[24] , _u0_ch21_csr[23] , _u0_ch21_csr[22] ,_u0_ch21_csr[21] , _u0_ch21_csr[20] , _u0_ch21_csr[19] ,_u0_ch21_csr[18] , _u0_ch21_csr[17] , _u0_ch21_csr[16] ,_u0_ch21_csr[15] , _u0_ch21_csr[14] , _u0_ch21_csr[13] ,_u0_ch21_csr[12] , _u0_ch21_csr[11] , _u0_ch21_csr[10] ,_u0_ch21_csr[9] , _u0_ch21_csr[8] , _u0_ch21_csr[7] ,_u0_ch21_csr[6] , _u0_ch21_csr[5] , _u0_ch21_csr[4] ,_u0_ch21_csr[3] , _u0_ch21_csr[2] , _u0_ch21_csr[1] ,_u0_ch21_csr[0] , _u0_ch21_txsz[31] , _u0_ch21_txsz[30] ,_u0_ch21_txsz[29] , _u0_ch21_txsz[28] , _u0_ch21_txsz[27] ,_u0_ch21_txsz[26] , _u0_ch21_txsz[25] , _u0_ch21_txsz[24] ,_u0_ch21_txsz[23] , _u0_ch21_txsz[22] , _u0_ch21_txsz[21] ,_u0_ch21_txsz[20] , _u0_ch21_txsz[19] , _u0_ch21_txsz[18] ,_u0_ch21_txsz[17] , _u0_ch21_txsz[16] , _u0_ch21_txsz[15] ,_u0_ch21_txsz[14] , _u0_ch21_txsz[13] , _u0_ch21_txsz[12] ,_u0_ch21_txsz[11] , _u0_ch21_txsz[10] , _u0_ch21_txsz[9] ,_u0_ch21_txsz[8] , _u0_ch21_txsz[7] , _u0_ch21_txsz[6] ,_u0_ch21_txsz[5] , _u0_ch21_txsz[4] , _u0_ch21_txsz[3] ,_u0_ch21_txsz[2] , _u0_ch21_txsz[1] , _u0_ch21_txsz[0] ,_u0_ch21_adr0[31] , _u0_ch21_adr0[30] , _u0_ch21_adr0[29] ,_u0_ch21_adr0[28] , _u0_ch21_adr0[27] , _u0_ch21_adr0[26] ,_u0_ch21_adr0[25] , _u0_ch21_adr0[24] , _u0_ch21_adr0[23] ,_u0_ch21_adr0[22] , _u0_ch21_adr0[21] , _u0_ch21_adr0[20] ,_u0_ch21_adr0[19] , _u0_ch21_adr0[18] , _u0_ch21_adr0[17] ,_u0_ch21_adr0[16] , _u0_ch21_adr0[15] , _u0_ch21_adr0[14] ,_u0_ch21_adr0[13] , _u0_ch21_adr0[12] , _u0_ch21_adr0[11] ,_u0_ch21_adr0[10] , _u0_ch21_adr0[9] , _u0_ch21_adr0[8] ,_u0_ch21_adr0[7] , _u0_ch21_adr0[6] , _u0_ch21_adr0[5] ,_u0_ch21_adr0[4] , _u0_ch21_adr0[3] , _u0_ch21_adr0[2] ,_u0_ch21_adr0[1] , _u0_ch21_adr0[0] , _u0_ch21_adr1[31] ,_u0_ch21_adr1[30] , _u0_ch21_adr1[29] , _u0_ch21_adr1[28] ,_u0_ch21_adr1[27] , _u0_ch21_adr1[26] , _u0_ch21_adr1[25] ,_u0_ch21_adr1[24] , _u0_ch21_adr1[23] , _u0_ch21_adr1[22] ,_u0_ch21_adr1[21] , _u0_ch21_adr1[20] , _u0_ch21_adr1[19] ,_u0_ch21_adr1[18] , _u0_ch21_adr1[17] , _u0_ch21_adr1[16] ,_u0_ch21_adr1[15] , _u0_ch21_adr1[14] , _u0_ch21_adr1[13] ,_u0_ch21_adr1[12] , _u0_ch21_adr1[11] , _u0_ch21_adr1[10] ,_u0_ch21_adr1[9] , _u0_ch21_adr1[8] , _u0_ch21_adr1[7] ,_u0_ch21_adr1[6] , _u0_ch21_adr1[5] , _u0_ch21_adr1[4] ,_u0_ch21_adr1[3] , _u0_ch21_adr1[2] , _u0_ch21_adr1[1] ,_u0_ch21_adr1[0] , _u0_ch21_am0[31] , _u0_ch21_am0[30] ,_u0_ch21_am0[29] , _u0_ch21_am0[28] , _u0_ch21_am0[27] ,_u0_ch21_am0[26] , _u0_ch21_am0[25] , _u0_ch21_am0[24] ,_u0_ch21_am0[23] , _u0_ch21_am0[22] , _u0_ch21_am0[21] ,_u0_ch21_am0[20] , _u0_ch21_am0[19] , _u0_ch21_am0[18] ,_u0_ch21_am0[17] , _u0_ch21_am0[16] , _u0_ch21_am0[15] ,_u0_ch21_am0[14] , _u0_ch21_am0[13] , _u0_ch21_am0[12] ,_u0_ch21_am0[11] , _u0_ch21_am0[10] , _u0_ch21_am0[9] ,_u0_ch21_am0[8] , _u0_ch21_am0[7] , _u0_ch21_am0[6] ,_u0_ch21_am0[5] , _u0_ch21_am0[4] , _u0_ch21_am0[3] ,_u0_ch21_am0[2] , _u0_ch21_am0[1] , _u0_ch21_am0[0] ,_u0_ch21_am1[31] , _u0_ch21_am1[30] , _u0_ch21_am1[29] ,_u0_ch21_am1[28] , _u0_ch21_am1[27] , _u0_ch21_am1[26] ,_u0_ch21_am1[25] , _u0_ch21_am1[24] , _u0_ch21_am1[23] ,_u0_ch21_am1[22] , _u0_ch21_am1[21] , _u0_ch21_am1[20] ,_u0_ch21_am1[19] , _u0_ch21_am1[18] , _u0_ch21_am1[17] ,_u0_ch21_am1[16] , _u0_ch21_am1[15] , _u0_ch21_am1[14] ,_u0_ch21_am1[13] , _u0_ch21_am1[12] , _u0_ch21_am1[11] ,_u0_ch21_am1[10] , _u0_ch21_am1[9] , _u0_ch21_am1[8] ,_u0_ch21_am1[7] , _u0_ch21_am1[6] , _u0_ch21_am1[5] ,_u0_ch21_am1[4] , _u0_ch21_am1[3] , _u0_ch21_am1[2] ,_u0_ch21_am1[1] , _u0_ch21_am1[0] , _u0_pointer22[31] ,_u0_pointer22[30] , _u0_pointer22[29] , _u0_pointer22[28] ,_u0_pointer22[27] , _u0_pointer22[26] , _u0_pointer22[25] ,_u0_pointer22[24] , _u0_pointer22[23] , _u0_pointer22[22] ,_u0_pointer22[21] , _u0_pointer22[20] , _u0_pointer22[19] ,_u0_pointer22[18] , _u0_pointer22[17] , _u0_pointer22[16] ,_u0_pointer22[15] , _u0_pointer22[14] , _u0_pointer22[13] ,_u0_pointer22[12] , _u0_pointer22[11] , _u0_pointer22[10] ,_u0_pointer22[9] , _u0_pointer22[8] , _u0_pointer22[7] ,_u0_pointer22[6] , _u0_pointer22[5] , _u0_pointer22[4] ,_u0_pointer22[3] , _u0_pointer22[2] , _u0_pointer22[1] ,_u0_pointer22[0] , _u0_pointer22_s[31] , _u0_pointer22_s[30] ,_u0_pointer22_s[29] , _u0_pointer22_s[28] , _u0_pointer22_s[27] ,_u0_pointer22_s[26] , _u0_pointer22_s[25] , _u0_pointer22_s[24] ,_u0_pointer22_s[23] , _u0_pointer22_s[22] , _u0_pointer22_s[21] ,_u0_pointer22_s[20] , _u0_pointer22_s[19] , _u0_pointer22_s[18] ,_u0_pointer22_s[17] , _u0_pointer22_s[16] , _u0_pointer22_s[15] ,_u0_pointer22_s[14] , _u0_pointer22_s[13] , _u0_pointer22_s[12] ,_u0_pointer22_s[11] , _u0_pointer22_s[10] , _u0_pointer22_s[9] ,_u0_pointer22_s[8] , _u0_pointer22_s[7] , _u0_pointer22_s[6] ,_u0_pointer22_s[5] , _u0_pointer22_s[4] , _u0_pointer22_s[3] ,_u0_pointer22_s[2] , _u0_pointer22_s[1] , _u0_pointer22_s[0] ,_u0_ch22_csr[31] , _u0_ch22_csr[30] , _u0_ch22_csr[29] ,_u0_ch22_csr[28] , _u0_ch22_csr[27] , _u0_ch22_csr[26] ,_u0_ch22_csr[25] , _u0_ch22_csr[24] , _u0_ch22_csr[23] ,_u0_ch22_csr[22] , _u0_ch22_csr[21] , _u0_ch22_csr[20] ,_u0_ch22_csr[19] , _u0_ch22_csr[18] , _u0_ch22_csr[17] ,_u0_ch22_csr[16] , _u0_ch22_csr[15] , _u0_ch22_csr[14] ,_u0_ch22_csr[13] , _u0_ch22_csr[12] , _u0_ch22_csr[11] ,_u0_ch22_csr[10] , _u0_ch22_csr[9] , _u0_ch22_csr[8] ,_u0_ch22_csr[7] , _u0_ch22_csr[6] , _u0_ch22_csr[5] ,_u0_ch22_csr[4] , _u0_ch22_csr[3] , _u0_ch22_csr[2] ,_u0_ch22_csr[1] , _u0_ch22_csr[0] , _u0_ch22_txsz[31] ,_u0_ch22_txsz[30] , _u0_ch22_txsz[29] , _u0_ch22_txsz[28] ,_u0_ch22_txsz[27] , _u0_ch22_txsz[26] , _u0_ch22_txsz[25] ,_u0_ch22_txsz[24] , _u0_ch22_txsz[23] , _u0_ch22_txsz[22] ,_u0_ch22_txsz[21] , _u0_ch22_txsz[20] , _u0_ch22_txsz[19] ,_u0_ch22_txsz[18] , _u0_ch22_txsz[17] , _u0_ch22_txsz[16] ,_u0_ch22_txsz[15] , _u0_ch22_txsz[14] , _u0_ch22_txsz[13] ,_u0_ch22_txsz[12] , _u0_ch22_txsz[11] , _u0_ch22_txsz[10] ,_u0_ch22_txsz[9] , _u0_ch22_txsz[8] , _u0_ch22_txsz[7] ,_u0_ch22_txsz[6] , _u0_ch22_txsz[5] , _u0_ch22_txsz[4] ,_u0_ch22_txsz[3] , _u0_ch22_txsz[2] , _u0_ch22_txsz[1] ,_u0_ch22_txsz[0] , _u0_ch22_adr0[31] , _u0_ch22_adr0[30] ,_u0_ch22_adr0[29] , _u0_ch22_adr0[28] , _u0_ch22_adr0[27] ,_u0_ch22_adr0[26] , _u0_ch22_adr0[25] , _u0_ch22_adr0[24] ,_u0_ch22_adr0[23] , _u0_ch22_adr0[22] , _u0_ch22_adr0[21] ,_u0_ch22_adr0[20] , _u0_ch22_adr0[19] , _u0_ch22_adr0[18] ,_u0_ch22_adr0[17] , _u0_ch22_adr0[16] , _u0_ch22_adr0[15] ,_u0_ch22_adr0[14] , _u0_ch22_adr0[13] , _u0_ch22_adr0[12] ,_u0_ch22_adr0[11] , _u0_ch22_adr0[10] , _u0_ch22_adr0[9] ,_u0_ch22_adr0[8] , _u0_ch22_adr0[7] , _u0_ch22_adr0[6] ,_u0_ch22_adr0[5] , _u0_ch22_adr0[4] , _u0_ch22_adr0[3] ,_u0_ch22_adr0[2] , _u0_ch22_adr0[1] , _u0_ch22_adr0[0] ,_u0_ch22_adr1[31] , _u0_ch22_adr1[30] , _u0_ch22_adr1[29] ,_u0_ch22_adr1[28] , _u0_ch22_adr1[27] , _u0_ch22_adr1[26] ,_u0_ch22_adr1[25] , _u0_ch22_adr1[24] , _u0_ch22_adr1[23] ,_u0_ch22_adr1[22] , _u0_ch22_adr1[21] , _u0_ch22_adr1[20] ,_u0_ch22_adr1[19] , _u0_ch22_adr1[18] , _u0_ch22_adr1[17] ,_u0_ch22_adr1[16] , _u0_ch22_adr1[15] , _u0_ch22_adr1[14] ,_u0_ch22_adr1[13] , _u0_ch22_adr1[12] , _u0_ch22_adr1[11] ,_u0_ch22_adr1[10] , _u0_ch22_adr1[9] , _u0_ch22_adr1[8] ,_u0_ch22_adr1[7] , _u0_ch22_adr1[6] , _u0_ch22_adr1[5] ,_u0_ch22_adr1[4] , _u0_ch22_adr1[3] , _u0_ch22_adr1[2] ,_u0_ch22_adr1[1] , _u0_ch22_adr1[0] , _u0_ch22_am0[31] ,_u0_ch22_am0[30] , _u0_ch22_am0[29] , _u0_ch22_am0[28] ,_u0_ch22_am0[27] , _u0_ch22_am0[26] , _u0_ch22_am0[25] ,_u0_ch22_am0[24] , _u0_ch22_am0[23] , _u0_ch22_am0[22] ,_u0_ch22_am0[21] , _u0_ch22_am0[20] , _u0_ch22_am0[19] ,_u0_ch22_am0[18] , _u0_ch22_am0[17] , _u0_ch22_am0[16] ,_u0_ch22_am0[15] , _u0_ch22_am0[14] , _u0_ch22_am0[13] ,_u0_ch22_am0[12] , _u0_ch22_am0[11] , _u0_ch22_am0[10] ,_u0_ch22_am0[9] , _u0_ch22_am0[8] , _u0_ch22_am0[7] ,_u0_ch22_am0[6] , _u0_ch22_am0[5] , _u0_ch22_am0[4] ,_u0_ch22_am0[3] , _u0_ch22_am0[2] , _u0_ch22_am0[1] ,_u0_ch22_am0[0] , _u0_ch22_am1[31] , _u0_ch22_am1[30] ,_u0_ch22_am1[29] , _u0_ch22_am1[28] , _u0_ch22_am1[27] ,_u0_ch22_am1[26] , _u0_ch22_am1[25] , _u0_ch22_am1[24] ,_u0_ch22_am1[23] , _u0_ch22_am1[22] , _u0_ch22_am1[21] ,_u0_ch22_am1[20] , _u0_ch22_am1[19] , _u0_ch22_am1[18] ,_u0_ch22_am1[17] , _u0_ch22_am1[16] , _u0_ch22_am1[15] ,_u0_ch22_am1[14] , _u0_ch22_am1[13] , _u0_ch22_am1[12] ,_u0_ch22_am1[11] , _u0_ch22_am1[10] , _u0_ch22_am1[9] ,_u0_ch22_am1[8] , _u0_ch22_am1[7] , _u0_ch22_am1[6] ,_u0_ch22_am1[5] , _u0_ch22_am1[4] , _u0_ch22_am1[3] ,_u0_ch22_am1[2] , _u0_ch22_am1[1] , _u0_ch22_am1[0] ,_u0_pointer23[31] , _u0_pointer23[30] , _u0_pointer23[29] ,_u0_pointer23[28] , _u0_pointer23[27] , _u0_pointer23[26] ,_u0_pointer23[25] , _u0_pointer23[24] , _u0_pointer23[23] ,_u0_pointer23[22] , _u0_pointer23[21] , _u0_pointer23[20] ,_u0_pointer23[19] , _u0_pointer23[18] , _u0_pointer23[17] ,_u0_pointer23[16] , _u0_pointer23[15] , _u0_pointer23[14] ,_u0_pointer23[13] , _u0_pointer23[12] , _u0_pointer23[11] ,_u0_pointer23[10] , _u0_pointer23[9] , _u0_pointer23[8] ,_u0_pointer23[7] , _u0_pointer23[6] , _u0_pointer23[5] ,_u0_pointer23[4] , _u0_pointer23[3] , _u0_pointer23[2] ,_u0_pointer23[1] , _u0_pointer23[0] , _u0_pointer23_s[31] ,_u0_pointer23_s[30] , _u0_pointer23_s[29] , _u0_pointer23_s[28] ,_u0_pointer23_s[27] , _u0_pointer23_s[26] , _u0_pointer23_s[25] ,_u0_pointer23_s[24] , _u0_pointer23_s[23] , _u0_pointer23_s[22] ,_u0_pointer23_s[21] , _u0_pointer23_s[20] , _u0_pointer23_s[19] ,_u0_pointer23_s[18] , _u0_pointer23_s[17] , _u0_pointer23_s[16] ,_u0_pointer23_s[15] , _u0_pointer23_s[14] , _u0_pointer23_s[13] ,_u0_pointer23_s[12] , _u0_pointer23_s[11] , _u0_pointer23_s[10] ,_u0_pointer23_s[9] , _u0_pointer23_s[8] , _u0_pointer23_s[7] ,_u0_pointer23_s[6] , _u0_pointer23_s[5] , _u0_pointer23_s[4] ,_u0_pointer23_s[3] , _u0_pointer23_s[2] , _u0_pointer23_s[1] ,_u0_pointer23_s[0] , _u0_ch23_csr[31] , _u0_ch23_csr[30] ,_u0_ch23_csr[29] , _u0_ch23_csr[28] , _u0_ch23_csr[27] ,_u0_ch23_csr[26] , _u0_ch23_csr[25] , _u0_ch23_csr[24] ,_u0_ch23_csr[23] , _u0_ch23_csr[22] , _u0_ch23_csr[21] ,_u0_ch23_csr[20] , _u0_ch23_csr[19] , _u0_ch23_csr[18] ,_u0_ch23_csr[17] , _u0_ch23_csr[16] , _u0_ch23_csr[15] ,_u0_ch23_csr[14] , _u0_ch23_csr[13] , _u0_ch23_csr[12] ,_u0_ch23_csr[11] , _u0_ch23_csr[10] , _u0_ch23_csr[9] ,_u0_ch23_csr[8] , _u0_ch23_csr[7] , _u0_ch23_csr[6] ,_u0_ch23_csr[5] , _u0_ch23_csr[4] , _u0_ch23_csr[3] ,_u0_ch23_csr[2] , _u0_ch23_csr[1] , _u0_ch23_csr[0] ,_u0_ch23_txsz[31] , _u0_ch23_txsz[30] , _u0_ch23_txsz[29] ,_u0_ch23_txsz[28] , _u0_ch23_txsz[27] , _u0_ch23_txsz[26] ,_u0_ch23_txsz[25] , _u0_ch23_txsz[24] , _u0_ch23_txsz[23] ,_u0_ch23_txsz[22] , _u0_ch23_txsz[21] , _u0_ch23_txsz[20] ,_u0_ch23_txsz[19] , _u0_ch23_txsz[18] , _u0_ch23_txsz[17] ,_u0_ch23_txsz[16] , _u0_ch23_txsz[15] , _u0_ch23_txsz[14] ,_u0_ch23_txsz[13] , _u0_ch23_txsz[12] , _u0_ch23_txsz[11] ,_u0_ch23_txsz[10] , _u0_ch23_txsz[9] , _u0_ch23_txsz[8] ,_u0_ch23_txsz[7] , _u0_ch23_txsz[6] , _u0_ch23_txsz[5] ,_u0_ch23_txsz[4] , _u0_ch23_txsz[3] , _u0_ch23_txsz[2] ,_u0_ch23_txsz[1] , _u0_ch23_txsz[0] , _u0_ch23_adr0[31] ,_u0_ch23_adr0[30] , _u0_ch23_adr0[29] , _u0_ch23_adr0[28] ,_u0_ch23_adr0[27] , _u0_ch23_adr0[26] , _u0_ch23_adr0[25] ,_u0_ch23_adr0[24] , _u0_ch23_adr0[23] , _u0_ch23_adr0[22] ,_u0_ch23_adr0[21] , _u0_ch23_adr0[20] , _u0_ch23_adr0[19] ,_u0_ch23_adr0[18] , _u0_ch23_adr0[17] , _u0_ch23_adr0[16] ,_u0_ch23_adr0[15] , _u0_ch23_adr0[14] , _u0_ch23_adr0[13] ,_u0_ch23_adr0[12] , _u0_ch23_adr0[11] , _u0_ch23_adr0[10] ,_u0_ch23_adr0[9] , _u0_ch23_adr0[8] , _u0_ch23_adr0[7] ,_u0_ch23_adr0[6] , _u0_ch23_adr0[5] , _u0_ch23_adr0[4] ,_u0_ch23_adr0[3] , _u0_ch23_adr0[2] , _u0_ch23_adr0[1] ,_u0_ch23_adr0[0] , _u0_ch23_adr1[31] , _u0_ch23_adr1[30] ,_u0_ch23_adr1[29] , _u0_ch23_adr1[28] , _u0_ch23_adr1[27] ,_u0_ch23_adr1[26] , _u0_ch23_adr1[25] , _u0_ch23_adr1[24] ,_u0_ch23_adr1[23] , _u0_ch23_adr1[22] , _u0_ch23_adr1[21] ,_u0_ch23_adr1[20] , _u0_ch23_adr1[19] , _u0_ch23_adr1[18] ,_u0_ch23_adr1[17] , _u0_ch23_adr1[16] , _u0_ch23_adr1[15] ,_u0_ch23_adr1[14] , _u0_ch23_adr1[13] , _u0_ch23_adr1[12] ,_u0_ch23_adr1[11] , _u0_ch23_adr1[10] , _u0_ch23_adr1[9] ,_u0_ch23_adr1[8] , _u0_ch23_adr1[7] , _u0_ch23_adr1[6] ,_u0_ch23_adr1[5] , _u0_ch23_adr1[4] , _u0_ch23_adr1[3] ,_u0_ch23_adr1[2] , _u0_ch23_adr1[1] , _u0_ch23_adr1[0] ,_u0_ch23_am0[31] , _u0_ch23_am0[30] , _u0_ch23_am0[29] ,_u0_ch23_am0[28] , _u0_ch23_am0[27] , _u0_ch23_am0[26] ,_u0_ch23_am0[25] , _u0_ch23_am0[24] , _u0_ch23_am0[23] ,_u0_ch23_am0[22] , _u0_ch23_am0[21] , _u0_ch23_am0[20] ,_u0_ch23_am0[19] , _u0_ch23_am0[18] , _u0_ch23_am0[17] ,_u0_ch23_am0[16] , _u0_ch23_am0[15] , _u0_ch23_am0[14] ,_u0_ch23_am0[13] , _u0_ch23_am0[12] , _u0_ch23_am0[11] ,_u0_ch23_am0[10] , _u0_ch23_am0[9] , _u0_ch23_am0[8] ,_u0_ch23_am0[7] , _u0_ch23_am0[6] , _u0_ch23_am0[5] ,_u0_ch23_am0[4] , _u0_ch23_am0[3] , _u0_ch23_am0[2] ,_u0_ch23_am0[1] , _u0_ch23_am0[0] , _u0_ch23_am1[31] ,_u0_ch23_am1[30] , _u0_ch23_am1[29] , _u0_ch23_am1[28] ,_u0_ch23_am1[27] , _u0_ch23_am1[26] , _u0_ch23_am1[25] ,_u0_ch23_am1[24] , _u0_ch23_am1[23] , _u0_ch23_am1[22] ,_u0_ch23_am1[21] , _u0_ch23_am1[20] , _u0_ch23_am1[19] ,_u0_ch23_am1[18] , _u0_ch23_am1[17] , _u0_ch23_am1[16] ,_u0_ch23_am1[15] , _u0_ch23_am1[14] , _u0_ch23_am1[13] ,_u0_ch23_am1[12] , _u0_ch23_am1[11] , _u0_ch23_am1[10] ,_u0_ch23_am1[9] , _u0_ch23_am1[8] , _u0_ch23_am1[7] ,_u0_ch23_am1[6] , _u0_ch23_am1[5] , _u0_ch23_am1[4] ,_u0_ch23_am1[3] , _u0_ch23_am1[2] , _u0_ch23_am1[1] ,_u0_ch23_am1[0] , _u0_pointer24[31] , _u0_pointer24[30] ,_u0_pointer24[29] , _u0_pointer24[28] , _u0_pointer24[27] ,_u0_pointer24[26] , _u0_pointer24[25] , _u0_pointer24[24] ,_u0_pointer24[23] , _u0_pointer24[22] , _u0_pointer24[21] ,_u0_pointer24[20] , _u0_pointer24[19] , _u0_pointer24[18] ,_u0_pointer24[17] , _u0_pointer24[16] , _u0_pointer24[15] ,_u0_pointer24[14] , _u0_pointer24[13] , _u0_pointer24[12] ,_u0_pointer24[11] , _u0_pointer24[10] , _u0_pointer24[9] ,_u0_pointer24[8] , _u0_pointer24[7] , _u0_pointer24[6] ,_u0_pointer24[5] , _u0_pointer24[4] , _u0_pointer24[3] ,_u0_pointer24[2] , _u0_pointer24[1] , _u0_pointer24[0] ,_u0_pointer24_s[31] , _u0_pointer24_s[30] , _u0_pointer24_s[29] ,_u0_pointer24_s[28] , _u0_pointer24_s[27] , _u0_pointer24_s[26] ,_u0_pointer24_s[25] , _u0_pointer24_s[24] , _u0_pointer24_s[23] ,_u0_pointer24_s[22] , _u0_pointer24_s[21] , _u0_pointer24_s[20] ,_u0_pointer24_s[19] , _u0_pointer24_s[18] , _u0_pointer24_s[17] ,_u0_pointer24_s[16] , _u0_pointer24_s[15] , _u0_pointer24_s[14] ,_u0_pointer24_s[13] , _u0_pointer24_s[12] , _u0_pointer24_s[11] ,_u0_pointer24_s[10] , _u0_pointer24_s[9] , _u0_pointer24_s[8] ,_u0_pointer24_s[7] , _u0_pointer24_s[6] , _u0_pointer24_s[5] ,_u0_pointer24_s[4] , _u0_pointer24_s[3] , _u0_pointer24_s[2] ,_u0_pointer24_s[1] , _u0_pointer24_s[0] , _u0_ch24_csr[31] ,_u0_ch24_csr[30] , _u0_ch24_csr[29] , _u0_ch24_csr[28] ,_u0_ch24_csr[27] , _u0_ch24_csr[26] , _u0_ch24_csr[25] ,_u0_ch24_csr[24] , _u0_ch24_csr[23] , _u0_ch24_csr[22] ,_u0_ch24_csr[21] , _u0_ch24_csr[20] , _u0_ch24_csr[19] ,_u0_ch24_csr[18] , _u0_ch24_csr[17] , _u0_ch24_csr[16] ,_u0_ch24_csr[15] , _u0_ch24_csr[14] , _u0_ch24_csr[13] ,_u0_ch24_csr[12] , _u0_ch24_csr[11] , _u0_ch24_csr[10] ,_u0_ch24_csr[9] , _u0_ch24_csr[8] , _u0_ch24_csr[7] ,_u0_ch24_csr[6] , _u0_ch24_csr[5] , _u0_ch24_csr[4] ,_u0_ch24_csr[3] , _u0_ch24_csr[2] , _u0_ch24_csr[1] ,_u0_ch24_csr[0] , _u0_ch24_txsz[31] , _u0_ch24_txsz[30] ,_u0_ch24_txsz[29] , _u0_ch24_txsz[28] , _u0_ch24_txsz[27] ,_u0_ch24_txsz[26] , _u0_ch24_txsz[25] , _u0_ch24_txsz[24] ,_u0_ch24_txsz[23] , _u0_ch24_txsz[22] , _u0_ch24_txsz[21] ,_u0_ch24_txsz[20] , _u0_ch24_txsz[19] , _u0_ch24_txsz[18] ,_u0_ch24_txsz[17] , _u0_ch24_txsz[16] , _u0_ch24_txsz[15] ,_u0_ch24_txsz[14] , _u0_ch24_txsz[13] , _u0_ch24_txsz[12] ,_u0_ch24_txsz[11] , _u0_ch24_txsz[10] , _u0_ch24_txsz[9] ,_u0_ch24_txsz[8] , _u0_ch24_txsz[7] , _u0_ch24_txsz[6] ,_u0_ch24_txsz[5] , _u0_ch24_txsz[4] , _u0_ch24_txsz[3] ,_u0_ch24_txsz[2] , _u0_ch24_txsz[1] , _u0_ch24_txsz[0] ,_u0_ch24_adr0[31] , _u0_ch24_adr0[30] , _u0_ch24_adr0[29] ,_u0_ch24_adr0[28] , _u0_ch24_adr0[27] , _u0_ch24_adr0[26] ,_u0_ch24_adr0[25] , _u0_ch24_adr0[24] , _u0_ch24_adr0[23] ,_u0_ch24_adr0[22] , _u0_ch24_adr0[21] , _u0_ch24_adr0[20] ,_u0_ch24_adr0[19] , _u0_ch24_adr0[18] , _u0_ch24_adr0[17] ,_u0_ch24_adr0[16] , _u0_ch24_adr0[15] , _u0_ch24_adr0[14] ,_u0_ch24_adr0[13] , _u0_ch24_adr0[12] , _u0_ch24_adr0[11] ,_u0_ch24_adr0[10] , _u0_ch24_adr0[9] , _u0_ch24_adr0[8] ,_u0_ch24_adr0[7] , _u0_ch24_adr0[6] , _u0_ch24_adr0[5] ,_u0_ch24_adr0[4] , _u0_ch24_adr0[3] , _u0_ch24_adr0[2] ,_u0_ch24_adr0[1] , _u0_ch24_adr0[0] , _u0_ch24_adr1[31] ,_u0_ch24_adr1[30] , _u0_ch24_adr1[29] , _u0_ch24_adr1[28] ,_u0_ch24_adr1[27] , _u0_ch24_adr1[26] , _u0_ch24_adr1[25] ,_u0_ch24_adr1[24] , _u0_ch24_adr1[23] , _u0_ch24_adr1[22] ,_u0_ch24_adr1[21] , _u0_ch24_adr1[20] , _u0_ch24_adr1[19] ,_u0_ch24_adr1[18] , _u0_ch24_adr1[17] , _u0_ch24_adr1[16] ,_u0_ch24_adr1[15] , _u0_ch24_adr1[14] , _u0_ch24_adr1[13] ,_u0_ch24_adr1[12] , _u0_ch24_adr1[11] , _u0_ch24_adr1[10] ,_u0_ch24_adr1[9] , _u0_ch24_adr1[8] , _u0_ch24_adr1[7] ,_u0_ch24_adr1[6] , _u0_ch24_adr1[5] , _u0_ch24_adr1[4] ,_u0_ch24_adr1[3] , _u0_ch24_adr1[2] , _u0_ch24_adr1[1] ,_u0_ch24_adr1[0] , _u0_ch24_am0[31] , _u0_ch24_am0[30] ,_u0_ch24_am0[29] , _u0_ch24_am0[28] , _u0_ch24_am0[27] ,_u0_ch24_am0[26] , _u0_ch24_am0[25] , _u0_ch24_am0[24] ,_u0_ch24_am0[23] , _u0_ch24_am0[22] , _u0_ch24_am0[21] ,_u0_ch24_am0[20] , _u0_ch24_am0[19] , _u0_ch24_am0[18] ,_u0_ch24_am0[17] , _u0_ch24_am0[16] , _u0_ch24_am0[15] ,_u0_ch24_am0[14] , _u0_ch24_am0[13] , _u0_ch24_am0[12] ,_u0_ch24_am0[11] , _u0_ch24_am0[10] , _u0_ch24_am0[9] ,_u0_ch24_am0[8] , _u0_ch24_am0[7] , _u0_ch24_am0[6] ,_u0_ch24_am0[5] , _u0_ch24_am0[4] , _u0_ch24_am0[3] ,_u0_ch24_am0[2] , _u0_ch24_am0[1] , _u0_ch24_am0[0] ,_u0_ch24_am1[31] , _u0_ch24_am1[30] , _u0_ch24_am1[29] ,_u0_ch24_am1[28] , _u0_ch24_am1[27] , _u0_ch24_am1[26] ,_u0_ch24_am1[25] , _u0_ch24_am1[24] , _u0_ch24_am1[23] ,_u0_ch24_am1[22] , _u0_ch24_am1[21] , _u0_ch24_am1[20] ,_u0_ch24_am1[19] , _u0_ch24_am1[18] , _u0_ch24_am1[17] ,_u0_ch24_am1[16] , _u0_ch24_am1[15] , _u0_ch24_am1[14] ,_u0_ch24_am1[13] , _u0_ch24_am1[12] , _u0_ch24_am1[11] ,_u0_ch24_am1[10] , _u0_ch24_am1[9] , _u0_ch24_am1[8] ,_u0_ch24_am1[7] , _u0_ch24_am1[6] , _u0_ch24_am1[5] ,_u0_ch24_am1[4] , _u0_ch24_am1[3] , _u0_ch24_am1[2] ,_u0_ch24_am1[1] , _u0_ch24_am1[0] , _u0_pointer25[31] ,_u0_pointer25[30] , _u0_pointer25[29] , _u0_pointer25[28] ,_u0_pointer25[27] , _u0_pointer25[26] , _u0_pointer25[25] ,_u0_pointer25[24] , _u0_pointer25[23] , _u0_pointer25[22] ,_u0_pointer25[21] , _u0_pointer25[20] , _u0_pointer25[19] ,_u0_pointer25[18] , _u0_pointer25[17] , _u0_pointer25[16] ,_u0_pointer25[15] , _u0_pointer25[14] , _u0_pointer25[13] ,_u0_pointer25[12] , _u0_pointer25[11] , _u0_pointer25[10] ,_u0_pointer25[9] , _u0_pointer25[8] , _u0_pointer25[7] ,_u0_pointer25[6] , _u0_pointer25[5] , _u0_pointer25[4] ,_u0_pointer25[3] , _u0_pointer25[2] , _u0_pointer25[1] ,_u0_pointer25[0] , _u0_pointer25_s[31] , _u0_pointer25_s[30] ,_u0_pointer25_s[29] , _u0_pointer25_s[28] , _u0_pointer25_s[27] ,_u0_pointer25_s[26] , _u0_pointer25_s[25] , _u0_pointer25_s[24] ,_u0_pointer25_s[23] , _u0_pointer25_s[22] , _u0_pointer25_s[21] ,_u0_pointer25_s[20] , _u0_pointer25_s[19] , _u0_pointer25_s[18] ,_u0_pointer25_s[17] , _u0_pointer25_s[16] , _u0_pointer25_s[15] ,_u0_pointer25_s[14] , _u0_pointer25_s[13] , _u0_pointer25_s[12] ,_u0_pointer25_s[11] , _u0_pointer25_s[10] , _u0_pointer25_s[9] ,_u0_pointer25_s[8] , _u0_pointer25_s[7] , _u0_pointer25_s[6] ,_u0_pointer25_s[5] , _u0_pointer25_s[4] , _u0_pointer25_s[3] ,_u0_pointer25_s[2] , _u0_pointer25_s[1] , _u0_pointer25_s[0] ,_u0_ch25_csr[31] , _u0_ch25_csr[30] , _u0_ch25_csr[29] ,_u0_ch25_csr[28] , _u0_ch25_csr[27] , _u0_ch25_csr[26] ,_u0_ch25_csr[25] , _u0_ch25_csr[24] , _u0_ch25_csr[23] ,_u0_ch25_csr[22] , _u0_ch25_csr[21] , _u0_ch25_csr[20] ,_u0_ch25_csr[19] , _u0_ch25_csr[18] , _u0_ch25_csr[17] ,_u0_ch25_csr[16] , _u0_ch25_csr[15] , _u0_ch25_csr[14] ,_u0_ch25_csr[13] , _u0_ch25_csr[12] , _u0_ch25_csr[11] ,_u0_ch25_csr[10] , _u0_ch25_csr[9] , _u0_ch25_csr[8] ,_u0_ch25_csr[7] , _u0_ch25_csr[6] , _u0_ch25_csr[5] ,_u0_ch25_csr[4] , _u0_ch25_csr[3] , _u0_ch25_csr[2] ,_u0_ch25_csr[1] , _u0_ch25_csr[0] , _u0_ch25_txsz[31] ,_u0_ch25_txsz[30] , _u0_ch25_txsz[29] , _u0_ch25_txsz[28] ,_u0_ch25_txsz[27] , _u0_ch25_txsz[26] , _u0_ch25_txsz[25] ,_u0_ch25_txsz[24] , _u0_ch25_txsz[23] , _u0_ch25_txsz[22] ,_u0_ch25_txsz[21] , _u0_ch25_txsz[20] , _u0_ch25_txsz[19] ,_u0_ch25_txsz[18] , _u0_ch25_txsz[17] , _u0_ch25_txsz[16] ,_u0_ch25_txsz[15] , _u0_ch25_txsz[14] , _u0_ch25_txsz[13] ,_u0_ch25_txsz[12] , _u0_ch25_txsz[11] , _u0_ch25_txsz[10] ,_u0_ch25_txsz[9] , _u0_ch25_txsz[8] , _u0_ch25_txsz[7] ,_u0_ch25_txsz[6] , _u0_ch25_txsz[5] , _u0_ch25_txsz[4] ,_u0_ch25_txsz[3] , _u0_ch25_txsz[2] , _u0_ch25_txsz[1] ,_u0_ch25_txsz[0] , _u0_ch25_adr0[31] , _u0_ch25_adr0[30] ,_u0_ch25_adr0[29] , _u0_ch25_adr0[28] , _u0_ch25_adr0[27] ,_u0_ch25_adr0[26] , _u0_ch25_adr0[25] , _u0_ch25_adr0[24] ,_u0_ch25_adr0[23] , _u0_ch25_adr0[22] , _u0_ch25_adr0[21] ,_u0_ch25_adr0[20] , _u0_ch25_adr0[19] , _u0_ch25_adr0[18] ,_u0_ch25_adr0[17] , _u0_ch25_adr0[16] , _u0_ch25_adr0[15] ,_u0_ch25_adr0[14] , _u0_ch25_adr0[13] , _u0_ch25_adr0[12] ,_u0_ch25_adr0[11] , _u0_ch25_adr0[10] , _u0_ch25_adr0[9] ,_u0_ch25_adr0[8] , _u0_ch25_adr0[7] , _u0_ch25_adr0[6] ,_u0_ch25_adr0[5] , _u0_ch25_adr0[4] , _u0_ch25_adr0[3] ,_u0_ch25_adr0[2] , _u0_ch25_adr0[1] , _u0_ch25_adr0[0] ,_u0_ch25_adr1[31] , _u0_ch25_adr1[30] , _u0_ch25_adr1[29] ,_u0_ch25_adr1[28] , _u0_ch25_adr1[27] , _u0_ch25_adr1[26] ,_u0_ch25_adr1[25] , _u0_ch25_adr1[24] , _u0_ch25_adr1[23] ,_u0_ch25_adr1[22] , _u0_ch25_adr1[21] , _u0_ch25_adr1[20] ,_u0_ch25_adr1[19] , _u0_ch25_adr1[18] , _u0_ch25_adr1[17] ,_u0_ch25_adr1[16] , _u0_ch25_adr1[15] , _u0_ch25_adr1[14] ,_u0_ch25_adr1[13] , _u0_ch25_adr1[12] , _u0_ch25_adr1[11] ,_u0_ch25_adr1[10] , _u0_ch25_adr1[9] , _u0_ch25_adr1[8] ,_u0_ch25_adr1[7] , _u0_ch25_adr1[6] , _u0_ch25_adr1[5] ,_u0_ch25_adr1[4] , _u0_ch25_adr1[3] , _u0_ch25_adr1[2] ,_u0_ch25_adr1[1] , _u0_ch25_adr1[0] , _u0_ch25_am0[31] ,_u0_ch25_am0[30] , _u0_ch25_am0[29] , _u0_ch25_am0[28] ,_u0_ch25_am0[27] , _u0_ch25_am0[26] , _u0_ch25_am0[25] ,_u0_ch25_am0[24] , _u0_ch25_am0[23] , _u0_ch25_am0[22] ,_u0_ch25_am0[21] , _u0_ch25_am0[20] , _u0_ch25_am0[19] ,_u0_ch25_am0[18] , _u0_ch25_am0[17] , _u0_ch25_am0[16] ,_u0_ch25_am0[15] , _u0_ch25_am0[14] , _u0_ch25_am0[13] ,_u0_ch25_am0[12] , _u0_ch25_am0[11] , _u0_ch25_am0[10] ,_u0_ch25_am0[9] , _u0_ch25_am0[8] , _u0_ch25_am0[7] ,_u0_ch25_am0[6] , _u0_ch25_am0[5] , _u0_ch25_am0[4] ,_u0_ch25_am0[3] , _u0_ch25_am0[2] , _u0_ch25_am0[1] ,_u0_ch25_am0[0] , _u0_ch25_am1[31] , _u0_ch25_am1[30] ,_u0_ch25_am1[29] , _u0_ch25_am1[28] , _u0_ch25_am1[27] ,_u0_ch25_am1[26] , _u0_ch25_am1[25] , _u0_ch25_am1[24] ,_u0_ch25_am1[23] , _u0_ch25_am1[22] , _u0_ch25_am1[21] ,_u0_ch25_am1[20] , _u0_ch25_am1[19] , _u0_ch25_am1[18] ,_u0_ch25_am1[17] , _u0_ch25_am1[16] , _u0_ch25_am1[15] ,_u0_ch25_am1[14] , _u0_ch25_am1[13] , _u0_ch25_am1[12] ,_u0_ch25_am1[11] , _u0_ch25_am1[10] , _u0_ch25_am1[9] ,_u0_ch25_am1[8] , _u0_ch25_am1[7] , _u0_ch25_am1[6] ,_u0_ch25_am1[5] , _u0_ch25_am1[4] , _u0_ch25_am1[3] ,_u0_ch25_am1[2] , _u0_ch25_am1[1] , _u0_ch25_am1[0] ,_u0_pointer26[31] , _u0_pointer26[30] , _u0_pointer26[29] ,_u0_pointer26[28] , _u0_pointer26[27] , _u0_pointer26[26] ,_u0_pointer26[25] , _u0_pointer26[24] , _u0_pointer26[23] ,_u0_pointer26[22] , _u0_pointer26[21] , _u0_pointer26[20] ,_u0_pointer26[19] , _u0_pointer26[18] , _u0_pointer26[17] ,_u0_pointer26[16] , _u0_pointer26[15] , _u0_pointer26[14] ,_u0_pointer26[13] , _u0_pointer26[12] , _u0_pointer26[11] ,_u0_pointer26[10] , _u0_pointer26[9] , _u0_pointer26[8] ,_u0_pointer26[7] , _u0_pointer26[6] , _u0_pointer26[5] ,_u0_pointer26[4] , _u0_pointer26[3] , _u0_pointer26[2] ,_u0_pointer26[1] , _u0_pointer26[0] , _u0_pointer26_s[31] ,_u0_pointer26_s[30] , _u0_pointer26_s[29] , _u0_pointer26_s[28] ,_u0_pointer26_s[27] , _u0_pointer26_s[26] , _u0_pointer26_s[25] ,_u0_pointer26_s[24] , _u0_pointer26_s[23] , _u0_pointer26_s[22] ,_u0_pointer26_s[21] , _u0_pointer26_s[20] , _u0_pointer26_s[19] ,_u0_pointer26_s[18] , _u0_pointer26_s[17] , _u0_pointer26_s[16] ,_u0_pointer26_s[15] , _u0_pointer26_s[14] , _u0_pointer26_s[13] ,_u0_pointer26_s[12] , _u0_pointer26_s[11] , _u0_pointer26_s[10] ,_u0_pointer26_s[9] , _u0_pointer26_s[8] , _u0_pointer26_s[7] ,_u0_pointer26_s[6] , _u0_pointer26_s[5] , _u0_pointer26_s[4] ,_u0_pointer26_s[3] , _u0_pointer26_s[2] , _u0_pointer26_s[1] ,_u0_pointer26_s[0] , _u0_ch26_csr[31] , _u0_ch26_csr[30] ,_u0_ch26_csr[29] , _u0_ch26_csr[28] , _u0_ch26_csr[27] ,_u0_ch26_csr[26] , _u0_ch26_csr[25] , _u0_ch26_csr[24] ,_u0_ch26_csr[23] , _u0_ch26_csr[22] , _u0_ch26_csr[21] ,_u0_ch26_csr[20] , _u0_ch26_csr[19] , _u0_ch26_csr[18] ,_u0_ch26_csr[17] , _u0_ch26_csr[16] , _u0_ch26_csr[15] ,_u0_ch26_csr[14] , _u0_ch26_csr[13] , _u0_ch26_csr[12] ,_u0_ch26_csr[11] , _u0_ch26_csr[10] , _u0_ch26_csr[9] ,_u0_ch26_csr[8] , _u0_ch26_csr[7] , _u0_ch26_csr[6] ,_u0_ch26_csr[5] , _u0_ch26_csr[4] , _u0_ch26_csr[3] ,_u0_ch26_csr[2] , _u0_ch26_csr[1] , _u0_ch26_csr[0] ,_u0_ch26_txsz[31] , _u0_ch26_txsz[30] , _u0_ch26_txsz[29] ,_u0_ch26_txsz[28] , _u0_ch26_txsz[27] , _u0_ch26_txsz[26] ,_u0_ch26_txsz[25] , _u0_ch26_txsz[24] , _u0_ch26_txsz[23] ,_u0_ch26_txsz[22] , _u0_ch26_txsz[21] , _u0_ch26_txsz[20] ,_u0_ch26_txsz[19] , _u0_ch26_txsz[18] , _u0_ch26_txsz[17] ,_u0_ch26_txsz[16] , _u0_ch26_txsz[15] , _u0_ch26_txsz[14] ,_u0_ch26_txsz[13] , _u0_ch26_txsz[12] , _u0_ch26_txsz[11] ,_u0_ch26_txsz[10] , _u0_ch26_txsz[9] , _u0_ch26_txsz[8] ,_u0_ch26_txsz[7] , _u0_ch26_txsz[6] , _u0_ch26_txsz[5] ,_u0_ch26_txsz[4] , _u0_ch26_txsz[3] , _u0_ch26_txsz[2] ,_u0_ch26_txsz[1] , _u0_ch26_txsz[0] , _u0_ch26_adr0[31] ,_u0_ch26_adr0[30] , _u0_ch26_adr0[29] , _u0_ch26_adr0[28] ,_u0_ch26_adr0[27] , _u0_ch26_adr0[26] , _u0_ch26_adr0[25] ,_u0_ch26_adr0[24] , _u0_ch26_adr0[23] , _u0_ch26_adr0[22] ,_u0_ch26_adr0[21] , _u0_ch26_adr0[20] , _u0_ch26_adr0[19] ,_u0_ch26_adr0[18] , _u0_ch26_adr0[17] , _u0_ch26_adr0[16] ,_u0_ch26_adr0[15] , _u0_ch26_adr0[14] , _u0_ch26_adr0[13] ,_u0_ch26_adr0[12] , _u0_ch26_adr0[11] , _u0_ch26_adr0[10] ,_u0_ch26_adr0[9] , _u0_ch26_adr0[8] , _u0_ch26_adr0[7] ,_u0_ch26_adr0[6] , _u0_ch26_adr0[5] , _u0_ch26_adr0[4] ,_u0_ch26_adr0[3] , _u0_ch26_adr0[2] , _u0_ch26_adr0[1] ,_u0_ch26_adr0[0] , _u0_ch26_adr1[31] , _u0_ch26_adr1[30] ,_u0_ch26_adr1[29] , _u0_ch26_adr1[28] , _u0_ch26_adr1[27] ,_u0_ch26_adr1[26] , _u0_ch26_adr1[25] , _u0_ch26_adr1[24] ,_u0_ch26_adr1[23] , _u0_ch26_adr1[22] , _u0_ch26_adr1[21] ,_u0_ch26_adr1[20] , _u0_ch26_adr1[19] , _u0_ch26_adr1[18] ,_u0_ch26_adr1[17] , _u0_ch26_adr1[16] , _u0_ch26_adr1[15] ,_u0_ch26_adr1[14] , _u0_ch26_adr1[13] , _u0_ch26_adr1[12] ,_u0_ch26_adr1[11] , _u0_ch26_adr1[10] , _u0_ch26_adr1[9] ,_u0_ch26_adr1[8] , _u0_ch26_adr1[7] , _u0_ch26_adr1[6] ,_u0_ch26_adr1[5] , _u0_ch26_adr1[4] , _u0_ch26_adr1[3] ,_u0_ch26_adr1[2] , _u0_ch26_adr1[1] , _u0_ch26_adr1[0] ,_u0_ch26_am0[31] , _u0_ch26_am0[30] , _u0_ch26_am0[29] ,_u0_ch26_am0[28] , _u0_ch26_am0[27] , _u0_ch26_am0[26] ,_u0_ch26_am0[25] , _u0_ch26_am0[24] , _u0_ch26_am0[23] ,_u0_ch26_am0[22] , _u0_ch26_am0[21] , _u0_ch26_am0[20] ,_u0_ch26_am0[19] , _u0_ch26_am0[18] , _u0_ch26_am0[17] ,_u0_ch26_am0[16] , _u0_ch26_am0[15] , _u0_ch26_am0[14] ,_u0_ch26_am0[13] , _u0_ch26_am0[12] , _u0_ch26_am0[11] ,_u0_ch26_am0[10] , _u0_ch26_am0[9] , _u0_ch26_am0[8] ,_u0_ch26_am0[7] , _u0_ch26_am0[6] , _u0_ch26_am0[5] ,_u0_ch26_am0[4] , _u0_ch26_am0[3] , _u0_ch26_am0[2] ,_u0_ch26_am0[1] , _u0_ch26_am0[0] , _u0_ch26_am1[31] ,_u0_ch26_am1[30] , _u0_ch26_am1[29] , _u0_ch26_am1[28] ,_u0_ch26_am1[27] , _u0_ch26_am1[26] , _u0_ch26_am1[25] ,_u0_ch26_am1[24] , _u0_ch26_am1[23] , _u0_ch26_am1[22] ,_u0_ch26_am1[21] , _u0_ch26_am1[20] , _u0_ch26_am1[19] ,_u0_ch26_am1[18] , _u0_ch26_am1[17] , _u0_ch26_am1[16] ,_u0_ch26_am1[15] , _u0_ch26_am1[14] , _u0_ch26_am1[13] ,_u0_ch26_am1[12] , _u0_ch26_am1[11] , _u0_ch26_am1[10] ,_u0_ch26_am1[9] , _u0_ch26_am1[8] , _u0_ch26_am1[7] ,_u0_ch26_am1[6] , _u0_ch26_am1[5] , _u0_ch26_am1[4] ,_u0_ch26_am1[3] , _u0_ch26_am1[2] , _u0_ch26_am1[1] ,_u0_ch26_am1[0] , _u0_pointer27[31] , _u0_pointer27[30] ,_u0_pointer27[29] , _u0_pointer27[28] , _u0_pointer27[27] ,_u0_pointer27[26] , _u0_pointer27[25] , _u0_pointer27[24] ,_u0_pointer27[23] , _u0_pointer27[22] , _u0_pointer27[21] ,_u0_pointer27[20] , _u0_pointer27[19] , _u0_pointer27[18] ,_u0_pointer27[17] , _u0_pointer27[16] , _u0_pointer27[15] ,_u0_pointer27[14] , _u0_pointer27[13] , _u0_pointer27[12] ,_u0_pointer27[11] , _u0_pointer27[10] , _u0_pointer27[9] ,_u0_pointer27[8] , _u0_pointer27[7] , _u0_pointer27[6] ,_u0_pointer27[5] , _u0_pointer27[4] , _u0_pointer27[3] ,_u0_pointer27[2] , _u0_pointer27[1] , _u0_pointer27[0] ,_u0_pointer27_s[31] , _u0_pointer27_s[30] , _u0_pointer27_s[29] ,_u0_pointer27_s[28] , _u0_pointer27_s[27] , _u0_pointer27_s[26] ,_u0_pointer27_s[25] , _u0_pointer27_s[24] , _u0_pointer27_s[23] ,_u0_pointer27_s[22] , _u0_pointer27_s[21] , _u0_pointer27_s[20] ,_u0_pointer27_s[19] , _u0_pointer27_s[18] , _u0_pointer27_s[17] ,_u0_pointer27_s[16] , _u0_pointer27_s[15] , _u0_pointer27_s[14] ,_u0_pointer27_s[13] , _u0_pointer27_s[12] , _u0_pointer27_s[11] ,_u0_pointer27_s[10] , _u0_pointer27_s[9] , _u0_pointer27_s[8] ,_u0_pointer27_s[7] , _u0_pointer27_s[6] , _u0_pointer27_s[5] ,_u0_pointer27_s[4] , _u0_pointer27_s[3] , _u0_pointer27_s[2] ,_u0_pointer27_s[1] , _u0_pointer27_s[0] , _u0_ch27_csr[31] ,_u0_ch27_csr[30] , _u0_ch27_csr[29] , _u0_ch27_csr[28] ,_u0_ch27_csr[27] , _u0_ch27_csr[26] , _u0_ch27_csr[25] ,_u0_ch27_csr[24] , _u0_ch27_csr[23] , _u0_ch27_csr[22] ,_u0_ch27_csr[21] , _u0_ch27_csr[20] , _u0_ch27_csr[19] ,_u0_ch27_csr[18] , _u0_ch27_csr[17] , _u0_ch27_csr[16] ,_u0_ch27_csr[15] , _u0_ch27_csr[14] , _u0_ch27_csr[13] ,_u0_ch27_csr[12] , _u0_ch27_csr[11] , _u0_ch27_csr[10] ,_u0_ch27_csr[9] , _u0_ch27_csr[8] , _u0_ch27_csr[7] ,_u0_ch27_csr[6] , _u0_ch27_csr[5] , _u0_ch27_csr[4] ,_u0_ch27_csr[3] , _u0_ch27_csr[2] , _u0_ch27_csr[1] ,_u0_ch27_csr[0] , _u0_ch27_txsz[31] , _u0_ch27_txsz[30] ,_u0_ch27_txsz[29] , _u0_ch27_txsz[28] , _u0_ch27_txsz[27] ,_u0_ch27_txsz[26] , _u0_ch27_txsz[25] , _u0_ch27_txsz[24] ,_u0_ch27_txsz[23] , _u0_ch27_txsz[22] , _u0_ch27_txsz[21] ,_u0_ch27_txsz[20] , _u0_ch27_txsz[19] , _u0_ch27_txsz[18] ,_u0_ch27_txsz[17] , _u0_ch27_txsz[16] , _u0_ch27_txsz[15] ,_u0_ch27_txsz[14] , _u0_ch27_txsz[13] , _u0_ch27_txsz[12] ,_u0_ch27_txsz[11] , _u0_ch27_txsz[10] , _u0_ch27_txsz[9] ,_u0_ch27_txsz[8] , _u0_ch27_txsz[7] , _u0_ch27_txsz[6] ,_u0_ch27_txsz[5] , _u0_ch27_txsz[4] , _u0_ch27_txsz[3] ,_u0_ch27_txsz[2] , _u0_ch27_txsz[1] , _u0_ch27_txsz[0] ,_u0_ch27_adr0[31] , _u0_ch27_adr0[30] , _u0_ch27_adr0[29] ,_u0_ch27_adr0[28] , _u0_ch27_adr0[27] , _u0_ch27_adr0[26] ,_u0_ch27_adr0[25] , _u0_ch27_adr0[24] , _u0_ch27_adr0[23] ,_u0_ch27_adr0[22] , _u0_ch27_adr0[21] , _u0_ch27_adr0[20] ,_u0_ch27_adr0[19] , _u0_ch27_adr0[18] , _u0_ch27_adr0[17] ,_u0_ch27_adr0[16] , _u0_ch27_adr0[15] , _u0_ch27_adr0[14] ,_u0_ch27_adr0[13] , _u0_ch27_adr0[12] , _u0_ch27_adr0[11] ,_u0_ch27_adr0[10] , _u0_ch27_adr0[9] , _u0_ch27_adr0[8] ,_u0_ch27_adr0[7] , _u0_ch27_adr0[6] , _u0_ch27_adr0[5] ,_u0_ch27_adr0[4] , _u0_ch27_adr0[3] , _u0_ch27_adr0[2] ,_u0_ch27_adr0[1] , _u0_ch27_adr0[0] , _u0_ch27_adr1[31] ,_u0_ch27_adr1[30] , _u0_ch27_adr1[29] , _u0_ch27_adr1[28] ,_u0_ch27_adr1[27] , _u0_ch27_adr1[26] , _u0_ch27_adr1[25] ,_u0_ch27_adr1[24] , _u0_ch27_adr1[23] , _u0_ch27_adr1[22] ,_u0_ch27_adr1[21] , _u0_ch27_adr1[20] , _u0_ch27_adr1[19] ,_u0_ch27_adr1[18] , _u0_ch27_adr1[17] , _u0_ch27_adr1[16] ,_u0_ch27_adr1[15] , _u0_ch27_adr1[14] , _u0_ch27_adr1[13] ,_u0_ch27_adr1[12] , _u0_ch27_adr1[11] , _u0_ch27_adr1[10] ,_u0_ch27_adr1[9] , _u0_ch27_adr1[8] , _u0_ch27_adr1[7] ,_u0_ch27_adr1[6] , _u0_ch27_adr1[5] , _u0_ch27_adr1[4] ,_u0_ch27_adr1[3] , _u0_ch27_adr1[2] , _u0_ch27_adr1[1] ,_u0_ch27_adr1[0] , _u0_ch27_am0[31] , _u0_ch27_am0[30] ,_u0_ch27_am0[29] , _u0_ch27_am0[28] , _u0_ch27_am0[27] ,_u0_ch27_am0[26] , _u0_ch27_am0[25] , _u0_ch27_am0[24] ,_u0_ch27_am0[23] , _u0_ch27_am0[22] , _u0_ch27_am0[21] ,_u0_ch27_am0[20] , _u0_ch27_am0[19] , _u0_ch27_am0[18] ,_u0_ch27_am0[17] , _u0_ch27_am0[16] , _u0_ch27_am0[15] ,_u0_ch27_am0[14] , _u0_ch27_am0[13] , _u0_ch27_am0[12] ,_u0_ch27_am0[11] , _u0_ch27_am0[10] , _u0_ch27_am0[9] ,_u0_ch27_am0[8] , _u0_ch27_am0[7] , _u0_ch27_am0[6] ,_u0_ch27_am0[5] , _u0_ch27_am0[4] , _u0_ch27_am0[3] ,_u0_ch27_am0[2] , _u0_ch27_am0[1] , _u0_ch27_am0[0] ,_u0_ch27_am1[31] , _u0_ch27_am1[30] , _u0_ch27_am1[29] ,_u0_ch27_am1[28] , _u0_ch27_am1[27] , _u0_ch27_am1[26] ,_u0_ch27_am1[25] , _u0_ch27_am1[24] , _u0_ch27_am1[23] ,_u0_ch27_am1[22] , _u0_ch27_am1[21] , _u0_ch27_am1[20] ,_u0_ch27_am1[19] , _u0_ch27_am1[18] , _u0_ch27_am1[17] ,_u0_ch27_am1[16] , _u0_ch27_am1[15] , _u0_ch27_am1[14] ,_u0_ch27_am1[13] , _u0_ch27_am1[12] , _u0_ch27_am1[11] ,_u0_ch27_am1[10] , _u0_ch27_am1[9] , _u0_ch27_am1[8] ,_u0_ch27_am1[7] , _u0_ch27_am1[6] , _u0_ch27_am1[5] ,_u0_ch27_am1[4] , _u0_ch27_am1[3] , _u0_ch27_am1[2] ,_u0_ch27_am1[1] , _u0_ch27_am1[0] , _u0_pointer28[31] ,_u0_pointer28[30] , _u0_pointer28[29] , _u0_pointer28[28] ,_u0_pointer28[27] , _u0_pointer28[26] , _u0_pointer28[25] ,_u0_pointer28[24] , _u0_pointer28[23] , _u0_pointer28[22] ,_u0_pointer28[21] , _u0_pointer28[20] , _u0_pointer28[19] ,_u0_pointer28[18] , _u0_pointer28[17] , _u0_pointer28[16] ,_u0_pointer28[15] , _u0_pointer28[14] , _u0_pointer28[13] ,_u0_pointer28[12] , _u0_pointer28[11] , _u0_pointer28[10] ,_u0_pointer28[9] , _u0_pointer28[8] , _u0_pointer28[7] ,_u0_pointer28[6] , _u0_pointer28[5] , _u0_pointer28[4] ,_u0_pointer28[3] , _u0_pointer28[2] , _u0_pointer28[1] ,_u0_pointer28[0] , _u0_pointer28_s[31] , _u0_pointer28_s[30] ,_u0_pointer28_s[29] , _u0_pointer28_s[28] , _u0_pointer28_s[27] ,_u0_pointer28_s[26] , _u0_pointer28_s[25] , _u0_pointer28_s[24] ,_u0_pointer28_s[23] , _u0_pointer28_s[22] , _u0_pointer28_s[21] ,_u0_pointer28_s[20] , _u0_pointer28_s[19] , _u0_pointer28_s[18] ,_u0_pointer28_s[17] , _u0_pointer28_s[16] , _u0_pointer28_s[15] ,_u0_pointer28_s[14] , _u0_pointer28_s[13] , _u0_pointer28_s[12] ,_u0_pointer28_s[11] , _u0_pointer28_s[10] , _u0_pointer28_s[9] ,_u0_pointer28_s[8] , _u0_pointer28_s[7] , _u0_pointer28_s[6] ,_u0_pointer28_s[5] , _u0_pointer28_s[4] , _u0_pointer28_s[3] ,_u0_pointer28_s[2] , _u0_pointer28_s[1] , _u0_pointer28_s[0] ,_u0_ch28_csr[31] , _u0_ch28_csr[30] , _u0_ch28_csr[29] ,_u0_ch28_csr[28] , _u0_ch28_csr[27] , _u0_ch28_csr[26] ,_u0_ch28_csr[25] , _u0_ch28_csr[24] , _u0_ch28_csr[23] ,_u0_ch28_csr[22] , _u0_ch28_csr[21] , _u0_ch28_csr[20] ,_u0_ch28_csr[19] , _u0_ch28_csr[18] , _u0_ch28_csr[17] ,_u0_ch28_csr[16] , _u0_ch28_csr[15] , _u0_ch28_csr[14] ,_u0_ch28_csr[13] , _u0_ch28_csr[12] , _u0_ch28_csr[11] ,_u0_ch28_csr[10] , _u0_ch28_csr[9] , _u0_ch28_csr[8] ,_u0_ch28_csr[7] , _u0_ch28_csr[6] , _u0_ch28_csr[5] ,_u0_ch28_csr[4] , _u0_ch28_csr[3] , _u0_ch28_csr[2] ,_u0_ch28_csr[1] , _u0_ch28_csr[0] , _u0_ch28_txsz[31] ,_u0_ch28_txsz[30] , _u0_ch28_txsz[29] , _u0_ch28_txsz[28] ,_u0_ch28_txsz[27] , _u0_ch28_txsz[26] , _u0_ch28_txsz[25] ,_u0_ch28_txsz[24] , _u0_ch28_txsz[23] , _u0_ch28_txsz[22] ,_u0_ch28_txsz[21] , _u0_ch28_txsz[20] , _u0_ch28_txsz[19] ,_u0_ch28_txsz[18] , _u0_ch28_txsz[17] , _u0_ch28_txsz[16] ,_u0_ch28_txsz[15] , _u0_ch28_txsz[14] , _u0_ch28_txsz[13] ,_u0_ch28_txsz[12] , _u0_ch28_txsz[11] , _u0_ch28_txsz[10] ,_u0_ch28_txsz[9] , _u0_ch28_txsz[8] , _u0_ch28_txsz[7] ,_u0_ch28_txsz[6] , _u0_ch28_txsz[5] , _u0_ch28_txsz[4] ,_u0_ch28_txsz[3] , _u0_ch28_txsz[2] , _u0_ch28_txsz[1] ,_u0_ch28_txsz[0] , _u0_ch28_adr0[31] , _u0_ch28_adr0[30] ,_u0_ch28_adr0[29] , _u0_ch28_adr0[28] , _u0_ch28_adr0[27] ,_u0_ch28_adr0[26] , _u0_ch28_adr0[25] , _u0_ch28_adr0[24] ,_u0_ch28_adr0[23] , _u0_ch28_adr0[22] , _u0_ch28_adr0[21] ,_u0_ch28_adr0[20] , _u0_ch28_adr0[19] , _u0_ch28_adr0[18] ,_u0_ch28_adr0[17] , _u0_ch28_adr0[16] , _u0_ch28_adr0[15] ,_u0_ch28_adr0[14] , _u0_ch28_adr0[13] , _u0_ch28_adr0[12] ,_u0_ch28_adr0[11] , _u0_ch28_adr0[10] , _u0_ch28_adr0[9] ,_u0_ch28_adr0[8] , _u0_ch28_adr0[7] , _u0_ch28_adr0[6] ,_u0_ch28_adr0[5] , _u0_ch28_adr0[4] , _u0_ch28_adr0[3] ,_u0_ch28_adr0[2] , _u0_ch28_adr0[1] , _u0_ch28_adr0[0] ,_u0_ch28_adr1[31] , _u0_ch28_adr1[30] , _u0_ch28_adr1[29] ,_u0_ch28_adr1[28] , _u0_ch28_adr1[27] , _u0_ch28_adr1[26] ,_u0_ch28_adr1[25] , _u0_ch28_adr1[24] , _u0_ch28_adr1[23] ,_u0_ch28_adr1[22] , _u0_ch28_adr1[21] , _u0_ch28_adr1[20] ,_u0_ch28_adr1[19] , _u0_ch28_adr1[18] , _u0_ch28_adr1[17] ,_u0_ch28_adr1[16] , _u0_ch28_adr1[15] , _u0_ch28_adr1[14] ,_u0_ch28_adr1[13] , _u0_ch28_adr1[12] , _u0_ch28_adr1[11] ,_u0_ch28_adr1[10] , _u0_ch28_adr1[9] , _u0_ch28_adr1[8] ,_u0_ch28_adr1[7] , _u0_ch28_adr1[6] , _u0_ch28_adr1[5] ,_u0_ch28_adr1[4] , _u0_ch28_adr1[3] , _u0_ch28_adr1[2] ,_u0_ch28_adr1[1] , _u0_ch28_adr1[0] , _u0_ch28_am0[31] ,_u0_ch28_am0[30] , _u0_ch28_am0[29] , _u0_ch28_am0[28] ,_u0_ch28_am0[27] , _u0_ch28_am0[26] , _u0_ch28_am0[25] ,_u0_ch28_am0[24] , _u0_ch28_am0[23] , _u0_ch28_am0[22] ,_u0_ch28_am0[21] , _u0_ch28_am0[20] , _u0_ch28_am0[19] ,_u0_ch28_am0[18] , _u0_ch28_am0[17] , _u0_ch28_am0[16] ,_u0_ch28_am0[15] , _u0_ch28_am0[14] , _u0_ch28_am0[13] ,_u0_ch28_am0[12] , _u0_ch28_am0[11] , _u0_ch28_am0[10] ,_u0_ch28_am0[9] , _u0_ch28_am0[8] , _u0_ch28_am0[7] ,_u0_ch28_am0[6] , _u0_ch28_am0[5] , _u0_ch28_am0[4] ,_u0_ch28_am0[3] , _u0_ch28_am0[2] , _u0_ch28_am0[1] ,_u0_ch28_am0[0] , _u0_ch28_am1[31] , _u0_ch28_am1[30] ,_u0_ch28_am1[29] , _u0_ch28_am1[28] , _u0_ch28_am1[27] ,_u0_ch28_am1[26] , _u0_ch28_am1[25] , _u0_ch28_am1[24] ,_u0_ch28_am1[23] , _u0_ch28_am1[22] , _u0_ch28_am1[21] ,_u0_ch28_am1[20] , _u0_ch28_am1[19] , _u0_ch28_am1[18] ,_u0_ch28_am1[17] , _u0_ch28_am1[16] , _u0_ch28_am1[15] ,_u0_ch28_am1[14] , _u0_ch28_am1[13] , _u0_ch28_am1[12] ,_u0_ch28_am1[11] , _u0_ch28_am1[10] , _u0_ch28_am1[9] ,_u0_ch28_am1[8] , _u0_ch28_am1[7] , _u0_ch28_am1[6] ,_u0_ch28_am1[5] , _u0_ch28_am1[4] , _u0_ch28_am1[3] ,_u0_ch28_am1[2] , _u0_ch28_am1[1] , _u0_ch28_am1[0] ,_u0_pointer29[31] , _u0_pointer29[30] , _u0_pointer29[29] ,_u0_pointer29[28] , _u0_pointer29[27] , _u0_pointer29[26] ,_u0_pointer29[25] , _u0_pointer29[24] , _u0_pointer29[23] ,_u0_pointer29[22] , _u0_pointer29[21] , _u0_pointer29[20] ,_u0_pointer29[19] , _u0_pointer29[18] , _u0_pointer29[17] ,_u0_pointer29[16] , _u0_pointer29[15] , _u0_pointer29[14] ,_u0_pointer29[13] , _u0_pointer29[12] , _u0_pointer29[11] ,_u0_pointer29[10] , _u0_pointer29[9] , _u0_pointer29[8] ,_u0_pointer29[7] , _u0_pointer29[6] , _u0_pointer29[5] ,_u0_pointer29[4] , _u0_pointer29[3] , _u0_pointer29[2] ,_u0_pointer29[1] , _u0_pointer29[0] , _u0_pointer29_s[31] ,_u0_pointer29_s[30] , _u0_pointer29_s[29] , _u0_pointer29_s[28] ,_u0_pointer29_s[27] , _u0_pointer29_s[26] , _u0_pointer29_s[25] ,_u0_pointer29_s[24] , _u0_pointer29_s[23] , _u0_pointer29_s[22] ,_u0_pointer29_s[21] , _u0_pointer29_s[20] , _u0_pointer29_s[19] ,_u0_pointer29_s[18] , _u0_pointer29_s[17] , _u0_pointer29_s[16] ,_u0_pointer29_s[15] , _u0_pointer29_s[14] , _u0_pointer29_s[13] ,_u0_pointer29_s[12] , _u0_pointer29_s[11] , _u0_pointer29_s[10] ,_u0_pointer29_s[9] , _u0_pointer29_s[8] , _u0_pointer29_s[7] ,_u0_pointer29_s[6] , _u0_pointer29_s[5] , _u0_pointer29_s[4] ,_u0_pointer29_s[3] , _u0_pointer29_s[2] , _u0_pointer29_s[1] ,_u0_pointer29_s[0] , _u0_ch29_csr[31] , _u0_ch29_csr[30] ,_u0_ch29_csr[29] , _u0_ch29_csr[28] , _u0_ch29_csr[27] ,_u0_ch29_csr[26] , _u0_ch29_csr[25] , _u0_ch29_csr[24] ,_u0_ch29_csr[23] , _u0_ch29_csr[22] , _u0_ch29_csr[21] ,_u0_ch29_csr[20] , _u0_ch29_csr[19] , _u0_ch29_csr[18] ,_u0_ch29_csr[17] , _u0_ch29_csr[16] , _u0_ch29_csr[15] ,_u0_ch29_csr[14] , _u0_ch29_csr[13] , _u0_ch29_csr[12] ,_u0_ch29_csr[11] , _u0_ch29_csr[10] , _u0_ch29_csr[9] ,_u0_ch29_csr[8] , _u0_ch29_csr[7] , _u0_ch29_csr[6] ,_u0_ch29_csr[5] , _u0_ch29_csr[4] , _u0_ch29_csr[3] ,_u0_ch29_csr[2] , _u0_ch29_csr[1] , _u0_ch29_csr[0] ,_u0_ch29_txsz[31] , _u0_ch29_txsz[30] , _u0_ch29_txsz[29] ,_u0_ch29_txsz[28] , _u0_ch29_txsz[27] , _u0_ch29_txsz[26] ,_u0_ch29_txsz[25] , _u0_ch29_txsz[24] , _u0_ch29_txsz[23] ,_u0_ch29_txsz[22] , _u0_ch29_txsz[21] , _u0_ch29_txsz[20] ,_u0_ch29_txsz[19] , _u0_ch29_txsz[18] , _u0_ch29_txsz[17] ,_u0_ch29_txsz[16] , _u0_ch29_txsz[15] , _u0_ch29_txsz[14] ,_u0_ch29_txsz[13] , _u0_ch29_txsz[12] , _u0_ch29_txsz[11] ,_u0_ch29_txsz[10] , _u0_ch29_txsz[9] , _u0_ch29_txsz[8] ,_u0_ch29_txsz[7] , _u0_ch29_txsz[6] , _u0_ch29_txsz[5] ,_u0_ch29_txsz[4] , _u0_ch29_txsz[3] , _u0_ch29_txsz[2] ,_u0_ch29_txsz[1] , _u0_ch29_txsz[0] , _u0_ch29_adr0[31] ,_u0_ch29_adr0[30] , _u0_ch29_adr0[29] , _u0_ch29_adr0[28] ,_u0_ch29_adr0[27] , _u0_ch29_adr0[26] , _u0_ch29_adr0[25] ,_u0_ch29_adr0[24] , _u0_ch29_adr0[23] , _u0_ch29_adr0[22] ,_u0_ch29_adr0[21] , _u0_ch29_adr0[20] , _u0_ch29_adr0[19] ,_u0_ch29_adr0[18] , _u0_ch29_adr0[17] , _u0_ch29_adr0[16] ,_u0_ch29_adr0[15] , _u0_ch29_adr0[14] , _u0_ch29_adr0[13] ,_u0_ch29_adr0[12] , _u0_ch29_adr0[11] , _u0_ch29_adr0[10] ,_u0_ch29_adr0[9] , _u0_ch29_adr0[8] , _u0_ch29_adr0[7] ,_u0_ch29_adr0[6] , _u0_ch29_adr0[5] , _u0_ch29_adr0[4] ,_u0_ch29_adr0[3] , _u0_ch29_adr0[2] , _u0_ch29_adr0[1] ,_u0_ch29_adr0[0] , _u0_ch29_adr1[31] , _u0_ch29_adr1[30] ,_u0_ch29_adr1[29] , _u0_ch29_adr1[28] , _u0_ch29_adr1[27] ,_u0_ch29_adr1[26] , _u0_ch29_adr1[25] , _u0_ch29_adr1[24] ,_u0_ch29_adr1[23] , _u0_ch29_adr1[22] , _u0_ch29_adr1[21] ,_u0_ch29_adr1[20] , _u0_ch29_adr1[19] , _u0_ch29_adr1[18] ,_u0_ch29_adr1[17] , _u0_ch29_adr1[16] , _u0_ch29_adr1[15] ,_u0_ch29_adr1[14] , _u0_ch29_adr1[13] , _u0_ch29_adr1[12] ,_u0_ch29_adr1[11] , _u0_ch29_adr1[10] , _u0_ch29_adr1[9] ,_u0_ch29_adr1[8] , _u0_ch29_adr1[7] , _u0_ch29_adr1[6] ,_u0_ch29_adr1[5] , _u0_ch29_adr1[4] , _u0_ch29_adr1[3] ,_u0_ch29_adr1[2] , _u0_ch29_adr1[1] , _u0_ch29_adr1[0] ,_u0_ch29_am0[31] , _u0_ch29_am0[30] , _u0_ch29_am0[29] ,_u0_ch29_am0[28] , _u0_ch29_am0[27] , _u0_ch29_am0[26] ,_u0_ch29_am0[25] , _u0_ch29_am0[24] , _u0_ch29_am0[23] ,_u0_ch29_am0[22] , _u0_ch29_am0[21] , _u0_ch29_am0[20] ,_u0_ch29_am0[19] , _u0_ch29_am0[18] , _u0_ch29_am0[17] ,_u0_ch29_am0[16] , _u0_ch29_am0[15] , _u0_ch29_am0[14] ,_u0_ch29_am0[13] , _u0_ch29_am0[12] , _u0_ch29_am0[11] ,_u0_ch29_am0[10] , _u0_ch29_am0[9] , _u0_ch29_am0[8] ,_u0_ch29_am0[7] , _u0_ch29_am0[6] , _u0_ch29_am0[5] ,_u0_ch29_am0[4] , _u0_ch29_am0[3] , _u0_ch29_am0[2] ,_u0_ch29_am0[1] , _u0_ch29_am0[0] , _u0_ch29_am1[31] ,_u0_ch29_am1[30] , _u0_ch29_am1[29] , _u0_ch29_am1[28] ,_u0_ch29_am1[27] , _u0_ch29_am1[26] , _u0_ch29_am1[25] ,_u0_ch29_am1[24] , _u0_ch29_am1[23] , _u0_ch29_am1[22] ,_u0_ch29_am1[21] , _u0_ch29_am1[20] , _u0_ch29_am1[19] ,_u0_ch29_am1[18] , _u0_ch29_am1[17] , _u0_ch29_am1[16] ,_u0_ch29_am1[15] , _u0_ch29_am1[14] , _u0_ch29_am1[13] ,_u0_ch29_am1[12] , _u0_ch29_am1[11] , _u0_ch29_am1[10] ,_u0_ch29_am1[9] , _u0_ch29_am1[8] , _u0_ch29_am1[7] ,_u0_ch29_am1[6] , _u0_ch29_am1[5] , _u0_ch29_am1[4] ,_u0_ch29_am1[3] , _u0_ch29_am1[2] , _u0_ch29_am1[1] ,_u0_ch29_am1[0] , _u0_pointer30[31] , _u0_pointer30[30] ,_u0_pointer30[29] , _u0_pointer30[28] , _u0_pointer30[27] ,_u0_pointer30[26] , _u0_pointer30[25] , _u0_pointer30[24] ,_u0_pointer30[23] , _u0_pointer30[22] , _u0_pointer30[21] ,_u0_pointer30[20] , _u0_pointer30[19] , _u0_pointer30[18] ,_u0_pointer30[17] , _u0_pointer30[16] , _u0_pointer30[15] ,_u0_pointer30[14] , _u0_pointer30[13] , _u0_pointer30[12] ,_u0_pointer30[11] , _u0_pointer30[10] , _u0_pointer30[9] ,_u0_pointer30[8] , _u0_pointer30[7] , _u0_pointer30[6] ,_u0_pointer30[5] , _u0_pointer30[4] , _u0_pointer30[3] ,_u0_pointer30[2] , _u0_pointer30[1] , _u0_pointer30[0] ,_u0_pointer30_s[31] , _u0_pointer30_s[30] , _u0_pointer30_s[29] ,_u0_pointer30_s[28] , _u0_pointer30_s[27] , _u0_pointer30_s[26] ,_u0_pointer30_s[25] , _u0_pointer30_s[24] , _u0_pointer30_s[23] ,_u0_pointer30_s[22] , _u0_pointer30_s[21] , _u0_pointer30_s[20] ,_u0_pointer30_s[19] , _u0_pointer30_s[18] , _u0_pointer30_s[17] ,_u0_pointer30_s[16] , _u0_pointer30_s[15] , _u0_pointer30_s[14] ,_u0_pointer30_s[13] , _u0_pointer30_s[12] , _u0_pointer30_s[11] ,_u0_pointer30_s[10] , _u0_pointer30_s[9] , _u0_pointer30_s[8] ,_u0_pointer30_s[7] , _u0_pointer30_s[6] , _u0_pointer30_s[5] ,_u0_pointer30_s[4] , _u0_pointer30_s[3] , _u0_pointer30_s[2] ,_u0_pointer30_s[1] , _u0_pointer30_s[0] , _u0_ch30_csr[31] ,_u0_ch30_csr[30] , _u0_ch30_csr[29] , _u0_ch30_csr[28] ,_u0_ch30_csr[27] , _u0_ch30_csr[26] , _u0_ch30_csr[25] ,_u0_ch30_csr[24] , _u0_ch30_csr[23] , _u0_ch30_csr[22] ,_u0_ch30_csr[21] , _u0_ch30_csr[20] , _u0_ch30_csr[19] ,_u0_ch30_csr[18] , _u0_ch30_csr[17] , _u0_ch30_csr[16] ,_u0_ch30_csr[15] , _u0_ch30_csr[14] , _u0_ch30_csr[13] ,_u0_ch30_csr[12] , _u0_ch30_csr[11] , _u0_ch30_csr[10] ,_u0_ch30_csr[9] , _u0_ch30_csr[8] , _u0_ch30_csr[7] ,_u0_ch30_csr[6] , _u0_ch30_csr[5] , _u0_ch30_csr[4] ,_u0_ch30_csr[3] , _u0_ch30_csr[2] , _u0_ch30_csr[1] ,_u0_ch30_csr[0] , _u0_ch30_txsz[31] , _u0_ch30_txsz[30] ,_u0_ch30_txsz[29] , _u0_ch30_txsz[28] , _u0_ch30_txsz[27] ,_u0_ch30_txsz[26] , _u0_ch30_txsz[25] , _u0_ch30_txsz[24] ,_u0_ch30_txsz[23] , _u0_ch30_txsz[22] , _u0_ch30_txsz[21] ,_u0_ch30_txsz[20] , _u0_ch30_txsz[19] , _u0_ch30_txsz[18] ,_u0_ch30_txsz[17] , _u0_ch30_txsz[16] , _u0_ch30_txsz[15] ,_u0_ch30_txsz[14] , _u0_ch30_txsz[13] , _u0_ch30_txsz[12] ,_u0_ch30_txsz[11] , _u0_ch30_txsz[10] , _u0_ch30_txsz[9] ,_u0_ch30_txsz[8] , _u0_ch30_txsz[7] , _u0_ch30_txsz[6] ,_u0_ch30_txsz[5] , _u0_ch30_txsz[4] , _u0_ch30_txsz[3] ,_u0_ch30_txsz[2] , _u0_ch30_txsz[1] , _u0_ch30_txsz[0] ,_u0_ch30_adr0[31] , _u0_ch30_adr0[30] , _u0_ch30_adr0[29] ,_u0_ch30_adr0[28] , _u0_ch30_adr0[27] , _u0_ch30_adr0[26] ,_u0_ch30_adr0[25] , _u0_ch30_adr0[24] , _u0_ch30_adr0[23] ,_u0_ch30_adr0[22] , _u0_ch30_adr0[21] , _u0_ch30_adr0[20] ,_u0_ch30_adr0[19] , _u0_ch30_adr0[18] , _u0_ch30_adr0[17] ,_u0_ch30_adr0[16] , _u0_ch30_adr0[15] , _u0_ch30_adr0[14] ,_u0_ch30_adr0[13] , _u0_ch30_adr0[12] , _u0_ch30_adr0[11] ,_u0_ch30_adr0[10] , _u0_ch30_adr0[9] , _u0_ch30_adr0[8] ,_u0_ch30_adr0[7] , _u0_ch30_adr0[6] , _u0_ch30_adr0[5] ,_u0_ch30_adr0[4] , _u0_ch30_adr0[3] , _u0_ch30_adr0[2] ,_u0_ch30_adr0[1] , _u0_ch30_adr0[0] , _u0_ch30_adr1[31] ,_u0_ch30_adr1[30] , _u0_ch30_adr1[29] , _u0_ch30_adr1[28] ,_u0_ch30_adr1[27] , _u0_ch30_adr1[26] , _u0_ch30_adr1[25] ,_u0_ch30_adr1[24] , _u0_ch30_adr1[23] , _u0_ch30_adr1[22] ,_u0_ch30_adr1[21] , _u0_ch30_adr1[20] , _u0_ch30_adr1[19] ,_u0_ch30_adr1[18] , _u0_ch30_adr1[17] , _u0_ch30_adr1[16] ,_u0_ch30_adr1[15] , _u0_ch30_adr1[14] , _u0_ch30_adr1[13] ,_u0_ch30_adr1[12] , _u0_ch30_adr1[11] , _u0_ch30_adr1[10] ,_u0_ch30_adr1[9] , _u0_ch30_adr1[8] , _u0_ch30_adr1[7] ,_u0_ch30_adr1[6] , _u0_ch30_adr1[5] , _u0_ch30_adr1[4] ,_u0_ch30_adr1[3] , _u0_ch30_adr1[2] , _u0_ch30_adr1[1] ,_u0_ch30_adr1[0] , _u0_ch30_am0[31] , _u0_ch30_am0[30] ,_u0_ch30_am0[29] , _u0_ch30_am0[28] , _u0_ch30_am0[27] ,_u0_ch30_am0[26] , _u0_ch30_am0[25] , _u0_ch30_am0[24] ,_u0_ch30_am0[23] , _u0_ch30_am0[22] , _u0_ch30_am0[21] ,_u0_ch30_am0[20] , _u0_ch30_am0[19] , _u0_ch30_am0[18] ,_u0_ch30_am0[17] , _u0_ch30_am0[16] , _u0_ch30_am0[15] ,_u0_ch30_am0[14] , _u0_ch30_am0[13] , _u0_ch30_am0[12] ,_u0_ch30_am0[11] , _u0_ch30_am0[10] , _u0_ch30_am0[9] ,_u0_ch30_am0[8] , _u0_ch30_am0[7] , _u0_ch30_am0[6] ,_u0_ch30_am0[5] , _u0_ch30_am0[4] , _u0_ch30_am0[3] ,_u0_ch30_am0[2] , _u0_ch30_am0[1] , _u0_ch30_am0[0] ,_u0_ch30_am1[31] , _u0_ch30_am1[30] , _u0_ch30_am1[29] ,_u0_ch30_am1[28] , _u0_ch30_am1[27] , _u0_ch30_am1[26] ,_u0_ch30_am1[25] , _u0_ch30_am1[24] , _u0_ch30_am1[23] ,_u0_ch30_am1[22] , _u0_ch30_am1[21] , _u0_ch30_am1[20] ,_u0_ch30_am1[19] , _u0_ch30_am1[18] , _u0_ch30_am1[17] ,_u0_ch30_am1[16] , _u0_ch30_am1[15] , _u0_ch30_am1[14] ,_u0_ch30_am1[13] , _u0_ch30_am1[12] , _u0_ch30_am1[11] ,_u0_ch30_am1[10] , _u0_ch30_am1[9] , _u0_ch30_am1[8] ,_u0_ch30_am1[7] , _u0_ch30_am1[6] , _u0_ch30_am1[5] ,_u0_ch30_am1[4] , _u0_ch30_am1[3] , _u0_ch30_am1[2] ,_u0_ch30_am1[1] , _u0_ch30_am1[0] , _u0_n453 , _u0_n915 , _u0_n914 ,_u0_n913 , _u0_n912 , _u0_n911 , _u0_n910 , _u0_n909 , _u0_n908 ,_u0_n907 , _u0_n906 , _u0_n905 , _u0_n904 , _u0_n903 , _u0_n902 ,_u0_n901 , _u0_n900 , _u0_n899 , _u0_n898 , _u0_n897 , _u0_n896 ,_u0_n895 , _u0_n894 , _u0_n893 , _u0_n892 , _u0_n891 , _u0_n890 ,_u0_n889 , _u0_n888 , _u0_n887 , _u0_n886 , _u0_n885 , _u0_n884 ,_u0_n883 , _u0_n882 , _u0_n881 , _u0_n880 , _u0_n879 , _u0_n878 ,_u0_n877 , _u0_n876 , _u0_n875 , _u0_n874 , _u0_n873 , _u0_n872 ,_u0_n871 , _u0_n870 , _u0_n869 , _u0_n868 , _u0_n867 , _u0_n866 ,_u0_n865 , _u0_n864 , _u0_n863 , _u0_n862 , _u0_n861 , _u0_n860 ,_u0_n859 , _u0_n858 , _u0_n857 , _u0_n856 , _u0_n855 , _u0_n854 ,_u0_n853 , _u0_N3078 , _u0_ch_int_0_ , _u0_N3074 , _u0_N3073 ,_u0_N3072 , _u0_N3071 , _u0_N3070 , _u0_N3069 , _u0_N3068 ,_u0_N3067 , _u0_N3066 , _u0_N3065 , _u0_N3064 , _u0_N3063 ,_u0_N3062 , _u0_N3061 , _u0_N3060 , _u0_N3059 , _u0_N3058 ,_u0_N3057 , _u0_N3056 , _u0_N3055 , _u0_N3054 , _u0_N3053 ,_u0_N3052 , _u0_N3051 , _u0_N3050 , _u0_N3049 , _u0_N3048 ,_u0_N3047 , _u0_N3046 , _u0_N3045 , _u0_N3044 , _u0_N3043 ,_u0_u0_n1026 , _u0_u0_n1025 , _u0_u0_n1024 , _u0_u0_n1023 ,_u0_u0_n1022 , _u0_u0_n1021 , _u0_u0_n1020 , _u0_u0_n1019 ,_u0_u0_n1018 , _u0_u0_n1017 , _u0_u0_n1016 , _u0_u0_n1015 ,_u0_u0_n1014 , _u0_u0_n1013 , _u0_u0_n1012 , _u0_u0_n1011 ,_u0_u0_n1010 , _u0_u0_n1009 , _u0_u0_n1008 , _u0_u0_n1007 ,_u0_u0_n1006 , _u0_u0_n1005 , _u0_u0_n1004 , _u0_u0_n1003 ,_u0_u0_n1002 , _u0_u0_n1001 , _u0_u0_n1000 , _u0_u0_n999 ,_u0_u0_n998 , _u0_u0_n997 , _u0_u0_n996 , _u0_u0_n995 , _u0_u0_n994 ,_u0_u0_n993 , _u0_u0_n992 , _u0_u0_n991 , _u0_u0_n990 , _u0_u0_n989 ,_u0_u0_n988 , _u0_u0_n987 , _u0_u0_n986 , _u0_u0_n985 , _u0_u0_n984 ,_u0_u0_n983 , _u0_u0_n982 , _u0_u0_n981 , _u0_u0_n980 , _u0_u0_n979 ,_u0_u0_n978 , _u0_u0_n977 , _u0_u0_n976 , _u0_u0_n975 , _u0_u0_n974 ,_u0_u0_n973 , _u0_u0_n972 , _u0_u0_n971 , _u0_u0_n970 , _u0_u0_n969 ,_u0_u0_n968 , _u0_u0_n967 , _u0_u0_n966 , _u0_u0_n965 , _u0_u0_n964 ,_u0_u0_n963 , _u0_u0_n962 , _u0_u0_n961 , _u0_u0_n960 , _u0_u0_n959 ,_u0_u0_n958 , _u0_u0_n957 , _u0_u0_n956 , _u0_u0_n955 , _u0_u0_n954 ,_u0_u0_n953 , _u0_u0_n952 , _u0_u0_n951 , _u0_u0_n950 , _u0_u0_n949 ,_u0_u0_n948 , _u0_u0_n947 , _u0_u0_n946 , _u0_u0_n945 , _u0_u0_n944 ,_u0_u0_n943 , _u0_u0_n942 , _u0_u0_n941 , _u0_u0_n940 , _u0_u0_n939 ,_u0_u0_n938 , _u0_u0_n937 , _u0_u0_n936 , _u0_u0_n935 , _u0_u0_n934 ,_u0_u0_n933 , _u0_u0_n932 , _u0_u0_n931 , _u0_u0_n930 , _u0_u0_n929 ,_u0_u0_n928 , _u0_u0_n927 , _u0_u0_n926 , _u0_u0_n925 , _u0_u0_n924 ,_u0_u0_n923 , _u0_u0_n922 , _u0_u0_n921 , _u0_u0_n920 , _u0_u0_n919 ,_u0_u0_n918 , _u0_u0_n917 , _u0_u0_n916 , _u0_u0_n915 , _u0_u0_n914 ,_u0_u0_n913 , _u0_u0_n912 , _u0_u0_n911 , _u0_u0_n910 , _u0_u0_n909 ,_u0_u0_n908 , _u0_u0_n907 , _u0_u0_n906 , _u0_u0_n905 , _u0_u0_n904 ,_u0_u0_n903 , _u0_u0_n902 , _u0_u0_n901 , _u0_u0_n900 , _u0_u0_n899 ,_u0_u0_n898 , _u0_u0_n897 , _u0_u0_n896 , _u0_u0_n895 , _u0_u0_n894 ,_u0_u0_n893 , _u0_u0_n892 , _u0_u0_n891 , _u0_u0_n890 , _u0_u0_n889 ,_u0_u0_n888 , _u0_u0_n887 , _u0_u0_n886 , _u0_u0_n885 , _u0_u0_n884 ,_u0_u0_n883 , _u0_u0_n882 , _u0_u0_n881 , _u0_u0_n880 , _u0_u0_n879 ,_u0_u0_n878 , _u0_u0_n877 , _u0_u0_n876 , _u0_u0_n875 , _u0_u0_n874 ,_u0_u0_n873 , _u0_u0_n872 , _u0_u0_n871 , _u0_u0_n870 , _u0_u0_n869 ,_u0_u0_n868 , _u0_u0_n867 , _u0_u0_n866 , _u0_u0_n865 , _u0_u0_n864 ,_u0_u0_n863 , _u0_u0_n862 , _u0_u0_n861 , _u0_u0_n860 , _u0_u0_n859 ,_u0_u0_n858 , _u0_u0_n857 , _u0_u0_n856 , _u0_u0_n855 , _u0_u0_n854 ,_u0_u0_n853 , _u0_u0_n852 , _u0_u0_n851 , _u0_u0_n850 , _u0_u0_n849 ,_u0_u0_n848 , _u0_u0_n847 , _u0_u0_n846 , _u0_u0_n845 , _u0_u0_n844 ,_u0_u0_n843 , _u0_u0_n842 , _u0_u0_n841 , _u0_u0_n840 , _u0_u0_n839 ,_u0_u0_n838 , _u0_u0_n837 , _u0_u0_n836 , _u0_u0_n835 , _u0_u0_n834 ,_u0_u0_n833 , _u0_u0_n832 , _u0_u0_n831 , _u0_u0_n830 , _u0_u0_n829 ,_u0_u0_n828 , _u0_u0_n827 , _u0_u0_n826 , _u0_u0_n825 , _u0_u0_n824 ,_u0_u0_n823 , _u0_u0_n822 , _u0_u0_n821 , _u0_u0_n820 , _u0_u0_n819 ,_u0_u0_n818 , _u0_u0_n817 , _u0_u0_n816 , _u0_u0_n815 , _u0_u0_n814 ,_u0_u0_n813 , _u0_u0_n812 , _u0_u0_n811 , _u0_u0_n810 , _u0_u0_n809 ,_u0_u0_n808 , _u0_u0_n807 , _u0_u0_n806 , _u0_u0_n805 , _u0_u0_n804 ,_u0_u0_n803 , _u0_u0_n802 , _u0_u0_n801 , _u0_u0_n800 , _u0_u0_n799 ,_u0_u0_n798 , _u0_u0_n797 , _u0_u0_n796 , _u0_u0_n795 , _u0_u0_n794 ,_u0_u0_n793 , _u0_u0_n792 , _u0_u0_n791 , _u0_u0_n790 , _u0_u0_n789 ,_u0_u0_n788 , _u0_u0_n787 , _u0_u0_n786 , _u0_u0_n785 , _u0_u0_n784 ,_u0_u0_n783 , _u0_u0_n782 , _u0_u0_n781 , _u0_u0_n780 , _u0_u0_n779 ,_u0_u0_n778 , _u0_u0_n777 , _u0_u0_n776 , _u0_u0_n775 , _u0_u0_n774 ,_u0_u0_n773 , _u0_u0_n772 , _u0_u0_n771 , _u0_u0_n770 , _u0_u0_n769 ,_u0_u0_n768 , _u0_u0_n767 , _u0_u0_n766 , _u0_u0_n765 , _u0_u0_n764 ,_u0_u0_n763 , _u0_u0_n762 , _u0_u0_n761 , _u0_u0_n760 , _u0_u0_n759 ,_u0_u0_n758 , _u0_u0_n757 , _u0_u0_n756 , _u0_u0_n755 , _u0_u0_n754 ,_u0_u0_n753 , _u0_u0_n752 , _u0_u0_n751 , _u0_u0_pointer[31] ,_u0_u0_pointer[30] , _u0_u0_pointer[29] , _u0_u0_pointer[28] ,_u0_u0_pointer[27] , _u0_u0_pointer[26] , _u0_u0_pointer[25] ,_u0_u0_pointer[24] , _u0_u0_pointer[23] , _u0_u0_pointer[22] ,_u0_u0_pointer[21] , _u0_u0_pointer[20] , _u0_u0_pointer[19] ,_u0_u0_pointer[18] , _u0_u0_pointer[17] , _u0_u0_pointer[16] ,_u0_u0_pointer[15] , _u0_u0_pointer[14] , _u0_u0_pointer[13] ,_u0_u0_pointer[12] , _u0_u0_pointer[11] , _u0_u0_pointer[10] ,_u0_u0_pointer[9] , _u0_u0_pointer[8] , _u0_u0_pointer[7] ,_u0_u0_pointer[6] , _u0_u0_pointer[5] , _u0_u0_pointer[4] ,_u0_u0_pointer[3] , _u0_u0_pointer[2] , _u0_u0_pointer[1] ,_u0_u0_pointer[0] , _u0_u0_pointer_s[31] , _u0_u0_pointer_s[30] ,_u0_u0_pointer_s[29] , _u0_u0_pointer_s[28] , _u0_u0_pointer_s[27] ,_u0_u0_pointer_s[26] , _u0_u0_pointer_s[25] , _u0_u0_pointer_s[24] ,_u0_u0_pointer_s[23] , _u0_u0_pointer_s[22] , _u0_u0_pointer_s[21] ,_u0_u0_pointer_s[20] , _u0_u0_pointer_s[19] , _u0_u0_pointer_s[18] ,_u0_u0_pointer_s[17] , _u0_u0_pointer_s[16] , _u0_u0_pointer_s[15] ,_u0_u0_pointer_s[14] , _u0_u0_pointer_s[13] , _u0_u0_pointer_s[12] ,_u0_u0_pointer_s[11] , _u0_u0_pointer_s[10] , _u0_u0_pointer_s[9] ,_u0_u0_pointer_s[8] , _u0_u0_pointer_s[7] , _u0_u0_pointer_s[6] ,_u0_u0_pointer_s[5] , _u0_u0_pointer_s[4] , _u0_u0_pointer_s[3] ,_u0_u0_pointer_s[2] , _u0_u0_pointer_s[1] , _u0_u0_pointer_s[0] ,_u0_u0_ch_csr[31] , _u0_u0_ch_csr[30] , _u0_u0_ch_csr[29] ,_u0_u0_ch_csr[28] , _u0_u0_ch_csr[27] , _u0_u0_ch_csr[26] ,_u0_u0_ch_csr[25] , _u0_u0_ch_csr[24] , _u0_u0_ch_csr[23] ,_u0_u0_ch_csr[9] , _u0_u0_ch_txsz[31] , _u0_u0_ch_txsz[30] ,_u0_u0_ch_txsz[29] , _u0_u0_ch_txsz[28] , _u0_u0_ch_txsz[27] ,_u0_u0_ch_txsz[14] , _u0_u0_ch_txsz[13] , _u0_u0_ch_txsz[12] ,_u0_u0_ch_adr0[1] , _u0_u0_ch_adr0[0] , _u0_u0_ch_adr1[1] ,_u0_u0_ch_adr1[0] , _u0_u0_ch_am0[31] , _u0_u0_ch_am0[30] ,_u0_u0_ch_am0[29] , _u0_u0_ch_am0[28] , _u0_u0_ch_am0[27] ,_u0_u0_ch_am0[26] , _u0_u0_ch_am0[25] , _u0_u0_ch_am0[24] ,_u0_u0_ch_am0[23] , _u0_u0_ch_am0[22] , _u0_u0_ch_am0[21] ,_u0_u0_ch_am0[20] , _u0_u0_ch_am0[19] , _u0_u0_ch_am0[18] ,_u0_u0_ch_am0[17] , _u0_u0_ch_am0[16] , _u0_u0_ch_am0[15] ,_u0_u0_ch_am0[14] , _u0_u0_ch_am0[13] , _u0_u0_ch_am0[12] ,_u0_u0_ch_am0[11] , _u0_u0_ch_am0[10] , _u0_u0_ch_am0[9] ,_u0_u0_ch_am0[8] , _u0_u0_ch_am0[7] , _u0_u0_ch_am0[6] ,_u0_u0_ch_am0[5] , _u0_u0_ch_am0[4] , _u0_u0_ch_am0[3] ,_u0_u0_ch_am0[2] , _u0_u0_ch_am0[1] , _u0_u0_ch_am0[0] ,_u0_u0_ch_am1[31] , _u0_u0_ch_am1[30] , _u0_u0_ch_am1[29] ,_u0_u0_ch_am1[28] , _u0_u0_ch_am1[27] , _u0_u0_ch_am1[26] ,_u0_u0_ch_am1[25] , _u0_u0_ch_am1[24] , _u0_u0_ch_am1[23] ,_u0_u0_ch_am1[22] , _u0_u0_ch_am1[21] , _u0_u0_ch_am1[20] ,_u0_u0_ch_am1[19] , _u0_u0_ch_am1[18] , _u0_u0_ch_am1[17] ,_u0_u0_ch_am1[16] , _u0_u0_ch_am1[15] , _u0_u0_ch_am1[14] ,_u0_u0_ch_am1[13] , _u0_u0_ch_am1[12] , _u0_u0_ch_am1[11] ,_u0_u0_ch_am1[10] , _u0_u0_ch_am1[9] , _u0_u0_ch_am1[8] ,_u0_u0_ch_am1[7] , _u0_u0_ch_am1[6] , _u0_u0_ch_am1[5] ,_u0_u0_ch_am1[4] , _u0_u0_ch_am1[3] , _u0_u0_ch_am1[2] ,_u0_u0_ch_am1[1] , _u0_u0_ch_am1[0] , _u0_u0_sw_pointer[31] ,_u0_u0_sw_pointer[30] , _u0_u0_sw_pointer[29] ,_u0_u0_sw_pointer[28] , _u0_u0_sw_pointer[27] ,_u0_u0_sw_pointer[26] , _u0_u0_sw_pointer[25] ,_u0_u0_sw_pointer[24] , _u0_u0_sw_pointer[23] ,_u0_u0_sw_pointer[22] , _u0_u0_sw_pointer[21] ,_u0_u0_sw_pointer[20] , _u0_u0_sw_pointer[19] ,_u0_u0_sw_pointer[18] , _u0_u0_sw_pointer[17] ,_u0_u0_sw_pointer[16] , _u0_u0_sw_pointer[15] ,_u0_u0_sw_pointer[14] , _u0_u0_sw_pointer[13] ,_u0_u0_sw_pointer[12] , _u0_u0_sw_pointer[11] ,_u0_u0_sw_pointer[10] , _u0_u0_sw_pointer[9] , _u0_u0_sw_pointer[8] ,_u0_u0_sw_pointer[7] , _u0_u0_sw_pointer[6] , _u0_u0_sw_pointer[5] ,_u0_u0_sw_pointer[4] , _u0_u0_sw_pointer[3] , _u0_u0_sw_pointer[2] ,_u0_u0_sw_pointer[1] , _u0_u0_sw_pointer[0] , _u0_u0_ch_dis ,_u0_u0_n439 , _u0_u0_n438 , _u0_u0_n437 , _u0_u0_n436 , _u0_u0_n435 ,_u0_u0_n434 , _u0_u0_n433 , _u0_u0_n432 , _u0_u0_n431 , _u0_u0_n430 ,_u0_u0_n429 , _u0_u0_n428 , _u0_u0_n427 , _u0_u0_n426 , _u0_u0_n425 ,_u0_u0_n424 , _u0_u0_n423 , _u0_u0_n422 , _u0_u0_n421 , _u0_u0_n420 ,_u0_u0_n419 , _u0_u0_n418 , _u0_u0_n417 , _u0_u0_n416 , _u0_u0_n415 ,_u0_u0_n414 , _u0_u0_n413 , _u0_u0_n412 , _u0_u0_n411 , _u0_u0_n410 ,_u0_u0_n409 , _u0_u0_n408 , _u0_u0_n407 , _u0_u0_n406 , _u0_u0_n405 ,_u0_u0_n404 , _u0_u0_n403 , _u0_u0_n402 , _u0_u0_n401 , _u0_u0_n400 ,_u0_u0_n399 , _u0_u0_n398 , _u0_u0_n397 , _u0_u0_n396 , _u0_u0_n395 ,_u0_u0_n394 , _u0_u0_n393 , _u0_u0_n392 , _u0_u0_n391 , _u0_u0_n390 ,_u0_u0_n389 , _u0_u0_n388 , _u0_u0_n387 , _u0_u0_n386 , _u0_u0_n385 ,_u0_u0_n384 , _u0_u0_n383 , _u0_u0_n382 , _u0_u0_n381 , _u0_u0_n380 ,_u0_u0_n379 , _u0_u0_n378 , _u0_u0_n377 , _u0_u0_n376 , _u0_u0_n375 ,_u0_u0_n374 , _u0_u0_n373 , _u0_u0_n372 , _u0_u0_n371 , _u0_u0_n370 ,_u0_u0_n369 , _u0_u0_n368 , _u0_u0_n367 , _u0_u0_n366 , _u0_u0_n365 ,_u0_u0_n364 , _u0_u0_n363 , _u0_u0_n362 , _u0_u0_n361 , _u0_u0_n360 ,_u0_u0_n359 , _u0_u0_n358 , _u0_u0_n357 , _u0_u0_n356 , _u0_u0_n355 ,_u0_u0_n354 , _u0_u0_n353 , _u0_u0_n352 , _u0_u0_n351 , _u0_u0_n350 ,_u0_u0_n349 , _u0_u0_n348 , _u0_u0_n347 , _u0_u0_n346 , _u0_u0_n345 ,_u0_u0_n344 , _u0_u0_n343 , _u0_u0_n342 , _u0_u0_n341 , _u0_u0_n340 ,_u0_u0_n339 , _u0_u0_n338 , _u0_u0_n337 , _u0_u0_n336 , _u0_u0_n335 ,_u0_u0_n334 , _u0_u0_n333 , _u0_u0_n326 , _u0_u0_N24 , _u0_u0_N23 ,_u0_u1_pointer[31] , _u0_u1_pointer[30] , _u0_u1_pointer[29] ,_u0_u1_pointer[28] , _u0_u1_pointer[27] , _u0_u1_pointer[26] ,_u0_u1_pointer[25] , _u0_u1_pointer[24] , _u0_u1_pointer[23] ,_u0_u1_pointer[22] , _u0_u1_pointer[21] , _u0_u1_pointer[20] ,_u0_u1_pointer[19] , _u0_u1_pointer[18] , _u0_u1_pointer[17] ,_u0_u1_pointer[16] , _u0_u1_pointer[15] , _u0_u1_pointer[14] ,_u0_u1_pointer[13] , _u0_u1_pointer[12] , _u0_u1_pointer[11] ,_u0_u1_pointer[10] , _u0_u1_pointer[9] , _u0_u1_pointer[8] ,_u0_u1_pointer[7] , _u0_u1_pointer[6] , _u0_u1_pointer[5] ,_u0_u1_pointer[4] , _u0_u1_pointer[3] , _u0_u1_pointer[2] ,_u0_u1_pointer[1] , _u0_u1_pointer[0] , _u0_u1_pointer_s[31] ,_u0_u1_pointer_s[30] , _u0_u1_pointer_s[29] , _u0_u1_pointer_s[28] ,_u0_u1_pointer_s[27] , _u0_u1_pointer_s[26] , _u0_u1_pointer_s[25] ,_u0_u1_pointer_s[24] , _u0_u1_pointer_s[23] , _u0_u1_pointer_s[22] ,_u0_u1_pointer_s[21] , _u0_u1_pointer_s[20] , _u0_u1_pointer_s[19] ,_u0_u1_pointer_s[18] , _u0_u1_pointer_s[17] , _u0_u1_pointer_s[16] ,_u0_u1_pointer_s[15] , _u0_u1_pointer_s[14] , _u0_u1_pointer_s[13] ,_u0_u1_pointer_s[12] , _u0_u1_pointer_s[11] , _u0_u1_pointer_s[10] ,_u0_u1_pointer_s[9] , _u0_u1_pointer_s[8] , _u0_u1_pointer_s[7] ,_u0_u1_pointer_s[6] , _u0_u1_pointer_s[5] , _u0_u1_pointer_s[4] ,_u0_u1_pointer_s[3] , _u0_u1_pointer_s[2] , _u0_u1_pointer_s[1] ,_u0_u1_pointer_s[0] , _u0_u1_ch_csr[31] , _u0_u1_ch_csr[30] ,_u0_u1_ch_csr[29] , _u0_u1_ch_csr[28] , _u0_u1_ch_csr[27] ,_u0_u1_ch_csr[26] , _u0_u1_ch_csr[25] , _u0_u1_ch_csr[24] ,_u0_u1_ch_csr[23] , _u0_u1_ch_csr[22] , _u0_u1_ch_csr[21] ,_u0_u1_ch_csr[20] , _u0_u1_ch_csr[19] , _u0_u1_ch_csr[18] ,_u0_u1_ch_csr[17] , _u0_u1_ch_csr[16] , _u0_u1_ch_csr[15] ,_u0_u1_ch_csr[14] , _u0_u1_ch_csr[13] , _u0_u1_ch_csr[12] ,_u0_u1_ch_csr[11] , _u0_u1_ch_csr[10] , _u0_u1_ch_csr[9] ,_u0_u1_ch_csr[8] , _u0_u1_ch_csr[7] , _u0_u1_ch_csr[6] ,_u0_u1_ch_csr[5] , _u0_u1_ch_csr[4] , _u0_u1_ch_csr[3] ,_u0_u1_ch_csr[2] , _u0_u1_ch_csr[1] , _u0_u1_ch_csr[0] ,_u0_u1_ch_txsz[31] , _u0_u1_ch_txsz[30] , _u0_u1_ch_txsz[29] ,_u0_u1_ch_txsz[28] , _u0_u1_ch_txsz[27] , _u0_u1_ch_txsz[26] ,_u0_u1_ch_txsz[25] , _u0_u1_ch_txsz[24] , _u0_u1_ch_txsz[23] ,_u0_u1_ch_txsz[22] , _u0_u1_ch_txsz[21] , _u0_u1_ch_txsz[20] ,_u0_u1_ch_txsz[19] , _u0_u1_ch_txsz[18] , _u0_u1_ch_txsz[17] ,_u0_u1_ch_txsz[16] , _u0_u1_ch_txsz[15] , _u0_u1_ch_txsz[14] ,_u0_u1_ch_txsz[13] , _u0_u1_ch_txsz[12] , _u0_u1_ch_txsz[11] ,_u0_u1_ch_txsz[10] , _u0_u1_ch_txsz[9] , _u0_u1_ch_txsz[8] ,_u0_u1_ch_txsz[7] , _u0_u1_ch_txsz[6] , _u0_u1_ch_txsz[5] ,_u0_u1_ch_txsz[4] , _u0_u1_ch_txsz[3] , _u0_u1_ch_txsz[2] ,_u0_u1_ch_txsz[1] , _u0_u1_ch_txsz[0] , _u0_u1_ch_adr0[31] ,_u0_u1_ch_adr0[30] , _u0_u1_ch_adr0[29] , _u0_u1_ch_adr0[28] ,_u0_u1_ch_adr0[27] , _u0_u1_ch_adr0[26] , _u0_u1_ch_adr0[25] ,_u0_u1_ch_adr0[24] , _u0_u1_ch_adr0[23] , _u0_u1_ch_adr0[22] ,_u0_u1_ch_adr0[21] , _u0_u1_ch_adr0[20] , _u0_u1_ch_adr0[19] ,_u0_u1_ch_adr0[18] , _u0_u1_ch_adr0[17] , _u0_u1_ch_adr0[16] ,_u0_u1_ch_adr0[15] , _u0_u1_ch_adr0[14] , _u0_u1_ch_adr0[13] ,_u0_u1_ch_adr0[12] , _u0_u1_ch_adr0[11] , _u0_u1_ch_adr0[10] ,_u0_u1_ch_adr0[9] , _u0_u1_ch_adr0[8] , _u0_u1_ch_adr0[7] ,_u0_u1_ch_adr0[6] , _u0_u1_ch_adr0[5] , _u0_u1_ch_adr0[4] ,_u0_u1_ch_adr0[3] , _u0_u1_ch_adr0[2] , _u0_u1_ch_adr0[1] ,_u0_u1_ch_adr0[0] , _u0_u1_ch_adr1[31] , _u0_u1_ch_adr1[30] ,_u0_u1_ch_adr1[29] , _u0_u1_ch_adr1[28] , _u0_u1_ch_adr1[27] ,_u0_u1_ch_adr1[26] , _u0_u1_ch_adr1[25] , _u0_u1_ch_adr1[24] ,_u0_u1_ch_adr1[23] , _u0_u1_ch_adr1[22] , _u0_u1_ch_adr1[21] ,_u0_u1_ch_adr1[20] , _u0_u1_ch_adr1[19] , _u0_u1_ch_adr1[18] ,_u0_u1_ch_adr1[17] , _u0_u1_ch_adr1[16] , _u0_u1_ch_adr1[15] ,_u0_u1_ch_adr1[14] , _u0_u1_ch_adr1[13] , _u0_u1_ch_adr1[12] ,_u0_u1_ch_adr1[11] , _u0_u1_ch_adr1[10] , _u0_u1_ch_adr1[9] ,_u0_u1_ch_adr1[8] , _u0_u1_ch_adr1[7] , _u0_u1_ch_adr1[6] ,_u0_u1_ch_adr1[5] , _u0_u1_ch_adr1[4] , _u0_u1_ch_adr1[3] ,_u0_u1_ch_adr1[2] , _u0_u1_ch_adr1[1] , _u0_u1_ch_adr1[0] ,_u0_u1_ch_am0[31] , _u0_u1_ch_am0[30] , _u0_u1_ch_am0[29] ,_u0_u1_ch_am0[28] , _u0_u1_ch_am0[27] , _u0_u1_ch_am0[26] ,_u0_u1_ch_am0[25] , _u0_u1_ch_am0[24] , _u0_u1_ch_am0[23] ,_u0_u1_ch_am0[22] , _u0_u1_ch_am0[21] , _u0_u1_ch_am0[20] ,_u0_u1_ch_am0[19] , _u0_u1_ch_am0[18] , _u0_u1_ch_am0[17] ,_u0_u1_ch_am0[16] , _u0_u1_ch_am0[15] , _u0_u1_ch_am0[14] ,_u0_u1_ch_am0[13] , _u0_u1_ch_am0[12] , _u0_u1_ch_am0[11] ,_u0_u1_ch_am0[10] , _u0_u1_ch_am0[9] , _u0_u1_ch_am0[8] ,_u0_u1_ch_am0[7] , _u0_u1_ch_am0[6] , _u0_u1_ch_am0[5] ,_u0_u1_ch_am0[4] , _u0_u1_ch_am0[3] , _u0_u1_ch_am0[2] ,_u0_u1_ch_am0[1] , _u0_u1_ch_am0[0] , _u0_u1_ch_am1[31] ,_u0_u1_ch_am1[30] , _u0_u1_ch_am1[29] , _u0_u1_ch_am1[28] ,_u0_u1_ch_am1[27] , _u0_u1_ch_am1[26] , _u0_u1_ch_am1[25] ,_u0_u1_ch_am1[24] , _u0_u1_ch_am1[23] , _u0_u1_ch_am1[22] ,_u0_u1_ch_am1[21] , _u0_u1_ch_am1[20] , _u0_u1_ch_am1[19] ,_u0_u1_ch_am1[18] , _u0_u1_ch_am1[17] , _u0_u1_ch_am1[16] ,_u0_u1_ch_am1[15] , _u0_u1_ch_am1[14] , _u0_u1_ch_am1[13] ,_u0_u1_ch_am1[12] , _u0_u1_ch_am1[11] , _u0_u1_ch_am1[10] ,_u0_u1_ch_am1[9] , _u0_u1_ch_am1[8] , _u0_u1_ch_am1[7] ,_u0_u1_ch_am1[6] , _u0_u1_ch_am1[5] , _u0_u1_ch_am1[4] ,_u0_u1_ch_am1[3] , _u0_u1_ch_am1[2] , _u0_u1_ch_am1[1] ,_u0_u1_ch_am1[0] , _u0_u1_sw_pointer[31] , _u0_u1_sw_pointer[30] ,_u0_u1_sw_pointer[29] , _u0_u1_sw_pointer[28] ,_u0_u1_sw_pointer[27] , _u0_u1_sw_pointer[26] ,_u0_u1_sw_pointer[25] , _u0_u1_sw_pointer[24] ,_u0_u1_sw_pointer[23] , _u0_u1_sw_pointer[22] ,_u0_u1_sw_pointer[21] , _u0_u1_sw_pointer[20] ,_u0_u1_sw_pointer[19] , _u0_u1_sw_pointer[18] ,_u0_u1_sw_pointer[17] , _u0_u1_sw_pointer[16] ,_u0_u1_sw_pointer[15] , _u0_u1_sw_pointer[14] ,_u0_u1_sw_pointer[13] , _u0_u1_sw_pointer[12] ,_u0_u1_sw_pointer[11] , _u0_u1_sw_pointer[10] , _u0_u1_sw_pointer[9] ,_u0_u1_sw_pointer[8] , _u0_u1_sw_pointer[7] , _u0_u1_sw_pointer[6] ,_u0_u1_sw_pointer[5] , _u0_u1_sw_pointer[4] , _u0_u1_sw_pointer[3] ,_u0_u1_sw_pointer[2] , _u0_u1_sw_pointer[1] , _u0_u1_sw_pointer[0] ,_u0_u1_ch_stop , _u0_u1_ch_dis , _u0_u1_int , _u0_u2_pointer[31] ,_u0_u2_pointer[30] , _u0_u2_pointer[29] , _u0_u2_pointer[28] ,_u0_u2_pointer[27] , _u0_u2_pointer[26] , _u0_u2_pointer[25] ,_u0_u2_pointer[24] , _u0_u2_pointer[23] , _u0_u2_pointer[22] ,_u0_u2_pointer[21] , _u0_u2_pointer[20] , _u0_u2_pointer[19] ,_u0_u2_pointer[18] , _u0_u2_pointer[17] , _u0_u2_pointer[16] ,_u0_u2_pointer[15] , _u0_u2_pointer[14] , _u0_u2_pointer[13] ,_u0_u2_pointer[12] , _u0_u2_pointer[11] , _u0_u2_pointer[10] ,_u0_u2_pointer[9] , _u0_u2_pointer[8] , _u0_u2_pointer[7] ,_u0_u2_pointer[6] , _u0_u2_pointer[5] , _u0_u2_pointer[4] ,_u0_u2_pointer[3] , _u0_u2_pointer[2] , _u0_u2_pointer[1] ,_u0_u2_pointer[0] , _u0_u2_pointer_s[31] , _u0_u2_pointer_s[30] ,_u0_u2_pointer_s[29] , _u0_u2_pointer_s[28] , _u0_u2_pointer_s[27] ,_u0_u2_pointer_s[26] , _u0_u2_pointer_s[25] , _u0_u2_pointer_s[24] ,_u0_u2_pointer_s[23] , _u0_u2_pointer_s[22] , _u0_u2_pointer_s[21] ,_u0_u2_pointer_s[20] , _u0_u2_pointer_s[19] , _u0_u2_pointer_s[18] ,_u0_u2_pointer_s[17] , _u0_u2_pointer_s[16] , _u0_u2_pointer_s[15] ,_u0_u2_pointer_s[14] , _u0_u2_pointer_s[13] , _u0_u2_pointer_s[12] ,_u0_u2_pointer_s[11] , _u0_u2_pointer_s[10] , _u0_u2_pointer_s[9] ,_u0_u2_pointer_s[8] , _u0_u2_pointer_s[7] , _u0_u2_pointer_s[6] ,_u0_u2_pointer_s[5] , _u0_u2_pointer_s[4] , _u0_u2_pointer_s[3] ,_u0_u2_pointer_s[2] , _u0_u2_pointer_s[1] , _u0_u2_pointer_s[0] ,_u0_u2_ch_csr[31] , _u0_u2_ch_csr[30] , _u0_u2_ch_csr[29] ,_u0_u2_ch_csr[28] , _u0_u2_ch_csr[27] , _u0_u2_ch_csr[26] ,_u0_u2_ch_csr[25] , _u0_u2_ch_csr[24] , _u0_u2_ch_csr[23] ,_u0_u2_ch_csr[22] , _u0_u2_ch_csr[21] , _u0_u2_ch_csr[20] ,_u0_u2_ch_csr[19] , _u0_u2_ch_csr[18] , _u0_u2_ch_csr[17] ,_u0_u2_ch_csr[16] , _u0_u2_ch_csr[15] , _u0_u2_ch_csr[14] ,_u0_u2_ch_csr[13] , _u0_u2_ch_csr[12] , _u0_u2_ch_csr[11] ,_u0_u2_ch_csr[10] , _u0_u2_ch_csr[9] , _u0_u2_ch_csr[8] ,_u0_u2_ch_csr[7] , _u0_u2_ch_csr[6] , _u0_u2_ch_csr[5] ,_u0_u2_ch_csr[4] , _u0_u2_ch_csr[3] , _u0_u2_ch_csr[2] ,_u0_u2_ch_csr[1] , _u0_u2_ch_csr[0] , _u0_u2_ch_txsz[31] ,_u0_u2_ch_txsz[30] , _u0_u2_ch_txsz[29] , _u0_u2_ch_txsz[28] ,_u0_u2_ch_txsz[27] , _u0_u2_ch_txsz[26] , _u0_u2_ch_txsz[25] ,_u0_u2_ch_txsz[24] , _u0_u2_ch_txsz[23] , _u0_u2_ch_txsz[22] ,_u0_u2_ch_txsz[21] , _u0_u2_ch_txsz[20] , _u0_u2_ch_txsz[19] ,_u0_u2_ch_txsz[18] , _u0_u2_ch_txsz[17] , _u0_u2_ch_txsz[16] ,_u0_u2_ch_txsz[15] , _u0_u2_ch_txsz[14] , _u0_u2_ch_txsz[13] ,_u0_u2_ch_txsz[12] , _u0_u2_ch_txsz[11] , _u0_u2_ch_txsz[10] ,_u0_u2_ch_txsz[9] , _u0_u2_ch_txsz[8] , _u0_u2_ch_txsz[7] ,_u0_u2_ch_txsz[6] , _u0_u2_ch_txsz[5] , _u0_u2_ch_txsz[4] ,_u0_u2_ch_txsz[3] , _u0_u2_ch_txsz[2] , _u0_u2_ch_txsz[1] ,_u0_u2_ch_txsz[0] , _u0_u2_ch_adr0[31] , _u0_u2_ch_adr0[30] ,_u0_u2_ch_adr0[29] , _u0_u2_ch_adr0[28] , _u0_u2_ch_adr0[27] ,_u0_u2_ch_adr0[26] , _u0_u2_ch_adr0[25] , _u0_u2_ch_adr0[24] ,_u0_u2_ch_adr0[23] , _u0_u2_ch_adr0[22] , _u0_u2_ch_adr0[21] ,_u0_u2_ch_adr0[20] , _u0_u2_ch_adr0[19] , _u0_u2_ch_adr0[18] ,_u0_u2_ch_adr0[17] , _u0_u2_ch_adr0[16] , _u0_u2_ch_adr0[15] ,_u0_u2_ch_adr0[14] , _u0_u2_ch_adr0[13] , _u0_u2_ch_adr0[12] ,_u0_u2_ch_adr0[11] , _u0_u2_ch_adr0[10] , _u0_u2_ch_adr0[9] ,_u0_u2_ch_adr0[8] , _u0_u2_ch_adr0[7] , _u0_u2_ch_adr0[6] ,_u0_u2_ch_adr0[5] , _u0_u2_ch_adr0[4] , _u0_u2_ch_adr0[3] ,_u0_u2_ch_adr0[2] , _u0_u2_ch_adr0[1] , _u0_u2_ch_adr0[0] ,_u0_u2_ch_adr1[31] , _u0_u2_ch_adr1[30] , _u0_u2_ch_adr1[29] ,_u0_u2_ch_adr1[28] , _u0_u2_ch_adr1[27] , _u0_u2_ch_adr1[26] ,_u0_u2_ch_adr1[25] , _u0_u2_ch_adr1[24] , _u0_u2_ch_adr1[23] ,_u0_u2_ch_adr1[22] , _u0_u2_ch_adr1[21] , _u0_u2_ch_adr1[20] ,_u0_u2_ch_adr1[19] , _u0_u2_ch_adr1[18] , _u0_u2_ch_adr1[17] ,_u0_u2_ch_adr1[16] , _u0_u2_ch_adr1[15] , _u0_u2_ch_adr1[14] ,_u0_u2_ch_adr1[13] , _u0_u2_ch_adr1[12] , _u0_u2_ch_adr1[11] ,_u0_u2_ch_adr1[10] , _u0_u2_ch_adr1[9] , _u0_u2_ch_adr1[8] ,_u0_u2_ch_adr1[7] , _u0_u2_ch_adr1[6] , _u0_u2_ch_adr1[5] ,_u0_u2_ch_adr1[4] , _u0_u2_ch_adr1[3] , _u0_u2_ch_adr1[2] ,_u0_u2_ch_adr1[1] , _u0_u2_ch_adr1[0] , _u0_u2_ch_am0[31] ,_u0_u2_ch_am0[30] , _u0_u2_ch_am0[29] , _u0_u2_ch_am0[28] ,_u0_u2_ch_am0[27] , _u0_u2_ch_am0[26] , _u0_u2_ch_am0[25] ,_u0_u2_ch_am0[24] , _u0_u2_ch_am0[23] , _u0_u2_ch_am0[22] ,_u0_u2_ch_am0[21] , _u0_u2_ch_am0[20] , _u0_u2_ch_am0[19] ,_u0_u2_ch_am0[18] , _u0_u2_ch_am0[17] , _u0_u2_ch_am0[16] ,_u0_u2_ch_am0[15] , _u0_u2_ch_am0[14] , _u0_u2_ch_am0[13] ,_u0_u2_ch_am0[12] , _u0_u2_ch_am0[11] , _u0_u2_ch_am0[10] ,_u0_u2_ch_am0[9] , _u0_u2_ch_am0[8] , _u0_u2_ch_am0[7] ,_u0_u2_ch_am0[6] , _u0_u2_ch_am0[5] , _u0_u2_ch_am0[4] ,_u0_u2_ch_am0[3] , _u0_u2_ch_am0[2] , _u0_u2_ch_am0[1] ,_u0_u2_ch_am0[0] , _u0_u2_ch_am1[31] , _u0_u2_ch_am1[30] ,_u0_u2_ch_am1[29] , _u0_u2_ch_am1[28] , _u0_u2_ch_am1[27] ,_u0_u2_ch_am1[26] , _u0_u2_ch_am1[25] , _u0_u2_ch_am1[24] ,_u0_u2_ch_am1[23] , _u0_u2_ch_am1[22] , _u0_u2_ch_am1[21] ,_u0_u2_ch_am1[20] , _u0_u2_ch_am1[19] , _u0_u2_ch_am1[18] ,_u0_u2_ch_am1[17] , _u0_u2_ch_am1[16] , _u0_u2_ch_am1[15] ,_u0_u2_ch_am1[14] , _u0_u2_ch_am1[13] , _u0_u2_ch_am1[12] ,_u0_u2_ch_am1[11] , _u0_u2_ch_am1[10] , _u0_u2_ch_am1[9] ,_u0_u2_ch_am1[8] , _u0_u2_ch_am1[7] , _u0_u2_ch_am1[6] ,_u0_u2_ch_am1[5] , _u0_u2_ch_am1[4] , _u0_u2_ch_am1[3] ,_u0_u2_ch_am1[2] , _u0_u2_ch_am1[1] , _u0_u2_ch_am1[0] ,_u0_u2_sw_pointer[31] , _u0_u2_sw_pointer[30] ,_u0_u2_sw_pointer[29] , _u0_u2_sw_pointer[28] ,_u0_u2_sw_pointer[27] , _u0_u2_sw_pointer[26] ,_u0_u2_sw_pointer[25] , _u0_u2_sw_pointer[24] ,_u0_u2_sw_pointer[23] , _u0_u2_sw_pointer[22] ,_u0_u2_sw_pointer[21] , _u0_u2_sw_pointer[20] ,_u0_u2_sw_pointer[19] , _u0_u2_sw_pointer[18] ,_u0_u2_sw_pointer[17] , _u0_u2_sw_pointer[16] ,_u0_u2_sw_pointer[15] , _u0_u2_sw_pointer[14] ,_u0_u2_sw_pointer[13] , _u0_u2_sw_pointer[12] ,_u0_u2_sw_pointer[11] , _u0_u2_sw_pointer[10] , _u0_u2_sw_pointer[9] ,_u0_u2_sw_pointer[8] , _u0_u2_sw_pointer[7] , _u0_u2_sw_pointer[6] ,_u0_u2_sw_pointer[5] , _u0_u2_sw_pointer[4] , _u0_u2_sw_pointer[3] ,_u0_u2_sw_pointer[2] , _u0_u2_sw_pointer[1] , _u0_u2_sw_pointer[0] ,_u0_u2_ch_stop , _u0_u2_ch_dis , _u0_u2_int , _u0_u3_pointer[31] ,_u0_u3_pointer[30] , _u0_u3_pointer[29] , _u0_u3_pointer[28] ,_u0_u3_pointer[27] , _u0_u3_pointer[26] , _u0_u3_pointer[25] ,_u0_u3_pointer[24] , _u0_u3_pointer[23] , _u0_u3_pointer[22] ,_u0_u3_pointer[21] , _u0_u3_pointer[20] , _u0_u3_pointer[19] ,_u0_u3_pointer[18] , _u0_u3_pointer[17] , _u0_u3_pointer[16] ,_u0_u3_pointer[15] , _u0_u3_pointer[14] , _u0_u3_pointer[13] ,_u0_u3_pointer[12] , _u0_u3_pointer[11] , _u0_u3_pointer[10] ,_u0_u3_pointer[9] , _u0_u3_pointer[8] , _u0_u3_pointer[7] ,_u0_u3_pointer[6] , _u0_u3_pointer[5] , _u0_u3_pointer[4] ,_u0_u3_pointer[3] , _u0_u3_pointer[2] , _u0_u3_pointer[1] ,_u0_u3_pointer[0] , _u0_u3_pointer_s[31] , _u0_u3_pointer_s[30] ,_u0_u3_pointer_s[29] , _u0_u3_pointer_s[28] , _u0_u3_pointer_s[27] ,_u0_u3_pointer_s[26] , _u0_u3_pointer_s[25] , _u0_u3_pointer_s[24] ,_u0_u3_pointer_s[23] , _u0_u3_pointer_s[22] , _u0_u3_pointer_s[21] ,_u0_u3_pointer_s[20] , _u0_u3_pointer_s[19] , _u0_u3_pointer_s[18] ,_u0_u3_pointer_s[17] , _u0_u3_pointer_s[16] , _u0_u3_pointer_s[15] ,_u0_u3_pointer_s[14] , _u0_u3_pointer_s[13] , _u0_u3_pointer_s[12] ,_u0_u3_pointer_s[11] , _u0_u3_pointer_s[10] , _u0_u3_pointer_s[9] ,_u0_u3_pointer_s[8] , _u0_u3_pointer_s[7] , _u0_u3_pointer_s[6] ,_u0_u3_pointer_s[5] , _u0_u3_pointer_s[4] , _u0_u3_pointer_s[3] ,_u0_u3_pointer_s[2] , _u0_u3_pointer_s[1] , _u0_u3_pointer_s[0] ,_u0_u3_ch_csr[31] , _u0_u3_ch_csr[30] , _u0_u3_ch_csr[29] ,_u0_u3_ch_csr[28] , _u0_u3_ch_csr[27] , _u0_u3_ch_csr[26] ,_u0_u3_ch_csr[25] , _u0_u3_ch_csr[24] , _u0_u3_ch_csr[23] ,_u0_u3_ch_csr[22] , _u0_u3_ch_csr[21] , _u0_u3_ch_csr[20] ,_u0_u3_ch_csr[19] , _u0_u3_ch_csr[18] , _u0_u3_ch_csr[17] ,_u0_u3_ch_csr[16] , _u0_u3_ch_csr[15] , _u0_u3_ch_csr[14] ,_u0_u3_ch_csr[13] , _u0_u3_ch_csr[12] , _u0_u3_ch_csr[11] ,_u0_u3_ch_csr[10] , _u0_u3_ch_csr[9] , _u0_u3_ch_csr[8] ,_u0_u3_ch_csr[7] , _u0_u3_ch_csr[6] , _u0_u3_ch_csr[5] ,_u0_u3_ch_csr[4] , _u0_u3_ch_csr[3] , _u0_u3_ch_csr[2] ,_u0_u3_ch_csr[1] , _u0_u3_ch_csr[0] , _u0_u3_ch_txsz[31] ,_u0_u3_ch_txsz[30] , _u0_u3_ch_txsz[29] , _u0_u3_ch_txsz[28] ,_u0_u3_ch_txsz[27] , _u0_u3_ch_txsz[26] , _u0_u3_ch_txsz[25] ,_u0_u3_ch_txsz[24] , _u0_u3_ch_txsz[23] , _u0_u3_ch_txsz[22] ,_u0_u3_ch_txsz[21] , _u0_u3_ch_txsz[20] , _u0_u3_ch_txsz[19] ,_u0_u3_ch_txsz[18] , _u0_u3_ch_txsz[17] , _u0_u3_ch_txsz[16] ,_u0_u3_ch_txsz[15] , _u0_u3_ch_txsz[14] , _u0_u3_ch_txsz[13] ,_u0_u3_ch_txsz[12] , _u0_u3_ch_txsz[11] , _u0_u3_ch_txsz[10] ,_u0_u3_ch_txsz[9] , _u0_u3_ch_txsz[8] , _u0_u3_ch_txsz[7] ,_u0_u3_ch_txsz[6] , _u0_u3_ch_txsz[5] , _u0_u3_ch_txsz[4] ,_u0_u3_ch_txsz[3] , _u0_u3_ch_txsz[2] , _u0_u3_ch_txsz[1] ,_u0_u3_ch_txsz[0] , _u0_u3_ch_adr0[31] , _u0_u3_ch_adr0[30] ,_u0_u3_ch_adr0[29] , _u0_u3_ch_adr0[28] , _u0_u3_ch_adr0[27] ,_u0_u3_ch_adr0[26] , _u0_u3_ch_adr0[25] , _u0_u3_ch_adr0[24] ,_u0_u3_ch_adr0[23] , _u0_u3_ch_adr0[22] , _u0_u3_ch_adr0[21] ,_u0_u3_ch_adr0[20] , _u0_u3_ch_adr0[19] , _u0_u3_ch_adr0[18] ,_u0_u3_ch_adr0[17] , _u0_u3_ch_adr0[16] , _u0_u3_ch_adr0[15] ,_u0_u3_ch_adr0[14] , _u0_u3_ch_adr0[13] , _u0_u3_ch_adr0[12] ,_u0_u3_ch_adr0[11] , _u0_u3_ch_adr0[10] , _u0_u3_ch_adr0[9] ,_u0_u3_ch_adr0[8] , _u0_u3_ch_adr0[7] , _u0_u3_ch_adr0[6] ,_u0_u3_ch_adr0[5] , _u0_u3_ch_adr0[4] , _u0_u3_ch_adr0[3] ,_u0_u3_ch_adr0[2] , _u0_u3_ch_adr0[1] , _u0_u3_ch_adr0[0] ,_u0_u3_ch_adr1[31] , _u0_u3_ch_adr1[30] , _u0_u3_ch_adr1[29] ,_u0_u3_ch_adr1[28] , _u0_u3_ch_adr1[27] , _u0_u3_ch_adr1[26] ,_u0_u3_ch_adr1[25] , _u0_u3_ch_adr1[24] , _u0_u3_ch_adr1[23] ,_u0_u3_ch_adr1[22] , _u0_u3_ch_adr1[21] , _u0_u3_ch_adr1[20] ,_u0_u3_ch_adr1[19] , _u0_u3_ch_adr1[18] , _u0_u3_ch_adr1[17] ,_u0_u3_ch_adr1[16] , _u0_u3_ch_adr1[15] , _u0_u3_ch_adr1[14] ,_u0_u3_ch_adr1[13] , _u0_u3_ch_adr1[12] , _u0_u3_ch_adr1[11] ,_u0_u3_ch_adr1[10] , _u0_u3_ch_adr1[9] , _u0_u3_ch_adr1[8] ,_u0_u3_ch_adr1[7] , _u0_u3_ch_adr1[6] , _u0_u3_ch_adr1[5] ,_u0_u3_ch_adr1[4] , _u0_u3_ch_adr1[3] , _u0_u3_ch_adr1[2] ,_u0_u3_ch_adr1[1] , _u0_u3_ch_adr1[0] , _u0_u3_ch_am0[31] ,_u0_u3_ch_am0[30] , _u0_u3_ch_am0[29] , _u0_u3_ch_am0[28] ,_u0_u3_ch_am0[27] , _u0_u3_ch_am0[26] , _u0_u3_ch_am0[25] ,_u0_u3_ch_am0[24] , _u0_u3_ch_am0[23] , _u0_u3_ch_am0[22] ,_u0_u3_ch_am0[21] , _u0_u3_ch_am0[20] , _u0_u3_ch_am0[19] ,_u0_u3_ch_am0[18] , _u0_u3_ch_am0[17] , _u0_u3_ch_am0[16] ,_u0_u3_ch_am0[15] , _u0_u3_ch_am0[14] , _u0_u3_ch_am0[13] ,_u0_u3_ch_am0[12] , _u0_u3_ch_am0[11] , _u0_u3_ch_am0[10] ,_u0_u3_ch_am0[9] , _u0_u3_ch_am0[8] , _u0_u3_ch_am0[7] ,_u0_u3_ch_am0[6] , _u0_u3_ch_am0[5] , _u0_u3_ch_am0[4] ,_u0_u3_ch_am0[3] , _u0_u3_ch_am0[2] , _u0_u3_ch_am0[1] ,_u0_u3_ch_am0[0] , _u0_u3_ch_am1[31] , _u0_u3_ch_am1[30] ,_u0_u3_ch_am1[29] , _u0_u3_ch_am1[28] , _u0_u3_ch_am1[27] ,_u0_u3_ch_am1[26] , _u0_u3_ch_am1[25] , _u0_u3_ch_am1[24] ,_u0_u3_ch_am1[23] , _u0_u3_ch_am1[22] , _u0_u3_ch_am1[21] ,_u0_u3_ch_am1[20] , _u0_u3_ch_am1[19] , _u0_u3_ch_am1[18] ,_u0_u3_ch_am1[17] , _u0_u3_ch_am1[16] , _u0_u3_ch_am1[15] ,_u0_u3_ch_am1[14] , _u0_u3_ch_am1[13] , _u0_u3_ch_am1[12] ,_u0_u3_ch_am1[11] , _u0_u3_ch_am1[10] , _u0_u3_ch_am1[9] ,_u0_u3_ch_am1[8] , _u0_u3_ch_am1[7] , _u0_u3_ch_am1[6] ,_u0_u3_ch_am1[5] , _u0_u3_ch_am1[4] , _u0_u3_ch_am1[3] ,_u0_u3_ch_am1[2] , _u0_u3_ch_am1[1] , _u0_u3_ch_am1[0] ,_u0_u3_sw_pointer[31] , _u0_u3_sw_pointer[30] ,_u0_u3_sw_pointer[29] , _u0_u3_sw_pointer[28] ,_u0_u3_sw_pointer[27] , _u0_u3_sw_pointer[26] ,_u0_u3_sw_pointer[25] , _u0_u3_sw_pointer[24] ,_u0_u3_sw_pointer[23] , _u0_u3_sw_pointer[22] ,_u0_u3_sw_pointer[21] , _u0_u3_sw_pointer[20] ,_u0_u3_sw_pointer[19] , _u0_u3_sw_pointer[18] ,_u0_u3_sw_pointer[17] , _u0_u3_sw_pointer[16] ,_u0_u3_sw_pointer[15] , _u0_u3_sw_pointer[14] ,_u0_u3_sw_pointer[13] , _u0_u3_sw_pointer[12] ,_u0_u3_sw_pointer[11] , _u0_u3_sw_pointer[10] , _u0_u3_sw_pointer[9] ,_u0_u3_sw_pointer[8] , _u0_u3_sw_pointer[7] , _u0_u3_sw_pointer[6] ,_u0_u3_sw_pointer[5] , _u0_u3_sw_pointer[4] , _u0_u3_sw_pointer[3] ,_u0_u3_sw_pointer[2] , _u0_u3_sw_pointer[1] , _u0_u3_sw_pointer[0] ,_u0_u3_ch_stop , _u0_u3_ch_dis , _u0_u3_int , _u0_u4_pointer[31] ,_u0_u4_pointer[30] , _u0_u4_pointer[29] , _u0_u4_pointer[28] ,_u0_u4_pointer[27] , _u0_u4_pointer[26] , _u0_u4_pointer[25] ,_u0_u4_pointer[24] , _u0_u4_pointer[23] , _u0_u4_pointer[22] ,_u0_u4_pointer[21] , _u0_u4_pointer[20] , _u0_u4_pointer[19] ,_u0_u4_pointer[18] , _u0_u4_pointer[17] , _u0_u4_pointer[16] ,_u0_u4_pointer[15] , _u0_u4_pointer[14] , _u0_u4_pointer[13] ,_u0_u4_pointer[12] , _u0_u4_pointer[11] , _u0_u4_pointer[10] ,_u0_u4_pointer[9] , _u0_u4_pointer[8] , _u0_u4_pointer[7] ,_u0_u4_pointer[6] , _u0_u4_pointer[5] , _u0_u4_pointer[4] ,_u0_u4_pointer[3] , _u0_u4_pointer[2] , _u0_u4_pointer[1] ,_u0_u4_pointer[0] , _u0_u4_pointer_s[31] , _u0_u4_pointer_s[30] ,_u0_u4_pointer_s[29] , _u0_u4_pointer_s[28] , _u0_u4_pointer_s[27] ,_u0_u4_pointer_s[26] , _u0_u4_pointer_s[25] , _u0_u4_pointer_s[24] ,_u0_u4_pointer_s[23] , _u0_u4_pointer_s[22] , _u0_u4_pointer_s[21] ,_u0_u4_pointer_s[20] , _u0_u4_pointer_s[19] , _u0_u4_pointer_s[18] ,_u0_u4_pointer_s[17] , _u0_u4_pointer_s[16] , _u0_u4_pointer_s[15] ,_u0_u4_pointer_s[14] , _u0_u4_pointer_s[13] , _u0_u4_pointer_s[12] ,_u0_u4_pointer_s[11] , _u0_u4_pointer_s[10] , _u0_u4_pointer_s[9] ,_u0_u4_pointer_s[8] , _u0_u4_pointer_s[7] , _u0_u4_pointer_s[6] ,_u0_u4_pointer_s[5] , _u0_u4_pointer_s[4] , _u0_u4_pointer_s[3] ,_u0_u4_pointer_s[2] , _u0_u4_pointer_s[1] , _u0_u4_pointer_s[0] ,_u0_u4_ch_csr[31] , _u0_u4_ch_csr[30] , _u0_u4_ch_csr[29] ,_u0_u4_ch_csr[28] , _u0_u4_ch_csr[27] , _u0_u4_ch_csr[26] ,_u0_u4_ch_csr[25] , _u0_u4_ch_csr[24] , _u0_u4_ch_csr[23] ,_u0_u4_ch_csr[22] , _u0_u4_ch_csr[21] , _u0_u4_ch_csr[20] ,_u0_u4_ch_csr[19] , _u0_u4_ch_csr[18] , _u0_u4_ch_csr[17] ,_u0_u4_ch_csr[16] , _u0_u4_ch_csr[15] , _u0_u4_ch_csr[14] ,_u0_u4_ch_csr[13] , _u0_u4_ch_csr[12] , _u0_u4_ch_csr[11] ,_u0_u4_ch_csr[10] , _u0_u4_ch_csr[9] , _u0_u4_ch_csr[8] ,_u0_u4_ch_csr[7] , _u0_u4_ch_csr[6] , _u0_u4_ch_csr[5] ,_u0_u4_ch_csr[4] , _u0_u4_ch_csr[3] , _u0_u4_ch_csr[2] ,_u0_u4_ch_csr[1] , _u0_u4_ch_csr[0] , _u0_u4_ch_txsz[31] ,_u0_u4_ch_txsz[30] , _u0_u4_ch_txsz[29] , _u0_u4_ch_txsz[28] ,_u0_u4_ch_txsz[27] , _u0_u4_ch_txsz[26] , _u0_u4_ch_txsz[25] ,_u0_u4_ch_txsz[24] , _u0_u4_ch_txsz[23] , _u0_u4_ch_txsz[22] ,_u0_u4_ch_txsz[21] , _u0_u4_ch_txsz[20] , _u0_u4_ch_txsz[19] ,_u0_u4_ch_txsz[18] , _u0_u4_ch_txsz[17] , _u0_u4_ch_txsz[16] ,_u0_u4_ch_txsz[15] , _u0_u4_ch_txsz[14] , _u0_u4_ch_txsz[13] ,_u0_u4_ch_txsz[12] , _u0_u4_ch_txsz[11] , _u0_u4_ch_txsz[10] ,_u0_u4_ch_txsz[9] , _u0_u4_ch_txsz[8] , _u0_u4_ch_txsz[7] ,_u0_u4_ch_txsz[6] , _u0_u4_ch_txsz[5] , _u0_u4_ch_txsz[4] ,_u0_u4_ch_txsz[3] , _u0_u4_ch_txsz[2] , _u0_u4_ch_txsz[1] ,_u0_u4_ch_txsz[0] , _u0_u4_ch_adr0[31] , _u0_u4_ch_adr0[30] ,_u0_u4_ch_adr0[29] , _u0_u4_ch_adr0[28] , _u0_u4_ch_adr0[27] ,_u0_u4_ch_adr0[26] , _u0_u4_ch_adr0[25] , _u0_u4_ch_adr0[24] ,_u0_u4_ch_adr0[23] , _u0_u4_ch_adr0[22] , _u0_u4_ch_adr0[21] ,_u0_u4_ch_adr0[20] , _u0_u4_ch_adr0[19] , _u0_u4_ch_adr0[18] ,_u0_u4_ch_adr0[17] , _u0_u4_ch_adr0[16] , _u0_u4_ch_adr0[15] ,_u0_u4_ch_adr0[14] , _u0_u4_ch_adr0[13] , _u0_u4_ch_adr0[12] ,_u0_u4_ch_adr0[11] , _u0_u4_ch_adr0[10] , _u0_u4_ch_adr0[9] ,_u0_u4_ch_adr0[8] , _u0_u4_ch_adr0[7] , _u0_u4_ch_adr0[6] ,_u0_u4_ch_adr0[5] , _u0_u4_ch_adr0[4] , _u0_u4_ch_adr0[3] ,_u0_u4_ch_adr0[2] , _u0_u4_ch_adr0[1] , _u0_u4_ch_adr0[0] ,_u0_u4_ch_adr1[31] , _u0_u4_ch_adr1[30] , _u0_u4_ch_adr1[29] ,_u0_u4_ch_adr1[28] , _u0_u4_ch_adr1[27] , _u0_u4_ch_adr1[26] ,_u0_u4_ch_adr1[25] , _u0_u4_ch_adr1[24] , _u0_u4_ch_adr1[23] ,_u0_u4_ch_adr1[22] , _u0_u4_ch_adr1[21] , _u0_u4_ch_adr1[20] ,_u0_u4_ch_adr1[19] , _u0_u4_ch_adr1[18] , _u0_u4_ch_adr1[17] ,_u0_u4_ch_adr1[16] , _u0_u4_ch_adr1[15] , _u0_u4_ch_adr1[14] ,_u0_u4_ch_adr1[13] , _u0_u4_ch_adr1[12] , _u0_u4_ch_adr1[11] ,_u0_u4_ch_adr1[10] , _u0_u4_ch_adr1[9] , _u0_u4_ch_adr1[8] ,_u0_u4_ch_adr1[7] , _u0_u4_ch_adr1[6] , _u0_u4_ch_adr1[5] ,_u0_u4_ch_adr1[4] , _u0_u4_ch_adr1[3] , _u0_u4_ch_adr1[2] ,_u0_u4_ch_adr1[1] , _u0_u4_ch_adr1[0] , _u0_u4_ch_am0[31] ,_u0_u4_ch_am0[30] , _u0_u4_ch_am0[29] , _u0_u4_ch_am0[28] ,_u0_u4_ch_am0[27] , _u0_u4_ch_am0[26] , _u0_u4_ch_am0[25] ,_u0_u4_ch_am0[24] , _u0_u4_ch_am0[23] , _u0_u4_ch_am0[22] ,_u0_u4_ch_am0[21] , _u0_u4_ch_am0[20] , _u0_u4_ch_am0[19] ,_u0_u4_ch_am0[18] , _u0_u4_ch_am0[17] , _u0_u4_ch_am0[16] ,_u0_u4_ch_am0[15] , _u0_u4_ch_am0[14] , _u0_u4_ch_am0[13] ,_u0_u4_ch_am0[12] , _u0_u4_ch_am0[11] , _u0_u4_ch_am0[10] ,_u0_u4_ch_am0[9] , _u0_u4_ch_am0[8] , _u0_u4_ch_am0[7] ,_u0_u4_ch_am0[6] , _u0_u4_ch_am0[5] , _u0_u4_ch_am0[4] ,_u0_u4_ch_am0[3] , _u0_u4_ch_am0[2] , _u0_u4_ch_am0[1] ,_u0_u4_ch_am0[0] , _u0_u4_ch_am1[31] , _u0_u4_ch_am1[30] ,_u0_u4_ch_am1[29] , _u0_u4_ch_am1[28] , _u0_u4_ch_am1[27] ,_u0_u4_ch_am1[26] , _u0_u4_ch_am1[25] , _u0_u4_ch_am1[24] ,_u0_u4_ch_am1[23] , _u0_u4_ch_am1[22] , _u0_u4_ch_am1[21] ,_u0_u4_ch_am1[20] , _u0_u4_ch_am1[19] , _u0_u4_ch_am1[18] ,_u0_u4_ch_am1[17] , _u0_u4_ch_am1[16] , _u0_u4_ch_am1[15] ,_u0_u4_ch_am1[14] , _u0_u4_ch_am1[13] , _u0_u4_ch_am1[12] ,_u0_u4_ch_am1[11] , _u0_u4_ch_am1[10] , _u0_u4_ch_am1[9] ,_u0_u4_ch_am1[8] , _u0_u4_ch_am1[7] , _u0_u4_ch_am1[6] ,_u0_u4_ch_am1[5] , _u0_u4_ch_am1[4] , _u0_u4_ch_am1[3] ,_u0_u4_ch_am1[2] , _u0_u4_ch_am1[1] , _u0_u4_ch_am1[0] ,_u0_u4_sw_pointer[31] , _u0_u4_sw_pointer[30] ,_u0_u4_sw_pointer[29] , _u0_u4_sw_pointer[28] ,_u0_u4_sw_pointer[27] , _u0_u4_sw_pointer[26] ,_u0_u4_sw_pointer[25] , _u0_u4_sw_pointer[24] ,_u0_u4_sw_pointer[23] , _u0_u4_sw_pointer[22] ,_u0_u4_sw_pointer[21] , _u0_u4_sw_pointer[20] ,_u0_u4_sw_pointer[19] , _u0_u4_sw_pointer[18] ,_u0_u4_sw_pointer[17] , _u0_u4_sw_pointer[16] ,_u0_u4_sw_pointer[15] , _u0_u4_sw_pointer[14] ,_u0_u4_sw_pointer[13] , _u0_u4_sw_pointer[12] ,_u0_u4_sw_pointer[11] , _u0_u4_sw_pointer[10] , _u0_u4_sw_pointer[9] ,_u0_u4_sw_pointer[8] , _u0_u4_sw_pointer[7] , _u0_u4_sw_pointer[6] ,_u0_u4_sw_pointer[5] , _u0_u4_sw_pointer[4] , _u0_u4_sw_pointer[3] ,_u0_u4_sw_pointer[2] , _u0_u4_sw_pointer[1] , _u0_u4_sw_pointer[0] ,_u0_u4_ch_stop , _u0_u4_ch_dis , _u0_u4_int , _u0_u5_pointer[31] ,_u0_u5_pointer[30] , _u0_u5_pointer[29] , _u0_u5_pointer[28] ,_u0_u5_pointer[27] , _u0_u5_pointer[26] , _u0_u5_pointer[25] ,_u0_u5_pointer[24] , _u0_u5_pointer[23] , _u0_u5_pointer[22] ,_u0_u5_pointer[21] , _u0_u5_pointer[20] , _u0_u5_pointer[19] ,_u0_u5_pointer[18] , _u0_u5_pointer[17] , _u0_u5_pointer[16] ,_u0_u5_pointer[15] , _u0_u5_pointer[14] , _u0_u5_pointer[13] ,_u0_u5_pointer[12] , _u0_u5_pointer[11] , _u0_u5_pointer[10] ,_u0_u5_pointer[9] , _u0_u5_pointer[8] , _u0_u5_pointer[7] ,_u0_u5_pointer[6] , _u0_u5_pointer[5] , _u0_u5_pointer[4] ,_u0_u5_pointer[3] , _u0_u5_pointer[2] , _u0_u5_pointer[1] ,_u0_u5_pointer[0] , _u0_u5_pointer_s[31] , _u0_u5_pointer_s[30] ,_u0_u5_pointer_s[29] , _u0_u5_pointer_s[28] , _u0_u5_pointer_s[27] ,_u0_u5_pointer_s[26] , _u0_u5_pointer_s[25] , _u0_u5_pointer_s[24] ,_u0_u5_pointer_s[23] , _u0_u5_pointer_s[22] , _u0_u5_pointer_s[21] ,_u0_u5_pointer_s[20] , _u0_u5_pointer_s[19] , _u0_u5_pointer_s[18] ,_u0_u5_pointer_s[17] , _u0_u5_pointer_s[16] , _u0_u5_pointer_s[15] ,_u0_u5_pointer_s[14] , _u0_u5_pointer_s[13] , _u0_u5_pointer_s[12] ,_u0_u5_pointer_s[11] , _u0_u5_pointer_s[10] , _u0_u5_pointer_s[9] ,_u0_u5_pointer_s[8] , _u0_u5_pointer_s[7] , _u0_u5_pointer_s[6] ,_u0_u5_pointer_s[5] , _u0_u5_pointer_s[4] , _u0_u5_pointer_s[3] ,_u0_u5_pointer_s[2] , _u0_u5_pointer_s[1] , _u0_u5_pointer_s[0] ,_u0_u5_ch_csr[31] , _u0_u5_ch_csr[30] , _u0_u5_ch_csr[29] ,_u0_u5_ch_csr[28] , _u0_u5_ch_csr[27] , _u0_u5_ch_csr[26] ,_u0_u5_ch_csr[25] , _u0_u5_ch_csr[24] , _u0_u5_ch_csr[23] ,_u0_u5_ch_csr[22] , _u0_u5_ch_csr[21] , _u0_u5_ch_csr[20] ,_u0_u5_ch_csr[19] , _u0_u5_ch_csr[18] , _u0_u5_ch_csr[17] ,_u0_u5_ch_csr[16] , _u0_u5_ch_csr[15] , _u0_u5_ch_csr[14] ,_u0_u5_ch_csr[13] , _u0_u5_ch_csr[12] , _u0_u5_ch_csr[11] ,_u0_u5_ch_csr[10] , _u0_u5_ch_csr[9] , _u0_u5_ch_csr[8] ,_u0_u5_ch_csr[7] , _u0_u5_ch_csr[6] , _u0_u5_ch_csr[5] ,_u0_u5_ch_csr[4] , _u0_u5_ch_csr[3] , _u0_u5_ch_csr[2] ,_u0_u5_ch_csr[1] , _u0_u5_ch_csr[0] , _u0_u5_ch_txsz[31] ,_u0_u5_ch_txsz[30] , _u0_u5_ch_txsz[29] , _u0_u5_ch_txsz[28] ,_u0_u5_ch_txsz[27] , _u0_u5_ch_txsz[26] , _u0_u5_ch_txsz[25] ,_u0_u5_ch_txsz[24] , _u0_u5_ch_txsz[23] , _u0_u5_ch_txsz[22] ,_u0_u5_ch_txsz[21] , _u0_u5_ch_txsz[20] , _u0_u5_ch_txsz[19] ,_u0_u5_ch_txsz[18] , _u0_u5_ch_txsz[17] , _u0_u5_ch_txsz[16] ,_u0_u5_ch_txsz[15] , _u0_u5_ch_txsz[14] , _u0_u5_ch_txsz[13] ,_u0_u5_ch_txsz[12] , _u0_u5_ch_txsz[11] , _u0_u5_ch_txsz[10] ,_u0_u5_ch_txsz[9] , _u0_u5_ch_txsz[8] , _u0_u5_ch_txsz[7] ,_u0_u5_ch_txsz[6] , _u0_u5_ch_txsz[5] , _u0_u5_ch_txsz[4] ,_u0_u5_ch_txsz[3] , _u0_u5_ch_txsz[2] , _u0_u5_ch_txsz[1] ,_u0_u5_ch_txsz[0] , _u0_u5_ch_adr0[31] , _u0_u5_ch_adr0[30] ,_u0_u5_ch_adr0[29] , _u0_u5_ch_adr0[28] , _u0_u5_ch_adr0[27] ,_u0_u5_ch_adr0[26] , _u0_u5_ch_adr0[25] , _u0_u5_ch_adr0[24] ,_u0_u5_ch_adr0[23] , _u0_u5_ch_adr0[22] , _u0_u5_ch_adr0[21] ,_u0_u5_ch_adr0[20] , _u0_u5_ch_adr0[19] , _u0_u5_ch_adr0[18] ,_u0_u5_ch_adr0[17] , _u0_u5_ch_adr0[16] , _u0_u5_ch_adr0[15] ,_u0_u5_ch_adr0[14] , _u0_u5_ch_adr0[13] , _u0_u5_ch_adr0[12] ,_u0_u5_ch_adr0[11] , _u0_u5_ch_adr0[10] , _u0_u5_ch_adr0[9] ,_u0_u5_ch_adr0[8] , _u0_u5_ch_adr0[7] , _u0_u5_ch_adr0[6] ,_u0_u5_ch_adr0[5] , _u0_u5_ch_adr0[4] , _u0_u5_ch_adr0[3] ,_u0_u5_ch_adr0[2] , _u0_u5_ch_adr0[1] , _u0_u5_ch_adr0[0] ,_u0_u5_ch_adr1[31] , _u0_u5_ch_adr1[30] , _u0_u5_ch_adr1[29] ,_u0_u5_ch_adr1[28] , _u0_u5_ch_adr1[27] , _u0_u5_ch_adr1[26] ,_u0_u5_ch_adr1[25] , _u0_u5_ch_adr1[24] , _u0_u5_ch_adr1[23] ,_u0_u5_ch_adr1[22] , _u0_u5_ch_adr1[21] , _u0_u5_ch_adr1[20] ,_u0_u5_ch_adr1[19] , _u0_u5_ch_adr1[18] , _u0_u5_ch_adr1[17] ,_u0_u5_ch_adr1[16] , _u0_u5_ch_adr1[15] , _u0_u5_ch_adr1[14] ,_u0_u5_ch_adr1[13] , _u0_u5_ch_adr1[12] , _u0_u5_ch_adr1[11] ,_u0_u5_ch_adr1[10] , _u0_u5_ch_adr1[9] , _u0_u5_ch_adr1[8] ,_u0_u5_ch_adr1[7] , _u0_u5_ch_adr1[6] , _u0_u5_ch_adr1[5] ,_u0_u5_ch_adr1[4] , _u0_u5_ch_adr1[3] , _u0_u5_ch_adr1[2] ,_u0_u5_ch_adr1[1] , _u0_u5_ch_adr1[0] , _u0_u5_ch_am0[31] ,_u0_u5_ch_am0[30] , _u0_u5_ch_am0[29] , _u0_u5_ch_am0[28] ,_u0_u5_ch_am0[27] , _u0_u5_ch_am0[26] , _u0_u5_ch_am0[25] ,_u0_u5_ch_am0[24] , _u0_u5_ch_am0[23] , _u0_u5_ch_am0[22] ,_u0_u5_ch_am0[21] , _u0_u5_ch_am0[20] , _u0_u5_ch_am0[19] ,_u0_u5_ch_am0[18] , _u0_u5_ch_am0[17] , _u0_u5_ch_am0[16] ,_u0_u5_ch_am0[15] , _u0_u5_ch_am0[14] , _u0_u5_ch_am0[13] ,_u0_u5_ch_am0[12] , _u0_u5_ch_am0[11] , _u0_u5_ch_am0[10] ,_u0_u5_ch_am0[9] , _u0_u5_ch_am0[8] , _u0_u5_ch_am0[7] ,_u0_u5_ch_am0[6] , _u0_u5_ch_am0[5] , _u0_u5_ch_am0[4] ,_u0_u5_ch_am0[3] , _u0_u5_ch_am0[2] , _u0_u5_ch_am0[1] ,_u0_u5_ch_am0[0] , _u0_u5_ch_am1[31] , _u0_u5_ch_am1[30] ,_u0_u5_ch_am1[29] , _u0_u5_ch_am1[28] , _u0_u5_ch_am1[27] ,_u0_u5_ch_am1[26] , _u0_u5_ch_am1[25] , _u0_u5_ch_am1[24] ,_u0_u5_ch_am1[23] , _u0_u5_ch_am1[22] , _u0_u5_ch_am1[21] ,_u0_u5_ch_am1[20] , _u0_u5_ch_am1[19] , _u0_u5_ch_am1[18] ,_u0_u5_ch_am1[17] , _u0_u5_ch_am1[16] , _u0_u5_ch_am1[15] ,_u0_u5_ch_am1[14] , _u0_u5_ch_am1[13] , _u0_u5_ch_am1[12] ,_u0_u5_ch_am1[11] , _u0_u5_ch_am1[10] , _u0_u5_ch_am1[9] ,_u0_u5_ch_am1[8] , _u0_u5_ch_am1[7] , _u0_u5_ch_am1[6] ,_u0_u5_ch_am1[5] , _u0_u5_ch_am1[4] , _u0_u5_ch_am1[3] ,_u0_u5_ch_am1[2] , _u0_u5_ch_am1[1] , _u0_u5_ch_am1[0] ,_u0_u5_sw_pointer[31] , _u0_u5_sw_pointer[30] ,_u0_u5_sw_pointer[29] , _u0_u5_sw_pointer[28] ,_u0_u5_sw_pointer[27] , _u0_u5_sw_pointer[26] ,_u0_u5_sw_pointer[25] , _u0_u5_sw_pointer[24] ,_u0_u5_sw_pointer[23] , _u0_u5_sw_pointer[22] ,_u0_u5_sw_pointer[21] , _u0_u5_sw_pointer[20] ,_u0_u5_sw_pointer[19] , _u0_u5_sw_pointer[18] ,_u0_u5_sw_pointer[17] , _u0_u5_sw_pointer[16] ,_u0_u5_sw_pointer[15] , _u0_u5_sw_pointer[14] ,_u0_u5_sw_pointer[13] , _u0_u5_sw_pointer[12] ,_u0_u5_sw_pointer[11] , _u0_u5_sw_pointer[10] , _u0_u5_sw_pointer[9] ,_u0_u5_sw_pointer[8] , _u0_u5_sw_pointer[7] , _u0_u5_sw_pointer[6] ,_u0_u5_sw_pointer[5] , _u0_u5_sw_pointer[4] , _u0_u5_sw_pointer[3] ,_u0_u5_sw_pointer[2] , _u0_u5_sw_pointer[1] , _u0_u5_sw_pointer[0] ,_u0_u5_ch_stop , _u0_u5_ch_dis , _u0_u5_int , _u0_u6_pointer[31] ,_u0_u6_pointer[30] , _u0_u6_pointer[29] , _u0_u6_pointer[28] ,_u0_u6_pointer[27] , _u0_u6_pointer[26] , _u0_u6_pointer[25] ,_u0_u6_pointer[24] , _u0_u6_pointer[23] , _u0_u6_pointer[22] ,_u0_u6_pointer[21] , _u0_u6_pointer[20] , _u0_u6_pointer[19] ,_u0_u6_pointer[18] , _u0_u6_pointer[17] , _u0_u6_pointer[16] ,_u0_u6_pointer[15] , _u0_u6_pointer[14] , _u0_u6_pointer[13] ,_u0_u6_pointer[12] , _u0_u6_pointer[11] , _u0_u6_pointer[10] ,_u0_u6_pointer[9] , _u0_u6_pointer[8] , _u0_u6_pointer[7] ,_u0_u6_pointer[6] , _u0_u6_pointer[5] , _u0_u6_pointer[4] ,_u0_u6_pointer[3] , _u0_u6_pointer[2] , _u0_u6_pointer[1] ,_u0_u6_pointer[0] , _u0_u6_pointer_s[31] , _u0_u6_pointer_s[30] ,_u0_u6_pointer_s[29] , _u0_u6_pointer_s[28] , _u0_u6_pointer_s[27] ,_u0_u6_pointer_s[26] , _u0_u6_pointer_s[25] , _u0_u6_pointer_s[24] ,_u0_u6_pointer_s[23] , _u0_u6_pointer_s[22] , _u0_u6_pointer_s[21] ,_u0_u6_pointer_s[20] , _u0_u6_pointer_s[19] , _u0_u6_pointer_s[18] ,_u0_u6_pointer_s[17] , _u0_u6_pointer_s[16] , _u0_u6_pointer_s[15] ,_u0_u6_pointer_s[14] , _u0_u6_pointer_s[13] , _u0_u6_pointer_s[12] ,_u0_u6_pointer_s[11] , _u0_u6_pointer_s[10] , _u0_u6_pointer_s[9] ,_u0_u6_pointer_s[8] , _u0_u6_pointer_s[7] , _u0_u6_pointer_s[6] ,_u0_u6_pointer_s[5] , _u0_u6_pointer_s[4] , _u0_u6_pointer_s[3] ,_u0_u6_pointer_s[2] , _u0_u6_pointer_s[1] , _u0_u6_pointer_s[0] ,_u0_u6_ch_csr[31] , _u0_u6_ch_csr[30] , _u0_u6_ch_csr[29] ,_u0_u6_ch_csr[28] , _u0_u6_ch_csr[27] , _u0_u6_ch_csr[26] ,_u0_u6_ch_csr[25] , _u0_u6_ch_csr[24] , _u0_u6_ch_csr[23] ,_u0_u6_ch_csr[22] , _u0_u6_ch_csr[21] , _u0_u6_ch_csr[20] ,_u0_u6_ch_csr[19] , _u0_u6_ch_csr[18] , _u0_u6_ch_csr[17] ,_u0_u6_ch_csr[16] , _u0_u6_ch_csr[15] , _u0_u6_ch_csr[14] ,_u0_u6_ch_csr[13] , _u0_u6_ch_csr[12] , _u0_u6_ch_csr[11] ,_u0_u6_ch_csr[10] , _u0_u6_ch_csr[9] , _u0_u6_ch_csr[8] ,_u0_u6_ch_csr[7] , _u0_u6_ch_csr[6] , _u0_u6_ch_csr[5] ,_u0_u6_ch_csr[4] , _u0_u6_ch_csr[3] , _u0_u6_ch_csr[2] ,_u0_u6_ch_csr[1] , _u0_u6_ch_csr[0] , _u0_u6_ch_txsz[31] ,_u0_u6_ch_txsz[30] , _u0_u6_ch_txsz[29] , _u0_u6_ch_txsz[28] ,_u0_u6_ch_txsz[27] , _u0_u6_ch_txsz[26] , _u0_u6_ch_txsz[25] ,_u0_u6_ch_txsz[24] , _u0_u6_ch_txsz[23] , _u0_u6_ch_txsz[22] ,_u0_u6_ch_txsz[21] , _u0_u6_ch_txsz[20] , _u0_u6_ch_txsz[19] ,_u0_u6_ch_txsz[18] , _u0_u6_ch_txsz[17] , _u0_u6_ch_txsz[16] ,_u0_u6_ch_txsz[15] , _u0_u6_ch_txsz[14] , _u0_u6_ch_txsz[13] ,_u0_u6_ch_txsz[12] , _u0_u6_ch_txsz[11] , _u0_u6_ch_txsz[10] ,_u0_u6_ch_txsz[9] , _u0_u6_ch_txsz[8] , _u0_u6_ch_txsz[7] ,_u0_u6_ch_txsz[6] , _u0_u6_ch_txsz[5] , _u0_u6_ch_txsz[4] ,_u0_u6_ch_txsz[3] , _u0_u6_ch_txsz[2] , _u0_u6_ch_txsz[1] ,_u0_u6_ch_txsz[0] , _u0_u6_ch_adr0[31] , _u0_u6_ch_adr0[30] ,_u0_u6_ch_adr0[29] , _u0_u6_ch_adr0[28] , _u0_u6_ch_adr0[27] ,_u0_u6_ch_adr0[26] , _u0_u6_ch_adr0[25] , _u0_u6_ch_adr0[24] ,_u0_u6_ch_adr0[23] , _u0_u6_ch_adr0[22] , _u0_u6_ch_adr0[21] ,_u0_u6_ch_adr0[20] , _u0_u6_ch_adr0[19] , _u0_u6_ch_adr0[18] ,_u0_u6_ch_adr0[17] , _u0_u6_ch_adr0[16] , _u0_u6_ch_adr0[15] ,_u0_u6_ch_adr0[14] , _u0_u6_ch_adr0[13] , _u0_u6_ch_adr0[12] ,_u0_u6_ch_adr0[11] , _u0_u6_ch_adr0[10] , _u0_u6_ch_adr0[9] ,_u0_u6_ch_adr0[8] , _u0_u6_ch_adr0[7] , _u0_u6_ch_adr0[6] ,_u0_u6_ch_adr0[5] , _u0_u6_ch_adr0[4] , _u0_u6_ch_adr0[3] ,_u0_u6_ch_adr0[2] , _u0_u6_ch_adr0[1] , _u0_u6_ch_adr0[0] ,_u0_u6_ch_adr1[31] , _u0_u6_ch_adr1[30] , _u0_u6_ch_adr1[29] ,_u0_u6_ch_adr1[28] , _u0_u6_ch_adr1[27] , _u0_u6_ch_adr1[26] ,_u0_u6_ch_adr1[25] , _u0_u6_ch_adr1[24] , _u0_u6_ch_adr1[23] ,_u0_u6_ch_adr1[22] , _u0_u6_ch_adr1[21] , _u0_u6_ch_adr1[20] ,_u0_u6_ch_adr1[19] , _u0_u6_ch_adr1[18] , _u0_u6_ch_adr1[17] ,_u0_u6_ch_adr1[16] , _u0_u6_ch_adr1[15] , _u0_u6_ch_adr1[14] ,_u0_u6_ch_adr1[13] , _u0_u6_ch_adr1[12] , _u0_u6_ch_adr1[11] ,_u0_u6_ch_adr1[10] , _u0_u6_ch_adr1[9] , _u0_u6_ch_adr1[8] ,_u0_u6_ch_adr1[7] , _u0_u6_ch_adr1[6] , _u0_u6_ch_adr1[5] ,_u0_u6_ch_adr1[4] , _u0_u6_ch_adr1[3] , _u0_u6_ch_adr1[2] ,_u0_u6_ch_adr1[1] , _u0_u6_ch_adr1[0] , _u0_u6_ch_am0[31] ,_u0_u6_ch_am0[30] , _u0_u6_ch_am0[29] , _u0_u6_ch_am0[28] ,_u0_u6_ch_am0[27] , _u0_u6_ch_am0[26] , _u0_u6_ch_am0[25] ,_u0_u6_ch_am0[24] , _u0_u6_ch_am0[23] , _u0_u6_ch_am0[22] ,_u0_u6_ch_am0[21] , _u0_u6_ch_am0[20] , _u0_u6_ch_am0[19] ,_u0_u6_ch_am0[18] , _u0_u6_ch_am0[17] , _u0_u6_ch_am0[16] ,_u0_u6_ch_am0[15] , _u0_u6_ch_am0[14] , _u0_u6_ch_am0[13] ,_u0_u6_ch_am0[12] , _u0_u6_ch_am0[11] , _u0_u6_ch_am0[10] ,_u0_u6_ch_am0[9] , _u0_u6_ch_am0[8] , _u0_u6_ch_am0[7] ,_u0_u6_ch_am0[6] , _u0_u6_ch_am0[5] , _u0_u6_ch_am0[4] ,_u0_u6_ch_am0[3] , _u0_u6_ch_am0[2] , _u0_u6_ch_am0[1] ,_u0_u6_ch_am0[0] , _u0_u6_ch_am1[31] , _u0_u6_ch_am1[30] ,_u0_u6_ch_am1[29] , _u0_u6_ch_am1[28] , _u0_u6_ch_am1[27] ,_u0_u6_ch_am1[26] , _u0_u6_ch_am1[25] , _u0_u6_ch_am1[24] ,_u0_u6_ch_am1[23] , _u0_u6_ch_am1[22] , _u0_u6_ch_am1[21] ,_u0_u6_ch_am1[20] , _u0_u6_ch_am1[19] , _u0_u6_ch_am1[18] ,_u0_u6_ch_am1[17] , _u0_u6_ch_am1[16] , _u0_u6_ch_am1[15] ,_u0_u6_ch_am1[14] , _u0_u6_ch_am1[13] , _u0_u6_ch_am1[12] ,_u0_u6_ch_am1[11] , _u0_u6_ch_am1[10] , _u0_u6_ch_am1[9] ,_u0_u6_ch_am1[8] , _u0_u6_ch_am1[7] , _u0_u6_ch_am1[6] ,_u0_u6_ch_am1[5] , _u0_u6_ch_am1[4] , _u0_u6_ch_am1[3] ,_u0_u6_ch_am1[2] , _u0_u6_ch_am1[1] , _u0_u6_ch_am1[0] ,_u0_u6_sw_pointer[31] , _u0_u6_sw_pointer[30] ,_u0_u6_sw_pointer[29] , _u0_u6_sw_pointer[28] ,_u0_u6_sw_pointer[27] , _u0_u6_sw_pointer[26] ,_u0_u6_sw_pointer[25] , _u0_u6_sw_pointer[24] ,_u0_u6_sw_pointer[23] , _u0_u6_sw_pointer[22] ,_u0_u6_sw_pointer[21] , _u0_u6_sw_pointer[20] ,_u0_u6_sw_pointer[19] , _u0_u6_sw_pointer[18] ,_u0_u6_sw_pointer[17] , _u0_u6_sw_pointer[16] ,_u0_u6_sw_pointer[15] , _u0_u6_sw_pointer[14] ,_u0_u6_sw_pointer[13] , _u0_u6_sw_pointer[12] ,_u0_u6_sw_pointer[11] , _u0_u6_sw_pointer[10] , _u0_u6_sw_pointer[9] ,_u0_u6_sw_pointer[8] , _u0_u6_sw_pointer[7] , _u0_u6_sw_pointer[6] ,_u0_u6_sw_pointer[5] , _u0_u6_sw_pointer[4] , _u0_u6_sw_pointer[3] ,_u0_u6_sw_pointer[2] , _u0_u6_sw_pointer[1] , _u0_u6_sw_pointer[0] ,_u0_u6_ch_stop , _u0_u6_ch_dis , _u0_u6_int , _u0_u7_pointer[31] ,_u0_u7_pointer[30] , _u0_u7_pointer[29] , _u0_u7_pointer[28] ,_u0_u7_pointer[27] , _u0_u7_pointer[26] , _u0_u7_pointer[25] ,_u0_u7_pointer[24] , _u0_u7_pointer[23] , _u0_u7_pointer[22] ,_u0_u7_pointer[21] , _u0_u7_pointer[20] , _u0_u7_pointer[19] ,_u0_u7_pointer[18] , _u0_u7_pointer[17] , _u0_u7_pointer[16] ,_u0_u7_pointer[15] , _u0_u7_pointer[14] , _u0_u7_pointer[13] ,_u0_u7_pointer[12] , _u0_u7_pointer[11] , _u0_u7_pointer[10] ,_u0_u7_pointer[9] , _u0_u7_pointer[8] , _u0_u7_pointer[7] ,_u0_u7_pointer[6] , _u0_u7_pointer[5] , _u0_u7_pointer[4] ,_u0_u7_pointer[3] , _u0_u7_pointer[2] , _u0_u7_pointer[1] ,_u0_u7_pointer[0] , _u0_u7_pointer_s[31] , _u0_u7_pointer_s[30] ,_u0_u7_pointer_s[29] , _u0_u7_pointer_s[28] , _u0_u7_pointer_s[27] ,_u0_u7_pointer_s[26] , _u0_u7_pointer_s[25] , _u0_u7_pointer_s[24] ,_u0_u7_pointer_s[23] , _u0_u7_pointer_s[22] , _u0_u7_pointer_s[21] ,_u0_u7_pointer_s[20] , _u0_u7_pointer_s[19] , _u0_u7_pointer_s[18] ,_u0_u7_pointer_s[17] , _u0_u7_pointer_s[16] , _u0_u7_pointer_s[15] ,_u0_u7_pointer_s[14] , _u0_u7_pointer_s[13] , _u0_u7_pointer_s[12] ,_u0_u7_pointer_s[11] , _u0_u7_pointer_s[10] , _u0_u7_pointer_s[9] ,_u0_u7_pointer_s[8] , _u0_u7_pointer_s[7] , _u0_u7_pointer_s[6] ,_u0_u7_pointer_s[5] , _u0_u7_pointer_s[4] , _u0_u7_pointer_s[3] ,_u0_u7_pointer_s[2] , _u0_u7_pointer_s[1] , _u0_u7_pointer_s[0] ,_u0_u7_ch_csr[31] , _u0_u7_ch_csr[30] , _u0_u7_ch_csr[29] ,_u0_u7_ch_csr[28] , _u0_u7_ch_csr[27] , _u0_u7_ch_csr[26] ,_u0_u7_ch_csr[25] , _u0_u7_ch_csr[24] , _u0_u7_ch_csr[23] ,_u0_u7_ch_csr[22] , _u0_u7_ch_csr[21] , _u0_u7_ch_csr[20] ,_u0_u7_ch_csr[19] , _u0_u7_ch_csr[18] , _u0_u7_ch_csr[17] ,_u0_u7_ch_csr[16] , _u0_u7_ch_csr[15] , _u0_u7_ch_csr[14] ,_u0_u7_ch_csr[13] , _u0_u7_ch_csr[12] , _u0_u7_ch_csr[11] ,_u0_u7_ch_csr[10] , _u0_u7_ch_csr[9] , _u0_u7_ch_csr[8] ,_u0_u7_ch_csr[7] , _u0_u7_ch_csr[6] , _u0_u7_ch_csr[5] ,_u0_u7_ch_csr[4] , _u0_u7_ch_csr[3] , _u0_u7_ch_csr[2] ,_u0_u7_ch_csr[1] , _u0_u7_ch_csr[0] , _u0_u7_ch_txsz[31] ,_u0_u7_ch_txsz[30] , _u0_u7_ch_txsz[29] , _u0_u7_ch_txsz[28] ,_u0_u7_ch_txsz[27] , _u0_u7_ch_txsz[26] , _u0_u7_ch_txsz[25] ,_u0_u7_ch_txsz[24] , _u0_u7_ch_txsz[23] , _u0_u7_ch_txsz[22] ,_u0_u7_ch_txsz[21] , _u0_u7_ch_txsz[20] , _u0_u7_ch_txsz[19] ,_u0_u7_ch_txsz[18] , _u0_u7_ch_txsz[17] , _u0_u7_ch_txsz[16] ,_u0_u7_ch_txsz[15] , _u0_u7_ch_txsz[14] , _u0_u7_ch_txsz[13] ,_u0_u7_ch_txsz[12] , _u0_u7_ch_txsz[11] , _u0_u7_ch_txsz[10] ,_u0_u7_ch_txsz[9] , _u0_u7_ch_txsz[8] , _u0_u7_ch_txsz[7] ,_u0_u7_ch_txsz[6] , _u0_u7_ch_txsz[5] , _u0_u7_ch_txsz[4] ,_u0_u7_ch_txsz[3] , _u0_u7_ch_txsz[2] , _u0_u7_ch_txsz[1] ,_u0_u7_ch_txsz[0] , _u0_u7_ch_adr0[31] , _u0_u7_ch_adr0[30] ,_u0_u7_ch_adr0[29] , _u0_u7_ch_adr0[28] , _u0_u7_ch_adr0[27] ,_u0_u7_ch_adr0[26] , _u0_u7_ch_adr0[25] , _u0_u7_ch_adr0[24] ,_u0_u7_ch_adr0[23] , _u0_u7_ch_adr0[22] , _u0_u7_ch_adr0[21] ,_u0_u7_ch_adr0[20] , _u0_u7_ch_adr0[19] , _u0_u7_ch_adr0[18] ,_u0_u7_ch_adr0[17] , _u0_u7_ch_adr0[16] , _u0_u7_ch_adr0[15] ,_u0_u7_ch_adr0[14] , _u0_u7_ch_adr0[13] , _u0_u7_ch_adr0[12] ,_u0_u7_ch_adr0[11] , _u0_u7_ch_adr0[10] , _u0_u7_ch_adr0[9] ,_u0_u7_ch_adr0[8] , _u0_u7_ch_adr0[7] , _u0_u7_ch_adr0[6] ,_u0_u7_ch_adr0[5] , _u0_u7_ch_adr0[4] , _u0_u7_ch_adr0[3] ,_u0_u7_ch_adr0[2] , _u0_u7_ch_adr0[1] , _u0_u7_ch_adr0[0] ,_u0_u7_ch_adr1[31] , _u0_u7_ch_adr1[30] , _u0_u7_ch_adr1[29] ,_u0_u7_ch_adr1[28] , _u0_u7_ch_adr1[27] , _u0_u7_ch_adr1[26] ,_u0_u7_ch_adr1[25] , _u0_u7_ch_adr1[24] , _u0_u7_ch_adr1[23] ,_u0_u7_ch_adr1[22] , _u0_u7_ch_adr1[21] , _u0_u7_ch_adr1[20] ,_u0_u7_ch_adr1[19] , _u0_u7_ch_adr1[18] , _u0_u7_ch_adr1[17] ,_u0_u7_ch_adr1[16] , _u0_u7_ch_adr1[15] , _u0_u7_ch_adr1[14] ,_u0_u7_ch_adr1[13] , _u0_u7_ch_adr1[12] , _u0_u7_ch_adr1[11] ,_u0_u7_ch_adr1[10] , _u0_u7_ch_adr1[9] , _u0_u7_ch_adr1[8] ,_u0_u7_ch_adr1[7] , _u0_u7_ch_adr1[6] , _u0_u7_ch_adr1[5] ,_u0_u7_ch_adr1[4] , _u0_u7_ch_adr1[3] , _u0_u7_ch_adr1[2] ,_u0_u7_ch_adr1[1] , _u0_u7_ch_adr1[0] , _u0_u7_ch_am0[31] ,_u0_u7_ch_am0[30] , _u0_u7_ch_am0[29] , _u0_u7_ch_am0[28] ,_u0_u7_ch_am0[27] , _u0_u7_ch_am0[26] , _u0_u7_ch_am0[25] ,_u0_u7_ch_am0[24] , _u0_u7_ch_am0[23] , _u0_u7_ch_am0[22] ,_u0_u7_ch_am0[21] , _u0_u7_ch_am0[20] , _u0_u7_ch_am0[19] ,_u0_u7_ch_am0[18] , _u0_u7_ch_am0[17] , _u0_u7_ch_am0[16] ,_u0_u7_ch_am0[15] , _u0_u7_ch_am0[14] , _u0_u7_ch_am0[13] ,_u0_u7_ch_am0[12] , _u0_u7_ch_am0[11] , _u0_u7_ch_am0[10] ,_u0_u7_ch_am0[9] , _u0_u7_ch_am0[8] , _u0_u7_ch_am0[7] ,_u0_u7_ch_am0[6] , _u0_u7_ch_am0[5] , _u0_u7_ch_am0[4] ,_u0_u7_ch_am0[3] , _u0_u7_ch_am0[2] , _u0_u7_ch_am0[1] ,_u0_u7_ch_am0[0] , _u0_u7_ch_am1[31] , _u0_u7_ch_am1[30] ,_u0_u7_ch_am1[29] , _u0_u7_ch_am1[28] , _u0_u7_ch_am1[27] ,_u0_u7_ch_am1[26] , _u0_u7_ch_am1[25] , _u0_u7_ch_am1[24] ,_u0_u7_ch_am1[23] , _u0_u7_ch_am1[22] , _u0_u7_ch_am1[21] ,_u0_u7_ch_am1[20] , _u0_u7_ch_am1[19] , _u0_u7_ch_am1[18] ,_u0_u7_ch_am1[17] , _u0_u7_ch_am1[16] , _u0_u7_ch_am1[15] ,_u0_u7_ch_am1[14] , _u0_u7_ch_am1[13] , _u0_u7_ch_am1[12] ,_u0_u7_ch_am1[11] , _u0_u7_ch_am1[10] , _u0_u7_ch_am1[9] ,_u0_u7_ch_am1[8] , _u0_u7_ch_am1[7] , _u0_u7_ch_am1[6] ,_u0_u7_ch_am1[5] , _u0_u7_ch_am1[4] , _u0_u7_ch_am1[3] ,_u0_u7_ch_am1[2] , _u0_u7_ch_am1[1] , _u0_u7_ch_am1[0] ,_u0_u7_sw_pointer[31] , _u0_u7_sw_pointer[30] ,_u0_u7_sw_pointer[29] , _u0_u7_sw_pointer[28] ,_u0_u7_sw_pointer[27] , _u0_u7_sw_pointer[26] ,_u0_u7_sw_pointer[25] , _u0_u7_sw_pointer[24] ,_u0_u7_sw_pointer[23] , _u0_u7_sw_pointer[22] ,_u0_u7_sw_pointer[21] , _u0_u7_sw_pointer[20] ,_u0_u7_sw_pointer[19] , _u0_u7_sw_pointer[18] ,_u0_u7_sw_pointer[17] , _u0_u7_sw_pointer[16] ,_u0_u7_sw_pointer[15] , _u0_u7_sw_pointer[14] ,_u0_u7_sw_pointer[13] , _u0_u7_sw_pointer[12] ,_u0_u7_sw_pointer[11] , _u0_u7_sw_pointer[10] , _u0_u7_sw_pointer[9] ,_u0_u7_sw_pointer[8] , _u0_u7_sw_pointer[7] , _u0_u7_sw_pointer[6] ,_u0_u7_sw_pointer[5] , _u0_u7_sw_pointer[4] , _u0_u7_sw_pointer[3] ,_u0_u7_sw_pointer[2] , _u0_u7_sw_pointer[1] , _u0_u7_sw_pointer[0] ,_u0_u7_ch_stop , _u0_u7_ch_dis , _u0_u7_int , _u0_u8_pointer[31] ,_u0_u8_pointer[30] , _u0_u8_pointer[29] , _u0_u8_pointer[28] ,_u0_u8_pointer[27] , _u0_u8_pointer[26] , _u0_u8_pointer[25] ,_u0_u8_pointer[24] , _u0_u8_pointer[23] , _u0_u8_pointer[22] ,_u0_u8_pointer[21] , _u0_u8_pointer[20] , _u0_u8_pointer[19] ,_u0_u8_pointer[18] , _u0_u8_pointer[17] , _u0_u8_pointer[16] ,_u0_u8_pointer[15] , _u0_u8_pointer[14] , _u0_u8_pointer[13] ,_u0_u8_pointer[12] , _u0_u8_pointer[11] , _u0_u8_pointer[10] ,_u0_u8_pointer[9] , _u0_u8_pointer[8] , _u0_u8_pointer[7] ,_u0_u8_pointer[6] , _u0_u8_pointer[5] , _u0_u8_pointer[4] ,_u0_u8_pointer[3] , _u0_u8_pointer[2] , _u0_u8_pointer[1] ,_u0_u8_pointer[0] , _u0_u8_pointer_s[31] , _u0_u8_pointer_s[30] ,_u0_u8_pointer_s[29] , _u0_u8_pointer_s[28] , _u0_u8_pointer_s[27] ,_u0_u8_pointer_s[26] , _u0_u8_pointer_s[25] , _u0_u8_pointer_s[24] ,_u0_u8_pointer_s[23] , _u0_u8_pointer_s[22] , _u0_u8_pointer_s[21] ,_u0_u8_pointer_s[20] , _u0_u8_pointer_s[19] , _u0_u8_pointer_s[18] ,_u0_u8_pointer_s[17] , _u0_u8_pointer_s[16] , _u0_u8_pointer_s[15] ,_u0_u8_pointer_s[14] , _u0_u8_pointer_s[13] , _u0_u8_pointer_s[12] ,_u0_u8_pointer_s[11] , _u0_u8_pointer_s[10] , _u0_u8_pointer_s[9] ,_u0_u8_pointer_s[8] , _u0_u8_pointer_s[7] , _u0_u8_pointer_s[6] ,_u0_u8_pointer_s[5] , _u0_u8_pointer_s[4] , _u0_u8_pointer_s[3] ,_u0_u8_pointer_s[2] , _u0_u8_pointer_s[1] , _u0_u8_pointer_s[0] ,_u0_u8_ch_csr[31] , _u0_u8_ch_csr[30] , _u0_u8_ch_csr[29] ,_u0_u8_ch_csr[28] , _u0_u8_ch_csr[27] , _u0_u8_ch_csr[26] ,_u0_u8_ch_csr[25] , _u0_u8_ch_csr[24] , _u0_u8_ch_csr[23] ,_u0_u8_ch_csr[22] , _u0_u8_ch_csr[21] , _u0_u8_ch_csr[20] ,_u0_u8_ch_csr[19] , _u0_u8_ch_csr[18] , _u0_u8_ch_csr[17] ,_u0_u8_ch_csr[16] , _u0_u8_ch_csr[15] , _u0_u8_ch_csr[14] ,_u0_u8_ch_csr[13] , _u0_u8_ch_csr[12] , _u0_u8_ch_csr[11] ,_u0_u8_ch_csr[10] , _u0_u8_ch_csr[9] , _u0_u8_ch_csr[8] ,_u0_u8_ch_csr[7] , _u0_u8_ch_csr[6] , _u0_u8_ch_csr[5] ,_u0_u8_ch_csr[4] , _u0_u8_ch_csr[3] , _u0_u8_ch_csr[2] ,_u0_u8_ch_csr[1] , _u0_u8_ch_csr[0] , _u0_u8_ch_txsz[31] ,_u0_u8_ch_txsz[30] , _u0_u8_ch_txsz[29] , _u0_u8_ch_txsz[28] ,_u0_u8_ch_txsz[27] , _u0_u8_ch_txsz[26] , _u0_u8_ch_txsz[25] ,_u0_u8_ch_txsz[24] , _u0_u8_ch_txsz[23] , _u0_u8_ch_txsz[22] ,_u0_u8_ch_txsz[21] , _u0_u8_ch_txsz[20] , _u0_u8_ch_txsz[19] ,_u0_u8_ch_txsz[18] , _u0_u8_ch_txsz[17] , _u0_u8_ch_txsz[16] ,_u0_u8_ch_txsz[15] , _u0_u8_ch_txsz[14] , _u0_u8_ch_txsz[13] ,_u0_u8_ch_txsz[12] , _u0_u8_ch_txsz[11] , _u0_u8_ch_txsz[10] ,_u0_u8_ch_txsz[9] , _u0_u8_ch_txsz[8] , _u0_u8_ch_txsz[7] ,_u0_u8_ch_txsz[6] , _u0_u8_ch_txsz[5] , _u0_u8_ch_txsz[4] ,_u0_u8_ch_txsz[3] , _u0_u8_ch_txsz[2] , _u0_u8_ch_txsz[1] ,_u0_u8_ch_txsz[0] , _u0_u8_ch_adr0[31] , _u0_u8_ch_adr0[30] ,_u0_u8_ch_adr0[29] , _u0_u8_ch_adr0[28] , _u0_u8_ch_adr0[27] ,_u0_u8_ch_adr0[26] , _u0_u8_ch_adr0[25] , _u0_u8_ch_adr0[24] ,_u0_u8_ch_adr0[23] , _u0_u8_ch_adr0[22] , _u0_u8_ch_adr0[21] ,_u0_u8_ch_adr0[20] , _u0_u8_ch_adr0[19] , _u0_u8_ch_adr0[18] ,_u0_u8_ch_adr0[17] , _u0_u8_ch_adr0[16] , _u0_u8_ch_adr0[15] ,_u0_u8_ch_adr0[14] , _u0_u8_ch_adr0[13] , _u0_u8_ch_adr0[12] ,_u0_u8_ch_adr0[11] , _u0_u8_ch_adr0[10] , _u0_u8_ch_adr0[9] ,_u0_u8_ch_adr0[8] , _u0_u8_ch_adr0[7] , _u0_u8_ch_adr0[6] ,_u0_u8_ch_adr0[5] , _u0_u8_ch_adr0[4] , _u0_u8_ch_adr0[3] ,_u0_u8_ch_adr0[2] , _u0_u8_ch_adr0[1] , _u0_u8_ch_adr0[0] ,_u0_u8_ch_adr1[31] , _u0_u8_ch_adr1[30] , _u0_u8_ch_adr1[29] ,_u0_u8_ch_adr1[28] , _u0_u8_ch_adr1[27] , _u0_u8_ch_adr1[26] ,_u0_u8_ch_adr1[25] , _u0_u8_ch_adr1[24] , _u0_u8_ch_adr1[23] ,_u0_u8_ch_adr1[22] , _u0_u8_ch_adr1[21] , _u0_u8_ch_adr1[20] ,_u0_u8_ch_adr1[19] , _u0_u8_ch_adr1[18] , _u0_u8_ch_adr1[17] ,_u0_u8_ch_adr1[16] , _u0_u8_ch_adr1[15] , _u0_u8_ch_adr1[14] ,_u0_u8_ch_adr1[13] , _u0_u8_ch_adr1[12] , _u0_u8_ch_adr1[11] ,_u0_u8_ch_adr1[10] , _u0_u8_ch_adr1[9] , _u0_u8_ch_adr1[8] ,_u0_u8_ch_adr1[7] , _u0_u8_ch_adr1[6] , _u0_u8_ch_adr1[5] ,_u0_u8_ch_adr1[4] , _u0_u8_ch_adr1[3] , _u0_u8_ch_adr1[2] ,_u0_u8_ch_adr1[1] , _u0_u8_ch_adr1[0] , _u0_u8_ch_am0[31] ,_u0_u8_ch_am0[30] , _u0_u8_ch_am0[29] , _u0_u8_ch_am0[28] ,_u0_u8_ch_am0[27] , _u0_u8_ch_am0[26] , _u0_u8_ch_am0[25] ,_u0_u8_ch_am0[24] , _u0_u8_ch_am0[23] , _u0_u8_ch_am0[22] ,_u0_u8_ch_am0[21] , _u0_u8_ch_am0[20] , _u0_u8_ch_am0[19] ,_u0_u8_ch_am0[18] , _u0_u8_ch_am0[17] , _u0_u8_ch_am0[16] ,_u0_u8_ch_am0[15] , _u0_u8_ch_am0[14] , _u0_u8_ch_am0[13] ,_u0_u8_ch_am0[12] , _u0_u8_ch_am0[11] , _u0_u8_ch_am0[10] ,_u0_u8_ch_am0[9] , _u0_u8_ch_am0[8] , _u0_u8_ch_am0[7] ,_u0_u8_ch_am0[6] , _u0_u8_ch_am0[5] , _u0_u8_ch_am0[4] ,_u0_u8_ch_am0[3] , _u0_u8_ch_am0[2] , _u0_u8_ch_am0[1] ,_u0_u8_ch_am0[0] , _u0_u8_ch_am1[31] , _u0_u8_ch_am1[30] ,_u0_u8_ch_am1[29] , _u0_u8_ch_am1[28] , _u0_u8_ch_am1[27] ,_u0_u8_ch_am1[26] , _u0_u8_ch_am1[25] , _u0_u8_ch_am1[24] ,_u0_u8_ch_am1[23] , _u0_u8_ch_am1[22] , _u0_u8_ch_am1[21] ,_u0_u8_ch_am1[20] , _u0_u8_ch_am1[19] , _u0_u8_ch_am1[18] ,_u0_u8_ch_am1[17] , _u0_u8_ch_am1[16] , _u0_u8_ch_am1[15] ,_u0_u8_ch_am1[14] , _u0_u8_ch_am1[13] , _u0_u8_ch_am1[12] ,_u0_u8_ch_am1[11] , _u0_u8_ch_am1[10] , _u0_u8_ch_am1[9] ,_u0_u8_ch_am1[8] , _u0_u8_ch_am1[7] , _u0_u8_ch_am1[6] ,_u0_u8_ch_am1[5] , _u0_u8_ch_am1[4] , _u0_u8_ch_am1[3] ,_u0_u8_ch_am1[2] , _u0_u8_ch_am1[1] , _u0_u8_ch_am1[0] ,_u0_u8_sw_pointer[31] , _u0_u8_sw_pointer[30] ,_u0_u8_sw_pointer[29] , _u0_u8_sw_pointer[28] ,_u0_u8_sw_pointer[27] , _u0_u8_sw_pointer[26] ,_u0_u8_sw_pointer[25] , _u0_u8_sw_pointer[24] ,_u0_u8_sw_pointer[23] , _u0_u8_sw_pointer[22] ,_u0_u8_sw_pointer[21] , _u0_u8_sw_pointer[20] ,_u0_u8_sw_pointer[19] , _u0_u8_sw_pointer[18] ,_u0_u8_sw_pointer[17] , _u0_u8_sw_pointer[16] ,_u0_u8_sw_pointer[15] , _u0_u8_sw_pointer[14] ,_u0_u8_sw_pointer[13] , _u0_u8_sw_pointer[12] ,_u0_u8_sw_pointer[11] , _u0_u8_sw_pointer[10] , _u0_u8_sw_pointer[9] ,_u0_u8_sw_pointer[8] , _u0_u8_sw_pointer[7] , _u0_u8_sw_pointer[6] ,_u0_u8_sw_pointer[5] , _u0_u8_sw_pointer[4] , _u0_u8_sw_pointer[3] ,_u0_u8_sw_pointer[2] , _u0_u8_sw_pointer[1] , _u0_u8_sw_pointer[0] ,_u0_u8_ch_stop , _u0_u8_ch_dis , _u0_u8_int , _u0_u9_pointer[31] ,_u0_u9_pointer[30] , _u0_u9_pointer[29] , _u0_u9_pointer[28] ,_u0_u9_pointer[27] , _u0_u9_pointer[26] , _u0_u9_pointer[25] ,_u0_u9_pointer[24] , _u0_u9_pointer[23] , _u0_u9_pointer[22] ,_u0_u9_pointer[21] , _u0_u9_pointer[20] , _u0_u9_pointer[19] ,_u0_u9_pointer[18] , _u0_u9_pointer[17] , _u0_u9_pointer[16] ,_u0_u9_pointer[15] , _u0_u9_pointer[14] , _u0_u9_pointer[13] ,_u0_u9_pointer[12] , _u0_u9_pointer[11] , _u0_u9_pointer[10] ,_u0_u9_pointer[9] , _u0_u9_pointer[8] , _u0_u9_pointer[7] ,_u0_u9_pointer[6] , _u0_u9_pointer[5] , _u0_u9_pointer[4] ,_u0_u9_pointer[3] , _u0_u9_pointer[2] , _u0_u9_pointer[1] ,_u0_u9_pointer[0] , _u0_u9_pointer_s[31] , _u0_u9_pointer_s[30] ,_u0_u9_pointer_s[29] , _u0_u9_pointer_s[28] , _u0_u9_pointer_s[27] ,_u0_u9_pointer_s[26] , _u0_u9_pointer_s[25] , _u0_u9_pointer_s[24] ,_u0_u9_pointer_s[23] , _u0_u9_pointer_s[22] , _u0_u9_pointer_s[21] ,_u0_u9_pointer_s[20] , _u0_u9_pointer_s[19] , _u0_u9_pointer_s[18] ,_u0_u9_pointer_s[17] , _u0_u9_pointer_s[16] , _u0_u9_pointer_s[15] ,_u0_u9_pointer_s[14] , _u0_u9_pointer_s[13] , _u0_u9_pointer_s[12] ,_u0_u9_pointer_s[11] , _u0_u9_pointer_s[10] , _u0_u9_pointer_s[9] ,_u0_u9_pointer_s[8] , _u0_u9_pointer_s[7] , _u0_u9_pointer_s[6] ,_u0_u9_pointer_s[5] , _u0_u9_pointer_s[4] , _u0_u9_pointer_s[3] ,_u0_u9_pointer_s[2] , _u0_u9_pointer_s[1] , _u0_u9_pointer_s[0] ,_u0_u9_ch_csr[31] , _u0_u9_ch_csr[30] , _u0_u9_ch_csr[29] ,_u0_u9_ch_csr[28] , _u0_u9_ch_csr[27] , _u0_u9_ch_csr[26] ,_u0_u9_ch_csr[25] , _u0_u9_ch_csr[24] , _u0_u9_ch_csr[23] ,_u0_u9_ch_csr[22] , _u0_u9_ch_csr[21] , _u0_u9_ch_csr[20] ,_u0_u9_ch_csr[19] , _u0_u9_ch_csr[18] , _u0_u9_ch_csr[17] ,_u0_u9_ch_csr[16] , _u0_u9_ch_csr[15] , _u0_u9_ch_csr[14] ,_u0_u9_ch_csr[13] , _u0_u9_ch_csr[12] , _u0_u9_ch_csr[11] ,_u0_u9_ch_csr[10] , _u0_u9_ch_csr[9] , _u0_u9_ch_csr[8] ,_u0_u9_ch_csr[7] , _u0_u9_ch_csr[6] , _u0_u9_ch_csr[5] ,_u0_u9_ch_csr[4] , _u0_u9_ch_csr[3] , _u0_u9_ch_csr[2] ,_u0_u9_ch_csr[1] , _u0_u9_ch_csr[0] , _u0_u9_ch_txsz[31] ,_u0_u9_ch_txsz[30] , _u0_u9_ch_txsz[29] , _u0_u9_ch_txsz[28] ,_u0_u9_ch_txsz[27] , _u0_u9_ch_txsz[26] , _u0_u9_ch_txsz[25] ,_u0_u9_ch_txsz[24] , _u0_u9_ch_txsz[23] , _u0_u9_ch_txsz[22] ,_u0_u9_ch_txsz[21] , _u0_u9_ch_txsz[20] , _u0_u9_ch_txsz[19] ,_u0_u9_ch_txsz[18] , _u0_u9_ch_txsz[17] , _u0_u9_ch_txsz[16] ,_u0_u9_ch_txsz[15] , _u0_u9_ch_txsz[14] , _u0_u9_ch_txsz[13] ,_u0_u9_ch_txsz[12] , _u0_u9_ch_txsz[11] , _u0_u9_ch_txsz[10] ,_u0_u9_ch_txsz[9] , _u0_u9_ch_txsz[8] , _u0_u9_ch_txsz[7] ,_u0_u9_ch_txsz[6] , _u0_u9_ch_txsz[5] , _u0_u9_ch_txsz[4] ,_u0_u9_ch_txsz[3] , _u0_u9_ch_txsz[2] , _u0_u9_ch_txsz[1] ,_u0_u9_ch_txsz[0] , _u0_u9_ch_adr0[31] , _u0_u9_ch_adr0[30] ,_u0_u9_ch_adr0[29] , _u0_u9_ch_adr0[28] , _u0_u9_ch_adr0[27] ,_u0_u9_ch_adr0[26] , _u0_u9_ch_adr0[25] , _u0_u9_ch_adr0[24] ,_u0_u9_ch_adr0[23] , _u0_u9_ch_adr0[22] , _u0_u9_ch_adr0[21] ,_u0_u9_ch_adr0[20] , _u0_u9_ch_adr0[19] , _u0_u9_ch_adr0[18] ,_u0_u9_ch_adr0[17] , _u0_u9_ch_adr0[16] , _u0_u9_ch_adr0[15] ,_u0_u9_ch_adr0[14] , _u0_u9_ch_adr0[13] , _u0_u9_ch_adr0[12] ,_u0_u9_ch_adr0[11] , _u0_u9_ch_adr0[10] , _u0_u9_ch_adr0[9] ,_u0_u9_ch_adr0[8] , _u0_u9_ch_adr0[7] , _u0_u9_ch_adr0[6] ,_u0_u9_ch_adr0[5] , _u0_u9_ch_adr0[4] , _u0_u9_ch_adr0[3] ,_u0_u9_ch_adr0[2] , _u0_u9_ch_adr0[1] , _u0_u9_ch_adr0[0] ,_u0_u9_ch_adr1[31] , _u0_u9_ch_adr1[30] , _u0_u9_ch_adr1[29] ,_u0_u9_ch_adr1[28] , _u0_u9_ch_adr1[27] , _u0_u9_ch_adr1[26] ,_u0_u9_ch_adr1[25] , _u0_u9_ch_adr1[24] , _u0_u9_ch_adr1[23] ,_u0_u9_ch_adr1[22] , _u0_u9_ch_adr1[21] , _u0_u9_ch_adr1[20] ,_u0_u9_ch_adr1[19] , _u0_u9_ch_adr1[18] , _u0_u9_ch_adr1[17] ,_u0_u9_ch_adr1[16] , _u0_u9_ch_adr1[15] , _u0_u9_ch_adr1[14] ,_u0_u9_ch_adr1[13] , _u0_u9_ch_adr1[12] , _u0_u9_ch_adr1[11] ,_u0_u9_ch_adr1[10] , _u0_u9_ch_adr1[9] , _u0_u9_ch_adr1[8] ,_u0_u9_ch_adr1[7] , _u0_u9_ch_adr1[6] , _u0_u9_ch_adr1[5] ,_u0_u9_ch_adr1[4] , _u0_u9_ch_adr1[3] , _u0_u9_ch_adr1[2] ,_u0_u9_ch_adr1[1] , _u0_u9_ch_adr1[0] , _u0_u9_ch_am0[31] ,_u0_u9_ch_am0[30] , _u0_u9_ch_am0[29] , _u0_u9_ch_am0[28] ,_u0_u9_ch_am0[27] , _u0_u9_ch_am0[26] , _u0_u9_ch_am0[25] ,_u0_u9_ch_am0[24] , _u0_u9_ch_am0[23] , _u0_u9_ch_am0[22] ,_u0_u9_ch_am0[21] , _u0_u9_ch_am0[20] , _u0_u9_ch_am0[19] ,_u0_u9_ch_am0[18] , _u0_u9_ch_am0[17] , _u0_u9_ch_am0[16] ,_u0_u9_ch_am0[15] , _u0_u9_ch_am0[14] , _u0_u9_ch_am0[13] ,_u0_u9_ch_am0[12] , _u0_u9_ch_am0[11] , _u0_u9_ch_am0[10] ,_u0_u9_ch_am0[9] , _u0_u9_ch_am0[8] , _u0_u9_ch_am0[7] ,_u0_u9_ch_am0[6] , _u0_u9_ch_am0[5] , _u0_u9_ch_am0[4] ,_u0_u9_ch_am0[3] , _u0_u9_ch_am0[2] , _u0_u9_ch_am0[1] ,_u0_u9_ch_am0[0] , _u0_u9_ch_am1[31] , _u0_u9_ch_am1[30] ,_u0_u9_ch_am1[29] , _u0_u9_ch_am1[28] , _u0_u9_ch_am1[27] ,_u0_u9_ch_am1[26] , _u0_u9_ch_am1[25] , _u0_u9_ch_am1[24] ,_u0_u9_ch_am1[23] , _u0_u9_ch_am1[22] , _u0_u9_ch_am1[21] ,_u0_u9_ch_am1[20] , _u0_u9_ch_am1[19] , _u0_u9_ch_am1[18] ,_u0_u9_ch_am1[17] , _u0_u9_ch_am1[16] , _u0_u9_ch_am1[15] ,_u0_u9_ch_am1[14] , _u0_u9_ch_am1[13] , _u0_u9_ch_am1[12] ,_u0_u9_ch_am1[11] , _u0_u9_ch_am1[10] , _u0_u9_ch_am1[9] ,_u0_u9_ch_am1[8] , _u0_u9_ch_am1[7] , _u0_u9_ch_am1[6] ,_u0_u9_ch_am1[5] , _u0_u9_ch_am1[4] , _u0_u9_ch_am1[3] ,_u0_u9_ch_am1[2] , _u0_u9_ch_am1[1] , _u0_u9_ch_am1[0] ,_u0_u9_sw_pointer[31] , _u0_u9_sw_pointer[30] ,_u0_u9_sw_pointer[29] , _u0_u9_sw_pointer[28] ,_u0_u9_sw_pointer[27] , _u0_u9_sw_pointer[26] ,_u0_u9_sw_pointer[25] , _u0_u9_sw_pointer[24] ,_u0_u9_sw_pointer[23] , _u0_u9_sw_pointer[22] ,_u0_u9_sw_pointer[21] , _u0_u9_sw_pointer[20] ,_u0_u9_sw_pointer[19] , _u0_u9_sw_pointer[18] ,_u0_u9_sw_pointer[17] , _u0_u9_sw_pointer[16] ,_u0_u9_sw_pointer[15] , _u0_u9_sw_pointer[14] ,_u0_u9_sw_pointer[13] , _u0_u9_sw_pointer[12] ,_u0_u9_sw_pointer[11] , _u0_u9_sw_pointer[10] , _u0_u9_sw_pointer[9] ,_u0_u9_sw_pointer[8] , _u0_u9_sw_pointer[7] , _u0_u9_sw_pointer[6] ,_u0_u9_sw_pointer[5] , _u0_u9_sw_pointer[4] , _u0_u9_sw_pointer[3] ,_u0_u9_sw_pointer[2] , _u0_u9_sw_pointer[1] , _u0_u9_sw_pointer[0] ,_u0_u9_ch_stop , _u0_u9_ch_dis , _u0_u9_int , _u0_u10_pointer[31] ,_u0_u10_pointer[30] , _u0_u10_pointer[29] , _u0_u10_pointer[28] ,_u0_u10_pointer[27] , _u0_u10_pointer[26] , _u0_u10_pointer[25] ,_u0_u10_pointer[24] , _u0_u10_pointer[23] , _u0_u10_pointer[22] ,_u0_u10_pointer[21] , _u0_u10_pointer[20] , _u0_u10_pointer[19] ,_u0_u10_pointer[18] , _u0_u10_pointer[17] , _u0_u10_pointer[16] ,_u0_u10_pointer[15] , _u0_u10_pointer[14] , _u0_u10_pointer[13] ,_u0_u10_pointer[12] , _u0_u10_pointer[11] , _u0_u10_pointer[10] ,_u0_u10_pointer[9] , _u0_u10_pointer[8] , _u0_u10_pointer[7] ,_u0_u10_pointer[6] , _u0_u10_pointer[5] , _u0_u10_pointer[4] ,_u0_u10_pointer[3] , _u0_u10_pointer[2] , _u0_u10_pointer[1] ,_u0_u10_pointer[0] , _u0_u10_pointer_s[31] , _u0_u10_pointer_s[30] ,_u0_u10_pointer_s[29] , _u0_u10_pointer_s[28] ,_u0_u10_pointer_s[27] , _u0_u10_pointer_s[26] ,_u0_u10_pointer_s[25] , _u0_u10_pointer_s[24] ,_u0_u10_pointer_s[23] , _u0_u10_pointer_s[22] ,_u0_u10_pointer_s[21] , _u0_u10_pointer_s[20] ,_u0_u10_pointer_s[19] , _u0_u10_pointer_s[18] ,_u0_u10_pointer_s[17] , _u0_u10_pointer_s[16] ,_u0_u10_pointer_s[15] , _u0_u10_pointer_s[14] ,_u0_u10_pointer_s[13] , _u0_u10_pointer_s[12] ,_u0_u10_pointer_s[11] , _u0_u10_pointer_s[10] , _u0_u10_pointer_s[9] ,_u0_u10_pointer_s[8] , _u0_u10_pointer_s[7] , _u0_u10_pointer_s[6] ,_u0_u10_pointer_s[5] , _u0_u10_pointer_s[4] , _u0_u10_pointer_s[3] ,_u0_u10_pointer_s[2] , _u0_u10_pointer_s[1] , _u0_u10_pointer_s[0] ,_u0_u10_ch_csr[31] , _u0_u10_ch_csr[30] , _u0_u10_ch_csr[29] ,_u0_u10_ch_csr[28] , _u0_u10_ch_csr[27] , _u0_u10_ch_csr[26] ,_u0_u10_ch_csr[25] , _u0_u10_ch_csr[24] , _u0_u10_ch_csr[23] ,_u0_u10_ch_csr[22] , _u0_u10_ch_csr[21] , _u0_u10_ch_csr[20] ,_u0_u10_ch_csr[19] , _u0_u10_ch_csr[18] , _u0_u10_ch_csr[17] ,_u0_u10_ch_csr[16] , _u0_u10_ch_csr[15] , _u0_u10_ch_csr[14] ,_u0_u10_ch_csr[13] , _u0_u10_ch_csr[12] , _u0_u10_ch_csr[11] ,_u0_u10_ch_csr[10] , _u0_u10_ch_csr[9] , _u0_u10_ch_csr[8] ,_u0_u10_ch_csr[7] , _u0_u10_ch_csr[6] , _u0_u10_ch_csr[5] ,_u0_u10_ch_csr[4] , _u0_u10_ch_csr[3] , _u0_u10_ch_csr[2] ,_u0_u10_ch_csr[1] , _u0_u10_ch_csr[0] , _u0_u10_ch_txsz[31] ,_u0_u10_ch_txsz[30] , _u0_u10_ch_txsz[29] , _u0_u10_ch_txsz[28] ,_u0_u10_ch_txsz[27] , _u0_u10_ch_txsz[26] , _u0_u10_ch_txsz[25] ,_u0_u10_ch_txsz[24] , _u0_u10_ch_txsz[23] , _u0_u10_ch_txsz[22] ,_u0_u10_ch_txsz[21] , _u0_u10_ch_txsz[20] , _u0_u10_ch_txsz[19] ,_u0_u10_ch_txsz[18] , _u0_u10_ch_txsz[17] , _u0_u10_ch_txsz[16] ,_u0_u10_ch_txsz[15] , _u0_u10_ch_txsz[14] , _u0_u10_ch_txsz[13] ,_u0_u10_ch_txsz[12] , _u0_u10_ch_txsz[11] , _u0_u10_ch_txsz[10] ,_u0_u10_ch_txsz[9] , _u0_u10_ch_txsz[8] , _u0_u10_ch_txsz[7] ,_u0_u10_ch_txsz[6] , _u0_u10_ch_txsz[5] , _u0_u10_ch_txsz[4] ,_u0_u10_ch_txsz[3] , _u0_u10_ch_txsz[2] , _u0_u10_ch_txsz[1] ,_u0_u10_ch_txsz[0] , _u0_u10_ch_adr0[31] , _u0_u10_ch_adr0[30] ,_u0_u10_ch_adr0[29] , _u0_u10_ch_adr0[28] , _u0_u10_ch_adr0[27] ,_u0_u10_ch_adr0[26] , _u0_u10_ch_adr0[25] , _u0_u10_ch_adr0[24] ,_u0_u10_ch_adr0[23] , _u0_u10_ch_adr0[22] , _u0_u10_ch_adr0[21] ,_u0_u10_ch_adr0[20] , _u0_u10_ch_adr0[19] , _u0_u10_ch_adr0[18] ,_u0_u10_ch_adr0[17] , _u0_u10_ch_adr0[16] , _u0_u10_ch_adr0[15] ,_u0_u10_ch_adr0[14] , _u0_u10_ch_adr0[13] , _u0_u10_ch_adr0[12] ,_u0_u10_ch_adr0[11] , _u0_u10_ch_adr0[10] , _u0_u10_ch_adr0[9] ,_u0_u10_ch_adr0[8] , _u0_u10_ch_adr0[7] , _u0_u10_ch_adr0[6] ,_u0_u10_ch_adr0[5] , _u0_u10_ch_adr0[4] , _u0_u10_ch_adr0[3] ,_u0_u10_ch_adr0[2] , _u0_u10_ch_adr0[1] , _u0_u10_ch_adr0[0] ,_u0_u10_ch_adr1[31] , _u0_u10_ch_adr1[30] , _u0_u10_ch_adr1[29] ,_u0_u10_ch_adr1[28] , _u0_u10_ch_adr1[27] , _u0_u10_ch_adr1[26] ,_u0_u10_ch_adr1[25] , _u0_u10_ch_adr1[24] , _u0_u10_ch_adr1[23] ,_u0_u10_ch_adr1[22] , _u0_u10_ch_adr1[21] , _u0_u10_ch_adr1[20] ,_u0_u10_ch_adr1[19] , _u0_u10_ch_adr1[18] , _u0_u10_ch_adr1[17] ,_u0_u10_ch_adr1[16] , _u0_u10_ch_adr1[15] , _u0_u10_ch_adr1[14] ,_u0_u10_ch_adr1[13] , _u0_u10_ch_adr1[12] , _u0_u10_ch_adr1[11] ,_u0_u10_ch_adr1[10] , _u0_u10_ch_adr1[9] , _u0_u10_ch_adr1[8] ,_u0_u10_ch_adr1[7] , _u0_u10_ch_adr1[6] , _u0_u10_ch_adr1[5] ,_u0_u10_ch_adr1[4] , _u0_u10_ch_adr1[3] , _u0_u10_ch_adr1[2] ,_u0_u10_ch_adr1[1] , _u0_u10_ch_adr1[0] , _u0_u10_ch_am0[31] ,_u0_u10_ch_am0[30] , _u0_u10_ch_am0[29] , _u0_u10_ch_am0[28] ,_u0_u10_ch_am0[27] , _u0_u10_ch_am0[26] , _u0_u10_ch_am0[25] ,_u0_u10_ch_am0[24] , _u0_u10_ch_am0[23] , _u0_u10_ch_am0[22] ,_u0_u10_ch_am0[21] , _u0_u10_ch_am0[20] , _u0_u10_ch_am0[19] ,_u0_u10_ch_am0[18] , _u0_u10_ch_am0[17] , _u0_u10_ch_am0[16] ,_u0_u10_ch_am0[15] , _u0_u10_ch_am0[14] , _u0_u10_ch_am0[13] ,_u0_u10_ch_am0[12] , _u0_u10_ch_am0[11] , _u0_u10_ch_am0[10] ,_u0_u10_ch_am0[9] , _u0_u10_ch_am0[8] , _u0_u10_ch_am0[7] ,_u0_u10_ch_am0[6] , _u0_u10_ch_am0[5] , _u0_u10_ch_am0[4] ,_u0_u10_ch_am0[3] , _u0_u10_ch_am0[2] , _u0_u10_ch_am0[1] ,_u0_u10_ch_am0[0] , _u0_u10_ch_am1[31] , _u0_u10_ch_am1[30] ,_u0_u10_ch_am1[29] , _u0_u10_ch_am1[28] , _u0_u10_ch_am1[27] ,_u0_u10_ch_am1[26] , _u0_u10_ch_am1[25] , _u0_u10_ch_am1[24] ,_u0_u10_ch_am1[23] , _u0_u10_ch_am1[22] , _u0_u10_ch_am1[21] ,_u0_u10_ch_am1[20] , _u0_u10_ch_am1[19] , _u0_u10_ch_am1[18] ,_u0_u10_ch_am1[17] , _u0_u10_ch_am1[16] , _u0_u10_ch_am1[15] ,_u0_u10_ch_am1[14] , _u0_u10_ch_am1[13] , _u0_u10_ch_am1[12] ,_u0_u10_ch_am1[11] , _u0_u10_ch_am1[10] , _u0_u10_ch_am1[9] ,_u0_u10_ch_am1[8] , _u0_u10_ch_am1[7] , _u0_u10_ch_am1[6] ,_u0_u10_ch_am1[5] , _u0_u10_ch_am1[4] , _u0_u10_ch_am1[3] ,_u0_u10_ch_am1[2] , _u0_u10_ch_am1[1] , _u0_u10_ch_am1[0] ,_u0_u10_sw_pointer[31] , _u0_u10_sw_pointer[30] ,_u0_u10_sw_pointer[29] , _u0_u10_sw_pointer[28] ,_u0_u10_sw_pointer[27] , _u0_u10_sw_pointer[26] ,_u0_u10_sw_pointer[25] , _u0_u10_sw_pointer[24] ,_u0_u10_sw_pointer[23] , _u0_u10_sw_pointer[22] ,_u0_u10_sw_pointer[21] , _u0_u10_sw_pointer[20] ,_u0_u10_sw_pointer[19] , _u0_u10_sw_pointer[18] ,_u0_u10_sw_pointer[17] , _u0_u10_sw_pointer[16] ,_u0_u10_sw_pointer[15] , _u0_u10_sw_pointer[14] ,_u0_u10_sw_pointer[13] , _u0_u10_sw_pointer[12] ,_u0_u10_sw_pointer[11] , _u0_u10_sw_pointer[10] ,_u0_u10_sw_pointer[9] , _u0_u10_sw_pointer[8] ,_u0_u10_sw_pointer[7] , _u0_u10_sw_pointer[6] ,_u0_u10_sw_pointer[5] , _u0_u10_sw_pointer[4] ,_u0_u10_sw_pointer[3] , _u0_u10_sw_pointer[2] ,_u0_u10_sw_pointer[1] , _u0_u10_sw_pointer[0] , _u0_u10_ch_stop ,_u0_u10_ch_dis , _u0_u10_int , _u0_u11_pointer[31] ,_u0_u11_pointer[30] , _u0_u11_pointer[29] , _u0_u11_pointer[28] ,_u0_u11_pointer[27] , _u0_u11_pointer[26] , _u0_u11_pointer[25] ,_u0_u11_pointer[24] , _u0_u11_pointer[23] , _u0_u11_pointer[22] ,_u0_u11_pointer[21] , _u0_u11_pointer[20] , _u0_u11_pointer[19] ,_u0_u11_pointer[18] , _u0_u11_pointer[17] , _u0_u11_pointer[16] ,_u0_u11_pointer[15] , _u0_u11_pointer[14] , _u0_u11_pointer[13] ,_u0_u11_pointer[12] , _u0_u11_pointer[11] , _u0_u11_pointer[10] ,_u0_u11_pointer[9] , _u0_u11_pointer[8] , _u0_u11_pointer[7] ,_u0_u11_pointer[6] , _u0_u11_pointer[5] , _u0_u11_pointer[4] ,_u0_u11_pointer[3] , _u0_u11_pointer[2] , _u0_u11_pointer[1] ,_u0_u11_pointer[0] , _u0_u11_pointer_s[31] , _u0_u11_pointer_s[30] ,_u0_u11_pointer_s[29] , _u0_u11_pointer_s[28] ,_u0_u11_pointer_s[27] , _u0_u11_pointer_s[26] ,_u0_u11_pointer_s[25] , _u0_u11_pointer_s[24] ,_u0_u11_pointer_s[23] , _u0_u11_pointer_s[22] ,_u0_u11_pointer_s[21] , _u0_u11_pointer_s[20] ,_u0_u11_pointer_s[19] , _u0_u11_pointer_s[18] ,_u0_u11_pointer_s[17] , _u0_u11_pointer_s[16] ,_u0_u11_pointer_s[15] , _u0_u11_pointer_s[14] ,_u0_u11_pointer_s[13] , _u0_u11_pointer_s[12] ,_u0_u11_pointer_s[11] , _u0_u11_pointer_s[10] , _u0_u11_pointer_s[9] ,_u0_u11_pointer_s[8] , _u0_u11_pointer_s[7] , _u0_u11_pointer_s[6] ,_u0_u11_pointer_s[5] , _u0_u11_pointer_s[4] , _u0_u11_pointer_s[3] ,_u0_u11_pointer_s[2] , _u0_u11_pointer_s[1] , _u0_u11_pointer_s[0] ,_u0_u11_ch_csr[31] , _u0_u11_ch_csr[30] , _u0_u11_ch_csr[29] ,_u0_u11_ch_csr[28] , _u0_u11_ch_csr[27] , _u0_u11_ch_csr[26] ,_u0_u11_ch_csr[25] , _u0_u11_ch_csr[24] , _u0_u11_ch_csr[23] ,_u0_u11_ch_csr[22] , _u0_u11_ch_csr[21] , _u0_u11_ch_csr[20] ,_u0_u11_ch_csr[19] , _u0_u11_ch_csr[18] , _u0_u11_ch_csr[17] ,_u0_u11_ch_csr[16] , _u0_u11_ch_csr[15] , _u0_u11_ch_csr[14] ,_u0_u11_ch_csr[13] , _u0_u11_ch_csr[12] , _u0_u11_ch_csr[11] ,_u0_u11_ch_csr[10] , _u0_u11_ch_csr[9] , _u0_u11_ch_csr[8] ,_u0_u11_ch_csr[7] , _u0_u11_ch_csr[6] , _u0_u11_ch_csr[5] ,_u0_u11_ch_csr[4] , _u0_u11_ch_csr[3] , _u0_u11_ch_csr[2] ,_u0_u11_ch_csr[1] , _u0_u11_ch_csr[0] , _u0_u11_ch_txsz[31] ,_u0_u11_ch_txsz[30] , _u0_u11_ch_txsz[29] , _u0_u11_ch_txsz[28] ,_u0_u11_ch_txsz[27] , _u0_u11_ch_txsz[26] , _u0_u11_ch_txsz[25] ,_u0_u11_ch_txsz[24] , _u0_u11_ch_txsz[23] , _u0_u11_ch_txsz[22] ,_u0_u11_ch_txsz[21] , _u0_u11_ch_txsz[20] , _u0_u11_ch_txsz[19] ,_u0_u11_ch_txsz[18] , _u0_u11_ch_txsz[17] , _u0_u11_ch_txsz[16] ,_u0_u11_ch_txsz[15] , _u0_u11_ch_txsz[14] , _u0_u11_ch_txsz[13] ,_u0_u11_ch_txsz[12] , _u0_u11_ch_txsz[11] , _u0_u11_ch_txsz[10] ,_u0_u11_ch_txsz[9] , _u0_u11_ch_txsz[8] , _u0_u11_ch_txsz[7] ,_u0_u11_ch_txsz[6] , _u0_u11_ch_txsz[5] , _u0_u11_ch_txsz[4] ,_u0_u11_ch_txsz[3] , _u0_u11_ch_txsz[2] , _u0_u11_ch_txsz[1] ,_u0_u11_ch_txsz[0] , _u0_u11_ch_adr0[31] , _u0_u11_ch_adr0[30] ,_u0_u11_ch_adr0[29] , _u0_u11_ch_adr0[28] , _u0_u11_ch_adr0[27] ,_u0_u11_ch_adr0[26] , _u0_u11_ch_adr0[25] , _u0_u11_ch_adr0[24] ,_u0_u11_ch_adr0[23] , _u0_u11_ch_adr0[22] , _u0_u11_ch_adr0[21] ,_u0_u11_ch_adr0[20] , _u0_u11_ch_adr0[19] , _u0_u11_ch_adr0[18] ,_u0_u11_ch_adr0[17] , _u0_u11_ch_adr0[16] , _u0_u11_ch_adr0[15] ,_u0_u11_ch_adr0[14] , _u0_u11_ch_adr0[13] , _u0_u11_ch_adr0[12] ,_u0_u11_ch_adr0[11] , _u0_u11_ch_adr0[10] , _u0_u11_ch_adr0[9] ,_u0_u11_ch_adr0[8] , _u0_u11_ch_adr0[7] , _u0_u11_ch_adr0[6] ,_u0_u11_ch_adr0[5] , _u0_u11_ch_adr0[4] , _u0_u11_ch_adr0[3] ,_u0_u11_ch_adr0[2] , _u0_u11_ch_adr0[1] , _u0_u11_ch_adr0[0] ,_u0_u11_ch_adr1[31] , _u0_u11_ch_adr1[30] , _u0_u11_ch_adr1[29] ,_u0_u11_ch_adr1[28] , _u0_u11_ch_adr1[27] , _u0_u11_ch_adr1[26] ,_u0_u11_ch_adr1[25] , _u0_u11_ch_adr1[24] , _u0_u11_ch_adr1[23] ,_u0_u11_ch_adr1[22] , _u0_u11_ch_adr1[21] , _u0_u11_ch_adr1[20] ,_u0_u11_ch_adr1[19] , _u0_u11_ch_adr1[18] , _u0_u11_ch_adr1[17] ,_u0_u11_ch_adr1[16] , _u0_u11_ch_adr1[15] , _u0_u11_ch_adr1[14] ,_u0_u11_ch_adr1[13] , _u0_u11_ch_adr1[12] , _u0_u11_ch_adr1[11] ,_u0_u11_ch_adr1[10] , _u0_u11_ch_adr1[9] , _u0_u11_ch_adr1[8] ,_u0_u11_ch_adr1[7] , _u0_u11_ch_adr1[6] , _u0_u11_ch_adr1[5] ,_u0_u11_ch_adr1[4] , _u0_u11_ch_adr1[3] , _u0_u11_ch_adr1[2] ,_u0_u11_ch_adr1[1] , _u0_u11_ch_adr1[0] , _u0_u11_ch_am0[31] ,_u0_u11_ch_am0[30] , _u0_u11_ch_am0[29] , _u0_u11_ch_am0[28] ,_u0_u11_ch_am0[27] , _u0_u11_ch_am0[26] , _u0_u11_ch_am0[25] ,_u0_u11_ch_am0[24] , _u0_u11_ch_am0[23] , _u0_u11_ch_am0[22] ,_u0_u11_ch_am0[21] , _u0_u11_ch_am0[20] , _u0_u11_ch_am0[19] ,_u0_u11_ch_am0[18] , _u0_u11_ch_am0[17] , _u0_u11_ch_am0[16] ,_u0_u11_ch_am0[15] , _u0_u11_ch_am0[14] , _u0_u11_ch_am0[13] ,_u0_u11_ch_am0[12] , _u0_u11_ch_am0[11] , _u0_u11_ch_am0[10] ,_u0_u11_ch_am0[9] , _u0_u11_ch_am0[8] , _u0_u11_ch_am0[7] ,_u0_u11_ch_am0[6] , _u0_u11_ch_am0[5] , _u0_u11_ch_am0[4] ,_u0_u11_ch_am0[3] , _u0_u11_ch_am0[2] , _u0_u11_ch_am0[1] ,_u0_u11_ch_am0[0] , _u0_u11_ch_am1[31] , _u0_u11_ch_am1[30] ,_u0_u11_ch_am1[29] , _u0_u11_ch_am1[28] , _u0_u11_ch_am1[27] ,_u0_u11_ch_am1[26] , _u0_u11_ch_am1[25] , _u0_u11_ch_am1[24] ,_u0_u11_ch_am1[23] , _u0_u11_ch_am1[22] , _u0_u11_ch_am1[21] ,_u0_u11_ch_am1[20] , _u0_u11_ch_am1[19] , _u0_u11_ch_am1[18] ,_u0_u11_ch_am1[17] , _u0_u11_ch_am1[16] , _u0_u11_ch_am1[15] ,_u0_u11_ch_am1[14] , _u0_u11_ch_am1[13] , _u0_u11_ch_am1[12] ,_u0_u11_ch_am1[11] , _u0_u11_ch_am1[10] , _u0_u11_ch_am1[9] ,_u0_u11_ch_am1[8] , _u0_u11_ch_am1[7] , _u0_u11_ch_am1[6] ,_u0_u11_ch_am1[5] , _u0_u11_ch_am1[4] , _u0_u11_ch_am1[3] ,_u0_u11_ch_am1[2] , _u0_u11_ch_am1[1] , _u0_u11_ch_am1[0] ,_u0_u11_sw_pointer[31] , _u0_u11_sw_pointer[30] ,_u0_u11_sw_pointer[29] , _u0_u11_sw_pointer[28] ,_u0_u11_sw_pointer[27] , _u0_u11_sw_pointer[26] ,_u0_u11_sw_pointer[25] , _u0_u11_sw_pointer[24] ,_u0_u11_sw_pointer[23] , _u0_u11_sw_pointer[22] ,_u0_u11_sw_pointer[21] , _u0_u11_sw_pointer[20] ,_u0_u11_sw_pointer[19] , _u0_u11_sw_pointer[18] ,_u0_u11_sw_pointer[17] , _u0_u11_sw_pointer[16] ,_u0_u11_sw_pointer[15] , _u0_u11_sw_pointer[14] ,_u0_u11_sw_pointer[13] , _u0_u11_sw_pointer[12] ,_u0_u11_sw_pointer[11] , _u0_u11_sw_pointer[10] ,_u0_u11_sw_pointer[9] , _u0_u11_sw_pointer[8] ,_u0_u11_sw_pointer[7] , _u0_u11_sw_pointer[6] ,_u0_u11_sw_pointer[5] , _u0_u11_sw_pointer[4] ,_u0_u11_sw_pointer[3] , _u0_u11_sw_pointer[2] ,_u0_u11_sw_pointer[1] , _u0_u11_sw_pointer[0] , _u0_u11_ch_stop ,_u0_u11_ch_dis , _u0_u11_int , _u0_u12_pointer[31] ,_u0_u12_pointer[30] , _u0_u12_pointer[29] , _u0_u12_pointer[28] ,_u0_u12_pointer[27] , _u0_u12_pointer[26] , _u0_u12_pointer[25] ,_u0_u12_pointer[24] , _u0_u12_pointer[23] , _u0_u12_pointer[22] ,_u0_u12_pointer[21] , _u0_u12_pointer[20] , _u0_u12_pointer[19] ,_u0_u12_pointer[18] , _u0_u12_pointer[17] , _u0_u12_pointer[16] ,_u0_u12_pointer[15] , _u0_u12_pointer[14] , _u0_u12_pointer[13] ,_u0_u12_pointer[12] , _u0_u12_pointer[11] , _u0_u12_pointer[10] ,_u0_u12_pointer[9] , _u0_u12_pointer[8] , _u0_u12_pointer[7] ,_u0_u12_pointer[6] , _u0_u12_pointer[5] , _u0_u12_pointer[4] ,_u0_u12_pointer[3] , _u0_u12_pointer[2] , _u0_u12_pointer[1] ,_u0_u12_pointer[0] , _u0_u12_pointer_s[31] , _u0_u12_pointer_s[30] ,_u0_u12_pointer_s[29] , _u0_u12_pointer_s[28] ,_u0_u12_pointer_s[27] , _u0_u12_pointer_s[26] ,_u0_u12_pointer_s[25] , _u0_u12_pointer_s[24] ,_u0_u12_pointer_s[23] , _u0_u12_pointer_s[22] ,_u0_u12_pointer_s[21] , _u0_u12_pointer_s[20] ,_u0_u12_pointer_s[19] , _u0_u12_pointer_s[18] ,_u0_u12_pointer_s[17] , _u0_u12_pointer_s[16] ,_u0_u12_pointer_s[15] , _u0_u12_pointer_s[14] ,_u0_u12_pointer_s[13] , _u0_u12_pointer_s[12] ,_u0_u12_pointer_s[11] , _u0_u12_pointer_s[10] , _u0_u12_pointer_s[9] ,_u0_u12_pointer_s[8] , _u0_u12_pointer_s[7] , _u0_u12_pointer_s[6] ,_u0_u12_pointer_s[5] , _u0_u12_pointer_s[4] , _u0_u12_pointer_s[3] ,_u0_u12_pointer_s[2] , _u0_u12_pointer_s[1] , _u0_u12_pointer_s[0] ,_u0_u12_ch_csr[31] , _u0_u12_ch_csr[30] , _u0_u12_ch_csr[29] ,_u0_u12_ch_csr[28] , _u0_u12_ch_csr[27] , _u0_u12_ch_csr[26] ,_u0_u12_ch_csr[25] , _u0_u12_ch_csr[24] , _u0_u12_ch_csr[23] ,_u0_u12_ch_csr[22] , _u0_u12_ch_csr[21] , _u0_u12_ch_csr[20] ,_u0_u12_ch_csr[19] , _u0_u12_ch_csr[18] , _u0_u12_ch_csr[17] ,_u0_u12_ch_csr[16] , _u0_u12_ch_csr[15] , _u0_u12_ch_csr[14] ,_u0_u12_ch_csr[13] , _u0_u12_ch_csr[12] , _u0_u12_ch_csr[11] ,_u0_u12_ch_csr[10] , _u0_u12_ch_csr[9] , _u0_u12_ch_csr[8] ,_u0_u12_ch_csr[7] , _u0_u12_ch_csr[6] , _u0_u12_ch_csr[5] ,_u0_u12_ch_csr[4] , _u0_u12_ch_csr[3] , _u0_u12_ch_csr[2] ,_u0_u12_ch_csr[1] , _u0_u12_ch_csr[0] , _u0_u12_ch_txsz[31] ,_u0_u12_ch_txsz[30] , _u0_u12_ch_txsz[29] , _u0_u12_ch_txsz[28] ,_u0_u12_ch_txsz[27] , _u0_u12_ch_txsz[26] , _u0_u12_ch_txsz[25] ,_u0_u12_ch_txsz[24] , _u0_u12_ch_txsz[23] , _u0_u12_ch_txsz[22] ,_u0_u12_ch_txsz[21] , _u0_u12_ch_txsz[20] , _u0_u12_ch_txsz[19] ,_u0_u12_ch_txsz[18] , _u0_u12_ch_txsz[17] , _u0_u12_ch_txsz[16] ,_u0_u12_ch_txsz[15] , _u0_u12_ch_txsz[14] , _u0_u12_ch_txsz[13] ,_u0_u12_ch_txsz[12] , _u0_u12_ch_txsz[11] , _u0_u12_ch_txsz[10] ,_u0_u12_ch_txsz[9] , _u0_u12_ch_txsz[8] , _u0_u12_ch_txsz[7] ,_u0_u12_ch_txsz[6] , _u0_u12_ch_txsz[5] , _u0_u12_ch_txsz[4] ,_u0_u12_ch_txsz[3] , _u0_u12_ch_txsz[2] , _u0_u12_ch_txsz[1] ,_u0_u12_ch_txsz[0] , _u0_u12_ch_adr0[31] , _u0_u12_ch_adr0[30] ,_u0_u12_ch_adr0[29] , _u0_u12_ch_adr0[28] , _u0_u12_ch_adr0[27] ,_u0_u12_ch_adr0[26] , _u0_u12_ch_adr0[25] , _u0_u12_ch_adr0[24] ,_u0_u12_ch_adr0[23] , _u0_u12_ch_adr0[22] , _u0_u12_ch_adr0[21] ,_u0_u12_ch_adr0[20] , _u0_u12_ch_adr0[19] , _u0_u12_ch_adr0[18] ,_u0_u12_ch_adr0[17] , _u0_u12_ch_adr0[16] , _u0_u12_ch_adr0[15] ,_u0_u12_ch_adr0[14] , _u0_u12_ch_adr0[13] , _u0_u12_ch_adr0[12] ,_u0_u12_ch_adr0[11] , _u0_u12_ch_adr0[10] , _u0_u12_ch_adr0[9] ,_u0_u12_ch_adr0[8] , _u0_u12_ch_adr0[7] , _u0_u12_ch_adr0[6] ,_u0_u12_ch_adr0[5] , _u0_u12_ch_adr0[4] , _u0_u12_ch_adr0[3] ,_u0_u12_ch_adr0[2] , _u0_u12_ch_adr0[1] , _u0_u12_ch_adr0[0] ,_u0_u12_ch_adr1[31] , _u0_u12_ch_adr1[30] , _u0_u12_ch_adr1[29] ,_u0_u12_ch_adr1[28] , _u0_u12_ch_adr1[27] , _u0_u12_ch_adr1[26] ,_u0_u12_ch_adr1[25] , _u0_u12_ch_adr1[24] , _u0_u12_ch_adr1[23] ,_u0_u12_ch_adr1[22] , _u0_u12_ch_adr1[21] , _u0_u12_ch_adr1[20] ,_u0_u12_ch_adr1[19] , _u0_u12_ch_adr1[18] , _u0_u12_ch_adr1[17] ,_u0_u12_ch_adr1[16] , _u0_u12_ch_adr1[15] , _u0_u12_ch_adr1[14] ,_u0_u12_ch_adr1[13] , _u0_u12_ch_adr1[12] , _u0_u12_ch_adr1[11] ,_u0_u12_ch_adr1[10] , _u0_u12_ch_adr1[9] , _u0_u12_ch_adr1[8] ,_u0_u12_ch_adr1[7] , _u0_u12_ch_adr1[6] , _u0_u12_ch_adr1[5] ,_u0_u12_ch_adr1[4] , _u0_u12_ch_adr1[3] , _u0_u12_ch_adr1[2] ,_u0_u12_ch_adr1[1] , _u0_u12_ch_adr1[0] , _u0_u12_ch_am0[31] ,_u0_u12_ch_am0[30] , _u0_u12_ch_am0[29] , _u0_u12_ch_am0[28] ,_u0_u12_ch_am0[27] , _u0_u12_ch_am0[26] , _u0_u12_ch_am0[25] ,_u0_u12_ch_am0[24] , _u0_u12_ch_am0[23] , _u0_u12_ch_am0[22] ,_u0_u12_ch_am0[21] , _u0_u12_ch_am0[20] , _u0_u12_ch_am0[19] ,_u0_u12_ch_am0[18] , _u0_u12_ch_am0[17] , _u0_u12_ch_am0[16] ,_u0_u12_ch_am0[15] , _u0_u12_ch_am0[14] , _u0_u12_ch_am0[13] ,_u0_u12_ch_am0[12] , _u0_u12_ch_am0[11] , _u0_u12_ch_am0[10] ,_u0_u12_ch_am0[9] , _u0_u12_ch_am0[8] , _u0_u12_ch_am0[7] ,_u0_u12_ch_am0[6] , _u0_u12_ch_am0[5] , _u0_u12_ch_am0[4] ,_u0_u12_ch_am0[3] , _u0_u12_ch_am0[2] , _u0_u12_ch_am0[1] ,_u0_u12_ch_am0[0] , _u0_u12_ch_am1[31] , _u0_u12_ch_am1[30] ,_u0_u12_ch_am1[29] , _u0_u12_ch_am1[28] , _u0_u12_ch_am1[27] ,_u0_u12_ch_am1[26] , _u0_u12_ch_am1[25] , _u0_u12_ch_am1[24] ,_u0_u12_ch_am1[23] , _u0_u12_ch_am1[22] , _u0_u12_ch_am1[21] ,_u0_u12_ch_am1[20] , _u0_u12_ch_am1[19] , _u0_u12_ch_am1[18] ,_u0_u12_ch_am1[17] , _u0_u12_ch_am1[16] , _u0_u12_ch_am1[15] ,_u0_u12_ch_am1[14] , _u0_u12_ch_am1[13] , _u0_u12_ch_am1[12] ,_u0_u12_ch_am1[11] , _u0_u12_ch_am1[10] , _u0_u12_ch_am1[9] ,_u0_u12_ch_am1[8] , _u0_u12_ch_am1[7] , _u0_u12_ch_am1[6] ,_u0_u12_ch_am1[5] , _u0_u12_ch_am1[4] , _u0_u12_ch_am1[3] ,_u0_u12_ch_am1[2] , _u0_u12_ch_am1[1] , _u0_u12_ch_am1[0] ,_u0_u12_sw_pointer[31] , _u0_u12_sw_pointer[30] ,_u0_u12_sw_pointer[29] , _u0_u12_sw_pointer[28] ,_u0_u12_sw_pointer[27] , _u0_u12_sw_pointer[26] ,_u0_u12_sw_pointer[25] , _u0_u12_sw_pointer[24] ,_u0_u12_sw_pointer[23] , _u0_u12_sw_pointer[22] ,_u0_u12_sw_pointer[21] , _u0_u12_sw_pointer[20] ,_u0_u12_sw_pointer[19] , _u0_u12_sw_pointer[18] ,_u0_u12_sw_pointer[17] , _u0_u12_sw_pointer[16] ,_u0_u12_sw_pointer[15] , _u0_u12_sw_pointer[14] ,_u0_u12_sw_pointer[13] , _u0_u12_sw_pointer[12] ,_u0_u12_sw_pointer[11] , _u0_u12_sw_pointer[10] ,_u0_u12_sw_pointer[9] , _u0_u12_sw_pointer[8] ,_u0_u12_sw_pointer[7] , _u0_u12_sw_pointer[6] ,_u0_u12_sw_pointer[5] , _u0_u12_sw_pointer[4] ,_u0_u12_sw_pointer[3] , _u0_u12_sw_pointer[2] ,_u0_u12_sw_pointer[1] , _u0_u12_sw_pointer[0] , _u0_u12_ch_stop ,_u0_u12_ch_dis , _u0_u12_int , _u0_u13_pointer[31] ,_u0_u13_pointer[30] , _u0_u13_pointer[29] , _u0_u13_pointer[28] ,_u0_u13_pointer[27] , _u0_u13_pointer[26] , _u0_u13_pointer[25] ,_u0_u13_pointer[24] , _u0_u13_pointer[23] , _u0_u13_pointer[22] ,_u0_u13_pointer[21] , _u0_u13_pointer[20] , _u0_u13_pointer[19] ,_u0_u13_pointer[18] , _u0_u13_pointer[17] , _u0_u13_pointer[16] ,_u0_u13_pointer[15] , _u0_u13_pointer[14] , _u0_u13_pointer[13] ,_u0_u13_pointer[12] , _u0_u13_pointer[11] , _u0_u13_pointer[10] ,_u0_u13_pointer[9] , _u0_u13_pointer[8] , _u0_u13_pointer[7] ,_u0_u13_pointer[6] , _u0_u13_pointer[5] , _u0_u13_pointer[4] ,_u0_u13_pointer[3] , _u0_u13_pointer[2] , _u0_u13_pointer[1] ,_u0_u13_pointer[0] , _u0_u13_pointer_s[31] , _u0_u13_pointer_s[30] ,_u0_u13_pointer_s[29] , _u0_u13_pointer_s[28] ,_u0_u13_pointer_s[27] , _u0_u13_pointer_s[26] ,_u0_u13_pointer_s[25] , _u0_u13_pointer_s[24] ,_u0_u13_pointer_s[23] , _u0_u13_pointer_s[22] ,_u0_u13_pointer_s[21] , _u0_u13_pointer_s[20] ,_u0_u13_pointer_s[19] , _u0_u13_pointer_s[18] ,_u0_u13_pointer_s[17] , _u0_u13_pointer_s[16] ,_u0_u13_pointer_s[15] , _u0_u13_pointer_s[14] ,_u0_u13_pointer_s[13] , _u0_u13_pointer_s[12] ,_u0_u13_pointer_s[11] , _u0_u13_pointer_s[10] , _u0_u13_pointer_s[9] ,_u0_u13_pointer_s[8] , _u0_u13_pointer_s[7] , _u0_u13_pointer_s[6] ,_u0_u13_pointer_s[5] , _u0_u13_pointer_s[4] , _u0_u13_pointer_s[3] ,_u0_u13_pointer_s[2] , _u0_u13_pointer_s[1] , _u0_u13_pointer_s[0] ,_u0_u13_ch_csr[31] , _u0_u13_ch_csr[30] , _u0_u13_ch_csr[29] ,_u0_u13_ch_csr[28] , _u0_u13_ch_csr[27] , _u0_u13_ch_csr[26] ,_u0_u13_ch_csr[25] , _u0_u13_ch_csr[24] , _u0_u13_ch_csr[23] ,_u0_u13_ch_csr[22] , _u0_u13_ch_csr[21] , _u0_u13_ch_csr[20] ,_u0_u13_ch_csr[19] , _u0_u13_ch_csr[18] , _u0_u13_ch_csr[17] ,_u0_u13_ch_csr[16] , _u0_u13_ch_csr[15] , _u0_u13_ch_csr[14] ,_u0_u13_ch_csr[13] , _u0_u13_ch_csr[12] , _u0_u13_ch_csr[11] ,_u0_u13_ch_csr[10] , _u0_u13_ch_csr[9] , _u0_u13_ch_csr[8] ,_u0_u13_ch_csr[7] , _u0_u13_ch_csr[6] , _u0_u13_ch_csr[5] ,_u0_u13_ch_csr[4] , _u0_u13_ch_csr[3] , _u0_u13_ch_csr[2] ,_u0_u13_ch_csr[1] , _u0_u13_ch_csr[0] , _u0_u13_ch_txsz[31] ,_u0_u13_ch_txsz[30] , _u0_u13_ch_txsz[29] , _u0_u13_ch_txsz[28] ,_u0_u13_ch_txsz[27] , _u0_u13_ch_txsz[26] , _u0_u13_ch_txsz[25] ,_u0_u13_ch_txsz[24] , _u0_u13_ch_txsz[23] , _u0_u13_ch_txsz[22] ,_u0_u13_ch_txsz[21] , _u0_u13_ch_txsz[20] , _u0_u13_ch_txsz[19] ,_u0_u13_ch_txsz[18] , _u0_u13_ch_txsz[17] , _u0_u13_ch_txsz[16] ,_u0_u13_ch_txsz[15] , _u0_u13_ch_txsz[14] , _u0_u13_ch_txsz[13] ,_u0_u13_ch_txsz[12] , _u0_u13_ch_txsz[11] , _u0_u13_ch_txsz[10] ,_u0_u13_ch_txsz[9] , _u0_u13_ch_txsz[8] , _u0_u13_ch_txsz[7] ,_u0_u13_ch_txsz[6] , _u0_u13_ch_txsz[5] , _u0_u13_ch_txsz[4] ,_u0_u13_ch_txsz[3] , _u0_u13_ch_txsz[2] , _u0_u13_ch_txsz[1] ,_u0_u13_ch_txsz[0] , _u0_u13_ch_adr0[31] , _u0_u13_ch_adr0[30] ,_u0_u13_ch_adr0[29] , _u0_u13_ch_adr0[28] , _u0_u13_ch_adr0[27] ,_u0_u13_ch_adr0[26] , _u0_u13_ch_adr0[25] , _u0_u13_ch_adr0[24] ,_u0_u13_ch_adr0[23] , _u0_u13_ch_adr0[22] , _u0_u13_ch_adr0[21] ,_u0_u13_ch_adr0[20] , _u0_u13_ch_adr0[19] , _u0_u13_ch_adr0[18] ,_u0_u13_ch_adr0[17] , _u0_u13_ch_adr0[16] , _u0_u13_ch_adr0[15] ,_u0_u13_ch_adr0[14] , _u0_u13_ch_adr0[13] , _u0_u13_ch_adr0[12] ,_u0_u13_ch_adr0[11] , _u0_u13_ch_adr0[10] , _u0_u13_ch_adr0[9] ,_u0_u13_ch_adr0[8] , _u0_u13_ch_adr0[7] , _u0_u13_ch_adr0[6] ,_u0_u13_ch_adr0[5] , _u0_u13_ch_adr0[4] , _u0_u13_ch_adr0[3] ,_u0_u13_ch_adr0[2] , _u0_u13_ch_adr0[1] , _u0_u13_ch_adr0[0] ,_u0_u13_ch_adr1[31] , _u0_u13_ch_adr1[30] , _u0_u13_ch_adr1[29] ,_u0_u13_ch_adr1[28] , _u0_u13_ch_adr1[27] , _u0_u13_ch_adr1[26] ,_u0_u13_ch_adr1[25] , _u0_u13_ch_adr1[24] , _u0_u13_ch_adr1[23] ,_u0_u13_ch_adr1[22] , _u0_u13_ch_adr1[21] , _u0_u13_ch_adr1[20] ,_u0_u13_ch_adr1[19] , _u0_u13_ch_adr1[18] , _u0_u13_ch_adr1[17] ,_u0_u13_ch_adr1[16] , _u0_u13_ch_adr1[15] , _u0_u13_ch_adr1[14] ,_u0_u13_ch_adr1[13] , _u0_u13_ch_adr1[12] , _u0_u13_ch_adr1[11] ,_u0_u13_ch_adr1[10] , _u0_u13_ch_adr1[9] , _u0_u13_ch_adr1[8] ,_u0_u13_ch_adr1[7] , _u0_u13_ch_adr1[6] , _u0_u13_ch_adr1[5] ,_u0_u13_ch_adr1[4] , _u0_u13_ch_adr1[3] , _u0_u13_ch_adr1[2] ,_u0_u13_ch_adr1[1] , _u0_u13_ch_adr1[0] , _u0_u13_ch_am0[31] ,_u0_u13_ch_am0[30] , _u0_u13_ch_am0[29] , _u0_u13_ch_am0[28] ,_u0_u13_ch_am0[27] , _u0_u13_ch_am0[26] , _u0_u13_ch_am0[25] ,_u0_u13_ch_am0[24] , _u0_u13_ch_am0[23] , _u0_u13_ch_am0[22] ,_u0_u13_ch_am0[21] , _u0_u13_ch_am0[20] , _u0_u13_ch_am0[19] ,_u0_u13_ch_am0[18] , _u0_u13_ch_am0[17] , _u0_u13_ch_am0[16] ,_u0_u13_ch_am0[15] , _u0_u13_ch_am0[14] , _u0_u13_ch_am0[13] ,_u0_u13_ch_am0[12] , _u0_u13_ch_am0[11] , _u0_u13_ch_am0[10] ,_u0_u13_ch_am0[9] , _u0_u13_ch_am0[8] , _u0_u13_ch_am0[7] ,_u0_u13_ch_am0[6] , _u0_u13_ch_am0[5] , _u0_u13_ch_am0[4] ,_u0_u13_ch_am0[3] , _u0_u13_ch_am0[2] , _u0_u13_ch_am0[1] ,_u0_u13_ch_am0[0] , _u0_u13_ch_am1[31] , _u0_u13_ch_am1[30] ,_u0_u13_ch_am1[29] , _u0_u13_ch_am1[28] , _u0_u13_ch_am1[27] ,_u0_u13_ch_am1[26] , _u0_u13_ch_am1[25] , _u0_u13_ch_am1[24] ,_u0_u13_ch_am1[23] , _u0_u13_ch_am1[22] , _u0_u13_ch_am1[21] ,_u0_u13_ch_am1[20] , _u0_u13_ch_am1[19] , _u0_u13_ch_am1[18] ,_u0_u13_ch_am1[17] , _u0_u13_ch_am1[16] , _u0_u13_ch_am1[15] ,_u0_u13_ch_am1[14] , _u0_u13_ch_am1[13] , _u0_u13_ch_am1[12] ,_u0_u13_ch_am1[11] , _u0_u13_ch_am1[10] , _u0_u13_ch_am1[9] ,_u0_u13_ch_am1[8] , _u0_u13_ch_am1[7] , _u0_u13_ch_am1[6] ,_u0_u13_ch_am1[5] , _u0_u13_ch_am1[4] , _u0_u13_ch_am1[3] ,_u0_u13_ch_am1[2] , _u0_u13_ch_am1[1] , _u0_u13_ch_am1[0] ,_u0_u13_sw_pointer[31] , _u0_u13_sw_pointer[30] ,_u0_u13_sw_pointer[29] , _u0_u13_sw_pointer[28] ,_u0_u13_sw_pointer[27] , _u0_u13_sw_pointer[26] ,_u0_u13_sw_pointer[25] , _u0_u13_sw_pointer[24] ,_u0_u13_sw_pointer[23] , _u0_u13_sw_pointer[22] ,_u0_u13_sw_pointer[21] , _u0_u13_sw_pointer[20] ,_u0_u13_sw_pointer[19] , _u0_u13_sw_pointer[18] ,_u0_u13_sw_pointer[17] , _u0_u13_sw_pointer[16] ,_u0_u13_sw_pointer[15] , _u0_u13_sw_pointer[14] ,_u0_u13_sw_pointer[13] , _u0_u13_sw_pointer[12] ,_u0_u13_sw_pointer[11] , _u0_u13_sw_pointer[10] ,_u0_u13_sw_pointer[9] , _u0_u13_sw_pointer[8] ,_u0_u13_sw_pointer[7] , _u0_u13_sw_pointer[6] ,_u0_u13_sw_pointer[5] , _u0_u13_sw_pointer[4] ,_u0_u13_sw_pointer[3] , _u0_u13_sw_pointer[2] ,_u0_u13_sw_pointer[1] , _u0_u13_sw_pointer[0] , _u0_u13_ch_stop ,_u0_u13_ch_dis , _u0_u13_int , _u0_u14_pointer[31] ,_u0_u14_pointer[30] , _u0_u14_pointer[29] , _u0_u14_pointer[28] ,_u0_u14_pointer[27] , _u0_u14_pointer[26] , _u0_u14_pointer[25] ,_u0_u14_pointer[24] , _u0_u14_pointer[23] , _u0_u14_pointer[22] ,_u0_u14_pointer[21] , _u0_u14_pointer[20] , _u0_u14_pointer[19] ,_u0_u14_pointer[18] , _u0_u14_pointer[17] , _u0_u14_pointer[16] ,_u0_u14_pointer[15] , _u0_u14_pointer[14] , _u0_u14_pointer[13] ,_u0_u14_pointer[12] , _u0_u14_pointer[11] , _u0_u14_pointer[10] ,_u0_u14_pointer[9] , _u0_u14_pointer[8] , _u0_u14_pointer[7] ,_u0_u14_pointer[6] , _u0_u14_pointer[5] , _u0_u14_pointer[4] ,_u0_u14_pointer[3] , _u0_u14_pointer[2] , _u0_u14_pointer[1] ,_u0_u14_pointer[0] , _u0_u14_pointer_s[31] , _u0_u14_pointer_s[30] ,_u0_u14_pointer_s[29] , _u0_u14_pointer_s[28] ,_u0_u14_pointer_s[27] , _u0_u14_pointer_s[26] ,_u0_u14_pointer_s[25] , _u0_u14_pointer_s[24] ,_u0_u14_pointer_s[23] , _u0_u14_pointer_s[22] ,_u0_u14_pointer_s[21] , _u0_u14_pointer_s[20] ,_u0_u14_pointer_s[19] , _u0_u14_pointer_s[18] ,_u0_u14_pointer_s[17] , _u0_u14_pointer_s[16] ,_u0_u14_pointer_s[15] , _u0_u14_pointer_s[14] ,_u0_u14_pointer_s[13] , _u0_u14_pointer_s[12] ,_u0_u14_pointer_s[11] , _u0_u14_pointer_s[10] , _u0_u14_pointer_s[9] ,_u0_u14_pointer_s[8] , _u0_u14_pointer_s[7] , _u0_u14_pointer_s[6] ,_u0_u14_pointer_s[5] , _u0_u14_pointer_s[4] , _u0_u14_pointer_s[3] ,_u0_u14_pointer_s[2] , _u0_u14_pointer_s[1] , _u0_u14_pointer_s[0] ,_u0_u14_ch_csr[31] , _u0_u14_ch_csr[30] , _u0_u14_ch_csr[29] ,_u0_u14_ch_csr[28] , _u0_u14_ch_csr[27] , _u0_u14_ch_csr[26] ,_u0_u14_ch_csr[25] , _u0_u14_ch_csr[24] , _u0_u14_ch_csr[23] ,_u0_u14_ch_csr[22] , _u0_u14_ch_csr[21] , _u0_u14_ch_csr[20] ,_u0_u14_ch_csr[19] , _u0_u14_ch_csr[18] , _u0_u14_ch_csr[17] ,_u0_u14_ch_csr[16] , _u0_u14_ch_csr[15] , _u0_u14_ch_csr[14] ,_u0_u14_ch_csr[13] , _u0_u14_ch_csr[12] , _u0_u14_ch_csr[11] ,_u0_u14_ch_csr[10] , _u0_u14_ch_csr[9] , _u0_u14_ch_csr[8] ,_u0_u14_ch_csr[7] , _u0_u14_ch_csr[6] , _u0_u14_ch_csr[5] ,_u0_u14_ch_csr[4] , _u0_u14_ch_csr[3] , _u0_u14_ch_csr[2] ,_u0_u14_ch_csr[1] , _u0_u14_ch_csr[0] , _u0_u14_ch_txsz[31] ,_u0_u14_ch_txsz[30] , _u0_u14_ch_txsz[29] , _u0_u14_ch_txsz[28] ,_u0_u14_ch_txsz[27] , _u0_u14_ch_txsz[26] , _u0_u14_ch_txsz[25] ,_u0_u14_ch_txsz[24] , _u0_u14_ch_txsz[23] , _u0_u14_ch_txsz[22] ,_u0_u14_ch_txsz[21] , _u0_u14_ch_txsz[20] , _u0_u14_ch_txsz[19] ,_u0_u14_ch_txsz[18] , _u0_u14_ch_txsz[17] , _u0_u14_ch_txsz[16] ,_u0_u14_ch_txsz[15] , _u0_u14_ch_txsz[14] , _u0_u14_ch_txsz[13] ,_u0_u14_ch_txsz[12] , _u0_u14_ch_txsz[11] , _u0_u14_ch_txsz[10] ,_u0_u14_ch_txsz[9] , _u0_u14_ch_txsz[8] , _u0_u14_ch_txsz[7] ,_u0_u14_ch_txsz[6] , _u0_u14_ch_txsz[5] , _u0_u14_ch_txsz[4] ,_u0_u14_ch_txsz[3] , _u0_u14_ch_txsz[2] , _u0_u14_ch_txsz[1] ,_u0_u14_ch_txsz[0] , _u0_u14_ch_adr0[31] , _u0_u14_ch_adr0[30] ,_u0_u14_ch_adr0[29] , _u0_u14_ch_adr0[28] , _u0_u14_ch_adr0[27] ,_u0_u14_ch_adr0[26] , _u0_u14_ch_adr0[25] , _u0_u14_ch_adr0[24] ,_u0_u14_ch_adr0[23] , _u0_u14_ch_adr0[22] , _u0_u14_ch_adr0[21] ,_u0_u14_ch_adr0[20] , _u0_u14_ch_adr0[19] , _u0_u14_ch_adr0[18] ,_u0_u14_ch_adr0[17] , _u0_u14_ch_adr0[16] , _u0_u14_ch_adr0[15] ,_u0_u14_ch_adr0[14] , _u0_u14_ch_adr0[13] , _u0_u14_ch_adr0[12] ,_u0_u14_ch_adr0[11] , _u0_u14_ch_adr0[10] , _u0_u14_ch_adr0[9] ,_u0_u14_ch_adr0[8] , _u0_u14_ch_adr0[7] , _u0_u14_ch_adr0[6] ,_u0_u14_ch_adr0[5] , _u0_u14_ch_adr0[4] , _u0_u14_ch_adr0[3] ,_u0_u14_ch_adr0[2] , _u0_u14_ch_adr0[1] , _u0_u14_ch_adr0[0] ,_u0_u14_ch_adr1[31] , _u0_u14_ch_adr1[30] , _u0_u14_ch_adr1[29] ,_u0_u14_ch_adr1[28] , _u0_u14_ch_adr1[27] , _u0_u14_ch_adr1[26] ,_u0_u14_ch_adr1[25] , _u0_u14_ch_adr1[24] , _u0_u14_ch_adr1[23] ,_u0_u14_ch_adr1[22] , _u0_u14_ch_adr1[21] , _u0_u14_ch_adr1[20] ,_u0_u14_ch_adr1[19] , _u0_u14_ch_adr1[18] , _u0_u14_ch_adr1[17] ,_u0_u14_ch_adr1[16] , _u0_u14_ch_adr1[15] , _u0_u14_ch_adr1[14] ,_u0_u14_ch_adr1[13] , _u0_u14_ch_adr1[12] , _u0_u14_ch_adr1[11] ,_u0_u14_ch_adr1[10] , _u0_u14_ch_adr1[9] , _u0_u14_ch_adr1[8] ,_u0_u14_ch_adr1[7] , _u0_u14_ch_adr1[6] , _u0_u14_ch_adr1[5] ,_u0_u14_ch_adr1[4] , _u0_u14_ch_adr1[3] , _u0_u14_ch_adr1[2] ,_u0_u14_ch_adr1[1] , _u0_u14_ch_adr1[0] , _u0_u14_ch_am0[31] ,_u0_u14_ch_am0[30] , _u0_u14_ch_am0[29] , _u0_u14_ch_am0[28] ,_u0_u14_ch_am0[27] , _u0_u14_ch_am0[26] , _u0_u14_ch_am0[25] ,_u0_u14_ch_am0[24] , _u0_u14_ch_am0[23] , _u0_u14_ch_am0[22] ,_u0_u14_ch_am0[21] , _u0_u14_ch_am0[20] , _u0_u14_ch_am0[19] ,_u0_u14_ch_am0[18] , _u0_u14_ch_am0[17] , _u0_u14_ch_am0[16] ,_u0_u14_ch_am0[15] , _u0_u14_ch_am0[14] , _u0_u14_ch_am0[13] ,_u0_u14_ch_am0[12] , _u0_u14_ch_am0[11] , _u0_u14_ch_am0[10] ,_u0_u14_ch_am0[9] , _u0_u14_ch_am0[8] , _u0_u14_ch_am0[7] ,_u0_u14_ch_am0[6] , _u0_u14_ch_am0[5] , _u0_u14_ch_am0[4] ,_u0_u14_ch_am0[3] , _u0_u14_ch_am0[2] , _u0_u14_ch_am0[1] ,_u0_u14_ch_am0[0] , _u0_u14_ch_am1[31] , _u0_u14_ch_am1[30] ,_u0_u14_ch_am1[29] , _u0_u14_ch_am1[28] , _u0_u14_ch_am1[27] ,_u0_u14_ch_am1[26] , _u0_u14_ch_am1[25] , _u0_u14_ch_am1[24] ,_u0_u14_ch_am1[23] , _u0_u14_ch_am1[22] , _u0_u14_ch_am1[21] ,_u0_u14_ch_am1[20] , _u0_u14_ch_am1[19] , _u0_u14_ch_am1[18] ,_u0_u14_ch_am1[17] , _u0_u14_ch_am1[16] , _u0_u14_ch_am1[15] ,_u0_u14_ch_am1[14] , _u0_u14_ch_am1[13] , _u0_u14_ch_am1[12] ,_u0_u14_ch_am1[11] , _u0_u14_ch_am1[10] , _u0_u14_ch_am1[9] ,_u0_u14_ch_am1[8] , _u0_u14_ch_am1[7] , _u0_u14_ch_am1[6] ,_u0_u14_ch_am1[5] , _u0_u14_ch_am1[4] , _u0_u14_ch_am1[3] ,_u0_u14_ch_am1[2] , _u0_u14_ch_am1[1] , _u0_u14_ch_am1[0] ,_u0_u14_sw_pointer[31] , _u0_u14_sw_pointer[30] ,_u0_u14_sw_pointer[29] , _u0_u14_sw_pointer[28] ,_u0_u14_sw_pointer[27] , _u0_u14_sw_pointer[26] ,_u0_u14_sw_pointer[25] , _u0_u14_sw_pointer[24] ,_u0_u14_sw_pointer[23] , _u0_u14_sw_pointer[22] ,_u0_u14_sw_pointer[21] , _u0_u14_sw_pointer[20] ,_u0_u14_sw_pointer[19] , _u0_u14_sw_pointer[18] ,_u0_u14_sw_pointer[17] , _u0_u14_sw_pointer[16] ,_u0_u14_sw_pointer[15] , _u0_u14_sw_pointer[14] ,_u0_u14_sw_pointer[13] , _u0_u14_sw_pointer[12] ,_u0_u14_sw_pointer[11] , _u0_u14_sw_pointer[10] ,_u0_u14_sw_pointer[9] , _u0_u14_sw_pointer[8] ,_u0_u14_sw_pointer[7] , _u0_u14_sw_pointer[6] ,_u0_u14_sw_pointer[5] , _u0_u14_sw_pointer[4] ,_u0_u14_sw_pointer[3] , _u0_u14_sw_pointer[2] ,_u0_u14_sw_pointer[1] , _u0_u14_sw_pointer[0] , _u0_u14_ch_stop ,_u0_u14_ch_dis , _u0_u14_int , _u0_u15_pointer[31] ,_u0_u15_pointer[30] , _u0_u15_pointer[29] , _u0_u15_pointer[28] ,_u0_u15_pointer[27] , _u0_u15_pointer[26] , _u0_u15_pointer[25] ,_u0_u15_pointer[24] , _u0_u15_pointer[23] , _u0_u15_pointer[22] ,_u0_u15_pointer[21] , _u0_u15_pointer[20] , _u0_u15_pointer[19] ,_u0_u15_pointer[18] , _u0_u15_pointer[17] , _u0_u15_pointer[16] ,_u0_u15_pointer[15] , _u0_u15_pointer[14] , _u0_u15_pointer[13] ,_u0_u15_pointer[12] , _u0_u15_pointer[11] , _u0_u15_pointer[10] ,_u0_u15_pointer[9] , _u0_u15_pointer[8] , _u0_u15_pointer[7] ,_u0_u15_pointer[6] , _u0_u15_pointer[5] , _u0_u15_pointer[4] ,_u0_u15_pointer[3] , _u0_u15_pointer[2] , _u0_u15_pointer[1] ,_u0_u15_pointer[0] , _u0_u15_pointer_s[31] , _u0_u15_pointer_s[30] ,_u0_u15_pointer_s[29] , _u0_u15_pointer_s[28] ,_u0_u15_pointer_s[27] , _u0_u15_pointer_s[26] ,_u0_u15_pointer_s[25] , _u0_u15_pointer_s[24] ,_u0_u15_pointer_s[23] , _u0_u15_pointer_s[22] ,_u0_u15_pointer_s[21] , _u0_u15_pointer_s[20] ,_u0_u15_pointer_s[19] , _u0_u15_pointer_s[18] ,_u0_u15_pointer_s[17] , _u0_u15_pointer_s[16] ,_u0_u15_pointer_s[15] , _u0_u15_pointer_s[14] ,_u0_u15_pointer_s[13] , _u0_u15_pointer_s[12] ,_u0_u15_pointer_s[11] , _u0_u15_pointer_s[10] , _u0_u15_pointer_s[9] ,_u0_u15_pointer_s[8] , _u0_u15_pointer_s[7] , _u0_u15_pointer_s[6] ,_u0_u15_pointer_s[5] , _u0_u15_pointer_s[4] , _u0_u15_pointer_s[3] ,_u0_u15_pointer_s[2] , _u0_u15_pointer_s[1] , _u0_u15_pointer_s[0] ,_u0_u15_ch_csr[31] , _u0_u15_ch_csr[30] , _u0_u15_ch_csr[29] ,_u0_u15_ch_csr[28] , _u0_u15_ch_csr[27] , _u0_u15_ch_csr[26] ,_u0_u15_ch_csr[25] , _u0_u15_ch_csr[24] , _u0_u15_ch_csr[23] ,_u0_u15_ch_csr[22] , _u0_u15_ch_csr[21] , _u0_u15_ch_csr[20] ,_u0_u15_ch_csr[19] , _u0_u15_ch_csr[18] , _u0_u15_ch_csr[17] ,_u0_u15_ch_csr[16] , _u0_u15_ch_csr[15] , _u0_u15_ch_csr[14] ,_u0_u15_ch_csr[13] , _u0_u15_ch_csr[12] , _u0_u15_ch_csr[11] ,_u0_u15_ch_csr[10] , _u0_u15_ch_csr[9] , _u0_u15_ch_csr[8] ,_u0_u15_ch_csr[7] , _u0_u15_ch_csr[6] , _u0_u15_ch_csr[5] ,_u0_u15_ch_csr[4] , _u0_u15_ch_csr[3] , _u0_u15_ch_csr[2] ,_u0_u15_ch_csr[1] , _u0_u15_ch_csr[0] , _u0_u15_ch_txsz[31] ,_u0_u15_ch_txsz[30] , _u0_u15_ch_txsz[29] , _u0_u15_ch_txsz[28] ,_u0_u15_ch_txsz[27] , _u0_u15_ch_txsz[26] , _u0_u15_ch_txsz[25] ,_u0_u15_ch_txsz[24] , _u0_u15_ch_txsz[23] , _u0_u15_ch_txsz[22] ,_u0_u15_ch_txsz[21] , _u0_u15_ch_txsz[20] , _u0_u15_ch_txsz[19] ,_u0_u15_ch_txsz[18] , _u0_u15_ch_txsz[17] , _u0_u15_ch_txsz[16] ,_u0_u15_ch_txsz[15] , _u0_u15_ch_txsz[14] , _u0_u15_ch_txsz[13] ,_u0_u15_ch_txsz[12] , _u0_u15_ch_txsz[11] , _u0_u15_ch_txsz[10] ,_u0_u15_ch_txsz[9] , _u0_u15_ch_txsz[8] , _u0_u15_ch_txsz[7] ,_u0_u15_ch_txsz[6] , _u0_u15_ch_txsz[5] , _u0_u15_ch_txsz[4] ,_u0_u15_ch_txsz[3] , _u0_u15_ch_txsz[2] , _u0_u15_ch_txsz[1] ,_u0_u15_ch_txsz[0] , _u0_u15_ch_adr0[31] , _u0_u15_ch_adr0[30] ,_u0_u15_ch_adr0[29] , _u0_u15_ch_adr0[28] , _u0_u15_ch_adr0[27] ,_u0_u15_ch_adr0[26] , _u0_u15_ch_adr0[25] , _u0_u15_ch_adr0[24] ,_u0_u15_ch_adr0[23] , _u0_u15_ch_adr0[22] , _u0_u15_ch_adr0[21] ,_u0_u15_ch_adr0[20] , _u0_u15_ch_adr0[19] , _u0_u15_ch_adr0[18] ,_u0_u15_ch_adr0[17] , _u0_u15_ch_adr0[16] , _u0_u15_ch_adr0[15] ,_u0_u15_ch_adr0[14] , _u0_u15_ch_adr0[13] , _u0_u15_ch_adr0[12] ,_u0_u15_ch_adr0[11] , _u0_u15_ch_adr0[10] , _u0_u15_ch_adr0[9] ,_u0_u15_ch_adr0[8] , _u0_u15_ch_adr0[7] , _u0_u15_ch_adr0[6] ,_u0_u15_ch_adr0[5] , _u0_u15_ch_adr0[4] , _u0_u15_ch_adr0[3] ,_u0_u15_ch_adr0[2] , _u0_u15_ch_adr0[1] , _u0_u15_ch_adr0[0] ,_u0_u15_ch_adr1[31] , _u0_u15_ch_adr1[30] , _u0_u15_ch_adr1[29] ,_u0_u15_ch_adr1[28] , _u0_u15_ch_adr1[27] , _u0_u15_ch_adr1[26] ,_u0_u15_ch_adr1[25] , _u0_u15_ch_adr1[24] , _u0_u15_ch_adr1[23] ,_u0_u15_ch_adr1[22] , _u0_u15_ch_adr1[21] , _u0_u15_ch_adr1[20] ,_u0_u15_ch_adr1[19] , _u0_u15_ch_adr1[18] , _u0_u15_ch_adr1[17] ,_u0_u15_ch_adr1[16] , _u0_u15_ch_adr1[15] , _u0_u15_ch_adr1[14] ,_u0_u15_ch_adr1[13] , _u0_u15_ch_adr1[12] , _u0_u15_ch_adr1[11] ,_u0_u15_ch_adr1[10] , _u0_u15_ch_adr1[9] , _u0_u15_ch_adr1[8] ,_u0_u15_ch_adr1[7] , _u0_u15_ch_adr1[6] , _u0_u15_ch_adr1[5] ,_u0_u15_ch_adr1[4] , _u0_u15_ch_adr1[3] , _u0_u15_ch_adr1[2] ,_u0_u15_ch_adr1[1] , _u0_u15_ch_adr1[0] , _u0_u15_ch_am0[31] ,_u0_u15_ch_am0[30] , _u0_u15_ch_am0[29] , _u0_u15_ch_am0[28] ,_u0_u15_ch_am0[27] , _u0_u15_ch_am0[26] , _u0_u15_ch_am0[25] ,_u0_u15_ch_am0[24] , _u0_u15_ch_am0[23] , _u0_u15_ch_am0[22] ,_u0_u15_ch_am0[21] , _u0_u15_ch_am0[20] , _u0_u15_ch_am0[19] ,_u0_u15_ch_am0[18] , _u0_u15_ch_am0[17] , _u0_u15_ch_am0[16] ,_u0_u15_ch_am0[15] , _u0_u15_ch_am0[14] , _u0_u15_ch_am0[13] ,_u0_u15_ch_am0[12] , _u0_u15_ch_am0[11] , _u0_u15_ch_am0[10] ,_u0_u15_ch_am0[9] , _u0_u15_ch_am0[8] , _u0_u15_ch_am0[7] ,_u0_u15_ch_am0[6] , _u0_u15_ch_am0[5] , _u0_u15_ch_am0[4] ,_u0_u15_ch_am0[3] , _u0_u15_ch_am0[2] , _u0_u15_ch_am0[1] ,_u0_u15_ch_am0[0] , _u0_u15_ch_am1[31] , _u0_u15_ch_am1[30] ,_u0_u15_ch_am1[29] , _u0_u15_ch_am1[28] , _u0_u15_ch_am1[27] ,_u0_u15_ch_am1[26] , _u0_u15_ch_am1[25] , _u0_u15_ch_am1[24] ,_u0_u15_ch_am1[23] , _u0_u15_ch_am1[22] , _u0_u15_ch_am1[21] ,_u0_u15_ch_am1[20] , _u0_u15_ch_am1[19] , _u0_u15_ch_am1[18] ,_u0_u15_ch_am1[17] , _u0_u15_ch_am1[16] , _u0_u15_ch_am1[15] ,_u0_u15_ch_am1[14] , _u0_u15_ch_am1[13] , _u0_u15_ch_am1[12] ,_u0_u15_ch_am1[11] , _u0_u15_ch_am1[10] , _u0_u15_ch_am1[9] ,_u0_u15_ch_am1[8] , _u0_u15_ch_am1[7] , _u0_u15_ch_am1[6] ,_u0_u15_ch_am1[5] , _u0_u15_ch_am1[4] , _u0_u15_ch_am1[3] ,_u0_u15_ch_am1[2] , _u0_u15_ch_am1[1] , _u0_u15_ch_am1[0] ,_u0_u15_sw_pointer[31] , _u0_u15_sw_pointer[30] ,_u0_u15_sw_pointer[29] , _u0_u15_sw_pointer[28] ,_u0_u15_sw_pointer[27] , _u0_u15_sw_pointer[26] ,_u0_u15_sw_pointer[25] , _u0_u15_sw_pointer[24] ,_u0_u15_sw_pointer[23] , _u0_u15_sw_pointer[22] ,_u0_u15_sw_pointer[21] , _u0_u15_sw_pointer[20] ,_u0_u15_sw_pointer[19] , _u0_u15_sw_pointer[18] ,_u0_u15_sw_pointer[17] , _u0_u15_sw_pointer[16] ,_u0_u15_sw_pointer[15] , _u0_u15_sw_pointer[14] ,_u0_u15_sw_pointer[13] , _u0_u15_sw_pointer[12] ,_u0_u15_sw_pointer[11] , _u0_u15_sw_pointer[10] ,_u0_u15_sw_pointer[9] , _u0_u15_sw_pointer[8] ,_u0_u15_sw_pointer[7] , _u0_u15_sw_pointer[6] ,_u0_u15_sw_pointer[5] , _u0_u15_sw_pointer[4] ,_u0_u15_sw_pointer[3] , _u0_u15_sw_pointer[2] ,_u0_u15_sw_pointer[1] , _u0_u15_sw_pointer[0] , _u0_u15_ch_stop ,_u0_u15_ch_dis , _u0_u15_int , _u0_u16_pointer[31] ,_u0_u16_pointer[30] , _u0_u16_pointer[29] , _u0_u16_pointer[28] ,_u0_u16_pointer[27] , _u0_u16_pointer[26] , _u0_u16_pointer[25] ,_u0_u16_pointer[24] , _u0_u16_pointer[23] , _u0_u16_pointer[22] ,_u0_u16_pointer[21] , _u0_u16_pointer[20] , _u0_u16_pointer[19] ,_u0_u16_pointer[18] , _u0_u16_pointer[17] , _u0_u16_pointer[16] ,_u0_u16_pointer[15] , _u0_u16_pointer[14] , _u0_u16_pointer[13] ,_u0_u16_pointer[12] , _u0_u16_pointer[11] , _u0_u16_pointer[10] ,_u0_u16_pointer[9] , _u0_u16_pointer[8] , _u0_u16_pointer[7] ,_u0_u16_pointer[6] , _u0_u16_pointer[5] , _u0_u16_pointer[4] ,_u0_u16_pointer[3] , _u0_u16_pointer[2] , _u0_u16_pointer[1] ,_u0_u16_pointer[0] , _u0_u16_pointer_s[31] , _u0_u16_pointer_s[30] ,_u0_u16_pointer_s[29] , _u0_u16_pointer_s[28] ,_u0_u16_pointer_s[27] , _u0_u16_pointer_s[26] ,_u0_u16_pointer_s[25] , _u0_u16_pointer_s[24] ,_u0_u16_pointer_s[23] , _u0_u16_pointer_s[22] ,_u0_u16_pointer_s[21] , _u0_u16_pointer_s[20] ,_u0_u16_pointer_s[19] , _u0_u16_pointer_s[18] ,_u0_u16_pointer_s[17] , _u0_u16_pointer_s[16] ,_u0_u16_pointer_s[15] , _u0_u16_pointer_s[14] ,_u0_u16_pointer_s[13] , _u0_u16_pointer_s[12] ,_u0_u16_pointer_s[11] , _u0_u16_pointer_s[10] , _u0_u16_pointer_s[9] ,_u0_u16_pointer_s[8] , _u0_u16_pointer_s[7] , _u0_u16_pointer_s[6] ,_u0_u16_pointer_s[5] , _u0_u16_pointer_s[4] , _u0_u16_pointer_s[3] ,_u0_u16_pointer_s[2] , _u0_u16_pointer_s[1] , _u0_u16_pointer_s[0] ,_u0_u16_ch_csr[31] , _u0_u16_ch_csr[30] , _u0_u16_ch_csr[29] ,_u0_u16_ch_csr[28] , _u0_u16_ch_csr[27] , _u0_u16_ch_csr[26] ,_u0_u16_ch_csr[25] , _u0_u16_ch_csr[24] , _u0_u16_ch_csr[23] ,_u0_u16_ch_csr[22] , _u0_u16_ch_csr[21] , _u0_u16_ch_csr[20] ,_u0_u16_ch_csr[19] , _u0_u16_ch_csr[18] , _u0_u16_ch_csr[17] ,_u0_u16_ch_csr[16] , _u0_u16_ch_csr[15] , _u0_u16_ch_csr[14] ,_u0_u16_ch_csr[13] , _u0_u16_ch_csr[12] , _u0_u16_ch_csr[11] ,_u0_u16_ch_csr[10] , _u0_u16_ch_csr[9] , _u0_u16_ch_csr[8] ,_u0_u16_ch_csr[7] , _u0_u16_ch_csr[6] , _u0_u16_ch_csr[5] ,_u0_u16_ch_csr[4] , _u0_u16_ch_csr[3] , _u0_u16_ch_csr[2] ,_u0_u16_ch_csr[1] , _u0_u16_ch_csr[0] , _u0_u16_ch_txsz[31] ,_u0_u16_ch_txsz[30] , _u0_u16_ch_txsz[29] , _u0_u16_ch_txsz[28] ,_u0_u16_ch_txsz[27] , _u0_u16_ch_txsz[26] , _u0_u16_ch_txsz[25] ,_u0_u16_ch_txsz[24] , _u0_u16_ch_txsz[23] , _u0_u16_ch_txsz[22] ,_u0_u16_ch_txsz[21] , _u0_u16_ch_txsz[20] , _u0_u16_ch_txsz[19] ,_u0_u16_ch_txsz[18] , _u0_u16_ch_txsz[17] , _u0_u16_ch_txsz[16] ,_u0_u16_ch_txsz[15] , _u0_u16_ch_txsz[14] , _u0_u16_ch_txsz[13] ,_u0_u16_ch_txsz[12] , _u0_u16_ch_txsz[11] , _u0_u16_ch_txsz[10] ,_u0_u16_ch_txsz[9] , _u0_u16_ch_txsz[8] , _u0_u16_ch_txsz[7] ,_u0_u16_ch_txsz[6] , _u0_u16_ch_txsz[5] , _u0_u16_ch_txsz[4] ,_u0_u16_ch_txsz[3] , _u0_u16_ch_txsz[2] , _u0_u16_ch_txsz[1] ,_u0_u16_ch_txsz[0] , _u0_u16_ch_adr0[31] , _u0_u16_ch_adr0[30] ,_u0_u16_ch_adr0[29] , _u0_u16_ch_adr0[28] , _u0_u16_ch_adr0[27] ,_u0_u16_ch_adr0[26] , _u0_u16_ch_adr0[25] , _u0_u16_ch_adr0[24] ,_u0_u16_ch_adr0[23] , _u0_u16_ch_adr0[22] , _u0_u16_ch_adr0[21] ,_u0_u16_ch_adr0[20] , _u0_u16_ch_adr0[19] , _u0_u16_ch_adr0[18] ,_u0_u16_ch_adr0[17] , _u0_u16_ch_adr0[16] , _u0_u16_ch_adr0[15] ,_u0_u16_ch_adr0[14] , _u0_u16_ch_adr0[13] , _u0_u16_ch_adr0[12] ,_u0_u16_ch_adr0[11] , _u0_u16_ch_adr0[10] , _u0_u16_ch_adr0[9] ,_u0_u16_ch_adr0[8] , _u0_u16_ch_adr0[7] , _u0_u16_ch_adr0[6] ,_u0_u16_ch_adr0[5] , _u0_u16_ch_adr0[4] , _u0_u16_ch_adr0[3] ,_u0_u16_ch_adr0[2] , _u0_u16_ch_adr0[1] , _u0_u16_ch_adr0[0] ,_u0_u16_ch_adr1[31] , _u0_u16_ch_adr1[30] , _u0_u16_ch_adr1[29] ,_u0_u16_ch_adr1[28] , _u0_u16_ch_adr1[27] , _u0_u16_ch_adr1[26] ,_u0_u16_ch_adr1[25] , _u0_u16_ch_adr1[24] , _u0_u16_ch_adr1[23] ,_u0_u16_ch_adr1[22] , _u0_u16_ch_adr1[21] , _u0_u16_ch_adr1[20] ,_u0_u16_ch_adr1[19] , _u0_u16_ch_adr1[18] , _u0_u16_ch_adr1[17] ,_u0_u16_ch_adr1[16] , _u0_u16_ch_adr1[15] , _u0_u16_ch_adr1[14] ,_u0_u16_ch_adr1[13] , _u0_u16_ch_adr1[12] , _u0_u16_ch_adr1[11] ,_u0_u16_ch_adr1[10] , _u0_u16_ch_adr1[9] , _u0_u16_ch_adr1[8] ,_u0_u16_ch_adr1[7] , _u0_u16_ch_adr1[6] , _u0_u16_ch_adr1[5] ,_u0_u16_ch_adr1[4] , _u0_u16_ch_adr1[3] , _u0_u16_ch_adr1[2] ,_u0_u16_ch_adr1[1] , _u0_u16_ch_adr1[0] , _u0_u16_ch_am0[31] ,_u0_u16_ch_am0[30] , _u0_u16_ch_am0[29] , _u0_u16_ch_am0[28] ,_u0_u16_ch_am0[27] , _u0_u16_ch_am0[26] , _u0_u16_ch_am0[25] ,_u0_u16_ch_am0[24] , _u0_u16_ch_am0[23] , _u0_u16_ch_am0[22] ,_u0_u16_ch_am0[21] , _u0_u16_ch_am0[20] , _u0_u16_ch_am0[19] ,_u0_u16_ch_am0[18] , _u0_u16_ch_am0[17] , _u0_u16_ch_am0[16] ,_u0_u16_ch_am0[15] , _u0_u16_ch_am0[14] , _u0_u16_ch_am0[13] ,_u0_u16_ch_am0[12] , _u0_u16_ch_am0[11] , _u0_u16_ch_am0[10] ,_u0_u16_ch_am0[9] , _u0_u16_ch_am0[8] , _u0_u16_ch_am0[7] ,_u0_u16_ch_am0[6] , _u0_u16_ch_am0[5] , _u0_u16_ch_am0[4] ,_u0_u16_ch_am0[3] , _u0_u16_ch_am0[2] , _u0_u16_ch_am0[1] ,_u0_u16_ch_am0[0] , _u0_u16_ch_am1[31] , _u0_u16_ch_am1[30] ,_u0_u16_ch_am1[29] , _u0_u16_ch_am1[28] , _u0_u16_ch_am1[27] ,_u0_u16_ch_am1[26] , _u0_u16_ch_am1[25] , _u0_u16_ch_am1[24] ,_u0_u16_ch_am1[23] , _u0_u16_ch_am1[22] , _u0_u16_ch_am1[21] ,_u0_u16_ch_am1[20] , _u0_u16_ch_am1[19] , _u0_u16_ch_am1[18] ,_u0_u16_ch_am1[17] , _u0_u16_ch_am1[16] , _u0_u16_ch_am1[15] ,_u0_u16_ch_am1[14] , _u0_u16_ch_am1[13] , _u0_u16_ch_am1[12] ,_u0_u16_ch_am1[11] , _u0_u16_ch_am1[10] , _u0_u16_ch_am1[9] ,_u0_u16_ch_am1[8] , _u0_u16_ch_am1[7] , _u0_u16_ch_am1[6] ,_u0_u16_ch_am1[5] , _u0_u16_ch_am1[4] , _u0_u16_ch_am1[3] ,_u0_u16_ch_am1[2] , _u0_u16_ch_am1[1] , _u0_u16_ch_am1[0] ,_u0_u16_sw_pointer[31] , _u0_u16_sw_pointer[30] ,_u0_u16_sw_pointer[29] , _u0_u16_sw_pointer[28] ,_u0_u16_sw_pointer[27] , _u0_u16_sw_pointer[26] ,_u0_u16_sw_pointer[25] , _u0_u16_sw_pointer[24] ,_u0_u16_sw_pointer[23] , _u0_u16_sw_pointer[22] ,_u0_u16_sw_pointer[21] , _u0_u16_sw_pointer[20] ,_u0_u16_sw_pointer[19] , _u0_u16_sw_pointer[18] ,_u0_u16_sw_pointer[17] , _u0_u16_sw_pointer[16] ,_u0_u16_sw_pointer[15] , _u0_u16_sw_pointer[14] ,_u0_u16_sw_pointer[13] , _u0_u16_sw_pointer[12] ,_u0_u16_sw_pointer[11] , _u0_u16_sw_pointer[10] ,_u0_u16_sw_pointer[9] , _u0_u16_sw_pointer[8] ,_u0_u16_sw_pointer[7] , _u0_u16_sw_pointer[6] ,_u0_u16_sw_pointer[5] , _u0_u16_sw_pointer[4] ,_u0_u16_sw_pointer[3] , _u0_u16_sw_pointer[2] ,_u0_u16_sw_pointer[1] , _u0_u16_sw_pointer[0] , _u0_u16_ch_stop ,_u0_u16_ch_dis , _u0_u16_int , _u0_u17_pointer[31] ,_u0_u17_pointer[30] , _u0_u17_pointer[29] , _u0_u17_pointer[28] ,_u0_u17_pointer[27] , _u0_u17_pointer[26] , _u0_u17_pointer[25] ,_u0_u17_pointer[24] , _u0_u17_pointer[23] , _u0_u17_pointer[22] ,_u0_u17_pointer[21] , _u0_u17_pointer[20] , _u0_u17_pointer[19] ,_u0_u17_pointer[18] , _u0_u17_pointer[17] , _u0_u17_pointer[16] ,_u0_u17_pointer[15] , _u0_u17_pointer[14] , _u0_u17_pointer[13] ,_u0_u17_pointer[12] , _u0_u17_pointer[11] , _u0_u17_pointer[10] ,_u0_u17_pointer[9] , _u0_u17_pointer[8] , _u0_u17_pointer[7] ,_u0_u17_pointer[6] , _u0_u17_pointer[5] , _u0_u17_pointer[4] ,_u0_u17_pointer[3] , _u0_u17_pointer[2] , _u0_u17_pointer[1] ,_u0_u17_pointer[0] , _u0_u17_pointer_s[31] , _u0_u17_pointer_s[30] ,_u0_u17_pointer_s[29] , _u0_u17_pointer_s[28] ,_u0_u17_pointer_s[27] , _u0_u17_pointer_s[26] ,_u0_u17_pointer_s[25] , _u0_u17_pointer_s[24] ,_u0_u17_pointer_s[23] , _u0_u17_pointer_s[22] ,_u0_u17_pointer_s[21] , _u0_u17_pointer_s[20] ,_u0_u17_pointer_s[19] , _u0_u17_pointer_s[18] ,_u0_u17_pointer_s[17] , _u0_u17_pointer_s[16] ,_u0_u17_pointer_s[15] , _u0_u17_pointer_s[14] ,_u0_u17_pointer_s[13] , _u0_u17_pointer_s[12] ,_u0_u17_pointer_s[11] , _u0_u17_pointer_s[10] , _u0_u17_pointer_s[9] ,_u0_u17_pointer_s[8] , _u0_u17_pointer_s[7] , _u0_u17_pointer_s[6] ,_u0_u17_pointer_s[5] , _u0_u17_pointer_s[4] , _u0_u17_pointer_s[3] ,_u0_u17_pointer_s[2] , _u0_u17_pointer_s[1] , _u0_u17_pointer_s[0] ,_u0_u17_ch_csr[31] , _u0_u17_ch_csr[30] , _u0_u17_ch_csr[29] ,_u0_u17_ch_csr[28] , _u0_u17_ch_csr[27] , _u0_u17_ch_csr[26] ,_u0_u17_ch_csr[25] , _u0_u17_ch_csr[24] , _u0_u17_ch_csr[23] ,_u0_u17_ch_csr[22] , _u0_u17_ch_csr[21] , _u0_u17_ch_csr[20] ,_u0_u17_ch_csr[19] , _u0_u17_ch_csr[18] , _u0_u17_ch_csr[17] ,_u0_u17_ch_csr[16] , _u0_u17_ch_csr[15] , _u0_u17_ch_csr[14] ,_u0_u17_ch_csr[13] , _u0_u17_ch_csr[12] , _u0_u17_ch_csr[11] ,_u0_u17_ch_csr[10] , _u0_u17_ch_csr[9] , _u0_u17_ch_csr[8] ,_u0_u17_ch_csr[7] , _u0_u17_ch_csr[6] , _u0_u17_ch_csr[5] ,_u0_u17_ch_csr[4] , _u0_u17_ch_csr[3] , _u0_u17_ch_csr[2] ,_u0_u17_ch_csr[1] , _u0_u17_ch_csr[0] , _u0_u17_ch_txsz[31] ,_u0_u17_ch_txsz[30] , _u0_u17_ch_txsz[29] , _u0_u17_ch_txsz[28] ,_u0_u17_ch_txsz[27] , _u0_u17_ch_txsz[26] , _u0_u17_ch_txsz[25] ,_u0_u17_ch_txsz[24] , _u0_u17_ch_txsz[23] , _u0_u17_ch_txsz[22] ,_u0_u17_ch_txsz[21] , _u0_u17_ch_txsz[20] , _u0_u17_ch_txsz[19] ,_u0_u17_ch_txsz[18] , _u0_u17_ch_txsz[17] , _u0_u17_ch_txsz[16] ,_u0_u17_ch_txsz[15] , _u0_u17_ch_txsz[14] , _u0_u17_ch_txsz[13] ,_u0_u17_ch_txsz[12] , _u0_u17_ch_txsz[11] , _u0_u17_ch_txsz[10] ,_u0_u17_ch_txsz[9] , _u0_u17_ch_txsz[8] , _u0_u17_ch_txsz[7] ,_u0_u17_ch_txsz[6] , _u0_u17_ch_txsz[5] , _u0_u17_ch_txsz[4] ,_u0_u17_ch_txsz[3] , _u0_u17_ch_txsz[2] , _u0_u17_ch_txsz[1] ,_u0_u17_ch_txsz[0] , _u0_u17_ch_adr0[31] , _u0_u17_ch_adr0[30] ,_u0_u17_ch_adr0[29] , _u0_u17_ch_adr0[28] , _u0_u17_ch_adr0[27] ,_u0_u17_ch_adr0[26] , _u0_u17_ch_adr0[25] , _u0_u17_ch_adr0[24] ,_u0_u17_ch_adr0[23] , _u0_u17_ch_adr0[22] , _u0_u17_ch_adr0[21] ,_u0_u17_ch_adr0[20] , _u0_u17_ch_adr0[19] , _u0_u17_ch_adr0[18] ,_u0_u17_ch_adr0[17] , _u0_u17_ch_adr0[16] , _u0_u17_ch_adr0[15] ,_u0_u17_ch_adr0[14] , _u0_u17_ch_adr0[13] , _u0_u17_ch_adr0[12] ,_u0_u17_ch_adr0[11] , _u0_u17_ch_adr0[10] , _u0_u17_ch_adr0[9] ,_u0_u17_ch_adr0[8] , _u0_u17_ch_adr0[7] , _u0_u17_ch_adr0[6] ,_u0_u17_ch_adr0[5] , _u0_u17_ch_adr0[4] , _u0_u17_ch_adr0[3] ,_u0_u17_ch_adr0[2] , _u0_u17_ch_adr0[1] , _u0_u17_ch_adr0[0] ,_u0_u17_ch_adr1[31] , _u0_u17_ch_adr1[30] , _u0_u17_ch_adr1[29] ,_u0_u17_ch_adr1[28] , _u0_u17_ch_adr1[27] , _u0_u17_ch_adr1[26] ,_u0_u17_ch_adr1[25] , _u0_u17_ch_adr1[24] , _u0_u17_ch_adr1[23] ,_u0_u17_ch_adr1[22] , _u0_u17_ch_adr1[21] , _u0_u17_ch_adr1[20] ,_u0_u17_ch_adr1[19] , _u0_u17_ch_adr1[18] , _u0_u17_ch_adr1[17] ,_u0_u17_ch_adr1[16] , _u0_u17_ch_adr1[15] , _u0_u17_ch_adr1[14] ,_u0_u17_ch_adr1[13] , _u0_u17_ch_adr1[12] , _u0_u17_ch_adr1[11] ,_u0_u17_ch_adr1[10] , _u0_u17_ch_adr1[9] , _u0_u17_ch_adr1[8] ,_u0_u17_ch_adr1[7] , _u0_u17_ch_adr1[6] , _u0_u17_ch_adr1[5] ,_u0_u17_ch_adr1[4] , _u0_u17_ch_adr1[3] , _u0_u17_ch_adr1[2] ,_u0_u17_ch_adr1[1] , _u0_u17_ch_adr1[0] , _u0_u17_ch_am0[31] ,_u0_u17_ch_am0[30] , _u0_u17_ch_am0[29] , _u0_u17_ch_am0[28] ,_u0_u17_ch_am0[27] , _u0_u17_ch_am0[26] , _u0_u17_ch_am0[25] ,_u0_u17_ch_am0[24] , _u0_u17_ch_am0[23] , _u0_u17_ch_am0[22] ,_u0_u17_ch_am0[21] , _u0_u17_ch_am0[20] , _u0_u17_ch_am0[19] ,_u0_u17_ch_am0[18] , _u0_u17_ch_am0[17] , _u0_u17_ch_am0[16] ,_u0_u17_ch_am0[15] , _u0_u17_ch_am0[14] , _u0_u17_ch_am0[13] ,_u0_u17_ch_am0[12] , _u0_u17_ch_am0[11] , _u0_u17_ch_am0[10] ,_u0_u17_ch_am0[9] , _u0_u17_ch_am0[8] , _u0_u17_ch_am0[7] ,_u0_u17_ch_am0[6] , _u0_u17_ch_am0[5] , _u0_u17_ch_am0[4] ,_u0_u17_ch_am0[3] , _u0_u17_ch_am0[2] , _u0_u17_ch_am0[1] ,_u0_u17_ch_am0[0] , _u0_u17_ch_am1[31] , _u0_u17_ch_am1[30] ,_u0_u17_ch_am1[29] , _u0_u17_ch_am1[28] , _u0_u17_ch_am1[27] ,_u0_u17_ch_am1[26] , _u0_u17_ch_am1[25] , _u0_u17_ch_am1[24] ,_u0_u17_ch_am1[23] , _u0_u17_ch_am1[22] , _u0_u17_ch_am1[21] ,_u0_u17_ch_am1[20] , _u0_u17_ch_am1[19] , _u0_u17_ch_am1[18] ,_u0_u17_ch_am1[17] , _u0_u17_ch_am1[16] , _u0_u17_ch_am1[15] ,_u0_u17_ch_am1[14] , _u0_u17_ch_am1[13] , _u0_u17_ch_am1[12] ,_u0_u17_ch_am1[11] , _u0_u17_ch_am1[10] , _u0_u17_ch_am1[9] ,_u0_u17_ch_am1[8] , _u0_u17_ch_am1[7] , _u0_u17_ch_am1[6] ,_u0_u17_ch_am1[5] , _u0_u17_ch_am1[4] , _u0_u17_ch_am1[3] ,_u0_u17_ch_am1[2] , _u0_u17_ch_am1[1] , _u0_u17_ch_am1[0] ,_u0_u17_sw_pointer[31] , _u0_u17_sw_pointer[30] ,_u0_u17_sw_pointer[29] , _u0_u17_sw_pointer[28] ,_u0_u17_sw_pointer[27] , _u0_u17_sw_pointer[26] ,_u0_u17_sw_pointer[25] , _u0_u17_sw_pointer[24] ,_u0_u17_sw_pointer[23] , _u0_u17_sw_pointer[22] ,_u0_u17_sw_pointer[21] , _u0_u17_sw_pointer[20] ,_u0_u17_sw_pointer[19] , _u0_u17_sw_pointer[18] ,_u0_u17_sw_pointer[17] , _u0_u17_sw_pointer[16] ,_u0_u17_sw_pointer[15] , _u0_u17_sw_pointer[14] ,_u0_u17_sw_pointer[13] , _u0_u17_sw_pointer[12] ,_u0_u17_sw_pointer[11] , _u0_u17_sw_pointer[10] ,_u0_u17_sw_pointer[9] , _u0_u17_sw_pointer[8] ,_u0_u17_sw_pointer[7] , _u0_u17_sw_pointer[6] ,_u0_u17_sw_pointer[5] , _u0_u17_sw_pointer[4] ,_u0_u17_sw_pointer[3] , _u0_u17_sw_pointer[2] ,_u0_u17_sw_pointer[1] , _u0_u17_sw_pointer[0] , _u0_u17_ch_stop ,_u0_u17_ch_dis , _u0_u17_int , _u0_u18_pointer[31] ,_u0_u18_pointer[30] , _u0_u18_pointer[29] , _u0_u18_pointer[28] ,_u0_u18_pointer[27] , _u0_u18_pointer[26] , _u0_u18_pointer[25] ,_u0_u18_pointer[24] , _u0_u18_pointer[23] , _u0_u18_pointer[22] ,_u0_u18_pointer[21] , _u0_u18_pointer[20] , _u0_u18_pointer[19] ,_u0_u18_pointer[18] , _u0_u18_pointer[17] , _u0_u18_pointer[16] ,_u0_u18_pointer[15] , _u0_u18_pointer[14] , _u0_u18_pointer[13] ,_u0_u18_pointer[12] , _u0_u18_pointer[11] , _u0_u18_pointer[10] ,_u0_u18_pointer[9] , _u0_u18_pointer[8] , _u0_u18_pointer[7] ,_u0_u18_pointer[6] , _u0_u18_pointer[5] , _u0_u18_pointer[4] ,_u0_u18_pointer[3] , _u0_u18_pointer[2] , _u0_u18_pointer[1] ,_u0_u18_pointer[0] , _u0_u18_pointer_s[31] , _u0_u18_pointer_s[30] ,_u0_u18_pointer_s[29] , _u0_u18_pointer_s[28] ,_u0_u18_pointer_s[27] , _u0_u18_pointer_s[26] ,_u0_u18_pointer_s[25] , _u0_u18_pointer_s[24] ,_u0_u18_pointer_s[23] , _u0_u18_pointer_s[22] ,_u0_u18_pointer_s[21] , _u0_u18_pointer_s[20] ,_u0_u18_pointer_s[19] , _u0_u18_pointer_s[18] ,_u0_u18_pointer_s[17] , _u0_u18_pointer_s[16] ,_u0_u18_pointer_s[15] , _u0_u18_pointer_s[14] ,_u0_u18_pointer_s[13] , _u0_u18_pointer_s[12] ,_u0_u18_pointer_s[11] , _u0_u18_pointer_s[10] , _u0_u18_pointer_s[9] ,_u0_u18_pointer_s[8] , _u0_u18_pointer_s[7] , _u0_u18_pointer_s[6] ,_u0_u18_pointer_s[5] , _u0_u18_pointer_s[4] , _u0_u18_pointer_s[3] ,_u0_u18_pointer_s[2] , _u0_u18_pointer_s[1] , _u0_u18_pointer_s[0] ,_u0_u18_ch_csr[31] , _u0_u18_ch_csr[30] , _u0_u18_ch_csr[29] ,_u0_u18_ch_csr[28] , _u0_u18_ch_csr[27] , _u0_u18_ch_csr[26] ,_u0_u18_ch_csr[25] , _u0_u18_ch_csr[24] , _u0_u18_ch_csr[23] ,_u0_u18_ch_csr[22] , _u0_u18_ch_csr[21] , _u0_u18_ch_csr[20] ,_u0_u18_ch_csr[19] , _u0_u18_ch_csr[18] , _u0_u18_ch_csr[17] ,_u0_u18_ch_csr[16] , _u0_u18_ch_csr[15] , _u0_u18_ch_csr[14] ,_u0_u18_ch_csr[13] , _u0_u18_ch_csr[12] , _u0_u18_ch_csr[11] ,_u0_u18_ch_csr[10] , _u0_u18_ch_csr[9] , _u0_u18_ch_csr[8] ,_u0_u18_ch_csr[7] , _u0_u18_ch_csr[6] , _u0_u18_ch_csr[5] ,_u0_u18_ch_csr[4] , _u0_u18_ch_csr[3] , _u0_u18_ch_csr[2] ,_u0_u18_ch_csr[1] , _u0_u18_ch_csr[0] , _u0_u18_ch_txsz[31] ,_u0_u18_ch_txsz[30] , _u0_u18_ch_txsz[29] , _u0_u18_ch_txsz[28] ,_u0_u18_ch_txsz[27] , _u0_u18_ch_txsz[26] , _u0_u18_ch_txsz[25] ,_u0_u18_ch_txsz[24] , _u0_u18_ch_txsz[23] , _u0_u18_ch_txsz[22] ,_u0_u18_ch_txsz[21] , _u0_u18_ch_txsz[20] , _u0_u18_ch_txsz[19] ,_u0_u18_ch_txsz[18] , _u0_u18_ch_txsz[17] , _u0_u18_ch_txsz[16] ,_u0_u18_ch_txsz[15] , _u0_u18_ch_txsz[14] , _u0_u18_ch_txsz[13] ,_u0_u18_ch_txsz[12] , _u0_u18_ch_txsz[11] , _u0_u18_ch_txsz[10] ,_u0_u18_ch_txsz[9] , _u0_u18_ch_txsz[8] , _u0_u18_ch_txsz[7] ,_u0_u18_ch_txsz[6] , _u0_u18_ch_txsz[5] , _u0_u18_ch_txsz[4] ,_u0_u18_ch_txsz[3] , _u0_u18_ch_txsz[2] , _u0_u18_ch_txsz[1] ,_u0_u18_ch_txsz[0] , _u0_u18_ch_adr0[31] , _u0_u18_ch_adr0[30] ,_u0_u18_ch_adr0[29] , _u0_u18_ch_adr0[28] , _u0_u18_ch_adr0[27] ,_u0_u18_ch_adr0[26] , _u0_u18_ch_adr0[25] , _u0_u18_ch_adr0[24] ,_u0_u18_ch_adr0[23] , _u0_u18_ch_adr0[22] , _u0_u18_ch_adr0[21] ,_u0_u18_ch_adr0[20] , _u0_u18_ch_adr0[19] , _u0_u18_ch_adr0[18] ,_u0_u18_ch_adr0[17] , _u0_u18_ch_adr0[16] , _u0_u18_ch_adr0[15] ,_u0_u18_ch_adr0[14] , _u0_u18_ch_adr0[13] , _u0_u18_ch_adr0[12] ,_u0_u18_ch_adr0[11] , _u0_u18_ch_adr0[10] , _u0_u18_ch_adr0[9] ,_u0_u18_ch_adr0[8] , _u0_u18_ch_adr0[7] , _u0_u18_ch_adr0[6] ,_u0_u18_ch_adr0[5] , _u0_u18_ch_adr0[4] , _u0_u18_ch_adr0[3] ,_u0_u18_ch_adr0[2] , _u0_u18_ch_adr0[1] , _u0_u18_ch_adr0[0] ,_u0_u18_ch_adr1[31] , _u0_u18_ch_adr1[30] , _u0_u18_ch_adr1[29] ,_u0_u18_ch_adr1[28] , _u0_u18_ch_adr1[27] , _u0_u18_ch_adr1[26] ,_u0_u18_ch_adr1[25] , _u0_u18_ch_adr1[24] , _u0_u18_ch_adr1[23] ,_u0_u18_ch_adr1[22] , _u0_u18_ch_adr1[21] , _u0_u18_ch_adr1[20] ,_u0_u18_ch_adr1[19] , _u0_u18_ch_adr1[18] , _u0_u18_ch_adr1[17] ,_u0_u18_ch_adr1[16] , _u0_u18_ch_adr1[15] , _u0_u18_ch_adr1[14] ,_u0_u18_ch_adr1[13] , _u0_u18_ch_adr1[12] , _u0_u18_ch_adr1[11] ,_u0_u18_ch_adr1[10] , _u0_u18_ch_adr1[9] , _u0_u18_ch_adr1[8] ,_u0_u18_ch_adr1[7] , _u0_u18_ch_adr1[6] , _u0_u18_ch_adr1[5] ,_u0_u18_ch_adr1[4] , _u0_u18_ch_adr1[3] , _u0_u18_ch_adr1[2] ,_u0_u18_ch_adr1[1] , _u0_u18_ch_adr1[0] , _u0_u18_ch_am0[31] ,_u0_u18_ch_am0[30] , _u0_u18_ch_am0[29] , _u0_u18_ch_am0[28] ,_u0_u18_ch_am0[27] , _u0_u18_ch_am0[26] , _u0_u18_ch_am0[25] ,_u0_u18_ch_am0[24] , _u0_u18_ch_am0[23] , _u0_u18_ch_am0[22] ,_u0_u18_ch_am0[21] , _u0_u18_ch_am0[20] , _u0_u18_ch_am0[19] ,_u0_u18_ch_am0[18] , _u0_u18_ch_am0[17] , _u0_u18_ch_am0[16] ,_u0_u18_ch_am0[15] , _u0_u18_ch_am0[14] , _u0_u18_ch_am0[13] ,_u0_u18_ch_am0[12] , _u0_u18_ch_am0[11] , _u0_u18_ch_am0[10] ,_u0_u18_ch_am0[9] , _u0_u18_ch_am0[8] , _u0_u18_ch_am0[7] ,_u0_u18_ch_am0[6] , _u0_u18_ch_am0[5] , _u0_u18_ch_am0[4] ,_u0_u18_ch_am0[3] , _u0_u18_ch_am0[2] , _u0_u18_ch_am0[1] ,_u0_u18_ch_am0[0] , _u0_u18_ch_am1[31] , _u0_u18_ch_am1[30] ,_u0_u18_ch_am1[29] , _u0_u18_ch_am1[28] , _u0_u18_ch_am1[27] ,_u0_u18_ch_am1[26] , _u0_u18_ch_am1[25] , _u0_u18_ch_am1[24] ,_u0_u18_ch_am1[23] , _u0_u18_ch_am1[22] , _u0_u18_ch_am1[21] ,_u0_u18_ch_am1[20] , _u0_u18_ch_am1[19] , _u0_u18_ch_am1[18] ,_u0_u18_ch_am1[17] , _u0_u18_ch_am1[16] , _u0_u18_ch_am1[15] ,_u0_u18_ch_am1[14] , _u0_u18_ch_am1[13] , _u0_u18_ch_am1[12] ,_u0_u18_ch_am1[11] , _u0_u18_ch_am1[10] , _u0_u18_ch_am1[9] ,_u0_u18_ch_am1[8] , _u0_u18_ch_am1[7] , _u0_u18_ch_am1[6] ,_u0_u18_ch_am1[5] , _u0_u18_ch_am1[4] , _u0_u18_ch_am1[3] ,_u0_u18_ch_am1[2] , _u0_u18_ch_am1[1] , _u0_u18_ch_am1[0] ,_u0_u18_sw_pointer[31] , _u0_u18_sw_pointer[30] ,_u0_u18_sw_pointer[29] , _u0_u18_sw_pointer[28] ,_u0_u18_sw_pointer[27] , _u0_u18_sw_pointer[26] ,_u0_u18_sw_pointer[25] , _u0_u18_sw_pointer[24] ,_u0_u18_sw_pointer[23] , _u0_u18_sw_pointer[22] ,_u0_u18_sw_pointer[21] , _u0_u18_sw_pointer[20] ,_u0_u18_sw_pointer[19] , _u0_u18_sw_pointer[18] ,_u0_u18_sw_pointer[17] , _u0_u18_sw_pointer[16] ,_u0_u18_sw_pointer[15] , _u0_u18_sw_pointer[14] ,_u0_u18_sw_pointer[13] , _u0_u18_sw_pointer[12] ,_u0_u18_sw_pointer[11] , _u0_u18_sw_pointer[10] ,_u0_u18_sw_pointer[9] , _u0_u18_sw_pointer[8] ,_u0_u18_sw_pointer[7] , _u0_u18_sw_pointer[6] ,_u0_u18_sw_pointer[5] , _u0_u18_sw_pointer[4] ,_u0_u18_sw_pointer[3] , _u0_u18_sw_pointer[2] ,_u0_u18_sw_pointer[1] , _u0_u18_sw_pointer[0] , _u0_u18_ch_stop ,_u0_u18_ch_dis , _u0_u18_int , _u0_u19_pointer[31] ,_u0_u19_pointer[30] , _u0_u19_pointer[29] , _u0_u19_pointer[28] ,_u0_u19_pointer[27] , _u0_u19_pointer[26] , _u0_u19_pointer[25] ,_u0_u19_pointer[24] , _u0_u19_pointer[23] , _u0_u19_pointer[22] ,_u0_u19_pointer[21] , _u0_u19_pointer[20] , _u0_u19_pointer[19] ,_u0_u19_pointer[18] , _u0_u19_pointer[17] , _u0_u19_pointer[16] ,_u0_u19_pointer[15] , _u0_u19_pointer[14] , _u0_u19_pointer[13] ,_u0_u19_pointer[12] , _u0_u19_pointer[11] , _u0_u19_pointer[10] ,_u0_u19_pointer[9] , _u0_u19_pointer[8] , _u0_u19_pointer[7] ,_u0_u19_pointer[6] , _u0_u19_pointer[5] , _u0_u19_pointer[4] ,_u0_u19_pointer[3] , _u0_u19_pointer[2] , _u0_u19_pointer[1] ,_u0_u19_pointer[0] , _u0_u19_pointer_s[31] , _u0_u19_pointer_s[30] ,_u0_u19_pointer_s[29] , _u0_u19_pointer_s[28] ,_u0_u19_pointer_s[27] , _u0_u19_pointer_s[26] ,_u0_u19_pointer_s[25] , _u0_u19_pointer_s[24] ,_u0_u19_pointer_s[23] , _u0_u19_pointer_s[22] ,_u0_u19_pointer_s[21] , _u0_u19_pointer_s[20] ,_u0_u19_pointer_s[19] , _u0_u19_pointer_s[18] ,_u0_u19_pointer_s[17] , _u0_u19_pointer_s[16] ,_u0_u19_pointer_s[15] , _u0_u19_pointer_s[14] ,_u0_u19_pointer_s[13] , _u0_u19_pointer_s[12] ,_u0_u19_pointer_s[11] , _u0_u19_pointer_s[10] , _u0_u19_pointer_s[9] ,_u0_u19_pointer_s[8] , _u0_u19_pointer_s[7] , _u0_u19_pointer_s[6] ,_u0_u19_pointer_s[5] , _u0_u19_pointer_s[4] , _u0_u19_pointer_s[3] ,_u0_u19_pointer_s[2] , _u0_u19_pointer_s[1] , _u0_u19_pointer_s[0] ,_u0_u19_ch_csr[31] , _u0_u19_ch_csr[30] , _u0_u19_ch_csr[29] ,_u0_u19_ch_csr[28] , _u0_u19_ch_csr[27] , _u0_u19_ch_csr[26] ,_u0_u19_ch_csr[25] , _u0_u19_ch_csr[24] , _u0_u19_ch_csr[23] ,_u0_u19_ch_csr[22] , _u0_u19_ch_csr[21] , _u0_u19_ch_csr[20] ,_u0_u19_ch_csr[19] , _u0_u19_ch_csr[18] , _u0_u19_ch_csr[17] ,_u0_u19_ch_csr[16] , _u0_u19_ch_csr[15] , _u0_u19_ch_csr[14] ,_u0_u19_ch_csr[13] , _u0_u19_ch_csr[12] , _u0_u19_ch_csr[11] ,_u0_u19_ch_csr[10] , _u0_u19_ch_csr[9] , _u0_u19_ch_csr[8] ,_u0_u19_ch_csr[7] , _u0_u19_ch_csr[6] , _u0_u19_ch_csr[5] ,_u0_u19_ch_csr[4] , _u0_u19_ch_csr[3] , _u0_u19_ch_csr[2] ,_u0_u19_ch_csr[1] , _u0_u19_ch_csr[0] , _u0_u19_ch_txsz[31] ,_u0_u19_ch_txsz[30] , _u0_u19_ch_txsz[29] , _u0_u19_ch_txsz[28] ,_u0_u19_ch_txsz[27] , _u0_u19_ch_txsz[26] , _u0_u19_ch_txsz[25] ,_u0_u19_ch_txsz[24] , _u0_u19_ch_txsz[23] , _u0_u19_ch_txsz[22] ,_u0_u19_ch_txsz[21] , _u0_u19_ch_txsz[20] , _u0_u19_ch_txsz[19] ,_u0_u19_ch_txsz[18] , _u0_u19_ch_txsz[17] , _u0_u19_ch_txsz[16] ,_u0_u19_ch_txsz[15] , _u0_u19_ch_txsz[14] , _u0_u19_ch_txsz[13] ,_u0_u19_ch_txsz[12] , _u0_u19_ch_txsz[11] , _u0_u19_ch_txsz[10] ,_u0_u19_ch_txsz[9] , _u0_u19_ch_txsz[8] , _u0_u19_ch_txsz[7] ,_u0_u19_ch_txsz[6] , _u0_u19_ch_txsz[5] , _u0_u19_ch_txsz[4] ,_u0_u19_ch_txsz[3] , _u0_u19_ch_txsz[2] , _u0_u19_ch_txsz[1] ,_u0_u19_ch_txsz[0] , _u0_u19_ch_adr0[31] , _u0_u19_ch_adr0[30] ,_u0_u19_ch_adr0[29] , _u0_u19_ch_adr0[28] , _u0_u19_ch_adr0[27] ,_u0_u19_ch_adr0[26] , _u0_u19_ch_adr0[25] , _u0_u19_ch_adr0[24] ,_u0_u19_ch_adr0[23] , _u0_u19_ch_adr0[22] , _u0_u19_ch_adr0[21] ,_u0_u19_ch_adr0[20] , _u0_u19_ch_adr0[19] , _u0_u19_ch_adr0[18] ,_u0_u19_ch_adr0[17] , _u0_u19_ch_adr0[16] , _u0_u19_ch_adr0[15] ,_u0_u19_ch_adr0[14] , _u0_u19_ch_adr0[13] , _u0_u19_ch_adr0[12] ,_u0_u19_ch_adr0[11] , _u0_u19_ch_adr0[10] , _u0_u19_ch_adr0[9] ,_u0_u19_ch_adr0[8] , _u0_u19_ch_adr0[7] , _u0_u19_ch_adr0[6] ,_u0_u19_ch_adr0[5] , _u0_u19_ch_adr0[4] , _u0_u19_ch_adr0[3] ,_u0_u19_ch_adr0[2] , _u0_u19_ch_adr0[1] , _u0_u19_ch_adr0[0] ,_u0_u19_ch_adr1[31] , _u0_u19_ch_adr1[30] , _u0_u19_ch_adr1[29] ,_u0_u19_ch_adr1[28] , _u0_u19_ch_adr1[27] , _u0_u19_ch_adr1[26] ,_u0_u19_ch_adr1[25] , _u0_u19_ch_adr1[24] , _u0_u19_ch_adr1[23] ,_u0_u19_ch_adr1[22] , _u0_u19_ch_adr1[21] , _u0_u19_ch_adr1[20] ,_u0_u19_ch_adr1[19] , _u0_u19_ch_adr1[18] , _u0_u19_ch_adr1[17] ,_u0_u19_ch_adr1[16] , _u0_u19_ch_adr1[15] , _u0_u19_ch_adr1[14] ,_u0_u19_ch_adr1[13] , _u0_u19_ch_adr1[12] , _u0_u19_ch_adr1[11] ,_u0_u19_ch_adr1[10] , _u0_u19_ch_adr1[9] , _u0_u19_ch_adr1[8] ,_u0_u19_ch_adr1[7] , _u0_u19_ch_adr1[6] , _u0_u19_ch_adr1[5] ,_u0_u19_ch_adr1[4] , _u0_u19_ch_adr1[3] , _u0_u19_ch_adr1[2] ,_u0_u19_ch_adr1[1] , _u0_u19_ch_adr1[0] , _u0_u19_ch_am0[31] ,_u0_u19_ch_am0[30] , _u0_u19_ch_am0[29] , _u0_u19_ch_am0[28] ,_u0_u19_ch_am0[27] , _u0_u19_ch_am0[26] , _u0_u19_ch_am0[25] ,_u0_u19_ch_am0[24] , _u0_u19_ch_am0[23] , _u0_u19_ch_am0[22] ,_u0_u19_ch_am0[21] , _u0_u19_ch_am0[20] , _u0_u19_ch_am0[19] ,_u0_u19_ch_am0[18] , _u0_u19_ch_am0[17] , _u0_u19_ch_am0[16] ,_u0_u19_ch_am0[15] , _u0_u19_ch_am0[14] , _u0_u19_ch_am0[13] ,_u0_u19_ch_am0[12] , _u0_u19_ch_am0[11] , _u0_u19_ch_am0[10] ,_u0_u19_ch_am0[9] , _u0_u19_ch_am0[8] , _u0_u19_ch_am0[7] ,_u0_u19_ch_am0[6] , _u0_u19_ch_am0[5] , _u0_u19_ch_am0[4] ,_u0_u19_ch_am0[3] , _u0_u19_ch_am0[2] , _u0_u19_ch_am0[1] ,_u0_u19_ch_am0[0] , _u0_u19_ch_am1[31] , _u0_u19_ch_am1[30] ,_u0_u19_ch_am1[29] , _u0_u19_ch_am1[28] , _u0_u19_ch_am1[27] ,_u0_u19_ch_am1[26] , _u0_u19_ch_am1[25] , _u0_u19_ch_am1[24] ,_u0_u19_ch_am1[23] , _u0_u19_ch_am1[22] , _u0_u19_ch_am1[21] ,_u0_u19_ch_am1[20] , _u0_u19_ch_am1[19] , _u0_u19_ch_am1[18] ,_u0_u19_ch_am1[17] , _u0_u19_ch_am1[16] , _u0_u19_ch_am1[15] ,_u0_u19_ch_am1[14] , _u0_u19_ch_am1[13] , _u0_u19_ch_am1[12] ,_u0_u19_ch_am1[11] , _u0_u19_ch_am1[10] , _u0_u19_ch_am1[9] ,_u0_u19_ch_am1[8] , _u0_u19_ch_am1[7] , _u0_u19_ch_am1[6] ,_u0_u19_ch_am1[5] , _u0_u19_ch_am1[4] , _u0_u19_ch_am1[3] ,_u0_u19_ch_am1[2] , _u0_u19_ch_am1[1] , _u0_u19_ch_am1[0] ,_u0_u19_sw_pointer[31] , _u0_u19_sw_pointer[30] ,_u0_u19_sw_pointer[29] , _u0_u19_sw_pointer[28] ,_u0_u19_sw_pointer[27] , _u0_u19_sw_pointer[26] ,_u0_u19_sw_pointer[25] , _u0_u19_sw_pointer[24] ,_u0_u19_sw_pointer[23] , _u0_u19_sw_pointer[22] ,_u0_u19_sw_pointer[21] , _u0_u19_sw_pointer[20] ,_u0_u19_sw_pointer[19] , _u0_u19_sw_pointer[18] ,_u0_u19_sw_pointer[17] , _u0_u19_sw_pointer[16] ,_u0_u19_sw_pointer[15] , _u0_u19_sw_pointer[14] ,_u0_u19_sw_pointer[13] , _u0_u19_sw_pointer[12] ,_u0_u19_sw_pointer[11] , _u0_u19_sw_pointer[10] ,_u0_u19_sw_pointer[9] , _u0_u19_sw_pointer[8] ,_u0_u19_sw_pointer[7] , _u0_u19_sw_pointer[6] ,_u0_u19_sw_pointer[5] , _u0_u19_sw_pointer[4] ,_u0_u19_sw_pointer[3] , _u0_u19_sw_pointer[2] ,_u0_u19_sw_pointer[1] , _u0_u19_sw_pointer[0] , _u0_u19_ch_stop ,_u0_u19_ch_dis , _u0_u19_int , _u0_u20_pointer[31] ,_u0_u20_pointer[30] , _u0_u20_pointer[29] , _u0_u20_pointer[28] ,_u0_u20_pointer[27] , _u0_u20_pointer[26] , _u0_u20_pointer[25] ,_u0_u20_pointer[24] , _u0_u20_pointer[23] , _u0_u20_pointer[22] ,_u0_u20_pointer[21] , _u0_u20_pointer[20] , _u0_u20_pointer[19] ,_u0_u20_pointer[18] , _u0_u20_pointer[17] , _u0_u20_pointer[16] ,_u0_u20_pointer[15] , _u0_u20_pointer[14] , _u0_u20_pointer[13] ,_u0_u20_pointer[12] , _u0_u20_pointer[11] , _u0_u20_pointer[10] ,_u0_u20_pointer[9] , _u0_u20_pointer[8] , _u0_u20_pointer[7] ,_u0_u20_pointer[6] , _u0_u20_pointer[5] , _u0_u20_pointer[4] ,_u0_u20_pointer[3] , _u0_u20_pointer[2] , _u0_u20_pointer[1] ,_u0_u20_pointer[0] , _u0_u20_pointer_s[31] , _u0_u20_pointer_s[30] ,_u0_u20_pointer_s[29] , _u0_u20_pointer_s[28] ,_u0_u20_pointer_s[27] , _u0_u20_pointer_s[26] ,_u0_u20_pointer_s[25] , _u0_u20_pointer_s[24] ,_u0_u20_pointer_s[23] , _u0_u20_pointer_s[22] ,_u0_u20_pointer_s[21] , _u0_u20_pointer_s[20] ,_u0_u20_pointer_s[19] , _u0_u20_pointer_s[18] ,_u0_u20_pointer_s[17] , _u0_u20_pointer_s[16] ,_u0_u20_pointer_s[15] , _u0_u20_pointer_s[14] ,_u0_u20_pointer_s[13] , _u0_u20_pointer_s[12] ,_u0_u20_pointer_s[11] , _u0_u20_pointer_s[10] , _u0_u20_pointer_s[9] ,_u0_u20_pointer_s[8] , _u0_u20_pointer_s[7] , _u0_u20_pointer_s[6] ,_u0_u20_pointer_s[5] , _u0_u20_pointer_s[4] , _u0_u20_pointer_s[3] ,_u0_u20_pointer_s[2] , _u0_u20_pointer_s[1] , _u0_u20_pointer_s[0] ,_u0_u20_ch_csr[31] , _u0_u20_ch_csr[30] , _u0_u20_ch_csr[29] ,_u0_u20_ch_csr[28] , _u0_u20_ch_csr[27] , _u0_u20_ch_csr[26] ,_u0_u20_ch_csr[25] , _u0_u20_ch_csr[24] , _u0_u20_ch_csr[23] ,_u0_u20_ch_csr[22] , _u0_u20_ch_csr[21] , _u0_u20_ch_csr[20] ,_u0_u20_ch_csr[19] , _u0_u20_ch_csr[18] , _u0_u20_ch_csr[17] ,_u0_u20_ch_csr[16] , _u0_u20_ch_csr[15] , _u0_u20_ch_csr[14] ,_u0_u20_ch_csr[13] , _u0_u20_ch_csr[12] , _u0_u20_ch_csr[11] ,_u0_u20_ch_csr[10] , _u0_u20_ch_csr[9] , _u0_u20_ch_csr[8] ,_u0_u20_ch_csr[7] , _u0_u20_ch_csr[6] , _u0_u20_ch_csr[5] ,_u0_u20_ch_csr[4] , _u0_u20_ch_csr[3] , _u0_u20_ch_csr[2] ,_u0_u20_ch_csr[1] , _u0_u20_ch_csr[0] , _u0_u20_ch_txsz[31] ,_u0_u20_ch_txsz[30] , _u0_u20_ch_txsz[29] , _u0_u20_ch_txsz[28] ,_u0_u20_ch_txsz[27] , _u0_u20_ch_txsz[26] , _u0_u20_ch_txsz[25] ,_u0_u20_ch_txsz[24] , _u0_u20_ch_txsz[23] , _u0_u20_ch_txsz[22] ,_u0_u20_ch_txsz[21] , _u0_u20_ch_txsz[20] , _u0_u20_ch_txsz[19] ,_u0_u20_ch_txsz[18] , _u0_u20_ch_txsz[17] , _u0_u20_ch_txsz[16] ,_u0_u20_ch_txsz[15] , _u0_u20_ch_txsz[14] , _u0_u20_ch_txsz[13] ,_u0_u20_ch_txsz[12] , _u0_u20_ch_txsz[11] , _u0_u20_ch_txsz[10] ,_u0_u20_ch_txsz[9] , _u0_u20_ch_txsz[8] , _u0_u20_ch_txsz[7] ,_u0_u20_ch_txsz[6] , _u0_u20_ch_txsz[5] , _u0_u20_ch_txsz[4] ,_u0_u20_ch_txsz[3] , _u0_u20_ch_txsz[2] , _u0_u20_ch_txsz[1] ,_u0_u20_ch_txsz[0] , _u0_u20_ch_adr0[31] , _u0_u20_ch_adr0[30] ,_u0_u20_ch_adr0[29] , _u0_u20_ch_adr0[28] , _u0_u20_ch_adr0[27] ,_u0_u20_ch_adr0[26] , _u0_u20_ch_adr0[25] , _u0_u20_ch_adr0[24] ,_u0_u20_ch_adr0[23] , _u0_u20_ch_adr0[22] , _u0_u20_ch_adr0[21] ,_u0_u20_ch_adr0[20] , _u0_u20_ch_adr0[19] , _u0_u20_ch_adr0[18] ,_u0_u20_ch_adr0[17] , _u0_u20_ch_adr0[16] , _u0_u20_ch_adr0[15] ,_u0_u20_ch_adr0[14] , _u0_u20_ch_adr0[13] , _u0_u20_ch_adr0[12] ,_u0_u20_ch_adr0[11] , _u0_u20_ch_adr0[10] , _u0_u20_ch_adr0[9] ,_u0_u20_ch_adr0[8] , _u0_u20_ch_adr0[7] , _u0_u20_ch_adr0[6] ,_u0_u20_ch_adr0[5] , _u0_u20_ch_adr0[4] , _u0_u20_ch_adr0[3] ,_u0_u20_ch_adr0[2] , _u0_u20_ch_adr0[1] , _u0_u20_ch_adr0[0] ,_u0_u20_ch_adr1[31] , _u0_u20_ch_adr1[30] , _u0_u20_ch_adr1[29] ,_u0_u20_ch_adr1[28] , _u0_u20_ch_adr1[27] , _u0_u20_ch_adr1[26] ,_u0_u20_ch_adr1[25] , _u0_u20_ch_adr1[24] , _u0_u20_ch_adr1[23] ,_u0_u20_ch_adr1[22] , _u0_u20_ch_adr1[21] , _u0_u20_ch_adr1[20] ,_u0_u20_ch_adr1[19] , _u0_u20_ch_adr1[18] , _u0_u20_ch_adr1[17] ,_u0_u20_ch_adr1[16] , _u0_u20_ch_adr1[15] , _u0_u20_ch_adr1[14] ,_u0_u20_ch_adr1[13] , _u0_u20_ch_adr1[12] , _u0_u20_ch_adr1[11] ,_u0_u20_ch_adr1[10] , _u0_u20_ch_adr1[9] , _u0_u20_ch_adr1[8] ,_u0_u20_ch_adr1[7] , _u0_u20_ch_adr1[6] , _u0_u20_ch_adr1[5] ,_u0_u20_ch_adr1[4] , _u0_u20_ch_adr1[3] , _u0_u20_ch_adr1[2] ,_u0_u20_ch_adr1[1] , _u0_u20_ch_adr1[0] , _u0_u20_ch_am0[31] ,_u0_u20_ch_am0[30] , _u0_u20_ch_am0[29] , _u0_u20_ch_am0[28] ,_u0_u20_ch_am0[27] , _u0_u20_ch_am0[26] , _u0_u20_ch_am0[25] ,_u0_u20_ch_am0[24] , _u0_u20_ch_am0[23] , _u0_u20_ch_am0[22] ,_u0_u20_ch_am0[21] , _u0_u20_ch_am0[20] , _u0_u20_ch_am0[19] ,_u0_u20_ch_am0[18] , _u0_u20_ch_am0[17] , _u0_u20_ch_am0[16] ,_u0_u20_ch_am0[15] , _u0_u20_ch_am0[14] , _u0_u20_ch_am0[13] ,_u0_u20_ch_am0[12] , _u0_u20_ch_am0[11] , _u0_u20_ch_am0[10] ,_u0_u20_ch_am0[9] , _u0_u20_ch_am0[8] , _u0_u20_ch_am0[7] ,_u0_u20_ch_am0[6] , _u0_u20_ch_am0[5] , _u0_u20_ch_am0[4] ,_u0_u20_ch_am0[3] , _u0_u20_ch_am0[2] , _u0_u20_ch_am0[1] ,_u0_u20_ch_am0[0] , _u0_u20_ch_am1[31] , _u0_u20_ch_am1[30] ,_u0_u20_ch_am1[29] , _u0_u20_ch_am1[28] , _u0_u20_ch_am1[27] ,_u0_u20_ch_am1[26] , _u0_u20_ch_am1[25] , _u0_u20_ch_am1[24] ,_u0_u20_ch_am1[23] , _u0_u20_ch_am1[22] , _u0_u20_ch_am1[21] ,_u0_u20_ch_am1[20] , _u0_u20_ch_am1[19] , _u0_u20_ch_am1[18] ,_u0_u20_ch_am1[17] , _u0_u20_ch_am1[16] , _u0_u20_ch_am1[15] ,_u0_u20_ch_am1[14] , _u0_u20_ch_am1[13] , _u0_u20_ch_am1[12] ,_u0_u20_ch_am1[11] , _u0_u20_ch_am1[10] , _u0_u20_ch_am1[9] ,_u0_u20_ch_am1[8] , _u0_u20_ch_am1[7] , _u0_u20_ch_am1[6] ,_u0_u20_ch_am1[5] , _u0_u20_ch_am1[4] , _u0_u20_ch_am1[3] ,_u0_u20_ch_am1[2] , _u0_u20_ch_am1[1] , _u0_u20_ch_am1[0] ,_u0_u20_sw_pointer[31] , _u0_u20_sw_pointer[30] ,_u0_u20_sw_pointer[29] , _u0_u20_sw_pointer[28] ,_u0_u20_sw_pointer[27] , _u0_u20_sw_pointer[26] ,_u0_u20_sw_pointer[25] , _u0_u20_sw_pointer[24] ,_u0_u20_sw_pointer[23] , _u0_u20_sw_pointer[22] ,_u0_u20_sw_pointer[21] , _u0_u20_sw_pointer[20] ,_u0_u20_sw_pointer[19] , _u0_u20_sw_pointer[18] ,_u0_u20_sw_pointer[17] , _u0_u20_sw_pointer[16] ,_u0_u20_sw_pointer[15] , _u0_u20_sw_pointer[14] ,_u0_u20_sw_pointer[13] , _u0_u20_sw_pointer[12] ,_u0_u20_sw_pointer[11] , _u0_u20_sw_pointer[10] ,_u0_u20_sw_pointer[9] , _u0_u20_sw_pointer[8] ,_u0_u20_sw_pointer[7] , _u0_u20_sw_pointer[6] ,_u0_u20_sw_pointer[5] , _u0_u20_sw_pointer[4] ,_u0_u20_sw_pointer[3] , _u0_u20_sw_pointer[2] ,_u0_u20_sw_pointer[1] , _u0_u20_sw_pointer[0] , _u0_u20_ch_stop ,_u0_u20_ch_dis , _u0_u20_int , _u0_u21_pointer[31] ,_u0_u21_pointer[30] , _u0_u21_pointer[29] , _u0_u21_pointer[28] ,_u0_u21_pointer[27] , _u0_u21_pointer[26] , _u0_u21_pointer[25] ,_u0_u21_pointer[24] , _u0_u21_pointer[23] , _u0_u21_pointer[22] ,_u0_u21_pointer[21] , _u0_u21_pointer[20] , _u0_u21_pointer[19] ,_u0_u21_pointer[18] , _u0_u21_pointer[17] , _u0_u21_pointer[16] ,_u0_u21_pointer[15] , _u0_u21_pointer[14] , _u0_u21_pointer[13] ,_u0_u21_pointer[12] , _u0_u21_pointer[11] , _u0_u21_pointer[10] ,_u0_u21_pointer[9] , _u0_u21_pointer[8] , _u0_u21_pointer[7] ,_u0_u21_pointer[6] , _u0_u21_pointer[5] , _u0_u21_pointer[4] ,_u0_u21_pointer[3] , _u0_u21_pointer[2] , _u0_u21_pointer[1] ,_u0_u21_pointer[0] , _u0_u21_pointer_s[31] , _u0_u21_pointer_s[30] ,_u0_u21_pointer_s[29] , _u0_u21_pointer_s[28] ,_u0_u21_pointer_s[27] , _u0_u21_pointer_s[26] ,_u0_u21_pointer_s[25] , _u0_u21_pointer_s[24] ,_u0_u21_pointer_s[23] , _u0_u21_pointer_s[22] ,_u0_u21_pointer_s[21] , _u0_u21_pointer_s[20] ,_u0_u21_pointer_s[19] , _u0_u21_pointer_s[18] ,_u0_u21_pointer_s[17] , _u0_u21_pointer_s[16] ,_u0_u21_pointer_s[15] , _u0_u21_pointer_s[14] ,_u0_u21_pointer_s[13] , _u0_u21_pointer_s[12] ,_u0_u21_pointer_s[11] , _u0_u21_pointer_s[10] , _u0_u21_pointer_s[9] ,_u0_u21_pointer_s[8] , _u0_u21_pointer_s[7] , _u0_u21_pointer_s[6] ,_u0_u21_pointer_s[5] , _u0_u21_pointer_s[4] , _u0_u21_pointer_s[3] ,_u0_u21_pointer_s[2] , _u0_u21_pointer_s[1] , _u0_u21_pointer_s[0] ,_u0_u21_ch_csr[31] , _u0_u21_ch_csr[30] , _u0_u21_ch_csr[29] ,_u0_u21_ch_csr[28] , _u0_u21_ch_csr[27] , _u0_u21_ch_csr[26] ,_u0_u21_ch_csr[25] , _u0_u21_ch_csr[24] , _u0_u21_ch_csr[23] ,_u0_u21_ch_csr[22] , _u0_u21_ch_csr[21] , _u0_u21_ch_csr[20] ,_u0_u21_ch_csr[19] , _u0_u21_ch_csr[18] , _u0_u21_ch_csr[17] ,_u0_u21_ch_csr[16] , _u0_u21_ch_csr[15] , _u0_u21_ch_csr[14] ,_u0_u21_ch_csr[13] , _u0_u21_ch_csr[12] , _u0_u21_ch_csr[11] ,_u0_u21_ch_csr[10] , _u0_u21_ch_csr[9] , _u0_u21_ch_csr[8] ,_u0_u21_ch_csr[7] , _u0_u21_ch_csr[6] , _u0_u21_ch_csr[5] ,_u0_u21_ch_csr[4] , _u0_u21_ch_csr[3] , _u0_u21_ch_csr[2] ,_u0_u21_ch_csr[1] , _u0_u21_ch_csr[0] , _u0_u21_ch_txsz[31] ,_u0_u21_ch_txsz[30] , _u0_u21_ch_txsz[29] , _u0_u21_ch_txsz[28] ,_u0_u21_ch_txsz[27] , _u0_u21_ch_txsz[26] , _u0_u21_ch_txsz[25] ,_u0_u21_ch_txsz[24] , _u0_u21_ch_txsz[23] , _u0_u21_ch_txsz[22] ,_u0_u21_ch_txsz[21] , _u0_u21_ch_txsz[20] , _u0_u21_ch_txsz[19] ,_u0_u21_ch_txsz[18] , _u0_u21_ch_txsz[17] , _u0_u21_ch_txsz[16] ,_u0_u21_ch_txsz[15] , _u0_u21_ch_txsz[14] , _u0_u21_ch_txsz[13] ,_u0_u21_ch_txsz[12] , _u0_u21_ch_txsz[11] , _u0_u21_ch_txsz[10] ,_u0_u21_ch_txsz[9] , _u0_u21_ch_txsz[8] , _u0_u21_ch_txsz[7] ,_u0_u21_ch_txsz[6] , _u0_u21_ch_txsz[5] , _u0_u21_ch_txsz[4] ,_u0_u21_ch_txsz[3] , _u0_u21_ch_txsz[2] , _u0_u21_ch_txsz[1] ,_u0_u21_ch_txsz[0] , _u0_u21_ch_adr0[31] , _u0_u21_ch_adr0[30] ,_u0_u21_ch_adr0[29] , _u0_u21_ch_adr0[28] , _u0_u21_ch_adr0[27] ,_u0_u21_ch_adr0[26] , _u0_u21_ch_adr0[25] , _u0_u21_ch_adr0[24] ,_u0_u21_ch_adr0[23] , _u0_u21_ch_adr0[22] , _u0_u21_ch_adr0[21] ,_u0_u21_ch_adr0[20] , _u0_u21_ch_adr0[19] , _u0_u21_ch_adr0[18] ,_u0_u21_ch_adr0[17] , _u0_u21_ch_adr0[16] , _u0_u21_ch_adr0[15] ,_u0_u21_ch_adr0[14] , _u0_u21_ch_adr0[13] , _u0_u21_ch_adr0[12] ,_u0_u21_ch_adr0[11] , _u0_u21_ch_adr0[10] , _u0_u21_ch_adr0[9] ,_u0_u21_ch_adr0[8] , _u0_u21_ch_adr0[7] , _u0_u21_ch_adr0[6] ,_u0_u21_ch_adr0[5] , _u0_u21_ch_adr0[4] , _u0_u21_ch_adr0[3] ,_u0_u21_ch_adr0[2] , _u0_u21_ch_adr0[1] , _u0_u21_ch_adr0[0] ,_u0_u21_ch_adr1[31] , _u0_u21_ch_adr1[30] , _u0_u21_ch_adr1[29] ,_u0_u21_ch_adr1[28] , _u0_u21_ch_adr1[27] , _u0_u21_ch_adr1[26] ,_u0_u21_ch_adr1[25] , _u0_u21_ch_adr1[24] , _u0_u21_ch_adr1[23] ,_u0_u21_ch_adr1[22] , _u0_u21_ch_adr1[21] , _u0_u21_ch_adr1[20] ,_u0_u21_ch_adr1[19] , _u0_u21_ch_adr1[18] , _u0_u21_ch_adr1[17] ,_u0_u21_ch_adr1[16] , _u0_u21_ch_adr1[15] , _u0_u21_ch_adr1[14] ,_u0_u21_ch_adr1[13] , _u0_u21_ch_adr1[12] , _u0_u21_ch_adr1[11] ,_u0_u21_ch_adr1[10] , _u0_u21_ch_adr1[9] , _u0_u21_ch_adr1[8] ,_u0_u21_ch_adr1[7] , _u0_u21_ch_adr1[6] , _u0_u21_ch_adr1[5] ,_u0_u21_ch_adr1[4] , _u0_u21_ch_adr1[3] , _u0_u21_ch_adr1[2] ,_u0_u21_ch_adr1[1] , _u0_u21_ch_adr1[0] , _u0_u21_ch_am0[31] ,_u0_u21_ch_am0[30] , _u0_u21_ch_am0[29] , _u0_u21_ch_am0[28] ,_u0_u21_ch_am0[27] , _u0_u21_ch_am0[26] , _u0_u21_ch_am0[25] ,_u0_u21_ch_am0[24] , _u0_u21_ch_am0[23] , _u0_u21_ch_am0[22] ,_u0_u21_ch_am0[21] , _u0_u21_ch_am0[20] , _u0_u21_ch_am0[19] ,_u0_u21_ch_am0[18] , _u0_u21_ch_am0[17] , _u0_u21_ch_am0[16] ,_u0_u21_ch_am0[15] , _u0_u21_ch_am0[14] , _u0_u21_ch_am0[13] ,_u0_u21_ch_am0[12] , _u0_u21_ch_am0[11] , _u0_u21_ch_am0[10] ,_u0_u21_ch_am0[9] , _u0_u21_ch_am0[8] , _u0_u21_ch_am0[7] ,_u0_u21_ch_am0[6] , _u0_u21_ch_am0[5] , _u0_u21_ch_am0[4] ,_u0_u21_ch_am0[3] , _u0_u21_ch_am0[2] , _u0_u21_ch_am0[1] ,_u0_u21_ch_am0[0] , _u0_u21_ch_am1[31] , _u0_u21_ch_am1[30] ,_u0_u21_ch_am1[29] , _u0_u21_ch_am1[28] , _u0_u21_ch_am1[27] ,_u0_u21_ch_am1[26] , _u0_u21_ch_am1[25] , _u0_u21_ch_am1[24] ,_u0_u21_ch_am1[23] , _u0_u21_ch_am1[22] , _u0_u21_ch_am1[21] ,_u0_u21_ch_am1[20] , _u0_u21_ch_am1[19] , _u0_u21_ch_am1[18] ,_u0_u21_ch_am1[17] , _u0_u21_ch_am1[16] , _u0_u21_ch_am1[15] ,_u0_u21_ch_am1[14] , _u0_u21_ch_am1[13] , _u0_u21_ch_am1[12] ,_u0_u21_ch_am1[11] , _u0_u21_ch_am1[10] , _u0_u21_ch_am1[9] ,_u0_u21_ch_am1[8] , _u0_u21_ch_am1[7] , _u0_u21_ch_am1[6] ,_u0_u21_ch_am1[5] , _u0_u21_ch_am1[4] , _u0_u21_ch_am1[3] ,_u0_u21_ch_am1[2] , _u0_u21_ch_am1[1] , _u0_u21_ch_am1[0] ,_u0_u21_sw_pointer[31] , _u0_u21_sw_pointer[30] ,_u0_u21_sw_pointer[29] , _u0_u21_sw_pointer[28] ,_u0_u21_sw_pointer[27] , _u0_u21_sw_pointer[26] ,_u0_u21_sw_pointer[25] , _u0_u21_sw_pointer[24] ,_u0_u21_sw_pointer[23] , _u0_u21_sw_pointer[22] ,_u0_u21_sw_pointer[21] , _u0_u21_sw_pointer[20] ,_u0_u21_sw_pointer[19] , _u0_u21_sw_pointer[18] ,_u0_u21_sw_pointer[17] , _u0_u21_sw_pointer[16] ,_u0_u21_sw_pointer[15] , _u0_u21_sw_pointer[14] ,_u0_u21_sw_pointer[13] , _u0_u21_sw_pointer[12] ,_u0_u21_sw_pointer[11] , _u0_u21_sw_pointer[10] ,_u0_u21_sw_pointer[9] , _u0_u21_sw_pointer[8] ,_u0_u21_sw_pointer[7] , _u0_u21_sw_pointer[6] ,_u0_u21_sw_pointer[5] , _u0_u21_sw_pointer[4] ,_u0_u21_sw_pointer[3] , _u0_u21_sw_pointer[2] ,_u0_u21_sw_pointer[1] , _u0_u21_sw_pointer[0] , _u0_u21_ch_stop ,_u0_u21_ch_dis , _u0_u21_int , _u0_u22_pointer[31] ,_u0_u22_pointer[30] , _u0_u22_pointer[29] , _u0_u22_pointer[28] ,_u0_u22_pointer[27] , _u0_u22_pointer[26] , _u0_u22_pointer[25] ,_u0_u22_pointer[24] , _u0_u22_pointer[23] , _u0_u22_pointer[22] ,_u0_u22_pointer[21] , _u0_u22_pointer[20] , _u0_u22_pointer[19] ,_u0_u22_pointer[18] , _u0_u22_pointer[17] , _u0_u22_pointer[16] ,_u0_u22_pointer[15] , _u0_u22_pointer[14] , _u0_u22_pointer[13] ,_u0_u22_pointer[12] , _u0_u22_pointer[11] , _u0_u22_pointer[10] ,_u0_u22_pointer[9] , _u0_u22_pointer[8] , _u0_u22_pointer[7] ,_u0_u22_pointer[6] , _u0_u22_pointer[5] , _u0_u22_pointer[4] ,_u0_u22_pointer[3] , _u0_u22_pointer[2] , _u0_u22_pointer[1] ,_u0_u22_pointer[0] , _u0_u22_pointer_s[31] , _u0_u22_pointer_s[30] ,_u0_u22_pointer_s[29] , _u0_u22_pointer_s[28] ,_u0_u22_pointer_s[27] , _u0_u22_pointer_s[26] ,_u0_u22_pointer_s[25] , _u0_u22_pointer_s[24] ,_u0_u22_pointer_s[23] , _u0_u22_pointer_s[22] ,_u0_u22_pointer_s[21] , _u0_u22_pointer_s[20] ,_u0_u22_pointer_s[19] , _u0_u22_pointer_s[18] ,_u0_u22_pointer_s[17] , _u0_u22_pointer_s[16] ,_u0_u22_pointer_s[15] , _u0_u22_pointer_s[14] ,_u0_u22_pointer_s[13] , _u0_u22_pointer_s[12] ,_u0_u22_pointer_s[11] , _u0_u22_pointer_s[10] , _u0_u22_pointer_s[9] ,_u0_u22_pointer_s[8] , _u0_u22_pointer_s[7] , _u0_u22_pointer_s[6] ,_u0_u22_pointer_s[5] , _u0_u22_pointer_s[4] , _u0_u22_pointer_s[3] ,_u0_u22_pointer_s[2] , _u0_u22_pointer_s[1] , _u0_u22_pointer_s[0] ,_u0_u22_ch_csr[31] , _u0_u22_ch_csr[30] , _u0_u22_ch_csr[29] ,_u0_u22_ch_csr[28] , _u0_u22_ch_csr[27] , _u0_u22_ch_csr[26] ,_u0_u22_ch_csr[25] , _u0_u22_ch_csr[24] , _u0_u22_ch_csr[23] ,_u0_u22_ch_csr[22] , _u0_u22_ch_csr[21] , _u0_u22_ch_csr[20] ,_u0_u22_ch_csr[19] , _u0_u22_ch_csr[18] , _u0_u22_ch_csr[17] ,_u0_u22_ch_csr[16] , _u0_u22_ch_csr[15] , _u0_u22_ch_csr[14] ,_u0_u22_ch_csr[13] , _u0_u22_ch_csr[12] , _u0_u22_ch_csr[11] ,_u0_u22_ch_csr[10] , _u0_u22_ch_csr[9] , _u0_u22_ch_csr[8] ,_u0_u22_ch_csr[7] , _u0_u22_ch_csr[6] , _u0_u22_ch_csr[5] ,_u0_u22_ch_csr[4] , _u0_u22_ch_csr[3] , _u0_u22_ch_csr[2] ,_u0_u22_ch_csr[1] , _u0_u22_ch_csr[0] , _u0_u22_ch_txsz[31] ,_u0_u22_ch_txsz[30] , _u0_u22_ch_txsz[29] , _u0_u22_ch_txsz[28] ,_u0_u22_ch_txsz[27] , _u0_u22_ch_txsz[26] , _u0_u22_ch_txsz[25] ,_u0_u22_ch_txsz[24] , _u0_u22_ch_txsz[23] , _u0_u22_ch_txsz[22] ,_u0_u22_ch_txsz[21] , _u0_u22_ch_txsz[20] , _u0_u22_ch_txsz[19] ,_u0_u22_ch_txsz[18] , _u0_u22_ch_txsz[17] , _u0_u22_ch_txsz[16] ,_u0_u22_ch_txsz[15] , _u0_u22_ch_txsz[14] , _u0_u22_ch_txsz[13] ,_u0_u22_ch_txsz[12] , _u0_u22_ch_txsz[11] , _u0_u22_ch_txsz[10] ,_u0_u22_ch_txsz[9] , _u0_u22_ch_txsz[8] , _u0_u22_ch_txsz[7] ,_u0_u22_ch_txsz[6] , _u0_u22_ch_txsz[5] , _u0_u22_ch_txsz[4] ,_u0_u22_ch_txsz[3] , _u0_u22_ch_txsz[2] , _u0_u22_ch_txsz[1] ,_u0_u22_ch_txsz[0] , _u0_u22_ch_adr0[31] , _u0_u22_ch_adr0[30] ,_u0_u22_ch_adr0[29] , _u0_u22_ch_adr0[28] , _u0_u22_ch_adr0[27] ,_u0_u22_ch_adr0[26] , _u0_u22_ch_adr0[25] , _u0_u22_ch_adr0[24] ,_u0_u22_ch_adr0[23] , _u0_u22_ch_adr0[22] , _u0_u22_ch_adr0[21] ,_u0_u22_ch_adr0[20] , _u0_u22_ch_adr0[19] , _u0_u22_ch_adr0[18] ,_u0_u22_ch_adr0[17] , _u0_u22_ch_adr0[16] , _u0_u22_ch_adr0[15] ,_u0_u22_ch_adr0[14] , _u0_u22_ch_adr0[13] , _u0_u22_ch_adr0[12] ,_u0_u22_ch_adr0[11] , _u0_u22_ch_adr0[10] , _u0_u22_ch_adr0[9] ,_u0_u22_ch_adr0[8] , _u0_u22_ch_adr0[7] , _u0_u22_ch_adr0[6] ,_u0_u22_ch_adr0[5] , _u0_u22_ch_adr0[4] , _u0_u22_ch_adr0[3] ,_u0_u22_ch_adr0[2] , _u0_u22_ch_adr0[1] , _u0_u22_ch_adr0[0] ,_u0_u22_ch_adr1[31] , _u0_u22_ch_adr1[30] , _u0_u22_ch_adr1[29] ,_u0_u22_ch_adr1[28] , _u0_u22_ch_adr1[27] , _u0_u22_ch_adr1[26] ,_u0_u22_ch_adr1[25] , _u0_u22_ch_adr1[24] , _u0_u22_ch_adr1[23] ,_u0_u22_ch_adr1[22] , _u0_u22_ch_adr1[21] , _u0_u22_ch_adr1[20] ,_u0_u22_ch_adr1[19] , _u0_u22_ch_adr1[18] , _u0_u22_ch_adr1[17] ,_u0_u22_ch_adr1[16] , _u0_u22_ch_adr1[15] , _u0_u22_ch_adr1[14] ,_u0_u22_ch_adr1[13] , _u0_u22_ch_adr1[12] , _u0_u22_ch_adr1[11] ,_u0_u22_ch_adr1[10] , _u0_u22_ch_adr1[9] , _u0_u22_ch_adr1[8] ,_u0_u22_ch_adr1[7] , _u0_u22_ch_adr1[6] , _u0_u22_ch_adr1[5] ,_u0_u22_ch_adr1[4] , _u0_u22_ch_adr1[3] , _u0_u22_ch_adr1[2] ,_u0_u22_ch_adr1[1] , _u0_u22_ch_adr1[0] , _u0_u22_ch_am0[31] ,_u0_u22_ch_am0[30] , _u0_u22_ch_am0[29] , _u0_u22_ch_am0[28] ,_u0_u22_ch_am0[27] , _u0_u22_ch_am0[26] , _u0_u22_ch_am0[25] ,_u0_u22_ch_am0[24] , _u0_u22_ch_am0[23] , _u0_u22_ch_am0[22] ,_u0_u22_ch_am0[21] , _u0_u22_ch_am0[20] , _u0_u22_ch_am0[19] ,_u0_u22_ch_am0[18] , _u0_u22_ch_am0[17] , _u0_u22_ch_am0[16] ,_u0_u22_ch_am0[15] , _u0_u22_ch_am0[14] , _u0_u22_ch_am0[13] ,_u0_u22_ch_am0[12] , _u0_u22_ch_am0[11] , _u0_u22_ch_am0[10] ,_u0_u22_ch_am0[9] , _u0_u22_ch_am0[8] , _u0_u22_ch_am0[7] ,_u0_u22_ch_am0[6] , _u0_u22_ch_am0[5] , _u0_u22_ch_am0[4] ,_u0_u22_ch_am0[3] , _u0_u22_ch_am0[2] , _u0_u22_ch_am0[1] ,_u0_u22_ch_am0[0] , _u0_u22_ch_am1[31] , _u0_u22_ch_am1[30] ,_u0_u22_ch_am1[29] , _u0_u22_ch_am1[28] , _u0_u22_ch_am1[27] ,_u0_u22_ch_am1[26] , _u0_u22_ch_am1[25] , _u0_u22_ch_am1[24] ,_u0_u22_ch_am1[23] , _u0_u22_ch_am1[22] , _u0_u22_ch_am1[21] ,_u0_u22_ch_am1[20] , _u0_u22_ch_am1[19] , _u0_u22_ch_am1[18] ,_u0_u22_ch_am1[17] , _u0_u22_ch_am1[16] , _u0_u22_ch_am1[15] ,_u0_u22_ch_am1[14] , _u0_u22_ch_am1[13] , _u0_u22_ch_am1[12] ,_u0_u22_ch_am1[11] , _u0_u22_ch_am1[10] , _u0_u22_ch_am1[9] ,_u0_u22_ch_am1[8] , _u0_u22_ch_am1[7] , _u0_u22_ch_am1[6] ,_u0_u22_ch_am1[5] , _u0_u22_ch_am1[4] , _u0_u22_ch_am1[3] ,_u0_u22_ch_am1[2] , _u0_u22_ch_am1[1] , _u0_u22_ch_am1[0] ,_u0_u22_sw_pointer[31] , _u0_u22_sw_pointer[30] ,_u0_u22_sw_pointer[29] , _u0_u22_sw_pointer[28] ,_u0_u22_sw_pointer[27] , _u0_u22_sw_pointer[26] ,_u0_u22_sw_pointer[25] , _u0_u22_sw_pointer[24] ,_u0_u22_sw_pointer[23] , _u0_u22_sw_pointer[22] ,_u0_u22_sw_pointer[21] , _u0_u22_sw_pointer[20] ,_u0_u22_sw_pointer[19] , _u0_u22_sw_pointer[18] ,_u0_u22_sw_pointer[17] , _u0_u22_sw_pointer[16] ,_u0_u22_sw_pointer[15] , _u0_u22_sw_pointer[14] ,_u0_u22_sw_pointer[13] , _u0_u22_sw_pointer[12] ,_u0_u22_sw_pointer[11] , _u0_u22_sw_pointer[10] ,_u0_u22_sw_pointer[9] , _u0_u22_sw_pointer[8] ,_u0_u22_sw_pointer[7] , _u0_u22_sw_pointer[6] ,_u0_u22_sw_pointer[5] , _u0_u22_sw_pointer[4] ,_u0_u22_sw_pointer[3] , _u0_u22_sw_pointer[2] ,_u0_u22_sw_pointer[1] , _u0_u22_sw_pointer[0] , _u0_u22_ch_stop ,_u0_u22_ch_dis , _u0_u22_int , _u0_u23_pointer[31] ,_u0_u23_pointer[30] , _u0_u23_pointer[29] , _u0_u23_pointer[28] ,_u0_u23_pointer[27] , _u0_u23_pointer[26] , _u0_u23_pointer[25] ,_u0_u23_pointer[24] , _u0_u23_pointer[23] , _u0_u23_pointer[22] ,_u0_u23_pointer[21] , _u0_u23_pointer[20] , _u0_u23_pointer[19] ,_u0_u23_pointer[18] , _u0_u23_pointer[17] , _u0_u23_pointer[16] ,_u0_u23_pointer[15] , _u0_u23_pointer[14] , _u0_u23_pointer[13] ,_u0_u23_pointer[12] , _u0_u23_pointer[11] , _u0_u23_pointer[10] ,_u0_u23_pointer[9] , _u0_u23_pointer[8] , _u0_u23_pointer[7] ,_u0_u23_pointer[6] , _u0_u23_pointer[5] , _u0_u23_pointer[4] ,_u0_u23_pointer[3] , _u0_u23_pointer[2] , _u0_u23_pointer[1] ,_u0_u23_pointer[0] , _u0_u23_pointer_s[31] , _u0_u23_pointer_s[30] ,_u0_u23_pointer_s[29] , _u0_u23_pointer_s[28] ,_u0_u23_pointer_s[27] , _u0_u23_pointer_s[26] ,_u0_u23_pointer_s[25] , _u0_u23_pointer_s[24] ,_u0_u23_pointer_s[23] , _u0_u23_pointer_s[22] ,_u0_u23_pointer_s[21] , _u0_u23_pointer_s[20] ,_u0_u23_pointer_s[19] , _u0_u23_pointer_s[18] ,_u0_u23_pointer_s[17] , _u0_u23_pointer_s[16] ,_u0_u23_pointer_s[15] , _u0_u23_pointer_s[14] ,_u0_u23_pointer_s[13] , _u0_u23_pointer_s[12] ,_u0_u23_pointer_s[11] , _u0_u23_pointer_s[10] , _u0_u23_pointer_s[9] ,_u0_u23_pointer_s[8] , _u0_u23_pointer_s[7] , _u0_u23_pointer_s[6] ,_u0_u23_pointer_s[5] , _u0_u23_pointer_s[4] , _u0_u23_pointer_s[3] ,_u0_u23_pointer_s[2] , _u0_u23_pointer_s[1] , _u0_u23_pointer_s[0] ,_u0_u23_ch_csr[31] , _u0_u23_ch_csr[30] , _u0_u23_ch_csr[29] ,_u0_u23_ch_csr[28] , _u0_u23_ch_csr[27] , _u0_u23_ch_csr[26] ,_u0_u23_ch_csr[25] , _u0_u23_ch_csr[24] , _u0_u23_ch_csr[23] ,_u0_u23_ch_csr[22] , _u0_u23_ch_csr[21] , _u0_u23_ch_csr[20] ,_u0_u23_ch_csr[19] , _u0_u23_ch_csr[18] , _u0_u23_ch_csr[17] ,_u0_u23_ch_csr[16] , _u0_u23_ch_csr[15] , _u0_u23_ch_csr[14] ,_u0_u23_ch_csr[13] , _u0_u23_ch_csr[12] , _u0_u23_ch_csr[11] ,_u0_u23_ch_csr[10] , _u0_u23_ch_csr[9] , _u0_u23_ch_csr[8] ,_u0_u23_ch_csr[7] , _u0_u23_ch_csr[6] , _u0_u23_ch_csr[5] ,_u0_u23_ch_csr[4] , _u0_u23_ch_csr[3] , _u0_u23_ch_csr[2] ,_u0_u23_ch_csr[1] , _u0_u23_ch_csr[0] , _u0_u23_ch_txsz[31] ,_u0_u23_ch_txsz[30] , _u0_u23_ch_txsz[29] , _u0_u23_ch_txsz[28] ,_u0_u23_ch_txsz[27] , _u0_u23_ch_txsz[26] , _u0_u23_ch_txsz[25] ,_u0_u23_ch_txsz[24] , _u0_u23_ch_txsz[23] , _u0_u23_ch_txsz[22] ,_u0_u23_ch_txsz[21] , _u0_u23_ch_txsz[20] , _u0_u23_ch_txsz[19] ,_u0_u23_ch_txsz[18] , _u0_u23_ch_txsz[17] , _u0_u23_ch_txsz[16] ,_u0_u23_ch_txsz[15] , _u0_u23_ch_txsz[14] , _u0_u23_ch_txsz[13] ,_u0_u23_ch_txsz[12] , _u0_u23_ch_txsz[11] , _u0_u23_ch_txsz[10] ,_u0_u23_ch_txsz[9] , _u0_u23_ch_txsz[8] , _u0_u23_ch_txsz[7] ,_u0_u23_ch_txsz[6] , _u0_u23_ch_txsz[5] , _u0_u23_ch_txsz[4] ,_u0_u23_ch_txsz[3] , _u0_u23_ch_txsz[2] , _u0_u23_ch_txsz[1] ,_u0_u23_ch_txsz[0] , _u0_u23_ch_adr0[31] , _u0_u23_ch_adr0[30] ,_u0_u23_ch_adr0[29] , _u0_u23_ch_adr0[28] , _u0_u23_ch_adr0[27] ,_u0_u23_ch_adr0[26] , _u0_u23_ch_adr0[25] , _u0_u23_ch_adr0[24] ,_u0_u23_ch_adr0[23] , _u0_u23_ch_adr0[22] , _u0_u23_ch_adr0[21] ,_u0_u23_ch_adr0[20] , _u0_u23_ch_adr0[19] , _u0_u23_ch_adr0[18] ,_u0_u23_ch_adr0[17] , _u0_u23_ch_adr0[16] , _u0_u23_ch_adr0[15] ,_u0_u23_ch_adr0[14] , _u0_u23_ch_adr0[13] , _u0_u23_ch_adr0[12] ,_u0_u23_ch_adr0[11] , _u0_u23_ch_adr0[10] , _u0_u23_ch_adr0[9] ,_u0_u23_ch_adr0[8] , _u0_u23_ch_adr0[7] , _u0_u23_ch_adr0[6] ,_u0_u23_ch_adr0[5] , _u0_u23_ch_adr0[4] , _u0_u23_ch_adr0[3] ,_u0_u23_ch_adr0[2] , _u0_u23_ch_adr0[1] , _u0_u23_ch_adr0[0] ,_u0_u23_ch_adr1[31] , _u0_u23_ch_adr1[30] , _u0_u23_ch_adr1[29] ,_u0_u23_ch_adr1[28] , _u0_u23_ch_adr1[27] , _u0_u23_ch_adr1[26] ,_u0_u23_ch_adr1[25] , _u0_u23_ch_adr1[24] , _u0_u23_ch_adr1[23] ,_u0_u23_ch_adr1[22] , _u0_u23_ch_adr1[21] , _u0_u23_ch_adr1[20] ,_u0_u23_ch_adr1[19] , _u0_u23_ch_adr1[18] , _u0_u23_ch_adr1[17] ,_u0_u23_ch_adr1[16] , _u0_u23_ch_adr1[15] , _u0_u23_ch_adr1[14] ,_u0_u23_ch_adr1[13] , _u0_u23_ch_adr1[12] , _u0_u23_ch_adr1[11] ,_u0_u23_ch_adr1[10] , _u0_u23_ch_adr1[9] , _u0_u23_ch_adr1[8] ,_u0_u23_ch_adr1[7] , _u0_u23_ch_adr1[6] , _u0_u23_ch_adr1[5] ,_u0_u23_ch_adr1[4] , _u0_u23_ch_adr1[3] , _u0_u23_ch_adr1[2] ,_u0_u23_ch_adr1[1] , _u0_u23_ch_adr1[0] , _u0_u23_ch_am0[31] ,_u0_u23_ch_am0[30] , _u0_u23_ch_am0[29] , _u0_u23_ch_am0[28] ,_u0_u23_ch_am0[27] , _u0_u23_ch_am0[26] , _u0_u23_ch_am0[25] ,_u0_u23_ch_am0[24] , _u0_u23_ch_am0[23] , _u0_u23_ch_am0[22] ,_u0_u23_ch_am0[21] , _u0_u23_ch_am0[20] , _u0_u23_ch_am0[19] ,_u0_u23_ch_am0[18] , _u0_u23_ch_am0[17] , _u0_u23_ch_am0[16] ,_u0_u23_ch_am0[15] , _u0_u23_ch_am0[14] , _u0_u23_ch_am0[13] ,_u0_u23_ch_am0[12] , _u0_u23_ch_am0[11] , _u0_u23_ch_am0[10] ,_u0_u23_ch_am0[9] , _u0_u23_ch_am0[8] , _u0_u23_ch_am0[7] ,_u0_u23_ch_am0[6] , _u0_u23_ch_am0[5] , _u0_u23_ch_am0[4] ,_u0_u23_ch_am0[3] , _u0_u23_ch_am0[2] , _u0_u23_ch_am0[1] ,_u0_u23_ch_am0[0] , _u0_u23_ch_am1[31] , _u0_u23_ch_am1[30] ,_u0_u23_ch_am1[29] , _u0_u23_ch_am1[28] , _u0_u23_ch_am1[27] ,_u0_u23_ch_am1[26] , _u0_u23_ch_am1[25] , _u0_u23_ch_am1[24] ,_u0_u23_ch_am1[23] , _u0_u23_ch_am1[22] , _u0_u23_ch_am1[21] ,_u0_u23_ch_am1[20] , _u0_u23_ch_am1[19] , _u0_u23_ch_am1[18] ,_u0_u23_ch_am1[17] , _u0_u23_ch_am1[16] , _u0_u23_ch_am1[15] ,_u0_u23_ch_am1[14] , _u0_u23_ch_am1[13] , _u0_u23_ch_am1[12] ,_u0_u23_ch_am1[11] , _u0_u23_ch_am1[10] , _u0_u23_ch_am1[9] ,_u0_u23_ch_am1[8] , _u0_u23_ch_am1[7] , _u0_u23_ch_am1[6] ,_u0_u23_ch_am1[5] , _u0_u23_ch_am1[4] , _u0_u23_ch_am1[3] ,_u0_u23_ch_am1[2] , _u0_u23_ch_am1[1] , _u0_u23_ch_am1[0] ,_u0_u23_sw_pointer[31] , _u0_u23_sw_pointer[30] ,_u0_u23_sw_pointer[29] , _u0_u23_sw_pointer[28] ,_u0_u23_sw_pointer[27] , _u0_u23_sw_pointer[26] ,_u0_u23_sw_pointer[25] , _u0_u23_sw_pointer[24] ,_u0_u23_sw_pointer[23] , _u0_u23_sw_pointer[22] ,_u0_u23_sw_pointer[21] , _u0_u23_sw_pointer[20] ,_u0_u23_sw_pointer[19] , _u0_u23_sw_pointer[18] ,_u0_u23_sw_pointer[17] , _u0_u23_sw_pointer[16] ,_u0_u23_sw_pointer[15] , _u0_u23_sw_pointer[14] ,_u0_u23_sw_pointer[13] , _u0_u23_sw_pointer[12] ,_u0_u23_sw_pointer[11] , _u0_u23_sw_pointer[10] ,_u0_u23_sw_pointer[9] , _u0_u23_sw_pointer[8] ,_u0_u23_sw_pointer[7] , _u0_u23_sw_pointer[6] ,_u0_u23_sw_pointer[5] , _u0_u23_sw_pointer[4] ,_u0_u23_sw_pointer[3] , _u0_u23_sw_pointer[2] ,_u0_u23_sw_pointer[1] , _u0_u23_sw_pointer[0] , _u0_u23_ch_stop ,_u0_u23_ch_dis , _u0_u23_int , _u0_u24_pointer[31] ,_u0_u24_pointer[30] , _u0_u24_pointer[29] , _u0_u24_pointer[28] ,_u0_u24_pointer[27] , _u0_u24_pointer[26] , _u0_u24_pointer[25] ,_u0_u24_pointer[24] , _u0_u24_pointer[23] , _u0_u24_pointer[22] ,_u0_u24_pointer[21] , _u0_u24_pointer[20] , _u0_u24_pointer[19] ,_u0_u24_pointer[18] , _u0_u24_pointer[17] , _u0_u24_pointer[16] ,_u0_u24_pointer[15] , _u0_u24_pointer[14] , _u0_u24_pointer[13] ,_u0_u24_pointer[12] , _u0_u24_pointer[11] , _u0_u24_pointer[10] ,_u0_u24_pointer[9] , _u0_u24_pointer[8] , _u0_u24_pointer[7] ,_u0_u24_pointer[6] , _u0_u24_pointer[5] , _u0_u24_pointer[4] ,_u0_u24_pointer[3] , _u0_u24_pointer[2] , _u0_u24_pointer[1] ,_u0_u24_pointer[0] , _u0_u24_pointer_s[31] , _u0_u24_pointer_s[30] ,_u0_u24_pointer_s[29] , _u0_u24_pointer_s[28] ,_u0_u24_pointer_s[27] , _u0_u24_pointer_s[26] ,_u0_u24_pointer_s[25] , _u0_u24_pointer_s[24] ,_u0_u24_pointer_s[23] , _u0_u24_pointer_s[22] ,_u0_u24_pointer_s[21] , _u0_u24_pointer_s[20] ,_u0_u24_pointer_s[19] , _u0_u24_pointer_s[18] ,_u0_u24_pointer_s[17] , _u0_u24_pointer_s[16] ,_u0_u24_pointer_s[15] , _u0_u24_pointer_s[14] ,_u0_u24_pointer_s[13] , _u0_u24_pointer_s[12] ,_u0_u24_pointer_s[11] , _u0_u24_pointer_s[10] , _u0_u24_pointer_s[9] ,_u0_u24_pointer_s[8] , _u0_u24_pointer_s[7] , _u0_u24_pointer_s[6] ,_u0_u24_pointer_s[5] , _u0_u24_pointer_s[4] , _u0_u24_pointer_s[3] ,_u0_u24_pointer_s[2] , _u0_u24_pointer_s[1] , _u0_u24_pointer_s[0] ,_u0_u24_ch_csr[31] , _u0_u24_ch_csr[30] , _u0_u24_ch_csr[29] ,_u0_u24_ch_csr[28] , _u0_u24_ch_csr[27] , _u0_u24_ch_csr[26] ,_u0_u24_ch_csr[25] , _u0_u24_ch_csr[24] , _u0_u24_ch_csr[23] ,_u0_u24_ch_csr[22] , _u0_u24_ch_csr[21] , _u0_u24_ch_csr[20] ,_u0_u24_ch_csr[19] , _u0_u24_ch_csr[18] , _u0_u24_ch_csr[17] ,_u0_u24_ch_csr[16] , _u0_u24_ch_csr[15] , _u0_u24_ch_csr[14] ,_u0_u24_ch_csr[13] , _u0_u24_ch_csr[12] , _u0_u24_ch_csr[11] ,_u0_u24_ch_csr[10] , _u0_u24_ch_csr[9] , _u0_u24_ch_csr[8] ,_u0_u24_ch_csr[7] , _u0_u24_ch_csr[6] , _u0_u24_ch_csr[5] ,_u0_u24_ch_csr[4] , _u0_u24_ch_csr[3] , _u0_u24_ch_csr[2] ,_u0_u24_ch_csr[1] , _u0_u24_ch_csr[0] , _u0_u24_ch_txsz[31] ,_u0_u24_ch_txsz[30] , _u0_u24_ch_txsz[29] , _u0_u24_ch_txsz[28] ,_u0_u24_ch_txsz[27] , _u0_u24_ch_txsz[26] , _u0_u24_ch_txsz[25] ,_u0_u24_ch_txsz[24] , _u0_u24_ch_txsz[23] , _u0_u24_ch_txsz[22] ,_u0_u24_ch_txsz[21] , _u0_u24_ch_txsz[20] , _u0_u24_ch_txsz[19] ,_u0_u24_ch_txsz[18] , _u0_u24_ch_txsz[17] , _u0_u24_ch_txsz[16] ,_u0_u24_ch_txsz[15] , _u0_u24_ch_txsz[14] , _u0_u24_ch_txsz[13] ,_u0_u24_ch_txsz[12] , _u0_u24_ch_txsz[11] , _u0_u24_ch_txsz[10] ,_u0_u24_ch_txsz[9] , _u0_u24_ch_txsz[8] , _u0_u24_ch_txsz[7] ,_u0_u24_ch_txsz[6] , _u0_u24_ch_txsz[5] , _u0_u24_ch_txsz[4] ,_u0_u24_ch_txsz[3] , _u0_u24_ch_txsz[2] , _u0_u24_ch_txsz[1] ,_u0_u24_ch_txsz[0] , _u0_u24_ch_adr0[31] , _u0_u24_ch_adr0[30] ,_u0_u24_ch_adr0[29] , _u0_u24_ch_adr0[28] , _u0_u24_ch_adr0[27] ,_u0_u24_ch_adr0[26] , _u0_u24_ch_adr0[25] , _u0_u24_ch_adr0[24] ,_u0_u24_ch_adr0[23] , _u0_u24_ch_adr0[22] , _u0_u24_ch_adr0[21] ,_u0_u24_ch_adr0[20] , _u0_u24_ch_adr0[19] , _u0_u24_ch_adr0[18] ,_u0_u24_ch_adr0[17] , _u0_u24_ch_adr0[16] , _u0_u24_ch_adr0[15] ,_u0_u24_ch_adr0[14] , _u0_u24_ch_adr0[13] , _u0_u24_ch_adr0[12] ,_u0_u24_ch_adr0[11] , _u0_u24_ch_adr0[10] , _u0_u24_ch_adr0[9] ,_u0_u24_ch_adr0[8] , _u0_u24_ch_adr0[7] , _u0_u24_ch_adr0[6] ,_u0_u24_ch_adr0[5] , _u0_u24_ch_adr0[4] , _u0_u24_ch_adr0[3] ,_u0_u24_ch_adr0[2] , _u0_u24_ch_adr0[1] , _u0_u24_ch_adr0[0] ,_u0_u24_ch_adr1[31] , _u0_u24_ch_adr1[30] , _u0_u24_ch_adr1[29] ,_u0_u24_ch_adr1[28] , _u0_u24_ch_adr1[27] , _u0_u24_ch_adr1[26] ,_u0_u24_ch_adr1[25] , _u0_u24_ch_adr1[24] , _u0_u24_ch_adr1[23] ,_u0_u24_ch_adr1[22] , _u0_u24_ch_adr1[21] , _u0_u24_ch_adr1[20] ,_u0_u24_ch_adr1[19] , _u0_u24_ch_adr1[18] , _u0_u24_ch_adr1[17] ,_u0_u24_ch_adr1[16] , _u0_u24_ch_adr1[15] , _u0_u24_ch_adr1[14] ,_u0_u24_ch_adr1[13] , _u0_u24_ch_adr1[12] , _u0_u24_ch_adr1[11] ,_u0_u24_ch_adr1[10] , _u0_u24_ch_adr1[9] , _u0_u24_ch_adr1[8] ,_u0_u24_ch_adr1[7] , _u0_u24_ch_adr1[6] , _u0_u24_ch_adr1[5] ,_u0_u24_ch_adr1[4] , _u0_u24_ch_adr1[3] , _u0_u24_ch_adr1[2] ,_u0_u24_ch_adr1[1] , _u0_u24_ch_adr1[0] , _u0_u24_ch_am0[31] ,_u0_u24_ch_am0[30] , _u0_u24_ch_am0[29] , _u0_u24_ch_am0[28] ,_u0_u24_ch_am0[27] , _u0_u24_ch_am0[26] , _u0_u24_ch_am0[25] ,_u0_u24_ch_am0[24] , _u0_u24_ch_am0[23] , _u0_u24_ch_am0[22] ,_u0_u24_ch_am0[21] , _u0_u24_ch_am0[20] , _u0_u24_ch_am0[19] ,_u0_u24_ch_am0[18] , _u0_u24_ch_am0[17] , _u0_u24_ch_am0[16] ,_u0_u24_ch_am0[15] , _u0_u24_ch_am0[14] , _u0_u24_ch_am0[13] ,_u0_u24_ch_am0[12] , _u0_u24_ch_am0[11] , _u0_u24_ch_am0[10] ,_u0_u24_ch_am0[9] , _u0_u24_ch_am0[8] , _u0_u24_ch_am0[7] ,_u0_u24_ch_am0[6] , _u0_u24_ch_am0[5] , _u0_u24_ch_am0[4] ,_u0_u24_ch_am0[3] , _u0_u24_ch_am0[2] , _u0_u24_ch_am0[1] ,_u0_u24_ch_am0[0] , _u0_u24_ch_am1[31] , _u0_u24_ch_am1[30] ,_u0_u24_ch_am1[29] , _u0_u24_ch_am1[28] , _u0_u24_ch_am1[27] ,_u0_u24_ch_am1[26] , _u0_u24_ch_am1[25] , _u0_u24_ch_am1[24] ,_u0_u24_ch_am1[23] , _u0_u24_ch_am1[22] , _u0_u24_ch_am1[21] ,_u0_u24_ch_am1[20] , _u0_u24_ch_am1[19] , _u0_u24_ch_am1[18] ,_u0_u24_ch_am1[17] , _u0_u24_ch_am1[16] , _u0_u24_ch_am1[15] ,_u0_u24_ch_am1[14] , _u0_u24_ch_am1[13] , _u0_u24_ch_am1[12] ,_u0_u24_ch_am1[11] , _u0_u24_ch_am1[10] , _u0_u24_ch_am1[9] ,_u0_u24_ch_am1[8] , _u0_u24_ch_am1[7] , _u0_u24_ch_am1[6] ,_u0_u24_ch_am1[5] , _u0_u24_ch_am1[4] , _u0_u24_ch_am1[3] ,_u0_u24_ch_am1[2] , _u0_u24_ch_am1[1] , _u0_u24_ch_am1[0] ,_u0_u24_sw_pointer[31] , _u0_u24_sw_pointer[30] ,_u0_u24_sw_pointer[29] , _u0_u24_sw_pointer[28] ,_u0_u24_sw_pointer[27] , _u0_u24_sw_pointer[26] ,_u0_u24_sw_pointer[25] , _u0_u24_sw_pointer[24] ,_u0_u24_sw_pointer[23] , _u0_u24_sw_pointer[22] ,_u0_u24_sw_pointer[21] , _u0_u24_sw_pointer[20] ,_u0_u24_sw_pointer[19] , _u0_u24_sw_pointer[18] ,_u0_u24_sw_pointer[17] , _u0_u24_sw_pointer[16] ,_u0_u24_sw_pointer[15] , _u0_u24_sw_pointer[14] ,_u0_u24_sw_pointer[13] , _u0_u24_sw_pointer[12] ,_u0_u24_sw_pointer[11] , _u0_u24_sw_pointer[10] ,_u0_u24_sw_pointer[9] , _u0_u24_sw_pointer[8] ,_u0_u24_sw_pointer[7] , _u0_u24_sw_pointer[6] ,_u0_u24_sw_pointer[5] , _u0_u24_sw_pointer[4] ,_u0_u24_sw_pointer[3] , _u0_u24_sw_pointer[2] ,_u0_u24_sw_pointer[1] , _u0_u24_sw_pointer[0] , _u0_u24_ch_stop ,_u0_u24_ch_dis , _u0_u24_int , _u0_u25_pointer[31] ,_u0_u25_pointer[30] , _u0_u25_pointer[29] , _u0_u25_pointer[28] ,_u0_u25_pointer[27] , _u0_u25_pointer[26] , _u0_u25_pointer[25] ,_u0_u25_pointer[24] , _u0_u25_pointer[23] , _u0_u25_pointer[22] ,_u0_u25_pointer[21] , _u0_u25_pointer[20] , _u0_u25_pointer[19] ,_u0_u25_pointer[18] , _u0_u25_pointer[17] , _u0_u25_pointer[16] ,_u0_u25_pointer[15] , _u0_u25_pointer[14] , _u0_u25_pointer[13] ,_u0_u25_pointer[12] , _u0_u25_pointer[11] , _u0_u25_pointer[10] ,_u0_u25_pointer[9] , _u0_u25_pointer[8] , _u0_u25_pointer[7] ,_u0_u25_pointer[6] , _u0_u25_pointer[5] , _u0_u25_pointer[4] ,_u0_u25_pointer[3] , _u0_u25_pointer[2] , _u0_u25_pointer[1] ,_u0_u25_pointer[0] , _u0_u25_pointer_s[31] , _u0_u25_pointer_s[30] ,_u0_u25_pointer_s[29] , _u0_u25_pointer_s[28] ,_u0_u25_pointer_s[27] , _u0_u25_pointer_s[26] ,_u0_u25_pointer_s[25] , _u0_u25_pointer_s[24] ,_u0_u25_pointer_s[23] , _u0_u25_pointer_s[22] ,_u0_u25_pointer_s[21] , _u0_u25_pointer_s[20] ,_u0_u25_pointer_s[19] , _u0_u25_pointer_s[18] ,_u0_u25_pointer_s[17] , _u0_u25_pointer_s[16] ,_u0_u25_pointer_s[15] , _u0_u25_pointer_s[14] ,_u0_u25_pointer_s[13] , _u0_u25_pointer_s[12] ,_u0_u25_pointer_s[11] , _u0_u25_pointer_s[10] , _u0_u25_pointer_s[9] ,_u0_u25_pointer_s[8] , _u0_u25_pointer_s[7] , _u0_u25_pointer_s[6] ,_u0_u25_pointer_s[5] , _u0_u25_pointer_s[4] , _u0_u25_pointer_s[3] ,_u0_u25_pointer_s[2] , _u0_u25_pointer_s[1] , _u0_u25_pointer_s[0] ,_u0_u25_ch_csr[31] , _u0_u25_ch_csr[30] , _u0_u25_ch_csr[29] ,_u0_u25_ch_csr[28] , _u0_u25_ch_csr[27] , _u0_u25_ch_csr[26] ,_u0_u25_ch_csr[25] , _u0_u25_ch_csr[24] , _u0_u25_ch_csr[23] ,_u0_u25_ch_csr[22] , _u0_u25_ch_csr[21] , _u0_u25_ch_csr[20] ,_u0_u25_ch_csr[19] , _u0_u25_ch_csr[18] , _u0_u25_ch_csr[17] ,_u0_u25_ch_csr[16] , _u0_u25_ch_csr[15] , _u0_u25_ch_csr[14] ,_u0_u25_ch_csr[13] , _u0_u25_ch_csr[12] , _u0_u25_ch_csr[11] ,_u0_u25_ch_csr[10] , _u0_u25_ch_csr[9] , _u0_u25_ch_csr[8] ,_u0_u25_ch_csr[7] , _u0_u25_ch_csr[6] , _u0_u25_ch_csr[5] ,_u0_u25_ch_csr[4] , _u0_u25_ch_csr[3] , _u0_u25_ch_csr[2] ,_u0_u25_ch_csr[1] , _u0_u25_ch_csr[0] , _u0_u25_ch_txsz[31] ,_u0_u25_ch_txsz[30] , _u0_u25_ch_txsz[29] , _u0_u25_ch_txsz[28] ,_u0_u25_ch_txsz[27] , _u0_u25_ch_txsz[26] , _u0_u25_ch_txsz[25] ,_u0_u25_ch_txsz[24] , _u0_u25_ch_txsz[23] , _u0_u25_ch_txsz[22] ,_u0_u25_ch_txsz[21] , _u0_u25_ch_txsz[20] , _u0_u25_ch_txsz[19] ,_u0_u25_ch_txsz[18] , _u0_u25_ch_txsz[17] , _u0_u25_ch_txsz[16] ,_u0_u25_ch_txsz[15] , _u0_u25_ch_txsz[14] , _u0_u25_ch_txsz[13] ,_u0_u25_ch_txsz[12] , _u0_u25_ch_txsz[11] , _u0_u25_ch_txsz[10] ,_u0_u25_ch_txsz[9] , _u0_u25_ch_txsz[8] , _u0_u25_ch_txsz[7] ,_u0_u25_ch_txsz[6] , _u0_u25_ch_txsz[5] , _u0_u25_ch_txsz[4] ,_u0_u25_ch_txsz[3] , _u0_u25_ch_txsz[2] , _u0_u25_ch_txsz[1] ,_u0_u25_ch_txsz[0] , _u0_u25_ch_adr0[31] , _u0_u25_ch_adr0[30] ,_u0_u25_ch_adr0[29] , _u0_u25_ch_adr0[28] , _u0_u25_ch_adr0[27] ,_u0_u25_ch_adr0[26] , _u0_u25_ch_adr0[25] , _u0_u25_ch_adr0[24] ,_u0_u25_ch_adr0[23] , _u0_u25_ch_adr0[22] , _u0_u25_ch_adr0[21] ,_u0_u25_ch_adr0[20] , _u0_u25_ch_adr0[19] , _u0_u25_ch_adr0[18] ,_u0_u25_ch_adr0[17] , _u0_u25_ch_adr0[16] , _u0_u25_ch_adr0[15] ,_u0_u25_ch_adr0[14] , _u0_u25_ch_adr0[13] , _u0_u25_ch_adr0[12] ,_u0_u25_ch_adr0[11] , _u0_u25_ch_adr0[10] , _u0_u25_ch_adr0[9] ,_u0_u25_ch_adr0[8] , _u0_u25_ch_adr0[7] , _u0_u25_ch_adr0[6] ,_u0_u25_ch_adr0[5] , _u0_u25_ch_adr0[4] , _u0_u25_ch_adr0[3] ,_u0_u25_ch_adr0[2] , _u0_u25_ch_adr0[1] , _u0_u25_ch_adr0[0] ,_u0_u25_ch_adr1[31] , _u0_u25_ch_adr1[30] , _u0_u25_ch_adr1[29] ,_u0_u25_ch_adr1[28] , _u0_u25_ch_adr1[27] , _u0_u25_ch_adr1[26] ,_u0_u25_ch_adr1[25] , _u0_u25_ch_adr1[24] , _u0_u25_ch_adr1[23] ,_u0_u25_ch_adr1[22] , _u0_u25_ch_adr1[21] , _u0_u25_ch_adr1[20] ,_u0_u25_ch_adr1[19] , _u0_u25_ch_adr1[18] , _u0_u25_ch_adr1[17] ,_u0_u25_ch_adr1[16] , _u0_u25_ch_adr1[15] , _u0_u25_ch_adr1[14] ,_u0_u25_ch_adr1[13] , _u0_u25_ch_adr1[12] , _u0_u25_ch_adr1[11] ,_u0_u25_ch_adr1[10] , _u0_u25_ch_adr1[9] , _u0_u25_ch_adr1[8] ,_u0_u25_ch_adr1[7] , _u0_u25_ch_adr1[6] , _u0_u25_ch_adr1[5] ,_u0_u25_ch_adr1[4] , _u0_u25_ch_adr1[3] , _u0_u25_ch_adr1[2] ,_u0_u25_ch_adr1[1] , _u0_u25_ch_adr1[0] , _u0_u25_ch_am0[31] ,_u0_u25_ch_am0[30] , _u0_u25_ch_am0[29] , _u0_u25_ch_am0[28] ,_u0_u25_ch_am0[27] , _u0_u25_ch_am0[26] , _u0_u25_ch_am0[25] ,_u0_u25_ch_am0[24] , _u0_u25_ch_am0[23] , _u0_u25_ch_am0[22] ,_u0_u25_ch_am0[21] , _u0_u25_ch_am0[20] , _u0_u25_ch_am0[19] ,_u0_u25_ch_am0[18] , _u0_u25_ch_am0[17] , _u0_u25_ch_am0[16] ,_u0_u25_ch_am0[15] , _u0_u25_ch_am0[14] , _u0_u25_ch_am0[13] ,_u0_u25_ch_am0[12] , _u0_u25_ch_am0[11] , _u0_u25_ch_am0[10] ,_u0_u25_ch_am0[9] , _u0_u25_ch_am0[8] , _u0_u25_ch_am0[7] ,_u0_u25_ch_am0[6] , _u0_u25_ch_am0[5] , _u0_u25_ch_am0[4] ,_u0_u25_ch_am0[3] , _u0_u25_ch_am0[2] , _u0_u25_ch_am0[1] ,_u0_u25_ch_am0[0] , _u0_u25_ch_am1[31] , _u0_u25_ch_am1[30] ,_u0_u25_ch_am1[29] , _u0_u25_ch_am1[28] , _u0_u25_ch_am1[27] ,_u0_u25_ch_am1[26] , _u0_u25_ch_am1[25] , _u0_u25_ch_am1[24] ,_u0_u25_ch_am1[23] , _u0_u25_ch_am1[22] , _u0_u25_ch_am1[21] ,_u0_u25_ch_am1[20] , _u0_u25_ch_am1[19] , _u0_u25_ch_am1[18] ,_u0_u25_ch_am1[17] , _u0_u25_ch_am1[16] , _u0_u25_ch_am1[15] ,_u0_u25_ch_am1[14] , _u0_u25_ch_am1[13] , _u0_u25_ch_am1[12] ,_u0_u25_ch_am1[11] , _u0_u25_ch_am1[10] , _u0_u25_ch_am1[9] ,_u0_u25_ch_am1[8] , _u0_u25_ch_am1[7] , _u0_u25_ch_am1[6] ,_u0_u25_ch_am1[5] , _u0_u25_ch_am1[4] , _u0_u25_ch_am1[3] ,_u0_u25_ch_am1[2] , _u0_u25_ch_am1[1] , _u0_u25_ch_am1[0] ,_u0_u25_sw_pointer[31] , _u0_u25_sw_pointer[30] ,_u0_u25_sw_pointer[29] , _u0_u25_sw_pointer[28] ,_u0_u25_sw_pointer[27] , _u0_u25_sw_pointer[26] ,_u0_u25_sw_pointer[25] , _u0_u25_sw_pointer[24] ,_u0_u25_sw_pointer[23] , _u0_u25_sw_pointer[22] ,_u0_u25_sw_pointer[21] , _u0_u25_sw_pointer[20] ,_u0_u25_sw_pointer[19] , _u0_u25_sw_pointer[18] ,_u0_u25_sw_pointer[17] , _u0_u25_sw_pointer[16] ,_u0_u25_sw_pointer[15] , _u0_u25_sw_pointer[14] ,_u0_u25_sw_pointer[13] , _u0_u25_sw_pointer[12] ,_u0_u25_sw_pointer[11] , _u0_u25_sw_pointer[10] ,_u0_u25_sw_pointer[9] , _u0_u25_sw_pointer[8] ,_u0_u25_sw_pointer[7] , _u0_u25_sw_pointer[6] ,_u0_u25_sw_pointer[5] , _u0_u25_sw_pointer[4] ,_u0_u25_sw_pointer[3] , _u0_u25_sw_pointer[2] ,_u0_u25_sw_pointer[1] , _u0_u25_sw_pointer[0] , _u0_u25_ch_stop ,_u0_u25_ch_dis , _u0_u25_int , _u0_u26_pointer[31] ,_u0_u26_pointer[30] , _u0_u26_pointer[29] , _u0_u26_pointer[28] ,_u0_u26_pointer[27] , _u0_u26_pointer[26] , _u0_u26_pointer[25] ,_u0_u26_pointer[24] , _u0_u26_pointer[23] , _u0_u26_pointer[22] ,_u0_u26_pointer[21] , _u0_u26_pointer[20] , _u0_u26_pointer[19] ,_u0_u26_pointer[18] , _u0_u26_pointer[17] , _u0_u26_pointer[16] ,_u0_u26_pointer[15] , _u0_u26_pointer[14] , _u0_u26_pointer[13] ,_u0_u26_pointer[12] , _u0_u26_pointer[11] , _u0_u26_pointer[10] ,_u0_u26_pointer[9] , _u0_u26_pointer[8] , _u0_u26_pointer[7] ,_u0_u26_pointer[6] , _u0_u26_pointer[5] , _u0_u26_pointer[4] ,_u0_u26_pointer[3] , _u0_u26_pointer[2] , _u0_u26_pointer[1] ,_u0_u26_pointer[0] , _u0_u26_pointer_s[31] , _u0_u26_pointer_s[30] ,_u0_u26_pointer_s[29] , _u0_u26_pointer_s[28] ,_u0_u26_pointer_s[27] , _u0_u26_pointer_s[26] ,_u0_u26_pointer_s[25] , _u0_u26_pointer_s[24] ,_u0_u26_pointer_s[23] , _u0_u26_pointer_s[22] ,_u0_u26_pointer_s[21] , _u0_u26_pointer_s[20] ,_u0_u26_pointer_s[19] , _u0_u26_pointer_s[18] ,_u0_u26_pointer_s[17] , _u0_u26_pointer_s[16] ,_u0_u26_pointer_s[15] , _u0_u26_pointer_s[14] ,_u0_u26_pointer_s[13] , _u0_u26_pointer_s[12] ,_u0_u26_pointer_s[11] , _u0_u26_pointer_s[10] , _u0_u26_pointer_s[9] ,_u0_u26_pointer_s[8] , _u0_u26_pointer_s[7] , _u0_u26_pointer_s[6] ,_u0_u26_pointer_s[5] , _u0_u26_pointer_s[4] , _u0_u26_pointer_s[3] ,_u0_u26_pointer_s[2] , _u0_u26_pointer_s[1] , _u0_u26_pointer_s[0] ,_u0_u26_ch_csr[31] , _u0_u26_ch_csr[30] , _u0_u26_ch_csr[29] ,_u0_u26_ch_csr[28] , _u0_u26_ch_csr[27] , _u0_u26_ch_csr[26] ,_u0_u26_ch_csr[25] , _u0_u26_ch_csr[24] , _u0_u26_ch_csr[23] ,_u0_u26_ch_csr[22] , _u0_u26_ch_csr[21] , _u0_u26_ch_csr[20] ,_u0_u26_ch_csr[19] , _u0_u26_ch_csr[18] , _u0_u26_ch_csr[17] ,_u0_u26_ch_csr[16] , _u0_u26_ch_csr[15] , _u0_u26_ch_csr[14] ,_u0_u26_ch_csr[13] , _u0_u26_ch_csr[12] , _u0_u26_ch_csr[11] ,_u0_u26_ch_csr[10] , _u0_u26_ch_csr[9] , _u0_u26_ch_csr[8] ,_u0_u26_ch_csr[7] , _u0_u26_ch_csr[6] , _u0_u26_ch_csr[5] ,_u0_u26_ch_csr[4] , _u0_u26_ch_csr[3] , _u0_u26_ch_csr[2] ,_u0_u26_ch_csr[1] , _u0_u26_ch_csr[0] , _u0_u26_ch_txsz[31] ,_u0_u26_ch_txsz[30] , _u0_u26_ch_txsz[29] , _u0_u26_ch_txsz[28] ,_u0_u26_ch_txsz[27] , _u0_u26_ch_txsz[26] , _u0_u26_ch_txsz[25] ,_u0_u26_ch_txsz[24] , _u0_u26_ch_txsz[23] , _u0_u26_ch_txsz[22] ,_u0_u26_ch_txsz[21] , _u0_u26_ch_txsz[20] , _u0_u26_ch_txsz[19] ,_u0_u26_ch_txsz[18] , _u0_u26_ch_txsz[17] , _u0_u26_ch_txsz[16] ,_u0_u26_ch_txsz[15] , _u0_u26_ch_txsz[14] , _u0_u26_ch_txsz[13] ,_u0_u26_ch_txsz[12] , _u0_u26_ch_txsz[11] , _u0_u26_ch_txsz[10] ,_u0_u26_ch_txsz[9] , _u0_u26_ch_txsz[8] , _u0_u26_ch_txsz[7] ,_u0_u26_ch_txsz[6] , _u0_u26_ch_txsz[5] , _u0_u26_ch_txsz[4] ,_u0_u26_ch_txsz[3] , _u0_u26_ch_txsz[2] , _u0_u26_ch_txsz[1] ,_u0_u26_ch_txsz[0] , _u0_u26_ch_adr0[31] , _u0_u26_ch_adr0[30] ,_u0_u26_ch_adr0[29] , _u0_u26_ch_adr0[28] , _u0_u26_ch_adr0[27] ,_u0_u26_ch_adr0[26] , _u0_u26_ch_adr0[25] , _u0_u26_ch_adr0[24] ,_u0_u26_ch_adr0[23] , _u0_u26_ch_adr0[22] , _u0_u26_ch_adr0[21] ,_u0_u26_ch_adr0[20] , _u0_u26_ch_adr0[19] , _u0_u26_ch_adr0[18] ,_u0_u26_ch_adr0[17] , _u0_u26_ch_adr0[16] , _u0_u26_ch_adr0[15] ,_u0_u26_ch_adr0[14] , _u0_u26_ch_adr0[13] , _u0_u26_ch_adr0[12] ,_u0_u26_ch_adr0[11] , _u0_u26_ch_adr0[10] , _u0_u26_ch_adr0[9] ,_u0_u26_ch_adr0[8] , _u0_u26_ch_adr0[7] , _u0_u26_ch_adr0[6] ,_u0_u26_ch_adr0[5] , _u0_u26_ch_adr0[4] , _u0_u26_ch_adr0[3] ,_u0_u26_ch_adr0[2] , _u0_u26_ch_adr0[1] , _u0_u26_ch_adr0[0] ,_u0_u26_ch_adr1[31] , _u0_u26_ch_adr1[30] , _u0_u26_ch_adr1[29] ,_u0_u26_ch_adr1[28] , _u0_u26_ch_adr1[27] , _u0_u26_ch_adr1[26] ,_u0_u26_ch_adr1[25] , _u0_u26_ch_adr1[24] , _u0_u26_ch_adr1[23] ,_u0_u26_ch_adr1[22] , _u0_u26_ch_adr1[21] , _u0_u26_ch_adr1[20] ,_u0_u26_ch_adr1[19] , _u0_u26_ch_adr1[18] , _u0_u26_ch_adr1[17] ,_u0_u26_ch_adr1[16] , _u0_u26_ch_adr1[15] , _u0_u26_ch_adr1[14] ,_u0_u26_ch_adr1[13] , _u0_u26_ch_adr1[12] , _u0_u26_ch_adr1[11] ,_u0_u26_ch_adr1[10] , _u0_u26_ch_adr1[9] , _u0_u26_ch_adr1[8] ,_u0_u26_ch_adr1[7] , _u0_u26_ch_adr1[6] , _u0_u26_ch_adr1[5] ,_u0_u26_ch_adr1[4] , _u0_u26_ch_adr1[3] , _u0_u26_ch_adr1[2] ,_u0_u26_ch_adr1[1] , _u0_u26_ch_adr1[0] , _u0_u26_ch_am0[31] ,_u0_u26_ch_am0[30] , _u0_u26_ch_am0[29] , _u0_u26_ch_am0[28] ,_u0_u26_ch_am0[27] , _u0_u26_ch_am0[26] , _u0_u26_ch_am0[25] ,_u0_u26_ch_am0[24] , _u0_u26_ch_am0[23] , _u0_u26_ch_am0[22] ,_u0_u26_ch_am0[21] , _u0_u26_ch_am0[20] , _u0_u26_ch_am0[19] ,_u0_u26_ch_am0[18] , _u0_u26_ch_am0[17] , _u0_u26_ch_am0[16] ,_u0_u26_ch_am0[15] , _u0_u26_ch_am0[14] , _u0_u26_ch_am0[13] ,_u0_u26_ch_am0[12] , _u0_u26_ch_am0[11] , _u0_u26_ch_am0[10] ,_u0_u26_ch_am0[9] , _u0_u26_ch_am0[8] , _u0_u26_ch_am0[7] ,_u0_u26_ch_am0[6] , _u0_u26_ch_am0[5] , _u0_u26_ch_am0[4] ,_u0_u26_ch_am0[3] , _u0_u26_ch_am0[2] , _u0_u26_ch_am0[1] ,_u0_u26_ch_am0[0] , _u0_u26_ch_am1[31] , _u0_u26_ch_am1[30] ,_u0_u26_ch_am1[29] , _u0_u26_ch_am1[28] , _u0_u26_ch_am1[27] ,_u0_u26_ch_am1[26] , _u0_u26_ch_am1[25] , _u0_u26_ch_am1[24] ,_u0_u26_ch_am1[23] , _u0_u26_ch_am1[22] , _u0_u26_ch_am1[21] ,_u0_u26_ch_am1[20] , _u0_u26_ch_am1[19] , _u0_u26_ch_am1[18] ,_u0_u26_ch_am1[17] , _u0_u26_ch_am1[16] , _u0_u26_ch_am1[15] ,_u0_u26_ch_am1[14] , _u0_u26_ch_am1[13] , _u0_u26_ch_am1[12] ,_u0_u26_ch_am1[11] , _u0_u26_ch_am1[10] , _u0_u26_ch_am1[9] ,_u0_u26_ch_am1[8] , _u0_u26_ch_am1[7] , _u0_u26_ch_am1[6] ,_u0_u26_ch_am1[5] , _u0_u26_ch_am1[4] , _u0_u26_ch_am1[3] ,_u0_u26_ch_am1[2] , _u0_u26_ch_am1[1] , _u0_u26_ch_am1[0] ,_u0_u26_sw_pointer[31] , _u0_u26_sw_pointer[30] ,_u0_u26_sw_pointer[29] , _u0_u26_sw_pointer[28] ,_u0_u26_sw_pointer[27] , _u0_u26_sw_pointer[26] ,_u0_u26_sw_pointer[25] , _u0_u26_sw_pointer[24] ,_u0_u26_sw_pointer[23] , _u0_u26_sw_pointer[22] ,_u0_u26_sw_pointer[21] , _u0_u26_sw_pointer[20] ,_u0_u26_sw_pointer[19] , _u0_u26_sw_pointer[18] ,_u0_u26_sw_pointer[17] , _u0_u26_sw_pointer[16] ,_u0_u26_sw_pointer[15] , _u0_u26_sw_pointer[14] ,_u0_u26_sw_pointer[13] , _u0_u26_sw_pointer[12] ,_u0_u26_sw_pointer[11] , _u0_u26_sw_pointer[10] ,_u0_u26_sw_pointer[9] , _u0_u26_sw_pointer[8] ,_u0_u26_sw_pointer[7] , _u0_u26_sw_pointer[6] ,_u0_u26_sw_pointer[5] , _u0_u26_sw_pointer[4] ,_u0_u26_sw_pointer[3] , _u0_u26_sw_pointer[2] ,_u0_u26_sw_pointer[1] , _u0_u26_sw_pointer[0] , _u0_u26_ch_stop ,_u0_u26_ch_dis , _u0_u26_int , _u0_u27_pointer[31] ,_u0_u27_pointer[30] , _u0_u27_pointer[29] , _u0_u27_pointer[28] ,_u0_u27_pointer[27] , _u0_u27_pointer[26] , _u0_u27_pointer[25] ,_u0_u27_pointer[24] , _u0_u27_pointer[23] , _u0_u27_pointer[22] ,_u0_u27_pointer[21] , _u0_u27_pointer[20] , _u0_u27_pointer[19] ,_u0_u27_pointer[18] , _u0_u27_pointer[17] , _u0_u27_pointer[16] ,_u0_u27_pointer[15] , _u0_u27_pointer[14] , _u0_u27_pointer[13] ,_u0_u27_pointer[12] , _u0_u27_pointer[11] , _u0_u27_pointer[10] ,_u0_u27_pointer[9] , _u0_u27_pointer[8] , _u0_u27_pointer[7] ,_u0_u27_pointer[6] , _u0_u27_pointer[5] , _u0_u27_pointer[4] ,_u0_u27_pointer[3] , _u0_u27_pointer[2] , _u0_u27_pointer[1] ,_u0_u27_pointer[0] , _u0_u27_pointer_s[31] , _u0_u27_pointer_s[30] ,_u0_u27_pointer_s[29] , _u0_u27_pointer_s[28] ,_u0_u27_pointer_s[27] , _u0_u27_pointer_s[26] ,_u0_u27_pointer_s[25] , _u0_u27_pointer_s[24] ,_u0_u27_pointer_s[23] , _u0_u27_pointer_s[22] ,_u0_u27_pointer_s[21] , _u0_u27_pointer_s[20] ,_u0_u27_pointer_s[19] , _u0_u27_pointer_s[18] ,_u0_u27_pointer_s[17] , _u0_u27_pointer_s[16] ,_u0_u27_pointer_s[15] , _u0_u27_pointer_s[14] ,_u0_u27_pointer_s[13] , _u0_u27_pointer_s[12] ,_u0_u27_pointer_s[11] , _u0_u27_pointer_s[10] , _u0_u27_pointer_s[9] ,_u0_u27_pointer_s[8] , _u0_u27_pointer_s[7] , _u0_u27_pointer_s[6] ,_u0_u27_pointer_s[5] , _u0_u27_pointer_s[4] , _u0_u27_pointer_s[3] ,_u0_u27_pointer_s[2] , _u0_u27_pointer_s[1] , _u0_u27_pointer_s[0] ,_u0_u27_ch_csr[31] , _u0_u27_ch_csr[30] , _u0_u27_ch_csr[29] ,_u0_u27_ch_csr[28] , _u0_u27_ch_csr[27] , _u0_u27_ch_csr[26] ,_u0_u27_ch_csr[25] , _u0_u27_ch_csr[24] , _u0_u27_ch_csr[23] ,_u0_u27_ch_csr[22] , _u0_u27_ch_csr[21] , _u0_u27_ch_csr[20] ,_u0_u27_ch_csr[19] , _u0_u27_ch_csr[18] , _u0_u27_ch_csr[17] ,_u0_u27_ch_csr[16] , _u0_u27_ch_csr[15] , _u0_u27_ch_csr[14] ,_u0_u27_ch_csr[13] , _u0_u27_ch_csr[12] , _u0_u27_ch_csr[11] ,_u0_u27_ch_csr[10] , _u0_u27_ch_csr[9] , _u0_u27_ch_csr[8] ,_u0_u27_ch_csr[7] , _u0_u27_ch_csr[6] , _u0_u27_ch_csr[5] ,_u0_u27_ch_csr[4] , _u0_u27_ch_csr[3] , _u0_u27_ch_csr[2] ,_u0_u27_ch_csr[1] , _u0_u27_ch_csr[0] , _u0_u27_ch_txsz[31] ,_u0_u27_ch_txsz[30] , _u0_u27_ch_txsz[29] , _u0_u27_ch_txsz[28] ,_u0_u27_ch_txsz[27] , _u0_u27_ch_txsz[26] , _u0_u27_ch_txsz[25] ,_u0_u27_ch_txsz[24] , _u0_u27_ch_txsz[23] , _u0_u27_ch_txsz[22] ,_u0_u27_ch_txsz[21] , _u0_u27_ch_txsz[20] , _u0_u27_ch_txsz[19] ,_u0_u27_ch_txsz[18] , _u0_u27_ch_txsz[17] , _u0_u27_ch_txsz[16] ,_u0_u27_ch_txsz[15] , _u0_u27_ch_txsz[14] , _u0_u27_ch_txsz[13] ,_u0_u27_ch_txsz[12] , _u0_u27_ch_txsz[11] , _u0_u27_ch_txsz[10] ,_u0_u27_ch_txsz[9] , _u0_u27_ch_txsz[8] , _u0_u27_ch_txsz[7] ,_u0_u27_ch_txsz[6] , _u0_u27_ch_txsz[5] , _u0_u27_ch_txsz[4] ,_u0_u27_ch_txsz[3] , _u0_u27_ch_txsz[2] , _u0_u27_ch_txsz[1] ,_u0_u27_ch_txsz[0] , _u0_u27_ch_adr0[31] , _u0_u27_ch_adr0[30] ,_u0_u27_ch_adr0[29] , _u0_u27_ch_adr0[28] , _u0_u27_ch_adr0[27] ,_u0_u27_ch_adr0[26] , _u0_u27_ch_adr0[25] , _u0_u27_ch_adr0[24] ,_u0_u27_ch_adr0[23] , _u0_u27_ch_adr0[22] , _u0_u27_ch_adr0[21] ,_u0_u27_ch_adr0[20] , _u0_u27_ch_adr0[19] , _u0_u27_ch_adr0[18] ,_u0_u27_ch_adr0[17] , _u0_u27_ch_adr0[16] , _u0_u27_ch_adr0[15] ,_u0_u27_ch_adr0[14] , _u0_u27_ch_adr0[13] , _u0_u27_ch_adr0[12] ,_u0_u27_ch_adr0[11] , _u0_u27_ch_adr0[10] , _u0_u27_ch_adr0[9] ,_u0_u27_ch_adr0[8] , _u0_u27_ch_adr0[7] , _u0_u27_ch_adr0[6] ,_u0_u27_ch_adr0[5] , _u0_u27_ch_adr0[4] , _u0_u27_ch_adr0[3] ,_u0_u27_ch_adr0[2] , _u0_u27_ch_adr0[1] , _u0_u27_ch_adr0[0] ,_u0_u27_ch_adr1[31] , _u0_u27_ch_adr1[30] , _u0_u27_ch_adr1[29] ,_u0_u27_ch_adr1[28] , _u0_u27_ch_adr1[27] , _u0_u27_ch_adr1[26] ,_u0_u27_ch_adr1[25] , _u0_u27_ch_adr1[24] , _u0_u27_ch_adr1[23] ,_u0_u27_ch_adr1[22] , _u0_u27_ch_adr1[21] , _u0_u27_ch_adr1[20] ,_u0_u27_ch_adr1[19] , _u0_u27_ch_adr1[18] , _u0_u27_ch_adr1[17] ,_u0_u27_ch_adr1[16] , _u0_u27_ch_adr1[15] , _u0_u27_ch_adr1[14] ,_u0_u27_ch_adr1[13] , _u0_u27_ch_adr1[12] , _u0_u27_ch_adr1[11] ,_u0_u27_ch_adr1[10] , _u0_u27_ch_adr1[9] , _u0_u27_ch_adr1[8] ,_u0_u27_ch_adr1[7] , _u0_u27_ch_adr1[6] , _u0_u27_ch_adr1[5] ,_u0_u27_ch_adr1[4] , _u0_u27_ch_adr1[3] , _u0_u27_ch_adr1[2] ,_u0_u27_ch_adr1[1] , _u0_u27_ch_adr1[0] , _u0_u27_ch_am0[31] ,_u0_u27_ch_am0[30] , _u0_u27_ch_am0[29] , _u0_u27_ch_am0[28] ,_u0_u27_ch_am0[27] , _u0_u27_ch_am0[26] , _u0_u27_ch_am0[25] ,_u0_u27_ch_am0[24] , _u0_u27_ch_am0[23] , _u0_u27_ch_am0[22] ,_u0_u27_ch_am0[21] , _u0_u27_ch_am0[20] , _u0_u27_ch_am0[19] ,_u0_u27_ch_am0[18] , _u0_u27_ch_am0[17] , _u0_u27_ch_am0[16] ,_u0_u27_ch_am0[15] , _u0_u27_ch_am0[14] , _u0_u27_ch_am0[13] ,_u0_u27_ch_am0[12] , _u0_u27_ch_am0[11] , _u0_u27_ch_am0[10] ,_u0_u27_ch_am0[9] , _u0_u27_ch_am0[8] , _u0_u27_ch_am0[7] ,_u0_u27_ch_am0[6] , _u0_u27_ch_am0[5] , _u0_u27_ch_am0[4] ,_u0_u27_ch_am0[3] , _u0_u27_ch_am0[2] , _u0_u27_ch_am0[1] ,_u0_u27_ch_am0[0] , _u0_u27_ch_am1[31] , _u0_u27_ch_am1[30] ,_u0_u27_ch_am1[29] , _u0_u27_ch_am1[28] , _u0_u27_ch_am1[27] ,_u0_u27_ch_am1[26] , _u0_u27_ch_am1[25] , _u0_u27_ch_am1[24] ,_u0_u27_ch_am1[23] , _u0_u27_ch_am1[22] , _u0_u27_ch_am1[21] ,_u0_u27_ch_am1[20] , _u0_u27_ch_am1[19] , _u0_u27_ch_am1[18] ,_u0_u27_ch_am1[17] , _u0_u27_ch_am1[16] , _u0_u27_ch_am1[15] ,_u0_u27_ch_am1[14] , _u0_u27_ch_am1[13] , _u0_u27_ch_am1[12] ,_u0_u27_ch_am1[11] , _u0_u27_ch_am1[10] , _u0_u27_ch_am1[9] ,_u0_u27_ch_am1[8] , _u0_u27_ch_am1[7] , _u0_u27_ch_am1[6] ,_u0_u27_ch_am1[5] , _u0_u27_ch_am1[4] , _u0_u27_ch_am1[3] ,_u0_u27_ch_am1[2] , _u0_u27_ch_am1[1] , _u0_u27_ch_am1[0] ,_u0_u27_sw_pointer[31] , _u0_u27_sw_pointer[30] ,_u0_u27_sw_pointer[29] , _u0_u27_sw_pointer[28] ,_u0_u27_sw_pointer[27] , _u0_u27_sw_pointer[26] ,_u0_u27_sw_pointer[25] , _u0_u27_sw_pointer[24] ,_u0_u27_sw_pointer[23] , _u0_u27_sw_pointer[22] ,_u0_u27_sw_pointer[21] , _u0_u27_sw_pointer[20] ,_u0_u27_sw_pointer[19] , _u0_u27_sw_pointer[18] ,_u0_u27_sw_pointer[17] , _u0_u27_sw_pointer[16] ,_u0_u27_sw_pointer[15] , _u0_u27_sw_pointer[14] ,_u0_u27_sw_pointer[13] , _u0_u27_sw_pointer[12] ,_u0_u27_sw_pointer[11] , _u0_u27_sw_pointer[10] ,_u0_u27_sw_pointer[9] , _u0_u27_sw_pointer[8] ,_u0_u27_sw_pointer[7] , _u0_u27_sw_pointer[6] ,_u0_u27_sw_pointer[5] , _u0_u27_sw_pointer[4] ,_u0_u27_sw_pointer[3] , _u0_u27_sw_pointer[2] ,_u0_u27_sw_pointer[1] , _u0_u27_sw_pointer[0] , _u0_u27_ch_stop ,_u0_u27_ch_dis , _u0_u27_int , _u0_u28_pointer[31] ,_u0_u28_pointer[30] , _u0_u28_pointer[29] , _u0_u28_pointer[28] ,_u0_u28_pointer[27] , _u0_u28_pointer[26] , _u0_u28_pointer[25] ,_u0_u28_pointer[24] , _u0_u28_pointer[23] , _u0_u28_pointer[22] ,_u0_u28_pointer[21] , _u0_u28_pointer[20] , _u0_u28_pointer[19] ,_u0_u28_pointer[18] , _u0_u28_pointer[17] , _u0_u28_pointer[16] ,_u0_u28_pointer[15] , _u0_u28_pointer[14] , _u0_u28_pointer[13] ,_u0_u28_pointer[12] , _u0_u28_pointer[11] , _u0_u28_pointer[10] ,_u0_u28_pointer[9] , _u0_u28_pointer[8] , _u0_u28_pointer[7] ,_u0_u28_pointer[6] , _u0_u28_pointer[5] , _u0_u28_pointer[4] ,_u0_u28_pointer[3] , _u0_u28_pointer[2] , _u0_u28_pointer[1] ,_u0_u28_pointer[0] , _u0_u28_pointer_s[31] , _u0_u28_pointer_s[30] ,_u0_u28_pointer_s[29] , _u0_u28_pointer_s[28] ,_u0_u28_pointer_s[27] , _u0_u28_pointer_s[26] ,_u0_u28_pointer_s[25] , _u0_u28_pointer_s[24] ,_u0_u28_pointer_s[23] , _u0_u28_pointer_s[22] ,_u0_u28_pointer_s[21] , _u0_u28_pointer_s[20] ,_u0_u28_pointer_s[19] , _u0_u28_pointer_s[18] ,_u0_u28_pointer_s[17] , _u0_u28_pointer_s[16] ,_u0_u28_pointer_s[15] , _u0_u28_pointer_s[14] ,_u0_u28_pointer_s[13] , _u0_u28_pointer_s[12] ,_u0_u28_pointer_s[11] , _u0_u28_pointer_s[10] , _u0_u28_pointer_s[9] ,_u0_u28_pointer_s[8] , _u0_u28_pointer_s[7] , _u0_u28_pointer_s[6] ,_u0_u28_pointer_s[5] , _u0_u28_pointer_s[4] , _u0_u28_pointer_s[3] ,_u0_u28_pointer_s[2] , _u0_u28_pointer_s[1] , _u0_u28_pointer_s[0] ,_u0_u28_ch_csr[31] , _u0_u28_ch_csr[30] , _u0_u28_ch_csr[29] ,_u0_u28_ch_csr[28] , _u0_u28_ch_csr[27] , _u0_u28_ch_csr[26] ,_u0_u28_ch_csr[25] , _u0_u28_ch_csr[24] , _u0_u28_ch_csr[23] ,_u0_u28_ch_csr[22] , _u0_u28_ch_csr[21] , _u0_u28_ch_csr[20] ,_u0_u28_ch_csr[19] , _u0_u28_ch_csr[18] , _u0_u28_ch_csr[17] ,_u0_u28_ch_csr[16] , _u0_u28_ch_csr[15] , _u0_u28_ch_csr[14] ,_u0_u28_ch_csr[13] , _u0_u28_ch_csr[12] , _u0_u28_ch_csr[11] ,_u0_u28_ch_csr[10] , _u0_u28_ch_csr[9] , _u0_u28_ch_csr[8] ,_u0_u28_ch_csr[7] , _u0_u28_ch_csr[6] , _u0_u28_ch_csr[5] ,_u0_u28_ch_csr[4] , _u0_u28_ch_csr[3] , _u0_u28_ch_csr[2] ,_u0_u28_ch_csr[1] , _u0_u28_ch_csr[0] , _u0_u28_ch_txsz[31] ,_u0_u28_ch_txsz[30] , _u0_u28_ch_txsz[29] , _u0_u28_ch_txsz[28] ,_u0_u28_ch_txsz[27] , _u0_u28_ch_txsz[26] , _u0_u28_ch_txsz[25] ,_u0_u28_ch_txsz[24] , _u0_u28_ch_txsz[23] , _u0_u28_ch_txsz[22] ,_u0_u28_ch_txsz[21] , _u0_u28_ch_txsz[20] , _u0_u28_ch_txsz[19] ,_u0_u28_ch_txsz[18] , _u0_u28_ch_txsz[17] , _u0_u28_ch_txsz[16] ,_u0_u28_ch_txsz[15] , _u0_u28_ch_txsz[14] , _u0_u28_ch_txsz[13] ,_u0_u28_ch_txsz[12] , _u0_u28_ch_txsz[11] , _u0_u28_ch_txsz[10] ,_u0_u28_ch_txsz[9] , _u0_u28_ch_txsz[8] , _u0_u28_ch_txsz[7] ,_u0_u28_ch_txsz[6] , _u0_u28_ch_txsz[5] , _u0_u28_ch_txsz[4] ,_u0_u28_ch_txsz[3] , _u0_u28_ch_txsz[2] , _u0_u28_ch_txsz[1] ,_u0_u28_ch_txsz[0] , _u0_u28_ch_adr0[31] , _u0_u28_ch_adr0[30] ,_u0_u28_ch_adr0[29] , _u0_u28_ch_adr0[28] , _u0_u28_ch_adr0[27] ,_u0_u28_ch_adr0[26] , _u0_u28_ch_adr0[25] , _u0_u28_ch_adr0[24] ,_u0_u28_ch_adr0[23] , _u0_u28_ch_adr0[22] , _u0_u28_ch_adr0[21] ,_u0_u28_ch_adr0[20] , _u0_u28_ch_adr0[19] , _u0_u28_ch_adr0[18] ,_u0_u28_ch_adr0[17] , _u0_u28_ch_adr0[16] , _u0_u28_ch_adr0[15] ,_u0_u28_ch_adr0[14] , _u0_u28_ch_adr0[13] , _u0_u28_ch_adr0[12] ,_u0_u28_ch_adr0[11] , _u0_u28_ch_adr0[10] , _u0_u28_ch_adr0[9] ,_u0_u28_ch_adr0[8] , _u0_u28_ch_adr0[7] , _u0_u28_ch_adr0[6] ,_u0_u28_ch_adr0[5] , _u0_u28_ch_adr0[4] , _u0_u28_ch_adr0[3] ,_u0_u28_ch_adr0[2] , _u0_u28_ch_adr0[1] , _u0_u28_ch_adr0[0] ,_u0_u28_ch_adr1[31] , _u0_u28_ch_adr1[30] , _u0_u28_ch_adr1[29] ,_u0_u28_ch_adr1[28] , _u0_u28_ch_adr1[27] , _u0_u28_ch_adr1[26] ,_u0_u28_ch_adr1[25] , _u0_u28_ch_adr1[24] , _u0_u28_ch_adr1[23] ,_u0_u28_ch_adr1[22] , _u0_u28_ch_adr1[21] , _u0_u28_ch_adr1[20] ,_u0_u28_ch_adr1[19] , _u0_u28_ch_adr1[18] , _u0_u28_ch_adr1[17] ,_u0_u28_ch_adr1[16] , _u0_u28_ch_adr1[15] , _u0_u28_ch_adr1[14] ,_u0_u28_ch_adr1[13] , _u0_u28_ch_adr1[12] , _u0_u28_ch_adr1[11] ,_u0_u28_ch_adr1[10] , _u0_u28_ch_adr1[9] , _u0_u28_ch_adr1[8] ,_u0_u28_ch_adr1[7] , _u0_u28_ch_adr1[6] , _u0_u28_ch_adr1[5] ,_u0_u28_ch_adr1[4] , _u0_u28_ch_adr1[3] , _u0_u28_ch_adr1[2] ,_u0_u28_ch_adr1[1] , _u0_u28_ch_adr1[0] , _u0_u28_ch_am0[31] ,_u0_u28_ch_am0[30] , _u0_u28_ch_am0[29] , _u0_u28_ch_am0[28] ,_u0_u28_ch_am0[27] , _u0_u28_ch_am0[26] , _u0_u28_ch_am0[25] ,_u0_u28_ch_am0[24] , _u0_u28_ch_am0[23] , _u0_u28_ch_am0[22] ,_u0_u28_ch_am0[21] , _u0_u28_ch_am0[20] , _u0_u28_ch_am0[19] ,_u0_u28_ch_am0[18] , _u0_u28_ch_am0[17] , _u0_u28_ch_am0[16] ,_u0_u28_ch_am0[15] , _u0_u28_ch_am0[14] , _u0_u28_ch_am0[13] ,_u0_u28_ch_am0[12] , _u0_u28_ch_am0[11] , _u0_u28_ch_am0[10] ,_u0_u28_ch_am0[9] , _u0_u28_ch_am0[8] , _u0_u28_ch_am0[7] ,_u0_u28_ch_am0[6] , _u0_u28_ch_am0[5] , _u0_u28_ch_am0[4] ,_u0_u28_ch_am0[3] , _u0_u28_ch_am0[2] , _u0_u28_ch_am0[1] ,_u0_u28_ch_am0[0] , _u0_u28_ch_am1[31] , _u0_u28_ch_am1[30] ,_u0_u28_ch_am1[29] , _u0_u28_ch_am1[28] , _u0_u28_ch_am1[27] ,_u0_u28_ch_am1[26] , _u0_u28_ch_am1[25] , _u0_u28_ch_am1[24] ,_u0_u28_ch_am1[23] , _u0_u28_ch_am1[22] , _u0_u28_ch_am1[21] ,_u0_u28_ch_am1[20] , _u0_u28_ch_am1[19] , _u0_u28_ch_am1[18] ,_u0_u28_ch_am1[17] , _u0_u28_ch_am1[16] , _u0_u28_ch_am1[15] ,_u0_u28_ch_am1[14] , _u0_u28_ch_am1[13] , _u0_u28_ch_am1[12] ,_u0_u28_ch_am1[11] , _u0_u28_ch_am1[10] , _u0_u28_ch_am1[9] ,_u0_u28_ch_am1[8] , _u0_u28_ch_am1[7] , _u0_u28_ch_am1[6] ,_u0_u28_ch_am1[5] , _u0_u28_ch_am1[4] , _u0_u28_ch_am1[3] ,_u0_u28_ch_am1[2] , _u0_u28_ch_am1[1] , _u0_u28_ch_am1[0] ,_u0_u28_sw_pointer[31] , _u0_u28_sw_pointer[30] ,_u0_u28_sw_pointer[29] , _u0_u28_sw_pointer[28] ,_u0_u28_sw_pointer[27] , _u0_u28_sw_pointer[26] ,_u0_u28_sw_pointer[25] , _u0_u28_sw_pointer[24] ,_u0_u28_sw_pointer[23] , _u0_u28_sw_pointer[22] ,_u0_u28_sw_pointer[21] , _u0_u28_sw_pointer[20] ,_u0_u28_sw_pointer[19] , _u0_u28_sw_pointer[18] ,_u0_u28_sw_pointer[17] , _u0_u28_sw_pointer[16] ,_u0_u28_sw_pointer[15] , _u0_u28_sw_pointer[14] ,_u0_u28_sw_pointer[13] , _u0_u28_sw_pointer[12] ,_u0_u28_sw_pointer[11] , _u0_u28_sw_pointer[10] ,_u0_u28_sw_pointer[9] , _u0_u28_sw_pointer[8] ,_u0_u28_sw_pointer[7] , _u0_u28_sw_pointer[6] ,_u0_u28_sw_pointer[5] , _u0_u28_sw_pointer[4] ,_u0_u28_sw_pointer[3] , _u0_u28_sw_pointer[2] ,_u0_u28_sw_pointer[1] , _u0_u28_sw_pointer[0] , _u0_u28_ch_stop ,_u0_u28_ch_dis , _u0_u28_int , _u0_u29_pointer[31] ,_u0_u29_pointer[30] , _u0_u29_pointer[29] , _u0_u29_pointer[28] ,_u0_u29_pointer[27] , _u0_u29_pointer[26] , _u0_u29_pointer[25] ,_u0_u29_pointer[24] , _u0_u29_pointer[23] , _u0_u29_pointer[22] ,_u0_u29_pointer[21] , _u0_u29_pointer[20] , _u0_u29_pointer[19] ,_u0_u29_pointer[18] , _u0_u29_pointer[17] , _u0_u29_pointer[16] ,_u0_u29_pointer[15] , _u0_u29_pointer[14] , _u0_u29_pointer[13] ,_u0_u29_pointer[12] , _u0_u29_pointer[11] , _u0_u29_pointer[10] ,_u0_u29_pointer[9] , _u0_u29_pointer[8] , _u0_u29_pointer[7] ,_u0_u29_pointer[6] , _u0_u29_pointer[5] , _u0_u29_pointer[4] ,_u0_u29_pointer[3] , _u0_u29_pointer[2] , _u0_u29_pointer[1] ,_u0_u29_pointer[0] , _u0_u29_pointer_s[31] , _u0_u29_pointer_s[30] ,_u0_u29_pointer_s[29] , _u0_u29_pointer_s[28] ,_u0_u29_pointer_s[27] , _u0_u29_pointer_s[26] ,_u0_u29_pointer_s[25] , _u0_u29_pointer_s[24] ,_u0_u29_pointer_s[23] , _u0_u29_pointer_s[22] ,_u0_u29_pointer_s[21] , _u0_u29_pointer_s[20] ,_u0_u29_pointer_s[19] , _u0_u29_pointer_s[18] ,_u0_u29_pointer_s[17] , _u0_u29_pointer_s[16] ,_u0_u29_pointer_s[15] , _u0_u29_pointer_s[14] ,_u0_u29_pointer_s[13] , _u0_u29_pointer_s[12] ,_u0_u29_pointer_s[11] , _u0_u29_pointer_s[10] , _u0_u29_pointer_s[9] ,_u0_u29_pointer_s[8] , _u0_u29_pointer_s[7] , _u0_u29_pointer_s[6] ,_u0_u29_pointer_s[5] , _u0_u29_pointer_s[4] , _u0_u29_pointer_s[3] ,_u0_u29_pointer_s[2] , _u0_u29_pointer_s[1] , _u0_u29_pointer_s[0] ,_u0_u29_ch_csr[31] , _u0_u29_ch_csr[30] , _u0_u29_ch_csr[29] ,_u0_u29_ch_csr[28] , _u0_u29_ch_csr[27] , _u0_u29_ch_csr[26] ,_u0_u29_ch_csr[25] , _u0_u29_ch_csr[24] , _u0_u29_ch_csr[23] ,_u0_u29_ch_csr[22] , _u0_u29_ch_csr[21] , _u0_u29_ch_csr[20] ,_u0_u29_ch_csr[19] , _u0_u29_ch_csr[18] , _u0_u29_ch_csr[17] ,_u0_u29_ch_csr[16] , _u0_u29_ch_csr[15] , _u0_u29_ch_csr[14] ,_u0_u29_ch_csr[13] , _u0_u29_ch_csr[12] , _u0_u29_ch_csr[11] ,_u0_u29_ch_csr[10] , _u0_u29_ch_csr[9] , _u0_u29_ch_csr[8] ,_u0_u29_ch_csr[7] , _u0_u29_ch_csr[6] , _u0_u29_ch_csr[5] ,_u0_u29_ch_csr[4] , _u0_u29_ch_csr[3] , _u0_u29_ch_csr[2] ,_u0_u29_ch_csr[1] , _u0_u29_ch_csr[0] , _u0_u29_ch_txsz[31] ,_u0_u29_ch_txsz[30] , _u0_u29_ch_txsz[29] , _u0_u29_ch_txsz[28] ,_u0_u29_ch_txsz[27] , _u0_u29_ch_txsz[26] , _u0_u29_ch_txsz[25] ,_u0_u29_ch_txsz[24] , _u0_u29_ch_txsz[23] , _u0_u29_ch_txsz[22] ,_u0_u29_ch_txsz[21] , _u0_u29_ch_txsz[20] , _u0_u29_ch_txsz[19] ,_u0_u29_ch_txsz[18] , _u0_u29_ch_txsz[17] , _u0_u29_ch_txsz[16] ,_u0_u29_ch_txsz[15] , _u0_u29_ch_txsz[14] , _u0_u29_ch_txsz[13] ,_u0_u29_ch_txsz[12] , _u0_u29_ch_txsz[11] , _u0_u29_ch_txsz[10] ,_u0_u29_ch_txsz[9] , _u0_u29_ch_txsz[8] , _u0_u29_ch_txsz[7] ,_u0_u29_ch_txsz[6] , _u0_u29_ch_txsz[5] , _u0_u29_ch_txsz[4] ,_u0_u29_ch_txsz[3] , _u0_u29_ch_txsz[2] , _u0_u29_ch_txsz[1] ,_u0_u29_ch_txsz[0] , _u0_u29_ch_adr0[31] , _u0_u29_ch_adr0[30] ,_u0_u29_ch_adr0[29] , _u0_u29_ch_adr0[28] , _u0_u29_ch_adr0[27] ,_u0_u29_ch_adr0[26] , _u0_u29_ch_adr0[25] , _u0_u29_ch_adr0[24] ,_u0_u29_ch_adr0[23] , _u0_u29_ch_adr0[22] , _u0_u29_ch_adr0[21] ,_u0_u29_ch_adr0[20] , _u0_u29_ch_adr0[19] , _u0_u29_ch_adr0[18] ,_u0_u29_ch_adr0[17] , _u0_u29_ch_adr0[16] , _u0_u29_ch_adr0[15] ,_u0_u29_ch_adr0[14] , _u0_u29_ch_adr0[13] , _u0_u29_ch_adr0[12] ,_u0_u29_ch_adr0[11] , _u0_u29_ch_adr0[10] , _u0_u29_ch_adr0[9] ,_u0_u29_ch_adr0[8] , _u0_u29_ch_adr0[7] , _u0_u29_ch_adr0[6] ,_u0_u29_ch_adr0[5] , _u0_u29_ch_adr0[4] , _u0_u29_ch_adr0[3] ,_u0_u29_ch_adr0[2] , _u0_u29_ch_adr0[1] , _u0_u29_ch_adr0[0] ,_u0_u29_ch_adr1[31] , _u0_u29_ch_adr1[30] , _u0_u29_ch_adr1[29] ,_u0_u29_ch_adr1[28] , _u0_u29_ch_adr1[27] , _u0_u29_ch_adr1[26] ,_u0_u29_ch_adr1[25] , _u0_u29_ch_adr1[24] , _u0_u29_ch_adr1[23] ,_u0_u29_ch_adr1[22] , _u0_u29_ch_adr1[21] , _u0_u29_ch_adr1[20] ,_u0_u29_ch_adr1[19] , _u0_u29_ch_adr1[18] , _u0_u29_ch_adr1[17] ,_u0_u29_ch_adr1[16] , _u0_u29_ch_adr1[15] , _u0_u29_ch_adr1[14] ,_u0_u29_ch_adr1[13] , _u0_u29_ch_adr1[12] , _u0_u29_ch_adr1[11] ,_u0_u29_ch_adr1[10] , _u0_u29_ch_adr1[9] , _u0_u29_ch_adr1[8] ,_u0_u29_ch_adr1[7] , _u0_u29_ch_adr1[6] , _u0_u29_ch_adr1[5] ,_u0_u29_ch_adr1[4] , _u0_u29_ch_adr1[3] , _u0_u29_ch_adr1[2] ,_u0_u29_ch_adr1[1] , _u0_u29_ch_adr1[0] , _u0_u29_ch_am0[31] ,_u0_u29_ch_am0[30] , _u0_u29_ch_am0[29] , _u0_u29_ch_am0[28] ,_u0_u29_ch_am0[27] , _u0_u29_ch_am0[26] , _u0_u29_ch_am0[25] ,_u0_u29_ch_am0[24] , _u0_u29_ch_am0[23] , _u0_u29_ch_am0[22] ,_u0_u29_ch_am0[21] , _u0_u29_ch_am0[20] , _u0_u29_ch_am0[19] ,_u0_u29_ch_am0[18] , _u0_u29_ch_am0[17] , _u0_u29_ch_am0[16] ,_u0_u29_ch_am0[15] , _u0_u29_ch_am0[14] , _u0_u29_ch_am0[13] ,_u0_u29_ch_am0[12] , _u0_u29_ch_am0[11] , _u0_u29_ch_am0[10] ,_u0_u29_ch_am0[9] , _u0_u29_ch_am0[8] , _u0_u29_ch_am0[7] ,_u0_u29_ch_am0[6] , _u0_u29_ch_am0[5] , _u0_u29_ch_am0[4] ,_u0_u29_ch_am0[3] , _u0_u29_ch_am0[2] , _u0_u29_ch_am0[1] ,_u0_u29_ch_am0[0] , _u0_u29_ch_am1[31] , _u0_u29_ch_am1[30] ,_u0_u29_ch_am1[29] , _u0_u29_ch_am1[28] , _u0_u29_ch_am1[27] ,_u0_u29_ch_am1[26] , _u0_u29_ch_am1[25] , _u0_u29_ch_am1[24] ,_u0_u29_ch_am1[23] , _u0_u29_ch_am1[22] , _u0_u29_ch_am1[21] ,_u0_u29_ch_am1[20] , _u0_u29_ch_am1[19] , _u0_u29_ch_am1[18] ,_u0_u29_ch_am1[17] , _u0_u29_ch_am1[16] , _u0_u29_ch_am1[15] ,_u0_u29_ch_am1[14] , _u0_u29_ch_am1[13] , _u0_u29_ch_am1[12] ,_u0_u29_ch_am1[11] , _u0_u29_ch_am1[10] , _u0_u29_ch_am1[9] ,_u0_u29_ch_am1[8] , _u0_u29_ch_am1[7] , _u0_u29_ch_am1[6] ,_u0_u29_ch_am1[5] , _u0_u29_ch_am1[4] , _u0_u29_ch_am1[3] ,_u0_u29_ch_am1[2] , _u0_u29_ch_am1[1] , _u0_u29_ch_am1[0] ,_u0_u29_sw_pointer[31] , _u0_u29_sw_pointer[30] ,_u0_u29_sw_pointer[29] , _u0_u29_sw_pointer[28] ,_u0_u29_sw_pointer[27] , _u0_u29_sw_pointer[26] ,_u0_u29_sw_pointer[25] , _u0_u29_sw_pointer[24] ,_u0_u29_sw_pointer[23] , _u0_u29_sw_pointer[22] ,_u0_u29_sw_pointer[21] , _u0_u29_sw_pointer[20] ,_u0_u29_sw_pointer[19] , _u0_u29_sw_pointer[18] ,_u0_u29_sw_pointer[17] , _u0_u29_sw_pointer[16] ,_u0_u29_sw_pointer[15] , _u0_u29_sw_pointer[14] ,_u0_u29_sw_pointer[13] , _u0_u29_sw_pointer[12] ,_u0_u29_sw_pointer[11] , _u0_u29_sw_pointer[10] ,_u0_u29_sw_pointer[9] , _u0_u29_sw_pointer[8] ,_u0_u29_sw_pointer[7] , _u0_u29_sw_pointer[6] ,_u0_u29_sw_pointer[5] , _u0_u29_sw_pointer[4] ,_u0_u29_sw_pointer[3] , _u0_u29_sw_pointer[2] ,_u0_u29_sw_pointer[1] , _u0_u29_sw_pointer[0] , _u0_u29_ch_stop ,_u0_u29_ch_dis , _u0_u29_int , _u0_u30_pointer[31] ,_u0_u30_pointer[30] , _u0_u30_pointer[29] , _u0_u30_pointer[28] ,_u0_u30_pointer[27] , _u0_u30_pointer[26] , _u0_u30_pointer[25] ,_u0_u30_pointer[24] , _u0_u30_pointer[23] , _u0_u30_pointer[22] ,_u0_u30_pointer[21] , _u0_u30_pointer[20] , _u0_u30_pointer[19] ,_u0_u30_pointer[18] , _u0_u30_pointer[17] , _u0_u30_pointer[16] ,_u0_u30_pointer[15] , _u0_u30_pointer[14] , _u0_u30_pointer[13] ,_u0_u30_pointer[12] , _u0_u30_pointer[11] , _u0_u30_pointer[10] ,_u0_u30_pointer[9] , _u0_u30_pointer[8] , _u0_u30_pointer[7] ,_u0_u30_pointer[6] , _u0_u30_pointer[5] , _u0_u30_pointer[4] ,_u0_u30_pointer[3] , _u0_u30_pointer[2] , _u0_u30_pointer[1] ,_u0_u30_pointer[0] , _u0_u30_pointer_s[31] , _u0_u30_pointer_s[30] ,_u0_u30_pointer_s[29] , _u0_u30_pointer_s[28] ,_u0_u30_pointer_s[27] , _u0_u30_pointer_s[26] ,_u0_u30_pointer_s[25] , _u0_u30_pointer_s[24] ,_u0_u30_pointer_s[23] , _u0_u30_pointer_s[22] ,_u0_u30_pointer_s[21] , _u0_u30_pointer_s[20] ,_u0_u30_pointer_s[19] , _u0_u30_pointer_s[18] ,_u0_u30_pointer_s[17] , _u0_u30_pointer_s[16] ,_u0_u30_pointer_s[15] , _u0_u30_pointer_s[14] ,_u0_u30_pointer_s[13] , _u0_u30_pointer_s[12] ,_u0_u30_pointer_s[11] , _u0_u30_pointer_s[10] , _u0_u30_pointer_s[9] ,_u0_u30_pointer_s[8] , _u0_u30_pointer_s[7] , _u0_u30_pointer_s[6] ,_u0_u30_pointer_s[5] , _u0_u30_pointer_s[4] , _u0_u30_pointer_s[3] ,_u0_u30_pointer_s[2] , _u0_u30_pointer_s[1] , _u0_u30_pointer_s[0] ,_u0_u30_ch_csr[31] , _u0_u30_ch_csr[30] , _u0_u30_ch_csr[29] ,_u0_u30_ch_csr[28] , _u0_u30_ch_csr[27] , _u0_u30_ch_csr[26] ,_u0_u30_ch_csr[25] , _u0_u30_ch_csr[24] , _u0_u30_ch_csr[23] ,_u0_u30_ch_csr[22] , _u0_u30_ch_csr[21] , _u0_u30_ch_csr[20] ,_u0_u30_ch_csr[19] , _u0_u30_ch_csr[18] , _u0_u30_ch_csr[17] ,_u0_u30_ch_csr[16] , _u0_u30_ch_csr[15] , _u0_u30_ch_csr[14] ,_u0_u30_ch_csr[13] , _u0_u30_ch_csr[12] , _u0_u30_ch_csr[11] ,_u0_u30_ch_csr[10] , _u0_u30_ch_csr[9] , _u0_u30_ch_csr[8] ,_u0_u30_ch_csr[7] , _u0_u30_ch_csr[6] , _u0_u30_ch_csr[5] ,_u0_u30_ch_csr[4] , _u0_u30_ch_csr[3] , _u0_u30_ch_csr[2] ,_u0_u30_ch_csr[1] , _u0_u30_ch_csr[0] , _u0_u30_ch_txsz[31] ,_u0_u30_ch_txsz[30] , _u0_u30_ch_txsz[29] , _u0_u30_ch_txsz[28] ,_u0_u30_ch_txsz[27] , _u0_u30_ch_txsz[26] , _u0_u30_ch_txsz[25] ,_u0_u30_ch_txsz[24] , _u0_u30_ch_txsz[23] , _u0_u30_ch_txsz[22] ,_u0_u30_ch_txsz[21] , _u0_u30_ch_txsz[20] , _u0_u30_ch_txsz[19] ,_u0_u30_ch_txsz[18] , _u0_u30_ch_txsz[17] , _u0_u30_ch_txsz[16] ,_u0_u30_ch_txsz[15] , _u0_u30_ch_txsz[14] , _u0_u30_ch_txsz[13] ,_u0_u30_ch_txsz[12] , _u0_u30_ch_txsz[11] , _u0_u30_ch_txsz[10] ,_u0_u30_ch_txsz[9] , _u0_u30_ch_txsz[8] , _u0_u30_ch_txsz[7] ,_u0_u30_ch_txsz[6] , _u0_u30_ch_txsz[5] , _u0_u30_ch_txsz[4] ,_u0_u30_ch_txsz[3] , _u0_u30_ch_txsz[2] , _u0_u30_ch_txsz[1] ,_u0_u30_ch_txsz[0] , _u0_u30_ch_adr0[31] , _u0_u30_ch_adr0[30] ,_u0_u30_ch_adr0[29] , _u0_u30_ch_adr0[28] , _u0_u30_ch_adr0[27] ,_u0_u30_ch_adr0[26] , _u0_u30_ch_adr0[25] , _u0_u30_ch_adr0[24] ,_u0_u30_ch_adr0[23] , _u0_u30_ch_adr0[22] , _u0_u30_ch_adr0[21] ,_u0_u30_ch_adr0[20] , _u0_u30_ch_adr0[19] , _u0_u30_ch_adr0[18] ,_u0_u30_ch_adr0[17] , _u0_u30_ch_adr0[16] , _u0_u30_ch_adr0[15] ,_u0_u30_ch_adr0[14] , _u0_u30_ch_adr0[13] , _u0_u30_ch_adr0[12] ,_u0_u30_ch_adr0[11] , _u0_u30_ch_adr0[10] , _u0_u30_ch_adr0[9] ,_u0_u30_ch_adr0[8] , _u0_u30_ch_adr0[7] , _u0_u30_ch_adr0[6] ,_u0_u30_ch_adr0[5] , _u0_u30_ch_adr0[4] , _u0_u30_ch_adr0[3] ,_u0_u30_ch_adr0[2] , _u0_u30_ch_adr0[1] , _u0_u30_ch_adr0[0] ,_u0_u30_ch_adr1[31] , _u0_u30_ch_adr1[30] , _u0_u30_ch_adr1[29] ,_u0_u30_ch_adr1[28] , _u0_u30_ch_adr1[27] , _u0_u30_ch_adr1[26] ,_u0_u30_ch_adr1[25] , _u0_u30_ch_adr1[24] , _u0_u30_ch_adr1[23] ,_u0_u30_ch_adr1[22] , _u0_u30_ch_adr1[21] , _u0_u30_ch_adr1[20] ,_u0_u30_ch_adr1[19] , _u0_u30_ch_adr1[18] , _u0_u30_ch_adr1[17] ,_u0_u30_ch_adr1[16] , _u0_u30_ch_adr1[15] , _u0_u30_ch_adr1[14] ,_u0_u30_ch_adr1[13] , _u0_u30_ch_adr1[12] , _u0_u30_ch_adr1[11] ,_u0_u30_ch_adr1[10] , _u0_u30_ch_adr1[9] , _u0_u30_ch_adr1[8] ,_u0_u30_ch_adr1[7] , _u0_u30_ch_adr1[6] , _u0_u30_ch_adr1[5] ,_u0_u30_ch_adr1[4] , _u0_u30_ch_adr1[3] , _u0_u30_ch_adr1[2] ,_u0_u30_ch_adr1[1] , _u0_u30_ch_adr1[0] , _u0_u30_ch_am0[31] ,_u0_u30_ch_am0[30] , _u0_u30_ch_am0[29] , _u0_u30_ch_am0[28] ,_u0_u30_ch_am0[27] , _u0_u30_ch_am0[26] , _u0_u30_ch_am0[25] ,_u0_u30_ch_am0[24] , _u0_u30_ch_am0[23] , _u0_u30_ch_am0[22] ,_u0_u30_ch_am0[21] , _u0_u30_ch_am0[20] , _u0_u30_ch_am0[19] ,_u0_u30_ch_am0[18] , _u0_u30_ch_am0[17] , _u0_u30_ch_am0[16] ,_u0_u30_ch_am0[15] , _u0_u30_ch_am0[14] , _u0_u30_ch_am0[13] ,_u0_u30_ch_am0[12] , _u0_u30_ch_am0[11] , _u0_u30_ch_am0[10] ,_u0_u30_ch_am0[9] , _u0_u30_ch_am0[8] , _u0_u30_ch_am0[7] ,_u0_u30_ch_am0[6] , _u0_u30_ch_am0[5] , _u0_u30_ch_am0[4] ,_u0_u30_ch_am0[3] , _u0_u30_ch_am0[2] , _u0_u30_ch_am0[1] ,_u0_u30_ch_am0[0] , _u0_u30_ch_am1[31] , _u0_u30_ch_am1[30] ,_u0_u30_ch_am1[29] , _u0_u30_ch_am1[28] , _u0_u30_ch_am1[27] ,_u0_u30_ch_am1[26] , _u0_u30_ch_am1[25] , _u0_u30_ch_am1[24] ,_u0_u30_ch_am1[23] , _u0_u30_ch_am1[22] , _u0_u30_ch_am1[21] ,_u0_u30_ch_am1[20] , _u0_u30_ch_am1[19] , _u0_u30_ch_am1[18] ,_u0_u30_ch_am1[17] , _u0_u30_ch_am1[16] , _u0_u30_ch_am1[15] ,_u0_u30_ch_am1[14] , _u0_u30_ch_am1[13] , _u0_u30_ch_am1[12] ,_u0_u30_ch_am1[11] , _u0_u30_ch_am1[10] , _u0_u30_ch_am1[9] ,_u0_u30_ch_am1[8] , _u0_u30_ch_am1[7] , _u0_u30_ch_am1[6] ,_u0_u30_ch_am1[5] , _u0_u30_ch_am1[4] , _u0_u30_ch_am1[3] ,_u0_u30_ch_am1[2] , _u0_u30_ch_am1[1] , _u0_u30_ch_am1[0] ,_u0_u30_sw_pointer[31] , _u0_u30_sw_pointer[30] ,_u0_u30_sw_pointer[29] , _u0_u30_sw_pointer[28] ,_u0_u30_sw_pointer[27] , _u0_u30_sw_pointer[26] ,_u0_u30_sw_pointer[25] , _u0_u30_sw_pointer[24] ,_u0_u30_sw_pointer[23] , _u0_u30_sw_pointer[22] ,_u0_u30_sw_pointer[21] , _u0_u30_sw_pointer[20] ,_u0_u30_sw_pointer[19] , _u0_u30_sw_pointer[18] ,_u0_u30_sw_pointer[17] , _u0_u30_sw_pointer[16] ,_u0_u30_sw_pointer[15] , _u0_u30_sw_pointer[14] ,_u0_u30_sw_pointer[13] , _u0_u30_sw_pointer[12] ,_u0_u30_sw_pointer[11] , _u0_u30_sw_pointer[10] ,_u0_u30_sw_pointer[9] , _u0_u30_sw_pointer[8] ,_u0_u30_sw_pointer[7] , _u0_u30_sw_pointer[6] ,_u0_u30_sw_pointer[5] , _u0_u30_sw_pointer[4] ,_u0_u30_sw_pointer[3] , _u0_u30_sw_pointer[2] ,_u0_u30_sw_pointer[1] , _u0_u30_sw_pointer[0] , _u0_u30_ch_stop ,_u0_u30_ch_dis , _u0_u30_int , _u10_SYNOPSYS_UNCONNECTED_38 ,_u10_SYNOPSYS_UNCONNECTED_37 , _u10_SYNOPSYS_UNCONNECTED_36 ,_u10_SYNOPSYS_UNCONNECTED_35 , _u10_SYNOPSYS_UNCONNECTED_34 ,_u10_SYNOPSYS_UNCONNECTED_33 , _u10_SYNOPSYS_UNCONNECTED_32 ,_u10_SYNOPSYS_UNCONNECTED_31 , _u10_SYNOPSYS_UNCONNECTED_30 ,_u10_SYNOPSYS_UNCONNECTED_29 , _u10_SYNOPSYS_UNCONNECTED_28 ,_u10_SYNOPSYS_UNCONNECTED_27 , _u10_SYNOPSYS_UNCONNECTED_26 ,_u10_SYNOPSYS_UNCONNECTED_25 , _u10_SYNOPSYS_UNCONNECTED_24 ,_u10_SYNOPSYS_UNCONNECTED_23 , _u10_SYNOPSYS_UNCONNECTED_22 ,_u10_SYNOPSYS_UNCONNECTED_21 , _u10_SYNOPSYS_UNCONNECTED_20 ,_u10_SYNOPSYS_UNCONNECTED_19 , _u10_SYNOPSYS_UNCONNECTED_18 ,_u10_SYNOPSYS_UNCONNECTED_17 , _u10_SYNOPSYS_UNCONNECTED_16 ,_u10_SYNOPSYS_UNCONNECTED_15 , _u10_SYNOPSYS_UNCONNECTED_14 ,_u10_SYNOPSYS_UNCONNECTED_13 , _u10_SYNOPSYS_UNCONNECTED_12 ,_u10_SYNOPSYS_UNCONNECTED_11 , _u10_SYNOPSYS_UNCONNECTED_10 ,_u10_SYNOPSYS_UNCONNECTED_9 , _u10_SYNOPSYS_UNCONNECTED_8 ,_u10_SYNOPSYS_UNCONNECTED_7 , _u10_SYNOPSYS_UNCONNECTED_6 ,_u10_SYNOPSYS_UNCONNECTED_5 , _u10_SYNOPSYS_UNCONNECTED_4 ,_u10_n23001 , _u10_n23000 , _u10_n22999 , _u10_n22998 , _u10_n22997 ,_u10_n22996 , _u10_n22995 , _u10_n22994 , _u10_n22993 , _u10_n22992 ,_u10_n22991 , _u10_n22990 , _u10_n22989 , _u10_n22988 , _u10_n22987 ,_u10_n22986 , _u10_n22985 , _u10_n22984 , _u10_n22983 , _u10_n22982 ,_u10_n22981 , _u10_n22980 , _u10_n22979 , _u10_n22978 , _u10_n22977 ,_u10_n22976 , _u10_n22975 , _u10_n22974 , _u10_n22973 , _u10_n22972 ,_u10_n22971 , _u10_n22970 , _u10_n22969 , _u10_n22968 , _u10_n22967 ,_u10_n22966 , _u10_n22965 , _u10_n22964 , _u10_n22963 , _u10_n22962 ,_u10_n22961 , _u10_n22960 , _u10_n22959 , _u10_n22958 , _u10_n22957 ,_u10_n22956 , _u10_n22955 , _u10_n22954 , _u10_n22953 , _u10_n22952 ,_u10_n22951 , _u10_n22950 , _u10_n22949 , _u10_n22948 , _u10_n22947 ,_u10_n22946 , _u10_n22945 , _u10_n22944 , _u10_n22943 , _u10_n22942 ,_u10_n22941 , _u10_n22940 , _u10_n22939 , _u10_n22938 , _u10_n22937 ,_u10_n22936 , _u10_n22935 , _u10_n22934 , _u10_n22933 , _u10_n22932 ,_u10_n22931 , _u10_n22930 , _u10_n22929 , _u10_n22928 , _u10_n22927 ,_u10_n22926 , _u10_n22925 , _u10_n22924 , _u10_n22923 , _u10_n22922 ,_u10_n22921 , _u10_n22920 , _u10_n22919 , _u10_n22918 , _u10_n22917 ,_u10_n22916 , _u10_n22915 , _u10_n22914 , _u10_n22913 , _u10_n22912 ,_u10_n22911 , _u10_n22910 , _u10_n22909 , _u10_n22908 , _u10_n22907 ,_u10_n22906 , _u10_n22905 , _u10_n22904 , _u10_n22903 , _u10_n22902 ,_u10_n22901 , _u10_n22900 , _u10_n22899 , _u10_n22898 , _u10_n22897 ,_u10_n22896 , _u10_n22895 , _u10_n22894 , _u10_n22893 , _u10_n22892 ,_u10_n22891 , _u10_n22890 , _u10_n22889 , _u10_n22888 , _u10_n22887 ,_u10_n22886 , _u10_n22885 , _u10_n22884 , _u10_n22883 , _u10_n22882 ,_u10_n22881 , _u10_n22880 , _u10_n22879 , _u10_n22878 , _u10_n22877 ,_u10_n22876 , _u10_n22875 , _u10_n22874 , _u10_n22873 , _u10_n22872 ,_u10_n22871 , _u10_n22870 , _u10_n22869 , _u10_n22868 , _u10_n22867 ,_u10_n22866 , _u10_n22865 , _u10_n22864 , _u10_n22863 , _u10_n22862 ,_u10_n22861 , _u10_n22860 , _u10_n22859 , _u10_n22858 , _u10_n22857 ,_u10_n22856 , _u10_n22855 , _u10_n22854 , _u10_n22853 , _u10_n22852 ,_u10_n22851 , _u10_n22850 , _u10_n22849 , _u10_n22848 , _u10_n22847 ,_u10_n22846 , _u10_n22845 , _u10_n22844 , _u10_n22843 , _u10_n22842 ,_u10_n22841 , _u10_n22840 , _u10_n22839 , _u10_n22838 , _u10_n22837 ,_u10_n22836 , _u10_n22835 , _u10_n22834 , _u10_n22833 , _u10_n22832 ,_u10_n22831 , _u10_n22830 , _u10_n22829 , _u10_n22828 , _u10_n22827 ,_u10_n22826 , _u10_n22825 , _u10_n22824 , _u10_n22823 , _u10_n22822 ,_u10_n22821 , _u10_n22820 , _u10_n22819 , _u10_n22818 , _u10_n22817 ,_u10_n22816 , _u10_n22815 , _u10_n22814 , _u10_n22813 , _u10_n22812 ,_u10_n22811 , _u10_n22810 , _u10_n22809 , _u10_n22808 , _u10_n22807 ,_u10_n22806 , _u10_n22805 , _u10_n22804 , _u10_n22803 , _u10_n22802 ,_u10_n22801 , _u10_n22800 , _u10_n22799 , _u10_n22798 , _u10_n22797 ,_u10_n22796 , _u10_n22795 , _u10_n22794 , _u10_n22793 , _u10_n22792 ,_u10_n22791 , _u10_n22790 , _u10_n22789 , _u10_n22788 , _u10_n22787 ,_u10_n22786 , _u10_n22785 , _u10_n22784 , _u10_n22783 , _u10_n22782 ,_u10_n22781 , _u10_n22780 , _u10_n22779 , _u10_n22778 , _u10_n22777 ,_u10_n22776 , _u10_n22775 , _u10_n22774 , _u10_n22773 , _u10_n22772 ,_u10_n22771 , _u10_n22770 , _u10_n22769 , _u10_n22768 , _u10_n22767 ,_u10_n22766 , _u10_n22765 , _u10_n22764 , _u10_n22763 , _u10_n22762 ,_u10_n22761 , _u10_n22760 , _u10_n22759 , _u10_n22758 , _u10_n22757 ,_u10_n22756 , _u10_n22755 , _u10_n22754 , _u10_n22753 , _u10_n22752 ,_u10_n22751 , _u10_n22750 , _u10_n22749 , _u10_n22748 , _u10_n22747 ,_u10_n22746 , _u10_n22745 , _u10_n22744 , _u10_n22743 , _u10_n22742 ,_u10_n22741 , _u10_n22740 , _u10_n22739 , _u10_n22738 , _u10_n22737 ,_u10_n22736 , _u10_n22735 , _u10_n22734 , _u10_n22733 , _u10_n22732 ,_u10_n22731 , _u10_n22730 , _u10_n22729 , _u10_n22728 , _u10_n22727 ,_u10_n22726 , _u10_n22725 , _u10_n22724 , _u10_n22723 , _u10_n22722 ,_u10_n22721 , _u10_n22720 , _u10_n22719 , _u10_n22718 , _u10_n22717 ,_u10_n22716 , _u10_n22715 , _u10_n22714 , _u10_n22713 , _u10_n22712 ,_u10_n22711 , _u10_n22710 , _u10_n22709 , _u10_n22708 , _u10_n22707 ,_u10_n22706 , _u10_n22705 , _u10_n22704 , _u10_n22703 , _u10_n22702 ,_u10_n22701 , _u10_n22700 , _u10_n22699 , _u10_n22698 , _u10_n22697 ,_u10_n22696 , _u10_n22695 , _u10_n22694 , _u10_n22693 , _u10_n22692 ,_u10_n22691 , _u10_n22690 , _u10_n22689 , _u10_n22688 , _u10_n22687 ,_u10_n22686 , _u10_n22685 , _u10_n22684 , _u10_n22683 , _u10_n22682 ,_u10_n22681 , _u10_n22680 , _u10_n22679 , _u10_n22678 , _u10_n22677 ,_u10_n22676 , _u10_n22675 , _u10_n22674 , _u10_n22673 , _u10_n22672 ,_u10_n22671 , _u10_n22670 , _u10_n22669 , _u10_n22668 , _u10_n22667 ,_u10_n22666 , _u10_n22665 , _u10_n22664 , _u10_n22663 , _u10_n22662 ,_u10_n22661 , _u10_n22660 , _u10_n22659 , _u10_n22658 , _u10_n22657 ,_u10_n22656 , _u10_n22655 , _u10_n22654 , _u10_n22653 , _u10_n22652 ,_u10_n22651 , _u10_n22650 , _u10_n22649 , _u10_n22648 , _u10_n22647 ,_u10_n22646 , _u10_n22645 , _u10_n22644 , _u10_n22643 , _u10_n22642 ,_u10_n22641 , _u10_n22640 , _u10_n22639 , _u10_n22638 , _u10_n22637 ,_u10_n22636 , _u10_n22635 , _u10_n22634 , _u10_n22633 , _u10_n22632 ,_u10_n22631 , _u10_n22630 , _u10_n22629 , _u10_n22628 , _u10_n22627 ,_u10_n22626 , _u10_n22625 , _u10_n22624 , _u10_n22623 , _u10_n22622 ,_u10_n22621 , _u10_n22620 , _u10_n22619 , _u10_n22618 , _u10_n22617 ,_u10_n22616 , _u10_n22615 , _u10_n22614 , _u10_n22613 , _u10_n22612 ,_u10_n22611 , _u10_n22610 , _u10_n22609 , _u10_n22608 , _u10_n22607 ,_u10_n22606 , _u10_n22605 , _u10_n22604 , _u10_n22603 , _u10_n22602 ,_u10_n22601 , _u10_n22600 , _u10_n22599 , _u10_n22598 , _u10_n22597 ,_u10_n22596 , _u10_n22595 , _u10_n22594 , _u10_n22593 , _u10_n22592 ,_u10_n22591 , _u10_n22590 , _u10_n22589 , _u10_n22588 , _u10_n22587 ,_u10_n22586 , _u10_n22585 , _u10_n22584 , _u10_n22583 , _u10_n22582 ,_u10_n22581 , _u10_n22580 , _u10_n22579 , _u10_n22578 , _u10_n22577 ,_u10_n22576 , _u10_n22575 , _u10_n22574 , _u10_n22573 , _u10_n22572 ,_u10_n22571 , _u10_n22570 , _u10_n22569 , _u10_n22568 , _u10_n22567 ,_u10_n22566 , _u10_n22565 , _u10_n22564 , _u10_n22563 , _u10_n22562 ,_u10_n22561 , _u10_n22560 , _u10_n22559 , _u10_n22558 , _u10_n22557 ,_u10_n22556 , _u10_n22555 , _u10_n22554 , _u10_n22553 , _u10_n22552 ,_u10_n22551 , _u10_n22550 , _u10_n22549 , _u10_n22548 , _u10_n22547 ,_u10_n22546 , _u10_n22545 , _u10_n22544 , _u10_n22543 , _u10_n22542 ,_u10_n22541 , _u10_n22540 , _u10_n22539 , _u10_n22538 , _u10_n22537 ,_u10_n22536 , _u10_n22535 , _u10_n22534 , _u10_n22533 , _u10_n22532 ,_u10_n22531 , _u10_n22530 , _u10_n22529 , _u10_n22528 , _u10_n22527 ,_u10_n22526 , _u10_n22525 , _u10_n22524 , _u10_n22523 , _u10_n22522 ,_u10_n22521 , _u10_n22520 , _u10_n22519 , _u10_n22518 , _u10_n22517 ,_u10_n22516 , _u10_n22515 , _u10_n22514 , _u10_n22513 , _u10_n22512 ,_u10_n22511 , _u10_n22510 , _u10_n22509 , _u10_n22508 , _u10_n22507 ,_u10_n22506 , _u10_n22505 , _u10_n22504 , _u10_n22503 , _u10_n22502 ,_u10_n22501 , _u10_n22500 , _u10_n22499 , _u10_n22498 , _u10_n22497 ,_u10_n22496 , _u10_n22495 , _u10_n22494 , _u10_n22493 , _u10_n22492 ,_u10_n22491 , _u10_n22490 , _u10_n22489 , _u10_n22488 , _u10_n22487 ,_u10_n22486 , _u10_n22485 , _u10_n22484 , _u10_n22483 , _u10_n22482 ,_u10_n22481 , _u10_n22480 , _u10_n22479 , _u10_n22478 , _u10_n22477 ,_u10_n22476 , _u10_n22475 , _u10_n22474 , _u10_n22473 , _u10_n22472 ,_u10_n22471 , _u10_n22470 , _u10_n22469 , _u10_n22468 , _u10_n22467 ,_u10_n22466 , _u10_n22465 , _u10_n22464 , _u10_n22463 , _u10_n22462 ,_u10_n22461 , _u10_n22460 , _u10_n22459 , _u10_n22458 , _u10_n22457 ,_u10_n22456 , _u10_n22455 , _u10_n22454 , _u10_n22453 , _u10_n22452 ,_u10_n22451 , _u10_n22450 , _u10_n22449 , _u10_n22448 , _u10_n22447 ,_u10_n22446 , _u10_n22445 , _u10_n22444 , _u10_n22443 , _u10_n22442 ,_u10_n22441 , _u10_n22440 , _u10_n22439 , _u10_n22438 , _u10_n22437 ,_u10_n22436 , _u10_n22435 , _u10_n22434 , _u10_n22433 , _u10_n22432 ,_u10_n22431 , _u10_n22430 , _u10_n22429 , _u10_n22428 , _u10_n22427 ,_u10_n22426 , _u10_n22425 , _u10_n22424 , _u10_n22423 , _u10_n22422 ,_u10_n22421 , _u10_n22420 , _u10_n22419 , _u10_n22418 , _u10_n22417 ,_u10_n22416 , _u10_n22415 , _u10_n22414 , _u10_n22413 , _u10_n22412 ,_u10_n22411 , _u10_n22410 , _u10_n22409 , _u10_n22408 , _u10_n22407 ,_u10_n22406 , _u10_n22405 , _u10_n22404 , _u10_n22403 , _u10_n22402 ,_u10_n22401 , _u10_n22400 , _u10_n22399 , _u10_n22398 , _u10_n22397 ,_u10_n22396 , _u10_n22395 , _u10_n22394 , _u10_n22393 , _u10_n22392 ,_u10_n22391 , _u10_n22390 , _u10_n22389 , _u10_n22388 , _u10_n22387 ,_u10_n22386 , _u10_n22385 , _u10_n22384 , _u10_n22383 , _u10_n22382 ,_u10_n22381 , _u10_n22380 , _u10_n22379 , _u10_n22378 , _u10_n22377 ,_u10_n22376 , _u10_n22375 , _u10_n22374 , _u10_n22373 , _u10_n22372 ,_u10_n22371 , _u10_n22370 , _u10_n22369 , _u10_n22368 , _u10_n22367 ,_u10_n22366 , _u10_n22365 , _u10_n22364 , _u10_n22363 , _u10_n22362 ,_u10_n22361 , _u10_n22360 , _u10_n22359 , _u10_n22358 , _u10_n22357 ,_u10_n22356 , _u10_n22355 , _u10_n22354 , _u10_n22353 , _u10_n22352 ,_u10_n22351 , _u10_n22350 , _u10_n22349 , _u10_n22348 , _u10_n22347 ,_u10_n22346 , _u10_n22345 , _u10_n22344 , _u10_n22343 , _u10_n22342 ,_u10_n22341 , _u10_n22340 , _u10_n22339 , _u10_n22338 , _u10_n22337 ,_u10_n22336 , _u10_n22335 , _u10_n22334 , _u10_n22333 , _u10_n22332 ,_u10_n22331 , _u10_n22330 , _u10_n22329 , _u10_n22328 , _u10_n22327 ,_u10_n22326 , _u10_n22325 , _u10_n22324 , _u10_n22323 , _u10_n22322 ,_u10_n22321 , _u10_n22320 , _u10_n22319 , _u10_n22318 , _u10_n22317 ,_u10_n22316 , _u10_n22315 , _u10_n22314 , _u10_n22313 , _u10_n22312 ,_u10_n22311 , _u10_n22310 , _u10_n22309 , _u10_n22308 , _u10_n22307 ,_u10_n22306 , _u10_n22305 , _u10_n22304 , _u10_n22303 , _u10_n22302 ,_u10_n22301 , _u10_n22300 , _u10_n22299 , _u10_n22298 , _u10_n22297 ,_u10_n22296 , _u10_n22295 , _u10_n22294 , _u10_n22293 , _u10_n22292 ,_u10_n22291 , _u10_n22290 , _u10_n22289 , _u10_n22288 , _u10_n22287 ,_u10_n22286 , _u10_n22285 , _u10_n22284 , _u10_n22283 , _u10_n22282 ,_u10_n22281 , _u10_n22280 , _u10_n22279 , _u10_n22278 , _u10_n22277 ,_u10_n22276 , _u10_n22275 , _u10_n22274 , _u10_n22273 , _u10_n22272 ,_u10_n22271 , _u10_n22270 , _u10_n22269 , _u10_n22268 , _u10_n22267 ,_u10_n22266 , _u10_n22265 , _u10_n22264 , _u10_n22263 , _u10_n22262 ,_u10_n22261 , _u10_n22260 , _u10_n22259 , _u10_n22258 , _u10_n22257 ,_u10_n22256 , _u10_n22255 , _u10_n22254 , _u10_n22253 , _u10_n22252 ,_u10_n22251 , _u10_n22250 , _u10_n22249 , _u10_n22248 , _u10_n22247 ,_u10_n22246 , _u10_n22245 , _u10_n22244 , _u10_n22243 , _u10_n22242 ,_u10_n22241 , _u10_n22240 , _u10_n22239 , _u10_n22238 , _u10_n22237 ,_u10_n22236 , _u10_n22235 , _u10_n22234 , _u10_n22233 , _u10_n22232 ,_u10_n22231 , _u10_n22230 , _u10_n22229 , _u10_n22228 , _u10_n22227 ,_u10_n22226 , _u10_n22225 , _u10_n22224 , _u10_n22223 , _u10_n22222 ,_u10_n22221 , _u10_n22220 , _u10_n22219 , _u10_n22218 , _u10_n22217 ,_u10_n22216 , _u10_n22215 , _u10_n22214 , _u10_n22213 , _u10_n22212 ,_u10_n22211 , _u10_n22210 , _u10_n22209 , _u10_n22208 , _u10_n22207 ,_u10_n22206 , _u10_n22205 , _u10_n22204 , _u10_n22203 , _u10_n22202 ,_u10_n22201 , _u10_n22200 , _u10_n22199 , _u10_n22198 , _u10_n22197 ,_u10_n22196 , _u10_n22195 , _u10_n22194 , _u10_n22193 , _u10_n22192 ,_u10_n22191 , _u10_n22190 , _u10_n22189 , _u10_n22188 , _u10_n22187 ,_u10_n22186 , _u10_n22185 , _u10_n22184 , _u10_n22183 , _u10_n22182 ,_u10_n22181 , _u10_n22180 , _u10_n22179 , _u10_n22178 , _u10_n22177 ,_u10_n22176 , _u10_n22175 , _u10_n22174 , _u10_n22173 , _u10_n22172 ,_u10_n22171 , _u10_n22170 , _u10_n22169 , _u10_n22168 , _u10_n22167 ,_u10_n22166 , _u10_n22165 , _u10_n22164 , _u10_n22163 , _u10_n22162 ,_u10_n22161 , _u10_n22160 , _u10_n22159 , _u10_n22158 , _u10_n22157 ,_u10_n22156 , _u10_n22155 , _u10_n22154 , _u10_n22153 , _u10_n22152 ,_u10_n22151 , _u10_n22150 , _u10_n22149 , _u10_n22148 , _u10_n22147 ,_u10_n22146 , _u10_n22145 , _u10_n22144 , _u10_n22143 , _u10_n22142 ,_u10_n22141 , _u10_n22140 , _u10_n22139 , _u10_n22138 , _u10_n22137 ,_u10_n22136 , _u10_n22135 , _u10_n22134 , _u10_n22133 , _u10_n22132 ,_u10_n22131 , _u10_n22130 , _u10_n22129 , _u10_n22128 , _u10_n22127 ,_u10_n22126 , _u10_n22125 , _u10_n22124 , _u10_n22123 , _u10_n22122 ,_u10_n22121 , _u10_n22120 , _u10_n22119 , _u10_n22118 , _u10_n22117 ,_u10_n22116 , _u10_n22115 , _u10_n22114 , _u10_n22113 , _u10_n22112 ,_u10_n22111 , _u10_n22110 , _u10_n22109 , _u10_n22108 , _u10_n22107 ,_u10_n22106 , _u10_n22105 , _u10_n22104 , _u10_n22103 , _u10_n22102 ,_u10_n22101 , _u10_n22100 , _u10_n22099 , _u10_n22098 , _u10_n22097 ,_u10_n22096 , _u10_n22095 , _u10_n22094 , _u10_n22093 , _u10_n22092 ,_u10_n22091 , _u10_n22090 , _u10_n22089 , _u10_n22088 , _u10_n22087 ,_u10_n22086 , _u10_n22085 , _u10_n22084 , _u10_n22083 , _u10_n22082 ,_u10_n22081 , _u10_n22080 , _u10_n22079 , _u10_n22078 , _u10_n22077 ,_u10_n22076 , _u10_n22075 , _u10_n22074 , _u10_n22073 , _u10_n22072 ,_u10_n22071 , _u10_n22070 , _u10_n22069 , _u10_n22068 , _u10_n22067 ,_u10_n22066 , _u10_n22065 , _u10_n22064 , _u10_n22063 , _u10_n22062 ,_u10_n22061 , _u10_n22060 , _u10_n22059 , _u10_n22058 , _u10_n22057 ,_u10_n22056 , _u10_n22055 , _u10_n22054 , _u10_n22053 , _u10_n22052 ,_u10_n22051 , _u10_n22050 , _u10_n22049 , _u10_n22048 , _u10_n22047 ,_u10_n22046 , _u10_n22045 , _u10_n22044 , _u10_n22043 , _u10_n22042 ,_u10_n22041 , _u10_n22040 , _u10_n22039 , _u10_n22038 , _u10_n22037 ,_u10_n22036 , _u10_n22035 , _u10_n22034 , _u10_n22033 , _u10_n22032 ,_u10_n22031 , _u10_n22030 , _u10_n22029 , _u10_n22028 , _u10_n22027 ,_u10_n22026 , _u10_n22025 , _u10_n22024 , _u10_n22023 , _u10_n22022 ,_u10_n22021 , _u10_n22020 , _u10_n22019 , _u10_n22018 , _u10_n22017 ,_u10_n22016 , _u10_n22015 , _u10_n22014 , _u10_n22013 , _u10_n22012 ,_u10_n22011 , _u10_n22010 , _u10_n22009 , _u10_n22008 , _u10_n22007 ,_u10_n22006 , _u10_n22005 , _u10_n22004 , _u10_n22003 , _u10_n22002 ,_u10_n22001 , _u10_n22000 , _u10_n21999 , _u10_n21998 , _u10_n21997 ,_u10_n21996 , _u10_n21995 , _u10_n21994 , _u10_n21993 , _u10_n21992 ,_u10_n21991 , _u10_n21990 , _u10_n21989 , _u10_n21988 , _u10_n21987 ,_u10_n21986 , _u10_n21985 , _u10_n21984 , _u10_n21983 , _u10_n21982 ,_u10_n21981 , _u10_n21980 , _u10_n21979 , _u10_n21978 , _u10_n21977 ,_u10_n21976 , _u10_n21975 , _u10_n21974 , _u10_n21973 , _u10_n21972 ,_u10_n21971 , _u10_n21970 , _u10_n21969 , _u10_n21968 , _u10_n21967 ,_u10_n21966 , _u10_n21965 , _u10_n21964 , _u10_n21963 , _u10_n21962 ,_u10_n21961 , _u10_n21960 , _u10_n21959 , _u10_n21958 , _u10_n21957 ,_u10_n21956 , _u10_n21955 , _u10_n21954 , _u10_n21953 , _u10_n21952 ,_u10_n21951 , _u10_n21950 , _u10_n21949 , _u10_n21948 , _u10_n21947 ,_u10_n21946 , _u10_n21945 , _u10_n21944 , _u10_n21943 , _u10_n21942 ,_u10_n21941 , _u10_n21940 , _u10_n21939 , _u10_n21938 , _u10_n21937 ,_u10_n21936 , _u10_n21935 , _u10_n21934 , _u10_n21933 , _u10_n21932 ,_u10_n21931 , _u10_n21930 , _u10_n21929 , _u10_n21928 , _u10_n21927 ,_u10_n21926 , _u10_n21925 , _u10_n21924 , _u10_n21923 , _u10_n21922 ,_u10_n21921 , _u10_n21920 , _u10_n21919 , _u10_n21918 , _u10_n21917 ,_u10_n21916 , _u10_n21915 , _u10_n21914 , _u10_n21913 , _u10_n21912 ,_u10_n21911 , _u10_n21910 , _u10_n21909 , _u10_n21908 , _u10_n21907 ,_u10_n21906 , _u10_n21905 , _u10_n21904 , _u10_n21903 , _u10_n21902 ,_u10_n21901 , _u10_n21900 , _u10_n21899 , _u10_n21898 , _u10_n21897 ,_u10_n21896 , _u10_n21895 , _u10_n21894 , _u10_n21893 , _u10_n21892 ,_u10_n21891 , _u10_n21890 , _u10_n21889 , _u10_n21888 , _u10_n21887 ,_u10_n21886 , _u10_n21885 , _u10_n21884 , _u10_n21883 , _u10_n21882 ,_u10_n21881 , _u10_n21880 , _u10_n21879 , _u10_n21878 , _u10_n21877 ,_u10_n21876 , _u10_n21875 , _u10_n21874 , _u10_n21873 , _u10_n21872 ,_u10_n21871 , _u10_n21870 , _u10_n21869 , _u10_n21868 , _u10_n21867 ,_u10_n21866 , _u10_n21865 , _u10_n21864 , _u10_n21863 , _u10_n21862 ,_u10_n21861 , _u10_n21860 , _u10_n21859 , _u10_n21858 , _u10_n21857 ,_u10_n21856 , _u10_n21855 , _u10_n21854 , _u10_n21853 , _u10_n21852 ,_u10_n21851 , _u10_n21850 , _u10_n21849 , _u10_n21848 , _u10_n21847 ,_u10_n21846 , _u10_n21845 , _u10_n21844 , _u10_n21843 , _u10_n21842 ,_u10_n21841 , _u10_n21840 , _u10_n21839 , _u10_n21838 , _u10_n21837 ,_u10_n21836 , _u10_n21835 , _u10_n21834 , _u10_n21833 , _u10_n21832 ,_u10_n21831 , _u10_n21830 , _u10_n21829 , _u10_n21828 , _u10_n21827 ,_u10_n21826 , _u10_n21825 , _u10_n21824 , _u10_n21823 , _u10_n21822 ,_u10_n21821 , _u10_n21820 , _u10_n21819 , _u10_n21818 , _u10_n21817 ,_u10_n21816 , _u10_n21815 , _u10_n21814 , _u10_n21813 , _u10_n21812 ,_u10_n21811 , _u10_n21810 , _u10_n21809 , _u10_n21808 , _u10_n21807 ,_u10_n21806 , _u10_n21805 , _u10_n21804 , _u10_n21803 , _u10_n21802 ,_u10_n21801 , _u10_n21800 , _u10_n21799 , _u10_n21798 , _u10_n21797 ,_u10_n21796 , _u10_n21795 , _u10_n21794 , _u10_n21793 , _u10_n21792 ,_u10_n21791 , _u10_n21790 , _u10_n21789 , _u10_n21788 , _u10_n21787 ,_u10_n21786 , _u10_n21785 , _u10_n21784 , _u10_n21783 , _u10_n21782 ,_u10_n21781 , _u10_n21780 , _u10_n21779 , _u10_n21778 , _u10_n21777 ,_u10_n21776 , _u10_n21775 , _u10_n21774 , _u10_n21773 , _u10_n21772 ,_u10_n21771 , _u10_n21770 , _u10_n21769 , _u10_n21768 , _u10_n21767 ,_u10_n21766 , _u10_n21765 , _u10_n21764 , _u10_n21763 , _u10_n21762 ,_u10_n21761 , _u10_n21760 , _u10_n21759 , _u10_n21758 , _u10_n21757 ,_u10_n21756 , _u10_n21755 , _u10_n21754 , _u10_n21753 , _u10_n21752 ,_u10_n21751 , _u10_n21750 , _u10_n21749 , _u10_n21748 , _u10_n21747 ,_u10_n21746 , _u10_n21745 , _u10_n21744 , _u10_n21743 , _u10_n21742 ,_u10_n21741 , _u10_n21740 , _u10_n21739 , _u10_n21738 , _u10_n21737 ,_u10_n21736 , _u10_n21735 , _u10_n21734 , _u10_n21733 , _u10_n21732 ,_u10_n21731 , _u10_n21730 , _u10_n21729 , _u10_n21728 , _u10_n21727 ,_u10_n21726 , _u10_n21725 , _u10_n21724 , _u10_n21723 , _u10_n21722 ,_u10_n21721 , _u10_n21720 , _u10_n21719 , _u10_n21718 , _u10_n21717 ,_u10_n21716 , _u10_n21715 , _u10_n21714 , _u10_n21713 , _u10_n21712 ,_u10_n21711 , _u10_n21710 , _u10_n21709 , _u10_n21708 , _u10_n21707 ,_u10_n21706 , _u10_n21705 , _u10_n21704 , _u10_n21703 , _u10_n21702 ,_u10_n21701 , _u10_n21700 , _u10_n21699 , _u10_n21698 , _u10_n21697 ,_u10_n21696 , _u10_n21695 , _u10_n21694 , _u10_n21693 , _u10_n21692 ,_u10_n21691 , _u10_n21690 , _u10_n21689 , _u10_n21688 , _u10_n21687 ,_u10_n21686 , _u10_n21685 , _u10_n21684 , _u10_n21683 , _u10_n21682 ,_u10_n21681 , _u10_n21680 , _u10_n21679 , _u10_n21678 , _u10_n21677 ,_u10_n21676 , _u10_n21675 , _u10_n21674 , _u10_n21673 , _u10_n21672 ,_u10_n21671 , _u10_n21670 , _u10_n21669 , _u10_n21668 , _u10_n21667 ,_u10_n21666 , _u10_n21665 , _u10_n21664 , _u10_n21663 , _u10_n21662 ,_u10_n21661 , _u10_n21660 , _u10_n21659 , _u10_n21658 , _u10_n21657 ,_u10_n21656 , _u10_n21655 , _u10_n21654 , _u10_n21653 , _u10_n21652 ,_u10_n21651 , _u10_n21650 , _u10_n21649 , _u10_n21648 , _u10_n21647 ,_u10_n21646 , _u10_n21645 , _u10_n21644 , _u10_n21643 , _u10_n21642 ,_u10_n21641 , _u10_n21640 , _u10_n21639 , _u10_n21638 , _u10_n21637 ,_u10_n21636 , _u10_n21635 , _u10_n21634 , _u10_n21633 , _u10_n21632 ,_u10_n21631 , _u10_n21630 , _u10_n21629 , _u10_n21628 , _u10_n21627 ,_u10_n21626 , _u10_n21625 , _u10_n21624 , _u10_n21623 , _u10_n21622 ,_u10_n21621 , _u10_n21620 , _u10_n21619 , _u10_n21618 , _u10_n21617 ,_u10_n21616 , _u10_n21615 , _u10_n21614 , _u10_n21613 , _u10_n21612 ,_u10_n21611 , _u10_n21610 , _u10_n21609 , _u10_n21608 , _u10_n21607 ,_u10_n21606 , _u10_n21605 , _u10_n21604 , _u10_n21603 , _u10_n21602 ,_u10_n21601 , _u10_n21600 , _u10_n21599 , _u10_n21598 , _u10_n21597 ,_u10_n21596 , _u10_n21595 , _u10_n21594 , _u10_n21593 , _u10_n21592 ,_u10_n21591 , _u10_n21590 , _u10_n21589 , _u10_n21588 , _u10_n21587 ,_u10_n21586 , _u10_n21585 , _u10_n21584 , _u10_n21583 , _u10_n21582 ,_u10_n21581 , _u10_n21580 , _u10_n21579 , _u10_n21578 , _u10_n21577 ,_u10_n21576 , _u10_n21575 , _u10_n21574 , _u10_n21573 , _u10_n21572 ,_u10_n21571 , _u10_n21570 , _u10_n21569 , _u10_n21568 , _u10_n21567 ,_u10_n21566 , _u10_n21565 , _u10_n21564 , _u10_n21563 , _u10_n21562 ,_u10_n21561 , _u10_n21560 , _u10_n21559 , _u10_n21558 , _u10_n21557 ,_u10_n21556 , _u10_n21555 , _u10_n21554 , _u10_n21553 , _u10_n21552 ,_u10_n21551 , _u10_n21550 , _u10_n21549 , _u10_n21548 , _u10_n21547 ,_u10_n21546 , _u10_n21545 , _u10_n21544 , _u10_n21543 , _u10_n21542 ,_u10_n21541 , _u10_n21540 , _u10_n21539 , _u10_n21538 , _u10_n21537 ,_u10_n21536 , _u10_n21535 , _u10_n21534 , _u10_n21533 , _u10_n21532 ,_u10_n21531 , _u10_n21530 , _u10_n21529 , _u10_n21528 , _u10_n21527 ,_u10_n21526 , _u10_n21525 , _u10_n21524 , _u10_n21523 , _u10_n21522 ,_u10_n21521 , _u10_n21520 , _u10_n21519 , _u10_n21518 , _u10_n21517 ,_u10_n21516 , _u10_n21515 , _u10_n21514 , _u10_n21513 , _u10_n21512 ,_u10_n21511 , _u10_n21510 , _u10_n21509 , _u10_n21508 , _u10_n21507 ,_u10_n21506 , _u10_n21505 , _u10_n21504 , _u10_n21503 , _u10_n21502 ,_u10_n21501 , _u10_n21500 , _u10_n21499 , _u10_n21498 , _u10_n21497 ,_u10_n21496 , _u10_n21495 , _u10_n21494 , _u10_n21493 , _u10_n21492 ,_u10_n21491 , _u10_n21490 , _u10_n21489 , _u10_n21488 , _u10_n21487 ,_u10_n21486 , _u10_n21485 , _u10_n21484 , _u10_n21483 , _u10_n21482 ,_u10_n21481 , _u10_n21480 , _u10_n21479 , _u10_n21478 , _u10_n21477 ,_u10_n21476 , _u10_n21475 , _u10_n21474 , _u10_n21473 , _u10_n21472 ,_u10_n21471 , _u10_n21470 , _u10_n21469 , _u10_n21468 , _u10_n21467 ,_u10_n21466 , _u10_n21465 , _u10_n21464 , _u10_n21463 , _u10_n21462 ,_u10_n21461 , _u10_n21460 , _u10_n21459 , _u10_n21458 , _u10_n21457 ,_u10_n21456 , _u10_n21455 , _u10_n21454 , _u10_n21453 , _u10_n21452 ,_u10_n21451 , _u10_n21450 , _u10_n21449 , _u10_n21448 , _u10_n21447 ,_u10_n21446 , _u10_n21445 , _u10_n21444 , _u10_n21443 , _u10_n21442 ,_u10_n21441 , _u10_n21440 , _u10_n21439 , _u10_n21438 , _u10_n21437 ,_u10_n21436 , _u10_n21435 , _u10_n21434 , _u10_n21433 , _u10_n21432 ,_u10_n21431 , _u10_n21430 , _u10_n21429 , _u10_n21428 , _u10_n21427 ,_u10_n21426 , _u10_n21425 , _u10_n21424 , _u10_n21423 , _u10_n21422 ,_u10_n21421 , _u10_n21420 , _u10_n21419 , _u10_n21418 , _u10_n21417 ,_u10_n21416 , _u10_n21415 , _u10_n21414 , _u10_n21413 , _u10_n21412 ,_u10_n21411 , _u10_n21410 , _u10_n21409 , _u10_n21408 , _u10_n21407 ,_u10_n21406 , _u10_n21405 , _u10_n21404 , _u10_n21403 , _u10_n21402 ,_u10_n21401 , _u10_n21400 , _u10_n21399 , _u10_n21398 , _u10_n21397 ,_u10_n21396 , _u10_n21395 , _u10_n21394 , _u10_n21393 , _u10_n21392 ,_u10_n21391 , _u10_n21390 , _u10_n21389 , _u10_n21388 , _u10_n21387 ,_u10_n21386 , _u10_n21385 , _u10_n21384 , _u10_n21383 , _u10_n21382 ,_u10_n21381 , _u10_n21380 , _u10_n21379 , _u10_n21378 , _u10_n21377 ,_u10_n21376 , _u10_n21375 , _u10_n21374 , _u10_n21373 , _u10_n21372 ,_u10_n21371 , _u10_n21370 , _u10_n21369 , _u10_n21368 , _u10_n21367 ,_u10_n21366 , _u10_n21365 , _u10_n21364 , _u10_n21363 , _u10_n21362 ,_u10_n21361 , _u10_n21360 , _u10_n21359 , _u10_n21358 , _u10_n21357 ,_u10_n21356 , _u10_n21355 , _u10_n21354 , _u10_n21353 , _u10_n21352 ,_u10_n21351 , _u10_n21350 , _u10_n21349 , _u10_n21348 , _u10_n21347 ,_u10_n21346 , _u10_n21345 , _u10_n21344 , _u10_n21343 , _u10_n21342 ,_u10_n21341 , _u10_n21340 , _u10_n21339 , _u10_n21338 , _u10_n21337 ,_u10_n21336 , _u10_n21335 , _u10_n21334 , _u10_n21333 , _u10_n21332 ,_u10_n21331 , _u10_n21330 , _u10_n21329 , _u10_n21328 , _u10_n21327 ,_u10_n21326 , _u10_n21325 , _u10_n21324 , _u10_n21323 , _u10_n21322 ,_u10_n21321 , _u10_n21320 , _u10_n21319 , _u10_n21318 , _u10_n21317 ,_u10_n21316 , _u10_n21315 , _u10_n21314 , _u10_n21313 , _u10_n21312 ,_u10_n21311 , _u10_n21310 , _u10_n21309 , _u10_n21308 , _u10_n21307 ,_u10_n21306 , _u10_n21305 , _u10_n21304 , _u10_n21303 , _u10_n21302 ,_u10_n21301 , _u10_n21300 , _u10_n21299 , _u10_n21298 , _u10_n21297 ,_u10_n21296 , _u10_n21295 , _u10_n21294 , _u10_n21293 , _u10_n21292 ,_u10_n21291 , _u10_n21290 , _u10_n21289 , _u10_n21288 , _u10_n21287 ,_u10_n21286 , _u10_n21285 , _u10_n21284 , _u10_n21283 , _u10_n21282 ,_u10_n21281 , _u10_n21280 , _u10_n21279 , _u10_n21278 , _u10_n21277 ,_u10_n21276 , _u10_n21275 , _u10_n21274 , _u10_n21273 , _u10_n21272 ,_u10_n21271 , _u10_n21270 , _u10_n21269 , _u10_n21268 , _u10_n21267 ,_u10_n21266 , _u10_n21265 , _u10_n21264 , _u10_n21263 , _u10_n21262 ,_u10_n21261 , _u10_n21260 , _u10_n21259 , _u10_n21258 , _u10_n21257 ,_u10_n21256 , _u10_n21255 , _u10_n21254 , _u10_n21253 , _u10_n21252 ,_u10_n21251 , _u10_n21250 , _u10_n21249 , _u10_n21248 , _u10_n21247 ,_u10_n21246 , _u10_n21245 , _u10_n21244 , _u10_n21243 , _u10_n21242 ,_u10_n21241 , _u10_n21240 , _u10_n21239 , _u10_n21238 , _u10_n21237 ,_u10_n21236 , _u10_n21235 , _u10_n21234 , _u10_n21233 , _u10_n21232 ,_u10_n21231 , _u10_n21230 , _u10_n21229 , _u10_n21228 , _u10_n21227 ,_u10_n21226 , _u10_n21225 , _u10_n21224 , _u10_n21223 , _u10_n21222 ,_u10_n21221 , _u10_n21220 , _u10_n21219 , _u10_n21218 , _u10_n21217 ,_u10_n21216 , _u10_n21215 , _u10_n21214 , _u10_n21213 , _u10_n21212 ,_u10_n21211 , _u10_n21210 , _u10_n21209 , _u10_n21208 , _u10_n21207 ,_u10_n21206 , _u10_n21205 , _u10_n21204 , _u10_n21203 , _u10_n21202 ,_u10_n21201 , _u10_n21200 , _u10_n21199 , _u10_n21198 , _u10_n21197 ,_u10_n21196 , _u10_n21195 , _u10_n21194 , _u10_n21193 , _u10_n21192 ,_u10_n21191 , _u10_n21190 , _u10_n21189 , _u10_n21188 , _u10_n21187 ,_u10_n21186 , _u10_n21185 , _u10_n21184 , _u10_n21183 , _u10_n21182 ,_u10_n21181 , _u10_n21180 , _u10_n21179 , _u10_n21178 , _u10_n21177 ,_u10_n21176 , _u10_n21175 , _u10_n21174 , _u10_n21173 , _u10_n21172 ,_u10_n21171 , _u10_n21170 , _u10_n21169 , _u10_n21168 , _u10_n21167 ,_u10_n21166 , _u10_n21165 , _u10_n21164 , _u10_n21163 , _u10_n21162 ,_u10_n21161 , _u10_n21160 , _u10_n21159 , _u10_n21158 , _u10_n21157 ,_u10_n21156 , _u10_n21155 , _u10_n21154 , _u10_n21153 , _u10_n21152 ,_u10_n21151 , _u10_n21150 , _u10_n21149 , _u10_n21148 , _u10_n21147 ,_u10_n21146 , _u10_n21145 , _u10_n21144 , _u10_n21143 , _u10_n21142 ,_u10_n21141 , _u10_n21140 , _u10_n21139 , _u10_n21138 , _u10_n21137 ,_u10_n21136 , _u10_n21135 , _u10_n21134 , _u10_n21133 , _u10_n21132 ,_u10_n21131 , _u10_n21130 , _u10_n21129 , _u10_n21128 , _u10_n21127 ,_u10_n21126 , _u10_n21125 , _u10_n21124 , _u10_n21123 , _u10_n21122 ,_u10_n21121 , _u10_n21120 , _u10_n21119 , _u10_n21118 , _u10_n21117 ,_u10_n21116 , _u10_n21115 , _u10_n21114 , _u10_n21113 , _u10_n21112 ,_u10_n21111 , _u10_n21110 , _u10_n21109 , _u10_n21108 , _u10_n21107 ,_u10_n21106 , _u10_n21105 , _u10_n21104 , _u10_n21103 , _u10_n21102 ,_u10_n21101 , _u10_n21100 , _u10_n21099 , _u10_n21098 , _u10_n21097 ,_u10_n21096 , _u10_n21095 , _u10_n21094 , _u10_n21093 , _u10_n21092 ,_u10_n21091 , _u10_n21090 , _u10_n21089 , _u10_n21088 , _u10_n21087 ,_u10_n21086 , _u10_n21085 , _u10_n21084 , _u10_n21083 , _u10_n21082 ,_u10_n21081 , _u10_n21080 , _u10_n21079 , _u10_n21078 , _u10_n21077 ,_u10_n21076 , _u10_n21075 , _u10_n21074 , _u10_n21073 , _u10_n21072 ,_u10_n21071 , _u10_n21070 , _u10_n21069 , _u10_n21068 , _u10_n21067 ,_u10_n21066 , _u10_n21065 , _u10_n21064 , _u10_n21063 , _u10_n21062 ,_u10_n21061 , _u10_n21060 , _u10_n21059 , _u10_n21058 , _u10_n21057 ,_u10_n21056 , _u10_n21055 , _u10_n21054 , _u10_n21053 , _u10_n21052 ,_u10_n21051 , _u10_n21050 , _u10_n21049 , _u10_n21048 , _u10_n21047 ,_u10_n21046 , _u10_n21045 , _u10_n21044 , _u10_n21043 , _u10_n21042 ,_u10_n21041 , _u10_n21040 , _u10_n21039 , _u10_n21038 , _u10_n21037 ,_u10_n21036 , _u10_n21035 , _u10_n21034 , _u10_n21033 , _u10_n21032 ,_u10_n21031 , _u10_n21030 , _u10_n21029 , _u10_n21028 , _u10_n21027 ,_u10_n21026 , _u10_n21025 , _u10_n21024 , _u10_n21023 , _u10_n21022 ,_u10_n21021 , _u10_n21020 , _u10_n21019 , _u10_n21018 , _u10_n21017 ,_u10_n21016 , _u10_n21015 , _u10_n21014 , _u10_n21013 , _u10_n21012 ,_u10_n21011 , _u10_n21010 , _u10_n21009 , _u10_n21008 , _u10_n21007 ,_u10_n21006 , _u10_n21005 , _u10_n21004 , _u10_n21003 , _u10_n21002 ,_u10_n21001 , _u10_n21000 , _u10_n20999 , _u10_n20998 , _u10_n20997 ,_u10_n20996 , _u10_n20995 , _u10_n20994 , _u10_n20993 , _u10_n20992 ,_u10_n20991 , _u10_n20990 , _u10_n20989 , _u10_n20988 , _u10_n20987 ,_u10_n20986 , _u10_n20985 , _u10_n20984 , _u10_n20983 , _u10_n20982 ,_u10_n20981 , _u10_n20980 , _u10_n20979 , _u10_n20978 , _u10_n20977 ,_u10_n20976 , _u10_n20975 , _u10_n20974 , _u10_n20973 , _u10_n20972 ,_u10_n20971 , _u10_n20970 , _u10_n20969 , _u10_n20968 , _u10_n20967 ,_u10_n20966 , _u10_n20965 , _u10_n20964 , _u10_n20963 , _u10_n20962 ,_u10_n20961 , _u10_n20960 , _u10_n20959 , _u10_n20958 , _u10_n20957 ,_u10_n20956 , _u10_n20955 , _u10_n20954 , _u10_n20953 , _u10_n20952 ,_u10_n20951 , _u10_n20950 , _u10_n20949 , _u10_n20948 , _u10_n20947 ,_u10_n20946 , _u10_n20945 , _u10_n20944 , _u10_n20943 , _u10_n20942 ,_u10_n20941 , _u10_n20940 , _u10_n20939 , _u10_n20938 , _u10_n20937 ,_u10_n20936 , _u10_n20935 , _u10_n20934 , _u10_n20933 , _u10_n20932 ,_u10_n20931 , _u10_n20930 , _u10_n20929 , _u10_n20928 , _u10_n20927 ,_u10_n20926 , _u10_n20925 , _u10_n20924 , _u10_n20923 , _u10_n20922 ,_u10_n20921 , _u10_n20920 , _u10_n20919 , _u10_n20918 , _u10_n20917 ,_u10_n20916 , _u10_n20915 , _u10_n20914 , _u10_n20913 , _u10_n20912 ,_u10_n20911 , _u10_n20910 , _u10_n20909 , _u10_n20908 , _u10_n20907 ,_u10_n20906 , _u10_n20905 , _u10_n20904 , _u10_n20903 , _u10_n20902 ,_u10_n20901 , _u10_n20900 , _u10_n20899 , _u10_n20898 , _u10_n20897 ,_u10_n20896 , _u10_n20895 , _u10_n20894 , _u10_n20893 , _u10_n20892 ,_u10_n20891 , _u10_n20890 , _u10_n20889 , _u10_n20888 , _u10_n20887 ,_u10_n20886 , _u10_n20885 , _u10_n20884 , _u10_n20883 , _u10_n20882 ,_u10_n20881 , _u10_n20880 , _u10_n20879 , _u10_n20878 , _u10_n20877 ,_u10_n20876 , _u10_n20875 , _u10_n20874 , _u10_n20873 , _u10_n20872 ,_u10_n20871 , _u10_n20870 , _u10_n20869 , _u10_n20868 , _u10_n20867 ,_u10_n20866 , _u10_n20865 , _u10_n20864 , _u10_n20863 , _u10_n20862 ,_u10_n20861 , _u10_n20860 , _u10_n20859 , _u10_n20858 , _u10_n20857 ,_u10_n20856 , _u10_n20855 , _u10_n20854 , _u10_n20853 , _u10_n20852 ,_u10_n20851 , _u10_n20850 , _u10_n20849 , _u10_n20848 , _u10_n20847 ,_u10_n20846 , _u10_n20845 , _u10_n20844 , _u10_n20843 , _u10_n20842 ,_u10_n20841 , _u10_n20840 , _u10_n20839 , _u10_n20838 , _u10_n20837 ,_u10_n20836 , _u10_n20835 , _u10_n20834 , _u10_n20833 , _u10_n20832 ,_u10_n20831 , _u10_n20830 , _u10_n20829 , _u10_n20828 , _u10_n20827 ,_u10_n20826 , _u10_n20825 , _u10_n20824 , _u10_n20823 , _u10_n20822 ,_u10_n20821 , _u10_n20820 , _u10_n20819 , _u10_n20818 , _u10_n20817 ,_u10_n20816 , _u10_n20815 , _u10_n20814 , _u10_n20813 , _u10_n20812 ,_u10_n20811 , _u10_n20810 , _u10_n20809 , _u10_n20808 , _u10_n20807 ,_u10_n20806 , _u10_n20805 , _u10_n20804 , _u10_n20803 , _u10_n20802 ,_u10_n20801 , _u10_n20800 , _u10_n20799 , _u10_n20798 , _u10_n20797 ,_u10_n20796 , _u10_n20795 , _u10_n20794 , _u10_n20793 , _u10_n20792 ,_u10_n20791 , _u10_n20790 , _u10_n20789 , _u10_n20788 , _u10_n20787 ,_u10_n20786 , _u10_n20785 , _u10_n20784 , _u10_n20783 , _u10_n20782 ,_u10_n20781 , _u10_n20780 , _u10_n20779 , _u10_n20778 , _u10_n20777 ,_u10_n20776 , _u10_n20775 , _u10_n20774 , _u10_n20773 , _u10_n20772 ,_u10_n20771 , _u10_n20770 , _u10_n20769 , _u10_n20768 , _u10_n20767 ,_u10_n20766 , _u10_n20765 , _u10_n20764 , _u10_n20763 , _u10_n20762 ,_u10_n20761 , _u10_n20760 , _u10_n20759 , _u10_n20758 , _u10_n20757 ,_u10_n20756 , _u10_n20755 , _u10_n20754 , _u10_n20753 , _u10_n20752 ,_u10_n20751 , _u10_n20750 , _u10_n20749 , _u10_n20748 , _u10_n20747 ,_u10_n20746 , _u10_n20745 , _u10_n20744 , _u10_n20743 , _u10_n20742 ,_u10_n20741 , _u10_n20740 , _u10_n20739 , _u10_n20738 , _u10_n20737 ,_u10_n20736 , _u10_n20735 , _u10_n20734 , _u10_n20733 , _u10_n20732 ,_u10_n20731 , _u10_n20730 , _u10_n20729 , _u10_n20728 , _u10_n20727 ,_u10_n20726 , _u10_n20725 , _u10_n20724 , _u10_n20723 , _u10_n20722 ,_u10_n20721 , _u10_n20720 , _u10_n20719 , _u10_n20718 , _u10_n20717 ,_u10_n20716 , _u10_n20715 , _u10_n20714 , _u10_n20713 , _u10_n20712 ,_u10_n20711 , _u10_n20710 , _u10_n20709 , _u10_n20708 , _u10_n20707 ,_u10_n20706 , _u10_n20705 , _u10_n20704 , _u10_n20703 , _u10_n20702 ,_u10_n20701 , _u10_n20700 , _u10_n20699 , _u10_n20698 , _u10_n20697 ,_u10_n20696 , _u10_n20695 , _u10_n20694 , _u10_n20693 , _u10_n20692 ,_u10_n20691 , _u10_n20690 , _u10_n20689 , _u10_n20688 , _u10_n20687 ,_u10_n20686 , _u10_n20685 , _u10_n20684 , _u10_n20683 , _u10_n20682 ,_u10_n20681 , _u10_n20680 , _u10_n20679 , _u10_n20678 , _u10_n20677 ,_u10_n20676 , _u10_n20675 , _u10_n20674 , _u10_n20673 , _u10_n20672 ,_u10_n20671 , _u10_n20670 , _u10_n20669 , _u10_n20668 , _u10_n20667 ,_u10_n20666 , _u10_n20665 , _u10_n20664 , _u10_n20663 , _u10_n20662 ,_u10_n20661 , _u10_n20660 , _u10_n20659 , _u10_n20658 , _u10_n20657 ,_u10_n20656 , _u10_n20655 , _u10_n20654 , _u10_n20653 , _u10_n20652 ,_u10_n20651 , _u10_n20650 , _u10_n20649 , _u10_n20648 , _u10_n20647 ,_u10_n20646 , _u10_n20645 , _u10_n20644 , _u10_n20643 , _u10_n20642 ,_u10_n20641 , _u10_n20640 , _u10_n20639 , _u10_n20638 , _u10_n20637 ,_u10_n20636 , _u10_n20635 , _u10_n20634 , _u10_n20633 , _u10_n20632 ,_u10_n20631 , _u10_n20630 , _u10_n20629 , _u10_n20628 , _u10_n20627 ,_u10_n20626 , _u10_n20625 , _u10_n20624 , _u10_n20623 , _u10_n20622 ,_u10_n20621 , _u10_n20620 , _u10_n20619 , _u10_n20618 , _u10_n20617 ,_u10_n20616 , _u10_n20615 , _u10_n20614 , _u10_n20613 , _u10_n20612 ,_u10_n20611 , _u10_n20610 , _u10_n20609 , _u10_n20608 , _u10_n20607 ,_u10_n20606 , _u10_n20605 , _u10_n20604 , _u10_n20603 , _u10_n20602 ,_u10_n20601 , _u10_n20600 , _u10_n20599 , _u10_n20598 , _u10_n20597 ,_u10_n20596 , _u10_n20595 , _u10_n20594 , _u10_n20593 , _u10_n20592 ,_u10_n20591 , _u10_n20590 , _u10_n20589 , _u10_n20588 , _u10_n20587 ,_u10_n20586 , _u10_n20585 , _u10_n20584 , _u10_n20583 , _u10_n20582 ,_u10_n20581 , _u10_n20580 , _u10_n20579 , _u10_n20578 , _u10_n20577 ,_u10_n20576 , _u10_n20575 , _u10_n20574 , _u10_n20573 , _u10_n20572 ,_u10_n20571 , _u10_n20570 , _u10_n20569 , _u10_n20568 , _u10_n20567 ,_u10_n20566 , _u10_n20565 , _u10_n20564 , _u10_n20563 , _u10_n20562 ,_u10_n20561 , _u10_n20560 , _u10_n20559 , _u10_n20558 , _u10_n20557 ,_u10_n20556 , _u10_n20555 , _u10_n20554 , _u10_n20553 , _u10_n20552 ,_u10_n20551 , _u10_n20550 , _u10_n20549 , _u10_n20548 , _u10_n20547 ,_u10_n20546 , _u10_n20545 , _u10_n20544 , _u10_n20543 , _u10_n20542 ,_u10_n20541 , _u10_n20540 , _u10_n20539 , _u10_n20538 , _u10_n20537 ,_u10_n20536 , _u10_n20535 , _u10_n20534 , _u10_n20533 , _u10_n20532 ,_u10_n20531 , _u10_n20530 , _u10_n20529 , _u10_n20528 , _u10_n20527 ,_u10_n20526 , _u10_n20525 , _u10_n20524 , _u10_n20523 , _u10_n20522 ,_u10_n20521 , _u10_n20520 , _u10_n20519 , _u10_n20518 , _u10_n20517 ,_u10_n20516 , _u10_n20515 , _u10_n20514 , _u10_n20513 , _u10_n20512 ,_u10_n20511 , _u10_n20510 , _u10_n20509 , _u10_n20508 , _u10_n20507 ,_u10_n20506 , _u10_n20505 , _u10_n20504 , _u10_n20503 , _u10_n20502 ,_u10_n20501 , _u10_n20500 , _u10_n20499 , _u10_n20498 , _u10_n20497 ,_u10_n20496 , _u10_n20495 , _u10_n20494 , _u10_n20493 , _u10_n20492 ,_u10_n20491 , _u10_n20490 , _u10_n20489 , _u10_n20488 , _u10_n20487 ,_u10_n20486 , _u10_n20485 , _u10_n20484 , _u10_n20483 , _u10_n20482 ,_u10_n20481 , _u10_n20480 , _u10_n20479 , _u10_n20478 , _u10_n20477 ,_u10_n20476 , _u10_n20475 , _u10_n20474 , _u10_n20473 , _u10_n20472 ,_u10_n20471 , _u10_n20470 , _u10_n20469 , _u10_n20468 , _u10_n20467 ,_u10_n20466 , _u10_n20465 , _u10_n20464 , _u10_n20463 , _u10_n20462 ,_u10_n20461 , _u10_n20460 , _u10_n20459 , _u10_n20458 , _u10_n20457 ,_u10_n20456 , _u10_n20455 , _u10_n20454 , _u10_n20453 , _u10_n20452 ,_u10_n20451 , _u10_n20450 , _u10_n20449 , _u10_n20448 , _u10_n20447 ,_u10_n20446 , _u10_n20445 , _u10_n20444 , _u10_n20443 , _u10_n20442 ,_u10_n20441 , _u10_n20440 , _u10_n20439 , _u10_n20438 , _u10_n20437 ,_u10_n20436 , _u10_n20435 , _u10_n20434 , _u10_n20433 , _u10_n20432 ,_u10_n20431 , _u10_n20430 , _u10_n20429 , _u10_n20428 , _u10_n20427 ,_u10_n20426 , _u10_n20425 , _u10_n20424 , _u10_n20423 , _u10_n20422 ,_u10_n20421 , _u10_n20420 , _u10_n20419 , _u10_n20418 , _u10_n20417 ,_u10_n20416 , _u10_n20415 , _u10_n20414 , _u10_n20413 , _u10_n20412 ,_u10_n20411 , _u10_n20410 , _u10_n20409 , _u10_n20408 , _u10_n20407 ,_u10_n20406 , _u10_n20405 , _u10_n20404 , _u10_n20403 , _u10_n20402 ,_u10_n20401 , _u10_n20400 , _u10_n20399 , _u10_n20398 , _u10_n20397 ,_u10_n20396 , _u10_n20395 , _u10_n20394 , _u10_n20393 , _u10_n20392 ,_u10_n20391 , _u10_n20390 , _u10_n20389 , _u10_n20388 , _u10_n20387 ,_u10_n20386 , _u10_n20385 , _u10_n20384 , _u10_n20383 , _u10_n20382 ,_u10_n20381 , _u10_n20380 , _u10_n20379 , _u10_n20378 , _u10_n20377 ,_u10_n20376 , _u10_n20375 , _u10_n20374 , _u10_n20373 , _u10_n20372 ,_u10_n20371 , _u10_n20370 , _u10_n20369 , _u10_n20368 , _u10_n20367 ,_u10_n20366 , _u10_n20365 , _u10_n20364 , _u10_n20363 , _u10_n20362 ,_u10_n20361 , _u10_n20360 , _u10_n20359 , _u10_n20358 , _u10_n20357 ,_u10_n20356 , _u10_n20355 , _u10_n20354 , _u10_n20353 , _u10_n20352 ,_u10_n20351 , _u10_n20350 , _u10_n20349 , _u10_n20348 , _u10_n20347 ,_u10_n20346 , _u10_n20345 , _u10_n20344 , _u10_n20343 , _u10_n20342 ,_u10_n20341 , _u10_n20340 , _u10_n20339 , _u10_n20338 , _u10_n20337 ,_u10_n20336 , _u10_n20335 , _u10_n20334 , _u10_n20333 , _u10_n20332 ,_u10_n20331 , _u10_n20330 , _u10_n20329 , _u10_n20328 , _u10_n20327 ,_u10_n20326 , _u10_n20325 , _u10_n20324 , _u10_n20323 , _u10_n20322 ,_u10_n20321 , _u10_n20320 , _u10_n20319 , _u10_n20318 , _u10_n20317 ,_u10_n20316 , _u10_n20315 , _u10_n20314 , _u10_n20313 , _u10_n20312 ,_u10_n20311 , _u10_n20310 , _u10_n20309 , _u10_n20308 , _u10_n20307 ,_u10_n20306 , _u10_n20305 , _u10_n20304 , _u10_n20303 , _u10_n20302 ,_u10_n20301 , _u10_n20300 , _u10_n20299 , _u10_n20298 , _u10_n20297 ,_u10_n20296 , _u10_n20295 , _u10_n20294 , _u10_n20293 , _u10_n20292 ,_u10_n20291 , _u10_n20290 , _u10_n20289 , _u10_n20288 , _u10_n20287 ,_u10_n20286 , _u10_n20285 , _u10_n20284 , _u10_n20283 , _u10_n20282 ,_u10_n20281 , _u10_n20280 , _u10_n20279 , _u10_n20278 , _u10_n20277 ,_u10_n20276 , _u10_n20275 , _u10_n20274 , _u10_n20273 , _u10_n20272 ,_u10_n20271 , _u10_n20270 , _u10_n20269 , _u10_n20268 , _u10_n20267 ,_u10_n20266 , _u10_n20265 , _u10_n20264 , _u10_n20263 , _u10_n20262 ,_u10_n20261 , _u10_n20260 , _u10_n20259 , _u10_n20258 , _u10_n20257 ,_u10_n20256 , _u10_n20255 , _u10_n20254 , _u10_n20253 , _u10_n20252 ,_u10_n20251 , _u10_n20250 , _u10_n20249 , _u10_n20248 , _u10_n20247 ,_u10_n20246 , _u10_n20245 , _u10_n20244 , _u10_n20243 , _u10_n20242 ,_u10_n20241 , _u10_n20240 , _u10_n20239 , _u10_n20238 , _u10_n20237 ,_u10_n20236 , _u10_n20235 , _u10_n20234 , _u10_n20233 , _u10_n20232 ,_u10_n20231 , _u10_n20230 , _u10_n20229 , _u10_n20228 , _u10_n20227 ,_u10_n20226 , _u10_n20225 , _u10_n20224 , _u10_n20223 , _u10_n20222 ,_u10_n20221 , _u10_n20220 , _u10_n20219 , _u10_n20218 , _u10_n20217 ,_u10_n20216 , _u10_n20215 , _u10_n20214 , _u10_n20213 , _u10_n20212 ,_u10_n20211 , _u10_n20210 , _u10_n20209 , _u10_n20208 , _u10_n20207 ,_u10_n20206 , _u10_n20205 , _u10_n20204 , _u10_n20203 , _u10_n20202 ,_u10_n20201 , _u10_n20200 , _u10_n20199 , _u10_n20198 , _u10_n20197 ,_u10_n20196 , _u10_n20195 , _u10_n20194 , _u10_n20193 , _u10_n20192 ,_u10_n20191 , _u10_n20190 , _u10_n20189 , _u10_n20188 , _u10_n20187 ,_u10_n20186 , _u10_n20185 , _u10_n20184 , _u10_n20183 , _u10_n20182 ,_u10_n20181 , _u10_n20180 , _u10_n20179 , _u10_n20178 , _u10_n20177 ,_u10_n20176 , _u10_n20175 , _u10_n20174 , _u10_n20173 , _u10_n20172 ,_u10_n20171 , _u10_n20170 , _u10_n20169 , _u10_n20168 , _u10_n20167 ,_u10_n20166 , _u10_n20165 , _u10_n20164 , _u10_n20163 , _u10_n20162 ,_u10_n20161 , _u10_n20160 , _u10_n20159 , _u10_n20158 , _u10_n20157 ,_u10_n20156 , _u10_n20155 , _u10_n20154 , _u10_n20153 , _u10_n20152 ,_u10_n20151 , _u10_n20150 , _u10_n20149 , _u10_n20148 , _u10_n20147 ,_u10_n20146 , _u10_n20145 , _u10_n20144 , _u10_n20143 , _u10_n20142 ,_u10_n20141 , _u10_n20140 , _u10_n20139 , _u10_n20138 , _u10_n20137 ,_u10_n20136 , _u10_n20135 , _u10_n20134 , _u10_n20133 , _u10_n20132 ,_u10_n20131 , _u10_n20130 , _u10_n20129 , _u10_n20128 , _u10_n20127 ,_u10_n20126 , _u10_n20125 , _u10_n20124 , _u10_n20123 , _u10_n20122 ,_u10_n20121 , _u10_n20120 , _u10_n20119 , _u10_n20118 , _u10_n20117 ,_u10_n20116 , _u10_n20115 , _u10_n20114 , _u10_n20113 , _u10_n20112 ,_u10_n20111 , _u10_n20110 , _u10_n20109 , _u10_n20108 , _u10_n20107 ,_u10_n20106 , _u10_n20105 , _u10_n20104 , _u10_n20103 , _u10_n20102 ,_u10_n20101 , _u10_n20100 , _u10_n20099 , _u10_n20098 , _u10_n20097 ,_u10_n20096 , _u10_n20095 , _u10_n20094 , _u10_n20093 , _u10_n20092 ,_u10_n20091 , _u10_n20090 , _u10_n20089 , _u10_n20088 , _u10_n20087 ,_u10_n20086 , _u10_n20085 , _u10_n20084 , _u10_n20083 , _u10_n20082 ,_u10_n20081 , _u10_n20080 , _u10_n20079 , _u10_n20078 , _u10_n20077 ,_u10_n20076 , _u10_n20075 , _u10_n20074 , _u10_n20073 , _u10_n20072 ,_u10_n20071 , _u10_n20070 , _u10_n20069 , _u10_n20068 , _u10_n20067 ,_u10_n20066 , _u10_n20065 , _u10_n20064 , _u10_n20063 , _u10_n20062 ,_u10_n20061 , _u10_n20060 , _u10_n20059 , _u10_n20058 , _u10_n20057 ,_u10_n20056 , _u10_n20055 , _u10_n20054 , _u10_n20053 , _u10_n20052 ,_u10_n20051 , _u10_n20050 , _u10_n20049 , _u10_n20048 , _u10_n20047 ,_u10_n20046 , _u10_n20045 , _u10_n20044 , _u10_n20043 , _u10_n20042 ,_u10_n20041 , _u10_n20040 , _u10_n20039 , _u10_n20038 , _u10_n20037 ,_u10_n20036 , _u10_n20035 , _u10_n20034 , _u10_n20033 , _u10_n20032 ,_u10_n20031 , _u10_n20030 , _u10_n20029 , _u10_n20028 , _u10_n20027 ,_u10_n20026 , _u10_n20025 , _u10_n20024 , _u10_n20023 , _u10_n20022 ,_u10_n20021 , _u10_n20020 , _u10_n20019 , _u10_n20018 , _u10_n20017 ,_u10_n20016 , _u10_n20015 , _u10_n20014 , _u10_n20013 , _u10_n20012 ,_u10_n20011 , _u10_n20010 , _u10_n20009 , _u10_n20008 , _u10_n20007 ,_u10_n20006 , _u10_n20005 , _u10_n20004 , _u10_n20003 , _u10_n20002 ,_u10_n20001 , _u10_n20000 , _u10_n19999 , _u10_n19998 , _u10_n19997 ,_u10_n19996 , _u10_n19995 , _u10_n19994 , _u10_n19993 , _u10_n19992 ,_u10_n19991 , _u10_n19990 , _u10_n19989 , _u10_n19988 , _u10_n19987 ,_u10_n19986 , _u10_n19985 , _u10_n19984 , _u10_n19983 , _u10_n19982 ,_u10_n19981 , _u10_n19980 , _u10_n19979 , _u10_n19978 , _u10_n19977 ,_u10_n19976 , _u10_n19975 , _u10_n19974 , _u10_n19973 , _u10_n19972 ,_u10_n19971 , _u10_n19970 , _u10_n19969 , _u10_n19968 , _u10_n19967 ,_u10_n19966 , _u10_n19965 , _u10_n19964 , _u10_n19963 , _u10_n19962 ,_u10_n19961 , _u10_n19960 , _u10_n19959 , _u10_n19958 , _u10_n19957 ,_u10_n19956 , _u10_n19955 , _u10_n19954 , _u10_n19953 , _u10_n19952 ,_u10_n19951 , _u10_n19950 , _u10_n19949 , _u10_n19948 , _u10_n19947 ,_u10_n19946 , _u10_n19945 , _u10_n19944 , _u10_n19943 , _u10_n19942 ,_u10_n19941 , _u10_n19940 , _u10_n19939 , _u10_n19938 , _u10_n19937 ,_u10_n19936 , _u10_n19935 , _u10_n19934 , _u10_n19933 , _u10_n19932 ,_u10_n19931 , _u10_n19930 , _u10_n19929 , _u10_n19928 , _u10_n19927 ,_u10_n19926 , _u10_n19925 , _u10_n19924 , _u10_n19923 , _u10_n19922 ,_u10_n19921 , _u10_n19920 , _u10_n19919 , _u10_n19918 , _u10_n19917 ,_u10_n19916 , _u10_n19915 , _u10_n19914 , _u10_n19913 , _u10_n19912 ,_u10_n19911 , _u10_n19910 , _u10_n19909 , _u10_n19908 , _u10_n19907 ,_u10_n19906 , _u10_n19905 , _u10_n19904 , _u10_n19903 , _u10_n19902 ,_u10_n19901 , _u10_n19900 , _u10_n19899 , _u10_n19898 , _u10_n19897 ,_u10_n19896 , _u10_n19895 , _u10_n19894 , _u10_n19893 , _u10_n19892 ,_u10_n19891 , _u10_n19890 , _u10_n19889 , _u10_n19888 , _u10_n19887 ,_u10_n19886 , _u10_n19885 , _u10_n19884 , _u10_n19883 , _u10_n19882 ,_u10_n19881 , _u10_n19880 , _u10_n19879 , _u10_n19878 , _u10_n19877 ,_u10_n19876 , _u10_n19875 , _u10_n19874 , _u10_n19873 , _u10_n19872 ,_u10_n19871 , _u10_n19870 , _u10_n19869 , _u10_n19868 , _u10_n19867 ,_u10_n19866 , _u10_n19865 , _u10_n19864 , _u10_n19863 , _u10_n19862 ,_u10_n19861 , _u10_n19860 , _u10_n19859 , _u10_n19858 , _u10_n19857 ,_u10_n19856 , _u10_n19855 , _u10_n19854 , _u10_n19853 , _u10_n19852 ,_u10_n19851 , _u10_n19850 , _u10_n19849 , _u10_n19848 , _u10_n19847 ,_u10_n19846 , _u10_n19845 , _u10_n19844 , _u10_n19843 , _u10_n19842 ,_u10_n19841 , _u10_n19840 , _u10_n19839 , _u10_n19838 , _u10_n19837 ,_u10_n19836 , _u10_n19835 , _u10_n19834 , _u10_n19833 , _u10_n19832 ,_u10_n19831 , _u10_n19830 , _u10_n19829 , _u10_n19828 , _u10_n19827 ,_u10_n19826 , _u10_n19825 , _u10_n19824 , _u10_n19823 , _u10_n19822 ,_u10_n19821 , _u10_n19820 , _u10_n19819 , _u10_n19818 , _u10_n19817 ,_u10_n19816 , _u10_n19815 , _u10_n19814 , _u10_n19813 , _u10_n19812 ,_u10_n19811 , _u10_n19810 , _u10_n19809 , _u10_n19808 , _u10_n19807 ,_u10_n19806 , _u10_n19805 , _u10_n19804 , _u10_n19803 , _u10_n19802 ,_u10_n19801 , _u10_n19800 , _u10_n19799 , _u10_n19798 , _u10_n19797 ,_u10_n19796 , _u10_n19795 , _u10_n19794 , _u10_n19793 , _u10_n19792 ,_u10_n19791 , _u10_n19790 , _u10_n19789 , _u10_n19788 , _u10_n19787 ,_u10_n19786 , _u10_n19785 , _u10_n19784 , _u10_n19783 , _u10_n19782 ,_u10_n19781 , _u10_n19780 , _u10_n19779 , _u10_n19778 , _u10_n19777 ,_u10_n19776 , _u10_n19775 , _u10_n19774 , _u10_n19773 , _u10_n19772 ,_u10_n19771 , _u10_n19770 , _u10_n19769 , _u10_n19768 , _u10_n19767 ,_u10_n19766 , _u10_n19765 , _u10_n19764 , _u10_n19763 , _u10_n19762 ,_u10_n19761 , _u10_n19760 , _u10_n19759 , _u10_n19758 , _u10_n19757 ,_u10_n19756 , _u10_n19755 , _u10_n19754 , _u10_n19753 , _u10_n19752 ,_u10_n19751 , _u10_n19750 , _u10_n19749 , _u10_n19748 , _u10_n19747 ,_u10_n19746 , _u10_n19745 , _u10_n19744 , _u10_n19743 , _u10_n19742 ,_u10_n19741 , _u10_n19740 , _u10_n19739 , _u10_n19738 , _u10_n19737 ,_u10_n19736 , _u10_n19735 , _u10_n19734 , _u10_n19733 , _u10_n19732 ,_u10_n19731 , _u10_n19730 , _u10_n19729 , _u10_n19728 , _u10_n19727 ,_u10_n19726 , _u10_n19725 , _u10_n19724 , _u10_n19723 , _u10_n19722 ,_u10_n19721 , _u10_n19720 , _u10_n19719 , _u10_n19718 , _u10_n19717 ,_u10_n19716 , _u10_n19715 , _u10_n19714 , _u10_n19713 , _u10_n19712 ,_u10_n19711 , _u10_n19710 , _u10_n19709 , _u10_n19708 , _u10_n19707 ,_u10_n19706 , _u10_n19705 , _u10_n19704 , _u10_n19703 , _u10_n19702 ,_u10_n19701 , _u10_n19700 , _u10_n19699 , _u10_n19698 , _u10_n19697 ,_u10_n19696 , _u10_n19695 , _u10_n19694 , _u10_n19693 , _u10_n19692 ,_u10_n19691 , _u10_n19690 , _u10_n19689 , _u10_n19688 , _u10_n19687 ,_u10_n19686 , _u10_n19685 , _u10_n19684 , _u10_n19683 , _u10_n19682 ,_u10_n19681 , _u10_n19680 , _u10_n19679 , _u10_n19678 , _u10_n19677 ,_u10_n19676 , _u10_n19675 , _u10_n19674 , _u10_n19673 , _u10_n19672 ,_u10_n19671 , _u10_n19670 , _u10_n19669 , _u10_n19668 , _u10_n19667 ,_u10_n19666 , _u10_n19665 , _u10_n19664 , _u10_n19663 , _u10_n19662 ,_u10_n19661 , _u10_n19660 , _u10_n19659 , _u10_n19658 , _u10_n19657 ,_u10_n19656 , _u10_n19655 , _u10_n19654 , _u10_n19653 , _u10_n19652 ,_u10_n19651 , _u10_n19650 , _u10_n19649 , _u10_n19648 , _u10_n19647 ,_u10_n19646 , _u10_n19645 , _u10_n19644 , _u10_n19643 , _u10_n19642 ,_u10_n19641 , _u10_n19640 , _u10_n19639 , _u10_n19638 , _u10_n19637 ,_u10_n19636 , _u10_n19635 , _u10_n19634 , _u10_n19633 , _u10_n19632 ,_u10_n19631 , _u10_n19630 , _u10_n19629 , _u10_n19628 , _u10_n19627 ,_u10_n19626 , _u10_n19625 , _u10_n19624 , _u10_n19623 , _u10_n19622 ,_u10_n19621 , _u10_n19620 , _u10_n19619 , _u10_n19618 , _u10_n19617 ,_u10_n19616 , _u10_n19615 , _u10_n19614 , _u10_n19613 , _u10_n19612 ,_u10_n19611 , _u10_n19610 , _u10_n19609 , _u10_n19608 , _u10_n19607 ,_u10_n19606 , _u10_n19605 , _u10_n19604 , _u10_n19603 , _u10_n19602 ,_u10_n19601 , _u10_n19600 , _u10_n19599 , _u10_n19598 , _u10_n19597 ,_u10_n19596 , _u10_n19595 , _u10_n19594 , _u10_n19593 , _u10_n19592 ,_u10_n19591 , _u10_n19590 , _u10_n19589 , _u10_n19588 , _u10_n19587 ,_u10_n19586 , _u10_n19585 , _u10_n19584 , _u10_n19583 , _u10_n19582 ,_u10_n19581 , _u10_n19580 , _u10_n19579 , _u10_n19578 , _u10_n19577 ,_u10_n19576 , _u10_n19575 , _u10_n19574 , _u10_n19573 , _u10_n19572 ,_u10_n19571 , _u10_n19570 , _u10_n19569 , _u10_n19568 , _u10_n19567 ,_u10_n19566 , _u10_n19565 , _u10_n19564 , _u10_n19563 , _u10_n19562 ,_u10_n19561 , _u10_n19560 , _u10_n19559 , _u10_n19558 , _u10_n19557 ,_u10_n19556 , _u10_n19555 , _u10_n19554 , _u10_n19553 , _u10_n19552 ,_u10_n19551 , _u10_n19550 , _u10_n19549 , _u10_n19548 , _u10_n19547 ,_u10_n19546 , _u10_n19545 , _u10_n19544 , _u10_n19543 , _u10_n19542 ,_u10_n19541 , _u10_n19540 , _u10_n19539 , _u10_n19538 , _u10_n19537 ,_u10_n19536 , _u10_n19535 , _u10_n19534 , _u10_n19533 , _u10_n19532 ,_u10_n19531 , _u10_n19530 , _u10_n19529 , _u10_n19528 , _u10_n19527 ,_u10_n19526 , _u10_n19525 , _u10_n19524 , _u10_n19523 , _u10_n19522 ,_u10_n19521 , _u10_n19520 , _u10_n19519 , _u10_n19518 , _u10_n19517 ,_u10_n19516 , _u10_n19515 , _u10_n19514 , _u10_n19513 , _u10_n19512 ,_u10_n19511 , _u10_n19510 , _u10_n19509 , _u10_n19508 , _u10_n19507 ,_u10_n19506 , _u10_n19505 , _u10_n19504 , _u10_n19503 , _u10_n19502 ,_u10_n19501 , _u10_n19500 , _u10_n19499 , _u10_n19498 , _u10_n19497 ,_u10_n19496 , _u10_n19495 , _u10_n19494 , _u10_n19493 , _u10_n19492 ,_u10_n19491 , _u10_n19490 , _u10_n19489 , _u10_n19488 , _u10_n19487 ,_u10_n19486 , _u10_n19485 , _u10_n19484 , _u10_n19483 , _u10_n19482 ,_u10_n19481 , _u10_n19480 , _u10_n19479 , _u10_n19478 , _u10_n19477 ,_u10_n19476 , _u10_n19475 , _u10_n19474 , _u10_n19473 , _u10_n19472 ,_u10_n19471 , _u10_n19470 , _u10_n19469 , _u10_n19468 , _u10_n19467 ,_u10_n19466 , _u10_n19465 , _u10_n19464 , _u10_n19463 , _u10_n19462 ,_u10_n19461 , _u10_n19460 , _u10_n19459 , _u10_n19458 , _u10_n19457 ,_u10_n19456 , _u10_n19455 , _u10_n19454 , _u10_n19453 , _u10_n19452 ,_u10_n19451 , _u10_n19450 , _u10_n19449 , _u10_n19448 , _u10_n19447 ,_u10_n19446 , _u10_n19445 , _u10_n19444 , _u10_n19443 , _u10_n19442 ,_u10_n19441 , _u10_n19440 , _u10_n19439 , _u10_n19438 , _u10_n19437 ,_u10_n19436 , _u10_n19435 , _u10_n19434 , _u10_n19433 , _u10_n19432 ,_u10_n19431 , _u10_n19430 , _u10_n19429 , _u10_n19428 , _u10_n19427 ,_u10_n19426 , _u10_n19425 , _u10_n19424 , _u10_n19423 , _u10_n19422 ,_u10_n19421 , _u10_n19420 , _u10_n19419 , _u10_n19418 , _u10_n19417 ,_u10_n19416 , _u10_n19415 , _u10_n19414 , _u10_n19413 , _u10_n19412 ,_u10_n19411 , _u10_n19410 , _u10_n19409 , _u10_n19408 , _u10_n19407 ,_u10_n19406 , _u10_n19405 , _u10_n19404 , _u10_n19403 , _u10_n19402 ,_u10_n19401 , _u10_n19400 , _u10_n19399 , _u10_n19398 , _u10_n19397 ,_u10_n19396 , _u10_n19395 , _u10_n19394 , _u10_n19393 , _u10_n19392 ,_u10_n19391 , _u10_n19390 , _u10_n19389 , _u10_n19388 , _u10_n19387 ,_u10_n19386 , _u10_n19385 , _u10_n19384 , _u10_n19383 , _u10_n19382 ,_u10_n19381 , _u10_n19380 , _u10_n19379 , _u10_n19378 , _u10_n19377 ,_u10_n19376 , _u10_n19375 , _u10_n19374 , _u10_n19373 , _u10_n19372 ,_u10_n19371 , _u10_n19370 , _u10_n19369 , _u10_n19368 , _u10_n19367 ,_u10_n19366 , _u10_n19365 , _u10_n19364 , _u10_n19363 , _u10_n19362 ,_u10_n19361 , _u10_n19360 , _u10_n19359 , _u10_n19358 , _u10_n19357 ,_u10_n19356 , _u10_n19355 , _u10_n19354 , _u10_n19353 , _u10_n19352 ,_u10_n19351 , _u10_n19350 , _u10_n19349 , _u10_n19348 , _u10_n19347 ,_u10_n19346 , _u10_n19345 , _u10_n19344 , _u10_n19343 , _u10_n19342 ,_u10_n19341 , _u10_n19340 , _u10_n19339 , _u10_n19338 , _u10_n19337 ,_u10_n19336 , _u10_n19335 , _u10_n19334 , _u10_n19333 , _u10_n19332 ,_u10_n19331 , _u10_n19330 , _u10_n19329 , _u10_n19328 , _u10_n19327 ,_u10_n19326 , _u10_n19325 , _u10_n19324 , _u10_n19323 , _u10_n19322 ,_u10_n19321 , _u10_n19320 , _u10_n19319 , _u10_n19318 , _u10_n19317 ,_u10_n19316 , _u10_n19315 , _u10_n19314 , _u10_n19313 , _u10_n19312 ,_u10_n19311 , _u10_n19310 , _u10_n19309 , _u10_n19308 , _u10_n19307 ,_u10_n19306 , _u10_n19305 , _u10_n19304 , _u10_n19303 , _u10_n19302 ,_u10_n19301 , _u10_n19300 , _u10_n19299 , _u10_n19298 , _u10_n19297 ,_u10_n19296 , _u10_n19295 , _u10_n19294 , _u10_n19293 , _u10_n19292 ,_u10_n19291 , _u10_n19290 , _u10_n19289 , _u10_n19288 , _u10_n19287 ,_u10_n19286 , _u10_n19285 , _u10_n19284 , _u10_n19283 , _u10_n19282 ,_u10_n19281 , _u10_n19280 , _u10_n19279 , _u10_n19278 , _u10_n19277 ,_u10_n19276 , _u10_n19275 , _u10_n19274 , _u10_n19273 , _u10_n19272 ,_u10_n19271 , _u10_n19270 , _u10_n19269 , _u10_n19268 , _u10_n19267 ,_u10_n19266 , _u10_n19265 , _u10_n19264 , _u10_n19263 , _u10_n19262 ,_u10_n19261 , _u10_n19260 , _u10_n19259 , _u10_n19258 , _u10_n19257 ,_u10_n19256 , _u10_n19255 , _u10_n19254 , _u10_n19253 , _u10_n19252 ,_u10_n19251 , _u10_n19250 , _u10_n19249 , _u10_n19248 , _u10_n19247 ,_u10_n19246 , _u10_n19245 , _u10_n19244 , _u10_n19243 , _u10_n19242 ,_u10_n19241 , _u10_n19240 , _u10_n19239 , _u10_n19238 , _u10_n19237 ,_u10_n19236 , _u10_n19235 , _u10_n19234 , _u10_n19233 , _u10_n19232 ,_u10_n19231 , _u10_n19230 , _u10_n19229 , _u10_n19228 , _u10_n19227 ,_u10_n19226 , _u10_n19225 , _u10_n19224 , _u10_n19223 , _u10_n19222 ,_u10_n19221 , _u10_n19220 , _u10_n19219 , _u10_n19218 , _u10_n19217 ,_u10_n19216 , _u10_n19215 , _u10_n19214 , _u10_n19213 , _u10_n19212 ,_u10_n19211 , _u10_n19210 , _u10_n19209 , _u10_n19208 , _u10_n19207 ,_u10_n19206 , _u10_n19205 , _u10_n19204 , _u10_n19203 , _u10_n19202 ,_u10_n19201 , _u10_n19200 , _u10_n19199 , _u10_n19198 , _u10_n19197 ,_u10_n19196 , _u10_n19195 , _u10_n19194 , _u10_n19193 , _u10_n19192 ,_u10_n19191 , _u10_n19190 , _u10_n19189 , _u10_n19188 , _u10_n19187 ,_u10_n19186 , _u10_n19185 , _u10_n19184 , _u10_n19183 , _u10_n19182 ,_u10_n19181 , _u10_n19180 , _u10_n19179 , _u10_n19178 , _u10_n19177 ,_u10_n19176 , _u10_n19175 , _u10_n19174 , _u10_n19173 , _u10_n19172 ,_u10_n19171 , _u10_n19170 , _u10_n19169 , _u10_n19168 , _u10_n19167 ,_u10_n19166 , _u10_n19165 , _u10_n19164 , _u10_n19163 , _u10_n19162 ,_u10_n19161 , _u10_n19160 , _u10_n19159 , _u10_n19158 , _u10_n19157 ,_u10_n19156 , _u10_n19155 , _u10_n19154 , _u10_n19153 , _u10_n19152 ,_u10_n19151 , _u10_n19150 , _u10_n19149 , _u10_n19148 , _u10_n19147 ,_u10_n19146 , _u10_n19145 , _u10_n19144 , _u10_n19143 , _u10_n19142 ,_u10_n19141 , _u10_n19140 , _u10_n19139 , _u10_n19138 , _u10_n19137 ,_u10_n19136 , _u10_n19135 , _u10_n19134 , _u10_n19133 , _u10_n19132 ,_u10_n19131 , _u10_n19130 , _u10_n19129 , _u10_n19128 , _u10_n19127 ,_u10_n19126 , _u10_n19125 , _u10_n19124 , _u10_n19123 , _u10_n19122 ,_u10_n19121 , _u10_n19120 , _u10_n19119 , _u10_n19118 , _u10_n19117 ,_u10_n19116 , _u10_n19115 , _u10_n19114 , _u10_n19113 , _u10_n19112 ,_u10_n19111 , _u10_n19110 , _u10_n19109 , _u10_n19108 , _u10_n19107 ,_u10_n19106 , _u10_n19105 , _u10_n19104 , _u10_n19103 , _u10_n19102 ,_u10_n19101 , _u10_n19100 , _u10_n19099 , _u10_n19098 , _u10_n19097 ,_u10_n19096 , _u10_n19095 , _u10_n19094 , _u10_n19093 , _u10_n19092 ,_u10_n19091 , _u10_n19090 , _u10_n19089 , _u10_n19088 , _u10_n19087 ,_u10_n19086 , _u10_n19085 , _u10_n19084 , _u10_n19083 , _u10_n19082 ,_u10_n19081 , _u10_n19080 , _u10_n19079 , _u10_n19078 , _u10_n19077 ,_u10_n19076 , _u10_n19075 , _u10_n19074 , _u10_n19073 , _u10_n19072 ,_u10_n19071 , _u10_n19070 , _u10_n19069 , _u10_n19068 , _u10_n19067 ,_u10_n19066 , _u10_n19065 , _u10_n19064 , _u10_n19063 , _u10_n19062 ,_u10_n19061 , _u10_n19060 , _u10_n19059 , _u10_n19058 , _u10_n19057 ,_u10_n19056 , _u10_n19055 , _u10_n19054 , _u10_n19053 , _u10_n19052 ,_u10_n19051 , _u10_n19050 , _u10_n19049 , _u10_n19048 , _u10_n19047 ,_u10_n19046 , _u10_n19045 , _u10_n19044 , _u10_n19043 , _u10_n19042 ,_u10_n19041 , _u10_n19040 , _u10_n19039 , _u10_n19038 , _u10_n19037 ,_u10_n19036 , _u10_n19035 , _u10_n19034 , _u10_n19033 , _u10_n19032 ,_u10_n19031 , _u10_n19030 , _u10_n19029 , _u10_n19028 , _u10_n19027 ,_u10_n19026 , _u10_n19025 , _u10_n19024 , _u10_n19023 , _u10_n19022 ,_u10_n19021 , _u10_n19020 , _u10_n19019 , _u10_n19018 , _u10_n19017 ,_u10_n19016 , _u10_n19015 , _u10_n19014 , _u10_n19013 , _u10_n19012 ,_u10_n19011 , _u10_n19010 , _u10_n19009 , _u10_n19008 , _u10_n19007 ,_u10_n19006 , _u10_n19005 , _u10_n19004 , _u10_n19003 , _u10_n19002 ,_u10_n19001 , _u10_n19000 , _u10_n18999 , _u10_n18998 , _u10_n18997 ,_u10_n18996 , _u10_n18995 , _u10_n18994 , _u10_n18993 , _u10_n18992 ,_u10_n18991 , _u10_n18990 , _u10_n18989 , _u10_n18988 , _u10_n18987 ,_u10_n18986 , _u10_n18985 , _u10_n18984 , _u10_n18983 , _u10_n18982 ,_u10_n18981 , _u10_n18980 , _u10_n18979 , _u10_n18978 , _u10_n18977 ,_u10_n18976 , _u10_n18975 , _u10_n18974 , _u10_n18973 , _u10_n18972 ,_u10_n18971 , _u10_n18970 , _u10_n18969 , _u10_n18968 , _u10_n18967 ,_u10_n18966 , _u10_n18965 , _u10_n18964 , _u10_n18963 , _u10_n18962 ,_u10_n18961 , _u10_n18960 , _u10_n18959 , _u10_n18958 , _u10_n18957 ,_u10_n18956 , _u10_n18955 , _u10_n18954 , _u10_n18953 , _u10_n18952 ,_u10_n18951 , _u10_n18950 , _u10_n18949 , _u10_n18948 , _u10_n18947 ,_u10_n18946 , _u10_n18945 , _u10_n18944 , _u10_n18943 , _u10_n18942 ,_u10_n18941 , _u10_n18940 , _u10_n18939 , _u10_n18938 , _u10_n18937 ,_u10_n18936 , _u10_n18935 , _u10_n18934 , _u10_n18933 , _u10_n18932 ,_u10_n18931 , _u10_n18930 , _u10_n18929 , _u10_n18928 , _u10_n18927 ,_u10_n18926 , _u10_n18925 , _u10_n18924 , _u10_n18923 , _u10_n18922 ,_u10_n18921 , _u10_n18920 , _u10_n18919 , _u10_n18918 , _u10_n18917 ,_u10_n18916 , _u10_n18915 , _u10_n18914 , _u10_n18913 , _u10_n18912 ,_u10_n18911 , _u10_n18910 , _u10_n18909 , _u10_n18908 , _u10_n18907 ,_u10_n18906 , _u10_n18905 , _u10_n18904 , _u10_n18903 , _u10_n18902 ,_u10_n18901 , _u10_n18900 , _u10_n18899 , _u10_n18898 , _u10_n18897 ,_u10_n18896 , _u10_n18895 , _u10_n18894 , _u10_n18893 , _u10_n18892 ,_u10_n18891 , _u10_n18890 , _u10_n18889 , _u10_n18888 , _u10_n18887 ,_u10_n18886 , _u10_n18885 , _u10_n18884 , _u10_n18883 , _u10_n18882 ,_u10_n18881 , _u10_n18880 , _u10_n18879 , _u10_n18878 , _u10_n18877 ,_u10_n18876 , _u10_n18875 , _u10_n18874 , _u10_n18873 , _u10_n18872 ,_u10_n18871 , _u10_n18870 , _u10_n18869 , _u10_n18868 , _u10_n18867 ,_u10_n18866 , _u10_n18865 , _u10_n18864 , _u10_n18863 , _u10_n18862 ,_u10_n18861 , _u10_n18860 , _u10_n18859 , _u10_n18858 , _u10_n18857 ,_u10_n18856 , _u10_n18855 , _u10_n18854 , _u10_n18853 , _u10_n18852 ,_u10_n18851 , _u10_n18850 , _u10_n18849 , _u10_n18848 , _u10_n18847 ,_u10_n18846 , _u10_n18845 , _u10_n18844 , _u10_n18843 , _u10_n18842 ,_u10_n18841 , _u10_n18840 , _u10_n18839 , _u10_n18838 , _u10_n18837 ,_u10_n18836 , _u10_n18835 , _u10_n18834 , _u10_n18833 , _u10_n18832 ,_u10_n18831 , _u10_n18830 , _u10_n18829 , _u10_n18828 , _u10_n18827 ,_u10_n18826 , _u10_n18825 , _u10_n18824 , _u10_n18823 , _u10_n18822 ,_u10_n18821 , _u10_n18820 , _u10_n18819 , _u10_n18818 , _u10_n18817 ,_u10_n18816 , _u10_n18815 , _u10_n18814 , _u10_n18813 , _u10_n18812 ,_u10_n18811 , _u10_n18810 , _u10_n18809 , _u10_n18808 , _u10_n18807 ,_u10_n18806 , _u10_n18805 , _u10_n18804 , _u10_n18803 , _u10_n18802 ,_u10_n18801 , _u10_n18800 , _u10_n18799 , _u10_n18798 , _u10_n18797 ,_u10_n18796 , _u10_n18795 , _u10_n18794 , _u10_n18793 , _u10_n18792 ,_u10_n18791 , _u10_n18790 , _u10_n18789 , _u10_n18788 , _u10_n18787 ,_u10_n18786 , _u10_n18785 , _u10_n18784 , _u10_n18783 , _u10_n18782 ,_u10_n18781 , _u10_n18780 , _u10_n18779 , _u10_n18778 , _u10_n18777 ,_u10_n18776 , _u10_n18775 , _u10_n18774 , _u10_n18773 , _u10_n18772 ,_u10_n18771 , _u10_n18770 , _u10_n18769 , _u10_n18768 , _u10_n18767 ,_u10_n18766 , _u10_n18765 , _u10_n18764 , _u10_n18763 , _u10_n18762 ,_u10_n18761 , _u10_n18760 , _u10_n18759 , _u10_n18758 , _u10_n18757 ,_u10_n18756 , _u10_n18755 , _u10_n18754 , _u10_n18753 , _u10_n18752 ,_u10_n18751 , _u10_n18750 , _u10_n18749 , _u10_n18748 , _u10_n18747 ,_u10_n18746 , _u10_n18745 , _u10_n18744 , _u10_n18743 , _u10_n18742 ,_u10_n18741 , _u10_n18740 , _u10_n18739 , _u10_n18738 , _u10_n18737 ,_u10_n18736 , _u10_n18735 , _u10_n18734 , _u10_n18733 , _u10_n18732 ,_u10_n18731 , _u10_n18730 , _u10_n18729 , _u10_n18728 , _u10_n18727 ,_u10_n18726 , _u10_n18725 , _u10_n18724 , _u10_n18723 , _u10_n18722 ,_u10_n18721 , _u10_n18720 , _u10_n18719 , _u10_n18718 , _u10_n18717 ,_u10_n18716 , _u10_n18715 , _u10_n18714 , _u10_n18713 , _u10_n18712 ,_u10_n18711 , _u10_n18710 , _u10_n18709 , _u10_n18708 , _u10_n18707 ,_u10_n18706 , _u10_n18705 , _u10_n18704 , _u10_n18703 , _u10_n18702 ,_u10_n18701 , _u10_n18700 , _u10_n18699 , _u10_n18698 , _u10_n18697 ,_u10_n18696 , _u10_n18695 , _u10_n18694 , _u10_n18693 , _u10_n18692 ,_u10_n18691 , _u10_n18690 , _u10_n18689 , _u10_n18688 , _u10_n18687 ,_u10_n18686 , _u10_n18685 , _u10_n18684 , _u10_n18683 , _u10_n18682 ,_u10_n18681 , _u10_n18680 , _u10_n18679 , _u10_n18678 , _u10_n18677 ,_u10_n18676 , _u10_n18675 , _u10_n18674 , _u10_n18673 , _u10_n18672 ,_u10_n18671 , _u10_n18670 , _u10_n18669 , _u10_n18668 , _u10_n18667 ,_u10_n18666 , _u10_n18665 , _u10_n18664 , _u10_n18663 , _u10_n18662 ,_u10_n18661 , _u10_n18660 , _u10_n18659 , _u10_n18658 , _u10_n18657 ,_u10_n18656 , _u10_n18655 , _u10_n18654 , _u10_n18653 , _u10_n18652 ,_u10_n18651 , _u10_n18650 , _u10_n18649 , _u10_n18648 , _u10_n18647 ,_u10_n18646 , _u10_n18645 , _u10_n18644 , _u10_n18643 , _u10_n18642 ,_u10_n18641 , _u10_n18640 , _u10_n18639 , _u10_n18638 , _u10_n18637 ,_u10_n18636 , _u10_n18635 , _u10_n18634 , _u10_n18633 , _u10_n18632 ,_u10_n18631 , _u10_n18630 , _u10_n18629 , _u10_n18628 , _u10_n18627 ,_u10_n18626 , _u10_n18625 , _u10_n18624 , _u10_n18623 , _u10_n18622 ,_u10_n18621 , _u10_n18620 , _u10_n18619 , _u10_n18618 , _u10_n18617 ,_u10_n18616 , _u10_n18615 , _u10_n18614 , _u10_n18613 , _u10_n18612 ,_u10_n18611 , _u10_n18610 , _u10_n18609 , _u10_n18608 , _u10_n18607 ,_u10_n18606 , _u10_n18605 , _u10_n18604 , _u10_n18603 , _u10_n18602 ,_u10_n18601 , _u10_n18600 , _u10_n18599 , _u10_n18598 , _u10_n18597 ,_u10_n18596 , _u10_n18595 , _u10_n18594 , _u10_n18593 , _u10_n18592 ,_u10_n18591 , _u10_n18590 , _u10_n18589 , _u10_n18588 , _u10_n18587 ,_u10_n18586 , _u10_n18585 , _u10_n18584 , _u10_n18583 , _u10_n18582 ,_u10_n18581 , _u10_n18580 , _u10_n18579 , _u10_n18578 , _u10_n18577 ,_u10_n18576 , _u10_n18575 , _u10_n18574 , _u10_n18573 , _u10_n18572 ,_u10_n18571 , _u10_n18570 , _u10_n18569 , _u10_n18568 , _u10_n18567 ,_u10_n18566 , _u10_n18565 , _u10_n18564 , _u10_n18563 , _u10_n18562 ,_u10_n18561 , _u10_n18560 , _u10_n18559 , _u10_n18558 , _u10_n18557 ,_u10_n18556 , _u10_n18555 , _u10_n18554 , _u10_n18553 , _u10_n18552 ,_u10_n18551 , _u10_n18550 , _u10_n18549 , _u10_n18548 , _u10_n18547 ,_u10_n18546 , _u10_n18545 , _u10_n18544 , _u10_n18543 , _u10_n18542 ,_u10_n18541 , _u10_n18540 , _u10_n18539 , _u10_n18538 , _u10_n18537 ,_u10_n18536 , _u10_n18535 , _u10_n18534 , _u10_n18533 , _u10_n18532 ,_u10_n18531 , _u10_n18530 , _u10_n18529 , _u10_n18528 , _u10_n18527 ,_u10_n18526 , _u10_n18525 , _u10_n18524 , _u10_n18523 , _u10_n18522 ,_u10_n18521 , _u10_n18520 , _u10_n18519 , _u10_n18518 , _u10_n18517 ,_u10_n18516 , _u10_n18515 , _u10_n18514 , _u10_n18513 , _u10_n18512 ,_u10_n18511 , _u10_n18510 , _u10_n18509 , _u10_n18508 , _u10_n18507 ,_u10_n18506 , _u10_n18505 , _u10_n18504 , _u10_n18503 , _u10_n18502 ,_u10_n18501 , _u10_n18500 , _u10_n18499 , _u10_n18498 , _u10_n18497 ,_u10_n18496 , _u10_n18495 , _u10_n18494 , _u10_n18493 , _u10_n18492 ,_u10_n18491 , _u10_n18490 , _u10_n18489 , _u10_n18488 , _u10_n18487 ,_u10_n18486 , _u10_n18485 , _u10_n18484 , _u10_n18483 , _u10_n18482 ,_u10_n18481 , _u10_n18480 , _u10_n18479 , _u10_n18478 , _u10_n18477 ,_u10_n18476 , _u10_n18475 , _u10_n18474 , _u10_n18473 , _u10_n18472 ,_u10_n18471 , _u10_n18470 , _u10_n18469 , _u10_n18468 , _u10_n18467 ,_u10_n18466 , _u10_n18465 , _u10_n18464 , _u10_n18463 , _u10_n18462 ,_u10_n18461 , _u10_n18460 , _u10_n18459 , _u10_n18458 , _u10_n18457 ,_u10_n18456 , _u10_n18455 , _u10_n18454 , _u10_n18453 , _u10_n18452 ,_u10_n18451 , _u10_n18450 , _u10_n18449 , _u10_n18448 , _u10_n18447 ,_u10_n18446 , _u10_n18445 , _u10_n18444 , _u10_n18443 , _u10_n18442 ,_u10_n18441 , _u10_n18440 , _u10_n18439 , _u10_n18438 , _u10_n18437 ,_u10_n18436 , _u10_n18435 , _u10_n18434 , _u10_n18433 , _u10_n18432 ,_u10_n18431 , _u10_n18430 , _u10_n18429 , _u10_n18428 , _u10_n18427 ,_u10_n18426 , _u10_n18425 , _u10_n18424 , _u10_n18423 , _u10_n18422 ,_u10_n18421 , _u10_n18420 , _u10_n18419 , _u10_n18418 , _u10_n18417 ,_u10_n18416 , _u10_n18415 , _u10_n18414 , _u10_n18413 , _u10_n18412 ,_u10_n18411 , _u10_n18410 , _u10_n18409 , _u10_n18408 , _u10_n18407 ,_u10_n18406 , _u10_n18405 , _u10_n18404 , _u10_n18403 , _u10_n18402 ,_u10_n18401 , _u10_n18400 , _u10_n18399 , _u10_n18398 , _u10_n18397 ,_u10_n18396 , _u10_n18395 , _u10_n18394 , _u10_n18393 , _u10_n18392 ,_u10_n18391 , _u10_n18390 , _u10_n18389 , _u10_n18388 , _u10_n18387 ,_u10_n18386 , _u10_n18385 , _u10_n18384 , _u10_n18383 , _u10_n18382 ,_u10_n18381 , _u10_n18380 , _u10_n18379 , _u10_n18378 , _u10_n18377 ,_u10_n18376 , _u10_n18375 , _u10_n18374 , _u10_n18373 , _u10_n18372 ,_u10_n18371 , _u10_n18370 , _u10_n18369 , _u10_n18368 , _u10_n18367 ,_u10_n18366 , _u10_n18365 , _u10_n18364 , _u10_n18363 , _u10_n18362 ,_u10_n18361 , _u10_n18360 , _u10_n18359 , _u10_n18358 , _u10_n18357 ,_u10_n18356 , _u10_n18355 , _u10_n18354 , _u10_n18353 , _u10_n18352 ,_u10_n18351 , _u10_n18350 , _u10_n18349 , _u10_n18348 , _u10_n18347 ,_u10_n18346 , _u10_n18345 , _u10_n18344 , _u10_n18343 , _u10_n18342 ,_u10_n18341 , _u10_n18340 , _u10_n18339 , _u10_n18338 , _u10_n18337 ,_u10_n18336 , _u10_n18335 , _u10_n18334 , _u10_n18333 , _u10_n18332 ,_u10_n18331 , _u10_n18330 , _u10_n18329 , _u10_n18328 , _u10_n18327 ,_u10_n18326 , _u10_n18325 , _u10_n18324 , _u10_n18323 , _u10_n18322 ,_u10_n18321 , _u10_n18320 , _u10_n18319 , _u10_n18318 , _u10_n18317 ,_u10_n18316 , _u10_n18315 , _u10_n18314 , _u10_n18313 , _u10_n18312 ,_u10_n18311 , _u10_n18310 , _u10_n18309 , _u10_n18308 , _u10_n18307 ,_u10_n18306 , _u10_n18305 , _u10_n18304 , _u10_n18303 , _u10_n18302 ,_u10_n18301 , _u10_n18300 , _u10_n18299 , _u10_n18298 , _u10_n18297 ,_u10_n18296 , _u10_n18295 , _u10_n18294 , _u10_n18293 , _u10_n18292 ,_u10_n18291 , _u10_n18290 , _u10_n18289 , _u10_n18288 , _u10_n18287 ,_u10_n18286 , _u10_n18285 , _u10_n18284 , _u10_n18283 , _u10_n18282 ,_u10_n18281 , _u10_n18280 , _u10_n18279 , _u10_n18278 , _u10_n18277 ,_u10_n18276 , _u10_n18275 , _u10_n18274 , _u10_n18273 , _u10_n18272 ,_u10_n18271 , _u10_n18270 , _u10_n18269 , _u10_n18268 , _u10_n18267 ,_u10_n18266 , _u10_n18265 , _u10_n18264 , _u10_n18263 , _u10_n18262 ,_u10_n18261 , _u10_n18260 , _u10_n18259 , _u10_n18258 , _u10_n18257 ,_u10_n18256 , _u10_n18255 , _u10_n18254 , _u10_n18253 , _u10_n18252 ,_u10_n18251 , _u10_n18250 , _u10_n18249 , _u10_n18248 , _u10_n18247 ,_u10_n18246 , _u10_n18245 , _u10_n18244 , _u10_n18243 , _u10_n18242 ,_u10_n18241 , _u10_n18240 , _u10_n18239 , _u10_n18238 , _u10_n18237 ,_u10_n18236 , _u10_n18235 , _u10_n18234 , _u10_n18233 , _u10_n18232 ,_u10_n18231 , _u10_n18230 , _u10_n18229 , _u10_n18228 , _u10_n18227 ,_u10_n18226 , _u10_n18225 , _u10_n18224 , _u10_n18223 , _u10_n18222 ,_u10_n18221 , _u10_n18220 , _u10_n18219 , _u10_n18218 , _u10_n18217 ,_u10_n18216 , _u10_n18215 , _u10_n18214 , _u10_n18213 , _u10_n18212 ,_u10_n18211 , _u10_n18210 , _u10_n18209 , _u10_n18208 , _u10_n18207 ,_u10_n18206 , _u10_n18205 , _u10_n18204 , _u10_n18203 , _u10_n18202 ,_u10_n18201 , _u10_n18200 , _u10_n18199 , _u10_n18198 , _u10_n18197 ,_u10_n18196 , _u10_n18195 , _u10_n18194 , _u10_n18193 , _u10_n18192 ,_u10_n18191 , _u10_n18190 , _u10_n18189 , _u10_n18188 , _u10_n18187 ,_u10_n18186 , _u10_n18185 , _u10_n18184 , _u10_n18183 , _u10_n18182 ,_u10_n18181 , _u10_n18180 , _u10_n18179 , _u10_n18178 , _u10_n18177 ,_u10_n18176 , _u10_n18175 , _u10_n18174 , _u10_n18173 , _u10_n18172 ,_u10_n18171 , _u10_n18170 , _u10_n18169 , _u10_n18168 , _u10_n18167 ,_u10_n18166 , _u10_n18165 , _u10_n18164 , _u10_n18163 , _u10_n18162 ,_u10_n18161 , _u10_n18160 , _u10_n18159 , _u10_n18158 , _u10_n18157 ,_u10_n18156 , _u10_n18155 , _u10_n18154 , _u10_n18153 , _u10_n18152 ,_u10_n18151 , _u10_n18150 , _u10_n18149 , _u10_n18148 , _u10_n18147 ,_u10_n18146 , _u10_n18145 , _u10_n18144 , _u10_n18143 , _u10_n18142 ,_u10_n18141 , _u10_n18140 , _u10_n18139 , _u10_n18138 , _u10_n18137 ,_u10_n18136 , _u10_n18135 , _u10_n18134 , _u10_n18133 , _u10_n18132 ,_u10_n18131 , _u10_n18130 , _u10_n18129 , _u10_n18128 , _u10_n18127 ,_u10_n18126 , _u10_n18125 , _u10_n18124 , _u10_n18123 , _u10_n18122 ,_u10_n18121 , _u10_n18120 , _u10_n18119 , _u10_n18118 , _u10_n18117 ,_u10_n18116 , _u10_n18115 , _u10_n18114 , _u10_n18113 , _u10_n18112 ,_u10_n18111 , _u10_n18110 , _u10_n18109 , _u10_n18108 , _u10_n18107 ,_u10_n18106 , _u10_n18105 , _u10_n18104 , _u10_n18103 , _u10_n18102 ,_u10_n18101 , _u10_n18100 , _u10_n18099 , _u10_n18098 , _u10_n18097 ,_u10_n18096 , _u10_n18095 , _u10_n18094 , _u10_n18093 , _u10_n18092 ,_u10_n18091 , _u10_n18090 , _u10_n18089 , _u10_n18088 , _u10_n18087 ,_u10_n18086 , _u10_n18085 , _u10_n18084 , _u10_n18083 , _u10_n18082 ,_u10_n18081 , _u10_n18080 , _u10_n18079 , _u10_n18078 , _u10_n18077 ,_u10_n18076 , _u10_n18075 , _u10_n18074 , _u10_n18073 , _u10_n18072 ,_u10_n18071 , _u10_n18070 , _u10_n18069 , _u10_n18068 , _u10_n18067 ,_u10_n18066 , _u10_n18065 , _u10_n18064 , _u10_n18063 , _u10_n18062 ,_u10_n18061 , _u10_n18060 , _u10_n18059 , _u10_n18058 , _u10_n18057 ,_u10_n18056 , _u10_n18055 , _u10_n18054 , _u10_n18053 , _u10_n18052 ,_u10_n18051 , _u10_n18050 , _u10_n18049 , _u10_n18048 , _u10_n18047 ,_u10_n18046 , _u10_n18045 , _u10_n18044 , _u10_n18043 , _u10_n18042 ,_u10_n18041 , _u10_n18040 , _u10_n18039 , _u10_n18038 , _u10_n18037 ,_u10_n18036 , _u10_n18035 , _u10_n18034 , _u10_n18033 , _u10_n18032 ,_u10_n18031 , _u10_n18030 , _u10_n18029 , _u10_n18028 , _u10_n18027 ,_u10_n18026 , _u10_n18025 , _u10_n18024 , _u10_n18023 , _u10_n18022 ,_u10_n18021 , _u10_n18020 , _u10_n18019 , _u10_n18018 , _u10_n18017 ,_u10_n18016 , _u10_n18015 , _u10_n18014 , _u10_n18013 , _u10_n18012 ,_u10_n18011 , _u10_n18010 , _u10_n18009 , _u10_n18008 , _u10_n18007 ,_u10_n18006 , _u10_n18005 , _u10_n18004 , _u10_n18003 , _u10_n18002 ,_u10_n18001 , _u10_n18000 , _u10_n17999 , _u10_n17998 , _u10_n17997 ,_u10_n17996 , _u10_n17995 , _u10_n17994 , _u10_n17993 , _u10_n17992 ,_u10_n17991 , _u10_n17990 , _u10_n17989 , _u10_n17988 , _u10_n17987 ,_u10_n17986 , _u10_n17985 , _u10_n17984 , _u10_n17983 , _u10_n17982 ,_u10_n17981 , _u10_n17980 , _u10_n17979 , _u10_n17978 , _u10_n17977 ,_u10_n17976 , _u10_n17975 , _u10_n17974 , _u10_n17973 , _u10_n17972 ,_u10_n17971 , _u10_n17970 , _u10_n17969 , _u10_n17968 , _u10_n17967 ,_u10_n17966 , _u10_n17965 , _u10_n17964 , _u10_n17963 , _u10_n17962 ,_u10_n17961 , _u10_n17960 , _u10_n17959 , _u10_n17958 , _u10_n17957 ,_u10_n17956 , _u10_n17955 , _u10_n17954 , _u10_n17953 , _u10_n17952 ,_u10_n17951 , _u10_n17950 , _u10_n17949 , _u10_n17948 , _u10_n17947 ,_u10_n17946 , _u10_n17945 , _u10_n17944 , _u10_n17943 , _u10_n17942 ,_u10_n17941 , _u10_n17940 , _u10_n17939 , _u10_n17938 , _u10_n17937 ,_u10_n17936 , _u10_n17935 , _u10_n17934 , _u10_n17933 , _u10_n17932 ,_u10_n17931 , _u10_n17930 , _u10_n17929 , _u10_n17928 , _u10_n17927 ,_u10_n17926 , _u10_n17925 , _u10_n17924 , _u10_n17923 , _u10_n17922 ,_u10_n17921 , _u10_n17920 , _u10_n17919 , _u10_n17918 , _u10_n17917 ,_u10_n17916 , _u10_n17915 , _u10_n17914 , _u10_n17913 , _u10_n17912 ,_u10_n17911 , _u10_n17910 , _u10_n17909 , _u10_n17908 , _u10_n17907 ,_u10_n17906 , _u10_n17905 , _u10_n17904 , _u10_n17903 , _u10_n17902 ,_u10_n17901 , _u10_n17900 , _u10_n17899 , _u10_n17898 , _u10_n17897 ,_u10_n17896 , _u10_n17895 , _u10_n17894 , _u10_n17893 , _u10_n17892 ,_u10_n17891 , _u10_n17890 , _u10_n17889 , _u10_n17888 , _u10_n17887 ,_u10_n17886 , _u10_n17885 , _u10_n17884 , _u10_n17883 , _u10_n17882 ,_u10_n17881 , _u10_n17880 , _u10_n17879 , _u10_n17878 , _u10_n17877 ,_u10_n17876 , _u10_n17875 , _u10_n17874 , _u10_n17873 , _u10_n17872 ,_u10_n17871 , _u10_n17870 , _u10_n17869 , _u10_n17868 , _u10_n17867 ,_u10_n17866 , _u10_n17865 , _u10_n17864 , _u10_n17863 , _u10_n17862 ,_u10_n17861 , _u10_n17860 , _u10_n17859 , _u10_n17858 , _u10_n17857 ,_u10_n17856 , _u10_n17855 , _u10_n17854 , _u10_n17853 , _u10_n17852 ,_u10_n17851 , _u10_n17850 , _u10_n17849 , _u10_n17848 , _u10_n17847 ,_u10_n17846 , _u10_n17845 , _u10_n17844 , _u10_n17843 , _u10_n17842 ,_u10_n17841 , _u10_n17840 , _u10_n17839 , _u10_n17838 , _u10_n17837 ,_u10_n17836 , _u10_n17835 , _u10_n17834 , _u10_n17833 , _u10_n17832 ,_u10_n17831 , _u10_n17830 , _u10_n17829 , _u10_n17828 , _u10_n17827 ,_u10_n17826 , _u10_n17825 , _u10_n17824 , _u10_n17823 , _u10_n17822 ,_u10_n17821 , _u10_n17820 , _u10_n17819 , _u10_n17818 , _u10_n17817 ,_u10_n17816 , _u10_n17815 , _u10_n17814 , _u10_n17813 , _u10_n17812 ,_u10_n17811 , _u10_n17810 , _u10_n17809 , _u10_n17808 , _u10_n17807 ,_u10_n17806 , _u10_n17805 , _u10_n17804 , _u10_n17803 , _u10_n17802 ,_u10_n17801 , _u10_n17800 , _u10_n17799 , _u10_n17798 , _u10_n17797 ,_u10_n17796 , _u10_n17795 , _u10_n17794 , _u10_n17793 , _u10_n17792 ,_u10_n17791 , _u10_n17790 , _u10_n17789 , _u10_n17788 , _u10_n17787 ,_u10_n17786 , _u10_n17785 , _u10_n17784 , _u10_n17783 , _u10_n17782 ,_u10_n17781 , _u10_n17780 , _u10_n17779 , _u10_n17778 , _u10_n17777 ,_u10_n17776 , _u10_n17775 , _u10_n17774 , _u10_n17773 , _u10_n17772 ,_u10_n17771 , _u10_n17770 , _u10_n17769 , _u10_n17768 , _u10_n17767 ,_u10_n17766 , _u10_n17765 , _u10_n17764 , _u10_n17763 , _u10_n17762 ,_u10_n17761 , _u10_n17760 , _u10_n17759 , _u10_n17758 , _u10_n17757 ,_u10_n17756 , _u10_n17755 , _u10_n17754 , _u10_n17753 , _u10_n17752 ,_u10_n17751 , _u10_n17750 , _u10_n17749 , _u10_n17748 , _u10_n17747 ,_u10_n17746 , _u10_n17745 , _u10_n17744 , _u10_n17743 , _u10_n17742 ,_u10_n17741 , _u10_n17740 , _u10_n17739 , _u10_n17738 , _u10_n17737 ,_u10_n17736 , _u10_n17735 , _u10_n17734 , _u10_n17733 , _u10_n17732 ,_u10_n17731 , _u10_n17730 , _u10_n17729 , _u10_n17728 , _u10_n17727 ,_u10_n17726 , _u10_n17725 , _u10_n17724 , _u10_n17723 , _u10_n17722 ,_u10_n17721 , _u10_n17720 , _u10_n17719 , _u10_n17718 , _u10_n17717 ,_u10_n17716 , _u10_n17715 , _u10_n17714 , _u10_n17713 , _u10_n17712 ,_u10_n17711 , _u10_n17710 , _u10_n17709 , _u10_n17708 , _u10_n17707 ,_u10_n17706 , _u10_n17705 , _u10_n17704 , _u10_n17703 , _u10_n17702 ,_u10_n17701 , _u10_n17700 , _u10_n17699 , _u10_n17698 , _u10_n17697 ,_u10_n17696 , _u10_n17695 , _u10_n17694 , _u10_n17693 , _u10_n17692 ,_u10_n17691 , _u10_n17690 , _u10_n17689 , _u10_n17688 , _u10_n17687 ,_u10_n17686 , _u10_n17685 , _u10_n17684 , _u10_n17683 , _u10_n17682 ,_u10_n17681 , _u10_n17680 , _u10_n17679 , _u10_n17678 , _u10_n17677 ,_u10_n17676 , _u10_n17675 , _u10_n17674 , _u10_n17673 , _u10_n17672 ,_u10_n17671 , _u10_n17670 , _u10_n17669 , _u10_n17668 , _u10_n17667 ,_u10_n17666 , _u10_n17665 , _u10_n17664 , _u10_n17663 , _u10_n17662 ,_u10_n17661 , _u10_n17660 , _u10_n17659 , _u10_n17658 , _u10_n17657 ,_u10_n17656 , _u10_n17655 , _u10_n17654 , _u10_n17653 , _u10_n17652 ,_u10_n17651 , _u10_n17650 , _u10_n17649 , _u10_n17648 , _u10_n17647 ,_u10_n17646 , _u10_n17645 , _u10_n17644 , _u10_n17643 , _u10_n17642 ,_u10_n17641 , _u10_n17640 , _u10_n17639 , _u10_n17638 , _u10_n17637 ,_u10_n17636 , _u10_n17635 , _u10_n17634 , _u10_n17633 , _u10_n17632 ,_u10_n17631 , _u10_n17630 , _u10_n17629 , _u10_n17628 , _u10_n17627 ,_u10_n17626 , _u10_n17625 , _u10_n17624 , _u10_n17623 , _u10_n17622 ,_u10_n17621 , _u10_n17620 , _u10_n17619 , _u10_n17618 , _u10_n17617 ,_u10_n17616 , _u10_n17615 , _u10_n17614 , _u10_n17613 , _u10_n17612 ,_u10_n17611 , _u10_n17610 , _u10_n17609 , _u10_n17608 , _u10_n17607 ,_u10_n17606 , _u10_n17605 , _u10_n17604 , _u10_n17603 , _u10_n17602 ,_u10_n17601 , _u10_n17600 , _u10_n17599 , _u10_n17598 , _u10_n17597 ,_u10_n17596 , _u10_n17595 , _u10_n17594 , _u10_n17593 , _u10_n17592 ,_u10_n17591 , _u10_n17590 , _u10_n17589 , _u10_n17588 , _u10_n17587 ,_u10_n17586 , _u10_n17585 , _u10_n17584 , _u10_n17583 , _u10_n17582 ,_u10_n17581 , _u10_n17580 , _u10_n17579 , _u10_n17578 , _u10_n17577 ,_u10_n17576 , _u10_n17575 , _u10_n17574 , _u10_n17573 , _u10_n17572 ,_u10_n17571 , _u10_n17570 , _u10_n17569 , _u10_n17568 , _u10_n17567 ,_u10_n17566 , _u10_n17565 , _u10_n17564 , _u10_n17563 , _u10_n17562 ,_u10_n17561 , _u10_n17560 , _u10_n17559 , _u10_n17558 , _u10_n17557 ,_u10_n17556 , _u10_n17555 , _u10_n17554 , _u10_n17553 , _u10_n17552 ,_u10_n17551 , _u10_n17550 , _u10_n17549 , _u10_n17548 , _u10_n17547 ,_u10_n17546 , _u10_n17545 , _u10_n17544 , _u10_n17543 , _u10_n17542 ,_u10_n17541 , _u10_n17540 , _u10_n17539 , _u10_n17538 , _u10_n17537 ,_u10_n17536 , _u10_n17535 , _u10_n17534 , _u10_n17533 , _u10_n17532 ,_u10_n17531 , _u10_n17530 , _u10_n17529 , _u10_n17528 , _u10_n17527 ,_u10_n17526 , _u10_n17525 , _u10_n17524 , _u10_n17523 , _u10_n17522 ,_u10_n17521 , _u10_n17520 , _u10_n17519 , _u10_n17518 , _u10_n17517 ,_u10_n17516 , _u10_n17515 , _u10_n17514 , _u10_n17513 , _u10_n17512 ,_u10_n17511 , _u10_n17510 , _u10_n17509 , _u10_n17508 , _u10_n17507 ,_u10_n17506 , _u10_n17505 , _u10_n17504 , _u10_n17503 , _u10_n17502 ,_u10_n17501 , _u10_n17500 , _u10_n17499 , _u10_n17498 , _u10_n17497 ,_u10_n17496 , _u10_n17495 , _u10_n17494 , _u10_n17493 , _u10_n17492 ,_u10_n17491 , _u10_n17490 , _u10_n17489 , _u10_n17488 , _u10_n17487 ,_u10_n17486 , _u10_n17485 , _u10_n17484 , _u10_n17483 , _u10_n17482 ,_u10_n17481 , _u10_n17480 , _u10_n17479 , _u10_n17478 , _u10_n17477 ,_u10_n17476 , _u10_n17475 , _u10_n17474 , _u10_n17473 , _u10_n17472 ,_u10_n17471 , _u10_n17470 , _u10_n17469 , _u10_n17468 , _u10_n17467 ,_u10_n17466 , _u10_n17465 , _u10_n17464 , _u10_n17463 , _u10_n17462 ,_u10_n17461 , _u10_n17460 , _u10_n17459 , _u10_n17458 , _u10_n17457 ,_u10_n17456 , _u10_n17455 , _u10_n17454 , _u10_n17453 , _u10_n17452 ,_u10_n17451 , _u10_n17450 , _u10_n17449 , _u10_n17448 , _u10_n17447 ,_u10_n17446 , _u10_n17445 , _u10_n17444 , _u10_n17443 , _u10_n17442 ,_u10_n17441 , _u10_n17440 , _u10_n17439 , _u10_n17438 , _u10_n17437 ,_u10_n17436 , _u10_n17435 , _u10_n17434 , _u10_n17433 , _u10_n17432 ,_u10_n17431 , _u10_n17430 , _u10_n17429 , _u10_n17428 , _u10_n17427 ,_u10_n17426 , _u10_n17425 , _u10_n17424 , _u10_n17423 , _u10_n17422 ,_u10_n17421 , _u10_n17420 , _u10_n17419 , _u10_n17418 , _u10_n17417 ,_u10_n17416 , _u10_n17415 , _u10_n17414 , _u10_n17413 , _u10_n17412 ,_u10_n17411 , _u10_n17410 , _u10_n17409 , _u10_n17408 , _u10_n17407 ,_u10_n17406 , _u10_n17405 , _u10_n17404 , _u10_n17403 , _u10_n17402 ,_u10_n17401 , _u10_n17400 , _u10_n17399 , _u10_n17398 , _u10_n17397 ,_u10_n17396 , _u10_n17395 , _u10_n17394 , _u10_n17393 , _u10_n17392 ,_u10_n17391 , _u10_n17390 , _u10_n17389 , _u10_n17388 , _u10_n17387 ,_u10_n17386 , _u10_n17385 , _u10_n17384 , _u10_n17383 , _u10_n17382 ,_u10_n17381 , _u10_n17380 , _u10_n17379 , _u10_n17378 , _u10_n17377 ,_u10_n17376 , _u10_n17375 , _u10_n17374 , _u10_n17373 , _u10_n17372 ,_u10_n17371 , _u10_n17370 , _u10_n17369 , _u10_n17368 , _u10_n17367 ,_u10_n17366 , _u10_n17365 , _u10_n17364 , _u10_n17363 , _u10_n17362 ,_u10_n17361 , _u10_n17360 , _u10_n17359 , _u10_n17358 , _u10_n17357 ,_u10_n17356 , _u10_n17355 , _u10_n17354 , _u10_n17353 , _u10_n17352 ,_u10_n17351 , _u10_n17350 , _u10_n17349 , _u10_n17348 , _u10_n17347 ,_u10_n17346 , _u10_n17345 , _u10_n17344 , _u10_n17343 , _u10_n17342 ,_u10_n17341 , _u10_n17340 , _u10_n17339 , _u10_n17338 , _u10_n17337 ,_u10_n17336 , _u10_n17335 , _u10_n17334 , _u10_n17333 , _u10_n17332 ,_u10_n17331 , _u10_n17330 , _u10_n17329 , _u10_n17328 , _u10_n17327 ,_u10_n17326 , _u10_n17325 , _u10_n17324 , _u10_n17323 , _u10_n17322 ,_u10_n17321 , _u10_n17320 , _u10_n17319 , _u10_n17318 , _u10_n17317 ,_u10_n17316 , _u10_n17315 , _u10_n17314 , _u10_n17313 , _u10_n17312 ,_u10_n17311 , _u10_n17310 , _u10_n17309 , _u10_n17308 , _u10_n17307 ,_u10_n17306 , _u10_n17305 , _u10_n17304 , _u10_n17303 , _u10_n17302 ,_u10_n17301 , _u10_n17300 , _u10_n17299 , _u10_n17298 , _u10_n17297 ,_u10_n17296 , _u10_n17295 , _u10_n17294 , _u10_n17293 , _u10_n17292 ,_u10_n17291 , _u10_n17290 , _u10_n17289 , _u10_n17288 , _u10_n17287 ,_u10_n17286 , _u10_n17285 , _u10_n17284 , _u10_n17283 , _u10_n17282 ,_u10_n17281 , _u10_n17280 , _u10_n17279 , _u10_n17278 , _u10_n17277 ,_u10_n17276 , _u10_n17275 , _u10_n17274 , _u10_n17273 , _u10_n17272 ,_u10_n17271 , _u10_n17270 , _u10_n17269 , _u10_n17268 , _u10_n17267 ,_u10_n17266 , _u10_n17265 , _u10_n17264 , _u10_n17263 , _u10_n17262 ,_u10_n17261 , _u10_n17260 , _u10_n17259 , _u10_n17258 , _u10_n17257 ,_u10_n17256 , _u10_n17255 , _u10_n17254 , _u10_n17253 , _u10_n17252 ,_u10_n17251 , _u10_n17250 , _u10_n17249 , _u10_n17248 , _u10_n17247 ,_u10_n17246 , _u10_n17245 , _u10_n17244 , _u10_n17243 , _u10_n17242 ,_u10_n17241 , _u10_n17240 , _u10_n17239 , _u10_n17238 , _u10_n17237 ,_u10_n17236 , _u10_n17235 , _u10_n17234 , _u10_n17233 , _u10_n17232 ,_u10_n17231 , _u10_n17230 , _u10_n17229 , _u10_n17228 , _u10_n17227 ,_u10_n17226 , _u10_n17225 , _u10_n17224 , _u10_n17223 , _u10_n17222 ,_u10_n17221 , _u10_n17220 , _u10_n17219 , _u10_n17218 , _u10_n17217 ,_u10_n17216 , _u10_n17215 , _u10_n17214 , _u10_n17213 , _u10_n17212 ,_u10_n17211 , _u10_n17210 , _u10_n17209 , _u10_n17208 , _u10_n17207 ,_u10_n17206 , _u10_n17205 , _u10_n17204 , _u10_n17203 , _u10_n17202 ,_u10_n17201 , _u10_n17200 , _u10_n17199 , _u10_n17198 , _u10_n17197 ,_u10_n17196 , _u10_n17195 , _u10_n17194 , _u10_n17193 , _u10_n17192 ,_u10_n17191 , _u10_n17190 , _u10_n17189 , _u10_n17188 , _u10_n17187 ,_u10_n17186 , _u10_n17185 , _u10_n17184 , _u10_n17183 , _u10_n17182 ,_u10_n17181 , _u10_n17180 , _u10_n17179 , _u10_n17178 , _u10_n17177 ,_u10_n17176 , _u10_n17175 , _u10_n17174 , _u10_n17173 , _u10_n17172 ,_u10_n17171 , _u10_n17170 , _u10_n17169 , _u10_n17168 , _u10_n17167 ,_u10_n17166 , _u10_n17165 , _u10_n17164 , _u10_n17163 , _u10_n17162 ,_u10_n17161 , _u10_n17160 , _u10_n17159 , _u10_n17158 , _u10_n17157 ,_u10_n17156 , _u10_n17155 , _u10_n17154 , _u10_n17153 , _u10_n17152 ,_u10_n17151 , _u10_n17150 , _u10_n17149 , _u10_n17148 , _u10_n17147 ,_u10_n17146 , _u10_n17145 , _u10_n17144 , _u10_n17143 , _u10_n17142 ,_u10_n17141 , _u10_n17140 , _u10_n17139 , _u10_n17138 , _u10_n17137 ,_u10_n17136 , _u10_n17135 , _u10_n17134 , _u10_n17133 , _u10_n17132 ,_u10_n17131 , _u10_n17130 , _u10_n17129 , _u10_n17128 , _u10_n17127 ,_u10_n17126 , _u10_n17125 , _u10_n17124 , _u10_n17123 , _u10_n17122 ,_u10_n17121 , _u10_n17120 , _u10_n17119 , _u10_n17118 , _u10_n17117 ,_u10_n17116 , _u10_n17115 , _u10_n17114 , _u10_n17113 , _u10_n17112 ,_u10_n17111 , _u10_n17110 , _u10_n17109 , _u10_n17108 , _u10_n17107 ,_u10_n17106 , _u10_n17105 , _u10_n17104 , _u10_n17103 , _u10_n17102 ,_u10_n17101 , _u10_n17100 , _u10_n17099 , _u10_n17098 , _u10_n17097 ,_u10_n17096 , _u10_n17095 , _u10_n17094 , _u10_n17093 , _u10_n17092 ,_u10_n17091 , _u10_n17090 , _u10_n17089 , _u10_n17088 , _u10_n17087 ,_u10_n17086 , _u10_n17085 , _u10_n17084 , _u10_n17083 , _u10_n17082 ,_u10_n17081 , _u10_n17080 , _u10_n17079 , _u10_n17078 , _u10_n17077 ,_u10_n17076 , _u10_n17075 , _u10_n17074 , _u10_n17073 , _u10_n17072 ,_u10_n17071 , _u10_n17070 , _u10_n17069 , _u10_n17068 , _u10_n17067 ,_u10_n17066 , _u10_n17065 , _u10_n17064 , _u10_n17063 , _u10_n17062 ,_u10_n17061 , _u10_n17060 , _u10_n17059 , _u10_n17058 , _u10_n17057 ,_u10_n17056 , _u10_n17055 , _u10_n17054 , _u10_n17053 , _u10_n17052 ,_u10_n17051 , _u10_n17050 , _u10_n17049 , _u10_n17048 , _u10_n17047 ,_u10_n17046 , _u10_n17045 , _u10_n17044 , _u10_n17043 , _u10_n17042 ,_u10_n17041 , _u10_n17040 , _u10_n17039 , _u10_n17038 , _u10_n17037 ,_u10_n17036 , _u10_n17035 , _u10_n17034 , _u10_n17033 , _u10_n17032 ,_u10_n17031 , _u10_n17030 , _u10_n17029 , _u10_n17028 , _u10_n17027 ,_u10_n17026 , _u10_n17025 , _u10_n17024 , _u10_n17023 , _u10_n17022 ,_u10_n17021 , _u10_n17020 , _u10_n17019 , _u10_n17018 , _u10_n17017 ,_u10_n17016 , _u10_n17015 , _u10_n17014 , _u10_n17013 , _u10_n17012 ,_u10_n17011 , _u10_n17010 , _u10_n17009 , _u10_n17008 , _u10_n17007 ,_u10_n17006 , _u10_n17005 , _u10_n17004 , _u10_n17003 , _u10_n17002 ,_u10_n17001 , _u10_n17000 , _u10_n16999 , _u10_n16998 , _u10_n16997 ,_u10_n16996 , _u10_n16995 , _u10_n16994 , _u10_n16993 , _u10_n16992 ,_u10_n16991 , _u10_n16990 , _u10_n16989 , _u10_n16988 , _u10_n16987 ,_u10_n16986 , _u10_n16985 , _u10_n16984 , _u10_n16983 , _u10_n16982 ,_u10_n16981 , _u10_n16980 , _u10_n16979 , _u10_n16978 , _u10_n16977 ,_u10_n16976 , _u10_n16975 , _u10_n16974 , _u10_n16973 , _u10_n16972 ,_u10_n16971 , _u10_n16970 , _u10_n16969 , _u10_n16968 , _u10_n16967 ,_u10_n16966 , _u10_n16965 , _u10_n16964 , _u10_n16963 , _u10_n16962 ,_u10_n16961 , _u10_n16960 , _u10_n16959 , _u10_n16958 , _u10_n16957 ,_u10_n16956 , _u10_n16955 , _u10_n16954 , _u10_n16953 , _u10_n16952 ,_u10_n16951 , _u10_n16950 , _u10_n16949 , _u10_n16948 , _u10_n16947 ,_u10_n16946 , _u10_n16945 , _u10_n16944 , _u10_n16943 , _u10_n16942 ,_u10_n16941 , _u10_n16940 , _u10_n16939 , _u10_n16938 , _u10_n16937 ,_u10_n16936 , _u10_n16935 , _u10_n16934 , _u10_n16933 , _u10_n16932 ,_u10_n16931 , _u10_n16930 , _u10_n16929 , _u10_n16928 , _u10_n16927 ,_u10_n16926 , _u10_n16925 , _u10_n16924 , _u10_n16923 , _u10_n16922 ,_u10_n16921 , _u10_n16920 , _u10_n16919 , _u10_n16918 , _u10_n16917 ,_u10_n16916 , _u10_n16915 , _u10_n16914 , _u10_n16913 , _u10_n16912 ,_u10_n16911 , _u10_n16910 , _u10_n16909 , _u10_n16908 , _u10_n16907 ,_u10_n16906 , _u10_n16905 , _u10_n16904 , _u10_n16903 , _u10_n16902 ,_u10_n16901 , _u10_n16900 , _u10_n16899 , _u10_n16898 , _u10_n16897 ,_u10_n16896 , _u10_n16895 , _u10_n16894 , _u10_n16893 , _u10_n16892 ,_u10_n16891 , _u10_n16890 , _u10_n16889 , _u10_n16888 , _u10_n16887 ,_u10_n16886 , _u10_n16885 , _u10_n16884 , _u10_n16883 , _u10_n16882 ,_u10_n16881 , _u10_n16880 , _u10_n16879 , _u10_n16878 , _u10_n16877 ,_u10_n16876 , _u10_n16875 , _u10_n16874 , _u10_n16873 , _u10_n16872 ,_u10_n16871 , _u10_n16870 , _u10_n16869 , _u10_n16868 , _u10_n16867 ,_u10_n16866 , _u10_n16865 , _u10_n16864 , _u10_n16863 , _u10_n16862 ,_u10_n16861 , _u10_n16860 , _u10_n16859 , _u10_n16858 , _u10_n16857 ,_u10_n16856 , _u10_n16855 , _u10_n16854 , _u10_n16853 , _u10_n16852 ,_u10_n16851 , _u10_n16850 , _u10_n16849 , _u10_n16848 , _u10_n16847 ,_u10_n16846 , _u10_n16845 , _u10_n16844 , _u10_n16843 , _u10_n16842 ,_u10_n16841 , _u10_n16840 , _u10_n16839 , _u10_n16838 , _u10_n16837 ,_u10_n16836 , _u10_n16835 , _u10_n16834 , _u10_n16833 , _u10_n16832 ,_u10_n16831 , _u10_n16830 , _u10_n16829 , _u10_n16828 , _u10_n16827 ,_u10_n16826 , _u10_n16825 , _u10_n16824 , _u10_n16823 , _u10_n16822 ,_u10_n16821 , _u10_n16820 , _u10_n16819 , _u10_n16818 , _u10_n16817 ,_u10_n16816 , _u10_n16815 , _u10_n16814 , _u10_n16813 , _u10_n16812 ,_u10_n16811 , _u10_n16810 , _u10_n16809 , _u10_n16808 , _u10_n16807 ,_u10_n16806 , _u10_n16805 , _u10_n16804 , _u10_n16803 , _u10_n16802 ,_u10_n16801 , _u10_n16800 , _u10_n16799 , _u10_n16798 , _u10_n16797 ,_u10_n16796 , _u10_n16795 , _u10_n16794 , _u10_n16793 , _u10_n16792 ,_u10_n16791 , _u10_n16790 , _u10_n16789 , _u10_n16788 , _u10_n16787 ,_u10_n16786 , _u10_n16785 , _u10_n16784 , _u10_n16783 , _u10_n16782 ,_u10_n16781 , _u10_n16780 , _u10_n16779 , _u10_n16778 , _u10_n16777 ,_u10_n16776 , _u10_n16775 , _u10_n16774 , _u10_n16773 , _u10_n16772 ,_u10_n16771 , _u10_n16770 , _u10_n16769 , _u10_n16768 , _u10_n16767 ,_u10_n16766 , _u10_n16765 , _u10_n16764 , _u10_n16763 , _u10_n16762 ,_u10_n16761 , _u10_n16760 , _u10_n16759 , _u10_n16758 , _u10_n16757 ,_u10_n16756 , _u10_n16755 , _u10_n16754 , _u10_n16753 , _u10_n16752 ,_u10_n16751 , _u10_n16750 , _u10_n16749 , _u10_n16748 , _u10_n16747 ,_u10_n16746 , _u10_n16745 , _u10_n16744 , _u10_n16743 , _u10_n16742 ,_u10_n16741 , _u10_n16740 , _u10_n16739 , _u10_n16738 , _u10_n16737 ,_u10_n16736 , _u10_n16735 , _u10_n16734 , _u10_n16733 , _u10_n16732 ,_u10_n16731 , _u10_n16730 , _u10_n16729 , _u10_n16728 , _u10_n16727 ,_u10_n16726 , _u10_n16725 , _u10_n16724 , _u10_n16723 , _u10_n16722 ,_u10_n16721 , _u10_n16720 , _u10_n16719 , _u10_n16718 , _u10_n16717 ,_u10_n16716 , _u10_n16715 , _u10_n16714 , _u10_n16713 , _u10_n16712 ,_u10_n16711 , _u10_n16710 , _u10_n16709 , _u10_n16708 , _u10_n16707 ,_u10_n16706 , _u10_n16705 , _u10_n16704 , _u10_n16703 , _u10_n16702 ,_u10_n16701 , _u10_n16700 , _u10_n16699 , _u10_n16698 , _u10_n16697 ,_u10_n16696 , _u10_n16695 , _u10_n16694 , _u10_n16693 , _u10_n16692 ,_u10_n16691 , _u10_n16690 , _u10_n16689 , _u10_n16688 , _u10_n16687 ,_u10_n16686 , _u10_n16685 , _u10_n16684 , _u10_n16683 , _u10_n16682 ,_u10_n16681 , _u10_n16680 , _u10_n16679 , _u10_n16678 , _u10_n16677 ,_u10_n16676 , _u10_n16675 , _u10_n16674 , _u10_n16673 , _u10_n16672 ,_u10_n16671 , _u10_n16670 , _u10_n16669 , _u10_n16668 , _u10_n16667 ,_u10_n16666 , _u10_n16665 , _u10_n16664 , _u10_n16663 , _u10_n16662 ,_u10_n16661 , _u10_n16660 , _u10_n16659 , _u10_n16658 , _u10_n16657 ,_u10_n16656 , _u10_n16655 , _u10_n16654 , _u10_n16653 , _u10_n16652 ,_u10_n16651 , _u10_n16650 , _u10_n16649 , _u10_n16648 , _u10_n16647 ,_u10_n16646 , _u10_n16645 , _u10_n16644 , _u10_n16643 , _u10_n16642 ,_u10_n16641 , _u10_n16640 , _u10_n16639 , _u10_n16638 , _u10_n16637 ,_u10_n16636 , _u10_n16635 , _u10_n16634 , _u10_n16633 , _u10_n16632 ,_u10_n16631 , _u10_n16630 , _u10_n16629 , _u10_n16628 , _u10_n16627 ,_u10_n16626 , _u10_n16625 , _u10_n16624 , _u10_n16623 , _u10_n16622 ,_u10_n16621 , _u10_n16620 , _u10_n16619 , _u10_n16618 , _u10_n16617 ,_u10_n16616 , _u10_n16615 , _u10_n16614 , _u10_n16613 , _u10_n16612 ,_u10_n16611 , _u10_n16610 , _u10_n16609 , _u10_n16608 , _u10_n16607 ,_u10_n16606 , _u10_n16605 , _u10_n16604 , _u10_n16603 , _u10_n16602 ,_u10_n16601 , _u10_n16600 , _u10_n16599 , _u10_n16598 , _u10_n16597 ,_u10_n16596 , _u10_n16595 , _u10_n16594 , _u10_n16593 , _u10_n16592 ,_u10_n16591 , _u10_n16590 , _u10_n16589 , _u10_n16588 , _u10_n16587 ,_u10_n16586 , _u10_n16585 , _u10_n16584 , _u10_n16583 , _u10_n16582 ,_u10_n16581 , _u10_n16580 , _u10_n16579 , _u10_n16578 , _u10_n16577 ,_u10_n16576 , _u10_n16575 , _u10_n16574 , _u10_n16573 , _u10_n16572 ,_u10_n16571 , _u10_n16570 , _u10_n16569 , _u10_n16568 , _u10_n16567 ,_u10_n16566 , _u10_n16565 , _u10_n16564 , _u10_n16563 , _u10_n16562 ,_u10_n16561 , _u10_n16560 , _u10_n16559 , _u10_n16558 , _u10_n16557 ,_u10_n16556 , _u10_n16555 , _u10_n16554 , _u10_n16553 , _u10_n16552 ,_u10_n16551 , _u10_n16550 , _u10_n16549 , _u10_n16548 , _u10_n16547 ,_u10_n16546 , _u10_n16545 , _u10_n16544 , _u10_n16543 , _u10_n16542 ,_u10_n16541 , _u10_n16540 , _u10_n16539 , _u10_n16538 , _u10_n16537 ,_u10_n16536 , _u10_n16535 , _u10_n16534 , _u10_n16533 , _u10_n16532 ,_u10_n16531 , _u10_n16530 , _u10_n16529 , _u10_n16528 , _u10_n16527 ,_u10_n16526 , _u10_n16525 , _u10_n16524 , _u10_n16523 , _u10_n16522 ,_u10_n16521 , _u10_n16520 , _u10_n16519 , _u10_n16518 , _u10_n16517 ,_u10_n16516 , _u10_n16515 , _u10_n16514 , _u10_n16513 , _u10_n16512 ,_u10_n16511 , _u10_n16510 , _u10_n16509 , _u10_n16508 , _u10_n16507 ,_u10_n16506 , _u10_n16505 , _u10_n16504 , _u10_n16503 , _u10_n16502 ,_u10_n16501 , _u10_n16500 , _u10_n16499 , _u10_n16498 , _u10_n16497 ,_u10_n16496 , _u10_n16495 , _u10_n16494 , _u10_n16493 , _u10_n16492 ,_u10_n16491 , _u10_n16490 , _u10_n16489 , _u10_n16488 , _u10_n16487 ,_u10_n16486 , _u10_n16485 , _u10_n16484 , _u10_n16483 , _u10_n16482 ,_u10_n16481 , _u10_n16480 , _u10_n16479 , _u10_n16478 , _u10_n16477 ,_u10_n16476 , _u10_n16475 , _u10_n16474 , _u10_n16473 , _u10_n16472 ,_u10_n16471 , _u10_n16470 , _u10_n16469 , _u10_n16468 , _u10_n16467 ,_u10_n16466 , _u10_n16465 , _u10_n16464 , _u10_n16463 , _u10_n16462 ,_u10_n16461 , _u10_n16460 , _u10_n16459 , _u10_n16458 , _u10_n16457 ,_u10_n16456 , _u10_n16455 , _u10_n16454 , _u10_n16453 , _u10_n16452 ,_u10_n16451 , _u10_n16450 , _u10_n16449 , _u10_n16448 , _u10_n16447 ,_u10_n16446 , _u10_n16445 , _u10_n16444 , _u10_n16443 , _u10_n16442 ,_u10_n16441 , _u10_n16440 , _u10_n16439 , _u10_n16438 , _u10_n16437 ,_u10_n16436 , _u10_n16435 , _u10_n16434 , _u10_n16433 , _u10_n16432 ,_u10_n16431 , _u10_n16430 , _u10_n16429 , _u10_n16428 , _u10_n16427 ,_u10_n16426 , _u10_n16425 , _u10_n16424 , _u10_n16423 , _u10_n16422 ,_u10_n16421 , _u10_n16420 , _u10_n16419 , _u10_n16418 , _u10_n16417 ,_u10_n16416 , _u10_n16415 , _u10_n16414 , _u10_n16413 , _u10_n16412 ,_u10_n16411 , _u10_n16410 , _u10_n16409 , _u10_n16408 , _u10_n16407 ,_u10_n16406 , _u10_n16405 , _u10_n16404 , _u10_n16403 , _u10_n16402 ,_u10_n16401 , _u10_n16400 , _u10_n16399 , _u10_n16398 , _u10_n16397 ,_u10_n16396 , _u10_n16395 , _u10_n16394 , _u10_n16393 , _u10_n16392 ,_u10_n16391 , _u10_n16390 , _u10_n16389 , _u10_n16388 , _u10_n16387 ,_u10_n16386 , _u10_n16385 , _u10_n16384 , _u10_n16383 , _u10_n16382 ,_u10_n16381 , _u10_n16380 , _u10_n16379 , _u10_n16378 , _u10_n16377 ,_u10_n16376 , _u10_n16375 , _u10_n16374 , _u10_n16373 , _u10_n16372 ,_u10_n16371 , _u10_n16370 , _u10_n16369 , _u10_n16368 , _u10_n16367 ,_u10_n16366 , _u10_n16365 , _u10_n16364 , _u10_n16363 , _u10_n16362 ,_u10_n16361 , _u10_n16360 , _u10_n16359 , _u10_n16358 , _u10_n16357 ,_u10_n16356 , _u10_n16355 , _u10_n16354 , _u10_n16353 , _u10_n16352 ,_u10_n16351 , _u10_n16350 , _u10_n16349 , _u10_n16348 , _u10_n16347 ,_u10_n16346 , _u10_n16345 , _u10_n16344 , _u10_n16343 , _u10_n16342 ,_u10_n16341 , _u10_n16340 , _u10_n16339 , _u10_n16338 , _u10_n16337 ,_u10_n16336 , _u10_n16335 , _u10_n16334 , _u10_n16333 , _u10_n16332 ,_u10_n16331 , _u10_n16330 , _u10_n16329 , _u10_n16328 , _u10_n16327 ,_u10_n16326 , _u10_n16325 , _u10_n16324 , _u10_n16323 , _u10_n16322 ,_u10_n16321 , _u10_n16320 , _u10_n16319 , _u10_n16318 , _u10_n16317 ,_u10_n16316 , _u10_n16315 , _u10_n16314 , _u10_n16313 , _u10_n16312 ,_u10_n16311 , _u10_n16310 , _u10_n16309 , _u10_n16308 , _u10_n16307 ,_u10_n16306 , _u10_n16305 , _u10_n16304 , _u10_n16303 , _u10_n16302 ,_u10_n16301 , _u10_n16300 , _u10_n16299 , _u10_n16298 , _u10_n16297 ,_u10_n16296 , _u10_n16295 , _u10_n16294 , _u10_n16293 , _u10_n16292 ,_u10_n16291 , _u10_n16290 , _u10_n16289 , _u10_n16288 , _u10_n16287 ,_u10_n16286 , _u10_n16285 , _u10_n16284 , _u10_n16283 , _u10_n16282 ,_u10_n16281 , _u10_n16280 , _u10_n16279 , _u10_n16278 , _u10_n16277 ,_u10_n16276 , _u10_n16275 , _u10_n16274 , _u10_n16273 , _u10_n16272 ,_u10_n16271 , _u10_n16270 , _u10_n16269 , _u10_n16268 , _u10_n16267 ,_u10_n16266 , _u10_n16265 , _u10_n16264 , _u10_n16263 , _u10_n16262 ,_u10_n16261 , _u10_n16260 , _u10_n16259 , _u10_n16258 , _u10_n16257 ,_u10_n16256 , _u10_n16255 , _u10_n16254 , _u10_n16253 , _u10_n16252 ,_u10_n16251 , _u10_n16250 , _u10_n16249 , _u10_n16248 , _u10_n16247 ,_u10_n16246 , _u10_n16245 , _u10_n16244 , _u10_n16243 , _u10_n16242 ,_u10_n16241 , _u10_n16240 , _u10_n16239 , _u10_n16238 , _u10_n16237 ,_u10_n16236 , _u10_n16235 , _u10_n16234 , _u10_n16233 , _u10_n16232 ,_u10_n16231 , _u10_n16230 , _u10_n16229 , _u10_n16228 , _u10_n16227 ,_u10_n16226 , _u10_n16225 , _u10_n16224 , _u10_n16223 , _u10_n16222 ,_u10_n16221 , _u10_n16220 , _u10_n16219 , _u10_n16218 , _u10_n16217 ,_u10_n16216 , _u10_n16215 , _u10_n16214 , _u10_n16213 , _u10_n16212 ,_u10_n16211 , _u10_n16210 , _u10_n16209 , _u10_n16208 , _u10_n16207 ,_u10_n16206 , _u10_n16205 , _u10_n16204 , _u10_n16203 , _u10_n16202 ,_u10_n16201 , _u10_n16200 , _u10_n16199 , _u10_n16198 , _u10_n16197 ,_u10_n16196 , _u10_n16195 , _u10_n16194 , _u10_n16193 , _u10_n16192 ,_u10_n16191 , _u10_n16190 , _u10_n16189 , _u10_n16188 , _u10_n16187 ,_u10_n16186 , _u10_n16185 , _u10_n16184 , _u10_n16183 , _u10_n16182 ,_u10_n16181 , _u10_n16180 , _u10_n16179 , _u10_n16178 , _u10_n16177 ,_u10_n16176 , _u10_n16175 , _u10_n16174 , _u10_n16173 , _u10_n16172 ,_u10_n16171 , _u10_n16170 , _u10_n16169 , _u10_n16168 , _u10_n16167 ,_u10_n16166 , _u10_n16165 , _u10_n16164 , _u10_n16163 , _u10_n16162 ,_u10_n16161 , _u10_n16160 , _u10_n16159 , _u10_n16158 , _u10_n16157 ,_u10_n16156 , _u10_n16155 , _u10_n16154 , _u10_n16153 , _u10_n16152 ,_u10_n16151 , _u10_n16150 , _u10_n16149 , _u10_n16148 , _u10_n16147 ,_u10_n16146 , _u10_n16145 , _u10_n16144 , _u10_n16143 , _u10_n16142 ,_u10_n16141 , _u10_n16140 , _u10_n16139 , _u10_n16138 , _u10_n16137 ,_u10_n16136 , _u10_n16135 , _u10_n16134 , _u10_n16133 , _u10_n16132 ,_u10_n16131 , _u10_n16130 , _u10_n16129 , _u10_n16128 , _u10_n16127 ,_u10_n16126 , _u10_n16125 , _u10_n16124 , _u10_n16123 , _u10_n16122 ,_u10_n16121 , _u10_n16120 , _u10_n16119 , _u10_n16118 , _u10_n16117 ,_u10_n16116 , _u10_n16115 , _u10_n16114 , _u10_n16113 , _u10_n16112 ,_u10_n16111 , _u10_n16110 , _u10_n16109 , _u10_n16108 , _u10_n16107 ,_u10_n16106 , _u10_n16105 , _u10_n16104 , _u10_n16103 , _u10_n16102 ,_u10_n16101 , _u10_n16100 , _u10_n16099 , _u10_n16098 , _u10_n16097 ,_u10_n16096 , _u10_n16095 , _u10_n16094 , _u10_n16093 , _u10_n16092 ,_u10_n16091 , _u10_n16090 , _u10_n16089 , _u10_n16088 , _u10_n16087 ,_u10_n16086 , _u10_n16085 , _u10_n16084 , _u10_n16083 , _u10_n16082 ,_u10_n16081 , _u10_n16080 , _u10_n16079 , _u10_n16078 , _u10_n16077 ,_u10_n16076 , _u10_n16075 , _u10_n16074 , _u10_n16073 , _u10_n16072 ,_u10_n16071 , _u10_n16070 , _u10_n16069 , _u10_n16068 , _u10_n16067 ,_u10_n16066 , _u10_n16065 , _u10_n16064 , _u10_n16063 , _u10_n16062 ,_u10_n16061 , _u10_n16060 , _u10_n16059 , _u10_n16058 , _u10_n16057 ,_u10_n16056 , _u10_n16055 , _u10_n16054 , _u10_n16053 , _u10_n16052 ,_u10_n16051 , _u10_n16050 , _u10_n16049 , _u10_n16048 , _u10_n16047 ,_u10_n16046 , _u10_n16045 , _u10_n16044 , _u10_n16043 , _u10_n16042 ,_u10_n16041 , _u10_n16040 , _u10_n16039 , _u10_n16038 , _u10_n16037 ,_u10_n16036 , _u10_n16035 , _u10_n16034 , _u10_n16033 , _u10_n16032 ,_u10_n16031 , _u10_n16030 , _u10_n16029 , _u10_n16028 , _u10_n16027 ,_u10_n16026 , _u10_n16025 , _u10_n16024 , _u10_n16023 , _u10_n16022 ,_u10_n16021 , _u10_n16020 , _u10_n16019 , _u10_n16018 , _u10_n16017 ,_u10_n16016 , _u10_n16015 , _u10_n16014 , _u10_n16013 , _u10_n16012 ,_u10_n16011 , _u10_n16010 , _u10_n16009 , _u10_n16008 , _u10_n16007 ,_u10_n16006 , _u10_n16005 , _u10_n16004 , _u10_n16003 , _u10_n16002 ,_u10_n16001 , _u10_n16000 , _u10_n15999 , _u10_n15998 , _u10_n15997 ,_u10_n15996 , _u10_n15995 , _u10_n15994 , _u10_n15993 , _u10_n15992 ,_u10_n15991 , _u10_n15990 , _u10_n15989 , _u10_n15988 , _u10_n15987 ,_u10_n15986 , _u10_n15985 , _u10_n15984 , _u10_n15983 , _u10_n15982 ,_u10_n15981 , _u10_n15980 , _u10_n15979 , _u10_n15978 , _u10_n15977 ,_u10_n15976 , _u10_n15975 , _u10_n15974 , _u10_n15973 , _u10_n15972 ,_u10_n15971 , _u10_n15970 , _u10_n15969 , _u10_n15968 , _u10_n15967 ,_u10_n15966 , _u10_n15965 , _u10_n15964 , _u10_n15963 , _u10_n15962 ,_u10_n15961 , _u10_n15960 , _u10_n15959 , _u10_n15958 , _u10_n15957 ,_u10_n15956 , _u10_n15955 , _u10_n15954 , _u10_n15953 , _u10_n15952 ,_u10_n15951 , _u10_n15950 , _u10_n15949 , _u10_n15948 , _u10_n15947 ,_u10_n15946 , _u10_n15945 , _u10_n15944 , _u10_n15943 , _u10_n15942 ,_u10_n15941 , _u10_n15940 , _u10_n15939 , _u10_n15938 , _u10_n15937 ,_u10_n15936 , _u10_n15935 , _u10_n15934 , _u10_n15933 , _u10_n15932 ,_u10_n15931 , _u10_n15930 , _u10_n15929 , _u10_n15928 , _u10_n15927 ,_u10_n15926 , _u10_n15925 , _u10_n15924 , _u10_n15923 , _u10_n15922 ,_u10_n15921 , _u10_n15920 , _u10_n15919 , _u10_n15918 , _u10_n15917 ,_u10_n15916 , _u10_n15915 , _u10_n15914 , _u10_n15913 , _u10_n15912 ,_u10_n15911 , _u10_n15910 , _u10_n15909 , _u10_n15908 , _u10_n15907 ,_u10_n15906 , _u10_n15905 , _u10_n15904 , _u10_n15903 , _u10_n15902 ,_u10_n15901 , _u10_n15900 , _u10_n15899 , _u10_n15898 , _u10_n15897 ,_u10_n15896 , _u10_n15895 , _u10_n15894 , _u10_n15893 , _u10_n15892 ,_u10_n15891 , _u10_n15890 , _u10_n15889 , _u10_n15888 , _u10_n15887 ,_u10_n15886 , _u10_n15885 , _u10_n15884 , _u10_n15883 , _u10_n15882 ,_u10_n15881 , _u10_n15880 , _u10_n15879 , _u10_n15878 , _u10_n15877 ,_u10_n15876 , _u10_n15875 , _u10_n15874 , _u10_n15873 , _u10_n15872 ,_u10_n15871 , _u10_n15870 , _u10_n15869 , _u10_n15868 , _u10_n15867 ,_u10_n15866 , _u10_n15865 , _u10_n15864 , _u10_n15863 , _u10_n15862 ,_u10_n15861 , _u10_n15860 , _u10_n15859 , _u10_n15858 , _u10_n15857 ,_u10_n15856 , _u10_n15855 , _u10_n15854 , _u10_n15853 , _u10_n15852 ,_u10_n15851 , _u10_n15850 , _u10_n15849 , _u10_n15848 , _u10_n15847 ,_u10_n15846 , _u10_n15845 , _u10_n15844 , _u10_n15843 , _u10_n15842 ,_u10_n15841 , _u10_n15840 , _u10_n15839 , _u10_n15838 , _u10_n15837 ,_u10_n15836 , _u10_n15835 , _u10_n15834 , _u10_n15833 , _u10_n15832 ,_u10_n15831 , _u10_n15830 , _u10_n15829 , _u10_n15828 , _u10_n15827 ,_u10_n15826 , _u10_n15825 , _u10_n15824 , _u10_n15823 , _u10_n15822 ,_u10_n15821 , _u10_n15820 , _u10_n15819 , _u10_n15818 , _u10_n15817 ,_u10_n15816 , _u10_n15815 , _u10_n15814 , _u10_n15813 , _u10_n15812 ,_u10_n15811 , _u10_n15810 , _u10_n15809 , _u10_n15808 , _u10_n15807 ,_u10_n15806 , _u10_n15805 , _u10_n15804 , _u10_n15803 , _u10_n15802 ,_u10_n15801 , _u10_n15800 , _u10_n15799 , _u10_n15798 , _u10_n15797 ,_u10_n15796 , _u10_n15795 , _u10_n15794 , _u10_n15793 , _u10_n15792 ,_u10_n15791 , _u10_n15790 , _u10_n15789 , _u10_n15788 , _u10_n15787 ,_u10_n15786 , _u10_n15785 , _u10_n15784 , _u10_n15783 , _u10_n15782 ,_u10_n15781 , _u10_n15780 , _u10_n15779 , _u10_n15778 , _u10_n15777 ,_u10_n15776 , _u10_n15775 , _u10_n15774 , _u10_n15773 , _u10_n15772 ,_u10_n15771 , _u10_n15770 , _u10_n15769 , _u10_n15768 , _u10_n15767 ,_u10_n15766 , _u10_n15765 , _u10_n15764 , _u10_n15763 , _u10_n15762 ,_u10_n15761 , _u10_n15760 , _u10_n15759 , _u10_n15758 , _u10_n15757 ,_u10_n15756 , _u10_n15755 , _u10_n15754 , _u10_n15753 , _u10_n15752 ,_u10_n15751 , _u10_n15750 , _u10_n15749 , _u10_n15748 , _u10_n15747 ,_u10_n15746 , _u10_n15745 , _u10_n15744 , _u10_n15743 , _u10_n15742 ,_u10_n15741 , _u10_n15740 , _u10_n15739 , _u10_n15738 , _u10_n15737 ,_u10_n15736 , _u10_n15735 , _u10_n15734 , _u10_n15733 , _u10_n15732 ,_u10_n15731 , _u10_n15730 , _u10_n15729 , _u10_n15728 , _u10_n15727 ,_u10_n15726 , _u10_n15725 , _u10_n15724 , _u10_n15723 , _u10_n15722 ,_u10_n15721 , _u10_n15720 , _u10_n15719 , _u10_n15718 , _u10_n15717 ,_u10_n15716 , _u10_n15715 , _u10_n15714 , _u10_n15713 , _u10_n15712 ,_u10_n15711 , _u10_n15710 , _u10_n15709 , _u10_n15708 , _u10_n15707 ,_u10_n15706 , _u10_n15705 , _u10_n15704 , _u10_n15703 , _u10_n15702 ,_u10_n15701 , _u10_n15700 , _u10_n15699 , _u10_n15698 , _u10_n15697 ,_u10_n15696 , _u10_n15695 , _u10_n15694 , _u10_n15693 , _u10_n15692 ,_u10_n15691 , _u10_n15690 , _u10_n15689 , _u10_n15688 , _u10_n15687 ,_u10_n15686 , _u10_n15685 , _u10_n15684 , _u10_n15683 , _u10_n15682 ,_u10_n15681 , _u10_n15680 , _u10_n15679 , _u10_n15678 , _u10_n15677 ,_u10_n15676 , _u10_n15675 , _u10_n15674 , _u10_n15673 , _u10_n15672 ,_u10_n15671 , _u10_n15670 , _u10_n15669 , _u10_n15668 , _u10_n15667 ,_u10_n15666 , _u10_n15665 , _u10_n15664 , _u10_n15663 , _u10_n15662 ,_u10_n15661 , _u10_n15660 , _u10_n15659 , _u10_n15658 , _u10_n15657 ,_u10_n15656 , _u10_n15655 , _u10_n15654 , _u10_n15653 , _u10_n15652 ,_u10_n15651 , _u10_n15650 , _u10_n15649 , _u10_n15648 , _u10_n15647 ,_u10_n15646 , _u10_n15645 , _u10_n15644 , _u10_n15643 , _u10_n15642 ,_u10_n15641 , _u10_n15640 , _u10_n15639 , _u10_n15638 , _u10_n15637 ,_u10_n15636 , _u10_n15635 , _u10_n15634 , _u10_n15633 , _u10_n15632 ,_u10_n15631 , _u10_n15630 , _u10_n15629 , _u10_n15628 , _u10_n15627 ,_u10_n15626 , _u10_n15625 , _u10_n15624 , _u10_n15623 , _u10_n15622 ,_u10_n15621 , _u10_n15620 , _u10_n15619 , _u10_n15618 , _u10_n15617 ,_u10_n15616 , _u10_n15615 , _u10_n15614 , _u10_n15613 , _u10_n15612 ,_u10_n15611 , _u10_n15610 , _u10_n15609 , _u10_n15608 , _u10_n15607 ,_u10_n15606 , _u10_n15605 , _u10_n15604 , _u10_n15603 , _u10_n15602 ,_u10_n15601 , _u10_n15600 , _u10_n15599 , _u10_n15598 , _u10_n15597 ,_u10_n15596 , _u10_n15595 , _u10_n15594 , _u10_n15593 , _u10_n15592 ,_u10_n15591 , _u10_n15590 , _u10_n15589 , _u10_n15588 , _u10_n15587 ,_u10_n15586 , _u10_n15585 , _u10_n15584 , _u10_n15583 , _u10_n15582 ,_u10_n15581 , _u10_n15580 , _u10_n15579 , _u10_n15578 , _u10_n15577 ,_u10_n15576 , _u10_n15575 , _u10_n15574 , _u10_n15573 , _u10_n15572 ,_u10_n15571 , _u10_n15570 , _u10_n15569 , _u10_n15568 , _u10_n15567 ,_u10_n15566 , _u10_n15565 , _u10_n15564 , _u10_n15563 , _u10_n15562 ,_u10_n15561 , _u10_n15560 , _u10_n15559 , _u10_n15558 , _u10_n15557 ,_u10_n15556 , _u10_n15555 , _u10_n15554 , _u10_n15553 , _u10_n15552 ,_u10_n15551 , _u10_n15550 , _u10_n15549 , _u10_n15548 , _u10_n15547 ,_u10_n15546 , _u10_n15545 , _u10_n15544 , _u10_n15543 , _u10_n15542 ,_u10_n15541 , _u10_n15540 , _u10_n15539 , _u10_n15538 , _u10_n15537 ,_u10_n15536 , _u10_n15535 , _u10_n15534 , _u10_n15533 , _u10_n15532 ,_u10_n15531 , _u10_n15530 , _u10_n15529 , _u10_n15528 , _u10_n15527 ,_u10_n15526 , _u10_n15525 , _u10_n15524 , _u10_n15523 , _u10_n15522 ,_u10_n15521 , _u10_n15520 , _u10_n15519 , _u10_n15518 , _u10_n15517 ,_u10_n15516 , _u10_n15515 , _u10_n15514 , _u10_n15513 , _u10_n15512 ,_u10_n15511 , _u10_n15510 , _u10_n15509 , _u10_n15508 , _u10_n15507 ,_u10_n15506 , _u10_n15505 , _u10_n15504 , _u10_n15503 , _u10_n15502 ,_u10_n15501 , _u10_n15500 , _u10_n15499 , _u10_n15498 , _u10_n15497 ,_u10_n15496 , _u10_n15495 , _u10_n15494 , _u10_n15493 , _u10_n15492 ,_u10_n15491 , _u10_n15490 , _u10_n15489 , _u10_n15488 , _u10_n15487 ,_u10_n15486 , _u10_n15485 , _u10_n15484 , _u10_n15483 , _u10_n15482 ,_u10_n15481 , _u10_n15480 , _u10_n15479 , _u10_n15478 , _u10_n15477 ,_u10_n15476 , _u10_n15475 , _u10_n15474 , _u10_n15473 , _u10_n15472 ,_u10_n15471 , _u10_n15470 , _u10_n15469 , _u10_n15468 , _u10_n15467 ,_u10_n15466 , _u10_n15465 , _u10_n15464 , _u10_n15463 , _u10_n15462 ,_u10_n15461 , _u10_n15460 , _u10_n15459 , _u10_n15458 , _u10_n15457 ,_u10_n15456 , _u10_n15455 , _u10_n15454 , _u10_n15453 , _u10_n15452 ,_u10_n15451 , _u10_n15450 , _u10_n15449 , _u10_n15448 , _u10_n15447 ,_u10_n15446 , _u10_n15445 , _u10_n15444 , _u10_n15443 , _u10_n15442 ,_u10_n15441 , _u10_n15440 , _u10_n15439 , _u10_n15438 , _u10_n15437 ,_u10_n15436 , _u10_n15435 , _u10_n15434 , _u10_n15433 , _u10_n15432 ,_u10_n15431 , _u10_n15430 , _u10_n15429 , _u10_n15428 , _u10_n15427 ,_u10_n15426 , _u10_n15425 , _u10_n15424 , _u10_n15423 , _u10_n15422 ,_u10_n15421 , _u10_n15420 , _u10_n15419 , _u10_n15418 , _u10_n15417 ,_u10_n15416 , _u10_n15415 , _u10_n15414 , _u10_n15413 , _u10_n15412 ,_u10_n15411 , _u10_n15410 , _u10_n15409 , _u10_n15408 , _u10_n15407 ,_u10_n15406 , _u10_n15405 , _u10_n15404 , _u10_n15403 , _u10_n15402 ,_u10_n15401 , _u10_n15400 , _u10_n15399 , _u10_n15398 , _u10_n15397 ,_u10_n15396 , _u10_n15395 , _u10_n15394 , _u10_n15393 , _u10_n15392 ,_u10_n15391 , _u10_n15390 , _u10_n15389 , _u10_n15388 , _u10_n15387 ,_u10_n15386 , _u10_n15385 , _u10_n15384 , _u10_n15383 , _u10_n15382 ,_u10_n15381 , _u10_n15380 , _u10_n15379 , _u10_n15378 , _u10_n15377 ,_u10_n15376 , _u10_n15375 , _u10_n15374 , _u10_n15373 , _u10_n15372 ,_u10_n15371 , _u10_n15370 , _u10_n15369 , _u10_n15368 , _u10_n15367 ,_u10_n15366 , _u10_n15365 , _u10_n15364 , _u10_n15363 , _u10_n15362 ,_u10_n15361 , _u10_n15360 , _u10_n15359 , _u10_n15358 , _u10_n15357 ,_u10_n15356 , _u10_n15355 , _u10_n15354 , _u10_n15353 , _u10_n15352 ,_u10_n15351 , _u10_n15350 , _u10_n15349 , _u10_n15348 , _u10_n15347 ,_u10_n15346 , _u10_n15345 , _u10_n15344 , _u10_n15343 , _u10_n15342 ,_u10_n15341 , _u10_n15340 , _u10_n15339 , _u10_n15338 , _u10_n15337 ,_u10_n15336 , _u10_n15335 , _u10_n15334 , _u10_n15333 , _u10_n15332 ,_u10_n15331 , _u10_n15330 , _u10_n15329 , _u10_n15328 , _u10_n15327 ,_u10_n15326 , _u10_n15325 , _u10_n15324 , _u10_n15323 , _u10_n15322 ,_u10_n15321 , _u10_n15320 , _u10_n15319 , _u10_n15318 , _u10_n15317 ,_u10_n15316 , _u10_n15315 , _u10_n15314 , _u10_n15313 , _u10_n15312 ,_u10_n15311 , _u10_n15310 , _u10_n15309 , _u10_n15308 , _u10_n15307 ,_u10_n15306 , _u10_n15305 , _u10_n15304 , _u10_n15303 , _u10_n15302 ,_u10_n15301 , _u10_n15300 , _u10_n15299 , _u10_n15298 , _u10_n15297 ,_u10_n15296 , _u10_n15295 , _u10_n15294 , _u10_n15293 , _u10_n15292 ,_u10_n15291 , _u10_n15290 , _u10_n15289 , _u10_n15288 , _u10_n15287 ,_u10_n15286 , _u10_n15285 , _u10_n15284 , _u10_n15283 , _u10_n15282 ,_u10_n15281 , _u10_n15280 , _u10_n15279 , _u10_n15278 , _u10_n15277 ,_u10_n15276 , _u10_n15275 , _u10_n15274 , _u10_n15273 , _u10_n15272 ,_u10_n15271 , _u10_n15270 , _u10_n15269 , _u10_n15268 , _u10_n15267 ,_u10_n15266 , _u10_n15265 , _u10_n15264 , _u10_n15263 , _u10_n15262 ,_u10_n15261 , _u10_n15260 , _u10_n15259 , _u10_n15258 , _u10_n15257 ,_u10_n15256 , _u10_n15255 , _u10_n15254 , _u10_n15253 , _u10_n15252 ,_u10_n15251 , _u10_n15250 , _u10_n15249 , _u10_n15248 , _u10_n15247 ,_u10_n15246 , _u10_n15245 , _u10_n15244 , _u10_n15243 , _u10_n15242 ,_u10_n15241 , _u10_n15240 , _u10_n15239 , _u10_n15238 , _u10_n15237 ,_u10_n15236 , _u10_n15235 , _u10_n15234 , _u10_n15233 , _u10_n15232 ,_u10_n15231 , _u10_n15230 , _u10_n15229 , _u10_n15228 , _u10_n15227 ,_u10_n15226 , _u10_n15225 , _u10_n15224 , _u10_n15223 , _u10_n15222 ,_u10_n15221 , _u10_n15220 , _u10_n15219 , _u10_n15218 , _u10_n15217 ,_u10_n15216 , _u10_n15215 , _u10_n15214 , _u10_n15213 , _u10_n15212 ,_u10_n15211 , _u10_n15210 , _u10_n15209 , _u10_n15208 , _u10_n15207 ,_u10_n15206 , _u10_n15205 , _u10_n15204 , _u10_n15203 , _u10_n15202 ,_u10_n15201 , _u10_n15200 , _u10_n15199 , _u10_n15198 , _u10_n15197 ,_u10_n15196 , _u10_n15195 , _u10_n15194 , _u10_n15193 , _u10_n15192 ,_u10_n15191 , _u10_n15190 , _u10_n15189 , _u10_n15188 , _u10_n15187 ,_u10_n15186 , _u10_n15185 , _u10_n15184 , _u10_n15183 , _u10_n15182 ,_u10_n15181 , _u10_n15180 , _u10_n15179 , _u10_n15178 , _u10_n15177 ,_u10_n15176 , _u10_n15175 , _u10_n15174 , _u10_n15173 , _u10_n15172 ,_u10_n15171 , _u10_n15170 , _u10_n15169 , _u10_n15168 , _u10_n15167 ,_u10_n15166 , _u10_n15165 , _u10_n15164 , _u10_n15163 , _u10_n15162 ,_u10_n15161 , _u10_n15160 , _u10_n15159 , _u10_n15158 , _u10_n15157 ,_u10_n15156 , _u10_n15155 , _u10_n15154 , _u10_n15153 , _u10_n15152 ,_u10_n15151 , _u10_n15150 , _u10_n15149 , _u10_n15148 , _u10_n15147 ,_u10_n15146 , _u10_n15145 , _u10_n15144 , _u10_n15143 , _u10_n15142 ,_u10_n15141 , _u10_n15140 , _u10_n15139 , _u10_n15138 , _u10_n15137 ,_u10_n15136 , _u10_n15135 , _u10_n15134 , _u10_n15133 , _u10_n15132 ,_u10_n15131 , _u10_n15130 , _u10_n15129 , _u10_n15128 , _u10_n15127 ,_u10_n15126 , _u10_n15125 , _u10_n15124 , _u10_n15123 , _u10_n15122 ,_u10_n15121 , _u10_n15120 , _u10_n15119 , _u10_n15118 , _u10_n15117 ,_u10_n15116 , _u10_n15115 , _u10_n15114 , _u10_n15113 , _u10_n15112 ,_u10_n15111 , _u10_n15110 , _u10_n15109 , _u10_n15108 , _u10_n15107 ,_u10_n15106 , _u10_n15105 , _u10_n15104 , _u10_n15103 , _u10_n15102 ,_u10_n15101 , _u10_n15100 , _u10_n15099 , _u10_n15098 , _u10_n15097 ,_u10_n15096 , _u10_n15095 , _u10_n15094 , _u10_n15093 , _u10_n15092 ,_u10_n15091 , _u10_n15090 , _u10_n15089 , _u10_n15088 , _u10_n15087 ,_u10_n15086 , _u10_n15085 , _u10_n15084 , _u10_n15083 , _u10_n15082 ,_u10_n15081 , _u10_n15080 , _u10_n15079 , _u10_n15078 , _u10_n15077 ,_u10_n15076 , _u10_n15075 , _u10_n15074 , _u10_n15073 , _u10_n15072 ,_u10_n15071 , _u10_n15070 , _u10_n15069 , _u10_n15068 , _u10_n15067 ,_u10_n15066 , _u10_n15065 , _u10_n15064 , _u10_n15063 , _u10_n15062 ,_u10_n15061 , _u10_n15060 , _u10_n15059 , _u10_n15058 , _u10_n15057 ,_u10_n15056 , _u10_n15055 , _u10_n15054 , _u10_n15053 , _u10_n15052 ,_u10_n15051 , _u10_n15050 , _u10_n15049 , _u10_n15048 , _u10_n15047 ,_u10_n15046 , _u10_n15045 , _u10_n15044 , _u10_n15043 , _u10_n15042 ,_u10_n15041 , _u10_n15040 , _u10_n15039 , _u10_n15038 , _u10_n15037 ,_u10_n15036 , _u10_n15035 , _u10_n15034 , _u10_n15033 , _u10_n15032 ,_u10_n15031 , _u10_n15030 , _u10_n15029 , _u10_n15028 , _u10_n15027 ,_u10_n15026 , _u10_n15025 , _u10_n15024 , _u10_n15023 , _u10_n15022 ,_u10_n15021 , _u10_n15020 , _u10_n15019 , _u10_n15018 , _u10_n15017 ,_u10_n15016 , _u10_n15015 , _u10_n15014 , _u10_n15013 , _u10_n15012 ,_u10_n15011 , _u10_n15010 , _u10_n15009 , _u10_n15008 , _u10_n15007 ,_u10_n15006 , _u10_n15005 , _u10_n15004 , _u10_n15003 , _u10_n15002 ,_u10_n15001 , _u10_n15000 , _u10_n14999 , _u10_n14998 , _u10_n14997 ,_u10_n14996 , _u10_n14995 , _u10_n14994 , _u10_n14993 , _u10_n14992 ,_u10_n14991 , _u10_n14990 , _u10_n14989 , _u10_n14988 , _u10_n14987 ,_u10_n14986 , _u10_n14985 , _u10_n14984 , _u10_n14983 , _u10_n14982 ,_u10_n14981 , _u10_n14980 , _u10_n14979 , _u10_n14978 , _u10_n14977 ,_u10_n14976 , _u10_n14975 , _u10_n14974 , _u10_n14973 , _u10_n14972 ,_u10_n14971 , _u10_n14970 , _u10_n14969 , _u10_n14968 , _u10_n14967 ,_u10_n14966 , _u10_n14965 , _u10_n14964 , _u10_n14963 , _u10_n14962 ,_u10_n14961 , _u10_n14960 , _u10_n14959 , _u10_n14958 , _u10_n14957 ,_u10_n14956 , _u10_n14955 , _u10_n14954 , _u10_n14953 , _u10_n14952 ,_u10_n14951 , _u10_n14950 , _u10_n14949 , _u10_n14948 , _u10_n14947 ,_u10_n14946 , _u10_n14945 , _u10_n14944 , _u10_n14943 , _u10_n14942 ,_u10_n14941 , _u10_n14940 , _u10_n14939 , _u10_n14938 , _u10_n14937 ,_u10_n14936 , _u10_n14935 , _u10_n14934 , _u10_n14933 , _u10_n14932 ,_u10_n14931 , _u10_n14930 , _u10_n14929 , _u10_n14928 , _u10_n14927 ,_u10_n14926 , _u10_n14925 , _u10_n14924 , _u10_n14923 , _u10_n14922 ,_u10_n14921 , _u10_n14920 , _u10_n14919 , _u10_n14918 , _u10_n14917 ,_u10_n14916 , _u10_n14915 , _u10_n14914 , _u10_n14913 , _u10_n14912 ,_u10_n14911 , _u10_n14910 , _u10_n14909 , _u10_n14908 , _u10_n14907 ,_u10_n14906 , _u10_n14905 , _u10_n14904 , _u10_n14903 , _u10_n14902 ,_u10_n14901 , _u10_n14900 , _u10_n14899 , _u10_n14898 , _u10_n14897 ,_u10_n14896 , _u10_n14895 , _u10_n14894 , _u10_n14893 , _u10_n14892 ,_u10_n14891 , _u10_n14890 , _u10_n14889 , _u10_n14888 , _u10_n14887 ,_u10_n14886 , _u10_n14885 , _u10_n14884 , _u10_n14883 , _u10_n14882 ,_u10_n14881 , _u10_n14880 , _u10_n14879 , _u10_n14878 , _u10_n14877 ,_u10_n14876 , _u10_n14875 , _u10_n14874 , _u10_n14873 , _u10_n14872 ,_u10_n14871 , _u10_n14870 , _u10_n14869 , _u10_n14868 , _u10_n14867 ,_u10_n14866 , _u10_n14865 , _u10_n14864 , _u10_n14863 , _u10_n14862 ,_u10_n14861 , _u10_n14860 , _u10_n14859 , _u10_n14858 , _u10_n14857 ,_u10_n14856 , _u10_n14855 , _u10_n14854 , _u10_n14853 , _u10_n14852 ,_u10_n14851 , _u10_n14850 , _u10_n14849 , _u10_n14848 , _u10_n14847 ,_u10_n14846 , _u10_n14845 , _u10_n14844 , _u10_n14843 , _u10_n14842 ,_u10_n14841 , _u10_n14840 , _u10_n14839 , _u10_n14838 , _u10_n14837 ,_u10_n14836 , _u10_n14835 , _u10_n14834 , _u10_n14833 , _u10_n14832 ,_u10_n14831 , _u10_n14830 , _u10_n14829 , _u10_n14828 , _u10_n14827 ,_u10_n14826 , _u10_n14825 , _u10_n14824 , _u10_n14823 , _u10_n14822 ,_u10_n14821 , _u10_n14820 , _u10_n14819 , _u10_n14818 , _u10_n14817 ,_u10_n14816 , _u10_n14815 , _u10_n14814 , _u10_n14813 , _u10_n14812 ,_u10_n14811 , _u10_n14810 , _u10_n14809 , _u10_n14808 , _u10_n14807 ,_u10_n14806 , _u10_n14805 , _u10_n14804 , _u10_n14803 , _u10_n14802 ,_u10_n14801 , _u10_n14800 , _u10_n14799 , _u10_n14798 , _u10_n14797 ,_u10_n14796 , _u10_n14795 , _u10_n14794 , _u10_n14793 , _u10_n14792 ,_u10_n14791 , _u10_n14790 , _u10_n14789 , _u10_n14788 , _u10_n14787 ,_u10_n14786 , _u10_n14785 , _u10_n14784 , _u10_n14783 , _u10_n14782 ,_u10_n14781 , _u10_n14780 , _u10_n14779 , _u10_n14778 , _u10_n14777 ,_u10_n14776 , _u10_n14775 , _u10_n14774 , _u10_n14773 , _u10_n14772 ,_u10_n14771 , _u10_n14770 , _u10_n14769 , _u10_n14768 , _u10_n14767 ,_u10_n14766 , _u10_n14765 , _u10_n14764 , _u10_n14763 , _u10_n14762 ,_u10_n14761 , _u10_n14760 , _u10_n14759 , _u10_n14758 , _u10_n14757 ,_u10_n14756 , _u10_n14755 , _u10_n14754 , _u10_n14753 , _u10_n14752 ,_u10_n14751 , _u10_n14750 , _u10_n14749 , _u10_n14748 , _u10_n14747 ,_u10_n14746 , _u10_n14745 , _u10_n14744 , _u10_n14743 , _u10_n14742 ,_u10_n14741 , _u10_n14740 , _u10_n14739 , _u10_n14738 , _u10_n14737 ,_u10_n14736 , _u10_n14735 , _u10_n14734 , _u10_n14733 , _u10_n14732 ,_u10_n14731 , _u10_n14730 , _u10_n14729 , _u10_n14728 , _u10_n14727 ,_u10_n14726 , _u10_n14725 , _u10_n14724 , _u10_n14723 , _u10_n14722 ,_u10_n14721 , _u10_n14720 , _u10_n14719 , _u10_n14718 , _u10_n14717 ,_u10_n14716 , _u10_n14715 , _u10_n14714 , _u10_n14713 , _u10_n14712 ,_u10_n14711 , _u10_n14710 , _u10_n14709 , _u10_n14708 , _u10_n14707 ,_u10_n14706 , _u10_n14705 , _u10_n14704 , _u10_n14703 , _u10_n14702 ,_u10_n14701 , _u10_n14700 , _u10_n14699 , _u10_n14698 , _u10_n14697 ,_u10_n14696 , _u10_n14695 , _u10_n14694 , _u10_n14693 , _u10_n14692 ,_u10_n14691 , _u10_n14690 , _u10_n14689 , _u10_n14688 , _u10_n14687 ,_u10_n14686 , _u10_n14685 , _u10_n14684 , _u10_n14683 , _u10_n14682 ,_u10_n14681 , _u10_n14680 , _u10_n14679 , _u10_n14678 , _u10_n14677 ,_u10_n14676 , _u10_n14675 , _u10_n14674 , _u10_n14673 , _u10_n14672 ,_u10_n14671 , _u10_n14670 , _u10_n14669 , _u10_n14668 , _u10_n14667 ,_u10_n14666 , _u10_n14665 , _u10_n14664 , _u10_n14663 , _u10_n14662 ,_u10_n14661 , _u10_n14660 , _u10_n14659 , _u10_n14658 , _u10_n14657 ,_u10_n14656 , _u10_n14655 , _u10_n14654 , _u10_n14653 , _u10_n14652 ,_u10_n14651 , _u10_n14650 , _u10_n14649 , _u10_n14648 , _u10_n14647 ,_u10_n14646 , _u10_n14645 , _u10_n14644 , _u10_n14643 , _u10_n14642 ,_u10_n14641 , _u10_n14640 , _u10_n14639 , _u10_n14638 , _u10_n14637 ,_u10_n14636 , _u10_n14635 , _u10_n14634 , _u10_n14633 , _u10_n14632 ,_u10_n14631 , _u10_n14630 , _u10_n14629 , _u10_n14628 , _u10_n14627 ,_u10_n14626 , _u10_n14625 , _u10_n14624 , _u10_n14623 , _u10_n14622 ,_u10_n14621 , _u10_n14620 , _u10_n14619 , _u10_n14618 , _u10_n14617 ,_u10_n14616 , _u10_n14615 , _u10_n14614 , _u10_n14613 , _u10_n14612 ,_u10_n14611 , _u10_n14610 , _u10_n14609 , _u10_n14608 , _u10_n14607 ,_u10_n14606 , _u10_n14605 , _u10_n14604 , _u10_n14603 , _u10_n14602 ,_u10_n14601 , _u10_n14600 , _u10_n14599 , _u10_n14598 , _u10_n14597 ,_u10_n14596 , _u10_n14595 , _u10_n14594 , _u10_n14593 , _u10_n14592 ,_u10_n14591 , _u10_n14590 , _u10_n14589 , _u10_n14588 , _u10_n14587 ,_u10_n14586 , _u10_n14585 , _u10_n14584 , _u10_n14583 , _u10_n14582 ,_u10_n14581 , _u10_n14580 , _u10_n14579 , _u10_n14578 , _u10_n14577 ,_u10_n14576 , _u10_n14575 , _u10_n14574 , _u10_n14573 , _u10_n14572 ,_u10_n14571 , _u10_n14570 , _u10_n14569 , _u10_n14568 , _u10_n14567 ,_u10_n14566 , _u10_n14565 , _u10_n14564 , _u10_n14563 , _u10_n14562 ,_u10_n14561 , _u10_n14560 , _u10_n14559 , _u10_n14558 , _u10_n14557 ,_u10_n14556 , _u10_n14555 , _u10_n14554 , _u10_n14553 , _u10_n14552 ,_u10_n14551 , _u10_n14550 , _u10_n14549 , _u10_n14548 , _u10_n14547 ,_u10_n14546 , _u10_n14545 , _u10_n14544 , _u10_n14543 , _u10_n14542 ,_u10_n14541 , _u10_n14540 , _u10_n14539 , _u10_n14538 , _u10_n14537 ,_u10_n14536 , _u10_n14535 , _u10_n14534 , _u10_n14533 , _u10_n14532 ,_u10_n14531 , _u10_n14530 , _u10_n14529 , _u10_n14528 , _u10_n14527 ,_u10_n14526 , _u10_n14525 , _u10_n14524 , _u10_n14523 , _u10_n14522 ,_u10_n14521 , _u10_n14520 , _u10_n14519 , _u10_n14518 , _u10_n14517 ,_u10_n14516 , _u10_n14515 , _u10_n14514 , _u10_n14513 , _u10_n14512 ,_u10_n14511 , _u10_n14510 , _u10_n14509 , _u10_n14508 , _u10_n14507 ,_u10_n14506 , _u10_n14505 , _u10_n14504 , _u10_n14503 , _u10_n14502 ,_u10_n14501 , _u10_n14500 , _u10_n14499 , _u10_n14498 , _u10_n14497 ,_u10_n14496 , _u10_n14495 , _u10_n14494 , _u10_n14493 , _u10_n14492 ,_u10_n14491 , _u10_n14490 , _u10_n14489 , _u10_n14488 , _u10_n14487 ,_u10_n14486 , _u10_n14485 , _u10_n14484 , _u10_n14483 , _u10_n14482 ,_u10_n14481 , _u10_n14480 , _u10_n14479 , _u10_n14478 , _u10_n14477 ,_u10_n14476 , _u10_n14475 , _u10_n14474 , _u10_n14473 , _u10_n14472 ,_u10_n14471 , _u10_n14470 , _u10_n14469 , _u10_n14468 , _u10_n14467 ,_u10_n14466 , _u10_n14465 , _u10_n14464 , _u10_n14463 , _u10_n14462 ,_u10_n14461 , _u10_n14460 , _u10_n14459 , _u10_n14458 , _u10_n14457 ,_u10_n14456 , _u10_n14455 , _u10_n14454 , _u10_n14453 , _u10_n14452 ,_u10_n14451 , _u10_n14450 , _u10_n14449 , _u10_n14448 , _u10_n14447 ,_u10_n14446 , _u10_n14445 , _u10_n14444 , _u10_n14443 , _u10_n14442 ,_u10_n14441 , _u10_n14440 , _u10_n14439 , _u10_n14438 , _u10_n14437 ,_u10_n14436 , _u10_n14435 , _u10_n14434 , _u10_n14433 , _u10_n14432 ,_u10_n14431 , _u10_n14430 , _u10_n14429 , _u10_n14428 , _u10_n14427 ,_u10_n14426 , _u10_n14425 , _u10_n14424 , _u10_n14423 , _u10_n14422 ,_u10_n14421 , _u10_n14420 , _u10_n14419 , _u10_n14418 , _u10_n14417 ,_u10_n14416 , _u10_n14415 , _u10_n14414 , _u10_n14413 , _u10_n14412 ,_u10_n14411 , _u10_n14410 , _u10_n14409 , _u10_n14408 , _u10_n14407 ,_u10_n14406 , _u10_n14405 , _u10_n14404 , _u10_n14403 , _u10_n14402 ,_u10_n14401 , _u10_n14400 , _u10_n14399 , _u10_n14398 , _u10_n14397 ,_u10_n14396 , _u10_n14395 , _u10_n14394 , _u10_n14393 , _u10_n14392 ,_u10_n14391 , _u10_n14390 , _u10_n14389 , _u10_n14388 , _u10_n14387 ,_u10_n14386 , _u10_n14385 , _u10_n14384 , _u10_n14383 , _u10_n14382 ,_u10_n14381 , _u10_n14380 , _u10_n14379 , _u10_n14378 , _u10_n14377 ,_u10_n14376 , _u10_n14375 , _u10_n14374 , _u10_n14373 , _u10_n14372 ,_u10_n14371 , _u10_n14370 , _u10_n14369 , _u10_n14368 , _u10_n14367 ,_u10_n14366 , _u10_n14365 , _u10_n14364 , _u10_n14363 , _u10_n14362 ,_u10_n14361 , _u10_n14360 , _u10_n14359 , _u10_n14358 , _u10_n14357 ,_u10_n14356 , _u10_n14355 , _u10_n14354 , _u10_n14353 , _u10_n14352 ,_u10_n14351 , _u10_n14350 , _u10_n14349 , _u10_n14348 , _u10_n14347 ,_u10_n14346 , _u10_n14345 , _u10_n14344 , _u10_n14343 , _u10_n14342 ,_u10_n14341 , _u10_n14340 , _u10_n14339 , _u10_n14338 , _u10_n14337 ,_u10_n14336 , _u10_n14335 , _u10_n14334 , _u10_n14333 , _u10_n14332 ,_u10_n14331 , _u10_n14330 , _u10_n14329 , _u10_n14328 , _u10_n14327 ,_u10_n14326 , _u10_n14325 , _u10_n14324 , _u10_n14323 , _u10_n14322 ,_u10_n14321 , _u10_n14320 , _u10_n14319 , _u10_n14318 , _u10_n14317 ,_u10_n14316 , _u10_n14315 , _u10_n14314 , _u10_n14313 , _u10_n14312 ,_u10_n14311 , _u10_n14310 , _u10_n14309 , _u10_n14308 , _u10_n14307 ,_u10_n14306 , _u10_n14305 , _u10_n14304 , _u10_n14303 , _u10_n14302 ,_u10_n14301 , _u10_n14300 , _u10_n14299 , _u10_n14298 , _u10_n14297 ,_u10_n14296 , _u10_n14295 , _u10_n14294 , _u10_n14293 , _u10_n14292 ,_u10_n14291 , _u10_n14290 , _u10_n14289 , _u10_n14288 , _u10_n14287 ,_u10_n14286 , _u10_n14285 , _u10_n14284 , _u10_n14283 , _u10_n14282 ,_u10_n14281 , _u10_n14280 , _u10_n14279 , _u10_n14278 , _u10_n14277 ,_u10_n14276 , _u10_n14275 , _u10_n14274 , _u10_n14273 , _u10_n14272 ,_u10_n14271 , _u10_n14270 , _u10_n14269 , _u10_n14268 , _u10_n14267 ,_u10_n14266 , _u10_n14265 , _u10_n14264 , _u10_n14263 , _u10_n14262 ,_u10_n14261 , _u10_n14260 , _u10_n14259 , _u10_n14258 , _u10_n14257 ,_u10_n14256 , _u10_n14255 , _u10_n14254 , _u10_n14253 , _u10_n14252 ,_u10_n14251 , _u10_n14250 , _u10_n14249 , _u10_n14248 , _u10_n14247 ,_u10_n14246 , _u10_n14245 , _u10_n14244 , _u10_n14243 , _u10_n14242 ,_u10_n14241 , _u10_n14240 , _u10_n14239 , _u10_n14238 , _u10_n14237 ,_u10_n14236 , _u10_n14235 , _u10_n14234 , _u10_n14233 , _u10_n14232 ,_u10_n14231 , _u10_n14230 , _u10_n14229 , _u10_n14228 , _u10_n14227 ,_u10_n14226 , _u10_n14225 , _u10_n14224 , _u10_n14223 , _u10_n14222 ,_u10_n14221 , _u10_n14220 , _u10_n14219 , _u10_n14218 , _u10_n14217 ,_u10_n14216 , _u10_n14215 , _u10_n14214 , _u10_n14213 , _u10_n14212 ,_u10_n14211 , _u10_n14210 , _u10_n14209 , _u10_n14208 , _u10_n14207 ,_u10_n14206 , _u10_n14205 , _u10_n14204 , _u10_n14203 , _u10_n14202 ,_u10_n14201 , _u10_n14200 , _u10_n14199 , _u10_n14198 , _u10_n14197 ,_u10_n14196 , _u10_n14195 , _u10_n14194 , _u10_n14193 , _u10_n14192 ,_u10_n14191 , _u10_n14190 , _u10_n14189 , _u10_n14188 , _u10_n14187 ,_u10_n14186 , _u10_n14185 , _u10_n14184 , _u10_n14183 , _u10_n14182 ,_u10_n14181 , _u10_n14180 , _u10_n14179 , _u10_n14178 , _u10_n14177 ,_u10_n14176 , _u10_n14175 , _u10_n14174 , _u10_n14173 , _u10_n14172 ,_u10_n14171 , _u10_n14170 , _u10_n14169 , _u10_n14168 , _u10_n14167 ,_u10_n14166 , _u10_n14165 , _u10_n14164 , _u10_n14163 , _u10_n14162 ,_u10_n14161 , _u10_n14160 , _u10_n14159 , _u10_n14158 , _u10_n14157 ,_u10_n14156 , _u10_n14155 , _u10_n14154 , _u10_n14153 , _u10_n14152 ,_u10_n14151 , _u10_n14150 , _u10_n14149 , _u10_n14148 , _u10_n14147 ,_u10_n14146 , _u10_n14145 , _u10_n14144 , _u10_n14143 , _u10_n14142 ,_u10_n14141 , _u10_n14140 , _u10_n14139 , _u10_n14138 , _u10_n14137 ,_u10_n14136 , _u10_n14135 , _u10_n14134 , _u10_n14133 , _u10_n14132 ,_u10_n14131 , _u10_n14130 , _u10_n14129 , _u10_n14128 , _u10_n14127 ,_u10_n14126 , _u10_n14125 , _u10_n14124 , _u10_n14123 , _u10_n14122 ,_u10_n14121 , _u10_n14120 , _u10_n14119 , _u10_n14118 , _u10_n14117 ,_u10_n14116 , _u10_n14115 , _u10_n14114 , _u10_n14113 , _u10_n14112 ,_u10_n14111 , _u10_n14110 , _u10_n14109 , _u10_n14108 , _u10_n14107 ,_u10_n14106 , _u10_n14105 , _u10_n14104 , _u10_n14103 , _u10_n14102 ,_u10_n14101 , _u10_n14100 , _u10_n14099 , _u10_n14098 , _u10_n14097 ,_u10_n14096 , _u10_n14095 , _u10_n14094 , _u10_n14093 , _u10_n14092 ,_u10_n14091 , _u10_n14090 , _u10_n14089 , _u10_n14088 , _u10_n14087 ,_u10_n14086 , _u10_n14085 , _u10_n14084 , _u10_n14083 , _u10_n14082 ,_u10_n14081 , _u10_n14080 , _u10_n14079 , _u10_n14078 , _u10_n14077 ,_u10_n14076 , _u10_n14075 , _u10_n14074 , _u10_n14073 , _u10_n14072 ,_u10_n14071 , _u10_n14070 , _u10_n14069 , _u10_n14068 , _u10_n14067 ,_u10_n14066 , _u10_n14065 , _u10_n14064 , _u10_n14063 , _u10_n14062 ,_u10_n14061 , _u10_n14060 , _u10_n14059 , _u10_n14058 , _u10_n14057 ,_u10_n14056 , _u10_n14055 , _u10_n14054 , _u10_n14053 , _u10_n14052 ,_u10_n14051 , _u10_n14050 , _u10_n14049 , _u10_n14048 , _u10_n14047 ,_u10_n14046 , _u10_n14045 , _u10_n14044 , _u10_n14043 , _u10_n14042 ,_u10_n14041 , _u10_n14040 , _u10_n14039 , _u10_n14038 , _u10_n14037 ,_u10_n14036 , _u10_n14035 , _u10_n14034 , _u10_n14033 , _u10_n14032 ,_u10_n14031 , _u10_n14030 , _u10_n14029 , _u10_n14028 , _u10_n14027 ,_u10_n14026 , _u10_n14025 , _u10_n14024 , _u10_n14023 , _u10_n14022 ,_u10_n14021 , _u10_n14020 , _u10_n14019 , _u10_n14018 , _u10_n14017 ,_u10_n14016 , _u10_n14015 , _u10_n14014 , _u10_n14013 , _u10_n14012 ,_u10_n14011 , _u10_n14010 , _u10_n14009 , _u10_n14008 , _u10_n14007 ,_u10_n14006 , _u10_n14005 , _u10_n14004 , _u10_n14003 , _u10_n14002 ,_u10_n14001 , _u10_n14000 , _u10_n13999 , _u10_n13998 , _u10_n13997 ,_u10_n13996 , _u10_n13995 , _u10_n13994 , _u10_n13993 , _u10_n13992 ,_u10_n13991 , _u10_n13990 , _u10_n13989 , _u10_n13988 , _u10_n13987 ,_u10_n13986 , _u10_n13985 , _u10_n13984 , _u10_n13983 , _u10_n13982 ,_u10_n13981 , _u10_n13980 , _u10_n13979 , _u10_n13978 , _u10_n13977 ,_u10_n13976 , _u10_n13975 , _u10_n13974 , _u10_n13973 , _u10_n13972 ,_u10_n13971 , _u10_n13970 , _u10_n13969 , _u10_n13968 , _u10_n13967 ,_u10_n13966 , _u10_n13965 , _u10_n13964 , _u10_n13963 , _u10_n13962 ,_u10_n13961 , _u10_n13960 , _u10_n13959 , _u10_n13958 , _u10_n13957 ,_u10_n13956 , _u10_n13955 , _u10_n13954 , _u10_n13953 , _u10_n13952 ,_u10_n13951 , _u10_n13950 , _u10_n13949 , _u10_n13948 , _u10_n13947 ,_u10_n13946 , _u10_n13945 , _u10_n13944 , _u10_n13943 , _u10_n13942 ,_u10_n13941 , _u10_n13940 , _u10_n13939 , _u10_n13938 , _u10_n13937 ,_u10_n13936 , _u10_n13935 , _u10_n13934 , _u10_n13933 , _u10_n13932 ,_u10_n13931 , _u10_n13930 , _u10_n13929 , _u10_n13928 , _u10_n13927 ,_u10_n13926 , _u10_n13925 , _u10_n13924 , _u10_n13923 , _u10_n13922 ,_u10_n13921 , _u10_n13920 , _u10_n13919 , _u10_n13918 , _u10_n13917 ,_u10_n13916 , _u10_n13915 , _u10_n13914 , _u10_n13913 , _u10_n13912 ,_u10_n13911 , _u10_n13910 , _u10_n13909 , _u10_n13908 , _u10_n13907 ,_u10_n13906 , _u10_n13905 , _u10_n13904 , _u10_n13903 , _u10_n13902 ,_u10_n13901 , _u10_n13900 , _u10_n13899 , _u10_n13898 , _u10_n13897 ,_u10_n13896 , _u10_n13895 , _u10_n13894 , _u10_n13893 , _u10_n13892 ,_u10_n13891 , _u10_n13890 , _u10_n13889 , _u10_n13888 , _u10_n13887 ,_u10_n13886 , _u10_n13885 , _u10_n13884 , _u10_n13883 , _u10_n13882 ,_u10_n13881 , _u10_n13880 , _u10_n13879 , _u10_n13878 , _u10_n13877 ,_u10_n13876 , _u10_n13875 , _u10_n13874 , _u10_n13873 , _u10_n13872 ,_u10_n13871 , _u10_n13870 , _u10_n13869 , _u10_n13868 , _u10_n13867 ,_u10_n13866 , _u10_n13865 , _u10_n13864 , _u10_n13863 , _u10_n13862 ,_u10_n13861 , _u10_n13860 , _u10_n13859 , _u10_n13858 , _u10_n13857 ,_u10_n13856 , _u10_n13855 , _u10_n13854 , _u10_n13853 , _u10_n13852 ,_u10_n13851 , _u10_n13850 , _u10_n13849 , _u10_n13848 , _u10_n13847 ,_u10_n13846 , _u10_n13845 , _u10_n13844 , _u10_n13843 , _u10_n13842 ,_u10_n13841 , _u10_n13840 , _u10_n13839 , _u10_n13838 , _u10_n13837 ,_u10_n13836 , _u10_n13835 , _u10_n13834 , _u10_n13833 , _u10_n13832 ,_u10_n13831 , _u10_n13830 , _u10_n13829 , _u10_n13828 , _u10_n13827 ,_u10_n13826 , _u10_n13825 , _u10_n13824 , _u10_n13823 , _u10_n13822 ,_u10_n13821 , _u10_n13820 , _u10_n13819 , _u10_n13818 , _u10_n13817 ,_u10_n13816 , _u10_n13815 , _u10_n13814 , _u10_n13813 , _u10_n13812 ,_u10_n13811 , _u10_n13810 , _u10_n13809 , _u10_n13808 , _u10_n13807 ,_u10_n13806 , _u10_n13805 , _u10_n13804 , _u10_n13803 , _u10_n13802 ,_u10_n13801 , _u10_n13800 , _u10_n13799 , _u10_n13798 , _u10_n13797 ,_u10_n13796 , _u10_n13795 , _u10_n13794 , _u10_n13793 , _u10_n13792 ,_u10_n13791 , _u10_n13790 , _u10_n13789 , _u10_n13788 , _u10_n13787 ,_u10_n13786 , _u10_n13785 , _u10_n13784 , _u10_n13783 , _u10_n13782 ,_u10_n13781 , _u10_n13780 , _u10_n13779 , _u10_n13778 , _u10_n13777 ,_u10_n13776 , _u10_n13775 , _u10_n13774 , _u10_n13773 , _u10_n13772 ,_u10_n13771 , _u10_n13770 , _u10_n13769 , _u10_n13768 , _u10_n13767 ,_u10_n13766 , _u10_n13765 , _u10_n13764 , _u10_n13763 , _u10_n13762 ,_u10_n13761 , _u10_n13760 , _u10_n13759 , _u10_n13758 , _u10_n13757 ,_u10_n13756 , _u10_n13755 , _u10_n13754 , _u10_n13753 , _u10_n13752 ,_u10_n13751 , _u10_n13750 , _u10_n13749 , _u10_n13748 , _u10_n13747 ,_u10_n13746 , _u10_n13745 , _u10_n13744 , _u10_n13743 , _u10_n13742 ,_u10_n13741 , _u10_n13740 , _u10_n13739 , _u10_n13738 , _u10_n13737 ,_u10_n13736 , _u10_n13735 , _u10_n13734 , _u10_n13733 , _u10_n13732 ,_u10_n13731 , _u10_n13730 , _u10_n13729 , _u10_n13728 , _u10_n13727 ,_u10_n13726 , _u10_n13725 , _u10_n13724 , _u10_n13723 , _u10_n13722 ,_u10_n13721 , _u10_n13720 , _u10_n13719 , _u10_n13718 , _u10_n13717 ,_u10_n13716 , _u10_n13715 , _u10_n13714 , _u10_n13713 , _u10_n13712 ,_u10_n13711 , _u10_n13710 , _u10_n13709 , _u10_n13708 , _u10_n13707 ,_u10_n13706 , _u10_n13705 , _u10_n13704 , _u10_n13703 , _u10_n13702 ,_u10_n13701 , _u10_n13700 , _u10_n13699 , _u10_n13698 , _u10_n13697 ,_u10_n13696 , _u10_n13695 , _u10_n13694 , _u10_n13693 , _u10_n13692 ,_u10_n13691 , _u10_n13690 , _u10_n13689 , _u10_n13688 , _u10_n13687 ,_u10_n13686 , _u10_n13685 , _u10_n13684 , _u10_n13683 , _u10_n13682 ,_u10_n13681 , _u10_n13680 , _u10_n13679 , _u10_n13678 , _u10_n13677 ,_u10_n13676 , _u10_n13675 , _u10_n13674 , _u10_n13673 , _u10_n13672 ,_u10_n13671 , _u10_n13670 , _u10_n13669 , _u10_n13668 , _u10_n13667 ,_u10_n13666 , _u10_n13665 , _u10_n13664 , _u10_n13663 , _u10_n13662 ,_u10_n13661 , _u10_n13660 , _u10_n13659 , _u10_n13658 , _u10_n13657 ,_u10_n13656 , _u10_n13655 , _u10_n13654 , _u10_n13653 , _u10_n13652 ,_u10_n13651 , _u10_n13650 , _u10_n13649 , _u10_n13648 , _u10_n13647 ,_u10_n13646 , _u10_n13645 , _u10_n13644 , _u10_n13643 , _u10_n13642 ,_u10_n13641 , _u10_n13640 , _u10_n13639 , _u10_n13638 , _u10_n13637 ,_u10_n13636 , _u10_n13635 , _u10_n13634 , _u10_n13633 , _u10_n13632 ,_u10_n13631 , _u10_n13630 , _u10_n13629 , _u10_n13628 , _u10_n13627 ,_u10_n13626 , _u10_n13625 , _u10_n13624 , _u10_n13623 , _u10_n13622 ,_u10_n13621 , _u10_n13620 , _u10_n13619 , _u10_n13618 , _u10_n13617 ,_u10_n13616 , _u10_n13615 , _u10_n13614 , _u10_n13613 , _u10_n13612 ,_u10_n13611 , _u10_n13610 , _u10_n13609 , _u10_n13608 , _u10_n13607 ,_u10_n13606 , _u10_n13605 , _u10_n13604 , _u10_n13603 , _u10_n13602 ,_u10_n13601 , _u10_n13600 , _u10_n13599 , _u10_n13598 , _u10_n13597 ,_u10_n13596 , _u10_n13595 , _u10_n13594 , _u10_n13593 , _u10_n13592 ,_u10_n13591 , _u10_n13590 , _u10_n13589 , _u10_n13588 , _u10_n13587 ,_u10_n13586 , _u10_n13585 , _u10_n13584 , _u10_n13583 , _u10_n13582 ,_u10_n13581 , _u10_n13580 , _u10_n13579 , _u10_n13578 , _u10_n13577 ,_u10_n13576 , _u10_n13575 , _u10_n13574 , _u10_n13573 , _u10_n13572 ,_u10_n13571 , _u10_n13570 , _u10_n13569 , _u10_n13568 , _u10_n13567 ,_u10_n13566 , _u10_n13565 , _u10_n13564 , _u10_n13563 , _u10_n13562 ,_u10_n13561 , _u10_n13560 , _u10_n13559 , _u10_n13558 , _u10_n13557 ,_u10_n13556 , _u10_n13555 , _u10_n13554 , _u10_n13553 , _u10_n13552 ,_u10_n13551 , _u10_n13550 , _u10_n13549 , _u10_n13548 , _u10_n13547 ,_u10_n13546 , _u10_n13545 , _u10_n13544 , _u10_n13543 , _u10_n13542 ,_u10_n13541 , _u10_n13540 , _u10_n13539 , _u10_n13538 , _u10_n13537 ,_u10_n13536 , _u10_n13535 , _u10_n13534 , _u10_n13533 , _u10_n13532 ,_u10_n13531 , _u10_n13530 , _u10_n13529 , _u10_n13528 , _u10_n13527 ,_u10_n13526 , _u10_n13525 , _u10_n13524 , _u10_n13523 , _u10_n13522 ,_u10_n13521 , _u10_n13520 , _u10_n13519 , _u10_n13518 , _u10_n13517 ,_u10_n13516 , _u10_n13515 , _u10_n13514 , _u10_n13513 , _u10_n13512 ,_u10_n13511 , _u10_n13510 , _u10_n13509 , _u10_n13508 , _u10_n13507 ,_u10_n13506 , _u10_n13505 , _u10_n13504 , _u10_n13503 , _u10_n13502 ,_u10_n13501 , _u10_n13500 , _u10_n13499 , _u10_n13498 , _u10_n13497 ,_u10_n13496 , _u10_n13495 , _u10_n13494 , _u10_n13493 , _u10_n13492 ,_u10_n13491 , _u10_n13490 , _u10_n13489 , _u10_n13488 , _u10_n13487 ,_u10_n13486 , _u10_n13485 , _u10_n13484 , _u10_n13483 , _u10_n13482 ,_u10_n13481 , _u10_n13480 , _u10_n13479 , _u10_n13478 , _u10_n13477 ,_u10_n13476 , _u10_n13475 , _u10_n13474 , _u10_n13473 , _u10_n13472 ,_u10_n13471 , _u10_n13470 , _u10_n13469 , _u10_n13468 , _u10_n13467 ,_u10_n13466 , _u10_n13465 , _u10_n13464 , _u10_n13463 , _u10_n13462 ,_u10_n13461 , _u10_n13460 , _u10_n13459 , _u10_n13458 , _u10_n13457 ,_u10_n13456 , _u10_n13455 , _u10_n13454 , _u10_n13453 , _u10_n13452 ,_u10_n13451 , _u10_n13450 , _u10_n13449 , _u10_n13448 , _u10_n13447 ,_u10_n13446 , _u10_n13445 , _u10_n13444 , _u10_n13443 , _u10_n13442 ,_u10_n13441 , _u10_n13440 , _u10_n13439 , _u10_n13438 , _u10_n13437 ,_u10_n13436 , _u10_n13435 , _u10_n13434 , _u10_n13433 , _u10_n13432 ,_u10_n13431 , _u10_n13430 , _u10_n13429 , _u10_n13428 , _u10_n13427 ,_u10_n13426 , _u10_n13425 , _u10_n13424 , _u10_n13423 , _u10_n13422 ,_u10_n13421 , _u10_n13420 , _u10_n13419 , _u10_n13418 , _u10_n13417 ,_u10_n13416 , _u10_n13415 , _u10_n13414 , _u10_n13413 , _u10_n13412 ,_u10_n13411 , _u10_n13410 , _u10_n13409 , _u10_n13408 , _u10_n13407 ,_u10_n13406 , _u10_n13405 , _u10_n13404 , _u10_n13403 , _u10_n13402 ,_u10_n13401 , _u10_n13400 , _u10_n13399 , _u10_n13398 , _u10_n13397 ,_u10_n13396 , _u10_n13395 , _u10_n13394 , _u10_n13393 , _u10_n13392 ,_u10_n13391 , _u10_n13390 , _u10_n13389 , _u10_n13388 , _u10_n13387 ,_u10_n13386 , _u10_n13385 , _u10_n13384 , _u10_n13383 , _u10_n13382 ,_u10_n13381 , _u10_n13380 , _u10_n13379 , _u10_n13378 , _u10_n13377 ,_u10_n13376 , _u10_n13375 , _u10_n13374 , _u10_n13373 , _u10_n13372 ,_u10_n13371 , _u10_n13370 , _u10_n13369 , _u10_n13368 , _u10_n13367 ,_u10_n13366 , _u10_n13365 , _u10_n13364 , _u10_n13363 , _u10_n13362 ,_u10_n13361 , _u10_n13360 , _u10_n13359 , _u10_n13358 , _u10_n13357 ,_u10_n13356 , _u10_n13355 , _u10_n13354 , _u10_n13353 , _u10_n13352 ,_u10_n13351 , _u10_n13350 , _u10_n13349 , _u10_n13348 , _u10_n13347 ,_u10_n13346 , _u10_n13345 , _u10_n13344 , _u10_n13343 , _u10_n13342 ,_u10_n13341 , _u10_n13340 , _u10_n13339 , _u10_n13338 , _u10_n13337 ,_u10_n13336 , _u10_n13335 , _u10_n13334 , _u10_n13333 , _u10_n13332 ,_u10_n13331 , _u10_n13330 , _u10_n13329 , _u10_n13328 , _u10_n13327 ,_u10_n13326 , _u10_n13325 , _u10_n13324 , _u10_n13323 , _u10_n13322 ,_u10_n13321 , _u10_n13320 , _u10_n13319 , _u10_n13318 , _u10_n13317 ,_u10_n13316 , _u10_n13315 , _u10_n13314 , _u10_n13313 , _u10_n13312 ,_u10_n13311 , _u10_n13310 , _u10_n13309 , _u10_n13308 , _u10_n13307 ,_u10_n13306 , _u10_n13305 , _u10_n13304 , _u10_n13303 , _u10_n13302 ,_u10_n13301 , _u10_n13300 , _u10_n13299 , _u10_n13298 , _u10_n13297 ,_u10_n13296 , _u10_n13295 , _u10_n13294 , _u10_n13293 , _u10_n13292 ,_u10_n13291 , _u10_n13290 , _u10_n13289 , _u10_n13288 , _u10_n13287 ,_u10_n13286 , _u10_n13285 , _u10_n13284 , _u10_n13283 , _u10_n13282 ,_u10_n13281 , _u10_n13280 , _u10_n13279 , _u10_n13278 , _u10_n13277 ,_u10_n13276 , _u10_n13275 , _u10_n13274 , _u10_n13273 , _u10_n13272 ,_u10_n13271 , _u10_n13270 , _u10_n13269 , _u10_n13268 , _u10_n13267 ,_u10_n13266 , _u10_n13265 , _u10_n13264 , _u10_n13263 , _u10_n13262 ,_u10_n13261 , _u10_n13260 , _u10_n13259 , _u10_n13258 , _u10_n13257 ,_u10_n13256 , _u10_n13255 , _u10_n13254 , _u10_n13253 , _u10_n13252 ,_u10_n13251 , _u10_n13250 , _u10_n13249 , _u10_n13248 , _u10_n13247 ,_u10_n13246 , _u10_n13245 , _u10_n13244 , _u10_n13243 , _u10_n13242 ,_u10_n13241 , _u10_n13240 , _u10_n13239 , _u10_n13238 , _u10_n13237 ,_u10_n13236 , _u10_n13235 , _u10_n13234 , _u10_n13233 , _u10_n13232 ,_u10_n13231 , _u10_n13230 , _u10_n13229 , _u10_n13228 , _u10_n13227 ,_u10_n13226 , _u10_n13225 , _u10_n13224 , _u10_n13223 , _u10_n13222 ,_u10_n13221 , _u10_n13220 , _u10_n13219 , _u10_n13218 , _u10_n13217 ,_u10_n13216 , _u10_n13215 , _u10_n13214 , _u10_n13213 , _u10_n13212 ,_u10_n13211 , _u10_n13210 , _u10_n13209 , _u10_n13208 , _u10_n13207 ,_u10_n13206 , _u10_n13205 , _u10_n13204 , _u10_n13203 , _u10_n13202 ,_u10_n13201 , _u10_n13200 , _u10_n13199 , _u10_n13198 , _u10_n13197 ,_u10_n13196 , _u10_n13195 , _u10_n13194 , _u10_n13193 , _u10_n13192 ,_u10_n13191 , _u10_n13190 , _u10_n13189 , _u10_n13188 , _u10_n13187 ,_u10_n13186 , _u10_n13185 , _u10_n13184 , _u10_n13183 , _u10_n13182 ,_u10_n13181 , _u10_n13180 , _u10_n13179 , _u10_n13178 , _u10_n13177 ,_u10_n13176 , _u10_n13175 , _u10_n13174 , _u10_n13173 , _u10_n13172 ,_u10_n13171 , _u10_n13170 , _u10_n13169 , _u10_n13168 , _u10_n13167 ,_u10_n13166 , _u10_n13165 , _u10_n13164 , _u10_n13163 , _u10_n13162 ,_u10_n13161 , _u10_n13160 , _u10_n13159 , _u10_n13158 , _u10_n13157 ,_u10_n13156 , _u10_n13155 , _u10_n13154 , _u10_n13153 , _u10_n13152 ,_u10_n13151 , _u10_n13150 , _u10_n13149 , _u10_n13148 , _u10_n13147 ,_u10_n13146 , _u10_n13145 , _u10_n13144 , _u10_n13143 , _u10_n13142 ,_u10_n13141 , _u10_n13140 , _u10_n13139 , _u10_n13138 , _u10_n13137 ,_u10_n13136 , _u10_n13135 , _u10_n13134 , _u10_n13133 , _u10_n13132 ,_u10_n13131 , _u10_n13130 , _u10_n13129 , _u10_n13128 , _u10_n13127 ,_u10_n13126 , _u10_n13125 , _u10_n13124 , _u10_n13123 , _u10_n13122 ,_u10_n13121 , _u10_n13120 , _u10_n13119 , _u10_n13118 , _u10_n13117 ,_u10_n13116 , _u10_n13115 , _u10_n13114 , _u10_n13113 , _u10_n13112 ,_u10_n13111 , _u10_n13110 , _u10_n13109 , _u10_n13108 , _u10_n13107 ,_u10_n13106 , _u10_n13105 , _u10_n13104 , _u10_n13103 , _u10_n13102 ,_u10_n13101 , _u10_n13100 , _u10_n13099 , _u10_n13098 , _u10_n13097 ,_u10_n13096 , _u10_n13095 , _u10_n13094 , _u10_n13093 , _u10_n13092 ,_u10_n13091 , _u10_n13090 , _u10_n13089 , _u10_n13088 , _u10_n13087 ,_u10_n13086 , _u10_n13085 , _u10_n13084 , _u10_n13083 , _u10_n13082 ,_u10_n13081 , _u10_n13080 , _u10_n13079 , _u10_n13078 , _u10_n13077 ,_u10_n13076 , _u10_n13075 , _u10_n13074 , _u10_n13073 , _u10_n13072 ,_u10_n13071 , _u10_n13070 , _u10_n13069 , _u10_n13068 , _u10_n13067 ,_u10_n13066 , _u10_n13065 , _u10_n13064 , _u10_n13063 , _u10_n13062 ,_u10_n13061 , _u10_n13060 , _u10_n13059 , _u10_n13058 , _u10_n13057 ,_u10_n13056 , _u10_n13055 , _u10_n13054 , _u10_n13053 , _u10_n13052 ,_u10_n13051 , _u10_n13050 , _u10_n13049 , _u10_n13048 , _u10_n13047 ,_u10_n13046 , _u10_n13045 , _u10_n13044 , _u10_n13043 , _u10_n13042 ,_u10_n13041 , _u10_n13040 , _u10_n13039 , _u10_n13038 , _u10_n13037 ,_u10_n13036 , _u10_n13035 , _u10_n13034 , _u10_n13033 , _u10_n13032 ,_u10_n13031 , _u10_n13030 , _u10_n13029 , _u10_n13028 , _u10_n13027 ,_u10_n13026 , _u10_n13025 , _u10_n13024 , _u10_n13023 , _u10_n13022 ,_u10_n13021 , _u10_n13020 , _u10_n13019 , _u10_n13018 , _u10_n13017 ,_u10_n13016 , _u10_n13015 , _u10_n13014 , _u10_n13013 , _u10_n13012 ,_u10_n13011 , _u10_n13010 , _u10_n13009 , _u10_n13008 , _u10_n13007 ,_u10_n13006 , _u10_n13005 , _u10_n13004 , _u10_n13003 , _u10_n13002 ,_u10_n13001 , _u10_n13000 , _u10_n12999 , _u10_n12998 , _u10_n12997 ,_u10_n12996 , _u10_n12995 , _u10_n12994 , _u10_n12993 , _u10_n12992 ,_u10_n12991 , _u10_n12990 , _u10_n12989 , _u10_n12988 , _u10_n12987 ,_u10_n12986 , _u10_n12985 , _u10_n12984 , _u10_n12983 , _u10_n12982 ,_u10_n12981 , _u10_n12980 , _u10_n12979 , _u10_n12978 , _u10_n12977 ,_u10_n12976 , _u10_n12975 , _u10_n12974 , _u10_n12973 , _u10_n12972 ,_u10_n12971 , _u10_n12970 , _u10_n12969 , _u10_n12968 , _u10_n12967 ,_u10_n12966 , _u10_n12965 , _u10_n12964 , _u10_n12963 , _u10_n12962 ,_u10_n12961 , _u10_n12960 , _u10_n12959 , _u10_n12958 , _u10_n12957 ,_u10_n12956 , _u10_n12955 , _u10_n12954 , _u10_n12953 , _u10_n12952 ,_u10_n12951 , _u10_n12950 , _u10_n12949 , _u10_n12948 , _u10_n12947 ,_u10_n12946 , _u10_n12945 , _u10_n12944 , _u10_n12943 , _u10_n12942 ,_u10_n12941 , _u10_n12940 , _u10_n12939 , _u10_n12938 , _u10_n12937 ,_u10_n12936 , _u10_n12935 , _u10_n12934 , _u10_n12933 , _u10_n12932 ,_u10_n12931 , _u10_n12930 , _u10_n12929 , _u10_n12928 , _u10_n12927 ,_u10_n12926 , _u10_n12925 , _u10_n12924 , _u10_n12923 , _u10_n12922 ,_u10_n12921 , _u10_n12920 , _u10_n12919 , _u10_n12918 , _u10_n12917 ,_u10_n12916 , _u10_n12915 , _u10_n12914 , _u10_n12913 , _u10_n12912 ,_u10_n12911 , _u10_n12910 , _u10_n12909 , _u10_n12908 , _u10_n12907 ,_u10_n12906 , _u10_n12905 , _u10_n12904 , _u10_n12903 , _u10_n12902 ,_u10_n12901 , _u10_n12900 , _u10_n12899 , _u10_n12898 , _u10_n12897 ,_u10_n12896 , _u10_n12895 , _u10_n12894 , _u10_n12893 , _u10_n12892 ,_u10_n12891 , _u10_n12890 , _u10_n12889 , _u10_n12888 , _u10_n12887 ,_u10_n12886 , _u10_n12885 , _u10_n12884 , _u10_n12883 , _u10_n12882 ,_u10_n12881 , _u10_n12880 , _u10_n12879 , _u10_n12878 , _u10_n12877 ,_u10_n12876 , _u10_n12875 , _u10_n12874 , _u10_n12873 , _u10_n12872 ,_u10_n12871 , _u10_n12870 , _u10_n12869 , _u10_n12868 , _u10_n12867 ,_u10_n12866 , _u10_n12865 , _u10_n12864 , _u10_n12863 , _u10_n12862 ,_u10_n12861 , _u10_n12860 , _u10_n12859 , _u10_n12858 , _u10_n12857 ,_u10_n12856 , _u10_n12855 , _u10_n12854 , _u10_n12853 , _u10_n12852 ,_u10_n12851 , _u10_n12850 , _u10_n12849 , _u10_n12848 , _u10_n12847 ,_u10_n12846 , _u10_n12845 , _u10_n12844 , _u10_n12843 , _u10_n12842 ,_u10_n12841 , _u10_n12840 , _u10_n12839 , _u10_n12838 , _u10_n12837 ,_u10_n12836 , _u10_n12835 , _u10_n12834 , _u10_n12833 , _u10_n12832 ,_u10_n12831 , _u10_n12830 , _u10_n12829 , _u10_n12828 , _u10_n12827 ,_u10_n12826 , _u10_n12825 , _u10_n12824 , _u10_n12823 , _u10_n12822 ,_u10_n12821 , _u10_n12820 , _u10_n12819 , _u10_n12818 , _u10_n12817 ,_u10_n12816 , _u10_n12815 , _u10_n12814 , _u10_n12813 , _u10_n12812 ,_u10_n12811 , _u10_n12810 , _u10_n12809 , _u10_n12808 , _u10_n12807 ,_u10_n12806 , _u10_n12805 , _u10_n12804 , _u10_n12803 , _u10_n12802 ,_u10_n12801 , _u10_n12800 , _u10_n12799 , _u10_n12798 , _u10_n12797 ,_u10_n12796 , _u10_n12795 , _u10_n12794 , _u10_n12793 , _u10_n12792 ,_u10_n12791 , _u10_n12790 , _u10_n12789 , _u10_n12788 , _u10_n12787 ,_u10_n12786 , _u10_n12785 , _u10_n12784 , _u10_n12783 , _u10_n12782 ,_u10_n12781 , _u10_n12780 , _u10_n12779 , _u10_n12778 , _u10_n12777 ,_u10_n12776 , _u10_n12775 , _u10_n12774 , _u10_n12773 , _u10_n12772 ,_u10_n12771 , _u10_n12770 , _u10_n12769 , _u10_n12768 , _u10_n12767 ,_u10_n12766 , _u10_n12765 , _u10_n12764 , _u10_n12763 , _u10_n12762 ,_u10_n12761 , _u10_n12760 , _u10_n12759 , _u10_n12758 , _u10_n12757 ,_u10_n12756 , _u10_n12755 , _u10_n12754 , _u10_n12753 , _u10_n12752 ,_u10_n12751 , _u10_n12750 , _u10_n12749 , _u10_n12748 , _u10_n12747 ,_u10_n12746 , _u10_n12745 , _u10_n12744 , _u10_n12743 , _u10_n12742 ,_u10_n12741 , _u10_n12740 , _u10_n12739 , _u10_n12738 , _u10_n12737 ,_u10_n12736 , _u10_n12735 , _u10_n12734 , _u10_n12733 , _u10_n12732 ,_u10_n12731 , _u10_n12730 , _u10_n12729 , _u10_n12728 , _u10_n12727 ,_u10_n12726 , _u10_n12725 , _u10_n12724 , _u10_n12723 , _u10_n12722 ,_u10_n12721 , _u10_n12720 , _u10_n12719 , _u10_n12718 , _u10_n12717 ,_u10_n12716 , _u10_n12715 , _u10_n12714 , _u10_n12713 , _u10_n12712 ,_u10_n12711 , _u10_n12710 , _u10_n12709 , _u10_n12708 , _u10_n12707 ,_u10_n12706 , _u10_n12705 , _u10_n12704 , _u10_n12703 , _u10_n12702 ,_u10_n12701 , _u10_n12700 , _u10_n12699 , _u10_n12698 , _u10_n12697 ,_u10_n12696 , _u10_n12695 , _u10_n12694 , _u10_n12693 , _u10_n12692 ,_u10_n12691 , _u10_n12690 , _u10_n12689 , _u10_n12688 , _u10_n12687 ,_u10_n12686 , _u10_n12685 , _u10_n12684 , _u10_n12683 , _u10_n12682 ,_u10_n12681 , _u10_n12680 , _u10_n12679 , _u10_n12678 , _u10_n12677 ,_u10_n12676 , _u10_n12675 , _u10_n12674 , _u10_n12673 , _u10_n12672 ,_u10_n12671 , _u10_n12670 , _u10_n12669 , _u10_n12668 , _u10_n12667 ,_u10_n12666 , _u10_n12665 , _u10_n12664 , _u10_n12663 , _u10_n12662 ,_u10_n12661 , _u10_n12660 , _u10_n12659 , _u10_n12658 , _u10_n12657 ,_u10_n12656 , _u10_n12655 , _u10_n12654 , _u10_n12653 , _u10_n12652 ,_u10_n12651 , _u10_n12650 , _u10_n12649 , _u10_n12648 , _u10_n12647 ,_u10_n12646 , _u10_n12645 , _u10_n12644 , _u10_n12643 , _u10_n12642 ,_u10_n12641 , _u10_n12640 , _u10_n12639 , _u10_n12638 , _u10_n12637 ,_u10_n12636 , _u10_n12635 , _u10_n12634 , _u10_n12633 , _u10_n12632 ,_u10_n12631 , _u10_n12630 , _u10_n12629 , _u10_n12628 , _u10_n12627 ,_u10_n12626 , _u10_n12625 , _u10_n12624 , _u10_n12623 , _u10_n12622 ,_u10_n12621 , _u10_n12620 , _u10_n12619 , _u10_n12618 , _u10_n12617 ,_u10_n12616 , _u10_n12615 , _u10_n12614 , _u10_n12613 , _u10_n12612 ,_u10_n12611 , _u10_n12610 , _u10_n12609 , _u10_n12608 , _u10_n12607 ,_u10_n12606 , _u10_n12605 , _u10_n12604 , _u10_n12603 , _u10_n12602 ,_u10_n12601 , _u10_n12600 , _u10_n12599 , _u10_n12598 , _u10_n12597 ,_u10_n12596 , _u10_n12595 , _u10_n12594 , _u10_n12593 , _u10_n12592 ,_u10_n12591 , _u10_n12590 , _u10_n12589 , _u10_n12588 , _u10_n12587 ,_u10_n12586 , _u10_n12585 , _u10_n12584 , _u10_n12583 , _u10_n12582 ,_u10_n12581 , _u10_n12580 , _u10_n12579 , _u10_n12578 , _u10_n12577 ,_u10_n12576 , _u10_n12575 , _u10_n12574 , _u10_n12573 , _u10_n12572 ,_u10_n12571 , _u10_n12570 , _u10_n12569 , _u10_n12568 , _u10_n12567 ,_u10_n12566 , _u10_n12565 , _u10_n12564 , _u10_n12563 , _u10_n12562 ,_u10_n12561 , _u10_n12560 , _u10_n12559 , _u10_n12558 , _u10_n12557 ,_u10_n12556 , _u10_n12555 , _u10_n12554 , _u10_n12553 , _u10_n12552 ,_u10_n12551 , _u10_n12550 , _u10_n12549 , _u10_n12548 , _u10_n12547 ,_u10_n12546 , _u10_n12545 , _u10_n12544 , _u10_n12543 , _u10_n12542 ,_u10_n12541 , _u10_n12540 , _u10_n12539 , _u10_n12538 , _u10_n12537 ,_u10_n12536 , _u10_n12535 , _u10_n12534 , _u10_n12533 , _u10_n12532 ,_u10_n12531 , _u10_n12530 , _u10_n12529 , _u10_n12528 , _u10_n12527 ,_u10_n12526 , _u10_n12525 , _u10_n12524 , _u10_n12523 , _u10_n12522 ,_u10_n12521 , _u10_n12520 , _u10_n12519 , _u10_n12518 , _u10_n12517 ,_u10_n12516 , _u10_n12515 , _u10_n12514 , _u10_n12513 , _u10_n12512 ,_u10_n12511 , _u10_n12510 , _u10_n12509 , _u10_n12508 , _u10_n12507 ,_u10_n12506 , _u10_n12505 , _u10_n12504 , _u10_n12503 , _u10_n12502 ,_u10_n12501 , _u10_n12500 , _u10_n12499 , _u10_n12498 , _u10_n12497 ,_u10_n12496 , _u10_n12495 , _u10_n12494 , _u10_n12493 , _u10_n12492 ,_u10_n12491 , _u10_n12490 , _u10_n12489 , _u10_n12488 , _u10_n12487 ,_u10_n12486 , _u10_n12485 , _u10_n12484 , _u10_n12483 , _u10_n12482 ,_u10_n12481 , _u10_n12480 , _u10_n12479 , _u10_n12478 , _u10_n12477 ,_u10_n12476 , _u10_n12475 , _u10_n12474 , _u10_n12473 , _u10_n12472 ,_u10_n12471 , _u10_n12470 , _u10_n12469 , _u10_n12468 , _u10_n12467 ,_u10_n12466 , _u10_n12465 , _u10_n12464 , _u10_n12463 , _u10_n12462 ,_u10_n12461 , _u10_n12460 , _u10_n12459 , _u10_n12458 , _u10_n12457 ,_u10_n12456 , _u10_n12455 , _u10_n12454 , _u10_n12453 , _u10_n12452 ,_u10_n12451 , _u10_n12450 , _u10_n12449 , _u10_n12448 , _u10_n12447 ,_u10_n12446 , _u10_n12445 , _u10_n12444 , _u10_n12443 , _u10_n12442 ,_u10_n12441 , _u10_n12440 , _u10_n12439 , _u10_n12438 , _u10_n12437 ,_u10_n12436 , _u10_n12435 , _u10_n12434 , _u10_n12433 , _u10_n12432 ,_u10_n12431 , _u10_n12430 , _u10_n12429 , _u10_n12428 , _u10_n12427 ,_u10_n12426 , _u10_n12425 , _u10_n12424 , _u10_n12423 , _u10_n12422 ,_u10_n12421 , _u10_n12420 , _u10_n12419 , _u10_n12418 , _u10_n12417 ,_u10_n12416 , _u10_n12415 , _u10_n12414 , _u10_n12413 , _u10_n12412 ,_u10_n12411 , _u10_n12410 , _u10_n12409 , _u10_n12408 , _u10_n12407 ,_u10_n12406 , _u10_n12405 , _u10_n12404 , _u10_n12403 , _u10_n12402 ,_u10_n12401 , _u10_n12400 , _u10_n12399 , _u10_n12398 , _u10_n12397 ,_u10_n12396 , _u10_n12395 , _u10_n12394 , _u10_n12393 , _u10_n12392 ,_u10_n12391 , _u10_n12390 , _u10_n12389 , _u10_n12388 , _u10_n12387 ,_u10_n12386 , _u10_n12385 , _u10_n12384 , _u10_n12383 , _u10_n12382 ,_u10_n12381 , _u10_n12380 , _u10_n12379 , _u10_n12378 , _u10_n12377 ,_u10_n12376 , _u10_n12375 , _u10_n12374 , _u10_n12373 , _u10_n12372 ,_u10_n12371 , _u10_n12370 , _u10_n12369 , _u10_n12368 , _u10_n12367 ,_u10_n12366 , _u10_n12365 , _u10_n12364 , _u10_n12363 , _u10_n12362 ,_u10_n12361 , _u10_n12360 , _u10_n12359 , _u10_n12358 , _u10_n12357 ,_u10_n12356 , _u10_n12355 , _u10_n12354 , _u10_n12353 , _u10_n12352 ,_u10_n12351 , _u10_n12350 , _u10_n12349 , _u10_n12348 , _u10_n12347 ,_u10_n12346 , _u10_n12345 , _u10_n12344 , _u10_n12343 , _u10_n12342 ,_u10_n12341 , _u10_n12340 , _u10_n12339 , _u10_n12338 , _u10_n12337 ,_u10_n12336 , _u10_n12335 , _u10_n12334 , _u10_n12333 , _u10_n12332 ,_u10_n12331 , _u10_n12330 , _u10_n12329 , _u10_n12328 , _u10_n12327 ,_u10_n12326 , _u10_n12325 , _u10_n12324 , _u10_n12323 , _u10_n12322 ,_u10_n12321 , _u10_n12320 , _u10_n12319 , _u10_n12318 , _u10_n12317 ,_u10_n12316 , _u10_n12315 , _u10_n12314 , _u10_n12313 , _u10_n12312 ,_u10_n12311 , _u10_n12310 , _u10_n12309 , _u10_n12308 , _u10_n12307 ,_u10_n12306 , _u10_n12305 , _u10_n12304 , _u10_n12303 , _u10_n12302 ,_u10_n12301 , _u10_n12300 , _u10_n12299 , _u10_n12298 , _u10_n12297 ,_u10_n12296 , _u10_n12295 , _u10_n12294 , _u10_n12293 , _u10_n12292 ,_u10_n12291 , _u10_n12290 , _u10_n12289 , _u10_n12288 , _u10_n12287 ,_u10_n12286 , _u10_n12285 , _u10_n12284 , _u10_n12283 , _u10_n12282 ,_u10_n12281 , _u10_n12280 , _u10_n12279 , _u10_n12278 , _u10_n12277 ,_u10_n12276 , _u10_n12275 , _u10_n12274 , _u10_n12273 , _u10_n12272 ,_u10_n12271 , _u10_n12270 , _u10_n12269 , _u10_n12268 , _u10_n12267 ,_u10_n12266 , _u10_n12265 , _u10_n12264 , _u10_n12263 , _u10_n12262 ,_u10_n12261 , _u10_n12260 , _u10_n12259 , _u10_n12258 , _u10_n12257 ,_u10_n12256 , _u10_n12255 , _u10_n12254 , _u10_n12253 , _u10_n12252 ,_u10_n12251 , _u10_n12250 , _u10_n12249 , _u10_n12248 , _u10_n12247 ,_u10_n12246 , _u10_n12245 , _u10_n12244 , _u10_n12243 , _u10_n12242 ,_u10_n12241 , _u10_n12240 , _u10_n12239 , _u10_n12238 , _u10_n12237 ,_u10_n12236 , _u10_n12235 , _u10_n12234 , _u10_n12233 , _u10_n12232 ,_u10_n12231 , _u10_n12230 , _u10_n12229 , _u10_n12228 , _u10_n12227 ,_u10_n12226 , _u10_n12225 , _u10_n12224 , _u10_n12223 , _u10_n12222 ,_u10_n12221 , _u10_n12220 , _u10_n12219 , _u10_n12218 , _u10_n12217 ,_u10_n12216 , _u10_n12215 , _u10_n12214 , _u10_n12213 , _u10_n12212 ,_u10_n12211 , _u10_n12210 , _u10_n12209 , _u10_n12208 , _u10_n12207 ,_u10_n12206 , _u10_n12205 , _u10_n12204 , _u10_n12203 , _u10_n12202 ,_u10_n12201 , _u10_n12200 , _u10_n12199 , _u10_n12198 , _u10_n12197 ,_u10_n12196 , _u10_n12195 , _u10_n12194 , _u10_n12193 , _u10_n12192 ,_u10_n12191 , _u10_n12190 , _u10_n12189 , _u10_n12188 , _u10_n12187 ,_u10_n12186 , _u10_n12185 , _u10_n12184 , _u10_n12183 , _u10_n12182 ,_u10_n12181 , _u10_n12180 , _u10_n12179 , _u10_n12178 , _u10_n12177 ,_u10_n12176 , _u10_n12175 , _u10_n12174 , _u10_n12173 , _u10_n12172 ,_u10_n12171 , _u10_n12170 , _u10_n12169 , _u10_n12168 , _u10_n12167 ,_u10_n12166 , _u10_n12165 , _u10_n12164 , _u10_n12163 , _u10_n12162 ,_u10_n12161 , _u10_n12160 , _u10_n12159 , _u10_n12158 , _u10_n12157 ,_u10_n12156 , _u10_n12155 , _u10_n12154 , _u10_n12153 , _u10_n12152 ,_u10_n12151 , _u10_n12150 , _u10_n12149 , _u10_n12148 , _u10_n12147 ,_u10_n12146 , _u10_n12145 , _u10_n12144 , _u10_n12143 , _u10_n12142 ,_u10_n12141 , _u10_n12140 , _u10_n12139 , _u10_n12138 , _u10_n12137 ,_u10_n12136 , _u10_n12135 , _u10_n12134 , _u10_n12133 , _u10_n12132 ,_u10_n12131 , _u10_n12130 , _u10_n12129 , _u10_n12128 , _u10_n12127 ,_u10_n12126 , _u10_n12125 , _u10_n12124 , _u10_n12123 , _u10_n12122 ,_u10_n12121 , _u10_n12120 , _u10_n12119 , _u10_n12118 , _u10_n12117 ,_u10_n12116 , _u10_n12115 , _u10_n12114 , _u10_n12113 , _u10_n12112 ,_u10_n12111 , _u10_n12110 , _u10_n12109 , _u10_n12108 , _u10_n12107 ,_u10_n12106 , _u10_n12105 , _u10_n12104 , _u10_n12103 , _u10_n12102 ,_u10_n12101 , _u10_n12100 , _u10_n12099 , _u10_n12098 , _u10_n12097 ,_u10_n12096 , _u10_n12095 , _u10_n12094 , _u10_n12093 , _u10_n12092 ,_u10_n12091 , _u10_n12090 , _u10_n12089 , _u10_n12088 , _u10_n12087 ,_u10_n12086 , _u10_n12085 , _u10_n12084 , _u10_n12083 , _u10_n12082 ,_u10_n12081 , _u10_n12080 , _u10_n12079 , _u10_n12078 , _u10_n12077 ,_u10_n12076 , _u10_n12075 , _u10_n12074 , _u10_n12073 , _u10_n12072 ,_u10_n12071 , _u10_n12070 , _u10_n12069 , _u10_n12068 , _u10_n12067 ,_u10_n12066 , _u10_n12065 , _u10_n12064 , _u10_n12063 , _u10_n12062 ,_u10_n12061 , _u10_n12060 , _u10_n12059 , _u10_n12058 , _u10_n12057 ,_u10_n12056 , _u10_n12055 , _u10_n12054 , _u10_n12053 , _u10_n12052 ,_u10_n12051 , _u10_n12050 , _u10_n12049 , _u10_n12048 , _u10_n12047 ,_u10_n12046 , _u10_n12045 , _u10_n12044 , _u10_n12043 , _u10_n12042 ,_u10_n12041 , _u10_n12040 , _u10_n12039 , _u10_n12038 , _u10_n12037 ,_u10_n12036 , _u10_n12035 , _u10_n12034 , _u10_n12033 , _u10_n12032 ,_u10_n12031 , _u10_n12030 , _u10_n12029 , _u10_n12028 , _u10_n12027 ,_u10_n12026 , _u10_n12025 , _u10_n12024 , _u10_n12023 , _u10_n12022 ,_u10_n12021 , _u10_n12020 , _u10_n12019 , _u10_n12018 , _u10_n12017 ,_u10_n12016 , _u10_n12015 , _u10_n12014 , _u10_n12013 , _u10_n12012 ,_u10_n12011 , _u10_n12010 , _u10_n12009 , _u10_n12008 , _u10_n12007 ,_u10_n12006 , _u10_n12005 , _u10_n12004 , _u10_n12003 , _u10_n12002 ,_u10_n12001 , _u10_n12000 , _u10_n11999 , _u10_n11998 , _u10_n11997 ,_u10_n11996 , _u10_n11995 , _u10_n11994 , _u10_n11993 , _u10_n11992 ,_u10_n11991 , _u10_n11990 , _u10_n11989 , _u10_n11988 , _u10_n11987 ,_u10_n11986 , _u10_n11985 , _u10_n11984 , _u10_n11983 , _u10_n11982 ,_u10_n11981 , _u10_n11980 , _u10_n11979 , _u10_n11978 , _u10_n11977 ,_u10_n11976 , _u10_n11975 , _u10_n11974 , _u10_n11973 , _u10_n11972 ,_u10_n11971 , _u10_n11970 , _u10_n11969 , _u10_n11968 , _u10_n11967 ,_u10_n11966 , _u10_n11965 , _u10_n11964 , _u10_n11963 , _u10_n11962 ,_u10_n11961 , _u10_n11960 , _u10_n11959 , _u10_n11958 , _u10_n11957 ,_u10_n11956 , _u10_n11955 , _u10_n11954 , _u10_n11953 , _u10_n11952 ,_u10_n11951 , _u10_n11950 , _u10_n11949 , _u10_n11948 , _u10_n11947 ,_u10_n11946 , _u10_n11945 , _u10_n11944 , _u10_n11943 , _u10_n11942 ,_u10_n11941 , _u10_n11940 , _u10_n11939 , _u10_n11938 , _u10_n11937 ,_u10_n11936 , _u10_n11935 , _u10_n11934 , _u10_n11933 , _u10_n11932 ,_u10_n11931 , _u10_n11930 , _u10_n11929 , _u10_n11928 , _u10_n11927 ,_u10_n11926 , _u10_n11925 , _u10_n11924 , _u10_n11923 , _u10_n11922 ,_u10_n11921 , _u10_n11920 , _u10_n11919 , _u10_n11918 , _u10_n11917 ,_u10_n11916 , _u10_n11915 , _u10_n11914 , _u10_n11913 , _u10_n11912 ,_u10_n11911 , _u10_n11910 , _u10_n11909 , _u10_n11908 , _u10_n11907 ,_u10_n11906 , _u10_n11905 , _u10_n11904 , _u10_n11903 , _u10_n11902 ,_u10_n11901 , _u10_n11900 , _u10_n11899 , _u10_n11898 , _u10_n11897 ,_u10_n11896 , _u10_n11895 , _u10_n11894 , _u10_n11893 , _u10_n11892 ,_u10_n11891 , _u10_n11890 , _u10_n11889 , _u10_n11888 , _u10_n11887 ,_u10_n11886 , _u10_n11885 , _u10_n11884 , _u10_n11883 , _u10_n11882 ,_u10_n11881 , _u10_n11880 , _u10_n11879 , _u10_n11878 , _u10_n11877 ,_u10_n11876 , _u10_n11875 , _u10_n11874 , _u10_n11873 , _u10_n11872 ,_u10_n11871 , _u10_n11870 , _u10_n11869 , _u10_n11868 , _u10_n11867 ,_u10_n11866 , _u10_n11865 , _u10_n11864 , _u10_n11863 , _u10_n11862 ,_u10_n11861 , _u10_n11860 , _u10_n11859 , _u10_n11858 , _u10_n11857 ,_u10_n11856 , _u10_n11855 , _u10_n11854 , _u10_n11853 , _u10_n11852 ,_u10_n11851 , _u10_n11850 , _u10_n11849 , _u10_n11848 , _u10_n11847 ,_u10_n11846 , _u10_n11845 , _u10_n11844 , _u10_n11843 , _u10_n11842 ,_u10_n11841 , _u10_n11840 , _u10_n11839 , _u10_n11838 , _u10_n11837 ,_u10_n11836 , _u10_n11835 , _u10_n11834 , _u10_n11833 , _u10_n11832 ,_u10_n11831 , _u10_n11830 , _u10_n11829 , _u10_n11828 , _u10_n11827 ,_u10_n11826 , _u10_n11825 , _u10_n11824 , _u10_n11823 , _u10_n11822 ,_u10_n11821 , _u10_n11820 , _u10_n11819 , _u10_n11818 , _u10_n11817 ,_u10_n11816 , _u10_n11815 , _u10_n11814 , _u10_n11813 , _u10_n11812 ,_u10_n11811 , _u10_n11810 , _u10_n11809 , _u10_n11808 , _u10_n11807 ,_u10_n11806 , _u10_n11805 , _u10_n11804 , _u10_n11803 , _u10_n11802 ,_u10_n11801 , _u10_n11800 , _u10_n11799 , _u10_n11798 , _u10_n11797 ,_u10_n11796 , _u10_n11795 , _u10_n11794 , _u10_n11793 , _u10_n11792 ,_u10_n11791 , _u10_n11790 , _u10_n11789 , _u10_n11788 , _u10_n11787 ,_u10_n11786 , _u10_n11785 , _u10_n11784 , _u10_n11783 , _u10_n11782 ,_u10_n11781 , _u10_n11780 , _u10_n11779 , _u10_n11778 , _u10_n11777 ,_u10_n11776 , _u10_n11775 , _u10_n11774 , _u10_n11773 , _u10_n11772 ,_u10_n11771 , _u10_n11770 , _u10_n11769 , _u10_n11768 , _u10_n11767 ,_u10_n11766 , _u10_n11765 , _u10_n11764 , _u10_n11763 , _u10_n11762 ,_u10_n11761 , _u10_n11760 , _u10_n11759 , _u10_n11758 , _u10_n11757 ,_u10_n11756 , _u10_n11755 , _u10_n11754 , _u10_n11753 , _u10_n11752 ,_u10_n11751 , _u10_n11750 , _u10_n11749 , _u10_n11748 , _u10_n11747 ,_u10_n11746 , _u10_n11745 , _u10_n11744 , _u10_n11743 , _u10_n11742 ,_u10_n11741 , _u10_n11740 , _u10_n11739 , _u10_n11738 , _u10_n11737 ,_u10_n11736 , _u10_n11735 , _u10_n11734 , _u10_n11733 , _u10_n11732 ,_u10_n11731 , _u10_n11730 , _u10_n11729 , _u10_n11728 , _u10_n11727 ,_u10_n11726 , _u10_n11725 , _u10_n11724 , _u10_n11723 , _u10_n11722 ,_u10_n11721 , _u10_n11720 , _u10_n11719 , _u10_n11718 , _u10_n11717 ,_u10_n11716 , _u10_n11715 , _u10_n11714 , _u10_n11713 , _u10_n11712 ,_u10_n11711 , _u10_n11710 , _u10_n11709 , _u10_n11708 , _u10_n11707 ,_u10_n11706 , _u10_n11705 , _u10_n11704 , _u10_n11703 , _u10_n11702 ,_u10_n11701 , _u10_n11700 , _u10_n11699 , _u10_n11698 , _u10_n11697 ,_u10_n11696 , _u10_n11695 , _u10_n11694 , _u10_n11693 , _u10_n11692 ,_u10_n11691 , _u10_n11690 , _u10_n11689 , _u10_n11688 , _u10_n11687 ,_u10_n11686 , _u10_n11685 , _u10_n11684 , _u10_n11683 , _u10_n11682 ,_u10_n11681 , _u10_n11680 , _u10_n11679 , _u10_n11678 , _u10_n11677 ,_u10_n11676 , _u10_n11675 , _u10_n11674 , _u10_n11673 , _u10_n11672 ,_u10_n11671 , _u10_n11670 , _u10_n11669 , _u10_n11668 , _u10_n11667 ,_u10_n11666 , _u10_n11665 , _u10_n11664 , _u10_n11663 , _u10_n11662 ,_u10_n11661 , _u10_n11660 , _u10_n11659 , _u10_n11658 , _u10_n11657 ,_u10_n11656 , _u10_n11655 , _u10_n11654 , _u10_n11653 , _u10_n11652 ,_u10_n11651 , _u10_n11650 , _u10_n11649 , _u10_n11648 , _u10_n11647 ,_u10_n11646 , _u10_n11645 , _u10_n11644 , _u10_n11643 , _u10_n11642 ,_u10_n11641 , _u10_n11640 , _u10_n11639 , _u10_n11638 , _u10_n11637 ,_u10_n11636 , _u10_n11635 , _u10_n11634 , _u10_n11633 , _u10_n11632 ,_u10_n11631 , _u10_n11630 , _u10_n11629 , _u10_n11628 , _u10_n11627 ,_u10_n11626 , _u10_n11625 , _u10_n11624 , _u10_n11623 , _u10_n11622 ,_u10_n11621 , _u10_n11620 , _u10_n11619 , _u10_n11618 , _u10_n11617 ,_u10_n11616 , _u10_ack_o[30] , _u10_ack_o[29] , _u10_ack_o[28] ,_u10_ack_o[27] , _u10_ack_o[26] , _u10_ack_o[25] , _u10_ack_o[24] ,_u10_ack_o[23] , _u10_ack_o[22] , _u10_ack_o[21] , _u10_ack_o[20] ,_u10_ack_o[19] , _u10_ack_o[18] , _u10_ack_o[17] , _u10_ack_o[16] ,_u10_ack_o[15] , _u10_ack_o[14] , _u10_ack_o[13] , _u10_ack_o[12] ,_u10_ack_o[11] , _u10_ack_o[10] , _u10_ack_o[9] , _u10_ack_o[8] ,_u10_ack_o[7] , _u10_ack_o[6] , _u10_ack_o[5] , _u10_ack_o[4] ,_u10_ack_o[3] , _u10_ack_o[2] , _u10_ack_o[1] , _u10_n10665 ,_u10_n10664 , _u10_n10663 , _u10_n10662 , _u10_n24 , _u10_n11552 ,_u10_n11551 , _u10_n11550 , _u10_n11543 , _u10_n11542 , _u10_n11539 ,_u10_n10676 , _u10_n10675 , _u10_n10674 , _u10_n10673 , _u10_n10672 ,_u10_n5 , _u10_gnt_p0_d[0] , _u10_gnt_p0_d[1] , _u10_gnt_p0_d[2] ,_u10_gnt_p0_d[3] , _u10_gnt_p0_d[4] , _u10_req_p1_0_ ,_u10_req_p0_0_ , _u10_N1034 , _u10_N1033 , _u10_N1032 , _u10_N1031 ,_u10_N1030 , _u10_N1029 , _u10_N1028 , _u10_N1027 , _u10_N1026 ,_u10_N1025 , _u10_N1024 , _u10_N1023 , _u10_N1022 , _u10_N1021 ,_u10_N1020 , _u10_N1019 , _u10_N1018 , _u10_N1017 , _u10_N1016 ,_u10_N1015 , _u10_N1014 , _u10_N1013 , _u10_N1012 , _u10_N1011 ,_u10_N1010 , _u10_N1009 , _u10_N1008 , _u10_N1007 , _u10_N1006 ,_u10_N1005 , _u10_N1004 , _u10_N1003 , _u10_N1002 , _u10_N1000 ,_u10_N999 , _u10_N998 , _u10_N997 , _u10_N996 , _u10_N995 ,_u10_N994 , _u10_N993 , _u10_N992 , _u10_N991 , _u10_N990 ,_u10_N989 , _u10_N988 , _u10_N987 , _u10_N986 , _u10_N985 ,_u10_N984 , _u10_N983 , _u10_N982 , _u10_N981 , _u10_N980 ,_u10_N979 , _u10_N978 , _u10_N977 , _u10_N976 , _u10_N975 ,_u10_N974 , _u10_N973 , _u10_N972 , _u10_N971 , _u10_req_r_0_ ,_u10_N967 , _u10_u0_pri_out[2] , _u10_u0_pri_out[1] ,_u10_u0_pri_out[0] , _u10_u0_u0_pri_out[7] , _u10_u0_u0_pri_out[6] ,_u10_u0_u0_pri_out[5] , _u10_u0_u0_pri_out[4] ,_u10_u0_u0_pri_out[3] , _u10_u0_u0_pri_out[2] ,_u10_u0_u0_pri_out[1] , _u10_u0_u0_pri_out[0] ,_u10_u0_u1_pri_out[7] , _u10_u0_u1_pri_out[6] ,_u10_u0_u1_pri_out[5] , _u10_u0_u1_pri_out[4] ,_u10_u0_u1_pri_out[3] , _u10_u0_u1_pri_out[2] ,_u10_u0_u1_pri_out[1] , _u10_u0_u1_pri_out[0] ,_u10_u0_u2_pri_out[7] , _u10_u0_u2_pri_out[6] ,_u10_u0_u2_pri_out[5] , _u10_u0_u2_pri_out[4] ,_u10_u0_u2_pri_out[3] , _u10_u0_u2_pri_out[2] ,_u10_u0_u2_pri_out[1] , _u10_u0_u2_pri_out[0] ,_u10_u0_u3_pri_out[7] , _u10_u0_u3_pri_out[6] ,_u10_u0_u3_pri_out[5] , _u10_u0_u3_pri_out[4] ,_u10_u0_u3_pri_out[3] , _u10_u0_u3_pri_out[2] ,_u10_u0_u3_pri_out[1] , _u10_u0_u3_pri_out[0] ,_u10_u0_u4_pri_out[7] , _u10_u0_u4_pri_out[6] ,_u10_u0_u4_pri_out[5] , _u10_u0_u4_pri_out[4] ,_u10_u0_u4_pri_out[3] , _u10_u0_u4_pri_out[2] ,_u10_u0_u4_pri_out[1] , _u10_u0_u4_pri_out[0] ,_u10_u0_u5_pri_out[7] , _u10_u0_u5_pri_out[6] ,_u10_u0_u5_pri_out[5] , _u10_u0_u5_pri_out[4] ,_u10_u0_u5_pri_out[3] , _u10_u0_u5_pri_out[2] ,_u10_u0_u5_pri_out[1] , _u10_u0_u5_pri_out[0] ,_u10_u0_u6_pri_out[7] , _u10_u0_u6_pri_out[6] ,_u10_u0_u6_pri_out[5] , _u10_u0_u6_pri_out[4] ,_u10_u0_u6_pri_out[3] , _u10_u0_u6_pri_out[2] ,_u10_u0_u6_pri_out[1] , _u10_u0_u6_pri_out[0] ,_u10_u0_u7_pri_out[7] , _u10_u0_u7_pri_out[6] ,_u10_u0_u7_pri_out[5] , _u10_u0_u7_pri_out[4] ,_u10_u0_u7_pri_out[3] , _u10_u0_u7_pri_out[2] ,_u10_u0_u7_pri_out[1] , _u10_u0_u7_pri_out[0] ,_u10_u0_u8_pri_out[7] , _u10_u0_u8_pri_out[6] ,_u10_u0_u8_pri_out[5] , _u10_u0_u8_pri_out[4] ,_u10_u0_u8_pri_out[3] , _u10_u0_u8_pri_out[2] ,_u10_u0_u8_pri_out[1] , _u10_u0_u8_pri_out[0] ,_u10_u0_u9_pri_out[7] , _u10_u0_u9_pri_out[6] ,_u10_u0_u9_pri_out[5] , _u10_u0_u9_pri_out[4] ,_u10_u0_u9_pri_out[3] , _u10_u0_u9_pri_out[2] ,_u10_u0_u9_pri_out[1] , _u10_u0_u9_pri_out[0] ,_u10_u0_u10_pri_out[7] , _u10_u0_u10_pri_out[6] ,_u10_u0_u10_pri_out[5] , _u10_u0_u10_pri_out[4] ,_u10_u0_u10_pri_out[3] , _u10_u0_u10_pri_out[2] ,_u10_u0_u10_pri_out[1] , _u10_u0_u10_pri_out[0] ,_u10_u0_u11_pri_out[7] , _u10_u0_u11_pri_out[6] ,_u10_u0_u11_pri_out[5] , _u10_u0_u11_pri_out[4] ,_u10_u0_u11_pri_out[3] , _u10_u0_u11_pri_out[2] ,_u10_u0_u11_pri_out[1] , _u10_u0_u11_pri_out[0] ,_u10_u0_u12_pri_out[7] , _u10_u0_u12_pri_out[6] ,_u10_u0_u12_pri_out[5] , _u10_u0_u12_pri_out[4] ,_u10_u0_u12_pri_out[3] , _u10_u0_u12_pri_out[2] ,_u10_u0_u12_pri_out[1] , _u10_u0_u12_pri_out[0] ,_u10_u0_u13_pri_out[7] , _u10_u0_u13_pri_out[6] ,_u10_u0_u13_pri_out[5] , _u10_u0_u13_pri_out[4] ,_u10_u0_u13_pri_out[3] , _u10_u0_u13_pri_out[2] ,_u10_u0_u13_pri_out[1] , _u10_u0_u13_pri_out[0] ,_u10_u0_u14_pri_out[7] , _u10_u0_u14_pri_out[6] ,_u10_u0_u14_pri_out[5] , _u10_u0_u14_pri_out[4] ,_u10_u0_u14_pri_out[3] , _u10_u0_u14_pri_out[2] ,_u10_u0_u14_pri_out[1] , _u10_u0_u14_pri_out[0] ,_u10_u0_u15_pri_out[7] , _u10_u0_u15_pri_out[6] ,_u10_u0_u15_pri_out[5] , _u10_u0_u15_pri_out[4] ,_u10_u0_u15_pri_out[3] , _u10_u0_u15_pri_out[2] ,_u10_u0_u15_pri_out[1] , _u10_u0_u15_pri_out[0] ,_u10_u0_u16_pri_out[7] , _u10_u0_u16_pri_out[6] ,_u10_u0_u16_pri_out[5] , _u10_u0_u16_pri_out[4] ,_u10_u0_u16_pri_out[3] , _u10_u0_u16_pri_out[2] ,_u10_u0_u16_pri_out[1] , _u10_u0_u16_pri_out[0] ,_u10_u0_u17_pri_out[7] , _u10_u0_u17_pri_out[6] ,_u10_u0_u17_pri_out[5] , _u10_u0_u17_pri_out[4] ,_u10_u0_u17_pri_out[3] , _u10_u0_u17_pri_out[2] ,_u10_u0_u17_pri_out[1] , _u10_u0_u17_pri_out[0] ,_u10_u0_u18_pri_out[7] , _u10_u0_u18_pri_out[6] ,_u10_u0_u18_pri_out[5] , _u10_u0_u18_pri_out[4] ,_u10_u0_u18_pri_out[3] , _u10_u0_u18_pri_out[2] ,_u10_u0_u18_pri_out[1] , _u10_u0_u18_pri_out[0] ,_u10_u0_u19_pri_out[7] , _u10_u0_u19_pri_out[6] ,_u10_u0_u19_pri_out[5] , _u10_u0_u19_pri_out[4] ,_u10_u0_u19_pri_out[3] , _u10_u0_u19_pri_out[2] ,_u10_u0_u19_pri_out[1] , _u10_u0_u19_pri_out[0] ,_u10_u0_u20_pri_out[7] , _u10_u0_u20_pri_out[6] ,_u10_u0_u20_pri_out[5] , _u10_u0_u20_pri_out[4] ,_u10_u0_u20_pri_out[3] , _u10_u0_u20_pri_out[2] ,_u10_u0_u20_pri_out[1] , _u10_u0_u20_pri_out[0] ,_u10_u0_u21_pri_out[7] , _u10_u0_u21_pri_out[6] ,_u10_u0_u21_pri_out[5] , _u10_u0_u21_pri_out[4] ,_u10_u0_u21_pri_out[3] , _u10_u0_u21_pri_out[2] ,_u10_u0_u21_pri_out[1] , _u10_u0_u21_pri_out[0] ,_u10_u0_u22_pri_out[7] , _u10_u0_u22_pri_out[6] ,_u10_u0_u22_pri_out[5] , _u10_u0_u22_pri_out[4] ,_u10_u0_u22_pri_out[3] , _u10_u0_u22_pri_out[2] ,_u10_u0_u22_pri_out[1] , _u10_u0_u22_pri_out[0] ,_u10_u0_u23_pri_out[7] , _u10_u0_u23_pri_out[6] ,_u10_u0_u23_pri_out[5] , _u10_u0_u23_pri_out[4] ,_u10_u0_u23_pri_out[3] , _u10_u0_u23_pri_out[2] ,_u10_u0_u23_pri_out[1] , _u10_u0_u23_pri_out[0] ,_u10_u0_u24_pri_out[7] , _u10_u0_u24_pri_out[6] ,_u10_u0_u24_pri_out[5] , _u10_u0_u24_pri_out[4] ,_u10_u0_u24_pri_out[3] , _u10_u0_u24_pri_out[2] ,_u10_u0_u24_pri_out[1] , _u10_u0_u24_pri_out[0] ,_u10_u0_u25_pri_out[7] , _u10_u0_u25_pri_out[6] ,_u10_u0_u25_pri_out[5] , _u10_u0_u25_pri_out[4] ,_u10_u0_u25_pri_out[3] , _u10_u0_u25_pri_out[2] ,_u10_u0_u25_pri_out[1] , _u10_u0_u25_pri_out[0] ,_u10_u0_u26_pri_out[7] , _u10_u0_u26_pri_out[6] ,_u10_u0_u26_pri_out[5] , _u10_u0_u26_pri_out[4] ,_u10_u0_u26_pri_out[3] , _u10_u0_u26_pri_out[2] ,_u10_u0_u26_pri_out[1] , _u10_u0_u26_pri_out[0] ,_u10_u0_u27_pri_out[7] , _u10_u0_u27_pri_out[6] ,_u10_u0_u27_pri_out[5] , _u10_u0_u27_pri_out[4] ,_u10_u0_u27_pri_out[3] , _u10_u0_u27_pri_out[2] ,_u10_u0_u27_pri_out[1] , _u10_u0_u27_pri_out[0] ,_u10_u0_u28_pri_out[7] , _u10_u0_u28_pri_out[6] ,_u10_u0_u28_pri_out[5] , _u10_u0_u28_pri_out[4] ,_u10_u0_u28_pri_out[3] , _u10_u0_u28_pri_out[2] ,_u10_u0_u28_pri_out[1] , _u10_u0_u28_pri_out[0] ,_u10_u0_u29_pri_out[7] , _u10_u0_u29_pri_out[6] ,_u10_u0_u29_pri_out[5] , _u10_u0_u29_pri_out[4] ,_u10_u0_u29_pri_out[3] , _u10_u0_u29_pri_out[2] ,_u10_u0_u29_pri_out[1] , _u10_u0_u29_pri_out[0] ,_u10_u0_u30_pri_out[7] , _u10_u0_u30_pri_out[6] ,_u10_u0_u30_pri_out[5] , _u10_u0_u30_pri_out[4] ,_u10_u0_u30_pri_out[3] , _u10_u0_u30_pri_out[2] ,_u10_u0_u30_pri_out[1] , _u10_u0_u30_pri_out[0] , _u10_u1_n3408 ,_u10_u1_n3407 , _u10_u1_n3406 , _u10_u1_n3405 , _u10_u1_n3404 ,_u10_u1_n3403 , _u10_u1_n3402 , _u10_u1_n3401 , _u10_u1_n3400 ,_u10_u1_n3399 , _u10_u1_n3398 , _u10_u1_n3397 , _u10_u1_n3396 ,_u10_u1_n3395 , _u10_u1_n3394 , _u10_u1_n3393 , _u10_u1_n3392 ,_u10_u1_n3391 , _u10_u1_n3390 , _u10_u1_n3389 , _u10_u1_n3388 ,_u10_u1_n3387 , _u10_u1_n3386 , _u10_u1_n3385 , _u10_u1_n3384 ,_u10_u1_n3383 , _u10_u1_n3382 , _u10_u1_n3381 , _u10_u1_n3380 ,_u10_u1_n3379 , _u10_u1_n3378 , _u10_u1_n3377 , _u10_u1_n3376 ,_u10_u1_n3375 , _u10_u1_n3374 , _u10_u1_n3373 , _u10_u1_n3372 ,_u10_u1_n3371 , _u10_u1_n3370 , _u10_u1_n3369 , _u10_u1_n3368 ,_u10_u1_n3367 , _u10_u1_n3366 , _u10_u1_n3365 , _u10_u1_n3364 ,_u10_u1_n3363 , _u10_u1_n3362 , _u10_u1_n3361 , _u10_u1_n3360 ,_u10_u1_n3359 , _u10_u1_n3358 , _u10_u1_n3357 , _u10_u1_n3356 ,_u10_u1_n3355 , _u10_u1_n3354 , _u10_u1_n3353 , _u10_u1_n3352 ,_u10_u1_n3351 , _u10_u1_n3350 , _u10_u1_n3349 , _u10_u1_n3348 ,_u10_u1_n3347 , _u10_u1_n3346 , _u10_u1_n3345 , _u10_u1_n3344 ,_u10_u1_n3343 , _u10_u1_n3342 , _u10_u1_n3341 , _u10_u1_n3340 ,_u10_u1_n3339 , _u10_u1_n3338 , _u10_u1_n3337 , _u10_u1_n3336 ,_u10_u1_n3335 , _u10_u1_n3334 , _u10_u1_n3333 , _u10_u1_n3332 ,_u10_u1_n3331 , _u10_u1_n3330 , _u10_u1_n3329 , _u10_u1_n3328 ,_u10_u1_n3327 , _u10_u1_n3326 , _u10_u1_n3325 , _u10_u1_n3324 ,_u10_u1_n3323 , _u10_u1_n3322 , _u10_u1_n3321 , _u10_u1_n3320 ,_u10_u1_n3319 , _u10_u1_n3318 , _u10_u1_n3317 , _u10_u1_n3316 ,_u10_u1_n3315 , _u10_u1_n3314 , _u10_u1_n3313 , _u10_u1_n3312 ,_u10_u1_n3311 , _u10_u1_n3310 , _u10_u1_n3309 , _u10_u1_n3308 ,_u10_u1_n3307 , _u10_u1_n3306 , _u10_u1_n3305 , _u10_u1_n3304 ,_u10_u1_n3303 , _u10_u1_n3302 , _u10_u1_n3301 , _u10_u1_n3300 ,_u10_u1_n3299 , _u10_u1_n3298 , _u10_u1_n3297 , _u10_u1_n3296 ,_u10_u1_n3295 , _u10_u1_n3294 , _u10_u1_n3293 , _u10_u1_n3292 ,_u10_u1_n3291 , _u10_u1_n3290 , _u10_u1_n3289 , _u10_u1_n3288 ,_u10_u1_n3287 , _u10_u1_n3286 , _u10_u1_n3285 , _u10_u1_n3284 ,_u10_u1_n3283 , _u10_u1_n3282 , _u10_u1_n3281 , _u10_u1_n3280 ,_u10_u1_n3279 , _u10_u1_n3278 , _u10_u1_n3277 , _u10_u1_n3276 ,_u10_u1_n3275 , _u10_u1_n3274 , _u10_u1_n3273 , _u10_u1_n3272 ,_u10_u1_n3271 , _u10_u1_n3270 , _u10_u1_n3269 , _u10_u1_n3268 ,_u10_u1_n3267 , _u10_u1_n3266 , _u10_u1_n3265 , _u10_u1_n3264 ,_u10_u1_n3263 , _u10_u1_n3262 , _u10_u1_n3261 , _u10_u1_n3260 ,_u10_u1_n3259 , _u10_u1_n3258 , _u10_u1_n3257 , _u10_u1_n3256 ,_u10_u1_n3255 , _u10_u1_n3254 , _u10_u1_n3253 , _u10_u1_n3252 ,_u10_u1_n3251 , _u10_u1_n3250 , _u10_u1_n3249 , _u10_u1_n3248 ,_u10_u1_n3247 , _u10_u1_n3246 , _u10_u1_n3245 , _u10_u1_n3244 ,_u10_u1_n3243 , _u10_u1_n3242 , _u10_u1_n3241 , _u10_u1_n3240 ,_u10_u1_n3239 , _u10_u1_n3238 , _u10_u1_n3237 , _u10_u1_n3236 ,_u10_u1_n3235 , _u10_u1_n3234 , _u10_u1_n3233 , _u10_u1_n3232 ,_u10_u1_n3231 , _u10_u1_n3230 , _u10_u1_n3229 , _u10_u1_n3228 ,_u10_u1_n3227 , _u10_u1_n3226 , _u10_u1_n3225 , _u10_u1_n3224 ,_u10_u1_n3223 , _u10_u1_n3222 , _u10_u1_n3221 , _u10_u1_n3220 ,_u10_u1_n3219 , _u10_u1_n3218 , _u10_u1_n3217 , _u10_u1_n3216 ,_u10_u1_n3215 , _u10_u1_n3214 , _u10_u1_n3213 , _u10_u1_n3212 ,_u10_u1_n3211 , _u10_u1_n3210 , _u10_u1_n3209 , _u10_u1_n3208 ,_u10_u1_n3207 , _u10_u1_n3206 , _u10_u1_n3205 , _u10_u1_n3204 ,_u10_u1_n3203 , _u10_u1_n3202 , _u10_u1_n3201 , _u10_u1_n3200 ,_u10_u1_n3199 , _u10_u1_n3198 , _u10_u1_n3197 , _u10_u1_n3196 ,_u10_u1_n3195 , _u10_u1_n3194 , _u10_u1_n3193 , _u10_u1_n3192 ,_u10_u1_n3191 , _u10_u1_n3190 , _u10_u1_n3189 , _u10_u1_n3188 ,_u10_u1_n3187 , _u10_u1_n3186 , _u10_u1_n3185 , _u10_u1_n3184 ,_u10_u1_n3183 , _u10_u1_n3182 , _u10_u1_n3181 , _u10_u1_n3180 ,_u10_u1_n3179 , _u10_u1_n3178 , _u10_u1_n3177 , _u10_u1_n3176 ,_u10_u1_n3175 , _u10_u1_n3174 , _u10_u1_n3173 , _u10_u1_n3172 ,_u10_u1_n3171 , _u10_u1_n3170 , _u10_u1_n3169 , _u10_u1_n3168 ,_u10_u1_n3167 , _u10_u1_n3166 , _u10_u1_n3165 , _u10_u1_n3164 ,_u10_u1_n3163 , _u10_u1_n3162 , _u10_u1_n3161 , _u10_u1_n3160 ,_u10_u1_n3159 , _u10_u1_n3158 , _u10_u1_n3157 , _u10_u1_n3156 ,_u10_u1_n3155 , _u10_u1_n3154 , _u10_u1_n3153 , _u10_u1_n3152 ,_u10_u1_n3151 , _u10_u1_n3150 , _u10_u1_n3149 , _u10_u1_n3148 ,_u10_u1_n3147 , _u10_u1_n3146 , _u10_u1_n3145 , _u10_u1_n3144 ,_u10_u1_n3143 , _u10_u1_n3142 , _u10_u1_n3141 , _u10_u1_n3140 ,_u10_u1_n3139 , _u10_u1_n3138 , _u10_u1_n3137 , _u10_u1_n3136 ,_u10_u1_n3135 , _u10_u1_n3134 , _u10_u1_n3133 , _u10_u1_n3132 ,_u10_u1_n3131 , _u10_u1_n3130 , _u10_u1_n3129 , _u10_u1_n3128 ,_u10_u1_n3127 , _u10_u1_n3126 , _u10_u1_n3125 , _u10_u1_n3124 ,_u10_u1_n3123 , _u10_u1_n3122 , _u10_u1_n3121 , _u10_u1_n3120 ,_u10_u1_n3119 , _u10_u1_n3118 , _u10_u1_n3117 , _u10_u1_n3116 ,_u10_u1_n3115 , _u10_u1_n3114 , _u10_u1_n3113 , _u10_u1_n3112 ,_u10_u1_n3111 , _u10_u1_n3110 , _u10_u1_n3109 , _u10_u1_n3108 ,_u10_u1_n3107 , _u10_u1_n3106 , _u10_u1_n3105 , _u10_u1_n3104 ,_u10_u1_n3103 , _u10_u1_n3102 , _u10_u1_n3101 , _u10_u1_n3100 ,_u10_u1_n3099 , _u10_u1_n3098 , _u10_u1_n3097 , _u10_u1_n3096 ,_u10_u1_n3095 , _u10_u1_n3094 , _u10_u1_n3093 , _u10_u1_n3092 ,_u10_u1_n3091 , _u10_u1_n3090 , _u10_u1_n3089 , _u10_u1_n3088 ,_u10_u1_n3087 , _u10_u1_n3086 , _u10_u1_n3085 , _u10_u1_n3084 ,_u10_u1_n3083 , _u10_u1_n3082 , _u10_u1_n3081 , _u10_u1_n3080 ,_u10_u1_n3079 , _u10_u1_n3078 , _u10_u1_n3077 , _u10_u1_n3076 ,_u10_u1_n3075 , _u10_u1_n3074 , _u10_u1_n3073 , _u10_u1_n3072 ,_u10_u1_n3071 , _u10_u1_n3070 , _u10_u1_n3069 , _u10_u1_n3068 ,_u10_u1_n3067 , _u10_u1_n3066 , _u10_u1_n3065 , _u10_u1_n3064 ,_u10_u1_n3063 , _u10_u1_n3062 , _u10_u1_n3061 , _u10_u1_n3060 ,_u10_u1_n3059 , _u10_u1_n3058 , _u10_u1_n3057 , _u10_u1_n3056 ,_u10_u1_n3055 , _u10_u1_n3054 , _u10_u1_n3053 , _u10_u1_n3052 ,_u10_u1_n3051 , _u10_u1_n3050 , _u10_u1_n3049 , _u10_u1_n3048 ,_u10_u1_n3047 , _u10_u1_n3046 , _u10_u1_n3045 , _u10_u1_n3044 ,_u10_u1_n3043 , _u10_u1_n3042 , _u10_u1_n3041 , _u10_u1_n3040 ,_u10_u1_n3039 , _u10_u1_n3038 , _u10_u1_n3037 , _u10_u1_n3036 ,_u10_u1_n3035 , _u10_u1_n3034 , _u10_u1_n3033 , _u10_u1_n3032 ,_u10_u1_n3031 , _u10_u1_n3030 , _u10_u1_n3029 , _u10_u1_n3028 ,_u10_u1_n3027 , _u10_u1_n3026 , _u10_u1_n3025 , _u10_u1_n3024 ,_u10_u1_n3023 , _u10_u1_n3022 , _u10_u1_n3021 , _u10_u1_n3020 ,_u10_u1_n3019 , _u10_u1_n3018 , _u10_u1_n3017 , _u10_u1_n3016 ,_u10_u1_n3015 , _u10_u1_n3014 , _u10_u1_n3013 , _u10_u1_n3012 ,_u10_u1_n3011 , _u10_u1_n3010 , _u10_u1_n3009 , _u10_u1_n3008 ,_u10_u1_n3007 , _u10_u1_n3006 , _u10_u1_n3005 , _u10_u1_n3004 ,_u10_u1_n3003 , _u10_u1_n3002 , _u10_u1_n3001 , _u10_u1_n3000 ,_u10_u1_n2999 , _u10_u1_n2998 , _u10_u1_n2997 , _u10_u1_n2996 ,_u10_u1_n2995 , _u10_u1_n2994 , _u10_u1_n2993 , _u10_u1_n2992 ,_u10_u1_n2991 , _u10_u1_n2990 , _u10_u1_n2989 , _u10_u1_n2988 ,_u10_u1_n2987 , _u10_u1_n2986 , _u10_u1_n2985 , _u10_u1_n2984 ,_u10_u1_n2983 , _u10_u1_n2982 , _u10_u1_n2981 , _u10_u1_n2980 ,_u10_u1_n2979 , _u10_u1_n2978 , _u10_u1_n2977 , _u10_u1_n2976 ,_u10_u1_n2975 , _u10_u1_n2974 , _u10_u1_n2973 , _u10_u1_n2972 ,_u10_u1_n2971 , _u10_u1_n2970 , _u10_u1_n2969 , _u10_u1_n2968 ,_u10_u1_n2967 , _u10_u1_n2966 , _u10_u1_n2965 , _u10_u1_n2964 ,_u10_u1_n2963 , _u10_u1_n2962 , _u10_u1_n2961 , _u10_u1_n2960 ,_u10_u1_n2959 , _u10_u1_n2958 , _u10_u1_n2957 , _u10_u1_n2956 ,_u10_u1_n2955 , _u10_u1_n2954 , _u10_u1_n2953 , _u10_u1_n2952 ,_u10_u1_n2951 , _u10_u1_n2950 , _u10_u1_n2949 , _u10_u1_n2948 ,_u10_u1_n2947 , _u10_u1_n2946 , _u10_u1_n2945 , _u10_u1_n2944 ,_u10_u1_n2943 , _u10_u1_n2942 , _u10_u1_n2941 , _u10_u1_n2940 ,_u10_u1_n2939 , _u10_u1_n2938 , _u10_u1_n2937 , _u10_u1_n2936 ,_u10_u1_n2935 , _u10_u1_n2934 , _u10_u1_n2933 , _u10_u1_n2932 ,_u10_u1_n2931 , _u10_u1_n2930 , _u10_u1_n2929 , _u10_u1_n2928 ,_u10_u1_n2927 , _u10_u1_n2926 , _u10_u1_n2925 , _u10_u1_n2924 ,_u10_u1_n2923 , _u10_u1_n2922 , _u10_u1_n2921 , _u10_u1_n2920 ,_u10_u1_n2919 , _u10_u1_n2918 , _u10_u1_n2917 , _u10_u1_n2916 ,_u10_u1_n2915 , _u10_u1_n2914 , _u10_u1_n2913 , _u10_u1_n2912 ,_u10_u1_n2911 , _u10_u1_n2910 , _u10_u1_n2909 , _u10_u1_n2908 ,_u10_u1_n2907 , _u10_u1_n2906 , _u10_u1_n2905 , _u10_u1_n2904 ,_u10_u1_n2903 , _u10_u1_n2902 , _u10_u1_n2901 , _u10_u1_n2900 ,_u10_u1_n2899 , _u10_u1_n2898 , _u10_u1_n2897 , _u10_u1_n2896 ,_u10_u1_n2895 , _u10_u1_n2894 , _u10_u1_n2893 , _u10_u1_n2892 ,_u10_u1_n2891 , _u10_u1_n2890 , _u10_u1_n2889 , _u10_u1_n2888 ,_u10_u1_n2887 , _u10_u1_n2886 , _u10_u1_n2885 , _u10_u1_n2884 ,_u10_u1_n2883 , _u10_u1_n2882 , _u10_u1_n2881 , _u10_u1_n2880 ,_u10_u1_n2879 , _u10_u1_n2878 , _u10_u1_n2877 , _u10_u1_n2876 ,_u10_u1_n2875 , _u10_u1_n2874 , _u10_u1_n2873 , _u10_u1_n2872 ,_u10_u1_n2871 , _u10_u1_n2870 , _u10_u1_n2869 , _u10_u1_n2868 ,_u10_u1_n2867 , _u10_u1_n2866 , _u10_u1_n2865 , _u10_u1_n2864 ,_u10_u1_n2863 , _u10_u1_n2862 , _u10_u1_n2861 , _u10_u1_n2860 ,_u10_u1_n2859 , _u10_u1_n2858 , _u10_u1_n2857 , _u10_u1_n2856 ,_u10_u1_n2855 , _u10_u1_n2854 , _u10_u1_n2853 , _u10_u1_n2852 ,_u10_u1_n2851 , _u10_u1_n2850 , _u10_u1_n2849 , _u10_u1_n2848 ,_u10_u1_n2847 , _u10_u1_n2846 , _u10_u1_n2845 , _u10_u1_n2844 ,_u10_u1_n2843 , _u10_u1_n2842 , _u10_u1_n2841 , _u10_u1_n2840 ,_u10_u1_n2839 , _u10_u1_n2838 , _u10_u1_n2837 , _u10_u1_n2836 ,_u10_u1_n2835 , _u10_u1_n2834 , _u10_u1_n2833 , _u10_u1_n2832 ,_u10_u1_n2831 , _u10_u1_n2830 , _u10_u1_n2829 , _u10_u1_n2828 ,_u10_u1_n2827 , _u10_u1_n2826 , _u10_u1_n2825 , _u10_u1_n2824 ,_u10_u1_n2823 , _u10_u1_n2822 , _u10_u1_n2821 , _u10_u1_n2820 ,_u10_u1_n2819 , _u10_u1_n2818 , _u10_u1_n2817 , _u10_u1_n2816 ,_u10_u1_n2815 , _u10_u1_n2814 , _u10_u1_n2813 , _u10_u1_n2812 ,_u10_u1_n2811 , _u10_u1_n2810 , _u10_u1_n2809 , _u10_u1_n2808 ,_u10_u1_n2807 , _u10_u1_n2806 , _u10_u1_n2805 , _u10_u1_n2804 ,_u10_u1_n2803 , _u10_u1_n2802 , _u10_u1_n2801 , _u10_u1_n2800 ,_u10_u1_n2799 , _u10_u1_n2798 , _u10_u1_n2797 , _u10_u1_n2796 ,_u10_u1_n2795 , _u10_u1_n2794 , _u10_u1_n2793 , _u10_u1_n2792 ,_u10_u1_n2791 , _u10_u1_n2790 , _u10_u1_n2789 , _u10_u1_n2788 ,_u10_u1_n2787 , _u10_u1_n2786 , _u10_u1_n2785 , _u10_u1_n2784 ,_u10_u1_n2783 , _u10_u1_n2782 , _u10_u1_n2781 , _u10_u1_n2780 ,_u10_u1_n2779 , _u10_u1_n2778 , _u10_u1_n2777 , _u10_u1_n2776 ,_u10_u1_n2775 , _u10_u1_n2774 , _u10_u1_n2773 , _u10_u1_n2772 ,_u10_u1_n2771 , _u10_u1_n2770 , _u10_u1_n2769 , _u10_u1_n2768 ,_u10_u1_n2767 , _u10_u1_n2766 , _u10_u1_n2765 , _u10_u1_n2764 ,_u10_u1_n2763 , _u10_u1_n2762 , _u10_u1_n2761 , _u10_u1_n2760 ,_u10_u1_n2759 , _u10_u1_n2758 , _u10_u1_n2757 , _u10_u1_n2756 ,_u10_u1_n2755 , _u10_u1_n2754 , _u10_u1_n2753 , _u10_u1_n2752 ,_u10_u1_n2751 , _u10_u1_n2750 , _u10_u1_n2749 , _u10_u1_n2748 ,_u10_u1_n2747 , _u10_u1_n2746 , _u10_u1_n2745 , _u10_u1_n2744 ,_u10_u1_n2743 , _u10_u1_n2742 , _u10_u1_n2741 , _u10_u1_n2740 ,_u10_u1_n2739 , _u10_u1_n2738 , _u10_u1_n2737 , _u10_u1_n2736 ,_u10_u1_n2735 , _u10_u1_n2734 , _u10_u1_n2733 , _u10_u1_n2732 ,_u10_u1_n2731 , _u10_u1_n2730 , _u10_u1_n2729 , _u10_u1_n2728 ,_u10_u1_n2727 , _u10_u1_n2726 , _u10_u1_n2725 , _u10_u1_n2724 ,_u10_u1_n2723 , _u10_u1_n2722 , _u10_u1_n2721 , _u10_u1_n2720 ,_u10_u1_n2719 , _u10_u1_n2718 , _u10_u1_n2717 , _u10_u1_n2716 ,_u10_u1_n2715 , _u10_u1_n2714 , _u10_u1_n2713 , _u10_u1_n2712 ,_u10_u1_n2711 , _u10_u1_n2710 , _u10_u1_n2709 , _u10_u1_n2708 ,_u10_u1_n2707 , _u10_u1_n2706 , _u10_u1_n2705 , _u10_u1_n2704 ,_u10_u1_n2703 , _u10_u1_n2702 , _u10_u1_n2701 , _u10_u1_n2700 ,_u10_u1_n2699 , _u10_u1_n2698 , _u10_u1_n2697 , _u10_u1_n2696 ,_u10_u1_n2695 , _u10_u1_n2694 , _u10_u1_n2693 , _u10_u1_n2692 ,_u10_u1_n2691 , _u10_u1_n2690 , _u10_u1_n2689 , _u10_u1_n2688 ,_u10_u1_n2687 , _u10_u1_n2686 , _u10_u1_n2685 , _u10_u1_n2684 ,_u10_u1_n2683 , _u10_u1_n2682 , _u10_u1_n2681 , _u10_u1_n2680 ,_u10_u1_n2679 , _u10_u1_n2678 , _u10_u1_n2677 , _u10_u1_n2676 ,_u10_u1_n2675 , _u10_u1_n2674 , _u10_u1_n2673 , _u10_u1_n2672 ,_u10_u1_n2671 , _u10_u1_n2670 , _u10_u1_n2669 , _u10_u1_n2668 ,_u10_u1_n2667 , _u10_u1_n2666 , _u10_u1_n2665 , _u10_u1_n2664 ,_u10_u1_n2663 , _u10_u1_n2662 , _u10_u1_n2661 , _u10_u1_n2660 ,_u10_u1_n2659 , _u10_u1_n2658 , _u10_u1_n2657 , _u10_u1_n2656 ,_u10_u1_n2655 , _u10_u1_n2654 , _u10_u1_n2653 , _u10_u1_n2652 ,_u10_u1_n2651 , _u10_u1_n2650 , _u10_u1_n2649 , _u10_u1_n2648 ,_u10_u1_n2647 , _u10_u1_n2646 , _u10_u1_n2645 , _u10_u1_n2644 ,_u10_u1_n2643 , _u10_u1_n2642 , _u10_u1_n2641 , _u10_u1_n2640 ,_u10_u1_n2639 , _u10_u1_n2638 , _u10_u1_n2637 , _u10_u1_n2636 ,_u10_u1_n2635 , _u10_u1_n2634 , _u10_u1_n2633 , _u10_u1_n2632 ,_u10_u1_n2631 , _u10_u1_n2630 , _u10_u1_n2629 , _u10_u1_n2628 ,_u10_u1_n2627 , _u10_u1_n2626 , _u10_u1_n2625 , _u10_u1_n2624 ,_u10_u1_n2623 , _u10_u1_n2622 , _u10_u1_n2621 , _u10_u1_n2620 ,_u10_u1_n2619 , _u10_u1_n2618 , _u10_u1_n2617 , _u10_u1_n2616 ,_u10_u1_n2615 , _u10_u1_n2614 , _u10_u1_n2613 , _u10_u1_n2612 ,_u10_u1_n2611 , _u10_u1_n2610 , _u10_u1_n2609 , _u10_u1_n2608 ,_u10_u1_n2607 , _u10_u1_n2606 , _u10_u1_n2605 , _u10_u1_n2604 ,_u10_u1_n2603 , _u10_u1_n2602 , _u10_u1_n2601 , _u10_u1_n2600 ,_u10_u1_n2599 , _u10_u1_n2598 , _u10_u1_n2597 , _u10_u1_n2596 ,_u10_u1_n2595 , _u10_u1_n2594 , _u10_u1_n2593 , _u10_u1_n2592 ,_u10_u1_n2591 , _u10_u1_n2590 , _u10_u1_n2589 , _u10_u1_n2588 ,_u10_u1_n2587 , _u10_u1_n2586 , _u10_u1_n2585 , _u10_u1_n2584 ,_u10_u1_n2583 , _u10_u1_n2582 , _u10_u1_n2581 , _u10_u1_n2580 ,_u10_u1_n2579 , _u10_u1_n2578 , _u10_u1_n2577 , _u10_u1_n2576 ,_u10_u1_n2575 , _u10_u1_n2574 , _u10_u1_n2573 , _u10_u1_n2572 ,_u10_u1_n2571 , _u10_u1_n2570 , _u10_u1_n2569 , _u10_u1_n2568 ,_u10_u1_n2567 , _u10_u1_n2566 , _u10_u1_n2565 , _u10_u1_n2564 ,_u10_u1_n2563 , _u10_u1_n2562 , _u10_u1_n2561 , _u10_u1_n2560 ,_u10_u1_n2559 , _u10_u1_n2558 , _u10_u1_n2557 , _u10_u1_n2556 ,_u10_u1_n2555 , _u10_u1_n2554 , _u10_u1_n2553 , _u10_u1_n2552 ,_u10_u1_n2551 , _u10_u1_n2550 , _u10_u1_n2549 , _u10_u1_n2548 ,_u10_u1_n2547 , _u10_u1_n2546 , _u10_u1_n2545 , _u10_u1_n2544 ,_u10_u1_n2543 , _u10_u1_n2542 , _u10_u1_n2541 , _u10_u1_n2540 ,_u10_u1_n2539 , _u10_u1_n2538 , _u10_u1_n2537 , _u10_u1_n2536 ,_u10_u1_n2535 , _u10_u1_n2534 , _u10_u1_n2533 , _u10_u1_n2532 ,_u10_u1_n2531 , _u10_u1_n2530 , _u10_u1_n2529 , _u10_u1_n2528 ,_u10_u1_n2527 , _u10_u1_n2526 , _u10_u1_n2525 , _u10_u1_n2524 ,_u10_u1_n2523 , _u10_u1_n2522 , _u10_u1_n2521 , _u10_u1_n2520 ,_u10_u1_n2519 , _u10_u1_n2518 , _u10_u1_n2517 , _u10_u1_n2516 ,_u10_u1_n2515 , _u10_u1_n2514 , _u10_u1_n2513 , _u10_u1_n2512 ,_u10_u1_n2511 , _u10_u1_n2510 , _u10_u1_n2509 , _u10_u1_n2508 ,_u10_u1_n2507 , _u10_u1_n2506 , _u10_u1_n2505 , _u10_u1_n2504 ,_u10_u1_n2503 , _u10_u1_n2502 , _u10_u1_n2501 , _u10_u1_n2500 ,_u10_u1_n2499 , _u10_u1_n2498 , _u10_u1_n2497 , _u10_u1_n2496 ,_u10_u1_n2495 , _u10_u1_n2494 , _u10_u1_n2493 , _u10_u1_n2492 ,_u10_u1_n2491 , _u10_u1_n2490 , _u10_u1_n2489 , _u10_u1_n2488 ,_u10_u1_n2487 , _u10_u1_n2486 , _u10_u1_n2485 , _u10_u1_n2484 ,_u10_u1_n2483 , _u10_u1_n2482 , _u10_u1_n2481 , _u10_u1_n2480 ,_u10_u1_n2479 , _u10_u1_n2478 , _u10_u1_n2477 , _u10_u1_n2476 ,_u10_u1_n2475 , _u10_u1_n2474 , _u10_u1_n2473 , _u10_u1_n2472 ,_u10_u1_n2471 , _u10_u1_n2470 , _u10_u1_n2469 , _u10_u1_n2468 ,_u10_u1_n2467 , _u10_u1_n2466 , _u10_u1_n2465 , _u10_u1_n2464 ,_u10_u1_n2463 , _u10_u1_n2462 , _u10_u1_n2461 , _u10_u1_n2460 ,_u10_u1_n2459 , _u10_u1_n2458 , _u10_u1_n2457 , _u10_u1_n2456 ,_u10_u1_n2455 , _u10_u1_n2454 , _u10_u1_n2453 , _u10_u1_n2452 ,_u10_u1_n2451 , _u10_u1_n2450 , _u10_u1_n2449 , _u10_u1_n2448 ,_u10_u1_n2447 , _u10_u1_n2446 , _u10_u1_n2445 , _u10_u1_n2444 ,_u10_u1_n2443 , _u10_u1_n2442 , _u10_u1_n2441 , _u10_u1_n2440 ,_u10_u1_n2439 , _u10_u1_n2438 , _u10_u1_n2437 , _u10_u1_n2436 ,_u10_u1_n2435 , _u10_u1_n2434 , _u10_u1_n2433 , _u10_u1_n2432 ,_u10_u1_n2431 , _u10_u1_n2430 , _u10_u1_n2429 , _u10_u1_n2428 ,_u10_u1_n2427 , _u10_u1_n2426 , _u10_u1_n2425 , _u10_u1_n2424 ,_u10_u1_n2423 , _u10_u1_n2422 , _u10_u1_n2421 , _u10_u1_n2420 ,_u10_u1_n2419 , _u10_u1_n2418 , _u10_u1_n2417 , _u10_u1_n2416 ,_u10_u1_n2415 , _u10_u1_n2414 , _u10_u1_n2413 , _u10_u1_n2412 ,_u10_u1_n2411 , _u10_u1_n2410 , _u10_u1_n2409 , _u10_u1_n2408 ,_u10_u1_n2407 , _u10_u1_n2406 , _u10_u1_n2405 , _u10_u1_n2404 ,_u10_u1_n2403 , _u10_u1_n2402 , _u10_u1_n2401 , _u10_u1_n2400 ,_u10_u1_n2399 , _u10_u1_n2398 , _u10_u1_n2397 , _u10_u1_n2396 ,_u10_u1_n2395 , _u10_u1_n2394 , _u10_u1_n2393 , _u10_u1_n2392 ,_u10_u1_n2391 , _u10_u1_n2390 , _u10_u1_n2389 , _u10_u1_n2388 ,_u10_u1_n2387 , _u10_u1_n2386 , _u10_u1_n2385 , _u10_u1_n2384 ,_u10_u1_n2383 , _u10_u1_n2382 , _u10_u1_n2381 , _u10_u1_n2380 ,_u10_u1_n2379 , _u10_u1_n2378 , _u10_u1_n2377 , _u10_u1_n2376 ,_u10_u1_n2375 , _u10_u1_n2374 , _u10_u1_n2373 , _u10_u1_n2372 ,_u10_u1_n2371 , _u10_u1_n2370 , _u10_u1_n2369 , _u10_u1_n2368 ,_u10_u1_n2367 , _u10_u1_n2366 , _u10_u1_n2365 , _u10_u1_n2364 ,_u10_u1_n2363 , _u10_u1_n2362 , _u10_u1_n2361 , _u10_u1_n2360 ,_u10_u1_n2359 , _u10_u1_n2358 , _u10_u1_n2357 , _u10_u1_n2356 ,_u10_u1_n2355 , _u10_u1_n2354 , _u10_u1_n2353 , _u10_u1_n2352 ,_u10_u1_n2351 , _u10_u1_n2350 , _u10_u1_n2349 , _u10_u1_n2348 ,_u10_u1_n2347 , _u10_u1_n2346 , _u10_u1_n2345 , _u10_u1_n2344 ,_u10_u1_n2343 , _u10_u1_n2342 , _u10_u1_n2341 , _u10_u1_n2340 ,_u10_u1_n2339 , _u10_u1_n2338 , _u10_u1_n2337 , _u10_u1_n2336 ,_u10_u1_n2335 , _u10_u1_n2334 , _u10_u1_n2333 , _u10_u1_n2332 ,_u10_u1_n2331 , _u10_u1_n2330 , _u10_u1_n2329 , _u10_u1_n2328 ,_u10_u1_n2327 , _u10_u1_n2326 , _u10_u1_n2325 , _u10_u1_n2324 ,_u10_u1_n2323 , _u10_u1_n2322 , _u10_u1_n2321 , _u10_u1_n2320 ,_u10_u1_n2319 , _u10_u1_n2318 , _u10_u1_n2317 , _u10_u1_n2316 ,_u10_u1_n2315 , _u10_u1_n2314 , _u10_u1_n2313 , _u10_u1_n2312 ,_u10_u1_n2311 , _u10_u1_n2310 , _u10_u1_n2309 , _u10_u1_n2308 ,_u10_u1_n2307 , _u10_u1_n2306 , _u10_u1_n2305 , _u10_u1_n2304 ,_u10_u1_n2303 , _u10_u1_n2302 , _u10_u1_n2301 , _u10_u1_n2300 ,_u10_u1_n2299 , _u10_u1_n2298 , _u10_u1_n2297 , _u10_u1_n2296 ,_u10_u1_n2295 , _u10_u1_n2294 , _u10_u1_n2293 , _u10_u1_n2292 ,_u10_u1_n2291 , _u10_u1_n2290 , _u10_u1_n2289 , _u10_u1_n2288 ,_u10_u1_n2287 , _u10_u1_n2286 , _u10_u1_n2285 , _u10_u1_n2284 ,_u10_u1_n2283 , _u10_u1_n2282 , _u10_u1_n2281 , _u10_u1_n2280 ,_u10_u1_n2279 , _u10_u1_n2278 , _u10_u1_n2277 , _u10_u1_n2276 ,_u10_u1_n2275 , _u10_u1_n2274 , _u10_u1_n2273 , _u10_u1_n2272 ,_u10_u1_n2271 , _u10_u1_n2270 , _u10_u1_n2269 , _u10_u1_n2268 ,_u10_u1_n2267 , _u10_u1_n2266 , _u10_u1_n2265 , _u10_u1_n2264 ,_u10_u1_n2263 , _u10_u1_n2262 , _u10_u1_n2261 , _u10_u1_n2260 ,_u10_u1_n2259 , _u10_u1_n2258 , _u10_u1_n2257 , _u10_u1_n2256 ,_u10_u1_n2255 , _u10_u1_n2254 , _u10_u1_n2253 , _u10_u1_n2252 ,_u10_u1_n2251 , _u10_u1_n2250 , _u10_u1_n2249 , _u10_u1_n2248 ,_u10_u1_n2247 , _u10_u1_n2246 , _u10_u1_n2245 , _u10_u1_n2244 ,_u10_u1_n2243 , _u10_u1_n2242 , _u10_u1_n2241 , _u10_u1_n2240 ,_u10_u1_n2239 , _u10_u1_n2238 , _u10_u1_n2237 , _u10_u1_n2236 ,_u10_u1_n2235 , _u10_u1_n2234 , _u10_u1_n2233 , _u10_u1_n2232 ,_u10_u1_n2231 , _u10_u1_n2230 , _u10_u1_n2229 , _u10_u1_n2228 ,_u10_u1_n2227 , _u10_u1_n2226 , _u10_u1_n2225 , _u10_u1_n2224 ,_u10_u1_n2223 , _u10_u1_n2222 , _u10_u1_n2221 , _u10_u1_n2220 ,_u10_u1_n2219 , _u10_u1_n2218 , _u10_u1_n2217 , _u10_u1_n2216 ,_u10_u1_n2215 , _u10_u1_n2214 , _u10_u1_n2213 , _u10_u1_n2212 ,_u10_u1_n2211 , _u10_u1_n2210 , _u10_u1_n2209 , _u10_u1_n2208 ,_u10_u1_n2207 , _u10_u1_n2206 , _u10_u1_n2205 , _u10_u1_n2204 ,_u10_u1_n2203 , _u10_u1_n2202 , _u10_u1_n2201 , _u10_u1_n2200 ,_u10_u1_n2199 , _u10_u1_n2198 , _u10_u1_n2197 , _u10_u1_n2196 ,_u10_u1_n2195 , _u10_u1_n2194 , _u10_u1_n2193 , _u10_u1_n2192 ,_u10_u1_n2191 , _u10_u1_n2190 , _u10_u1_n2189 , _u10_u1_n2188 ,_u10_u1_n2187 , _u10_u1_n2186 , _u10_u1_n2185 , _u10_u1_n2184 ,_u10_u1_n2183 , _u10_u1_n2182 , _u10_u1_n2181 , _u10_u1_n2180 ,_u10_u1_n2179 , _u10_u1_n2178 , _u10_u1_n2177 , _u10_u1_n2176 ,_u10_u1_n2175 , _u10_u1_n2174 , _u10_u1_n2173 , _u10_u1_n2172 ,_u10_u1_n2171 , _u10_u1_n2170 , _u10_u1_n2169 , _u10_u1_n2168 ,_u10_u1_n2167 , _u10_u1_n2166 , _u10_u1_n2165 , _u10_u1_n2164 ,_u10_u1_n2163 , _u10_u1_n2162 , _u10_u1_n2161 , _u10_u1_n2160 ,_u10_u1_n2159 , _u10_u1_n2158 , _u10_u1_n2157 , _u10_u1_n2156 ,_u10_u1_n2155 , _u10_u1_n2154 , _u10_u1_n2153 , _u10_u1_n2152 ,_u10_u1_n2151 , _u10_u1_n2150 , _u10_u1_n2149 , _u10_u1_n2148 ,_u10_u1_n2147 , _u10_u1_n2146 , _u10_u1_n2145 , _u10_u1_n2144 ,_u10_u1_n2143 , _u10_u1_n2142 , _u10_u1_n2141 , _u10_u1_n2140 ,_u10_u1_n2139 , _u10_u1_n2138 , _u10_u1_n2137 , _u10_u1_n2136 ,_u10_u1_n2135 , _u10_u1_n2134 , _u10_u1_n2133 , _u10_u1_n2132 ,_u10_u1_n2131 , _u10_u1_n2130 , _u10_u1_n2129 , _u10_u1_n2128 ,_u10_u1_n2127 , _u10_u1_n2126 , _u10_u1_n2125 , _u10_u1_n2124 ,_u10_u1_n2123 , _u10_u1_n2122 , _u10_u1_n2121 , _u10_u1_n2120 ,_u10_u1_n2119 , _u10_u1_n2118 , _u10_u1_n2117 , _u10_u1_n2116 ,_u10_u1_n2115 , _u10_u1_n2114 , _u10_u1_n2113 , _u10_u1_n2112 ,_u10_u1_n2111 , _u10_u1_n2110 , _u10_u1_n2109 , _u10_u1_n2108 ,_u10_u1_n2107 , _u10_u1_n2106 , _u10_u1_n2105 , _u10_u1_n2104 ,_u10_u1_n2103 , _u10_u1_n2102 , _u10_u1_n2101 , _u10_u1_n2100 ,_u10_u1_n2099 , _u10_u1_n2098 , _u10_u1_n2097 , _u10_u1_n2096 ,_u10_u1_n2095 , _u10_u1_n2094 , _u10_u1_n2093 , _u10_u1_n2092 ,_u10_u1_n2091 , _u10_u1_n2090 , _u10_u1_n2089 , _u10_u1_n2088 ,_u10_u1_n2087 , _u10_u1_n2086 , _u10_u1_n2085 , _u10_u1_n2084 ,_u10_u1_n2083 , _u10_u1_n2082 , _u10_u1_n2081 , _u10_u1_n2080 ,_u10_u1_n2079 , _u10_u1_n2078 , _u10_u1_n2077 , _u10_u1_n2076 ,_u10_u1_n2075 , _u10_u1_n2074 , _u10_u1_n2073 , _u10_u1_n2072 ,_u10_u1_n2071 , _u10_u1_n2070 , _u10_u1_n2069 , _u10_u1_n2068 ,_u10_u1_n2067 , _u10_u1_n2066 , _u10_u1_n2065 , _u10_u1_n2064 ,_u10_u1_n2063 , _u10_u1_n2062 , _u10_u1_n2061 , _u10_u1_n2060 ,_u10_u1_n2059 , _u10_u1_n2058 , _u10_u1_n2057 , _u10_u1_n2056 ,_u10_u1_n2055 , _u10_u1_n2054 , _u10_u1_n2053 , _u10_u1_n2052 ,_u10_u1_n2051 , _u10_u1_n2050 , _u10_u1_n2049 , _u10_u1_n2048 ,_u10_u1_n2047 , _u10_u1_n2046 , _u10_u1_n2045 , _u10_u1_n2044 ,_u10_u1_n2043 , _u10_u1_n2042 , _u10_u1_n2041 , _u10_u1_n2040 ,_u10_u1_n2039 , _u10_u1_n2038 , _u10_u1_n2037 , _u10_u1_n2036 ,_u10_u1_n2035 , _u10_u1_n2034 , _u10_u1_n2033 , _u10_u1_n2032 ,_u10_u1_n2031 , _u10_u1_n2030 , _u10_u1_n2029 , _u10_u1_n2028 ,_u10_u1_n2027 , _u10_u1_n2026 , _u10_u1_n2025 , _u10_u1_n2024 ,_u10_u1_n2023 , _u10_u1_n2022 , _u10_u1_n2021 , _u10_u1_n2020 ,_u10_u1_n2019 , _u10_u1_n2018 , _u10_u1_n2017 , _u10_u1_n2016 ,_u10_u1_n2015 , _u10_u1_n2014 , _u10_u1_n2013 , _u10_u1_n2012 ,_u10_u1_n2011 , _u10_u1_n2010 , _u10_u1_n2009 , _u10_u1_n2008 ,_u10_u1_n2007 , _u10_u1_n2006 , _u10_u1_n2005 , _u10_u1_n2004 ,_u10_u1_n2003 , _u10_u1_n1997 , _u10_u1_n1996 , _u10_u1_n1995 ,_u10_u1_n1994 , _u10_u1_n1993 , _u10_u1_n1992 , _u10_u1_n1991 ,_u10_u1_n1990 , _u10_u1_n1989 , _u10_u1_n1988 , _u10_u1_n1987 ,_u10_u1_n1986 , _u10_u1_n1985 , _u10_u1_n1984 , _u10_u1_n1983 ,_u10_u1_n1982 , _u10_u1_n1981 , _u10_u1_n1980 , _u10_u1_n1979 ,_u10_u1_n1978 , _u10_u1_n1977 , _u10_u1_n1976 , _u10_u1_n1975 ,_u10_u1_n1974 , _u10_u1_n1973 , _u10_u1_n1972 , _u10_u1_n1971 ,_u10_u1_n1970 , _u10_u1_n1969 , _u10_u1_n1968 , _u10_u1_n1967 ,_u10_u1_n1966 , _u10_u1_n1965 , _u10_u1_n1964 , _u10_u1_n1963 ,_u10_u1_n1962 , _u10_u1_n1961 , _u10_u1_n1960 , _u10_u1_n1959 ,_u10_u1_n1958 , _u10_u1_n1957 , _u10_u1_n1956 , _u10_u1_n1955 ,_u10_u1_n1954 , _u10_u1_n1953 , _u10_u1_n1952 , _u10_u1_n1951 ,_u10_u1_n1950 , _u10_u1_n1949 , _u10_u1_n1948 , _u10_u1_n1947 ,_u10_u1_n1946 , _u10_u1_n1945 , _u10_u1_n1944 , _u10_u1_n1943 ,_u10_u1_n1942 , _u10_u1_n1941 , _u10_u1_n1940 , _u10_u1_n1939 ,_u10_u1_n1938 , _u10_u1_n1937 , _u10_u1_n1936 , _u10_u1_n1935 ,_u10_u1_n1934 , _u10_u1_n1933 , _u10_u1_n1932 , _u10_u1_n1931 ,_u10_u1_n1930 , _u10_u1_n1929 , _u10_u1_n1928 , _u10_u1_n1927 ,_u10_u1_n1926 , _u10_u1_n1925 , _u10_u1_n1924 , _u10_u1_n1923 ,_u10_u1_n1922 , _u10_u1_n1921 , _u10_u1_n1920 , _u10_u1_n1919 ,_u10_u1_n1918 , _u10_u1_n1917 , _u10_u1_n1916 , _u10_u1_n1915 ,_u10_u1_n1914 , _u10_u1_n1913 , _u10_u1_n1912 , _u10_u1_n1911 ,_u10_u1_n1910 , _u10_u1_n1909 , _u10_u1_n1908 , _u10_u1_n1907 ,_u10_u1_n1906 , _u10_u1_n1905 , _u10_u1_n1904 , _u10_u1_n1903 ,_u10_u1_n1902 , _u10_u1_n1901 , _u10_u1_n1900 , _u10_u1_n1899 ,_u10_u1_n1898 , _u10_u1_n1897 , _u10_u1_n1896 , _u10_u1_n1895 ,_u10_u1_n1894 , _u10_u1_n1893 , _u10_u1_n1892 , _u10_u1_n1891 ,_u10_u1_n1890 , _u10_u1_n1889 , _u10_u1_n1888 , _u10_u1_n1887 ,_u10_u1_n1886 , _u10_u1_n1885 , _u10_u1_n1884 , _u10_u1_n1883 ,_u10_u1_n1882 , _u10_u1_n1881 , _u10_u1_n1880 , _u10_u1_n1879 ,_u10_u1_n1878 , _u10_u1_n1877 , _u10_u1_n1876 , _u10_u1_n1875 ,_u10_u1_n1874 , _u10_u1_n1873 , _u10_u1_n1872 , _u10_u1_n1871 ,_u10_u1_n1870 , _u10_u1_n1869 , _u10_u1_n1868 , _u10_u1_n1867 ,_u10_u1_n1866 , _u10_u1_n1865 , _u10_u1_n1864 , _u10_u1_n1863 ,_u10_u1_n1862 , _u10_u1_n1861 , _u10_u1_n1860 , _u10_u1_n1859 ,_u10_u1_n1858 , _u10_u1_n1857 , _u10_u1_n1856 , _u10_u1_n1855 ,_u10_u1_n1854 , _u10_u1_n1853 , _u10_u1_n1852 , _u10_u1_n1851 ,_u10_u1_n1850 , _u10_u1_n1849 , _u10_u1_n1848 , _u10_u1_n1847 ,_u10_u1_n1846 , _u10_u1_n1845 , _u10_u1_n1844 , _u10_u1_n1843 ,_u10_u1_n1842 , _u10_u1_n1841 , _u10_u1_n1840 , _u10_u1_n1839 ,_u10_u1_n1838 , _u10_u1_n1837 , _u10_u1_n1836 , _u10_u1_n1835 ,_u10_u1_n1834 , _u10_u1_n1833 , _u10_u1_n1832 , _u10_u1_n1831 ,_u10_u1_n1830 , _u10_u1_n1829 , _u10_u1_n1828 , _u10_u1_n1827 ,_u10_u1_n1826 , _u10_u1_n1825 , _u10_u1_n1824 , _u10_u1_n1823 ,_u10_u1_n1822 , _u10_u1_n1821 , _u10_u1_n1820 , _u10_u1_n1819 ,_u10_u1_n1818 , _u10_u1_n1817 , _u10_u1_n1816 , _u10_u1_n1815 ,_u10_u1_n1814 , _u10_u1_n1813 , _u10_u1_n1812 , _u10_u1_n1811 ,_u10_u1_n1810 , _u10_u1_n1809 , _u10_u1_n1808 , _u10_u1_n2002 ,_u10_u1_n2001 , _u10_u1_n2000 , _u10_u1_n1999 , _u10_u1_n1998 ,_u10_u1_n15 , _u10_u1_n14 , _u10_u1_n13 , _u10_u1_n12 , _u10_u1_n10 ,_u10_u20_n3416 , _u10_u20_n3415 , _u10_u20_n3414 , _u10_u20_n3413 ,_u10_u20_n3412 , _u10_u20_n3411 , _u10_u20_n3410 , _u10_u20_n3409 ,_u10_u20_n3408 , _u10_u20_n3407 , _u10_u20_n3406 , _u10_u20_n3405 ,_u10_u20_n3404 , _u10_u20_n3403 , _u10_u20_n3402 , _u10_u20_n3401 ,_u10_u20_n3400 , _u10_u20_n3399 , _u10_u20_n3398 , _u10_u20_n3397 ,_u10_u20_n3396 , _u10_u20_n3395 , _u10_u20_n3394 , _u10_u20_n3393 ,_u10_u20_n3392 , _u10_u20_n3391 , _u10_u20_n3390 , _u10_u20_n3389 ,_u10_u20_n3388 , _u10_u20_n3387 , _u10_u20_n3386 , _u10_u20_n3385 ,_u10_u20_n3384 , _u10_u20_n3383 , _u10_u20_n3382 , _u10_u20_n3381 ,_u10_u20_n3380 , _u10_u20_n3379 , _u10_u20_n3378 , _u10_u20_n3377 ,_u10_u20_n3376 , _u10_u20_n3375 , _u10_u20_n3374 , _u10_u20_n3373 ,_u10_u20_n3372 , _u10_u20_n3371 , _u10_u20_n3370 , _u10_u20_n3369 ,_u10_u20_n3368 , _u10_u20_n3367 , _u10_u20_n3366 , _u10_u20_n3365 ,_u10_u20_n3364 , _u10_u20_n3363 , _u10_u20_n3362 , _u10_u20_n3361 ,_u10_u20_n3360 , _u10_u20_n3359 , _u10_u20_n3358 , _u10_u20_n3357 ,_u10_u20_n3356 , _u10_u20_n3355 , _u10_u20_n3354 , _u10_u20_n3353 ,_u10_u20_n3352 , _u10_u20_n3351 , _u10_u20_n3350 , _u10_u20_n3349 ,_u10_u20_n3348 , _u10_u20_n3347 , _u10_u20_n3346 , _u10_u20_n3345 ,_u10_u20_n3344 , _u10_u20_n3343 , _u10_u20_n3342 , _u10_u20_n3341 ,_u10_u20_n3340 , _u10_u20_n3339 , _u10_u20_n3338 , _u10_u20_n3337 ,_u10_u20_n3336 , _u10_u20_n3335 , _u10_u20_n3334 , _u10_u20_n3333 ,_u10_u20_n3332 , _u10_u20_n3331 , _u10_u20_n3330 , _u10_u20_n3329 ,_u10_u20_n3328 , _u10_u20_n3327 , _u10_u20_n3326 , _u10_u20_n3325 ,_u10_u20_n3324 , _u10_u20_n3323 , _u10_u20_n3322 , _u10_u20_n3321 ,_u10_u20_n3320 , _u10_u20_n3319 , _u10_u20_n3318 , _u10_u20_n3317 ,_u10_u20_n3316 , _u10_u20_n3315 , _u10_u20_n3314 , _u10_u20_n3313 ,_u10_u20_n3312 , _u10_u20_n3311 , _u10_u20_n3310 , _u10_u20_n3309 ,_u10_u20_n3308 , _u10_u20_n3307 , _u10_u20_n3306 , _u10_u20_n3305 ,_u10_u20_n3304 , _u10_u20_n3303 , _u10_u20_n3302 , _u10_u20_n3301 ,_u10_u20_n3300 , _u10_u20_n3299 , _u10_u20_n3298 , _u10_u20_n3297 ,_u10_u20_n3296 , _u10_u20_n3295 , _u10_u20_n3294 , _u10_u20_n3293 ,_u10_u20_n3292 , _u10_u20_n3291 , _u10_u20_n3290 , _u10_u20_n3289 ,_u10_u20_n3288 , _u10_u20_n3287 , _u10_u20_n3286 , _u10_u20_n3285 ,_u10_u20_n3284 , _u10_u20_n3283 , _u10_u20_n3282 , _u10_u20_n3281 ,_u10_u20_n3280 , _u10_u20_n3279 , _u10_u20_n3278 , _u10_u20_n3277 ,_u10_u20_n3276 , _u10_u20_n3275 , _u10_u20_n3274 , _u10_u20_n3273 ,_u10_u20_n3272 , _u10_u20_n3271 , _u10_u20_n3270 , _u10_u20_n3269 ,_u10_u20_n3268 , _u10_u20_n3267 , _u10_u20_n3266 , _u10_u20_n3265 ,_u10_u20_n3264 , _u10_u20_n3263 , _u10_u20_n3262 , _u10_u20_n3261 ,_u10_u20_n3260 , _u10_u20_n3259 , _u10_u20_n3258 , _u10_u20_n3257 ,_u10_u20_n3256 , _u10_u20_n3255 , _u10_u20_n3254 , _u10_u20_n3253 ,_u10_u20_n3252 , _u10_u20_n3251 , _u10_u20_n3250 , _u10_u20_n3249 ,_u10_u20_n3248 , _u10_u20_n3247 , _u10_u20_n3246 , _u10_u20_n3245 ,_u10_u20_n3244 , _u10_u20_n3243 , _u10_u20_n3242 , _u10_u20_n3241 ,_u10_u20_n3240 , _u10_u20_n3239 , _u10_u20_n3238 , _u10_u20_n3237 ,_u10_u20_n3236 , _u10_u20_n3235 , _u10_u20_n3234 , _u10_u20_n3233 ,_u10_u20_n3232 , _u10_u20_n3231 , _u10_u20_n3230 , _u10_u20_n3229 ,_u10_u20_n3228 , _u10_u20_n3227 , _u10_u20_n3226 , _u10_u20_n3225 ,_u10_u20_n3224 , _u10_u20_n3223 , _u10_u20_n3222 , _u10_u20_n3221 ,_u10_u20_n3220 , _u10_u20_n3219 , _u10_u20_n3218 , _u10_u20_n3217 ,_u10_u20_n3216 , _u10_u20_n3215 , _u10_u20_n3214 , _u10_u20_n3213 ,_u10_u20_n3212 , _u10_u20_n3211 , _u10_u20_n3210 , _u10_u20_n3209 ,_u10_u20_n3208 , _u10_u20_n3207 , _u10_u20_n3206 , _u10_u20_n3205 ,_u10_u20_n3204 , _u10_u20_n3203 , _u10_u20_n3202 , _u10_u20_n3201 ,_u10_u20_n3200 , _u10_u20_n3199 , _u10_u20_n3198 , _u10_u20_n3197 ,_u10_u20_n3196 , _u10_u20_n3195 , _u10_u20_n3194 , _u10_u20_n3193 ,_u10_u20_n3192 , _u10_u20_n3191 , _u10_u20_n3190 , _u10_u20_n3189 ,_u10_u20_n3188 , _u10_u20_n3187 , _u10_u20_n3186 , _u10_u20_n3185 ,_u10_u20_n3184 , _u10_u20_n3183 , _u10_u20_n3182 , _u10_u20_n3181 ,_u10_u20_n3180 , _u10_u20_n3179 , _u10_u20_n3178 , _u10_u20_n3177 ,_u10_u20_n3176 , _u10_u20_n3175 , _u10_u20_n3174 , _u10_u20_n3173 ,_u10_u20_n3172 , _u10_u20_n3171 , _u10_u20_n3170 , _u10_u20_n3169 ,_u10_u20_n3168 , _u10_u20_n3167 , _u10_u20_n3166 , _u10_u20_n3165 ,_u10_u20_n3164 , _u10_u20_n3163 , _u10_u20_n3162 , _u10_u20_n3161 ,_u10_u20_n3160 , _u10_u20_n3159 , _u10_u20_n3158 , _u10_u20_n3157 ,_u10_u20_n3156 , _u10_u20_n3155 , _u10_u20_n3154 , _u10_u20_n3153 ,_u10_u20_n3152 , _u10_u20_n3151 , _u10_u20_n3150 , _u10_u20_n3149 ,_u10_u20_n3148 , _u10_u20_n3147 , _u10_u20_n3146 , _u10_u20_n3145 ,_u10_u20_n3144 , _u10_u20_n3143 , _u10_u20_n3142 , _u10_u20_n3141 ,_u10_u20_n3140 , _u10_u20_n3139 , _u10_u20_n3138 , _u10_u20_n3137 ,_u10_u20_n3136 , _u10_u20_n3135 , _u10_u20_n3134 , _u10_u20_n3133 ,_u10_u20_n3132 , _u10_u20_n3131 , _u10_u20_n3130 , _u10_u20_n3129 ,_u10_u20_n3128 , _u10_u20_n3127 , _u10_u20_n3126 , _u10_u20_n3125 ,_u10_u20_n3124 , _u10_u20_n3123 , _u10_u20_n3122 , _u10_u20_n3121 ,_u10_u20_n3120 , _u10_u20_n3119 , _u10_u20_n3118 , _u10_u20_n3117 ,_u10_u20_n3116 , _u10_u20_n3115 , _u10_u20_n3114 , _u10_u20_n3113 ,_u10_u20_n3112 , _u10_u20_n3111 , _u10_u20_n3110 , _u10_u20_n3109 ,_u10_u20_n3108 , _u10_u20_n3107 , _u10_u20_n3106 , _u10_u20_n3105 ,_u10_u20_n3104 , _u10_u20_n3103 , _u10_u20_n3102 , _u10_u20_n3101 ,_u10_u20_n3100 , _u10_u20_n3099 , _u10_u20_n3098 , _u10_u20_n3097 ,_u10_u20_n3096 , _u10_u20_n3095 , _u10_u20_n3094 , _u10_u20_n3093 ,_u10_u20_n3092 , _u10_u20_n3091 , _u10_u20_n3090 , _u10_u20_n3089 ,_u10_u20_n3088 , _u10_u20_n3087 , _u10_u20_n3086 , _u10_u20_n3085 ,_u10_u20_n3084 , _u10_u20_n3083 , _u10_u20_n3082 , _u10_u20_n3081 ,_u10_u20_n3080 , _u10_u20_n3079 , _u10_u20_n3078 , _u10_u20_n3077 ,_u10_u20_n3076 , _u10_u20_n3075 , _u10_u20_n3074 , _u10_u20_n3073 ,_u10_u20_n3072 , _u10_u20_n3071 , _u10_u20_n3070 , _u10_u20_n3069 ,_u10_u20_n3068 , _u10_u20_n3067 , _u10_u20_n3066 , _u10_u20_n3065 ,_u10_u20_n3064 , _u10_u20_n3063 , _u10_u20_n3062 , _u10_u20_n3061 ,_u10_u20_n3060 , _u10_u20_n3059 , _u10_u20_n3058 , _u10_u20_n3057 ,_u10_u20_n3056 , _u10_u20_n3055 , _u10_u20_n3054 , _u10_u20_n3053 ,_u10_u20_n3052 , _u10_u20_n3051 , _u10_u20_n3050 , _u10_u20_n3049 ,_u10_u20_n3048 , _u10_u20_n3047 , _u10_u20_n3046 , _u10_u20_n3045 ,_u10_u20_n3044 , _u10_u20_n3043 , _u10_u20_n3042 , _u10_u20_n3041 ,_u10_u20_n3040 , _u10_u20_n3039 , _u10_u20_n3038 , _u10_u20_n3037 ,_u10_u20_n3036 , _u10_u20_n3035 , _u10_u20_n3034 , _u10_u20_n3033 ,_u10_u20_n3032 , _u10_u20_n3031 , _u10_u20_n3030 , _u10_u20_n3029 ,_u10_u20_n3028 , _u10_u20_n3027 , _u10_u20_n3026 , _u10_u20_n3025 ,_u10_u20_n3024 , _u10_u20_n3023 , _u10_u20_n3022 , _u10_u20_n3021 ,_u10_u20_n3020 , _u10_u20_n3019 , _u10_u20_n3018 , _u10_u20_n3017 ,_u10_u20_n3016 , _u10_u20_n3015 , _u10_u20_n3014 , _u10_u20_n3013 ,_u10_u20_n3012 , _u10_u20_n3011 , _u10_u20_n3010 , _u10_u20_n3009 ,_u10_u20_n3008 , _u10_u20_n3007 , _u10_u20_n3006 , _u10_u20_n3005 ,_u10_u20_n3004 , _u10_u20_n3003 , _u10_u20_n3002 , _u10_u20_n3001 ,_u10_u20_n3000 , _u10_u20_n2999 , _u10_u20_n2998 , _u10_u20_n2997 ,_u10_u20_n2996 , _u10_u20_n2995 , _u10_u20_n2994 , _u10_u20_n2993 ,_u10_u20_n2992 , _u10_u20_n2991 , _u10_u20_n2990 , _u10_u20_n2989 ,_u10_u20_n2988 , _u10_u20_n2987 , _u10_u20_n2986 , _u10_u20_n2985 ,_u10_u20_n2984 , _u10_u20_n2983 , _u10_u20_n2982 , _u10_u20_n2981 ,_u10_u20_n2980 , _u10_u20_n2979 , _u10_u20_n2978 , _u10_u20_n2977 ,_u10_u20_n2976 , _u10_u20_n2975 , _u10_u20_n2974 , _u10_u20_n2973 ,_u10_u20_n2972 , _u10_u20_n2971 , _u10_u20_n2970 , _u10_u20_n2969 ,_u10_u20_n2968 , _u10_u20_n2967 , _u10_u20_n2966 , _u10_u20_n2965 ,_u10_u20_n2964 , _u10_u20_n2963 , _u10_u20_n2962 , _u10_u20_n2961 ,_u10_u20_n2960 , _u10_u20_n2959 , _u10_u20_n2958 , _u10_u20_n2957 ,_u10_u20_n2956 , _u10_u20_n2955 , _u10_u20_n2954 , _u10_u20_n2953 ,_u10_u20_n2952 , _u10_u20_n2951 , _u10_u20_n2950 , _u10_u20_n2949 ,_u10_u20_n2948 , _u10_u20_n2947 , _u10_u20_n2946 , _u10_u20_n2945 ,_u10_u20_n2944 , _u10_u20_n2943 , _u10_u20_n2942 , _u10_u20_n2941 ,_u10_u20_n2940 , _u10_u20_n2939 , _u10_u20_n2938 , _u10_u20_n2937 ,_u10_u20_n2936 , _u10_u20_n2935 , _u10_u20_n2934 , _u10_u20_n2933 ,_u10_u20_n2932 , _u10_u20_n2931 , _u10_u20_n2930 , _u10_u20_n2929 ,_u10_u20_n2928 , _u10_u20_n2927 , _u10_u20_n2926 , _u10_u20_n2925 ,_u10_u20_n2924 , _u10_u20_n2923 , _u10_u20_n2922 , _u10_u20_n2921 ,_u10_u20_n2920 , _u10_u20_n2919 , _u10_u20_n2918 , _u10_u20_n2917 ,_u10_u20_n2916 , _u10_u20_n2915 , _u10_u20_n2914 , _u10_u20_n2913 ,_u10_u20_n2912 , _u10_u20_n2911 , _u10_u20_n2910 , _u10_u20_n2909 ,_u10_u20_n2908 , _u10_u20_n2907 , _u10_u20_n2906 , _u10_u20_n2905 ,_u10_u20_n2904 , _u10_u20_n2903 , _u10_u20_n2902 , _u10_u20_n2901 ,_u10_u20_n2900 , _u10_u20_n2899 , _u10_u20_n2898 , _u10_u20_n2897 ,_u10_u20_n2896 , _u10_u20_n2895 , _u10_u20_n2894 , _u10_u20_n2893 ,_u10_u20_n2892 , _u10_u20_n2891 , _u10_u20_n2890 , _u10_u20_n2889 ,_u10_u20_n2888 , _u10_u20_n2887 , _u10_u20_n2886 , _u10_u20_n2885 ,_u10_u20_n2884 , _u10_u20_n2883 , _u10_u20_n2882 , _u10_u20_n2881 ,_u10_u20_n2880 , _u10_u20_n2879 , _u10_u20_n2878 , _u10_u20_n2877 ,_u10_u20_n2876 , _u10_u20_n2875 , _u10_u20_n2874 , _u10_u20_n2873 ,_u10_u20_n2872 , _u10_u20_n2871 , _u10_u20_n2870 , _u10_u20_n2869 ,_u10_u20_n2868 , _u10_u20_n2867 , _u10_u20_n2866 , _u10_u20_n2865 ,_u10_u20_n2864 , _u10_u20_n2863 , _u10_u20_n2862 , _u10_u20_n2861 ,_u10_u20_n2860 , _u10_u20_n2859 , _u10_u20_n2858 , _u10_u20_n2857 ,_u10_u20_n2856 , _u10_u20_n2855 , _u10_u20_n2854 , _u10_u20_n2853 ,_u10_u20_n2852 , _u10_u20_n2851 , _u10_u20_n2850 , _u10_u20_n2849 ,_u10_u20_n2848 , _u10_u20_n2847 , _u10_u20_n2846 , _u10_u20_n2845 ,_u10_u20_n2844 , _u10_u20_n2843 , _u10_u20_n2842 , _u10_u20_n2841 ,_u10_u20_n2840 , _u10_u20_n2839 , _u10_u20_n2838 , _u10_u20_n2837 ,_u10_u20_n2836 , _u10_u20_n2835 , _u10_u20_n2834 , _u10_u20_n2833 ,_u10_u20_n2832 , _u10_u20_n2831 , _u10_u20_n2830 , _u10_u20_n2829 ,_u10_u20_n2828 , _u10_u20_n2827 , _u10_u20_n2826 , _u10_u20_n2825 ,_u10_u20_n2824 , _u10_u20_n2823 , _u10_u20_n2822 , _u10_u20_n2821 ,_u10_u20_n2820 , _u10_u20_n2819 , _u10_u20_n2818 , _u10_u20_n2817 ,_u10_u20_n2816 , _u10_u20_n2815 , _u10_u20_n2814 , _u10_u20_n2813 ,_u10_u20_n2812 , _u10_u20_n2811 , _u10_u20_n2810 , _u10_u20_n2809 ,_u10_u20_n2808 , _u10_u20_n2807 , _u10_u20_n2806 , _u10_u20_n2805 ,_u10_u20_n2804 , _u10_u20_n2803 , _u10_u20_n2802 , _u10_u20_n2801 ,_u10_u20_n2800 , _u10_u20_n2799 , _u10_u20_n2798 , _u10_u20_n2797 ,_u10_u20_n2796 , _u10_u20_n2795 , _u10_u20_n2794 , _u10_u20_n2793 ,_u10_u20_n2792 , _u10_u20_n2791 , _u10_u20_n2790 , _u10_u20_n2789 ,_u10_u20_n2788 , _u10_u20_n2787 , _u10_u20_n2786 , _u10_u20_n2785 ,_u10_u20_n2784 , _u10_u20_n2783 , _u10_u20_n2782 , _u10_u20_n2781 ,_u10_u20_n2780 , _u10_u20_n2779 , _u10_u20_n2778 , _u10_u20_n2777 ,_u10_u20_n2776 , _u10_u20_n2775 , _u10_u20_n2774 , _u10_u20_n2773 ,_u10_u20_n2772 , _u10_u20_n2771 , _u10_u20_n2770 , _u10_u20_n2769 ,_u10_u20_n2768 , _u10_u20_n2767 , _u10_u20_n2766 , _u10_u20_n2765 ,_u10_u20_n2764 , _u10_u20_n2763 , _u10_u20_n2762 , _u10_u20_n2761 ,_u10_u20_n2760 , _u10_u20_n2759 , _u10_u20_n2758 , _u10_u20_n2757 ,_u10_u20_n2756 , _u10_u20_n2755 , _u10_u20_n2754 , _u10_u20_n2753 ,_u10_u20_n2752 , _u10_u20_n2751 , _u10_u20_n2750 , _u10_u20_n2749 ,_u10_u20_n2748 , _u10_u20_n2747 , _u10_u20_n2746 , _u10_u20_n2745 ,_u10_u20_n2744 , _u10_u20_n2743 , _u10_u20_n2742 , _u10_u20_n2741 ,_u10_u20_n2740 , _u10_u20_n2739 , _u10_u20_n2738 , _u10_u20_n2737 ,_u10_u20_n2736 , _u10_u20_n2735 , _u10_u20_n2734 , _u10_u20_n2733 ,_u10_u20_n2732 , _u10_u20_n2731 , _u10_u20_n2730 , _u10_u20_n2729 ,_u10_u20_n2728 , _u10_u20_n2727 , _u10_u20_n2726 , _u10_u20_n2725 ,_u10_u20_n2724 , _u10_u20_n2723 , _u10_u20_n2722 , _u10_u20_n2721 ,_u10_u20_n2720 , _u10_u20_n2719 , _u10_u20_n2718 , _u10_u20_n2717 ,_u10_u20_n2716 , _u10_u20_n2715 , _u10_u20_n2714 , _u10_u20_n2713 ,_u10_u20_n2712 , _u10_u20_n2711 , _u10_u20_n2710 , _u10_u20_n2709 ,_u10_u20_n2708 , _u10_u20_n2707 , _u10_u20_n2706 , _u10_u20_n2705 ,_u10_u20_n2704 , _u10_u20_n2703 , _u10_u20_n2702 , _u10_u20_n2701 ,_u10_u20_n2700 , _u10_u20_n2699 , _u10_u20_n2698 , _u10_u20_n2697 ,_u10_u20_n2696 , _u10_u20_n2695 , _u10_u20_n2694 , _u10_u20_n2693 ,_u10_u20_n2692 , _u10_u20_n2691 , _u10_u20_n2690 , _u10_u20_n2689 ,_u10_u20_n2688 , _u10_u20_n2687 , _u10_u20_n2686 , _u10_u20_n2685 ,_u10_u20_n2684 , _u10_u20_n2683 , _u10_u20_n2682 , _u10_u20_n2681 ,_u10_u20_n2680 , _u10_u20_n2679 , _u10_u20_n2678 , _u10_u20_n2677 ,_u10_u20_n2676 , _u10_u20_n2675 , _u10_u20_n2674 , _u10_u20_n2673 ,_u10_u20_n2672 , _u10_u20_n2671 , _u10_u20_n2670 , _u10_u20_n2669 ,_u10_u20_n2668 , _u10_u20_n2667 , _u10_u20_n2666 , _u10_u20_n2665 ,_u10_u20_n2664 , _u10_u20_n2663 , _u10_u20_n2662 , _u10_u20_n2661 ,_u10_u20_n2660 , _u10_u20_n2659 , _u10_u20_n2658 , _u10_u20_n2657 ,_u10_u20_n2656 , _u10_u20_n2655 , _u10_u20_n2654 , _u10_u20_n2653 ,_u10_u20_n2652 , _u10_u20_n2651 , _u10_u20_n2650 , _u10_u20_n2649 ,_u10_u20_n2648 , _u10_u20_n2647 , _u10_u20_n2646 , _u10_u20_n2645 ,_u10_u20_n2644 , _u10_u20_n2643 , _u10_u20_n2642 , _u10_u20_n2641 ,_u10_u20_n2640 , _u10_u20_n2639 , _u10_u20_n2638 , _u10_u20_n2637 ,_u10_u20_n2636 , _u10_u20_n2635 , _u10_u20_n2634 , _u10_u20_n2633 ,_u10_u20_n2632 , _u10_u20_n2631 , _u10_u20_n2630 , _u10_u20_n2629 ,_u10_u20_n2628 , _u10_u20_n2627 , _u10_u20_n2626 , _u10_u20_n2625 ,_u10_u20_n2624 , _u10_u20_n2623 , _u10_u20_n2622 , _u10_u20_n2621 ,_u10_u20_n2620 , _u10_u20_n2619 , _u10_u20_n2618 , _u10_u20_n2617 ,_u10_u20_n2616 , _u10_u20_n2615 , _u10_u20_n2614 , _u10_u20_n2613 ,_u10_u20_n2612 , _u10_u20_n2611 , _u10_u20_n2610 , _u10_u20_n2609 ,_u10_u20_n2608 , _u10_u20_n2607 , _u10_u20_n2606 , _u10_u20_n2605 ,_u10_u20_n2604 , _u10_u20_n2603 , _u10_u20_n2602 , _u10_u20_n2601 ,_u10_u20_n2600 , _u10_u20_n2599 , _u10_u20_n2598 , _u10_u20_n2597 ,_u10_u20_n2596 , _u10_u20_n2595 , _u10_u20_n2594 , _u10_u20_n2593 ,_u10_u20_n2592 , _u10_u20_n2591 , _u10_u20_n2590 , _u10_u20_n2589 ,_u10_u20_n2588 , _u10_u20_n2587 , _u10_u20_n2586 , _u10_u20_n2585 ,_u10_u20_n2584 , _u10_u20_n2583 , _u10_u20_n2582 , _u10_u20_n2581 ,_u10_u20_n2580 , _u10_u20_n2579 , _u10_u20_n2578 , _u10_u20_n2577 ,_u10_u20_n2576 , _u10_u20_n2575 , _u10_u20_n2574 , _u10_u20_n2573 ,_u10_u20_n2572 , _u10_u20_n2571 , _u10_u20_n2570 , _u10_u20_n2569 ,_u10_u20_n2568 , _u10_u20_n2567 , _u10_u20_n2566 , _u10_u20_n2565 ,_u10_u20_n2564 , _u10_u20_n2563 , _u10_u20_n2562 , _u10_u20_n2561 ,_u10_u20_n2560 , _u10_u20_n2559 , _u10_u20_n2558 , _u10_u20_n2557 ,_u10_u20_n2556 , _u10_u20_n2555 , _u10_u20_n2554 , _u10_u20_n2553 ,_u10_u20_n2552 , _u10_u20_n2551 , _u10_u20_n2550 , _u10_u20_n2549 ,_u10_u20_n2548 , _u10_u20_n2547 , _u10_u20_n2546 , _u10_u20_n2545 ,_u10_u20_n2544 , _u10_u20_n2543 , _u10_u20_n2542 , _u10_u20_n2541 ,_u10_u20_n2540 , _u10_u20_n2539 , _u10_u20_n2538 , _u10_u20_n2537 ,_u10_u20_n2536 , _u10_u20_n2535 , _u10_u20_n2534 , _u10_u20_n2533 ,_u10_u20_n2532 , _u10_u20_n2531 , _u10_u20_n2530 , _u10_u20_n2529 ,_u10_u20_n2528 , _u10_u20_n2527 , _u10_u20_n2526 , _u10_u20_n2525 ,_u10_u20_n2524 , _u10_u20_n2523 , _u10_u20_n2522 , _u10_u20_n2521 ,_u10_u20_n2520 , _u10_u20_n2519 , _u10_u20_n2518 , _u10_u20_n2517 ,_u10_u20_n2516 , _u10_u20_n2515 , _u10_u20_n2514 , _u10_u20_n2513 ,_u10_u20_n2512 , _u10_u20_n2511 , _u10_u20_n2510 , _u10_u20_n2509 ,_u10_u20_n2508 , _u10_u20_n2507 , _u10_u20_n2506 , _u10_u20_n2505 ,_u10_u20_n2504 , _u10_u20_n2503 , _u10_u20_n2502 , _u10_u20_n2501 ,_u10_u20_n2500 , _u10_u20_n2499 , _u10_u20_n2498 , _u10_u20_n2497 ,_u10_u20_n2496 , _u10_u20_n2495 , _u10_u20_n2494 , _u10_u20_n2493 ,_u10_u20_n2492 , _u10_u20_n2491 , _u10_u20_n2490 , _u10_u20_n2489 ,_u10_u20_n2488 , _u10_u20_n2487 , _u10_u20_n2486 , _u10_u20_n2485 ,_u10_u20_n2484 , _u10_u20_n2483 , _u10_u20_n2482 , _u10_u20_n2481 ,_u10_u20_n2480 , _u10_u20_n2479 , _u10_u20_n2478 , _u10_u20_n2477 ,_u10_u20_n2476 , _u10_u20_n2475 , _u10_u20_n2474 , _u10_u20_n2473 ,_u10_u20_n2472 , _u10_u20_n2471 , _u10_u20_n2470 , _u10_u20_n2469 ,_u10_u20_n2468 , _u10_u20_n2467 , _u10_u20_n2466 , _u10_u20_n2465 ,_u10_u20_n2464 , _u10_u20_n2463 , _u10_u20_n2462 , _u10_u20_n2461 ,_u10_u20_n2460 , _u10_u20_n2459 , _u10_u20_n2458 , _u10_u20_n2457 ,_u10_u20_n2456 , _u10_u20_n2455 , _u10_u20_n2454 , _u10_u20_n2453 ,_u10_u20_n2452 , _u10_u20_n2451 , _u10_u20_n2450 , _u10_u20_n2449 ,_u10_u20_n2448 , _u10_u20_n2447 , _u10_u20_n2446 , _u10_u20_n2445 ,_u10_u20_n2444 , _u10_u20_n2443 , _u10_u20_n2442 , _u10_u20_n2441 ,_u10_u20_n2440 , _u10_u20_n2439 , _u10_u20_n2438 , _u10_u20_n2437 ,_u10_u20_n2436 , _u10_u20_n2435 , _u10_u20_n2434 , _u10_u20_n2433 ,_u10_u20_n2432 , _u10_u20_n2431 , _u10_u20_n2430 , _u10_u20_n2429 ,_u10_u20_n2428 , _u10_u20_n2427 , _u10_u20_n2426 , _u10_u20_n2425 ,_u10_u20_n2424 , _u10_u20_n2423 , _u10_u20_n2422 , _u10_u20_n2421 ,_u10_u20_n2420 , _u10_u20_n2419 , _u10_u20_n2418 , _u10_u20_n2417 ,_u10_u20_n2416 , _u10_u20_n2415 , _u10_u20_n2414 , _u10_u20_n2413 ,_u10_u20_n2412 , _u10_u20_n2411 , _u10_u20_n2410 , _u10_u20_n2409 ,_u10_u20_n2408 , _u10_u20_n2407 , _u10_u20_n2406 , _u10_u20_n2405 ,_u10_u20_n2404 , _u10_u20_n2403 , _u10_u20_n2402 , _u10_u20_n2401 ,_u10_u20_n2400 , _u10_u20_n2399 , _u10_u20_n2398 , _u10_u20_n2397 ,_u10_u20_n2396 , _u10_u20_n2395 , _u10_u20_n2394 , _u10_u20_n2393 ,_u10_u20_n2392 , _u10_u20_n2391 , _u10_u20_n2390 , _u10_u20_n2389 ,_u10_u20_n2388 , _u10_u20_n2387 , _u10_u20_n2386 , _u10_u20_n2385 ,_u10_u20_n2384 , _u10_u20_n2383 , _u10_u20_n2382 , _u10_u20_n2381 ,_u10_u20_n2380 , _u10_u20_n2379 , _u10_u20_n2378 , _u10_u20_n2377 ,_u10_u20_n2376 , _u10_u20_n2375 , _u10_u20_n2374 , _u10_u20_n2373 ,_u10_u20_n2372 , _u10_u20_n2371 , _u10_u20_n2370 , _u10_u20_n2369 ,_u10_u20_n2368 , _u10_u20_n2367 , _u10_u20_n2366 , _u10_u20_n2365 ,_u10_u20_n2364 , _u10_u20_n2363 , _u10_u20_n2362 , _u10_u20_n2361 ,_u10_u20_n2360 , _u10_u20_n2359 , _u10_u20_n2358 , _u10_u20_n2357 ,_u10_u20_n2356 , _u10_u20_n2355 , _u10_u20_n2354 , _u10_u20_n2353 ,_u10_u20_n2352 , _u10_u20_n2351 , _u10_u20_n2350 , _u10_u20_n2349 ,_u10_u20_n2348 , _u10_u20_n2347 , _u10_u20_n2346 , _u10_u20_n2345 ,_u10_u20_n2344 , _u10_u20_n2343 , _u10_u20_n2342 , _u10_u20_n2341 ,_u10_u20_n2340 , _u10_u20_n2339 , _u10_u20_n2338 , _u10_u20_n2337 ,_u10_u20_n2336 , _u10_u20_n2335 , _u10_u20_n2334 , _u10_u20_n2333 ,_u10_u20_n2332 , _u10_u20_n2331 , _u10_u20_n2330 , _u10_u20_n2329 ,_u10_u20_n2328 , _u10_u20_n2327 , _u10_u20_n2326 , _u10_u20_n2325 ,_u10_u20_n2324 , _u10_u20_n2323 , _u10_u20_n2322 , _u10_u20_n2321 ,_u10_u20_n2320 , _u10_u20_n2319 , _u10_u20_n2318 , _u10_u20_n2317 ,_u10_u20_n2316 , _u10_u20_n2315 , _u10_u20_n2314 , _u10_u20_n2313 ,_u10_u20_n2312 , _u10_u20_n2311 , _u10_u20_n2310 , _u10_u20_n2309 ,_u10_u20_n2308 , _u10_u20_n2307 , _u10_u20_n2306 , _u10_u20_n2305 ,_u10_u20_n2304 , _u10_u20_n2303 , _u10_u20_n2302 , _u10_u20_n2301 ,_u10_u20_n2300 , _u10_u20_n2299 , _u10_u20_n2298 , _u10_u20_n2297 ,_u10_u20_n2296 , _u10_u20_n2295 , _u10_u20_n2294 , _u10_u20_n2293 ,_u10_u20_n2292 , _u10_u20_n2291 , _u10_u20_n2290 , _u10_u20_n2289 ,_u10_u20_n2288 , _u10_u20_n2287 , _u10_u20_n2286 , _u10_u20_n2285 ,_u10_u20_n2284 , _u10_u20_n2283 , _u10_u20_n2282 , _u10_u20_n2281 ,_u10_u20_n2280 , _u10_u20_n2279 , _u10_u20_n2278 , _u10_u20_n2277 ,_u10_u20_n2276 , _u10_u20_n2275 , _u10_u20_n2274 , _u10_u20_n2273 ,_u10_u20_n2272 , _u10_u20_n2271 , _u10_u20_n2270 , _u10_u20_n2269 ,_u10_u20_n2268 , _u10_u20_n2267 , _u10_u20_n2266 , _u10_u20_n2265 ,_u10_u20_n2264 , _u10_u20_n2263 , _u10_u20_n2262 , _u10_u20_n2261 ,_u10_u20_n2260 , _u10_u20_n2259 , _u10_u20_n2258 , _u10_u20_n2257 ,_u10_u20_n2256 , _u10_u20_n2255 , _u10_u20_n2254 , _u10_u20_n2253 ,_u10_u20_n2252 , _u10_u20_n2251 , _u10_u20_n2250 , _u10_u20_n2249 ,_u10_u20_n2248 , _u10_u20_n2247 , _u10_u20_n2246 , _u10_u20_n2245 ,_u10_u20_n2244 , _u10_u20_n2243 , _u10_u20_n2242 , _u10_u20_n2241 ,_u10_u20_n2240 , _u10_u20_n2239 , _u10_u20_n2238 , _u10_u20_n2237 ,_u10_u20_n2236 , _u10_u20_n2235 , _u10_u20_n2234 , _u10_u20_n2233 ,_u10_u20_n2232 , _u10_u20_n2231 , _u10_u20_n2230 , _u10_u20_n2229 ,_u10_u20_n2228 , _u10_u20_n2227 , _u10_u20_n2226 , _u10_u20_n2225 ,_u10_u20_n2224 , _u10_u20_n2223 , _u10_u20_n2222 , _u10_u20_n2221 ,_u10_u20_n2220 , _u10_u20_n2219 , _u10_u20_n2218 , _u10_u20_n2217 ,_u10_u20_n2216 , _u10_u20_n2215 , _u10_u20_n2214 , _u10_u20_n2213 ,_u10_u20_n2212 , _u10_u20_n2211 , _u10_u20_n2210 , _u10_u20_n2209 ,_u10_u20_n2208 , _u10_u20_n2207 , _u10_u20_n2206 , _u10_u20_n2205 ,_u10_u20_n2204 , _u10_u20_n2203 , _u10_u20_n2202 , _u10_u20_n2201 ,_u10_u20_n2200 , _u10_u20_n2199 , _u10_u20_n2198 , _u10_u20_n2197 ,_u10_u20_n2196 , _u10_u20_n2195 , _u10_u20_n2194 , _u10_u20_n2193 ,_u10_u20_n2192 , _u10_u20_n2191 , _u10_u20_n2190 , _u10_u20_n2189 ,_u10_u20_n2188 , _u10_u20_n2187 , _u10_u20_n2186 , _u10_u20_n2185 ,_u10_u20_n2184 , _u10_u20_n2183 , _u10_u20_n2182 , _u10_u20_n2181 ,_u10_u20_n2180 , _u10_u20_n2179 , _u10_u20_n2178 , _u10_u20_n2177 ,_u10_u20_n2176 , _u10_u20_n2175 , _u10_u20_n2174 , _u10_u20_n2173 ,_u10_u20_n2172 , _u10_u20_n2171 , _u10_u20_n2170 , _u10_u20_n2169 ,_u10_u20_n2168 , _u10_u20_n2167 , _u10_u20_n2166 , _u10_u20_n2165 ,_u10_u20_n2164 , _u10_u20_n2163 , _u10_u20_n2162 , _u10_u20_n2161 ,_u10_u20_n2160 , _u10_u20_n2159 , _u10_u20_n2158 , _u10_u20_n2157 ,_u10_u20_n2156 , _u10_u20_n2155 , _u10_u20_n2154 , _u10_u20_n2153 ,_u10_u20_n2152 , _u10_u20_n2151 , _u10_u20_n2150 , _u10_u20_n2149 ,_u10_u20_n2148 , _u10_u20_n2147 , _u10_u20_n2146 , _u10_u20_n2145 ,_u10_u20_n2144 , _u10_u20_n2143 , _u10_u20_n2142 , _u10_u20_n2141 ,_u10_u20_n2140 , _u10_u20_n2139 , _u10_u20_n2138 , _u10_u20_n2137 ,_u10_u20_n2136 , _u10_u20_n2135 , _u10_u20_n2134 , _u10_u20_n2133 ,_u10_u20_n2132 , _u10_u20_n2131 , _u10_u20_n2130 , _u10_u20_n2129 ,_u10_u20_n2128 , _u10_u20_n2127 , _u10_u20_n2126 , _u10_u20_n2125 ,_u10_u20_n2124 , _u10_u20_n2123 , _u10_u20_n2122 , _u10_u20_n2121 ,_u10_u20_n2120 , _u10_u20_n2119 , _u10_u20_n2118 , _u10_u20_n2117 ,_u10_u20_n2116 , _u10_u20_n2115 , _u10_u20_n2114 , _u10_u20_n2113 ,_u10_u20_n2112 , _u10_u20_n2111 , _u10_u20_n2110 , _u10_u20_n2109 ,_u10_u20_n2108 , _u10_u20_n2107 , _u10_u20_n2106 , _u10_u20_n2105 ,_u10_u20_n2104 , _u10_u20_n2103 , _u10_u20_n2102 , _u10_u20_n2101 ,_u10_u20_n2100 , _u10_u20_n2099 , _u10_u20_n2098 , _u10_u20_n2097 ,_u10_u20_n2096 , _u10_u20_n2095 , _u10_u20_n2094 , _u10_u20_n2093 ,_u10_u20_n2092 , _u10_u20_n2091 , _u10_u20_n2090 , _u10_u20_n2089 ,_u10_u20_n2088 , _u10_u20_n2087 , _u10_u20_n2086 , _u10_u20_n2085 ,_u10_u20_n2084 , _u10_u20_n2083 , _u10_u20_n2082 , _u10_u20_n2081 ,_u10_u20_n2080 , _u10_u20_n2079 , _u10_u20_n2078 , _u10_u20_n2077 ,_u10_u20_n2076 , _u10_u20_n2075 , _u10_u20_n2074 , _u10_u20_n2073 ,_u10_u20_n2072 , _u10_u20_n2071 , _u10_u20_n2070 , _u10_u20_n2069 ,_u10_u20_n2068 , _u10_u20_n2067 , _u10_u20_n2066 , _u10_u20_n2065 ,_u10_u20_n2064 , _u10_u20_n2063 , _u10_u20_n2062 , _u10_u20_n2061 ,_u10_u20_n2060 , _u10_u20_n2059 , _u10_u20_n2058 , _u10_u20_n2057 ,_u10_u20_n2056 , _u10_u20_n2055 , _u10_u20_n2054 , _u10_u20_n2053 ,_u10_u20_n2052 , _u10_u20_n2051 , _u10_u20_n2050 , _u10_u20_n2049 ,_u10_u20_n2048 , _u10_u20_n2047 , _u10_u20_n2046 , _u10_u20_n2045 ,_u10_u20_n2044 , _u10_u20_n2043 , _u10_u20_n2042 , _u10_u20_n2041 ,_u10_u20_n2040 , _u10_u20_n2039 , _u10_u20_n2038 , _u10_u20_n2037 ,_u10_u20_n2036 , _u10_u20_n2035 , _u10_u20_n2034 , _u10_u20_n2033 ,_u10_u20_n2032 , _u10_u20_n2031 , _u10_u20_n2030 , _u10_u20_n2029 ,_u10_u20_n2028 , _u10_u20_n2027 , _u10_u20_n2026 , _u10_u20_n2025 ,_u10_u20_n2024 , _u10_u20_n2023 , _u10_u20_n2022 , _u10_u20_n2021 ,_u10_u20_n2020 , _u10_u20_n2019 , _u10_u20_n2018 , _u10_u20_n2017 ,_u10_u20_n2016 , _u10_u20_n2015 , _u10_u20_n2014 , _u10_u20_n2013 ,_u10_u20_n2012 , _u10_u20_n2011 , _u10_u20_n2010 , _u10_u20_n2009 ,_u10_u20_n2008 , _u10_u20_n2007 , _u10_u20_n2006 , _u10_u20_n2005 ,_u10_u20_n2004 , _u10_u20_n2003 , _u10_u20_n2002 , _u10_u20_n2001 ,_u10_u20_n2000 , _u10_u20_n1999 , _u10_u20_n1998 , _u10_u20_n1997 ,_u10_u20_n1996 , _u10_u20_n1995 , _u10_u20_n1994 , _u10_u20_n1993 ,_u10_u20_n1992 , _u10_u20_n1991 , _u10_u20_n1990 , _u10_u20_n1989 ,_u10_u20_n1988 , _u10_u20_n1987 , _u10_u20_n1986 , _u10_u20_n1985 ,_u10_u20_n1984 , _u10_u20_n1983 , _u10_u20_n1982 , _u10_u20_n1981 ,_u10_u20_n1980 , _u10_u20_n1979 , _u10_u20_n1978 , _u10_u20_n1977 ,_u10_u20_n1976 , _u10_u20_n1975 , _u10_u20_n1974 , _u10_u20_n1973 ,_u10_u20_n1972 , _u10_u20_n1971 , _u10_u20_n1970 , _u10_u20_n1969 ,_u10_u20_n1968 , _u10_u20_n1967 , _u10_u20_n1966 , _u10_u20_n1965 ,_u10_u20_n1964 , _u10_u20_n1963 , _u10_u20_n1962 , _u10_u20_n1961 ,_u10_u20_n1960 , _u10_u20_n1959 , _u10_u20_n1958 , _u10_u20_n1957 ,_u10_u20_n1956 , _u10_u20_n1955 , _u10_u20_n1954 , _u10_u20_n1953 ,_u10_u20_n1952 , _u10_u20_n1951 , _u10_u20_n1950 , _u10_u20_n1949 ,_u10_u20_n1948 , _u10_u20_n1947 , _u10_u20_n1946 , _u10_u20_n1945 ,_u10_u20_n1944 , _u10_u20_n1943 , _u10_u20_n1942 , _u10_u20_n1941 ,_u10_u20_n1940 , _u10_u20_n1939 , _u10_u20_n1938 , _u10_u20_n1937 ,_u10_u20_n1936 , _u10_u20_n1935 , _u10_u20_n1934 , _u10_u20_n1933 ,_u10_u20_n1932 , _u10_u20_n1931 , _u10_u20_n1930 , _u10_u20_n1929 ,_u10_u20_n1928 , _u10_u20_n1927 , _u10_u20_n1926 , _u10_u20_n1925 ,_u10_u20_n1924 , _u10_u20_n1923 , _u10_u20_n1922 , _u10_u20_n1921 ,_u10_u20_n1920 , _u10_u20_n1919 , _u10_u20_n1918 , _u10_u20_n1917 ,_u10_u20_n1916 , _u10_u20_n1915 , _u10_u20_n1914 , _u10_u20_n1913 ,_u10_u20_n1912 , _u10_u20_n1911 , _u10_u20_n1910 , _u10_u20_n1909 ,_u10_u20_n1908 , _u10_u20_n1907 , _u10_u20_n1906 , _u10_u20_n1905 ,_u10_u20_n1904 , _u10_u20_n1903 , _u10_u20_n1902 , _u10_u20_n1901 ,_u10_u20_n1900 , _u10_u20_n1899 , _u10_u20_n1898 , _u10_u20_n1897 ,_u10_u20_n1896 , _u10_u20_n1895 , _u10_u20_n1894 , _u10_u20_n1893 ,_u10_u20_n1892 , _u10_u20_n1891 , _u10_u20_n1890 , _u10_u20_n1889 ,_u10_u20_n1888 , _u10_u20_n1887 , _u10_u20_n1886 , _u10_u20_n1885 ,_u10_u20_n1884 , _u10_u20_n1883 , _u10_u20_n1882 , _u10_u20_n1881 ,_u10_u20_n1880 , _u10_u20_n1879 , _u10_u20_n1878 , _u10_u20_n1877 ,_u10_u20_n1876 , _u10_u20_n1875 , _u10_u20_n1874 , _u10_u20_n1873 ,_u10_u20_n1872 , _u10_u20_n1871 , _u10_u20_n1870 , _u10_u20_n1869 ,_u10_u20_n1868 , _u10_u20_n1867 , _u10_u20_n1866 , _u10_u20_n1865 ,_u10_u20_n1864 , _u10_u20_n1863 , _u10_u20_n1862 , _u10_u20_n1861 ,_u10_u20_n1860 , _u10_u20_n1859 , _u10_u20_n1858 , _u10_u20_n1857 ,_u10_u20_n1856 , _u10_u20_n1855 , _u10_u20_n1854 , _u10_u20_n1853 ,_u10_u20_n1852 , _u10_u20_n1851 , _u10_u20_n1850 , _u10_u20_n1849 ,_u10_u20_n1848 , _u10_u20_n1847 , _u10_u20_n1846 , _u10_u20_n1845 ,_u10_u20_n1844 , _u10_u20_n1843 , _u10_u20_n1842 , _u10_u20_n1841 ,_u10_u20_n1840 , _u10_u20_n1839 , _u10_u20_n1838 , _u10_u20_n1837 ,_u10_u20_n1836 , _u10_u20_n1835 , _u10_u20_n1834 , _u10_u20_n1833 ,_u10_u20_n1832 , _u10_u20_n1831 , _u10_u20_n1830 , _u10_u20_n1829 ,_u10_u20_n1828 , _u10_u20_n1827 , _u10_u20_n1826 , _u10_u20_n1825 ,_u10_u20_n1824 , _u10_u20_n1823 , _u10_u20_n1822 , _u10_u20_n1821 ,_u10_u20_n1820 , _u10_u20_n1819 , _u10_u20_n1818 , _u10_u20_n1817 ,_u10_u20_n1816 , _u10_u20_n1815 , _u10_u20_n1814 , _u10_u20_n1813 ,_u10_u20_n1812 , _u10_u20_n1811 , _u10_u20_n1810 , _u10_u20_n1809 ,_u10_u20_n1808 , _u10_u3_n3416 , _u10_u3_n3415 , _u10_u3_n3414 ,_u10_u3_n3413 , _u10_u3_n3412 , _u10_u3_n3411 , _u10_u3_n3410 ,_u10_u3_n3409 , _u10_u3_n3408 , _u10_u3_n3407 , _u10_u3_n3406 ,_u10_u3_n3405 , _u10_u3_n3404 , _u10_u3_n3403 , _u10_u3_n3402 ,_u10_u3_n3401 , _u10_u3_n3400 , _u10_u3_n3399 , _u10_u3_n3398 ,_u10_u3_n3397 , _u10_u3_n3396 , _u10_u3_n3395 , _u10_u3_n3394 ,_u10_u3_n3393 , _u10_u3_n3392 , _u10_u3_n3391 , _u10_u3_n3390 ,_u10_u3_n3389 , _u10_u3_n3388 , _u10_u3_n3387 , _u10_u3_n3386 ,_u10_u3_n3385 , _u10_u3_n3384 , _u10_u3_n3383 , _u10_u3_n3382 ,_u10_u3_n3381 , _u10_u3_n3380 , _u10_u3_n3379 , _u10_u3_n3378 ,_u10_u3_n3377 , _u10_u3_n3376 , _u10_u3_n3375 , _u10_u3_n3374 ,_u10_u3_n3373 , _u10_u3_n3372 , _u10_u3_n3371 , _u10_u3_n3370 ,_u10_u3_n3369 , _u10_u3_n3368 , _u10_u3_n3367 , _u10_u3_n3366 ,_u10_u3_n3365 , _u10_u3_n3364 , _u10_u3_n3363 , _u10_u3_n3362 ,_u10_u3_n3361 , _u10_u3_n3360 , _u10_u3_n3359 , _u10_u3_n3358 ,_u10_u3_n3357 , _u10_u3_n3356 , _u10_u3_n3355 , _u10_u3_n3354 ,_u10_u3_n3353 , _u10_u3_n3352 , _u10_u3_n3351 , _u10_u3_n3350 ,_u10_u3_n3349 , _u10_u3_n3348 , _u10_u3_n3347 , _u10_u3_n3346 ,_u10_u3_n3345 , _u10_u3_n3344 , _u10_u3_n3343 , _u10_u3_n3342 ,_u10_u3_n3341 , _u10_u3_n3340 , _u10_u3_n3339 , _u10_u3_n3338 ,_u10_u3_n3337 , _u10_u3_n3336 , _u10_u3_n3335 , _u10_u3_n3334 ,_u10_u3_n3333 , _u10_u3_n3332 , _u10_u3_n3331 , _u10_u3_n3330 ,_u10_u3_n3329 , _u10_u3_n3328 , _u10_u3_n3327 , _u10_u3_n3326 ,_u10_u3_n3325 , _u10_u3_n3324 , _u10_u3_n3323 , _u10_u3_n3322 ,_u10_u3_n3321 , _u10_u3_n3320 , _u10_u3_n3319 , _u10_u3_n3318 ,_u10_u3_n3317 , _u10_u3_n3316 , _u10_u3_n3315 , _u10_u3_n3314 ,_u10_u3_n3313 , _u10_u3_n3312 , _u10_u3_n3311 , _u10_u3_n3310 ,_u10_u3_n3309 , _u10_u3_n3308 , _u10_u3_n3307 , _u10_u3_n3306 ,_u10_u3_n3305 , _u10_u3_n3304 , _u10_u3_n3303 , _u10_u3_n3302 ,_u10_u3_n3301 , _u10_u3_n3300 , _u10_u3_n3299 , _u10_u3_n3298 ,_u10_u3_n3297 , _u10_u3_n3296 , _u10_u3_n3295 , _u10_u3_n3294 ,_u10_u3_n3293 , _u10_u3_n3292 , _u10_u3_n3291 , _u10_u3_n3290 ,_u10_u3_n3289 , _u10_u3_n3288 , _u10_u3_n3287 , _u10_u3_n3286 ,_u10_u3_n3285 , _u10_u3_n3284 , _u10_u3_n3283 , _u10_u3_n3282 ,_u10_u3_n3281 , _u10_u3_n3280 , _u10_u3_n3279 , _u10_u3_n3278 ,_u10_u3_n3277 , _u10_u3_n3276 , _u10_u3_n3275 , _u10_u3_n3274 ,_u10_u3_n3273 , _u10_u3_n3272 , _u10_u3_n3271 , _u10_u3_n3270 ,_u10_u3_n3269 , _u10_u3_n3268 , _u10_u3_n3267 , _u10_u3_n3266 ,_u10_u3_n3265 , _u10_u3_n3264 , _u10_u3_n3263 , _u10_u3_n3262 ,_u10_u3_n3261 , _u10_u3_n3260 , _u10_u3_n3259 , _u10_u3_n3258 ,_u10_u3_n3257 , _u10_u3_n3256 , _u10_u3_n3255 , _u10_u3_n3254 ,_u10_u3_n3253 , _u10_u3_n3252 , _u10_u3_n3251 , _u10_u3_n3250 ,_u10_u3_n3249 , _u10_u3_n3248 , _u10_u3_n3247 , _u10_u3_n3246 ,_u10_u3_n3245 , _u10_u3_n3244 , _u10_u3_n3243 , _u10_u3_n3242 ,_u10_u3_n3241 , _u10_u3_n3240 , _u10_u3_n3239 , _u10_u3_n3238 ,_u10_u3_n3237 , _u10_u3_n3236 , _u10_u3_n3235 , _u10_u3_n3234 ,_u10_u3_n3233 , _u10_u3_n3232 , _u10_u3_n3231 , _u10_u3_n3230 ,_u10_u3_n3229 , _u10_u3_n3228 , _u10_u3_n3227 , _u10_u3_n3226 ,_u10_u3_n3225 , _u10_u3_n3224 , _u10_u3_n3223 , _u10_u3_n3222 ,_u10_u3_n3221 , _u10_u3_n3220 , _u10_u3_n3219 , _u10_u3_n3218 ,_u10_u3_n3217 , _u10_u3_n3216 , _u10_u3_n3215 , _u10_u3_n3214 ,_u10_u3_n3213 , _u10_u3_n3212 , _u10_u3_n3211 , _u10_u3_n3210 ,_u10_u3_n3209 , _u10_u3_n3208 , _u10_u3_n3207 , _u10_u3_n3206 ,_u10_u3_n3205 , _u10_u3_n3204 , _u10_u3_n3203 , _u10_u3_n3202 ,_u10_u3_n3201 , _u10_u3_n3200 , _u10_u3_n3199 , _u10_u3_n3198 ,_u10_u3_n3197 , _u10_u3_n3196 , _u10_u3_n3195 , _u10_u3_n3194 ,_u10_u3_n3193 , _u10_u3_n3192 , _u10_u3_n3191 , _u10_u3_n3190 ,_u10_u3_n3189 , _u10_u3_n3188 , _u10_u3_n3187 , _u10_u3_n3186 ,_u10_u3_n3185 , _u10_u3_n3184 , _u10_u3_n3183 , _u10_u3_n3182 ,_u10_u3_n3181 , _u10_u3_n3180 , _u10_u3_n3179 , _u10_u3_n3178 ,_u10_u3_n3177 , _u10_u3_n3176 , _u10_u3_n3175 , _u10_u3_n3174 ,_u10_u3_n3173 , _u10_u3_n3172 , _u10_u3_n3171 , _u10_u3_n3170 ,_u10_u3_n3169 , _u10_u3_n3168 , _u10_u3_n3167 , _u10_u3_n3166 ,_u10_u3_n3165 , _u10_u3_n3164 , _u10_u3_n3163 , _u10_u3_n3162 ,_u10_u3_n3161 , _u10_u3_n3160 , _u10_u3_n3159 , _u10_u3_n3158 ,_u10_u3_n3157 , _u10_u3_n3156 , _u10_u3_n3155 , _u10_u3_n3154 ,_u10_u3_n3153 , _u10_u3_n3152 , _u10_u3_n3151 , _u10_u3_n3150 ,_u10_u3_n3149 , _u10_u3_n3148 , _u10_u3_n3147 , _u10_u3_n3146 ,_u10_u3_n3145 , _u10_u3_n3144 , _u10_u3_n3143 , _u10_u3_n3142 ,_u10_u3_n3141 , _u10_u3_n3140 , _u10_u3_n3139 , _u10_u3_n3138 ,_u10_u3_n3137 , _u10_u3_n3136 , _u10_u3_n3135 , _u10_u3_n3134 ,_u10_u3_n3133 , _u10_u3_n3132 , _u10_u3_n3131 , _u10_u3_n3130 ,_u10_u3_n3129 , _u10_u3_n3128 , _u10_u3_n3127 , _u10_u3_n3126 ,_u10_u3_n3125 , _u10_u3_n3124 , _u10_u3_n3123 , _u10_u3_n3122 ,_u10_u3_n3121 , _u10_u3_n3120 , _u10_u3_n3119 , _u10_u3_n3118 ,_u10_u3_n3117 , _u10_u3_n3116 , _u10_u3_n3115 , _u10_u3_n3114 ,_u10_u3_n3113 , _u10_u3_n3112 , _u10_u3_n3111 , _u10_u3_n3110 ,_u10_u3_n3109 , _u10_u3_n3108 , _u10_u3_n3107 , _u10_u3_n3106 ,_u10_u3_n3105 , _u10_u3_n3104 , _u10_u3_n3103 , _u10_u3_n3102 ,_u10_u3_n3101 , _u10_u3_n3100 , _u10_u3_n3099 , _u10_u3_n3098 ,_u10_u3_n3097 , _u10_u3_n3096 , _u10_u3_n3095 , _u10_u3_n3094 ,_u10_u3_n3093 , _u10_u3_n3092 , _u10_u3_n3091 , _u10_u3_n3090 ,_u10_u3_n3089 , _u10_u3_n3088 , _u10_u3_n3087 , _u10_u3_n3086 ,_u10_u3_n3085 , _u10_u3_n3084 , _u10_u3_n3083 , _u10_u3_n3082 ,_u10_u3_n3081 , _u10_u3_n3080 , _u10_u3_n3079 , _u10_u3_n3078 ,_u10_u3_n3077 , _u10_u3_n3076 , _u10_u3_n3075 , _u10_u3_n3074 ,_u10_u3_n3073 , _u10_u3_n3072 , _u10_u3_n3071 , _u10_u3_n3070 ,_u10_u3_n3069 , _u10_u3_n3068 , _u10_u3_n3067 , _u10_u3_n3066 ,_u10_u3_n3065 , _u10_u3_n3064 , _u10_u3_n3063 , _u10_u3_n3062 ,_u10_u3_n3061 , _u10_u3_n3060 , _u10_u3_n3059 , _u10_u3_n3058 ,_u10_u3_n3057 , _u10_u3_n3056 , _u10_u3_n3055 , _u10_u3_n3054 ,_u10_u3_n3053 , _u10_u3_n3052 , _u10_u3_n3051 , _u10_u3_n3050 ,_u10_u3_n3049 , _u10_u3_n3048 , _u10_u3_n3047 , _u10_u3_n3046 ,_u10_u3_n3045 , _u10_u3_n3044 , _u10_u3_n3043 , _u10_u3_n3042 ,_u10_u3_n3041 , _u10_u3_n3040 , _u10_u3_n3039 , _u10_u3_n3038 ,_u10_u3_n3037 , _u10_u3_n3036 , _u10_u3_n3035 , _u10_u3_n3034 ,_u10_u3_n3033 , _u10_u3_n3032 , _u10_u3_n3031 , _u10_u3_n3030 ,_u10_u3_n3029 , _u10_u3_n3028 , _u10_u3_n3027 , _u10_u3_n3026 ,_u10_u3_n3025 , _u10_u3_n3024 , _u10_u3_n3023 , _u10_u3_n3022 ,_u10_u3_n3021 , _u10_u3_n3020 , _u10_u3_n3019 , _u10_u3_n3018 ,_u10_u3_n3017 , _u10_u3_n3016 , _u10_u3_n3015 , _u10_u3_n3014 ,_u10_u3_n3013 , _u10_u3_n3012 , _u10_u3_n3011 , _u10_u3_n3010 ,_u10_u3_n3009 , _u10_u3_n3008 , _u10_u3_n3007 , _u10_u3_n3006 ,_u10_u3_n3005 , _u10_u3_n3004 , _u10_u3_n3003 , _u10_u3_n3002 ,_u10_u3_n3001 , _u10_u3_n3000 , _u10_u3_n2999 , _u10_u3_n2998 ,_u10_u3_n2997 , _u10_u3_n2996 , _u10_u3_n2995 , _u10_u3_n2994 ,_u10_u3_n2993 , _u10_u3_n2992 , _u10_u3_n2991 , _u10_u3_n2990 ,_u10_u3_n2989 , _u10_u3_n2988 , _u10_u3_n2987 , _u10_u3_n2986 ,_u10_u3_n2985 , _u10_u3_n2984 , _u10_u3_n2983 , _u10_u3_n2982 ,_u10_u3_n2981 , _u10_u3_n2980 , _u10_u3_n2979 , _u10_u3_n2978 ,_u10_u3_n2977 , _u10_u3_n2976 , _u10_u3_n2975 , _u10_u3_n2974 ,_u10_u3_n2973 , _u10_u3_n2972 , _u10_u3_n2971 , _u10_u3_n2970 ,_u10_u3_n2969 , _u10_u3_n2968 , _u10_u3_n2967 , _u10_u3_n2966 ,_u10_u3_n2965 , _u10_u3_n2964 , _u10_u3_n2963 , _u10_u3_n2962 ,_u10_u3_n2961 , _u10_u3_n2960 , _u10_u3_n2959 , _u10_u3_n2958 ,_u10_u3_n2957 , _u10_u3_n2956 , _u10_u3_n2955 , _u10_u3_n2954 ,_u10_u3_n2953 , _u10_u3_n2952 , _u10_u3_n2951 , _u10_u3_n2950 ,_u10_u3_n2949 , _u10_u3_n2948 , _u10_u3_n2947 , _u10_u3_n2946 ,_u10_u3_n2945 , _u10_u3_n2944 , _u10_u3_n2943 , _u10_u3_n2942 ,_u10_u3_n2941 , _u10_u3_n2940 , _u10_u3_n2939 , _u10_u3_n2938 ,_u10_u3_n2937 , _u10_u3_n2936 , _u10_u3_n2935 , _u10_u3_n2934 ,_u10_u3_n2933 , _u10_u3_n2932 , _u10_u3_n2931 , _u10_u3_n2930 ,_u10_u3_n2929 , _u10_u3_n2928 , _u10_u3_n2927 , _u10_u3_n2926 ,_u10_u3_n2925 , _u10_u3_n2924 , _u10_u3_n2923 , _u10_u3_n2922 ,_u10_u3_n2921 , _u10_u3_n2920 , _u10_u3_n2919 , _u10_u3_n2918 ,_u10_u3_n2917 , _u10_u3_n2916 , _u10_u3_n2915 , _u10_u3_n2914 ,_u10_u3_n2913 , _u10_u3_n2912 , _u10_u3_n2911 , _u10_u3_n2910 ,_u10_u3_n2909 , _u10_u3_n2908 , _u10_u3_n2907 , _u10_u3_n2906 ,_u10_u3_n2905 , _u10_u3_n2904 , _u10_u3_n2903 , _u10_u3_n2902 ,_u10_u3_n2901 , _u10_u3_n2900 , _u10_u3_n2899 , _u10_u3_n2898 ,_u10_u3_n2897 , _u10_u3_n2896 , _u10_u3_n2895 , _u10_u3_n2894 ,_u10_u3_n2893 , _u10_u3_n2892 , _u10_u3_n2891 , _u10_u3_n2890 ,_u10_u3_n2889 , _u10_u3_n2888 , _u10_u3_n2887 , _u10_u3_n2886 ,_u10_u3_n2885 , _u10_u3_n2884 , _u10_u3_n2883 , _u10_u3_n2882 ,_u10_u3_n2881 , _u10_u3_n2880 , _u10_u3_n2879 , _u10_u3_n2878 ,_u10_u3_n2877 , _u10_u3_n2876 , _u10_u3_n2875 , _u10_u3_n2874 ,_u10_u3_n2873 , _u10_u3_n2872 , _u10_u3_n2871 , _u10_u3_n2870 ,_u10_u3_n2869 , _u10_u3_n2868 , _u10_u3_n2867 , _u10_u3_n2866 ,_u10_u3_n2865 , _u10_u3_n2864 , _u10_u3_n2863 , _u10_u3_n2862 ,_u10_u3_n2861 , _u10_u3_n2860 , _u10_u3_n2859 , _u10_u3_n2858 ,_u10_u3_n2857 , _u10_u3_n2856 , _u10_u3_n2855 , _u10_u3_n2854 ,_u10_u3_n2853 , _u10_u3_n2852 , _u10_u3_n2851 , _u10_u3_n2850 ,_u10_u3_n2849 , _u10_u3_n2848 , _u10_u3_n2847 , _u10_u3_n2846 ,_u10_u3_n2845 , _u10_u3_n2844 , _u10_u3_n2843 , _u10_u3_n2842 ,_u10_u3_n2841 , _u10_u3_n2840 , _u10_u3_n2839 , _u10_u3_n2838 ,_u10_u3_n2837 , _u10_u3_n2836 , _u10_u3_n2835 , _u10_u3_n2834 ,_u10_u3_n2833 , _u10_u3_n2832 , _u10_u3_n2831 , _u10_u3_n2830 ,_u10_u3_n2829 , _u10_u3_n2828 , _u10_u3_n2827 , _u10_u3_n2826 ,_u10_u3_n2825 , _u10_u3_n2824 , _u10_u3_n2823 , _u10_u3_n2822 ,_u10_u3_n2821 , _u10_u3_n2820 , _u10_u3_n2819 , _u10_u3_n2818 ,_u10_u3_n2817 , _u10_u3_n2816 , _u10_u3_n2815 , _u10_u3_n2814 ,_u10_u3_n2813 , _u10_u3_n2812 , _u10_u3_n2811 , _u10_u3_n2810 ,_u10_u3_n2809 , _u10_u3_n2808 , _u10_u3_n2807 , _u10_u3_n2806 ,_u10_u3_n2805 , _u10_u3_n2804 , _u10_u3_n2803 , _u10_u3_n2802 ,_u10_u3_n2801 , _u10_u3_n2800 , _u10_u3_n2799 , _u10_u3_n2798 ,_u10_u3_n2797 , _u10_u3_n2796 , _u10_u3_n2795 , _u10_u3_n2794 ,_u10_u3_n2793 , _u10_u3_n2792 , _u10_u3_n2791 , _u10_u3_n2790 ,_u10_u3_n2789 , _u10_u3_n2788 , _u10_u3_n2787 , _u10_u3_n2786 ,_u10_u3_n2785 , _u10_u3_n2784 , _u10_u3_n2783 , _u10_u3_n2782 ,_u10_u3_n2781 , _u10_u3_n2780 , _u10_u3_n2779 , _u10_u3_n2778 ,_u10_u3_n2777 , _u10_u3_n2776 , _u10_u3_n2775 , _u10_u3_n2774 ,_u10_u3_n2773 , _u10_u3_n2772 , _u10_u3_n2771 , _u10_u3_n2770 ,_u10_u3_n2769 , _u10_u3_n2768 , _u10_u3_n2767 , _u10_u3_n2766 ,_u10_u3_n2765 , _u10_u3_n2764 , _u10_u3_n2763 , _u10_u3_n2762 ,_u10_u3_n2761 , _u10_u3_n2760 , _u10_u3_n2759 , _u10_u3_n2758 ,_u10_u3_n2757 , _u10_u3_n2756 , _u10_u3_n2755 , _u10_u3_n2754 ,_u10_u3_n2753 , _u10_u3_n2752 , _u10_u3_n2751 , _u10_u3_n2750 ,_u10_u3_n2749 , _u10_u3_n2748 , _u10_u3_n2747 , _u10_u3_n2746 ,_u10_u3_n2745 , _u10_u3_n2744 , _u10_u3_n2743 , _u10_u3_n2742 ,_u10_u3_n2741 , _u10_u3_n2740 , _u10_u3_n2739 , _u10_u3_n2738 ,_u10_u3_n2737 , _u10_u3_n2736 , _u10_u3_n2735 , _u10_u3_n2734 ,_u10_u3_n2733 , _u10_u3_n2732 , _u10_u3_n2731 , _u10_u3_n2730 ,_u10_u3_n2729 , _u10_u3_n2728 , _u10_u3_n2727 , _u10_u3_n2726 ,_u10_u3_n2725 , _u10_u3_n2724 , _u10_u3_n2723 , _u10_u3_n2722 ,_u10_u3_n2721 , _u10_u3_n2720 , _u10_u3_n2719 , _u10_u3_n2718 ,_u10_u3_n2717 , _u10_u3_n2716 , _u10_u3_n2715 , _u10_u3_n2714 ,_u10_u3_n2713 , _u10_u3_n2712 , _u10_u3_n2711 , _u10_u3_n2710 ,_u10_u3_n2709 , _u10_u3_n2708 , _u10_u3_n2707 , _u10_u3_n2706 ,_u10_u3_n2705 , _u10_u3_n2704 , _u10_u3_n2703 , _u10_u3_n2702 ,_u10_u3_n2701 , _u10_u3_n2700 , _u10_u3_n2699 , _u10_u3_n2698 ,_u10_u3_n2697 , _u10_u3_n2696 , _u10_u3_n2695 , _u10_u3_n2694 ,_u10_u3_n2693 , _u10_u3_n2692 , _u10_u3_n2691 , _u10_u3_n2690 ,_u10_u3_n2689 , _u10_u3_n2688 , _u10_u3_n2687 , _u10_u3_n2686 ,_u10_u3_n2685 , _u10_u3_n2684 , _u10_u3_n2683 , _u10_u3_n2682 ,_u10_u3_n2681 , _u10_u3_n2680 , _u10_u3_n2679 , _u10_u3_n2678 ,_u10_u3_n2677 , _u10_u3_n2676 , _u10_u3_n2675 , _u10_u3_n2674 ,_u10_u3_n2673 , _u10_u3_n2672 , _u10_u3_n2671 , _u10_u3_n2670 ,_u10_u3_n2669 , _u10_u3_n2668 , _u10_u3_n2667 , _u10_u3_n2666 ,_u10_u3_n2665 , _u10_u3_n2664 , _u10_u3_n2663 , _u10_u3_n2662 ,_u10_u3_n2661 , _u10_u3_n2660 , _u10_u3_n2659 , _u10_u3_n2658 ,_u10_u3_n2657 , _u10_u3_n2656 , _u10_u3_n2655 , _u10_u3_n2654 ,_u10_u3_n2653 , _u10_u3_n2652 , _u10_u3_n2651 , _u10_u3_n2650 ,_u10_u3_n2649 , _u10_u3_n2648 , _u10_u3_n2647 , _u10_u3_n2646 ,_u10_u3_n2645 , _u10_u3_n2644 , _u10_u3_n2643 , _u10_u3_n2642 ,_u10_u3_n2641 , _u10_u3_n2640 , _u10_u3_n2639 , _u10_u3_n2638 ,_u10_u3_n2637 , _u10_u3_n2636 , _u10_u3_n2635 , _u10_u3_n2634 ,_u10_u3_n2633 , _u10_u3_n2632 , _u10_u3_n2631 , _u10_u3_n2630 ,_u10_u3_n2629 , _u10_u3_n2628 , _u10_u3_n2627 , _u10_u3_n2626 ,_u10_u3_n2625 , _u10_u3_n2624 , _u10_u3_n2623 , _u10_u3_n2622 ,_u10_u3_n2621 , _u10_u3_n2620 , _u10_u3_n2619 , _u10_u3_n2618 ,_u10_u3_n2617 , _u10_u3_n2616 , _u10_u3_n2615 , _u10_u3_n2614 ,_u10_u3_n2613 , _u10_u3_n2612 , _u10_u3_n2611 , _u10_u3_n2610 ,_u10_u3_n2609 , _u10_u3_n2608 , _u10_u3_n2607 , _u10_u3_n2606 ,_u10_u3_n2605 , _u10_u3_n2604 , _u10_u3_n2603 , _u10_u3_n2602 ,_u10_u3_n2601 , _u10_u3_n2600 , _u10_u3_n2599 , _u10_u3_n2598 ,_u10_u3_n2597 , _u10_u3_n2596 , _u10_u3_n2595 , _u10_u3_n2594 ,_u10_u3_n2593 , _u10_u3_n2592 , _u10_u3_n2591 , _u10_u3_n2590 ,_u10_u3_n2589 , _u10_u3_n2588 , _u10_u3_n2587 , _u10_u3_n2586 ,_u10_u3_n2585 , _u10_u3_n2584 , _u10_u3_n2583 , _u10_u3_n2582 ,_u10_u3_n2581 , _u10_u3_n2580 , _u10_u3_n2579 , _u10_u3_n2578 ,_u10_u3_n2577 , _u10_u3_n2576 , _u10_u3_n2575 , _u10_u3_n2574 ,_u10_u3_n2573 , _u10_u3_n2572 , _u10_u3_n2571 , _u10_u3_n2570 ,_u10_u3_n2569 , _u10_u3_n2568 , _u10_u3_n2567 , _u10_u3_n2566 ,_u10_u3_n2565 , _u10_u3_n2564 , _u10_u3_n2563 , _u10_u3_n2562 ,_u10_u3_n2561 , _u10_u3_n2560 , _u10_u3_n2559 , _u10_u3_n2558 ,_u10_u3_n2557 , _u10_u3_n2556 , _u10_u3_n2555 , _u10_u3_n2554 ,_u10_u3_n2553 , _u10_u3_n2552 , _u10_u3_n2551 , _u10_u3_n2550 ,_u10_u3_n2549 , _u10_u3_n2548 , _u10_u3_n2547 , _u10_u3_n2546 ,_u10_u3_n2545 , _u10_u3_n2544 , _u10_u3_n2543 , _u10_u3_n2542 ,_u10_u3_n2541 , _u10_u3_n2540 , _u10_u3_n2539 , _u10_u3_n2538 ,_u10_u3_n2537 , _u10_u3_n2536 , _u10_u3_n2535 , _u10_u3_n2534 ,_u10_u3_n2533 , _u10_u3_n2532 , _u10_u3_n2531 , _u10_u3_n2530 ,_u10_u3_n2529 , _u10_u3_n2528 , _u10_u3_n2527 , _u10_u3_n2526 ,_u10_u3_n2525 , _u10_u3_n2524 , _u10_u3_n2523 , _u10_u3_n2522 ,_u10_u3_n2521 , _u10_u3_n2520 , _u10_u3_n2519 , _u10_u3_n2518 ,_u10_u3_n2517 , _u10_u3_n2516 , _u10_u3_n2515 , _u10_u3_n2514 ,_u10_u3_n2513 , _u10_u3_n2512 , _u10_u3_n2511 , _u10_u3_n2510 ,_u10_u3_n2509 , _u10_u3_n2508 , _u10_u3_n2507 , _u10_u3_n2506 ,_u10_u3_n2505 , _u10_u3_n2504 , _u10_u3_n2503 , _u10_u3_n2502 ,_u10_u3_n2501 , _u10_u3_n2500 , _u10_u3_n2499 , _u10_u3_n2498 ,_u10_u3_n2497 , _u10_u3_n2496 , _u10_u3_n2495 , _u10_u3_n2494 ,_u10_u3_n2493 , _u10_u3_n2492 , _u10_u3_n2491 , _u10_u3_n2490 ,_u10_u3_n2489 , _u10_u3_n2488 , _u10_u3_n2487 , _u10_u3_n2486 ,_u10_u3_n2485 , _u10_u3_n2484 , _u10_u3_n2483 , _u10_u3_n2482 ,_u10_u3_n2481 , _u10_u3_n2480 , _u10_u3_n2479 , _u10_u3_n2478 ,_u10_u3_n2477 , _u10_u3_n2476 , _u10_u3_n2475 , _u10_u3_n2474 ,_u10_u3_n2473 , _u10_u3_n2472 , _u10_u3_n2471 , _u10_u3_n2470 ,_u10_u3_n2469 , _u10_u3_n2468 , _u10_u3_n2467 , _u10_u3_n2466 ,_u10_u3_n2465 , _u10_u3_n2464 , _u10_u3_n2463 , _u10_u3_n2462 ,_u10_u3_n2461 , _u10_u3_n2460 , _u10_u3_n2459 , _u10_u3_n2458 ,_u10_u3_n2457 , _u10_u3_n2456 , _u10_u3_n2455 , _u10_u3_n2454 ,_u10_u3_n2453 , _u10_u3_n2452 , _u10_u3_n2451 , _u10_u3_n2450 ,_u10_u3_n2449 , _u10_u3_n2448 , _u10_u3_n2447 , _u10_u3_n2446 ,_u10_u3_n2445 , _u10_u3_n2444 , _u10_u3_n2443 , _u10_u3_n2442 ,_u10_u3_n2441 , _u10_u3_n2440 , _u10_u3_n2439 , _u10_u3_n2438 ,_u10_u3_n2437 , _u10_u3_n2436 , _u10_u3_n2435 , _u10_u3_n2434 ,_u10_u3_n2433 , _u10_u3_n2432 , _u10_u3_n2431 , _u10_u3_n2430 ,_u10_u3_n2429 , _u10_u3_n2428 , _u10_u3_n2427 , _u10_u3_n2426 ,_u10_u3_n2425 , _u10_u3_n2424 , _u10_u3_n2423 , _u10_u3_n2422 ,_u10_u3_n2421 , _u10_u3_n2420 , _u10_u3_n2419 , _u10_u3_n2418 ,_u10_u3_n2417 , _u10_u3_n2416 , _u10_u3_n2415 , _u10_u3_n2414 ,_u10_u3_n2413 , _u10_u3_n2412 , _u10_u3_n2411 , _u10_u3_n2410 ,_u10_u3_n2409 , _u10_u3_n2408 , _u10_u3_n2407 , _u10_u3_n2406 ,_u10_u3_n2405 , _u10_u3_n2404 , _u10_u3_n2403 , _u10_u3_n2402 ,_u10_u3_n2401 , _u10_u3_n2400 , _u10_u3_n2399 , _u10_u3_n2398 ,_u10_u3_n2397 , _u10_u3_n2396 , _u10_u3_n2395 , _u10_u3_n2394 ,_u10_u3_n2393 , _u10_u3_n2392 , _u10_u3_n2391 , _u10_u3_n2390 ,_u10_u3_n2389 , _u10_u3_n2388 , _u10_u3_n2387 , _u10_u3_n2386 ,_u10_u3_n2385 , _u10_u3_n2384 , _u10_u3_n2383 , _u10_u3_n2382 ,_u10_u3_n2381 , _u10_u3_n2380 , _u10_u3_n2379 , _u10_u3_n2378 ,_u10_u3_n2377 , _u10_u3_n2376 , _u10_u3_n2375 , _u10_u3_n2374 ,_u10_u3_n2373 , _u10_u3_n2372 , _u10_u3_n2371 , _u10_u3_n2370 ,_u10_u3_n2369 , _u10_u3_n2368 , _u10_u3_n2367 , _u10_u3_n2366 ,_u10_u3_n2365 , _u10_u3_n2364 , _u10_u3_n2363 , _u10_u3_n2362 ,_u10_u3_n2361 , _u10_u3_n2360 , _u10_u3_n2359 , _u10_u3_n2358 ,_u10_u3_n2357 , _u10_u3_n2356 , _u10_u3_n2355 , _u10_u3_n2354 ,_u10_u3_n2353 , _u10_u3_n2352 , _u10_u3_n2351 , _u10_u3_n2350 ,_u10_u3_n2349 , _u10_u3_n2348 , _u10_u3_n2347 , _u10_u3_n2346 ,_u10_u3_n2345 , _u10_u3_n2344 , _u10_u3_n2343 , _u10_u3_n2342 ,_u10_u3_n2341 , _u10_u3_n2340 , _u10_u3_n2339 , _u10_u3_n2338 ,_u10_u3_n2337 , _u10_u3_n2336 , _u10_u3_n2335 , _u10_u3_n2334 ,_u10_u3_n2333 , _u10_u3_n2332 , _u10_u3_n2331 , _u10_u3_n2330 ,_u10_u3_n2329 , _u10_u3_n2328 , _u10_u3_n2327 , _u10_u3_n2326 ,_u10_u3_n2325 , _u10_u3_n2324 , _u10_u3_n2323 , _u10_u3_n2322 ,_u10_u3_n2321 , _u10_u3_n2320 , _u10_u3_n2319 , _u10_u3_n2318 ,_u10_u3_n2317 , _u10_u3_n2316 , _u10_u3_n2315 , _u10_u3_n2314 ,_u10_u3_n2313 , _u10_u3_n2312 , _u10_u3_n2311 , _u10_u3_n2310 ,_u10_u3_n2309 , _u10_u3_n2308 , _u10_u3_n2307 , _u10_u3_n2306 ,_u10_u3_n2305 , _u10_u3_n2304 , _u10_u3_n2303 , _u10_u3_n2302 ,_u10_u3_n2301 , _u10_u3_n2300 , _u10_u3_n2299 , _u10_u3_n2298 ,_u10_u3_n2297 , _u10_u3_n2296 , _u10_u3_n2295 , _u10_u3_n2294 ,_u10_u3_n2293 , _u10_u3_n2292 , _u10_u3_n2291 , _u10_u3_n2290 ,_u10_u3_n2289 , _u10_u3_n2288 , _u10_u3_n2287 , _u10_u3_n2286 ,_u10_u3_n2285 , _u10_u3_n2284 , _u10_u3_n2283 , _u10_u3_n2282 ,_u10_u3_n2281 , _u10_u3_n2280 , _u10_u3_n2279 , _u10_u3_n2278 ,_u10_u3_n2277 , _u10_u3_n2276 , _u10_u3_n2275 , _u10_u3_n2274 ,_u10_u3_n2273 , _u10_u3_n2272 , _u10_u3_n2271 , _u10_u3_n2270 ,_u10_u3_n2269 , _u10_u3_n2268 , _u10_u3_n2267 , _u10_u3_n2266 ,_u10_u3_n2265 , _u10_u3_n2264 , _u10_u3_n2263 , _u10_u3_n2262 ,_u10_u3_n2261 , _u10_u3_n2260 , _u10_u3_n2259 , _u10_u3_n2258 ,_u10_u3_n2257 , _u10_u3_n2256 , _u10_u3_n2255 , _u10_u3_n2254 ,_u10_u3_n2253 , _u10_u3_n2252 , _u10_u3_n2251 , _u10_u3_n2250 ,_u10_u3_n2249 , _u10_u3_n2248 , _u10_u3_n2247 , _u10_u3_n2246 ,_u10_u3_n2245 , _u10_u3_n2244 , _u10_u3_n2243 , _u10_u3_n2242 ,_u10_u3_n2241 , _u10_u3_n2240 , _u10_u3_n2239 , _u10_u3_n2238 ,_u10_u3_n2237 , _u10_u3_n2236 , _u10_u3_n2235 , _u10_u3_n2234 ,_u10_u3_n2233 , _u10_u3_n2232 , _u10_u3_n2231 , _u10_u3_n2230 ,_u10_u3_n2229 , _u10_u3_n2228 , _u10_u3_n2227 , _u10_u3_n2226 ,_u10_u3_n2225 , _u10_u3_n2224 , _u10_u3_n2223 , _u10_u3_n2222 ,_u10_u3_n2221 , _u10_u3_n2220 , _u10_u3_n2219 , _u10_u3_n2218 ,_u10_u3_n2217 , _u10_u3_n2216 , _u10_u3_n2215 , _u10_u3_n2214 ,_u10_u3_n2213 , _u10_u3_n2212 , _u10_u3_n2211 , _u10_u3_n2210 ,_u10_u3_n2209 , _u10_u3_n2208 , _u10_u3_n2207 , _u10_u3_n2206 ,_u10_u3_n2205 , _u10_u3_n2204 , _u10_u3_n2203 , _u10_u3_n2202 ,_u10_u3_n2201 , _u10_u3_n2200 , _u10_u3_n2199 , _u10_u3_n2198 ,_u10_u3_n2197 , _u10_u3_n2196 , _u10_u3_n2195 , _u10_u3_n2194 ,_u10_u3_n2193 , _u10_u3_n2192 , _u10_u3_n2191 , _u10_u3_n2190 ,_u10_u3_n2189 , _u10_u3_n2188 , _u10_u3_n2187 , _u10_u3_n2186 ,_u10_u3_n2185 , _u10_u3_n2184 , _u10_u3_n2183 , _u10_u3_n2182 ,_u10_u3_n2181 , _u10_u3_n2180 , _u10_u3_n2179 , _u10_u3_n2178 ,_u10_u3_n2177 , _u10_u3_n2176 , _u10_u3_n2175 , _u10_u3_n2174 ,_u10_u3_n2173 , _u10_u3_n2172 , _u10_u3_n2171 , _u10_u3_n2170 ,_u10_u3_n2169 , _u10_u3_n2168 , _u10_u3_n2167 , _u10_u3_n2166 ,_u10_u3_n2165 , _u10_u3_n2164 , _u10_u3_n2163 , _u10_u3_n2162 ,_u10_u3_n2161 , _u10_u3_n2160 , _u10_u3_n2159 , _u10_u3_n2158 ,_u10_u3_n2157 , _u10_u3_n2156 , _u10_u3_n2155 , _u10_u3_n2154 ,_u10_u3_n2153 , _u10_u3_n2152 , _u10_u3_n2151 , _u10_u3_n2150 ,_u10_u3_n2149 , _u10_u3_n2148 , _u10_u3_n2147 , _u10_u3_n2146 ,_u10_u3_n2145 , _u10_u3_n2144 , _u10_u3_n2143 , _u10_u3_n2142 ,_u10_u3_n2141 , _u10_u3_n2140 , _u10_u3_n2139 , _u10_u3_n2138 ,_u10_u3_n2137 , _u10_u3_n2136 , _u10_u3_n2135 , _u10_u3_n2134 ,_u10_u3_n2133 , _u10_u3_n2132 , _u10_u3_n2131 , _u10_u3_n2130 ,_u10_u3_n2129 , _u10_u3_n2128 , _u10_u3_n2127 , _u10_u3_n2126 ,_u10_u3_n2125 , _u10_u3_n2124 , _u10_u3_n2123 , _u10_u3_n2122 ,_u10_u3_n2121 , _u10_u3_n2120 , _u10_u3_n2119 , _u10_u3_n2118 ,_u10_u3_n2117 , _u10_u3_n2116 , _u10_u3_n2115 , _u10_u3_n2114 ,_u10_u3_n2113 , _u10_u3_n2112 , _u10_u3_n2111 , _u10_u3_n2110 ,_u10_u3_n2109 , _u10_u3_n2108 , _u10_u3_n2107 , _u10_u3_n2106 ,_u10_u3_n2105 , _u10_u3_n2104 , _u10_u3_n2103 , _u10_u3_n2102 ,_u10_u3_n2101 , _u10_u3_n2100 , _u10_u3_n2099 , _u10_u3_n2098 ,_u10_u3_n2097 , _u10_u3_n2096 , _u10_u3_n2095 , _u10_u3_n2094 ,_u10_u3_n2093 , _u10_u3_n2092 , _u10_u3_n2091 , _u10_u3_n2090 ,_u10_u3_n2089 , _u10_u3_n2088 , _u10_u3_n2087 , _u10_u3_n2086 ,_u10_u3_n2085 , _u10_u3_n2084 , _u10_u3_n2083 , _u10_u3_n2082 ,_u10_u3_n2081 , _u10_u3_n2080 , _u10_u3_n2079 , _u10_u3_n2078 ,_u10_u3_n2077 , _u10_u3_n2076 , _u10_u3_n2075 , _u10_u3_n2074 ,_u10_u3_n2073 , _u10_u3_n2072 , _u10_u3_n2071 , _u10_u3_n2070 ,_u10_u3_n2069 , _u10_u3_n2068 , _u10_u3_n2067 , _u10_u3_n2066 ,_u10_u3_n2065 , _u10_u3_n2064 , _u10_u3_n2063 , _u10_u3_n2062 ,_u10_u3_n2061 , _u10_u3_n2060 , _u10_u3_n2059 , _u10_u3_n2058 ,_u10_u3_n2057 , _u10_u3_n2056 , _u10_u3_n2055 , _u10_u3_n2054 ,_u10_u3_n2053 , _u10_u3_n2052 , _u10_u3_n2051 , _u10_u3_n2050 ,_u10_u3_n2049 , _u10_u3_n2048 , _u10_u3_n2047 , _u10_u3_n2046 ,_u10_u3_n2045 , _u10_u3_n2044 , _u10_u3_n2043 , _u10_u3_n2042 ,_u10_u3_n2041 , _u10_u3_n2040 , _u10_u3_n2039 , _u10_u3_n2038 ,_u10_u3_n2037 , _u10_u3_n2036 , _u10_u3_n2035 , _u10_u3_n2034 ,_u10_u3_n2033 , _u10_u3_n2032 , _u10_u3_n2031 , _u10_u3_n2030 ,_u10_u3_n2029 , _u10_u3_n2028 , _u10_u3_n2027 , _u10_u3_n2026 ,_u10_u3_n2025 , _u10_u3_n2024 , _u10_u3_n2023 , _u10_u3_n2022 ,_u10_u3_n2021 , _u10_u3_n2020 , _u10_u3_n2019 , _u10_u3_n2018 ,_u10_u3_n2017 , _u10_u3_n2016 , _u10_u3_n2015 , _u10_u3_n2014 ,_u10_u3_n2013 , _u10_u3_n2012 , _u10_u3_n2011 , _u10_u3_n2010 ,_u10_u3_n2009 , _u10_u3_n2008 , _u10_u3_n2007 , _u10_u3_n2006 ,_u10_u3_n2005 , _u10_u3_n2004 , _u10_u3_n2003 , _u10_u3_n2002 ,_u10_u3_n2001 , _u10_u3_n2000 , _u10_u3_n1999 , _u10_u3_n1998 ,_u10_u3_n1997 , _u10_u3_n1996 , _u10_u3_n1995 , _u10_u3_n1994 ,_u10_u3_n1993 , _u10_u3_n1992 , _u10_u3_n1991 , _u10_u3_n1990 ,_u10_u3_n1989 , _u10_u3_n1988 , _u10_u3_n1987 , _u10_u3_n1986 ,_u10_u3_n1985 , _u10_u3_n1984 , _u10_u3_n1983 , _u10_u3_n1982 ,_u10_u3_n1981 , _u10_u3_n1980 , _u10_u3_n1979 , _u10_u3_n1978 ,_u10_u3_n1977 , _u10_u3_n1976 , _u10_u3_n1975 , _u10_u3_n1974 ,_u10_u3_n1973 , _u10_u3_n1972 , _u10_u3_n1971 , _u10_u3_n1970 ,_u10_u3_n1969 , _u10_u3_n1968 , _u10_u3_n1967 , _u10_u3_n1966 ,_u10_u3_n1965 , _u10_u3_n1964 , _u10_u3_n1963 , _u10_u3_n1962 ,_u10_u3_n1961 , _u10_u3_n1960 , _u10_u3_n1959 , _u10_u3_n1958 ,_u10_u3_n1957 , _u10_u3_n1956 , _u10_u3_n1955 , _u10_u3_n1954 ,_u10_u3_n1953 , _u10_u3_n1952 , _u10_u3_n1951 , _u10_u3_n1950 ,_u10_u3_n1949 , _u10_u3_n1948 , _u10_u3_n1947 , _u10_u3_n1946 ,_u10_u3_n1945 , _u10_u3_n1944 , _u10_u3_n1943 , _u10_u3_n1942 ,_u10_u3_n1941 , _u10_u3_n1940 , _u10_u3_n1939 , _u10_u3_n1938 ,_u10_u3_n1937 , _u10_u3_n1936 , _u10_u3_n1935 , _u10_u3_n1934 ,_u10_u3_n1933 , _u10_u3_n1932 , _u10_u3_n1931 , _u10_u3_n1930 ,_u10_u3_n1929 , _u10_u3_n1928 , _u10_u3_n1927 , _u10_u3_n1926 ,_u10_u3_n1925 , _u10_u3_n1924 , _u10_u3_n1923 , _u10_u3_n1922 ,_u10_u3_n1921 , _u10_u3_n1920 , _u10_u3_n1919 , _u10_u3_n1918 ,_u10_u3_n1917 , _u10_u3_n1916 , _u10_u3_n1915 , _u10_u3_n1914 ,_u10_u3_n1913 , _u10_u3_n1912 , _u10_u3_n1911 , _u10_u3_n1910 ,_u10_u3_n1909 , _u10_u3_n1908 , _u10_u3_n1907 , _u10_u3_n1906 ,_u10_u3_n1905 , _u10_u3_n1904 , _u10_u3_n1903 , _u10_u3_n1902 ,_u10_u3_n1901 , _u10_u3_n1900 , _u10_u3_n1899 , _u10_u3_n1898 ,_u10_u3_n1897 , _u10_u3_n1896 , _u10_u3_n1895 , _u10_u3_n1894 ,_u10_u3_n1893 , _u10_u3_n1892 , _u10_u3_n1891 , _u10_u3_n1890 ,_u10_u3_n1889 , _u10_u3_n1888 , _u10_u3_n1887 , _u10_u3_n1886 ,_u10_u3_n1885 , _u10_u3_n1884 , _u10_u3_n1883 , _u10_u3_n1882 ,_u10_u3_n1881 , _u10_u3_n1880 , _u10_u3_n1879 , _u10_u3_n1878 ,_u10_u3_n1877 , _u10_u3_n1876 , _u10_u3_n1875 , _u10_u3_n1874 ,_u10_u3_n1873 , _u10_u3_n1872 , _u10_u3_n1871 , _u10_u3_n1870 ,_u10_u3_n1869 , _u10_u3_n1868 , _u10_u3_n1867 , _u10_u3_n1866 ,_u10_u3_n1865 , _u10_u3_n1864 , _u10_u3_n1863 , _u10_u3_n1862 ,_u10_u3_n1861 , _u10_u3_n1860 , _u10_u3_n1859 , _u10_u3_n1858 ,_u10_u3_n1857 , _u10_u3_n1856 , _u10_u3_n1855 , _u10_u3_n1854 ,_u10_u3_n1853 , _u10_u3_n1852 , _u10_u3_n1851 , _u10_u3_n1850 ,_u10_u3_n1849 , _u10_u3_n1848 , _u10_u3_n1847 , _u10_u3_n1846 ,_u10_u3_n1845 , _u10_u3_n1844 , _u10_u3_n1843 , _u10_u3_n1842 ,_u10_u3_n1841 , _u10_u3_n1840 , _u10_u3_n1839 , _u10_u3_n1838 ,_u10_u3_n1837 , _u10_u3_n1836 , _u10_u3_n1835 , _u10_u3_n1834 ,_u10_u3_n1833 , _u10_u3_n1832 , _u10_u3_n1831 , _u10_u3_n1830 ,_u10_u3_n1829 , _u10_u3_n1828 , _u10_u3_n1827 , _u10_u3_n1826 ,_u10_u3_n1825 , _u10_u3_n1824 , _u10_u3_n1823 , _u10_u3_n1822 ,_u10_u3_n1821 , _u10_u3_n1820 , _u10_u3_n1819 , _u10_u3_n1818 ,_u10_u3_n1817 , _u10_u3_n1816 , _u10_u3_n1815 , _u10_u3_n1814 ,_u10_u3_n1813 , _u10_u3_n1812 , _u10_u3_n1811 , _u10_u3_n1810 ,_u10_u3_n1809 , _u10_u3_n1808 , _u10_u4_n3416 , _u10_u4_n3415 ,_u10_u4_n3414 , _u10_u4_n3413 , _u10_u4_n3412 , _u10_u4_n3411 ,_u10_u4_n3410 , _u10_u4_n3409 , _u10_u4_n3408 , _u10_u4_n3407 ,_u10_u4_n3406 , _u10_u4_n3405 , _u10_u4_n3404 , _u10_u4_n3403 ,_u10_u4_n3402 , _u10_u4_n3401 , _u10_u4_n3400 , _u10_u4_n3399 ,_u10_u4_n3398 , _u10_u4_n3397 , _u10_u4_n3396 , _u10_u4_n3395 ,_u10_u4_n3394 , _u10_u4_n3393 , _u10_u4_n3392 , _u10_u4_n3391 ,_u10_u4_n3390 , _u10_u4_n3389 , _u10_u4_n3388 , _u10_u4_n3387 ,_u10_u4_n3386 , _u10_u4_n3385 , _u10_u4_n3384 , _u10_u4_n3383 ,_u10_u4_n3382 , _u10_u4_n3381 , _u10_u4_n3380 , _u10_u4_n3379 ,_u10_u4_n3378 , _u10_u4_n3377 , _u10_u4_n3376 , _u10_u4_n3375 ,_u10_u4_n3374 , _u10_u4_n3373 , _u10_u4_n3372 , _u10_u4_n3371 ,_u10_u4_n3370 , _u10_u4_n3369 , _u10_u4_n3368 , _u10_u4_n3367 ,_u10_u4_n3366 , _u10_u4_n3365 , _u10_u4_n3364 , _u10_u4_n3363 ,_u10_u4_n3362 , _u10_u4_n3361 , _u10_u4_n3360 , _u10_u4_n3359 ,_u10_u4_n3358 , _u10_u4_n3357 , _u10_u4_n3356 , _u10_u4_n3355 ,_u10_u4_n3354 , _u10_u4_n3353 , _u10_u4_n3352 , _u10_u4_n3351 ,_u10_u4_n3350 , _u10_u4_n3349 , _u10_u4_n3348 , _u10_u4_n3347 ,_u10_u4_n3346 , _u10_u4_n3345 , _u10_u4_n3344 , _u10_u4_n3343 ,_u10_u4_n3342 , _u10_u4_n3341 , _u10_u4_n3340 , _u10_u4_n3339 ,_u10_u4_n3338 , _u10_u4_n3337 , _u10_u4_n3336 , _u10_u4_n3335 ,_u10_u4_n3334 , _u10_u4_n3333 , _u10_u4_n3332 , _u10_u4_n3331 ,_u10_u4_n3330 , _u10_u4_n3329 , _u10_u4_n3328 , _u10_u4_n3327 ,_u10_u4_n3326 , _u10_u4_n3325 , _u10_u4_n3324 , _u10_u4_n3323 ,_u10_u4_n3322 , _u10_u4_n3321 , _u10_u4_n3320 , _u10_u4_n3319 ,_u10_u4_n3318 , _u10_u4_n3317 , _u10_u4_n3316 , _u10_u4_n3315 ,_u10_u4_n3314 , _u10_u4_n3313 , _u10_u4_n3312 , _u10_u4_n3311 ,_u10_u4_n3310 , _u10_u4_n3309 , _u10_u4_n3308 , _u10_u4_n3307 ,_u10_u4_n3306 , _u10_u4_n3305 , _u10_u4_n3304 , _u10_u4_n3303 ,_u10_u4_n3302 , _u10_u4_n3301 , _u10_u4_n3300 , _u10_u4_n3299 ,_u10_u4_n3298 , _u10_u4_n3297 , _u10_u4_n3296 , _u10_u4_n3295 ,_u10_u4_n3294 , _u10_u4_n3293 , _u10_u4_n3292 , _u10_u4_n3291 ,_u10_u4_n3290 , _u10_u4_n3289 , _u10_u4_n3288 , _u10_u4_n3287 ,_u10_u4_n3286 , _u10_u4_n3285 , _u10_u4_n3284 , _u10_u4_n3283 ,_u10_u4_n3282 , _u10_u4_n3281 , _u10_u4_n3280 , _u10_u4_n3279 ,_u10_u4_n3278 , _u10_u4_n3277 , _u10_u4_n3276 , _u10_u4_n3275 ,_u10_u4_n3274 , _u10_u4_n3273 , _u10_u4_n3272 , _u10_u4_n3271 ,_u10_u4_n3270 , _u10_u4_n3269 , _u10_u4_n3268 , _u10_u4_n3267 ,_u10_u4_n3266 , _u10_u4_n3265 , _u10_u4_n3264 , _u10_u4_n3263 ,_u10_u4_n3262 , _u10_u4_n3261 , _u10_u4_n3260 , _u10_u4_n3259 ,_u10_u4_n3258 , _u10_u4_n3257 , _u10_u4_n3256 , _u10_u4_n3255 ,_u10_u4_n3254 , _u10_u4_n3253 , _u10_u4_n3252 , _u10_u4_n3251 ,_u10_u4_n3250 , _u10_u4_n3249 , _u10_u4_n3248 , _u10_u4_n3247 ,_u10_u4_n3246 , _u10_u4_n3245 , _u10_u4_n3244 , _u10_u4_n3243 ,_u10_u4_n3242 , _u10_u4_n3241 , _u10_u4_n3240 , _u10_u4_n3239 ,_u10_u4_n3238 , _u10_u4_n3237 , _u10_u4_n3236 , _u10_u4_n3235 ,_u10_u4_n3234 , _u10_u4_n3233 , _u10_u4_n3232 , _u10_u4_n3231 ,_u10_u4_n3230 , _u10_u4_n3229 , _u10_u4_n3228 , _u10_u4_n3227 ,_u10_u4_n3226 , _u10_u4_n3225 , _u10_u4_n3224 , _u10_u4_n3223 ,_u10_u4_n3222 , _u10_u4_n3221 , _u10_u4_n3220 , _u10_u4_n3219 ,_u10_u4_n3218 , _u10_u4_n3217 , _u10_u4_n3216 , _u10_u4_n3215 ,_u10_u4_n3214 , _u10_u4_n3213 , _u10_u4_n3212 , _u10_u4_n3211 ,_u10_u4_n3210 , _u10_u4_n3209 , _u10_u4_n3208 , _u10_u4_n3207 ,_u10_u4_n3206 , _u10_u4_n3205 , _u10_u4_n3204 , _u10_u4_n3203 ,_u10_u4_n3202 , _u10_u4_n3201 , _u10_u4_n3200 , _u10_u4_n3199 ,_u10_u4_n3198 , _u10_u4_n3197 , _u10_u4_n3196 , _u10_u4_n3195 ,_u10_u4_n3194 , _u10_u4_n3193 , _u10_u4_n3192 , _u10_u4_n3191 ,_u10_u4_n3190 , _u10_u4_n3189 , _u10_u4_n3188 , _u10_u4_n3187 ,_u10_u4_n3186 , _u10_u4_n3185 , _u10_u4_n3184 , _u10_u4_n3183 ,_u10_u4_n3182 , _u10_u4_n3181 , _u10_u4_n3180 , _u10_u4_n3179 ,_u10_u4_n3178 , _u10_u4_n3177 , _u10_u4_n3176 , _u10_u4_n3175 ,_u10_u4_n3174 , _u10_u4_n3173 , _u10_u4_n3172 , _u10_u4_n3171 ,_u10_u4_n3170 , _u10_u4_n3169 , _u10_u4_n3168 , _u10_u4_n3167 ,_u10_u4_n3166 , _u10_u4_n3165 , _u10_u4_n3164 , _u10_u4_n3163 ,_u10_u4_n3162 , _u10_u4_n3161 , _u10_u4_n3160 , _u10_u4_n3159 ,_u10_u4_n3158 , _u10_u4_n3157 , _u10_u4_n3156 , _u10_u4_n3155 ,_u10_u4_n3154 , _u10_u4_n3153 , _u10_u4_n3152 , _u10_u4_n3151 ,_u10_u4_n3150 , _u10_u4_n3149 , _u10_u4_n3148 , _u10_u4_n3147 ,_u10_u4_n3146 , _u10_u4_n3145 , _u10_u4_n3144 , _u10_u4_n3143 ,_u10_u4_n3142 , _u10_u4_n3141 , _u10_u4_n3140 , _u10_u4_n3139 ,_u10_u4_n3138 , _u10_u4_n3137 , _u10_u4_n3136 , _u10_u4_n3135 ,_u10_u4_n3134 , _u10_u4_n3133 , _u10_u4_n3132 , _u10_u4_n3131 ,_u10_u4_n3130 , _u10_u4_n3129 , _u10_u4_n3128 , _u10_u4_n3127 ,_u10_u4_n3126 , _u10_u4_n3125 , _u10_u4_n3124 , _u10_u4_n3123 ,_u10_u4_n3122 , _u10_u4_n3121 , _u10_u4_n3120 , _u10_u4_n3119 ,_u10_u4_n3118 , _u10_u4_n3117 , _u10_u4_n3116 , _u10_u4_n3115 ,_u10_u4_n3114 , _u10_u4_n3113 , _u10_u4_n3112 , _u10_u4_n3111 ,_u10_u4_n3110 , _u10_u4_n3109 , _u10_u4_n3108 , _u10_u4_n3107 ,_u10_u4_n3106 , _u10_u4_n3105 , _u10_u4_n3104 , _u10_u4_n3103 ,_u10_u4_n3102 , _u10_u4_n3101 , _u10_u4_n3100 , _u10_u4_n3099 ,_u10_u4_n3098 , _u10_u4_n3097 , _u10_u4_n3096 , _u10_u4_n3095 ,_u10_u4_n3094 , _u10_u4_n3093 , _u10_u4_n3092 , _u10_u4_n3091 ,_u10_u4_n3090 , _u10_u4_n3089 , _u10_u4_n3088 , _u10_u4_n3087 ,_u10_u4_n3086 , _u10_u4_n3085 , _u10_u4_n3084 , _u10_u4_n3083 ,_u10_u4_n3082 , _u10_u4_n3081 , _u10_u4_n3080 , _u10_u4_n3079 ,_u10_u4_n3078 , _u10_u4_n3077 , _u10_u4_n3076 , _u10_u4_n3075 ,_u10_u4_n3074 , _u10_u4_n3073 , _u10_u4_n3072 , _u10_u4_n3071 ,_u10_u4_n3070 , _u10_u4_n3069 , _u10_u4_n3068 , _u10_u4_n3067 ,_u10_u4_n3066 , _u10_u4_n3065 , _u10_u4_n3064 , _u10_u4_n3063 ,_u10_u4_n3062 , _u10_u4_n3061 , _u10_u4_n3060 , _u10_u4_n3059 ,_u10_u4_n3058 , _u10_u4_n3057 , _u10_u4_n3056 , _u10_u4_n3055 ,_u10_u4_n3054 , _u10_u4_n3053 , _u10_u4_n3052 , _u10_u4_n3051 ,_u10_u4_n3050 , _u10_u4_n3049 , _u10_u4_n3048 , _u10_u4_n3047 ,_u10_u4_n3046 , _u10_u4_n3045 , _u10_u4_n3044 , _u10_u4_n3043 ,_u10_u4_n3042 , _u10_u4_n3041 , _u10_u4_n3040 , _u10_u4_n3039 ,_u10_u4_n3038 , _u10_u4_n3037 , _u10_u4_n3036 , _u10_u4_n3035 ,_u10_u4_n3034 , _u10_u4_n3033 , _u10_u4_n3032 , _u10_u4_n3031 ,_u10_u4_n3030 , _u10_u4_n3029 , _u10_u4_n3028 , _u10_u4_n3027 ,_u10_u4_n3026 , _u10_u4_n3025 , _u10_u4_n3024 , _u10_u4_n3023 ,_u10_u4_n3022 , _u10_u4_n3021 , _u10_u4_n3020 , _u10_u4_n3019 ,_u10_u4_n3018 , _u10_u4_n3017 , _u10_u4_n3016 , _u10_u4_n3015 ,_u10_u4_n3014 , _u10_u4_n3013 , _u10_u4_n3012 , _u10_u4_n3011 ,_u10_u4_n3010 , _u10_u4_n3009 , _u10_u4_n3008 , _u10_u4_n3007 ,_u10_u4_n3006 , _u10_u4_n3005 , _u10_u4_n3004 , _u10_u4_n3003 ,_u10_u4_n3002 , _u10_u4_n3001 , _u10_u4_n3000 , _u10_u4_n2999 ,_u10_u4_n2998 , _u10_u4_n2997 , _u10_u4_n2996 , _u10_u4_n2995 ,_u10_u4_n2994 , _u10_u4_n2993 , _u10_u4_n2992 , _u10_u4_n2991 ,_u10_u4_n2990 , _u10_u4_n2989 , _u10_u4_n2988 , _u10_u4_n2987 ,_u10_u4_n2986 , _u10_u4_n2985 , _u10_u4_n2984 , _u10_u4_n2983 ,_u10_u4_n2982 , _u10_u4_n2981 , _u10_u4_n2980 , _u10_u4_n2979 ,_u10_u4_n2978 , _u10_u4_n2977 , _u10_u4_n2976 , _u10_u4_n2975 ,_u10_u4_n2974 , _u10_u4_n2973 , _u10_u4_n2972 , _u10_u4_n2971 ,_u10_u4_n2970 , _u10_u4_n2969 , _u10_u4_n2968 , _u10_u4_n2967 ,_u10_u4_n2966 , _u10_u4_n2965 , _u10_u4_n2964 , _u10_u4_n2963 ,_u10_u4_n2962 , _u10_u4_n2961 , _u10_u4_n2960 , _u10_u4_n2959 ,_u10_u4_n2958 , _u10_u4_n2957 , _u10_u4_n2956 , _u10_u4_n2955 ,_u10_u4_n2954 , _u10_u4_n2953 , _u10_u4_n2952 , _u10_u4_n2951 ,_u10_u4_n2950 , _u10_u4_n2949 , _u10_u4_n2948 , _u10_u4_n2947 ,_u10_u4_n2946 , _u10_u4_n2945 , _u10_u4_n2944 , _u10_u4_n2943 ,_u10_u4_n2942 , _u10_u4_n2941 , _u10_u4_n2940 , _u10_u4_n2939 ,_u10_u4_n2938 , _u10_u4_n2937 , _u10_u4_n2936 , _u10_u4_n2935 ,_u10_u4_n2934 , _u10_u4_n2933 , _u10_u4_n2932 , _u10_u4_n2931 ,_u10_u4_n2930 , _u10_u4_n2929 , _u10_u4_n2928 , _u10_u4_n2927 ,_u10_u4_n2926 , _u10_u4_n2925 , _u10_u4_n2924 , _u10_u4_n2923 ,_u10_u4_n2922 , _u10_u4_n2921 , _u10_u4_n2920 , _u10_u4_n2919 ,_u10_u4_n2918 , _u10_u4_n2917 , _u10_u4_n2916 , _u10_u4_n2915 ,_u10_u4_n2914 , _u10_u4_n2913 , _u10_u4_n2912 , _u10_u4_n2911 ,_u10_u4_n2910 , _u10_u4_n2909 , _u10_u4_n2908 , _u10_u4_n2907 ,_u10_u4_n2906 , _u10_u4_n2905 , _u10_u4_n2904 , _u10_u4_n2903 ,_u10_u4_n2902 , _u10_u4_n2901 , _u10_u4_n2900 , _u10_u4_n2899 ,_u10_u4_n2898 , _u10_u4_n2897 , _u10_u4_n2896 , _u10_u4_n2895 ,_u10_u4_n2894 , _u10_u4_n2893 , _u10_u4_n2892 , _u10_u4_n2891 ,_u10_u4_n2890 , _u10_u4_n2889 , _u10_u4_n2888 , _u10_u4_n2887 ,_u10_u4_n2886 , _u10_u4_n2885 , _u10_u4_n2884 , _u10_u4_n2883 ,_u10_u4_n2882 , _u10_u4_n2881 , _u10_u4_n2880 , _u10_u4_n2879 ,_u10_u4_n2878 , _u10_u4_n2877 , _u10_u4_n2876 , _u10_u4_n2875 ,_u10_u4_n2874 , _u10_u4_n2873 , _u10_u4_n2872 , _u10_u4_n2871 ,_u10_u4_n2870 , _u10_u4_n2869 , _u10_u4_n2868 , _u10_u4_n2867 ,_u10_u4_n2866 , _u10_u4_n2865 , _u10_u4_n2864 , _u10_u4_n2863 ,_u10_u4_n2862 , _u10_u4_n2861 , _u10_u4_n2860 , _u10_u4_n2859 ,_u10_u4_n2858 , _u10_u4_n2857 , _u10_u4_n2856 , _u10_u4_n2855 ,_u10_u4_n2854 , _u10_u4_n2853 , _u10_u4_n2852 , _u10_u4_n2851 ,_u10_u4_n2850 , _u10_u4_n2849 , _u10_u4_n2848 , _u10_u4_n2847 ,_u10_u4_n2846 , _u10_u4_n2845 , _u10_u4_n2844 , _u10_u4_n2843 ,_u10_u4_n2842 , _u10_u4_n2841 , _u10_u4_n2840 , _u10_u4_n2839 ,_u10_u4_n2838 , _u10_u4_n2837 , _u10_u4_n2836 , _u10_u4_n2835 ,_u10_u4_n2834 , _u10_u4_n2833 , _u10_u4_n2832 , _u10_u4_n2831 ,_u10_u4_n2830 , _u10_u4_n2829 , _u10_u4_n2828 , _u10_u4_n2827 ,_u10_u4_n2826 , _u10_u4_n2825 , _u10_u4_n2824 , _u10_u4_n2823 ,_u10_u4_n2822 , _u10_u4_n2821 , _u10_u4_n2820 , _u10_u4_n2819 ,_u10_u4_n2818 , _u10_u4_n2817 , _u10_u4_n2816 , _u10_u4_n2815 ,_u10_u4_n2814 , _u10_u4_n2813 , _u10_u4_n2812 , _u10_u4_n2811 ,_u10_u4_n2810 , _u10_u4_n2809 , _u10_u4_n2808 , _u10_u4_n2807 ,_u10_u4_n2806 , _u10_u4_n2805 , _u10_u4_n2804 , _u10_u4_n2803 ,_u10_u4_n2802 , _u10_u4_n2801 , _u10_u4_n2800 , _u10_u4_n2799 ,_u10_u4_n2798 , _u10_u4_n2797 , _u10_u4_n2796 , _u10_u4_n2795 ,_u10_u4_n2794 , _u10_u4_n2793 , _u10_u4_n2792 , _u10_u4_n2791 ,_u10_u4_n2790 , _u10_u4_n2789 , _u10_u4_n2788 , _u10_u4_n2787 ,_u10_u4_n2786 , _u10_u4_n2785 , _u10_u4_n2784 , _u10_u4_n2783 ,_u10_u4_n2782 , _u10_u4_n2781 , _u10_u4_n2780 , _u10_u4_n2779 ,_u10_u4_n2778 , _u10_u4_n2777 , _u10_u4_n2776 , _u10_u4_n2775 ,_u10_u4_n2774 , _u10_u4_n2773 , _u10_u4_n2772 , _u10_u4_n2771 ,_u10_u4_n2770 , _u10_u4_n2769 , _u10_u4_n2768 , _u10_u4_n2767 ,_u10_u4_n2766 , _u10_u4_n2765 , _u10_u4_n2764 , _u10_u4_n2763 ,_u10_u4_n2762 , _u10_u4_n2761 , _u10_u4_n2760 , _u10_u4_n2759 ,_u10_u4_n2758 , _u10_u4_n2757 , _u10_u4_n2756 , _u10_u4_n2755 ,_u10_u4_n2754 , _u10_u4_n2753 , _u10_u4_n2752 , _u10_u4_n2751 ,_u10_u4_n2750 , _u10_u4_n2749 , _u10_u4_n2748 , _u10_u4_n2747 ,_u10_u4_n2746 , _u10_u4_n2745 , _u10_u4_n2744 , _u10_u4_n2743 ,_u10_u4_n2742 , _u10_u4_n2741 , _u10_u4_n2740 , _u10_u4_n2739 ,_u10_u4_n2738 , _u10_u4_n2737 , _u10_u4_n2736 , _u10_u4_n2735 ,_u10_u4_n2734 , _u10_u4_n2733 , _u10_u4_n2732 , _u10_u4_n2731 ,_u10_u4_n2730 , _u10_u4_n2729 , _u10_u4_n2728 , _u10_u4_n2727 ,_u10_u4_n2726 , _u10_u4_n2725 , _u10_u4_n2724 , _u10_u4_n2723 ,_u10_u4_n2722 , _u10_u4_n2721 , _u10_u4_n2720 , _u10_u4_n2719 ,_u10_u4_n2718 , _u10_u4_n2717 , _u10_u4_n2716 , _u10_u4_n2715 ,_u10_u4_n2714 , _u10_u4_n2713 , _u10_u4_n2712 , _u10_u4_n2711 ,_u10_u4_n2710 , _u10_u4_n2709 , _u10_u4_n2708 , _u10_u4_n2707 ,_u10_u4_n2706 , _u10_u4_n2705 , _u10_u4_n2704 , _u10_u4_n2703 ,_u10_u4_n2702 , _u10_u4_n2701 , _u10_u4_n2700 , _u10_u4_n2699 ,_u10_u4_n2698 , _u10_u4_n2697 , _u10_u4_n2696 , _u10_u4_n2695 ,_u10_u4_n2694 , _u10_u4_n2693 , _u10_u4_n2692 , _u10_u4_n2691 ,_u10_u4_n2690 , _u10_u4_n2689 , _u10_u4_n2688 , _u10_u4_n2687 ,_u10_u4_n2686 , _u10_u4_n2685 , _u10_u4_n2684 , _u10_u4_n2683 ,_u10_u4_n2682 , _u10_u4_n2681 , _u10_u4_n2680 , _u10_u4_n2679 ,_u10_u4_n2678 , _u10_u4_n2677 , _u10_u4_n2676 , _u10_u4_n2675 ,_u10_u4_n2674 , _u10_u4_n2673 , _u10_u4_n2672 , _u10_u4_n2671 ,_u10_u4_n2670 , _u10_u4_n2669 , _u10_u4_n2668 , _u10_u4_n2667 ,_u10_u4_n2666 , _u10_u4_n2665 , _u10_u4_n2664 , _u10_u4_n2663 ,_u10_u4_n2662 , _u10_u4_n2661 , _u10_u4_n2660 , _u10_u4_n2659 ,_u10_u4_n2658 , _u10_u4_n2657 , _u10_u4_n2656 , _u10_u4_n2655 ,_u10_u4_n2654 , _u10_u4_n2653 , _u10_u4_n2652 , _u10_u4_n2651 ,_u10_u4_n2650 , _u10_u4_n2649 , _u10_u4_n2648 , _u10_u4_n2647 ,_u10_u4_n2646 , _u10_u4_n2645 , _u10_u4_n2644 , _u10_u4_n2643 ,_u10_u4_n2642 , _u10_u4_n2641 , _u10_u4_n2640 , _u10_u4_n2639 ,_u10_u4_n2638 , _u10_u4_n2637 , _u10_u4_n2636 , _u10_u4_n2635 ,_u10_u4_n2634 , _u10_u4_n2633 , _u10_u4_n2632 , _u10_u4_n2631 ,_u10_u4_n2630 , _u10_u4_n2629 , _u10_u4_n2628 , _u10_u4_n2627 ,_u10_u4_n2626 , _u10_u4_n2625 , _u10_u4_n2624 , _u10_u4_n2623 ,_u10_u4_n2622 , _u10_u4_n2621 , _u10_u4_n2620 , _u10_u4_n2619 ,_u10_u4_n2618 , _u10_u4_n2617 , _u10_u4_n2616 , _u10_u4_n2615 ,_u10_u4_n2614 , _u10_u4_n2613 , _u10_u4_n2612 , _u10_u4_n2611 ,_u10_u4_n2610 , _u10_u4_n2609 , _u10_u4_n2608 , _u10_u4_n2607 ,_u10_u4_n2606 , _u10_u4_n2605 , _u10_u4_n2604 , _u10_u4_n2603 ,_u10_u4_n2602 , _u10_u4_n2601 , _u10_u4_n2600 , _u10_u4_n2599 ,_u10_u4_n2598 , _u10_u4_n2597 , _u10_u4_n2596 , _u10_u4_n2595 ,_u10_u4_n2594 , _u10_u4_n2593 , _u10_u4_n2592 , _u10_u4_n2591 ,_u10_u4_n2590 , _u10_u4_n2589 , _u10_u4_n2588 , _u10_u4_n2587 ,_u10_u4_n2586 , _u10_u4_n2585 , _u10_u4_n2584 , _u10_u4_n2583 ,_u10_u4_n2582 , _u10_u4_n2581 , _u10_u4_n2580 , _u10_u4_n2579 ,_u10_u4_n2578 , _u10_u4_n2577 , _u10_u4_n2576 , _u10_u4_n2575 ,_u10_u4_n2574 , _u10_u4_n2573 , _u10_u4_n2572 , _u10_u4_n2571 ,_u10_u4_n2570 , _u10_u4_n2569 , _u10_u4_n2568 , _u10_u4_n2567 ,_u10_u4_n2566 , _u10_u4_n2565 , _u10_u4_n2564 , _u10_u4_n2563 ,_u10_u4_n2562 , _u10_u4_n2561 , _u10_u4_n2560 , _u10_u4_n2559 ,_u10_u4_n2558 , _u10_u4_n2557 , _u10_u4_n2556 , _u10_u4_n2555 ,_u10_u4_n2554 , _u10_u4_n2553 , _u10_u4_n2552 , _u10_u4_n2551 ,_u10_u4_n2550 , _u10_u4_n2549 , _u10_u4_n2548 , _u10_u4_n2547 ,_u10_u4_n2546 , _u10_u4_n2545 , _u10_u4_n2544 , _u10_u4_n2543 ,_u10_u4_n2542 , _u10_u4_n2541 , _u10_u4_n2540 , _u10_u4_n2539 ,_u10_u4_n2538 , _u10_u4_n2537 , _u10_u4_n2536 , _u10_u4_n2535 ,_u10_u4_n2534 , _u10_u4_n2533 , _u10_u4_n2532 , _u10_u4_n2531 ,_u10_u4_n2530 , _u10_u4_n2529 , _u10_u4_n2528 , _u10_u4_n2527 ,_u10_u4_n2526 , _u10_u4_n2525 , _u10_u4_n2524 , _u10_u4_n2523 ,_u10_u4_n2522 , _u10_u4_n2521 , _u10_u4_n2520 , _u10_u4_n2519 ,_u10_u4_n2518 , _u10_u4_n2517 , _u10_u4_n2516 , _u10_u4_n2515 ,_u10_u4_n2514 , _u10_u4_n2513 , _u10_u4_n2512 , _u10_u4_n2511 ,_u10_u4_n2510 , _u10_u4_n2509 , _u10_u4_n2508 , _u10_u4_n2507 ,_u10_u4_n2506 , _u10_u4_n2505 , _u10_u4_n2504 , _u10_u4_n2503 ,_u10_u4_n2502 , _u10_u4_n2501 , _u10_u4_n2500 , _u10_u4_n2499 ,_u10_u4_n2498 , _u10_u4_n2497 , _u10_u4_n2496 , _u10_u4_n2495 ,_u10_u4_n2494 , _u10_u4_n2493 , _u10_u4_n2492 , _u10_u4_n2491 ,_u10_u4_n2490 , _u10_u4_n2489 , _u10_u4_n2488 , _u10_u4_n2487 ,_u10_u4_n2486 , _u10_u4_n2485 , _u10_u4_n2484 , _u10_u4_n2483 ,_u10_u4_n2482 , _u10_u4_n2481 , _u10_u4_n2480 , _u10_u4_n2479 ,_u10_u4_n2478 , _u10_u4_n2477 , _u10_u4_n2476 , _u10_u4_n2475 ,_u10_u4_n2474 , _u10_u4_n2473 , _u10_u4_n2472 , _u10_u4_n2471 ,_u10_u4_n2470 , _u10_u4_n2469 , _u10_u4_n2468 , _u10_u4_n2467 ,_u10_u4_n2466 , _u10_u4_n2465 , _u10_u4_n2464 , _u10_u4_n2463 ,_u10_u4_n2462 , _u10_u4_n2461 , _u10_u4_n2460 , _u10_u4_n2459 ,_u10_u4_n2458 , _u10_u4_n2457 , _u10_u4_n2456 , _u10_u4_n2455 ,_u10_u4_n2454 , _u10_u4_n2453 , _u10_u4_n2452 , _u10_u4_n2451 ,_u10_u4_n2450 , _u10_u4_n2449 , _u10_u4_n2448 , _u10_u4_n2447 ,_u10_u4_n2446 , _u10_u4_n2445 , _u10_u4_n2444 , _u10_u4_n2443 ,_u10_u4_n2442 , _u10_u4_n2441 , _u10_u4_n2440 , _u10_u4_n2439 ,_u10_u4_n2438 , _u10_u4_n2437 , _u10_u4_n2436 , _u10_u4_n2435 ,_u10_u4_n2434 , _u10_u4_n2433 , _u10_u4_n2432 , _u10_u4_n2431 ,_u10_u4_n2430 , _u10_u4_n2429 , _u10_u4_n2428 , _u10_u4_n2427 ,_u10_u4_n2426 , _u10_u4_n2425 , _u10_u4_n2424 , _u10_u4_n2423 ,_u10_u4_n2422 , _u10_u4_n2421 , _u10_u4_n2420 , _u10_u4_n2419 ,_u10_u4_n2418 , _u10_u4_n2417 , _u10_u4_n2416 , _u10_u4_n2415 ,_u10_u4_n2414 , _u10_u4_n2413 , _u10_u4_n2412 , _u10_u4_n2411 ,_u10_u4_n2410 , _u10_u4_n2409 , _u10_u4_n2408 , _u10_u4_n2407 ,_u10_u4_n2406 , _u10_u4_n2405 , _u10_u4_n2404 , _u10_u4_n2403 ,_u10_u4_n2402 , _u10_u4_n2401 , _u10_u4_n2400 , _u10_u4_n2399 ,_u10_u4_n2398 , _u10_u4_n2397 , _u10_u4_n2396 , _u10_u4_n2395 ,_u10_u4_n2394 , _u10_u4_n2393 , _u10_u4_n2392 , _u10_u4_n2391 ,_u10_u4_n2390 , _u10_u4_n2389 , _u10_u4_n2388 , _u10_u4_n2387 ,_u10_u4_n2386 , _u10_u4_n2385 , _u10_u4_n2384 , _u10_u4_n2383 ,_u10_u4_n2382 , _u10_u4_n2381 , _u10_u4_n2380 , _u10_u4_n2379 ,_u10_u4_n2378 , _u10_u4_n2377 , _u10_u4_n2376 , _u10_u4_n2375 ,_u10_u4_n2374 , _u10_u4_n2373 , _u10_u4_n2372 , _u10_u4_n2371 ,_u10_u4_n2370 , _u10_u4_n2369 , _u10_u4_n2368 , _u10_u4_n2367 ,_u10_u4_n2366 , _u10_u4_n2365 , _u10_u4_n2364 , _u10_u4_n2363 ,_u10_u4_n2362 , _u10_u4_n2361 , _u10_u4_n2360 , _u10_u4_n2359 ,_u10_u4_n2358 , _u10_u4_n2357 , _u10_u4_n2356 , _u10_u4_n2355 ,_u10_u4_n2354 , _u10_u4_n2353 , _u10_u4_n2352 , _u10_u4_n2351 ,_u10_u4_n2350 , _u10_u4_n2349 , _u10_u4_n2348 , _u10_u4_n2347 ,_u10_u4_n2346 , _u10_u4_n2345 , _u10_u4_n2344 , _u10_u4_n2343 ,_u10_u4_n2342 , _u10_u4_n2341 , _u10_u4_n2340 , _u10_u4_n2339 ,_u10_u4_n2338 , _u10_u4_n2337 , _u10_u4_n2336 , _u10_u4_n2335 ,_u10_u4_n2334 , _u10_u4_n2333 , _u10_u4_n2332 , _u10_u4_n2331 ,_u10_u4_n2330 , _u10_u4_n2329 , _u10_u4_n2328 , _u10_u4_n2327 ,_u10_u4_n2326 , _u10_u4_n2325 , _u10_u4_n2324 , _u10_u4_n2323 ,_u10_u4_n2322 , _u10_u4_n2321 , _u10_u4_n2320 , _u10_u4_n2319 ,_u10_u4_n2318 , _u10_u4_n2317 , _u10_u4_n2316 , _u10_u4_n2315 ,_u10_u4_n2314 , _u10_u4_n2313 , _u10_u4_n2312 , _u10_u4_n2311 ,_u10_u4_n2310 , _u10_u4_n2309 , _u10_u4_n2308 , _u10_u4_n2307 ,_u10_u4_n2306 , _u10_u4_n2305 , _u10_u4_n2304 , _u10_u4_n2303 ,_u10_u4_n2302 , _u10_u4_n2301 , _u10_u4_n2300 , _u10_u4_n2299 ,_u10_u4_n2298 , _u10_u4_n2297 , _u10_u4_n2296 , _u10_u4_n2295 ,_u10_u4_n2294 , _u10_u4_n2293 , _u10_u4_n2292 , _u10_u4_n2291 ,_u10_u4_n2290 , _u10_u4_n2289 , _u10_u4_n2288 , _u10_u4_n2287 ,_u10_u4_n2286 , _u10_u4_n2285 , _u10_u4_n2284 , _u10_u4_n2283 ,_u10_u4_n2282 , _u10_u4_n2281 , _u10_u4_n2280 , _u10_u4_n2279 ,_u10_u4_n2278 , _u10_u4_n2277 , _u10_u4_n2276 , _u10_u4_n2275 ,_u10_u4_n2274 , _u10_u4_n2273 , _u10_u4_n2272 , _u10_u4_n2271 ,_u10_u4_n2270 , _u10_u4_n2269 , _u10_u4_n2268 , _u10_u4_n2267 ,_u10_u4_n2266 , _u10_u4_n2265 , _u10_u4_n2264 , _u10_u4_n2263 ,_u10_u4_n2262 , _u10_u4_n2261 , _u10_u4_n2260 , _u10_u4_n2259 ,_u10_u4_n2258 , _u10_u4_n2257 , _u10_u4_n2256 , _u10_u4_n2255 ,_u10_u4_n2254 , _u10_u4_n2253 , _u10_u4_n2252 , _u10_u4_n2251 ,_u10_u4_n2250 , _u10_u4_n2249 , _u10_u4_n2248 , _u10_u4_n2247 ,_u10_u4_n2246 , _u10_u4_n2245 , _u10_u4_n2244 , _u10_u4_n2243 ,_u10_u4_n2242 , _u10_u4_n2241 , _u10_u4_n2240 , _u10_u4_n2239 ,_u10_u4_n2238 , _u10_u4_n2237 , _u10_u4_n2236 , _u10_u4_n2235 ,_u10_u4_n2234 , _u10_u4_n2233 , _u10_u4_n2232 , _u10_u4_n2231 ,_u10_u4_n2230 , _u10_u4_n2229 , _u10_u4_n2228 , _u10_u4_n2227 ,_u10_u4_n2226 , _u10_u4_n2225 , _u10_u4_n2224 , _u10_u4_n2223 ,_u10_u4_n2222 , _u10_u4_n2221 , _u10_u4_n2220 , _u10_u4_n2219 ,_u10_u4_n2218 , _u10_u4_n2217 , _u10_u4_n2216 , _u10_u4_n2215 ,_u10_u4_n2214 , _u10_u4_n2213 , _u10_u4_n2212 , _u10_u4_n2211 ,_u10_u4_n2210 , _u10_u4_n2209 , _u10_u4_n2208 , _u10_u4_n2207 ,_u10_u4_n2206 , _u10_u4_n2205 , _u10_u4_n2204 , _u10_u4_n2203 ,_u10_u4_n2202 , _u10_u4_n2201 , _u10_u4_n2200 , _u10_u4_n2199 ,_u10_u4_n2198 , _u10_u4_n2197 , _u10_u4_n2196 , _u10_u4_n2195 ,_u10_u4_n2194 , _u10_u4_n2193 , _u10_u4_n2192 , _u10_u4_n2191 ,_u10_u4_n2190 , _u10_u4_n2189 , _u10_u4_n2188 , _u10_u4_n2187 ,_u10_u4_n2186 , _u10_u4_n2185 , _u10_u4_n2184 , _u10_u4_n2183 ,_u10_u4_n2182 , _u10_u4_n2181 , _u10_u4_n2180 , _u10_u4_n2179 ,_u10_u4_n2178 , _u10_u4_n2177 , _u10_u4_n2176 , _u10_u4_n2175 ,_u10_u4_n2174 , _u10_u4_n2173 , _u10_u4_n2172 , _u10_u4_n2171 ,_u10_u4_n2170 , _u10_u4_n2169 , _u10_u4_n2168 , _u10_u4_n2167 ,_u10_u4_n2166 , _u10_u4_n2165 , _u10_u4_n2164 , _u10_u4_n2163 ,_u10_u4_n2162 , _u10_u4_n2161 , _u10_u4_n2160 , _u10_u4_n2159 ,_u10_u4_n2158 , _u10_u4_n2157 , _u10_u4_n2156 , _u10_u4_n2155 ,_u10_u4_n2154 , _u10_u4_n2153 , _u10_u4_n2152 , _u10_u4_n2151 ,_u10_u4_n2150 , _u10_u4_n2149 , _u10_u4_n2148 , _u10_u4_n2147 ,_u10_u4_n2146 , _u10_u4_n2145 , _u10_u4_n2144 , _u10_u4_n2143 ,_u10_u4_n2142 , _u10_u4_n2141 , _u10_u4_n2140 , _u10_u4_n2139 ,_u10_u4_n2138 , _u10_u4_n2137 , _u10_u4_n2136 , _u10_u4_n2135 ,_u10_u4_n2134 , _u10_u4_n2133 , _u10_u4_n2132 , _u10_u4_n2131 ,_u10_u4_n2130 , _u10_u4_n2129 , _u10_u4_n2128 , _u10_u4_n2127 ,_u10_u4_n2126 , _u10_u4_n2125 , _u10_u4_n2124 , _u10_u4_n2123 ,_u10_u4_n2122 , _u10_u4_n2121 , _u10_u4_n2120 , _u10_u4_n2119 ,_u10_u4_n2118 , _u10_u4_n2117 , _u10_u4_n2116 , _u10_u4_n2115 ,_u10_u4_n2114 , _u10_u4_n2113 , _u10_u4_n2112 , _u10_u4_n2111 ,_u10_u4_n2110 , _u10_u4_n2109 , _u10_u4_n2108 , _u10_u4_n2107 ,_u10_u4_n2106 , _u10_u4_n2105 , _u10_u4_n2104 , _u10_u4_n2103 ,_u10_u4_n2102 , _u10_u4_n2101 , _u10_u4_n2100 , _u10_u4_n2099 ,_u10_u4_n2098 , _u10_u4_n2097 , _u10_u4_n2096 , _u10_u4_n2095 ,_u10_u4_n2094 , _u10_u4_n2093 , _u10_u4_n2092 , _u10_u4_n2091 ,_u10_u4_n2090 , _u10_u4_n2089 , _u10_u4_n2088 , _u10_u4_n2087 ,_u10_u4_n2086 , _u10_u4_n2085 , _u10_u4_n2084 , _u10_u4_n2083 ,_u10_u4_n2082 , _u10_u4_n2081 , _u10_u4_n2080 , _u10_u4_n2079 ,_u10_u4_n2078 , _u10_u4_n2077 , _u10_u4_n2076 , _u10_u4_n2075 ,_u10_u4_n2074 , _u10_u4_n2073 , _u10_u4_n2072 , _u10_u4_n2071 ,_u10_u4_n2070 , _u10_u4_n2069 , _u10_u4_n2068 , _u10_u4_n2067 ,_u10_u4_n2066 , _u10_u4_n2065 , _u10_u4_n2064 , _u10_u4_n2063 ,_u10_u4_n2062 , _u10_u4_n2061 , _u10_u4_n2060 , _u10_u4_n2059 ,_u10_u4_n2058 , _u10_u4_n2057 , _u10_u4_n2056 , _u10_u4_n2055 ,_u10_u4_n2054 , _u10_u4_n2053 , _u10_u4_n2052 , _u10_u4_n2051 ,_u10_u4_n2050 , _u10_u4_n2049 , _u10_u4_n2048 , _u10_u4_n2047 ,_u10_u4_n2046 , _u10_u4_n2045 , _u10_u4_n2044 , _u10_u4_n2043 ,_u10_u4_n2042 , _u10_u4_n2041 , _u10_u4_n2040 , _u10_u4_n2039 ,_u10_u4_n2038 , _u10_u4_n2037 , _u10_u4_n2036 , _u10_u4_n2035 ,_u10_u4_n2034 , _u10_u4_n2033 , _u10_u4_n2032 , _u10_u4_n2031 ,_u10_u4_n2030 , _u10_u4_n2029 , _u10_u4_n2028 , _u10_u4_n2027 ,_u10_u4_n2026 , _u10_u4_n2025 , _u10_u4_n2024 , _u10_u4_n2023 ,_u10_u4_n2022 , _u10_u4_n2021 , _u10_u4_n2020 , _u10_u4_n2019 ,_u10_u4_n2018 , _u10_u4_n2017 , _u10_u4_n2016 , _u10_u4_n2015 ,_u10_u4_n2014 , _u10_u4_n2013 , _u10_u4_n2012 , _u10_u4_n2011 ,_u10_u4_n2010 , _u10_u4_n2009 , _u10_u4_n2008 , _u10_u4_n2007 ,_u10_u4_n2006 , _u10_u4_n2005 , _u10_u4_n2004 , _u10_u4_n2003 ,_u10_u4_n2002 , _u10_u4_n2001 , _u10_u4_n2000 , _u10_u4_n1999 ,_u10_u4_n1998 , _u10_u4_n1997 , _u10_u4_n1996 , _u10_u4_n1995 ,_u10_u4_n1994 , _u10_u4_n1993 , _u10_u4_n1992 , _u10_u4_n1991 ,_u10_u4_n1990 , _u10_u4_n1989 , _u10_u4_n1988 , _u10_u4_n1987 ,_u10_u4_n1986 , _u10_u4_n1985 , _u10_u4_n1984 , _u10_u4_n1983 ,_u10_u4_n1982 , _u10_u4_n1981 , _u10_u4_n1980 , _u10_u4_n1979 ,_u10_u4_n1978 , _u10_u4_n1977 , _u10_u4_n1976 , _u10_u4_n1975 ,_u10_u4_n1974 , _u10_u4_n1973 , _u10_u4_n1972 , _u10_u4_n1971 ,_u10_u4_n1970 , _u10_u4_n1969 , _u10_u4_n1968 , _u10_u4_n1967 ,_u10_u4_n1966 , _u10_u4_n1965 , _u10_u4_n1964 , _u10_u4_n1963 ,_u10_u4_n1962 , _u10_u4_n1961 , _u10_u4_n1960 , _u10_u4_n1959 ,_u10_u4_n1958 , _u10_u4_n1957 , _u10_u4_n1956 , _u10_u4_n1955 ,_u10_u4_n1954 , _u10_u4_n1953 , _u10_u4_n1952 , _u10_u4_n1951 ,_u10_u4_n1950 , _u10_u4_n1949 , _u10_u4_n1948 , _u10_u4_n1947 ,_u10_u4_n1946 , _u10_u4_n1945 , _u10_u4_n1944 , _u10_u4_n1943 ,_u10_u4_n1942 , _u10_u4_n1941 , _u10_u4_n1940 , _u10_u4_n1939 ,_u10_u4_n1938 , _u10_u4_n1937 , _u10_u4_n1936 , _u10_u4_n1935 ,_u10_u4_n1934 , _u10_u4_n1933 , _u10_u4_n1932 , _u10_u4_n1931 ,_u10_u4_n1930 , _u10_u4_n1929 , _u10_u4_n1928 , _u10_u4_n1927 ,_u10_u4_n1926 , _u10_u4_n1925 , _u10_u4_n1924 , _u10_u4_n1923 ,_u10_u4_n1922 , _u10_u4_n1921 , _u10_u4_n1920 , _u10_u4_n1919 ,_u10_u4_n1918 , _u10_u4_n1917 , _u10_u4_n1916 , _u10_u4_n1915 ,_u10_u4_n1914 , _u10_u4_n1913 , _u10_u4_n1912 , _u10_u4_n1911 ,_u10_u4_n1910 , _u10_u4_n1909 , _u10_u4_n1908 , _u10_u4_n1907 ,_u10_u4_n1906 , _u10_u4_n1905 , _u10_u4_n1904 , _u10_u4_n1903 ,_u10_u4_n1902 , _u10_u4_n1901 , _u10_u4_n1900 , _u10_u4_n1899 ,_u10_u4_n1898 , _u10_u4_n1897 , _u10_u4_n1896 , _u10_u4_n1895 ,_u10_u4_n1894 , _u10_u4_n1893 , _u10_u4_n1892 , _u10_u4_n1891 ,_u10_u4_n1890 , _u10_u4_n1889 , _u10_u4_n1888 , _u10_u4_n1887 ,_u10_u4_n1886 , _u10_u4_n1885 , _u10_u4_n1884 , _u10_u4_n1883 ,_u10_u4_n1882 , _u10_u4_n1881 , _u10_u4_n1880 , _u10_u4_n1879 ,_u10_u4_n1878 , _u10_u4_n1877 , _u10_u4_n1876 , _u10_u4_n1875 ,_u10_u4_n1874 , _u10_u4_n1873 , _u10_u4_n1872 , _u10_u4_n1871 ,_u10_u4_n1870 , _u10_u4_n1869 , _u10_u4_n1868 , _u10_u4_n1867 ,_u10_u4_n1866 , _u10_u4_n1865 , _u10_u4_n1864 , _u10_u4_n1863 ,_u10_u4_n1862 , _u10_u4_n1861 , _u10_u4_n1860 , _u10_u4_n1859 ,_u10_u4_n1858 , _u10_u4_n1857 , _u10_u4_n1856 , _u10_u4_n1855 ,_u10_u4_n1854 , _u10_u4_n1853 , _u10_u4_n1852 , _u10_u4_n1851 ,_u10_u4_n1850 , _u10_u4_n1849 , _u10_u4_n1848 , _u10_u4_n1847 ,_u10_u4_n1846 , _u10_u4_n1845 , _u10_u4_n1844 , _u10_u4_n1843 ,_u10_u4_n1842 , _u10_u4_n1841 , _u10_u4_n1840 , _u10_u4_n1839 ,_u10_u4_n1838 , _u10_u4_n1837 , _u10_u4_n1836 , _u10_u4_n1835 ,_u10_u4_n1834 , _u10_u4_n1833 , _u10_u4_n1832 , _u10_u4_n1831 ,_u10_u4_n1830 , _u10_u4_n1829 , _u10_u4_n1828 , _u10_u4_n1827 ,_u10_u4_n1826 , _u10_u4_n1825 , _u10_u4_n1824 , _u10_u4_n1823 ,_u10_u4_n1822 , _u10_u4_n1821 , _u10_u4_n1820 , _u10_u4_n1819 ,_u10_u4_n1818 , _u10_u4_n1817 , _u10_u4_n1816 , _u10_u4_n1815 ,_u10_u4_n1814 , _u10_u4_n1813 , _u10_u4_n1812 , _u10_u4_n1811 ,_u10_u4_n1810 , _u10_u4_n1809 , _u10_u4_n1808 , _u10_u5_n3416 ,_u10_u5_n3415 , _u10_u5_n3414 , _u10_u5_n3413 , _u10_u5_n3412 ,_u10_u5_n3411 , _u10_u5_n3410 , _u10_u5_n3409 , _u10_u5_n3408 ,_u10_u5_n3407 , _u10_u5_n3406 , _u10_u5_n3405 , _u10_u5_n3404 ,_u10_u5_n3403 , _u10_u5_n3402 , _u10_u5_n3401 , _u10_u5_n3400 ,_u10_u5_n3399 , _u10_u5_n3398 , _u10_u5_n3397 , _u10_u5_n3396 ,_u10_u5_n3395 , _u10_u5_n3394 , _u10_u5_n3393 , _u10_u5_n3392 ,_u10_u5_n3391 , _u10_u5_n3390 , _u10_u5_n3389 , _u10_u5_n3388 ,_u10_u5_n3387 , _u10_u5_n3386 , _u10_u5_n3385 , _u10_u5_n3384 ,_u10_u5_n3383 , _u10_u5_n3382 , _u10_u5_n3381 , _u10_u5_n3380 ,_u10_u5_n3379 , _u10_u5_n3378 , _u10_u5_n3377 , _u10_u5_n3376 ,_u10_u5_n3375 , _u10_u5_n3374 , _u10_u5_n3373 , _u10_u5_n3372 ,_u10_u5_n3371 , _u10_u5_n3370 , _u10_u5_n3369 , _u10_u5_n3368 ,_u10_u5_n3367 , _u10_u5_n3366 , _u10_u5_n3365 , _u10_u5_n3364 ,_u10_u5_n3363 , _u10_u5_n3362 , _u10_u5_n3361 , _u10_u5_n3360 ,_u10_u5_n3359 , _u10_u5_n3358 , _u10_u5_n3357 , _u10_u5_n3356 ,_u10_u5_n3355 , _u10_u5_n3354 , _u10_u5_n3353 , _u10_u5_n3352 ,_u10_u5_n3351 , _u10_u5_n3350 , _u10_u5_n3349 , _u10_u5_n3348 ,_u10_u5_n3347 , _u10_u5_n3346 , _u10_u5_n3345 , _u10_u5_n3344 ,_u10_u5_n3343 , _u10_u5_n3342 , _u10_u5_n3341 , _u10_u5_n3340 ,_u10_u5_n3339 , _u10_u5_n3338 , _u10_u5_n3337 , _u10_u5_n3336 ,_u10_u5_n3335 , _u10_u5_n3334 , _u10_u5_n3333 , _u10_u5_n3332 ,_u10_u5_n3331 , _u10_u5_n3330 , _u10_u5_n3329 , _u10_u5_n3328 ,_u10_u5_n3327 , _u10_u5_n3326 , _u10_u5_n3325 , _u10_u5_n3324 ,_u10_u5_n3323 , _u10_u5_n3322 , _u10_u5_n3321 , _u10_u5_n3320 ,_u10_u5_n3319 , _u10_u5_n3318 , _u10_u5_n3317 , _u10_u5_n3316 ,_u10_u5_n3315 , _u10_u5_n3314 , _u10_u5_n3313 , _u10_u5_n3312 ,_u10_u5_n3311 , _u10_u5_n3310 , _u10_u5_n3309 , _u10_u5_n3308 ,_u10_u5_n3307 , _u10_u5_n3306 , _u10_u5_n3305 , _u10_u5_n3304 ,_u10_u5_n3303 , _u10_u5_n3302 , _u10_u5_n3301 , _u10_u5_n3300 ,_u10_u5_n3299 , _u10_u5_n3298 , _u10_u5_n3297 , _u10_u5_n3296 ,_u10_u5_n3295 , _u10_u5_n3294 , _u10_u5_n3293 , _u10_u5_n3292 ,_u10_u5_n3291 , _u10_u5_n3290 , _u10_u5_n3289 , _u10_u5_n3288 ,_u10_u5_n3287 , _u10_u5_n3286 , _u10_u5_n3285 , _u10_u5_n3284 ,_u10_u5_n3283 , _u10_u5_n3282 , _u10_u5_n3281 , _u10_u5_n3280 ,_u10_u5_n3279 , _u10_u5_n3278 , _u10_u5_n3277 , _u10_u5_n3276 ,_u10_u5_n3275 , _u10_u5_n3274 , _u10_u5_n3273 , _u10_u5_n3272 ,_u10_u5_n3271 , _u10_u5_n3270 , _u10_u5_n3269 , _u10_u5_n3268 ,_u10_u5_n3267 , _u10_u5_n3266 , _u10_u5_n3265 , _u10_u5_n3264 ,_u10_u5_n3263 , _u10_u5_n3262 , _u10_u5_n3261 , _u10_u5_n3260 ,_u10_u5_n3259 , _u10_u5_n3258 , _u10_u5_n3257 , _u10_u5_n3256 ,_u10_u5_n3255 , _u10_u5_n3254 , _u10_u5_n3253 , _u10_u5_n3252 ,_u10_u5_n3251 , _u10_u5_n3250 , _u10_u5_n3249 , _u10_u5_n3248 ,_u10_u5_n3247 , _u10_u5_n3246 , _u10_u5_n3245 , _u10_u5_n3244 ,_u10_u5_n3243 , _u10_u5_n3242 , _u10_u5_n3241 , _u10_u5_n3240 ,_u10_u5_n3239 , _u10_u5_n3238 , _u10_u5_n3237 , _u10_u5_n3236 ,_u10_u5_n3235 , _u10_u5_n3234 , _u10_u5_n3233 , _u10_u5_n3232 ,_u10_u5_n3231 , _u10_u5_n3230 , _u10_u5_n3229 , _u10_u5_n3228 ,_u10_u5_n3227 , _u10_u5_n3226 , _u10_u5_n3225 , _u10_u5_n3224 ,_u10_u5_n3223 , _u10_u5_n3222 , _u10_u5_n3221 , _u10_u5_n3220 ,_u10_u5_n3219 , _u10_u5_n3218 , _u10_u5_n3217 , _u10_u5_n3216 ,_u10_u5_n3215 , _u10_u5_n3214 , _u10_u5_n3213 , _u10_u5_n3212 ,_u10_u5_n3211 , _u10_u5_n3210 , _u10_u5_n3209 , _u10_u5_n3208 ,_u10_u5_n3207 , _u10_u5_n3206 , _u10_u5_n3205 , _u10_u5_n3204 ,_u10_u5_n3203 , _u10_u5_n3202 , _u10_u5_n3201 , _u10_u5_n3200 ,_u10_u5_n3199 , _u10_u5_n3198 , _u10_u5_n3197 , _u10_u5_n3196 ,_u10_u5_n3195 , _u10_u5_n3194 , _u10_u5_n3193 , _u10_u5_n3192 ,_u10_u5_n3191 , _u10_u5_n3190 , _u10_u5_n3189 , _u10_u5_n3188 ,_u10_u5_n3187 , _u10_u5_n3186 , _u10_u5_n3185 , _u10_u5_n3184 ,_u10_u5_n3183 , _u10_u5_n3182 , _u10_u5_n3181 , _u10_u5_n3180 ,_u10_u5_n3179 , _u10_u5_n3178 , _u10_u5_n3177 , _u10_u5_n3176 ,_u10_u5_n3175 , _u10_u5_n3174 , _u10_u5_n3173 , _u10_u5_n3172 ,_u10_u5_n3171 , _u10_u5_n3170 , _u10_u5_n3169 , _u10_u5_n3168 ,_u10_u5_n3167 , _u10_u5_n3166 , _u10_u5_n3165 , _u10_u5_n3164 ,_u10_u5_n3163 , _u10_u5_n3162 , _u10_u5_n3161 , _u10_u5_n3160 ,_u10_u5_n3159 , _u10_u5_n3158 , _u10_u5_n3157 , _u10_u5_n3156 ,_u10_u5_n3155 , _u10_u5_n3154 , _u10_u5_n3153 , _u10_u5_n3152 ,_u10_u5_n3151 , _u10_u5_n3150 , _u10_u5_n3149 , _u10_u5_n3148 ,_u10_u5_n3147 , _u10_u5_n3146 , _u10_u5_n3145 , _u10_u5_n3144 ,_u10_u5_n3143 , _u10_u5_n3142 , _u10_u5_n3141 , _u10_u5_n3140 ,_u10_u5_n3139 , _u10_u5_n3138 , _u10_u5_n3137 , _u10_u5_n3136 ,_u10_u5_n3135 , _u10_u5_n3134 , _u10_u5_n3133 , _u10_u5_n3132 ,_u10_u5_n3131 , _u10_u5_n3130 , _u10_u5_n3129 , _u10_u5_n3128 ,_u10_u5_n3127 , _u10_u5_n3126 , _u10_u5_n3125 , _u10_u5_n3124 ,_u10_u5_n3123 , _u10_u5_n3122 , _u10_u5_n3121 , _u10_u5_n3120 ,_u10_u5_n3119 , _u10_u5_n3118 , _u10_u5_n3117 , _u10_u5_n3116 ,_u10_u5_n3115 , _u10_u5_n3114 , _u10_u5_n3113 , _u10_u5_n3112 ,_u10_u5_n3111 , _u10_u5_n3110 , _u10_u5_n3109 , _u10_u5_n3108 ,_u10_u5_n3107 , _u10_u5_n3106 , _u10_u5_n3105 , _u10_u5_n3104 ,_u10_u5_n3103 , _u10_u5_n3102 , _u10_u5_n3101 , _u10_u5_n3100 ,_u10_u5_n3099 , _u10_u5_n3098 , _u10_u5_n3097 , _u10_u5_n3096 ,_u10_u5_n3095 , _u10_u5_n3094 , _u10_u5_n3093 , _u10_u5_n3092 ,_u10_u5_n3091 , _u10_u5_n3090 , _u10_u5_n3089 , _u10_u5_n3088 ,_u10_u5_n3087 , _u10_u5_n3086 , _u10_u5_n3085 , _u10_u5_n3084 ,_u10_u5_n3083 , _u10_u5_n3082 , _u10_u5_n3081 , _u10_u5_n3080 ,_u10_u5_n3079 , _u10_u5_n3078 , _u10_u5_n3077 , _u10_u5_n3076 ,_u10_u5_n3075 , _u10_u5_n3074 , _u10_u5_n3073 , _u10_u5_n3072 ,_u10_u5_n3071 , _u10_u5_n3070 , _u10_u5_n3069 , _u10_u5_n3068 ,_u10_u5_n3067 , _u10_u5_n3066 , _u10_u5_n3065 , _u10_u5_n3064 ,_u10_u5_n3063 , _u10_u5_n3062 , _u10_u5_n3061 , _u10_u5_n3060 ,_u10_u5_n3059 , _u10_u5_n3058 , _u10_u5_n3057 , _u10_u5_n3056 ,_u10_u5_n3055 , _u10_u5_n3054 , _u10_u5_n3053 , _u10_u5_n3052 ,_u10_u5_n3051 , _u10_u5_n3050 , _u10_u5_n3049 , _u10_u5_n3048 ,_u10_u5_n3047 , _u10_u5_n3046 , _u10_u5_n3045 , _u10_u5_n3044 ,_u10_u5_n3043 , _u10_u5_n3042 , _u10_u5_n3041 , _u10_u5_n3040 ,_u10_u5_n3039 , _u10_u5_n3038 , _u10_u5_n3037 , _u10_u5_n3036 ,_u10_u5_n3035 , _u10_u5_n3034 , _u10_u5_n3033 , _u10_u5_n3032 ,_u10_u5_n3031 , _u10_u5_n3030 , _u10_u5_n3029 , _u10_u5_n3028 ,_u10_u5_n3027 , _u10_u5_n3026 , _u10_u5_n3025 , _u10_u5_n3024 ,_u10_u5_n3023 , _u10_u5_n3022 , _u10_u5_n3021 , _u10_u5_n3020 ,_u10_u5_n3019 , _u10_u5_n3018 , _u10_u5_n3017 , _u10_u5_n3016 ,_u10_u5_n3015 , _u10_u5_n3014 , _u10_u5_n3013 , _u10_u5_n3012 ,_u10_u5_n3011 , _u10_u5_n3010 , _u10_u5_n3009 , _u10_u5_n3008 ,_u10_u5_n3007 , _u10_u5_n3006 , _u10_u5_n3005 , _u10_u5_n3004 ,_u10_u5_n3003 , _u10_u5_n3002 , _u10_u5_n3001 , _u10_u5_n3000 ,_u10_u5_n2999 , _u10_u5_n2998 , _u10_u5_n2997 , _u10_u5_n2996 ,_u10_u5_n2995 , _u10_u5_n2994 , _u10_u5_n2993 , _u10_u5_n2992 ,_u10_u5_n2991 , _u10_u5_n2990 , _u10_u5_n2989 , _u10_u5_n2988 ,_u10_u5_n2987 , _u10_u5_n2986 , _u10_u5_n2985 , _u10_u5_n2984 ,_u10_u5_n2983 , _u10_u5_n2982 , _u10_u5_n2981 , _u10_u5_n2980 ,_u10_u5_n2979 , _u10_u5_n2978 , _u10_u5_n2977 , _u10_u5_n2976 ,_u10_u5_n2975 , _u10_u5_n2974 , _u10_u5_n2973 , _u10_u5_n2972 ,_u10_u5_n2971 , _u10_u5_n2970 , _u10_u5_n2969 , _u10_u5_n2968 ,_u10_u5_n2967 , _u10_u5_n2966 , _u10_u5_n2965 , _u10_u5_n2964 ,_u10_u5_n2963 , _u10_u5_n2962 , _u10_u5_n2961 , _u10_u5_n2960 ,_u10_u5_n2959 , _u10_u5_n2958 , _u10_u5_n2957 , _u10_u5_n2956 ,_u10_u5_n2955 , _u10_u5_n2954 , _u10_u5_n2953 , _u10_u5_n2952 ,_u10_u5_n2951 , _u10_u5_n2950 , _u10_u5_n2949 , _u10_u5_n2948 ,_u10_u5_n2947 , _u10_u5_n2946 , _u10_u5_n2945 , _u10_u5_n2944 ,_u10_u5_n2943 , _u10_u5_n2942 , _u10_u5_n2941 , _u10_u5_n2940 ,_u10_u5_n2939 , _u10_u5_n2938 , _u10_u5_n2937 , _u10_u5_n2936 ,_u10_u5_n2935 , _u10_u5_n2934 , _u10_u5_n2933 , _u10_u5_n2932 ,_u10_u5_n2931 , _u10_u5_n2930 , _u10_u5_n2929 , _u10_u5_n2928 ,_u10_u5_n2927 , _u10_u5_n2926 , _u10_u5_n2925 , _u10_u5_n2924 ,_u10_u5_n2923 , _u10_u5_n2922 , _u10_u5_n2921 , _u10_u5_n2920 ,_u10_u5_n2919 , _u10_u5_n2918 , _u10_u5_n2917 , _u10_u5_n2916 ,_u10_u5_n2915 , _u10_u5_n2914 , _u10_u5_n2913 , _u10_u5_n2912 ,_u10_u5_n2911 , _u10_u5_n2910 , _u10_u5_n2909 , _u10_u5_n2908 ,_u10_u5_n2907 , _u10_u5_n2906 , _u10_u5_n2905 , _u10_u5_n2904 ,_u10_u5_n2903 , _u10_u5_n2902 , _u10_u5_n2901 , _u10_u5_n2900 ,_u10_u5_n2899 , _u10_u5_n2898 , _u10_u5_n2897 , _u10_u5_n2896 ,_u10_u5_n2895 , _u10_u5_n2894 , _u10_u5_n2893 , _u10_u5_n2892 ,_u10_u5_n2891 , _u10_u5_n2890 , _u10_u5_n2889 , _u10_u5_n2888 ,_u10_u5_n2887 , _u10_u5_n2886 , _u10_u5_n2885 , _u10_u5_n2884 ,_u10_u5_n2883 , _u10_u5_n2882 , _u10_u5_n2881 , _u10_u5_n2880 ,_u10_u5_n2879 , _u10_u5_n2878 , _u10_u5_n2877 , _u10_u5_n2876 ,_u10_u5_n2875 , _u10_u5_n2874 , _u10_u5_n2873 , _u10_u5_n2872 ,_u10_u5_n2871 , _u10_u5_n2870 , _u10_u5_n2869 , _u10_u5_n2868 ,_u10_u5_n2867 , _u10_u5_n2866 , _u10_u5_n2865 , _u10_u5_n2864 ,_u10_u5_n2863 , _u10_u5_n2862 , _u10_u5_n2861 , _u10_u5_n2860 ,_u10_u5_n2859 , _u10_u5_n2858 , _u10_u5_n2857 , _u10_u5_n2856 ,_u10_u5_n2855 , _u10_u5_n2854 , _u10_u5_n2853 , _u10_u5_n2852 ,_u10_u5_n2851 , _u10_u5_n2850 , _u10_u5_n2849 , _u10_u5_n2848 ,_u10_u5_n2847 , _u10_u5_n2846 , _u10_u5_n2845 , _u10_u5_n2844 ,_u10_u5_n2843 , _u10_u5_n2842 , _u10_u5_n2841 , _u10_u5_n2840 ,_u10_u5_n2839 , _u10_u5_n2838 , _u10_u5_n2837 , _u10_u5_n2836 ,_u10_u5_n2835 , _u10_u5_n2834 , _u10_u5_n2833 , _u10_u5_n2832 ,_u10_u5_n2831 , _u10_u5_n2830 , _u10_u5_n2829 , _u10_u5_n2828 ,_u10_u5_n2827 , _u10_u5_n2826 , _u10_u5_n2825 , _u10_u5_n2824 ,_u10_u5_n2823 , _u10_u5_n2822 , _u10_u5_n2821 , _u10_u5_n2820 ,_u10_u5_n2819 , _u10_u5_n2818 , _u10_u5_n2817 , _u10_u5_n2816 ,_u10_u5_n2815 , _u10_u5_n2814 , _u10_u5_n2813 , _u10_u5_n2812 ,_u10_u5_n2811 , _u10_u5_n2810 , _u10_u5_n2809 , _u10_u5_n2808 ,_u10_u5_n2807 , _u10_u5_n2806 , _u10_u5_n2805 , _u10_u5_n2804 ,_u10_u5_n2803 , _u10_u5_n2802 , _u10_u5_n2801 , _u10_u5_n2800 ,_u10_u5_n2799 , _u10_u5_n2798 , _u10_u5_n2797 , _u10_u5_n2796 ,_u10_u5_n2795 , _u10_u5_n2794 , _u10_u5_n2793 , _u10_u5_n2792 ,_u10_u5_n2791 , _u10_u5_n2790 , _u10_u5_n2789 , _u10_u5_n2788 ,_u10_u5_n2787 , _u10_u5_n2786 , _u10_u5_n2785 , _u10_u5_n2784 ,_u10_u5_n2783 , _u10_u5_n2782 , _u10_u5_n2781 , _u10_u5_n2780 ,_u10_u5_n2779 , _u10_u5_n2778 , _u10_u5_n2777 , _u10_u5_n2776 ,_u10_u5_n2775 , _u10_u5_n2774 , _u10_u5_n2773 , _u10_u5_n2772 ,_u10_u5_n2771 , _u10_u5_n2770 , _u10_u5_n2769 , _u10_u5_n2768 ,_u10_u5_n2767 , _u10_u5_n2766 , _u10_u5_n2765 , _u10_u5_n2764 ,_u10_u5_n2763 , _u10_u5_n2762 , _u10_u5_n2761 , _u10_u5_n2760 ,_u10_u5_n2759 , _u10_u5_n2758 , _u10_u5_n2757 , _u10_u5_n2756 ,_u10_u5_n2755 , _u10_u5_n2754 , _u10_u5_n2753 , _u10_u5_n2752 ,_u10_u5_n2751 , _u10_u5_n2750 , _u10_u5_n2749 , _u10_u5_n2748 ,_u10_u5_n2747 , _u10_u5_n2746 , _u10_u5_n2745 , _u10_u5_n2744 ,_u10_u5_n2743 , _u10_u5_n2742 , _u10_u5_n2741 , _u10_u5_n2740 ,_u10_u5_n2739 , _u10_u5_n2738 , _u10_u5_n2737 , _u10_u5_n2736 ,_u10_u5_n2735 , _u10_u5_n2734 , _u10_u5_n2733 , _u10_u5_n2732 ,_u10_u5_n2731 , _u10_u5_n2730 , _u10_u5_n2729 , _u10_u5_n2728 ,_u10_u5_n2727 , _u10_u5_n2726 , _u10_u5_n2725 , _u10_u5_n2724 ,_u10_u5_n2723 , _u10_u5_n2722 , _u10_u5_n2721 , _u10_u5_n2720 ,_u10_u5_n2719 , _u10_u5_n2718 , _u10_u5_n2717 , _u10_u5_n2716 ,_u10_u5_n2715 , _u10_u5_n2714 , _u10_u5_n2713 , _u10_u5_n2712 ,_u10_u5_n2711 , _u10_u5_n2710 , _u10_u5_n2709 , _u10_u5_n2708 ,_u10_u5_n2707 , _u10_u5_n2706 , _u10_u5_n2705 , _u10_u5_n2704 ,_u10_u5_n2703 , _u10_u5_n2702 , _u10_u5_n2701 , _u10_u5_n2700 ,_u10_u5_n2699 , _u10_u5_n2698 , _u10_u5_n2697 , _u10_u5_n2696 ,_u10_u5_n2695 , _u10_u5_n2694 , _u10_u5_n2693 , _u10_u5_n2692 ,_u10_u5_n2691 , _u10_u5_n2690 , _u10_u5_n2689 , _u10_u5_n2688 ,_u10_u5_n2687 , _u10_u5_n2686 , _u10_u5_n2685 , _u10_u5_n2684 ,_u10_u5_n2683 , _u10_u5_n2682 , _u10_u5_n2681 , _u10_u5_n2680 ,_u10_u5_n2679 , _u10_u5_n2678 , _u10_u5_n2677 , _u10_u5_n2676 ,_u10_u5_n2675 , _u10_u5_n2674 , _u10_u5_n2673 , _u10_u5_n2672 ,_u10_u5_n2671 , _u10_u5_n2670 , _u10_u5_n2669 , _u10_u5_n2668 ,_u10_u5_n2667 , _u10_u5_n2666 , _u10_u5_n2665 , _u10_u5_n2664 ,_u10_u5_n2663 , _u10_u5_n2662 , _u10_u5_n2661 , _u10_u5_n2660 ,_u10_u5_n2659 , _u10_u5_n2658 , _u10_u5_n2657 , _u10_u5_n2656 ,_u10_u5_n2655 , _u10_u5_n2654 , _u10_u5_n2653 , _u10_u5_n2652 ,_u10_u5_n2651 , _u10_u5_n2650 , _u10_u5_n2649 , _u10_u5_n2648 ,_u10_u5_n2647 , _u10_u5_n2646 , _u10_u5_n2645 , _u10_u5_n2644 ,_u10_u5_n2643 , _u10_u5_n2642 , _u10_u5_n2641 , _u10_u5_n2640 ,_u10_u5_n2639 , _u10_u5_n2638 , _u10_u5_n2637 , _u10_u5_n2636 ,_u10_u5_n2635 , _u10_u5_n2634 , _u10_u5_n2633 , _u10_u5_n2632 ,_u10_u5_n2631 , _u10_u5_n2630 , _u10_u5_n2629 , _u10_u5_n2628 ,_u10_u5_n2627 , _u10_u5_n2626 , _u10_u5_n2625 , _u10_u5_n2624 ,_u10_u5_n2623 , _u10_u5_n2622 , _u10_u5_n2621 , _u10_u5_n2620 ,_u10_u5_n2619 , _u10_u5_n2618 , _u10_u5_n2617 , _u10_u5_n2616 ,_u10_u5_n2615 , _u10_u5_n2614 , _u10_u5_n2613 , _u10_u5_n2612 ,_u10_u5_n2611 , _u10_u5_n2610 , _u10_u5_n2609 , _u10_u5_n2608 ,_u10_u5_n2607 , _u10_u5_n2606 , _u10_u5_n2605 , _u10_u5_n2604 ,_u10_u5_n2603 , _u10_u5_n2602 , _u10_u5_n2601 , _u10_u5_n2600 ,_u10_u5_n2599 , _u10_u5_n2598 , _u10_u5_n2597 , _u10_u5_n2596 ,_u10_u5_n2595 , _u10_u5_n2594 , _u10_u5_n2593 , _u10_u5_n2592 ,_u10_u5_n2591 , _u10_u5_n2590 , _u10_u5_n2589 , _u10_u5_n2588 ,_u10_u5_n2587 , _u10_u5_n2586 , _u10_u5_n2585 , _u10_u5_n2584 ,_u10_u5_n2583 , _u10_u5_n2582 , _u10_u5_n2581 , _u10_u5_n2580 ,_u10_u5_n2579 , _u10_u5_n2578 , _u10_u5_n2577 , _u10_u5_n2576 ,_u10_u5_n2575 , _u10_u5_n2574 , _u10_u5_n2573 , _u10_u5_n2572 ,_u10_u5_n2571 , _u10_u5_n2570 , _u10_u5_n2569 , _u10_u5_n2568 ,_u10_u5_n2567 , _u10_u5_n2566 , _u10_u5_n2565 , _u10_u5_n2564 ,_u10_u5_n2563 , _u10_u5_n2562 , _u10_u5_n2561 , _u10_u5_n2560 ,_u10_u5_n2559 , _u10_u5_n2558 , _u10_u5_n2557 , _u10_u5_n2556 ,_u10_u5_n2555 , _u10_u5_n2554 , _u10_u5_n2553 , _u10_u5_n2552 ,_u10_u5_n2551 , _u10_u5_n2550 , _u10_u5_n2549 , _u10_u5_n2548 ,_u10_u5_n2547 , _u10_u5_n2546 , _u10_u5_n2545 , _u10_u5_n2544 ,_u10_u5_n2543 , _u10_u5_n2542 , _u10_u5_n2541 , _u10_u5_n2540 ,_u10_u5_n2539 , _u10_u5_n2538 , _u10_u5_n2537 , _u10_u5_n2536 ,_u10_u5_n2535 , _u10_u5_n2534 , _u10_u5_n2533 , _u10_u5_n2532 ,_u10_u5_n2531 , _u10_u5_n2530 , _u10_u5_n2529 , _u10_u5_n2528 ,_u10_u5_n2527 , _u10_u5_n2526 , _u10_u5_n2525 , _u10_u5_n2524 ,_u10_u5_n2523 , _u10_u5_n2522 , _u10_u5_n2521 , _u10_u5_n2520 ,_u10_u5_n2519 , _u10_u5_n2518 , _u10_u5_n2517 , _u10_u5_n2516 ,_u10_u5_n2515 , _u10_u5_n2514 , _u10_u5_n2513 , _u10_u5_n2512 ,_u10_u5_n2511 , _u10_u5_n2510 , _u10_u5_n2509 , _u10_u5_n2508 ,_u10_u5_n2507 , _u10_u5_n2506 , _u10_u5_n2505 , _u10_u5_n2504 ,_u10_u5_n2503 , _u10_u5_n2502 , _u10_u5_n2501 , _u10_u5_n2500 ,_u10_u5_n2499 , _u10_u5_n2498 , _u10_u5_n2497 , _u10_u5_n2496 ,_u10_u5_n2495 , _u10_u5_n2494 , _u10_u5_n2493 , _u10_u5_n2492 ,_u10_u5_n2491 , _u10_u5_n2490 , _u10_u5_n2489 , _u10_u5_n2488 ,_u10_u5_n2487 , _u10_u5_n2486 , _u10_u5_n2485 , _u10_u5_n2484 ,_u10_u5_n2483 , _u10_u5_n2482 , _u10_u5_n2481 , _u10_u5_n2480 ,_u10_u5_n2479 , _u10_u5_n2478 , _u10_u5_n2477 , _u10_u5_n2476 ,_u10_u5_n2475 , _u10_u5_n2474 , _u10_u5_n2473 , _u10_u5_n2472 ,_u10_u5_n2471 , _u10_u5_n2470 , _u10_u5_n2469 , _u10_u5_n2468 ,_u10_u5_n2467 , _u10_u5_n2466 , _u10_u5_n2465 , _u10_u5_n2464 ,_u10_u5_n2463 , _u10_u5_n2462 , _u10_u5_n2461 , _u10_u5_n2460 ,_u10_u5_n2459 , _u10_u5_n2458 , _u10_u5_n2457 , _u10_u5_n2456 ,_u10_u5_n2455 , _u10_u5_n2454 , _u10_u5_n2453 , _u10_u5_n2452 ,_u10_u5_n2451 , _u10_u5_n2450 , _u10_u5_n2449 , _u10_u5_n2448 ,_u10_u5_n2447 , _u10_u5_n2446 , _u10_u5_n2445 , _u10_u5_n2444 ,_u10_u5_n2443 , _u10_u5_n2442 , _u10_u5_n2441 , _u10_u5_n2440 ,_u10_u5_n2439 , _u10_u5_n2438 , _u10_u5_n2437 , _u10_u5_n2436 ,_u10_u5_n2435 , _u10_u5_n2434 , _u10_u5_n2433 , _u10_u5_n2432 ,_u10_u5_n2431 , _u10_u5_n2430 , _u10_u5_n2429 , _u10_u5_n2428 ,_u10_u5_n2427 , _u10_u5_n2426 , _u10_u5_n2425 , _u10_u5_n2424 ,_u10_u5_n2423 , _u10_u5_n2422 , _u10_u5_n2421 , _u10_u5_n2420 ,_u10_u5_n2419 , _u10_u5_n2418 , _u10_u5_n2417 , _u10_u5_n2416 ,_u10_u5_n2415 , _u10_u5_n2414 , _u10_u5_n2413 , _u10_u5_n2412 ,_u10_u5_n2411 , _u10_u5_n2410 , _u10_u5_n2409 , _u10_u5_n2408 ,_u10_u5_n2407 , _u10_u5_n2406 , _u10_u5_n2405 , _u10_u5_n2404 ,_u10_u5_n2403 , _u10_u5_n2402 , _u10_u5_n2401 , _u10_u5_n2400 ,_u10_u5_n2399 , _u10_u5_n2398 , _u10_u5_n2397 , _u10_u5_n2396 ,_u10_u5_n2395 , _u10_u5_n2394 , _u10_u5_n2393 , _u10_u5_n2392 ,_u10_u5_n2391 , _u10_u5_n2390 , _u10_u5_n2389 , _u10_u5_n2388 ,_u10_u5_n2387 , _u10_u5_n2386 , _u10_u5_n2385 , _u10_u5_n2384 ,_u10_u5_n2383 , _u10_u5_n2382 , _u10_u5_n2381 , _u10_u5_n2380 ,_u10_u5_n2379 , _u10_u5_n2378 , _u10_u5_n2377 , _u10_u5_n2376 ,_u10_u5_n2375 , _u10_u5_n2374 , _u10_u5_n2373 , _u10_u5_n2372 ,_u10_u5_n2371 , _u10_u5_n2370 , _u10_u5_n2369 , _u10_u5_n2368 ,_u10_u5_n2367 , _u10_u5_n2366 , _u10_u5_n2365 , _u10_u5_n2364 ,_u10_u5_n2363 , _u10_u5_n2362 , _u10_u5_n2361 , _u10_u5_n2360 ,_u10_u5_n2359 , _u10_u5_n2358 , _u10_u5_n2357 , _u10_u5_n2356 ,_u10_u5_n2355 , _u10_u5_n2354 , _u10_u5_n2353 , _u10_u5_n2352 ,_u10_u5_n2351 , _u10_u5_n2350 , _u10_u5_n2349 , _u10_u5_n2348 ,_u10_u5_n2347 , _u10_u5_n2346 , _u10_u5_n2345 , _u10_u5_n2344 ,_u10_u5_n2343 , _u10_u5_n2342 , _u10_u5_n2341 , _u10_u5_n2340 ,_u10_u5_n2339 , _u10_u5_n2338 , _u10_u5_n2337 , _u10_u5_n2336 ,_u10_u5_n2335 , _u10_u5_n2334 , _u10_u5_n2333 , _u10_u5_n2332 ,_u10_u5_n2331 , _u10_u5_n2330 , _u10_u5_n2329 , _u10_u5_n2328 ,_u10_u5_n2327 , _u10_u5_n2326 , _u10_u5_n2325 , _u10_u5_n2324 ,_u10_u5_n2323 , _u10_u5_n2322 , _u10_u5_n2321 , _u10_u5_n2320 ,_u10_u5_n2319 , _u10_u5_n2318 , _u10_u5_n2317 , _u10_u5_n2316 ,_u10_u5_n2315 , _u10_u5_n2314 , _u10_u5_n2313 , _u10_u5_n2312 ,_u10_u5_n2311 , _u10_u5_n2310 , _u10_u5_n2309 , _u10_u5_n2308 ,_u10_u5_n2307 , _u10_u5_n2306 , _u10_u5_n2305 , _u10_u5_n2304 ,_u10_u5_n2303 , _u10_u5_n2302 , _u10_u5_n2301 , _u10_u5_n2300 ,_u10_u5_n2299 , _u10_u5_n2298 , _u10_u5_n2297 , _u10_u5_n2296 ,_u10_u5_n2295 , _u10_u5_n2294 , _u10_u5_n2293 , _u10_u5_n2292 ,_u10_u5_n2291 , _u10_u5_n2290 , _u10_u5_n2289 , _u10_u5_n2288 ,_u10_u5_n2287 , _u10_u5_n2286 , _u10_u5_n2285 , _u10_u5_n2284 ,_u10_u5_n2283 , _u10_u5_n2282 , _u10_u5_n2281 , _u10_u5_n2280 ,_u10_u5_n2279 , _u10_u5_n2278 , _u10_u5_n2277 , _u10_u5_n2276 ,_u10_u5_n2275 , _u10_u5_n2274 , _u10_u5_n2273 , _u10_u5_n2272 ,_u10_u5_n2271 , _u10_u5_n2270 , _u10_u5_n2269 , _u10_u5_n2268 ,_u10_u5_n2267 , _u10_u5_n2266 , _u10_u5_n2265 , _u10_u5_n2264 ,_u10_u5_n2263 , _u10_u5_n2262 , _u10_u5_n2261 , _u10_u5_n2260 ,_u10_u5_n2259 , _u10_u5_n2258 , _u10_u5_n2257 , _u10_u5_n2256 ,_u10_u5_n2255 , _u10_u5_n2254 , _u10_u5_n2253 , _u10_u5_n2252 ,_u10_u5_n2251 , _u10_u5_n2250 , _u10_u5_n2249 , _u10_u5_n2248 ,_u10_u5_n2247 , _u10_u5_n2246 , _u10_u5_n2245 , _u10_u5_n2244 ,_u10_u5_n2243 , _u10_u5_n2242 , _u10_u5_n2241 , _u10_u5_n2240 ,_u10_u5_n2239 , _u10_u5_n2238 , _u10_u5_n2237 , _u10_u5_n2236 ,_u10_u5_n2235 , _u10_u5_n2234 , _u10_u5_n2233 , _u10_u5_n2232 ,_u10_u5_n2231 , _u10_u5_n2230 , _u10_u5_n2229 , _u10_u5_n2228 ,_u10_u5_n2227 , _u10_u5_n2226 , _u10_u5_n2225 , _u10_u5_n2224 ,_u10_u5_n2223 , _u10_u5_n2222 , _u10_u5_n2221 , _u10_u5_n2220 ,_u10_u5_n2219 , _u10_u5_n2218 , _u10_u5_n2217 , _u10_u5_n2216 ,_u10_u5_n2215 , _u10_u5_n2214 , _u10_u5_n2213 , _u10_u5_n2212 ,_u10_u5_n2211 , _u10_u5_n2210 , _u10_u5_n2209 , _u10_u5_n2208 ,_u10_u5_n2207 , _u10_u5_n2206 , _u10_u5_n2205 , _u10_u5_n2204 ,_u10_u5_n2203 , _u10_u5_n2202 , _u10_u5_n2201 , _u10_u5_n2200 ,_u10_u5_n2199 , _u10_u5_n2198 , _u10_u5_n2197 , _u10_u5_n2196 ,_u10_u5_n2195 , _u10_u5_n2194 , _u10_u5_n2193 , _u10_u5_n2192 ,_u10_u5_n2191 , _u10_u5_n2190 , _u10_u5_n2189 , _u10_u5_n2188 ,_u10_u5_n2187 , _u10_u5_n2186 , _u10_u5_n2185 , _u10_u5_n2184 ,_u10_u5_n2183 , _u10_u5_n2182 , _u10_u5_n2181 , _u10_u5_n2180 ,_u10_u5_n2179 , _u10_u5_n2178 , _u10_u5_n2177 , _u10_u5_n2176 ,_u10_u5_n2175 , _u10_u5_n2174 , _u10_u5_n2173 , _u10_u5_n2172 ,_u10_u5_n2171 , _u10_u5_n2170 , _u10_u5_n2169 , _u10_u5_n2168 ,_u10_u5_n2167 , _u10_u5_n2166 , _u10_u5_n2165 , _u10_u5_n2164 ,_u10_u5_n2163 , _u10_u5_n2162 , _u10_u5_n2161 , _u10_u5_n2160 ,_u10_u5_n2159 , _u10_u5_n2158 , _u10_u5_n2157 , _u10_u5_n2156 ,_u10_u5_n2155 , _u10_u5_n2154 , _u10_u5_n2153 , _u10_u5_n2152 ,_u10_u5_n2151 , _u10_u5_n2150 , _u10_u5_n2149 , _u10_u5_n2148 ,_u10_u5_n2147 , _u10_u5_n2146 , _u10_u5_n2145 , _u10_u5_n2144 ,_u10_u5_n2143 , _u10_u5_n2142 , _u10_u5_n2141 , _u10_u5_n2140 ,_u10_u5_n2139 , _u10_u5_n2138 , _u10_u5_n2137 , _u10_u5_n2136 ,_u10_u5_n2135 , _u10_u5_n2134 , _u10_u5_n2133 , _u10_u5_n2132 ,_u10_u5_n2131 , _u10_u5_n2130 , _u10_u5_n2129 , _u10_u5_n2128 ,_u10_u5_n2127 , _u10_u5_n2126 , _u10_u5_n2125 , _u10_u5_n2124 ,_u10_u5_n2123 , _u10_u5_n2122 , _u10_u5_n2121 , _u10_u5_n2120 ,_u10_u5_n2119 , _u10_u5_n2118 , _u10_u5_n2117 , _u10_u5_n2116 ,_u10_u5_n2115 , _u10_u5_n2114 , _u10_u5_n2113 , _u10_u5_n2112 ,_u10_u5_n2111 , _u10_u5_n2110 , _u10_u5_n2109 , _u10_u5_n2108 ,_u10_u5_n2107 , _u10_u5_n2106 , _u10_u5_n2105 , _u10_u5_n2104 ,_u10_u5_n2103 , _u10_u5_n2102 , _u10_u5_n2101 , _u10_u5_n2100 ,_u10_u5_n2099 , _u10_u5_n2098 , _u10_u5_n2097 , _u10_u5_n2096 ,_u10_u5_n2095 , _u10_u5_n2094 , _u10_u5_n2093 , _u10_u5_n2092 ,_u10_u5_n2091 , _u10_u5_n2090 , _u10_u5_n2089 , _u10_u5_n2088 ,_u10_u5_n2087 , _u10_u5_n2086 , _u10_u5_n2085 , _u10_u5_n2084 ,_u10_u5_n2083 , _u10_u5_n2082 , _u10_u5_n2081 , _u10_u5_n2080 ,_u10_u5_n2079 , _u10_u5_n2078 , _u10_u5_n2077 , _u10_u5_n2076 ,_u10_u5_n2075 , _u10_u5_n2074 , _u10_u5_n2073 , _u10_u5_n2072 ,_u10_u5_n2071 , _u10_u5_n2070 , _u10_u5_n2069 , _u10_u5_n2068 ,_u10_u5_n2067 , _u10_u5_n2066 , _u10_u5_n2065 , _u10_u5_n2064 ,_u10_u5_n2063 , _u10_u5_n2062 , _u10_u5_n2061 , _u10_u5_n2060 ,_u10_u5_n2059 , _u10_u5_n2058 , _u10_u5_n2057 , _u10_u5_n2056 ,_u10_u5_n2055 , _u10_u5_n2054 , _u10_u5_n2053 , _u10_u5_n2052 ,_u10_u5_n2051 , _u10_u5_n2050 , _u10_u5_n2049 , _u10_u5_n2048 ,_u10_u5_n2047 , _u10_u5_n2046 , _u10_u5_n2045 , _u10_u5_n2044 ,_u10_u5_n2043 , _u10_u5_n2042 , _u10_u5_n2041 , _u10_u5_n2040 ,_u10_u5_n2039 , _u10_u5_n2038 , _u10_u5_n2037 , _u10_u5_n2036 ,_u10_u5_n2035 , _u10_u5_n2034 , _u10_u5_n2033 , _u10_u5_n2032 ,_u10_u5_n2031 , _u10_u5_n2030 , _u10_u5_n2029 , _u10_u5_n2028 ,_u10_u5_n2027 , _u10_u5_n2026 , _u10_u5_n2025 , _u10_u5_n2024 ,_u10_u5_n2023 , _u10_u5_n2022 , _u10_u5_n2021 , _u10_u5_n2020 ,_u10_u5_n2019 , _u10_u5_n2018 , _u10_u5_n2017 , _u10_u5_n2016 ,_u10_u5_n2015 , _u10_u5_n2014 , _u10_u5_n2013 , _u10_u5_n2012 ,_u10_u5_n2011 , _u10_u5_n2010 , _u10_u5_n2009 , _u10_u5_n2008 ,_u10_u5_n2007 , _u10_u5_n2006 , _u10_u5_n2005 , _u10_u5_n2004 ,_u10_u5_n2003 , _u10_u5_n2002 , _u10_u5_n2001 , _u10_u5_n2000 ,_u10_u5_n1999 , _u10_u5_n1998 , _u10_u5_n1997 , _u10_u5_n1996 ,_u10_u5_n1995 , _u10_u5_n1994 , _u10_u5_n1993 , _u10_u5_n1992 ,_u10_u5_n1991 , _u10_u5_n1990 , _u10_u5_n1989 , _u10_u5_n1988 ,_u10_u5_n1987 , _u10_u5_n1986 , _u10_u5_n1985 , _u10_u5_n1984 ,_u10_u5_n1983 , _u10_u5_n1982 , _u10_u5_n1981 , _u10_u5_n1980 ,_u10_u5_n1979 , _u10_u5_n1978 , _u10_u5_n1977 , _u10_u5_n1976 ,_u10_u5_n1975 , _u10_u5_n1974 , _u10_u5_n1973 , _u10_u5_n1972 ,_u10_u5_n1971 , _u10_u5_n1970 , _u10_u5_n1969 , _u10_u5_n1968 ,_u10_u5_n1967 , _u10_u5_n1966 , _u10_u5_n1965 , _u10_u5_n1964 ,_u10_u5_n1963 , _u10_u5_n1962 , _u10_u5_n1961 , _u10_u5_n1960 ,_u10_u5_n1959 , _u10_u5_n1958 , _u10_u5_n1957 , _u10_u5_n1956 ,_u10_u5_n1955 , _u10_u5_n1954 , _u10_u5_n1953 , _u10_u5_n1952 ,_u10_u5_n1951 , _u10_u5_n1950 , _u10_u5_n1949 , _u10_u5_n1948 ,_u10_u5_n1947 , _u10_u5_n1946 , _u10_u5_n1945 , _u10_u5_n1944 ,_u10_u5_n1943 , _u10_u5_n1942 , _u10_u5_n1941 , _u10_u5_n1940 ,_u10_u5_n1939 , _u10_u5_n1938 , _u10_u5_n1937 , _u10_u5_n1936 ,_u10_u5_n1935 , _u10_u5_n1934 , _u10_u5_n1933 , _u10_u5_n1932 ,_u10_u5_n1931 , _u10_u5_n1930 , _u10_u5_n1929 , _u10_u5_n1928 ,_u10_u5_n1927 , _u10_u5_n1926 , _u10_u5_n1925 , _u10_u5_n1924 ,_u10_u5_n1923 , _u10_u5_n1922 , _u10_u5_n1921 , _u10_u5_n1920 ,_u10_u5_n1919 , _u10_u5_n1918 , _u10_u5_n1917 , _u10_u5_n1916 ,_u10_u5_n1915 , _u10_u5_n1914 , _u10_u5_n1913 , _u10_u5_n1912 ,_u10_u5_n1911 , _u10_u5_n1910 , _u10_u5_n1909 , _u10_u5_n1908 ,_u10_u5_n1907 , _u10_u5_n1906 , _u10_u5_n1905 , _u10_u5_n1904 ,_u10_u5_n1903 , _u10_u5_n1902 , _u10_u5_n1901 , _u10_u5_n1900 ,_u10_u5_n1899 , _u10_u5_n1898 , _u10_u5_n1897 , _u10_u5_n1896 ,_u10_u5_n1895 , _u10_u5_n1894 , _u10_u5_n1893 , _u10_u5_n1892 ,_u10_u5_n1891 , _u10_u5_n1890 , _u10_u5_n1889 , _u10_u5_n1888 ,_u10_u5_n1887 , _u10_u5_n1886 , _u10_u5_n1885 , _u10_u5_n1884 ,_u10_u5_n1883 , _u10_u5_n1882 , _u10_u5_n1881 , _u10_u5_n1880 ,_u10_u5_n1879 , _u10_u5_n1878 , _u10_u5_n1877 , _u10_u5_n1876 ,_u10_u5_n1875 , _u10_u5_n1874 , _u10_u5_n1873 , _u10_u5_n1872 ,_u10_u5_n1871 , _u10_u5_n1870 , _u10_u5_n1869 , _u10_u5_n1868 ,_u10_u5_n1867 , _u10_u5_n1866 , _u10_u5_n1865 , _u10_u5_n1864 ,_u10_u5_n1863 , _u10_u5_n1862 , _u10_u5_n1861 , _u10_u5_n1860 ,_u10_u5_n1859 , _u10_u5_n1858 , _u10_u5_n1857 , _u10_u5_n1856 ,_u10_u5_n1855 , _u10_u5_n1854 , _u10_u5_n1853 , _u10_u5_n1852 ,_u10_u5_n1851 , _u10_u5_n1850 , _u10_u5_n1849 , _u10_u5_n1848 ,_u10_u5_n1847 , _u10_u5_n1846 , _u10_u5_n1845 , _u10_u5_n1844 ,_u10_u5_n1843 , _u10_u5_n1842 , _u10_u5_n1841 , _u10_u5_n1840 ,_u10_u5_n1839 , _u10_u5_n1838 , _u10_u5_n1837 , _u10_u5_n1836 ,_u10_u5_n1835 , _u10_u5_n1834 , _u10_u5_n1833 , _u10_u5_n1832 ,_u10_u5_n1831 , _u10_u5_n1830 , _u10_u5_n1829 , _u10_u5_n1828 ,_u10_u5_n1827 , _u10_u5_n1826 , _u10_u5_n1825 , _u10_u5_n1824 ,_u10_u5_n1823 , _u10_u5_n1822 , _u10_u5_n1821 , _u10_u5_n1820 ,_u10_u5_n1819 , _u10_u5_n1818 , _u10_u5_n1817 , _u10_u5_n1816 ,_u10_u5_n1815 , _u10_u5_n1814 , _u10_u5_n1813 , _u10_u5_n1812 ,_u10_u5_n1811 , _u10_u5_n1810 , _u10_u5_n1809 , _u10_u5_n1808 ,_u10_u6_n3416 , _u10_u6_n3415 , _u10_u6_n3414 , _u10_u6_n3413 ,_u10_u6_n3412 , _u10_u6_n3411 , _u10_u6_n3410 , _u10_u6_n3409 ,_u10_u6_n3408 , _u10_u6_n3407 , _u10_u6_n3406 , _u10_u6_n3405 ,_u10_u6_n3404 , _u10_u6_n3403 , _u10_u6_n3402 , _u10_u6_n3401 ,_u10_u6_n3400 , _u10_u6_n3399 , _u10_u6_n3398 , _u10_u6_n3397 ,_u10_u6_n3396 , _u10_u6_n3395 , _u10_u6_n3394 , _u10_u6_n3393 ,_u10_u6_n3392 , _u10_u6_n3391 , _u10_u6_n3390 , _u10_u6_n3389 ,_u10_u6_n3388 , _u10_u6_n3387 , _u10_u6_n3386 , _u10_u6_n3385 ,_u10_u6_n3384 , _u10_u6_n3383 , _u10_u6_n3382 , _u10_u6_n3381 ,_u10_u6_n3380 , _u10_u6_n3379 , _u10_u6_n3378 , _u10_u6_n3377 ,_u10_u6_n3376 , _u10_u6_n3375 , _u10_u6_n3374 , _u10_u6_n3373 ,_u10_u6_n3372 , _u10_u6_n3371 , _u10_u6_n3370 , _u10_u6_n3369 ,_u10_u6_n3368 , _u10_u6_n3367 , _u10_u6_n3366 , _u10_u6_n3365 ,_u10_u6_n3364 , _u10_u6_n3363 , _u10_u6_n3362 , _u10_u6_n3361 ,_u10_u6_n3360 , _u10_u6_n3359 , _u10_u6_n3358 , _u10_u6_n3357 ,_u10_u6_n3356 , _u10_u6_n3355 , _u10_u6_n3354 , _u10_u6_n3353 ,_u10_u6_n3352 , _u10_u6_n3351 , _u10_u6_n3350 , _u10_u6_n3349 ,_u10_u6_n3348 , _u10_u6_n3347 , _u10_u6_n3346 , _u10_u6_n3345 ,_u10_u6_n3344 , _u10_u6_n3343 , _u10_u6_n3342 , _u10_u6_n3341 ,_u10_u6_n3340 , _u10_u6_n3339 , _u10_u6_n3338 , _u10_u6_n3337 ,_u10_u6_n3336 , _u10_u6_n3335 , _u10_u6_n3334 , _u10_u6_n3333 ,_u10_u6_n3332 , _u10_u6_n3331 , _u10_u6_n3330 , _u10_u6_n3329 ,_u10_u6_n3328 , _u10_u6_n3327 , _u10_u6_n3326 , _u10_u6_n3325 ,_u10_u6_n3324 , _u10_u6_n3323 , _u10_u6_n3322 , _u10_u6_n3321 ,_u10_u6_n3320 , _u10_u6_n3319 , _u10_u6_n3318 , _u10_u6_n3317 ,_u10_u6_n3316 , _u10_u6_n3315 , _u10_u6_n3314 , _u10_u6_n3313 ,_u10_u6_n3312 , _u10_u6_n3311 , _u10_u6_n3310 , _u10_u6_n3309 ,_u10_u6_n3308 , _u10_u6_n3307 , _u10_u6_n3306 , _u10_u6_n3305 ,_u10_u6_n3304 , _u10_u6_n3303 , _u10_u6_n3302 , _u10_u6_n3301 ,_u10_u6_n3300 , _u10_u6_n3299 , _u10_u6_n3298 , _u10_u6_n3297 ,_u10_u6_n3296 , _u10_u6_n3295 , _u10_u6_n3294 , _u10_u6_n3293 ,_u10_u6_n3292 , _u10_u6_n3291 , _u10_u6_n3290 , _u10_u6_n3289 ,_u10_u6_n3288 , _u10_u6_n3287 , _u10_u6_n3286 , _u10_u6_n3285 ,_u10_u6_n3284 , _u10_u6_n3283 , _u10_u6_n3282 , _u10_u6_n3281 ,_u10_u6_n3280 , _u10_u6_n3279 , _u10_u6_n3278 , _u10_u6_n3277 ,_u10_u6_n3276 , _u10_u6_n3275 , _u10_u6_n3274 , _u10_u6_n3273 ,_u10_u6_n3272 , _u10_u6_n3271 , _u10_u6_n3270 , _u10_u6_n3269 ,_u10_u6_n3268 , _u10_u6_n3267 , _u10_u6_n3266 , _u10_u6_n3265 ,_u10_u6_n3264 , _u10_u6_n3263 , _u10_u6_n3262 , _u10_u6_n3261 ,_u10_u6_n3260 , _u10_u6_n3259 , _u10_u6_n3258 , _u10_u6_n3257 ,_u10_u6_n3256 , _u10_u6_n3255 , _u10_u6_n3254 , _u10_u6_n3253 ,_u10_u6_n3252 , _u10_u6_n3251 , _u10_u6_n3250 , _u10_u6_n3249 ,_u10_u6_n3248 , _u10_u6_n3247 , _u10_u6_n3246 , _u10_u6_n3245 ,_u10_u6_n3244 , _u10_u6_n3243 , _u10_u6_n3242 , _u10_u6_n3241 ,_u10_u6_n3240 , _u10_u6_n3239 , _u10_u6_n3238 , _u10_u6_n3237 ,_u10_u6_n3236 , _u10_u6_n3235 , _u10_u6_n3234 , _u10_u6_n3233 ,_u10_u6_n3232 , _u10_u6_n3231 , _u10_u6_n3230 , _u10_u6_n3229 ,_u10_u6_n3228 , _u10_u6_n3227 , _u10_u6_n3226 , _u10_u6_n3225 ,_u10_u6_n3224 , _u10_u6_n3223 , _u10_u6_n3222 , _u10_u6_n3221 ,_u10_u6_n3220 , _u10_u6_n3219 , _u10_u6_n3218 , _u10_u6_n3217 ,_u10_u6_n3216 , _u10_u6_n3215 , _u10_u6_n3214 , _u10_u6_n3213 ,_u10_u6_n3212 , _u10_u6_n3211 , _u10_u6_n3210 , _u10_u6_n3209 ,_u10_u6_n3208 , _u10_u6_n3207 , _u10_u6_n3206 , _u10_u6_n3205 ,_u10_u6_n3204 , _u10_u6_n3203 , _u10_u6_n3202 , _u10_u6_n3201 ,_u10_u6_n3200 , _u10_u6_n3199 , _u10_u6_n3198 , _u10_u6_n3197 ,_u10_u6_n3196 , _u10_u6_n3195 , _u10_u6_n3194 , _u10_u6_n3193 ,_u10_u6_n3192 , _u10_u6_n3191 , _u10_u6_n3190 , _u10_u6_n3189 ,_u10_u6_n3188 , _u10_u6_n3187 , _u10_u6_n3186 , _u10_u6_n3185 ,_u10_u6_n3184 , _u10_u6_n3183 , _u10_u6_n3182 , _u10_u6_n3181 ,_u10_u6_n3180 , _u10_u6_n3179 , _u10_u6_n3178 , _u10_u6_n3177 ,_u10_u6_n3176 , _u10_u6_n3175 , _u10_u6_n3174 , _u10_u6_n3173 ,_u10_u6_n3172 , _u10_u6_n3171 , _u10_u6_n3170 , _u10_u6_n3169 ,_u10_u6_n3168 , _u10_u6_n3167 , _u10_u6_n3166 , _u10_u6_n3165 ,_u10_u6_n3164 , _u10_u6_n3163 , _u10_u6_n3162 , _u10_u6_n3161 ,_u10_u6_n3160 , _u10_u6_n3159 , _u10_u6_n3158 , _u10_u6_n3157 ,_u10_u6_n3156 , _u10_u6_n3155 , _u10_u6_n3154 , _u10_u6_n3153 ,_u10_u6_n3152 , _u10_u6_n3151 , _u10_u6_n3150 , _u10_u6_n3149 ,_u10_u6_n3148 , _u10_u6_n3147 , _u10_u6_n3146 , _u10_u6_n3145 ,_u10_u6_n3144 , _u10_u6_n3143 , _u10_u6_n3142 , _u10_u6_n3141 ,_u10_u6_n3140 , _u10_u6_n3139 , _u10_u6_n3138 , _u10_u6_n3137 ,_u10_u6_n3136 , _u10_u6_n3135 , _u10_u6_n3134 , _u10_u6_n3133 ,_u10_u6_n3132 , _u10_u6_n3131 , _u10_u6_n3130 , _u10_u6_n3129 ,_u10_u6_n3128 , _u10_u6_n3127 , _u10_u6_n3126 , _u10_u6_n3125 ,_u10_u6_n3124 , _u10_u6_n3123 , _u10_u6_n3122 , _u10_u6_n3121 ,_u10_u6_n3120 , _u10_u6_n3119 , _u10_u6_n3118 , _u10_u6_n3117 ,_u10_u6_n3116 , _u10_u6_n3115 , _u10_u6_n3114 , _u10_u6_n3113 ,_u10_u6_n3112 , _u10_u6_n3111 , _u10_u6_n3110 , _u10_u6_n3109 ,_u10_u6_n3108 , _u10_u6_n3107 , _u10_u6_n3106 , _u10_u6_n3105 ,_u10_u6_n3104 , _u10_u6_n3103 , _u10_u6_n3102 , _u10_u6_n3101 ,_u10_u6_n3100 , _u10_u6_n3099 , _u10_u6_n3098 , _u10_u6_n3097 ,_u10_u6_n3096 , _u10_u6_n3095 , _u10_u6_n3094 , _u10_u6_n3093 ,_u10_u6_n3092 , _u10_u6_n3091 , _u10_u6_n3090 , _u10_u6_n3089 ,_u10_u6_n3088 , _u10_u6_n3087 , _u10_u6_n3086 , _u10_u6_n3085 ,_u10_u6_n3084 , _u10_u6_n3083 , _u10_u6_n3082 , _u10_u6_n3081 ,_u10_u6_n3080 , _u10_u6_n3079 , _u10_u6_n3078 , _u10_u6_n3077 ,_u10_u6_n3076 , _u10_u6_n3075 , _u10_u6_n3074 , _u10_u6_n3073 ,_u10_u6_n3072 , _u10_u6_n3071 , _u10_u6_n3070 , _u10_u6_n3069 ,_u10_u6_n3068 , _u10_u6_n3067 , _u10_u6_n3066 , _u10_u6_n3065 ,_u10_u6_n3064 , _u10_u6_n3063 , _u10_u6_n3062 , _u10_u6_n3061 ,_u10_u6_n3060 , _u10_u6_n3059 , _u10_u6_n3058 , _u10_u6_n3057 ,_u10_u6_n3056 , _u10_u6_n3055 , _u10_u6_n3054 , _u10_u6_n3053 ,_u10_u6_n3052 , _u10_u6_n3051 , _u10_u6_n3050 , _u10_u6_n3049 ,_u10_u6_n3048 , _u10_u6_n3047 , _u10_u6_n3046 , _u10_u6_n3045 ,_u10_u6_n3044 , _u10_u6_n3043 , _u10_u6_n3042 , _u10_u6_n3041 ,_u10_u6_n3040 , _u10_u6_n3039 , _u10_u6_n3038 , _u10_u6_n3037 ,_u10_u6_n3036 , _u10_u6_n3035 , _u10_u6_n3034 , _u10_u6_n3033 ,_u10_u6_n3032 , _u10_u6_n3031 , _u10_u6_n3030 , _u10_u6_n3029 ,_u10_u6_n3028 , _u10_u6_n3027 , _u10_u6_n3026 , _u10_u6_n3025 ,_u10_u6_n3024 , _u10_u6_n3023 , _u10_u6_n3022 , _u10_u6_n3021 ,_u10_u6_n3020 , _u10_u6_n3019 , _u10_u6_n3018 , _u10_u6_n3017 ,_u10_u6_n3016 , _u10_u6_n3015 , _u10_u6_n3014 , _u10_u6_n3013 ,_u10_u6_n3012 , _u10_u6_n3011 , _u10_u6_n3010 , _u10_u6_n3009 ,_u10_u6_n3008 , _u10_u6_n3007 , _u10_u6_n3006 , _u10_u6_n3005 ,_u10_u6_n3004 , _u10_u6_n3003 , _u10_u6_n3002 , _u10_u6_n3001 ,_u10_u6_n3000 , _u10_u6_n2999 , _u10_u6_n2998 , _u10_u6_n2997 ,_u10_u6_n2996 , _u10_u6_n2995 , _u10_u6_n2994 , _u10_u6_n2993 ,_u10_u6_n2992 , _u10_u6_n2991 , _u10_u6_n2990 , _u10_u6_n2989 ,_u10_u6_n2988 , _u10_u6_n2987 , _u10_u6_n2986 , _u10_u6_n2985 ,_u10_u6_n2984 , _u10_u6_n2983 , _u10_u6_n2982 , _u10_u6_n2981 ,_u10_u6_n2980 , _u10_u6_n2979 , _u10_u6_n2978 , _u10_u6_n2977 ,_u10_u6_n2976 , _u10_u6_n2975 , _u10_u6_n2974 , _u10_u6_n2973 ,_u10_u6_n2972 , _u10_u6_n2971 , _u10_u6_n2970 , _u10_u6_n2969 ,_u10_u6_n2968 , _u10_u6_n2967 , _u10_u6_n2966 , _u10_u6_n2965 ,_u10_u6_n2964 , _u10_u6_n2963 , _u10_u6_n2962 , _u10_u6_n2961 ,_u10_u6_n2960 , _u10_u6_n2959 , _u10_u6_n2958 , _u10_u6_n2957 ,_u10_u6_n2956 , _u10_u6_n2955 , _u10_u6_n2954 , _u10_u6_n2953 ,_u10_u6_n2952 , _u10_u6_n2951 , _u10_u6_n2950 , _u10_u6_n2949 ,_u10_u6_n2948 , _u10_u6_n2947 , _u10_u6_n2946 , _u10_u6_n2945 ,_u10_u6_n2944 , _u10_u6_n2943 , _u10_u6_n2942 , _u10_u6_n2941 ,_u10_u6_n2940 , _u10_u6_n2939 , _u10_u6_n2938 , _u10_u6_n2937 ,_u10_u6_n2936 , _u10_u6_n2935 , _u10_u6_n2934 , _u10_u6_n2933 ,_u10_u6_n2932 , _u10_u6_n2931 , _u10_u6_n2930 , _u10_u6_n2929 ,_u10_u6_n2928 , _u10_u6_n2927 , _u10_u6_n2926 , _u10_u6_n2925 ,_u10_u6_n2924 , _u10_u6_n2923 , _u10_u6_n2922 , _u10_u6_n2921 ,_u10_u6_n2920 , _u10_u6_n2919 , _u10_u6_n2918 , _u10_u6_n2917 ,_u10_u6_n2916 , _u10_u6_n2915 , _u10_u6_n2914 , _u10_u6_n2913 ,_u10_u6_n2912 , _u10_u6_n2911 , _u10_u6_n2910 , _u10_u6_n2909 ,_u10_u6_n2908 , _u10_u6_n2907 , _u10_u6_n2906 , _u10_u6_n2905 ,_u10_u6_n2904 , _u10_u6_n2903 , _u10_u6_n2902 , _u10_u6_n2901 ,_u10_u6_n2900 , _u10_u6_n2899 , _u10_u6_n2898 , _u10_u6_n2897 ,_u10_u6_n2896 , _u10_u6_n2895 , _u10_u6_n2894 , _u10_u6_n2893 ,_u10_u6_n2892 , _u10_u6_n2891 , _u10_u6_n2890 , _u10_u6_n2889 ,_u10_u6_n2888 , _u10_u6_n2887 , _u10_u6_n2886 , _u10_u6_n2885 ,_u10_u6_n2884 , _u10_u6_n2883 , _u10_u6_n2882 , _u10_u6_n2881 ,_u10_u6_n2880 , _u10_u6_n2879 , _u10_u6_n2878 , _u10_u6_n2877 ,_u10_u6_n2876 , _u10_u6_n2875 , _u10_u6_n2874 , _u10_u6_n2873 ,_u10_u6_n2872 , _u10_u6_n2871 , _u10_u6_n2870 , _u10_u6_n2869 ,_u10_u6_n2868 , _u10_u6_n2867 , _u10_u6_n2866 , _u10_u6_n2865 ,_u10_u6_n2864 , _u10_u6_n2863 , _u10_u6_n2862 , _u10_u6_n2861 ,_u10_u6_n2860 , _u10_u6_n2859 , _u10_u6_n2858 , _u10_u6_n2857 ,_u10_u6_n2856 , _u10_u6_n2855 , _u10_u6_n2854 , _u10_u6_n2853 ,_u10_u6_n2852 , _u10_u6_n2851 , _u10_u6_n2850 , _u10_u6_n2849 ,_u10_u6_n2848 , _u10_u6_n2847 , _u10_u6_n2846 , _u10_u6_n2845 ,_u10_u6_n2844 , _u10_u6_n2843 , _u10_u6_n2842 , _u10_u6_n2841 ,_u10_u6_n2840 , _u10_u6_n2839 , _u10_u6_n2838 , _u10_u6_n2837 ,_u10_u6_n2836 , _u10_u6_n2835 , _u10_u6_n2834 , _u10_u6_n2833 ,_u10_u6_n2832 , _u10_u6_n2831 , _u10_u6_n2830 , _u10_u6_n2829 ,_u10_u6_n2828 , _u10_u6_n2827 , _u10_u6_n2826 , _u10_u6_n2825 ,_u10_u6_n2824 , _u10_u6_n2823 , _u10_u6_n2822 , _u10_u6_n2821 ,_u10_u6_n2820 , _u10_u6_n2819 , _u10_u6_n2818 , _u10_u6_n2817 ,_u10_u6_n2816 , _u10_u6_n2815 , _u10_u6_n2814 , _u10_u6_n2813 ,_u10_u6_n2812 , _u10_u6_n2811 , _u10_u6_n2810 , _u10_u6_n2809 ,_u10_u6_n2808 , _u10_u6_n2807 , _u10_u6_n2806 , _u10_u6_n2805 ,_u10_u6_n2804 , _u10_u6_n2803 , _u10_u6_n2802 , _u10_u6_n2801 ,_u10_u6_n2800 , _u10_u6_n2799 , _u10_u6_n2798 , _u10_u6_n2797 ,_u10_u6_n2796 , _u10_u6_n2795 , _u10_u6_n2794 , _u10_u6_n2793 ,_u10_u6_n2792 , _u10_u6_n2791 , _u10_u6_n2790 , _u10_u6_n2789 ,_u10_u6_n2788 , _u10_u6_n2787 , _u10_u6_n2786 , _u10_u6_n2785 ,_u10_u6_n2784 , _u10_u6_n2783 , _u10_u6_n2782 , _u10_u6_n2781 ,_u10_u6_n2780 , _u10_u6_n2779 , _u10_u6_n2778 , _u10_u6_n2777 ,_u10_u6_n2776 , _u10_u6_n2775 , _u10_u6_n2774 , _u10_u6_n2773 ,_u10_u6_n2772 , _u10_u6_n2771 , _u10_u6_n2770 , _u10_u6_n2769 ,_u10_u6_n2768 , _u10_u6_n2767 , _u10_u6_n2766 , _u10_u6_n2765 ,_u10_u6_n2764 , _u10_u6_n2763 , _u10_u6_n2762 , _u10_u6_n2761 ,_u10_u6_n2760 , _u10_u6_n2759 , _u10_u6_n2758 , _u10_u6_n2757 ,_u10_u6_n2756 , _u10_u6_n2755 , _u10_u6_n2754 , _u10_u6_n2753 ,_u10_u6_n2752 , _u10_u6_n2751 , _u10_u6_n2750 , _u10_u6_n2749 ,_u10_u6_n2748 , _u10_u6_n2747 , _u10_u6_n2746 , _u10_u6_n2745 ,_u10_u6_n2744 , _u10_u6_n2743 , _u10_u6_n2742 , _u10_u6_n2741 ,_u10_u6_n2740 , _u10_u6_n2739 , _u10_u6_n2738 , _u10_u6_n2737 ,_u10_u6_n2736 , _u10_u6_n2735 , _u10_u6_n2734 , _u10_u6_n2733 ,_u10_u6_n2732 , _u10_u6_n2731 , _u10_u6_n2730 , _u10_u6_n2729 ,_u10_u6_n2728 , _u10_u6_n2727 , _u10_u6_n2726 , _u10_u6_n2725 ,_u10_u6_n2724 , _u10_u6_n2723 , _u10_u6_n2722 , _u10_u6_n2721 ,_u10_u6_n2720 , _u10_u6_n2719 , _u10_u6_n2718 , _u10_u6_n2717 ,_u10_u6_n2716 , _u10_u6_n2715 , _u10_u6_n2714 , _u10_u6_n2713 ,_u10_u6_n2712 , _u10_u6_n2711 , _u10_u6_n2710 , _u10_u6_n2709 ,_u10_u6_n2708 , _u10_u6_n2707 , _u10_u6_n2706 , _u10_u6_n2705 ,_u10_u6_n2704 , _u10_u6_n2703 , _u10_u6_n2702 , _u10_u6_n2701 ,_u10_u6_n2700 , _u10_u6_n2699 , _u10_u6_n2698 , _u10_u6_n2697 ,_u10_u6_n2696 , _u10_u6_n2695 , _u10_u6_n2694 , _u10_u6_n2693 ,_u10_u6_n2692 , _u10_u6_n2691 , _u10_u6_n2690 , _u10_u6_n2689 ,_u10_u6_n2688 , _u10_u6_n2687 , _u10_u6_n2686 , _u10_u6_n2685 ,_u10_u6_n2684 , _u10_u6_n2683 , _u10_u6_n2682 , _u10_u6_n2681 ,_u10_u6_n2680 , _u10_u6_n2679 , _u10_u6_n2678 , _u10_u6_n2677 ,_u10_u6_n2676 , _u10_u6_n2675 , _u10_u6_n2674 , _u10_u6_n2673 ,_u10_u6_n2672 , _u10_u6_n2671 , _u10_u6_n2670 , _u10_u6_n2669 ,_u10_u6_n2668 , _u10_u6_n2667 , _u10_u6_n2666 , _u10_u6_n2665 ,_u10_u6_n2664 , _u10_u6_n2663 , _u10_u6_n2662 , _u10_u6_n2661 ,_u10_u6_n2660 , _u10_u6_n2659 , _u10_u6_n2658 , _u10_u6_n2657 ,_u10_u6_n2656 , _u10_u6_n2655 , _u10_u6_n2654 , _u10_u6_n2653 ,_u10_u6_n2652 , _u10_u6_n2651 , _u10_u6_n2650 , _u10_u6_n2649 ,_u10_u6_n2648 , _u10_u6_n2647 , _u10_u6_n2646 , _u10_u6_n2645 ,_u10_u6_n2644 , _u10_u6_n2643 , _u10_u6_n2642 , _u10_u6_n2641 ,_u10_u6_n2640 , _u10_u6_n2639 , _u10_u6_n2638 , _u10_u6_n2637 ,_u10_u6_n2636 , _u10_u6_n2635 , _u10_u6_n2634 , _u10_u6_n2633 ,_u10_u6_n2632 , _u10_u6_n2631 , _u10_u6_n2630 , _u10_u6_n2629 ,_u10_u6_n2628 , _u10_u6_n2627 , _u10_u6_n2626 , _u10_u6_n2625 ,_u10_u6_n2624 , _u10_u6_n2623 , _u10_u6_n2622 , _u10_u6_n2621 ,_u10_u6_n2620 , _u10_u6_n2619 , _u10_u6_n2618 , _u10_u6_n2617 ,_u10_u6_n2616 , _u10_u6_n2615 , _u10_u6_n2614 , _u10_u6_n2613 ,_u10_u6_n2612 , _u10_u6_n2611 , _u10_u6_n2610 , _u10_u6_n2609 ,_u10_u6_n2608 , _u10_u6_n2607 , _u10_u6_n2606 , _u10_u6_n2605 ,_u10_u6_n2604 , _u10_u6_n2603 , _u10_u6_n2602 , _u10_u6_n2601 ,_u10_u6_n2600 , _u10_u6_n2599 , _u10_u6_n2598 , _u10_u6_n2597 ,_u10_u6_n2596 , _u10_u6_n2595 , _u10_u6_n2594 , _u10_u6_n2593 ,_u10_u6_n2592 , _u10_u6_n2591 , _u10_u6_n2590 , _u10_u6_n2589 ,_u10_u6_n2588 , _u10_u6_n2587 , _u10_u6_n2586 , _u10_u6_n2585 ,_u10_u6_n2584 , _u10_u6_n2583 , _u10_u6_n2582 , _u10_u6_n2581 ,_u10_u6_n2580 , _u10_u6_n2579 , _u10_u6_n2578 , _u10_u6_n2577 ,_u10_u6_n2576 , _u10_u6_n2575 , _u10_u6_n2574 , _u10_u6_n2573 ,_u10_u6_n2572 , _u10_u6_n2571 , _u10_u6_n2570 , _u10_u6_n2569 ,_u10_u6_n2568 , _u10_u6_n2567 , _u10_u6_n2566 , _u10_u6_n2565 ,_u10_u6_n2564 , _u10_u6_n2563 , _u10_u6_n2562 , _u10_u6_n2561 ,_u10_u6_n2560 , _u10_u6_n2559 , _u10_u6_n2558 , _u10_u6_n2557 ,_u10_u6_n2556 , _u10_u6_n2555 , _u10_u6_n2554 , _u10_u6_n2553 ,_u10_u6_n2552 , _u10_u6_n2551 , _u10_u6_n2550 , _u10_u6_n2549 ,_u10_u6_n2548 , _u10_u6_n2547 , _u10_u6_n2546 , _u10_u6_n2545 ,_u10_u6_n2544 , _u10_u6_n2543 , _u10_u6_n2542 , _u10_u6_n2541 ,_u10_u6_n2540 , _u10_u6_n2539 , _u10_u6_n2538 , _u10_u6_n2537 ,_u10_u6_n2536 , _u10_u6_n2535 , _u10_u6_n2534 , _u10_u6_n2533 ,_u10_u6_n2532 , _u10_u6_n2531 , _u10_u6_n2530 , _u10_u6_n2529 ,_u10_u6_n2528 , _u10_u6_n2527 , _u10_u6_n2526 , _u10_u6_n2525 ,_u10_u6_n2524 , _u10_u6_n2523 , _u10_u6_n2522 , _u10_u6_n2521 ,_u10_u6_n2520 , _u10_u6_n2519 , _u10_u6_n2518 , _u10_u6_n2517 ,_u10_u6_n2516 , _u10_u6_n2515 , _u10_u6_n2514 , _u10_u6_n2513 ,_u10_u6_n2512 , _u10_u6_n2511 , _u10_u6_n2510 , _u10_u6_n2509 ,_u10_u6_n2508 , _u10_u6_n2507 , _u10_u6_n2506 , _u10_u6_n2505 ,_u10_u6_n2504 , _u10_u6_n2503 , _u10_u6_n2502 , _u10_u6_n2501 ,_u10_u6_n2500 , _u10_u6_n2499 , _u10_u6_n2498 , _u10_u6_n2497 ,_u10_u6_n2496 , _u10_u6_n2495 , _u10_u6_n2494 , _u10_u6_n2493 ,_u10_u6_n2492 , _u10_u6_n2491 , _u10_u6_n2490 , _u10_u6_n2489 ,_u10_u6_n2488 , _u10_u6_n2487 , _u10_u6_n2486 , _u10_u6_n2485 ,_u10_u6_n2484 , _u10_u6_n2483 , _u10_u6_n2482 , _u10_u6_n2481 ,_u10_u6_n2480 , _u10_u6_n2479 , _u10_u6_n2478 , _u10_u6_n2477 ,_u10_u6_n2476 , _u10_u6_n2475 , _u10_u6_n2474 , _u10_u6_n2473 ,_u10_u6_n2472 , _u10_u6_n2471 , _u10_u6_n2470 , _u10_u6_n2469 ,_u10_u6_n2468 , _u10_u6_n2467 , _u10_u6_n2466 , _u10_u6_n2465 ,_u10_u6_n2464 , _u10_u6_n2463 , _u10_u6_n2462 , _u10_u6_n2461 ,_u10_u6_n2460 , _u10_u6_n2459 , _u10_u6_n2458 , _u10_u6_n2457 ,_u10_u6_n2456 , _u10_u6_n2455 , _u10_u6_n2454 , _u10_u6_n2453 ,_u10_u6_n2452 , _u10_u6_n2451 , _u10_u6_n2450 , _u10_u6_n2449 ,_u10_u6_n2448 , _u10_u6_n2447 , _u10_u6_n2446 , _u10_u6_n2445 ,_u10_u6_n2444 , _u10_u6_n2443 , _u10_u6_n2442 , _u10_u6_n2441 ,_u10_u6_n2440 , _u10_u6_n2439 , _u10_u6_n2438 , _u10_u6_n2437 ,_u10_u6_n2436 , _u10_u6_n2435 , _u10_u6_n2434 , _u10_u6_n2433 ,_u10_u6_n2432 , _u10_u6_n2431 , _u10_u6_n2430 , _u10_u6_n2429 ,_u10_u6_n2428 , _u10_u6_n2427 , _u10_u6_n2426 , _u10_u6_n2425 ,_u10_u6_n2424 , _u10_u6_n2423 , _u10_u6_n2422 , _u10_u6_n2421 ,_u10_u6_n2420 , _u10_u6_n2419 , _u10_u6_n2418 , _u10_u6_n2417 ,_u10_u6_n2416 , _u10_u6_n2415 , _u10_u6_n2414 , _u10_u6_n2413 ,_u10_u6_n2412 , _u10_u6_n2411 , _u10_u6_n2410 , _u10_u6_n2409 ,_u10_u6_n2408 , _u10_u6_n2407 , _u10_u6_n2406 , _u10_u6_n2405 ,_u10_u6_n2404 , _u10_u6_n2403 , _u10_u6_n2402 , _u10_u6_n2401 ,_u10_u6_n2400 , _u10_u6_n2399 , _u10_u6_n2398 , _u10_u6_n2397 ,_u10_u6_n2396 , _u10_u6_n2395 , _u10_u6_n2394 , _u10_u6_n2393 ,_u10_u6_n2392 , _u10_u6_n2391 , _u10_u6_n2390 , _u10_u6_n2389 ,_u10_u6_n2388 , _u10_u6_n2387 , _u10_u6_n2386 , _u10_u6_n2385 ,_u10_u6_n2384 , _u10_u6_n2383 , _u10_u6_n2382 , _u10_u6_n2381 ,_u10_u6_n2380 , _u10_u6_n2379 , _u10_u6_n2378 , _u10_u6_n2377 ,_u10_u6_n2376 , _u10_u6_n2375 , _u10_u6_n2374 , _u10_u6_n2373 ,_u10_u6_n2372 , _u10_u6_n2371 , _u10_u6_n2370 , _u10_u6_n2369 ,_u10_u6_n2368 , _u10_u6_n2367 , _u10_u6_n2366 , _u10_u6_n2365 ,_u10_u6_n2364 , _u10_u6_n2363 , _u10_u6_n2362 , _u10_u6_n2361 ,_u10_u6_n2360 , _u10_u6_n2359 , _u10_u6_n2358 , _u10_u6_n2357 ,_u10_u6_n2356 , _u10_u6_n2355 , _u10_u6_n2354 , _u10_u6_n2353 ,_u10_u6_n2352 , _u10_u6_n2351 , _u10_u6_n2350 , _u10_u6_n2349 ,_u10_u6_n2348 , _u10_u6_n2347 , _u10_u6_n2346 , _u10_u6_n2345 ,_u10_u6_n2344 , _u10_u6_n2343 , _u10_u6_n2342 , _u10_u6_n2341 ,_u10_u6_n2340 , _u10_u6_n2339 , _u10_u6_n2338 , _u10_u6_n2337 ,_u10_u6_n2336 , _u10_u6_n2335 , _u10_u6_n2334 , _u10_u6_n2333 ,_u10_u6_n2332 , _u10_u6_n2331 , _u10_u6_n2330 , _u10_u6_n2329 ,_u10_u6_n2328 , _u10_u6_n2327 , _u10_u6_n2326 , _u10_u6_n2325 ,_u10_u6_n2324 , _u10_u6_n2323 , _u10_u6_n2322 , _u10_u6_n2321 ,_u10_u6_n2320 , _u10_u6_n2319 , _u10_u6_n2318 , _u10_u6_n2317 ,_u10_u6_n2316 , _u10_u6_n2315 , _u10_u6_n2314 , _u10_u6_n2313 ,_u10_u6_n2312 , _u10_u6_n2311 , _u10_u6_n2310 , _u10_u6_n2309 ,_u10_u6_n2308 , _u10_u6_n2307 , _u10_u6_n2306 , _u10_u6_n2305 ,_u10_u6_n2304 , _u10_u6_n2303 , _u10_u6_n2302 , _u10_u6_n2301 ,_u10_u6_n2300 , _u10_u6_n2299 , _u10_u6_n2298 , _u10_u6_n2297 ,_u10_u6_n2296 , _u10_u6_n2295 , _u10_u6_n2294 , _u10_u6_n2293 ,_u10_u6_n2292 , _u10_u6_n2291 , _u10_u6_n2290 , _u10_u6_n2289 ,_u10_u6_n2288 , _u10_u6_n2287 , _u10_u6_n2286 , _u10_u6_n2285 ,_u10_u6_n2284 , _u10_u6_n2283 , _u10_u6_n2282 , _u10_u6_n2281 ,_u10_u6_n2280 , _u10_u6_n2279 , _u10_u6_n2278 , _u10_u6_n2277 ,_u10_u6_n2276 , _u10_u6_n2275 , _u10_u6_n2274 , _u10_u6_n2273 ,_u10_u6_n2272 , _u10_u6_n2271 , _u10_u6_n2270 , _u10_u6_n2269 ,_u10_u6_n2268 , _u10_u6_n2267 , _u10_u6_n2266 , _u10_u6_n2265 ,_u10_u6_n2264 , _u10_u6_n2263 , _u10_u6_n2262 , _u10_u6_n2261 ,_u10_u6_n2260 , _u10_u6_n2259 , _u10_u6_n2258 , _u10_u6_n2257 ,_u10_u6_n2256 , _u10_u6_n2255 , _u10_u6_n2254 , _u10_u6_n2253 ,_u10_u6_n2252 , _u10_u6_n2251 , _u10_u6_n2250 , _u10_u6_n2249 ,_u10_u6_n2248 , _u10_u6_n2247 , _u10_u6_n2246 , _u10_u6_n2245 ,_u10_u6_n2244 , _u10_u6_n2243 , _u10_u6_n2242 , _u10_u6_n2241 ,_u10_u6_n2240 , _u10_u6_n2239 , _u10_u6_n2238 , _u10_u6_n2237 ,_u10_u6_n2236 , _u10_u6_n2235 , _u10_u6_n2234 , _u10_u6_n2233 ,_u10_u6_n2232 , _u10_u6_n2231 , _u10_u6_n2230 , _u10_u6_n2229 ,_u10_u6_n2228 , _u10_u6_n2227 , _u10_u6_n2226 , _u10_u6_n2225 ,_u10_u6_n2224 , _u10_u6_n2223 , _u10_u6_n2222 , _u10_u6_n2221 ,_u10_u6_n2220 , _u10_u6_n2219 , _u10_u6_n2218 , _u10_u6_n2217 ,_u10_u6_n2216 , _u10_u6_n2215 , _u10_u6_n2214 , _u10_u6_n2213 ,_u10_u6_n2212 , _u10_u6_n2211 , _u10_u6_n2210 , _u10_u6_n2209 ,_u10_u6_n2208 , _u10_u6_n2207 , _u10_u6_n2206 , _u10_u6_n2205 ,_u10_u6_n2204 , _u10_u6_n2203 , _u10_u6_n2202 , _u10_u6_n2201 ,_u10_u6_n2200 , _u10_u6_n2199 , _u10_u6_n2198 , _u10_u6_n2197 ,_u10_u6_n2196 , _u10_u6_n2195 , _u10_u6_n2194 , _u10_u6_n2193 ,_u10_u6_n2192 , _u10_u6_n2191 , _u10_u6_n2190 , _u10_u6_n2189 ,_u10_u6_n2188 , _u10_u6_n2187 , _u10_u6_n2186 , _u10_u6_n2185 ,_u10_u6_n2184 , _u10_u6_n2183 , _u10_u6_n2182 , _u10_u6_n2181 ,_u10_u6_n2180 , _u10_u6_n2179 , _u10_u6_n2178 , _u10_u6_n2177 ,_u10_u6_n2176 , _u10_u6_n2175 , _u10_u6_n2174 , _u10_u6_n2173 ,_u10_u6_n2172 , _u10_u6_n2171 , _u10_u6_n2170 , _u10_u6_n2169 ,_u10_u6_n2168 , _u10_u6_n2167 , _u10_u6_n2166 , _u10_u6_n2165 ,_u10_u6_n2164 , _u10_u6_n2163 , _u10_u6_n2162 , _u10_u6_n2161 ,_u10_u6_n2160 , _u10_u6_n2159 , _u10_u6_n2158 , _u10_u6_n2157 ,_u10_u6_n2156 , _u10_u6_n2155 , _u10_u6_n2154 , _u10_u6_n2153 ,_u10_u6_n2152 , _u10_u6_n2151 , _u10_u6_n2150 , _u10_u6_n2149 ,_u10_u6_n2148 , _u10_u6_n2147 , _u10_u6_n2146 , _u10_u6_n2145 ,_u10_u6_n2144 , _u10_u6_n2143 , _u10_u6_n2142 , _u10_u6_n2141 ,_u10_u6_n2140 , _u10_u6_n2139 , _u10_u6_n2138 , _u10_u6_n2137 ,_u10_u6_n2136 , _u10_u6_n2135 , _u10_u6_n2134 , _u10_u6_n2133 ,_u10_u6_n2132 , _u10_u6_n2131 , _u10_u6_n2130 , _u10_u6_n2129 ,_u10_u6_n2128 , _u10_u6_n2127 , _u10_u6_n2126 , _u10_u6_n2125 ,_u10_u6_n2124 , _u10_u6_n2123 , _u10_u6_n2122 , _u10_u6_n2121 ,_u10_u6_n2120 , _u10_u6_n2119 , _u10_u6_n2118 , _u10_u6_n2117 ,_u10_u6_n2116 , _u10_u6_n2115 , _u10_u6_n2114 , _u10_u6_n2113 ,_u10_u6_n2112 , _u10_u6_n2111 , _u10_u6_n2110 , _u10_u6_n2109 ,_u10_u6_n2108 , _u10_u6_n2107 , _u10_u6_n2106 , _u10_u6_n2105 ,_u10_u6_n2104 , _u10_u6_n2103 , _u10_u6_n2102 , _u10_u6_n2101 ,_u10_u6_n2100 , _u10_u6_n2099 , _u10_u6_n2098 , _u10_u6_n2097 ,_u10_u6_n2096 , _u10_u6_n2095 , _u10_u6_n2094 , _u10_u6_n2093 ,_u10_u6_n2092 , _u10_u6_n2091 , _u10_u6_n2090 , _u10_u6_n2089 ,_u10_u6_n2088 , _u10_u6_n2087 , _u10_u6_n2086 , _u10_u6_n2085 ,_u10_u6_n2084 , _u10_u6_n2083 , _u10_u6_n2082 , _u10_u6_n2081 ,_u10_u6_n2080 , _u10_u6_n2079 , _u10_u6_n2078 , _u10_u6_n2077 ,_u10_u6_n2076 , _u10_u6_n2075 , _u10_u6_n2074 , _u10_u6_n2073 ,_u10_u6_n2072 , _u10_u6_n2071 , _u10_u6_n2070 , _u10_u6_n2069 ,_u10_u6_n2068 , _u10_u6_n2067 , _u10_u6_n2066 , _u10_u6_n2065 ,_u10_u6_n2064 , _u10_u6_n2063 , _u10_u6_n2062 , _u10_u6_n2061 ,_u10_u6_n2060 , _u10_u6_n2059 , _u10_u6_n2058 , _u10_u6_n2057 ,_u10_u6_n2056 , _u10_u6_n2055 , _u10_u6_n2054 , _u10_u6_n2053 ,_u10_u6_n2052 , _u10_u6_n2051 , _u10_u6_n2050 , _u10_u6_n2049 ,_u10_u6_n2048 , _u10_u6_n2047 , _u10_u6_n2046 , _u10_u6_n2045 ,_u10_u6_n2044 , _u10_u6_n2043 , _u10_u6_n2042 , _u10_u6_n2041 ,_u10_u6_n2040 , _u10_u6_n2039 , _u10_u6_n2038 , _u10_u6_n2037 ,_u10_u6_n2036 , _u10_u6_n2035 , _u10_u6_n2034 , _u10_u6_n2033 ,_u10_u6_n2032 , _u10_u6_n2031 , _u10_u6_n2030 , _u10_u6_n2029 ,_u10_u6_n2028 , _u10_u6_n2027 , _u10_u6_n2026 , _u10_u6_n2025 ,_u10_u6_n2024 , _u10_u6_n2023 , _u10_u6_n2022 , _u10_u6_n2021 ,_u10_u6_n2020 , _u10_u6_n2019 , _u10_u6_n2018 , _u10_u6_n2017 ,_u10_u6_n2016 , _u10_u6_n2015 , _u10_u6_n2014 , _u10_u6_n2013 ,_u10_u6_n2012 , _u10_u6_n2011 , _u10_u6_n2010 , _u10_u6_n2009 ,_u10_u6_n2008 , _u10_u6_n2007 , _u10_u6_n2006 , _u10_u6_n2005 ,_u10_u6_n2004 , _u10_u6_n2003 , _u10_u6_n2002 , _u10_u6_n2001 ,_u10_u6_n2000 , _u10_u6_n1999 , _u10_u6_n1998 , _u10_u6_n1997 ,_u10_u6_n1996 , _u10_u6_n1995 , _u10_u6_n1994 , _u10_u6_n1993 ,_u10_u6_n1992 , _u10_u6_n1991 , _u10_u6_n1990 , _u10_u6_n1989 ,_u10_u6_n1988 , _u10_u6_n1987 , _u10_u6_n1986 , _u10_u6_n1985 ,_u10_u6_n1984 , _u10_u6_n1983 , _u10_u6_n1982 , _u10_u6_n1981 ,_u10_u6_n1980 , _u10_u6_n1979 , _u10_u6_n1978 , _u10_u6_n1977 ,_u10_u6_n1976 , _u10_u6_n1975 , _u10_u6_n1974 , _u10_u6_n1973 ,_u10_u6_n1972 , _u10_u6_n1971 , _u10_u6_n1970 , _u10_u6_n1969 ,_u10_u6_n1968 , _u10_u6_n1967 , _u10_u6_n1966 , _u10_u6_n1965 ,_u10_u6_n1964 , _u10_u6_n1963 , _u10_u6_n1962 , _u10_u6_n1961 ,_u10_u6_n1960 , _u10_u6_n1959 , _u10_u6_n1958 , _u10_u6_n1957 ,_u10_u6_n1956 , _u10_u6_n1955 , _u10_u6_n1954 , _u10_u6_n1953 ,_u10_u6_n1952 , _u10_u6_n1951 , _u10_u6_n1950 , _u10_u6_n1949 ,_u10_u6_n1948 , _u10_u6_n1947 , _u10_u6_n1946 , _u10_u6_n1945 ,_u10_u6_n1944 , _u10_u6_n1943 , _u10_u6_n1942 , _u10_u6_n1941 ,_u10_u6_n1940 , _u10_u6_n1939 , _u10_u6_n1938 , _u10_u6_n1937 ,_u10_u6_n1936 , _u10_u6_n1935 , _u10_u6_n1934 , _u10_u6_n1933 ,_u10_u6_n1932 , _u10_u6_n1931 , _u10_u6_n1930 , _u10_u6_n1929 ,_u10_u6_n1928 , _u10_u6_n1927 , _u10_u6_n1926 , _u10_u6_n1925 ,_u10_u6_n1924 , _u10_u6_n1923 , _u10_u6_n1922 , _u10_u6_n1921 ,_u10_u6_n1920 , _u10_u6_n1919 , _u10_u6_n1918 , _u10_u6_n1917 ,_u10_u6_n1916 , _u10_u6_n1915 , _u10_u6_n1914 , _u10_u6_n1913 ,_u10_u6_n1912 , _u10_u6_n1911 , _u10_u6_n1910 , _u10_u6_n1909 ,_u10_u6_n1908 , _u10_u6_n1907 , _u10_u6_n1906 , _u10_u6_n1905 ,_u10_u6_n1904 , _u10_u6_n1903 , _u10_u6_n1902 , _u10_u6_n1901 ,_u10_u6_n1900 , _u10_u6_n1899 , _u10_u6_n1898 , _u10_u6_n1897 ,_u10_u6_n1896 , _u10_u6_n1895 , _u10_u6_n1894 , _u10_u6_n1893 ,_u10_u6_n1892 , _u10_u6_n1891 , _u10_u6_n1890 , _u10_u6_n1889 ,_u10_u6_n1888 , _u10_u6_n1887 , _u10_u6_n1886 , _u10_u6_n1885 ,_u10_u6_n1884 , _u10_u6_n1883 , _u10_u6_n1882 , _u10_u6_n1881 ,_u10_u6_n1880 , _u10_u6_n1879 , _u10_u6_n1878 , _u10_u6_n1877 ,_u10_u6_n1876 , _u10_u6_n1875 , _u10_u6_n1874 , _u10_u6_n1873 ,_u10_u6_n1872 , _u10_u6_n1871 , _u10_u6_n1870 , _u10_u6_n1869 ,_u10_u6_n1868 , _u10_u6_n1867 , _u10_u6_n1866 , _u10_u6_n1865 ,_u10_u6_n1864 , _u10_u6_n1863 , _u10_u6_n1862 , _u10_u6_n1861 ,_u10_u6_n1860 , _u10_u6_n1859 , _u10_u6_n1858 , _u10_u6_n1857 ,_u10_u6_n1856 , _u10_u6_n1855 , _u10_u6_n1854 , _u10_u6_n1853 ,_u10_u6_n1852 , _u10_u6_n1851 , _u10_u6_n1850 , _u10_u6_n1849 ,_u10_u6_n1848 , _u10_u6_n1847 , _u10_u6_n1846 , _u10_u6_n1845 ,_u10_u6_n1844 , _u10_u6_n1843 , _u10_u6_n1842 , _u10_u6_n1841 ,_u10_u6_n1840 , _u10_u6_n1839 , _u10_u6_n1838 , _u10_u6_n1837 ,_u10_u6_n1836 , _u10_u6_n1835 , _u10_u6_n1834 , _u10_u6_n1833 ,_u10_u6_n1832 , _u10_u6_n1831 , _u10_u6_n1830 , _u10_u6_n1829 ,_u10_u6_n1828 , _u10_u6_n1827 , _u10_u6_n1826 , _u10_u6_n1825 ,_u10_u6_n1824 , _u10_u6_n1823 , _u10_u6_n1822 , _u10_u6_n1821 ,_u10_u6_n1820 , _u10_u6_n1819 , _u10_u6_n1818 , _u10_u6_n1817 ,_u10_u6_n1816 , _u10_u6_n1815 , _u10_u6_n1814 , _u10_u6_n1813 ,_u10_u6_n1812 , _u10_u6_n1811 , _u10_u6_n1810 , _u10_u6_n1809 ,_u10_u6_n1808 , _u10_u7_n3416 , _u10_u7_n3415 , _u10_u7_n3414 ,_u10_u7_n3413 , _u10_u7_n3412 , _u10_u7_n3411 , _u10_u7_n3410 ,_u10_u7_n3409 , _u10_u7_n3408 , _u10_u7_n3407 , _u10_u7_n3406 ,_u10_u7_n3405 , _u10_u7_n3404 , _u10_u7_n3403 , _u10_u7_n3402 ,_u10_u7_n3401 , _u10_u7_n3400 , _u10_u7_n3399 , _u10_u7_n3398 ,_u10_u7_n3397 , _u10_u7_n3396 , _u10_u7_n3395 , _u10_u7_n3394 ,_u10_u7_n3393 , _u10_u7_n3392 , _u10_u7_n3391 , _u10_u7_n3390 ,_u10_u7_n3389 , _u10_u7_n3388 , _u10_u7_n3387 , _u10_u7_n3386 ,_u10_u7_n3385 , _u10_u7_n3384 , _u10_u7_n3383 , _u10_u7_n3382 ,_u10_u7_n3381 , _u10_u7_n3380 , _u10_u7_n3379 , _u10_u7_n3378 ,_u10_u7_n3377 , _u10_u7_n3376 , _u10_u7_n3375 , _u10_u7_n3374 ,_u10_u7_n3373 , _u10_u7_n3372 , _u10_u7_n3371 , _u10_u7_n3370 ,_u10_u7_n3369 , _u10_u7_n3368 , _u10_u7_n3367 , _u10_u7_n3366 ,_u10_u7_n3365 , _u10_u7_n3364 , _u10_u7_n3363 , _u10_u7_n3362 ,_u10_u7_n3361 , _u10_u7_n3360 , _u10_u7_n3359 , _u10_u7_n3358 ,_u10_u7_n3357 , _u10_u7_n3356 , _u10_u7_n3355 , _u10_u7_n3354 ,_u10_u7_n3353 , _u10_u7_n3352 , _u10_u7_n3351 , _u10_u7_n3350 ,_u10_u7_n3349 , _u10_u7_n3348 , _u10_u7_n3347 , _u10_u7_n3346 ,_u10_u7_n3345 , _u10_u7_n3344 , _u10_u7_n3343 , _u10_u7_n3342 ,_u10_u7_n3341 , _u10_u7_n3340 , _u10_u7_n3339 , _u10_u7_n3338 ,_u10_u7_n3337 , _u10_u7_n3336 , _u10_u7_n3335 , _u10_u7_n3334 ,_u10_u7_n3333 , _u10_u7_n3332 , _u10_u7_n3331 , _u10_u7_n3330 ,_u10_u7_n3329 , _u10_u7_n3328 , _u10_u7_n3327 , _u10_u7_n3326 ,_u10_u7_n3325 , _u10_u7_n3324 , _u10_u7_n3323 , _u10_u7_n3322 ,_u10_u7_n3321 , _u10_u7_n3320 , _u10_u7_n3319 , _u10_u7_n3318 ,_u10_u7_n3317 , _u10_u7_n3316 , _u10_u7_n3315 , _u10_u7_n3314 ,_u10_u7_n3313 , _u10_u7_n3312 , _u10_u7_n3311 , _u10_u7_n3310 ,_u10_u7_n3309 , _u10_u7_n3308 , _u10_u7_n3307 , _u10_u7_n3306 ,_u10_u7_n3305 , _u10_u7_n3304 , _u10_u7_n3303 , _u10_u7_n3302 ,_u10_u7_n3301 , _u10_u7_n3300 , _u10_u7_n3299 , _u10_u7_n3298 ,_u10_u7_n3297 , _u10_u7_n3296 , _u10_u7_n3295 , _u10_u7_n3294 ,_u10_u7_n3293 , _u10_u7_n3292 , _u10_u7_n3291 , _u10_u7_n3290 ,_u10_u7_n3289 , _u10_u7_n3288 , _u10_u7_n3287 , _u10_u7_n3286 ,_u10_u7_n3285 , _u10_u7_n3284 , _u10_u7_n3283 , _u10_u7_n3282 ,_u10_u7_n3281 , _u10_u7_n3280 , _u10_u7_n3279 , _u10_u7_n3278 ,_u10_u7_n3277 , _u10_u7_n3276 , _u10_u7_n3275 , _u10_u7_n3274 ,_u10_u7_n3273 , _u10_u7_n3272 , _u10_u7_n3271 , _u10_u7_n3270 ,_u10_u7_n3269 , _u10_u7_n3268 , _u10_u7_n3267 , _u10_u7_n3266 ,_u10_u7_n3265 , _u10_u7_n3264 , _u10_u7_n3263 , _u10_u7_n3262 ,_u10_u7_n3261 , _u10_u7_n3260 , _u10_u7_n3259 , _u10_u7_n3258 ,_u10_u7_n3257 , _u10_u7_n3256 , _u10_u7_n3255 , _u10_u7_n3254 ,_u10_u7_n3253 , _u10_u7_n3252 , _u10_u7_n3251 , _u10_u7_n3250 ,_u10_u7_n3249 , _u10_u7_n3248 , _u10_u7_n3247 , _u10_u7_n3246 ,_u10_u7_n3245 , _u10_u7_n3244 , _u10_u7_n3243 , _u10_u7_n3242 ,_u10_u7_n3241 , _u10_u7_n3240 , _u10_u7_n3239 , _u10_u7_n3238 ,_u10_u7_n3237 , _u10_u7_n3236 , _u10_u7_n3235 , _u10_u7_n3234 ,_u10_u7_n3233 , _u10_u7_n3232 , _u10_u7_n3231 , _u10_u7_n3230 ,_u10_u7_n3229 , _u10_u7_n3228 , _u10_u7_n3227 , _u10_u7_n3226 ,_u10_u7_n3225 , _u10_u7_n3224 , _u10_u7_n3223 , _u10_u7_n3222 ,_u10_u7_n3221 , _u10_u7_n3220 , _u10_u7_n3219 , _u10_u7_n3218 ,_u10_u7_n3217 , _u10_u7_n3216 , _u10_u7_n3215 , _u10_u7_n3214 ,_u10_u7_n3213 , _u10_u7_n3212 , _u10_u7_n3211 , _u10_u7_n3210 ,_u10_u7_n3209 , _u10_u7_n3208 , _u10_u7_n3207 , _u10_u7_n3206 ,_u10_u7_n3205 , _u10_u7_n3204 , _u10_u7_n3203 , _u10_u7_n3202 ,_u10_u7_n3201 , _u10_u7_n3200 , _u10_u7_n3199 , _u10_u7_n3198 ,_u10_u7_n3197 , _u10_u7_n3196 , _u10_u7_n3195 , _u10_u7_n3194 ,_u10_u7_n3193 , _u10_u7_n3192 , _u10_u7_n3191 , _u10_u7_n3190 ,_u10_u7_n3189 , _u10_u7_n3188 , _u10_u7_n3187 , _u10_u7_n3186 ,_u10_u7_n3185 , _u10_u7_n3184 , _u10_u7_n3183 , _u10_u7_n3182 ,_u10_u7_n3181 , _u10_u7_n3180 , _u10_u7_n3179 , _u10_u7_n3178 ,_u10_u7_n3177 , _u10_u7_n3176 , _u10_u7_n3175 , _u10_u7_n3174 ,_u10_u7_n3173 , _u10_u7_n3172 , _u10_u7_n3171 , _u10_u7_n3170 ,_u10_u7_n3169 , _u10_u7_n3168 , _u10_u7_n3167 , _u10_u7_n3166 ,_u10_u7_n3165 , _u10_u7_n3164 , _u10_u7_n3163 , _u10_u7_n3162 ,_u10_u7_n3161 , _u10_u7_n3160 , _u10_u7_n3159 , _u10_u7_n3158 ,_u10_u7_n3157 , _u10_u7_n3156 , _u10_u7_n3155 , _u10_u7_n3154 ,_u10_u7_n3153 , _u10_u7_n3152 , _u10_u7_n3151 , _u10_u7_n3150 ,_u10_u7_n3149 , _u10_u7_n3148 , _u10_u7_n3147 , _u10_u7_n3146 ,_u10_u7_n3145 , _u10_u7_n3144 , _u10_u7_n3143 , _u10_u7_n3142 ,_u10_u7_n3141 , _u10_u7_n3140 , _u10_u7_n3139 , _u10_u7_n3138 ,_u10_u7_n3137 , _u10_u7_n3136 , _u10_u7_n3135 , _u10_u7_n3134 ,_u10_u7_n3133 , _u10_u7_n3132 , _u10_u7_n3131 , _u10_u7_n3130 ,_u10_u7_n3129 , _u10_u7_n3128 , _u10_u7_n3127 , _u10_u7_n3126 ,_u10_u7_n3125 , _u10_u7_n3124 , _u10_u7_n3123 , _u10_u7_n3122 ,_u10_u7_n3121 , _u10_u7_n3120 , _u10_u7_n3119 , _u10_u7_n3118 ,_u10_u7_n3117 , _u10_u7_n3116 , _u10_u7_n3115 , _u10_u7_n3114 ,_u10_u7_n3113 , _u10_u7_n3112 , _u10_u7_n3111 , _u10_u7_n3110 ,_u10_u7_n3109 , _u10_u7_n3108 , _u10_u7_n3107 , _u10_u7_n3106 ,_u10_u7_n3105 , _u10_u7_n3104 , _u10_u7_n3103 , _u10_u7_n3102 ,_u10_u7_n3101 , _u10_u7_n3100 , _u10_u7_n3099 , _u10_u7_n3098 ,_u10_u7_n3097 , _u10_u7_n3096 , _u10_u7_n3095 , _u10_u7_n3094 ,_u10_u7_n3093 , _u10_u7_n3092 , _u10_u7_n3091 , _u10_u7_n3090 ,_u10_u7_n3089 , _u10_u7_n3088 , _u10_u7_n3087 , _u10_u7_n3086 ,_u10_u7_n3085 , _u10_u7_n3084 , _u10_u7_n3083 , _u10_u7_n3082 ,_u10_u7_n3081 , _u10_u7_n3080 , _u10_u7_n3079 , _u10_u7_n3078 ,_u10_u7_n3077 , _u10_u7_n3076 , _u10_u7_n3075 , _u10_u7_n3074 ,_u10_u7_n3073 , _u10_u7_n3072 , _u10_u7_n3071 , _u10_u7_n3070 ,_u10_u7_n3069 , _u10_u7_n3068 , _u10_u7_n3067 , _u10_u7_n3066 ,_u10_u7_n3065 , _u10_u7_n3064 , _u10_u7_n3063 , _u10_u7_n3062 ,_u10_u7_n3061 , _u10_u7_n3060 , _u10_u7_n3059 , _u10_u7_n3058 ,_u10_u7_n3057 , _u10_u7_n3056 , _u10_u7_n3055 , _u10_u7_n3054 ,_u10_u7_n3053 , _u10_u7_n3052 , _u10_u7_n3051 , _u10_u7_n3050 ,_u10_u7_n3049 , _u10_u7_n3048 , _u10_u7_n3047 , _u10_u7_n3046 ,_u10_u7_n3045 , _u10_u7_n3044 , _u10_u7_n3043 , _u10_u7_n3042 ,_u10_u7_n3041 , _u10_u7_n3040 , _u10_u7_n3039 , _u10_u7_n3038 ,_u10_u7_n3037 , _u10_u7_n3036 , _u10_u7_n3035 , _u10_u7_n3034 ,_u10_u7_n3033 , _u10_u7_n3032 , _u10_u7_n3031 , _u10_u7_n3030 ,_u10_u7_n3029 , _u10_u7_n3028 , _u10_u7_n3027 , _u10_u7_n3026 ,_u10_u7_n3025 , _u10_u7_n3024 , _u10_u7_n3023 , _u10_u7_n3022 ,_u10_u7_n3021 , _u10_u7_n3020 , _u10_u7_n3019 , _u10_u7_n3018 ,_u10_u7_n3017 , _u10_u7_n3016 , _u10_u7_n3015 , _u10_u7_n3014 ,_u10_u7_n3013 , _u10_u7_n3012 , _u10_u7_n3011 , _u10_u7_n3010 ,_u10_u7_n3009 , _u10_u7_n3008 , _u10_u7_n3007 , _u10_u7_n3006 ,_u10_u7_n3005 , _u10_u7_n3004 , _u10_u7_n3003 , _u10_u7_n3002 ,_u10_u7_n3001 , _u10_u7_n3000 , _u10_u7_n2999 , _u10_u7_n2998 ,_u10_u7_n2997 , _u10_u7_n2996 , _u10_u7_n2995 , _u10_u7_n2994 ,_u10_u7_n2993 , _u10_u7_n2992 , _u10_u7_n2991 , _u10_u7_n2990 ,_u10_u7_n2989 , _u10_u7_n2988 , _u10_u7_n2987 , _u10_u7_n2986 ,_u10_u7_n2985 , _u10_u7_n2984 , _u10_u7_n2983 , _u10_u7_n2982 ,_u10_u7_n2981 , _u10_u7_n2980 , _u10_u7_n2979 , _u10_u7_n2978 ,_u10_u7_n2977 , _u10_u7_n2976 , _u10_u7_n2975 , _u10_u7_n2974 ,_u10_u7_n2973 , _u10_u7_n2972 , _u10_u7_n2971 , _u10_u7_n2970 ,_u10_u7_n2969 , _u10_u7_n2968 , _u10_u7_n2967 , _u10_u7_n2966 ,_u10_u7_n2965 , _u10_u7_n2964 , _u10_u7_n2963 , _u10_u7_n2962 ,_u10_u7_n2961 , _u10_u7_n2960 , _u10_u7_n2959 , _u10_u7_n2958 ,_u10_u7_n2957 , _u10_u7_n2956 , _u10_u7_n2955 , _u10_u7_n2954 ,_u10_u7_n2953 , _u10_u7_n2952 , _u10_u7_n2951 , _u10_u7_n2950 ,_u10_u7_n2949 , _u10_u7_n2948 , _u10_u7_n2947 , _u10_u7_n2946 ,_u10_u7_n2945 , _u10_u7_n2944 , _u10_u7_n2943 , _u10_u7_n2942 ,_u10_u7_n2941 , _u10_u7_n2940 , _u10_u7_n2939 , _u10_u7_n2938 ,_u10_u7_n2937 , _u10_u7_n2936 , _u10_u7_n2935 , _u10_u7_n2934 ,_u10_u7_n2933 , _u10_u7_n2932 , _u10_u7_n2931 , _u10_u7_n2930 ,_u10_u7_n2929 , _u10_u7_n2928 , _u10_u7_n2927 , _u10_u7_n2926 ,_u10_u7_n2925 , _u10_u7_n2924 , _u10_u7_n2923 , _u10_u7_n2922 ,_u10_u7_n2921 , _u10_u7_n2920 , _u10_u7_n2919 , _u10_u7_n2918 ,_u10_u7_n2917 , _u10_u7_n2916 , _u10_u7_n2915 , _u10_u7_n2914 ,_u10_u7_n2913 , _u10_u7_n2912 , _u10_u7_n2911 , _u10_u7_n2910 ,_u10_u7_n2909 , _u10_u7_n2908 , _u10_u7_n2907 , _u10_u7_n2906 ,_u10_u7_n2905 , _u10_u7_n2904 , _u10_u7_n2903 , _u10_u7_n2902 ,_u10_u7_n2901 , _u10_u7_n2900 , _u10_u7_n2899 , _u10_u7_n2898 ,_u10_u7_n2897 , _u10_u7_n2896 , _u10_u7_n2895 , _u10_u7_n2894 ,_u10_u7_n2893 , _u10_u7_n2892 , _u10_u7_n2891 , _u10_u7_n2890 ,_u10_u7_n2889 , _u10_u7_n2888 , _u10_u7_n2887 , _u10_u7_n2886 ,_u10_u7_n2885 , _u10_u7_n2884 , _u10_u7_n2883 , _u10_u7_n2882 ,_u10_u7_n2881 , _u10_u7_n2880 , _u10_u7_n2879 , _u10_u7_n2878 ,_u10_u7_n2877 , _u10_u7_n2876 , _u10_u7_n2875 , _u10_u7_n2874 ,_u10_u7_n2873 , _u10_u7_n2872 , _u10_u7_n2871 , _u10_u7_n2870 ,_u10_u7_n2869 , _u10_u7_n2868 , _u10_u7_n2867 , _u10_u7_n2866 ,_u10_u7_n2865 , _u10_u7_n2864 , _u10_u7_n2863 , _u10_u7_n2862 ,_u10_u7_n2861 , _u10_u7_n2860 , _u10_u7_n2859 , _u10_u7_n2858 ,_u10_u7_n2857 , _u10_u7_n2856 , _u10_u7_n2855 , _u10_u7_n2854 ,_u10_u7_n2853 , _u10_u7_n2852 , _u10_u7_n2851 , _u10_u7_n2850 ,_u10_u7_n2849 , _u10_u7_n2848 , _u10_u7_n2847 , _u10_u7_n2846 ,_u10_u7_n2845 , _u10_u7_n2844 , _u10_u7_n2843 , _u10_u7_n2842 ,_u10_u7_n2841 , _u10_u7_n2840 , _u10_u7_n2839 , _u10_u7_n2838 ,_u10_u7_n2837 , _u10_u7_n2836 , _u10_u7_n2835 , _u10_u7_n2834 ,_u10_u7_n2833 , _u10_u7_n2832 , _u10_u7_n2831 , _u10_u7_n2830 ,_u10_u7_n2829 , _u10_u7_n2828 , _u10_u7_n2827 , _u10_u7_n2826 ,_u10_u7_n2825 , _u10_u7_n2824 , _u10_u7_n2823 , _u10_u7_n2822 ,_u10_u7_n2821 , _u10_u7_n2820 , _u10_u7_n2819 , _u10_u7_n2818 ,_u10_u7_n2817 , _u10_u7_n2816 , _u10_u7_n2815 , _u10_u7_n2814 ,_u10_u7_n2813 , _u10_u7_n2812 , _u10_u7_n2811 , _u10_u7_n2810 ,_u10_u7_n2809 , _u10_u7_n2808 , _u10_u7_n2807 , _u10_u7_n2806 ,_u10_u7_n2805 , _u10_u7_n2804 , _u10_u7_n2803 , _u10_u7_n2802 ,_u10_u7_n2801 , _u10_u7_n2800 , _u10_u7_n2799 , _u10_u7_n2798 ,_u10_u7_n2797 , _u10_u7_n2796 , _u10_u7_n2795 , _u10_u7_n2794 ,_u10_u7_n2793 , _u10_u7_n2792 , _u10_u7_n2791 , _u10_u7_n2790 ,_u10_u7_n2789 , _u10_u7_n2788 , _u10_u7_n2787 , _u10_u7_n2786 ,_u10_u7_n2785 , _u10_u7_n2784 , _u10_u7_n2783 , _u10_u7_n2782 ,_u10_u7_n2781 , _u10_u7_n2780 , _u10_u7_n2779 , _u10_u7_n2778 ,_u10_u7_n2777 , _u10_u7_n2776 , _u10_u7_n2775 , _u10_u7_n2774 ,_u10_u7_n2773 , _u10_u7_n2772 , _u10_u7_n2771 , _u10_u7_n2770 ,_u10_u7_n2769 , _u10_u7_n2768 , _u10_u7_n2767 , _u10_u7_n2766 ,_u10_u7_n2765 , _u10_u7_n2764 , _u10_u7_n2763 , _u10_u7_n2762 ,_u10_u7_n2761 , _u10_u7_n2760 , _u10_u7_n2759 , _u10_u7_n2758 ,_u10_u7_n2757 , _u10_u7_n2756 , _u10_u7_n2755 , _u10_u7_n2754 ,_u10_u7_n2753 , _u10_u7_n2752 , _u10_u7_n2751 , _u10_u7_n2750 ,_u10_u7_n2749 , _u10_u7_n2748 , _u10_u7_n2747 , _u10_u7_n2746 ,_u10_u7_n2745 , _u10_u7_n2744 , _u10_u7_n2743 , _u10_u7_n2742 ,_u10_u7_n2741 , _u10_u7_n2740 , _u10_u7_n2739 , _u10_u7_n2738 ,_u10_u7_n2737 , _u10_u7_n2736 , _u10_u7_n2735 , _u10_u7_n2734 ,_u10_u7_n2733 , _u10_u7_n2732 , _u10_u7_n2731 , _u10_u7_n2730 ,_u10_u7_n2729 , _u10_u7_n2728 , _u10_u7_n2727 , _u10_u7_n2726 ,_u10_u7_n2725 , _u10_u7_n2724 , _u10_u7_n2723 , _u10_u7_n2722 ,_u10_u7_n2721 , _u10_u7_n2720 , _u10_u7_n2719 , _u10_u7_n2718 ,_u10_u7_n2717 , _u10_u7_n2716 , _u10_u7_n2715 , _u10_u7_n2714 ,_u10_u7_n2713 , _u10_u7_n2712 , _u10_u7_n2711 , _u10_u7_n2710 ,_u10_u7_n2709 , _u10_u7_n2708 , _u10_u7_n2707 , _u10_u7_n2706 ,_u10_u7_n2705 , _u10_u7_n2704 , _u10_u7_n2703 , _u10_u7_n2702 ,_u10_u7_n2701 , _u10_u7_n2700 , _u10_u7_n2699 , _u10_u7_n2698 ,_u10_u7_n2697 , _u10_u7_n2696 , _u10_u7_n2695 , _u10_u7_n2694 ,_u10_u7_n2693 , _u10_u7_n2692 , _u10_u7_n2691 , _u10_u7_n2690 ,_u10_u7_n2689 , _u10_u7_n2688 , _u10_u7_n2687 , _u10_u7_n2686 ,_u10_u7_n2685 , _u10_u7_n2684 , _u10_u7_n2683 , _u10_u7_n2682 ,_u10_u7_n2681 , _u10_u7_n2680 , _u10_u7_n2679 , _u10_u7_n2678 ,_u10_u7_n2677 , _u10_u7_n2676 , _u10_u7_n2675 , _u10_u7_n2674 ,_u10_u7_n2673 , _u10_u7_n2672 , _u10_u7_n2671 , _u10_u7_n2670 ,_u10_u7_n2669 , _u10_u7_n2668 , _u10_u7_n2667 , _u10_u7_n2666 ,_u10_u7_n2665 , _u10_u7_n2664 , _u10_u7_n2663 , _u10_u7_n2662 ,_u10_u7_n2661 , _u10_u7_n2660 , _u10_u7_n2659 , _u10_u7_n2658 ,_u10_u7_n2657 , _u10_u7_n2656 , _u10_u7_n2655 , _u10_u7_n2654 ,_u10_u7_n2653 , _u10_u7_n2652 , _u10_u7_n2651 , _u10_u7_n2650 ,_u10_u7_n2649 , _u10_u7_n2648 , _u10_u7_n2647 , _u10_u7_n2646 ,_u10_u7_n2645 , _u10_u7_n2644 , _u10_u7_n2643 , _u10_u7_n2642 ,_u10_u7_n2641 , _u10_u7_n2640 , _u10_u7_n2639 , _u10_u7_n2638 ,_u10_u7_n2637 , _u10_u7_n2636 , _u10_u7_n2635 , _u10_u7_n2634 ,_u10_u7_n2633 , _u10_u7_n2632 , _u10_u7_n2631 , _u10_u7_n2630 ,_u10_u7_n2629 , _u10_u7_n2628 , _u10_u7_n2627 , _u10_u7_n2626 ,_u10_u7_n2625 , _u10_u7_n2624 , _u10_u7_n2623 , _u10_u7_n2622 ,_u10_u7_n2621 , _u10_u7_n2620 , _u10_u7_n2619 , _u10_u7_n2618 ,_u10_u7_n2617 , _u10_u7_n2616 , _u10_u7_n2615 , _u10_u7_n2614 ,_u10_u7_n2613 , _u10_u7_n2612 , _u10_u7_n2611 , _u10_u7_n2610 ,_u10_u7_n2609 , _u10_u7_n2608 , _u10_u7_n2607 , _u10_u7_n2606 ,_u10_u7_n2605 , _u10_u7_n2604 , _u10_u7_n2603 , _u10_u7_n2602 ,_u10_u7_n2601 , _u10_u7_n2600 , _u10_u7_n2599 , _u10_u7_n2598 ,_u10_u7_n2597 , _u10_u7_n2596 , _u10_u7_n2595 , _u10_u7_n2594 ,_u10_u7_n2593 , _u10_u7_n2592 , _u10_u7_n2591 , _u10_u7_n2590 ,_u10_u7_n2589 , _u10_u7_n2588 , _u10_u7_n2587 , _u10_u7_n2586 ,_u10_u7_n2585 , _u10_u7_n2584 , _u10_u7_n2583 , _u10_u7_n2582 ,_u10_u7_n2581 , _u10_u7_n2580 , _u10_u7_n2579 , _u10_u7_n2578 ,_u10_u7_n2577 , _u10_u7_n2576 , _u10_u7_n2575 , _u10_u7_n2574 ,_u10_u7_n2573 , _u10_u7_n2572 , _u10_u7_n2571 , _u10_u7_n2570 ,_u10_u7_n2569 , _u10_u7_n2568 , _u10_u7_n2567 , _u10_u7_n2566 ,_u10_u7_n2565 , _u10_u7_n2564 , _u10_u7_n2563 , _u10_u7_n2562 ,_u10_u7_n2561 , _u10_u7_n2560 , _u10_u7_n2559 , _u10_u7_n2558 ,_u10_u7_n2557 , _u10_u7_n2556 , _u10_u7_n2555 , _u10_u7_n2554 ,_u10_u7_n2553 , _u10_u7_n2552 , _u10_u7_n2551 , _u10_u7_n2550 ,_u10_u7_n2549 , _u10_u7_n2548 , _u10_u7_n2547 , _u10_u7_n2546 ,_u10_u7_n2545 , _u10_u7_n2544 , _u10_u7_n2543 , _u10_u7_n2542 ,_u10_u7_n2541 , _u10_u7_n2540 , _u10_u7_n2539 , _u10_u7_n2538 ,_u10_u7_n2537 , _u10_u7_n2536 , _u10_u7_n2535 , _u10_u7_n2534 ,_u10_u7_n2533 , _u10_u7_n2532 , _u10_u7_n2531 , _u10_u7_n2530 ,_u10_u7_n2529 , _u10_u7_n2528 , _u10_u7_n2527 , _u10_u7_n2526 ,_u10_u7_n2525 , _u10_u7_n2524 , _u10_u7_n2523 , _u10_u7_n2522 ,_u10_u7_n2521 , _u10_u7_n2520 , _u10_u7_n2519 , _u10_u7_n2518 ,_u10_u7_n2517 , _u10_u7_n2516 , _u10_u7_n2515 , _u10_u7_n2514 ,_u10_u7_n2513 , _u10_u7_n2512 , _u10_u7_n2511 , _u10_u7_n2510 ,_u10_u7_n2509 , _u10_u7_n2508 , _u10_u7_n2507 , _u10_u7_n2506 ,_u10_u7_n2505 , _u10_u7_n2504 , _u10_u7_n2503 , _u10_u7_n2502 ,_u10_u7_n2501 , _u10_u7_n2500 , _u10_u7_n2499 , _u10_u7_n2498 ,_u10_u7_n2497 , _u10_u7_n2496 , _u10_u7_n2495 , _u10_u7_n2494 ,_u10_u7_n2493 , _u10_u7_n2492 , _u10_u7_n2491 , _u10_u7_n2490 ,_u10_u7_n2489 , _u10_u7_n2488 , _u10_u7_n2487 , _u10_u7_n2486 ,_u10_u7_n2485 , _u10_u7_n2484 , _u10_u7_n2483 , _u10_u7_n2482 ,_u10_u7_n2481 , _u10_u7_n2480 , _u10_u7_n2479 , _u10_u7_n2478 ,_u10_u7_n2477 , _u10_u7_n2476 , _u10_u7_n2475 , _u10_u7_n2474 ,_u10_u7_n2473 , _u10_u7_n2472 , _u10_u7_n2471 , _u10_u7_n2470 ,_u10_u7_n2469 , _u10_u7_n2468 , _u10_u7_n2467 , _u10_u7_n2466 ,_u10_u7_n2465 , _u10_u7_n2464 , _u10_u7_n2463 , _u10_u7_n2462 ,_u10_u7_n2461 , _u10_u7_n2460 , _u10_u7_n2459 , _u10_u7_n2458 ,_u10_u7_n2457 , _u10_u7_n2456 , _u10_u7_n2455 , _u10_u7_n2454 ,_u10_u7_n2453 , _u10_u7_n2452 , _u10_u7_n2451 , _u10_u7_n2450 ,_u10_u7_n2449 , _u10_u7_n2448 , _u10_u7_n2447 , _u10_u7_n2446 ,_u10_u7_n2445 , _u10_u7_n2444 , _u10_u7_n2443 , _u10_u7_n2442 ,_u10_u7_n2441 , _u10_u7_n2440 , _u10_u7_n2439 , _u10_u7_n2438 ,_u10_u7_n2437 , _u10_u7_n2436 , _u10_u7_n2435 , _u10_u7_n2434 ,_u10_u7_n2433 , _u10_u7_n2432 , _u10_u7_n2431 , _u10_u7_n2430 ,_u10_u7_n2429 , _u10_u7_n2428 , _u10_u7_n2427 , _u10_u7_n2426 ,_u10_u7_n2425 , _u10_u7_n2424 , _u10_u7_n2423 , _u10_u7_n2422 ,_u10_u7_n2421 , _u10_u7_n2420 , _u10_u7_n2419 , _u10_u7_n2418 ,_u10_u7_n2417 , _u10_u7_n2416 , _u10_u7_n2415 , _u10_u7_n2414 ,_u10_u7_n2413 , _u10_u7_n2412 , _u10_u7_n2411 , _u10_u7_n2410 ,_u10_u7_n2409 , _u10_u7_n2408 , _u10_u7_n2407 , _u10_u7_n2406 ,_u10_u7_n2405 , _u10_u7_n2404 , _u10_u7_n2403 , _u10_u7_n2402 ,_u10_u7_n2401 , _u10_u7_n2400 , _u10_u7_n2399 , _u10_u7_n2398 ,_u10_u7_n2397 , _u10_u7_n2396 , _u10_u7_n2395 , _u10_u7_n2394 ,_u10_u7_n2393 , _u10_u7_n2392 , _u10_u7_n2391 , _u10_u7_n2390 ,_u10_u7_n2389 , _u10_u7_n2388 , _u10_u7_n2387 , _u10_u7_n2386 ,_u10_u7_n2385 , _u10_u7_n2384 , _u10_u7_n2383 , _u10_u7_n2382 ,_u10_u7_n2381 , _u10_u7_n2380 , _u10_u7_n2379 , _u10_u7_n2378 ,_u10_u7_n2377 , _u10_u7_n2376 , _u10_u7_n2375 , _u10_u7_n2374 ,_u10_u7_n2373 , _u10_u7_n2372 , _u10_u7_n2371 , _u10_u7_n2370 ,_u10_u7_n2369 , _u10_u7_n2368 , _u10_u7_n2367 , _u10_u7_n2366 ,_u10_u7_n2365 , _u10_u7_n2364 , _u10_u7_n2363 , _u10_u7_n2362 ,_u10_u7_n2361 , _u10_u7_n2360 , _u10_u7_n2359 , _u10_u7_n2358 ,_u10_u7_n2357 , _u10_u7_n2356 , _u10_u7_n2355 , _u10_u7_n2354 ,_u10_u7_n2353 , _u10_u7_n2352 , _u10_u7_n2351 , _u10_u7_n2350 ,_u10_u7_n2349 , _u10_u7_n2348 , _u10_u7_n2347 , _u10_u7_n2346 ,_u10_u7_n2345 , _u10_u7_n2344 , _u10_u7_n2343 , _u10_u7_n2342 ,_u10_u7_n2341 , _u10_u7_n2340 , _u10_u7_n2339 , _u10_u7_n2338 ,_u10_u7_n2337 , _u10_u7_n2336 , _u10_u7_n2335 , _u10_u7_n2334 ,_u10_u7_n2333 , _u10_u7_n2332 , _u10_u7_n2331 , _u10_u7_n2330 ,_u10_u7_n2329 , _u10_u7_n2328 , _u10_u7_n2327 , _u10_u7_n2326 ,_u10_u7_n2325 , _u10_u7_n2324 , _u10_u7_n2323 , _u10_u7_n2322 ,_u10_u7_n2321 , _u10_u7_n2320 , _u10_u7_n2319 , _u10_u7_n2318 ,_u10_u7_n2317 , _u10_u7_n2316 , _u10_u7_n2315 , _u10_u7_n2314 ,_u10_u7_n2313 , _u10_u7_n2312 , _u10_u7_n2311 , _u10_u7_n2310 ,_u10_u7_n2309 , _u10_u7_n2308 , _u10_u7_n2307 , _u10_u7_n2306 ,_u10_u7_n2305 , _u10_u7_n2304 , _u10_u7_n2303 , _u10_u7_n2302 ,_u10_u7_n2301 , _u10_u7_n2300 , _u10_u7_n2299 , _u10_u7_n2298 ,_u10_u7_n2297 , _u10_u7_n2296 , _u10_u7_n2295 , _u10_u7_n2294 ,_u10_u7_n2293 , _u10_u7_n2292 , _u10_u7_n2291 , _u10_u7_n2290 ,_u10_u7_n2289 , _u10_u7_n2288 , _u10_u7_n2287 , _u10_u7_n2286 ,_u10_u7_n2285 , _u10_u7_n2284 , _u10_u7_n2283 , _u10_u7_n2282 ,_u10_u7_n2281 , _u10_u7_n2280 , _u10_u7_n2279 , _u10_u7_n2278 ,_u10_u7_n2277 , _u10_u7_n2276 , _u10_u7_n2275 , _u10_u7_n2274 ,_u10_u7_n2273 , _u10_u7_n2272 , _u10_u7_n2271 , _u10_u7_n2270 ,_u10_u7_n2269 , _u10_u7_n2268 , _u10_u7_n2267 , _u10_u7_n2266 ,_u10_u7_n2265 , _u10_u7_n2264 , _u10_u7_n2263 , _u10_u7_n2262 ,_u10_u7_n2261 , _u10_u7_n2260 , _u10_u7_n2259 , _u10_u7_n2258 ,_u10_u7_n2257 , _u10_u7_n2256 , _u10_u7_n2255 , _u10_u7_n2254 ,_u10_u7_n2253 , _u10_u7_n2252 , _u10_u7_n2251 , _u10_u7_n2250 ,_u10_u7_n2249 , _u10_u7_n2248 , _u10_u7_n2247 , _u10_u7_n2246 ,_u10_u7_n2245 , _u10_u7_n2244 , _u10_u7_n2243 , _u10_u7_n2242 ,_u10_u7_n2241 , _u10_u7_n2240 , _u10_u7_n2239 , _u10_u7_n2238 ,_u10_u7_n2237 , _u10_u7_n2236 , _u10_u7_n2235 , _u10_u7_n2234 ,_u10_u7_n2233 , _u10_u7_n2232 , _u10_u7_n2231 , _u10_u7_n2230 ,_u10_u7_n2229 , _u10_u7_n2228 , _u10_u7_n2227 , _u10_u7_n2226 ,_u10_u7_n2225 , _u10_u7_n2224 , _u10_u7_n2223 , _u10_u7_n2222 ,_u10_u7_n2221 , _u10_u7_n2220 , _u10_u7_n2219 , _u10_u7_n2218 ,_u10_u7_n2217 , _u10_u7_n2216 , _u10_u7_n2215 , _u10_u7_n2214 ,_u10_u7_n2213 , _u10_u7_n2212 , _u10_u7_n2211 , _u10_u7_n2210 ,_u10_u7_n2209 , _u10_u7_n2208 , _u10_u7_n2207 , _u10_u7_n2206 ,_u10_u7_n2205 , _u10_u7_n2204 , _u10_u7_n2203 , _u10_u7_n2202 ,_u10_u7_n2201 , _u10_u7_n2200 , _u10_u7_n2199 , _u10_u7_n2198 ,_u10_u7_n2197 , _u10_u7_n2196 , _u10_u7_n2195 , _u10_u7_n2194 ,_u10_u7_n2193 , _u10_u7_n2192 , _u10_u7_n2191 , _u10_u7_n2190 ,_u10_u7_n2189 , _u10_u7_n2188 , _u10_u7_n2187 , _u10_u7_n2186 ,_u10_u7_n2185 , _u10_u7_n2184 , _u10_u7_n2183 , _u10_u7_n2182 ,_u10_u7_n2181 , _u10_u7_n2180 , _u10_u7_n2179 , _u10_u7_n2178 ,_u10_u7_n2177 , _u10_u7_n2176 , _u10_u7_n2175 , _u10_u7_n2174 ,_u10_u7_n2173 , _u10_u7_n2172 , _u10_u7_n2171 , _u10_u7_n2170 ,_u10_u7_n2169 , _u10_u7_n2168 , _u10_u7_n2167 , _u10_u7_n2166 ,_u10_u7_n2165 , _u10_u7_n2164 , _u10_u7_n2163 , _u10_u7_n2162 ,_u10_u7_n2161 , _u10_u7_n2160 , _u10_u7_n2159 , _u10_u7_n2158 ,_u10_u7_n2157 , _u10_u7_n2156 , _u10_u7_n2155 , _u10_u7_n2154 ,_u10_u7_n2153 , _u10_u7_n2152 , _u10_u7_n2151 , _u10_u7_n2150 ,_u10_u7_n2149 , _u10_u7_n2148 , _u10_u7_n2147 , _u10_u7_n2146 ,_u10_u7_n2145 , _u10_u7_n2144 , _u10_u7_n2143 , _u10_u7_n2142 ,_u10_u7_n2141 , _u10_u7_n2140 , _u10_u7_n2139 , _u10_u7_n2138 ,_u10_u7_n2137 , _u10_u7_n2136 , _u10_u7_n2135 , _u10_u7_n2134 ,_u10_u7_n2133 , _u10_u7_n2132 , _u10_u7_n2131 , _u10_u7_n2130 ,_u10_u7_n2129 , _u10_u7_n2128 , _u10_u7_n2127 , _u10_u7_n2126 ,_u10_u7_n2125 , _u10_u7_n2124 , _u10_u7_n2123 , _u10_u7_n2122 ,_u10_u7_n2121 , _u10_u7_n2120 , _u10_u7_n2119 , _u10_u7_n2118 ,_u10_u7_n2117 , _u10_u7_n2116 , _u10_u7_n2115 , _u10_u7_n2114 ,_u10_u7_n2113 , _u10_u7_n2112 , _u10_u7_n2111 , _u10_u7_n2110 ,_u10_u7_n2109 , _u10_u7_n2108 , _u10_u7_n2107 , _u10_u7_n2106 ,_u10_u7_n2105 , _u10_u7_n2104 , _u10_u7_n2103 , _u10_u7_n2102 ,_u10_u7_n2101 , _u10_u7_n2100 , _u10_u7_n2099 , _u10_u7_n2098 ,_u10_u7_n2097 , _u10_u7_n2096 , _u10_u7_n2095 , _u10_u7_n2094 ,_u10_u7_n2093 , _u10_u7_n2092 , _u10_u7_n2091 , _u10_u7_n2090 ,_u10_u7_n2089 , _u10_u7_n2088 , _u10_u7_n2087 , _u10_u7_n2086 ,_u10_u7_n2085 , _u10_u7_n2084 , _u10_u7_n2083 , _u10_u7_n2082 ,_u10_u7_n2081 , _u10_u7_n2080 , _u10_u7_n2079 , _u10_u7_n2078 ,_u10_u7_n2077 , _u10_u7_n2076 , _u10_u7_n2075 , _u10_u7_n2074 ,_u10_u7_n2073 , _u10_u7_n2072 , _u10_u7_n2071 , _u10_u7_n2070 ,_u10_u7_n2069 , _u10_u7_n2068 , _u10_u7_n2067 , _u10_u7_n2066 ,_u10_u7_n2065 , _u10_u7_n2064 , _u10_u7_n2063 , _u10_u7_n2062 ,_u10_u7_n2061 , _u10_u7_n2060 , _u10_u7_n2059 , _u10_u7_n2058 ,_u10_u7_n2057 , _u10_u7_n2056 , _u10_u7_n2055 , _u10_u7_n2054 ,_u10_u7_n2053 , _u10_u7_n2052 , _u10_u7_n2051 , _u10_u7_n2050 ,_u10_u7_n2049 , _u10_u7_n2048 , _u10_u7_n2047 , _u10_u7_n2046 ,_u10_u7_n2045 , _u10_u7_n2044 , _u10_u7_n2043 , _u10_u7_n2042 ,_u10_u7_n2041 , _u10_u7_n2040 , _u10_u7_n2039 , _u10_u7_n2038 ,_u10_u7_n2037 , _u10_u7_n2036 , _u10_u7_n2035 , _u10_u7_n2034 ,_u10_u7_n2033 , _u10_u7_n2032 , _u10_u7_n2031 , _u10_u7_n2030 ,_u10_u7_n2029 , _u10_u7_n2028 , _u10_u7_n2027 , _u10_u7_n2026 ,_u10_u7_n2025 , _u10_u7_n2024 , _u10_u7_n2023 , _u10_u7_n2022 ,_u10_u7_n2021 , _u10_u7_n2020 , _u10_u7_n2019 , _u10_u7_n2018 ,_u10_u7_n2017 , _u10_u7_n2016 , _u10_u7_n2015 , _u10_u7_n2014 ,_u10_u7_n2013 , _u10_u7_n2012 , _u10_u7_n2011 , _u10_u7_n2010 ,_u10_u7_n2009 , _u10_u7_n2008 , _u10_u7_n2007 , _u10_u7_n2006 ,_u10_u7_n2005 , _u10_u7_n2004 , _u10_u7_n2003 , _u10_u7_n2002 ,_u10_u7_n2001 , _u10_u7_n2000 , _u10_u7_n1999 , _u10_u7_n1998 ,_u10_u7_n1997 , _u10_u7_n1996 , _u10_u7_n1995 , _u10_u7_n1994 ,_u10_u7_n1993 , _u10_u7_n1992 , _u10_u7_n1991 , _u10_u7_n1990 ,_u10_u7_n1989 , _u10_u7_n1988 , _u10_u7_n1987 , _u10_u7_n1986 ,_u10_u7_n1985 , _u10_u7_n1984 , _u10_u7_n1983 , _u10_u7_n1982 ,_u10_u7_n1981 , _u10_u7_n1980 , _u10_u7_n1979 , _u10_u7_n1978 ,_u10_u7_n1977 , _u10_u7_n1976 , _u10_u7_n1975 , _u10_u7_n1974 ,_u10_u7_n1973 , _u10_u7_n1972 , _u10_u7_n1971 , _u10_u7_n1970 ,_u10_u7_n1969 , _u10_u7_n1968 , _u10_u7_n1967 , _u10_u7_n1966 ,_u10_u7_n1965 , _u10_u7_n1964 , _u10_u7_n1963 , _u10_u7_n1962 ,_u10_u7_n1961 , _u10_u7_n1960 , _u10_u7_n1959 , _u10_u7_n1958 ,_u10_u7_n1957 , _u10_u7_n1956 , _u10_u7_n1955 , _u10_u7_n1954 ,_u10_u7_n1953 , _u10_u7_n1952 , _u10_u7_n1951 , _u10_u7_n1950 ,_u10_u7_n1949 , _u10_u7_n1948 , _u10_u7_n1947 , _u10_u7_n1946 ,_u10_u7_n1945 , _u10_u7_n1944 , _u10_u7_n1943 , _u10_u7_n1942 ,_u10_u7_n1941 , _u10_u7_n1940 , _u10_u7_n1939 , _u10_u7_n1938 ,_u10_u7_n1937 , _u10_u7_n1936 , _u10_u7_n1935 , _u10_u7_n1934 ,_u10_u7_n1933 , _u10_u7_n1932 , _u10_u7_n1931 , _u10_u7_n1930 ,_u10_u7_n1929 , _u10_u7_n1928 , _u10_u7_n1927 , _u10_u7_n1926 ,_u10_u7_n1925 , _u10_u7_n1924 , _u10_u7_n1923 , _u10_u7_n1922 ,_u10_u7_n1921 , _u10_u7_n1920 , _u10_u7_n1919 , _u10_u7_n1918 ,_u10_u7_n1917 , _u10_u7_n1916 , _u10_u7_n1915 , _u10_u7_n1914 ,_u10_u7_n1913 , _u10_u7_n1912 , _u10_u7_n1911 , _u10_u7_n1910 ,_u10_u7_n1909 , _u10_u7_n1908 , _u10_u7_n1907 , _u10_u7_n1906 ,_u10_u7_n1905 , _u10_u7_n1904 , _u10_u7_n1903 , _u10_u7_n1902 ,_u10_u7_n1901 , _u10_u7_n1900 , _u10_u7_n1899 , _u10_u7_n1898 ,_u10_u7_n1897 , _u10_u7_n1896 , _u10_u7_n1895 , _u10_u7_n1894 ,_u10_u7_n1893 , _u10_u7_n1892 , _u10_u7_n1891 , _u10_u7_n1890 ,_u10_u7_n1889 , _u10_u7_n1888 , _u10_u7_n1887 , _u10_u7_n1886 ,_u10_u7_n1885 , _u10_u7_n1884 , _u10_u7_n1883 , _u10_u7_n1882 ,_u10_u7_n1881 , _u10_u7_n1880 , _u10_u7_n1879 , _u10_u7_n1878 ,_u10_u7_n1877 , _u10_u7_n1876 , _u10_u7_n1875 , _u10_u7_n1874 ,_u10_u7_n1873 , _u10_u7_n1872 , _u10_u7_n1871 , _u10_u7_n1870 ,_u10_u7_n1869 , _u10_u7_n1868 , _u10_u7_n1867 , _u10_u7_n1866 ,_u10_u7_n1865 , _u10_u7_n1864 , _u10_u7_n1863 , _u10_u7_n1862 ,_u10_u7_n1861 , _u10_u7_n1860 , _u10_u7_n1859 , _u10_u7_n1858 ,_u10_u7_n1857 , _u10_u7_n1856 , _u10_u7_n1855 , _u10_u7_n1854 ,_u10_u7_n1853 , _u10_u7_n1852 , _u10_u7_n1851 , _u10_u7_n1850 ,_u10_u7_n1849 , _u10_u7_n1848 , _u10_u7_n1847 , _u10_u7_n1846 ,_u10_u7_n1845 , _u10_u7_n1844 , _u10_u7_n1843 , _u10_u7_n1842 ,_u10_u7_n1841 , _u10_u7_n1840 , _u10_u7_n1839 , _u10_u7_n1838 ,_u10_u7_n1837 , _u10_u7_n1836 , _u10_u7_n1835 , _u10_u7_n1834 ,_u10_u7_n1833 , _u10_u7_n1832 , _u10_u7_n1831 , _u10_u7_n1830 ,_u10_u7_n1829 , _u10_u7_n1828 , _u10_u7_n1827 , _u10_u7_n1826 ,_u10_u7_n1825 , _u10_u7_n1824 , _u10_u7_n1823 , _u10_u7_n1822 ,_u10_u7_n1821 , _u10_u7_n1820 , _u10_u7_n1819 , _u10_u7_n1818 ,_u10_u7_n1817 , _u10_u7_n1816 , _u10_u7_n1815 , _u10_u7_n1814 ,_u10_u7_n1813 , _u10_u7_n1812 , _u10_u7_n1811 , _u10_u7_n1810 ,_u10_u7_n1809 , _u10_u7_n1808 , _u10_u8_n3416 , _u10_u8_n3415 ,_u10_u8_n3414 , _u10_u8_n3413 , _u10_u8_n3412 , _u10_u8_n3411 ,_u10_u8_n3410 , _u10_u8_n3409 , _u10_u8_n3408 , _u10_u8_n3407 ,_u10_u8_n3406 , _u10_u8_n3405 , _u10_u8_n3404 , _u10_u8_n3403 ,_u10_u8_n3402 , _u10_u8_n3401 , _u10_u8_n3400 , _u10_u8_n3399 ,_u10_u8_n3398 , _u10_u8_n3397 , _u10_u8_n3396 , _u10_u8_n3395 ,_u10_u8_n3394 , _u10_u8_n3393 , _u10_u8_n3392 , _u10_u8_n3391 ,_u10_u8_n3390 , _u10_u8_n3389 , _u10_u8_n3388 , _u10_u8_n3387 ,_u10_u8_n3386 , _u10_u8_n3385 , _u10_u8_n3384 , _u10_u8_n3383 ,_u10_u8_n3382 , _u10_u8_n3381 , _u10_u8_n3380 , _u10_u8_n3379 ,_u10_u8_n3378 , _u10_u8_n3377 , _u10_u8_n3376 , _u10_u8_n3375 ,_u10_u8_n3374 , _u10_u8_n3373 , _u10_u8_n3372 , _u10_u8_n3371 ,_u10_u8_n3370 , _u10_u8_n3369 , _u10_u8_n3368 , _u10_u8_n3367 ,_u10_u8_n3366 , _u10_u8_n3365 , _u10_u8_n3364 , _u10_u8_n3363 ,_u10_u8_n3362 , _u10_u8_n3361 , _u10_u8_n3360 , _u10_u8_n3359 ,_u10_u8_n3358 , _u10_u8_n3357 , _u10_u8_n3356 , _u10_u8_n3355 ,_u10_u8_n3354 , _u10_u8_n3353 , _u10_u8_n3352 , _u10_u8_n3351 ,_u10_u8_n3350 , _u10_u8_n3349 , _u10_u8_n3348 , _u10_u8_n3347 ,_u10_u8_n3346 , _u10_u8_n3345 , _u10_u8_n3344 , _u10_u8_n3343 ,_u10_u8_n3342 , _u10_u8_n3341 , _u10_u8_n3340 , _u10_u8_n3339 ,_u10_u8_n3338 , _u10_u8_n3337 , _u10_u8_n3336 , _u10_u8_n3335 ,_u10_u8_n3334 , _u10_u8_n3333 , _u10_u8_n3332 , _u10_u8_n3331 ,_u10_u8_n3330 , _u10_u8_n3329 , _u10_u8_n3328 , _u10_u8_n3327 ,_u10_u8_n3326 , _u10_u8_n3325 , _u10_u8_n3324 , _u10_u8_n3323 ,_u10_u8_n3322 , _u10_u8_n3321 , _u10_u8_n3320 , _u10_u8_n3319 ,_u10_u8_n3318 , _u10_u8_n3317 , _u10_u8_n3316 , _u10_u8_n3315 ,_u10_u8_n3314 , _u10_u8_n3313 , _u10_u8_n3312 , _u10_u8_n3311 ,_u10_u8_n3310 , _u10_u8_n3309 , _u10_u8_n3308 , _u10_u8_n3307 ,_u10_u8_n3306 , _u10_u8_n3305 , _u10_u8_n3304 , _u10_u8_n3303 ,_u10_u8_n3302 , _u10_u8_n3301 , _u10_u8_n3300 , _u10_u8_n3299 ,_u10_u8_n3298 , _u10_u8_n3297 , _u10_u8_n3296 , _u10_u8_n3295 ,_u10_u8_n3294 , _u10_u8_n3293 , _u10_u8_n3292 , _u10_u8_n3291 ,_u10_u8_n3290 , _u10_u8_n3289 , _u10_u8_n3288 , _u10_u8_n3287 ,_u10_u8_n3286 , _u10_u8_n3285 , _u10_u8_n3284 , _u10_u8_n3283 ,_u10_u8_n3282 , _u10_u8_n3281 , _u10_u8_n3280 , _u10_u8_n3279 ,_u10_u8_n3278 , _u10_u8_n3277 , _u10_u8_n3276 , _u10_u8_n3275 ,_u10_u8_n3274 , _u10_u8_n3273 , _u10_u8_n3272 , _u10_u8_n3271 ,_u10_u8_n3270 , _u10_u8_n3269 , _u10_u8_n3268 , _u10_u8_n3267 ,_u10_u8_n3266 , _u10_u8_n3265 , _u10_u8_n3264 , _u10_u8_n3263 ,_u10_u8_n3262 , _u10_u8_n3261 , _u10_u8_n3260 , _u10_u8_n3259 ,_u10_u8_n3258 , _u10_u8_n3257 , _u10_u8_n3256 , _u10_u8_n3255 ,_u10_u8_n3254 , _u10_u8_n3253 , _u10_u8_n3252 , _u10_u8_n3251 ,_u10_u8_n3250 , _u10_u8_n3249 , _u10_u8_n3248 , _u10_u8_n3247 ,_u10_u8_n3246 , _u10_u8_n3245 , _u10_u8_n3244 , _u10_u8_n3243 ,_u10_u8_n3242 , _u10_u8_n3241 , _u10_u8_n3240 , _u10_u8_n3239 ,_u10_u8_n3238 , _u10_u8_n3237 , _u10_u8_n3236 , _u10_u8_n3235 ,_u10_u8_n3234 , _u10_u8_n3233 , _u10_u8_n3232 , _u10_u8_n3231 ,_u10_u8_n3230 , _u10_u8_n3229 , _u10_u8_n3228 , _u10_u8_n3227 ,_u10_u8_n3226 , _u10_u8_n3225 , _u10_u8_n3224 , _u10_u8_n3223 ,_u10_u8_n3222 , _u10_u8_n3221 , _u10_u8_n3220 , _u10_u8_n3219 ,_u10_u8_n3218 , _u10_u8_n3217 , _u10_u8_n3216 , _u10_u8_n3215 ,_u10_u8_n3214 , _u10_u8_n3213 , _u10_u8_n3212 , _u10_u8_n3211 ,_u10_u8_n3210 , _u10_u8_n3209 , _u10_u8_n3208 , _u10_u8_n3207 ,_u10_u8_n3206 , _u10_u8_n3205 , _u10_u8_n3204 , _u10_u8_n3203 ,_u10_u8_n3202 , _u10_u8_n3201 , _u10_u8_n3200 , _u10_u8_n3199 ,_u10_u8_n3198 , _u10_u8_n3197 , _u10_u8_n3196 , _u10_u8_n3195 ,_u10_u8_n3194 , _u10_u8_n3193 , _u10_u8_n3192 , _u10_u8_n3191 ,_u10_u8_n3190 , _u10_u8_n3189 , _u10_u8_n3188 , _u10_u8_n3187 ,_u10_u8_n3186 , _u10_u8_n3185 , _u10_u8_n3184 , _u10_u8_n3183 ,_u10_u8_n3182 , _u10_u8_n3181 , _u10_u8_n3180 , _u10_u8_n3179 ,_u10_u8_n3178 , _u10_u8_n3177 , _u10_u8_n3176 , _u10_u8_n3175 ,_u10_u8_n3174 , _u10_u8_n3173 , _u10_u8_n3172 , _u10_u8_n3171 ,_u10_u8_n3170 , _u10_u8_n3169 , _u10_u8_n3168 , _u10_u8_n3167 ,_u10_u8_n3166 , _u10_u8_n3165 , _u10_u8_n3164 , _u10_u8_n3163 ,_u10_u8_n3162 , _u10_u8_n3161 , _u10_u8_n3160 , _u10_u8_n3159 ,_u10_u8_n3158 , _u10_u8_n3157 , _u10_u8_n3156 , _u10_u8_n3155 ,_u10_u8_n3154 , _u10_u8_n3153 , _u10_u8_n3152 , _u10_u8_n3151 ,_u10_u8_n3150 , _u10_u8_n3149 , _u10_u8_n3148 , _u10_u8_n3147 ,_u10_u8_n3146 , _u10_u8_n3145 , _u10_u8_n3144 , _u10_u8_n3143 ,_u10_u8_n3142 , _u10_u8_n3141 , _u10_u8_n3140 , _u10_u8_n3139 ,_u10_u8_n3138 , _u10_u8_n3137 , _u10_u8_n3136 , _u10_u8_n3135 ,_u10_u8_n3134 , _u10_u8_n3133 , _u10_u8_n3132 , _u10_u8_n3131 ,_u10_u8_n3130 , _u10_u8_n3129 , _u10_u8_n3128 , _u10_u8_n3127 ,_u10_u8_n3126 , _u10_u8_n3125 , _u10_u8_n3124 , _u10_u8_n3123 ,_u10_u8_n3122 , _u10_u8_n3121 , _u10_u8_n3120 , _u10_u8_n3119 ,_u10_u8_n3118 , _u10_u8_n3117 , _u10_u8_n3116 , _u10_u8_n3115 ,_u10_u8_n3114 , _u10_u8_n3113 , _u10_u8_n3112 , _u10_u8_n3111 ,_u10_u8_n3110 , _u10_u8_n3109 , _u10_u8_n3108 , _u10_u8_n3107 ,_u10_u8_n3106 , _u10_u8_n3105 , _u10_u8_n3104 , _u10_u8_n3103 ,_u10_u8_n3102 , _u10_u8_n3101 , _u10_u8_n3100 , _u10_u8_n3099 ,_u10_u8_n3098 , _u10_u8_n3097 , _u10_u8_n3096 , _u10_u8_n3095 ,_u10_u8_n3094 , _u10_u8_n3093 , _u10_u8_n3092 , _u10_u8_n3091 ,_u10_u8_n3090 , _u10_u8_n3089 , _u10_u8_n3088 , _u10_u8_n3087 ,_u10_u8_n3086 , _u10_u8_n3085 , _u10_u8_n3084 , _u10_u8_n3083 ,_u10_u8_n3082 , _u10_u8_n3081 , _u10_u8_n3080 , _u10_u8_n3079 ,_u10_u8_n3078 , _u10_u8_n3077 , _u10_u8_n3076 , _u10_u8_n3075 ,_u10_u8_n3074 , _u10_u8_n3073 , _u10_u8_n3072 , _u10_u8_n3071 ,_u10_u8_n3070 , _u10_u8_n3069 , _u10_u8_n3068 , _u10_u8_n3067 ,_u10_u8_n3066 , _u10_u8_n3065 , _u10_u8_n3064 , _u10_u8_n3063 ,_u10_u8_n3062 , _u10_u8_n3061 , _u10_u8_n3060 , _u10_u8_n3059 ,_u10_u8_n3058 , _u10_u8_n3057 , _u10_u8_n3056 , _u10_u8_n3055 ,_u10_u8_n3054 , _u10_u8_n3053 , _u10_u8_n3052 , _u10_u8_n3051 ,_u10_u8_n3050 , _u10_u8_n3049 , _u10_u8_n3048 , _u10_u8_n3047 ,_u10_u8_n3046 , _u10_u8_n3045 , _u10_u8_n3044 , _u10_u8_n3043 ,_u10_u8_n3042 , _u10_u8_n3041 , _u10_u8_n3040 , _u10_u8_n3039 ,_u10_u8_n3038 , _u10_u8_n3037 , _u10_u8_n3036 , _u10_u8_n3035 ,_u10_u8_n3034 , _u10_u8_n3033 , _u10_u8_n3032 , _u10_u8_n3031 ,_u10_u8_n3030 , _u10_u8_n3029 , _u10_u8_n3028 , _u10_u8_n3027 ,_u10_u8_n3026 , _u10_u8_n3025 , _u10_u8_n3024 , _u10_u8_n3023 ,_u10_u8_n3022 , _u10_u8_n3021 , _u10_u8_n3020 , _u10_u8_n3019 ,_u10_u8_n3018 , _u10_u8_n3017 , _u10_u8_n3016 , _u10_u8_n3015 ,_u10_u8_n3014 , _u10_u8_n3013 , _u10_u8_n3012 , _u10_u8_n3011 ,_u10_u8_n3010 , _u10_u8_n3009 , _u10_u8_n3008 , _u10_u8_n3007 ,_u10_u8_n3006 , _u10_u8_n3005 , _u10_u8_n3004 , _u10_u8_n3003 ,_u10_u8_n3002 , _u10_u8_n3001 , _u10_u8_n3000 , _u10_u8_n2999 ,_u10_u8_n2998 , _u10_u8_n2997 , _u10_u8_n2996 , _u10_u8_n2995 ,_u10_u8_n2994 , _u10_u8_n2993 , _u10_u8_n2992 , _u10_u8_n2991 ,_u10_u8_n2990 , _u10_u8_n2989 , _u10_u8_n2988 , _u10_u8_n2987 ,_u10_u8_n2986 , _u10_u8_n2985 , _u10_u8_n2984 , _u10_u8_n2983 ,_u10_u8_n2982 , _u10_u8_n2981 , _u10_u8_n2980 , _u10_u8_n2979 ,_u10_u8_n2978 , _u10_u8_n2977 , _u10_u8_n2976 , _u10_u8_n2975 ,_u10_u8_n2974 , _u10_u8_n2973 , _u10_u8_n2972 , _u10_u8_n2971 ,_u10_u8_n2970 , _u10_u8_n2969 , _u10_u8_n2968 , _u10_u8_n2967 ,_u10_u8_n2966 , _u10_u8_n2965 , _u10_u8_n2964 , _u10_u8_n2963 ,_u10_u8_n2962 , _u10_u8_n2961 , _u10_u8_n2960 , _u10_u8_n2959 ,_u10_u8_n2958 , _u10_u8_n2957 , _u10_u8_n2956 , _u10_u8_n2955 ,_u10_u8_n2954 , _u10_u8_n2953 , _u10_u8_n2952 , _u10_u8_n2951 ,_u10_u8_n2950 , _u10_u8_n2949 , _u10_u8_n2948 , _u10_u8_n2947 ,_u10_u8_n2946 , _u10_u8_n2945 , _u10_u8_n2944 , _u10_u8_n2943 ,_u10_u8_n2942 , _u10_u8_n2941 , _u10_u8_n2940 , _u10_u8_n2939 ,_u10_u8_n2938 , _u10_u8_n2937 , _u10_u8_n2936 , _u10_u8_n2935 ,_u10_u8_n2934 , _u10_u8_n2933 , _u10_u8_n2932 , _u10_u8_n2931 ,_u10_u8_n2930 , _u10_u8_n2929 , _u10_u8_n2928 , _u10_u8_n2927 ,_u10_u8_n2926 , _u10_u8_n2925 , _u10_u8_n2924 , _u10_u8_n2923 ,_u10_u8_n2922 , _u10_u8_n2921 , _u10_u8_n2920 , _u10_u8_n2919 ,_u10_u8_n2918 , _u10_u8_n2917 , _u10_u8_n2916 , _u10_u8_n2915 ,_u10_u8_n2914 , _u10_u8_n2913 , _u10_u8_n2912 , _u10_u8_n2911 ,_u10_u8_n2910 , _u10_u8_n2909 , _u10_u8_n2908 , _u10_u8_n2907 ,_u10_u8_n2906 , _u10_u8_n2905 , _u10_u8_n2904 , _u10_u8_n2903 ,_u10_u8_n2902 , _u10_u8_n2901 , _u10_u8_n2900 , _u10_u8_n2899 ,_u10_u8_n2898 , _u10_u8_n2897 , _u10_u8_n2896 , _u10_u8_n2895 ,_u10_u8_n2894 , _u10_u8_n2893 , _u10_u8_n2892 , _u10_u8_n2891 ,_u10_u8_n2890 , _u10_u8_n2889 , _u10_u8_n2888 , _u10_u8_n2887 ,_u10_u8_n2886 , _u10_u8_n2885 , _u10_u8_n2884 , _u10_u8_n2883 ,_u10_u8_n2882 , _u10_u8_n2881 , _u10_u8_n2880 , _u10_u8_n2879 ,_u10_u8_n2878 , _u10_u8_n2877 , _u10_u8_n2876 , _u10_u8_n2875 ,_u10_u8_n2874 , _u10_u8_n2873 , _u10_u8_n2872 , _u10_u8_n2871 ,_u10_u8_n2870 , _u10_u8_n2869 , _u10_u8_n2868 , _u10_u8_n2867 ,_u10_u8_n2866 , _u10_u8_n2865 , _u10_u8_n2864 , _u10_u8_n2863 ,_u10_u8_n2862 , _u10_u8_n2861 , _u10_u8_n2860 , _u10_u8_n2859 ,_u10_u8_n2858 , _u10_u8_n2857 , _u10_u8_n2856 , _u10_u8_n2855 ,_u10_u8_n2854 , _u10_u8_n2853 , _u10_u8_n2852 , _u10_u8_n2851 ,_u10_u8_n2850 , _u10_u8_n2849 , _u10_u8_n2848 , _u10_u8_n2847 ,_u10_u8_n2846 , _u10_u8_n2845 , _u10_u8_n2844 , _u10_u8_n2843 ,_u10_u8_n2842 , _u10_u8_n2841 , _u10_u8_n2840 , _u10_u8_n2839 ,_u10_u8_n2838 , _u10_u8_n2837 , _u10_u8_n2836 , _u10_u8_n2835 ,_u10_u8_n2834 , _u10_u8_n2833 , _u10_u8_n2832 , _u10_u8_n2831 ,_u10_u8_n2830 , _u10_u8_n2829 , _u10_u8_n2828 , _u10_u8_n2827 ,_u10_u8_n2826 , _u10_u8_n2825 , _u10_u8_n2824 , _u10_u8_n2823 ,_u10_u8_n2822 , _u10_u8_n2821 , _u10_u8_n2820 , _u10_u8_n2819 ,_u10_u8_n2818 , _u10_u8_n2817 , _u10_u8_n2816 , _u10_u8_n2815 ,_u10_u8_n2814 , _u10_u8_n2813 , _u10_u8_n2812 , _u10_u8_n2811 ,_u10_u8_n2810 , _u10_u8_n2809 , _u10_u8_n2808 , _u10_u8_n2807 ,_u10_u8_n2806 , _u10_u8_n2805 , _u10_u8_n2804 , _u10_u8_n2803 ,_u10_u8_n2802 , _u10_u8_n2801 , _u10_u8_n2800 , _u10_u8_n2799 ,_u10_u8_n2798 , _u10_u8_n2797 , _u10_u8_n2796 , _u10_u8_n2795 ,_u10_u8_n2794 , _u10_u8_n2793 , _u10_u8_n2792 , _u10_u8_n2791 ,_u10_u8_n2790 , _u10_u8_n2789 , _u10_u8_n2788 , _u10_u8_n2787 ,_u10_u8_n2786 , _u10_u8_n2785 , _u10_u8_n2784 , _u10_u8_n2783 ,_u10_u8_n2782 , _u10_u8_n2781 , _u10_u8_n2780 , _u10_u8_n2779 ,_u10_u8_n2778 , _u10_u8_n2777 , _u10_u8_n2776 , _u10_u8_n2775 ,_u10_u8_n2774 , _u10_u8_n2773 , _u10_u8_n2772 , _u10_u8_n2771 ,_u10_u8_n2770 , _u10_u8_n2769 , _u10_u8_n2768 , _u10_u8_n2767 ,_u10_u8_n2766 , _u10_u8_n2765 , _u10_u8_n2764 , _u10_u8_n2763 ,_u10_u8_n2762 , _u10_u8_n2761 , _u10_u8_n2760 , _u10_u8_n2759 ,_u10_u8_n2758 , _u10_u8_n2757 , _u10_u8_n2756 , _u10_u8_n2755 ,_u10_u8_n2754 , _u10_u8_n2753 , _u10_u8_n2752 , _u10_u8_n2751 ,_u10_u8_n2750 , _u10_u8_n2749 , _u10_u8_n2748 , _u10_u8_n2747 ,_u10_u8_n2746 , _u10_u8_n2745 , _u10_u8_n2744 , _u10_u8_n2743 ,_u10_u8_n2742 , _u10_u8_n2741 , _u10_u8_n2740 , _u10_u8_n2739 ,_u10_u8_n2738 , _u10_u8_n2737 , _u10_u8_n2736 , _u10_u8_n2735 ,_u10_u8_n2734 , _u10_u8_n2733 , _u10_u8_n2732 , _u10_u8_n2731 ,_u10_u8_n2730 , _u10_u8_n2729 , _u10_u8_n2728 , _u10_u8_n2727 ,_u10_u8_n2726 , _u10_u8_n2725 , _u10_u8_n2724 , _u10_u8_n2723 ,_u10_u8_n2722 , _u10_u8_n2721 , _u10_u8_n2720 , _u10_u8_n2719 ,_u10_u8_n2718 , _u10_u8_n2717 , _u10_u8_n2716 , _u10_u8_n2715 ,_u10_u8_n2714 , _u10_u8_n2713 , _u10_u8_n2712 , _u10_u8_n2711 ,_u10_u8_n2710 , _u10_u8_n2709 , _u10_u8_n2708 , _u10_u8_n2707 ,_u10_u8_n2706 , _u10_u8_n2705 , _u10_u8_n2704 , _u10_u8_n2703 ,_u10_u8_n2702 , _u10_u8_n2701 , _u10_u8_n2700 , _u10_u8_n2699 ,_u10_u8_n2698 , _u10_u8_n2697 , _u10_u8_n2696 , _u10_u8_n2695 ,_u10_u8_n2694 , _u10_u8_n2693 , _u10_u8_n2692 , _u10_u8_n2691 ,_u10_u8_n2690 , _u10_u8_n2689 , _u10_u8_n2688 , _u10_u8_n2687 ,_u10_u8_n2686 , _u10_u8_n2685 , _u10_u8_n2684 , _u10_u8_n2683 ,_u10_u8_n2682 , _u10_u8_n2681 , _u10_u8_n2680 , _u10_u8_n2679 ,_u10_u8_n2678 , _u10_u8_n2677 , _u10_u8_n2676 , _u10_u8_n2675 ,_u10_u8_n2674 , _u10_u8_n2673 , _u10_u8_n2672 , _u10_u8_n2671 ,_u10_u8_n2670 , _u10_u8_n2669 , _u10_u8_n2668 , _u10_u8_n2667 ,_u10_u8_n2666 , _u10_u8_n2665 , _u10_u8_n2664 , _u10_u8_n2663 ,_u10_u8_n2662 , _u10_u8_n2661 , _u10_u8_n2660 , _u10_u8_n2659 ,_u10_u8_n2658 , _u10_u8_n2657 , _u10_u8_n2656 , _u10_u8_n2655 ,_u10_u8_n2654 , _u10_u8_n2653 , _u10_u8_n2652 , _u10_u8_n2651 ,_u10_u8_n2650 , _u10_u8_n2649 , _u10_u8_n2648 , _u10_u8_n2647 ,_u10_u8_n2646 , _u10_u8_n2645 , _u10_u8_n2644 , _u10_u8_n2643 ,_u10_u8_n2642 , _u10_u8_n2641 , _u10_u8_n2640 , _u10_u8_n2639 ,_u10_u8_n2638 , _u10_u8_n2637 , _u10_u8_n2636 , _u10_u8_n2635 ,_u10_u8_n2634 , _u10_u8_n2633 , _u10_u8_n2632 , _u10_u8_n2631 ,_u10_u8_n2630 , _u10_u8_n2629 , _u10_u8_n2628 , _u10_u8_n2627 ,_u10_u8_n2626 , _u10_u8_n2625 , _u10_u8_n2624 , _u10_u8_n2623 ,_u10_u8_n2622 , _u10_u8_n2621 , _u10_u8_n2620 , _u10_u8_n2619 ,_u10_u8_n2618 , _u10_u8_n2617 , _u10_u8_n2616 , _u10_u8_n2615 ,_u10_u8_n2614 , _u10_u8_n2613 , _u10_u8_n2612 , _u10_u8_n2611 ,_u10_u8_n2610 , _u10_u8_n2609 , _u10_u8_n2608 , _u10_u8_n2607 ,_u10_u8_n2606 , _u10_u8_n2605 , _u10_u8_n2604 , _u10_u8_n2603 ,_u10_u8_n2602 , _u10_u8_n2601 , _u10_u8_n2600 , _u10_u8_n2599 ,_u10_u8_n2598 , _u10_u8_n2597 , _u10_u8_n2596 , _u10_u8_n2595 ,_u10_u8_n2594 , _u10_u8_n2593 , _u10_u8_n2592 , _u10_u8_n2591 ,_u10_u8_n2590 , _u10_u8_n2589 , _u10_u8_n2588 , _u10_u8_n2587 ,_u10_u8_n2586 , _u10_u8_n2585 , _u10_u8_n2584 , _u10_u8_n2583 ,_u10_u8_n2582 , _u10_u8_n2581 , _u10_u8_n2580 , _u10_u8_n2579 ,_u10_u8_n2578 , _u10_u8_n2577 , _u10_u8_n2576 , _u10_u8_n2575 ,_u10_u8_n2574 , _u10_u8_n2573 , _u10_u8_n2572 , _u10_u8_n2571 ,_u10_u8_n2570 , _u10_u8_n2569 , _u10_u8_n2568 , _u10_u8_n2567 ,_u10_u8_n2566 , _u10_u8_n2565 , _u10_u8_n2564 , _u10_u8_n2563 ,_u10_u8_n2562 , _u10_u8_n2561 , _u10_u8_n2560 , _u10_u8_n2559 ,_u10_u8_n2558 , _u10_u8_n2557 , _u10_u8_n2556 , _u10_u8_n2555 ,_u10_u8_n2554 , _u10_u8_n2553 , _u10_u8_n2552 , _u10_u8_n2551 ,_u10_u8_n2550 , _u10_u8_n2549 , _u10_u8_n2548 , _u10_u8_n2547 ,_u10_u8_n2546 , _u10_u8_n2545 , _u10_u8_n2544 , _u10_u8_n2543 ,_u10_u8_n2542 , _u10_u8_n2541 , _u10_u8_n2540 , _u10_u8_n2539 ,_u10_u8_n2538 , _u10_u8_n2537 , _u10_u8_n2536 , _u10_u8_n2535 ,_u10_u8_n2534 , _u10_u8_n2533 , _u10_u8_n2532 , _u10_u8_n2531 ,_u10_u8_n2530 , _u10_u8_n2529 , _u10_u8_n2528 , _u10_u8_n2527 ,_u10_u8_n2526 , _u10_u8_n2525 , _u10_u8_n2524 , _u10_u8_n2523 ,_u10_u8_n2522 , _u10_u8_n2521 , _u10_u8_n2520 , _u10_u8_n2519 ,_u10_u8_n2518 , _u10_u8_n2517 , _u10_u8_n2516 , _u10_u8_n2515 ,_u10_u8_n2514 , _u10_u8_n2513 , _u10_u8_n2512 , _u10_u8_n2511 ,_u10_u8_n2510 , _u10_u8_n2509 , _u10_u8_n2508 , _u10_u8_n2507 ,_u10_u8_n2506 , _u10_u8_n2505 , _u10_u8_n2504 , _u10_u8_n2503 ,_u10_u8_n2502 , _u10_u8_n2501 , _u10_u8_n2500 , _u10_u8_n2499 ,_u10_u8_n2498 , _u10_u8_n2497 , _u10_u8_n2496 , _u10_u8_n2495 ,_u10_u8_n2494 , _u10_u8_n2493 , _u10_u8_n2492 , _u10_u8_n2491 ,_u10_u8_n2490 , _u10_u8_n2489 , _u10_u8_n2488 , _u10_u8_n2487 ,_u10_u8_n2486 , _u10_u8_n2485 , _u10_u8_n2484 , _u10_u8_n2483 ,_u10_u8_n2482 , _u10_u8_n2481 , _u10_u8_n2480 , _u10_u8_n2479 ,_u10_u8_n2478 , _u10_u8_n2477 , _u10_u8_n2476 , _u10_u8_n2475 ,_u10_u8_n2474 , _u10_u8_n2473 , _u10_u8_n2472 , _u10_u8_n2471 ,_u10_u8_n2470 , _u10_u8_n2469 , _u10_u8_n2468 , _u10_u8_n2467 ,_u10_u8_n2466 , _u10_u8_n2465 , _u10_u8_n2464 , _u10_u8_n2463 ,_u10_u8_n2462 , _u10_u8_n2461 , _u10_u8_n2460 , _u10_u8_n2459 ,_u10_u8_n2458 , _u10_u8_n2457 , _u10_u8_n2456 , _u10_u8_n2455 ,_u10_u8_n2454 , _u10_u8_n2453 , _u10_u8_n2452 , _u10_u8_n2451 ,_u10_u8_n2450 , _u10_u8_n2449 , _u10_u8_n2448 , _u10_u8_n2447 ,_u10_u8_n2446 , _u10_u8_n2445 , _u10_u8_n2444 , _u10_u8_n2443 ,_u10_u8_n2442 , _u10_u8_n2441 , _u10_u8_n2440 , _u10_u8_n2439 ,_u10_u8_n2438 , _u10_u8_n2437 , _u10_u8_n2436 , _u10_u8_n2435 ,_u10_u8_n2434 , _u10_u8_n2433 , _u10_u8_n2432 , _u10_u8_n2431 ,_u10_u8_n2430 , _u10_u8_n2429 , _u10_u8_n2428 , _u10_u8_n2427 ,_u10_u8_n2426 , _u10_u8_n2425 , _u10_u8_n2424 , _u10_u8_n2423 ,_u10_u8_n2422 , _u10_u8_n2421 , _u10_u8_n2420 , _u10_u8_n2419 ,_u10_u8_n2418 , _u10_u8_n2417 , _u10_u8_n2416 , _u10_u8_n2415 ,_u10_u8_n2414 , _u10_u8_n2413 , _u10_u8_n2412 , _u10_u8_n2411 ,_u10_u8_n2410 , _u10_u8_n2409 , _u10_u8_n2408 , _u10_u8_n2407 ,_u10_u8_n2406 , _u10_u8_n2405 , _u10_u8_n2404 , _u10_u8_n2403 ,_u10_u8_n2402 , _u10_u8_n2401 , _u10_u8_n2400 , _u10_u8_n2399 ,_u10_u8_n2398 , _u10_u8_n2397 , _u10_u8_n2396 , _u10_u8_n2395 ,_u10_u8_n2394 , _u10_u8_n2393 , _u10_u8_n2392 , _u10_u8_n2391 ,_u10_u8_n2390 , _u10_u8_n2389 , _u10_u8_n2388 , _u10_u8_n2387 ,_u10_u8_n2386 , _u10_u8_n2385 , _u10_u8_n2384 , _u10_u8_n2383 ,_u10_u8_n2382 , _u10_u8_n2381 , _u10_u8_n2380 , _u10_u8_n2379 ,_u10_u8_n2378 , _u10_u8_n2377 , _u10_u8_n2376 , _u10_u8_n2375 ,_u10_u8_n2374 , _u10_u8_n2373 , _u10_u8_n2372 , _u10_u8_n2371 ,_u10_u8_n2370 , _u10_u8_n2369 , _u10_u8_n2368 , _u10_u8_n2367 ,_u10_u8_n2366 , _u10_u8_n2365 , _u10_u8_n2364 , _u10_u8_n2363 ,_u10_u8_n2362 , _u10_u8_n2361 , _u10_u8_n2360 , _u10_u8_n2359 ,_u10_u8_n2358 , _u10_u8_n2357 , _u10_u8_n2356 , _u10_u8_n2355 ,_u10_u8_n2354 , _u10_u8_n2353 , _u10_u8_n2352 , _u10_u8_n2351 ,_u10_u8_n2350 , _u10_u8_n2349 , _u10_u8_n2348 , _u10_u8_n2347 ,_u10_u8_n2346 , _u10_u8_n2345 , _u10_u8_n2344 , _u10_u8_n2343 ,_u10_u8_n2342 , _u10_u8_n2341 , _u10_u8_n2340 , _u10_u8_n2339 ,_u10_u8_n2338 , _u10_u8_n2337 , _u10_u8_n2336 , _u10_u8_n2335 ,_u10_u8_n2334 , _u10_u8_n2333 , _u10_u8_n2332 , _u10_u8_n2331 ,_u10_u8_n2330 , _u10_u8_n2329 , _u10_u8_n2328 , _u10_u8_n2327 ,_u10_u8_n2326 , _u10_u8_n2325 , _u10_u8_n2324 , _u10_u8_n2323 ,_u10_u8_n2322 , _u10_u8_n2321 , _u10_u8_n2320 , _u10_u8_n2319 ,_u10_u8_n2318 , _u10_u8_n2317 , _u10_u8_n2316 , _u10_u8_n2315 ,_u10_u8_n2314 , _u10_u8_n2313 , _u10_u8_n2312 , _u10_u8_n2311 ,_u10_u8_n2310 , _u10_u8_n2309 , _u10_u8_n2308 , _u10_u8_n2307 ,_u10_u8_n2306 , _u10_u8_n2305 , _u10_u8_n2304 , _u10_u8_n2303 ,_u10_u8_n2302 , _u10_u8_n2301 , _u10_u8_n2300 , _u10_u8_n2299 ,_u10_u8_n2298 , _u10_u8_n2297 , _u10_u8_n2296 , _u10_u8_n2295 ,_u10_u8_n2294 , _u10_u8_n2293 , _u10_u8_n2292 , _u10_u8_n2291 ,_u10_u8_n2290 , _u10_u8_n2289 , _u10_u8_n2288 , _u10_u8_n2287 ,_u10_u8_n2286 , _u10_u8_n2285 , _u10_u8_n2284 , _u10_u8_n2283 ,_u10_u8_n2282 , _u10_u8_n2281 , _u10_u8_n2280 , _u10_u8_n2279 ,_u10_u8_n2278 , _u10_u8_n2277 , _u10_u8_n2276 , _u10_u8_n2275 ,_u10_u8_n2274 , _u10_u8_n2273 , _u10_u8_n2272 , _u10_u8_n2271 ,_u10_u8_n2270 , _u10_u8_n2269 , _u10_u8_n2268 , _u10_u8_n2267 ,_u10_u8_n2266 , _u10_u8_n2265 , _u10_u8_n2264 , _u10_u8_n2263 ,_u10_u8_n2262 , _u10_u8_n2261 , _u10_u8_n2260 , _u10_u8_n2259 ,_u10_u8_n2258 , _u10_u8_n2257 , _u10_u8_n2256 , _u10_u8_n2255 ,_u10_u8_n2254 , _u10_u8_n2253 , _u10_u8_n2252 , _u10_u8_n2251 ,_u10_u8_n2250 , _u10_u8_n2249 , _u10_u8_n2248 , _u10_u8_n2247 ,_u10_u8_n2246 , _u10_u8_n2245 , _u10_u8_n2244 , _u10_u8_n2243 ,_u10_u8_n2242 , _u10_u8_n2241 , _u10_u8_n2240 , _u10_u8_n2239 ,_u10_u8_n2238 , _u10_u8_n2237 , _u10_u8_n2236 , _u10_u8_n2235 ,_u10_u8_n2234 , _u10_u8_n2233 , _u10_u8_n2232 , _u10_u8_n2231 ,_u10_u8_n2230 , _u10_u8_n2229 , _u10_u8_n2228 , _u10_u8_n2227 ,_u10_u8_n2226 , _u10_u8_n2225 , _u10_u8_n2224 , _u10_u8_n2223 ,_u10_u8_n2222 , _u10_u8_n2221 , _u10_u8_n2220 , _u10_u8_n2219 ,_u10_u8_n2218 , _u10_u8_n2217 , _u10_u8_n2216 , _u10_u8_n2215 ,_u10_u8_n2214 , _u10_u8_n2213 , _u10_u8_n2212 , _u10_u8_n2211 ,_u10_u8_n2210 , _u10_u8_n2209 , _u10_u8_n2208 , _u10_u8_n2207 ,_u10_u8_n2206 , _u10_u8_n2205 , _u10_u8_n2204 , _u10_u8_n2203 ,_u10_u8_n2202 , _u10_u8_n2201 , _u10_u8_n2200 , _u10_u8_n2199 ,_u10_u8_n2198 , _u10_u8_n2197 , _u10_u8_n2196 , _u10_u8_n2195 ,_u10_u8_n2194 , _u10_u8_n2193 , _u10_u8_n2192 , _u10_u8_n2191 ,_u10_u8_n2190 , _u10_u8_n2189 , _u10_u8_n2188 , _u10_u8_n2187 ,_u10_u8_n2186 , _u10_u8_n2185 , _u10_u8_n2184 , _u10_u8_n2183 ,_u10_u8_n2182 , _u10_u8_n2181 , _u10_u8_n2180 , _u10_u8_n2179 ,_u10_u8_n2178 , _u10_u8_n2177 , _u10_u8_n2176 , _u10_u8_n2175 ,_u10_u8_n2174 , _u10_u8_n2173 , _u10_u8_n2172 , _u10_u8_n2171 ,_u10_u8_n2170 , _u10_u8_n2169 , _u10_u8_n2168 , _u10_u8_n2167 ,_u10_u8_n2166 , _u10_u8_n2165 , _u10_u8_n2164 , _u10_u8_n2163 ,_u10_u8_n2162 , _u10_u8_n2161 , _u10_u8_n2160 , _u10_u8_n2159 ,_u10_u8_n2158 , _u10_u8_n2157 , _u10_u8_n2156 , _u10_u8_n2155 ,_u10_u8_n2154 , _u10_u8_n2153 , _u10_u8_n2152 , _u10_u8_n2151 ,_u10_u8_n2150 , _u10_u8_n2149 , _u10_u8_n2148 , _u10_u8_n2147 ,_u10_u8_n2146 , _u10_u8_n2145 , _u10_u8_n2144 , _u10_u8_n2143 ,_u10_u8_n2142 , _u10_u8_n2141 , _u10_u8_n2140 , _u10_u8_n2139 ,_u10_u8_n2138 , _u10_u8_n2137 , _u10_u8_n2136 , _u10_u8_n2135 ,_u10_u8_n2134 , _u10_u8_n2133 , _u10_u8_n2132 , _u10_u8_n2131 ,_u10_u8_n2130 , _u10_u8_n2129 , _u10_u8_n2128 , _u10_u8_n2127 ,_u10_u8_n2126 , _u10_u8_n2125 , _u10_u8_n2124 , _u10_u8_n2123 ,_u10_u8_n2122 , _u10_u8_n2121 , _u10_u8_n2120 , _u10_u8_n2119 ,_u10_u8_n2118 , _u10_u8_n2117 , _u10_u8_n2116 , _u10_u8_n2115 ,_u10_u8_n2114 , _u10_u8_n2113 , _u10_u8_n2112 , _u10_u8_n2111 ,_u10_u8_n2110 , _u10_u8_n2109 , _u10_u8_n2108 , _u10_u8_n2107 ,_u10_u8_n2106 , _u10_u8_n2105 , _u10_u8_n2104 , _u10_u8_n2103 ,_u10_u8_n2102 , _u10_u8_n2101 , _u10_u8_n2100 , _u10_u8_n2099 ,_u10_u8_n2098 , _u10_u8_n2097 , _u10_u8_n2096 , _u10_u8_n2095 ,_u10_u8_n2094 , _u10_u8_n2093 , _u10_u8_n2092 , _u10_u8_n2091 ,_u10_u8_n2090 , _u10_u8_n2089 , _u10_u8_n2088 , _u10_u8_n2087 ,_u10_u8_n2086 , _u10_u8_n2085 , _u10_u8_n2084 , _u10_u8_n2083 ,_u10_u8_n2082 , _u10_u8_n2081 , _u10_u8_n2080 , _u10_u8_n2079 ,_u10_u8_n2078 , _u10_u8_n2077 , _u10_u8_n2076 , _u10_u8_n2075 ,_u10_u8_n2074 , _u10_u8_n2073 , _u10_u8_n2072 , _u10_u8_n2071 ,_u10_u8_n2070 , _u10_u8_n2069 , _u10_u8_n2068 , _u10_u8_n2067 ,_u10_u8_n2066 , _u10_u8_n2065 , _u10_u8_n2064 , _u10_u8_n2063 ,_u10_u8_n2062 , _u10_u8_n2061 , _u10_u8_n2060 , _u10_u8_n2059 ,_u10_u8_n2058 , _u10_u8_n2057 , _u10_u8_n2056 , _u10_u8_n2055 ,_u10_u8_n2054 , _u10_u8_n2053 , _u10_u8_n2052 , _u10_u8_n2051 ,_u10_u8_n2050 , _u10_u8_n2049 , _u10_u8_n2048 , _u10_u8_n2047 ,_u10_u8_n2046 , _u10_u8_n2045 , _u10_u8_n2044 , _u10_u8_n2043 ,_u10_u8_n2042 , _u10_u8_n2041 , _u10_u8_n2040 , _u10_u8_n2039 ,_u10_u8_n2038 , _u10_u8_n2037 , _u10_u8_n2036 , _u10_u8_n2035 ,_u10_u8_n2034 , _u10_u8_n2033 , _u10_u8_n2032 , _u10_u8_n2031 ,_u10_u8_n2030 , _u10_u8_n2029 , _u10_u8_n2028 , _u10_u8_n2027 ,_u10_u8_n2026 , _u10_u8_n2025 , _u10_u8_n2024 , _u10_u8_n2023 ,_u10_u8_n2022 , _u10_u8_n2021 , _u10_u8_n2020 , _u10_u8_n2019 ,_u10_u8_n2018 , _u10_u8_n2017 , _u10_u8_n2016 , _u10_u8_n2015 ,_u10_u8_n2014 , _u10_u8_n2013 , _u10_u8_n2012 , _u10_u8_n2011 ,_u10_u8_n2010 , _u10_u8_n2009 , _u10_u8_n2008 , _u10_u8_n2007 ,_u10_u8_n2006 , _u10_u8_n2005 , _u10_u8_n2004 , _u10_u8_n2003 ,_u10_u8_n2002 , _u10_u8_n2001 , _u10_u8_n2000 , _u10_u8_n1999 ,_u10_u8_n1998 , _u10_u8_n1997 , _u10_u8_n1996 , _u10_u8_n1995 ,_u10_u8_n1994 , _u10_u8_n1993 , _u10_u8_n1992 , _u10_u8_n1991 ,_u10_u8_n1990 , _u10_u8_n1989 , _u10_u8_n1988 , _u10_u8_n1987 ,_u10_u8_n1986 , _u10_u8_n1985 , _u10_u8_n1984 , _u10_u8_n1983 ,_u10_u8_n1982 , _u10_u8_n1981 , _u10_u8_n1980 , _u10_u8_n1979 ,_u10_u8_n1978 , _u10_u8_n1977 , _u10_u8_n1976 , _u10_u8_n1975 ,_u10_u8_n1974 , _u10_u8_n1973 , _u10_u8_n1972 , _u10_u8_n1971 ,_u10_u8_n1970 , _u10_u8_n1969 , _u10_u8_n1968 , _u10_u8_n1967 ,_u10_u8_n1966 , _u10_u8_n1965 , _u10_u8_n1964 , _u10_u8_n1963 ,_u10_u8_n1962 , _u10_u8_n1961 , _u10_u8_n1960 , _u10_u8_n1959 ,_u10_u8_n1958 , _u10_u8_n1957 , _u10_u8_n1956 , _u10_u8_n1955 ,_u10_u8_n1954 , _u10_u8_n1953 , _u10_u8_n1952 , _u10_u8_n1951 ,_u10_u8_n1950 , _u10_u8_n1949 , _u10_u8_n1948 , _u10_u8_n1947 ,_u10_u8_n1946 , _u10_u8_n1945 , _u10_u8_n1944 , _u10_u8_n1943 ,_u10_u8_n1942 , _u10_u8_n1941 , _u10_u8_n1940 , _u10_u8_n1939 ,_u10_u8_n1938 , _u10_u8_n1937 , _u10_u8_n1936 , _u10_u8_n1935 ,_u10_u8_n1934 , _u10_u8_n1933 , _u10_u8_n1932 , _u10_u8_n1931 ,_u10_u8_n1930 , _u10_u8_n1929 , _u10_u8_n1928 , _u10_u8_n1927 ,_u10_u8_n1926 , _u10_u8_n1925 , _u10_u8_n1924 , _u10_u8_n1923 ,_u10_u8_n1922 , _u10_u8_n1921 , _u10_u8_n1920 , _u10_u8_n1919 ,_u10_u8_n1918 , _u10_u8_n1917 , _u10_u8_n1916 , _u10_u8_n1915 ,_u10_u8_n1914 , _u10_u8_n1913 , _u10_u8_n1912 , _u10_u8_n1911 ,_u10_u8_n1910 , _u10_u8_n1909 , _u10_u8_n1908 , _u10_u8_n1907 ,_u10_u8_n1906 , _u10_u8_n1905 , _u10_u8_n1904 , _u10_u8_n1903 ,_u10_u8_n1902 , _u10_u8_n1901 , _u10_u8_n1900 , _u10_u8_n1899 ,_u10_u8_n1898 , _u10_u8_n1897 , _u10_u8_n1896 , _u10_u8_n1895 ,_u10_u8_n1894 , _u10_u8_n1893 , _u10_u8_n1892 , _u10_u8_n1891 ,_u10_u8_n1890 , _u10_u8_n1889 , _u10_u8_n1888 , _u10_u8_n1887 ,_u10_u8_n1886 , _u10_u8_n1885 , _u10_u8_n1884 , _u10_u8_n1883 ,_u10_u8_n1882 , _u10_u8_n1881 , _u10_u8_n1880 , _u10_u8_n1879 ,_u10_u8_n1878 , _u10_u8_n1877 , _u10_u8_n1876 , _u10_u8_n1875 ,_u10_u8_n1874 , _u10_u8_n1873 , _u10_u8_n1872 , _u10_u8_n1871 ,_u10_u8_n1870 , _u10_u8_n1869 , _u10_u8_n1868 , _u10_u8_n1867 ,_u10_u8_n1866 , _u10_u8_n1865 , _u10_u8_n1864 , _u10_u8_n1863 ,_u10_u8_n1862 , _u10_u8_n1861 , _u10_u8_n1860 , _u10_u8_n1859 ,_u10_u8_n1858 , _u10_u8_n1857 , _u10_u8_n1856 , _u10_u8_n1855 ,_u10_u8_n1854 , _u10_u8_n1853 , _u10_u8_n1852 , _u10_u8_n1851 ,_u10_u8_n1850 , _u10_u8_n1849 , _u10_u8_n1848 , _u10_u8_n1847 ,_u10_u8_n1846 , _u10_u8_n1845 , _u10_u8_n1844 , _u10_u8_n1843 ,_u10_u8_n1842 , _u10_u8_n1841 , _u10_u8_n1840 , _u10_u8_n1839 ,_u10_u8_n1838 , _u10_u8_n1837 , _u10_u8_n1836 , _u10_u8_n1835 ,_u10_u8_n1834 , _u10_u8_n1833 , _u10_u8_n1832 , _u10_u8_n1831 ,_u10_u8_n1830 , _u10_u8_n1829 , _u10_u8_n1828 , _u10_u8_n1827 ,_u10_u8_n1826 , _u10_u8_n1825 , _u10_u8_n1824 , _u10_u8_n1823 ,_u10_u8_n1822 , _u10_u8_n1821 , _u10_u8_n1820 , _u10_u8_n1819 ,_u10_u8_n1818 , _u10_u8_n1817 , _u10_u8_n1816 , _u10_u8_n1815 ,_u10_u8_n1814 , _u10_u8_n1813 , _u10_u8_n1812 , _u10_u8_n1811 ,_u10_u8_n1810 , _u10_u8_n1809 , _u10_u8_n1808 , _u2_n1566 ,_u2_n1565 , _u2_n1564 , _u2_n1563 , _u2_n1562 , _u2_n1561 ,_u2_n1560 , _u2_n1559 , _u2_n1558 , _u2_n1557 , _u2_n1556 ,_u2_n1555 , _u2_n1554 , _u2_n1553 , _u2_n1552 , _u2_n1551 ,_u2_n1550 , _u2_n1549 , _u2_n1548 , _u2_n1547 , _u2_n1546 ,_u2_n1545 , _u2_n1544 , _u2_n1543 , _u2_n1542 , _u2_n1541 ,_u2_n1540 , _u2_n1539 , _u2_n1538 , _u2_n1537 , _u2_n1536 ,_u2_n1535 , _u2_n1534 , _u2_n1533 , _u2_n1532 , _u2_n1531 ,_u2_n1530 , _u2_n1529 , _u2_n1528 , _u2_n1527 , _u2_n1526 ,_u2_n1525 , _u2_n1524 , _u2_n1523 , _u2_n1522 , _u2_n1521 ,_u2_n1520 , _u2_n1519 , _u2_n1518 , _u2_n1517 , _u2_n1516 ,_u2_n1515 , _u2_n1514 , _u2_n1513 , _u2_n1512 , _u2_n1511 ,_u2_n1510 , _u2_n1509 , _u2_n1508 , _u2_n1507 , _u2_n1506 ,_u2_n1505 , _u2_n1504 , _u2_n1503 , _u2_n1502 , _u2_n1501 ,_u2_n1500 , _u2_n1499 , _u2_n1498 , _u2_n1497 , _u2_n1496 ,_u2_n1495 , _u2_n1494 , _u2_n1493 , _u2_n1492 , _u2_n1491 ,_u2_n1490 , _u2_n1489 , _u2_n1488 , _u2_n1487 , _u2_n1486 ,_u2_n1485 , _u2_n1484 , _u2_n1483 , _u2_n1482 , _u2_n1481 ,_u2_n1480 , _u2_n1479 , _u2_n1478 , _u2_n1477 , _u2_n1476 ,_u2_n1475 , _u2_n1474 , _u2_n1473 , _u2_n1472 , _u2_n1471 ,_u2_n1470 , _u2_n1469 , _u2_n1468 , _u2_n1467 , _u2_n1466 ,_u2_n1465 , _u2_n1464 , _u2_n1463 , _u2_n1462 , _u2_n1461 ,_u2_n1460 , _u2_n1459 , _u2_n1458 , _u2_n1457 , _u2_n1456 ,_u2_n1455 , _u2_n1454 , _u2_n1453 , _u2_n1452 , _u2_n1451 ,_u2_n1450 , _u2_n1449 , _u2_n1448 , _u2_n1447 , _u2_n1446 ,_u2_n1445 , _u2_n1444 , _u2_n1443 , _u2_n1442 , _u2_n1441 ,_u2_n1440 , _u2_n1439 , _u2_n1438 , _u2_n1437 , _u2_n1436 ,_u2_n1435 , _u2_n1434 , _u2_n1433 , _u2_n1432 , _u2_n1431 ,_u2_n1430 , _u2_n1429 , _u2_n1428 , _u2_n1427 , _u2_n1426 ,_u2_n1425 , _u2_n1424 , _u2_n1423 , _u2_n1422 , _u2_n1421 ,_u2_n1420 , _u2_n1419 , _u2_n1418 , _u2_n1417 , _u2_n1416 ,_u2_n1415 , _u2_n1414 , _u2_n1413 , _u2_n1412 , _u2_n1411 ,_u2_n1410 , _u2_n1409 , _u2_n1408 , _u2_n1407 , _u2_n1406 ,_u2_n1405 , _u2_n1404 , _u2_n1403 , _u2_n1402 , _u2_n1401 ,_u2_n1400 , _u2_n1399 , _u2_n1398 , _u2_n1397 , _u2_n1396 ,_u2_n1395 , _u2_n1394 , _u2_n1393 , _u2_n1392 , _u2_n1391 ,_u2_n1390 , _u2_n1389 , _u2_n1388 , _u2_n1387 , _u2_n1386 ,_u2_n1385 , _u2_n1384 , _u2_n1383 , _u2_n1382 , _u2_n1381 ,_u2_n1380 , _u2_n1379 , _u2_n1378 , _u2_n1377 , _u2_n1376 ,_u2_n1375 , _u2_n1374 , _u2_n1373 , _u2_n1372 , _u2_n1371 ,_u2_n1370 , _u2_n1369 , _u2_n1368 , _u2_n1367 , _u2_n1366 ,_u2_n1365 , _u2_n1364 , _u2_n1363 , _u2_n1362 , _u2_n1361 ,_u2_n1360 , _u2_n1359 , _u2_n1358 , _u2_n1357 , _u2_n1356 ,_u2_n1355 , _u2_n1354 , _u2_n1353 , _u2_n1352 , _u2_n1351 ,_u2_n1350 , _u2_n1349 , _u2_n1348 , _u2_n1347 , _u2_n1346 ,_u2_n1345 , _u2_n1344 , _u2_n1343 , _u2_n1342 , _u2_n1341 ,_u2_n1340 , _u2_n1339 , _u2_n1338 , _u2_n1337 , _u2_n1336 ,_u2_n1335 , _u2_n1334 , _u2_n1333 , _u2_n1332 , _u2_n1331 ,_u2_n1330 , _u2_n1329 , _u2_n1328 , _u2_n1327 , _u2_n1326 ,_u2_n1325 , _u2_n1324 , _u2_n1323 , _u2_n1322 , _u2_n1321 ,_u2_n1320 , _u2_n1319 , _u2_n1318 , _u2_n1317 , _u2_n1316 ,_u2_n1315 , _u2_n1314 , _u2_n1313 , _u2_n1312 , _u2_n1311 ,_u2_n1310 , _u2_n1309 , _u2_n1308 , _u2_n1307 , _u2_n1306 ,_u2_n1305 , _u2_n1304 , _u2_n1303 , _u2_n1302 , _u2_n1301 ,_u2_n1300 , _u2_n1299 , _u2_n1298 , _u2_n1297 , _u2_n1296 ,_u2_n1295 , _u2_n1294 , _u2_n1293 , _u2_n1292 , _u2_n1291 ,_u2_n1290 , _u2_n1289 , _u2_n1288 , _u2_n1287 , _u2_n1286 ,_u2_n1285 , _u2_n1284 , _u2_n1283 , _u2_n1282 , _u2_n1281 ,_u2_n1280 , _u2_n1279 , _u2_n1278 , _u2_n1277 , _u2_n1276 ,_u2_n1275 , _u2_n1274 , _u2_n1273 , _u2_n1272 , _u2_n1271 ,_u2_n1270 , _u2_n1269 , _u2_n1268 , _u2_n1267 , _u2_n1266 ,_u2_n1265 , _u2_n1264 , _u2_n1263 , _u2_n1262 , _u2_n1261 ,_u2_n1260 , _u2_n1259 , _u2_n1258 , _u2_n1257 , _u2_n1256 ,_u2_n1255 , _u2_n1254 , _u2_n1253 , _u2_n1252 , _u2_n1251 ,_u2_n1250 , _u2_n1249 , _u2_n1248 , _u2_n1247 , _u2_n1246 ,_u2_n1245 , _u2_n1244 , _u2_n1243 , _u2_n1242 , _u2_n1241 ,_u2_n1240 , _u2_n1239 , _u2_n1238 , _u2_n1237 , _u2_n1236 ,_u2_n1235 , _u2_n1234 , _u2_n1233 , _u2_n1232 , _u2_n1231 ,_u2_n1230 , _u2_n1229 , _u2_n1228 , _u2_n1227 , _u2_n1226 ,_u2_n1225 , _u2_n1224 , _u2_n1223 , _u2_n1222 , _u2_n1221 ,_u2_n1220 , _u2_n1219 , _u2_n1218 , _u2_n1217 , _u2_n1216 ,_u2_n1215 , _u2_n1214 , _u2_n1213 , _u2_n1212 , _u2_n1211 ,_u2_n1210 , _u2_n1209 , _u2_n1208 , _u2_n1207 , _u2_n1206 ,_u2_n1205 , _u2_n1204 , _u2_n1203 , _u2_n1202 , _u2_n1201 ,_u2_n1200 , _u2_n1199 , _u2_n1198 , _u2_n1197 , _u2_n1196 ,_u2_n1195 , _u2_n1194 , _u2_n1193 , _u2_n1192 , _u2_n1191 ,_u2_n1190 , _u2_n1189 , _u2_n1188 , _u2_n1187 , _u2_n1186 ,_u2_n1185 , _u2_n1184 , _u2_n1183 , _u2_n1182 , _u2_n1181 ,_u2_n1180 , _u2_n1179 , _u2_n1178 , _u2_n1177 , _u2_n1176 ,_u2_n1175 , _u2_n1174 , _u2_n1173 , _u2_n1172 , _u2_n1171 ,_u2_n1170 , _u2_n1169 , _u2_n1168 , _u2_n1167 , _u2_n1166 ,_u2_n1165 , _u2_n1164 , _u2_n1163 , _u2_n1162 , _u2_n1161 ,_u2_n1160 , _u2_n1159 , _u2_n1158 , _u2_n1157 , _u2_n1156 ,_u2_n1155 , _u2_n1154 , _u2_n1153 , _u2_n1152 , _u2_n1151 ,_u2_n1150 , _u2_n1149 , _u2_n1148 , _u2_n1147 , _u2_n1146 ,_u2_n1145 , _u2_n1144 , _u2_n1143 , _u2_n1142 , _u2_n1141 ,_u2_n1140 , _u2_n1139 , _u2_n1138 , _u2_n1137 , _u2_n1136 ,_u2_n1135 , _u2_n1134 , _u2_n1133 , _u2_n1132 , _u2_n1131 ,_u2_n1130 , _u2_n1129 , _u2_n1128 , _u2_n1127 , _u2_n1126 ,_u2_n1125 , _u2_n1124 , _u2_n1123 , _u2_n1122 , _u2_n1121 ,_u2_n1120 , _u2_n1119 , _u2_n1118 , _u2_n1117 , _u2_n1116 ,_u2_n1115 , _u2_n1114 , _u2_n1113 , _u2_n1112 , _u2_n1111 ,_u2_n1110 , _u2_n1109 , _u2_n1108 , _u2_n1107 , _u2_n1106 ,_u2_n1105 , _u2_n1104 , _u2_n1103 , _u2_n1102 , _u2_n1101 ,_u2_n1100 , _u2_n1099 , _u2_n1098 , _u2_n1097 , _u2_n1096 ,_u2_n1095 , _u2_n1094 , _u2_n1093 , _u2_n1092 , _u2_n1091 ,_u2_n1090 , _u2_n1089 , _u2_n1088 , _u2_n1087 , _u2_n1086 ,_u2_n1085 , _u2_n1084 , _u2_n1083 , _u2_n1082 , _u2_n1081 ,_u2_n1080 , _u2_n1079 , _u2_n1078 , _u2_n1077 , _u2_n1076 ,_u2_n1075 , _u2_n1074 , _u2_n1073 , _u2_n1072 , _u2_n1071 ,_u2_n1070 , _u2_n1069 , _u2_n1068 , _u2_n1067 , _u2_n1066 ,_u2_n1065 , _u2_n1064 , _u2_n1063 , _u2_n1062 , _u2_n1061 ,_u2_n1060 , _u2_n1059 , _u2_n1058 , _u2_n1057 , _u2_n1056 ,_u2_n1055 , _u2_n1054 , _u2_n1051 , _u2_n1050 , _u2_n1049 ,_u2_n1048 , _u2_n1047 , _u2_n1046 , _u2_n1043 , _u2_n1010 ,_u2_n1009 , _u2_n1008 , _u2_n1007 , _u2_n1005 , _u2_n943 , _u2_n942 ,_u2_n941 , _u2_n940 , _u2_n939 , _u2_n938 , _u2_n937 , _u2_n936 ,_u2_n935 , _u2_n933 , _u2_n932 , _u2_n930 , _u2_n929 , _u2_n928 ,_u2_n927 , _u2_n926 , _u2_n925 , _u2_n924 , _u2_n923 , _u2_n922 ,_u2_n921 , _u2_n920 , _u2_n919 , _u2_n918 , _u2_n917 , _u2_n916 ,_u2_n915 , _u2_n914 , _u2_n913 , _u2_n912 , _u2_n911 , _u2_n910 ,_u2_n909 , _u2_n908 , _u2_n907 , _u2_n906 , _u2_n905 , _u2_n904 ,_u2_n903 , _u2_n902 , _u2_n901 , _u2_n900 , _u2_n899 , _u2_n898 ,_u2_n897 , _u2_n896 , _u2_n895 , _u2_n894 , _u2_n893 , _u2_n892 ,_u2_n891 , _u2_n890 , _u2_n889 , _u2_n888 , _u2_n887 , _u2_n886 ,_u2_n885 , _u2_n884 , _u2_n883 , _u2_n882 , _u2_n881 , _u2_n880 ,_u2_n879 , _u2_n878 , _u2_n877 , _u2_n876 , _u2_n875 , _u2_n874 ,_u2_n873 , _u2_n872 , _u2_n871 , _u2_n870 , _u2_n869 , _u2_n868 ,_u2_n867 , _u2_n866 , _u2_n865 , _u2_n864 , _u2_n863 , _u2_n862 ,_u2_n861 , _u2_n860 , _u2_n859 , _u2_n858 , _u2_n857 , _u2_n856 ,_u2_n855 , _u2_n854 , _u2_n853 , _u2_n852 , _u2_n851 , _u2_n850 ,_u2_n849 , _u2_n848 , _u2_n847 , _u2_n846 , _u2_n845 , _u2_n844 ,_u2_n843 , _u2_n842 , _u2_n841 , _u2_n840 , _u2_n839 , _u2_n838 ,_u2_n837 , _u2_n836 , _u2_n835 , _u2_n834 , _u2_n833 , _u2_n832 ,_u2_n831 , _u2_n830 , _u2_n829 , _u2_n828 , _u2_n827 , _u2_n826 ,_u2_n825 , _u2_n824 , _u2_n823 , _u2_n822 , _u2_n821 , _u2_n820 ,_u2_n819 , _u2_n818 , _u2_n817 , _u2_n816 , _u2_n815 , _u2_n814 ,_u2_n813 , _u2_n812 , _u2_n811 , _u2_n810 , _u2_n809 , _u2_n808 ,_u2_n807 , _u2_n806 , _u2_n805 , _u2_n804 , _u2_n803 , _u2_n802 ,_u2_n801 , _u2_n800 , _u2_n799 , _u2_n798 , _u2_n797 , _u2_n796 ,_u2_n795 , _u2_n794 , _u2_n793 , _u2_n792 , _u2_n791 , _u2_n790 ,_u2_n789 , _u2_n788 , _u2_n787 , _u2_n786 , _u2_n785 , _u2_n784 ,_u2_n783 , _u2_n782 , _u2_n781 , _u2_n780 , _u2_n779 , _u2_n778 ,_u2_n777 , _u2_n776 , _u2_n775 , _u2_n774 , _u2_n773 , _u2_n772 ,_u2_n771 , _u2_n770 , _u2_n769 , _u2_n768 , _u2_n767 , _u2_n766 ,_u2_n765 , _u2_n729 , _u2_n728 , _u2_n727 , _u2_n726 , _u2_n725 ,_u2_n724 , _u2_n723 , _u2_n722 , _u2_n721 , _u2_n720 , _u2_n719 ,_u2_n718 , _u2_mast1_adr[1] , _u2_mast1_adr[0] , _u2_n1053 ,_u2_n1052 , _u2_n1045 , _u2_n1044 , _u2_n1042 , _u2_n1041 ,_u2_n1040 , _u2_n1039 , _u2_n1038 , _u2_n1037 , _u2_n1036 ,_u2_n1035 , _u2_n1034 , _u2_n1033 , _u2_n1032 , _u2_n1031 ,_u2_n1030 , _u2_n1029 , _u2_n1028 , _u2_n1027 , _u2_n1026 ,_u2_n1025 , _u2_n1024 , _u2_n1023 , _u2_n1022 , _u2_n1021 ,_u2_n1020 , _u2_n1019 , _u2_n1018 , _u2_n1017 , _u2_n1016 ,_u2_n1015 , _u2_n1014 , _u2_n1013 , _u2_n1012 , _u2_n1011 ,_u2_n1006 , _u2_n1004 , _u2_n1003 , _u2_n1002 , _u2_n1001 ,_u2_n1000 , _u2_n999 , _u2_n998 , _u2_n997 , _u2_n996 , _u2_n995 ,_u2_n994 , _u2_n993 , _u2_n992 , _u2_n991 , _u2_n990 , _u2_n989 ,_u2_n988 , _u2_n987 , _u2_n986 , _u2_n985 , _u2_n984 , _u2_n983 ,_u2_n982 , _u2_n981 , _u2_n980 , _u2_n979 , _u2_n978 , _u2_n977 ,_u2_n976 , _u2_n975 , _u2_n974 , _u2_n973 , _u2_n972 , _u2_n971 ,_u2_n970 , _u2_n969 , _u2_n968 , _u2_n967 , _u2_n966 , _u2_n965 ,_u2_n964 , _u2_n963 , _u2_n962 , _u2_n961 , _u2_n960 , _u2_n959 ,_u2_n958 , _u2_n957 , _u2_n956 , _u2_n955 , _u2_n954 , _u2_n953 ,_u2_n952 , _u2_n951 , _u2_n950 , _u2_n949 , _u2_n948 , _u2_n947 ,_u2_n946 , _u2_n945 , _u2_n944 , _u2_n934 , _u2_n931 , _u2_N342 ,_u2_write_hold_r , _u2_N341 , _u2_N340 , _u2_N339 , _u2_N338 ,_u2_N337 , _u2_N336 , _u2_N335 , _u2_N334 , _u2_N333 , _u2_N332 ,_u2_N331 , _u2_N330 , _u2_N329 , _u2_N328 , _u2_N327 , _u2_N326 ,_u2_N325 , _u2_N324 , _u2_N323 , _u2_N322 , _u2_N321 , _u2_N320 ,_u2_N319 , _u2_N318 , _u2_N317 , _u2_N316 , _u2_N315 , _u2_N314 ,_u2_N313 , _u2_N312 , _u2_N308 , _u2_N307 , _u2_N306 , _u2_N305 ,_u2_N304 , _u2_N303 , _u2_N302 , _u2_N301 , _u2_N300 , _u2_N299 ,_u2_N298 , _u2_N297 , _u2_N296 , _u2_N295 , _u2_N294 , _u2_N293 ,_u2_N292 , _u2_N291 , _u2_N290 , _u2_N289 , _u2_N288 , _u2_N287 ,_u2_N286 , _u2_N285 , _u2_N284 , _u2_N283 , _u2_N282 , _u2_N281 ,_u2_N280 , _u2_N279 , _u2_N278 , _u2_N277 , _u2_state_0_ ,_u2_state_1_ , _u2_state_2_ , _u2_state_3_ , _u2_state_4_ ,_u2_state_5_ , _u2_state_6_ , _u2_state_7_ , _u2_state_9_ , _u2_N236 ,_u2_N232 , _u2_read_r , _u2_read , _u2_N215 , _u2_N214 , _u2_N213 ,_u2_N212 , _u2_N211 , _u2_N210 , _u2_N209 , _u2_N208 , _u2_N207 ,_u2_N206 , _u2_N205 , _u2_N204 , _u2_tsz_cnt[0] , _u2_tsz_cnt[1] ,_u2_tsz_cnt[2] , _u2_tsz_cnt[3] , _u2_tsz_cnt[4] , _u2_tsz_cnt[5] ,_u2_tsz_cnt[6] , _u2_tsz_cnt[7] , _u2_tsz_cnt[8] , _u2_tsz_cnt[9] ,_u2_tsz_cnt[10] , _u2_tsz_cnt[11] , _u2_tsz_cnt_is_0_r , _u2_N188 ,_u2_N187 , _u2_N186 , _u2_N185 , _u2_N184 , _u2_N183 , _u2_N182 ,_u2_N181 , _u2_N180 , _u2_chunk_cnt[0] , _u2_chunk_cnt[1] ,_u2_chunk_cnt[2] , _u2_chunk_cnt[3] , _u2_chunk_cnt[4] ,_u2_chunk_cnt[5] , _u2_chunk_cnt[6] , _u2_chunk_cnt[7] ,_u2_chunk_cnt[8] , _u2_chunk_dec , _u2_adr1_cnt[0] , _u2_adr1_cnt[1] ,_u2_adr1_cnt[2] , _u2_adr1_cnt[3] , _u2_adr1_cnt[4] ,_u2_adr1_cnt[5] , _u2_adr1_cnt[6] , _u2_adr1_cnt[7] ,_u2_adr1_cnt[8] , _u2_adr1_cnt[9] , _u2_adr1_cnt[10] ,_u2_adr1_cnt[11] , _u2_adr1_cnt[12] , _u2_adr1_cnt[13] ,_u2_adr1_cnt[14] , _u2_adr1_cnt[15] , _u2_adr1_cnt[16] ,_u2_adr1_cnt[17] , _u2_adr1_cnt[18] , _u2_adr1_cnt[19] ,_u2_adr1_cnt[20] , _u2_adr1_cnt[21] , _u2_adr1_cnt[22] ,_u2_adr1_cnt[23] , _u2_adr1_cnt[24] , _u2_adr1_cnt[25] ,_u2_adr1_cnt[26] , _u2_adr1_cnt[27] , _u2_adr1_cnt[28] ,_u2_adr1_cnt[29] , _u2_adr0_cnt[0] , _u2_adr0_cnt[1] ,_u2_adr0_cnt[2] , _u2_adr0_cnt[3] , _u2_adr0_cnt[4] ,_u2_adr0_cnt[5] , _u2_adr0_cnt[6] , _u2_adr0_cnt[7] ,_u2_adr0_cnt[8] , _u2_adr0_cnt[9] , _u2_adr0_cnt[10] ,_u2_adr0_cnt[11] , _u2_adr0_cnt[12] , _u2_adr0_cnt[13] ,_u2_adr0_cnt[14] , _u2_adr0_cnt[15] , _u2_adr0_cnt[16] ,_u2_adr0_cnt[17] , _u2_adr0_cnt[18] , _u2_adr0_cnt[19] ,_u2_adr0_cnt[20] , _u2_adr0_cnt[21] , _u2_adr0_cnt[22] ,_u2_adr0_cnt[23] , _u2_adr0_cnt[24] , _u2_adr0_cnt[25] ,_u2_adr0_cnt[26] , _u2_adr0_cnt[27] , _u2_adr0_cnt[28] ,_u2_adr0_cnt[29] , _u2_sub_360_S2_n39 , _u2_sub_360_S2_n38 ,_u2_sub_360_S2_n37 , _u2_sub_360_S2_n36 , _u2_sub_360_S2_n35 ,_u2_sub_360_S2_n34 , _u2_sub_360_S2_n33 , _u2_sub_360_S2_n32 ,_u2_sub_360_S2_n31 , _u2_sub_360_S2_n30 , _u2_sub_360_S2_n29 ,_u2_sub_360_S2_n28 , _u2_sub_360_S2_n27 , _u2_sub_360_S2_n26 ,_u2_sub_360_S2_n25 , _u2_sub_360_S2_n24 , _u2_sub_360_S2_n23 ,_u2_sub_360_S2_n22 , _u2_sub_360_S2_n21 , _u2_sub_349_S2_n27 ,_u2_sub_349_S2_n26 , _u2_sub_349_S2_n25 , _u2_sub_349_S2_n24 ,_u2_sub_349_S2_n23 , _u2_sub_349_S2_n22 , _u2_sub_349_S2_n21 ,_u2_sub_349_S2_n20 , _u2_sub_349_S2_n19 , _u2_sub_349_S2_n18 ,_u2_sub_349_S2_n17 , _u2_sub_349_S2_n16 , _u2_sub_349_S2_n15 ,_u3_u0_n42 , _u3_u0_n41 , _u3_u0_n6 , _u3_u0_n233 , _u3_u0_n232 ,_u3_u0_n231 , _u3_u0_n230 , _u3_u0_n229 , _u3_u0_n228 , _u3_u0_n227 ,_u3_u0_n226 , _u3_u0_n225 , _u3_u0_n224 , _u3_u0_n223 , _u3_u0_n222 ,_u3_u0_n221 , _u3_u0_n220 , _u3_u0_n219 , _u3_u0_n218 , _u3_u0_n217 ,_u3_u0_n216 , _u3_u0_n215 , _u3_u0_n214 , _u3_u0_n213 , _u3_u0_n212 ,_u3_u0_n211 , _u3_u0_n210 , _u3_u0_n209 , _u3_u0_n208 , _u3_u0_n207 ,_u3_u0_n206 , _u3_u0_n205 , _u3_u0_n204 , _u3_u0_n203 , _u3_u0_n202 ,_u3_u0_N3 , _u3_u0_mast_stb , _u3_u0_mast_cyc , _u3_u0_mast_we_r ,_u3_u1_n91 , _u3_u1_n90 , _u3_u1_n89 , _u3_u1_n88 , _u3_u1_n16 ,_u3_u1_n15 , _u3_u1_n14 , _u3_u1_n12 , _u3_u1_n11 , _u3_u1_N5 ,_u3_u1_N4 , _u3_u1_N3 , _u3_u1_rf_ack , _u40_slv_we , _u40_slv_re ,_u40_u0_n74 , _u40_u0_n73 , _u40_u0_n38 , _u40_u0_n34 , _u40_u0_n33 ,_u40_u0_n32 , _u40_u0_n31 , _u40_u0_n301 , _u40_u0_n29 , _u40_u0_n28 ,_u40_u0_n27 , _u40_u0_n26 , _u40_u0_n25 , _u40_u0_n24 , _u40_u0_n23 ,_u40_u0_n22 , _u40_u0_n21 , _u40_u0_n20 , _u40_u0_n19 , _u40_u0_n18 ,_u40_u0_n17 , _u40_u0_n16 , _u40_u0_n15 , _u40_u0_n14 , _u40_u0_n13 ,_u40_u0_n12 , _u40_u0_n11 , _u40_u0_n10 , _u40_u0_n9 , _u40_u0_n8 ,_u40_u0_n7 , _u40_u0_n6 , _u40_u0_n5 , _u40_u0_n4 , _u40_u0_n300 ,_u40_u0_N3 , _u40_u0_mast_stb , _u40_u0_mast_cyc , _u40_u0_mast_we_r ,_u40_u1_n91 , _u40_u1_n90 , _u40_u1_n89 , _u40_u1_n88 , _u40_u1_n16 ,_u40_u1_n15 , _u40_u1_n14 , _u40_u1_n12 , _u40_u1_n11 , _u40_u1_N5 ,_u40_u1_N4 , _u40_u1_N3 , _u40_u1_rf_ack;
wire  [30:1] dma_req;
wire  [30:1] dma_nd;
wire  [30:1] dma_rest;
wire  [70:0] mast1_pt_in;
wire  [34:0] slv0_pt_in;
wire  [70:0] mast0_pt_in;
wire  [34:0] slv1_pt_in;
wire  [9:2] slv0_adr;
wire  [31:0] slv0_dout;
wire  [31:0] slv0_din;
wire  [22:0] ch0_csr;
wire  [26:0] ch0_txsz;
wire  [31:2] ch0_adr0;
wire  [31:2] ch0_adr1;
wire  [4:0] ch_sel;
wire  [30:0] ndnr;
wire  [31:0] de_csr;
wire  [11:0] de_txsz;
wire  [31:0] de_adr0;
wire  [31:0] de_adr1;
wire  [31:0] csr;
wire  [31:0] pointer;
wire  [31:0] txsz;
wire  [31:0] adr0;
wire  [31:0] adr1;
wire  [31:0] am0;
wire  [31:0] am1;
wire  [31:0] pointer_s;
wire  [31:0] mast0_adr;
wire  [31:0] mast0_dout;
wire  [31:0] mast0_din;
wire  [31:0] mast1_adr;
wire  [31:0] mast1_dout;
wire  [31:0] mast1_din;
wire  [30:15] _u10_ndr_r;
input  [29:0] _u2_adr1_cnt_next1;
input  [29:0] _u2_adr0_cnt_next1;
INV_X4 U8 ( .A(rst_i), .ZN(n5) );
NOR4_X1 _u0_U23819  ( .A1(slv0_adr[7]), .A2(slv0_adr[6]), .A3(slv0_adr[9]),.A4(slv0_adr[8]), .ZN(_u0_n16233 ) );
INV_X1 _u0_U23818  ( .A(slv0_adr[4]), .ZN(_u0_n16029 ) );
AND3_X1 _u0_U23817  ( .A1(_u0_n16233 ), .A2(_u0_n16029 ), .A3(slv0_adr[5]),.ZN(_u0_n16214 ) );
NOR2_X1 _u0_U23816  ( .A1(slv0_adr[2]), .A2(slv0_adr[3]), .ZN(_u0_n16021 ));
AND2_X1 _u0_U23815  ( .A1(_u0_n16214 ), .A2(_u0_n16021 ), .ZN(_u0_n16090 ));
NAND2_X1 _u0_U23814  ( .A1(ch0_csr[0]), .A2(_u0_n16090 ), .ZN(_u0_n16238 ));
INV_X1 _u0_U23813  ( .A(_u0_n16233 ), .ZN(_u0_n16217 ) );
NOR2_X1 _u0_U23812  ( .A1(_u0_n16217 ), .A2(slv0_adr[5]), .ZN(_u0_n16022 ));
NAND2_X1 _u0_U23811  ( .A1(_u0_ch_int_0_ ), .A2(_u0_n16276 ), .ZN(_u0_n16030 ) );
NAND2_X1 _u0_U23810  ( .A1(paused), .A2(_u0_n16021 ), .ZN(_u0_n16247 ) );
MUX2_X1 _u0_U23809  ( .A(_u0_n16030 ), .B(_u0_n16247 ), .S(_u0_n16029 ), .Z(_u0_n16245 ) );
AND2_X1 _u0_U23808  ( .A1(_u0_ch_int_0_ ), .A2(_u0_n16293 ), .ZN(_u0_N3078 ));
NAND2_X1 _u0_U23807  ( .A1(_u0_N3078 ), .A2(slv0_adr[2]), .ZN(_u0_n16246 ));
NAND2_X1 _u0_U23806  ( .A1(_u0_n16245 ), .A2(_u0_n16246 ), .ZN(_u0_n16244 ));
NAND2_X1 _u0_U23805  ( .A1(_u0_n16022 ), .A2(_u0_n16244 ), .ZN(_u0_n16239 ));
INV_X1 _u0_U23804  ( .A(slv0_adr[3]), .ZN(_u0_n16216 ) );
NAND3_X1 _u0_U23803  ( .A1(_u0_n16022 ), .A2(_u0_n16216 ), .A3(slv0_adr[2]),.ZN(_u0_n16026 ) );
NAND2_X1 _u0_U23802  ( .A1(_u0_n16293 ), .A2(_u0_n16042 ), .ZN(_u0_n16240 ));
INV_X1 _u0_U23801  ( .A(slv0_adr[2]), .ZN(_u0_n16232 ) );
NAND3_X1 _u0_U23800  ( .A1(_u0_n16022 ), .A2(_u0_n16232 ), .A3(slv0_adr[3]),.ZN(_u0_n16028 ) );
AND2_X1 _u0_U23799  ( .A1(_u0_n16041 ), .A2(_u0_n16276 ), .ZN(_u0_n16242 ));
AND2_X1 _u0_U23798  ( .A1(ch0_txsz[0]), .A2(_u0_n16064 ), .ZN(_u0_n16243 ));
NOR2_X1 _u0_U23797  ( .A1(_u0_n16242 ), .A2(_u0_n16243 ), .ZN(_u0_n16241 ));
NAND4_X1 _u0_U23796  ( .A1(_u0_n16238 ), .A2(_u0_n16239 ), .A3(_u0_n16240 ),.A4(_u0_n16241 ), .ZN(_u0_N3043 ) );
NAND2_X1 _u0_U23795  ( .A1(ch0_txsz[1]), .A2(_u0_n16064 ), .ZN(_u0_n16234 ));
NAND2_X1 _u0_U23794  ( .A1(_u0_n16277 ), .A2(_u0_n16041 ), .ZN(_u0_n16235 ));
NAND2_X1 _u0_U23793  ( .A1(_u0_n16294 ), .A2(_u0_n16042 ), .ZN(_u0_n16236 ));
NAND2_X1 _u0_U23792  ( .A1(ch0_csr[1]), .A2(_u0_n16090 ), .ZN(_u0_n16237 ));
NAND4_X1 _u0_U23791  ( .A1(_u0_n16234 ), .A2(_u0_n16235 ), .A3(_u0_n16236 ),.A4(_u0_n16237 ), .ZN(_u0_N3044 ) );
NAND2_X1 _u0_U23790  ( .A1(ch0_adr1[2]), .A2(_u0_n16034 ), .ZN(_u0_n16225 ));
NAND2_X1 _u0_U23789  ( .A1(ch0_adr0[2]), .A2(_u0_n16035 ), .ZN(_u0_n16226 ));
NAND2_X1 _u0_U23788  ( .A1(ch0_csr[2]), .A2(_u0_n16090 ), .ZN(_u0_n16227 ));
AND2_X1 _u0_U23787  ( .A1(ch0_txsz[2]), .A2(_u0_n16064 ), .ZN(_u0_n16229 ));
AND2_X1 _u0_U23786  ( .A1(_u0_n16042 ), .A2(_u0_n16274 ), .ZN(_u0_n16230 ));
AND2_X1 _u0_U23785  ( .A1(_u0_n16041 ), .A2(_u0_n16275 ), .ZN(_u0_n16231 ));
NOR3_X1 _u0_U23784  ( .A1(_u0_n16229 ), .A2(_u0_n16230 ), .A3(_u0_n16231 ),.ZN(_u0_n16228 ) );
NAND4_X1 _u0_U23783  ( .A1(_u0_n16225 ), .A2(_u0_n16226 ), .A3(_u0_n16227 ),.A4(_u0_n16228 ), .ZN(_u0_N3045 ) );
NAND2_X1 _u0_U23782  ( .A1(ch0_adr1[3]), .A2(_u0_n16034 ), .ZN(_u0_n16218 ));
NAND2_X1 _u0_U23781  ( .A1(ch0_adr0[3]), .A2(_u0_n16035 ), .ZN(_u0_n16219 ));
NAND2_X1 _u0_U23780  ( .A1(ch0_csr[3]), .A2(_u0_n16090 ), .ZN(_u0_n16220 ));
AND2_X1 _u0_U23779  ( .A1(ch0_txsz[3]), .A2(_u0_n16064 ), .ZN(_u0_n16222 ));
AND2_X1 _u0_U23778  ( .A1(_u0_n16042 ), .A2(_u0_n16272 ), .ZN(_u0_n16223 ));
AND2_X1 _u0_U23777  ( .A1(_u0_n16041 ), .A2(_u0_n16273 ), .ZN(_u0_n16224 ));
NOR3_X1 _u0_U23776  ( .A1(_u0_n16222 ), .A2(_u0_n16223 ), .A3(_u0_n16224 ),.ZN(_u0_n16221 ) );
NAND4_X1 _u0_U23775  ( .A1(_u0_n16218 ), .A2(_u0_n16219 ), .A3(_u0_n16220 ),.A4(_u0_n16221 ), .ZN(_u0_N3046 ) );
NAND2_X1 _u0_U23774  ( .A1(_u0_n16278 ), .A2(_u0_n16041 ), .ZN(_u0_n16206 ));
NAND2_X1 _u0_U23773  ( .A1(_u0_n16295 ), .A2(_u0_n16042 ), .ZN(_u0_n16207 ));
NAND2_X1 _u0_U23772  ( .A1(ch0_txsz[4]), .A2(_u0_n16064 ), .ZN(_u0_n16208 ));
NAND2_X1 _u0_U23771  ( .A1(ch0_csr[4]), .A2(_u0_n16090 ), .ZN(_u0_n16210 ));
NAND2_X1 _u0_U23770  ( .A1(ch0_adr1[4]), .A2(_u0_n16034 ), .ZN(_u0_n16211 ));
NAND2_X1 _u0_U23769  ( .A1(ch0_adr0[4]), .A2(_u0_n16035 ), .ZN(_u0_n16212 ));
NOR2_X1 _u0_U23768  ( .A1(_u0_n16217 ), .A2(_u0_n16029 ), .ZN(_u0_n16215 ));
MUX2_X1 _u0_U23767  ( .A(_u0_n16214 ), .B(_u0_n16215 ), .S(_u0_n16216 ), .Z(_u0_n16213 ) );
AND4_X1 _u0_U23766  ( .A1(_u0_n16210 ), .A2(_u0_n16211 ), .A3(_u0_n16212 ),.A4(_u0_n16032 ), .ZN(_u0_n16209 ) );
NAND4_X1 _u0_U23765  ( .A1(_u0_n16206 ), .A2(_u0_n16207 ), .A3(_u0_n16208 ),.A4(_u0_n16209 ), .ZN(_u0_N3047 ) );
NAND2_X1 _u0_U23764  ( .A1(_u0_n16279 ), .A2(_u0_n16041 ), .ZN(_u0_n16199 ));
NAND2_X1 _u0_U23763  ( .A1(_u0_n16296 ), .A2(_u0_n16042 ), .ZN(_u0_n16200 ));
NAND2_X1 _u0_U23762  ( .A1(ch0_txsz[5]), .A2(_u0_n16064 ), .ZN(_u0_n16201 ));
NAND2_X1 _u0_U23761  ( .A1(ch0_csr[5]), .A2(_u0_n16090 ), .ZN(_u0_n16203 ));
NAND2_X1 _u0_U23760  ( .A1(ch0_adr1[5]), .A2(_u0_n16034 ), .ZN(_u0_n16204 ));
NAND2_X1 _u0_U23759  ( .A1(ch0_adr0[5]), .A2(_u0_n16035 ), .ZN(_u0_n16205 ));
AND4_X1 _u0_U23758  ( .A1(_u0_n16203 ), .A2(_u0_n16204 ), .A3(_u0_n16205 ),.A4(_u0_n16032 ), .ZN(_u0_n16202 ) );
NAND4_X1 _u0_U23757  ( .A1(_u0_n16199 ), .A2(_u0_n16200 ), .A3(_u0_n16201 ),.A4(_u0_n16202 ), .ZN(_u0_N3048 ) );
NAND2_X1 _u0_U23756  ( .A1(_u0_n16280 ), .A2(_u0_n16041 ), .ZN(_u0_n16192 ));
NAND2_X1 _u0_U23755  ( .A1(_u0_n16297 ), .A2(_u0_n16042 ), .ZN(_u0_n16193 ));
NAND2_X1 _u0_U23754  ( .A1(ch0_txsz[6]), .A2(_u0_n16064 ), .ZN(_u0_n16194 ));
NAND2_X1 _u0_U23753  ( .A1(ch0_csr[6]), .A2(_u0_n16090 ), .ZN(_u0_n16196 ));
NAND2_X1 _u0_U23752  ( .A1(ch0_adr1[6]), .A2(_u0_n16034 ), .ZN(_u0_n16197 ));
NAND2_X1 _u0_U23751  ( .A1(ch0_adr0[6]), .A2(_u0_n16035 ), .ZN(_u0_n16198 ));
AND4_X1 _u0_U23750  ( .A1(_u0_n16196 ), .A2(_u0_n16197 ), .A3(_u0_n16198 ),.A4(_u0_n16032 ), .ZN(_u0_n16195 ) );
NAND4_X1 _u0_U23749  ( .A1(_u0_n16192 ), .A2(_u0_n16193 ), .A3(_u0_n16194 ),.A4(_u0_n16195 ), .ZN(_u0_N3049 ) );
NAND2_X1 _u0_U23748  ( .A1(_u0_n16281 ), .A2(_u0_n16041 ), .ZN(_u0_n16185 ));
NAND2_X1 _u0_U23747  ( .A1(_u0_n16298 ), .A2(_u0_n16042 ), .ZN(_u0_n16186 ));
NAND2_X1 _u0_U23746  ( .A1(ch0_txsz[7]), .A2(_u0_n16064 ), .ZN(_u0_n16187 ));
NAND2_X1 _u0_U23745  ( .A1(ch0_csr[7]), .A2(_u0_n16090 ), .ZN(_u0_n16189 ));
NAND2_X1 _u0_U23744  ( .A1(ch0_adr1[7]), .A2(_u0_n16034 ), .ZN(_u0_n16190 ));
NAND2_X1 _u0_U23743  ( .A1(ch0_adr0[7]), .A2(_u0_n16035 ), .ZN(_u0_n16191 ));
AND4_X1 _u0_U23742  ( .A1(_u0_n16189 ), .A2(_u0_n16190 ), .A3(_u0_n16191 ),.A4(_u0_n16032 ), .ZN(_u0_n16188 ) );
NAND4_X1 _u0_U23741  ( .A1(_u0_n16185 ), .A2(_u0_n16186 ), .A3(_u0_n16187 ),.A4(_u0_n16188 ), .ZN(_u0_N3050 ) );
NAND2_X1 _u0_U23740  ( .A1(_u0_n16282 ), .A2(_u0_n16041 ), .ZN(_u0_n16178 ));
NAND2_X1 _u0_U23739  ( .A1(_u0_n16299 ), .A2(_u0_n16042 ), .ZN(_u0_n16179 ));
NAND2_X1 _u0_U23738  ( .A1(ch0_txsz[8]), .A2(_u0_n16064 ), .ZN(_u0_n16180 ));
NAND2_X1 _u0_U23737  ( .A1(ch0_csr[8]), .A2(_u0_n16090 ), .ZN(_u0_n16182 ));
NAND2_X1 _u0_U23736  ( .A1(ch0_adr1[8]), .A2(_u0_n16034 ), .ZN(_u0_n16183 ));
NAND2_X1 _u0_U23735  ( .A1(ch0_adr0[8]), .A2(_u0_n16035 ), .ZN(_u0_n16184 ));
AND4_X1 _u0_U23734  ( .A1(_u0_n16182 ), .A2(_u0_n16183 ), .A3(_u0_n16184 ),.A4(_u0_n16032 ), .ZN(_u0_n16181 ) );
NAND4_X1 _u0_U23733  ( .A1(_u0_n16178 ), .A2(_u0_n16179 ), .A3(_u0_n16180 ),.A4(_u0_n16181 ), .ZN(_u0_N3051 ) );
NAND2_X1 _u0_U23732  ( .A1(ch0_adr0[9]), .A2(_u0_n16035 ), .ZN(_u0_n16172 ));
NAND2_X1 _u0_U23731  ( .A1(ch0_adr1[9]), .A2(_u0_n16034 ), .ZN(_u0_n16173 ));
AND2_X1 _u0_U23730  ( .A1(ch0_txsz[9]), .A2(_u0_n16064 ), .ZN(_u0_n16175 ));
AND2_X1 _u0_U23729  ( .A1(_u0_n16042 ), .A2(_u0_n16271 ), .ZN(_u0_n16176 ));
AND2_X1 _u0_U23728  ( .A1(_u0_n16041 ), .A2(_u0_n16270 ), .ZN(_u0_n16177 ));
NOR3_X1 _u0_U23727  ( .A1(_u0_n16175 ), .A2(_u0_n16176 ), .A3(_u0_n16177 ),.ZN(_u0_n16174 ) );
NAND4_X1 _u0_U23726  ( .A1(_u0_n16172 ), .A2(_u0_n16032 ), .A3(_u0_n16173 ),.A4(_u0_n16174 ), .ZN(_u0_N3052 ) );
NAND2_X1 _u0_U23725  ( .A1(_u0_n16283 ), .A2(_u0_n16041 ), .ZN(_u0_n16165 ));
NAND2_X1 _u0_U23724  ( .A1(_u0_n16300 ), .A2(_u0_n16042 ), .ZN(_u0_n16166 ));
NAND2_X1 _u0_U23723  ( .A1(ch0_txsz[10]), .A2(_u0_n16064 ), .ZN(_u0_n16167 ));
NAND2_X1 _u0_U23722  ( .A1(ch0_csr[10]), .A2(_u0_n16090 ), .ZN(_u0_n16169 ));
NAND2_X1 _u0_U23721  ( .A1(ch0_adr1[10]), .A2(_u0_n16034 ), .ZN(_u0_n16170 ));
NAND2_X1 _u0_U23720  ( .A1(ch0_adr0[10]), .A2(_u0_n16035 ), .ZN(_u0_n16171 ));
AND4_X1 _u0_U23719  ( .A1(_u0_n16169 ), .A2(_u0_n16170 ), .A3(_u0_n16171 ),.A4(_u0_n16032 ), .ZN(_u0_n16168 ) );
NAND4_X1 _u0_U23718  ( .A1(_u0_n16165 ), .A2(_u0_n16166 ), .A3(_u0_n16167 ),.A4(_u0_n16168 ), .ZN(_u0_N3053 ) );
NAND2_X1 _u0_U23717  ( .A1(_u0_n16284 ), .A2(_u0_n16041 ), .ZN(_u0_n16158 ));
NAND2_X1 _u0_U23716  ( .A1(_u0_n16301 ), .A2(_u0_n16042 ), .ZN(_u0_n16159 ));
NAND2_X1 _u0_U23715  ( .A1(ch0_txsz[11]), .A2(_u0_n16064 ), .ZN(_u0_n16160 ));
NAND2_X1 _u0_U23714  ( .A1(ch0_csr[11]), .A2(_u0_n16090 ), .ZN(_u0_n16162 ));
NAND2_X1 _u0_U23713  ( .A1(ch0_adr1[11]), .A2(_u0_n16034 ), .ZN(_u0_n16163 ));
NAND2_X1 _u0_U23712  ( .A1(ch0_adr0[11]), .A2(_u0_n16035 ), .ZN(_u0_n16164 ));
AND4_X1 _u0_U23711  ( .A1(_u0_n16162 ), .A2(_u0_n16163 ), .A3(_u0_n16164 ),.A4(_u0_n16032 ), .ZN(_u0_n16161 ) );
NAND4_X1 _u0_U23710  ( .A1(_u0_n16158 ), .A2(_u0_n16159 ), .A3(_u0_n16160 ),.A4(_u0_n16161 ), .ZN(_u0_N3054 ) );
NAND2_X1 _u0_U23709  ( .A1(ch0_adr0[12]), .A2(_u0_n16035 ), .ZN(_u0_n16152 ));
NAND2_X1 _u0_U23708  ( .A1(ch0_adr1[12]), .A2(_u0_n16034 ), .ZN(_u0_n16153 ));
AND2_X1 _u0_U23707  ( .A1(_u0_n16041 ), .A2(_u0_n16269 ), .ZN(_u0_n16155 ));
AND2_X1 _u0_U23706  ( .A1(ch0_csr[12]), .A2(_u0_n16090 ), .ZN(_u0_n16156 ));
AND2_X1 _u0_U23705  ( .A1(_u0_n16042 ), .A2(_u0_n16268 ), .ZN(_u0_n16157 ));
NOR3_X1 _u0_U23704  ( .A1(_u0_n16155 ), .A2(_u0_n16156 ), .A3(_u0_n16157 ),.ZN(_u0_n16154 ) );
NAND4_X1 _u0_U23703  ( .A1(_u0_n16152 ), .A2(_u0_n16032 ), .A3(_u0_n16153 ),.A4(_u0_n16154 ), .ZN(_u0_N3055 ) );
NAND2_X1 _u0_U23702  ( .A1(ch0_adr0[13]), .A2(_u0_n16035 ), .ZN(_u0_n16146 ));
NAND2_X1 _u0_U23701  ( .A1(ch0_adr1[13]), .A2(_u0_n16034 ), .ZN(_u0_n16147 ));
AND2_X1 _u0_U23700  ( .A1(_u0_n16041 ), .A2(_u0_n16267 ), .ZN(_u0_n16149 ));
AND2_X1 _u0_U23699  ( .A1(ch0_csr[13]), .A2(_u0_n16090 ), .ZN(_u0_n16150 ));
AND2_X1 _u0_U23698  ( .A1(_u0_n16042 ), .A2(_u0_n16266 ), .ZN(_u0_n16151 ));
NOR3_X1 _u0_U23697  ( .A1(_u0_n16149 ), .A2(_u0_n16150 ), .A3(_u0_n16151 ),.ZN(_u0_n16148 ) );
NAND4_X1 _u0_U23696  ( .A1(_u0_n16146 ), .A2(_u0_n16032 ), .A3(_u0_n16147 ),.A4(_u0_n16148 ), .ZN(_u0_N3056 ) );
NAND2_X1 _u0_U23695  ( .A1(ch0_adr0[14]), .A2(_u0_n16035 ), .ZN(_u0_n16140 ));
NAND2_X1 _u0_U23694  ( .A1(ch0_adr1[14]), .A2(_u0_n16034 ), .ZN(_u0_n16141 ));
AND2_X1 _u0_U23693  ( .A1(_u0_n16041 ), .A2(_u0_n16265 ), .ZN(_u0_n16143 ));
AND2_X1 _u0_U23692  ( .A1(ch0_csr[14]), .A2(_u0_n16090 ), .ZN(_u0_n16144 ));
AND2_X1 _u0_U23691  ( .A1(_u0_n16042 ), .A2(_u0_n16264 ), .ZN(_u0_n16145 ));
NOR3_X1 _u0_U23690  ( .A1(_u0_n16143 ), .A2(_u0_n16144 ), .A3(_u0_n16145 ),.ZN(_u0_n16142 ) );
NAND4_X1 _u0_U23689  ( .A1(_u0_n16140 ), .A2(_u0_n16032 ), .A3(_u0_n16141 ),.A4(_u0_n16142 ), .ZN(_u0_N3057 ) );
NAND2_X1 _u0_U23688  ( .A1(_u0_n16285 ), .A2(_u0_n16041 ), .ZN(_u0_n16133 ));
NAND2_X1 _u0_U23687  ( .A1(_u0_n16302 ), .A2(_u0_n16042 ), .ZN(_u0_n16134 ));
NAND2_X1 _u0_U23686  ( .A1(ch0_txsz[15]), .A2(_u0_n16064 ), .ZN(_u0_n16135 ));
NAND2_X1 _u0_U23685  ( .A1(ch0_csr[15]), .A2(_u0_n16090 ), .ZN(_u0_n16137 ));
NAND2_X1 _u0_U23684  ( .A1(ch0_adr1[15]), .A2(_u0_n16034 ), .ZN(_u0_n16138 ));
NAND2_X1 _u0_U23683  ( .A1(ch0_adr0[15]), .A2(_u0_n16035 ), .ZN(_u0_n16139 ));
AND4_X1 _u0_U23682  ( .A1(_u0_n16137 ), .A2(_u0_n16138 ), .A3(_u0_n16139 ),.A4(_u0_n16032 ), .ZN(_u0_n16136 ) );
NAND4_X1 _u0_U23681  ( .A1(_u0_n16133 ), .A2(_u0_n16134 ), .A3(_u0_n16135 ),.A4(_u0_n16136 ), .ZN(_u0_N3058 ) );
NAND2_X1 _u0_U23680  ( .A1(_u0_n16286 ), .A2(_u0_n16041 ), .ZN(_u0_n16126 ));
NAND2_X1 _u0_U23679  ( .A1(_u0_n16303 ), .A2(_u0_n16042 ), .ZN(_u0_n16127 ));
NAND2_X1 _u0_U23678  ( .A1(ch0_txsz[16]), .A2(_u0_n16064 ), .ZN(_u0_n16128 ));
NAND2_X1 _u0_U23677  ( .A1(ch0_csr[16]), .A2(_u0_n16090 ), .ZN(_u0_n16130 ));
NAND2_X1 _u0_U23676  ( .A1(ch0_adr1[16]), .A2(_u0_n16034 ), .ZN(_u0_n16131 ));
NAND2_X1 _u0_U23675  ( .A1(ch0_adr0[16]), .A2(_u0_n16035 ), .ZN(_u0_n16132 ));
AND4_X1 _u0_U23674  ( .A1(_u0_n16130 ), .A2(_u0_n16131 ), .A3(_u0_n16132 ),.A4(_u0_n16032 ), .ZN(_u0_n16129 ) );
NAND4_X1 _u0_U23673  ( .A1(_u0_n16126 ), .A2(_u0_n16127 ), .A3(_u0_n16128 ),.A4(_u0_n16129 ), .ZN(_u0_N3059 ) );
NAND2_X1 _u0_U23672  ( .A1(_u0_n16287 ), .A2(_u0_n16041 ), .ZN(_u0_n16119 ));
NAND2_X1 _u0_U23671  ( .A1(_u0_n16304 ), .A2(_u0_n16042 ), .ZN(_u0_n16120 ));
NAND2_X1 _u0_U23670  ( .A1(ch0_txsz[17]), .A2(_u0_n16064 ), .ZN(_u0_n16121 ));
NAND2_X1 _u0_U23669  ( .A1(ch0_csr[17]), .A2(_u0_n16090 ), .ZN(_u0_n16123 ));
NAND2_X1 _u0_U23668  ( .A1(ch0_adr1[17]), .A2(_u0_n16034 ), .ZN(_u0_n16124 ));
NAND2_X1 _u0_U23667  ( .A1(ch0_adr0[17]), .A2(_u0_n16035 ), .ZN(_u0_n16125 ));
AND4_X1 _u0_U23666  ( .A1(_u0_n16123 ), .A2(_u0_n16124 ), .A3(_u0_n16125 ),.A4(_u0_n16032 ), .ZN(_u0_n16122 ) );
NAND4_X1 _u0_U23665  ( .A1(_u0_n16119 ), .A2(_u0_n16120 ), .A3(_u0_n16121 ),.A4(_u0_n16122 ), .ZN(_u0_N3060 ) );
NAND2_X1 _u0_U23664  ( .A1(_u0_n16288 ), .A2(_u0_n16041 ), .ZN(_u0_n16112 ));
NAND2_X1 _u0_U23663  ( .A1(_u0_n16305 ), .A2(_u0_n16042 ), .ZN(_u0_n16113 ));
NAND2_X1 _u0_U23662  ( .A1(ch0_txsz[18]), .A2(_u0_n16064 ), .ZN(_u0_n16114 ));
NAND2_X1 _u0_U23661  ( .A1(ch0_csr[18]), .A2(_u0_n16090 ), .ZN(_u0_n16116 ));
NAND2_X1 _u0_U23660  ( .A1(ch0_adr1[18]), .A2(_u0_n16034 ), .ZN(_u0_n16117 ));
NAND2_X1 _u0_U23659  ( .A1(ch0_adr0[18]), .A2(_u0_n16035 ), .ZN(_u0_n16118 ));
AND4_X1 _u0_U23658  ( .A1(_u0_n16116 ), .A2(_u0_n16117 ), .A3(_u0_n16118 ),.A4(_u0_n16032 ), .ZN(_u0_n16115 ) );
NAND4_X1 _u0_U23657  ( .A1(_u0_n16112 ), .A2(_u0_n16113 ), .A3(_u0_n16114 ),.A4(_u0_n16115 ), .ZN(_u0_N3061 ) );
NAND2_X1 _u0_U23656  ( .A1(_u0_n16289 ), .A2(_u0_n16041 ), .ZN(_u0_n16105 ));
NAND2_X1 _u0_U23655  ( .A1(_u0_n16306 ), .A2(_u0_n16042 ), .ZN(_u0_n16106 ));
NAND2_X1 _u0_U23654  ( .A1(ch0_txsz[19]), .A2(_u0_n16064 ), .ZN(_u0_n16107 ));
NAND2_X1 _u0_U23653  ( .A1(ch0_csr[19]), .A2(_u0_n16090 ), .ZN(_u0_n16109 ));
NAND2_X1 _u0_U23652  ( .A1(ch0_adr1[19]), .A2(_u0_n16034 ), .ZN(_u0_n16110 ));
NAND2_X1 _u0_U23651  ( .A1(ch0_adr0[19]), .A2(_u0_n16035 ), .ZN(_u0_n16111 ));
AND4_X1 _u0_U23650  ( .A1(_u0_n16109 ), .A2(_u0_n16110 ), .A3(_u0_n16111 ),.A4(_u0_n16032 ), .ZN(_u0_n16108 ) );
NAND4_X1 _u0_U23649  ( .A1(_u0_n16105 ), .A2(_u0_n16106 ), .A3(_u0_n16107 ),.A4(_u0_n16108 ), .ZN(_u0_N3062 ) );
NAND2_X1 _u0_U23648  ( .A1(_u0_n16290 ), .A2(_u0_n16041 ), .ZN(_u0_n16098 ));
NAND2_X1 _u0_U23647  ( .A1(_u0_n16307 ), .A2(_u0_n16042 ), .ZN(_u0_n16099 ));
NAND2_X1 _u0_U23646  ( .A1(ch0_txsz[20]), .A2(_u0_n16064 ), .ZN(_u0_n16100 ));
NAND2_X1 _u0_U23645  ( .A1(ch0_csr[20]), .A2(_u0_n16090 ), .ZN(_u0_n16102 ));
NAND2_X1 _u0_U23644  ( .A1(ch0_adr1[20]), .A2(_u0_n16034 ), .ZN(_u0_n16103 ));
NAND2_X1 _u0_U23643  ( .A1(ch0_adr0[20]), .A2(_u0_n16035 ), .ZN(_u0_n16104 ));
AND4_X1 _u0_U23642  ( .A1(_u0_n16102 ), .A2(_u0_n16103 ), .A3(_u0_n16104 ),.A4(_u0_n16032 ), .ZN(_u0_n16101 ) );
NAND4_X1 _u0_U23641  ( .A1(_u0_n16098 ), .A2(_u0_n16099 ), .A3(_u0_n16100 ),.A4(_u0_n16101 ), .ZN(_u0_N3063 ) );
NAND2_X1 _u0_U23640  ( .A1(_u0_n16291 ), .A2(_u0_n16041 ), .ZN(_u0_n16091 ));
NAND2_X1 _u0_U23639  ( .A1(_u0_n16308 ), .A2(_u0_n16042 ), .ZN(_u0_n16092 ));
NAND2_X1 _u0_U23638  ( .A1(ch0_txsz[21]), .A2(_u0_n16064 ), .ZN(_u0_n16093 ));
NAND2_X1 _u0_U23637  ( .A1(ch0_csr[21]), .A2(_u0_n16090 ), .ZN(_u0_n16095 ));
NAND2_X1 _u0_U23636  ( .A1(ch0_adr1[21]), .A2(_u0_n16034 ), .ZN(_u0_n16096 ));
NAND2_X1 _u0_U23635  ( .A1(ch0_adr0[21]), .A2(_u0_n16035 ), .ZN(_u0_n16097 ));
AND4_X1 _u0_U23634  ( .A1(_u0_n16095 ), .A2(_u0_n16096 ), .A3(_u0_n16097 ),.A4(_u0_n16032 ), .ZN(_u0_n16094 ) );
NAND4_X1 _u0_U23633  ( .A1(_u0_n16091 ), .A2(_u0_n16092 ), .A3(_u0_n16093 ),.A4(_u0_n16094 ), .ZN(_u0_N3064 ) );
NAND2_X1 _u0_U23632  ( .A1(_u0_n16292 ), .A2(_u0_n16041 ), .ZN(_u0_n16083 ));
NAND2_X1 _u0_U23631  ( .A1(_u0_n16309 ), .A2(_u0_n16042 ), .ZN(_u0_n16084 ));
NAND2_X1 _u0_U23630  ( .A1(ch0_txsz[22]), .A2(_u0_n16064 ), .ZN(_u0_n16085 ));
NAND2_X1 _u0_U23629  ( .A1(ch0_csr[22]), .A2(_u0_n16090 ), .ZN(_u0_n16087 ));
NAND2_X1 _u0_U23628  ( .A1(ch0_adr1[22]), .A2(_u0_n16034 ), .ZN(_u0_n16088 ));
NAND2_X1 _u0_U23627  ( .A1(ch0_adr0[22]), .A2(_u0_n16035 ), .ZN(_u0_n16089 ));
AND4_X1 _u0_U23626  ( .A1(_u0_n16087 ), .A2(_u0_n16088 ), .A3(_u0_n16089 ),.A4(_u0_n16032 ), .ZN(_u0_n16086 ) );
NAND4_X1 _u0_U23625  ( .A1(_u0_n16083 ), .A2(_u0_n16084 ), .A3(_u0_n16085 ),.A4(_u0_n16086 ), .ZN(_u0_N3065 ) );
NAND2_X1 _u0_U23624  ( .A1(ch0_adr0[23]), .A2(_u0_n16035 ), .ZN(_u0_n16077 ));
NAND2_X1 _u0_U23623  ( .A1(ch0_adr1[23]), .A2(_u0_n16034 ), .ZN(_u0_n16078 ));
AND2_X1 _u0_U23622  ( .A1(ch0_txsz[23]), .A2(_u0_n16064 ), .ZN(_u0_n16080 ));
AND2_X1 _u0_U23621  ( .A1(_u0_n16042 ), .A2(_u0_n16263 ), .ZN(_u0_n16081 ));
AND2_X1 _u0_U23620  ( .A1(_u0_n16041 ), .A2(_u0_n16262 ), .ZN(_u0_n16082 ));
NOR3_X1 _u0_U23619  ( .A1(_u0_n16080 ), .A2(_u0_n16081 ), .A3(_u0_n16082 ),.ZN(_u0_n16079 ) );
NAND4_X1 _u0_U23618  ( .A1(_u0_n16077 ), .A2(_u0_n16032 ), .A3(_u0_n16078 ),.A4(_u0_n16079 ), .ZN(_u0_N3066 ) );
NAND2_X1 _u0_U23617  ( .A1(ch0_adr0[24]), .A2(_u0_n16035 ), .ZN(_u0_n16071 ));
NAND2_X1 _u0_U23616  ( .A1(ch0_adr1[24]), .A2(_u0_n16034 ), .ZN(_u0_n16072 ));
AND2_X1 _u0_U23615  ( .A1(ch0_txsz[24]), .A2(_u0_n16064 ), .ZN(_u0_n16074 ));
AND2_X1 _u0_U23614  ( .A1(_u0_n16042 ), .A2(_u0_n16261 ), .ZN(_u0_n16075 ));
AND2_X1 _u0_U23613  ( .A1(_u0_n16041 ), .A2(_u0_n16260 ), .ZN(_u0_n16076 ));
NOR3_X1 _u0_U23612  ( .A1(_u0_n16074 ), .A2(_u0_n16075 ), .A3(_u0_n16076 ),.ZN(_u0_n16073 ) );
NAND4_X1 _u0_U23611  ( .A1(_u0_n16071 ), .A2(_u0_n16032 ), .A3(_u0_n16072 ),.A4(_u0_n16073 ), .ZN(_u0_N3067 ) );
NAND2_X1 _u0_U23610  ( .A1(ch0_adr0[25]), .A2(_u0_n16035 ), .ZN(_u0_n16065 ));
NAND2_X1 _u0_U23609  ( .A1(ch0_adr1[25]), .A2(_u0_n16034 ), .ZN(_u0_n16066 ));
AND2_X1 _u0_U23608  ( .A1(ch0_txsz[25]), .A2(_u0_n16064 ), .ZN(_u0_n16068 ));
AND2_X1 _u0_U23607  ( .A1(_u0_n16042 ), .A2(_u0_n16259 ), .ZN(_u0_n16069 ));
AND2_X1 _u0_U23606  ( .A1(_u0_n16041 ), .A2(_u0_n16258 ), .ZN(_u0_n16070 ));
NOR3_X1 _u0_U23605  ( .A1(_u0_n16068 ), .A2(_u0_n16069 ), .A3(_u0_n16070 ),.ZN(_u0_n16067 ) );
NAND4_X1 _u0_U23604  ( .A1(_u0_n16065 ), .A2(_u0_n16032 ), .A3(_u0_n16066 ),.A4(_u0_n16067 ), .ZN(_u0_N3068 ) );
NAND2_X1 _u0_U23603  ( .A1(ch0_adr0[26]), .A2(_u0_n16035 ), .ZN(_u0_n16058 ));
NAND2_X1 _u0_U23602  ( .A1(ch0_adr1[26]), .A2(_u0_n16034 ), .ZN(_u0_n16059 ));
AND2_X1 _u0_U23601  ( .A1(ch0_txsz[26]), .A2(_u0_n16064 ), .ZN(_u0_n16061 ));
AND2_X1 _u0_U23600  ( .A1(_u0_n16042 ), .A2(_u0_n16257 ), .ZN(_u0_n16062 ));
AND2_X1 _u0_U23599  ( .A1(_u0_n16041 ), .A2(_u0_n16256 ), .ZN(_u0_n16063 ));
NOR3_X1 _u0_U23598  ( .A1(_u0_n16061 ), .A2(_u0_n16062 ), .A3(_u0_n16063 ),.ZN(_u0_n16060 ) );
NAND4_X1 _u0_U23597  ( .A1(_u0_n16058 ), .A2(_u0_n16032 ), .A3(_u0_n16059 ),.A4(_u0_n16060 ), .ZN(_u0_N3069 ) );
NAND2_X1 _u0_U23596  ( .A1(ch0_adr0[27]), .A2(_u0_n16035 ), .ZN(_u0_n16053 ));
NAND2_X1 _u0_U23595  ( .A1(ch0_adr1[27]), .A2(_u0_n16034 ), .ZN(_u0_n16054 ));
AND2_X1 _u0_U23594  ( .A1(_u0_n16042 ), .A2(_u0_n16254 ), .ZN(_u0_n16056 ));
AND2_X1 _u0_U23593  ( .A1(_u0_n16041 ), .A2(_u0_n16255 ), .ZN(_u0_n16057 ));
NOR2_X1 _u0_U23592  ( .A1(_u0_n16056 ), .A2(_u0_n16057 ), .ZN(_u0_n16055 ));
NAND4_X1 _u0_U23591  ( .A1(_u0_n16053 ), .A2(_u0_n16032 ), .A3(_u0_n16054 ),.A4(_u0_n16055 ), .ZN(_u0_N3070 ) );
NAND2_X1 _u0_U23590  ( .A1(ch0_adr0[28]), .A2(_u0_n16035 ), .ZN(_u0_n16048 ));
NAND2_X1 _u0_U23589  ( .A1(ch0_adr1[28]), .A2(_u0_n16034 ), .ZN(_u0_n16049 ));
AND2_X1 _u0_U23588  ( .A1(_u0_n16042 ), .A2(_u0_n16252 ), .ZN(_u0_n16051 ));
AND2_X1 _u0_U23587  ( .A1(_u0_n16041 ), .A2(_u0_n16253 ), .ZN(_u0_n16052 ));
NOR2_X1 _u0_U23586  ( .A1(_u0_n16051 ), .A2(_u0_n16052 ), .ZN(_u0_n16050 ));
NAND4_X1 _u0_U23585  ( .A1(_u0_n16048 ), .A2(_u0_n16032 ), .A3(_u0_n16049 ),.A4(_u0_n16050 ), .ZN(_u0_N3071 ) );
NAND2_X1 _u0_U23584  ( .A1(ch0_adr0[29]), .A2(_u0_n16035 ), .ZN(_u0_n16043 ));
NAND2_X1 _u0_U23583  ( .A1(ch0_adr1[29]), .A2(_u0_n16034 ), .ZN(_u0_n16044 ));
AND2_X1 _u0_U23582  ( .A1(_u0_n16042 ), .A2(_u0_n16250 ), .ZN(_u0_n16046 ));
AND2_X1 _u0_U23581  ( .A1(_u0_n16041 ), .A2(_u0_n16251 ), .ZN(_u0_n16047 ));
NOR2_X1 _u0_U23580  ( .A1(_u0_n16046 ), .A2(_u0_n16047 ), .ZN(_u0_n16045 ));
NAND4_X1 _u0_U23579  ( .A1(_u0_n16043 ), .A2(_u0_n16032 ), .A3(_u0_n16044 ),.A4(_u0_n16045 ), .ZN(_u0_N3072 ) );
NAND2_X1 _u0_U23578  ( .A1(ch0_adr0[30]), .A2(_u0_n16035 ), .ZN(_u0_n16036 ));
NAND2_X1 _u0_U23577  ( .A1(ch0_adr1[30]), .A2(_u0_n16034 ), .ZN(_u0_n16037 ));
AND2_X1 _u0_U23576  ( .A1(_u0_n16042 ), .A2(_u0_n16248 ), .ZN(_u0_n16039 ));
AND2_X1 _u0_U23575  ( .A1(_u0_n16041 ), .A2(_u0_n16249 ), .ZN(_u0_n16040 ));
NOR2_X1 _u0_U23574  ( .A1(_u0_n16039 ), .A2(_u0_n16040 ), .ZN(_u0_n16038 ));
NAND4_X1 _u0_U23573  ( .A1(_u0_n16036 ), .A2(_u0_n16032 ), .A3(_u0_n16037 ),.A4(_u0_n16038 ), .ZN(_u0_N3073 ) );
NAND2_X1 _u0_U23572  ( .A1(ch0_adr0[31]), .A2(_u0_n16035 ), .ZN(_u0_n16031 ));
NAND2_X1 _u0_U23571  ( .A1(ch0_adr1[31]), .A2(_u0_n16034 ), .ZN(_u0_n16033 ));
NAND3_X1 _u0_U23570  ( .A1(_u0_n16031 ), .A2(_u0_n16032 ), .A3(_u0_n16033 ),.ZN(_u0_N3074 ) );
INV_X1 _u0_U23569  ( .A(_u0_n16030 ), .ZN(_u0_n453 ) );
NAND2_X1 _u0_U23568  ( .A1(slv0_we), .A2(_u0_n16029 ), .ZN(_u0_n16024 ) );
MUX2_X1 _u0_U23567  ( .A(_u0_n16276 ), .B(slv0_dout[0]), .S(_u0_n16027 ),.Z(_u0_n853 ) );
MUX2_X1 _u0_U23566  ( .A(_u0_n16277 ), .B(slv0_dout[1]), .S(_u0_n16027 ),.Z(_u0_n854 ) );
MUX2_X1 _u0_U23565  ( .A(_u0_n16275 ), .B(slv0_dout[2]), .S(_u0_n16027 ),.Z(_u0_n855 ) );
MUX2_X1 _u0_U23564  ( .A(_u0_n16273 ), .B(slv0_dout[3]), .S(_u0_n16027 ),.Z(_u0_n856 ) );
MUX2_X1 _u0_U23563  ( .A(_u0_n16278 ), .B(slv0_dout[4]), .S(_u0_n16027 ),.Z(_u0_n857 ) );
MUX2_X1 _u0_U23562  ( .A(_u0_n16279 ), .B(slv0_dout[5]), .S(_u0_n16027 ),.Z(_u0_n858 ) );
MUX2_X1 _u0_U23561  ( .A(_u0_n16280 ), .B(slv0_dout[6]), .S(_u0_n16027 ),.Z(_u0_n859 ) );
MUX2_X1 _u0_U23560  ( .A(_u0_n16281 ), .B(slv0_dout[7]), .S(_u0_n16027 ),.Z(_u0_n860 ) );
MUX2_X1 _u0_U23559  ( .A(_u0_n16282 ), .B(slv0_dout[8]), .S(_u0_n16027 ),.Z(_u0_n861 ) );
MUX2_X1 _u0_U23558  ( .A(_u0_n16270 ), .B(slv0_dout[9]), .S(_u0_n16027 ),.Z(_u0_n862 ) );
MUX2_X1 _u0_U23557  ( .A(_u0_n16283 ), .B(slv0_dout[10]), .S(_u0_n16027 ),.Z(_u0_n863 ) );
MUX2_X1 _u0_U23556  ( .A(_u0_n16284 ), .B(slv0_dout[11]), .S(_u0_n16027 ),.Z(_u0_n864 ) );
MUX2_X1 _u0_U23555  ( .A(_u0_n16269 ), .B(slv0_dout[12]), .S(_u0_n16027 ),.Z(_u0_n865 ) );
MUX2_X1 _u0_U23554  ( .A(_u0_n16267 ), .B(slv0_dout[13]), .S(_u0_n16027 ),.Z(_u0_n866 ) );
MUX2_X1 _u0_U23553  ( .A(_u0_n16265 ), .B(slv0_dout[14]), .S(_u0_n16027 ),.Z(_u0_n867 ) );
MUX2_X1 _u0_U23552  ( .A(_u0_n16285 ), .B(slv0_dout[15]), .S(_u0_n16027 ),.Z(_u0_n868 ) );
MUX2_X1 _u0_U23551  ( .A(_u0_n16286 ), .B(slv0_dout[16]), .S(_u0_n16027 ),.Z(_u0_n869 ) );
MUX2_X1 _u0_U23550  ( .A(_u0_n16287 ), .B(slv0_dout[17]), .S(_u0_n16027 ),.Z(_u0_n870 ) );
MUX2_X1 _u0_U23549  ( .A(_u0_n16288 ), .B(slv0_dout[18]), .S(_u0_n16027 ),.Z(_u0_n871 ) );
MUX2_X1 _u0_U23548  ( .A(_u0_n16289 ), .B(slv0_dout[19]), .S(_u0_n16027 ),.Z(_u0_n872 ) );
MUX2_X1 _u0_U23547  ( .A(_u0_n16290 ), .B(slv0_dout[20]), .S(_u0_n16027 ),.Z(_u0_n873 ) );
MUX2_X1 _u0_U23546  ( .A(_u0_n16291 ), .B(slv0_dout[21]), .S(_u0_n16027 ),.Z(_u0_n874 ) );
MUX2_X1 _u0_U23545  ( .A(_u0_n16292 ), .B(slv0_dout[22]), .S(_u0_n16027 ),.Z(_u0_n875 ) );
MUX2_X1 _u0_U23544  ( .A(_u0_n16262 ), .B(slv0_dout[23]), .S(_u0_n16027 ),.Z(_u0_n876 ) );
MUX2_X1 _u0_U23543  ( .A(_u0_n16260 ), .B(slv0_dout[24]), .S(_u0_n16027 ),.Z(_u0_n877 ) );
MUX2_X1 _u0_U23542  ( .A(_u0_n16258 ), .B(slv0_dout[25]), .S(_u0_n16027 ),.Z(_u0_n878 ) );
MUX2_X1 _u0_U23541  ( .A(_u0_n16256 ), .B(slv0_dout[26]), .S(_u0_n16027 ),.Z(_u0_n879 ) );
MUX2_X1 _u0_U23540  ( .A(_u0_n16255 ), .B(slv0_dout[27]), .S(_u0_n16027 ),.Z(_u0_n880 ) );
MUX2_X1 _u0_U23539  ( .A(_u0_n16253 ), .B(slv0_dout[28]), .S(_u0_n16027 ),.Z(_u0_n881 ) );
MUX2_X1 _u0_U23538  ( .A(_u0_n16251 ), .B(slv0_dout[29]), .S(_u0_n16027 ),.Z(_u0_n882 ) );
MUX2_X1 _u0_U23537  ( .A(_u0_n16249 ), .B(slv0_dout[30]), .S(_u0_n16027 ),.Z(_u0_n883 ) );
MUX2_X1 _u0_U23536  ( .A(_u0_n16293 ), .B(slv0_dout[0]), .S(_u0_n16025 ),.Z(_u0_n884 ) );
MUX2_X1 _u0_U23535  ( .A(_u0_n16294 ), .B(slv0_dout[1]), .S(_u0_n16025 ),.Z(_u0_n885 ) );
MUX2_X1 _u0_U23534  ( .A(_u0_n16274 ), .B(slv0_dout[2]), .S(_u0_n16025 ),.Z(_u0_n886 ) );
MUX2_X1 _u0_U23533  ( .A(_u0_n16272 ), .B(slv0_dout[3]), .S(_u0_n16025 ),.Z(_u0_n887 ) );
MUX2_X1 _u0_U23532  ( .A(_u0_n16295 ), .B(slv0_dout[4]), .S(_u0_n16025 ),.Z(_u0_n888 ) );
MUX2_X1 _u0_U23531  ( .A(_u0_n16296 ), .B(slv0_dout[5]), .S(_u0_n16025 ),.Z(_u0_n889 ) );
MUX2_X1 _u0_U23530  ( .A(_u0_n16297 ), .B(slv0_dout[6]), .S(_u0_n16025 ),.Z(_u0_n890 ) );
MUX2_X1 _u0_U23529  ( .A(_u0_n16298 ), .B(slv0_dout[7]), .S(_u0_n16025 ),.Z(_u0_n891 ) );
MUX2_X1 _u0_U23528  ( .A(_u0_n16299 ), .B(slv0_dout[8]), .S(_u0_n16025 ),.Z(_u0_n892 ) );
MUX2_X1 _u0_U23527  ( .A(_u0_n16271 ), .B(slv0_dout[9]), .S(_u0_n16025 ),.Z(_u0_n893 ) );
MUX2_X1 _u0_U23526  ( .A(_u0_n16300 ), .B(slv0_dout[10]), .S(_u0_n16025 ),.Z(_u0_n894 ) );
MUX2_X1 _u0_U23525  ( .A(_u0_n16301 ), .B(slv0_dout[11]), .S(_u0_n16025 ),.Z(_u0_n895 ) );
MUX2_X1 _u0_U23524  ( .A(_u0_n16268 ), .B(slv0_dout[12]), .S(_u0_n16025 ),.Z(_u0_n896 ) );
MUX2_X1 _u0_U23523  ( .A(_u0_n16266 ), .B(slv0_dout[13]), .S(_u0_n16025 ),.Z(_u0_n897 ) );
MUX2_X1 _u0_U23522  ( .A(_u0_n16264 ), .B(slv0_dout[14]), .S(_u0_n16025 ),.Z(_u0_n898 ) );
MUX2_X1 _u0_U23521  ( .A(_u0_n16302 ), .B(slv0_dout[15]), .S(_u0_n16025 ),.Z(_u0_n899 ) );
MUX2_X1 _u0_U23520  ( .A(_u0_n16303 ), .B(slv0_dout[16]), .S(_u0_n16025 ),.Z(_u0_n900 ) );
MUX2_X1 _u0_U23519  ( .A(_u0_n16304 ), .B(slv0_dout[17]), .S(_u0_n16025 ),.Z(_u0_n901 ) );
MUX2_X1 _u0_U23518  ( .A(_u0_n16305 ), .B(slv0_dout[18]), .S(_u0_n16025 ),.Z(_u0_n902 ) );
MUX2_X1 _u0_U23517  ( .A(_u0_n16306 ), .B(slv0_dout[19]), .S(_u0_n16025 ),.Z(_u0_n903 ) );
MUX2_X1 _u0_U23516  ( .A(_u0_n16307 ), .B(slv0_dout[20]), .S(_u0_n16025 ),.Z(_u0_n904 ) );
MUX2_X1 _u0_U23515  ( .A(_u0_n16308 ), .B(slv0_dout[21]), .S(_u0_n16025 ),.Z(_u0_n905 ) );
MUX2_X1 _u0_U23514  ( .A(_u0_n16309 ), .B(slv0_dout[22]), .S(_u0_n16025 ),.Z(_u0_n906 ) );
MUX2_X1 _u0_U23513  ( .A(_u0_n16263 ), .B(slv0_dout[23]), .S(_u0_n16025 ),.Z(_u0_n907 ) );
MUX2_X1 _u0_U23512  ( .A(_u0_n16261 ), .B(slv0_dout[24]), .S(_u0_n16025 ),.Z(_u0_n908 ) );
MUX2_X1 _u0_U23511  ( .A(_u0_n16259 ), .B(slv0_dout[25]), .S(_u0_n16025 ),.Z(_u0_n909 ) );
MUX2_X1 _u0_U23510  ( .A(_u0_n16257 ), .B(slv0_dout[26]), .S(_u0_n16025 ),.Z(_u0_n910 ) );
MUX2_X1 _u0_U23509  ( .A(_u0_n16254 ), .B(slv0_dout[27]), .S(_u0_n16025 ),.Z(_u0_n911 ) );
MUX2_X1 _u0_U23508  ( .A(_u0_n16252 ), .B(slv0_dout[28]), .S(_u0_n16025 ),.Z(_u0_n912 ) );
MUX2_X1 _u0_U23507  ( .A(_u0_n16250 ), .B(slv0_dout[29]), .S(_u0_n16025 ),.Z(_u0_n913 ) );
MUX2_X1 _u0_U23506  ( .A(_u0_n16248 ), .B(slv0_dout[30]), .S(_u0_n16025 ),.Z(_u0_n914 ) );
INV_X1 _u0_U23505  ( .A(_u0_n16024 ), .ZN(_u0_n16023 ) );
AND3_X1 _u0_U23504  ( .A1(_u0_n16021 ), .A2(_u0_n16022 ), .A3(_u0_n16023 ),.ZN(_u0_n16020 ) );
MUX2_X1 _u0_U23503  ( .A(pause_req), .B(slv0_dout[0]), .S(_u0_n16020 ), .Z(_u0_n915 ) );
INV_X4 _u0_U23502  ( .A(n5), .ZN(_u0_n16019 ) );
INV_X8 _u0_U23501  ( .A(_u0_n16019 ), .ZN(_u0_n16018 ) );
NOR2_X4 _u0_U23500  ( .A1(_u0_n16028 ), .A2(_u0_n16024 ), .ZN(_u0_n16027 ));
INV_X4 _u0_U23499  ( .A(_u0_n16026 ), .ZN(_u0_n16042 ) );
NAND2_X2 _u0_U23498  ( .A1(_u0_n16213 ), .A2(slv0_adr[2]), .ZN(_u0_n16032 ));
NOR2_X4 _u0_U23497  ( .A1(_u0_n16026 ), .A2(_u0_n16024 ), .ZN(_u0_n16025 ));
INV_X4 _u0_U23496  ( .A(_u0_n16028 ), .ZN(_u0_n16041 ) );
AND4_X4 _u0_U23495  ( .A1(slv0_adr[5]), .A2(slv0_adr[4]), .A3(_u0_n16021 ),.A4(_u0_n16233 ), .ZN(_u0_n16034 ) );
AND3_X4 _u0_U23494  ( .A1(slv0_adr[2]), .A2(_u0_n16216 ), .A3(_u0_n16214 ),.ZN(_u0_n16064 ) );
AND3_X4 _u0_U23493  ( .A1(slv0_adr[3]), .A2(_u0_n16232 ), .A3(_u0_n16214 ),.ZN(_u0_n16035 ) );
INV_X4 _u0_U23491  ( .A(1'b1), .ZN(_u0_pointer0[31] ) );
INV_X4 _u0_U23489  ( .A(1'b1), .ZN(_u0_pointer0[30] ) );
INV_X4 _u0_U23487  ( .A(1'b1), .ZN(_u0_pointer0[29] ) );
INV_X4 _u0_U23485  ( .A(1'b1), .ZN(_u0_pointer0[28] ) );
INV_X4 _u0_U23483  ( .A(1'b1), .ZN(_u0_pointer0[27] ) );
INV_X4 _u0_U23481  ( .A(1'b1), .ZN(_u0_pointer0[26] ) );
INV_X4 _u0_U23479  ( .A(1'b1), .ZN(_u0_pointer0[25] ) );
INV_X4 _u0_U23477  ( .A(1'b1), .ZN(_u0_pointer0[24] ) );
INV_X4 _u0_U23475  ( .A(1'b1), .ZN(_u0_pointer0[23] ) );
INV_X4 _u0_U23473  ( .A(1'b1), .ZN(_u0_pointer0[22] ) );
INV_X4 _u0_U23471  ( .A(1'b1), .ZN(_u0_pointer0[21] ) );
INV_X4 _u0_U23469  ( .A(1'b1), .ZN(_u0_pointer0[20] ) );
INV_X4 _u0_U23467  ( .A(1'b1), .ZN(_u0_pointer0[19] ) );
INV_X4 _u0_U23465  ( .A(1'b1), .ZN(_u0_pointer0[18] ) );
INV_X4 _u0_U23463  ( .A(1'b1), .ZN(_u0_pointer0[17] ) );
INV_X4 _u0_U23461  ( .A(1'b1), .ZN(_u0_pointer0[16] ) );
INV_X4 _u0_U23459  ( .A(1'b1), .ZN(_u0_pointer0[15] ) );
INV_X4 _u0_U23457  ( .A(1'b1), .ZN(_u0_pointer0[14] ) );
INV_X4 _u0_U23455  ( .A(1'b1), .ZN(_u0_pointer0[13] ) );
INV_X4 _u0_U23453  ( .A(1'b1), .ZN(_u0_pointer0[12] ) );
INV_X4 _u0_U23451  ( .A(1'b1), .ZN(_u0_pointer0[11] ) );
INV_X4 _u0_U23449  ( .A(1'b1), .ZN(_u0_pointer0[10] ) );
INV_X4 _u0_U23447  ( .A(1'b1), .ZN(_u0_pointer0[9] ) );
INV_X4 _u0_U23445  ( .A(1'b1), .ZN(_u0_pointer0[8] ) );
INV_X4 _u0_U23443  ( .A(1'b1), .ZN(_u0_pointer0[7] ) );
INV_X4 _u0_U23441  ( .A(1'b1), .ZN(_u0_pointer0[6] ) );
INV_X4 _u0_U23439  ( .A(1'b1), .ZN(_u0_pointer0[5] ) );
INV_X4 _u0_U23437  ( .A(1'b1), .ZN(_u0_pointer0[4] ) );
INV_X4 _u0_U23435  ( .A(1'b1), .ZN(_u0_pointer0[3] ) );
INV_X4 _u0_U23433  ( .A(1'b1), .ZN(_u0_pointer0[2] ) );
INV_X4 _u0_U23431  ( .A(1'b1), .ZN(_u0_pointer0[1] ) );
INV_X4 _u0_U23429  ( .A(1'b1), .ZN(_u0_pointer0[0] ) );
INV_X4 _u0_U23427  ( .A(1'b1), .ZN(_u0_pointer0_s[31] ) );
INV_X4 _u0_U23425  ( .A(1'b1), .ZN(_u0_pointer0_s[30] ) );
INV_X4 _u0_U23423  ( .A(1'b1), .ZN(_u0_pointer0_s[29] ) );
INV_X4 _u0_U23421  ( .A(1'b1), .ZN(_u0_pointer0_s[28] ) );
INV_X4 _u0_U23419  ( .A(1'b1), .ZN(_u0_pointer0_s[27] ) );
INV_X4 _u0_U23417  ( .A(1'b1), .ZN(_u0_pointer0_s[26] ) );
INV_X4 _u0_U23415  ( .A(1'b1), .ZN(_u0_pointer0_s[25] ) );
INV_X4 _u0_U23413  ( .A(1'b1), .ZN(_u0_pointer0_s[24] ) );
INV_X4 _u0_U23411  ( .A(1'b1), .ZN(_u0_pointer0_s[23] ) );
INV_X4 _u0_U23409  ( .A(1'b1), .ZN(_u0_pointer0_s[22] ) );
INV_X4 _u0_U23407  ( .A(1'b1), .ZN(_u0_pointer0_s[21] ) );
INV_X4 _u0_U23405  ( .A(1'b1), .ZN(_u0_pointer0_s[20] ) );
INV_X4 _u0_U23403  ( .A(1'b1), .ZN(_u0_pointer0_s[19] ) );
INV_X4 _u0_U23401  ( .A(1'b1), .ZN(_u0_pointer0_s[18] ) );
INV_X4 _u0_U23399  ( .A(1'b1), .ZN(_u0_pointer0_s[17] ) );
INV_X4 _u0_U23397  ( .A(1'b1), .ZN(_u0_pointer0_s[16] ) );
INV_X4 _u0_U23395  ( .A(1'b1), .ZN(_u0_pointer0_s[15] ) );
INV_X4 _u0_U23393  ( .A(1'b1), .ZN(_u0_pointer0_s[14] ) );
INV_X4 _u0_U23391  ( .A(1'b1), .ZN(_u0_pointer0_s[13] ) );
INV_X4 _u0_U23389  ( .A(1'b1), .ZN(_u0_pointer0_s[12] ) );
INV_X4 _u0_U23387  ( .A(1'b1), .ZN(_u0_pointer0_s[11] ) );
INV_X4 _u0_U23385  ( .A(1'b1), .ZN(_u0_pointer0_s[10] ) );
INV_X4 _u0_U23383  ( .A(1'b1), .ZN(_u0_pointer0_s[9] ) );
INV_X4 _u0_U23381  ( .A(1'b1), .ZN(_u0_pointer0_s[8] ) );
INV_X4 _u0_U23379  ( .A(1'b1), .ZN(_u0_pointer0_s[7] ) );
INV_X4 _u0_U23377  ( .A(1'b1), .ZN(_u0_pointer0_s[6] ) );
INV_X4 _u0_U23375  ( .A(1'b1), .ZN(_u0_pointer0_s[5] ) );
INV_X4 _u0_U23373  ( .A(1'b1), .ZN(_u0_pointer0_s[4] ) );
INV_X4 _u0_U23371  ( .A(1'b1), .ZN(_u0_pointer0_s[3] ) );
INV_X4 _u0_U23369  ( .A(1'b1), .ZN(_u0_pointer0_s[2] ) );
INV_X4 _u0_U23367  ( .A(1'b1), .ZN(_u0_pointer0_s[1] ) );
INV_X4 _u0_U23365  ( .A(1'b1), .ZN(_u0_pointer0_s[0] ) );
INV_X4 _u0_U23363  ( .A(1'b1), .ZN(_u0_ch0_csr[31] ) );
INV_X4 _u0_U23361  ( .A(1'b1), .ZN(_u0_ch0_csr[30] ) );
INV_X4 _u0_U23359  ( .A(1'b1), .ZN(_u0_ch0_csr[29] ) );
INV_X4 _u0_U23357  ( .A(1'b1), .ZN(_u0_ch0_csr[28] ) );
INV_X4 _u0_U23355  ( .A(1'b1), .ZN(_u0_ch0_csr[27] ) );
INV_X4 _u0_U23353  ( .A(1'b1), .ZN(_u0_ch0_csr[26] ) );
INV_X4 _u0_U23351  ( .A(1'b1), .ZN(_u0_ch0_csr[25] ) );
INV_X4 _u0_U23349  ( .A(1'b1), .ZN(_u0_ch0_csr[24] ) );
INV_X4 _u0_U23347  ( .A(1'b1), .ZN(_u0_ch0_csr[23] ) );
INV_X4 _u0_U23345  ( .A(1'b1), .ZN(_u0_ch0_csr[9] ) );
INV_X4 _u0_U23343  ( .A(1'b1), .ZN(_u0_ch0_txsz[31] ) );
INV_X4 _u0_U23341  ( .A(1'b1), .ZN(_u0_ch0_txsz[30] ) );
INV_X4 _u0_U23339  ( .A(1'b1), .ZN(_u0_ch0_txsz[29] ) );
INV_X4 _u0_U23337  ( .A(1'b1), .ZN(_u0_ch0_txsz[28] ) );
INV_X4 _u0_U23335  ( .A(1'b1), .ZN(_u0_ch0_txsz[27] ) );
INV_X4 _u0_U23333  ( .A(1'b1), .ZN(_u0_ch0_txsz[14] ) );
INV_X4 _u0_U23331  ( .A(1'b1), .ZN(_u0_ch0_txsz[13] ) );
INV_X4 _u0_U23329  ( .A(1'b1), .ZN(_u0_ch0_txsz[12] ) );
INV_X4 _u0_U23327  ( .A(1'b1), .ZN(_u0_ch0_adr0[1] ) );
INV_X4 _u0_U23325  ( .A(1'b1), .ZN(_u0_ch0_adr0[0] ) );
INV_X4 _u0_U23323  ( .A(1'b1), .ZN(_u0_ch0_adr1[1] ) );
INV_X4 _u0_U23321  ( .A(1'b1), .ZN(_u0_ch0_adr1[0] ) );
INV_X4 _u0_U23319  ( .A(1'b0), .ZN(_u0_ch0_am0[31] ) );
INV_X4 _u0_U23317  ( .A(1'b0), .ZN(_u0_ch0_am0[30] ) );
INV_X4 _u0_U23315  ( .A(1'b0), .ZN(_u0_ch0_am0[29] ) );
INV_X4 _u0_U23313  ( .A(1'b0), .ZN(_u0_ch0_am0[28] ) );
INV_X4 _u0_U23311  ( .A(1'b0), .ZN(_u0_ch0_am0[27] ) );
INV_X4 _u0_U23309  ( .A(1'b0), .ZN(_u0_ch0_am0[26] ) );
INV_X4 _u0_U23307  ( .A(1'b0), .ZN(_u0_ch0_am0[25] ) );
INV_X4 _u0_U23305  ( .A(1'b0), .ZN(_u0_ch0_am0[24] ) );
INV_X4 _u0_U23303  ( .A(1'b0), .ZN(_u0_ch0_am0[23] ) );
INV_X4 _u0_U23301  ( .A(1'b0), .ZN(_u0_ch0_am0[22] ) );
INV_X4 _u0_U23299  ( .A(1'b0), .ZN(_u0_ch0_am0[21] ) );
INV_X4 _u0_U23297  ( .A(1'b0), .ZN(_u0_ch0_am0[20] ) );
INV_X4 _u0_U23295  ( .A(1'b0), .ZN(_u0_ch0_am0[19] ) );
INV_X4 _u0_U23293  ( .A(1'b0), .ZN(_u0_ch0_am0[18] ) );
INV_X4 _u0_U23291  ( .A(1'b0), .ZN(_u0_ch0_am0[17] ) );
INV_X4 _u0_U23289  ( .A(1'b0), .ZN(_u0_ch0_am0[16] ) );
INV_X4 _u0_U23287  ( .A(1'b0), .ZN(_u0_ch0_am0[15] ) );
INV_X4 _u0_U23285  ( .A(1'b0), .ZN(_u0_ch0_am0[14] ) );
INV_X4 _u0_U23283  ( .A(1'b0), .ZN(_u0_ch0_am0[13] ) );
INV_X4 _u0_U23281  ( .A(1'b0), .ZN(_u0_ch0_am0[12] ) );
INV_X4 _u0_U23279  ( .A(1'b0), .ZN(_u0_ch0_am0[11] ) );
INV_X4 _u0_U23277  ( .A(1'b0), .ZN(_u0_ch0_am0[10] ) );
INV_X4 _u0_U23275  ( .A(1'b0), .ZN(_u0_ch0_am0[9] ) );
INV_X4 _u0_U23273  ( .A(1'b0), .ZN(_u0_ch0_am0[8] ) );
INV_X4 _u0_U23271  ( .A(1'b0), .ZN(_u0_ch0_am0[7] ) );
INV_X4 _u0_U23269  ( .A(1'b0), .ZN(_u0_ch0_am0[6] ) );
INV_X4 _u0_U23267  ( .A(1'b0), .ZN(_u0_ch0_am0[5] ) );
INV_X4 _u0_U23265  ( .A(1'b0), .ZN(_u0_ch0_am0[4] ) );
INV_X4 _u0_U23263  ( .A(1'b1), .ZN(_u0_ch0_am0[3] ) );
INV_X4 _u0_U23261  ( .A(1'b1), .ZN(_u0_ch0_am0[2] ) );
INV_X4 _u0_U23259  ( .A(1'b1), .ZN(_u0_ch0_am0[1] ) );
INV_X4 _u0_U23257  ( .A(1'b1), .ZN(_u0_ch0_am0[0] ) );
INV_X4 _u0_U23255  ( .A(1'b0), .ZN(_u0_ch0_am1[31] ) );
INV_X4 _u0_U23253  ( .A(1'b0), .ZN(_u0_ch0_am1[30] ) );
INV_X4 _u0_U23251  ( .A(1'b0), .ZN(_u0_ch0_am1[29] ) );
INV_X4 _u0_U23249  ( .A(1'b0), .ZN(_u0_ch0_am1[28] ) );
INV_X4 _u0_U23247  ( .A(1'b0), .ZN(_u0_ch0_am1[27] ) );
INV_X4 _u0_U23245  ( .A(1'b0), .ZN(_u0_ch0_am1[26] ) );
INV_X4 _u0_U23243  ( .A(1'b0), .ZN(_u0_ch0_am1[25] ) );
INV_X4 _u0_U23241  ( .A(1'b0), .ZN(_u0_ch0_am1[24] ) );
INV_X4 _u0_U23239  ( .A(1'b0), .ZN(_u0_ch0_am1[23] ) );
INV_X4 _u0_U23237  ( .A(1'b0), .ZN(_u0_ch0_am1[22] ) );
INV_X4 _u0_U23235  ( .A(1'b0), .ZN(_u0_ch0_am1[21] ) );
INV_X4 _u0_U23233  ( .A(1'b0), .ZN(_u0_ch0_am1[20] ) );
INV_X4 _u0_U23231  ( .A(1'b0), .ZN(_u0_ch0_am1[19] ) );
INV_X4 _u0_U23229  ( .A(1'b0), .ZN(_u0_ch0_am1[18] ) );
INV_X4 _u0_U23227  ( .A(1'b0), .ZN(_u0_ch0_am1[17] ) );
INV_X4 _u0_U23225  ( .A(1'b0), .ZN(_u0_ch0_am1[16] ) );
INV_X4 _u0_U23223  ( .A(1'b0), .ZN(_u0_ch0_am1[15] ) );
INV_X4 _u0_U23221  ( .A(1'b0), .ZN(_u0_ch0_am1[14] ) );
INV_X4 _u0_U23219  ( .A(1'b0), .ZN(_u0_ch0_am1[13] ) );
INV_X4 _u0_U23217  ( .A(1'b0), .ZN(_u0_ch0_am1[12] ) );
INV_X4 _u0_U23215  ( .A(1'b0), .ZN(_u0_ch0_am1[11] ) );
INV_X4 _u0_U23213  ( .A(1'b0), .ZN(_u0_ch0_am1[10] ) );
INV_X4 _u0_U23211  ( .A(1'b0), .ZN(_u0_ch0_am1[9] ) );
INV_X4 _u0_U23209  ( .A(1'b0), .ZN(_u0_ch0_am1[8] ) );
INV_X4 _u0_U23207  ( .A(1'b0), .ZN(_u0_ch0_am1[7] ) );
INV_X4 _u0_U23205  ( .A(1'b0), .ZN(_u0_ch0_am1[6] ) );
INV_X4 _u0_U23203  ( .A(1'b0), .ZN(_u0_ch0_am1[5] ) );
INV_X4 _u0_U23201  ( .A(1'b0), .ZN(_u0_ch0_am1[4] ) );
INV_X4 _u0_U23199  ( .A(1'b1), .ZN(_u0_ch0_am1[3] ) );
INV_X4 _u0_U23197  ( .A(1'b1), .ZN(_u0_ch0_am1[2] ) );
INV_X4 _u0_U23195  ( .A(1'b1), .ZN(_u0_ch0_am1[1] ) );
INV_X4 _u0_U23193  ( .A(1'b1), .ZN(_u0_ch0_am1[0] ) );
INV_X4 _u0_U23191  ( .A(1'b1), .ZN(_u0_pointer1[31] ) );
INV_X4 _u0_U23189  ( .A(1'b1), .ZN(_u0_pointer1[30] ) );
INV_X4 _u0_U23187  ( .A(1'b1), .ZN(_u0_pointer1[29] ) );
INV_X4 _u0_U23185  ( .A(1'b1), .ZN(_u0_pointer1[28] ) );
INV_X4 _u0_U23183  ( .A(1'b1), .ZN(_u0_pointer1[27] ) );
INV_X4 _u0_U23181  ( .A(1'b1), .ZN(_u0_pointer1[26] ) );
INV_X4 _u0_U23179  ( .A(1'b1), .ZN(_u0_pointer1[25] ) );
INV_X4 _u0_U23177  ( .A(1'b1), .ZN(_u0_pointer1[24] ) );
INV_X4 _u0_U23175  ( .A(1'b1), .ZN(_u0_pointer1[23] ) );
INV_X4 _u0_U23173  ( .A(1'b1), .ZN(_u0_pointer1[22] ) );
INV_X4 _u0_U23171  ( .A(1'b1), .ZN(_u0_pointer1[21] ) );
INV_X4 _u0_U23169  ( .A(1'b1), .ZN(_u0_pointer1[20] ) );
INV_X4 _u0_U23167  ( .A(1'b1), .ZN(_u0_pointer1[19] ) );
INV_X4 _u0_U23165  ( .A(1'b1), .ZN(_u0_pointer1[18] ) );
INV_X4 _u0_U23163  ( .A(1'b1), .ZN(_u0_pointer1[17] ) );
INV_X4 _u0_U23161  ( .A(1'b1), .ZN(_u0_pointer1[16] ) );
INV_X4 _u0_U23159  ( .A(1'b1), .ZN(_u0_pointer1[15] ) );
INV_X4 _u0_U23157  ( .A(1'b1), .ZN(_u0_pointer1[14] ) );
INV_X4 _u0_U23155  ( .A(1'b1), .ZN(_u0_pointer1[13] ) );
INV_X4 _u0_U23153  ( .A(1'b1), .ZN(_u0_pointer1[12] ) );
INV_X4 _u0_U23151  ( .A(1'b1), .ZN(_u0_pointer1[11] ) );
INV_X4 _u0_U23149  ( .A(1'b1), .ZN(_u0_pointer1[10] ) );
INV_X4 _u0_U23147  ( .A(1'b1), .ZN(_u0_pointer1[9] ) );
INV_X4 _u0_U23145  ( .A(1'b1), .ZN(_u0_pointer1[8] ) );
INV_X4 _u0_U23143  ( .A(1'b1), .ZN(_u0_pointer1[7] ) );
INV_X4 _u0_U23141  ( .A(1'b1), .ZN(_u0_pointer1[6] ) );
INV_X4 _u0_U23139  ( .A(1'b1), .ZN(_u0_pointer1[5] ) );
INV_X4 _u0_U23137  ( .A(1'b1), .ZN(_u0_pointer1[4] ) );
INV_X4 _u0_U23135  ( .A(1'b1), .ZN(_u0_pointer1[3] ) );
INV_X4 _u0_U23133  ( .A(1'b1), .ZN(_u0_pointer1[2] ) );
INV_X4 _u0_U23131  ( .A(1'b1), .ZN(_u0_pointer1[1] ) );
INV_X4 _u0_U23129  ( .A(1'b1), .ZN(_u0_pointer1[0] ) );
INV_X4 _u0_U23127  ( .A(1'b1), .ZN(_u0_pointer1_s[31] ) );
INV_X4 _u0_U23125  ( .A(1'b1), .ZN(_u0_pointer1_s[30] ) );
INV_X4 _u0_U23123  ( .A(1'b1), .ZN(_u0_pointer1_s[29] ) );
INV_X4 _u0_U23121  ( .A(1'b1), .ZN(_u0_pointer1_s[28] ) );
INV_X4 _u0_U23119  ( .A(1'b1), .ZN(_u0_pointer1_s[27] ) );
INV_X4 _u0_U23117  ( .A(1'b1), .ZN(_u0_pointer1_s[26] ) );
INV_X4 _u0_U23115  ( .A(1'b1), .ZN(_u0_pointer1_s[25] ) );
INV_X4 _u0_U23113  ( .A(1'b1), .ZN(_u0_pointer1_s[24] ) );
INV_X4 _u0_U23111  ( .A(1'b1), .ZN(_u0_pointer1_s[23] ) );
INV_X4 _u0_U23109  ( .A(1'b1), .ZN(_u0_pointer1_s[22] ) );
INV_X4 _u0_U23107  ( .A(1'b1), .ZN(_u0_pointer1_s[21] ) );
INV_X4 _u0_U23105  ( .A(1'b1), .ZN(_u0_pointer1_s[20] ) );
INV_X4 _u0_U23103  ( .A(1'b1), .ZN(_u0_pointer1_s[19] ) );
INV_X4 _u0_U23101  ( .A(1'b1), .ZN(_u0_pointer1_s[18] ) );
INV_X4 _u0_U23099  ( .A(1'b1), .ZN(_u0_pointer1_s[17] ) );
INV_X4 _u0_U23097  ( .A(1'b1), .ZN(_u0_pointer1_s[16] ) );
INV_X4 _u0_U23095  ( .A(1'b1), .ZN(_u0_pointer1_s[15] ) );
INV_X4 _u0_U23093  ( .A(1'b1), .ZN(_u0_pointer1_s[14] ) );
INV_X4 _u0_U23091  ( .A(1'b1), .ZN(_u0_pointer1_s[13] ) );
INV_X4 _u0_U23089  ( .A(1'b1), .ZN(_u0_pointer1_s[12] ) );
INV_X4 _u0_U23087  ( .A(1'b1), .ZN(_u0_pointer1_s[11] ) );
INV_X4 _u0_U23085  ( .A(1'b1), .ZN(_u0_pointer1_s[10] ) );
INV_X4 _u0_U23083  ( .A(1'b1), .ZN(_u0_pointer1_s[9] ) );
INV_X4 _u0_U23081  ( .A(1'b1), .ZN(_u0_pointer1_s[8] ) );
INV_X4 _u0_U23079  ( .A(1'b1), .ZN(_u0_pointer1_s[7] ) );
INV_X4 _u0_U23077  ( .A(1'b1), .ZN(_u0_pointer1_s[6] ) );
INV_X4 _u0_U23075  ( .A(1'b1), .ZN(_u0_pointer1_s[5] ) );
INV_X4 _u0_U23073  ( .A(1'b1), .ZN(_u0_pointer1_s[4] ) );
INV_X4 _u0_U23071  ( .A(1'b1), .ZN(_u0_pointer1_s[3] ) );
INV_X4 _u0_U23069  ( .A(1'b1), .ZN(_u0_pointer1_s[2] ) );
INV_X4 _u0_U23067  ( .A(1'b1), .ZN(_u0_pointer1_s[1] ) );
INV_X4 _u0_U23065  ( .A(1'b1), .ZN(_u0_pointer1_s[0] ) );
INV_X4 _u0_U23063  ( .A(1'b1), .ZN(_u0_ch1_csr[31] ) );
INV_X4 _u0_U23061  ( .A(1'b1), .ZN(_u0_ch1_csr[30] ) );
INV_X4 _u0_U23059  ( .A(1'b1), .ZN(_u0_ch1_csr[29] ) );
INV_X4 _u0_U23057  ( .A(1'b1), .ZN(_u0_ch1_csr[28] ) );
INV_X4 _u0_U23055  ( .A(1'b1), .ZN(_u0_ch1_csr[27] ) );
INV_X4 _u0_U23053  ( .A(1'b1), .ZN(_u0_ch1_csr[26] ) );
INV_X4 _u0_U23051  ( .A(1'b1), .ZN(_u0_ch1_csr[25] ) );
INV_X4 _u0_U23049  ( .A(1'b1), .ZN(_u0_ch1_csr[24] ) );
INV_X4 _u0_U23047  ( .A(1'b1), .ZN(_u0_ch1_csr[23] ) );
INV_X4 _u0_U23045  ( .A(1'b1), .ZN(_u0_ch1_csr[22] ) );
INV_X4 _u0_U23043  ( .A(1'b1), .ZN(_u0_ch1_csr[21] ) );
INV_X4 _u0_U23041  ( .A(1'b1), .ZN(_u0_ch1_csr[20] ) );
INV_X4 _u0_U23039  ( .A(1'b1), .ZN(_u0_ch1_csr[19] ) );
INV_X4 _u0_U23037  ( .A(1'b1), .ZN(_u0_ch1_csr[18] ) );
INV_X4 _u0_U23035  ( .A(1'b1), .ZN(_u0_ch1_csr[17] ) );
INV_X4 _u0_U23033  ( .A(1'b1), .ZN(_u0_ch1_csr[16] ) );
INV_X4 _u0_U23031  ( .A(1'b1), .ZN(_u0_ch1_csr[15] ) );
INV_X4 _u0_U23029  ( .A(1'b1), .ZN(_u0_ch1_csr[14] ) );
INV_X4 _u0_U23027  ( .A(1'b1), .ZN(_u0_ch1_csr[13] ) );
INV_X4 _u0_U23025  ( .A(1'b1), .ZN(_u0_ch1_csr[12] ) );
INV_X4 _u0_U23023  ( .A(1'b1), .ZN(_u0_ch1_csr[11] ) );
INV_X4 _u0_U23021  ( .A(1'b1), .ZN(_u0_ch1_csr[10] ) );
INV_X4 _u0_U23019  ( .A(1'b1), .ZN(_u0_ch1_csr[9] ) );
INV_X4 _u0_U23017  ( .A(1'b1), .ZN(_u0_ch1_csr[8] ) );
INV_X4 _u0_U23015  ( .A(1'b1), .ZN(_u0_ch1_csr[7] ) );
INV_X4 _u0_U23013  ( .A(1'b1), .ZN(_u0_ch1_csr[6] ) );
INV_X4 _u0_U23011  ( .A(1'b1), .ZN(_u0_ch1_csr[5] ) );
INV_X4 _u0_U23009  ( .A(1'b1), .ZN(_u0_ch1_csr[4] ) );
INV_X4 _u0_U23007  ( .A(1'b1), .ZN(_u0_ch1_csr[3] ) );
INV_X4 _u0_U23005  ( .A(1'b1), .ZN(_u0_ch1_csr[2] ) );
INV_X4 _u0_U23003  ( .A(1'b1), .ZN(_u0_ch1_csr[1] ) );
INV_X4 _u0_U23001  ( .A(1'b1), .ZN(_u0_ch1_csr[0] ) );
INV_X4 _u0_U22999  ( .A(1'b1), .ZN(_u0_ch1_txsz[31] ) );
INV_X4 _u0_U22997  ( .A(1'b1), .ZN(_u0_ch1_txsz[30] ) );
INV_X4 _u0_U22995  ( .A(1'b1), .ZN(_u0_ch1_txsz[29] ) );
INV_X4 _u0_U22993  ( .A(1'b1), .ZN(_u0_ch1_txsz[28] ) );
INV_X4 _u0_U22991  ( .A(1'b1), .ZN(_u0_ch1_txsz[27] ) );
INV_X4 _u0_U22989  ( .A(1'b1), .ZN(_u0_ch1_txsz[26] ) );
INV_X4 _u0_U22987  ( .A(1'b1), .ZN(_u0_ch1_txsz[25] ) );
INV_X4 _u0_U22985  ( .A(1'b1), .ZN(_u0_ch1_txsz[24] ) );
INV_X4 _u0_U22983  ( .A(1'b1), .ZN(_u0_ch1_txsz[23] ) );
INV_X4 _u0_U22981  ( .A(1'b1), .ZN(_u0_ch1_txsz[22] ) );
INV_X4 _u0_U22979  ( .A(1'b1), .ZN(_u0_ch1_txsz[21] ) );
INV_X4 _u0_U22977  ( .A(1'b1), .ZN(_u0_ch1_txsz[20] ) );
INV_X4 _u0_U22975  ( .A(1'b1), .ZN(_u0_ch1_txsz[19] ) );
INV_X4 _u0_U22973  ( .A(1'b1), .ZN(_u0_ch1_txsz[18] ) );
INV_X4 _u0_U22971  ( .A(1'b1), .ZN(_u0_ch1_txsz[17] ) );
INV_X4 _u0_U22969  ( .A(1'b1), .ZN(_u0_ch1_txsz[16] ) );
INV_X4 _u0_U22967  ( .A(1'b1), .ZN(_u0_ch1_txsz[15] ) );
INV_X4 _u0_U22965  ( .A(1'b1), .ZN(_u0_ch1_txsz[14] ) );
INV_X4 _u0_U22963  ( .A(1'b1), .ZN(_u0_ch1_txsz[13] ) );
INV_X4 _u0_U22961  ( .A(1'b1), .ZN(_u0_ch1_txsz[12] ) );
INV_X4 _u0_U22959  ( .A(1'b1), .ZN(_u0_ch1_txsz[11] ) );
INV_X4 _u0_U22957  ( .A(1'b1), .ZN(_u0_ch1_txsz[10] ) );
INV_X4 _u0_U22955  ( .A(1'b1), .ZN(_u0_ch1_txsz[9] ) );
INV_X4 _u0_U22953  ( .A(1'b1), .ZN(_u0_ch1_txsz[8] ) );
INV_X4 _u0_U22951  ( .A(1'b1), .ZN(_u0_ch1_txsz[7] ) );
INV_X4 _u0_U22949  ( .A(1'b1), .ZN(_u0_ch1_txsz[6] ) );
INV_X4 _u0_U22947  ( .A(1'b1), .ZN(_u0_ch1_txsz[5] ) );
INV_X4 _u0_U22945  ( .A(1'b1), .ZN(_u0_ch1_txsz[4] ) );
INV_X4 _u0_U22943  ( .A(1'b1), .ZN(_u0_ch1_txsz[3] ) );
INV_X4 _u0_U22941  ( .A(1'b1), .ZN(_u0_ch1_txsz[2] ) );
INV_X4 _u0_U22939  ( .A(1'b1), .ZN(_u0_ch1_txsz[1] ) );
INV_X4 _u0_U22937  ( .A(1'b1), .ZN(_u0_ch1_txsz[0] ) );
INV_X4 _u0_U22935  ( .A(1'b1), .ZN(_u0_ch1_adr0[31] ) );
INV_X4 _u0_U22933  ( .A(1'b1), .ZN(_u0_ch1_adr0[30] ) );
INV_X4 _u0_U22931  ( .A(1'b1), .ZN(_u0_ch1_adr0[29] ) );
INV_X4 _u0_U22929  ( .A(1'b1), .ZN(_u0_ch1_adr0[28] ) );
INV_X4 _u0_U22927  ( .A(1'b1), .ZN(_u0_ch1_adr0[27] ) );
INV_X4 _u0_U22925  ( .A(1'b1), .ZN(_u0_ch1_adr0[26] ) );
INV_X4 _u0_U22923  ( .A(1'b1), .ZN(_u0_ch1_adr0[25] ) );
INV_X4 _u0_U22921  ( .A(1'b1), .ZN(_u0_ch1_adr0[24] ) );
INV_X4 _u0_U22919  ( .A(1'b1), .ZN(_u0_ch1_adr0[23] ) );
INV_X4 _u0_U22917  ( .A(1'b1), .ZN(_u0_ch1_adr0[22] ) );
INV_X4 _u0_U22915  ( .A(1'b1), .ZN(_u0_ch1_adr0[21] ) );
INV_X4 _u0_U22913  ( .A(1'b1), .ZN(_u0_ch1_adr0[20] ) );
INV_X4 _u0_U22911  ( .A(1'b1), .ZN(_u0_ch1_adr0[19] ) );
INV_X4 _u0_U22909  ( .A(1'b1), .ZN(_u0_ch1_adr0[18] ) );
INV_X4 _u0_U22907  ( .A(1'b1), .ZN(_u0_ch1_adr0[17] ) );
INV_X4 _u0_U22905  ( .A(1'b1), .ZN(_u0_ch1_adr0[16] ) );
INV_X4 _u0_U22903  ( .A(1'b1), .ZN(_u0_ch1_adr0[15] ) );
INV_X4 _u0_U22901  ( .A(1'b1), .ZN(_u0_ch1_adr0[14] ) );
INV_X4 _u0_U22899  ( .A(1'b1), .ZN(_u0_ch1_adr0[13] ) );
INV_X4 _u0_U22897  ( .A(1'b1), .ZN(_u0_ch1_adr0[12] ) );
INV_X4 _u0_U22895  ( .A(1'b1), .ZN(_u0_ch1_adr0[11] ) );
INV_X4 _u0_U22893  ( .A(1'b1), .ZN(_u0_ch1_adr0[10] ) );
INV_X4 _u0_U22891  ( .A(1'b1), .ZN(_u0_ch1_adr0[9] ) );
INV_X4 _u0_U22889  ( .A(1'b1), .ZN(_u0_ch1_adr0[8] ) );
INV_X4 _u0_U22887  ( .A(1'b1), .ZN(_u0_ch1_adr0[7] ) );
INV_X4 _u0_U22885  ( .A(1'b1), .ZN(_u0_ch1_adr0[6] ) );
INV_X4 _u0_U22883  ( .A(1'b1), .ZN(_u0_ch1_adr0[5] ) );
INV_X4 _u0_U22881  ( .A(1'b1), .ZN(_u0_ch1_adr0[4] ) );
INV_X4 _u0_U22879  ( .A(1'b1), .ZN(_u0_ch1_adr0[3] ) );
INV_X4 _u0_U22877  ( .A(1'b1), .ZN(_u0_ch1_adr0[2] ) );
INV_X4 _u0_U22875  ( .A(1'b1), .ZN(_u0_ch1_adr0[1] ) );
INV_X4 _u0_U22873  ( .A(1'b1), .ZN(_u0_ch1_adr0[0] ) );
INV_X4 _u0_U22871  ( .A(1'b1), .ZN(_u0_ch1_adr1[31] ) );
INV_X4 _u0_U22869  ( .A(1'b1), .ZN(_u0_ch1_adr1[30] ) );
INV_X4 _u0_U22867  ( .A(1'b1), .ZN(_u0_ch1_adr1[29] ) );
INV_X4 _u0_U22865  ( .A(1'b1), .ZN(_u0_ch1_adr1[28] ) );
INV_X4 _u0_U22863  ( .A(1'b1), .ZN(_u0_ch1_adr1[27] ) );
INV_X4 _u0_U22861  ( .A(1'b1), .ZN(_u0_ch1_adr1[26] ) );
INV_X4 _u0_U22859  ( .A(1'b1), .ZN(_u0_ch1_adr1[25] ) );
INV_X4 _u0_U22857  ( .A(1'b1), .ZN(_u0_ch1_adr1[24] ) );
INV_X4 _u0_U22855  ( .A(1'b1), .ZN(_u0_ch1_adr1[23] ) );
INV_X4 _u0_U22853  ( .A(1'b1), .ZN(_u0_ch1_adr1[22] ) );
INV_X4 _u0_U22851  ( .A(1'b1), .ZN(_u0_ch1_adr1[21] ) );
INV_X4 _u0_U22849  ( .A(1'b1), .ZN(_u0_ch1_adr1[20] ) );
INV_X4 _u0_U22847  ( .A(1'b1), .ZN(_u0_ch1_adr1[19] ) );
INV_X4 _u0_U22845  ( .A(1'b1), .ZN(_u0_ch1_adr1[18] ) );
INV_X4 _u0_U22843  ( .A(1'b1), .ZN(_u0_ch1_adr1[17] ) );
INV_X4 _u0_U22841  ( .A(1'b1), .ZN(_u0_ch1_adr1[16] ) );
INV_X4 _u0_U22839  ( .A(1'b1), .ZN(_u0_ch1_adr1[15] ) );
INV_X4 _u0_U22837  ( .A(1'b1), .ZN(_u0_ch1_adr1[14] ) );
INV_X4 _u0_U22835  ( .A(1'b1), .ZN(_u0_ch1_adr1[13] ) );
INV_X4 _u0_U22833  ( .A(1'b1), .ZN(_u0_ch1_adr1[12] ) );
INV_X4 _u0_U22831  ( .A(1'b1), .ZN(_u0_ch1_adr1[11] ) );
INV_X4 _u0_U22829  ( .A(1'b1), .ZN(_u0_ch1_adr1[10] ) );
INV_X4 _u0_U22827  ( .A(1'b1), .ZN(_u0_ch1_adr1[9] ) );
INV_X4 _u0_U22825  ( .A(1'b1), .ZN(_u0_ch1_adr1[8] ) );
INV_X4 _u0_U22823  ( .A(1'b1), .ZN(_u0_ch1_adr1[7] ) );
INV_X4 _u0_U22821  ( .A(1'b1), .ZN(_u0_ch1_adr1[6] ) );
INV_X4 _u0_U22819  ( .A(1'b1), .ZN(_u0_ch1_adr1[5] ) );
INV_X4 _u0_U22817  ( .A(1'b1), .ZN(_u0_ch1_adr1[4] ) );
INV_X4 _u0_U22815  ( .A(1'b1), .ZN(_u0_ch1_adr1[3] ) );
INV_X4 _u0_U22813  ( .A(1'b1), .ZN(_u0_ch1_adr1[2] ) );
INV_X4 _u0_U22811  ( .A(1'b1), .ZN(_u0_ch1_adr1[1] ) );
INV_X4 _u0_U22809  ( .A(1'b1), .ZN(_u0_ch1_adr1[0] ) );
INV_X4 _u0_U22807  ( .A(1'b0), .ZN(_u0_ch1_am0[31] ) );
INV_X4 _u0_U22805  ( .A(1'b0), .ZN(_u0_ch1_am0[30] ) );
INV_X4 _u0_U22803  ( .A(1'b0), .ZN(_u0_ch1_am0[29] ) );
INV_X4 _u0_U22801  ( .A(1'b0), .ZN(_u0_ch1_am0[28] ) );
INV_X4 _u0_U22799  ( .A(1'b0), .ZN(_u0_ch1_am0[27] ) );
INV_X4 _u0_U22797  ( .A(1'b0), .ZN(_u0_ch1_am0[26] ) );
INV_X4 _u0_U22795  ( .A(1'b0), .ZN(_u0_ch1_am0[25] ) );
INV_X4 _u0_U22793  ( .A(1'b0), .ZN(_u0_ch1_am0[24] ) );
INV_X4 _u0_U22791  ( .A(1'b0), .ZN(_u0_ch1_am0[23] ) );
INV_X4 _u0_U22789  ( .A(1'b0), .ZN(_u0_ch1_am0[22] ) );
INV_X4 _u0_U22787  ( .A(1'b0), .ZN(_u0_ch1_am0[21] ) );
INV_X4 _u0_U22785  ( .A(1'b0), .ZN(_u0_ch1_am0[20] ) );
INV_X4 _u0_U22783  ( .A(1'b0), .ZN(_u0_ch1_am0[19] ) );
INV_X4 _u0_U22781  ( .A(1'b0), .ZN(_u0_ch1_am0[18] ) );
INV_X4 _u0_U22779  ( .A(1'b0), .ZN(_u0_ch1_am0[17] ) );
INV_X4 _u0_U22777  ( .A(1'b0), .ZN(_u0_ch1_am0[16] ) );
INV_X4 _u0_U22775  ( .A(1'b0), .ZN(_u0_ch1_am0[15] ) );
INV_X4 _u0_U22773  ( .A(1'b0), .ZN(_u0_ch1_am0[14] ) );
INV_X4 _u0_U22771  ( .A(1'b0), .ZN(_u0_ch1_am0[13] ) );
INV_X4 _u0_U22769  ( .A(1'b0), .ZN(_u0_ch1_am0[12] ) );
INV_X4 _u0_U22767  ( .A(1'b0), .ZN(_u0_ch1_am0[11] ) );
INV_X4 _u0_U22765  ( .A(1'b0), .ZN(_u0_ch1_am0[10] ) );
INV_X4 _u0_U22763  ( .A(1'b0), .ZN(_u0_ch1_am0[9] ) );
INV_X4 _u0_U22761  ( .A(1'b0), .ZN(_u0_ch1_am0[8] ) );
INV_X4 _u0_U22759  ( .A(1'b0), .ZN(_u0_ch1_am0[7] ) );
INV_X4 _u0_U22757  ( .A(1'b0), .ZN(_u0_ch1_am0[6] ) );
INV_X4 _u0_U22755  ( .A(1'b0), .ZN(_u0_ch1_am0[5] ) );
INV_X4 _u0_U22753  ( .A(1'b0), .ZN(_u0_ch1_am0[4] ) );
INV_X4 _u0_U22751  ( .A(1'b1), .ZN(_u0_ch1_am0[3] ) );
INV_X4 _u0_U22749  ( .A(1'b1), .ZN(_u0_ch1_am0[2] ) );
INV_X4 _u0_U22747  ( .A(1'b1), .ZN(_u0_ch1_am0[1] ) );
INV_X4 _u0_U22745  ( .A(1'b1), .ZN(_u0_ch1_am0[0] ) );
INV_X4 _u0_U22743  ( .A(1'b0), .ZN(_u0_ch1_am1[31] ) );
INV_X4 _u0_U22741  ( .A(1'b0), .ZN(_u0_ch1_am1[30] ) );
INV_X4 _u0_U22739  ( .A(1'b0), .ZN(_u0_ch1_am1[29] ) );
INV_X4 _u0_U22737  ( .A(1'b0), .ZN(_u0_ch1_am1[28] ) );
INV_X4 _u0_U22735  ( .A(1'b0), .ZN(_u0_ch1_am1[27] ) );
INV_X4 _u0_U22733  ( .A(1'b0), .ZN(_u0_ch1_am1[26] ) );
INV_X4 _u0_U22731  ( .A(1'b0), .ZN(_u0_ch1_am1[25] ) );
INV_X4 _u0_U22729  ( .A(1'b0), .ZN(_u0_ch1_am1[24] ) );
INV_X4 _u0_U22727  ( .A(1'b0), .ZN(_u0_ch1_am1[23] ) );
INV_X4 _u0_U22725  ( .A(1'b0), .ZN(_u0_ch1_am1[22] ) );
INV_X4 _u0_U22723  ( .A(1'b0), .ZN(_u0_ch1_am1[21] ) );
INV_X4 _u0_U22721  ( .A(1'b0), .ZN(_u0_ch1_am1[20] ) );
INV_X4 _u0_U22719  ( .A(1'b0), .ZN(_u0_ch1_am1[19] ) );
INV_X4 _u0_U22717  ( .A(1'b0), .ZN(_u0_ch1_am1[18] ) );
INV_X4 _u0_U22715  ( .A(1'b0), .ZN(_u0_ch1_am1[17] ) );
INV_X4 _u0_U22713  ( .A(1'b0), .ZN(_u0_ch1_am1[16] ) );
INV_X4 _u0_U22711  ( .A(1'b0), .ZN(_u0_ch1_am1[15] ) );
INV_X4 _u0_U22709  ( .A(1'b0), .ZN(_u0_ch1_am1[14] ) );
INV_X4 _u0_U22707  ( .A(1'b0), .ZN(_u0_ch1_am1[13] ) );
INV_X4 _u0_U22705  ( .A(1'b0), .ZN(_u0_ch1_am1[12] ) );
INV_X4 _u0_U22703  ( .A(1'b0), .ZN(_u0_ch1_am1[11] ) );
INV_X4 _u0_U22701  ( .A(1'b0), .ZN(_u0_ch1_am1[10] ) );
INV_X4 _u0_U22699  ( .A(1'b0), .ZN(_u0_ch1_am1[9] ) );
INV_X4 _u0_U22697  ( .A(1'b0), .ZN(_u0_ch1_am1[8] ) );
INV_X4 _u0_U22695  ( .A(1'b0), .ZN(_u0_ch1_am1[7] ) );
INV_X4 _u0_U22693  ( .A(1'b0), .ZN(_u0_ch1_am1[6] ) );
INV_X4 _u0_U22691  ( .A(1'b0), .ZN(_u0_ch1_am1[5] ) );
INV_X4 _u0_U22689  ( .A(1'b0), .ZN(_u0_ch1_am1[4] ) );
INV_X4 _u0_U22687  ( .A(1'b1), .ZN(_u0_ch1_am1[3] ) );
INV_X4 _u0_U22685  ( .A(1'b1), .ZN(_u0_ch1_am1[2] ) );
INV_X4 _u0_U22683  ( .A(1'b1), .ZN(_u0_ch1_am1[1] ) );
INV_X4 _u0_U22681  ( .A(1'b1), .ZN(_u0_ch1_am1[0] ) );
INV_X4 _u0_U22679  ( .A(1'b1), .ZN(_u0_pointer2[31] ) );
INV_X4 _u0_U22677  ( .A(1'b1), .ZN(_u0_pointer2[30] ) );
INV_X4 _u0_U22675  ( .A(1'b1), .ZN(_u0_pointer2[29] ) );
INV_X4 _u0_U22673  ( .A(1'b1), .ZN(_u0_pointer2[28] ) );
INV_X4 _u0_U22671  ( .A(1'b1), .ZN(_u0_pointer2[27] ) );
INV_X4 _u0_U22669  ( .A(1'b1), .ZN(_u0_pointer2[26] ) );
INV_X4 _u0_U22667  ( .A(1'b1), .ZN(_u0_pointer2[25] ) );
INV_X4 _u0_U22665  ( .A(1'b1), .ZN(_u0_pointer2[24] ) );
INV_X4 _u0_U22663  ( .A(1'b1), .ZN(_u0_pointer2[23] ) );
INV_X4 _u0_U22661  ( .A(1'b1), .ZN(_u0_pointer2[22] ) );
INV_X4 _u0_U22659  ( .A(1'b1), .ZN(_u0_pointer2[21] ) );
INV_X4 _u0_U22657  ( .A(1'b1), .ZN(_u0_pointer2[20] ) );
INV_X4 _u0_U22655  ( .A(1'b1), .ZN(_u0_pointer2[19] ) );
INV_X4 _u0_U22653  ( .A(1'b1), .ZN(_u0_pointer2[18] ) );
INV_X4 _u0_U22651  ( .A(1'b1), .ZN(_u0_pointer2[17] ) );
INV_X4 _u0_U22649  ( .A(1'b1), .ZN(_u0_pointer2[16] ) );
INV_X4 _u0_U22647  ( .A(1'b1), .ZN(_u0_pointer2[15] ) );
INV_X4 _u0_U22645  ( .A(1'b1), .ZN(_u0_pointer2[14] ) );
INV_X4 _u0_U22643  ( .A(1'b1), .ZN(_u0_pointer2[13] ) );
INV_X4 _u0_U22641  ( .A(1'b1), .ZN(_u0_pointer2[12] ) );
INV_X4 _u0_U22639  ( .A(1'b1), .ZN(_u0_pointer2[11] ) );
INV_X4 _u0_U22637  ( .A(1'b1), .ZN(_u0_pointer2[10] ) );
INV_X4 _u0_U22635  ( .A(1'b1), .ZN(_u0_pointer2[9] ) );
INV_X4 _u0_U22633  ( .A(1'b1), .ZN(_u0_pointer2[8] ) );
INV_X4 _u0_U22631  ( .A(1'b1), .ZN(_u0_pointer2[7] ) );
INV_X4 _u0_U22629  ( .A(1'b1), .ZN(_u0_pointer2[6] ) );
INV_X4 _u0_U22627  ( .A(1'b1), .ZN(_u0_pointer2[5] ) );
INV_X4 _u0_U22625  ( .A(1'b1), .ZN(_u0_pointer2[4] ) );
INV_X4 _u0_U22623  ( .A(1'b1), .ZN(_u0_pointer2[3] ) );
INV_X4 _u0_U22621  ( .A(1'b1), .ZN(_u0_pointer2[2] ) );
INV_X4 _u0_U22619  ( .A(1'b1), .ZN(_u0_pointer2[1] ) );
INV_X4 _u0_U22617  ( .A(1'b1), .ZN(_u0_pointer2[0] ) );
INV_X4 _u0_U22615  ( .A(1'b1), .ZN(_u0_pointer2_s[31] ) );
INV_X4 _u0_U22613  ( .A(1'b1), .ZN(_u0_pointer2_s[30] ) );
INV_X4 _u0_U22611  ( .A(1'b1), .ZN(_u0_pointer2_s[29] ) );
INV_X4 _u0_U22609  ( .A(1'b1), .ZN(_u0_pointer2_s[28] ) );
INV_X4 _u0_U22607  ( .A(1'b1), .ZN(_u0_pointer2_s[27] ) );
INV_X4 _u0_U22605  ( .A(1'b1), .ZN(_u0_pointer2_s[26] ) );
INV_X4 _u0_U22603  ( .A(1'b1), .ZN(_u0_pointer2_s[25] ) );
INV_X4 _u0_U22601  ( .A(1'b1), .ZN(_u0_pointer2_s[24] ) );
INV_X4 _u0_U22599  ( .A(1'b1), .ZN(_u0_pointer2_s[23] ) );
INV_X4 _u0_U22597  ( .A(1'b1), .ZN(_u0_pointer2_s[22] ) );
INV_X4 _u0_U22595  ( .A(1'b1), .ZN(_u0_pointer2_s[21] ) );
INV_X4 _u0_U22593  ( .A(1'b1), .ZN(_u0_pointer2_s[20] ) );
INV_X4 _u0_U22591  ( .A(1'b1), .ZN(_u0_pointer2_s[19] ) );
INV_X4 _u0_U22589  ( .A(1'b1), .ZN(_u0_pointer2_s[18] ) );
INV_X4 _u0_U22587  ( .A(1'b1), .ZN(_u0_pointer2_s[17] ) );
INV_X4 _u0_U22585  ( .A(1'b1), .ZN(_u0_pointer2_s[16] ) );
INV_X4 _u0_U22583  ( .A(1'b1), .ZN(_u0_pointer2_s[15] ) );
INV_X4 _u0_U22581  ( .A(1'b1), .ZN(_u0_pointer2_s[14] ) );
INV_X4 _u0_U22579  ( .A(1'b1), .ZN(_u0_pointer2_s[13] ) );
INV_X4 _u0_U22577  ( .A(1'b1), .ZN(_u0_pointer2_s[12] ) );
INV_X4 _u0_U22575  ( .A(1'b1), .ZN(_u0_pointer2_s[11] ) );
INV_X4 _u0_U22573  ( .A(1'b1), .ZN(_u0_pointer2_s[10] ) );
INV_X4 _u0_U22571  ( .A(1'b1), .ZN(_u0_pointer2_s[9] ) );
INV_X4 _u0_U22569  ( .A(1'b1), .ZN(_u0_pointer2_s[8] ) );
INV_X4 _u0_U22567  ( .A(1'b1), .ZN(_u0_pointer2_s[7] ) );
INV_X4 _u0_U22565  ( .A(1'b1), .ZN(_u0_pointer2_s[6] ) );
INV_X4 _u0_U22563  ( .A(1'b1), .ZN(_u0_pointer2_s[5] ) );
INV_X4 _u0_U22561  ( .A(1'b1), .ZN(_u0_pointer2_s[4] ) );
INV_X4 _u0_U22559  ( .A(1'b1), .ZN(_u0_pointer2_s[3] ) );
INV_X4 _u0_U22557  ( .A(1'b1), .ZN(_u0_pointer2_s[2] ) );
INV_X4 _u0_U22555  ( .A(1'b1), .ZN(_u0_pointer2_s[1] ) );
INV_X4 _u0_U22553  ( .A(1'b1), .ZN(_u0_pointer2_s[0] ) );
INV_X4 _u0_U22551  ( .A(1'b1), .ZN(_u0_ch2_csr[31] ) );
INV_X4 _u0_U22549  ( .A(1'b1), .ZN(_u0_ch2_csr[30] ) );
INV_X4 _u0_U22547  ( .A(1'b1), .ZN(_u0_ch2_csr[29] ) );
INV_X4 _u0_U22545  ( .A(1'b1), .ZN(_u0_ch2_csr[28] ) );
INV_X4 _u0_U22543  ( .A(1'b1), .ZN(_u0_ch2_csr[27] ) );
INV_X4 _u0_U22541  ( .A(1'b1), .ZN(_u0_ch2_csr[26] ) );
INV_X4 _u0_U22539  ( .A(1'b1), .ZN(_u0_ch2_csr[25] ) );
INV_X4 _u0_U22537  ( .A(1'b1), .ZN(_u0_ch2_csr[24] ) );
INV_X4 _u0_U22535  ( .A(1'b1), .ZN(_u0_ch2_csr[23] ) );
INV_X4 _u0_U22533  ( .A(1'b1), .ZN(_u0_ch2_csr[22] ) );
INV_X4 _u0_U22531  ( .A(1'b1), .ZN(_u0_ch2_csr[21] ) );
INV_X4 _u0_U22529  ( .A(1'b1), .ZN(_u0_ch2_csr[20] ) );
INV_X4 _u0_U22527  ( .A(1'b1), .ZN(_u0_ch2_csr[19] ) );
INV_X4 _u0_U22525  ( .A(1'b1), .ZN(_u0_ch2_csr[18] ) );
INV_X4 _u0_U22523  ( .A(1'b1), .ZN(_u0_ch2_csr[17] ) );
INV_X4 _u0_U22521  ( .A(1'b1), .ZN(_u0_ch2_csr[16] ) );
INV_X4 _u0_U22519  ( .A(1'b1), .ZN(_u0_ch2_csr[15] ) );
INV_X4 _u0_U22517  ( .A(1'b1), .ZN(_u0_ch2_csr[14] ) );
INV_X4 _u0_U22515  ( .A(1'b1), .ZN(_u0_ch2_csr[13] ) );
INV_X4 _u0_U22513  ( .A(1'b1), .ZN(_u0_ch2_csr[12] ) );
INV_X4 _u0_U22511  ( .A(1'b1), .ZN(_u0_ch2_csr[11] ) );
INV_X4 _u0_U22509  ( .A(1'b1), .ZN(_u0_ch2_csr[10] ) );
INV_X4 _u0_U22507  ( .A(1'b1), .ZN(_u0_ch2_csr[9] ) );
INV_X4 _u0_U22505  ( .A(1'b1), .ZN(_u0_ch2_csr[8] ) );
INV_X4 _u0_U22503  ( .A(1'b1), .ZN(_u0_ch2_csr[7] ) );
INV_X4 _u0_U22501  ( .A(1'b1), .ZN(_u0_ch2_csr[6] ) );
INV_X4 _u0_U22499  ( .A(1'b1), .ZN(_u0_ch2_csr[5] ) );
INV_X4 _u0_U22497  ( .A(1'b1), .ZN(_u0_ch2_csr[4] ) );
INV_X4 _u0_U22495  ( .A(1'b1), .ZN(_u0_ch2_csr[3] ) );
INV_X4 _u0_U22493  ( .A(1'b1), .ZN(_u0_ch2_csr[2] ) );
INV_X4 _u0_U22491  ( .A(1'b1), .ZN(_u0_ch2_csr[1] ) );
INV_X4 _u0_U22489  ( .A(1'b1), .ZN(_u0_ch2_csr[0] ) );
INV_X4 _u0_U22487  ( .A(1'b1), .ZN(_u0_ch2_txsz[31] ) );
INV_X4 _u0_U22485  ( .A(1'b1), .ZN(_u0_ch2_txsz[30] ) );
INV_X4 _u0_U22483  ( .A(1'b1), .ZN(_u0_ch2_txsz[29] ) );
INV_X4 _u0_U22481  ( .A(1'b1), .ZN(_u0_ch2_txsz[28] ) );
INV_X4 _u0_U22479  ( .A(1'b1), .ZN(_u0_ch2_txsz[27] ) );
INV_X4 _u0_U22477  ( .A(1'b1), .ZN(_u0_ch2_txsz[26] ) );
INV_X4 _u0_U22475  ( .A(1'b1), .ZN(_u0_ch2_txsz[25] ) );
INV_X4 _u0_U22473  ( .A(1'b1), .ZN(_u0_ch2_txsz[24] ) );
INV_X4 _u0_U22471  ( .A(1'b1), .ZN(_u0_ch2_txsz[23] ) );
INV_X4 _u0_U22469  ( .A(1'b1), .ZN(_u0_ch2_txsz[22] ) );
INV_X4 _u0_U22467  ( .A(1'b1), .ZN(_u0_ch2_txsz[21] ) );
INV_X4 _u0_U22465  ( .A(1'b1), .ZN(_u0_ch2_txsz[20] ) );
INV_X4 _u0_U22463  ( .A(1'b1), .ZN(_u0_ch2_txsz[19] ) );
INV_X4 _u0_U22461  ( .A(1'b1), .ZN(_u0_ch2_txsz[18] ) );
INV_X4 _u0_U22459  ( .A(1'b1), .ZN(_u0_ch2_txsz[17] ) );
INV_X4 _u0_U22457  ( .A(1'b1), .ZN(_u0_ch2_txsz[16] ) );
INV_X4 _u0_U22455  ( .A(1'b1), .ZN(_u0_ch2_txsz[15] ) );
INV_X4 _u0_U22453  ( .A(1'b1), .ZN(_u0_ch2_txsz[14] ) );
INV_X4 _u0_U22451  ( .A(1'b1), .ZN(_u0_ch2_txsz[13] ) );
INV_X4 _u0_U22449  ( .A(1'b1), .ZN(_u0_ch2_txsz[12] ) );
INV_X4 _u0_U22447  ( .A(1'b1), .ZN(_u0_ch2_txsz[11] ) );
INV_X4 _u0_U22445  ( .A(1'b1), .ZN(_u0_ch2_txsz[10] ) );
INV_X4 _u0_U22443  ( .A(1'b1), .ZN(_u0_ch2_txsz[9] ) );
INV_X4 _u0_U22441  ( .A(1'b1), .ZN(_u0_ch2_txsz[8] ) );
INV_X4 _u0_U22439  ( .A(1'b1), .ZN(_u0_ch2_txsz[7] ) );
INV_X4 _u0_U22437  ( .A(1'b1), .ZN(_u0_ch2_txsz[6] ) );
INV_X4 _u0_U22435  ( .A(1'b1), .ZN(_u0_ch2_txsz[5] ) );
INV_X4 _u0_U22433  ( .A(1'b1), .ZN(_u0_ch2_txsz[4] ) );
INV_X4 _u0_U22431  ( .A(1'b1), .ZN(_u0_ch2_txsz[3] ) );
INV_X4 _u0_U22429  ( .A(1'b1), .ZN(_u0_ch2_txsz[2] ) );
INV_X4 _u0_U22427  ( .A(1'b1), .ZN(_u0_ch2_txsz[1] ) );
INV_X4 _u0_U22425  ( .A(1'b1), .ZN(_u0_ch2_txsz[0] ) );
INV_X4 _u0_U22423  ( .A(1'b1), .ZN(_u0_ch2_adr0[31] ) );
INV_X4 _u0_U22421  ( .A(1'b1), .ZN(_u0_ch2_adr0[30] ) );
INV_X4 _u0_U22419  ( .A(1'b1), .ZN(_u0_ch2_adr0[29] ) );
INV_X4 _u0_U22417  ( .A(1'b1), .ZN(_u0_ch2_adr0[28] ) );
INV_X4 _u0_U22415  ( .A(1'b1), .ZN(_u0_ch2_adr0[27] ) );
INV_X4 _u0_U22413  ( .A(1'b1), .ZN(_u0_ch2_adr0[26] ) );
INV_X4 _u0_U22411  ( .A(1'b1), .ZN(_u0_ch2_adr0[25] ) );
INV_X4 _u0_U22409  ( .A(1'b1), .ZN(_u0_ch2_adr0[24] ) );
INV_X4 _u0_U22407  ( .A(1'b1), .ZN(_u0_ch2_adr0[23] ) );
INV_X4 _u0_U22405  ( .A(1'b1), .ZN(_u0_ch2_adr0[22] ) );
INV_X4 _u0_U22403  ( .A(1'b1), .ZN(_u0_ch2_adr0[21] ) );
INV_X4 _u0_U22401  ( .A(1'b1), .ZN(_u0_ch2_adr0[20] ) );
INV_X4 _u0_U22399  ( .A(1'b1), .ZN(_u0_ch2_adr0[19] ) );
INV_X4 _u0_U22397  ( .A(1'b1), .ZN(_u0_ch2_adr0[18] ) );
INV_X4 _u0_U22395  ( .A(1'b1), .ZN(_u0_ch2_adr0[17] ) );
INV_X4 _u0_U22393  ( .A(1'b1), .ZN(_u0_ch2_adr0[16] ) );
INV_X4 _u0_U22391  ( .A(1'b1), .ZN(_u0_ch2_adr0[15] ) );
INV_X4 _u0_U22389  ( .A(1'b1), .ZN(_u0_ch2_adr0[14] ) );
INV_X4 _u0_U22387  ( .A(1'b1), .ZN(_u0_ch2_adr0[13] ) );
INV_X4 _u0_U22385  ( .A(1'b1), .ZN(_u0_ch2_adr0[12] ) );
INV_X4 _u0_U22383  ( .A(1'b1), .ZN(_u0_ch2_adr0[11] ) );
INV_X4 _u0_U22381  ( .A(1'b1), .ZN(_u0_ch2_adr0[10] ) );
INV_X4 _u0_U22379  ( .A(1'b1), .ZN(_u0_ch2_adr0[9] ) );
INV_X4 _u0_U22377  ( .A(1'b1), .ZN(_u0_ch2_adr0[8] ) );
INV_X4 _u0_U22375  ( .A(1'b1), .ZN(_u0_ch2_adr0[7] ) );
INV_X4 _u0_U22373  ( .A(1'b1), .ZN(_u0_ch2_adr0[6] ) );
INV_X4 _u0_U22371  ( .A(1'b1), .ZN(_u0_ch2_adr0[5] ) );
INV_X4 _u0_U22369  ( .A(1'b1), .ZN(_u0_ch2_adr0[4] ) );
INV_X4 _u0_U22367  ( .A(1'b1), .ZN(_u0_ch2_adr0[3] ) );
INV_X4 _u0_U22365  ( .A(1'b1), .ZN(_u0_ch2_adr0[2] ) );
INV_X4 _u0_U22363  ( .A(1'b1), .ZN(_u0_ch2_adr0[1] ) );
INV_X4 _u0_U22361  ( .A(1'b1), .ZN(_u0_ch2_adr0[0] ) );
INV_X4 _u0_U22359  ( .A(1'b1), .ZN(_u0_ch2_adr1[31] ) );
INV_X4 _u0_U22357  ( .A(1'b1), .ZN(_u0_ch2_adr1[30] ) );
INV_X4 _u0_U22355  ( .A(1'b1), .ZN(_u0_ch2_adr1[29] ) );
INV_X4 _u0_U22353  ( .A(1'b1), .ZN(_u0_ch2_adr1[28] ) );
INV_X4 _u0_U22351  ( .A(1'b1), .ZN(_u0_ch2_adr1[27] ) );
INV_X4 _u0_U22349  ( .A(1'b1), .ZN(_u0_ch2_adr1[26] ) );
INV_X4 _u0_U22347  ( .A(1'b1), .ZN(_u0_ch2_adr1[25] ) );
INV_X4 _u0_U22345  ( .A(1'b1), .ZN(_u0_ch2_adr1[24] ) );
INV_X4 _u0_U22343  ( .A(1'b1), .ZN(_u0_ch2_adr1[23] ) );
INV_X4 _u0_U22341  ( .A(1'b1), .ZN(_u0_ch2_adr1[22] ) );
INV_X4 _u0_U22339  ( .A(1'b1), .ZN(_u0_ch2_adr1[21] ) );
INV_X4 _u0_U22337  ( .A(1'b1), .ZN(_u0_ch2_adr1[20] ) );
INV_X4 _u0_U22335  ( .A(1'b1), .ZN(_u0_ch2_adr1[19] ) );
INV_X4 _u0_U22333  ( .A(1'b1), .ZN(_u0_ch2_adr1[18] ) );
INV_X4 _u0_U22331  ( .A(1'b1), .ZN(_u0_ch2_adr1[17] ) );
INV_X4 _u0_U22329  ( .A(1'b1), .ZN(_u0_ch2_adr1[16] ) );
INV_X4 _u0_U22327  ( .A(1'b1), .ZN(_u0_ch2_adr1[15] ) );
INV_X4 _u0_U22325  ( .A(1'b1), .ZN(_u0_ch2_adr1[14] ) );
INV_X4 _u0_U22323  ( .A(1'b1), .ZN(_u0_ch2_adr1[13] ) );
INV_X4 _u0_U22321  ( .A(1'b1), .ZN(_u0_ch2_adr1[12] ) );
INV_X4 _u0_U22319  ( .A(1'b1), .ZN(_u0_ch2_adr1[11] ) );
INV_X4 _u0_U22317  ( .A(1'b1), .ZN(_u0_ch2_adr1[10] ) );
INV_X4 _u0_U22315  ( .A(1'b1), .ZN(_u0_ch2_adr1[9] ) );
INV_X4 _u0_U22313  ( .A(1'b1), .ZN(_u0_ch2_adr1[8] ) );
INV_X4 _u0_U22311  ( .A(1'b1), .ZN(_u0_ch2_adr1[7] ) );
INV_X4 _u0_U22309  ( .A(1'b1), .ZN(_u0_ch2_adr1[6] ) );
INV_X4 _u0_U22307  ( .A(1'b1), .ZN(_u0_ch2_adr1[5] ) );
INV_X4 _u0_U22305  ( .A(1'b1), .ZN(_u0_ch2_adr1[4] ) );
INV_X4 _u0_U22303  ( .A(1'b1), .ZN(_u0_ch2_adr1[3] ) );
INV_X4 _u0_U22301  ( .A(1'b1), .ZN(_u0_ch2_adr1[2] ) );
INV_X4 _u0_U22299  ( .A(1'b1), .ZN(_u0_ch2_adr1[1] ) );
INV_X4 _u0_U22297  ( .A(1'b1), .ZN(_u0_ch2_adr1[0] ) );
INV_X4 _u0_U22295  ( .A(1'b0), .ZN(_u0_ch2_am0[31] ) );
INV_X4 _u0_U22293  ( .A(1'b0), .ZN(_u0_ch2_am0[30] ) );
INV_X4 _u0_U22291  ( .A(1'b0), .ZN(_u0_ch2_am0[29] ) );
INV_X4 _u0_U22289  ( .A(1'b0), .ZN(_u0_ch2_am0[28] ) );
INV_X4 _u0_U22287  ( .A(1'b0), .ZN(_u0_ch2_am0[27] ) );
INV_X4 _u0_U22285  ( .A(1'b0), .ZN(_u0_ch2_am0[26] ) );
INV_X4 _u0_U22283  ( .A(1'b0), .ZN(_u0_ch2_am0[25] ) );
INV_X4 _u0_U22281  ( .A(1'b0), .ZN(_u0_ch2_am0[24] ) );
INV_X4 _u0_U22279  ( .A(1'b0), .ZN(_u0_ch2_am0[23] ) );
INV_X4 _u0_U22277  ( .A(1'b0), .ZN(_u0_ch2_am0[22] ) );
INV_X4 _u0_U22275  ( .A(1'b0), .ZN(_u0_ch2_am0[21] ) );
INV_X4 _u0_U22273  ( .A(1'b0), .ZN(_u0_ch2_am0[20] ) );
INV_X4 _u0_U22271  ( .A(1'b0), .ZN(_u0_ch2_am0[19] ) );
INV_X4 _u0_U22269  ( .A(1'b0), .ZN(_u0_ch2_am0[18] ) );
INV_X4 _u0_U22267  ( .A(1'b0), .ZN(_u0_ch2_am0[17] ) );
INV_X4 _u0_U22265  ( .A(1'b0), .ZN(_u0_ch2_am0[16] ) );
INV_X4 _u0_U22263  ( .A(1'b0), .ZN(_u0_ch2_am0[15] ) );
INV_X4 _u0_U22261  ( .A(1'b0), .ZN(_u0_ch2_am0[14] ) );
INV_X4 _u0_U22259  ( .A(1'b0), .ZN(_u0_ch2_am0[13] ) );
INV_X4 _u0_U22257  ( .A(1'b0), .ZN(_u0_ch2_am0[12] ) );
INV_X4 _u0_U22255  ( .A(1'b0), .ZN(_u0_ch2_am0[11] ) );
INV_X4 _u0_U22253  ( .A(1'b0), .ZN(_u0_ch2_am0[10] ) );
INV_X4 _u0_U22251  ( .A(1'b0), .ZN(_u0_ch2_am0[9] ) );
INV_X4 _u0_U22249  ( .A(1'b0), .ZN(_u0_ch2_am0[8] ) );
INV_X4 _u0_U22247  ( .A(1'b0), .ZN(_u0_ch2_am0[7] ) );
INV_X4 _u0_U22245  ( .A(1'b0), .ZN(_u0_ch2_am0[6] ) );
INV_X4 _u0_U22243  ( .A(1'b0), .ZN(_u0_ch2_am0[5] ) );
INV_X4 _u0_U22241  ( .A(1'b0), .ZN(_u0_ch2_am0[4] ) );
INV_X4 _u0_U22239  ( .A(1'b1), .ZN(_u0_ch2_am0[3] ) );
INV_X4 _u0_U22237  ( .A(1'b1), .ZN(_u0_ch2_am0[2] ) );
INV_X4 _u0_U22235  ( .A(1'b1), .ZN(_u0_ch2_am0[1] ) );
INV_X4 _u0_U22233  ( .A(1'b1), .ZN(_u0_ch2_am0[0] ) );
INV_X4 _u0_U22231  ( .A(1'b0), .ZN(_u0_ch2_am1[31] ) );
INV_X4 _u0_U22229  ( .A(1'b0), .ZN(_u0_ch2_am1[30] ) );
INV_X4 _u0_U22227  ( .A(1'b0), .ZN(_u0_ch2_am1[29] ) );
INV_X4 _u0_U22225  ( .A(1'b0), .ZN(_u0_ch2_am1[28] ) );
INV_X4 _u0_U22223  ( .A(1'b0), .ZN(_u0_ch2_am1[27] ) );
INV_X4 _u0_U22221  ( .A(1'b0), .ZN(_u0_ch2_am1[26] ) );
INV_X4 _u0_U22219  ( .A(1'b0), .ZN(_u0_ch2_am1[25] ) );
INV_X4 _u0_U22217  ( .A(1'b0), .ZN(_u0_ch2_am1[24] ) );
INV_X4 _u0_U22215  ( .A(1'b0), .ZN(_u0_ch2_am1[23] ) );
INV_X4 _u0_U22213  ( .A(1'b0), .ZN(_u0_ch2_am1[22] ) );
INV_X4 _u0_U22211  ( .A(1'b0), .ZN(_u0_ch2_am1[21] ) );
INV_X4 _u0_U22209  ( .A(1'b0), .ZN(_u0_ch2_am1[20] ) );
INV_X4 _u0_U22207  ( .A(1'b0), .ZN(_u0_ch2_am1[19] ) );
INV_X4 _u0_U22205  ( .A(1'b0), .ZN(_u0_ch2_am1[18] ) );
INV_X4 _u0_U22203  ( .A(1'b0), .ZN(_u0_ch2_am1[17] ) );
INV_X4 _u0_U22201  ( .A(1'b0), .ZN(_u0_ch2_am1[16] ) );
INV_X4 _u0_U22199  ( .A(1'b0), .ZN(_u0_ch2_am1[15] ) );
INV_X4 _u0_U22197  ( .A(1'b0), .ZN(_u0_ch2_am1[14] ) );
INV_X4 _u0_U22195  ( .A(1'b0), .ZN(_u0_ch2_am1[13] ) );
INV_X4 _u0_U22193  ( .A(1'b0), .ZN(_u0_ch2_am1[12] ) );
INV_X4 _u0_U22191  ( .A(1'b0), .ZN(_u0_ch2_am1[11] ) );
INV_X4 _u0_U22189  ( .A(1'b0), .ZN(_u0_ch2_am1[10] ) );
INV_X4 _u0_U22187  ( .A(1'b0), .ZN(_u0_ch2_am1[9] ) );
INV_X4 _u0_U22185  ( .A(1'b0), .ZN(_u0_ch2_am1[8] ) );
INV_X4 _u0_U22183  ( .A(1'b0), .ZN(_u0_ch2_am1[7] ) );
INV_X4 _u0_U22181  ( .A(1'b0), .ZN(_u0_ch2_am1[6] ) );
INV_X4 _u0_U22179  ( .A(1'b0), .ZN(_u0_ch2_am1[5] ) );
INV_X4 _u0_U22177  ( .A(1'b0), .ZN(_u0_ch2_am1[4] ) );
INV_X4 _u0_U22175  ( .A(1'b1), .ZN(_u0_ch2_am1[3] ) );
INV_X4 _u0_U22173  ( .A(1'b1), .ZN(_u0_ch2_am1[2] ) );
INV_X4 _u0_U22171  ( .A(1'b1), .ZN(_u0_ch2_am1[1] ) );
INV_X4 _u0_U22169  ( .A(1'b1), .ZN(_u0_ch2_am1[0] ) );
INV_X4 _u0_U22167  ( .A(1'b1), .ZN(_u0_pointer3[31] ) );
INV_X4 _u0_U22165  ( .A(1'b1), .ZN(_u0_pointer3[30] ) );
INV_X4 _u0_U22163  ( .A(1'b1), .ZN(_u0_pointer3[29] ) );
INV_X4 _u0_U22161  ( .A(1'b1), .ZN(_u0_pointer3[28] ) );
INV_X4 _u0_U22159  ( .A(1'b1), .ZN(_u0_pointer3[27] ) );
INV_X4 _u0_U22157  ( .A(1'b1), .ZN(_u0_pointer3[26] ) );
INV_X4 _u0_U22155  ( .A(1'b1), .ZN(_u0_pointer3[25] ) );
INV_X4 _u0_U22153  ( .A(1'b1), .ZN(_u0_pointer3[24] ) );
INV_X4 _u0_U22151  ( .A(1'b1), .ZN(_u0_pointer3[23] ) );
INV_X4 _u0_U22149  ( .A(1'b1), .ZN(_u0_pointer3[22] ) );
INV_X4 _u0_U22147  ( .A(1'b1), .ZN(_u0_pointer3[21] ) );
INV_X4 _u0_U22145  ( .A(1'b1), .ZN(_u0_pointer3[20] ) );
INV_X4 _u0_U22143  ( .A(1'b1), .ZN(_u0_pointer3[19] ) );
INV_X4 _u0_U22141  ( .A(1'b1), .ZN(_u0_pointer3[18] ) );
INV_X4 _u0_U22139  ( .A(1'b1), .ZN(_u0_pointer3[17] ) );
INV_X4 _u0_U22137  ( .A(1'b1), .ZN(_u0_pointer3[16] ) );
INV_X4 _u0_U22135  ( .A(1'b1), .ZN(_u0_pointer3[15] ) );
INV_X4 _u0_U22133  ( .A(1'b1), .ZN(_u0_pointer3[14] ) );
INV_X4 _u0_U22131  ( .A(1'b1), .ZN(_u0_pointer3[13] ) );
INV_X4 _u0_U22129  ( .A(1'b1), .ZN(_u0_pointer3[12] ) );
INV_X4 _u0_U22127  ( .A(1'b1), .ZN(_u0_pointer3[11] ) );
INV_X4 _u0_U22125  ( .A(1'b1), .ZN(_u0_pointer3[10] ) );
INV_X4 _u0_U22123  ( .A(1'b1), .ZN(_u0_pointer3[9] ) );
INV_X4 _u0_U22121  ( .A(1'b1), .ZN(_u0_pointer3[8] ) );
INV_X4 _u0_U22119  ( .A(1'b1), .ZN(_u0_pointer3[7] ) );
INV_X4 _u0_U22117  ( .A(1'b1), .ZN(_u0_pointer3[6] ) );
INV_X4 _u0_U22115  ( .A(1'b1), .ZN(_u0_pointer3[5] ) );
INV_X4 _u0_U22113  ( .A(1'b1), .ZN(_u0_pointer3[4] ) );
INV_X4 _u0_U22111  ( .A(1'b1), .ZN(_u0_pointer3[3] ) );
INV_X4 _u0_U22109  ( .A(1'b1), .ZN(_u0_pointer3[2] ) );
INV_X4 _u0_U22107  ( .A(1'b1), .ZN(_u0_pointer3[1] ) );
INV_X4 _u0_U22105  ( .A(1'b1), .ZN(_u0_pointer3[0] ) );
INV_X4 _u0_U22103  ( .A(1'b1), .ZN(_u0_pointer3_s[31] ) );
INV_X4 _u0_U22101  ( .A(1'b1), .ZN(_u0_pointer3_s[30] ) );
INV_X4 _u0_U22099  ( .A(1'b1), .ZN(_u0_pointer3_s[29] ) );
INV_X4 _u0_U22097  ( .A(1'b1), .ZN(_u0_pointer3_s[28] ) );
INV_X4 _u0_U22095  ( .A(1'b1), .ZN(_u0_pointer3_s[27] ) );
INV_X4 _u0_U22093  ( .A(1'b1), .ZN(_u0_pointer3_s[26] ) );
INV_X4 _u0_U22091  ( .A(1'b1), .ZN(_u0_pointer3_s[25] ) );
INV_X4 _u0_U22089  ( .A(1'b1), .ZN(_u0_pointer3_s[24] ) );
INV_X4 _u0_U22087  ( .A(1'b1), .ZN(_u0_pointer3_s[23] ) );
INV_X4 _u0_U22085  ( .A(1'b1), .ZN(_u0_pointer3_s[22] ) );
INV_X4 _u0_U22083  ( .A(1'b1), .ZN(_u0_pointer3_s[21] ) );
INV_X4 _u0_U22081  ( .A(1'b1), .ZN(_u0_pointer3_s[20] ) );
INV_X4 _u0_U22079  ( .A(1'b1), .ZN(_u0_pointer3_s[19] ) );
INV_X4 _u0_U22077  ( .A(1'b1), .ZN(_u0_pointer3_s[18] ) );
INV_X4 _u0_U22075  ( .A(1'b1), .ZN(_u0_pointer3_s[17] ) );
INV_X4 _u0_U22073  ( .A(1'b1), .ZN(_u0_pointer3_s[16] ) );
INV_X4 _u0_U22071  ( .A(1'b1), .ZN(_u0_pointer3_s[15] ) );
INV_X4 _u0_U22069  ( .A(1'b1), .ZN(_u0_pointer3_s[14] ) );
INV_X4 _u0_U22067  ( .A(1'b1), .ZN(_u0_pointer3_s[13] ) );
INV_X4 _u0_U22065  ( .A(1'b1), .ZN(_u0_pointer3_s[12] ) );
INV_X4 _u0_U22063  ( .A(1'b1), .ZN(_u0_pointer3_s[11] ) );
INV_X4 _u0_U22061  ( .A(1'b1), .ZN(_u0_pointer3_s[10] ) );
INV_X4 _u0_U22059  ( .A(1'b1), .ZN(_u0_pointer3_s[9] ) );
INV_X4 _u0_U22057  ( .A(1'b1), .ZN(_u0_pointer3_s[8] ) );
INV_X4 _u0_U22055  ( .A(1'b1), .ZN(_u0_pointer3_s[7] ) );
INV_X4 _u0_U22053  ( .A(1'b1), .ZN(_u0_pointer3_s[6] ) );
INV_X4 _u0_U22051  ( .A(1'b1), .ZN(_u0_pointer3_s[5] ) );
INV_X4 _u0_U22049  ( .A(1'b1), .ZN(_u0_pointer3_s[4] ) );
INV_X4 _u0_U22047  ( .A(1'b1), .ZN(_u0_pointer3_s[3] ) );
INV_X4 _u0_U22045  ( .A(1'b1), .ZN(_u0_pointer3_s[2] ) );
INV_X4 _u0_U22043  ( .A(1'b1), .ZN(_u0_pointer3_s[1] ) );
INV_X4 _u0_U22041  ( .A(1'b1), .ZN(_u0_pointer3_s[0] ) );
INV_X4 _u0_U22039  ( .A(1'b1), .ZN(_u0_ch3_csr[31] ) );
INV_X4 _u0_U22037  ( .A(1'b1), .ZN(_u0_ch3_csr[30] ) );
INV_X4 _u0_U22035  ( .A(1'b1), .ZN(_u0_ch3_csr[29] ) );
INV_X4 _u0_U22033  ( .A(1'b1), .ZN(_u0_ch3_csr[28] ) );
INV_X4 _u0_U22031  ( .A(1'b1), .ZN(_u0_ch3_csr[27] ) );
INV_X4 _u0_U22029  ( .A(1'b1), .ZN(_u0_ch3_csr[26] ) );
INV_X4 _u0_U22027  ( .A(1'b1), .ZN(_u0_ch3_csr[25] ) );
INV_X4 _u0_U22025  ( .A(1'b1), .ZN(_u0_ch3_csr[24] ) );
INV_X4 _u0_U22023  ( .A(1'b1), .ZN(_u0_ch3_csr[23] ) );
INV_X4 _u0_U22021  ( .A(1'b1), .ZN(_u0_ch3_csr[22] ) );
INV_X4 _u0_U22019  ( .A(1'b1), .ZN(_u0_ch3_csr[21] ) );
INV_X4 _u0_U22017  ( .A(1'b1), .ZN(_u0_ch3_csr[20] ) );
INV_X4 _u0_U22015  ( .A(1'b1), .ZN(_u0_ch3_csr[19] ) );
INV_X4 _u0_U22013  ( .A(1'b1), .ZN(_u0_ch3_csr[18] ) );
INV_X4 _u0_U22011  ( .A(1'b1), .ZN(_u0_ch3_csr[17] ) );
INV_X4 _u0_U22009  ( .A(1'b1), .ZN(_u0_ch3_csr[16] ) );
INV_X4 _u0_U22007  ( .A(1'b1), .ZN(_u0_ch3_csr[15] ) );
INV_X4 _u0_U22005  ( .A(1'b1), .ZN(_u0_ch3_csr[14] ) );
INV_X4 _u0_U22003  ( .A(1'b1), .ZN(_u0_ch3_csr[13] ) );
INV_X4 _u0_U22001  ( .A(1'b1), .ZN(_u0_ch3_csr[12] ) );
INV_X4 _u0_U21999  ( .A(1'b1), .ZN(_u0_ch3_csr[11] ) );
INV_X4 _u0_U21997  ( .A(1'b1), .ZN(_u0_ch3_csr[10] ) );
INV_X4 _u0_U21995  ( .A(1'b1), .ZN(_u0_ch3_csr[9] ) );
INV_X4 _u0_U21993  ( .A(1'b1), .ZN(_u0_ch3_csr[8] ) );
INV_X4 _u0_U21991  ( .A(1'b1), .ZN(_u0_ch3_csr[7] ) );
INV_X4 _u0_U21989  ( .A(1'b1), .ZN(_u0_ch3_csr[6] ) );
INV_X4 _u0_U21987  ( .A(1'b1), .ZN(_u0_ch3_csr[5] ) );
INV_X4 _u0_U21985  ( .A(1'b1), .ZN(_u0_ch3_csr[4] ) );
INV_X4 _u0_U21983  ( .A(1'b1), .ZN(_u0_ch3_csr[3] ) );
INV_X4 _u0_U21981  ( .A(1'b1), .ZN(_u0_ch3_csr[2] ) );
INV_X4 _u0_U21979  ( .A(1'b1), .ZN(_u0_ch3_csr[1] ) );
INV_X4 _u0_U21977  ( .A(1'b1), .ZN(_u0_ch3_csr[0] ) );
INV_X4 _u0_U21975  ( .A(1'b1), .ZN(_u0_ch3_txsz[31] ) );
INV_X4 _u0_U21973  ( .A(1'b1), .ZN(_u0_ch3_txsz[30] ) );
INV_X4 _u0_U21971  ( .A(1'b1), .ZN(_u0_ch3_txsz[29] ) );
INV_X4 _u0_U21969  ( .A(1'b1), .ZN(_u0_ch3_txsz[28] ) );
INV_X4 _u0_U21967  ( .A(1'b1), .ZN(_u0_ch3_txsz[27] ) );
INV_X4 _u0_U21965  ( .A(1'b1), .ZN(_u0_ch3_txsz[26] ) );
INV_X4 _u0_U21963  ( .A(1'b1), .ZN(_u0_ch3_txsz[25] ) );
INV_X4 _u0_U21961  ( .A(1'b1), .ZN(_u0_ch3_txsz[24] ) );
INV_X4 _u0_U21959  ( .A(1'b1), .ZN(_u0_ch3_txsz[23] ) );
INV_X4 _u0_U21957  ( .A(1'b1), .ZN(_u0_ch3_txsz[22] ) );
INV_X4 _u0_U21955  ( .A(1'b1), .ZN(_u0_ch3_txsz[21] ) );
INV_X4 _u0_U21953  ( .A(1'b1), .ZN(_u0_ch3_txsz[20] ) );
INV_X4 _u0_U21951  ( .A(1'b1), .ZN(_u0_ch3_txsz[19] ) );
INV_X4 _u0_U21949  ( .A(1'b1), .ZN(_u0_ch3_txsz[18] ) );
INV_X4 _u0_U21947  ( .A(1'b1), .ZN(_u0_ch3_txsz[17] ) );
INV_X4 _u0_U21945  ( .A(1'b1), .ZN(_u0_ch3_txsz[16] ) );
INV_X4 _u0_U21943  ( .A(1'b1), .ZN(_u0_ch3_txsz[15] ) );
INV_X4 _u0_U21941  ( .A(1'b1), .ZN(_u0_ch3_txsz[14] ) );
INV_X4 _u0_U21939  ( .A(1'b1), .ZN(_u0_ch3_txsz[13] ) );
INV_X4 _u0_U21937  ( .A(1'b1), .ZN(_u0_ch3_txsz[12] ) );
INV_X4 _u0_U21935  ( .A(1'b1), .ZN(_u0_ch3_txsz[11] ) );
INV_X4 _u0_U21933  ( .A(1'b1), .ZN(_u0_ch3_txsz[10] ) );
INV_X4 _u0_U21931  ( .A(1'b1), .ZN(_u0_ch3_txsz[9] ) );
INV_X4 _u0_U21929  ( .A(1'b1), .ZN(_u0_ch3_txsz[8] ) );
INV_X4 _u0_U21927  ( .A(1'b1), .ZN(_u0_ch3_txsz[7] ) );
INV_X4 _u0_U21925  ( .A(1'b1), .ZN(_u0_ch3_txsz[6] ) );
INV_X4 _u0_U21923  ( .A(1'b1), .ZN(_u0_ch3_txsz[5] ) );
INV_X4 _u0_U21921  ( .A(1'b1), .ZN(_u0_ch3_txsz[4] ) );
INV_X4 _u0_U21919  ( .A(1'b1), .ZN(_u0_ch3_txsz[3] ) );
INV_X4 _u0_U21917  ( .A(1'b1), .ZN(_u0_ch3_txsz[2] ) );
INV_X4 _u0_U21915  ( .A(1'b1), .ZN(_u0_ch3_txsz[1] ) );
INV_X4 _u0_U21913  ( .A(1'b1), .ZN(_u0_ch3_txsz[0] ) );
INV_X4 _u0_U21911  ( .A(1'b1), .ZN(_u0_ch3_adr0[31] ) );
INV_X4 _u0_U21909  ( .A(1'b1), .ZN(_u0_ch3_adr0[30] ) );
INV_X4 _u0_U21907  ( .A(1'b1), .ZN(_u0_ch3_adr0[29] ) );
INV_X4 _u0_U21905  ( .A(1'b1), .ZN(_u0_ch3_adr0[28] ) );
INV_X4 _u0_U21903  ( .A(1'b1), .ZN(_u0_ch3_adr0[27] ) );
INV_X4 _u0_U21901  ( .A(1'b1), .ZN(_u0_ch3_adr0[26] ) );
INV_X4 _u0_U21899  ( .A(1'b1), .ZN(_u0_ch3_adr0[25] ) );
INV_X4 _u0_U21897  ( .A(1'b1), .ZN(_u0_ch3_adr0[24] ) );
INV_X4 _u0_U21895  ( .A(1'b1), .ZN(_u0_ch3_adr0[23] ) );
INV_X4 _u0_U21893  ( .A(1'b1), .ZN(_u0_ch3_adr0[22] ) );
INV_X4 _u0_U21891  ( .A(1'b1), .ZN(_u0_ch3_adr0[21] ) );
INV_X4 _u0_U21889  ( .A(1'b1), .ZN(_u0_ch3_adr0[20] ) );
INV_X4 _u0_U21887  ( .A(1'b1), .ZN(_u0_ch3_adr0[19] ) );
INV_X4 _u0_U21885  ( .A(1'b1), .ZN(_u0_ch3_adr0[18] ) );
INV_X4 _u0_U21883  ( .A(1'b1), .ZN(_u0_ch3_adr0[17] ) );
INV_X4 _u0_U21881  ( .A(1'b1), .ZN(_u0_ch3_adr0[16] ) );
INV_X4 _u0_U21879  ( .A(1'b1), .ZN(_u0_ch3_adr0[15] ) );
INV_X4 _u0_U21877  ( .A(1'b1), .ZN(_u0_ch3_adr0[14] ) );
INV_X4 _u0_U21875  ( .A(1'b1), .ZN(_u0_ch3_adr0[13] ) );
INV_X4 _u0_U21873  ( .A(1'b1), .ZN(_u0_ch3_adr0[12] ) );
INV_X4 _u0_U21871  ( .A(1'b1), .ZN(_u0_ch3_adr0[11] ) );
INV_X4 _u0_U21869  ( .A(1'b1), .ZN(_u0_ch3_adr0[10] ) );
INV_X4 _u0_U21867  ( .A(1'b1), .ZN(_u0_ch3_adr0[9] ) );
INV_X4 _u0_U21865  ( .A(1'b1), .ZN(_u0_ch3_adr0[8] ) );
INV_X4 _u0_U21863  ( .A(1'b1), .ZN(_u0_ch3_adr0[7] ) );
INV_X4 _u0_U21861  ( .A(1'b1), .ZN(_u0_ch3_adr0[6] ) );
INV_X4 _u0_U21859  ( .A(1'b1), .ZN(_u0_ch3_adr0[5] ) );
INV_X4 _u0_U21857  ( .A(1'b1), .ZN(_u0_ch3_adr0[4] ) );
INV_X4 _u0_U21855  ( .A(1'b1), .ZN(_u0_ch3_adr0[3] ) );
INV_X4 _u0_U21853  ( .A(1'b1), .ZN(_u0_ch3_adr0[2] ) );
INV_X4 _u0_U21851  ( .A(1'b1), .ZN(_u0_ch3_adr0[1] ) );
INV_X4 _u0_U21849  ( .A(1'b1), .ZN(_u0_ch3_adr0[0] ) );
INV_X4 _u0_U21847  ( .A(1'b1), .ZN(_u0_ch3_adr1[31] ) );
INV_X4 _u0_U21845  ( .A(1'b1), .ZN(_u0_ch3_adr1[30] ) );
INV_X4 _u0_U21843  ( .A(1'b1), .ZN(_u0_ch3_adr1[29] ) );
INV_X4 _u0_U21841  ( .A(1'b1), .ZN(_u0_ch3_adr1[28] ) );
INV_X4 _u0_U21839  ( .A(1'b1), .ZN(_u0_ch3_adr1[27] ) );
INV_X4 _u0_U21837  ( .A(1'b1), .ZN(_u0_ch3_adr1[26] ) );
INV_X4 _u0_U21835  ( .A(1'b1), .ZN(_u0_ch3_adr1[25] ) );
INV_X4 _u0_U21833  ( .A(1'b1), .ZN(_u0_ch3_adr1[24] ) );
INV_X4 _u0_U21831  ( .A(1'b1), .ZN(_u0_ch3_adr1[23] ) );
INV_X4 _u0_U21829  ( .A(1'b1), .ZN(_u0_ch3_adr1[22] ) );
INV_X4 _u0_U21827  ( .A(1'b1), .ZN(_u0_ch3_adr1[21] ) );
INV_X4 _u0_U21825  ( .A(1'b1), .ZN(_u0_ch3_adr1[20] ) );
INV_X4 _u0_U21823  ( .A(1'b1), .ZN(_u0_ch3_adr1[19] ) );
INV_X4 _u0_U21821  ( .A(1'b1), .ZN(_u0_ch3_adr1[18] ) );
INV_X4 _u0_U21819  ( .A(1'b1), .ZN(_u0_ch3_adr1[17] ) );
INV_X4 _u0_U21817  ( .A(1'b1), .ZN(_u0_ch3_adr1[16] ) );
INV_X4 _u0_U21815  ( .A(1'b1), .ZN(_u0_ch3_adr1[15] ) );
INV_X4 _u0_U21813  ( .A(1'b1), .ZN(_u0_ch3_adr1[14] ) );
INV_X4 _u0_U21811  ( .A(1'b1), .ZN(_u0_ch3_adr1[13] ) );
INV_X4 _u0_U21809  ( .A(1'b1), .ZN(_u0_ch3_adr1[12] ) );
INV_X4 _u0_U21807  ( .A(1'b1), .ZN(_u0_ch3_adr1[11] ) );
INV_X4 _u0_U21805  ( .A(1'b1), .ZN(_u0_ch3_adr1[10] ) );
INV_X4 _u0_U21803  ( .A(1'b1), .ZN(_u0_ch3_adr1[9] ) );
INV_X4 _u0_U21801  ( .A(1'b1), .ZN(_u0_ch3_adr1[8] ) );
INV_X4 _u0_U21799  ( .A(1'b1), .ZN(_u0_ch3_adr1[7] ) );
INV_X4 _u0_U21797  ( .A(1'b1), .ZN(_u0_ch3_adr1[6] ) );
INV_X4 _u0_U21795  ( .A(1'b1), .ZN(_u0_ch3_adr1[5] ) );
INV_X4 _u0_U21793  ( .A(1'b1), .ZN(_u0_ch3_adr1[4] ) );
INV_X4 _u0_U21791  ( .A(1'b1), .ZN(_u0_ch3_adr1[3] ) );
INV_X4 _u0_U21789  ( .A(1'b1), .ZN(_u0_ch3_adr1[2] ) );
INV_X4 _u0_U21787  ( .A(1'b1), .ZN(_u0_ch3_adr1[1] ) );
INV_X4 _u0_U21785  ( .A(1'b1), .ZN(_u0_ch3_adr1[0] ) );
INV_X4 _u0_U21783  ( .A(1'b0), .ZN(_u0_ch3_am0[31] ) );
INV_X4 _u0_U21781  ( .A(1'b0), .ZN(_u0_ch3_am0[30] ) );
INV_X4 _u0_U21779  ( .A(1'b0), .ZN(_u0_ch3_am0[29] ) );
INV_X4 _u0_U21777  ( .A(1'b0), .ZN(_u0_ch3_am0[28] ) );
INV_X4 _u0_U21775  ( .A(1'b0), .ZN(_u0_ch3_am0[27] ) );
INV_X4 _u0_U21773  ( .A(1'b0), .ZN(_u0_ch3_am0[26] ) );
INV_X4 _u0_U21771  ( .A(1'b0), .ZN(_u0_ch3_am0[25] ) );
INV_X4 _u0_U21769  ( .A(1'b0), .ZN(_u0_ch3_am0[24] ) );
INV_X4 _u0_U21767  ( .A(1'b0), .ZN(_u0_ch3_am0[23] ) );
INV_X4 _u0_U21765  ( .A(1'b0), .ZN(_u0_ch3_am0[22] ) );
INV_X4 _u0_U21763  ( .A(1'b0), .ZN(_u0_ch3_am0[21] ) );
INV_X4 _u0_U21761  ( .A(1'b0), .ZN(_u0_ch3_am0[20] ) );
INV_X4 _u0_U21759  ( .A(1'b0), .ZN(_u0_ch3_am0[19] ) );
INV_X4 _u0_U21757  ( .A(1'b0), .ZN(_u0_ch3_am0[18] ) );
INV_X4 _u0_U21755  ( .A(1'b0), .ZN(_u0_ch3_am0[17] ) );
INV_X4 _u0_U21753  ( .A(1'b0), .ZN(_u0_ch3_am0[16] ) );
INV_X4 _u0_U21751  ( .A(1'b0), .ZN(_u0_ch3_am0[15] ) );
INV_X4 _u0_U21749  ( .A(1'b0), .ZN(_u0_ch3_am0[14] ) );
INV_X4 _u0_U21747  ( .A(1'b0), .ZN(_u0_ch3_am0[13] ) );
INV_X4 _u0_U21745  ( .A(1'b0), .ZN(_u0_ch3_am0[12] ) );
INV_X4 _u0_U21743  ( .A(1'b0), .ZN(_u0_ch3_am0[11] ) );
INV_X4 _u0_U21741  ( .A(1'b0), .ZN(_u0_ch3_am0[10] ) );
INV_X4 _u0_U21739  ( .A(1'b0), .ZN(_u0_ch3_am0[9] ) );
INV_X4 _u0_U21737  ( .A(1'b0), .ZN(_u0_ch3_am0[8] ) );
INV_X4 _u0_U21735  ( .A(1'b0), .ZN(_u0_ch3_am0[7] ) );
INV_X4 _u0_U21733  ( .A(1'b0), .ZN(_u0_ch3_am0[6] ) );
INV_X4 _u0_U21731  ( .A(1'b0), .ZN(_u0_ch3_am0[5] ) );
INV_X4 _u0_U21729  ( .A(1'b0), .ZN(_u0_ch3_am0[4] ) );
INV_X4 _u0_U21727  ( .A(1'b1), .ZN(_u0_ch3_am0[3] ) );
INV_X4 _u0_U21725  ( .A(1'b1), .ZN(_u0_ch3_am0[2] ) );
INV_X4 _u0_U21723  ( .A(1'b1), .ZN(_u0_ch3_am0[1] ) );
INV_X4 _u0_U21721  ( .A(1'b1), .ZN(_u0_ch3_am0[0] ) );
INV_X4 _u0_U21719  ( .A(1'b0), .ZN(_u0_ch3_am1[31] ) );
INV_X4 _u0_U21717  ( .A(1'b0), .ZN(_u0_ch3_am1[30] ) );
INV_X4 _u0_U21715  ( .A(1'b0), .ZN(_u0_ch3_am1[29] ) );
INV_X4 _u0_U21713  ( .A(1'b0), .ZN(_u0_ch3_am1[28] ) );
INV_X4 _u0_U21711  ( .A(1'b0), .ZN(_u0_ch3_am1[27] ) );
INV_X4 _u0_U21709  ( .A(1'b0), .ZN(_u0_ch3_am1[26] ) );
INV_X4 _u0_U21707  ( .A(1'b0), .ZN(_u0_ch3_am1[25] ) );
INV_X4 _u0_U21705  ( .A(1'b0), .ZN(_u0_ch3_am1[24] ) );
INV_X4 _u0_U21703  ( .A(1'b0), .ZN(_u0_ch3_am1[23] ) );
INV_X4 _u0_U21701  ( .A(1'b0), .ZN(_u0_ch3_am1[22] ) );
INV_X4 _u0_U21699  ( .A(1'b0), .ZN(_u0_ch3_am1[21] ) );
INV_X4 _u0_U21697  ( .A(1'b0), .ZN(_u0_ch3_am1[20] ) );
INV_X4 _u0_U21695  ( .A(1'b0), .ZN(_u0_ch3_am1[19] ) );
INV_X4 _u0_U21693  ( .A(1'b0), .ZN(_u0_ch3_am1[18] ) );
INV_X4 _u0_U21691  ( .A(1'b0), .ZN(_u0_ch3_am1[17] ) );
INV_X4 _u0_U21689  ( .A(1'b0), .ZN(_u0_ch3_am1[16] ) );
INV_X4 _u0_U21687  ( .A(1'b0), .ZN(_u0_ch3_am1[15] ) );
INV_X4 _u0_U21685  ( .A(1'b0), .ZN(_u0_ch3_am1[14] ) );
INV_X4 _u0_U21683  ( .A(1'b0), .ZN(_u0_ch3_am1[13] ) );
INV_X4 _u0_U21681  ( .A(1'b0), .ZN(_u0_ch3_am1[12] ) );
INV_X4 _u0_U21679  ( .A(1'b0), .ZN(_u0_ch3_am1[11] ) );
INV_X4 _u0_U21677  ( .A(1'b0), .ZN(_u0_ch3_am1[10] ) );
INV_X4 _u0_U21675  ( .A(1'b0), .ZN(_u0_ch3_am1[9] ) );
INV_X4 _u0_U21673  ( .A(1'b0), .ZN(_u0_ch3_am1[8] ) );
INV_X4 _u0_U21671  ( .A(1'b0), .ZN(_u0_ch3_am1[7] ) );
INV_X4 _u0_U21669  ( .A(1'b0), .ZN(_u0_ch3_am1[6] ) );
INV_X4 _u0_U21667  ( .A(1'b0), .ZN(_u0_ch3_am1[5] ) );
INV_X4 _u0_U21665  ( .A(1'b0), .ZN(_u0_ch3_am1[4] ) );
INV_X4 _u0_U21663  ( .A(1'b1), .ZN(_u0_ch3_am1[3] ) );
INV_X4 _u0_U21661  ( .A(1'b1), .ZN(_u0_ch3_am1[2] ) );
INV_X4 _u0_U21659  ( .A(1'b1), .ZN(_u0_ch3_am1[1] ) );
INV_X4 _u0_U21657  ( .A(1'b1), .ZN(_u0_ch3_am1[0] ) );
INV_X4 _u0_U21655  ( .A(1'b1), .ZN(_u0_pointer4[31] ) );
INV_X4 _u0_U21653  ( .A(1'b1), .ZN(_u0_pointer4[30] ) );
INV_X4 _u0_U21651  ( .A(1'b1), .ZN(_u0_pointer4[29] ) );
INV_X4 _u0_U21649  ( .A(1'b1), .ZN(_u0_pointer4[28] ) );
INV_X4 _u0_U21647  ( .A(1'b1), .ZN(_u0_pointer4[27] ) );
INV_X4 _u0_U21645  ( .A(1'b1), .ZN(_u0_pointer4[26] ) );
INV_X4 _u0_U21643  ( .A(1'b1), .ZN(_u0_pointer4[25] ) );
INV_X4 _u0_U21641  ( .A(1'b1), .ZN(_u0_pointer4[24] ) );
INV_X4 _u0_U21639  ( .A(1'b1), .ZN(_u0_pointer4[23] ) );
INV_X4 _u0_U21637  ( .A(1'b1), .ZN(_u0_pointer4[22] ) );
INV_X4 _u0_U21635  ( .A(1'b1), .ZN(_u0_pointer4[21] ) );
INV_X4 _u0_U21633  ( .A(1'b1), .ZN(_u0_pointer4[20] ) );
INV_X4 _u0_U21631  ( .A(1'b1), .ZN(_u0_pointer4[19] ) );
INV_X4 _u0_U21629  ( .A(1'b1), .ZN(_u0_pointer4[18] ) );
INV_X4 _u0_U21627  ( .A(1'b1), .ZN(_u0_pointer4[17] ) );
INV_X4 _u0_U21625  ( .A(1'b1), .ZN(_u0_pointer4[16] ) );
INV_X4 _u0_U21623  ( .A(1'b1), .ZN(_u0_pointer4[15] ) );
INV_X4 _u0_U21621  ( .A(1'b1), .ZN(_u0_pointer4[14] ) );
INV_X4 _u0_U21619  ( .A(1'b1), .ZN(_u0_pointer4[13] ) );
INV_X4 _u0_U21617  ( .A(1'b1), .ZN(_u0_pointer4[12] ) );
INV_X4 _u0_U21615  ( .A(1'b1), .ZN(_u0_pointer4[11] ) );
INV_X4 _u0_U21613  ( .A(1'b1), .ZN(_u0_pointer4[10] ) );
INV_X4 _u0_U21611  ( .A(1'b1), .ZN(_u0_pointer4[9] ) );
INV_X4 _u0_U21609  ( .A(1'b1), .ZN(_u0_pointer4[8] ) );
INV_X4 _u0_U21607  ( .A(1'b1), .ZN(_u0_pointer4[7] ) );
INV_X4 _u0_U21605  ( .A(1'b1), .ZN(_u0_pointer4[6] ) );
INV_X4 _u0_U21603  ( .A(1'b1), .ZN(_u0_pointer4[5] ) );
INV_X4 _u0_U21601  ( .A(1'b1), .ZN(_u0_pointer4[4] ) );
INV_X4 _u0_U21599  ( .A(1'b1), .ZN(_u0_pointer4[3] ) );
INV_X4 _u0_U21597  ( .A(1'b1), .ZN(_u0_pointer4[2] ) );
INV_X4 _u0_U21595  ( .A(1'b1), .ZN(_u0_pointer4[1] ) );
INV_X4 _u0_U21593  ( .A(1'b1), .ZN(_u0_pointer4[0] ) );
INV_X4 _u0_U21591  ( .A(1'b1), .ZN(_u0_pointer4_s[31] ) );
INV_X4 _u0_U21589  ( .A(1'b1), .ZN(_u0_pointer4_s[30] ) );
INV_X4 _u0_U21587  ( .A(1'b1), .ZN(_u0_pointer4_s[29] ) );
INV_X4 _u0_U21585  ( .A(1'b1), .ZN(_u0_pointer4_s[28] ) );
INV_X4 _u0_U21583  ( .A(1'b1), .ZN(_u0_pointer4_s[27] ) );
INV_X4 _u0_U21581  ( .A(1'b1), .ZN(_u0_pointer4_s[26] ) );
INV_X4 _u0_U21579  ( .A(1'b1), .ZN(_u0_pointer4_s[25] ) );
INV_X4 _u0_U21577  ( .A(1'b1), .ZN(_u0_pointer4_s[24] ) );
INV_X4 _u0_U21575  ( .A(1'b1), .ZN(_u0_pointer4_s[23] ) );
INV_X4 _u0_U21573  ( .A(1'b1), .ZN(_u0_pointer4_s[22] ) );
INV_X4 _u0_U21571  ( .A(1'b1), .ZN(_u0_pointer4_s[21] ) );
INV_X4 _u0_U21569  ( .A(1'b1), .ZN(_u0_pointer4_s[20] ) );
INV_X4 _u0_U21567  ( .A(1'b1), .ZN(_u0_pointer4_s[19] ) );
INV_X4 _u0_U21565  ( .A(1'b1), .ZN(_u0_pointer4_s[18] ) );
INV_X4 _u0_U21563  ( .A(1'b1), .ZN(_u0_pointer4_s[17] ) );
INV_X4 _u0_U21561  ( .A(1'b1), .ZN(_u0_pointer4_s[16] ) );
INV_X4 _u0_U21559  ( .A(1'b1), .ZN(_u0_pointer4_s[15] ) );
INV_X4 _u0_U21557  ( .A(1'b1), .ZN(_u0_pointer4_s[14] ) );
INV_X4 _u0_U21555  ( .A(1'b1), .ZN(_u0_pointer4_s[13] ) );
INV_X4 _u0_U21553  ( .A(1'b1), .ZN(_u0_pointer4_s[12] ) );
INV_X4 _u0_U21551  ( .A(1'b1), .ZN(_u0_pointer4_s[11] ) );
INV_X4 _u0_U21549  ( .A(1'b1), .ZN(_u0_pointer4_s[10] ) );
INV_X4 _u0_U21547  ( .A(1'b1), .ZN(_u0_pointer4_s[9] ) );
INV_X4 _u0_U21545  ( .A(1'b1), .ZN(_u0_pointer4_s[8] ) );
INV_X4 _u0_U21543  ( .A(1'b1), .ZN(_u0_pointer4_s[7] ) );
INV_X4 _u0_U21541  ( .A(1'b1), .ZN(_u0_pointer4_s[6] ) );
INV_X4 _u0_U21539  ( .A(1'b1), .ZN(_u0_pointer4_s[5] ) );
INV_X4 _u0_U21537  ( .A(1'b1), .ZN(_u0_pointer4_s[4] ) );
INV_X4 _u0_U21535  ( .A(1'b1), .ZN(_u0_pointer4_s[3] ) );
INV_X4 _u0_U21533  ( .A(1'b1), .ZN(_u0_pointer4_s[2] ) );
INV_X4 _u0_U21531  ( .A(1'b1), .ZN(_u0_pointer4_s[1] ) );
INV_X4 _u0_U21529  ( .A(1'b1), .ZN(_u0_pointer4_s[0] ) );
INV_X4 _u0_U21527  ( .A(1'b1), .ZN(_u0_ch4_csr[31] ) );
INV_X4 _u0_U21525  ( .A(1'b1), .ZN(_u0_ch4_csr[30] ) );
INV_X4 _u0_U21523  ( .A(1'b1), .ZN(_u0_ch4_csr[29] ) );
INV_X4 _u0_U21521  ( .A(1'b1), .ZN(_u0_ch4_csr[28] ) );
INV_X4 _u0_U21519  ( .A(1'b1), .ZN(_u0_ch4_csr[27] ) );
INV_X4 _u0_U21517  ( .A(1'b1), .ZN(_u0_ch4_csr[26] ) );
INV_X4 _u0_U21515  ( .A(1'b1), .ZN(_u0_ch4_csr[25] ) );
INV_X4 _u0_U21513  ( .A(1'b1), .ZN(_u0_ch4_csr[24] ) );
INV_X4 _u0_U21511  ( .A(1'b1), .ZN(_u0_ch4_csr[23] ) );
INV_X4 _u0_U21509  ( .A(1'b1), .ZN(_u0_ch4_csr[22] ) );
INV_X4 _u0_U21507  ( .A(1'b1), .ZN(_u0_ch4_csr[21] ) );
INV_X4 _u0_U21505  ( .A(1'b1), .ZN(_u0_ch4_csr[20] ) );
INV_X4 _u0_U21503  ( .A(1'b1), .ZN(_u0_ch4_csr[19] ) );
INV_X4 _u0_U21501  ( .A(1'b1), .ZN(_u0_ch4_csr[18] ) );
INV_X4 _u0_U21499  ( .A(1'b1), .ZN(_u0_ch4_csr[17] ) );
INV_X4 _u0_U21497  ( .A(1'b1), .ZN(_u0_ch4_csr[16] ) );
INV_X4 _u0_U21495  ( .A(1'b1), .ZN(_u0_ch4_csr[15] ) );
INV_X4 _u0_U21493  ( .A(1'b1), .ZN(_u0_ch4_csr[14] ) );
INV_X4 _u0_U21491  ( .A(1'b1), .ZN(_u0_ch4_csr[13] ) );
INV_X4 _u0_U21489  ( .A(1'b1), .ZN(_u0_ch4_csr[12] ) );
INV_X4 _u0_U21487  ( .A(1'b1), .ZN(_u0_ch4_csr[11] ) );
INV_X4 _u0_U21485  ( .A(1'b1), .ZN(_u0_ch4_csr[10] ) );
INV_X4 _u0_U21483  ( .A(1'b1), .ZN(_u0_ch4_csr[9] ) );
INV_X4 _u0_U21481  ( .A(1'b1), .ZN(_u0_ch4_csr[8] ) );
INV_X4 _u0_U21479  ( .A(1'b1), .ZN(_u0_ch4_csr[7] ) );
INV_X4 _u0_U21477  ( .A(1'b1), .ZN(_u0_ch4_csr[6] ) );
INV_X4 _u0_U21475  ( .A(1'b1), .ZN(_u0_ch4_csr[5] ) );
INV_X4 _u0_U21473  ( .A(1'b1), .ZN(_u0_ch4_csr[4] ) );
INV_X4 _u0_U21471  ( .A(1'b1), .ZN(_u0_ch4_csr[3] ) );
INV_X4 _u0_U21469  ( .A(1'b1), .ZN(_u0_ch4_csr[2] ) );
INV_X4 _u0_U21467  ( .A(1'b1), .ZN(_u0_ch4_csr[1] ) );
INV_X4 _u0_U21465  ( .A(1'b1), .ZN(_u0_ch4_csr[0] ) );
INV_X4 _u0_U21463  ( .A(1'b1), .ZN(_u0_ch4_txsz[31] ) );
INV_X4 _u0_U21461  ( .A(1'b1), .ZN(_u0_ch4_txsz[30] ) );
INV_X4 _u0_U21459  ( .A(1'b1), .ZN(_u0_ch4_txsz[29] ) );
INV_X4 _u0_U21457  ( .A(1'b1), .ZN(_u0_ch4_txsz[28] ) );
INV_X4 _u0_U21455  ( .A(1'b1), .ZN(_u0_ch4_txsz[27] ) );
INV_X4 _u0_U21453  ( .A(1'b1), .ZN(_u0_ch4_txsz[26] ) );
INV_X4 _u0_U21451  ( .A(1'b1), .ZN(_u0_ch4_txsz[25] ) );
INV_X4 _u0_U21449  ( .A(1'b1), .ZN(_u0_ch4_txsz[24] ) );
INV_X4 _u0_U21447  ( .A(1'b1), .ZN(_u0_ch4_txsz[23] ) );
INV_X4 _u0_U21445  ( .A(1'b1), .ZN(_u0_ch4_txsz[22] ) );
INV_X4 _u0_U21443  ( .A(1'b1), .ZN(_u0_ch4_txsz[21] ) );
INV_X4 _u0_U21441  ( .A(1'b1), .ZN(_u0_ch4_txsz[20] ) );
INV_X4 _u0_U21439  ( .A(1'b1), .ZN(_u0_ch4_txsz[19] ) );
INV_X4 _u0_U21437  ( .A(1'b1), .ZN(_u0_ch4_txsz[18] ) );
INV_X4 _u0_U21435  ( .A(1'b1), .ZN(_u0_ch4_txsz[17] ) );
INV_X4 _u0_U21433  ( .A(1'b1), .ZN(_u0_ch4_txsz[16] ) );
INV_X4 _u0_U21431  ( .A(1'b1), .ZN(_u0_ch4_txsz[15] ) );
INV_X4 _u0_U21429  ( .A(1'b1), .ZN(_u0_ch4_txsz[14] ) );
INV_X4 _u0_U21427  ( .A(1'b1), .ZN(_u0_ch4_txsz[13] ) );
INV_X4 _u0_U21425  ( .A(1'b1), .ZN(_u0_ch4_txsz[12] ) );
INV_X4 _u0_U21423  ( .A(1'b1), .ZN(_u0_ch4_txsz[11] ) );
INV_X4 _u0_U21421  ( .A(1'b1), .ZN(_u0_ch4_txsz[10] ) );
INV_X4 _u0_U21419  ( .A(1'b1), .ZN(_u0_ch4_txsz[9] ) );
INV_X4 _u0_U21417  ( .A(1'b1), .ZN(_u0_ch4_txsz[8] ) );
INV_X4 _u0_U21415  ( .A(1'b1), .ZN(_u0_ch4_txsz[7] ) );
INV_X4 _u0_U21413  ( .A(1'b1), .ZN(_u0_ch4_txsz[6] ) );
INV_X4 _u0_U21411  ( .A(1'b1), .ZN(_u0_ch4_txsz[5] ) );
INV_X4 _u0_U21409  ( .A(1'b1), .ZN(_u0_ch4_txsz[4] ) );
INV_X4 _u0_U21407  ( .A(1'b1), .ZN(_u0_ch4_txsz[3] ) );
INV_X4 _u0_U21405  ( .A(1'b1), .ZN(_u0_ch4_txsz[2] ) );
INV_X4 _u0_U21403  ( .A(1'b1), .ZN(_u0_ch4_txsz[1] ) );
INV_X4 _u0_U21401  ( .A(1'b1), .ZN(_u0_ch4_txsz[0] ) );
INV_X4 _u0_U21399  ( .A(1'b1), .ZN(_u0_ch4_adr0[31] ) );
INV_X4 _u0_U21397  ( .A(1'b1), .ZN(_u0_ch4_adr0[30] ) );
INV_X4 _u0_U21395  ( .A(1'b1), .ZN(_u0_ch4_adr0[29] ) );
INV_X4 _u0_U21393  ( .A(1'b1), .ZN(_u0_ch4_adr0[28] ) );
INV_X4 _u0_U21391  ( .A(1'b1), .ZN(_u0_ch4_adr0[27] ) );
INV_X4 _u0_U21389  ( .A(1'b1), .ZN(_u0_ch4_adr0[26] ) );
INV_X4 _u0_U21387  ( .A(1'b1), .ZN(_u0_ch4_adr0[25] ) );
INV_X4 _u0_U21385  ( .A(1'b1), .ZN(_u0_ch4_adr0[24] ) );
INV_X4 _u0_U21383  ( .A(1'b1), .ZN(_u0_ch4_adr0[23] ) );
INV_X4 _u0_U21381  ( .A(1'b1), .ZN(_u0_ch4_adr0[22] ) );
INV_X4 _u0_U21379  ( .A(1'b1), .ZN(_u0_ch4_adr0[21] ) );
INV_X4 _u0_U21377  ( .A(1'b1), .ZN(_u0_ch4_adr0[20] ) );
INV_X4 _u0_U21375  ( .A(1'b1), .ZN(_u0_ch4_adr0[19] ) );
INV_X4 _u0_U21373  ( .A(1'b1), .ZN(_u0_ch4_adr0[18] ) );
INV_X4 _u0_U21371  ( .A(1'b1), .ZN(_u0_ch4_adr0[17] ) );
INV_X4 _u0_U21369  ( .A(1'b1), .ZN(_u0_ch4_adr0[16] ) );
INV_X4 _u0_U21367  ( .A(1'b1), .ZN(_u0_ch4_adr0[15] ) );
INV_X4 _u0_U21365  ( .A(1'b1), .ZN(_u0_ch4_adr0[14] ) );
INV_X4 _u0_U21363  ( .A(1'b1), .ZN(_u0_ch4_adr0[13] ) );
INV_X4 _u0_U21361  ( .A(1'b1), .ZN(_u0_ch4_adr0[12] ) );
INV_X4 _u0_U21359  ( .A(1'b1), .ZN(_u0_ch4_adr0[11] ) );
INV_X4 _u0_U21357  ( .A(1'b1), .ZN(_u0_ch4_adr0[10] ) );
INV_X4 _u0_U21355  ( .A(1'b1), .ZN(_u0_ch4_adr0[9] ) );
INV_X4 _u0_U21353  ( .A(1'b1), .ZN(_u0_ch4_adr0[8] ) );
INV_X4 _u0_U21351  ( .A(1'b1), .ZN(_u0_ch4_adr0[7] ) );
INV_X4 _u0_U21349  ( .A(1'b1), .ZN(_u0_ch4_adr0[6] ) );
INV_X4 _u0_U21347  ( .A(1'b1), .ZN(_u0_ch4_adr0[5] ) );
INV_X4 _u0_U21345  ( .A(1'b1), .ZN(_u0_ch4_adr0[4] ) );
INV_X4 _u0_U21343  ( .A(1'b1), .ZN(_u0_ch4_adr0[3] ) );
INV_X4 _u0_U21341  ( .A(1'b1), .ZN(_u0_ch4_adr0[2] ) );
INV_X4 _u0_U21339  ( .A(1'b1), .ZN(_u0_ch4_adr0[1] ) );
INV_X4 _u0_U21337  ( .A(1'b1), .ZN(_u0_ch4_adr0[0] ) );
INV_X4 _u0_U21335  ( .A(1'b1), .ZN(_u0_ch4_adr1[31] ) );
INV_X4 _u0_U21333  ( .A(1'b1), .ZN(_u0_ch4_adr1[30] ) );
INV_X4 _u0_U21331  ( .A(1'b1), .ZN(_u0_ch4_adr1[29] ) );
INV_X4 _u0_U21329  ( .A(1'b1), .ZN(_u0_ch4_adr1[28] ) );
INV_X4 _u0_U21327  ( .A(1'b1), .ZN(_u0_ch4_adr1[27] ) );
INV_X4 _u0_U21325  ( .A(1'b1), .ZN(_u0_ch4_adr1[26] ) );
INV_X4 _u0_U21323  ( .A(1'b1), .ZN(_u0_ch4_adr1[25] ) );
INV_X4 _u0_U21321  ( .A(1'b1), .ZN(_u0_ch4_adr1[24] ) );
INV_X4 _u0_U21319  ( .A(1'b1), .ZN(_u0_ch4_adr1[23] ) );
INV_X4 _u0_U21317  ( .A(1'b1), .ZN(_u0_ch4_adr1[22] ) );
INV_X4 _u0_U21315  ( .A(1'b1), .ZN(_u0_ch4_adr1[21] ) );
INV_X4 _u0_U21313  ( .A(1'b1), .ZN(_u0_ch4_adr1[20] ) );
INV_X4 _u0_U21311  ( .A(1'b1), .ZN(_u0_ch4_adr1[19] ) );
INV_X4 _u0_U21309  ( .A(1'b1), .ZN(_u0_ch4_adr1[18] ) );
INV_X4 _u0_U21307  ( .A(1'b1), .ZN(_u0_ch4_adr1[17] ) );
INV_X4 _u0_U21305  ( .A(1'b1), .ZN(_u0_ch4_adr1[16] ) );
INV_X4 _u0_U21303  ( .A(1'b1), .ZN(_u0_ch4_adr1[15] ) );
INV_X4 _u0_U21301  ( .A(1'b1), .ZN(_u0_ch4_adr1[14] ) );
INV_X4 _u0_U21299  ( .A(1'b1), .ZN(_u0_ch4_adr1[13] ) );
INV_X4 _u0_U21297  ( .A(1'b1), .ZN(_u0_ch4_adr1[12] ) );
INV_X4 _u0_U21295  ( .A(1'b1), .ZN(_u0_ch4_adr1[11] ) );
INV_X4 _u0_U21293  ( .A(1'b1), .ZN(_u0_ch4_adr1[10] ) );
INV_X4 _u0_U21291  ( .A(1'b1), .ZN(_u0_ch4_adr1[9] ) );
INV_X4 _u0_U21289  ( .A(1'b1), .ZN(_u0_ch4_adr1[8] ) );
INV_X4 _u0_U21287  ( .A(1'b1), .ZN(_u0_ch4_adr1[7] ) );
INV_X4 _u0_U21285  ( .A(1'b1), .ZN(_u0_ch4_adr1[6] ) );
INV_X4 _u0_U21283  ( .A(1'b1), .ZN(_u0_ch4_adr1[5] ) );
INV_X4 _u0_U21281  ( .A(1'b1), .ZN(_u0_ch4_adr1[4] ) );
INV_X4 _u0_U21279  ( .A(1'b1), .ZN(_u0_ch4_adr1[3] ) );
INV_X4 _u0_U21277  ( .A(1'b1), .ZN(_u0_ch4_adr1[2] ) );
INV_X4 _u0_U21275  ( .A(1'b1), .ZN(_u0_ch4_adr1[1] ) );
INV_X4 _u0_U21273  ( .A(1'b1), .ZN(_u0_ch4_adr1[0] ) );
INV_X4 _u0_U21271  ( .A(1'b0), .ZN(_u0_ch4_am0[31] ) );
INV_X4 _u0_U21269  ( .A(1'b0), .ZN(_u0_ch4_am0[30] ) );
INV_X4 _u0_U21267  ( .A(1'b0), .ZN(_u0_ch4_am0[29] ) );
INV_X4 _u0_U21265  ( .A(1'b0), .ZN(_u0_ch4_am0[28] ) );
INV_X4 _u0_U21263  ( .A(1'b0), .ZN(_u0_ch4_am0[27] ) );
INV_X4 _u0_U21261  ( .A(1'b0), .ZN(_u0_ch4_am0[26] ) );
INV_X4 _u0_U21259  ( .A(1'b0), .ZN(_u0_ch4_am0[25] ) );
INV_X4 _u0_U21257  ( .A(1'b0), .ZN(_u0_ch4_am0[24] ) );
INV_X4 _u0_U21255  ( .A(1'b0), .ZN(_u0_ch4_am0[23] ) );
INV_X4 _u0_U21253  ( .A(1'b0), .ZN(_u0_ch4_am0[22] ) );
INV_X4 _u0_U21251  ( .A(1'b0), .ZN(_u0_ch4_am0[21] ) );
INV_X4 _u0_U21249  ( .A(1'b0), .ZN(_u0_ch4_am0[20] ) );
INV_X4 _u0_U21247  ( .A(1'b0), .ZN(_u0_ch4_am0[19] ) );
INV_X4 _u0_U21245  ( .A(1'b0), .ZN(_u0_ch4_am0[18] ) );
INV_X4 _u0_U21243  ( .A(1'b0), .ZN(_u0_ch4_am0[17] ) );
INV_X4 _u0_U21241  ( .A(1'b0), .ZN(_u0_ch4_am0[16] ) );
INV_X4 _u0_U21239  ( .A(1'b0), .ZN(_u0_ch4_am0[15] ) );
INV_X4 _u0_U21237  ( .A(1'b0), .ZN(_u0_ch4_am0[14] ) );
INV_X4 _u0_U21235  ( .A(1'b0), .ZN(_u0_ch4_am0[13] ) );
INV_X4 _u0_U21233  ( .A(1'b0), .ZN(_u0_ch4_am0[12] ) );
INV_X4 _u0_U21231  ( .A(1'b0), .ZN(_u0_ch4_am0[11] ) );
INV_X4 _u0_U21229  ( .A(1'b0), .ZN(_u0_ch4_am0[10] ) );
INV_X4 _u0_U21227  ( .A(1'b0), .ZN(_u0_ch4_am0[9] ) );
INV_X4 _u0_U21225  ( .A(1'b0), .ZN(_u0_ch4_am0[8] ) );
INV_X4 _u0_U21223  ( .A(1'b0), .ZN(_u0_ch4_am0[7] ) );
INV_X4 _u0_U21221  ( .A(1'b0), .ZN(_u0_ch4_am0[6] ) );
INV_X4 _u0_U21219  ( .A(1'b0), .ZN(_u0_ch4_am0[5] ) );
INV_X4 _u0_U21217  ( .A(1'b0), .ZN(_u0_ch4_am0[4] ) );
INV_X4 _u0_U21215  ( .A(1'b1), .ZN(_u0_ch4_am0[3] ) );
INV_X4 _u0_U21213  ( .A(1'b1), .ZN(_u0_ch4_am0[2] ) );
INV_X4 _u0_U21211  ( .A(1'b1), .ZN(_u0_ch4_am0[1] ) );
INV_X4 _u0_U21209  ( .A(1'b1), .ZN(_u0_ch4_am0[0] ) );
INV_X4 _u0_U21207  ( .A(1'b0), .ZN(_u0_ch4_am1[31] ) );
INV_X4 _u0_U21205  ( .A(1'b0), .ZN(_u0_ch4_am1[30] ) );
INV_X4 _u0_U21203  ( .A(1'b0), .ZN(_u0_ch4_am1[29] ) );
INV_X4 _u0_U21201  ( .A(1'b0), .ZN(_u0_ch4_am1[28] ) );
INV_X4 _u0_U21199  ( .A(1'b0), .ZN(_u0_ch4_am1[27] ) );
INV_X4 _u0_U21197  ( .A(1'b0), .ZN(_u0_ch4_am1[26] ) );
INV_X4 _u0_U21195  ( .A(1'b0), .ZN(_u0_ch4_am1[25] ) );
INV_X4 _u0_U21193  ( .A(1'b0), .ZN(_u0_ch4_am1[24] ) );
INV_X4 _u0_U21191  ( .A(1'b0), .ZN(_u0_ch4_am1[23] ) );
INV_X4 _u0_U21189  ( .A(1'b0), .ZN(_u0_ch4_am1[22] ) );
INV_X4 _u0_U21187  ( .A(1'b0), .ZN(_u0_ch4_am1[21] ) );
INV_X4 _u0_U21185  ( .A(1'b0), .ZN(_u0_ch4_am1[20] ) );
INV_X4 _u0_U21183  ( .A(1'b0), .ZN(_u0_ch4_am1[19] ) );
INV_X4 _u0_U21181  ( .A(1'b0), .ZN(_u0_ch4_am1[18] ) );
INV_X4 _u0_U21179  ( .A(1'b0), .ZN(_u0_ch4_am1[17] ) );
INV_X4 _u0_U21177  ( .A(1'b0), .ZN(_u0_ch4_am1[16] ) );
INV_X4 _u0_U21175  ( .A(1'b0), .ZN(_u0_ch4_am1[15] ) );
INV_X4 _u0_U21173  ( .A(1'b0), .ZN(_u0_ch4_am1[14] ) );
INV_X4 _u0_U21171  ( .A(1'b0), .ZN(_u0_ch4_am1[13] ) );
INV_X4 _u0_U21169  ( .A(1'b0), .ZN(_u0_ch4_am1[12] ) );
INV_X4 _u0_U21167  ( .A(1'b0), .ZN(_u0_ch4_am1[11] ) );
INV_X4 _u0_U21165  ( .A(1'b0), .ZN(_u0_ch4_am1[10] ) );
INV_X4 _u0_U21163  ( .A(1'b0), .ZN(_u0_ch4_am1[9] ) );
INV_X4 _u0_U21161  ( .A(1'b0), .ZN(_u0_ch4_am1[8] ) );
INV_X4 _u0_U21159  ( .A(1'b0), .ZN(_u0_ch4_am1[7] ) );
INV_X4 _u0_U21157  ( .A(1'b0), .ZN(_u0_ch4_am1[6] ) );
INV_X4 _u0_U21155  ( .A(1'b0), .ZN(_u0_ch4_am1[5] ) );
INV_X4 _u0_U21153  ( .A(1'b0), .ZN(_u0_ch4_am1[4] ) );
INV_X4 _u0_U21151  ( .A(1'b1), .ZN(_u0_ch4_am1[3] ) );
INV_X4 _u0_U21149  ( .A(1'b1), .ZN(_u0_ch4_am1[2] ) );
INV_X4 _u0_U21147  ( .A(1'b1), .ZN(_u0_ch4_am1[1] ) );
INV_X4 _u0_U21145  ( .A(1'b1), .ZN(_u0_ch4_am1[0] ) );
INV_X4 _u0_U21143  ( .A(1'b1), .ZN(_u0_pointer5[31] ) );
INV_X4 _u0_U21141  ( .A(1'b1), .ZN(_u0_pointer5[30] ) );
INV_X4 _u0_U21139  ( .A(1'b1), .ZN(_u0_pointer5[29] ) );
INV_X4 _u0_U21137  ( .A(1'b1), .ZN(_u0_pointer5[28] ) );
INV_X4 _u0_U21135  ( .A(1'b1), .ZN(_u0_pointer5[27] ) );
INV_X4 _u0_U21133  ( .A(1'b1), .ZN(_u0_pointer5[26] ) );
INV_X4 _u0_U21131  ( .A(1'b1), .ZN(_u0_pointer5[25] ) );
INV_X4 _u0_U21129  ( .A(1'b1), .ZN(_u0_pointer5[24] ) );
INV_X4 _u0_U21127  ( .A(1'b1), .ZN(_u0_pointer5[23] ) );
INV_X4 _u0_U21125  ( .A(1'b1), .ZN(_u0_pointer5[22] ) );
INV_X4 _u0_U21123  ( .A(1'b1), .ZN(_u0_pointer5[21] ) );
INV_X4 _u0_U21121  ( .A(1'b1), .ZN(_u0_pointer5[20] ) );
INV_X4 _u0_U21119  ( .A(1'b1), .ZN(_u0_pointer5[19] ) );
INV_X4 _u0_U21117  ( .A(1'b1), .ZN(_u0_pointer5[18] ) );
INV_X4 _u0_U21115  ( .A(1'b1), .ZN(_u0_pointer5[17] ) );
INV_X4 _u0_U21113  ( .A(1'b1), .ZN(_u0_pointer5[16] ) );
INV_X4 _u0_U21111  ( .A(1'b1), .ZN(_u0_pointer5[15] ) );
INV_X4 _u0_U21109  ( .A(1'b1), .ZN(_u0_pointer5[14] ) );
INV_X4 _u0_U21107  ( .A(1'b1), .ZN(_u0_pointer5[13] ) );
INV_X4 _u0_U21105  ( .A(1'b1), .ZN(_u0_pointer5[12] ) );
INV_X4 _u0_U21103  ( .A(1'b1), .ZN(_u0_pointer5[11] ) );
INV_X4 _u0_U21101  ( .A(1'b1), .ZN(_u0_pointer5[10] ) );
INV_X4 _u0_U21099  ( .A(1'b1), .ZN(_u0_pointer5[9] ) );
INV_X4 _u0_U21097  ( .A(1'b1), .ZN(_u0_pointer5[8] ) );
INV_X4 _u0_U21095  ( .A(1'b1), .ZN(_u0_pointer5[7] ) );
INV_X4 _u0_U21093  ( .A(1'b1), .ZN(_u0_pointer5[6] ) );
INV_X4 _u0_U21091  ( .A(1'b1), .ZN(_u0_pointer5[5] ) );
INV_X4 _u0_U21089  ( .A(1'b1), .ZN(_u0_pointer5[4] ) );
INV_X4 _u0_U21087  ( .A(1'b1), .ZN(_u0_pointer5[3] ) );
INV_X4 _u0_U21085  ( .A(1'b1), .ZN(_u0_pointer5[2] ) );
INV_X4 _u0_U21083  ( .A(1'b1), .ZN(_u0_pointer5[1] ) );
INV_X4 _u0_U21081  ( .A(1'b1), .ZN(_u0_pointer5[0] ) );
INV_X4 _u0_U21079  ( .A(1'b1), .ZN(_u0_pointer5_s[31] ) );
INV_X4 _u0_U21077  ( .A(1'b1), .ZN(_u0_pointer5_s[30] ) );
INV_X4 _u0_U21075  ( .A(1'b1), .ZN(_u0_pointer5_s[29] ) );
INV_X4 _u0_U21073  ( .A(1'b1), .ZN(_u0_pointer5_s[28] ) );
INV_X4 _u0_U21071  ( .A(1'b1), .ZN(_u0_pointer5_s[27] ) );
INV_X4 _u0_U21069  ( .A(1'b1), .ZN(_u0_pointer5_s[26] ) );
INV_X4 _u0_U21067  ( .A(1'b1), .ZN(_u0_pointer5_s[25] ) );
INV_X4 _u0_U21065  ( .A(1'b1), .ZN(_u0_pointer5_s[24] ) );
INV_X4 _u0_U21063  ( .A(1'b1), .ZN(_u0_pointer5_s[23] ) );
INV_X4 _u0_U21061  ( .A(1'b1), .ZN(_u0_pointer5_s[22] ) );
INV_X4 _u0_U21059  ( .A(1'b1), .ZN(_u0_pointer5_s[21] ) );
INV_X4 _u0_U21057  ( .A(1'b1), .ZN(_u0_pointer5_s[20] ) );
INV_X4 _u0_U21055  ( .A(1'b1), .ZN(_u0_pointer5_s[19] ) );
INV_X4 _u0_U21053  ( .A(1'b1), .ZN(_u0_pointer5_s[18] ) );
INV_X4 _u0_U21051  ( .A(1'b1), .ZN(_u0_pointer5_s[17] ) );
INV_X4 _u0_U21049  ( .A(1'b1), .ZN(_u0_pointer5_s[16] ) );
INV_X4 _u0_U21047  ( .A(1'b1), .ZN(_u0_pointer5_s[15] ) );
INV_X4 _u0_U21045  ( .A(1'b1), .ZN(_u0_pointer5_s[14] ) );
INV_X4 _u0_U21043  ( .A(1'b1), .ZN(_u0_pointer5_s[13] ) );
INV_X4 _u0_U21041  ( .A(1'b1), .ZN(_u0_pointer5_s[12] ) );
INV_X4 _u0_U21039  ( .A(1'b1), .ZN(_u0_pointer5_s[11] ) );
INV_X4 _u0_U21037  ( .A(1'b1), .ZN(_u0_pointer5_s[10] ) );
INV_X4 _u0_U21035  ( .A(1'b1), .ZN(_u0_pointer5_s[9] ) );
INV_X4 _u0_U21033  ( .A(1'b1), .ZN(_u0_pointer5_s[8] ) );
INV_X4 _u0_U21031  ( .A(1'b1), .ZN(_u0_pointer5_s[7] ) );
INV_X4 _u0_U21029  ( .A(1'b1), .ZN(_u0_pointer5_s[6] ) );
INV_X4 _u0_U21027  ( .A(1'b1), .ZN(_u0_pointer5_s[5] ) );
INV_X4 _u0_U21025  ( .A(1'b1), .ZN(_u0_pointer5_s[4] ) );
INV_X4 _u0_U21023  ( .A(1'b1), .ZN(_u0_pointer5_s[3] ) );
INV_X4 _u0_U21021  ( .A(1'b1), .ZN(_u0_pointer5_s[2] ) );
INV_X4 _u0_U21019  ( .A(1'b1), .ZN(_u0_pointer5_s[1] ) );
INV_X4 _u0_U21017  ( .A(1'b1), .ZN(_u0_pointer5_s[0] ) );
INV_X4 _u0_U21015  ( .A(1'b1), .ZN(_u0_ch5_csr[31] ) );
INV_X4 _u0_U21013  ( .A(1'b1), .ZN(_u0_ch5_csr[30] ) );
INV_X4 _u0_U21011  ( .A(1'b1), .ZN(_u0_ch5_csr[29] ) );
INV_X4 _u0_U21009  ( .A(1'b1), .ZN(_u0_ch5_csr[28] ) );
INV_X4 _u0_U21007  ( .A(1'b1), .ZN(_u0_ch5_csr[27] ) );
INV_X4 _u0_U21005  ( .A(1'b1), .ZN(_u0_ch5_csr[26] ) );
INV_X4 _u0_U21003  ( .A(1'b1), .ZN(_u0_ch5_csr[25] ) );
INV_X4 _u0_U21001  ( .A(1'b1), .ZN(_u0_ch5_csr[24] ) );
INV_X4 _u0_U20999  ( .A(1'b1), .ZN(_u0_ch5_csr[23] ) );
INV_X4 _u0_U20997  ( .A(1'b1), .ZN(_u0_ch5_csr[22] ) );
INV_X4 _u0_U20995  ( .A(1'b1), .ZN(_u0_ch5_csr[21] ) );
INV_X4 _u0_U20993  ( .A(1'b1), .ZN(_u0_ch5_csr[20] ) );
INV_X4 _u0_U20991  ( .A(1'b1), .ZN(_u0_ch5_csr[19] ) );
INV_X4 _u0_U20989  ( .A(1'b1), .ZN(_u0_ch5_csr[18] ) );
INV_X4 _u0_U20987  ( .A(1'b1), .ZN(_u0_ch5_csr[17] ) );
INV_X4 _u0_U20985  ( .A(1'b1), .ZN(_u0_ch5_csr[16] ) );
INV_X4 _u0_U20983  ( .A(1'b1), .ZN(_u0_ch5_csr[15] ) );
INV_X4 _u0_U20981  ( .A(1'b1), .ZN(_u0_ch5_csr[14] ) );
INV_X4 _u0_U20979  ( .A(1'b1), .ZN(_u0_ch5_csr[13] ) );
INV_X4 _u0_U20977  ( .A(1'b1), .ZN(_u0_ch5_csr[12] ) );
INV_X4 _u0_U20975  ( .A(1'b1), .ZN(_u0_ch5_csr[11] ) );
INV_X4 _u0_U20973  ( .A(1'b1), .ZN(_u0_ch5_csr[10] ) );
INV_X4 _u0_U20971  ( .A(1'b1), .ZN(_u0_ch5_csr[9] ) );
INV_X4 _u0_U20969  ( .A(1'b1), .ZN(_u0_ch5_csr[8] ) );
INV_X4 _u0_U20967  ( .A(1'b1), .ZN(_u0_ch5_csr[7] ) );
INV_X4 _u0_U20965  ( .A(1'b1), .ZN(_u0_ch5_csr[6] ) );
INV_X4 _u0_U20963  ( .A(1'b1), .ZN(_u0_ch5_csr[5] ) );
INV_X4 _u0_U20961  ( .A(1'b1), .ZN(_u0_ch5_csr[4] ) );
INV_X4 _u0_U20959  ( .A(1'b1), .ZN(_u0_ch5_csr[3] ) );
INV_X4 _u0_U20957  ( .A(1'b1), .ZN(_u0_ch5_csr[2] ) );
INV_X4 _u0_U20955  ( .A(1'b1), .ZN(_u0_ch5_csr[1] ) );
INV_X4 _u0_U20953  ( .A(1'b1), .ZN(_u0_ch5_csr[0] ) );
INV_X4 _u0_U20951  ( .A(1'b1), .ZN(_u0_ch5_txsz[31] ) );
INV_X4 _u0_U20949  ( .A(1'b1), .ZN(_u0_ch5_txsz[30] ) );
INV_X4 _u0_U20947  ( .A(1'b1), .ZN(_u0_ch5_txsz[29] ) );
INV_X4 _u0_U20945  ( .A(1'b1), .ZN(_u0_ch5_txsz[28] ) );
INV_X4 _u0_U20943  ( .A(1'b1), .ZN(_u0_ch5_txsz[27] ) );
INV_X4 _u0_U20941  ( .A(1'b1), .ZN(_u0_ch5_txsz[26] ) );
INV_X4 _u0_U20939  ( .A(1'b1), .ZN(_u0_ch5_txsz[25] ) );
INV_X4 _u0_U20937  ( .A(1'b1), .ZN(_u0_ch5_txsz[24] ) );
INV_X4 _u0_U20935  ( .A(1'b1), .ZN(_u0_ch5_txsz[23] ) );
INV_X4 _u0_U20933  ( .A(1'b1), .ZN(_u0_ch5_txsz[22] ) );
INV_X4 _u0_U20931  ( .A(1'b1), .ZN(_u0_ch5_txsz[21] ) );
INV_X4 _u0_U20929  ( .A(1'b1), .ZN(_u0_ch5_txsz[20] ) );
INV_X4 _u0_U20927  ( .A(1'b1), .ZN(_u0_ch5_txsz[19] ) );
INV_X4 _u0_U20925  ( .A(1'b1), .ZN(_u0_ch5_txsz[18] ) );
INV_X4 _u0_U20923  ( .A(1'b1), .ZN(_u0_ch5_txsz[17] ) );
INV_X4 _u0_U20921  ( .A(1'b1), .ZN(_u0_ch5_txsz[16] ) );
INV_X4 _u0_U20919  ( .A(1'b1), .ZN(_u0_ch5_txsz[15] ) );
INV_X4 _u0_U20917  ( .A(1'b1), .ZN(_u0_ch5_txsz[14] ) );
INV_X4 _u0_U20915  ( .A(1'b1), .ZN(_u0_ch5_txsz[13] ) );
INV_X4 _u0_U20913  ( .A(1'b1), .ZN(_u0_ch5_txsz[12] ) );
INV_X4 _u0_U20911  ( .A(1'b1), .ZN(_u0_ch5_txsz[11] ) );
INV_X4 _u0_U20909  ( .A(1'b1), .ZN(_u0_ch5_txsz[10] ) );
INV_X4 _u0_U20907  ( .A(1'b1), .ZN(_u0_ch5_txsz[9] ) );
INV_X4 _u0_U20905  ( .A(1'b1), .ZN(_u0_ch5_txsz[8] ) );
INV_X4 _u0_U20903  ( .A(1'b1), .ZN(_u0_ch5_txsz[7] ) );
INV_X4 _u0_U20901  ( .A(1'b1), .ZN(_u0_ch5_txsz[6] ) );
INV_X4 _u0_U20899  ( .A(1'b1), .ZN(_u0_ch5_txsz[5] ) );
INV_X4 _u0_U20897  ( .A(1'b1), .ZN(_u0_ch5_txsz[4] ) );
INV_X4 _u0_U20895  ( .A(1'b1), .ZN(_u0_ch5_txsz[3] ) );
INV_X4 _u0_U20893  ( .A(1'b1), .ZN(_u0_ch5_txsz[2] ) );
INV_X4 _u0_U20891  ( .A(1'b1), .ZN(_u0_ch5_txsz[1] ) );
INV_X4 _u0_U20889  ( .A(1'b1), .ZN(_u0_ch5_txsz[0] ) );
INV_X4 _u0_U20887  ( .A(1'b1), .ZN(_u0_ch5_adr0[31] ) );
INV_X4 _u0_U20885  ( .A(1'b1), .ZN(_u0_ch5_adr0[30] ) );
INV_X4 _u0_U20883  ( .A(1'b1), .ZN(_u0_ch5_adr0[29] ) );
INV_X4 _u0_U20881  ( .A(1'b1), .ZN(_u0_ch5_adr0[28] ) );
INV_X4 _u0_U20879  ( .A(1'b1), .ZN(_u0_ch5_adr0[27] ) );
INV_X4 _u0_U20877  ( .A(1'b1), .ZN(_u0_ch5_adr0[26] ) );
INV_X4 _u0_U20875  ( .A(1'b1), .ZN(_u0_ch5_adr0[25] ) );
INV_X4 _u0_U20873  ( .A(1'b1), .ZN(_u0_ch5_adr0[24] ) );
INV_X4 _u0_U20871  ( .A(1'b1), .ZN(_u0_ch5_adr0[23] ) );
INV_X4 _u0_U20869  ( .A(1'b1), .ZN(_u0_ch5_adr0[22] ) );
INV_X4 _u0_U20867  ( .A(1'b1), .ZN(_u0_ch5_adr0[21] ) );
INV_X4 _u0_U20865  ( .A(1'b1), .ZN(_u0_ch5_adr0[20] ) );
INV_X4 _u0_U20863  ( .A(1'b1), .ZN(_u0_ch5_adr0[19] ) );
INV_X4 _u0_U20861  ( .A(1'b1), .ZN(_u0_ch5_adr0[18] ) );
INV_X4 _u0_U20859  ( .A(1'b1), .ZN(_u0_ch5_adr0[17] ) );
INV_X4 _u0_U20857  ( .A(1'b1), .ZN(_u0_ch5_adr0[16] ) );
INV_X4 _u0_U20855  ( .A(1'b1), .ZN(_u0_ch5_adr0[15] ) );
INV_X4 _u0_U20853  ( .A(1'b1), .ZN(_u0_ch5_adr0[14] ) );
INV_X4 _u0_U20851  ( .A(1'b1), .ZN(_u0_ch5_adr0[13] ) );
INV_X4 _u0_U20849  ( .A(1'b1), .ZN(_u0_ch5_adr0[12] ) );
INV_X4 _u0_U20847  ( .A(1'b1), .ZN(_u0_ch5_adr0[11] ) );
INV_X4 _u0_U20845  ( .A(1'b1), .ZN(_u0_ch5_adr0[10] ) );
INV_X4 _u0_U20843  ( .A(1'b1), .ZN(_u0_ch5_adr0[9] ) );
INV_X4 _u0_U20841  ( .A(1'b1), .ZN(_u0_ch5_adr0[8] ) );
INV_X4 _u0_U20839  ( .A(1'b1), .ZN(_u0_ch5_adr0[7] ) );
INV_X4 _u0_U20837  ( .A(1'b1), .ZN(_u0_ch5_adr0[6] ) );
INV_X4 _u0_U20835  ( .A(1'b1), .ZN(_u0_ch5_adr0[5] ) );
INV_X4 _u0_U20833  ( .A(1'b1), .ZN(_u0_ch5_adr0[4] ) );
INV_X4 _u0_U20831  ( .A(1'b1), .ZN(_u0_ch5_adr0[3] ) );
INV_X4 _u0_U20829  ( .A(1'b1), .ZN(_u0_ch5_adr0[2] ) );
INV_X4 _u0_U20827  ( .A(1'b1), .ZN(_u0_ch5_adr0[1] ) );
INV_X4 _u0_U20825  ( .A(1'b1), .ZN(_u0_ch5_adr0[0] ) );
INV_X4 _u0_U20823  ( .A(1'b1), .ZN(_u0_ch5_adr1[31] ) );
INV_X4 _u0_U20821  ( .A(1'b1), .ZN(_u0_ch5_adr1[30] ) );
INV_X4 _u0_U20819  ( .A(1'b1), .ZN(_u0_ch5_adr1[29] ) );
INV_X4 _u0_U20817  ( .A(1'b1), .ZN(_u0_ch5_adr1[28] ) );
INV_X4 _u0_U20815  ( .A(1'b1), .ZN(_u0_ch5_adr1[27] ) );
INV_X4 _u0_U20813  ( .A(1'b1), .ZN(_u0_ch5_adr1[26] ) );
INV_X4 _u0_U20811  ( .A(1'b1), .ZN(_u0_ch5_adr1[25] ) );
INV_X4 _u0_U20809  ( .A(1'b1), .ZN(_u0_ch5_adr1[24] ) );
INV_X4 _u0_U20807  ( .A(1'b1), .ZN(_u0_ch5_adr1[23] ) );
INV_X4 _u0_U20805  ( .A(1'b1), .ZN(_u0_ch5_adr1[22] ) );
INV_X4 _u0_U20803  ( .A(1'b1), .ZN(_u0_ch5_adr1[21] ) );
INV_X4 _u0_U20801  ( .A(1'b1), .ZN(_u0_ch5_adr1[20] ) );
INV_X4 _u0_U20799  ( .A(1'b1), .ZN(_u0_ch5_adr1[19] ) );
INV_X4 _u0_U20797  ( .A(1'b1), .ZN(_u0_ch5_adr1[18] ) );
INV_X4 _u0_U20795  ( .A(1'b1), .ZN(_u0_ch5_adr1[17] ) );
INV_X4 _u0_U20793  ( .A(1'b1), .ZN(_u0_ch5_adr1[16] ) );
INV_X4 _u0_U20791  ( .A(1'b1), .ZN(_u0_ch5_adr1[15] ) );
INV_X4 _u0_U20789  ( .A(1'b1), .ZN(_u0_ch5_adr1[14] ) );
INV_X4 _u0_U20787  ( .A(1'b1), .ZN(_u0_ch5_adr1[13] ) );
INV_X4 _u0_U20785  ( .A(1'b1), .ZN(_u0_ch5_adr1[12] ) );
INV_X4 _u0_U20783  ( .A(1'b1), .ZN(_u0_ch5_adr1[11] ) );
INV_X4 _u0_U20781  ( .A(1'b1), .ZN(_u0_ch5_adr1[10] ) );
INV_X4 _u0_U20779  ( .A(1'b1), .ZN(_u0_ch5_adr1[9] ) );
INV_X4 _u0_U20777  ( .A(1'b1), .ZN(_u0_ch5_adr1[8] ) );
INV_X4 _u0_U20775  ( .A(1'b1), .ZN(_u0_ch5_adr1[7] ) );
INV_X4 _u0_U20773  ( .A(1'b1), .ZN(_u0_ch5_adr1[6] ) );
INV_X4 _u0_U20771  ( .A(1'b1), .ZN(_u0_ch5_adr1[5] ) );
INV_X4 _u0_U20769  ( .A(1'b1), .ZN(_u0_ch5_adr1[4] ) );
INV_X4 _u0_U20767  ( .A(1'b1), .ZN(_u0_ch5_adr1[3] ) );
INV_X4 _u0_U20765  ( .A(1'b1), .ZN(_u0_ch5_adr1[2] ) );
INV_X4 _u0_U20763  ( .A(1'b1), .ZN(_u0_ch5_adr1[1] ) );
INV_X4 _u0_U20761  ( .A(1'b1), .ZN(_u0_ch5_adr1[0] ) );
INV_X4 _u0_U20759  ( .A(1'b0), .ZN(_u0_ch5_am0[31] ) );
INV_X4 _u0_U20757  ( .A(1'b0), .ZN(_u0_ch5_am0[30] ) );
INV_X4 _u0_U20755  ( .A(1'b0), .ZN(_u0_ch5_am0[29] ) );
INV_X4 _u0_U20753  ( .A(1'b0), .ZN(_u0_ch5_am0[28] ) );
INV_X4 _u0_U20751  ( .A(1'b0), .ZN(_u0_ch5_am0[27] ) );
INV_X4 _u0_U20749  ( .A(1'b0), .ZN(_u0_ch5_am0[26] ) );
INV_X4 _u0_U20747  ( .A(1'b0), .ZN(_u0_ch5_am0[25] ) );
INV_X4 _u0_U20745  ( .A(1'b0), .ZN(_u0_ch5_am0[24] ) );
INV_X4 _u0_U20743  ( .A(1'b0), .ZN(_u0_ch5_am0[23] ) );
INV_X4 _u0_U20741  ( .A(1'b0), .ZN(_u0_ch5_am0[22] ) );
INV_X4 _u0_U20739  ( .A(1'b0), .ZN(_u0_ch5_am0[21] ) );
INV_X4 _u0_U20737  ( .A(1'b0), .ZN(_u0_ch5_am0[20] ) );
INV_X4 _u0_U20735  ( .A(1'b0), .ZN(_u0_ch5_am0[19] ) );
INV_X4 _u0_U20733  ( .A(1'b0), .ZN(_u0_ch5_am0[18] ) );
INV_X4 _u0_U20731  ( .A(1'b0), .ZN(_u0_ch5_am0[17] ) );
INV_X4 _u0_U20729  ( .A(1'b0), .ZN(_u0_ch5_am0[16] ) );
INV_X4 _u0_U20727  ( .A(1'b0), .ZN(_u0_ch5_am0[15] ) );
INV_X4 _u0_U20725  ( .A(1'b0), .ZN(_u0_ch5_am0[14] ) );
INV_X4 _u0_U20723  ( .A(1'b0), .ZN(_u0_ch5_am0[13] ) );
INV_X4 _u0_U20721  ( .A(1'b0), .ZN(_u0_ch5_am0[12] ) );
INV_X4 _u0_U20719  ( .A(1'b0), .ZN(_u0_ch5_am0[11] ) );
INV_X4 _u0_U20717  ( .A(1'b0), .ZN(_u0_ch5_am0[10] ) );
INV_X4 _u0_U20715  ( .A(1'b0), .ZN(_u0_ch5_am0[9] ) );
INV_X4 _u0_U20713  ( .A(1'b0), .ZN(_u0_ch5_am0[8] ) );
INV_X4 _u0_U20711  ( .A(1'b0), .ZN(_u0_ch5_am0[7] ) );
INV_X4 _u0_U20709  ( .A(1'b0), .ZN(_u0_ch5_am0[6] ) );
INV_X4 _u0_U20707  ( .A(1'b0), .ZN(_u0_ch5_am0[5] ) );
INV_X4 _u0_U20705  ( .A(1'b0), .ZN(_u0_ch5_am0[4] ) );
INV_X4 _u0_U20703  ( .A(1'b1), .ZN(_u0_ch5_am0[3] ) );
INV_X4 _u0_U20701  ( .A(1'b1), .ZN(_u0_ch5_am0[2] ) );
INV_X4 _u0_U20699  ( .A(1'b1), .ZN(_u0_ch5_am0[1] ) );
INV_X4 _u0_U20697  ( .A(1'b1), .ZN(_u0_ch5_am0[0] ) );
INV_X4 _u0_U20695  ( .A(1'b0), .ZN(_u0_ch5_am1[31] ) );
INV_X4 _u0_U20693  ( .A(1'b0), .ZN(_u0_ch5_am1[30] ) );
INV_X4 _u0_U20691  ( .A(1'b0), .ZN(_u0_ch5_am1[29] ) );
INV_X4 _u0_U20689  ( .A(1'b0), .ZN(_u0_ch5_am1[28] ) );
INV_X4 _u0_U20687  ( .A(1'b0), .ZN(_u0_ch5_am1[27] ) );
INV_X4 _u0_U20685  ( .A(1'b0), .ZN(_u0_ch5_am1[26] ) );
INV_X4 _u0_U20683  ( .A(1'b0), .ZN(_u0_ch5_am1[25] ) );
INV_X4 _u0_U20681  ( .A(1'b0), .ZN(_u0_ch5_am1[24] ) );
INV_X4 _u0_U20679  ( .A(1'b0), .ZN(_u0_ch5_am1[23] ) );
INV_X4 _u0_U20677  ( .A(1'b0), .ZN(_u0_ch5_am1[22] ) );
INV_X4 _u0_U20675  ( .A(1'b0), .ZN(_u0_ch5_am1[21] ) );
INV_X4 _u0_U20673  ( .A(1'b0), .ZN(_u0_ch5_am1[20] ) );
INV_X4 _u0_U20671  ( .A(1'b0), .ZN(_u0_ch5_am1[19] ) );
INV_X4 _u0_U20669  ( .A(1'b0), .ZN(_u0_ch5_am1[18] ) );
INV_X4 _u0_U20667  ( .A(1'b0), .ZN(_u0_ch5_am1[17] ) );
INV_X4 _u0_U20665  ( .A(1'b0), .ZN(_u0_ch5_am1[16] ) );
INV_X4 _u0_U20663  ( .A(1'b0), .ZN(_u0_ch5_am1[15] ) );
INV_X4 _u0_U20661  ( .A(1'b0), .ZN(_u0_ch5_am1[14] ) );
INV_X4 _u0_U20659  ( .A(1'b0), .ZN(_u0_ch5_am1[13] ) );
INV_X4 _u0_U20657  ( .A(1'b0), .ZN(_u0_ch5_am1[12] ) );
INV_X4 _u0_U20655  ( .A(1'b0), .ZN(_u0_ch5_am1[11] ) );
INV_X4 _u0_U20653  ( .A(1'b0), .ZN(_u0_ch5_am1[10] ) );
INV_X4 _u0_U20651  ( .A(1'b0), .ZN(_u0_ch5_am1[9] ) );
INV_X4 _u0_U20649  ( .A(1'b0), .ZN(_u0_ch5_am1[8] ) );
INV_X4 _u0_U20647  ( .A(1'b0), .ZN(_u0_ch5_am1[7] ) );
INV_X4 _u0_U20645  ( .A(1'b0), .ZN(_u0_ch5_am1[6] ) );
INV_X4 _u0_U20643  ( .A(1'b0), .ZN(_u0_ch5_am1[5] ) );
INV_X4 _u0_U20641  ( .A(1'b0), .ZN(_u0_ch5_am1[4] ) );
INV_X4 _u0_U20639  ( .A(1'b1), .ZN(_u0_ch5_am1[3] ) );
INV_X4 _u0_U20637  ( .A(1'b1), .ZN(_u0_ch5_am1[2] ) );
INV_X4 _u0_U20635  ( .A(1'b1), .ZN(_u0_ch5_am1[1] ) );
INV_X4 _u0_U20633  ( .A(1'b1), .ZN(_u0_ch5_am1[0] ) );
INV_X4 _u0_U20631  ( .A(1'b1), .ZN(_u0_pointer6[31] ) );
INV_X4 _u0_U20629  ( .A(1'b1), .ZN(_u0_pointer6[30] ) );
INV_X4 _u0_U20627  ( .A(1'b1), .ZN(_u0_pointer6[29] ) );
INV_X4 _u0_U20625  ( .A(1'b1), .ZN(_u0_pointer6[28] ) );
INV_X4 _u0_U20623  ( .A(1'b1), .ZN(_u0_pointer6[27] ) );
INV_X4 _u0_U20621  ( .A(1'b1), .ZN(_u0_pointer6[26] ) );
INV_X4 _u0_U20619  ( .A(1'b1), .ZN(_u0_pointer6[25] ) );
INV_X4 _u0_U20617  ( .A(1'b1), .ZN(_u0_pointer6[24] ) );
INV_X4 _u0_U20615  ( .A(1'b1), .ZN(_u0_pointer6[23] ) );
INV_X4 _u0_U20613  ( .A(1'b1), .ZN(_u0_pointer6[22] ) );
INV_X4 _u0_U20611  ( .A(1'b1), .ZN(_u0_pointer6[21] ) );
INV_X4 _u0_U20609  ( .A(1'b1), .ZN(_u0_pointer6[20] ) );
INV_X4 _u0_U20607  ( .A(1'b1), .ZN(_u0_pointer6[19] ) );
INV_X4 _u0_U20605  ( .A(1'b1), .ZN(_u0_pointer6[18] ) );
INV_X4 _u0_U20603  ( .A(1'b1), .ZN(_u0_pointer6[17] ) );
INV_X4 _u0_U20601  ( .A(1'b1), .ZN(_u0_pointer6[16] ) );
INV_X4 _u0_U20599  ( .A(1'b1), .ZN(_u0_pointer6[15] ) );
INV_X4 _u0_U20597  ( .A(1'b1), .ZN(_u0_pointer6[14] ) );
INV_X4 _u0_U20595  ( .A(1'b1), .ZN(_u0_pointer6[13] ) );
INV_X4 _u0_U20593  ( .A(1'b1), .ZN(_u0_pointer6[12] ) );
INV_X4 _u0_U20591  ( .A(1'b1), .ZN(_u0_pointer6[11] ) );
INV_X4 _u0_U20589  ( .A(1'b1), .ZN(_u0_pointer6[10] ) );
INV_X4 _u0_U20587  ( .A(1'b1), .ZN(_u0_pointer6[9] ) );
INV_X4 _u0_U20585  ( .A(1'b1), .ZN(_u0_pointer6[8] ) );
INV_X4 _u0_U20583  ( .A(1'b1), .ZN(_u0_pointer6[7] ) );
INV_X4 _u0_U20581  ( .A(1'b1), .ZN(_u0_pointer6[6] ) );
INV_X4 _u0_U20579  ( .A(1'b1), .ZN(_u0_pointer6[5] ) );
INV_X4 _u0_U20577  ( .A(1'b1), .ZN(_u0_pointer6[4] ) );
INV_X4 _u0_U20575  ( .A(1'b1), .ZN(_u0_pointer6[3] ) );
INV_X4 _u0_U20573  ( .A(1'b1), .ZN(_u0_pointer6[2] ) );
INV_X4 _u0_U20571  ( .A(1'b1), .ZN(_u0_pointer6[1] ) );
INV_X4 _u0_U20569  ( .A(1'b1), .ZN(_u0_pointer6[0] ) );
INV_X4 _u0_U20567  ( .A(1'b1), .ZN(_u0_pointer6_s[31] ) );
INV_X4 _u0_U20565  ( .A(1'b1), .ZN(_u0_pointer6_s[30] ) );
INV_X4 _u0_U20563  ( .A(1'b1), .ZN(_u0_pointer6_s[29] ) );
INV_X4 _u0_U20561  ( .A(1'b1), .ZN(_u0_pointer6_s[28] ) );
INV_X4 _u0_U20559  ( .A(1'b1), .ZN(_u0_pointer6_s[27] ) );
INV_X4 _u0_U20557  ( .A(1'b1), .ZN(_u0_pointer6_s[26] ) );
INV_X4 _u0_U20555  ( .A(1'b1), .ZN(_u0_pointer6_s[25] ) );
INV_X4 _u0_U20553  ( .A(1'b1), .ZN(_u0_pointer6_s[24] ) );
INV_X4 _u0_U20551  ( .A(1'b1), .ZN(_u0_pointer6_s[23] ) );
INV_X4 _u0_U20549  ( .A(1'b1), .ZN(_u0_pointer6_s[22] ) );
INV_X4 _u0_U20547  ( .A(1'b1), .ZN(_u0_pointer6_s[21] ) );
INV_X4 _u0_U20545  ( .A(1'b1), .ZN(_u0_pointer6_s[20] ) );
INV_X4 _u0_U20543  ( .A(1'b1), .ZN(_u0_pointer6_s[19] ) );
INV_X4 _u0_U20541  ( .A(1'b1), .ZN(_u0_pointer6_s[18] ) );
INV_X4 _u0_U20539  ( .A(1'b1), .ZN(_u0_pointer6_s[17] ) );
INV_X4 _u0_U20537  ( .A(1'b1), .ZN(_u0_pointer6_s[16] ) );
INV_X4 _u0_U20535  ( .A(1'b1), .ZN(_u0_pointer6_s[15] ) );
INV_X4 _u0_U20533  ( .A(1'b1), .ZN(_u0_pointer6_s[14] ) );
INV_X4 _u0_U20531  ( .A(1'b1), .ZN(_u0_pointer6_s[13] ) );
INV_X4 _u0_U20529  ( .A(1'b1), .ZN(_u0_pointer6_s[12] ) );
INV_X4 _u0_U20527  ( .A(1'b1), .ZN(_u0_pointer6_s[11] ) );
INV_X4 _u0_U20525  ( .A(1'b1), .ZN(_u0_pointer6_s[10] ) );
INV_X4 _u0_U20523  ( .A(1'b1), .ZN(_u0_pointer6_s[9] ) );
INV_X4 _u0_U20521  ( .A(1'b1), .ZN(_u0_pointer6_s[8] ) );
INV_X4 _u0_U20519  ( .A(1'b1), .ZN(_u0_pointer6_s[7] ) );
INV_X4 _u0_U20517  ( .A(1'b1), .ZN(_u0_pointer6_s[6] ) );
INV_X4 _u0_U20515  ( .A(1'b1), .ZN(_u0_pointer6_s[5] ) );
INV_X4 _u0_U20513  ( .A(1'b1), .ZN(_u0_pointer6_s[4] ) );
INV_X4 _u0_U20511  ( .A(1'b1), .ZN(_u0_pointer6_s[3] ) );
INV_X4 _u0_U20509  ( .A(1'b1), .ZN(_u0_pointer6_s[2] ) );
INV_X4 _u0_U20507  ( .A(1'b1), .ZN(_u0_pointer6_s[1] ) );
INV_X4 _u0_U20505  ( .A(1'b1), .ZN(_u0_pointer6_s[0] ) );
INV_X4 _u0_U20503  ( .A(1'b1), .ZN(_u0_ch6_csr[31] ) );
INV_X4 _u0_U20501  ( .A(1'b1), .ZN(_u0_ch6_csr[30] ) );
INV_X4 _u0_U20499  ( .A(1'b1), .ZN(_u0_ch6_csr[29] ) );
INV_X4 _u0_U20497  ( .A(1'b1), .ZN(_u0_ch6_csr[28] ) );
INV_X4 _u0_U20495  ( .A(1'b1), .ZN(_u0_ch6_csr[27] ) );
INV_X4 _u0_U20493  ( .A(1'b1), .ZN(_u0_ch6_csr[26] ) );
INV_X4 _u0_U20491  ( .A(1'b1), .ZN(_u0_ch6_csr[25] ) );
INV_X4 _u0_U20489  ( .A(1'b1), .ZN(_u0_ch6_csr[24] ) );
INV_X4 _u0_U20487  ( .A(1'b1), .ZN(_u0_ch6_csr[23] ) );
INV_X4 _u0_U20485  ( .A(1'b1), .ZN(_u0_ch6_csr[22] ) );
INV_X4 _u0_U20483  ( .A(1'b1), .ZN(_u0_ch6_csr[21] ) );
INV_X4 _u0_U20481  ( .A(1'b1), .ZN(_u0_ch6_csr[20] ) );
INV_X4 _u0_U20479  ( .A(1'b1), .ZN(_u0_ch6_csr[19] ) );
INV_X4 _u0_U20477  ( .A(1'b1), .ZN(_u0_ch6_csr[18] ) );
INV_X4 _u0_U20475  ( .A(1'b1), .ZN(_u0_ch6_csr[17] ) );
INV_X4 _u0_U20473  ( .A(1'b1), .ZN(_u0_ch6_csr[16] ) );
INV_X4 _u0_U20471  ( .A(1'b1), .ZN(_u0_ch6_csr[15] ) );
INV_X4 _u0_U20469  ( .A(1'b1), .ZN(_u0_ch6_csr[14] ) );
INV_X4 _u0_U20467  ( .A(1'b1), .ZN(_u0_ch6_csr[13] ) );
INV_X4 _u0_U20465  ( .A(1'b1), .ZN(_u0_ch6_csr[12] ) );
INV_X4 _u0_U20463  ( .A(1'b1), .ZN(_u0_ch6_csr[11] ) );
INV_X4 _u0_U20461  ( .A(1'b1), .ZN(_u0_ch6_csr[10] ) );
INV_X4 _u0_U20459  ( .A(1'b1), .ZN(_u0_ch6_csr[9] ) );
INV_X4 _u0_U20457  ( .A(1'b1), .ZN(_u0_ch6_csr[8] ) );
INV_X4 _u0_U20455  ( .A(1'b1), .ZN(_u0_ch6_csr[7] ) );
INV_X4 _u0_U20453  ( .A(1'b1), .ZN(_u0_ch6_csr[6] ) );
INV_X4 _u0_U20451  ( .A(1'b1), .ZN(_u0_ch6_csr[5] ) );
INV_X4 _u0_U20449  ( .A(1'b1), .ZN(_u0_ch6_csr[4] ) );
INV_X4 _u0_U20447  ( .A(1'b1), .ZN(_u0_ch6_csr[3] ) );
INV_X4 _u0_U20445  ( .A(1'b1), .ZN(_u0_ch6_csr[2] ) );
INV_X4 _u0_U20443  ( .A(1'b1), .ZN(_u0_ch6_csr[1] ) );
INV_X4 _u0_U20441  ( .A(1'b1), .ZN(_u0_ch6_csr[0] ) );
INV_X4 _u0_U20439  ( .A(1'b1), .ZN(_u0_ch6_txsz[31] ) );
INV_X4 _u0_U20437  ( .A(1'b1), .ZN(_u0_ch6_txsz[30] ) );
INV_X4 _u0_U20435  ( .A(1'b1), .ZN(_u0_ch6_txsz[29] ) );
INV_X4 _u0_U20433  ( .A(1'b1), .ZN(_u0_ch6_txsz[28] ) );
INV_X4 _u0_U20431  ( .A(1'b1), .ZN(_u0_ch6_txsz[27] ) );
INV_X4 _u0_U20429  ( .A(1'b1), .ZN(_u0_ch6_txsz[26] ) );
INV_X4 _u0_U20427  ( .A(1'b1), .ZN(_u0_ch6_txsz[25] ) );
INV_X4 _u0_U20425  ( .A(1'b1), .ZN(_u0_ch6_txsz[24] ) );
INV_X4 _u0_U20423  ( .A(1'b1), .ZN(_u0_ch6_txsz[23] ) );
INV_X4 _u0_U20421  ( .A(1'b1), .ZN(_u0_ch6_txsz[22] ) );
INV_X4 _u0_U20419  ( .A(1'b1), .ZN(_u0_ch6_txsz[21] ) );
INV_X4 _u0_U20417  ( .A(1'b1), .ZN(_u0_ch6_txsz[20] ) );
INV_X4 _u0_U20415  ( .A(1'b1), .ZN(_u0_ch6_txsz[19] ) );
INV_X4 _u0_U20413  ( .A(1'b1), .ZN(_u0_ch6_txsz[18] ) );
INV_X4 _u0_U20411  ( .A(1'b1), .ZN(_u0_ch6_txsz[17] ) );
INV_X4 _u0_U20409  ( .A(1'b1), .ZN(_u0_ch6_txsz[16] ) );
INV_X4 _u0_U20407  ( .A(1'b1), .ZN(_u0_ch6_txsz[15] ) );
INV_X4 _u0_U20405  ( .A(1'b1), .ZN(_u0_ch6_txsz[14] ) );
INV_X4 _u0_U20403  ( .A(1'b1), .ZN(_u0_ch6_txsz[13] ) );
INV_X4 _u0_U20401  ( .A(1'b1), .ZN(_u0_ch6_txsz[12] ) );
INV_X4 _u0_U20399  ( .A(1'b1), .ZN(_u0_ch6_txsz[11] ) );
INV_X4 _u0_U20397  ( .A(1'b1), .ZN(_u0_ch6_txsz[10] ) );
INV_X4 _u0_U20395  ( .A(1'b1), .ZN(_u0_ch6_txsz[9] ) );
INV_X4 _u0_U20393  ( .A(1'b1), .ZN(_u0_ch6_txsz[8] ) );
INV_X4 _u0_U20391  ( .A(1'b1), .ZN(_u0_ch6_txsz[7] ) );
INV_X4 _u0_U20389  ( .A(1'b1), .ZN(_u0_ch6_txsz[6] ) );
INV_X4 _u0_U20387  ( .A(1'b1), .ZN(_u0_ch6_txsz[5] ) );
INV_X4 _u0_U20385  ( .A(1'b1), .ZN(_u0_ch6_txsz[4] ) );
INV_X4 _u0_U20383  ( .A(1'b1), .ZN(_u0_ch6_txsz[3] ) );
INV_X4 _u0_U20381  ( .A(1'b1), .ZN(_u0_ch6_txsz[2] ) );
INV_X4 _u0_U20379  ( .A(1'b1), .ZN(_u0_ch6_txsz[1] ) );
INV_X4 _u0_U20377  ( .A(1'b1), .ZN(_u0_ch6_txsz[0] ) );
INV_X4 _u0_U20375  ( .A(1'b1), .ZN(_u0_ch6_adr0[31] ) );
INV_X4 _u0_U20373  ( .A(1'b1), .ZN(_u0_ch6_adr0[30] ) );
INV_X4 _u0_U20371  ( .A(1'b1), .ZN(_u0_ch6_adr0[29] ) );
INV_X4 _u0_U20369  ( .A(1'b1), .ZN(_u0_ch6_adr0[28] ) );
INV_X4 _u0_U20367  ( .A(1'b1), .ZN(_u0_ch6_adr0[27] ) );
INV_X4 _u0_U20365  ( .A(1'b1), .ZN(_u0_ch6_adr0[26] ) );
INV_X4 _u0_U20363  ( .A(1'b1), .ZN(_u0_ch6_adr0[25] ) );
INV_X4 _u0_U20361  ( .A(1'b1), .ZN(_u0_ch6_adr0[24] ) );
INV_X4 _u0_U20359  ( .A(1'b1), .ZN(_u0_ch6_adr0[23] ) );
INV_X4 _u0_U20357  ( .A(1'b1), .ZN(_u0_ch6_adr0[22] ) );
INV_X4 _u0_U20355  ( .A(1'b1), .ZN(_u0_ch6_adr0[21] ) );
INV_X4 _u0_U20353  ( .A(1'b1), .ZN(_u0_ch6_adr0[20] ) );
INV_X4 _u0_U20351  ( .A(1'b1), .ZN(_u0_ch6_adr0[19] ) );
INV_X4 _u0_U20349  ( .A(1'b1), .ZN(_u0_ch6_adr0[18] ) );
INV_X4 _u0_U20347  ( .A(1'b1), .ZN(_u0_ch6_adr0[17] ) );
INV_X4 _u0_U20345  ( .A(1'b1), .ZN(_u0_ch6_adr0[16] ) );
INV_X4 _u0_U20343  ( .A(1'b1), .ZN(_u0_ch6_adr0[15] ) );
INV_X4 _u0_U20341  ( .A(1'b1), .ZN(_u0_ch6_adr0[14] ) );
INV_X4 _u0_U20339  ( .A(1'b1), .ZN(_u0_ch6_adr0[13] ) );
INV_X4 _u0_U20337  ( .A(1'b1), .ZN(_u0_ch6_adr0[12] ) );
INV_X4 _u0_U20335  ( .A(1'b1), .ZN(_u0_ch6_adr0[11] ) );
INV_X4 _u0_U20333  ( .A(1'b1), .ZN(_u0_ch6_adr0[10] ) );
INV_X4 _u0_U20331  ( .A(1'b1), .ZN(_u0_ch6_adr0[9] ) );
INV_X4 _u0_U20329  ( .A(1'b1), .ZN(_u0_ch6_adr0[8] ) );
INV_X4 _u0_U20327  ( .A(1'b1), .ZN(_u0_ch6_adr0[7] ) );
INV_X4 _u0_U20325  ( .A(1'b1), .ZN(_u0_ch6_adr0[6] ) );
INV_X4 _u0_U20323  ( .A(1'b1), .ZN(_u0_ch6_adr0[5] ) );
INV_X4 _u0_U20321  ( .A(1'b1), .ZN(_u0_ch6_adr0[4] ) );
INV_X4 _u0_U20319  ( .A(1'b1), .ZN(_u0_ch6_adr0[3] ) );
INV_X4 _u0_U20317  ( .A(1'b1), .ZN(_u0_ch6_adr0[2] ) );
INV_X4 _u0_U20315  ( .A(1'b1), .ZN(_u0_ch6_adr0[1] ) );
INV_X4 _u0_U20313  ( .A(1'b1), .ZN(_u0_ch6_adr0[0] ) );
INV_X4 _u0_U20311  ( .A(1'b1), .ZN(_u0_ch6_adr1[31] ) );
INV_X4 _u0_U20309  ( .A(1'b1), .ZN(_u0_ch6_adr1[30] ) );
INV_X4 _u0_U20307  ( .A(1'b1), .ZN(_u0_ch6_adr1[29] ) );
INV_X4 _u0_U20305  ( .A(1'b1), .ZN(_u0_ch6_adr1[28] ) );
INV_X4 _u0_U20303  ( .A(1'b1), .ZN(_u0_ch6_adr1[27] ) );
INV_X4 _u0_U20301  ( .A(1'b1), .ZN(_u0_ch6_adr1[26] ) );
INV_X4 _u0_U20299  ( .A(1'b1), .ZN(_u0_ch6_adr1[25] ) );
INV_X4 _u0_U20297  ( .A(1'b1), .ZN(_u0_ch6_adr1[24] ) );
INV_X4 _u0_U20295  ( .A(1'b1), .ZN(_u0_ch6_adr1[23] ) );
INV_X4 _u0_U20293  ( .A(1'b1), .ZN(_u0_ch6_adr1[22] ) );
INV_X4 _u0_U20291  ( .A(1'b1), .ZN(_u0_ch6_adr1[21] ) );
INV_X4 _u0_U20289  ( .A(1'b1), .ZN(_u0_ch6_adr1[20] ) );
INV_X4 _u0_U20287  ( .A(1'b1), .ZN(_u0_ch6_adr1[19] ) );
INV_X4 _u0_U20285  ( .A(1'b1), .ZN(_u0_ch6_adr1[18] ) );
INV_X4 _u0_U20283  ( .A(1'b1), .ZN(_u0_ch6_adr1[17] ) );
INV_X4 _u0_U20281  ( .A(1'b1), .ZN(_u0_ch6_adr1[16] ) );
INV_X4 _u0_U20279  ( .A(1'b1), .ZN(_u0_ch6_adr1[15] ) );
INV_X4 _u0_U20277  ( .A(1'b1), .ZN(_u0_ch6_adr1[14] ) );
INV_X4 _u0_U20275  ( .A(1'b1), .ZN(_u0_ch6_adr1[13] ) );
INV_X4 _u0_U20273  ( .A(1'b1), .ZN(_u0_ch6_adr1[12] ) );
INV_X4 _u0_U20271  ( .A(1'b1), .ZN(_u0_ch6_adr1[11] ) );
INV_X4 _u0_U20269  ( .A(1'b1), .ZN(_u0_ch6_adr1[10] ) );
INV_X4 _u0_U20267  ( .A(1'b1), .ZN(_u0_ch6_adr1[9] ) );
INV_X4 _u0_U20265  ( .A(1'b1), .ZN(_u0_ch6_adr1[8] ) );
INV_X4 _u0_U20263  ( .A(1'b1), .ZN(_u0_ch6_adr1[7] ) );
INV_X4 _u0_U20261  ( .A(1'b1), .ZN(_u0_ch6_adr1[6] ) );
INV_X4 _u0_U20259  ( .A(1'b1), .ZN(_u0_ch6_adr1[5] ) );
INV_X4 _u0_U20257  ( .A(1'b1), .ZN(_u0_ch6_adr1[4] ) );
INV_X4 _u0_U20255  ( .A(1'b1), .ZN(_u0_ch6_adr1[3] ) );
INV_X4 _u0_U20253  ( .A(1'b1), .ZN(_u0_ch6_adr1[2] ) );
INV_X4 _u0_U20251  ( .A(1'b1), .ZN(_u0_ch6_adr1[1] ) );
INV_X4 _u0_U20249  ( .A(1'b1), .ZN(_u0_ch6_adr1[0] ) );
INV_X4 _u0_U20247  ( .A(1'b0), .ZN(_u0_ch6_am0[31] ) );
INV_X4 _u0_U20245  ( .A(1'b0), .ZN(_u0_ch6_am0[30] ) );
INV_X4 _u0_U20243  ( .A(1'b0), .ZN(_u0_ch6_am0[29] ) );
INV_X4 _u0_U20241  ( .A(1'b0), .ZN(_u0_ch6_am0[28] ) );
INV_X4 _u0_U20239  ( .A(1'b0), .ZN(_u0_ch6_am0[27] ) );
INV_X4 _u0_U20237  ( .A(1'b0), .ZN(_u0_ch6_am0[26] ) );
INV_X4 _u0_U20235  ( .A(1'b0), .ZN(_u0_ch6_am0[25] ) );
INV_X4 _u0_U20233  ( .A(1'b0), .ZN(_u0_ch6_am0[24] ) );
INV_X4 _u0_U20231  ( .A(1'b0), .ZN(_u0_ch6_am0[23] ) );
INV_X4 _u0_U20229  ( .A(1'b0), .ZN(_u0_ch6_am0[22] ) );
INV_X4 _u0_U20227  ( .A(1'b0), .ZN(_u0_ch6_am0[21] ) );
INV_X4 _u0_U20225  ( .A(1'b0), .ZN(_u0_ch6_am0[20] ) );
INV_X4 _u0_U20223  ( .A(1'b0), .ZN(_u0_ch6_am0[19] ) );
INV_X4 _u0_U20221  ( .A(1'b0), .ZN(_u0_ch6_am0[18] ) );
INV_X4 _u0_U20219  ( .A(1'b0), .ZN(_u0_ch6_am0[17] ) );
INV_X4 _u0_U20217  ( .A(1'b0), .ZN(_u0_ch6_am0[16] ) );
INV_X4 _u0_U20215  ( .A(1'b0), .ZN(_u0_ch6_am0[15] ) );
INV_X4 _u0_U20213  ( .A(1'b0), .ZN(_u0_ch6_am0[14] ) );
INV_X4 _u0_U20211  ( .A(1'b0), .ZN(_u0_ch6_am0[13] ) );
INV_X4 _u0_U20209  ( .A(1'b0), .ZN(_u0_ch6_am0[12] ) );
INV_X4 _u0_U20207  ( .A(1'b0), .ZN(_u0_ch6_am0[11] ) );
INV_X4 _u0_U20205  ( .A(1'b0), .ZN(_u0_ch6_am0[10] ) );
INV_X4 _u0_U20203  ( .A(1'b0), .ZN(_u0_ch6_am0[9] ) );
INV_X4 _u0_U20201  ( .A(1'b0), .ZN(_u0_ch6_am0[8] ) );
INV_X4 _u0_U20199  ( .A(1'b0), .ZN(_u0_ch6_am0[7] ) );
INV_X4 _u0_U20197  ( .A(1'b0), .ZN(_u0_ch6_am0[6] ) );
INV_X4 _u0_U20195  ( .A(1'b0), .ZN(_u0_ch6_am0[5] ) );
INV_X4 _u0_U20193  ( .A(1'b0), .ZN(_u0_ch6_am0[4] ) );
INV_X4 _u0_U20191  ( .A(1'b1), .ZN(_u0_ch6_am0[3] ) );
INV_X4 _u0_U20189  ( .A(1'b1), .ZN(_u0_ch6_am0[2] ) );
INV_X4 _u0_U20187  ( .A(1'b1), .ZN(_u0_ch6_am0[1] ) );
INV_X4 _u0_U20185  ( .A(1'b1), .ZN(_u0_ch6_am0[0] ) );
INV_X4 _u0_U20183  ( .A(1'b0), .ZN(_u0_ch6_am1[31] ) );
INV_X4 _u0_U20181  ( .A(1'b0), .ZN(_u0_ch6_am1[30] ) );
INV_X4 _u0_U20179  ( .A(1'b0), .ZN(_u0_ch6_am1[29] ) );
INV_X4 _u0_U20177  ( .A(1'b0), .ZN(_u0_ch6_am1[28] ) );
INV_X4 _u0_U20175  ( .A(1'b0), .ZN(_u0_ch6_am1[27] ) );
INV_X4 _u0_U20173  ( .A(1'b0), .ZN(_u0_ch6_am1[26] ) );
INV_X4 _u0_U20171  ( .A(1'b0), .ZN(_u0_ch6_am1[25] ) );
INV_X4 _u0_U20169  ( .A(1'b0), .ZN(_u0_ch6_am1[24] ) );
INV_X4 _u0_U20167  ( .A(1'b0), .ZN(_u0_ch6_am1[23] ) );
INV_X4 _u0_U20165  ( .A(1'b0), .ZN(_u0_ch6_am1[22] ) );
INV_X4 _u0_U20163  ( .A(1'b0), .ZN(_u0_ch6_am1[21] ) );
INV_X4 _u0_U20161  ( .A(1'b0), .ZN(_u0_ch6_am1[20] ) );
INV_X4 _u0_U20159  ( .A(1'b0), .ZN(_u0_ch6_am1[19] ) );
INV_X4 _u0_U20157  ( .A(1'b0), .ZN(_u0_ch6_am1[18] ) );
INV_X4 _u0_U20155  ( .A(1'b0), .ZN(_u0_ch6_am1[17] ) );
INV_X4 _u0_U20153  ( .A(1'b0), .ZN(_u0_ch6_am1[16] ) );
INV_X4 _u0_U20151  ( .A(1'b0), .ZN(_u0_ch6_am1[15] ) );
INV_X4 _u0_U20149  ( .A(1'b0), .ZN(_u0_ch6_am1[14] ) );
INV_X4 _u0_U20147  ( .A(1'b0), .ZN(_u0_ch6_am1[13] ) );
INV_X4 _u0_U20145  ( .A(1'b0), .ZN(_u0_ch6_am1[12] ) );
INV_X4 _u0_U20143  ( .A(1'b0), .ZN(_u0_ch6_am1[11] ) );
INV_X4 _u0_U20141  ( .A(1'b0), .ZN(_u0_ch6_am1[10] ) );
INV_X4 _u0_U20139  ( .A(1'b0), .ZN(_u0_ch6_am1[9] ) );
INV_X4 _u0_U20137  ( .A(1'b0), .ZN(_u0_ch6_am1[8] ) );
INV_X4 _u0_U20135  ( .A(1'b0), .ZN(_u0_ch6_am1[7] ) );
INV_X4 _u0_U20133  ( .A(1'b0), .ZN(_u0_ch6_am1[6] ) );
INV_X4 _u0_U20131  ( .A(1'b0), .ZN(_u0_ch6_am1[5] ) );
INV_X4 _u0_U20129  ( .A(1'b0), .ZN(_u0_ch6_am1[4] ) );
INV_X4 _u0_U20127  ( .A(1'b1), .ZN(_u0_ch6_am1[3] ) );
INV_X4 _u0_U20125  ( .A(1'b1), .ZN(_u0_ch6_am1[2] ) );
INV_X4 _u0_U20123  ( .A(1'b1), .ZN(_u0_ch6_am1[1] ) );
INV_X4 _u0_U20121  ( .A(1'b1), .ZN(_u0_ch6_am1[0] ) );
INV_X4 _u0_U20119  ( .A(1'b1), .ZN(_u0_pointer7[31] ) );
INV_X4 _u0_U20117  ( .A(1'b1), .ZN(_u0_pointer7[30] ) );
INV_X4 _u0_U20115  ( .A(1'b1), .ZN(_u0_pointer7[29] ) );
INV_X4 _u0_U20113  ( .A(1'b1), .ZN(_u0_pointer7[28] ) );
INV_X4 _u0_U20111  ( .A(1'b1), .ZN(_u0_pointer7[27] ) );
INV_X4 _u0_U20109  ( .A(1'b1), .ZN(_u0_pointer7[26] ) );
INV_X4 _u0_U20107  ( .A(1'b1), .ZN(_u0_pointer7[25] ) );
INV_X4 _u0_U20105  ( .A(1'b1), .ZN(_u0_pointer7[24] ) );
INV_X4 _u0_U20103  ( .A(1'b1), .ZN(_u0_pointer7[23] ) );
INV_X4 _u0_U20101  ( .A(1'b1), .ZN(_u0_pointer7[22] ) );
INV_X4 _u0_U20099  ( .A(1'b1), .ZN(_u0_pointer7[21] ) );
INV_X4 _u0_U20097  ( .A(1'b1), .ZN(_u0_pointer7[20] ) );
INV_X4 _u0_U20095  ( .A(1'b1), .ZN(_u0_pointer7[19] ) );
INV_X4 _u0_U20093  ( .A(1'b1), .ZN(_u0_pointer7[18] ) );
INV_X4 _u0_U20091  ( .A(1'b1), .ZN(_u0_pointer7[17] ) );
INV_X4 _u0_U20089  ( .A(1'b1), .ZN(_u0_pointer7[16] ) );
INV_X4 _u0_U20087  ( .A(1'b1), .ZN(_u0_pointer7[15] ) );
INV_X4 _u0_U20085  ( .A(1'b1), .ZN(_u0_pointer7[14] ) );
INV_X4 _u0_U20083  ( .A(1'b1), .ZN(_u0_pointer7[13] ) );
INV_X4 _u0_U20081  ( .A(1'b1), .ZN(_u0_pointer7[12] ) );
INV_X4 _u0_U20079  ( .A(1'b1), .ZN(_u0_pointer7[11] ) );
INV_X4 _u0_U20077  ( .A(1'b1), .ZN(_u0_pointer7[10] ) );
INV_X4 _u0_U20075  ( .A(1'b1), .ZN(_u0_pointer7[9] ) );
INV_X4 _u0_U20073  ( .A(1'b1), .ZN(_u0_pointer7[8] ) );
INV_X4 _u0_U20071  ( .A(1'b1), .ZN(_u0_pointer7[7] ) );
INV_X4 _u0_U20069  ( .A(1'b1), .ZN(_u0_pointer7[6] ) );
INV_X4 _u0_U20067  ( .A(1'b1), .ZN(_u0_pointer7[5] ) );
INV_X4 _u0_U20065  ( .A(1'b1), .ZN(_u0_pointer7[4] ) );
INV_X4 _u0_U20063  ( .A(1'b1), .ZN(_u0_pointer7[3] ) );
INV_X4 _u0_U20061  ( .A(1'b1), .ZN(_u0_pointer7[2] ) );
INV_X4 _u0_U20059  ( .A(1'b1), .ZN(_u0_pointer7[1] ) );
INV_X4 _u0_U20057  ( .A(1'b1), .ZN(_u0_pointer7[0] ) );
INV_X4 _u0_U20055  ( .A(1'b1), .ZN(_u0_pointer7_s[31] ) );
INV_X4 _u0_U20053  ( .A(1'b1), .ZN(_u0_pointer7_s[30] ) );
INV_X4 _u0_U20051  ( .A(1'b1), .ZN(_u0_pointer7_s[29] ) );
INV_X4 _u0_U20049  ( .A(1'b1), .ZN(_u0_pointer7_s[28] ) );
INV_X4 _u0_U20047  ( .A(1'b1), .ZN(_u0_pointer7_s[27] ) );
INV_X4 _u0_U20045  ( .A(1'b1), .ZN(_u0_pointer7_s[26] ) );
INV_X4 _u0_U20043  ( .A(1'b1), .ZN(_u0_pointer7_s[25] ) );
INV_X4 _u0_U20041  ( .A(1'b1), .ZN(_u0_pointer7_s[24] ) );
INV_X4 _u0_U20039  ( .A(1'b1), .ZN(_u0_pointer7_s[23] ) );
INV_X4 _u0_U20037  ( .A(1'b1), .ZN(_u0_pointer7_s[22] ) );
INV_X4 _u0_U20035  ( .A(1'b1), .ZN(_u0_pointer7_s[21] ) );
INV_X4 _u0_U20033  ( .A(1'b1), .ZN(_u0_pointer7_s[20] ) );
INV_X4 _u0_U20031  ( .A(1'b1), .ZN(_u0_pointer7_s[19] ) );
INV_X4 _u0_U20029  ( .A(1'b1), .ZN(_u0_pointer7_s[18] ) );
INV_X4 _u0_U20027  ( .A(1'b1), .ZN(_u0_pointer7_s[17] ) );
INV_X4 _u0_U20025  ( .A(1'b1), .ZN(_u0_pointer7_s[16] ) );
INV_X4 _u0_U20023  ( .A(1'b1), .ZN(_u0_pointer7_s[15] ) );
INV_X4 _u0_U20021  ( .A(1'b1), .ZN(_u0_pointer7_s[14] ) );
INV_X4 _u0_U20019  ( .A(1'b1), .ZN(_u0_pointer7_s[13] ) );
INV_X4 _u0_U20017  ( .A(1'b1), .ZN(_u0_pointer7_s[12] ) );
INV_X4 _u0_U20015  ( .A(1'b1), .ZN(_u0_pointer7_s[11] ) );
INV_X4 _u0_U20013  ( .A(1'b1), .ZN(_u0_pointer7_s[10] ) );
INV_X4 _u0_U20011  ( .A(1'b1), .ZN(_u0_pointer7_s[9] ) );
INV_X4 _u0_U20009  ( .A(1'b1), .ZN(_u0_pointer7_s[8] ) );
INV_X4 _u0_U20007  ( .A(1'b1), .ZN(_u0_pointer7_s[7] ) );
INV_X4 _u0_U20005  ( .A(1'b1), .ZN(_u0_pointer7_s[6] ) );
INV_X4 _u0_U20003  ( .A(1'b1), .ZN(_u0_pointer7_s[5] ) );
INV_X4 _u0_U20001  ( .A(1'b1), .ZN(_u0_pointer7_s[4] ) );
INV_X4 _u0_U19999  ( .A(1'b1), .ZN(_u0_pointer7_s[3] ) );
INV_X4 _u0_U19997  ( .A(1'b1), .ZN(_u0_pointer7_s[2] ) );
INV_X4 _u0_U19995  ( .A(1'b1), .ZN(_u0_pointer7_s[1] ) );
INV_X4 _u0_U19993  ( .A(1'b1), .ZN(_u0_pointer7_s[0] ) );
INV_X4 _u0_U19991  ( .A(1'b1), .ZN(_u0_ch7_csr[31] ) );
INV_X4 _u0_U19989  ( .A(1'b1), .ZN(_u0_ch7_csr[30] ) );
INV_X4 _u0_U19987  ( .A(1'b1), .ZN(_u0_ch7_csr[29] ) );
INV_X4 _u0_U19985  ( .A(1'b1), .ZN(_u0_ch7_csr[28] ) );
INV_X4 _u0_U19983  ( .A(1'b1), .ZN(_u0_ch7_csr[27] ) );
INV_X4 _u0_U19981  ( .A(1'b1), .ZN(_u0_ch7_csr[26] ) );
INV_X4 _u0_U19979  ( .A(1'b1), .ZN(_u0_ch7_csr[25] ) );
INV_X4 _u0_U19977  ( .A(1'b1), .ZN(_u0_ch7_csr[24] ) );
INV_X4 _u0_U19975  ( .A(1'b1), .ZN(_u0_ch7_csr[23] ) );
INV_X4 _u0_U19973  ( .A(1'b1), .ZN(_u0_ch7_csr[22] ) );
INV_X4 _u0_U19971  ( .A(1'b1), .ZN(_u0_ch7_csr[21] ) );
INV_X4 _u0_U19969  ( .A(1'b1), .ZN(_u0_ch7_csr[20] ) );
INV_X4 _u0_U19967  ( .A(1'b1), .ZN(_u0_ch7_csr[19] ) );
INV_X4 _u0_U19965  ( .A(1'b1), .ZN(_u0_ch7_csr[18] ) );
INV_X4 _u0_U19963  ( .A(1'b1), .ZN(_u0_ch7_csr[17] ) );
INV_X4 _u0_U19961  ( .A(1'b1), .ZN(_u0_ch7_csr[16] ) );
INV_X4 _u0_U19959  ( .A(1'b1), .ZN(_u0_ch7_csr[15] ) );
INV_X4 _u0_U19957  ( .A(1'b1), .ZN(_u0_ch7_csr[14] ) );
INV_X4 _u0_U19955  ( .A(1'b1), .ZN(_u0_ch7_csr[13] ) );
INV_X4 _u0_U19953  ( .A(1'b1), .ZN(_u0_ch7_csr[12] ) );
INV_X4 _u0_U19951  ( .A(1'b1), .ZN(_u0_ch7_csr[11] ) );
INV_X4 _u0_U19949  ( .A(1'b1), .ZN(_u0_ch7_csr[10] ) );
INV_X4 _u0_U19947  ( .A(1'b1), .ZN(_u0_ch7_csr[9] ) );
INV_X4 _u0_U19945  ( .A(1'b1), .ZN(_u0_ch7_csr[8] ) );
INV_X4 _u0_U19943  ( .A(1'b1), .ZN(_u0_ch7_csr[7] ) );
INV_X4 _u0_U19941  ( .A(1'b1), .ZN(_u0_ch7_csr[6] ) );
INV_X4 _u0_U19939  ( .A(1'b1), .ZN(_u0_ch7_csr[5] ) );
INV_X4 _u0_U19937  ( .A(1'b1), .ZN(_u0_ch7_csr[4] ) );
INV_X4 _u0_U19935  ( .A(1'b1), .ZN(_u0_ch7_csr[3] ) );
INV_X4 _u0_U19933  ( .A(1'b1), .ZN(_u0_ch7_csr[2] ) );
INV_X4 _u0_U19931  ( .A(1'b1), .ZN(_u0_ch7_csr[1] ) );
INV_X4 _u0_U19929  ( .A(1'b1), .ZN(_u0_ch7_csr[0] ) );
INV_X4 _u0_U19927  ( .A(1'b1), .ZN(_u0_ch7_txsz[31] ) );
INV_X4 _u0_U19925  ( .A(1'b1), .ZN(_u0_ch7_txsz[30] ) );
INV_X4 _u0_U19923  ( .A(1'b1), .ZN(_u0_ch7_txsz[29] ) );
INV_X4 _u0_U19921  ( .A(1'b1), .ZN(_u0_ch7_txsz[28] ) );
INV_X4 _u0_U19919  ( .A(1'b1), .ZN(_u0_ch7_txsz[27] ) );
INV_X4 _u0_U19917  ( .A(1'b1), .ZN(_u0_ch7_txsz[26] ) );
INV_X4 _u0_U19915  ( .A(1'b1), .ZN(_u0_ch7_txsz[25] ) );
INV_X4 _u0_U19913  ( .A(1'b1), .ZN(_u0_ch7_txsz[24] ) );
INV_X4 _u0_U19911  ( .A(1'b1), .ZN(_u0_ch7_txsz[23] ) );
INV_X4 _u0_U19909  ( .A(1'b1), .ZN(_u0_ch7_txsz[22] ) );
INV_X4 _u0_U19907  ( .A(1'b1), .ZN(_u0_ch7_txsz[21] ) );
INV_X4 _u0_U19905  ( .A(1'b1), .ZN(_u0_ch7_txsz[20] ) );
INV_X4 _u0_U19903  ( .A(1'b1), .ZN(_u0_ch7_txsz[19] ) );
INV_X4 _u0_U19901  ( .A(1'b1), .ZN(_u0_ch7_txsz[18] ) );
INV_X4 _u0_U19899  ( .A(1'b1), .ZN(_u0_ch7_txsz[17] ) );
INV_X4 _u0_U19897  ( .A(1'b1), .ZN(_u0_ch7_txsz[16] ) );
INV_X4 _u0_U19895  ( .A(1'b1), .ZN(_u0_ch7_txsz[15] ) );
INV_X4 _u0_U19893  ( .A(1'b1), .ZN(_u0_ch7_txsz[14] ) );
INV_X4 _u0_U19891  ( .A(1'b1), .ZN(_u0_ch7_txsz[13] ) );
INV_X4 _u0_U19889  ( .A(1'b1), .ZN(_u0_ch7_txsz[12] ) );
INV_X4 _u0_U19887  ( .A(1'b1), .ZN(_u0_ch7_txsz[11] ) );
INV_X4 _u0_U19885  ( .A(1'b1), .ZN(_u0_ch7_txsz[10] ) );
INV_X4 _u0_U19883  ( .A(1'b1), .ZN(_u0_ch7_txsz[9] ) );
INV_X4 _u0_U19881  ( .A(1'b1), .ZN(_u0_ch7_txsz[8] ) );
INV_X4 _u0_U19879  ( .A(1'b1), .ZN(_u0_ch7_txsz[7] ) );
INV_X4 _u0_U19877  ( .A(1'b1), .ZN(_u0_ch7_txsz[6] ) );
INV_X4 _u0_U19875  ( .A(1'b1), .ZN(_u0_ch7_txsz[5] ) );
INV_X4 _u0_U19873  ( .A(1'b1), .ZN(_u0_ch7_txsz[4] ) );
INV_X4 _u0_U19871  ( .A(1'b1), .ZN(_u0_ch7_txsz[3] ) );
INV_X4 _u0_U19869  ( .A(1'b1), .ZN(_u0_ch7_txsz[2] ) );
INV_X4 _u0_U19867  ( .A(1'b1), .ZN(_u0_ch7_txsz[1] ) );
INV_X4 _u0_U19865  ( .A(1'b1), .ZN(_u0_ch7_txsz[0] ) );
INV_X4 _u0_U19863  ( .A(1'b1), .ZN(_u0_ch7_adr0[31] ) );
INV_X4 _u0_U19861  ( .A(1'b1), .ZN(_u0_ch7_adr0[30] ) );
INV_X4 _u0_U19859  ( .A(1'b1), .ZN(_u0_ch7_adr0[29] ) );
INV_X4 _u0_U19857  ( .A(1'b1), .ZN(_u0_ch7_adr0[28] ) );
INV_X4 _u0_U19855  ( .A(1'b1), .ZN(_u0_ch7_adr0[27] ) );
INV_X4 _u0_U19853  ( .A(1'b1), .ZN(_u0_ch7_adr0[26] ) );
INV_X4 _u0_U19851  ( .A(1'b1), .ZN(_u0_ch7_adr0[25] ) );
INV_X4 _u0_U19849  ( .A(1'b1), .ZN(_u0_ch7_adr0[24] ) );
INV_X4 _u0_U19847  ( .A(1'b1), .ZN(_u0_ch7_adr0[23] ) );
INV_X4 _u0_U19845  ( .A(1'b1), .ZN(_u0_ch7_adr0[22] ) );
INV_X4 _u0_U19843  ( .A(1'b1), .ZN(_u0_ch7_adr0[21] ) );
INV_X4 _u0_U19841  ( .A(1'b1), .ZN(_u0_ch7_adr0[20] ) );
INV_X4 _u0_U19839  ( .A(1'b1), .ZN(_u0_ch7_adr0[19] ) );
INV_X4 _u0_U19837  ( .A(1'b1), .ZN(_u0_ch7_adr0[18] ) );
INV_X4 _u0_U19835  ( .A(1'b1), .ZN(_u0_ch7_adr0[17] ) );
INV_X4 _u0_U19833  ( .A(1'b1), .ZN(_u0_ch7_adr0[16] ) );
INV_X4 _u0_U19831  ( .A(1'b1), .ZN(_u0_ch7_adr0[15] ) );
INV_X4 _u0_U19829  ( .A(1'b1), .ZN(_u0_ch7_adr0[14] ) );
INV_X4 _u0_U19827  ( .A(1'b1), .ZN(_u0_ch7_adr0[13] ) );
INV_X4 _u0_U19825  ( .A(1'b1), .ZN(_u0_ch7_adr0[12] ) );
INV_X4 _u0_U19823  ( .A(1'b1), .ZN(_u0_ch7_adr0[11] ) );
INV_X4 _u0_U19821  ( .A(1'b1), .ZN(_u0_ch7_adr0[10] ) );
INV_X4 _u0_U19819  ( .A(1'b1), .ZN(_u0_ch7_adr0[9] ) );
INV_X4 _u0_U19817  ( .A(1'b1), .ZN(_u0_ch7_adr0[8] ) );
INV_X4 _u0_U19815  ( .A(1'b1), .ZN(_u0_ch7_adr0[7] ) );
INV_X4 _u0_U19813  ( .A(1'b1), .ZN(_u0_ch7_adr0[6] ) );
INV_X4 _u0_U19811  ( .A(1'b1), .ZN(_u0_ch7_adr0[5] ) );
INV_X4 _u0_U19809  ( .A(1'b1), .ZN(_u0_ch7_adr0[4] ) );
INV_X4 _u0_U19807  ( .A(1'b1), .ZN(_u0_ch7_adr0[3] ) );
INV_X4 _u0_U19805  ( .A(1'b1), .ZN(_u0_ch7_adr0[2] ) );
INV_X4 _u0_U19803  ( .A(1'b1), .ZN(_u0_ch7_adr0[1] ) );
INV_X4 _u0_U19801  ( .A(1'b1), .ZN(_u0_ch7_adr0[0] ) );
INV_X4 _u0_U19799  ( .A(1'b1), .ZN(_u0_ch7_adr1[31] ) );
INV_X4 _u0_U19797  ( .A(1'b1), .ZN(_u0_ch7_adr1[30] ) );
INV_X4 _u0_U19795  ( .A(1'b1), .ZN(_u0_ch7_adr1[29] ) );
INV_X4 _u0_U19793  ( .A(1'b1), .ZN(_u0_ch7_adr1[28] ) );
INV_X4 _u0_U19791  ( .A(1'b1), .ZN(_u0_ch7_adr1[27] ) );
INV_X4 _u0_U19789  ( .A(1'b1), .ZN(_u0_ch7_adr1[26] ) );
INV_X4 _u0_U19787  ( .A(1'b1), .ZN(_u0_ch7_adr1[25] ) );
INV_X4 _u0_U19785  ( .A(1'b1), .ZN(_u0_ch7_adr1[24] ) );
INV_X4 _u0_U19783  ( .A(1'b1), .ZN(_u0_ch7_adr1[23] ) );
INV_X4 _u0_U19781  ( .A(1'b1), .ZN(_u0_ch7_adr1[22] ) );
INV_X4 _u0_U19779  ( .A(1'b1), .ZN(_u0_ch7_adr1[21] ) );
INV_X4 _u0_U19777  ( .A(1'b1), .ZN(_u0_ch7_adr1[20] ) );
INV_X4 _u0_U19775  ( .A(1'b1), .ZN(_u0_ch7_adr1[19] ) );
INV_X4 _u0_U19773  ( .A(1'b1), .ZN(_u0_ch7_adr1[18] ) );
INV_X4 _u0_U19771  ( .A(1'b1), .ZN(_u0_ch7_adr1[17] ) );
INV_X4 _u0_U19769  ( .A(1'b1), .ZN(_u0_ch7_adr1[16] ) );
INV_X4 _u0_U19767  ( .A(1'b1), .ZN(_u0_ch7_adr1[15] ) );
INV_X4 _u0_U19765  ( .A(1'b1), .ZN(_u0_ch7_adr1[14] ) );
INV_X4 _u0_U19763  ( .A(1'b1), .ZN(_u0_ch7_adr1[13] ) );
INV_X4 _u0_U19761  ( .A(1'b1), .ZN(_u0_ch7_adr1[12] ) );
INV_X4 _u0_U19759  ( .A(1'b1), .ZN(_u0_ch7_adr1[11] ) );
INV_X4 _u0_U19757  ( .A(1'b1), .ZN(_u0_ch7_adr1[10] ) );
INV_X4 _u0_U19755  ( .A(1'b1), .ZN(_u0_ch7_adr1[9] ) );
INV_X4 _u0_U19753  ( .A(1'b1), .ZN(_u0_ch7_adr1[8] ) );
INV_X4 _u0_U19751  ( .A(1'b1), .ZN(_u0_ch7_adr1[7] ) );
INV_X4 _u0_U19749  ( .A(1'b1), .ZN(_u0_ch7_adr1[6] ) );
INV_X4 _u0_U19747  ( .A(1'b1), .ZN(_u0_ch7_adr1[5] ) );
INV_X4 _u0_U19745  ( .A(1'b1), .ZN(_u0_ch7_adr1[4] ) );
INV_X4 _u0_U19743  ( .A(1'b1), .ZN(_u0_ch7_adr1[3] ) );
INV_X4 _u0_U19741  ( .A(1'b1), .ZN(_u0_ch7_adr1[2] ) );
INV_X4 _u0_U19739  ( .A(1'b1), .ZN(_u0_ch7_adr1[1] ) );
INV_X4 _u0_U19737  ( .A(1'b1), .ZN(_u0_ch7_adr1[0] ) );
INV_X4 _u0_U19735  ( .A(1'b0), .ZN(_u0_ch7_am0[31] ) );
INV_X4 _u0_U19733  ( .A(1'b0), .ZN(_u0_ch7_am0[30] ) );
INV_X4 _u0_U19731  ( .A(1'b0), .ZN(_u0_ch7_am0[29] ) );
INV_X4 _u0_U19729  ( .A(1'b0), .ZN(_u0_ch7_am0[28] ) );
INV_X4 _u0_U19727  ( .A(1'b0), .ZN(_u0_ch7_am0[27] ) );
INV_X4 _u0_U19725  ( .A(1'b0), .ZN(_u0_ch7_am0[26] ) );
INV_X4 _u0_U19723  ( .A(1'b0), .ZN(_u0_ch7_am0[25] ) );
INV_X4 _u0_U19721  ( .A(1'b0), .ZN(_u0_ch7_am0[24] ) );
INV_X4 _u0_U19719  ( .A(1'b0), .ZN(_u0_ch7_am0[23] ) );
INV_X4 _u0_U19717  ( .A(1'b0), .ZN(_u0_ch7_am0[22] ) );
INV_X4 _u0_U19715  ( .A(1'b0), .ZN(_u0_ch7_am0[21] ) );
INV_X4 _u0_U19713  ( .A(1'b0), .ZN(_u0_ch7_am0[20] ) );
INV_X4 _u0_U19711  ( .A(1'b0), .ZN(_u0_ch7_am0[19] ) );
INV_X4 _u0_U19709  ( .A(1'b0), .ZN(_u0_ch7_am0[18] ) );
INV_X4 _u0_U19707  ( .A(1'b0), .ZN(_u0_ch7_am0[17] ) );
INV_X4 _u0_U19705  ( .A(1'b0), .ZN(_u0_ch7_am0[16] ) );
INV_X4 _u0_U19703  ( .A(1'b0), .ZN(_u0_ch7_am0[15] ) );
INV_X4 _u0_U19701  ( .A(1'b0), .ZN(_u0_ch7_am0[14] ) );
INV_X4 _u0_U19699  ( .A(1'b0), .ZN(_u0_ch7_am0[13] ) );
INV_X4 _u0_U19697  ( .A(1'b0), .ZN(_u0_ch7_am0[12] ) );
INV_X4 _u0_U19695  ( .A(1'b0), .ZN(_u0_ch7_am0[11] ) );
INV_X4 _u0_U19693  ( .A(1'b0), .ZN(_u0_ch7_am0[10] ) );
INV_X4 _u0_U19691  ( .A(1'b0), .ZN(_u0_ch7_am0[9] ) );
INV_X4 _u0_U19689  ( .A(1'b0), .ZN(_u0_ch7_am0[8] ) );
INV_X4 _u0_U19687  ( .A(1'b0), .ZN(_u0_ch7_am0[7] ) );
INV_X4 _u0_U19685  ( .A(1'b0), .ZN(_u0_ch7_am0[6] ) );
INV_X4 _u0_U19683  ( .A(1'b0), .ZN(_u0_ch7_am0[5] ) );
INV_X4 _u0_U19681  ( .A(1'b0), .ZN(_u0_ch7_am0[4] ) );
INV_X4 _u0_U19679  ( .A(1'b1), .ZN(_u0_ch7_am0[3] ) );
INV_X4 _u0_U19677  ( .A(1'b1), .ZN(_u0_ch7_am0[2] ) );
INV_X4 _u0_U19675  ( .A(1'b1), .ZN(_u0_ch7_am0[1] ) );
INV_X4 _u0_U19673  ( .A(1'b1), .ZN(_u0_ch7_am0[0] ) );
INV_X4 _u0_U19671  ( .A(1'b0), .ZN(_u0_ch7_am1[31] ) );
INV_X4 _u0_U19669  ( .A(1'b0), .ZN(_u0_ch7_am1[30] ) );
INV_X4 _u0_U19667  ( .A(1'b0), .ZN(_u0_ch7_am1[29] ) );
INV_X4 _u0_U19665  ( .A(1'b0), .ZN(_u0_ch7_am1[28] ) );
INV_X4 _u0_U19663  ( .A(1'b0), .ZN(_u0_ch7_am1[27] ) );
INV_X4 _u0_U19661  ( .A(1'b0), .ZN(_u0_ch7_am1[26] ) );
INV_X4 _u0_U19659  ( .A(1'b0), .ZN(_u0_ch7_am1[25] ) );
INV_X4 _u0_U19657  ( .A(1'b0), .ZN(_u0_ch7_am1[24] ) );
INV_X4 _u0_U19655  ( .A(1'b0), .ZN(_u0_ch7_am1[23] ) );
INV_X4 _u0_U19653  ( .A(1'b0), .ZN(_u0_ch7_am1[22] ) );
INV_X4 _u0_U19651  ( .A(1'b0), .ZN(_u0_ch7_am1[21] ) );
INV_X4 _u0_U19649  ( .A(1'b0), .ZN(_u0_ch7_am1[20] ) );
INV_X4 _u0_U19647  ( .A(1'b0), .ZN(_u0_ch7_am1[19] ) );
INV_X4 _u0_U19645  ( .A(1'b0), .ZN(_u0_ch7_am1[18] ) );
INV_X4 _u0_U19643  ( .A(1'b0), .ZN(_u0_ch7_am1[17] ) );
INV_X4 _u0_U19641  ( .A(1'b0), .ZN(_u0_ch7_am1[16] ) );
INV_X4 _u0_U19639  ( .A(1'b0), .ZN(_u0_ch7_am1[15] ) );
INV_X4 _u0_U19637  ( .A(1'b0), .ZN(_u0_ch7_am1[14] ) );
INV_X4 _u0_U19635  ( .A(1'b0), .ZN(_u0_ch7_am1[13] ) );
INV_X4 _u0_U19633  ( .A(1'b0), .ZN(_u0_ch7_am1[12] ) );
INV_X4 _u0_U19631  ( .A(1'b0), .ZN(_u0_ch7_am1[11] ) );
INV_X4 _u0_U19629  ( .A(1'b0), .ZN(_u0_ch7_am1[10] ) );
INV_X4 _u0_U19627  ( .A(1'b0), .ZN(_u0_ch7_am1[9] ) );
INV_X4 _u0_U19625  ( .A(1'b0), .ZN(_u0_ch7_am1[8] ) );
INV_X4 _u0_U19623  ( .A(1'b0), .ZN(_u0_ch7_am1[7] ) );
INV_X4 _u0_U19621  ( .A(1'b0), .ZN(_u0_ch7_am1[6] ) );
INV_X4 _u0_U19619  ( .A(1'b0), .ZN(_u0_ch7_am1[5] ) );
INV_X4 _u0_U19617  ( .A(1'b0), .ZN(_u0_ch7_am1[4] ) );
INV_X4 _u0_U19615  ( .A(1'b1), .ZN(_u0_ch7_am1[3] ) );
INV_X4 _u0_U19613  ( .A(1'b1), .ZN(_u0_ch7_am1[2] ) );
INV_X4 _u0_U19611  ( .A(1'b1), .ZN(_u0_ch7_am1[1] ) );
INV_X4 _u0_U19609  ( .A(1'b1), .ZN(_u0_ch7_am1[0] ) );
INV_X4 _u0_U19607  ( .A(1'b1), .ZN(_u0_pointer8[31] ) );
INV_X4 _u0_U19605  ( .A(1'b1), .ZN(_u0_pointer8[30] ) );
INV_X4 _u0_U19603  ( .A(1'b1), .ZN(_u0_pointer8[29] ) );
INV_X4 _u0_U19601  ( .A(1'b1), .ZN(_u0_pointer8[28] ) );
INV_X4 _u0_U19599  ( .A(1'b1), .ZN(_u0_pointer8[27] ) );
INV_X4 _u0_U19597  ( .A(1'b1), .ZN(_u0_pointer8[26] ) );
INV_X4 _u0_U19595  ( .A(1'b1), .ZN(_u0_pointer8[25] ) );
INV_X4 _u0_U19593  ( .A(1'b1), .ZN(_u0_pointer8[24] ) );
INV_X4 _u0_U19591  ( .A(1'b1), .ZN(_u0_pointer8[23] ) );
INV_X4 _u0_U19589  ( .A(1'b1), .ZN(_u0_pointer8[22] ) );
INV_X4 _u0_U19587  ( .A(1'b1), .ZN(_u0_pointer8[21] ) );
INV_X4 _u0_U19585  ( .A(1'b1), .ZN(_u0_pointer8[20] ) );
INV_X4 _u0_U19583  ( .A(1'b1), .ZN(_u0_pointer8[19] ) );
INV_X4 _u0_U19581  ( .A(1'b1), .ZN(_u0_pointer8[18] ) );
INV_X4 _u0_U19579  ( .A(1'b1), .ZN(_u0_pointer8[17] ) );
INV_X4 _u0_U19577  ( .A(1'b1), .ZN(_u0_pointer8[16] ) );
INV_X4 _u0_U19575  ( .A(1'b1), .ZN(_u0_pointer8[15] ) );
INV_X4 _u0_U19573  ( .A(1'b1), .ZN(_u0_pointer8[14] ) );
INV_X4 _u0_U19571  ( .A(1'b1), .ZN(_u0_pointer8[13] ) );
INV_X4 _u0_U19569  ( .A(1'b1), .ZN(_u0_pointer8[12] ) );
INV_X4 _u0_U19567  ( .A(1'b1), .ZN(_u0_pointer8[11] ) );
INV_X4 _u0_U19565  ( .A(1'b1), .ZN(_u0_pointer8[10] ) );
INV_X4 _u0_U19563  ( .A(1'b1), .ZN(_u0_pointer8[9] ) );
INV_X4 _u0_U19561  ( .A(1'b1), .ZN(_u0_pointer8[8] ) );
INV_X4 _u0_U19559  ( .A(1'b1), .ZN(_u0_pointer8[7] ) );
INV_X4 _u0_U19557  ( .A(1'b1), .ZN(_u0_pointer8[6] ) );
INV_X4 _u0_U19555  ( .A(1'b1), .ZN(_u0_pointer8[5] ) );
INV_X4 _u0_U19553  ( .A(1'b1), .ZN(_u0_pointer8[4] ) );
INV_X4 _u0_U19551  ( .A(1'b1), .ZN(_u0_pointer8[3] ) );
INV_X4 _u0_U19549  ( .A(1'b1), .ZN(_u0_pointer8[2] ) );
INV_X4 _u0_U19547  ( .A(1'b1), .ZN(_u0_pointer8[1] ) );
INV_X4 _u0_U19545  ( .A(1'b1), .ZN(_u0_pointer8[0] ) );
INV_X4 _u0_U19543  ( .A(1'b1), .ZN(_u0_pointer8_s[31] ) );
INV_X4 _u0_U19541  ( .A(1'b1), .ZN(_u0_pointer8_s[30] ) );
INV_X4 _u0_U19539  ( .A(1'b1), .ZN(_u0_pointer8_s[29] ) );
INV_X4 _u0_U19537  ( .A(1'b1), .ZN(_u0_pointer8_s[28] ) );
INV_X4 _u0_U19535  ( .A(1'b1), .ZN(_u0_pointer8_s[27] ) );
INV_X4 _u0_U19533  ( .A(1'b1), .ZN(_u0_pointer8_s[26] ) );
INV_X4 _u0_U19531  ( .A(1'b1), .ZN(_u0_pointer8_s[25] ) );
INV_X4 _u0_U19529  ( .A(1'b1), .ZN(_u0_pointer8_s[24] ) );
INV_X4 _u0_U19527  ( .A(1'b1), .ZN(_u0_pointer8_s[23] ) );
INV_X4 _u0_U19525  ( .A(1'b1), .ZN(_u0_pointer8_s[22] ) );
INV_X4 _u0_U19523  ( .A(1'b1), .ZN(_u0_pointer8_s[21] ) );
INV_X4 _u0_U19521  ( .A(1'b1), .ZN(_u0_pointer8_s[20] ) );
INV_X4 _u0_U19519  ( .A(1'b1), .ZN(_u0_pointer8_s[19] ) );
INV_X4 _u0_U19517  ( .A(1'b1), .ZN(_u0_pointer8_s[18] ) );
INV_X4 _u0_U19515  ( .A(1'b1), .ZN(_u0_pointer8_s[17] ) );
INV_X4 _u0_U19513  ( .A(1'b1), .ZN(_u0_pointer8_s[16] ) );
INV_X4 _u0_U19511  ( .A(1'b1), .ZN(_u0_pointer8_s[15] ) );
INV_X4 _u0_U19509  ( .A(1'b1), .ZN(_u0_pointer8_s[14] ) );
INV_X4 _u0_U19507  ( .A(1'b1), .ZN(_u0_pointer8_s[13] ) );
INV_X4 _u0_U19505  ( .A(1'b1), .ZN(_u0_pointer8_s[12] ) );
INV_X4 _u0_U19503  ( .A(1'b1), .ZN(_u0_pointer8_s[11] ) );
INV_X4 _u0_U19501  ( .A(1'b1), .ZN(_u0_pointer8_s[10] ) );
INV_X4 _u0_U19499  ( .A(1'b1), .ZN(_u0_pointer8_s[9] ) );
INV_X4 _u0_U19497  ( .A(1'b1), .ZN(_u0_pointer8_s[8] ) );
INV_X4 _u0_U19495  ( .A(1'b1), .ZN(_u0_pointer8_s[7] ) );
INV_X4 _u0_U19493  ( .A(1'b1), .ZN(_u0_pointer8_s[6] ) );
INV_X4 _u0_U19491  ( .A(1'b1), .ZN(_u0_pointer8_s[5] ) );
INV_X4 _u0_U19489  ( .A(1'b1), .ZN(_u0_pointer8_s[4] ) );
INV_X4 _u0_U19487  ( .A(1'b1), .ZN(_u0_pointer8_s[3] ) );
INV_X4 _u0_U19485  ( .A(1'b1), .ZN(_u0_pointer8_s[2] ) );
INV_X4 _u0_U19483  ( .A(1'b1), .ZN(_u0_pointer8_s[1] ) );
INV_X4 _u0_U19481  ( .A(1'b1), .ZN(_u0_pointer8_s[0] ) );
INV_X4 _u0_U19479  ( .A(1'b1), .ZN(_u0_ch8_csr[31] ) );
INV_X4 _u0_U19477  ( .A(1'b1), .ZN(_u0_ch8_csr[30] ) );
INV_X4 _u0_U19475  ( .A(1'b1), .ZN(_u0_ch8_csr[29] ) );
INV_X4 _u0_U19473  ( .A(1'b1), .ZN(_u0_ch8_csr[28] ) );
INV_X4 _u0_U19471  ( .A(1'b1), .ZN(_u0_ch8_csr[27] ) );
INV_X4 _u0_U19469  ( .A(1'b1), .ZN(_u0_ch8_csr[26] ) );
INV_X4 _u0_U19467  ( .A(1'b1), .ZN(_u0_ch8_csr[25] ) );
INV_X4 _u0_U19465  ( .A(1'b1), .ZN(_u0_ch8_csr[24] ) );
INV_X4 _u0_U19463  ( .A(1'b1), .ZN(_u0_ch8_csr[23] ) );
INV_X4 _u0_U19461  ( .A(1'b1), .ZN(_u0_ch8_csr[22] ) );
INV_X4 _u0_U19459  ( .A(1'b1), .ZN(_u0_ch8_csr[21] ) );
INV_X4 _u0_U19457  ( .A(1'b1), .ZN(_u0_ch8_csr[20] ) );
INV_X4 _u0_U19455  ( .A(1'b1), .ZN(_u0_ch8_csr[19] ) );
INV_X4 _u0_U19453  ( .A(1'b1), .ZN(_u0_ch8_csr[18] ) );
INV_X4 _u0_U19451  ( .A(1'b1), .ZN(_u0_ch8_csr[17] ) );
INV_X4 _u0_U19449  ( .A(1'b1), .ZN(_u0_ch8_csr[16] ) );
INV_X4 _u0_U19447  ( .A(1'b1), .ZN(_u0_ch8_csr[15] ) );
INV_X4 _u0_U19445  ( .A(1'b1), .ZN(_u0_ch8_csr[14] ) );
INV_X4 _u0_U19443  ( .A(1'b1), .ZN(_u0_ch8_csr[13] ) );
INV_X4 _u0_U19441  ( .A(1'b1), .ZN(_u0_ch8_csr[12] ) );
INV_X4 _u0_U19439  ( .A(1'b1), .ZN(_u0_ch8_csr[11] ) );
INV_X4 _u0_U19437  ( .A(1'b1), .ZN(_u0_ch8_csr[10] ) );
INV_X4 _u0_U19435  ( .A(1'b1), .ZN(_u0_ch8_csr[9] ) );
INV_X4 _u0_U19433  ( .A(1'b1), .ZN(_u0_ch8_csr[8] ) );
INV_X4 _u0_U19431  ( .A(1'b1), .ZN(_u0_ch8_csr[7] ) );
INV_X4 _u0_U19429  ( .A(1'b1), .ZN(_u0_ch8_csr[6] ) );
INV_X4 _u0_U19427  ( .A(1'b1), .ZN(_u0_ch8_csr[5] ) );
INV_X4 _u0_U19425  ( .A(1'b1), .ZN(_u0_ch8_csr[4] ) );
INV_X4 _u0_U19423  ( .A(1'b1), .ZN(_u0_ch8_csr[3] ) );
INV_X4 _u0_U19421  ( .A(1'b1), .ZN(_u0_ch8_csr[2] ) );
INV_X4 _u0_U19419  ( .A(1'b1), .ZN(_u0_ch8_csr[1] ) );
INV_X4 _u0_U19417  ( .A(1'b1), .ZN(_u0_ch8_csr[0] ) );
INV_X4 _u0_U19415  ( .A(1'b1), .ZN(_u0_ch8_txsz[31] ) );
INV_X4 _u0_U19413  ( .A(1'b1), .ZN(_u0_ch8_txsz[30] ) );
INV_X4 _u0_U19411  ( .A(1'b1), .ZN(_u0_ch8_txsz[29] ) );
INV_X4 _u0_U19409  ( .A(1'b1), .ZN(_u0_ch8_txsz[28] ) );
INV_X4 _u0_U19407  ( .A(1'b1), .ZN(_u0_ch8_txsz[27] ) );
INV_X4 _u0_U19405  ( .A(1'b1), .ZN(_u0_ch8_txsz[26] ) );
INV_X4 _u0_U19403  ( .A(1'b1), .ZN(_u0_ch8_txsz[25] ) );
INV_X4 _u0_U19401  ( .A(1'b1), .ZN(_u0_ch8_txsz[24] ) );
INV_X4 _u0_U19399  ( .A(1'b1), .ZN(_u0_ch8_txsz[23] ) );
INV_X4 _u0_U19397  ( .A(1'b1), .ZN(_u0_ch8_txsz[22] ) );
INV_X4 _u0_U19395  ( .A(1'b1), .ZN(_u0_ch8_txsz[21] ) );
INV_X4 _u0_U19393  ( .A(1'b1), .ZN(_u0_ch8_txsz[20] ) );
INV_X4 _u0_U19391  ( .A(1'b1), .ZN(_u0_ch8_txsz[19] ) );
INV_X4 _u0_U19389  ( .A(1'b1), .ZN(_u0_ch8_txsz[18] ) );
INV_X4 _u0_U19387  ( .A(1'b1), .ZN(_u0_ch8_txsz[17] ) );
INV_X4 _u0_U19385  ( .A(1'b1), .ZN(_u0_ch8_txsz[16] ) );
INV_X4 _u0_U19383  ( .A(1'b1), .ZN(_u0_ch8_txsz[15] ) );
INV_X4 _u0_U19381  ( .A(1'b1), .ZN(_u0_ch8_txsz[14] ) );
INV_X4 _u0_U19379  ( .A(1'b1), .ZN(_u0_ch8_txsz[13] ) );
INV_X4 _u0_U19377  ( .A(1'b1), .ZN(_u0_ch8_txsz[12] ) );
INV_X4 _u0_U19375  ( .A(1'b1), .ZN(_u0_ch8_txsz[11] ) );
INV_X4 _u0_U19373  ( .A(1'b1), .ZN(_u0_ch8_txsz[10] ) );
INV_X4 _u0_U19371  ( .A(1'b1), .ZN(_u0_ch8_txsz[9] ) );
INV_X4 _u0_U19369  ( .A(1'b1), .ZN(_u0_ch8_txsz[8] ) );
INV_X4 _u0_U19367  ( .A(1'b1), .ZN(_u0_ch8_txsz[7] ) );
INV_X4 _u0_U19365  ( .A(1'b1), .ZN(_u0_ch8_txsz[6] ) );
INV_X4 _u0_U19363  ( .A(1'b1), .ZN(_u0_ch8_txsz[5] ) );
INV_X4 _u0_U19361  ( .A(1'b1), .ZN(_u0_ch8_txsz[4] ) );
INV_X4 _u0_U19359  ( .A(1'b1), .ZN(_u0_ch8_txsz[3] ) );
INV_X4 _u0_U19357  ( .A(1'b1), .ZN(_u0_ch8_txsz[2] ) );
INV_X4 _u0_U19355  ( .A(1'b1), .ZN(_u0_ch8_txsz[1] ) );
INV_X4 _u0_U19353  ( .A(1'b1), .ZN(_u0_ch8_txsz[0] ) );
INV_X4 _u0_U19351  ( .A(1'b1), .ZN(_u0_ch8_adr0[31] ) );
INV_X4 _u0_U19349  ( .A(1'b1), .ZN(_u0_ch8_adr0[30] ) );
INV_X4 _u0_U19347  ( .A(1'b1), .ZN(_u0_ch8_adr0[29] ) );
INV_X4 _u0_U19345  ( .A(1'b1), .ZN(_u0_ch8_adr0[28] ) );
INV_X4 _u0_U19343  ( .A(1'b1), .ZN(_u0_ch8_adr0[27] ) );
INV_X4 _u0_U19341  ( .A(1'b1), .ZN(_u0_ch8_adr0[26] ) );
INV_X4 _u0_U19339  ( .A(1'b1), .ZN(_u0_ch8_adr0[25] ) );
INV_X4 _u0_U19337  ( .A(1'b1), .ZN(_u0_ch8_adr0[24] ) );
INV_X4 _u0_U19335  ( .A(1'b1), .ZN(_u0_ch8_adr0[23] ) );
INV_X4 _u0_U19333  ( .A(1'b1), .ZN(_u0_ch8_adr0[22] ) );
INV_X4 _u0_U19331  ( .A(1'b1), .ZN(_u0_ch8_adr0[21] ) );
INV_X4 _u0_U19329  ( .A(1'b1), .ZN(_u0_ch8_adr0[20] ) );
INV_X4 _u0_U19327  ( .A(1'b1), .ZN(_u0_ch8_adr0[19] ) );
INV_X4 _u0_U19325  ( .A(1'b1), .ZN(_u0_ch8_adr0[18] ) );
INV_X4 _u0_U19323  ( .A(1'b1), .ZN(_u0_ch8_adr0[17] ) );
INV_X4 _u0_U19321  ( .A(1'b1), .ZN(_u0_ch8_adr0[16] ) );
INV_X4 _u0_U19319  ( .A(1'b1), .ZN(_u0_ch8_adr0[15] ) );
INV_X4 _u0_U19317  ( .A(1'b1), .ZN(_u0_ch8_adr0[14] ) );
INV_X4 _u0_U19315  ( .A(1'b1), .ZN(_u0_ch8_adr0[13] ) );
INV_X4 _u0_U19313  ( .A(1'b1), .ZN(_u0_ch8_adr0[12] ) );
INV_X4 _u0_U19311  ( .A(1'b1), .ZN(_u0_ch8_adr0[11] ) );
INV_X4 _u0_U19309  ( .A(1'b1), .ZN(_u0_ch8_adr0[10] ) );
INV_X4 _u0_U19307  ( .A(1'b1), .ZN(_u0_ch8_adr0[9] ) );
INV_X4 _u0_U19305  ( .A(1'b1), .ZN(_u0_ch8_adr0[8] ) );
INV_X4 _u0_U19303  ( .A(1'b1), .ZN(_u0_ch8_adr0[7] ) );
INV_X4 _u0_U19301  ( .A(1'b1), .ZN(_u0_ch8_adr0[6] ) );
INV_X4 _u0_U19299  ( .A(1'b1), .ZN(_u0_ch8_adr0[5] ) );
INV_X4 _u0_U19297  ( .A(1'b1), .ZN(_u0_ch8_adr0[4] ) );
INV_X4 _u0_U19295  ( .A(1'b1), .ZN(_u0_ch8_adr0[3] ) );
INV_X4 _u0_U19293  ( .A(1'b1), .ZN(_u0_ch8_adr0[2] ) );
INV_X4 _u0_U19291  ( .A(1'b1), .ZN(_u0_ch8_adr0[1] ) );
INV_X4 _u0_U19289  ( .A(1'b1), .ZN(_u0_ch8_adr0[0] ) );
INV_X4 _u0_U19287  ( .A(1'b1), .ZN(_u0_ch8_adr1[31] ) );
INV_X4 _u0_U19285  ( .A(1'b1), .ZN(_u0_ch8_adr1[30] ) );
INV_X4 _u0_U19283  ( .A(1'b1), .ZN(_u0_ch8_adr1[29] ) );
INV_X4 _u0_U19281  ( .A(1'b1), .ZN(_u0_ch8_adr1[28] ) );
INV_X4 _u0_U19279  ( .A(1'b1), .ZN(_u0_ch8_adr1[27] ) );
INV_X4 _u0_U19277  ( .A(1'b1), .ZN(_u0_ch8_adr1[26] ) );
INV_X4 _u0_U19275  ( .A(1'b1), .ZN(_u0_ch8_adr1[25] ) );
INV_X4 _u0_U19273  ( .A(1'b1), .ZN(_u0_ch8_adr1[24] ) );
INV_X4 _u0_U19271  ( .A(1'b1), .ZN(_u0_ch8_adr1[23] ) );
INV_X4 _u0_U19269  ( .A(1'b1), .ZN(_u0_ch8_adr1[22] ) );
INV_X4 _u0_U19267  ( .A(1'b1), .ZN(_u0_ch8_adr1[21] ) );
INV_X4 _u0_U19265  ( .A(1'b1), .ZN(_u0_ch8_adr1[20] ) );
INV_X4 _u0_U19263  ( .A(1'b1), .ZN(_u0_ch8_adr1[19] ) );
INV_X4 _u0_U19261  ( .A(1'b1), .ZN(_u0_ch8_adr1[18] ) );
INV_X4 _u0_U19259  ( .A(1'b1), .ZN(_u0_ch8_adr1[17] ) );
INV_X4 _u0_U19257  ( .A(1'b1), .ZN(_u0_ch8_adr1[16] ) );
INV_X4 _u0_U19255  ( .A(1'b1), .ZN(_u0_ch8_adr1[15] ) );
INV_X4 _u0_U19253  ( .A(1'b1), .ZN(_u0_ch8_adr1[14] ) );
INV_X4 _u0_U19251  ( .A(1'b1), .ZN(_u0_ch8_adr1[13] ) );
INV_X4 _u0_U19249  ( .A(1'b1), .ZN(_u0_ch8_adr1[12] ) );
INV_X4 _u0_U19247  ( .A(1'b1), .ZN(_u0_ch8_adr1[11] ) );
INV_X4 _u0_U19245  ( .A(1'b1), .ZN(_u0_ch8_adr1[10] ) );
INV_X4 _u0_U19243  ( .A(1'b1), .ZN(_u0_ch8_adr1[9] ) );
INV_X4 _u0_U19241  ( .A(1'b1), .ZN(_u0_ch8_adr1[8] ) );
INV_X4 _u0_U19239  ( .A(1'b1), .ZN(_u0_ch8_adr1[7] ) );
INV_X4 _u0_U19237  ( .A(1'b1), .ZN(_u0_ch8_adr1[6] ) );
INV_X4 _u0_U19235  ( .A(1'b1), .ZN(_u0_ch8_adr1[5] ) );
INV_X4 _u0_U19233  ( .A(1'b1), .ZN(_u0_ch8_adr1[4] ) );
INV_X4 _u0_U19231  ( .A(1'b1), .ZN(_u0_ch8_adr1[3] ) );
INV_X4 _u0_U19229  ( .A(1'b1), .ZN(_u0_ch8_adr1[2] ) );
INV_X4 _u0_U19227  ( .A(1'b1), .ZN(_u0_ch8_adr1[1] ) );
INV_X4 _u0_U19225  ( .A(1'b1), .ZN(_u0_ch8_adr1[0] ) );
INV_X4 _u0_U19223  ( .A(1'b0), .ZN(_u0_ch8_am0[31] ) );
INV_X4 _u0_U19221  ( .A(1'b0), .ZN(_u0_ch8_am0[30] ) );
INV_X4 _u0_U19219  ( .A(1'b0), .ZN(_u0_ch8_am0[29] ) );
INV_X4 _u0_U19217  ( .A(1'b0), .ZN(_u0_ch8_am0[28] ) );
INV_X4 _u0_U19215  ( .A(1'b0), .ZN(_u0_ch8_am0[27] ) );
INV_X4 _u0_U19213  ( .A(1'b0), .ZN(_u0_ch8_am0[26] ) );
INV_X4 _u0_U19211  ( .A(1'b0), .ZN(_u0_ch8_am0[25] ) );
INV_X4 _u0_U19209  ( .A(1'b0), .ZN(_u0_ch8_am0[24] ) );
INV_X4 _u0_U19207  ( .A(1'b0), .ZN(_u0_ch8_am0[23] ) );
INV_X4 _u0_U19205  ( .A(1'b0), .ZN(_u0_ch8_am0[22] ) );
INV_X4 _u0_U19203  ( .A(1'b0), .ZN(_u0_ch8_am0[21] ) );
INV_X4 _u0_U19201  ( .A(1'b0), .ZN(_u0_ch8_am0[20] ) );
INV_X4 _u0_U19199  ( .A(1'b0), .ZN(_u0_ch8_am0[19] ) );
INV_X4 _u0_U19197  ( .A(1'b0), .ZN(_u0_ch8_am0[18] ) );
INV_X4 _u0_U19195  ( .A(1'b0), .ZN(_u0_ch8_am0[17] ) );
INV_X4 _u0_U19193  ( .A(1'b0), .ZN(_u0_ch8_am0[16] ) );
INV_X4 _u0_U19191  ( .A(1'b0), .ZN(_u0_ch8_am0[15] ) );
INV_X4 _u0_U19189  ( .A(1'b0), .ZN(_u0_ch8_am0[14] ) );
INV_X4 _u0_U19187  ( .A(1'b0), .ZN(_u0_ch8_am0[13] ) );
INV_X4 _u0_U19185  ( .A(1'b0), .ZN(_u0_ch8_am0[12] ) );
INV_X4 _u0_U19183  ( .A(1'b0), .ZN(_u0_ch8_am0[11] ) );
INV_X4 _u0_U19181  ( .A(1'b0), .ZN(_u0_ch8_am0[10] ) );
INV_X4 _u0_U19179  ( .A(1'b0), .ZN(_u0_ch8_am0[9] ) );
INV_X4 _u0_U19177  ( .A(1'b0), .ZN(_u0_ch8_am0[8] ) );
INV_X4 _u0_U19175  ( .A(1'b0), .ZN(_u0_ch8_am0[7] ) );
INV_X4 _u0_U19173  ( .A(1'b0), .ZN(_u0_ch8_am0[6] ) );
INV_X4 _u0_U19171  ( .A(1'b0), .ZN(_u0_ch8_am0[5] ) );
INV_X4 _u0_U19169  ( .A(1'b0), .ZN(_u0_ch8_am0[4] ) );
INV_X4 _u0_U19167  ( .A(1'b1), .ZN(_u0_ch8_am0[3] ) );
INV_X4 _u0_U19165  ( .A(1'b1), .ZN(_u0_ch8_am0[2] ) );
INV_X4 _u0_U19163  ( .A(1'b1), .ZN(_u0_ch8_am0[1] ) );
INV_X4 _u0_U19161  ( .A(1'b1), .ZN(_u0_ch8_am0[0] ) );
INV_X4 _u0_U19159  ( .A(1'b0), .ZN(_u0_ch8_am1[31] ) );
INV_X4 _u0_U19157  ( .A(1'b0), .ZN(_u0_ch8_am1[30] ) );
INV_X4 _u0_U19155  ( .A(1'b0), .ZN(_u0_ch8_am1[29] ) );
INV_X4 _u0_U19153  ( .A(1'b0), .ZN(_u0_ch8_am1[28] ) );
INV_X4 _u0_U19151  ( .A(1'b0), .ZN(_u0_ch8_am1[27] ) );
INV_X4 _u0_U19149  ( .A(1'b0), .ZN(_u0_ch8_am1[26] ) );
INV_X4 _u0_U19147  ( .A(1'b0), .ZN(_u0_ch8_am1[25] ) );
INV_X4 _u0_U19145  ( .A(1'b0), .ZN(_u0_ch8_am1[24] ) );
INV_X4 _u0_U19143  ( .A(1'b0), .ZN(_u0_ch8_am1[23] ) );
INV_X4 _u0_U19141  ( .A(1'b0), .ZN(_u0_ch8_am1[22] ) );
INV_X4 _u0_U19139  ( .A(1'b0), .ZN(_u0_ch8_am1[21] ) );
INV_X4 _u0_U19137  ( .A(1'b0), .ZN(_u0_ch8_am1[20] ) );
INV_X4 _u0_U19135  ( .A(1'b0), .ZN(_u0_ch8_am1[19] ) );
INV_X4 _u0_U19133  ( .A(1'b0), .ZN(_u0_ch8_am1[18] ) );
INV_X4 _u0_U19131  ( .A(1'b0), .ZN(_u0_ch8_am1[17] ) );
INV_X4 _u0_U19129  ( .A(1'b0), .ZN(_u0_ch8_am1[16] ) );
INV_X4 _u0_U19127  ( .A(1'b0), .ZN(_u0_ch8_am1[15] ) );
INV_X4 _u0_U19125  ( .A(1'b0), .ZN(_u0_ch8_am1[14] ) );
INV_X4 _u0_U19123  ( .A(1'b0), .ZN(_u0_ch8_am1[13] ) );
INV_X4 _u0_U19121  ( .A(1'b0), .ZN(_u0_ch8_am1[12] ) );
INV_X4 _u0_U19119  ( .A(1'b0), .ZN(_u0_ch8_am1[11] ) );
INV_X4 _u0_U19117  ( .A(1'b0), .ZN(_u0_ch8_am1[10] ) );
INV_X4 _u0_U19115  ( .A(1'b0), .ZN(_u0_ch8_am1[9] ) );
INV_X4 _u0_U19113  ( .A(1'b0), .ZN(_u0_ch8_am1[8] ) );
INV_X4 _u0_U19111  ( .A(1'b0), .ZN(_u0_ch8_am1[7] ) );
INV_X4 _u0_U19109  ( .A(1'b0), .ZN(_u0_ch8_am1[6] ) );
INV_X4 _u0_U19107  ( .A(1'b0), .ZN(_u0_ch8_am1[5] ) );
INV_X4 _u0_U19105  ( .A(1'b0), .ZN(_u0_ch8_am1[4] ) );
INV_X4 _u0_U19103  ( .A(1'b1), .ZN(_u0_ch8_am1[3] ) );
INV_X4 _u0_U19101  ( .A(1'b1), .ZN(_u0_ch8_am1[2] ) );
INV_X4 _u0_U19099  ( .A(1'b1), .ZN(_u0_ch8_am1[1] ) );
INV_X4 _u0_U19097  ( .A(1'b1), .ZN(_u0_ch8_am1[0] ) );
INV_X4 _u0_U19095  ( .A(1'b1), .ZN(_u0_pointer9[31] ) );
INV_X4 _u0_U19093  ( .A(1'b1), .ZN(_u0_pointer9[30] ) );
INV_X4 _u0_U19091  ( .A(1'b1), .ZN(_u0_pointer9[29] ) );
INV_X4 _u0_U19089  ( .A(1'b1), .ZN(_u0_pointer9[28] ) );
INV_X4 _u0_U19087  ( .A(1'b1), .ZN(_u0_pointer9[27] ) );
INV_X4 _u0_U19085  ( .A(1'b1), .ZN(_u0_pointer9[26] ) );
INV_X4 _u0_U19083  ( .A(1'b1), .ZN(_u0_pointer9[25] ) );
INV_X4 _u0_U19081  ( .A(1'b1), .ZN(_u0_pointer9[24] ) );
INV_X4 _u0_U19079  ( .A(1'b1), .ZN(_u0_pointer9[23] ) );
INV_X4 _u0_U19077  ( .A(1'b1), .ZN(_u0_pointer9[22] ) );
INV_X4 _u0_U19075  ( .A(1'b1), .ZN(_u0_pointer9[21] ) );
INV_X4 _u0_U19073  ( .A(1'b1), .ZN(_u0_pointer9[20] ) );
INV_X4 _u0_U19071  ( .A(1'b1), .ZN(_u0_pointer9[19] ) );
INV_X4 _u0_U19069  ( .A(1'b1), .ZN(_u0_pointer9[18] ) );
INV_X4 _u0_U19067  ( .A(1'b1), .ZN(_u0_pointer9[17] ) );
INV_X4 _u0_U19065  ( .A(1'b1), .ZN(_u0_pointer9[16] ) );
INV_X4 _u0_U19063  ( .A(1'b1), .ZN(_u0_pointer9[15] ) );
INV_X4 _u0_U19061  ( .A(1'b1), .ZN(_u0_pointer9[14] ) );
INV_X4 _u0_U19059  ( .A(1'b1), .ZN(_u0_pointer9[13] ) );
INV_X4 _u0_U19057  ( .A(1'b1), .ZN(_u0_pointer9[12] ) );
INV_X4 _u0_U19055  ( .A(1'b1), .ZN(_u0_pointer9[11] ) );
INV_X4 _u0_U19053  ( .A(1'b1), .ZN(_u0_pointer9[10] ) );
INV_X4 _u0_U19051  ( .A(1'b1), .ZN(_u0_pointer9[9] ) );
INV_X4 _u0_U19049  ( .A(1'b1), .ZN(_u0_pointer9[8] ) );
INV_X4 _u0_U19047  ( .A(1'b1), .ZN(_u0_pointer9[7] ) );
INV_X4 _u0_U19045  ( .A(1'b1), .ZN(_u0_pointer9[6] ) );
INV_X4 _u0_U19043  ( .A(1'b1), .ZN(_u0_pointer9[5] ) );
INV_X4 _u0_U19041  ( .A(1'b1), .ZN(_u0_pointer9[4] ) );
INV_X4 _u0_U19039  ( .A(1'b1), .ZN(_u0_pointer9[3] ) );
INV_X4 _u0_U19037  ( .A(1'b1), .ZN(_u0_pointer9[2] ) );
INV_X4 _u0_U19035  ( .A(1'b1), .ZN(_u0_pointer9[1] ) );
INV_X4 _u0_U19033  ( .A(1'b1), .ZN(_u0_pointer9[0] ) );
INV_X4 _u0_U19031  ( .A(1'b1), .ZN(_u0_pointer9_s[31] ) );
INV_X4 _u0_U19029  ( .A(1'b1), .ZN(_u0_pointer9_s[30] ) );
INV_X4 _u0_U19027  ( .A(1'b1), .ZN(_u0_pointer9_s[29] ) );
INV_X4 _u0_U19025  ( .A(1'b1), .ZN(_u0_pointer9_s[28] ) );
INV_X4 _u0_U19023  ( .A(1'b1), .ZN(_u0_pointer9_s[27] ) );
INV_X4 _u0_U19021  ( .A(1'b1), .ZN(_u0_pointer9_s[26] ) );
INV_X4 _u0_U19019  ( .A(1'b1), .ZN(_u0_pointer9_s[25] ) );
INV_X4 _u0_U19017  ( .A(1'b1), .ZN(_u0_pointer9_s[24] ) );
INV_X4 _u0_U19015  ( .A(1'b1), .ZN(_u0_pointer9_s[23] ) );
INV_X4 _u0_U19013  ( .A(1'b1), .ZN(_u0_pointer9_s[22] ) );
INV_X4 _u0_U19011  ( .A(1'b1), .ZN(_u0_pointer9_s[21] ) );
INV_X4 _u0_U19009  ( .A(1'b1), .ZN(_u0_pointer9_s[20] ) );
INV_X4 _u0_U19007  ( .A(1'b1), .ZN(_u0_pointer9_s[19] ) );
INV_X4 _u0_U19005  ( .A(1'b1), .ZN(_u0_pointer9_s[18] ) );
INV_X4 _u0_U19003  ( .A(1'b1), .ZN(_u0_pointer9_s[17] ) );
INV_X4 _u0_U19001  ( .A(1'b1), .ZN(_u0_pointer9_s[16] ) );
INV_X4 _u0_U18999  ( .A(1'b1), .ZN(_u0_pointer9_s[15] ) );
INV_X4 _u0_U18997  ( .A(1'b1), .ZN(_u0_pointer9_s[14] ) );
INV_X4 _u0_U18995  ( .A(1'b1), .ZN(_u0_pointer9_s[13] ) );
INV_X4 _u0_U18993  ( .A(1'b1), .ZN(_u0_pointer9_s[12] ) );
INV_X4 _u0_U18991  ( .A(1'b1), .ZN(_u0_pointer9_s[11] ) );
INV_X4 _u0_U18989  ( .A(1'b1), .ZN(_u0_pointer9_s[10] ) );
INV_X4 _u0_U18987  ( .A(1'b1), .ZN(_u0_pointer9_s[9] ) );
INV_X4 _u0_U18985  ( .A(1'b1), .ZN(_u0_pointer9_s[8] ) );
INV_X4 _u0_U18983  ( .A(1'b1), .ZN(_u0_pointer9_s[7] ) );
INV_X4 _u0_U18981  ( .A(1'b1), .ZN(_u0_pointer9_s[6] ) );
INV_X4 _u0_U18979  ( .A(1'b1), .ZN(_u0_pointer9_s[5] ) );
INV_X4 _u0_U18977  ( .A(1'b1), .ZN(_u0_pointer9_s[4] ) );
INV_X4 _u0_U18975  ( .A(1'b1), .ZN(_u0_pointer9_s[3] ) );
INV_X4 _u0_U18973  ( .A(1'b1), .ZN(_u0_pointer9_s[2] ) );
INV_X4 _u0_U18971  ( .A(1'b1), .ZN(_u0_pointer9_s[1] ) );
INV_X4 _u0_U18969  ( .A(1'b1), .ZN(_u0_pointer9_s[0] ) );
INV_X4 _u0_U18967  ( .A(1'b1), .ZN(_u0_ch9_csr[31] ) );
INV_X4 _u0_U18965  ( .A(1'b1), .ZN(_u0_ch9_csr[30] ) );
INV_X4 _u0_U18963  ( .A(1'b1), .ZN(_u0_ch9_csr[29] ) );
INV_X4 _u0_U18961  ( .A(1'b1), .ZN(_u0_ch9_csr[28] ) );
INV_X4 _u0_U18959  ( .A(1'b1), .ZN(_u0_ch9_csr[27] ) );
INV_X4 _u0_U18957  ( .A(1'b1), .ZN(_u0_ch9_csr[26] ) );
INV_X4 _u0_U18955  ( .A(1'b1), .ZN(_u0_ch9_csr[25] ) );
INV_X4 _u0_U18953  ( .A(1'b1), .ZN(_u0_ch9_csr[24] ) );
INV_X4 _u0_U18951  ( .A(1'b1), .ZN(_u0_ch9_csr[23] ) );
INV_X4 _u0_U18949  ( .A(1'b1), .ZN(_u0_ch9_csr[22] ) );
INV_X4 _u0_U18947  ( .A(1'b1), .ZN(_u0_ch9_csr[21] ) );
INV_X4 _u0_U18945  ( .A(1'b1), .ZN(_u0_ch9_csr[20] ) );
INV_X4 _u0_U18943  ( .A(1'b1), .ZN(_u0_ch9_csr[19] ) );
INV_X4 _u0_U18941  ( .A(1'b1), .ZN(_u0_ch9_csr[18] ) );
INV_X4 _u0_U18939  ( .A(1'b1), .ZN(_u0_ch9_csr[17] ) );
INV_X4 _u0_U18937  ( .A(1'b1), .ZN(_u0_ch9_csr[16] ) );
INV_X4 _u0_U18935  ( .A(1'b1), .ZN(_u0_ch9_csr[15] ) );
INV_X4 _u0_U18933  ( .A(1'b1), .ZN(_u0_ch9_csr[14] ) );
INV_X4 _u0_U18931  ( .A(1'b1), .ZN(_u0_ch9_csr[13] ) );
INV_X4 _u0_U18929  ( .A(1'b1), .ZN(_u0_ch9_csr[12] ) );
INV_X4 _u0_U18927  ( .A(1'b1), .ZN(_u0_ch9_csr[11] ) );
INV_X4 _u0_U18925  ( .A(1'b1), .ZN(_u0_ch9_csr[10] ) );
INV_X4 _u0_U18923  ( .A(1'b1), .ZN(_u0_ch9_csr[9] ) );
INV_X4 _u0_U18921  ( .A(1'b1), .ZN(_u0_ch9_csr[8] ) );
INV_X4 _u0_U18919  ( .A(1'b1), .ZN(_u0_ch9_csr[7] ) );
INV_X4 _u0_U18917  ( .A(1'b1), .ZN(_u0_ch9_csr[6] ) );
INV_X4 _u0_U18915  ( .A(1'b1), .ZN(_u0_ch9_csr[5] ) );
INV_X4 _u0_U18913  ( .A(1'b1), .ZN(_u0_ch9_csr[4] ) );
INV_X4 _u0_U18911  ( .A(1'b1), .ZN(_u0_ch9_csr[3] ) );
INV_X4 _u0_U18909  ( .A(1'b1), .ZN(_u0_ch9_csr[2] ) );
INV_X4 _u0_U18907  ( .A(1'b1), .ZN(_u0_ch9_csr[1] ) );
INV_X4 _u0_U18905  ( .A(1'b1), .ZN(_u0_ch9_csr[0] ) );
INV_X4 _u0_U18903  ( .A(1'b1), .ZN(_u0_ch9_txsz[31] ) );
INV_X4 _u0_U18901  ( .A(1'b1), .ZN(_u0_ch9_txsz[30] ) );
INV_X4 _u0_U18899  ( .A(1'b1), .ZN(_u0_ch9_txsz[29] ) );
INV_X4 _u0_U18897  ( .A(1'b1), .ZN(_u0_ch9_txsz[28] ) );
INV_X4 _u0_U18895  ( .A(1'b1), .ZN(_u0_ch9_txsz[27] ) );
INV_X4 _u0_U18893  ( .A(1'b1), .ZN(_u0_ch9_txsz[26] ) );
INV_X4 _u0_U18891  ( .A(1'b1), .ZN(_u0_ch9_txsz[25] ) );
INV_X4 _u0_U18889  ( .A(1'b1), .ZN(_u0_ch9_txsz[24] ) );
INV_X4 _u0_U18887  ( .A(1'b1), .ZN(_u0_ch9_txsz[23] ) );
INV_X4 _u0_U18885  ( .A(1'b1), .ZN(_u0_ch9_txsz[22] ) );
INV_X4 _u0_U18883  ( .A(1'b1), .ZN(_u0_ch9_txsz[21] ) );
INV_X4 _u0_U18881  ( .A(1'b1), .ZN(_u0_ch9_txsz[20] ) );
INV_X4 _u0_U18879  ( .A(1'b1), .ZN(_u0_ch9_txsz[19] ) );
INV_X4 _u0_U18877  ( .A(1'b1), .ZN(_u0_ch9_txsz[18] ) );
INV_X4 _u0_U18875  ( .A(1'b1), .ZN(_u0_ch9_txsz[17] ) );
INV_X4 _u0_U18873  ( .A(1'b1), .ZN(_u0_ch9_txsz[16] ) );
INV_X4 _u0_U18871  ( .A(1'b1), .ZN(_u0_ch9_txsz[15] ) );
INV_X4 _u0_U18869  ( .A(1'b1), .ZN(_u0_ch9_txsz[14] ) );
INV_X4 _u0_U18867  ( .A(1'b1), .ZN(_u0_ch9_txsz[13] ) );
INV_X4 _u0_U18865  ( .A(1'b1), .ZN(_u0_ch9_txsz[12] ) );
INV_X4 _u0_U18863  ( .A(1'b1), .ZN(_u0_ch9_txsz[11] ) );
INV_X4 _u0_U18861  ( .A(1'b1), .ZN(_u0_ch9_txsz[10] ) );
INV_X4 _u0_U18859  ( .A(1'b1), .ZN(_u0_ch9_txsz[9] ) );
INV_X4 _u0_U18857  ( .A(1'b1), .ZN(_u0_ch9_txsz[8] ) );
INV_X4 _u0_U18855  ( .A(1'b1), .ZN(_u0_ch9_txsz[7] ) );
INV_X4 _u0_U18853  ( .A(1'b1), .ZN(_u0_ch9_txsz[6] ) );
INV_X4 _u0_U18851  ( .A(1'b1), .ZN(_u0_ch9_txsz[5] ) );
INV_X4 _u0_U18849  ( .A(1'b1), .ZN(_u0_ch9_txsz[4] ) );
INV_X4 _u0_U18847  ( .A(1'b1), .ZN(_u0_ch9_txsz[3] ) );
INV_X4 _u0_U18845  ( .A(1'b1), .ZN(_u0_ch9_txsz[2] ) );
INV_X4 _u0_U18843  ( .A(1'b1), .ZN(_u0_ch9_txsz[1] ) );
INV_X4 _u0_U18841  ( .A(1'b1), .ZN(_u0_ch9_txsz[0] ) );
INV_X4 _u0_U18839  ( .A(1'b1), .ZN(_u0_ch9_adr0[31] ) );
INV_X4 _u0_U18837  ( .A(1'b1), .ZN(_u0_ch9_adr0[30] ) );
INV_X4 _u0_U18835  ( .A(1'b1), .ZN(_u0_ch9_adr0[29] ) );
INV_X4 _u0_U18833  ( .A(1'b1), .ZN(_u0_ch9_adr0[28] ) );
INV_X4 _u0_U18831  ( .A(1'b1), .ZN(_u0_ch9_adr0[27] ) );
INV_X4 _u0_U18829  ( .A(1'b1), .ZN(_u0_ch9_adr0[26] ) );
INV_X4 _u0_U18827  ( .A(1'b1), .ZN(_u0_ch9_adr0[25] ) );
INV_X4 _u0_U18825  ( .A(1'b1), .ZN(_u0_ch9_adr0[24] ) );
INV_X4 _u0_U18823  ( .A(1'b1), .ZN(_u0_ch9_adr0[23] ) );
INV_X4 _u0_U18821  ( .A(1'b1), .ZN(_u0_ch9_adr0[22] ) );
INV_X4 _u0_U18819  ( .A(1'b1), .ZN(_u0_ch9_adr0[21] ) );
INV_X4 _u0_U18817  ( .A(1'b1), .ZN(_u0_ch9_adr0[20] ) );
INV_X4 _u0_U18815  ( .A(1'b1), .ZN(_u0_ch9_adr0[19] ) );
INV_X4 _u0_U18813  ( .A(1'b1), .ZN(_u0_ch9_adr0[18] ) );
INV_X4 _u0_U18811  ( .A(1'b1), .ZN(_u0_ch9_adr0[17] ) );
INV_X4 _u0_U18809  ( .A(1'b1), .ZN(_u0_ch9_adr0[16] ) );
INV_X4 _u0_U18807  ( .A(1'b1), .ZN(_u0_ch9_adr0[15] ) );
INV_X4 _u0_U18805  ( .A(1'b1), .ZN(_u0_ch9_adr0[14] ) );
INV_X4 _u0_U18803  ( .A(1'b1), .ZN(_u0_ch9_adr0[13] ) );
INV_X4 _u0_U18801  ( .A(1'b1), .ZN(_u0_ch9_adr0[12] ) );
INV_X4 _u0_U18799  ( .A(1'b1), .ZN(_u0_ch9_adr0[11] ) );
INV_X4 _u0_U18797  ( .A(1'b1), .ZN(_u0_ch9_adr0[10] ) );
INV_X4 _u0_U18795  ( .A(1'b1), .ZN(_u0_ch9_adr0[9] ) );
INV_X4 _u0_U18793  ( .A(1'b1), .ZN(_u0_ch9_adr0[8] ) );
INV_X4 _u0_U18791  ( .A(1'b1), .ZN(_u0_ch9_adr0[7] ) );
INV_X4 _u0_U18789  ( .A(1'b1), .ZN(_u0_ch9_adr0[6] ) );
INV_X4 _u0_U18787  ( .A(1'b1), .ZN(_u0_ch9_adr0[5] ) );
INV_X4 _u0_U18785  ( .A(1'b1), .ZN(_u0_ch9_adr0[4] ) );
INV_X4 _u0_U18783  ( .A(1'b1), .ZN(_u0_ch9_adr0[3] ) );
INV_X4 _u0_U18781  ( .A(1'b1), .ZN(_u0_ch9_adr0[2] ) );
INV_X4 _u0_U18779  ( .A(1'b1), .ZN(_u0_ch9_adr0[1] ) );
INV_X4 _u0_U18777  ( .A(1'b1), .ZN(_u0_ch9_adr0[0] ) );
INV_X4 _u0_U18775  ( .A(1'b1), .ZN(_u0_ch9_adr1[31] ) );
INV_X4 _u0_U18773  ( .A(1'b1), .ZN(_u0_ch9_adr1[30] ) );
INV_X4 _u0_U18771  ( .A(1'b1), .ZN(_u0_ch9_adr1[29] ) );
INV_X4 _u0_U18769  ( .A(1'b1), .ZN(_u0_ch9_adr1[28] ) );
INV_X4 _u0_U18767  ( .A(1'b1), .ZN(_u0_ch9_adr1[27] ) );
INV_X4 _u0_U18765  ( .A(1'b1), .ZN(_u0_ch9_adr1[26] ) );
INV_X4 _u0_U18763  ( .A(1'b1), .ZN(_u0_ch9_adr1[25] ) );
INV_X4 _u0_U18761  ( .A(1'b1), .ZN(_u0_ch9_adr1[24] ) );
INV_X4 _u0_U18759  ( .A(1'b1), .ZN(_u0_ch9_adr1[23] ) );
INV_X4 _u0_U18757  ( .A(1'b1), .ZN(_u0_ch9_adr1[22] ) );
INV_X4 _u0_U18755  ( .A(1'b1), .ZN(_u0_ch9_adr1[21] ) );
INV_X4 _u0_U18753  ( .A(1'b1), .ZN(_u0_ch9_adr1[20] ) );
INV_X4 _u0_U18751  ( .A(1'b1), .ZN(_u0_ch9_adr1[19] ) );
INV_X4 _u0_U18749  ( .A(1'b1), .ZN(_u0_ch9_adr1[18] ) );
INV_X4 _u0_U18747  ( .A(1'b1), .ZN(_u0_ch9_adr1[17] ) );
INV_X4 _u0_U18745  ( .A(1'b1), .ZN(_u0_ch9_adr1[16] ) );
INV_X4 _u0_U18743  ( .A(1'b1), .ZN(_u0_ch9_adr1[15] ) );
INV_X4 _u0_U18741  ( .A(1'b1), .ZN(_u0_ch9_adr1[14] ) );
INV_X4 _u0_U18739  ( .A(1'b1), .ZN(_u0_ch9_adr1[13] ) );
INV_X4 _u0_U18737  ( .A(1'b1), .ZN(_u0_ch9_adr1[12] ) );
INV_X4 _u0_U18735  ( .A(1'b1), .ZN(_u0_ch9_adr1[11] ) );
INV_X4 _u0_U18733  ( .A(1'b1), .ZN(_u0_ch9_adr1[10] ) );
INV_X4 _u0_U18731  ( .A(1'b1), .ZN(_u0_ch9_adr1[9] ) );
INV_X4 _u0_U18729  ( .A(1'b1), .ZN(_u0_ch9_adr1[8] ) );
INV_X4 _u0_U18727  ( .A(1'b1), .ZN(_u0_ch9_adr1[7] ) );
INV_X4 _u0_U18725  ( .A(1'b1), .ZN(_u0_ch9_adr1[6] ) );
INV_X4 _u0_U18723  ( .A(1'b1), .ZN(_u0_ch9_adr1[5] ) );
INV_X4 _u0_U18721  ( .A(1'b1), .ZN(_u0_ch9_adr1[4] ) );
INV_X4 _u0_U18719  ( .A(1'b1), .ZN(_u0_ch9_adr1[3] ) );
INV_X4 _u0_U18717  ( .A(1'b1), .ZN(_u0_ch9_adr1[2] ) );
INV_X4 _u0_U18715  ( .A(1'b1), .ZN(_u0_ch9_adr1[1] ) );
INV_X4 _u0_U18713  ( .A(1'b1), .ZN(_u0_ch9_adr1[0] ) );
INV_X4 _u0_U18711  ( .A(1'b0), .ZN(_u0_ch9_am0[31] ) );
INV_X4 _u0_U18709  ( .A(1'b0), .ZN(_u0_ch9_am0[30] ) );
INV_X4 _u0_U18707  ( .A(1'b0), .ZN(_u0_ch9_am0[29] ) );
INV_X4 _u0_U18705  ( .A(1'b0), .ZN(_u0_ch9_am0[28] ) );
INV_X4 _u0_U18703  ( .A(1'b0), .ZN(_u0_ch9_am0[27] ) );
INV_X4 _u0_U18701  ( .A(1'b0), .ZN(_u0_ch9_am0[26] ) );
INV_X4 _u0_U18699  ( .A(1'b0), .ZN(_u0_ch9_am0[25] ) );
INV_X4 _u0_U18697  ( .A(1'b0), .ZN(_u0_ch9_am0[24] ) );
INV_X4 _u0_U18695  ( .A(1'b0), .ZN(_u0_ch9_am0[23] ) );
INV_X4 _u0_U18693  ( .A(1'b0), .ZN(_u0_ch9_am0[22] ) );
INV_X4 _u0_U18691  ( .A(1'b0), .ZN(_u0_ch9_am0[21] ) );
INV_X4 _u0_U18689  ( .A(1'b0), .ZN(_u0_ch9_am0[20] ) );
INV_X4 _u0_U18687  ( .A(1'b0), .ZN(_u0_ch9_am0[19] ) );
INV_X4 _u0_U18685  ( .A(1'b0), .ZN(_u0_ch9_am0[18] ) );
INV_X4 _u0_U18683  ( .A(1'b0), .ZN(_u0_ch9_am0[17] ) );
INV_X4 _u0_U18681  ( .A(1'b0), .ZN(_u0_ch9_am0[16] ) );
INV_X4 _u0_U18679  ( .A(1'b0), .ZN(_u0_ch9_am0[15] ) );
INV_X4 _u0_U18677  ( .A(1'b0), .ZN(_u0_ch9_am0[14] ) );
INV_X4 _u0_U18675  ( .A(1'b0), .ZN(_u0_ch9_am0[13] ) );
INV_X4 _u0_U18673  ( .A(1'b0), .ZN(_u0_ch9_am0[12] ) );
INV_X4 _u0_U18671  ( .A(1'b0), .ZN(_u0_ch9_am0[11] ) );
INV_X4 _u0_U18669  ( .A(1'b0), .ZN(_u0_ch9_am0[10] ) );
INV_X4 _u0_U18667  ( .A(1'b0), .ZN(_u0_ch9_am0[9] ) );
INV_X4 _u0_U18665  ( .A(1'b0), .ZN(_u0_ch9_am0[8] ) );
INV_X4 _u0_U18663  ( .A(1'b0), .ZN(_u0_ch9_am0[7] ) );
INV_X4 _u0_U18661  ( .A(1'b0), .ZN(_u0_ch9_am0[6] ) );
INV_X4 _u0_U18659  ( .A(1'b0), .ZN(_u0_ch9_am0[5] ) );
INV_X4 _u0_U18657  ( .A(1'b0), .ZN(_u0_ch9_am0[4] ) );
INV_X4 _u0_U18655  ( .A(1'b1), .ZN(_u0_ch9_am0[3] ) );
INV_X4 _u0_U18653  ( .A(1'b1), .ZN(_u0_ch9_am0[2] ) );
INV_X4 _u0_U18651  ( .A(1'b1), .ZN(_u0_ch9_am0[1] ) );
INV_X4 _u0_U18649  ( .A(1'b1), .ZN(_u0_ch9_am0[0] ) );
INV_X4 _u0_U18647  ( .A(1'b0), .ZN(_u0_ch9_am1[31] ) );
INV_X4 _u0_U18645  ( .A(1'b0), .ZN(_u0_ch9_am1[30] ) );
INV_X4 _u0_U18643  ( .A(1'b0), .ZN(_u0_ch9_am1[29] ) );
INV_X4 _u0_U18641  ( .A(1'b0), .ZN(_u0_ch9_am1[28] ) );
INV_X4 _u0_U18639  ( .A(1'b0), .ZN(_u0_ch9_am1[27] ) );
INV_X4 _u0_U18637  ( .A(1'b0), .ZN(_u0_ch9_am1[26] ) );
INV_X4 _u0_U18635  ( .A(1'b0), .ZN(_u0_ch9_am1[25] ) );
INV_X4 _u0_U18633  ( .A(1'b0), .ZN(_u0_ch9_am1[24] ) );
INV_X4 _u0_U18631  ( .A(1'b0), .ZN(_u0_ch9_am1[23] ) );
INV_X4 _u0_U18629  ( .A(1'b0), .ZN(_u0_ch9_am1[22] ) );
INV_X4 _u0_U18627  ( .A(1'b0), .ZN(_u0_ch9_am1[21] ) );
INV_X4 _u0_U18625  ( .A(1'b0), .ZN(_u0_ch9_am1[20] ) );
INV_X4 _u0_U18623  ( .A(1'b0), .ZN(_u0_ch9_am1[19] ) );
INV_X4 _u0_U18621  ( .A(1'b0), .ZN(_u0_ch9_am1[18] ) );
INV_X4 _u0_U18619  ( .A(1'b0), .ZN(_u0_ch9_am1[17] ) );
INV_X4 _u0_U18617  ( .A(1'b0), .ZN(_u0_ch9_am1[16] ) );
INV_X4 _u0_U18615  ( .A(1'b0), .ZN(_u0_ch9_am1[15] ) );
INV_X4 _u0_U18613  ( .A(1'b0), .ZN(_u0_ch9_am1[14] ) );
INV_X4 _u0_U18611  ( .A(1'b0), .ZN(_u0_ch9_am1[13] ) );
INV_X4 _u0_U18609  ( .A(1'b0), .ZN(_u0_ch9_am1[12] ) );
INV_X4 _u0_U18607  ( .A(1'b0), .ZN(_u0_ch9_am1[11] ) );
INV_X4 _u0_U18605  ( .A(1'b0), .ZN(_u0_ch9_am1[10] ) );
INV_X4 _u0_U18603  ( .A(1'b0), .ZN(_u0_ch9_am1[9] ) );
INV_X4 _u0_U18601  ( .A(1'b0), .ZN(_u0_ch9_am1[8] ) );
INV_X4 _u0_U18599  ( .A(1'b0), .ZN(_u0_ch9_am1[7] ) );
INV_X4 _u0_U18597  ( .A(1'b0), .ZN(_u0_ch9_am1[6] ) );
INV_X4 _u0_U18595  ( .A(1'b0), .ZN(_u0_ch9_am1[5] ) );
INV_X4 _u0_U18593  ( .A(1'b0), .ZN(_u0_ch9_am1[4] ) );
INV_X4 _u0_U18591  ( .A(1'b1), .ZN(_u0_ch9_am1[3] ) );
INV_X4 _u0_U18589  ( .A(1'b1), .ZN(_u0_ch9_am1[2] ) );
INV_X4 _u0_U18587  ( .A(1'b1), .ZN(_u0_ch9_am1[1] ) );
INV_X4 _u0_U18585  ( .A(1'b1), .ZN(_u0_ch9_am1[0] ) );
INV_X4 _u0_U18583  ( .A(1'b1), .ZN(_u0_pointer10[31] ) );
INV_X4 _u0_U18581  ( .A(1'b1), .ZN(_u0_pointer10[30] ) );
INV_X4 _u0_U18579  ( .A(1'b1), .ZN(_u0_pointer10[29] ) );
INV_X4 _u0_U18577  ( .A(1'b1), .ZN(_u0_pointer10[28] ) );
INV_X4 _u0_U18575  ( .A(1'b1), .ZN(_u0_pointer10[27] ) );
INV_X4 _u0_U18573  ( .A(1'b1), .ZN(_u0_pointer10[26] ) );
INV_X4 _u0_U18571  ( .A(1'b1), .ZN(_u0_pointer10[25] ) );
INV_X4 _u0_U18569  ( .A(1'b1), .ZN(_u0_pointer10[24] ) );
INV_X4 _u0_U18567  ( .A(1'b1), .ZN(_u0_pointer10[23] ) );
INV_X4 _u0_U18565  ( .A(1'b1), .ZN(_u0_pointer10[22] ) );
INV_X4 _u0_U18563  ( .A(1'b1), .ZN(_u0_pointer10[21] ) );
INV_X4 _u0_U18561  ( .A(1'b1), .ZN(_u0_pointer10[20] ) );
INV_X4 _u0_U18559  ( .A(1'b1), .ZN(_u0_pointer10[19] ) );
INV_X4 _u0_U18557  ( .A(1'b1), .ZN(_u0_pointer10[18] ) );
INV_X4 _u0_U18555  ( .A(1'b1), .ZN(_u0_pointer10[17] ) );
INV_X4 _u0_U18553  ( .A(1'b1), .ZN(_u0_pointer10[16] ) );
INV_X4 _u0_U18551  ( .A(1'b1), .ZN(_u0_pointer10[15] ) );
INV_X4 _u0_U18549  ( .A(1'b1), .ZN(_u0_pointer10[14] ) );
INV_X4 _u0_U18547  ( .A(1'b1), .ZN(_u0_pointer10[13] ) );
INV_X4 _u0_U18545  ( .A(1'b1), .ZN(_u0_pointer10[12] ) );
INV_X4 _u0_U18543  ( .A(1'b1), .ZN(_u0_pointer10[11] ) );
INV_X4 _u0_U18541  ( .A(1'b1), .ZN(_u0_pointer10[10] ) );
INV_X4 _u0_U18539  ( .A(1'b1), .ZN(_u0_pointer10[9] ) );
INV_X4 _u0_U18537  ( .A(1'b1), .ZN(_u0_pointer10[8] ) );
INV_X4 _u0_U18535  ( .A(1'b1), .ZN(_u0_pointer10[7] ) );
INV_X4 _u0_U18533  ( .A(1'b1), .ZN(_u0_pointer10[6] ) );
INV_X4 _u0_U18531  ( .A(1'b1), .ZN(_u0_pointer10[5] ) );
INV_X4 _u0_U18529  ( .A(1'b1), .ZN(_u0_pointer10[4] ) );
INV_X4 _u0_U18527  ( .A(1'b1), .ZN(_u0_pointer10[3] ) );
INV_X4 _u0_U18525  ( .A(1'b1), .ZN(_u0_pointer10[2] ) );
INV_X4 _u0_U18523  ( .A(1'b1), .ZN(_u0_pointer10[1] ) );
INV_X4 _u0_U18521  ( .A(1'b1), .ZN(_u0_pointer10[0] ) );
INV_X4 _u0_U18519  ( .A(1'b1), .ZN(_u0_pointer10_s[31] ) );
INV_X4 _u0_U18517  ( .A(1'b1), .ZN(_u0_pointer10_s[30] ) );
INV_X4 _u0_U18515  ( .A(1'b1), .ZN(_u0_pointer10_s[29] ) );
INV_X4 _u0_U18513  ( .A(1'b1), .ZN(_u0_pointer10_s[28] ) );
INV_X4 _u0_U18511  ( .A(1'b1), .ZN(_u0_pointer10_s[27] ) );
INV_X4 _u0_U18509  ( .A(1'b1), .ZN(_u0_pointer10_s[26] ) );
INV_X4 _u0_U18507  ( .A(1'b1), .ZN(_u0_pointer10_s[25] ) );
INV_X4 _u0_U18505  ( .A(1'b1), .ZN(_u0_pointer10_s[24] ) );
INV_X4 _u0_U18503  ( .A(1'b1), .ZN(_u0_pointer10_s[23] ) );
INV_X4 _u0_U18501  ( .A(1'b1), .ZN(_u0_pointer10_s[22] ) );
INV_X4 _u0_U18499  ( .A(1'b1), .ZN(_u0_pointer10_s[21] ) );
INV_X4 _u0_U18497  ( .A(1'b1), .ZN(_u0_pointer10_s[20] ) );
INV_X4 _u0_U18495  ( .A(1'b1), .ZN(_u0_pointer10_s[19] ) );
INV_X4 _u0_U18493  ( .A(1'b1), .ZN(_u0_pointer10_s[18] ) );
INV_X4 _u0_U18491  ( .A(1'b1), .ZN(_u0_pointer10_s[17] ) );
INV_X4 _u0_U18489  ( .A(1'b1), .ZN(_u0_pointer10_s[16] ) );
INV_X4 _u0_U18487  ( .A(1'b1), .ZN(_u0_pointer10_s[15] ) );
INV_X4 _u0_U18485  ( .A(1'b1), .ZN(_u0_pointer10_s[14] ) );
INV_X4 _u0_U18483  ( .A(1'b1), .ZN(_u0_pointer10_s[13] ) );
INV_X4 _u0_U18481  ( .A(1'b1), .ZN(_u0_pointer10_s[12] ) );
INV_X4 _u0_U18479  ( .A(1'b1), .ZN(_u0_pointer10_s[11] ) );
INV_X4 _u0_U18477  ( .A(1'b1), .ZN(_u0_pointer10_s[10] ) );
INV_X4 _u0_U18475  ( .A(1'b1), .ZN(_u0_pointer10_s[9] ) );
INV_X4 _u0_U18473  ( .A(1'b1), .ZN(_u0_pointer10_s[8] ) );
INV_X4 _u0_U18471  ( .A(1'b1), .ZN(_u0_pointer10_s[7] ) );
INV_X4 _u0_U18469  ( .A(1'b1), .ZN(_u0_pointer10_s[6] ) );
INV_X4 _u0_U18467  ( .A(1'b1), .ZN(_u0_pointer10_s[5] ) );
INV_X4 _u0_U18465  ( .A(1'b1), .ZN(_u0_pointer10_s[4] ) );
INV_X4 _u0_U18463  ( .A(1'b1), .ZN(_u0_pointer10_s[3] ) );
INV_X4 _u0_U18461  ( .A(1'b1), .ZN(_u0_pointer10_s[2] ) );
INV_X4 _u0_U18459  ( .A(1'b1), .ZN(_u0_pointer10_s[1] ) );
INV_X4 _u0_U18457  ( .A(1'b1), .ZN(_u0_pointer10_s[0] ) );
INV_X4 _u0_U18455  ( .A(1'b1), .ZN(_u0_ch10_csr[31] ) );
INV_X4 _u0_U18453  ( .A(1'b1), .ZN(_u0_ch10_csr[30] ) );
INV_X4 _u0_U18451  ( .A(1'b1), .ZN(_u0_ch10_csr[29] ) );
INV_X4 _u0_U18449  ( .A(1'b1), .ZN(_u0_ch10_csr[28] ) );
INV_X4 _u0_U18447  ( .A(1'b1), .ZN(_u0_ch10_csr[27] ) );
INV_X4 _u0_U18445  ( .A(1'b1), .ZN(_u0_ch10_csr[26] ) );
INV_X4 _u0_U18443  ( .A(1'b1), .ZN(_u0_ch10_csr[25] ) );
INV_X4 _u0_U18441  ( .A(1'b1), .ZN(_u0_ch10_csr[24] ) );
INV_X4 _u0_U18439  ( .A(1'b1), .ZN(_u0_ch10_csr[23] ) );
INV_X4 _u0_U18437  ( .A(1'b1), .ZN(_u0_ch10_csr[22] ) );
INV_X4 _u0_U18435  ( .A(1'b1), .ZN(_u0_ch10_csr[21] ) );
INV_X4 _u0_U18433  ( .A(1'b1), .ZN(_u0_ch10_csr[20] ) );
INV_X4 _u0_U18431  ( .A(1'b1), .ZN(_u0_ch10_csr[19] ) );
INV_X4 _u0_U18429  ( .A(1'b1), .ZN(_u0_ch10_csr[18] ) );
INV_X4 _u0_U18427  ( .A(1'b1), .ZN(_u0_ch10_csr[17] ) );
INV_X4 _u0_U18425  ( .A(1'b1), .ZN(_u0_ch10_csr[16] ) );
INV_X4 _u0_U18423  ( .A(1'b1), .ZN(_u0_ch10_csr[15] ) );
INV_X4 _u0_U18421  ( .A(1'b1), .ZN(_u0_ch10_csr[14] ) );
INV_X4 _u0_U18419  ( .A(1'b1), .ZN(_u0_ch10_csr[13] ) );
INV_X4 _u0_U18417  ( .A(1'b1), .ZN(_u0_ch10_csr[12] ) );
INV_X4 _u0_U18415  ( .A(1'b1), .ZN(_u0_ch10_csr[11] ) );
INV_X4 _u0_U18413  ( .A(1'b1), .ZN(_u0_ch10_csr[10] ) );
INV_X4 _u0_U18411  ( .A(1'b1), .ZN(_u0_ch10_csr[9] ) );
INV_X4 _u0_U18409  ( .A(1'b1), .ZN(_u0_ch10_csr[8] ) );
INV_X4 _u0_U18407  ( .A(1'b1), .ZN(_u0_ch10_csr[7] ) );
INV_X4 _u0_U18405  ( .A(1'b1), .ZN(_u0_ch10_csr[6] ) );
INV_X4 _u0_U18403  ( .A(1'b1), .ZN(_u0_ch10_csr[5] ) );
INV_X4 _u0_U18401  ( .A(1'b1), .ZN(_u0_ch10_csr[4] ) );
INV_X4 _u0_U18399  ( .A(1'b1), .ZN(_u0_ch10_csr[3] ) );
INV_X4 _u0_U18397  ( .A(1'b1), .ZN(_u0_ch10_csr[2] ) );
INV_X4 _u0_U18395  ( .A(1'b1), .ZN(_u0_ch10_csr[1] ) );
INV_X4 _u0_U18393  ( .A(1'b1), .ZN(_u0_ch10_csr[0] ) );
INV_X4 _u0_U18391  ( .A(1'b1), .ZN(_u0_ch10_txsz[31] ) );
INV_X4 _u0_U18389  ( .A(1'b1), .ZN(_u0_ch10_txsz[30] ) );
INV_X4 _u0_U18387  ( .A(1'b1), .ZN(_u0_ch10_txsz[29] ) );
INV_X4 _u0_U18385  ( .A(1'b1), .ZN(_u0_ch10_txsz[28] ) );
INV_X4 _u0_U18383  ( .A(1'b1), .ZN(_u0_ch10_txsz[27] ) );
INV_X4 _u0_U18381  ( .A(1'b1), .ZN(_u0_ch10_txsz[26] ) );
INV_X4 _u0_U18379  ( .A(1'b1), .ZN(_u0_ch10_txsz[25] ) );
INV_X4 _u0_U18377  ( .A(1'b1), .ZN(_u0_ch10_txsz[24] ) );
INV_X4 _u0_U18375  ( .A(1'b1), .ZN(_u0_ch10_txsz[23] ) );
INV_X4 _u0_U18373  ( .A(1'b1), .ZN(_u0_ch10_txsz[22] ) );
INV_X4 _u0_U18371  ( .A(1'b1), .ZN(_u0_ch10_txsz[21] ) );
INV_X4 _u0_U18369  ( .A(1'b1), .ZN(_u0_ch10_txsz[20] ) );
INV_X4 _u0_U18367  ( .A(1'b1), .ZN(_u0_ch10_txsz[19] ) );
INV_X4 _u0_U18365  ( .A(1'b1), .ZN(_u0_ch10_txsz[18] ) );
INV_X4 _u0_U18363  ( .A(1'b1), .ZN(_u0_ch10_txsz[17] ) );
INV_X4 _u0_U18361  ( .A(1'b1), .ZN(_u0_ch10_txsz[16] ) );
INV_X4 _u0_U18359  ( .A(1'b1), .ZN(_u0_ch10_txsz[15] ) );
INV_X4 _u0_U18357  ( .A(1'b1), .ZN(_u0_ch10_txsz[14] ) );
INV_X4 _u0_U18355  ( .A(1'b1), .ZN(_u0_ch10_txsz[13] ) );
INV_X4 _u0_U18353  ( .A(1'b1), .ZN(_u0_ch10_txsz[12] ) );
INV_X4 _u0_U18351  ( .A(1'b1), .ZN(_u0_ch10_txsz[11] ) );
INV_X4 _u0_U18349  ( .A(1'b1), .ZN(_u0_ch10_txsz[10] ) );
INV_X4 _u0_U18347  ( .A(1'b1), .ZN(_u0_ch10_txsz[9] ) );
INV_X4 _u0_U18345  ( .A(1'b1), .ZN(_u0_ch10_txsz[8] ) );
INV_X4 _u0_U18343  ( .A(1'b1), .ZN(_u0_ch10_txsz[7] ) );
INV_X4 _u0_U18341  ( .A(1'b1), .ZN(_u0_ch10_txsz[6] ) );
INV_X4 _u0_U18339  ( .A(1'b1), .ZN(_u0_ch10_txsz[5] ) );
INV_X4 _u0_U18337  ( .A(1'b1), .ZN(_u0_ch10_txsz[4] ) );
INV_X4 _u0_U18335  ( .A(1'b1), .ZN(_u0_ch10_txsz[3] ) );
INV_X4 _u0_U18333  ( .A(1'b1), .ZN(_u0_ch10_txsz[2] ) );
INV_X4 _u0_U18331  ( .A(1'b1), .ZN(_u0_ch10_txsz[1] ) );
INV_X4 _u0_U18329  ( .A(1'b1), .ZN(_u0_ch10_txsz[0] ) );
INV_X4 _u0_U18327  ( .A(1'b1), .ZN(_u0_ch10_adr0[31] ) );
INV_X4 _u0_U18325  ( .A(1'b1), .ZN(_u0_ch10_adr0[30] ) );
INV_X4 _u0_U18323  ( .A(1'b1), .ZN(_u0_ch10_adr0[29] ) );
INV_X4 _u0_U18321  ( .A(1'b1), .ZN(_u0_ch10_adr0[28] ) );
INV_X4 _u0_U18319  ( .A(1'b1), .ZN(_u0_ch10_adr0[27] ) );
INV_X4 _u0_U18317  ( .A(1'b1), .ZN(_u0_ch10_adr0[26] ) );
INV_X4 _u0_U18315  ( .A(1'b1), .ZN(_u0_ch10_adr0[25] ) );
INV_X4 _u0_U18313  ( .A(1'b1), .ZN(_u0_ch10_adr0[24] ) );
INV_X4 _u0_U18311  ( .A(1'b1), .ZN(_u0_ch10_adr0[23] ) );
INV_X4 _u0_U18309  ( .A(1'b1), .ZN(_u0_ch10_adr0[22] ) );
INV_X4 _u0_U18307  ( .A(1'b1), .ZN(_u0_ch10_adr0[21] ) );
INV_X4 _u0_U18305  ( .A(1'b1), .ZN(_u0_ch10_adr0[20] ) );
INV_X4 _u0_U18303  ( .A(1'b1), .ZN(_u0_ch10_adr0[19] ) );
INV_X4 _u0_U18301  ( .A(1'b1), .ZN(_u0_ch10_adr0[18] ) );
INV_X4 _u0_U18299  ( .A(1'b1), .ZN(_u0_ch10_adr0[17] ) );
INV_X4 _u0_U18297  ( .A(1'b1), .ZN(_u0_ch10_adr0[16] ) );
INV_X4 _u0_U18295  ( .A(1'b1), .ZN(_u0_ch10_adr0[15] ) );
INV_X4 _u0_U18293  ( .A(1'b1), .ZN(_u0_ch10_adr0[14] ) );
INV_X4 _u0_U18291  ( .A(1'b1), .ZN(_u0_ch10_adr0[13] ) );
INV_X4 _u0_U18289  ( .A(1'b1), .ZN(_u0_ch10_adr0[12] ) );
INV_X4 _u0_U18287  ( .A(1'b1), .ZN(_u0_ch10_adr0[11] ) );
INV_X4 _u0_U18285  ( .A(1'b1), .ZN(_u0_ch10_adr0[10] ) );
INV_X4 _u0_U18283  ( .A(1'b1), .ZN(_u0_ch10_adr0[9] ) );
INV_X4 _u0_U18281  ( .A(1'b1), .ZN(_u0_ch10_adr0[8] ) );
INV_X4 _u0_U18279  ( .A(1'b1), .ZN(_u0_ch10_adr0[7] ) );
INV_X4 _u0_U18277  ( .A(1'b1), .ZN(_u0_ch10_adr0[6] ) );
INV_X4 _u0_U18275  ( .A(1'b1), .ZN(_u0_ch10_adr0[5] ) );
INV_X4 _u0_U18273  ( .A(1'b1), .ZN(_u0_ch10_adr0[4] ) );
INV_X4 _u0_U18271  ( .A(1'b1), .ZN(_u0_ch10_adr0[3] ) );
INV_X4 _u0_U18269  ( .A(1'b1), .ZN(_u0_ch10_adr0[2] ) );
INV_X4 _u0_U18267  ( .A(1'b1), .ZN(_u0_ch10_adr0[1] ) );
INV_X4 _u0_U18265  ( .A(1'b1), .ZN(_u0_ch10_adr0[0] ) );
INV_X4 _u0_U18263  ( .A(1'b1), .ZN(_u0_ch10_adr1[31] ) );
INV_X4 _u0_U18261  ( .A(1'b1), .ZN(_u0_ch10_adr1[30] ) );
INV_X4 _u0_U18259  ( .A(1'b1), .ZN(_u0_ch10_adr1[29] ) );
INV_X4 _u0_U18257  ( .A(1'b1), .ZN(_u0_ch10_adr1[28] ) );
INV_X4 _u0_U18255  ( .A(1'b1), .ZN(_u0_ch10_adr1[27] ) );
INV_X4 _u0_U18253  ( .A(1'b1), .ZN(_u0_ch10_adr1[26] ) );
INV_X4 _u0_U18251  ( .A(1'b1), .ZN(_u0_ch10_adr1[25] ) );
INV_X4 _u0_U18249  ( .A(1'b1), .ZN(_u0_ch10_adr1[24] ) );
INV_X4 _u0_U18247  ( .A(1'b1), .ZN(_u0_ch10_adr1[23] ) );
INV_X4 _u0_U18245  ( .A(1'b1), .ZN(_u0_ch10_adr1[22] ) );
INV_X4 _u0_U18243  ( .A(1'b1), .ZN(_u0_ch10_adr1[21] ) );
INV_X4 _u0_U18241  ( .A(1'b1), .ZN(_u0_ch10_adr1[20] ) );
INV_X4 _u0_U18239  ( .A(1'b1), .ZN(_u0_ch10_adr1[19] ) );
INV_X4 _u0_U18237  ( .A(1'b1), .ZN(_u0_ch10_adr1[18] ) );
INV_X4 _u0_U18235  ( .A(1'b1), .ZN(_u0_ch10_adr1[17] ) );
INV_X4 _u0_U18233  ( .A(1'b1), .ZN(_u0_ch10_adr1[16] ) );
INV_X4 _u0_U18231  ( .A(1'b1), .ZN(_u0_ch10_adr1[15] ) );
INV_X4 _u0_U18229  ( .A(1'b1), .ZN(_u0_ch10_adr1[14] ) );
INV_X4 _u0_U18227  ( .A(1'b1), .ZN(_u0_ch10_adr1[13] ) );
INV_X4 _u0_U18225  ( .A(1'b1), .ZN(_u0_ch10_adr1[12] ) );
INV_X4 _u0_U18223  ( .A(1'b1), .ZN(_u0_ch10_adr1[11] ) );
INV_X4 _u0_U18221  ( .A(1'b1), .ZN(_u0_ch10_adr1[10] ) );
INV_X4 _u0_U18219  ( .A(1'b1), .ZN(_u0_ch10_adr1[9] ) );
INV_X4 _u0_U18217  ( .A(1'b1), .ZN(_u0_ch10_adr1[8] ) );
INV_X4 _u0_U18215  ( .A(1'b1), .ZN(_u0_ch10_adr1[7] ) );
INV_X4 _u0_U18213  ( .A(1'b1), .ZN(_u0_ch10_adr1[6] ) );
INV_X4 _u0_U18211  ( .A(1'b1), .ZN(_u0_ch10_adr1[5] ) );
INV_X4 _u0_U18209  ( .A(1'b1), .ZN(_u0_ch10_adr1[4] ) );
INV_X4 _u0_U18207  ( .A(1'b1), .ZN(_u0_ch10_adr1[3] ) );
INV_X4 _u0_U18205  ( .A(1'b1), .ZN(_u0_ch10_adr1[2] ) );
INV_X4 _u0_U18203  ( .A(1'b1), .ZN(_u0_ch10_adr1[1] ) );
INV_X4 _u0_U18201  ( .A(1'b1), .ZN(_u0_ch10_adr1[0] ) );
INV_X4 _u0_U18199  ( .A(1'b0), .ZN(_u0_ch10_am0[31] ) );
INV_X4 _u0_U18197  ( .A(1'b0), .ZN(_u0_ch10_am0[30] ) );
INV_X4 _u0_U18195  ( .A(1'b0), .ZN(_u0_ch10_am0[29] ) );
INV_X4 _u0_U18193  ( .A(1'b0), .ZN(_u0_ch10_am0[28] ) );
INV_X4 _u0_U18191  ( .A(1'b0), .ZN(_u0_ch10_am0[27] ) );
INV_X4 _u0_U18189  ( .A(1'b0), .ZN(_u0_ch10_am0[26] ) );
INV_X4 _u0_U18187  ( .A(1'b0), .ZN(_u0_ch10_am0[25] ) );
INV_X4 _u0_U18185  ( .A(1'b0), .ZN(_u0_ch10_am0[24] ) );
INV_X4 _u0_U18183  ( .A(1'b0), .ZN(_u0_ch10_am0[23] ) );
INV_X4 _u0_U18181  ( .A(1'b0), .ZN(_u0_ch10_am0[22] ) );
INV_X4 _u0_U18179  ( .A(1'b0), .ZN(_u0_ch10_am0[21] ) );
INV_X4 _u0_U18177  ( .A(1'b0), .ZN(_u0_ch10_am0[20] ) );
INV_X4 _u0_U18175  ( .A(1'b0), .ZN(_u0_ch10_am0[19] ) );
INV_X4 _u0_U18173  ( .A(1'b0), .ZN(_u0_ch10_am0[18] ) );
INV_X4 _u0_U18171  ( .A(1'b0), .ZN(_u0_ch10_am0[17] ) );
INV_X4 _u0_U18169  ( .A(1'b0), .ZN(_u0_ch10_am0[16] ) );
INV_X4 _u0_U18167  ( .A(1'b0), .ZN(_u0_ch10_am0[15] ) );
INV_X4 _u0_U18165  ( .A(1'b0), .ZN(_u0_ch10_am0[14] ) );
INV_X4 _u0_U18163  ( .A(1'b0), .ZN(_u0_ch10_am0[13] ) );
INV_X4 _u0_U18161  ( .A(1'b0), .ZN(_u0_ch10_am0[12] ) );
INV_X4 _u0_U18159  ( .A(1'b0), .ZN(_u0_ch10_am0[11] ) );
INV_X4 _u0_U18157  ( .A(1'b0), .ZN(_u0_ch10_am0[10] ) );
INV_X4 _u0_U18155  ( .A(1'b0), .ZN(_u0_ch10_am0[9] ) );
INV_X4 _u0_U18153  ( .A(1'b0), .ZN(_u0_ch10_am0[8] ) );
INV_X4 _u0_U18151  ( .A(1'b0), .ZN(_u0_ch10_am0[7] ) );
INV_X4 _u0_U18149  ( .A(1'b0), .ZN(_u0_ch10_am0[6] ) );
INV_X4 _u0_U18147  ( .A(1'b0), .ZN(_u0_ch10_am0[5] ) );
INV_X4 _u0_U18145  ( .A(1'b0), .ZN(_u0_ch10_am0[4] ) );
INV_X4 _u0_U18143  ( .A(1'b1), .ZN(_u0_ch10_am0[3] ) );
INV_X4 _u0_U18141  ( .A(1'b1), .ZN(_u0_ch10_am0[2] ) );
INV_X4 _u0_U18139  ( .A(1'b1), .ZN(_u0_ch10_am0[1] ) );
INV_X4 _u0_U18137  ( .A(1'b1), .ZN(_u0_ch10_am0[0] ) );
INV_X4 _u0_U18135  ( .A(1'b0), .ZN(_u0_ch10_am1[31] ) );
INV_X4 _u0_U18133  ( .A(1'b0), .ZN(_u0_ch10_am1[30] ) );
INV_X4 _u0_U18131  ( .A(1'b0), .ZN(_u0_ch10_am1[29] ) );
INV_X4 _u0_U18129  ( .A(1'b0), .ZN(_u0_ch10_am1[28] ) );
INV_X4 _u0_U18127  ( .A(1'b0), .ZN(_u0_ch10_am1[27] ) );
INV_X4 _u0_U18125  ( .A(1'b0), .ZN(_u0_ch10_am1[26] ) );
INV_X4 _u0_U18123  ( .A(1'b0), .ZN(_u0_ch10_am1[25] ) );
INV_X4 _u0_U18121  ( .A(1'b0), .ZN(_u0_ch10_am1[24] ) );
INV_X4 _u0_U18119  ( .A(1'b0), .ZN(_u0_ch10_am1[23] ) );
INV_X4 _u0_U18117  ( .A(1'b0), .ZN(_u0_ch10_am1[22] ) );
INV_X4 _u0_U18115  ( .A(1'b0), .ZN(_u0_ch10_am1[21] ) );
INV_X4 _u0_U18113  ( .A(1'b0), .ZN(_u0_ch10_am1[20] ) );
INV_X4 _u0_U18111  ( .A(1'b0), .ZN(_u0_ch10_am1[19] ) );
INV_X4 _u0_U18109  ( .A(1'b0), .ZN(_u0_ch10_am1[18] ) );
INV_X4 _u0_U18107  ( .A(1'b0), .ZN(_u0_ch10_am1[17] ) );
INV_X4 _u0_U18105  ( .A(1'b0), .ZN(_u0_ch10_am1[16] ) );
INV_X4 _u0_U18103  ( .A(1'b0), .ZN(_u0_ch10_am1[15] ) );
INV_X4 _u0_U18101  ( .A(1'b0), .ZN(_u0_ch10_am1[14] ) );
INV_X4 _u0_U18099  ( .A(1'b0), .ZN(_u0_ch10_am1[13] ) );
INV_X4 _u0_U18097  ( .A(1'b0), .ZN(_u0_ch10_am1[12] ) );
INV_X4 _u0_U18095  ( .A(1'b0), .ZN(_u0_ch10_am1[11] ) );
INV_X4 _u0_U18093  ( .A(1'b0), .ZN(_u0_ch10_am1[10] ) );
INV_X4 _u0_U18091  ( .A(1'b0), .ZN(_u0_ch10_am1[9] ) );
INV_X4 _u0_U18089  ( .A(1'b0), .ZN(_u0_ch10_am1[8] ) );
INV_X4 _u0_U18087  ( .A(1'b0), .ZN(_u0_ch10_am1[7] ) );
INV_X4 _u0_U18085  ( .A(1'b0), .ZN(_u0_ch10_am1[6] ) );
INV_X4 _u0_U18083  ( .A(1'b0), .ZN(_u0_ch10_am1[5] ) );
INV_X4 _u0_U18081  ( .A(1'b0), .ZN(_u0_ch10_am1[4] ) );
INV_X4 _u0_U18079  ( .A(1'b1), .ZN(_u0_ch10_am1[3] ) );
INV_X4 _u0_U18077  ( .A(1'b1), .ZN(_u0_ch10_am1[2] ) );
INV_X4 _u0_U18075  ( .A(1'b1), .ZN(_u0_ch10_am1[1] ) );
INV_X4 _u0_U18073  ( .A(1'b1), .ZN(_u0_ch10_am1[0] ) );
INV_X4 _u0_U18071  ( .A(1'b1), .ZN(_u0_pointer11[31] ) );
INV_X4 _u0_U18069  ( .A(1'b1), .ZN(_u0_pointer11[30] ) );
INV_X4 _u0_U18067  ( .A(1'b1), .ZN(_u0_pointer11[29] ) );
INV_X4 _u0_U18065  ( .A(1'b1), .ZN(_u0_pointer11[28] ) );
INV_X4 _u0_U18063  ( .A(1'b1), .ZN(_u0_pointer11[27] ) );
INV_X4 _u0_U18061  ( .A(1'b1), .ZN(_u0_pointer11[26] ) );
INV_X4 _u0_U18059  ( .A(1'b1), .ZN(_u0_pointer11[25] ) );
INV_X4 _u0_U18057  ( .A(1'b1), .ZN(_u0_pointer11[24] ) );
INV_X4 _u0_U18055  ( .A(1'b1), .ZN(_u0_pointer11[23] ) );
INV_X4 _u0_U18053  ( .A(1'b1), .ZN(_u0_pointer11[22] ) );
INV_X4 _u0_U18051  ( .A(1'b1), .ZN(_u0_pointer11[21] ) );
INV_X4 _u0_U18049  ( .A(1'b1), .ZN(_u0_pointer11[20] ) );
INV_X4 _u0_U18047  ( .A(1'b1), .ZN(_u0_pointer11[19] ) );
INV_X4 _u0_U18045  ( .A(1'b1), .ZN(_u0_pointer11[18] ) );
INV_X4 _u0_U18043  ( .A(1'b1), .ZN(_u0_pointer11[17] ) );
INV_X4 _u0_U18041  ( .A(1'b1), .ZN(_u0_pointer11[16] ) );
INV_X4 _u0_U18039  ( .A(1'b1), .ZN(_u0_pointer11[15] ) );
INV_X4 _u0_U18037  ( .A(1'b1), .ZN(_u0_pointer11[14] ) );
INV_X4 _u0_U18035  ( .A(1'b1), .ZN(_u0_pointer11[13] ) );
INV_X4 _u0_U18033  ( .A(1'b1), .ZN(_u0_pointer11[12] ) );
INV_X4 _u0_U18031  ( .A(1'b1), .ZN(_u0_pointer11[11] ) );
INV_X4 _u0_U18029  ( .A(1'b1), .ZN(_u0_pointer11[10] ) );
INV_X4 _u0_U18027  ( .A(1'b1), .ZN(_u0_pointer11[9] ) );
INV_X4 _u0_U18025  ( .A(1'b1), .ZN(_u0_pointer11[8] ) );
INV_X4 _u0_U18023  ( .A(1'b1), .ZN(_u0_pointer11[7] ) );
INV_X4 _u0_U18021  ( .A(1'b1), .ZN(_u0_pointer11[6] ) );
INV_X4 _u0_U18019  ( .A(1'b1), .ZN(_u0_pointer11[5] ) );
INV_X4 _u0_U18017  ( .A(1'b1), .ZN(_u0_pointer11[4] ) );
INV_X4 _u0_U18015  ( .A(1'b1), .ZN(_u0_pointer11[3] ) );
INV_X4 _u0_U18013  ( .A(1'b1), .ZN(_u0_pointer11[2] ) );
INV_X4 _u0_U18011  ( .A(1'b1), .ZN(_u0_pointer11[1] ) );
INV_X4 _u0_U18009  ( .A(1'b1), .ZN(_u0_pointer11[0] ) );
INV_X4 _u0_U18007  ( .A(1'b1), .ZN(_u0_pointer11_s[31] ) );
INV_X4 _u0_U18005  ( .A(1'b1), .ZN(_u0_pointer11_s[30] ) );
INV_X4 _u0_U18003  ( .A(1'b1), .ZN(_u0_pointer11_s[29] ) );
INV_X4 _u0_U18001  ( .A(1'b1), .ZN(_u0_pointer11_s[28] ) );
INV_X4 _u0_U17999  ( .A(1'b1), .ZN(_u0_pointer11_s[27] ) );
INV_X4 _u0_U17997  ( .A(1'b1), .ZN(_u0_pointer11_s[26] ) );
INV_X4 _u0_U17995  ( .A(1'b1), .ZN(_u0_pointer11_s[25] ) );
INV_X4 _u0_U17993  ( .A(1'b1), .ZN(_u0_pointer11_s[24] ) );
INV_X4 _u0_U17991  ( .A(1'b1), .ZN(_u0_pointer11_s[23] ) );
INV_X4 _u0_U17989  ( .A(1'b1), .ZN(_u0_pointer11_s[22] ) );
INV_X4 _u0_U17987  ( .A(1'b1), .ZN(_u0_pointer11_s[21] ) );
INV_X4 _u0_U17985  ( .A(1'b1), .ZN(_u0_pointer11_s[20] ) );
INV_X4 _u0_U17983  ( .A(1'b1), .ZN(_u0_pointer11_s[19] ) );
INV_X4 _u0_U17981  ( .A(1'b1), .ZN(_u0_pointer11_s[18] ) );
INV_X4 _u0_U17979  ( .A(1'b1), .ZN(_u0_pointer11_s[17] ) );
INV_X4 _u0_U17977  ( .A(1'b1), .ZN(_u0_pointer11_s[16] ) );
INV_X4 _u0_U17975  ( .A(1'b1), .ZN(_u0_pointer11_s[15] ) );
INV_X4 _u0_U17973  ( .A(1'b1), .ZN(_u0_pointer11_s[14] ) );
INV_X4 _u0_U17971  ( .A(1'b1), .ZN(_u0_pointer11_s[13] ) );
INV_X4 _u0_U17969  ( .A(1'b1), .ZN(_u0_pointer11_s[12] ) );
INV_X4 _u0_U17967  ( .A(1'b1), .ZN(_u0_pointer11_s[11] ) );
INV_X4 _u0_U17965  ( .A(1'b1), .ZN(_u0_pointer11_s[10] ) );
INV_X4 _u0_U17963  ( .A(1'b1), .ZN(_u0_pointer11_s[9] ) );
INV_X4 _u0_U17961  ( .A(1'b1), .ZN(_u0_pointer11_s[8] ) );
INV_X4 _u0_U17959  ( .A(1'b1), .ZN(_u0_pointer11_s[7] ) );
INV_X4 _u0_U17957  ( .A(1'b1), .ZN(_u0_pointer11_s[6] ) );
INV_X4 _u0_U17955  ( .A(1'b1), .ZN(_u0_pointer11_s[5] ) );
INV_X4 _u0_U17953  ( .A(1'b1), .ZN(_u0_pointer11_s[4] ) );
INV_X4 _u0_U17951  ( .A(1'b1), .ZN(_u0_pointer11_s[3] ) );
INV_X4 _u0_U17949  ( .A(1'b1), .ZN(_u0_pointer11_s[2] ) );
INV_X4 _u0_U17947  ( .A(1'b1), .ZN(_u0_pointer11_s[1] ) );
INV_X4 _u0_U17945  ( .A(1'b1), .ZN(_u0_pointer11_s[0] ) );
INV_X4 _u0_U17943  ( .A(1'b1), .ZN(_u0_ch11_csr[31] ) );
INV_X4 _u0_U17941  ( .A(1'b1), .ZN(_u0_ch11_csr[30] ) );
INV_X4 _u0_U17939  ( .A(1'b1), .ZN(_u0_ch11_csr[29] ) );
INV_X4 _u0_U17937  ( .A(1'b1), .ZN(_u0_ch11_csr[28] ) );
INV_X4 _u0_U17935  ( .A(1'b1), .ZN(_u0_ch11_csr[27] ) );
INV_X4 _u0_U17933  ( .A(1'b1), .ZN(_u0_ch11_csr[26] ) );
INV_X4 _u0_U17931  ( .A(1'b1), .ZN(_u0_ch11_csr[25] ) );
INV_X4 _u0_U17929  ( .A(1'b1), .ZN(_u0_ch11_csr[24] ) );
INV_X4 _u0_U17927  ( .A(1'b1), .ZN(_u0_ch11_csr[23] ) );
INV_X4 _u0_U17925  ( .A(1'b1), .ZN(_u0_ch11_csr[22] ) );
INV_X4 _u0_U17923  ( .A(1'b1), .ZN(_u0_ch11_csr[21] ) );
INV_X4 _u0_U17921  ( .A(1'b1), .ZN(_u0_ch11_csr[20] ) );
INV_X4 _u0_U17919  ( .A(1'b1), .ZN(_u0_ch11_csr[19] ) );
INV_X4 _u0_U17917  ( .A(1'b1), .ZN(_u0_ch11_csr[18] ) );
INV_X4 _u0_U17915  ( .A(1'b1), .ZN(_u0_ch11_csr[17] ) );
INV_X4 _u0_U17913  ( .A(1'b1), .ZN(_u0_ch11_csr[16] ) );
INV_X4 _u0_U17911  ( .A(1'b1), .ZN(_u0_ch11_csr[15] ) );
INV_X4 _u0_U17909  ( .A(1'b1), .ZN(_u0_ch11_csr[14] ) );
INV_X4 _u0_U17907  ( .A(1'b1), .ZN(_u0_ch11_csr[13] ) );
INV_X4 _u0_U17905  ( .A(1'b1), .ZN(_u0_ch11_csr[12] ) );
INV_X4 _u0_U17903  ( .A(1'b1), .ZN(_u0_ch11_csr[11] ) );
INV_X4 _u0_U17901  ( .A(1'b1), .ZN(_u0_ch11_csr[10] ) );
INV_X4 _u0_U17899  ( .A(1'b1), .ZN(_u0_ch11_csr[9] ) );
INV_X4 _u0_U17897  ( .A(1'b1), .ZN(_u0_ch11_csr[8] ) );
INV_X4 _u0_U17895  ( .A(1'b1), .ZN(_u0_ch11_csr[7] ) );
INV_X4 _u0_U17893  ( .A(1'b1), .ZN(_u0_ch11_csr[6] ) );
INV_X4 _u0_U17891  ( .A(1'b1), .ZN(_u0_ch11_csr[5] ) );
INV_X4 _u0_U17889  ( .A(1'b1), .ZN(_u0_ch11_csr[4] ) );
INV_X4 _u0_U17887  ( .A(1'b1), .ZN(_u0_ch11_csr[3] ) );
INV_X4 _u0_U17885  ( .A(1'b1), .ZN(_u0_ch11_csr[2] ) );
INV_X4 _u0_U17883  ( .A(1'b1), .ZN(_u0_ch11_csr[1] ) );
INV_X4 _u0_U17881  ( .A(1'b1), .ZN(_u0_ch11_csr[0] ) );
INV_X4 _u0_U17879  ( .A(1'b1), .ZN(_u0_ch11_txsz[31] ) );
INV_X4 _u0_U17877  ( .A(1'b1), .ZN(_u0_ch11_txsz[30] ) );
INV_X4 _u0_U17875  ( .A(1'b1), .ZN(_u0_ch11_txsz[29] ) );
INV_X4 _u0_U17873  ( .A(1'b1), .ZN(_u0_ch11_txsz[28] ) );
INV_X4 _u0_U17871  ( .A(1'b1), .ZN(_u0_ch11_txsz[27] ) );
INV_X4 _u0_U17869  ( .A(1'b1), .ZN(_u0_ch11_txsz[26] ) );
INV_X4 _u0_U17867  ( .A(1'b1), .ZN(_u0_ch11_txsz[25] ) );
INV_X4 _u0_U17865  ( .A(1'b1), .ZN(_u0_ch11_txsz[24] ) );
INV_X4 _u0_U17863  ( .A(1'b1), .ZN(_u0_ch11_txsz[23] ) );
INV_X4 _u0_U17861  ( .A(1'b1), .ZN(_u0_ch11_txsz[22] ) );
INV_X4 _u0_U17859  ( .A(1'b1), .ZN(_u0_ch11_txsz[21] ) );
INV_X4 _u0_U17857  ( .A(1'b1), .ZN(_u0_ch11_txsz[20] ) );
INV_X4 _u0_U17855  ( .A(1'b1), .ZN(_u0_ch11_txsz[19] ) );
INV_X4 _u0_U17853  ( .A(1'b1), .ZN(_u0_ch11_txsz[18] ) );
INV_X4 _u0_U17851  ( .A(1'b1), .ZN(_u0_ch11_txsz[17] ) );
INV_X4 _u0_U17849  ( .A(1'b1), .ZN(_u0_ch11_txsz[16] ) );
INV_X4 _u0_U17847  ( .A(1'b1), .ZN(_u0_ch11_txsz[15] ) );
INV_X4 _u0_U17845  ( .A(1'b1), .ZN(_u0_ch11_txsz[14] ) );
INV_X4 _u0_U17843  ( .A(1'b1), .ZN(_u0_ch11_txsz[13] ) );
INV_X4 _u0_U17841  ( .A(1'b1), .ZN(_u0_ch11_txsz[12] ) );
INV_X4 _u0_U17839  ( .A(1'b1), .ZN(_u0_ch11_txsz[11] ) );
INV_X4 _u0_U17837  ( .A(1'b1), .ZN(_u0_ch11_txsz[10] ) );
INV_X4 _u0_U17835  ( .A(1'b1), .ZN(_u0_ch11_txsz[9] ) );
INV_X4 _u0_U17833  ( .A(1'b1), .ZN(_u0_ch11_txsz[8] ) );
INV_X4 _u0_U17831  ( .A(1'b1), .ZN(_u0_ch11_txsz[7] ) );
INV_X4 _u0_U17829  ( .A(1'b1), .ZN(_u0_ch11_txsz[6] ) );
INV_X4 _u0_U17827  ( .A(1'b1), .ZN(_u0_ch11_txsz[5] ) );
INV_X4 _u0_U17825  ( .A(1'b1), .ZN(_u0_ch11_txsz[4] ) );
INV_X4 _u0_U17823  ( .A(1'b1), .ZN(_u0_ch11_txsz[3] ) );
INV_X4 _u0_U17821  ( .A(1'b1), .ZN(_u0_ch11_txsz[2] ) );
INV_X4 _u0_U17819  ( .A(1'b1), .ZN(_u0_ch11_txsz[1] ) );
INV_X4 _u0_U17817  ( .A(1'b1), .ZN(_u0_ch11_txsz[0] ) );
INV_X4 _u0_U17815  ( .A(1'b1), .ZN(_u0_ch11_adr0[31] ) );
INV_X4 _u0_U17813  ( .A(1'b1), .ZN(_u0_ch11_adr0[30] ) );
INV_X4 _u0_U17811  ( .A(1'b1), .ZN(_u0_ch11_adr0[29] ) );
INV_X4 _u0_U17809  ( .A(1'b1), .ZN(_u0_ch11_adr0[28] ) );
INV_X4 _u0_U17807  ( .A(1'b1), .ZN(_u0_ch11_adr0[27] ) );
INV_X4 _u0_U17805  ( .A(1'b1), .ZN(_u0_ch11_adr0[26] ) );
INV_X4 _u0_U17803  ( .A(1'b1), .ZN(_u0_ch11_adr0[25] ) );
INV_X4 _u0_U17801  ( .A(1'b1), .ZN(_u0_ch11_adr0[24] ) );
INV_X4 _u0_U17799  ( .A(1'b1), .ZN(_u0_ch11_adr0[23] ) );
INV_X4 _u0_U17797  ( .A(1'b1), .ZN(_u0_ch11_adr0[22] ) );
INV_X4 _u0_U17795  ( .A(1'b1), .ZN(_u0_ch11_adr0[21] ) );
INV_X4 _u0_U17793  ( .A(1'b1), .ZN(_u0_ch11_adr0[20] ) );
INV_X4 _u0_U17791  ( .A(1'b1), .ZN(_u0_ch11_adr0[19] ) );
INV_X4 _u0_U17789  ( .A(1'b1), .ZN(_u0_ch11_adr0[18] ) );
INV_X4 _u0_U17787  ( .A(1'b1), .ZN(_u0_ch11_adr0[17] ) );
INV_X4 _u0_U17785  ( .A(1'b1), .ZN(_u0_ch11_adr0[16] ) );
INV_X4 _u0_U17783  ( .A(1'b1), .ZN(_u0_ch11_adr0[15] ) );
INV_X4 _u0_U17781  ( .A(1'b1), .ZN(_u0_ch11_adr0[14] ) );
INV_X4 _u0_U17779  ( .A(1'b1), .ZN(_u0_ch11_adr0[13] ) );
INV_X4 _u0_U17777  ( .A(1'b1), .ZN(_u0_ch11_adr0[12] ) );
INV_X4 _u0_U17775  ( .A(1'b1), .ZN(_u0_ch11_adr0[11] ) );
INV_X4 _u0_U17773  ( .A(1'b1), .ZN(_u0_ch11_adr0[10] ) );
INV_X4 _u0_U17771  ( .A(1'b1), .ZN(_u0_ch11_adr0[9] ) );
INV_X4 _u0_U17769  ( .A(1'b1), .ZN(_u0_ch11_adr0[8] ) );
INV_X4 _u0_U17767  ( .A(1'b1), .ZN(_u0_ch11_adr0[7] ) );
INV_X4 _u0_U17765  ( .A(1'b1), .ZN(_u0_ch11_adr0[6] ) );
INV_X4 _u0_U17763  ( .A(1'b1), .ZN(_u0_ch11_adr0[5] ) );
INV_X4 _u0_U17761  ( .A(1'b1), .ZN(_u0_ch11_adr0[4] ) );
INV_X4 _u0_U17759  ( .A(1'b1), .ZN(_u0_ch11_adr0[3] ) );
INV_X4 _u0_U17757  ( .A(1'b1), .ZN(_u0_ch11_adr0[2] ) );
INV_X4 _u0_U17755  ( .A(1'b1), .ZN(_u0_ch11_adr0[1] ) );
INV_X4 _u0_U17753  ( .A(1'b1), .ZN(_u0_ch11_adr0[0] ) );
INV_X4 _u0_U17751  ( .A(1'b1), .ZN(_u0_ch11_adr1[31] ) );
INV_X4 _u0_U17749  ( .A(1'b1), .ZN(_u0_ch11_adr1[30] ) );
INV_X4 _u0_U17747  ( .A(1'b1), .ZN(_u0_ch11_adr1[29] ) );
INV_X4 _u0_U17745  ( .A(1'b1), .ZN(_u0_ch11_adr1[28] ) );
INV_X4 _u0_U17743  ( .A(1'b1), .ZN(_u0_ch11_adr1[27] ) );
INV_X4 _u0_U17741  ( .A(1'b1), .ZN(_u0_ch11_adr1[26] ) );
INV_X4 _u0_U17739  ( .A(1'b1), .ZN(_u0_ch11_adr1[25] ) );
INV_X4 _u0_U17737  ( .A(1'b1), .ZN(_u0_ch11_adr1[24] ) );
INV_X4 _u0_U17735  ( .A(1'b1), .ZN(_u0_ch11_adr1[23] ) );
INV_X4 _u0_U17733  ( .A(1'b1), .ZN(_u0_ch11_adr1[22] ) );
INV_X4 _u0_U17731  ( .A(1'b1), .ZN(_u0_ch11_adr1[21] ) );
INV_X4 _u0_U17729  ( .A(1'b1), .ZN(_u0_ch11_adr1[20] ) );
INV_X4 _u0_U17727  ( .A(1'b1), .ZN(_u0_ch11_adr1[19] ) );
INV_X4 _u0_U17725  ( .A(1'b1), .ZN(_u0_ch11_adr1[18] ) );
INV_X4 _u0_U17723  ( .A(1'b1), .ZN(_u0_ch11_adr1[17] ) );
INV_X4 _u0_U17721  ( .A(1'b1), .ZN(_u0_ch11_adr1[16] ) );
INV_X4 _u0_U17719  ( .A(1'b1), .ZN(_u0_ch11_adr1[15] ) );
INV_X4 _u0_U17717  ( .A(1'b1), .ZN(_u0_ch11_adr1[14] ) );
INV_X4 _u0_U17715  ( .A(1'b1), .ZN(_u0_ch11_adr1[13] ) );
INV_X4 _u0_U17713  ( .A(1'b1), .ZN(_u0_ch11_adr1[12] ) );
INV_X4 _u0_U17711  ( .A(1'b1), .ZN(_u0_ch11_adr1[11] ) );
INV_X4 _u0_U17709  ( .A(1'b1), .ZN(_u0_ch11_adr1[10] ) );
INV_X4 _u0_U17707  ( .A(1'b1), .ZN(_u0_ch11_adr1[9] ) );
INV_X4 _u0_U17705  ( .A(1'b1), .ZN(_u0_ch11_adr1[8] ) );
INV_X4 _u0_U17703  ( .A(1'b1), .ZN(_u0_ch11_adr1[7] ) );
INV_X4 _u0_U17701  ( .A(1'b1), .ZN(_u0_ch11_adr1[6] ) );
INV_X4 _u0_U17699  ( .A(1'b1), .ZN(_u0_ch11_adr1[5] ) );
INV_X4 _u0_U17697  ( .A(1'b1), .ZN(_u0_ch11_adr1[4] ) );
INV_X4 _u0_U17695  ( .A(1'b1), .ZN(_u0_ch11_adr1[3] ) );
INV_X4 _u0_U17693  ( .A(1'b1), .ZN(_u0_ch11_adr1[2] ) );
INV_X4 _u0_U17691  ( .A(1'b1), .ZN(_u0_ch11_adr1[1] ) );
INV_X4 _u0_U17689  ( .A(1'b1), .ZN(_u0_ch11_adr1[0] ) );
INV_X4 _u0_U17687  ( .A(1'b0), .ZN(_u0_ch11_am0[31] ) );
INV_X4 _u0_U17685  ( .A(1'b0), .ZN(_u0_ch11_am0[30] ) );
INV_X4 _u0_U17683  ( .A(1'b0), .ZN(_u0_ch11_am0[29] ) );
INV_X4 _u0_U17681  ( .A(1'b0), .ZN(_u0_ch11_am0[28] ) );
INV_X4 _u0_U17679  ( .A(1'b0), .ZN(_u0_ch11_am0[27] ) );
INV_X4 _u0_U17677  ( .A(1'b0), .ZN(_u0_ch11_am0[26] ) );
INV_X4 _u0_U17675  ( .A(1'b0), .ZN(_u0_ch11_am0[25] ) );
INV_X4 _u0_U17673  ( .A(1'b0), .ZN(_u0_ch11_am0[24] ) );
INV_X4 _u0_U17671  ( .A(1'b0), .ZN(_u0_ch11_am0[23] ) );
INV_X4 _u0_U17669  ( .A(1'b0), .ZN(_u0_ch11_am0[22] ) );
INV_X4 _u0_U17667  ( .A(1'b0), .ZN(_u0_ch11_am0[21] ) );
INV_X4 _u0_U17665  ( .A(1'b0), .ZN(_u0_ch11_am0[20] ) );
INV_X4 _u0_U17663  ( .A(1'b0), .ZN(_u0_ch11_am0[19] ) );
INV_X4 _u0_U17661  ( .A(1'b0), .ZN(_u0_ch11_am0[18] ) );
INV_X4 _u0_U17659  ( .A(1'b0), .ZN(_u0_ch11_am0[17] ) );
INV_X4 _u0_U17657  ( .A(1'b0), .ZN(_u0_ch11_am0[16] ) );
INV_X4 _u0_U17655  ( .A(1'b0), .ZN(_u0_ch11_am0[15] ) );
INV_X4 _u0_U17653  ( .A(1'b0), .ZN(_u0_ch11_am0[14] ) );
INV_X4 _u0_U17651  ( .A(1'b0), .ZN(_u0_ch11_am0[13] ) );
INV_X4 _u0_U17649  ( .A(1'b0), .ZN(_u0_ch11_am0[12] ) );
INV_X4 _u0_U17647  ( .A(1'b0), .ZN(_u0_ch11_am0[11] ) );
INV_X4 _u0_U17645  ( .A(1'b0), .ZN(_u0_ch11_am0[10] ) );
INV_X4 _u0_U17643  ( .A(1'b0), .ZN(_u0_ch11_am0[9] ) );
INV_X4 _u0_U17641  ( .A(1'b0), .ZN(_u0_ch11_am0[8] ) );
INV_X4 _u0_U17639  ( .A(1'b0), .ZN(_u0_ch11_am0[7] ) );
INV_X4 _u0_U17637  ( .A(1'b0), .ZN(_u0_ch11_am0[6] ) );
INV_X4 _u0_U17635  ( .A(1'b0), .ZN(_u0_ch11_am0[5] ) );
INV_X4 _u0_U17633  ( .A(1'b0), .ZN(_u0_ch11_am0[4] ) );
INV_X4 _u0_U17631  ( .A(1'b1), .ZN(_u0_ch11_am0[3] ) );
INV_X4 _u0_U17629  ( .A(1'b1), .ZN(_u0_ch11_am0[2] ) );
INV_X4 _u0_U17627  ( .A(1'b1), .ZN(_u0_ch11_am0[1] ) );
INV_X4 _u0_U17625  ( .A(1'b1), .ZN(_u0_ch11_am0[0] ) );
INV_X4 _u0_U17623  ( .A(1'b0), .ZN(_u0_ch11_am1[31] ) );
INV_X4 _u0_U17621  ( .A(1'b0), .ZN(_u0_ch11_am1[30] ) );
INV_X4 _u0_U17619  ( .A(1'b0), .ZN(_u0_ch11_am1[29] ) );
INV_X4 _u0_U17617  ( .A(1'b0), .ZN(_u0_ch11_am1[28] ) );
INV_X4 _u0_U17615  ( .A(1'b0), .ZN(_u0_ch11_am1[27] ) );
INV_X4 _u0_U17613  ( .A(1'b0), .ZN(_u0_ch11_am1[26] ) );
INV_X4 _u0_U17611  ( .A(1'b0), .ZN(_u0_ch11_am1[25] ) );
INV_X4 _u0_U17609  ( .A(1'b0), .ZN(_u0_ch11_am1[24] ) );
INV_X4 _u0_U17607  ( .A(1'b0), .ZN(_u0_ch11_am1[23] ) );
INV_X4 _u0_U17605  ( .A(1'b0), .ZN(_u0_ch11_am1[22] ) );
INV_X4 _u0_U17603  ( .A(1'b0), .ZN(_u0_ch11_am1[21] ) );
INV_X4 _u0_U17601  ( .A(1'b0), .ZN(_u0_ch11_am1[20] ) );
INV_X4 _u0_U17599  ( .A(1'b0), .ZN(_u0_ch11_am1[19] ) );
INV_X4 _u0_U17597  ( .A(1'b0), .ZN(_u0_ch11_am1[18] ) );
INV_X4 _u0_U17595  ( .A(1'b0), .ZN(_u0_ch11_am1[17] ) );
INV_X4 _u0_U17593  ( .A(1'b0), .ZN(_u0_ch11_am1[16] ) );
INV_X4 _u0_U17591  ( .A(1'b0), .ZN(_u0_ch11_am1[15] ) );
INV_X4 _u0_U17589  ( .A(1'b0), .ZN(_u0_ch11_am1[14] ) );
INV_X4 _u0_U17587  ( .A(1'b0), .ZN(_u0_ch11_am1[13] ) );
INV_X4 _u0_U17585  ( .A(1'b0), .ZN(_u0_ch11_am1[12] ) );
INV_X4 _u0_U17583  ( .A(1'b0), .ZN(_u0_ch11_am1[11] ) );
INV_X4 _u0_U17581  ( .A(1'b0), .ZN(_u0_ch11_am1[10] ) );
INV_X4 _u0_U17579  ( .A(1'b0), .ZN(_u0_ch11_am1[9] ) );
INV_X4 _u0_U17577  ( .A(1'b0), .ZN(_u0_ch11_am1[8] ) );
INV_X4 _u0_U17575  ( .A(1'b0), .ZN(_u0_ch11_am1[7] ) );
INV_X4 _u0_U17573  ( .A(1'b0), .ZN(_u0_ch11_am1[6] ) );
INV_X4 _u0_U17571  ( .A(1'b0), .ZN(_u0_ch11_am1[5] ) );
INV_X4 _u0_U17569  ( .A(1'b0), .ZN(_u0_ch11_am1[4] ) );
INV_X4 _u0_U17567  ( .A(1'b1), .ZN(_u0_ch11_am1[3] ) );
INV_X4 _u0_U17565  ( .A(1'b1), .ZN(_u0_ch11_am1[2] ) );
INV_X4 _u0_U17563  ( .A(1'b1), .ZN(_u0_ch11_am1[1] ) );
INV_X4 _u0_U17561  ( .A(1'b1), .ZN(_u0_ch11_am1[0] ) );
INV_X4 _u0_U17559  ( .A(1'b1), .ZN(_u0_pointer12[31] ) );
INV_X4 _u0_U17557  ( .A(1'b1), .ZN(_u0_pointer12[30] ) );
INV_X4 _u0_U17555  ( .A(1'b1), .ZN(_u0_pointer12[29] ) );
INV_X4 _u0_U17553  ( .A(1'b1), .ZN(_u0_pointer12[28] ) );
INV_X4 _u0_U17551  ( .A(1'b1), .ZN(_u0_pointer12[27] ) );
INV_X4 _u0_U17549  ( .A(1'b1), .ZN(_u0_pointer12[26] ) );
INV_X4 _u0_U17547  ( .A(1'b1), .ZN(_u0_pointer12[25] ) );
INV_X4 _u0_U17545  ( .A(1'b1), .ZN(_u0_pointer12[24] ) );
INV_X4 _u0_U17543  ( .A(1'b1), .ZN(_u0_pointer12[23] ) );
INV_X4 _u0_U17541  ( .A(1'b1), .ZN(_u0_pointer12[22] ) );
INV_X4 _u0_U17539  ( .A(1'b1), .ZN(_u0_pointer12[21] ) );
INV_X4 _u0_U17537  ( .A(1'b1), .ZN(_u0_pointer12[20] ) );
INV_X4 _u0_U17535  ( .A(1'b1), .ZN(_u0_pointer12[19] ) );
INV_X4 _u0_U17533  ( .A(1'b1), .ZN(_u0_pointer12[18] ) );
INV_X4 _u0_U17531  ( .A(1'b1), .ZN(_u0_pointer12[17] ) );
INV_X4 _u0_U17529  ( .A(1'b1), .ZN(_u0_pointer12[16] ) );
INV_X4 _u0_U17527  ( .A(1'b1), .ZN(_u0_pointer12[15] ) );
INV_X4 _u0_U17525  ( .A(1'b1), .ZN(_u0_pointer12[14] ) );
INV_X4 _u0_U17523  ( .A(1'b1), .ZN(_u0_pointer12[13] ) );
INV_X4 _u0_U17521  ( .A(1'b1), .ZN(_u0_pointer12[12] ) );
INV_X4 _u0_U17519  ( .A(1'b1), .ZN(_u0_pointer12[11] ) );
INV_X4 _u0_U17517  ( .A(1'b1), .ZN(_u0_pointer12[10] ) );
INV_X4 _u0_U17515  ( .A(1'b1), .ZN(_u0_pointer12[9] ) );
INV_X4 _u0_U17513  ( .A(1'b1), .ZN(_u0_pointer12[8] ) );
INV_X4 _u0_U17511  ( .A(1'b1), .ZN(_u0_pointer12[7] ) );
INV_X4 _u0_U17509  ( .A(1'b1), .ZN(_u0_pointer12[6] ) );
INV_X4 _u0_U17507  ( .A(1'b1), .ZN(_u0_pointer12[5] ) );
INV_X4 _u0_U17505  ( .A(1'b1), .ZN(_u0_pointer12[4] ) );
INV_X4 _u0_U17503  ( .A(1'b1), .ZN(_u0_pointer12[3] ) );
INV_X4 _u0_U17501  ( .A(1'b1), .ZN(_u0_pointer12[2] ) );
INV_X4 _u0_U17499  ( .A(1'b1), .ZN(_u0_pointer12[1] ) );
INV_X4 _u0_U17497  ( .A(1'b1), .ZN(_u0_pointer12[0] ) );
INV_X4 _u0_U17495  ( .A(1'b1), .ZN(_u0_pointer12_s[31] ) );
INV_X4 _u0_U17493  ( .A(1'b1), .ZN(_u0_pointer12_s[30] ) );
INV_X4 _u0_U17491  ( .A(1'b1), .ZN(_u0_pointer12_s[29] ) );
INV_X4 _u0_U17489  ( .A(1'b1), .ZN(_u0_pointer12_s[28] ) );
INV_X4 _u0_U17487  ( .A(1'b1), .ZN(_u0_pointer12_s[27] ) );
INV_X4 _u0_U17485  ( .A(1'b1), .ZN(_u0_pointer12_s[26] ) );
INV_X4 _u0_U17483  ( .A(1'b1), .ZN(_u0_pointer12_s[25] ) );
INV_X4 _u0_U17481  ( .A(1'b1), .ZN(_u0_pointer12_s[24] ) );
INV_X4 _u0_U17479  ( .A(1'b1), .ZN(_u0_pointer12_s[23] ) );
INV_X4 _u0_U17477  ( .A(1'b1), .ZN(_u0_pointer12_s[22] ) );
INV_X4 _u0_U17475  ( .A(1'b1), .ZN(_u0_pointer12_s[21] ) );
INV_X4 _u0_U17473  ( .A(1'b1), .ZN(_u0_pointer12_s[20] ) );
INV_X4 _u0_U17471  ( .A(1'b1), .ZN(_u0_pointer12_s[19] ) );
INV_X4 _u0_U17469  ( .A(1'b1), .ZN(_u0_pointer12_s[18] ) );
INV_X4 _u0_U17467  ( .A(1'b1), .ZN(_u0_pointer12_s[17] ) );
INV_X4 _u0_U17465  ( .A(1'b1), .ZN(_u0_pointer12_s[16] ) );
INV_X4 _u0_U17463  ( .A(1'b1), .ZN(_u0_pointer12_s[15] ) );
INV_X4 _u0_U17461  ( .A(1'b1), .ZN(_u0_pointer12_s[14] ) );
INV_X4 _u0_U17459  ( .A(1'b1), .ZN(_u0_pointer12_s[13] ) );
INV_X4 _u0_U17457  ( .A(1'b1), .ZN(_u0_pointer12_s[12] ) );
INV_X4 _u0_U17455  ( .A(1'b1), .ZN(_u0_pointer12_s[11] ) );
INV_X4 _u0_U17453  ( .A(1'b1), .ZN(_u0_pointer12_s[10] ) );
INV_X4 _u0_U17451  ( .A(1'b1), .ZN(_u0_pointer12_s[9] ) );
INV_X4 _u0_U17449  ( .A(1'b1), .ZN(_u0_pointer12_s[8] ) );
INV_X4 _u0_U17447  ( .A(1'b1), .ZN(_u0_pointer12_s[7] ) );
INV_X4 _u0_U17445  ( .A(1'b1), .ZN(_u0_pointer12_s[6] ) );
INV_X4 _u0_U17443  ( .A(1'b1), .ZN(_u0_pointer12_s[5] ) );
INV_X4 _u0_U17441  ( .A(1'b1), .ZN(_u0_pointer12_s[4] ) );
INV_X4 _u0_U17439  ( .A(1'b1), .ZN(_u0_pointer12_s[3] ) );
INV_X4 _u0_U17437  ( .A(1'b1), .ZN(_u0_pointer12_s[2] ) );
INV_X4 _u0_U17435  ( .A(1'b1), .ZN(_u0_pointer12_s[1] ) );
INV_X4 _u0_U17433  ( .A(1'b1), .ZN(_u0_pointer12_s[0] ) );
INV_X4 _u0_U17431  ( .A(1'b1), .ZN(_u0_ch12_csr[31] ) );
INV_X4 _u0_U17429  ( .A(1'b1), .ZN(_u0_ch12_csr[30] ) );
INV_X4 _u0_U17427  ( .A(1'b1), .ZN(_u0_ch12_csr[29] ) );
INV_X4 _u0_U17425  ( .A(1'b1), .ZN(_u0_ch12_csr[28] ) );
INV_X4 _u0_U17423  ( .A(1'b1), .ZN(_u0_ch12_csr[27] ) );
INV_X4 _u0_U17421  ( .A(1'b1), .ZN(_u0_ch12_csr[26] ) );
INV_X4 _u0_U17419  ( .A(1'b1), .ZN(_u0_ch12_csr[25] ) );
INV_X4 _u0_U17417  ( .A(1'b1), .ZN(_u0_ch12_csr[24] ) );
INV_X4 _u0_U17415  ( .A(1'b1), .ZN(_u0_ch12_csr[23] ) );
INV_X4 _u0_U17413  ( .A(1'b1), .ZN(_u0_ch12_csr[22] ) );
INV_X4 _u0_U17411  ( .A(1'b1), .ZN(_u0_ch12_csr[21] ) );
INV_X4 _u0_U17409  ( .A(1'b1), .ZN(_u0_ch12_csr[20] ) );
INV_X4 _u0_U17407  ( .A(1'b1), .ZN(_u0_ch12_csr[19] ) );
INV_X4 _u0_U17405  ( .A(1'b1), .ZN(_u0_ch12_csr[18] ) );
INV_X4 _u0_U17403  ( .A(1'b1), .ZN(_u0_ch12_csr[17] ) );
INV_X4 _u0_U17401  ( .A(1'b1), .ZN(_u0_ch12_csr[16] ) );
INV_X4 _u0_U17399  ( .A(1'b1), .ZN(_u0_ch12_csr[15] ) );
INV_X4 _u0_U17397  ( .A(1'b1), .ZN(_u0_ch12_csr[14] ) );
INV_X4 _u0_U17395  ( .A(1'b1), .ZN(_u0_ch12_csr[13] ) );
INV_X4 _u0_U17393  ( .A(1'b1), .ZN(_u0_ch12_csr[12] ) );
INV_X4 _u0_U17391  ( .A(1'b1), .ZN(_u0_ch12_csr[11] ) );
INV_X4 _u0_U17389  ( .A(1'b1), .ZN(_u0_ch12_csr[10] ) );
INV_X4 _u0_U17387  ( .A(1'b1), .ZN(_u0_ch12_csr[9] ) );
INV_X4 _u0_U17385  ( .A(1'b1), .ZN(_u0_ch12_csr[8] ) );
INV_X4 _u0_U17383  ( .A(1'b1), .ZN(_u0_ch12_csr[7] ) );
INV_X4 _u0_U17381  ( .A(1'b1), .ZN(_u0_ch12_csr[6] ) );
INV_X4 _u0_U17379  ( .A(1'b1), .ZN(_u0_ch12_csr[5] ) );
INV_X4 _u0_U17377  ( .A(1'b1), .ZN(_u0_ch12_csr[4] ) );
INV_X4 _u0_U17375  ( .A(1'b1), .ZN(_u0_ch12_csr[3] ) );
INV_X4 _u0_U17373  ( .A(1'b1), .ZN(_u0_ch12_csr[2] ) );
INV_X4 _u0_U17371  ( .A(1'b1), .ZN(_u0_ch12_csr[1] ) );
INV_X4 _u0_U17369  ( .A(1'b1), .ZN(_u0_ch12_csr[0] ) );
INV_X4 _u0_U17367  ( .A(1'b1), .ZN(_u0_ch12_txsz[31] ) );
INV_X4 _u0_U17365  ( .A(1'b1), .ZN(_u0_ch12_txsz[30] ) );
INV_X4 _u0_U17363  ( .A(1'b1), .ZN(_u0_ch12_txsz[29] ) );
INV_X4 _u0_U17361  ( .A(1'b1), .ZN(_u0_ch12_txsz[28] ) );
INV_X4 _u0_U17359  ( .A(1'b1), .ZN(_u0_ch12_txsz[27] ) );
INV_X4 _u0_U17357  ( .A(1'b1), .ZN(_u0_ch12_txsz[26] ) );
INV_X4 _u0_U17355  ( .A(1'b1), .ZN(_u0_ch12_txsz[25] ) );
INV_X4 _u0_U17353  ( .A(1'b1), .ZN(_u0_ch12_txsz[24] ) );
INV_X4 _u0_U17351  ( .A(1'b1), .ZN(_u0_ch12_txsz[23] ) );
INV_X4 _u0_U17349  ( .A(1'b1), .ZN(_u0_ch12_txsz[22] ) );
INV_X4 _u0_U17347  ( .A(1'b1), .ZN(_u0_ch12_txsz[21] ) );
INV_X4 _u0_U17345  ( .A(1'b1), .ZN(_u0_ch12_txsz[20] ) );
INV_X4 _u0_U17343  ( .A(1'b1), .ZN(_u0_ch12_txsz[19] ) );
INV_X4 _u0_U17341  ( .A(1'b1), .ZN(_u0_ch12_txsz[18] ) );
INV_X4 _u0_U17339  ( .A(1'b1), .ZN(_u0_ch12_txsz[17] ) );
INV_X4 _u0_U17337  ( .A(1'b1), .ZN(_u0_ch12_txsz[16] ) );
INV_X4 _u0_U17335  ( .A(1'b1), .ZN(_u0_ch12_txsz[15] ) );
INV_X4 _u0_U17333  ( .A(1'b1), .ZN(_u0_ch12_txsz[14] ) );
INV_X4 _u0_U17331  ( .A(1'b1), .ZN(_u0_ch12_txsz[13] ) );
INV_X4 _u0_U17329  ( .A(1'b1), .ZN(_u0_ch12_txsz[12] ) );
INV_X4 _u0_U17327  ( .A(1'b1), .ZN(_u0_ch12_txsz[11] ) );
INV_X4 _u0_U17325  ( .A(1'b1), .ZN(_u0_ch12_txsz[10] ) );
INV_X4 _u0_U17323  ( .A(1'b1), .ZN(_u0_ch12_txsz[9] ) );
INV_X4 _u0_U17321  ( .A(1'b1), .ZN(_u0_ch12_txsz[8] ) );
INV_X4 _u0_U17319  ( .A(1'b1), .ZN(_u0_ch12_txsz[7] ) );
INV_X4 _u0_U17317  ( .A(1'b1), .ZN(_u0_ch12_txsz[6] ) );
INV_X4 _u0_U17315  ( .A(1'b1), .ZN(_u0_ch12_txsz[5] ) );
INV_X4 _u0_U17313  ( .A(1'b1), .ZN(_u0_ch12_txsz[4] ) );
INV_X4 _u0_U17311  ( .A(1'b1), .ZN(_u0_ch12_txsz[3] ) );
INV_X4 _u0_U17309  ( .A(1'b1), .ZN(_u0_ch12_txsz[2] ) );
INV_X4 _u0_U17307  ( .A(1'b1), .ZN(_u0_ch12_txsz[1] ) );
INV_X4 _u0_U17305  ( .A(1'b1), .ZN(_u0_ch12_txsz[0] ) );
INV_X4 _u0_U17303  ( .A(1'b1), .ZN(_u0_ch12_adr0[31] ) );
INV_X4 _u0_U17301  ( .A(1'b1), .ZN(_u0_ch12_adr0[30] ) );
INV_X4 _u0_U17299  ( .A(1'b1), .ZN(_u0_ch12_adr0[29] ) );
INV_X4 _u0_U17297  ( .A(1'b1), .ZN(_u0_ch12_adr0[28] ) );
INV_X4 _u0_U17295  ( .A(1'b1), .ZN(_u0_ch12_adr0[27] ) );
INV_X4 _u0_U17293  ( .A(1'b1), .ZN(_u0_ch12_adr0[26] ) );
INV_X4 _u0_U17291  ( .A(1'b1), .ZN(_u0_ch12_adr0[25] ) );
INV_X4 _u0_U17289  ( .A(1'b1), .ZN(_u0_ch12_adr0[24] ) );
INV_X4 _u0_U17287  ( .A(1'b1), .ZN(_u0_ch12_adr0[23] ) );
INV_X4 _u0_U17285  ( .A(1'b1), .ZN(_u0_ch12_adr0[22] ) );
INV_X4 _u0_U17283  ( .A(1'b1), .ZN(_u0_ch12_adr0[21] ) );
INV_X4 _u0_U17281  ( .A(1'b1), .ZN(_u0_ch12_adr0[20] ) );
INV_X4 _u0_U17279  ( .A(1'b1), .ZN(_u0_ch12_adr0[19] ) );
INV_X4 _u0_U17277  ( .A(1'b1), .ZN(_u0_ch12_adr0[18] ) );
INV_X4 _u0_U17275  ( .A(1'b1), .ZN(_u0_ch12_adr0[17] ) );
INV_X4 _u0_U17273  ( .A(1'b1), .ZN(_u0_ch12_adr0[16] ) );
INV_X4 _u0_U17271  ( .A(1'b1), .ZN(_u0_ch12_adr0[15] ) );
INV_X4 _u0_U17269  ( .A(1'b1), .ZN(_u0_ch12_adr0[14] ) );
INV_X4 _u0_U17267  ( .A(1'b1), .ZN(_u0_ch12_adr0[13] ) );
INV_X4 _u0_U17265  ( .A(1'b1), .ZN(_u0_ch12_adr0[12] ) );
INV_X4 _u0_U17263  ( .A(1'b1), .ZN(_u0_ch12_adr0[11] ) );
INV_X4 _u0_U17261  ( .A(1'b1), .ZN(_u0_ch12_adr0[10] ) );
INV_X4 _u0_U17259  ( .A(1'b1), .ZN(_u0_ch12_adr0[9] ) );
INV_X4 _u0_U17257  ( .A(1'b1), .ZN(_u0_ch12_adr0[8] ) );
INV_X4 _u0_U17255  ( .A(1'b1), .ZN(_u0_ch12_adr0[7] ) );
INV_X4 _u0_U17253  ( .A(1'b1), .ZN(_u0_ch12_adr0[6] ) );
INV_X4 _u0_U17251  ( .A(1'b1), .ZN(_u0_ch12_adr0[5] ) );
INV_X4 _u0_U17249  ( .A(1'b1), .ZN(_u0_ch12_adr0[4] ) );
INV_X4 _u0_U17247  ( .A(1'b1), .ZN(_u0_ch12_adr0[3] ) );
INV_X4 _u0_U17245  ( .A(1'b1), .ZN(_u0_ch12_adr0[2] ) );
INV_X4 _u0_U17243  ( .A(1'b1), .ZN(_u0_ch12_adr0[1] ) );
INV_X4 _u0_U17241  ( .A(1'b1), .ZN(_u0_ch12_adr0[0] ) );
INV_X4 _u0_U17239  ( .A(1'b1), .ZN(_u0_ch12_adr1[31] ) );
INV_X4 _u0_U17237  ( .A(1'b1), .ZN(_u0_ch12_adr1[30] ) );
INV_X4 _u0_U17235  ( .A(1'b1), .ZN(_u0_ch12_adr1[29] ) );
INV_X4 _u0_U17233  ( .A(1'b1), .ZN(_u0_ch12_adr1[28] ) );
INV_X4 _u0_U17231  ( .A(1'b1), .ZN(_u0_ch12_adr1[27] ) );
INV_X4 _u0_U17229  ( .A(1'b1), .ZN(_u0_ch12_adr1[26] ) );
INV_X4 _u0_U17227  ( .A(1'b1), .ZN(_u0_ch12_adr1[25] ) );
INV_X4 _u0_U17225  ( .A(1'b1), .ZN(_u0_ch12_adr1[24] ) );
INV_X4 _u0_U17223  ( .A(1'b1), .ZN(_u0_ch12_adr1[23] ) );
INV_X4 _u0_U17221  ( .A(1'b1), .ZN(_u0_ch12_adr1[22] ) );
INV_X4 _u0_U17219  ( .A(1'b1), .ZN(_u0_ch12_adr1[21] ) );
INV_X4 _u0_U17217  ( .A(1'b1), .ZN(_u0_ch12_adr1[20] ) );
INV_X4 _u0_U17215  ( .A(1'b1), .ZN(_u0_ch12_adr1[19] ) );
INV_X4 _u0_U17213  ( .A(1'b1), .ZN(_u0_ch12_adr1[18] ) );
INV_X4 _u0_U17211  ( .A(1'b1), .ZN(_u0_ch12_adr1[17] ) );
INV_X4 _u0_U17209  ( .A(1'b1), .ZN(_u0_ch12_adr1[16] ) );
INV_X4 _u0_U17207  ( .A(1'b1), .ZN(_u0_ch12_adr1[15] ) );
INV_X4 _u0_U17205  ( .A(1'b1), .ZN(_u0_ch12_adr1[14] ) );
INV_X4 _u0_U17203  ( .A(1'b1), .ZN(_u0_ch12_adr1[13] ) );
INV_X4 _u0_U17201  ( .A(1'b1), .ZN(_u0_ch12_adr1[12] ) );
INV_X4 _u0_U17199  ( .A(1'b1), .ZN(_u0_ch12_adr1[11] ) );
INV_X4 _u0_U17197  ( .A(1'b1), .ZN(_u0_ch12_adr1[10] ) );
INV_X4 _u0_U17195  ( .A(1'b1), .ZN(_u0_ch12_adr1[9] ) );
INV_X4 _u0_U17193  ( .A(1'b1), .ZN(_u0_ch12_adr1[8] ) );
INV_X4 _u0_U17191  ( .A(1'b1), .ZN(_u0_ch12_adr1[7] ) );
INV_X4 _u0_U17189  ( .A(1'b1), .ZN(_u0_ch12_adr1[6] ) );
INV_X4 _u0_U17187  ( .A(1'b1), .ZN(_u0_ch12_adr1[5] ) );
INV_X4 _u0_U17185  ( .A(1'b1), .ZN(_u0_ch12_adr1[4] ) );
INV_X4 _u0_U17183  ( .A(1'b1), .ZN(_u0_ch12_adr1[3] ) );
INV_X4 _u0_U17181  ( .A(1'b1), .ZN(_u0_ch12_adr1[2] ) );
INV_X4 _u0_U17179  ( .A(1'b1), .ZN(_u0_ch12_adr1[1] ) );
INV_X4 _u0_U17177  ( .A(1'b1), .ZN(_u0_ch12_adr1[0] ) );
INV_X4 _u0_U17175  ( .A(1'b0), .ZN(_u0_ch12_am0[31] ) );
INV_X4 _u0_U17173  ( .A(1'b0), .ZN(_u0_ch12_am0[30] ) );
INV_X4 _u0_U17171  ( .A(1'b0), .ZN(_u0_ch12_am0[29] ) );
INV_X4 _u0_U17169  ( .A(1'b0), .ZN(_u0_ch12_am0[28] ) );
INV_X4 _u0_U17167  ( .A(1'b0), .ZN(_u0_ch12_am0[27] ) );
INV_X4 _u0_U17165  ( .A(1'b0), .ZN(_u0_ch12_am0[26] ) );
INV_X4 _u0_U17163  ( .A(1'b0), .ZN(_u0_ch12_am0[25] ) );
INV_X4 _u0_U17161  ( .A(1'b0), .ZN(_u0_ch12_am0[24] ) );
INV_X4 _u0_U17159  ( .A(1'b0), .ZN(_u0_ch12_am0[23] ) );
INV_X4 _u0_U17157  ( .A(1'b0), .ZN(_u0_ch12_am0[22] ) );
INV_X4 _u0_U17155  ( .A(1'b0), .ZN(_u0_ch12_am0[21] ) );
INV_X4 _u0_U17153  ( .A(1'b0), .ZN(_u0_ch12_am0[20] ) );
INV_X4 _u0_U17151  ( .A(1'b0), .ZN(_u0_ch12_am0[19] ) );
INV_X4 _u0_U17149  ( .A(1'b0), .ZN(_u0_ch12_am0[18] ) );
INV_X4 _u0_U17147  ( .A(1'b0), .ZN(_u0_ch12_am0[17] ) );
INV_X4 _u0_U17145  ( .A(1'b0), .ZN(_u0_ch12_am0[16] ) );
INV_X4 _u0_U17143  ( .A(1'b0), .ZN(_u0_ch12_am0[15] ) );
INV_X4 _u0_U17141  ( .A(1'b0), .ZN(_u0_ch12_am0[14] ) );
INV_X4 _u0_U17139  ( .A(1'b0), .ZN(_u0_ch12_am0[13] ) );
INV_X4 _u0_U17137  ( .A(1'b0), .ZN(_u0_ch12_am0[12] ) );
INV_X4 _u0_U17135  ( .A(1'b0), .ZN(_u0_ch12_am0[11] ) );
INV_X4 _u0_U17133  ( .A(1'b0), .ZN(_u0_ch12_am0[10] ) );
INV_X4 _u0_U17131  ( .A(1'b0), .ZN(_u0_ch12_am0[9] ) );
INV_X4 _u0_U17129  ( .A(1'b0), .ZN(_u0_ch12_am0[8] ) );
INV_X4 _u0_U17127  ( .A(1'b0), .ZN(_u0_ch12_am0[7] ) );
INV_X4 _u0_U17125  ( .A(1'b0), .ZN(_u0_ch12_am0[6] ) );
INV_X4 _u0_U17123  ( .A(1'b0), .ZN(_u0_ch12_am0[5] ) );
INV_X4 _u0_U17121  ( .A(1'b0), .ZN(_u0_ch12_am0[4] ) );
INV_X4 _u0_U17119  ( .A(1'b1), .ZN(_u0_ch12_am0[3] ) );
INV_X4 _u0_U17117  ( .A(1'b1), .ZN(_u0_ch12_am0[2] ) );
INV_X4 _u0_U17115  ( .A(1'b1), .ZN(_u0_ch12_am0[1] ) );
INV_X4 _u0_U17113  ( .A(1'b1), .ZN(_u0_ch12_am0[0] ) );
INV_X4 _u0_U17111  ( .A(1'b0), .ZN(_u0_ch12_am1[31] ) );
INV_X4 _u0_U17109  ( .A(1'b0), .ZN(_u0_ch12_am1[30] ) );
INV_X4 _u0_U17107  ( .A(1'b0), .ZN(_u0_ch12_am1[29] ) );
INV_X4 _u0_U17105  ( .A(1'b0), .ZN(_u0_ch12_am1[28] ) );
INV_X4 _u0_U17103  ( .A(1'b0), .ZN(_u0_ch12_am1[27] ) );
INV_X4 _u0_U17101  ( .A(1'b0), .ZN(_u0_ch12_am1[26] ) );
INV_X4 _u0_U17099  ( .A(1'b0), .ZN(_u0_ch12_am1[25] ) );
INV_X4 _u0_U17097  ( .A(1'b0), .ZN(_u0_ch12_am1[24] ) );
INV_X4 _u0_U17095  ( .A(1'b0), .ZN(_u0_ch12_am1[23] ) );
INV_X4 _u0_U17093  ( .A(1'b0), .ZN(_u0_ch12_am1[22] ) );
INV_X4 _u0_U17091  ( .A(1'b0), .ZN(_u0_ch12_am1[21] ) );
INV_X4 _u0_U17089  ( .A(1'b0), .ZN(_u0_ch12_am1[20] ) );
INV_X4 _u0_U17087  ( .A(1'b0), .ZN(_u0_ch12_am1[19] ) );
INV_X4 _u0_U17085  ( .A(1'b0), .ZN(_u0_ch12_am1[18] ) );
INV_X4 _u0_U17083  ( .A(1'b0), .ZN(_u0_ch12_am1[17] ) );
INV_X4 _u0_U17081  ( .A(1'b0), .ZN(_u0_ch12_am1[16] ) );
INV_X4 _u0_U17079  ( .A(1'b0), .ZN(_u0_ch12_am1[15] ) );
INV_X4 _u0_U17077  ( .A(1'b0), .ZN(_u0_ch12_am1[14] ) );
INV_X4 _u0_U17075  ( .A(1'b0), .ZN(_u0_ch12_am1[13] ) );
INV_X4 _u0_U17073  ( .A(1'b0), .ZN(_u0_ch12_am1[12] ) );
INV_X4 _u0_U17071  ( .A(1'b0), .ZN(_u0_ch12_am1[11] ) );
INV_X4 _u0_U17069  ( .A(1'b0), .ZN(_u0_ch12_am1[10] ) );
INV_X4 _u0_U17067  ( .A(1'b0), .ZN(_u0_ch12_am1[9] ) );
INV_X4 _u0_U17065  ( .A(1'b0), .ZN(_u0_ch12_am1[8] ) );
INV_X4 _u0_U17063  ( .A(1'b0), .ZN(_u0_ch12_am1[7] ) );
INV_X4 _u0_U17061  ( .A(1'b0), .ZN(_u0_ch12_am1[6] ) );
INV_X4 _u0_U17059  ( .A(1'b0), .ZN(_u0_ch12_am1[5] ) );
INV_X4 _u0_U17057  ( .A(1'b0), .ZN(_u0_ch12_am1[4] ) );
INV_X4 _u0_U17055  ( .A(1'b1), .ZN(_u0_ch12_am1[3] ) );
INV_X4 _u0_U17053  ( .A(1'b1), .ZN(_u0_ch12_am1[2] ) );
INV_X4 _u0_U17051  ( .A(1'b1), .ZN(_u0_ch12_am1[1] ) );
INV_X4 _u0_U17049  ( .A(1'b1), .ZN(_u0_ch12_am1[0] ) );
INV_X4 _u0_U17047  ( .A(1'b1), .ZN(_u0_pointer13[31] ) );
INV_X4 _u0_U17045  ( .A(1'b1), .ZN(_u0_pointer13[30] ) );
INV_X4 _u0_U17043  ( .A(1'b1), .ZN(_u0_pointer13[29] ) );
INV_X4 _u0_U17041  ( .A(1'b1), .ZN(_u0_pointer13[28] ) );
INV_X4 _u0_U17039  ( .A(1'b1), .ZN(_u0_pointer13[27] ) );
INV_X4 _u0_U17037  ( .A(1'b1), .ZN(_u0_pointer13[26] ) );
INV_X4 _u0_U17035  ( .A(1'b1), .ZN(_u0_pointer13[25] ) );
INV_X4 _u0_U17033  ( .A(1'b1), .ZN(_u0_pointer13[24] ) );
INV_X4 _u0_U17031  ( .A(1'b1), .ZN(_u0_pointer13[23] ) );
INV_X4 _u0_U17029  ( .A(1'b1), .ZN(_u0_pointer13[22] ) );
INV_X4 _u0_U17027  ( .A(1'b1), .ZN(_u0_pointer13[21] ) );
INV_X4 _u0_U17025  ( .A(1'b1), .ZN(_u0_pointer13[20] ) );
INV_X4 _u0_U17023  ( .A(1'b1), .ZN(_u0_pointer13[19] ) );
INV_X4 _u0_U17021  ( .A(1'b1), .ZN(_u0_pointer13[18] ) );
INV_X4 _u0_U17019  ( .A(1'b1), .ZN(_u0_pointer13[17] ) );
INV_X4 _u0_U17017  ( .A(1'b1), .ZN(_u0_pointer13[16] ) );
INV_X4 _u0_U17015  ( .A(1'b1), .ZN(_u0_pointer13[15] ) );
INV_X4 _u0_U17013  ( .A(1'b1), .ZN(_u0_pointer13[14] ) );
INV_X4 _u0_U17011  ( .A(1'b1), .ZN(_u0_pointer13[13] ) );
INV_X4 _u0_U17009  ( .A(1'b1), .ZN(_u0_pointer13[12] ) );
INV_X4 _u0_U17007  ( .A(1'b1), .ZN(_u0_pointer13[11] ) );
INV_X4 _u0_U17005  ( .A(1'b1), .ZN(_u0_pointer13[10] ) );
INV_X4 _u0_U17003  ( .A(1'b1), .ZN(_u0_pointer13[9] ) );
INV_X4 _u0_U17001  ( .A(1'b1), .ZN(_u0_pointer13[8] ) );
INV_X4 _u0_U16999  ( .A(1'b1), .ZN(_u0_pointer13[7] ) );
INV_X4 _u0_U16997  ( .A(1'b1), .ZN(_u0_pointer13[6] ) );
INV_X4 _u0_U16995  ( .A(1'b1), .ZN(_u0_pointer13[5] ) );
INV_X4 _u0_U16993  ( .A(1'b1), .ZN(_u0_pointer13[4] ) );
INV_X4 _u0_U16991  ( .A(1'b1), .ZN(_u0_pointer13[3] ) );
INV_X4 _u0_U16989  ( .A(1'b1), .ZN(_u0_pointer13[2] ) );
INV_X4 _u0_U16987  ( .A(1'b1), .ZN(_u0_pointer13[1] ) );
INV_X4 _u0_U16985  ( .A(1'b1), .ZN(_u0_pointer13[0] ) );
INV_X4 _u0_U16983  ( .A(1'b1), .ZN(_u0_pointer13_s[31] ) );
INV_X4 _u0_U16981  ( .A(1'b1), .ZN(_u0_pointer13_s[30] ) );
INV_X4 _u0_U16979  ( .A(1'b1), .ZN(_u0_pointer13_s[29] ) );
INV_X4 _u0_U16977  ( .A(1'b1), .ZN(_u0_pointer13_s[28] ) );
INV_X4 _u0_U16975  ( .A(1'b1), .ZN(_u0_pointer13_s[27] ) );
INV_X4 _u0_U16973  ( .A(1'b1), .ZN(_u0_pointer13_s[26] ) );
INV_X4 _u0_U16971  ( .A(1'b1), .ZN(_u0_pointer13_s[25] ) );
INV_X4 _u0_U16969  ( .A(1'b1), .ZN(_u0_pointer13_s[24] ) );
INV_X4 _u0_U16967  ( .A(1'b1), .ZN(_u0_pointer13_s[23] ) );
INV_X4 _u0_U16965  ( .A(1'b1), .ZN(_u0_pointer13_s[22] ) );
INV_X4 _u0_U16963  ( .A(1'b1), .ZN(_u0_pointer13_s[21] ) );
INV_X4 _u0_U16961  ( .A(1'b1), .ZN(_u0_pointer13_s[20] ) );
INV_X4 _u0_U16959  ( .A(1'b1), .ZN(_u0_pointer13_s[19] ) );
INV_X4 _u0_U16957  ( .A(1'b1), .ZN(_u0_pointer13_s[18] ) );
INV_X4 _u0_U16955  ( .A(1'b1), .ZN(_u0_pointer13_s[17] ) );
INV_X4 _u0_U16953  ( .A(1'b1), .ZN(_u0_pointer13_s[16] ) );
INV_X4 _u0_U16951  ( .A(1'b1), .ZN(_u0_pointer13_s[15] ) );
INV_X4 _u0_U16949  ( .A(1'b1), .ZN(_u0_pointer13_s[14] ) );
INV_X4 _u0_U16947  ( .A(1'b1), .ZN(_u0_pointer13_s[13] ) );
INV_X4 _u0_U16945  ( .A(1'b1), .ZN(_u0_pointer13_s[12] ) );
INV_X4 _u0_U16943  ( .A(1'b1), .ZN(_u0_pointer13_s[11] ) );
INV_X4 _u0_U16941  ( .A(1'b1), .ZN(_u0_pointer13_s[10] ) );
INV_X4 _u0_U16939  ( .A(1'b1), .ZN(_u0_pointer13_s[9] ) );
INV_X4 _u0_U16937  ( .A(1'b1), .ZN(_u0_pointer13_s[8] ) );
INV_X4 _u0_U16935  ( .A(1'b1), .ZN(_u0_pointer13_s[7] ) );
INV_X4 _u0_U16933  ( .A(1'b1), .ZN(_u0_pointer13_s[6] ) );
INV_X4 _u0_U16931  ( .A(1'b1), .ZN(_u0_pointer13_s[5] ) );
INV_X4 _u0_U16929  ( .A(1'b1), .ZN(_u0_pointer13_s[4] ) );
INV_X4 _u0_U16927  ( .A(1'b1), .ZN(_u0_pointer13_s[3] ) );
INV_X4 _u0_U16925  ( .A(1'b1), .ZN(_u0_pointer13_s[2] ) );
INV_X4 _u0_U16923  ( .A(1'b1), .ZN(_u0_pointer13_s[1] ) );
INV_X4 _u0_U16921  ( .A(1'b1), .ZN(_u0_pointer13_s[0] ) );
INV_X4 _u0_U16919  ( .A(1'b1), .ZN(_u0_ch13_csr[31] ) );
INV_X4 _u0_U16917  ( .A(1'b1), .ZN(_u0_ch13_csr[30] ) );
INV_X4 _u0_U16915  ( .A(1'b1), .ZN(_u0_ch13_csr[29] ) );
INV_X4 _u0_U16913  ( .A(1'b1), .ZN(_u0_ch13_csr[28] ) );
INV_X4 _u0_U16911  ( .A(1'b1), .ZN(_u0_ch13_csr[27] ) );
INV_X4 _u0_U16909  ( .A(1'b1), .ZN(_u0_ch13_csr[26] ) );
INV_X4 _u0_U16907  ( .A(1'b1), .ZN(_u0_ch13_csr[25] ) );
INV_X4 _u0_U16905  ( .A(1'b1), .ZN(_u0_ch13_csr[24] ) );
INV_X4 _u0_U16903  ( .A(1'b1), .ZN(_u0_ch13_csr[23] ) );
INV_X4 _u0_U16901  ( .A(1'b1), .ZN(_u0_ch13_csr[22] ) );
INV_X4 _u0_U16899  ( .A(1'b1), .ZN(_u0_ch13_csr[21] ) );
INV_X4 _u0_U16897  ( .A(1'b1), .ZN(_u0_ch13_csr[20] ) );
INV_X4 _u0_U16895  ( .A(1'b1), .ZN(_u0_ch13_csr[19] ) );
INV_X4 _u0_U16893  ( .A(1'b1), .ZN(_u0_ch13_csr[18] ) );
INV_X4 _u0_U16891  ( .A(1'b1), .ZN(_u0_ch13_csr[17] ) );
INV_X4 _u0_U16889  ( .A(1'b1), .ZN(_u0_ch13_csr[16] ) );
INV_X4 _u0_U16887  ( .A(1'b1), .ZN(_u0_ch13_csr[15] ) );
INV_X4 _u0_U16885  ( .A(1'b1), .ZN(_u0_ch13_csr[14] ) );
INV_X4 _u0_U16883  ( .A(1'b1), .ZN(_u0_ch13_csr[13] ) );
INV_X4 _u0_U16881  ( .A(1'b1), .ZN(_u0_ch13_csr[12] ) );
INV_X4 _u0_U16879  ( .A(1'b1), .ZN(_u0_ch13_csr[11] ) );
INV_X4 _u0_U16877  ( .A(1'b1), .ZN(_u0_ch13_csr[10] ) );
INV_X4 _u0_U16875  ( .A(1'b1), .ZN(_u0_ch13_csr[9] ) );
INV_X4 _u0_U16873  ( .A(1'b1), .ZN(_u0_ch13_csr[8] ) );
INV_X4 _u0_U16871  ( .A(1'b1), .ZN(_u0_ch13_csr[7] ) );
INV_X4 _u0_U16869  ( .A(1'b1), .ZN(_u0_ch13_csr[6] ) );
INV_X4 _u0_U16867  ( .A(1'b1), .ZN(_u0_ch13_csr[5] ) );
INV_X4 _u0_U16865  ( .A(1'b1), .ZN(_u0_ch13_csr[4] ) );
INV_X4 _u0_U16863  ( .A(1'b1), .ZN(_u0_ch13_csr[3] ) );
INV_X4 _u0_U16861  ( .A(1'b1), .ZN(_u0_ch13_csr[2] ) );
INV_X4 _u0_U16859  ( .A(1'b1), .ZN(_u0_ch13_csr[1] ) );
INV_X4 _u0_U16857  ( .A(1'b1), .ZN(_u0_ch13_csr[0] ) );
INV_X4 _u0_U16855  ( .A(1'b1), .ZN(_u0_ch13_txsz[31] ) );
INV_X4 _u0_U16853  ( .A(1'b1), .ZN(_u0_ch13_txsz[30] ) );
INV_X4 _u0_U16851  ( .A(1'b1), .ZN(_u0_ch13_txsz[29] ) );
INV_X4 _u0_U16849  ( .A(1'b1), .ZN(_u0_ch13_txsz[28] ) );
INV_X4 _u0_U16847  ( .A(1'b1), .ZN(_u0_ch13_txsz[27] ) );
INV_X4 _u0_U16845  ( .A(1'b1), .ZN(_u0_ch13_txsz[26] ) );
INV_X4 _u0_U16843  ( .A(1'b1), .ZN(_u0_ch13_txsz[25] ) );
INV_X4 _u0_U16841  ( .A(1'b1), .ZN(_u0_ch13_txsz[24] ) );
INV_X4 _u0_U16839  ( .A(1'b1), .ZN(_u0_ch13_txsz[23] ) );
INV_X4 _u0_U16837  ( .A(1'b1), .ZN(_u0_ch13_txsz[22] ) );
INV_X4 _u0_U16835  ( .A(1'b1), .ZN(_u0_ch13_txsz[21] ) );
INV_X4 _u0_U16833  ( .A(1'b1), .ZN(_u0_ch13_txsz[20] ) );
INV_X4 _u0_U16831  ( .A(1'b1), .ZN(_u0_ch13_txsz[19] ) );
INV_X4 _u0_U16829  ( .A(1'b1), .ZN(_u0_ch13_txsz[18] ) );
INV_X4 _u0_U16827  ( .A(1'b1), .ZN(_u0_ch13_txsz[17] ) );
INV_X4 _u0_U16825  ( .A(1'b1), .ZN(_u0_ch13_txsz[16] ) );
INV_X4 _u0_U16823  ( .A(1'b1), .ZN(_u0_ch13_txsz[15] ) );
INV_X4 _u0_U16821  ( .A(1'b1), .ZN(_u0_ch13_txsz[14] ) );
INV_X4 _u0_U16819  ( .A(1'b1), .ZN(_u0_ch13_txsz[13] ) );
INV_X4 _u0_U16817  ( .A(1'b1), .ZN(_u0_ch13_txsz[12] ) );
INV_X4 _u0_U16815  ( .A(1'b1), .ZN(_u0_ch13_txsz[11] ) );
INV_X4 _u0_U16813  ( .A(1'b1), .ZN(_u0_ch13_txsz[10] ) );
INV_X4 _u0_U16811  ( .A(1'b1), .ZN(_u0_ch13_txsz[9] ) );
INV_X4 _u0_U16809  ( .A(1'b1), .ZN(_u0_ch13_txsz[8] ) );
INV_X4 _u0_U16807  ( .A(1'b1), .ZN(_u0_ch13_txsz[7] ) );
INV_X4 _u0_U16805  ( .A(1'b1), .ZN(_u0_ch13_txsz[6] ) );
INV_X4 _u0_U16803  ( .A(1'b1), .ZN(_u0_ch13_txsz[5] ) );
INV_X4 _u0_U16801  ( .A(1'b1), .ZN(_u0_ch13_txsz[4] ) );
INV_X4 _u0_U16799  ( .A(1'b1), .ZN(_u0_ch13_txsz[3] ) );
INV_X4 _u0_U16797  ( .A(1'b1), .ZN(_u0_ch13_txsz[2] ) );
INV_X4 _u0_U16795  ( .A(1'b1), .ZN(_u0_ch13_txsz[1] ) );
INV_X4 _u0_U16793  ( .A(1'b1), .ZN(_u0_ch13_txsz[0] ) );
INV_X4 _u0_U16791  ( .A(1'b1), .ZN(_u0_ch13_adr0[31] ) );
INV_X4 _u0_U16789  ( .A(1'b1), .ZN(_u0_ch13_adr0[30] ) );
INV_X4 _u0_U16787  ( .A(1'b1), .ZN(_u0_ch13_adr0[29] ) );
INV_X4 _u0_U16785  ( .A(1'b1), .ZN(_u0_ch13_adr0[28] ) );
INV_X4 _u0_U16783  ( .A(1'b1), .ZN(_u0_ch13_adr0[27] ) );
INV_X4 _u0_U16781  ( .A(1'b1), .ZN(_u0_ch13_adr0[26] ) );
INV_X4 _u0_U16779  ( .A(1'b1), .ZN(_u0_ch13_adr0[25] ) );
INV_X4 _u0_U16777  ( .A(1'b1), .ZN(_u0_ch13_adr0[24] ) );
INV_X4 _u0_U16775  ( .A(1'b1), .ZN(_u0_ch13_adr0[23] ) );
INV_X4 _u0_U16773  ( .A(1'b1), .ZN(_u0_ch13_adr0[22] ) );
INV_X4 _u0_U16771  ( .A(1'b1), .ZN(_u0_ch13_adr0[21] ) );
INV_X4 _u0_U16769  ( .A(1'b1), .ZN(_u0_ch13_adr0[20] ) );
INV_X4 _u0_U16767  ( .A(1'b1), .ZN(_u0_ch13_adr0[19] ) );
INV_X4 _u0_U16765  ( .A(1'b1), .ZN(_u0_ch13_adr0[18] ) );
INV_X4 _u0_U16763  ( .A(1'b1), .ZN(_u0_ch13_adr0[17] ) );
INV_X4 _u0_U16761  ( .A(1'b1), .ZN(_u0_ch13_adr0[16] ) );
INV_X4 _u0_U16759  ( .A(1'b1), .ZN(_u0_ch13_adr0[15] ) );
INV_X4 _u0_U16757  ( .A(1'b1), .ZN(_u0_ch13_adr0[14] ) );
INV_X4 _u0_U16755  ( .A(1'b1), .ZN(_u0_ch13_adr0[13] ) );
INV_X4 _u0_U16753  ( .A(1'b1), .ZN(_u0_ch13_adr0[12] ) );
INV_X4 _u0_U16751  ( .A(1'b1), .ZN(_u0_ch13_adr0[11] ) );
INV_X4 _u0_U16749  ( .A(1'b1), .ZN(_u0_ch13_adr0[10] ) );
INV_X4 _u0_U16747  ( .A(1'b1), .ZN(_u0_ch13_adr0[9] ) );
INV_X4 _u0_U16745  ( .A(1'b1), .ZN(_u0_ch13_adr0[8] ) );
INV_X4 _u0_U16743  ( .A(1'b1), .ZN(_u0_ch13_adr0[7] ) );
INV_X4 _u0_U16741  ( .A(1'b1), .ZN(_u0_ch13_adr0[6] ) );
INV_X4 _u0_U16739  ( .A(1'b1), .ZN(_u0_ch13_adr0[5] ) );
INV_X4 _u0_U16737  ( .A(1'b1), .ZN(_u0_ch13_adr0[4] ) );
INV_X4 _u0_U16735  ( .A(1'b1), .ZN(_u0_ch13_adr0[3] ) );
INV_X4 _u0_U16733  ( .A(1'b1), .ZN(_u0_ch13_adr0[2] ) );
INV_X4 _u0_U16731  ( .A(1'b1), .ZN(_u0_ch13_adr0[1] ) );
INV_X4 _u0_U16729  ( .A(1'b1), .ZN(_u0_ch13_adr0[0] ) );
INV_X4 _u0_U16727  ( .A(1'b1), .ZN(_u0_ch13_adr1[31] ) );
INV_X4 _u0_U16725  ( .A(1'b1), .ZN(_u0_ch13_adr1[30] ) );
INV_X4 _u0_U16723  ( .A(1'b1), .ZN(_u0_ch13_adr1[29] ) );
INV_X4 _u0_U16721  ( .A(1'b1), .ZN(_u0_ch13_adr1[28] ) );
INV_X4 _u0_U16719  ( .A(1'b1), .ZN(_u0_ch13_adr1[27] ) );
INV_X4 _u0_U16717  ( .A(1'b1), .ZN(_u0_ch13_adr1[26] ) );
INV_X4 _u0_U16715  ( .A(1'b1), .ZN(_u0_ch13_adr1[25] ) );
INV_X4 _u0_U16713  ( .A(1'b1), .ZN(_u0_ch13_adr1[24] ) );
INV_X4 _u0_U16711  ( .A(1'b1), .ZN(_u0_ch13_adr1[23] ) );
INV_X4 _u0_U16709  ( .A(1'b1), .ZN(_u0_ch13_adr1[22] ) );
INV_X4 _u0_U16707  ( .A(1'b1), .ZN(_u0_ch13_adr1[21] ) );
INV_X4 _u0_U16705  ( .A(1'b1), .ZN(_u0_ch13_adr1[20] ) );
INV_X4 _u0_U16703  ( .A(1'b1), .ZN(_u0_ch13_adr1[19] ) );
INV_X4 _u0_U16701  ( .A(1'b1), .ZN(_u0_ch13_adr1[18] ) );
INV_X4 _u0_U16699  ( .A(1'b1), .ZN(_u0_ch13_adr1[17] ) );
INV_X4 _u0_U16697  ( .A(1'b1), .ZN(_u0_ch13_adr1[16] ) );
INV_X4 _u0_U16695  ( .A(1'b1), .ZN(_u0_ch13_adr1[15] ) );
INV_X4 _u0_U16693  ( .A(1'b1), .ZN(_u0_ch13_adr1[14] ) );
INV_X4 _u0_U16691  ( .A(1'b1), .ZN(_u0_ch13_adr1[13] ) );
INV_X4 _u0_U16689  ( .A(1'b1), .ZN(_u0_ch13_adr1[12] ) );
INV_X4 _u0_U16687  ( .A(1'b1), .ZN(_u0_ch13_adr1[11] ) );
INV_X4 _u0_U16685  ( .A(1'b1), .ZN(_u0_ch13_adr1[10] ) );
INV_X4 _u0_U16683  ( .A(1'b1), .ZN(_u0_ch13_adr1[9] ) );
INV_X4 _u0_U16681  ( .A(1'b1), .ZN(_u0_ch13_adr1[8] ) );
INV_X4 _u0_U16679  ( .A(1'b1), .ZN(_u0_ch13_adr1[7] ) );
INV_X4 _u0_U16677  ( .A(1'b1), .ZN(_u0_ch13_adr1[6] ) );
INV_X4 _u0_U16675  ( .A(1'b1), .ZN(_u0_ch13_adr1[5] ) );
INV_X4 _u0_U16673  ( .A(1'b1), .ZN(_u0_ch13_adr1[4] ) );
INV_X4 _u0_U16671  ( .A(1'b1), .ZN(_u0_ch13_adr1[3] ) );
INV_X4 _u0_U16669  ( .A(1'b1), .ZN(_u0_ch13_adr1[2] ) );
INV_X4 _u0_U16667  ( .A(1'b1), .ZN(_u0_ch13_adr1[1] ) );
INV_X4 _u0_U16665  ( .A(1'b1), .ZN(_u0_ch13_adr1[0] ) );
INV_X4 _u0_U16663  ( .A(1'b0), .ZN(_u0_ch13_am0[31] ) );
INV_X4 _u0_U16661  ( .A(1'b0), .ZN(_u0_ch13_am0[30] ) );
INV_X4 _u0_U16659  ( .A(1'b0), .ZN(_u0_ch13_am0[29] ) );
INV_X4 _u0_U16657  ( .A(1'b0), .ZN(_u0_ch13_am0[28] ) );
INV_X4 _u0_U16655  ( .A(1'b0), .ZN(_u0_ch13_am0[27] ) );
INV_X4 _u0_U16653  ( .A(1'b0), .ZN(_u0_ch13_am0[26] ) );
INV_X4 _u0_U16651  ( .A(1'b0), .ZN(_u0_ch13_am0[25] ) );
INV_X4 _u0_U16649  ( .A(1'b0), .ZN(_u0_ch13_am0[24] ) );
INV_X4 _u0_U16647  ( .A(1'b0), .ZN(_u0_ch13_am0[23] ) );
INV_X4 _u0_U16645  ( .A(1'b0), .ZN(_u0_ch13_am0[22] ) );
INV_X4 _u0_U16643  ( .A(1'b0), .ZN(_u0_ch13_am0[21] ) );
INV_X4 _u0_U16641  ( .A(1'b0), .ZN(_u0_ch13_am0[20] ) );
INV_X4 _u0_U16639  ( .A(1'b0), .ZN(_u0_ch13_am0[19] ) );
INV_X4 _u0_U16637  ( .A(1'b0), .ZN(_u0_ch13_am0[18] ) );
INV_X4 _u0_U16635  ( .A(1'b0), .ZN(_u0_ch13_am0[17] ) );
INV_X4 _u0_U16633  ( .A(1'b0), .ZN(_u0_ch13_am0[16] ) );
INV_X4 _u0_U16631  ( .A(1'b0), .ZN(_u0_ch13_am0[15] ) );
INV_X4 _u0_U16629  ( .A(1'b0), .ZN(_u0_ch13_am0[14] ) );
INV_X4 _u0_U16627  ( .A(1'b0), .ZN(_u0_ch13_am0[13] ) );
INV_X4 _u0_U16625  ( .A(1'b0), .ZN(_u0_ch13_am0[12] ) );
INV_X4 _u0_U16623  ( .A(1'b0), .ZN(_u0_ch13_am0[11] ) );
INV_X4 _u0_U16621  ( .A(1'b0), .ZN(_u0_ch13_am0[10] ) );
INV_X4 _u0_U16619  ( .A(1'b0), .ZN(_u0_ch13_am0[9] ) );
INV_X4 _u0_U16617  ( .A(1'b0), .ZN(_u0_ch13_am0[8] ) );
INV_X4 _u0_U16615  ( .A(1'b0), .ZN(_u0_ch13_am0[7] ) );
INV_X4 _u0_U16613  ( .A(1'b0), .ZN(_u0_ch13_am0[6] ) );
INV_X4 _u0_U16611  ( .A(1'b0), .ZN(_u0_ch13_am0[5] ) );
INV_X4 _u0_U16609  ( .A(1'b0), .ZN(_u0_ch13_am0[4] ) );
INV_X4 _u0_U16607  ( .A(1'b1), .ZN(_u0_ch13_am0[3] ) );
INV_X4 _u0_U16605  ( .A(1'b1), .ZN(_u0_ch13_am0[2] ) );
INV_X4 _u0_U16603  ( .A(1'b1), .ZN(_u0_ch13_am0[1] ) );
INV_X4 _u0_U16601  ( .A(1'b1), .ZN(_u0_ch13_am0[0] ) );
INV_X4 _u0_U16599  ( .A(1'b0), .ZN(_u0_ch13_am1[31] ) );
INV_X4 _u0_U16597  ( .A(1'b0), .ZN(_u0_ch13_am1[30] ) );
INV_X4 _u0_U16595  ( .A(1'b0), .ZN(_u0_ch13_am1[29] ) );
INV_X4 _u0_U16593  ( .A(1'b0), .ZN(_u0_ch13_am1[28] ) );
INV_X4 _u0_U16591  ( .A(1'b0), .ZN(_u0_ch13_am1[27] ) );
INV_X4 _u0_U16589  ( .A(1'b0), .ZN(_u0_ch13_am1[26] ) );
INV_X4 _u0_U16587  ( .A(1'b0), .ZN(_u0_ch13_am1[25] ) );
INV_X4 _u0_U16585  ( .A(1'b0), .ZN(_u0_ch13_am1[24] ) );
INV_X4 _u0_U16583  ( .A(1'b0), .ZN(_u0_ch13_am1[23] ) );
INV_X4 _u0_U16581  ( .A(1'b0), .ZN(_u0_ch13_am1[22] ) );
INV_X4 _u0_U16579  ( .A(1'b0), .ZN(_u0_ch13_am1[21] ) );
INV_X4 _u0_U16577  ( .A(1'b0), .ZN(_u0_ch13_am1[20] ) );
INV_X4 _u0_U16575  ( .A(1'b0), .ZN(_u0_ch13_am1[19] ) );
INV_X4 _u0_U16573  ( .A(1'b0), .ZN(_u0_ch13_am1[18] ) );
INV_X4 _u0_U16571  ( .A(1'b0), .ZN(_u0_ch13_am1[17] ) );
INV_X4 _u0_U16569  ( .A(1'b0), .ZN(_u0_ch13_am1[16] ) );
INV_X4 _u0_U16567  ( .A(1'b0), .ZN(_u0_ch13_am1[15] ) );
INV_X4 _u0_U16565  ( .A(1'b0), .ZN(_u0_ch13_am1[14] ) );
INV_X4 _u0_U16563  ( .A(1'b0), .ZN(_u0_ch13_am1[13] ) );
INV_X4 _u0_U16561  ( .A(1'b0), .ZN(_u0_ch13_am1[12] ) );
INV_X4 _u0_U16559  ( .A(1'b0), .ZN(_u0_ch13_am1[11] ) );
INV_X4 _u0_U16557  ( .A(1'b0), .ZN(_u0_ch13_am1[10] ) );
INV_X4 _u0_U16555  ( .A(1'b0), .ZN(_u0_ch13_am1[9] ) );
INV_X4 _u0_U16553  ( .A(1'b0), .ZN(_u0_ch13_am1[8] ) );
INV_X4 _u0_U16551  ( .A(1'b0), .ZN(_u0_ch13_am1[7] ) );
INV_X4 _u0_U16549  ( .A(1'b0), .ZN(_u0_ch13_am1[6] ) );
INV_X4 _u0_U16547  ( .A(1'b0), .ZN(_u0_ch13_am1[5] ) );
INV_X4 _u0_U16545  ( .A(1'b0), .ZN(_u0_ch13_am1[4] ) );
INV_X4 _u0_U16543  ( .A(1'b1), .ZN(_u0_ch13_am1[3] ) );
INV_X4 _u0_U16541  ( .A(1'b1), .ZN(_u0_ch13_am1[2] ) );
INV_X4 _u0_U16539  ( .A(1'b1), .ZN(_u0_ch13_am1[1] ) );
INV_X4 _u0_U16537  ( .A(1'b1), .ZN(_u0_ch13_am1[0] ) );
INV_X4 _u0_U16535  ( .A(1'b1), .ZN(_u0_pointer14[31] ) );
INV_X4 _u0_U16533  ( .A(1'b1), .ZN(_u0_pointer14[30] ) );
INV_X4 _u0_U16531  ( .A(1'b1), .ZN(_u0_pointer14[29] ) );
INV_X4 _u0_U16529  ( .A(1'b1), .ZN(_u0_pointer14[28] ) );
INV_X4 _u0_U16527  ( .A(1'b1), .ZN(_u0_pointer14[27] ) );
INV_X4 _u0_U16525  ( .A(1'b1), .ZN(_u0_pointer14[26] ) );
INV_X4 _u0_U16523  ( .A(1'b1), .ZN(_u0_pointer14[25] ) );
INV_X4 _u0_U16521  ( .A(1'b1), .ZN(_u0_pointer14[24] ) );
INV_X4 _u0_U16519  ( .A(1'b1), .ZN(_u0_pointer14[23] ) );
INV_X4 _u0_U16517  ( .A(1'b1), .ZN(_u0_pointer14[22] ) );
INV_X4 _u0_U16515  ( .A(1'b1), .ZN(_u0_pointer14[21] ) );
INV_X4 _u0_U16513  ( .A(1'b1), .ZN(_u0_pointer14[20] ) );
INV_X4 _u0_U16511  ( .A(1'b1), .ZN(_u0_pointer14[19] ) );
INV_X4 _u0_U16509  ( .A(1'b1), .ZN(_u0_pointer14[18] ) );
INV_X4 _u0_U16507  ( .A(1'b1), .ZN(_u0_pointer14[17] ) );
INV_X4 _u0_U16505  ( .A(1'b1), .ZN(_u0_pointer14[16] ) );
INV_X4 _u0_U16503  ( .A(1'b1), .ZN(_u0_pointer14[15] ) );
INV_X4 _u0_U16501  ( .A(1'b1), .ZN(_u0_pointer14[14] ) );
INV_X4 _u0_U16499  ( .A(1'b1), .ZN(_u0_pointer14[13] ) );
INV_X4 _u0_U16497  ( .A(1'b1), .ZN(_u0_pointer14[12] ) );
INV_X4 _u0_U16495  ( .A(1'b1), .ZN(_u0_pointer14[11] ) );
INV_X4 _u0_U16493  ( .A(1'b1), .ZN(_u0_pointer14[10] ) );
INV_X4 _u0_U16491  ( .A(1'b1), .ZN(_u0_pointer14[9] ) );
INV_X4 _u0_U16489  ( .A(1'b1), .ZN(_u0_pointer14[8] ) );
INV_X4 _u0_U16487  ( .A(1'b1), .ZN(_u0_pointer14[7] ) );
INV_X4 _u0_U16485  ( .A(1'b1), .ZN(_u0_pointer14[6] ) );
INV_X4 _u0_U16483  ( .A(1'b1), .ZN(_u0_pointer14[5] ) );
INV_X4 _u0_U16481  ( .A(1'b1), .ZN(_u0_pointer14[4] ) );
INV_X4 _u0_U16479  ( .A(1'b1), .ZN(_u0_pointer14[3] ) );
INV_X4 _u0_U16477  ( .A(1'b1), .ZN(_u0_pointer14[2] ) );
INV_X4 _u0_U16475  ( .A(1'b1), .ZN(_u0_pointer14[1] ) );
INV_X4 _u0_U16473  ( .A(1'b1), .ZN(_u0_pointer14[0] ) );
INV_X4 _u0_U16471  ( .A(1'b1), .ZN(_u0_pointer14_s[31] ) );
INV_X4 _u0_U16469  ( .A(1'b1), .ZN(_u0_pointer14_s[30] ) );
INV_X4 _u0_U16467  ( .A(1'b1), .ZN(_u0_pointer14_s[29] ) );
INV_X4 _u0_U16465  ( .A(1'b1), .ZN(_u0_pointer14_s[28] ) );
INV_X4 _u0_U16463  ( .A(1'b1), .ZN(_u0_pointer14_s[27] ) );
INV_X4 _u0_U16461  ( .A(1'b1), .ZN(_u0_pointer14_s[26] ) );
INV_X4 _u0_U16459  ( .A(1'b1), .ZN(_u0_pointer14_s[25] ) );
INV_X4 _u0_U16457  ( .A(1'b1), .ZN(_u0_pointer14_s[24] ) );
INV_X4 _u0_U16455  ( .A(1'b1), .ZN(_u0_pointer14_s[23] ) );
INV_X4 _u0_U16453  ( .A(1'b1), .ZN(_u0_pointer14_s[22] ) );
INV_X4 _u0_U16451  ( .A(1'b1), .ZN(_u0_pointer14_s[21] ) );
INV_X4 _u0_U16449  ( .A(1'b1), .ZN(_u0_pointer14_s[20] ) );
INV_X4 _u0_U16447  ( .A(1'b1), .ZN(_u0_pointer14_s[19] ) );
INV_X4 _u0_U16445  ( .A(1'b1), .ZN(_u0_pointer14_s[18] ) );
INV_X4 _u0_U16443  ( .A(1'b1), .ZN(_u0_pointer14_s[17] ) );
INV_X4 _u0_U16441  ( .A(1'b1), .ZN(_u0_pointer14_s[16] ) );
INV_X4 _u0_U16439  ( .A(1'b1), .ZN(_u0_pointer14_s[15] ) );
INV_X4 _u0_U16437  ( .A(1'b1), .ZN(_u0_pointer14_s[14] ) );
INV_X4 _u0_U16435  ( .A(1'b1), .ZN(_u0_pointer14_s[13] ) );
INV_X4 _u0_U16433  ( .A(1'b1), .ZN(_u0_pointer14_s[12] ) );
INV_X4 _u0_U16431  ( .A(1'b1), .ZN(_u0_pointer14_s[11] ) );
INV_X4 _u0_U16429  ( .A(1'b1), .ZN(_u0_pointer14_s[10] ) );
INV_X4 _u0_U16427  ( .A(1'b1), .ZN(_u0_pointer14_s[9] ) );
INV_X4 _u0_U16425  ( .A(1'b1), .ZN(_u0_pointer14_s[8] ) );
INV_X4 _u0_U16423  ( .A(1'b1), .ZN(_u0_pointer14_s[7] ) );
INV_X4 _u0_U16421  ( .A(1'b1), .ZN(_u0_pointer14_s[6] ) );
INV_X4 _u0_U16419  ( .A(1'b1), .ZN(_u0_pointer14_s[5] ) );
INV_X4 _u0_U16417  ( .A(1'b1), .ZN(_u0_pointer14_s[4] ) );
INV_X4 _u0_U16415  ( .A(1'b1), .ZN(_u0_pointer14_s[3] ) );
INV_X4 _u0_U16413  ( .A(1'b1), .ZN(_u0_pointer14_s[2] ) );
INV_X4 _u0_U16411  ( .A(1'b1), .ZN(_u0_pointer14_s[1] ) );
INV_X4 _u0_U16409  ( .A(1'b1), .ZN(_u0_pointer14_s[0] ) );
INV_X4 _u0_U16407  ( .A(1'b1), .ZN(_u0_ch14_csr[31] ) );
INV_X4 _u0_U16405  ( .A(1'b1), .ZN(_u0_ch14_csr[30] ) );
INV_X4 _u0_U16403  ( .A(1'b1), .ZN(_u0_ch14_csr[29] ) );
INV_X4 _u0_U16401  ( .A(1'b1), .ZN(_u0_ch14_csr[28] ) );
INV_X4 _u0_U16399  ( .A(1'b1), .ZN(_u0_ch14_csr[27] ) );
INV_X4 _u0_U16397  ( .A(1'b1), .ZN(_u0_ch14_csr[26] ) );
INV_X4 _u0_U16395  ( .A(1'b1), .ZN(_u0_ch14_csr[25] ) );
INV_X4 _u0_U16393  ( .A(1'b1), .ZN(_u0_ch14_csr[24] ) );
INV_X4 _u0_U16391  ( .A(1'b1), .ZN(_u0_ch14_csr[23] ) );
INV_X4 _u0_U16389  ( .A(1'b1), .ZN(_u0_ch14_csr[22] ) );
INV_X4 _u0_U16387  ( .A(1'b1), .ZN(_u0_ch14_csr[21] ) );
INV_X4 _u0_U16385  ( .A(1'b1), .ZN(_u0_ch14_csr[20] ) );
INV_X4 _u0_U16383  ( .A(1'b1), .ZN(_u0_ch14_csr[19] ) );
INV_X4 _u0_U16381  ( .A(1'b1), .ZN(_u0_ch14_csr[18] ) );
INV_X4 _u0_U16379  ( .A(1'b1), .ZN(_u0_ch14_csr[17] ) );
INV_X4 _u0_U16377  ( .A(1'b1), .ZN(_u0_ch14_csr[16] ) );
INV_X4 _u0_U16375  ( .A(1'b1), .ZN(_u0_ch14_csr[15] ) );
INV_X4 _u0_U16373  ( .A(1'b1), .ZN(_u0_ch14_csr[14] ) );
INV_X4 _u0_U16371  ( .A(1'b1), .ZN(_u0_ch14_csr[13] ) );
INV_X4 _u0_U16369  ( .A(1'b1), .ZN(_u0_ch14_csr[12] ) );
INV_X4 _u0_U16367  ( .A(1'b1), .ZN(_u0_ch14_csr[11] ) );
INV_X4 _u0_U16365  ( .A(1'b1), .ZN(_u0_ch14_csr[10] ) );
INV_X4 _u0_U16363  ( .A(1'b1), .ZN(_u0_ch14_csr[9] ) );
INV_X4 _u0_U16361  ( .A(1'b1), .ZN(_u0_ch14_csr[8] ) );
INV_X4 _u0_U16359  ( .A(1'b1), .ZN(_u0_ch14_csr[7] ) );
INV_X4 _u0_U16357  ( .A(1'b1), .ZN(_u0_ch14_csr[6] ) );
INV_X4 _u0_U16355  ( .A(1'b1), .ZN(_u0_ch14_csr[5] ) );
INV_X4 _u0_U16353  ( .A(1'b1), .ZN(_u0_ch14_csr[4] ) );
INV_X4 _u0_U16351  ( .A(1'b1), .ZN(_u0_ch14_csr[3] ) );
INV_X4 _u0_U16349  ( .A(1'b1), .ZN(_u0_ch14_csr[2] ) );
INV_X4 _u0_U16347  ( .A(1'b1), .ZN(_u0_ch14_csr[1] ) );
INV_X4 _u0_U16345  ( .A(1'b1), .ZN(_u0_ch14_csr[0] ) );
INV_X4 _u0_U16343  ( .A(1'b1), .ZN(_u0_ch14_txsz[31] ) );
INV_X4 _u0_U16341  ( .A(1'b1), .ZN(_u0_ch14_txsz[30] ) );
INV_X4 _u0_U16339  ( .A(1'b1), .ZN(_u0_ch14_txsz[29] ) );
INV_X4 _u0_U16337  ( .A(1'b1), .ZN(_u0_ch14_txsz[28] ) );
INV_X4 _u0_U16335  ( .A(1'b1), .ZN(_u0_ch14_txsz[27] ) );
INV_X4 _u0_U16333  ( .A(1'b1), .ZN(_u0_ch14_txsz[26] ) );
INV_X4 _u0_U16331  ( .A(1'b1), .ZN(_u0_ch14_txsz[25] ) );
INV_X4 _u0_U16329  ( .A(1'b1), .ZN(_u0_ch14_txsz[24] ) );
INV_X4 _u0_U16327  ( .A(1'b1), .ZN(_u0_ch14_txsz[23] ) );
INV_X4 _u0_U16325  ( .A(1'b1), .ZN(_u0_ch14_txsz[22] ) );
INV_X4 _u0_U16323  ( .A(1'b1), .ZN(_u0_ch14_txsz[21] ) );
INV_X4 _u0_U16321  ( .A(1'b1), .ZN(_u0_ch14_txsz[20] ) );
INV_X4 _u0_U16319  ( .A(1'b1), .ZN(_u0_ch14_txsz[19] ) );
INV_X4 _u0_U16317  ( .A(1'b1), .ZN(_u0_ch14_txsz[18] ) );
INV_X4 _u0_U16315  ( .A(1'b1), .ZN(_u0_ch14_txsz[17] ) );
INV_X4 _u0_U16313  ( .A(1'b1), .ZN(_u0_ch14_txsz[16] ) );
INV_X4 _u0_U16311  ( .A(1'b1), .ZN(_u0_ch14_txsz[15] ) );
INV_X4 _u0_U16309  ( .A(1'b1), .ZN(_u0_ch14_txsz[14] ) );
INV_X4 _u0_U16307  ( .A(1'b1), .ZN(_u0_ch14_txsz[13] ) );
INV_X4 _u0_U16305  ( .A(1'b1), .ZN(_u0_ch14_txsz[12] ) );
INV_X4 _u0_U16303  ( .A(1'b1), .ZN(_u0_ch14_txsz[11] ) );
INV_X4 _u0_U16301  ( .A(1'b1), .ZN(_u0_ch14_txsz[10] ) );
INV_X4 _u0_U16299  ( .A(1'b1), .ZN(_u0_ch14_txsz[9] ) );
INV_X4 _u0_U16297  ( .A(1'b1), .ZN(_u0_ch14_txsz[8] ) );
INV_X4 _u0_U16295  ( .A(1'b1), .ZN(_u0_ch14_txsz[7] ) );
INV_X4 _u0_U16293  ( .A(1'b1), .ZN(_u0_ch14_txsz[6] ) );
INV_X4 _u0_U16291  ( .A(1'b1), .ZN(_u0_ch14_txsz[5] ) );
INV_X4 _u0_U16289  ( .A(1'b1), .ZN(_u0_ch14_txsz[4] ) );
INV_X4 _u0_U16287  ( .A(1'b1), .ZN(_u0_ch14_txsz[3] ) );
INV_X4 _u0_U16285  ( .A(1'b1), .ZN(_u0_ch14_txsz[2] ) );
INV_X4 _u0_U16283  ( .A(1'b1), .ZN(_u0_ch14_txsz[1] ) );
INV_X4 _u0_U16281  ( .A(1'b1), .ZN(_u0_ch14_txsz[0] ) );
INV_X4 _u0_U16279  ( .A(1'b1), .ZN(_u0_ch14_adr0[31] ) );
INV_X4 _u0_U16277  ( .A(1'b1), .ZN(_u0_ch14_adr0[30] ) );
INV_X4 _u0_U16275  ( .A(1'b1), .ZN(_u0_ch14_adr0[29] ) );
INV_X4 _u0_U16273  ( .A(1'b1), .ZN(_u0_ch14_adr0[28] ) );
INV_X4 _u0_U16271  ( .A(1'b1), .ZN(_u0_ch14_adr0[27] ) );
INV_X4 _u0_U16269  ( .A(1'b1), .ZN(_u0_ch14_adr0[26] ) );
INV_X4 _u0_U16267  ( .A(1'b1), .ZN(_u0_ch14_adr0[25] ) );
INV_X4 _u0_U16265  ( .A(1'b1), .ZN(_u0_ch14_adr0[24] ) );
INV_X4 _u0_U16263  ( .A(1'b1), .ZN(_u0_ch14_adr0[23] ) );
INV_X4 _u0_U16261  ( .A(1'b1), .ZN(_u0_ch14_adr0[22] ) );
INV_X4 _u0_U16259  ( .A(1'b1), .ZN(_u0_ch14_adr0[21] ) );
INV_X4 _u0_U16257  ( .A(1'b1), .ZN(_u0_ch14_adr0[20] ) );
INV_X4 _u0_U16255  ( .A(1'b1), .ZN(_u0_ch14_adr0[19] ) );
INV_X4 _u0_U16253  ( .A(1'b1), .ZN(_u0_ch14_adr0[18] ) );
INV_X4 _u0_U16251  ( .A(1'b1), .ZN(_u0_ch14_adr0[17] ) );
INV_X4 _u0_U16249  ( .A(1'b1), .ZN(_u0_ch14_adr0[16] ) );
INV_X4 _u0_U16247  ( .A(1'b1), .ZN(_u0_ch14_adr0[15] ) );
INV_X4 _u0_U16245  ( .A(1'b1), .ZN(_u0_ch14_adr0[14] ) );
INV_X4 _u0_U16243  ( .A(1'b1), .ZN(_u0_ch14_adr0[13] ) );
INV_X4 _u0_U16241  ( .A(1'b1), .ZN(_u0_ch14_adr0[12] ) );
INV_X4 _u0_U16239  ( .A(1'b1), .ZN(_u0_ch14_adr0[11] ) );
INV_X4 _u0_U16237  ( .A(1'b1), .ZN(_u0_ch14_adr0[10] ) );
INV_X4 _u0_U16235  ( .A(1'b1), .ZN(_u0_ch14_adr0[9] ) );
INV_X4 _u0_U16233  ( .A(1'b1), .ZN(_u0_ch14_adr0[8] ) );
INV_X4 _u0_U16231  ( .A(1'b1), .ZN(_u0_ch14_adr0[7] ) );
INV_X4 _u0_U16229  ( .A(1'b1), .ZN(_u0_ch14_adr0[6] ) );
INV_X4 _u0_U16227  ( .A(1'b1), .ZN(_u0_ch14_adr0[5] ) );
INV_X4 _u0_U16225  ( .A(1'b1), .ZN(_u0_ch14_adr0[4] ) );
INV_X4 _u0_U16223  ( .A(1'b1), .ZN(_u0_ch14_adr0[3] ) );
INV_X4 _u0_U16221  ( .A(1'b1), .ZN(_u0_ch14_adr0[2] ) );
INV_X4 _u0_U16219  ( .A(1'b1), .ZN(_u0_ch14_adr0[1] ) );
INV_X4 _u0_U16217  ( .A(1'b1), .ZN(_u0_ch14_adr0[0] ) );
INV_X4 _u0_U16215  ( .A(1'b1), .ZN(_u0_ch14_adr1[31] ) );
INV_X4 _u0_U16213  ( .A(1'b1), .ZN(_u0_ch14_adr1[30] ) );
INV_X4 _u0_U16211  ( .A(1'b1), .ZN(_u0_ch14_adr1[29] ) );
INV_X4 _u0_U16209  ( .A(1'b1), .ZN(_u0_ch14_adr1[28] ) );
INV_X4 _u0_U16207  ( .A(1'b1), .ZN(_u0_ch14_adr1[27] ) );
INV_X4 _u0_U16205  ( .A(1'b1), .ZN(_u0_ch14_adr1[26] ) );
INV_X4 _u0_U16203  ( .A(1'b1), .ZN(_u0_ch14_adr1[25] ) );
INV_X4 _u0_U16201  ( .A(1'b1), .ZN(_u0_ch14_adr1[24] ) );
INV_X4 _u0_U16199  ( .A(1'b1), .ZN(_u0_ch14_adr1[23] ) );
INV_X4 _u0_U16197  ( .A(1'b1), .ZN(_u0_ch14_adr1[22] ) );
INV_X4 _u0_U16195  ( .A(1'b1), .ZN(_u0_ch14_adr1[21] ) );
INV_X4 _u0_U16193  ( .A(1'b1), .ZN(_u0_ch14_adr1[20] ) );
INV_X4 _u0_U16191  ( .A(1'b1), .ZN(_u0_ch14_adr1[19] ) );
INV_X4 _u0_U16189  ( .A(1'b1), .ZN(_u0_ch14_adr1[18] ) );
INV_X4 _u0_U16187  ( .A(1'b1), .ZN(_u0_ch14_adr1[17] ) );
INV_X4 _u0_U16185  ( .A(1'b1), .ZN(_u0_ch14_adr1[16] ) );
INV_X4 _u0_U16183  ( .A(1'b1), .ZN(_u0_ch14_adr1[15] ) );
INV_X4 _u0_U16181  ( .A(1'b1), .ZN(_u0_ch14_adr1[14] ) );
INV_X4 _u0_U16179  ( .A(1'b1), .ZN(_u0_ch14_adr1[13] ) );
INV_X4 _u0_U16177  ( .A(1'b1), .ZN(_u0_ch14_adr1[12] ) );
INV_X4 _u0_U16175  ( .A(1'b1), .ZN(_u0_ch14_adr1[11] ) );
INV_X4 _u0_U16173  ( .A(1'b1), .ZN(_u0_ch14_adr1[10] ) );
INV_X4 _u0_U16171  ( .A(1'b1), .ZN(_u0_ch14_adr1[9] ) );
INV_X4 _u0_U16169  ( .A(1'b1), .ZN(_u0_ch14_adr1[8] ) );
INV_X4 _u0_U16167  ( .A(1'b1), .ZN(_u0_ch14_adr1[7] ) );
INV_X4 _u0_U16165  ( .A(1'b1), .ZN(_u0_ch14_adr1[6] ) );
INV_X4 _u0_U16163  ( .A(1'b1), .ZN(_u0_ch14_adr1[5] ) );
INV_X4 _u0_U16161  ( .A(1'b1), .ZN(_u0_ch14_adr1[4] ) );
INV_X4 _u0_U16159  ( .A(1'b1), .ZN(_u0_ch14_adr1[3] ) );
INV_X4 _u0_U16157  ( .A(1'b1), .ZN(_u0_ch14_adr1[2] ) );
INV_X4 _u0_U16155  ( .A(1'b1), .ZN(_u0_ch14_adr1[1] ) );
INV_X4 _u0_U16153  ( .A(1'b1), .ZN(_u0_ch14_adr1[0] ) );
INV_X4 _u0_U16151  ( .A(1'b0), .ZN(_u0_ch14_am0[31] ) );
INV_X4 _u0_U16149  ( .A(1'b0), .ZN(_u0_ch14_am0[30] ) );
INV_X4 _u0_U16147  ( .A(1'b0), .ZN(_u0_ch14_am0[29] ) );
INV_X4 _u0_U16145  ( .A(1'b0), .ZN(_u0_ch14_am0[28] ) );
INV_X4 _u0_U16143  ( .A(1'b0), .ZN(_u0_ch14_am0[27] ) );
INV_X4 _u0_U16141  ( .A(1'b0), .ZN(_u0_ch14_am0[26] ) );
INV_X4 _u0_U16139  ( .A(1'b0), .ZN(_u0_ch14_am0[25] ) );
INV_X4 _u0_U16137  ( .A(1'b0), .ZN(_u0_ch14_am0[24] ) );
INV_X4 _u0_U16135  ( .A(1'b0), .ZN(_u0_ch14_am0[23] ) );
INV_X4 _u0_U16133  ( .A(1'b0), .ZN(_u0_ch14_am0[22] ) );
INV_X4 _u0_U16131  ( .A(1'b0), .ZN(_u0_ch14_am0[21] ) );
INV_X4 _u0_U16129  ( .A(1'b0), .ZN(_u0_ch14_am0[20] ) );
INV_X4 _u0_U16127  ( .A(1'b0), .ZN(_u0_ch14_am0[19] ) );
INV_X4 _u0_U16125  ( .A(1'b0), .ZN(_u0_ch14_am0[18] ) );
INV_X4 _u0_U16123  ( .A(1'b0), .ZN(_u0_ch14_am0[17] ) );
INV_X4 _u0_U16121  ( .A(1'b0), .ZN(_u0_ch14_am0[16] ) );
INV_X4 _u0_U16119  ( .A(1'b0), .ZN(_u0_ch14_am0[15] ) );
INV_X4 _u0_U16117  ( .A(1'b0), .ZN(_u0_ch14_am0[14] ) );
INV_X4 _u0_U16115  ( .A(1'b0), .ZN(_u0_ch14_am0[13] ) );
INV_X4 _u0_U16113  ( .A(1'b0), .ZN(_u0_ch14_am0[12] ) );
INV_X4 _u0_U16111  ( .A(1'b0), .ZN(_u0_ch14_am0[11] ) );
INV_X4 _u0_U16109  ( .A(1'b0), .ZN(_u0_ch14_am0[10] ) );
INV_X4 _u0_U16107  ( .A(1'b0), .ZN(_u0_ch14_am0[9] ) );
INV_X4 _u0_U16105  ( .A(1'b0), .ZN(_u0_ch14_am0[8] ) );
INV_X4 _u0_U16103  ( .A(1'b0), .ZN(_u0_ch14_am0[7] ) );
INV_X4 _u0_U16101  ( .A(1'b0), .ZN(_u0_ch14_am0[6] ) );
INV_X4 _u0_U16099  ( .A(1'b0), .ZN(_u0_ch14_am0[5] ) );
INV_X4 _u0_U16097  ( .A(1'b0), .ZN(_u0_ch14_am0[4] ) );
INV_X4 _u0_U16095  ( .A(1'b1), .ZN(_u0_ch14_am0[3] ) );
INV_X4 _u0_U16093  ( .A(1'b1), .ZN(_u0_ch14_am0[2] ) );
INV_X4 _u0_U16091  ( .A(1'b1), .ZN(_u0_ch14_am0[1] ) );
INV_X4 _u0_U16089  ( .A(1'b1), .ZN(_u0_ch14_am0[0] ) );
INV_X4 _u0_U16087  ( .A(1'b0), .ZN(_u0_ch14_am1[31] ) );
INV_X4 _u0_U16085  ( .A(1'b0), .ZN(_u0_ch14_am1[30] ) );
INV_X4 _u0_U16083  ( .A(1'b0), .ZN(_u0_ch14_am1[29] ) );
INV_X4 _u0_U16081  ( .A(1'b0), .ZN(_u0_ch14_am1[28] ) );
INV_X4 _u0_U16079  ( .A(1'b0), .ZN(_u0_ch14_am1[27] ) );
INV_X4 _u0_U16077  ( .A(1'b0), .ZN(_u0_ch14_am1[26] ) );
INV_X4 _u0_U16075  ( .A(1'b0), .ZN(_u0_ch14_am1[25] ) );
INV_X4 _u0_U16073  ( .A(1'b0), .ZN(_u0_ch14_am1[24] ) );
INV_X4 _u0_U16071  ( .A(1'b0), .ZN(_u0_ch14_am1[23] ) );
INV_X4 _u0_U16069  ( .A(1'b0), .ZN(_u0_ch14_am1[22] ) );
INV_X4 _u0_U16067  ( .A(1'b0), .ZN(_u0_ch14_am1[21] ) );
INV_X4 _u0_U16065  ( .A(1'b0), .ZN(_u0_ch14_am1[20] ) );
INV_X4 _u0_U16063  ( .A(1'b0), .ZN(_u0_ch14_am1[19] ) );
INV_X4 _u0_U16061  ( .A(1'b0), .ZN(_u0_ch14_am1[18] ) );
INV_X4 _u0_U16059  ( .A(1'b0), .ZN(_u0_ch14_am1[17] ) );
INV_X4 _u0_U16057  ( .A(1'b0), .ZN(_u0_ch14_am1[16] ) );
INV_X4 _u0_U16055  ( .A(1'b0), .ZN(_u0_ch14_am1[15] ) );
INV_X4 _u0_U16053  ( .A(1'b0), .ZN(_u0_ch14_am1[14] ) );
INV_X4 _u0_U16051  ( .A(1'b0), .ZN(_u0_ch14_am1[13] ) );
INV_X4 _u0_U16049  ( .A(1'b0), .ZN(_u0_ch14_am1[12] ) );
INV_X4 _u0_U16047  ( .A(1'b0), .ZN(_u0_ch14_am1[11] ) );
INV_X4 _u0_U16045  ( .A(1'b0), .ZN(_u0_ch14_am1[10] ) );
INV_X4 _u0_U16043  ( .A(1'b0), .ZN(_u0_ch14_am1[9] ) );
INV_X4 _u0_U16041  ( .A(1'b0), .ZN(_u0_ch14_am1[8] ) );
INV_X4 _u0_U16039  ( .A(1'b0), .ZN(_u0_ch14_am1[7] ) );
INV_X4 _u0_U16037  ( .A(1'b0), .ZN(_u0_ch14_am1[6] ) );
INV_X4 _u0_U16035  ( .A(1'b0), .ZN(_u0_ch14_am1[5] ) );
INV_X4 _u0_U16033  ( .A(1'b0), .ZN(_u0_ch14_am1[4] ) );
INV_X4 _u0_U16031  ( .A(1'b1), .ZN(_u0_ch14_am1[3] ) );
INV_X4 _u0_U16029  ( .A(1'b1), .ZN(_u0_ch14_am1[2] ) );
INV_X4 _u0_U16027  ( .A(1'b1), .ZN(_u0_ch14_am1[1] ) );
INV_X4 _u0_U16025  ( .A(1'b1), .ZN(_u0_ch14_am1[0] ) );
INV_X4 _u0_U16023  ( .A(1'b1), .ZN(_u0_pointer15[31] ) );
INV_X4 _u0_U16021  ( .A(1'b1), .ZN(_u0_pointer15[30] ) );
INV_X4 _u0_U16019  ( .A(1'b1), .ZN(_u0_pointer15[29] ) );
INV_X4 _u0_U16017  ( .A(1'b1), .ZN(_u0_pointer15[28] ) );
INV_X4 _u0_U16015  ( .A(1'b1), .ZN(_u0_pointer15[27] ) );
INV_X4 _u0_U16013  ( .A(1'b1), .ZN(_u0_pointer15[26] ) );
INV_X4 _u0_U16011  ( .A(1'b1), .ZN(_u0_pointer15[25] ) );
INV_X4 _u0_U16009  ( .A(1'b1), .ZN(_u0_pointer15[24] ) );
INV_X4 _u0_U16007  ( .A(1'b1), .ZN(_u0_pointer15[23] ) );
INV_X4 _u0_U16005  ( .A(1'b1), .ZN(_u0_pointer15[22] ) );
INV_X4 _u0_U16003  ( .A(1'b1), .ZN(_u0_pointer15[21] ) );
INV_X4 _u0_U16001  ( .A(1'b1), .ZN(_u0_pointer15[20] ) );
INV_X4 _u0_U15999  ( .A(1'b1), .ZN(_u0_pointer15[19] ) );
INV_X4 _u0_U15997  ( .A(1'b1), .ZN(_u0_pointer15[18] ) );
INV_X4 _u0_U15995  ( .A(1'b1), .ZN(_u0_pointer15[17] ) );
INV_X4 _u0_U15993  ( .A(1'b1), .ZN(_u0_pointer15[16] ) );
INV_X4 _u0_U15991  ( .A(1'b1), .ZN(_u0_pointer15[15] ) );
INV_X4 _u0_U15989  ( .A(1'b1), .ZN(_u0_pointer15[14] ) );
INV_X4 _u0_U15987  ( .A(1'b1), .ZN(_u0_pointer15[13] ) );
INV_X4 _u0_U15985  ( .A(1'b1), .ZN(_u0_pointer15[12] ) );
INV_X4 _u0_U15983  ( .A(1'b1), .ZN(_u0_pointer15[11] ) );
INV_X4 _u0_U15981  ( .A(1'b1), .ZN(_u0_pointer15[10] ) );
INV_X4 _u0_U15979  ( .A(1'b1), .ZN(_u0_pointer15[9] ) );
INV_X4 _u0_U15977  ( .A(1'b1), .ZN(_u0_pointer15[8] ) );
INV_X4 _u0_U15975  ( .A(1'b1), .ZN(_u0_pointer15[7] ) );
INV_X4 _u0_U15973  ( .A(1'b1), .ZN(_u0_pointer15[6] ) );
INV_X4 _u0_U15971  ( .A(1'b1), .ZN(_u0_pointer15[5] ) );
INV_X4 _u0_U15969  ( .A(1'b1), .ZN(_u0_pointer15[4] ) );
INV_X4 _u0_U15967  ( .A(1'b1), .ZN(_u0_pointer15[3] ) );
INV_X4 _u0_U15965  ( .A(1'b1), .ZN(_u0_pointer15[2] ) );
INV_X4 _u0_U15963  ( .A(1'b1), .ZN(_u0_pointer15[1] ) );
INV_X4 _u0_U15961  ( .A(1'b1), .ZN(_u0_pointer15[0] ) );
INV_X4 _u0_U15959  ( .A(1'b1), .ZN(_u0_pointer15_s[31] ) );
INV_X4 _u0_U15957  ( .A(1'b1), .ZN(_u0_pointer15_s[30] ) );
INV_X4 _u0_U15955  ( .A(1'b1), .ZN(_u0_pointer15_s[29] ) );
INV_X4 _u0_U15953  ( .A(1'b1), .ZN(_u0_pointer15_s[28] ) );
INV_X4 _u0_U15951  ( .A(1'b1), .ZN(_u0_pointer15_s[27] ) );
INV_X4 _u0_U15949  ( .A(1'b1), .ZN(_u0_pointer15_s[26] ) );
INV_X4 _u0_U15947  ( .A(1'b1), .ZN(_u0_pointer15_s[25] ) );
INV_X4 _u0_U15945  ( .A(1'b1), .ZN(_u0_pointer15_s[24] ) );
INV_X4 _u0_U15943  ( .A(1'b1), .ZN(_u0_pointer15_s[23] ) );
INV_X4 _u0_U15941  ( .A(1'b1), .ZN(_u0_pointer15_s[22] ) );
INV_X4 _u0_U15939  ( .A(1'b1), .ZN(_u0_pointer15_s[21] ) );
INV_X4 _u0_U15937  ( .A(1'b1), .ZN(_u0_pointer15_s[20] ) );
INV_X4 _u0_U15935  ( .A(1'b1), .ZN(_u0_pointer15_s[19] ) );
INV_X4 _u0_U15933  ( .A(1'b1), .ZN(_u0_pointer15_s[18] ) );
INV_X4 _u0_U15931  ( .A(1'b1), .ZN(_u0_pointer15_s[17] ) );
INV_X4 _u0_U15929  ( .A(1'b1), .ZN(_u0_pointer15_s[16] ) );
INV_X4 _u0_U15927  ( .A(1'b1), .ZN(_u0_pointer15_s[15] ) );
INV_X4 _u0_U15925  ( .A(1'b1), .ZN(_u0_pointer15_s[14] ) );
INV_X4 _u0_U15923  ( .A(1'b1), .ZN(_u0_pointer15_s[13] ) );
INV_X4 _u0_U15921  ( .A(1'b1), .ZN(_u0_pointer15_s[12] ) );
INV_X4 _u0_U15919  ( .A(1'b1), .ZN(_u0_pointer15_s[11] ) );
INV_X4 _u0_U15917  ( .A(1'b1), .ZN(_u0_pointer15_s[10] ) );
INV_X4 _u0_U15915  ( .A(1'b1), .ZN(_u0_pointer15_s[9] ) );
INV_X4 _u0_U15913  ( .A(1'b1), .ZN(_u0_pointer15_s[8] ) );
INV_X4 _u0_U15911  ( .A(1'b1), .ZN(_u0_pointer15_s[7] ) );
INV_X4 _u0_U15909  ( .A(1'b1), .ZN(_u0_pointer15_s[6] ) );
INV_X4 _u0_U15907  ( .A(1'b1), .ZN(_u0_pointer15_s[5] ) );
INV_X4 _u0_U15905  ( .A(1'b1), .ZN(_u0_pointer15_s[4] ) );
INV_X4 _u0_U15903  ( .A(1'b1), .ZN(_u0_pointer15_s[3] ) );
INV_X4 _u0_U15901  ( .A(1'b1), .ZN(_u0_pointer15_s[2] ) );
INV_X4 _u0_U15899  ( .A(1'b1), .ZN(_u0_pointer15_s[1] ) );
INV_X4 _u0_U15897  ( .A(1'b1), .ZN(_u0_pointer15_s[0] ) );
INV_X4 _u0_U15895  ( .A(1'b1), .ZN(_u0_ch15_csr[31] ) );
INV_X4 _u0_U15893  ( .A(1'b1), .ZN(_u0_ch15_csr[30] ) );
INV_X4 _u0_U15891  ( .A(1'b1), .ZN(_u0_ch15_csr[29] ) );
INV_X4 _u0_U15889  ( .A(1'b1), .ZN(_u0_ch15_csr[28] ) );
INV_X4 _u0_U15887  ( .A(1'b1), .ZN(_u0_ch15_csr[27] ) );
INV_X4 _u0_U15885  ( .A(1'b1), .ZN(_u0_ch15_csr[26] ) );
INV_X4 _u0_U15883  ( .A(1'b1), .ZN(_u0_ch15_csr[25] ) );
INV_X4 _u0_U15881  ( .A(1'b1), .ZN(_u0_ch15_csr[24] ) );
INV_X4 _u0_U15879  ( .A(1'b1), .ZN(_u0_ch15_csr[23] ) );
INV_X4 _u0_U15877  ( .A(1'b1), .ZN(_u0_ch15_csr[22] ) );
INV_X4 _u0_U15875  ( .A(1'b1), .ZN(_u0_ch15_csr[21] ) );
INV_X4 _u0_U15873  ( .A(1'b1), .ZN(_u0_ch15_csr[20] ) );
INV_X4 _u0_U15871  ( .A(1'b1), .ZN(_u0_ch15_csr[19] ) );
INV_X4 _u0_U15869  ( .A(1'b1), .ZN(_u0_ch15_csr[18] ) );
INV_X4 _u0_U15867  ( .A(1'b1), .ZN(_u0_ch15_csr[17] ) );
INV_X4 _u0_U15865  ( .A(1'b1), .ZN(_u0_ch15_csr[16] ) );
INV_X4 _u0_U15863  ( .A(1'b1), .ZN(_u0_ch15_csr[15] ) );
INV_X4 _u0_U15861  ( .A(1'b1), .ZN(_u0_ch15_csr[14] ) );
INV_X4 _u0_U15859  ( .A(1'b1), .ZN(_u0_ch15_csr[13] ) );
INV_X4 _u0_U15857  ( .A(1'b1), .ZN(_u0_ch15_csr[12] ) );
INV_X4 _u0_U15855  ( .A(1'b1), .ZN(_u0_ch15_csr[11] ) );
INV_X4 _u0_U15853  ( .A(1'b1), .ZN(_u0_ch15_csr[10] ) );
INV_X4 _u0_U15851  ( .A(1'b1), .ZN(_u0_ch15_csr[9] ) );
INV_X4 _u0_U15849  ( .A(1'b1), .ZN(_u0_ch15_csr[8] ) );
INV_X4 _u0_U15847  ( .A(1'b1), .ZN(_u0_ch15_csr[7] ) );
INV_X4 _u0_U15845  ( .A(1'b1), .ZN(_u0_ch15_csr[6] ) );
INV_X4 _u0_U15843  ( .A(1'b1), .ZN(_u0_ch15_csr[5] ) );
INV_X4 _u0_U15841  ( .A(1'b1), .ZN(_u0_ch15_csr[4] ) );
INV_X4 _u0_U15839  ( .A(1'b1), .ZN(_u0_ch15_csr[3] ) );
INV_X4 _u0_U15837  ( .A(1'b1), .ZN(_u0_ch15_csr[2] ) );
INV_X4 _u0_U15835  ( .A(1'b1), .ZN(_u0_ch15_csr[1] ) );
INV_X4 _u0_U15833  ( .A(1'b1), .ZN(_u0_ch15_csr[0] ) );
INV_X4 _u0_U15831  ( .A(1'b1), .ZN(_u0_ch15_txsz[31] ) );
INV_X4 _u0_U15829  ( .A(1'b1), .ZN(_u0_ch15_txsz[30] ) );
INV_X4 _u0_U15827  ( .A(1'b1), .ZN(_u0_ch15_txsz[29] ) );
INV_X4 _u0_U15825  ( .A(1'b1), .ZN(_u0_ch15_txsz[28] ) );
INV_X4 _u0_U15823  ( .A(1'b1), .ZN(_u0_ch15_txsz[27] ) );
INV_X4 _u0_U15821  ( .A(1'b1), .ZN(_u0_ch15_txsz[26] ) );
INV_X4 _u0_U15819  ( .A(1'b1), .ZN(_u0_ch15_txsz[25] ) );
INV_X4 _u0_U15817  ( .A(1'b1), .ZN(_u0_ch15_txsz[24] ) );
INV_X4 _u0_U15815  ( .A(1'b1), .ZN(_u0_ch15_txsz[23] ) );
INV_X4 _u0_U15813  ( .A(1'b1), .ZN(_u0_ch15_txsz[22] ) );
INV_X4 _u0_U15811  ( .A(1'b1), .ZN(_u0_ch15_txsz[21] ) );
INV_X4 _u0_U15809  ( .A(1'b1), .ZN(_u0_ch15_txsz[20] ) );
INV_X4 _u0_U15807  ( .A(1'b1), .ZN(_u0_ch15_txsz[19] ) );
INV_X4 _u0_U15805  ( .A(1'b1), .ZN(_u0_ch15_txsz[18] ) );
INV_X4 _u0_U15803  ( .A(1'b1), .ZN(_u0_ch15_txsz[17] ) );
INV_X4 _u0_U15801  ( .A(1'b1), .ZN(_u0_ch15_txsz[16] ) );
INV_X4 _u0_U15799  ( .A(1'b1), .ZN(_u0_ch15_txsz[15] ) );
INV_X4 _u0_U15797  ( .A(1'b1), .ZN(_u0_ch15_txsz[14] ) );
INV_X4 _u0_U15795  ( .A(1'b1), .ZN(_u0_ch15_txsz[13] ) );
INV_X4 _u0_U15793  ( .A(1'b1), .ZN(_u0_ch15_txsz[12] ) );
INV_X4 _u0_U15791  ( .A(1'b1), .ZN(_u0_ch15_txsz[11] ) );
INV_X4 _u0_U15789  ( .A(1'b1), .ZN(_u0_ch15_txsz[10] ) );
INV_X4 _u0_U15787  ( .A(1'b1), .ZN(_u0_ch15_txsz[9] ) );
INV_X4 _u0_U15785  ( .A(1'b1), .ZN(_u0_ch15_txsz[8] ) );
INV_X4 _u0_U15783  ( .A(1'b1), .ZN(_u0_ch15_txsz[7] ) );
INV_X4 _u0_U15781  ( .A(1'b1), .ZN(_u0_ch15_txsz[6] ) );
INV_X4 _u0_U15779  ( .A(1'b1), .ZN(_u0_ch15_txsz[5] ) );
INV_X4 _u0_U15777  ( .A(1'b1), .ZN(_u0_ch15_txsz[4] ) );
INV_X4 _u0_U15775  ( .A(1'b1), .ZN(_u0_ch15_txsz[3] ) );
INV_X4 _u0_U15773  ( .A(1'b1), .ZN(_u0_ch15_txsz[2] ) );
INV_X4 _u0_U15771  ( .A(1'b1), .ZN(_u0_ch15_txsz[1] ) );
INV_X4 _u0_U15769  ( .A(1'b1), .ZN(_u0_ch15_txsz[0] ) );
INV_X4 _u0_U15767  ( .A(1'b1), .ZN(_u0_ch15_adr0[31] ) );
INV_X4 _u0_U15765  ( .A(1'b1), .ZN(_u0_ch15_adr0[30] ) );
INV_X4 _u0_U15763  ( .A(1'b1), .ZN(_u0_ch15_adr0[29] ) );
INV_X4 _u0_U15761  ( .A(1'b1), .ZN(_u0_ch15_adr0[28] ) );
INV_X4 _u0_U15759  ( .A(1'b1), .ZN(_u0_ch15_adr0[27] ) );
INV_X4 _u0_U15757  ( .A(1'b1), .ZN(_u0_ch15_adr0[26] ) );
INV_X4 _u0_U15755  ( .A(1'b1), .ZN(_u0_ch15_adr0[25] ) );
INV_X4 _u0_U15753  ( .A(1'b1), .ZN(_u0_ch15_adr0[24] ) );
INV_X4 _u0_U15751  ( .A(1'b1), .ZN(_u0_ch15_adr0[23] ) );
INV_X4 _u0_U15749  ( .A(1'b1), .ZN(_u0_ch15_adr0[22] ) );
INV_X4 _u0_U15747  ( .A(1'b1), .ZN(_u0_ch15_adr0[21] ) );
INV_X4 _u0_U15745  ( .A(1'b1), .ZN(_u0_ch15_adr0[20] ) );
INV_X4 _u0_U15743  ( .A(1'b1), .ZN(_u0_ch15_adr0[19] ) );
INV_X4 _u0_U15741  ( .A(1'b1), .ZN(_u0_ch15_adr0[18] ) );
INV_X4 _u0_U15739  ( .A(1'b1), .ZN(_u0_ch15_adr0[17] ) );
INV_X4 _u0_U15737  ( .A(1'b1), .ZN(_u0_ch15_adr0[16] ) );
INV_X4 _u0_U15735  ( .A(1'b1), .ZN(_u0_ch15_adr0[15] ) );
INV_X4 _u0_U15733  ( .A(1'b1), .ZN(_u0_ch15_adr0[14] ) );
INV_X4 _u0_U15731  ( .A(1'b1), .ZN(_u0_ch15_adr0[13] ) );
INV_X4 _u0_U15729  ( .A(1'b1), .ZN(_u0_ch15_adr0[12] ) );
INV_X4 _u0_U15727  ( .A(1'b1), .ZN(_u0_ch15_adr0[11] ) );
INV_X4 _u0_U15725  ( .A(1'b1), .ZN(_u0_ch15_adr0[10] ) );
INV_X4 _u0_U15723  ( .A(1'b1), .ZN(_u0_ch15_adr0[9] ) );
INV_X4 _u0_U15721  ( .A(1'b1), .ZN(_u0_ch15_adr0[8] ) );
INV_X4 _u0_U15719  ( .A(1'b1), .ZN(_u0_ch15_adr0[7] ) );
INV_X4 _u0_U15717  ( .A(1'b1), .ZN(_u0_ch15_adr0[6] ) );
INV_X4 _u0_U15715  ( .A(1'b1), .ZN(_u0_ch15_adr0[5] ) );
INV_X4 _u0_U15713  ( .A(1'b1), .ZN(_u0_ch15_adr0[4] ) );
INV_X4 _u0_U15711  ( .A(1'b1), .ZN(_u0_ch15_adr0[3] ) );
INV_X4 _u0_U15709  ( .A(1'b1), .ZN(_u0_ch15_adr0[2] ) );
INV_X4 _u0_U15707  ( .A(1'b1), .ZN(_u0_ch15_adr0[1] ) );
INV_X4 _u0_U15705  ( .A(1'b1), .ZN(_u0_ch15_adr0[0] ) );
INV_X4 _u0_U15703  ( .A(1'b1), .ZN(_u0_ch15_adr1[31] ) );
INV_X4 _u0_U15701  ( .A(1'b1), .ZN(_u0_ch15_adr1[30] ) );
INV_X4 _u0_U15699  ( .A(1'b1), .ZN(_u0_ch15_adr1[29] ) );
INV_X4 _u0_U15697  ( .A(1'b1), .ZN(_u0_ch15_adr1[28] ) );
INV_X4 _u0_U15695  ( .A(1'b1), .ZN(_u0_ch15_adr1[27] ) );
INV_X4 _u0_U15693  ( .A(1'b1), .ZN(_u0_ch15_adr1[26] ) );
INV_X4 _u0_U15691  ( .A(1'b1), .ZN(_u0_ch15_adr1[25] ) );
INV_X4 _u0_U15689  ( .A(1'b1), .ZN(_u0_ch15_adr1[24] ) );
INV_X4 _u0_U15687  ( .A(1'b1), .ZN(_u0_ch15_adr1[23] ) );
INV_X4 _u0_U15685  ( .A(1'b1), .ZN(_u0_ch15_adr1[22] ) );
INV_X4 _u0_U15683  ( .A(1'b1), .ZN(_u0_ch15_adr1[21] ) );
INV_X4 _u0_U15681  ( .A(1'b1), .ZN(_u0_ch15_adr1[20] ) );
INV_X4 _u0_U15679  ( .A(1'b1), .ZN(_u0_ch15_adr1[19] ) );
INV_X4 _u0_U15677  ( .A(1'b1), .ZN(_u0_ch15_adr1[18] ) );
INV_X4 _u0_U15675  ( .A(1'b1), .ZN(_u0_ch15_adr1[17] ) );
INV_X4 _u0_U15673  ( .A(1'b1), .ZN(_u0_ch15_adr1[16] ) );
INV_X4 _u0_U15671  ( .A(1'b1), .ZN(_u0_ch15_adr1[15] ) );
INV_X4 _u0_U15669  ( .A(1'b1), .ZN(_u0_ch15_adr1[14] ) );
INV_X4 _u0_U15667  ( .A(1'b1), .ZN(_u0_ch15_adr1[13] ) );
INV_X4 _u0_U15665  ( .A(1'b1), .ZN(_u0_ch15_adr1[12] ) );
INV_X4 _u0_U15663  ( .A(1'b1), .ZN(_u0_ch15_adr1[11] ) );
INV_X4 _u0_U15661  ( .A(1'b1), .ZN(_u0_ch15_adr1[10] ) );
INV_X4 _u0_U15659  ( .A(1'b1), .ZN(_u0_ch15_adr1[9] ) );
INV_X4 _u0_U15657  ( .A(1'b1), .ZN(_u0_ch15_adr1[8] ) );
INV_X4 _u0_U15655  ( .A(1'b1), .ZN(_u0_ch15_adr1[7] ) );
INV_X4 _u0_U15653  ( .A(1'b1), .ZN(_u0_ch15_adr1[6] ) );
INV_X4 _u0_U15651  ( .A(1'b1), .ZN(_u0_ch15_adr1[5] ) );
INV_X4 _u0_U15649  ( .A(1'b1), .ZN(_u0_ch15_adr1[4] ) );
INV_X4 _u0_U15647  ( .A(1'b1), .ZN(_u0_ch15_adr1[3] ) );
INV_X4 _u0_U15645  ( .A(1'b1), .ZN(_u0_ch15_adr1[2] ) );
INV_X4 _u0_U15643  ( .A(1'b1), .ZN(_u0_ch15_adr1[1] ) );
INV_X4 _u0_U15641  ( .A(1'b1), .ZN(_u0_ch15_adr1[0] ) );
INV_X4 _u0_U15639  ( .A(1'b0), .ZN(_u0_ch15_am0[31] ) );
INV_X4 _u0_U15637  ( .A(1'b0), .ZN(_u0_ch15_am0[30] ) );
INV_X4 _u0_U15635  ( .A(1'b0), .ZN(_u0_ch15_am0[29] ) );
INV_X4 _u0_U15633  ( .A(1'b0), .ZN(_u0_ch15_am0[28] ) );
INV_X4 _u0_U15631  ( .A(1'b0), .ZN(_u0_ch15_am0[27] ) );
INV_X4 _u0_U15629  ( .A(1'b0), .ZN(_u0_ch15_am0[26] ) );
INV_X4 _u0_U15627  ( .A(1'b0), .ZN(_u0_ch15_am0[25] ) );
INV_X4 _u0_U15625  ( .A(1'b0), .ZN(_u0_ch15_am0[24] ) );
INV_X4 _u0_U15623  ( .A(1'b0), .ZN(_u0_ch15_am0[23] ) );
INV_X4 _u0_U15621  ( .A(1'b0), .ZN(_u0_ch15_am0[22] ) );
INV_X4 _u0_U15619  ( .A(1'b0), .ZN(_u0_ch15_am0[21] ) );
INV_X4 _u0_U15617  ( .A(1'b0), .ZN(_u0_ch15_am0[20] ) );
INV_X4 _u0_U15615  ( .A(1'b0), .ZN(_u0_ch15_am0[19] ) );
INV_X4 _u0_U15613  ( .A(1'b0), .ZN(_u0_ch15_am0[18] ) );
INV_X4 _u0_U15611  ( .A(1'b0), .ZN(_u0_ch15_am0[17] ) );
INV_X4 _u0_U15609  ( .A(1'b0), .ZN(_u0_ch15_am0[16] ) );
INV_X4 _u0_U15607  ( .A(1'b0), .ZN(_u0_ch15_am0[15] ) );
INV_X4 _u0_U15605  ( .A(1'b0), .ZN(_u0_ch15_am0[14] ) );
INV_X4 _u0_U15603  ( .A(1'b0), .ZN(_u0_ch15_am0[13] ) );
INV_X4 _u0_U15601  ( .A(1'b0), .ZN(_u0_ch15_am0[12] ) );
INV_X4 _u0_U15599  ( .A(1'b0), .ZN(_u0_ch15_am0[11] ) );
INV_X4 _u0_U15597  ( .A(1'b0), .ZN(_u0_ch15_am0[10] ) );
INV_X4 _u0_U15595  ( .A(1'b0), .ZN(_u0_ch15_am0[9] ) );
INV_X4 _u0_U15593  ( .A(1'b0), .ZN(_u0_ch15_am0[8] ) );
INV_X4 _u0_U15591  ( .A(1'b0), .ZN(_u0_ch15_am0[7] ) );
INV_X4 _u0_U15589  ( .A(1'b0), .ZN(_u0_ch15_am0[6] ) );
INV_X4 _u0_U15587  ( .A(1'b0), .ZN(_u0_ch15_am0[5] ) );
INV_X4 _u0_U15585  ( .A(1'b0), .ZN(_u0_ch15_am0[4] ) );
INV_X4 _u0_U15583  ( .A(1'b1), .ZN(_u0_ch15_am0[3] ) );
INV_X4 _u0_U15581  ( .A(1'b1), .ZN(_u0_ch15_am0[2] ) );
INV_X4 _u0_U15579  ( .A(1'b1), .ZN(_u0_ch15_am0[1] ) );
INV_X4 _u0_U15577  ( .A(1'b1), .ZN(_u0_ch15_am0[0] ) );
INV_X4 _u0_U15575  ( .A(1'b0), .ZN(_u0_ch15_am1[31] ) );
INV_X4 _u0_U15573  ( .A(1'b0), .ZN(_u0_ch15_am1[30] ) );
INV_X4 _u0_U15571  ( .A(1'b0), .ZN(_u0_ch15_am1[29] ) );
INV_X4 _u0_U15569  ( .A(1'b0), .ZN(_u0_ch15_am1[28] ) );
INV_X4 _u0_U15567  ( .A(1'b0), .ZN(_u0_ch15_am1[27] ) );
INV_X4 _u0_U15565  ( .A(1'b0), .ZN(_u0_ch15_am1[26] ) );
INV_X4 _u0_U15563  ( .A(1'b0), .ZN(_u0_ch15_am1[25] ) );
INV_X4 _u0_U15561  ( .A(1'b0), .ZN(_u0_ch15_am1[24] ) );
INV_X4 _u0_U15559  ( .A(1'b0), .ZN(_u0_ch15_am1[23] ) );
INV_X4 _u0_U15557  ( .A(1'b0), .ZN(_u0_ch15_am1[22] ) );
INV_X4 _u0_U15555  ( .A(1'b0), .ZN(_u0_ch15_am1[21] ) );
INV_X4 _u0_U15553  ( .A(1'b0), .ZN(_u0_ch15_am1[20] ) );
INV_X4 _u0_U15551  ( .A(1'b0), .ZN(_u0_ch15_am1[19] ) );
INV_X4 _u0_U15549  ( .A(1'b0), .ZN(_u0_ch15_am1[18] ) );
INV_X4 _u0_U15547  ( .A(1'b0), .ZN(_u0_ch15_am1[17] ) );
INV_X4 _u0_U15545  ( .A(1'b0), .ZN(_u0_ch15_am1[16] ) );
INV_X4 _u0_U15543  ( .A(1'b0), .ZN(_u0_ch15_am1[15] ) );
INV_X4 _u0_U15541  ( .A(1'b0), .ZN(_u0_ch15_am1[14] ) );
INV_X4 _u0_U15539  ( .A(1'b0), .ZN(_u0_ch15_am1[13] ) );
INV_X4 _u0_U15537  ( .A(1'b0), .ZN(_u0_ch15_am1[12] ) );
INV_X4 _u0_U15535  ( .A(1'b0), .ZN(_u0_ch15_am1[11] ) );
INV_X4 _u0_U15533  ( .A(1'b0), .ZN(_u0_ch15_am1[10] ) );
INV_X4 _u0_U15531  ( .A(1'b0), .ZN(_u0_ch15_am1[9] ) );
INV_X4 _u0_U15529  ( .A(1'b0), .ZN(_u0_ch15_am1[8] ) );
INV_X4 _u0_U15527  ( .A(1'b0), .ZN(_u0_ch15_am1[7] ) );
INV_X4 _u0_U15525  ( .A(1'b0), .ZN(_u0_ch15_am1[6] ) );
INV_X4 _u0_U15523  ( .A(1'b0), .ZN(_u0_ch15_am1[5] ) );
INV_X4 _u0_U15521  ( .A(1'b0), .ZN(_u0_ch15_am1[4] ) );
INV_X4 _u0_U15519  ( .A(1'b1), .ZN(_u0_ch15_am1[3] ) );
INV_X4 _u0_U15517  ( .A(1'b1), .ZN(_u0_ch15_am1[2] ) );
INV_X4 _u0_U15515  ( .A(1'b1), .ZN(_u0_ch15_am1[1] ) );
INV_X4 _u0_U15513  ( .A(1'b1), .ZN(_u0_ch15_am1[0] ) );
INV_X4 _u0_U15511  ( .A(1'b1), .ZN(_u0_pointer16[31] ) );
INV_X4 _u0_U15509  ( .A(1'b1), .ZN(_u0_pointer16[30] ) );
INV_X4 _u0_U15507  ( .A(1'b1), .ZN(_u0_pointer16[29] ) );
INV_X4 _u0_U15505  ( .A(1'b1), .ZN(_u0_pointer16[28] ) );
INV_X4 _u0_U15503  ( .A(1'b1), .ZN(_u0_pointer16[27] ) );
INV_X4 _u0_U15501  ( .A(1'b1), .ZN(_u0_pointer16[26] ) );
INV_X4 _u0_U15499  ( .A(1'b1), .ZN(_u0_pointer16[25] ) );
INV_X4 _u0_U15497  ( .A(1'b1), .ZN(_u0_pointer16[24] ) );
INV_X4 _u0_U15495  ( .A(1'b1), .ZN(_u0_pointer16[23] ) );
INV_X4 _u0_U15493  ( .A(1'b1), .ZN(_u0_pointer16[22] ) );
INV_X4 _u0_U15491  ( .A(1'b1), .ZN(_u0_pointer16[21] ) );
INV_X4 _u0_U15489  ( .A(1'b1), .ZN(_u0_pointer16[20] ) );
INV_X4 _u0_U15487  ( .A(1'b1), .ZN(_u0_pointer16[19] ) );
INV_X4 _u0_U15485  ( .A(1'b1), .ZN(_u0_pointer16[18] ) );
INV_X4 _u0_U15483  ( .A(1'b1), .ZN(_u0_pointer16[17] ) );
INV_X4 _u0_U15481  ( .A(1'b1), .ZN(_u0_pointer16[16] ) );
INV_X4 _u0_U15479  ( .A(1'b1), .ZN(_u0_pointer16[15] ) );
INV_X4 _u0_U15477  ( .A(1'b1), .ZN(_u0_pointer16[14] ) );
INV_X4 _u0_U15475  ( .A(1'b1), .ZN(_u0_pointer16[13] ) );
INV_X4 _u0_U15473  ( .A(1'b1), .ZN(_u0_pointer16[12] ) );
INV_X4 _u0_U15471  ( .A(1'b1), .ZN(_u0_pointer16[11] ) );
INV_X4 _u0_U15469  ( .A(1'b1), .ZN(_u0_pointer16[10] ) );
INV_X4 _u0_U15467  ( .A(1'b1), .ZN(_u0_pointer16[9] ) );
INV_X4 _u0_U15465  ( .A(1'b1), .ZN(_u0_pointer16[8] ) );
INV_X4 _u0_U15463  ( .A(1'b1), .ZN(_u0_pointer16[7] ) );
INV_X4 _u0_U15461  ( .A(1'b1), .ZN(_u0_pointer16[6] ) );
INV_X4 _u0_U15459  ( .A(1'b1), .ZN(_u0_pointer16[5] ) );
INV_X4 _u0_U15457  ( .A(1'b1), .ZN(_u0_pointer16[4] ) );
INV_X4 _u0_U15455  ( .A(1'b1), .ZN(_u0_pointer16[3] ) );
INV_X4 _u0_U15453  ( .A(1'b1), .ZN(_u0_pointer16[2] ) );
INV_X4 _u0_U15451  ( .A(1'b1), .ZN(_u0_pointer16[1] ) );
INV_X4 _u0_U15449  ( .A(1'b1), .ZN(_u0_pointer16[0] ) );
INV_X4 _u0_U15447  ( .A(1'b1), .ZN(_u0_pointer16_s[31] ) );
INV_X4 _u0_U15445  ( .A(1'b1), .ZN(_u0_pointer16_s[30] ) );
INV_X4 _u0_U15443  ( .A(1'b1), .ZN(_u0_pointer16_s[29] ) );
INV_X4 _u0_U15441  ( .A(1'b1), .ZN(_u0_pointer16_s[28] ) );
INV_X4 _u0_U15439  ( .A(1'b1), .ZN(_u0_pointer16_s[27] ) );
INV_X4 _u0_U15437  ( .A(1'b1), .ZN(_u0_pointer16_s[26] ) );
INV_X4 _u0_U15435  ( .A(1'b1), .ZN(_u0_pointer16_s[25] ) );
INV_X4 _u0_U15433  ( .A(1'b1), .ZN(_u0_pointer16_s[24] ) );
INV_X4 _u0_U15431  ( .A(1'b1), .ZN(_u0_pointer16_s[23] ) );
INV_X4 _u0_U15429  ( .A(1'b1), .ZN(_u0_pointer16_s[22] ) );
INV_X4 _u0_U15427  ( .A(1'b1), .ZN(_u0_pointer16_s[21] ) );
INV_X4 _u0_U15425  ( .A(1'b1), .ZN(_u0_pointer16_s[20] ) );
INV_X4 _u0_U15423  ( .A(1'b1), .ZN(_u0_pointer16_s[19] ) );
INV_X4 _u0_U15421  ( .A(1'b1), .ZN(_u0_pointer16_s[18] ) );
INV_X4 _u0_U15419  ( .A(1'b1), .ZN(_u0_pointer16_s[17] ) );
INV_X4 _u0_U15417  ( .A(1'b1), .ZN(_u0_pointer16_s[16] ) );
INV_X4 _u0_U15415  ( .A(1'b1), .ZN(_u0_pointer16_s[15] ) );
INV_X4 _u0_U15413  ( .A(1'b1), .ZN(_u0_pointer16_s[14] ) );
INV_X4 _u0_U15411  ( .A(1'b1), .ZN(_u0_pointer16_s[13] ) );
INV_X4 _u0_U15409  ( .A(1'b1), .ZN(_u0_pointer16_s[12] ) );
INV_X4 _u0_U15407  ( .A(1'b1), .ZN(_u0_pointer16_s[11] ) );
INV_X4 _u0_U15405  ( .A(1'b1), .ZN(_u0_pointer16_s[10] ) );
INV_X4 _u0_U15403  ( .A(1'b1), .ZN(_u0_pointer16_s[9] ) );
INV_X4 _u0_U15401  ( .A(1'b1), .ZN(_u0_pointer16_s[8] ) );
INV_X4 _u0_U15399  ( .A(1'b1), .ZN(_u0_pointer16_s[7] ) );
INV_X4 _u0_U15397  ( .A(1'b1), .ZN(_u0_pointer16_s[6] ) );
INV_X4 _u0_U15395  ( .A(1'b1), .ZN(_u0_pointer16_s[5] ) );
INV_X4 _u0_U15393  ( .A(1'b1), .ZN(_u0_pointer16_s[4] ) );
INV_X4 _u0_U15391  ( .A(1'b1), .ZN(_u0_pointer16_s[3] ) );
INV_X4 _u0_U15389  ( .A(1'b1), .ZN(_u0_pointer16_s[2] ) );
INV_X4 _u0_U15387  ( .A(1'b1), .ZN(_u0_pointer16_s[1] ) );
INV_X4 _u0_U15385  ( .A(1'b1), .ZN(_u0_pointer16_s[0] ) );
INV_X4 _u0_U15383  ( .A(1'b1), .ZN(_u0_ch16_csr[31] ) );
INV_X4 _u0_U15381  ( .A(1'b1), .ZN(_u0_ch16_csr[30] ) );
INV_X4 _u0_U15379  ( .A(1'b1), .ZN(_u0_ch16_csr[29] ) );
INV_X4 _u0_U15377  ( .A(1'b1), .ZN(_u0_ch16_csr[28] ) );
INV_X4 _u0_U15375  ( .A(1'b1), .ZN(_u0_ch16_csr[27] ) );
INV_X4 _u0_U15373  ( .A(1'b1), .ZN(_u0_ch16_csr[26] ) );
INV_X4 _u0_U15371  ( .A(1'b1), .ZN(_u0_ch16_csr[25] ) );
INV_X4 _u0_U15369  ( .A(1'b1), .ZN(_u0_ch16_csr[24] ) );
INV_X4 _u0_U15367  ( .A(1'b1), .ZN(_u0_ch16_csr[23] ) );
INV_X4 _u0_U15365  ( .A(1'b1), .ZN(_u0_ch16_csr[22] ) );
INV_X4 _u0_U15363  ( .A(1'b1), .ZN(_u0_ch16_csr[21] ) );
INV_X4 _u0_U15361  ( .A(1'b1), .ZN(_u0_ch16_csr[20] ) );
INV_X4 _u0_U15359  ( .A(1'b1), .ZN(_u0_ch16_csr[19] ) );
INV_X4 _u0_U15357  ( .A(1'b1), .ZN(_u0_ch16_csr[18] ) );
INV_X4 _u0_U15355  ( .A(1'b1), .ZN(_u0_ch16_csr[17] ) );
INV_X4 _u0_U15353  ( .A(1'b1), .ZN(_u0_ch16_csr[16] ) );
INV_X4 _u0_U15351  ( .A(1'b1), .ZN(_u0_ch16_csr[15] ) );
INV_X4 _u0_U15349  ( .A(1'b1), .ZN(_u0_ch16_csr[14] ) );
INV_X4 _u0_U15347  ( .A(1'b1), .ZN(_u0_ch16_csr[13] ) );
INV_X4 _u0_U15345  ( .A(1'b1), .ZN(_u0_ch16_csr[12] ) );
INV_X4 _u0_U15343  ( .A(1'b1), .ZN(_u0_ch16_csr[11] ) );
INV_X4 _u0_U15341  ( .A(1'b1), .ZN(_u0_ch16_csr[10] ) );
INV_X4 _u0_U15339  ( .A(1'b1), .ZN(_u0_ch16_csr[9] ) );
INV_X4 _u0_U15337  ( .A(1'b1), .ZN(_u0_ch16_csr[8] ) );
INV_X4 _u0_U15335  ( .A(1'b1), .ZN(_u0_ch16_csr[7] ) );
INV_X4 _u0_U15333  ( .A(1'b1), .ZN(_u0_ch16_csr[6] ) );
INV_X4 _u0_U15331  ( .A(1'b1), .ZN(_u0_ch16_csr[5] ) );
INV_X4 _u0_U15329  ( .A(1'b1), .ZN(_u0_ch16_csr[4] ) );
INV_X4 _u0_U15327  ( .A(1'b1), .ZN(_u0_ch16_csr[3] ) );
INV_X4 _u0_U15325  ( .A(1'b1), .ZN(_u0_ch16_csr[2] ) );
INV_X4 _u0_U15323  ( .A(1'b1), .ZN(_u0_ch16_csr[1] ) );
INV_X4 _u0_U15321  ( .A(1'b1), .ZN(_u0_ch16_csr[0] ) );
INV_X4 _u0_U15319  ( .A(1'b1), .ZN(_u0_ch16_txsz[31] ) );
INV_X4 _u0_U15317  ( .A(1'b1), .ZN(_u0_ch16_txsz[30] ) );
INV_X4 _u0_U15315  ( .A(1'b1), .ZN(_u0_ch16_txsz[29] ) );
INV_X4 _u0_U15313  ( .A(1'b1), .ZN(_u0_ch16_txsz[28] ) );
INV_X4 _u0_U15311  ( .A(1'b1), .ZN(_u0_ch16_txsz[27] ) );
INV_X4 _u0_U15309  ( .A(1'b1), .ZN(_u0_ch16_txsz[26] ) );
INV_X4 _u0_U15307  ( .A(1'b1), .ZN(_u0_ch16_txsz[25] ) );
INV_X4 _u0_U15305  ( .A(1'b1), .ZN(_u0_ch16_txsz[24] ) );
INV_X4 _u0_U15303  ( .A(1'b1), .ZN(_u0_ch16_txsz[23] ) );
INV_X4 _u0_U15301  ( .A(1'b1), .ZN(_u0_ch16_txsz[22] ) );
INV_X4 _u0_U15299  ( .A(1'b1), .ZN(_u0_ch16_txsz[21] ) );
INV_X4 _u0_U15297  ( .A(1'b1), .ZN(_u0_ch16_txsz[20] ) );
INV_X4 _u0_U15295  ( .A(1'b1), .ZN(_u0_ch16_txsz[19] ) );
INV_X4 _u0_U15293  ( .A(1'b1), .ZN(_u0_ch16_txsz[18] ) );
INV_X4 _u0_U15291  ( .A(1'b1), .ZN(_u0_ch16_txsz[17] ) );
INV_X4 _u0_U15289  ( .A(1'b1), .ZN(_u0_ch16_txsz[16] ) );
INV_X4 _u0_U15287  ( .A(1'b1), .ZN(_u0_ch16_txsz[15] ) );
INV_X4 _u0_U15285  ( .A(1'b1), .ZN(_u0_ch16_txsz[14] ) );
INV_X4 _u0_U15283  ( .A(1'b1), .ZN(_u0_ch16_txsz[13] ) );
INV_X4 _u0_U15281  ( .A(1'b1), .ZN(_u0_ch16_txsz[12] ) );
INV_X4 _u0_U15279  ( .A(1'b1), .ZN(_u0_ch16_txsz[11] ) );
INV_X4 _u0_U15277  ( .A(1'b1), .ZN(_u0_ch16_txsz[10] ) );
INV_X4 _u0_U15275  ( .A(1'b1), .ZN(_u0_ch16_txsz[9] ) );
INV_X4 _u0_U15273  ( .A(1'b1), .ZN(_u0_ch16_txsz[8] ) );
INV_X4 _u0_U15271  ( .A(1'b1), .ZN(_u0_ch16_txsz[7] ) );
INV_X4 _u0_U15269  ( .A(1'b1), .ZN(_u0_ch16_txsz[6] ) );
INV_X4 _u0_U15267  ( .A(1'b1), .ZN(_u0_ch16_txsz[5] ) );
INV_X4 _u0_U15265  ( .A(1'b1), .ZN(_u0_ch16_txsz[4] ) );
INV_X4 _u0_U15263  ( .A(1'b1), .ZN(_u0_ch16_txsz[3] ) );
INV_X4 _u0_U15261  ( .A(1'b1), .ZN(_u0_ch16_txsz[2] ) );
INV_X4 _u0_U15259  ( .A(1'b1), .ZN(_u0_ch16_txsz[1] ) );
INV_X4 _u0_U15257  ( .A(1'b1), .ZN(_u0_ch16_txsz[0] ) );
INV_X4 _u0_U15255  ( .A(1'b1), .ZN(_u0_ch16_adr0[31] ) );
INV_X4 _u0_U15253  ( .A(1'b1), .ZN(_u0_ch16_adr0[30] ) );
INV_X4 _u0_U15251  ( .A(1'b1), .ZN(_u0_ch16_adr0[29] ) );
INV_X4 _u0_U15249  ( .A(1'b1), .ZN(_u0_ch16_adr0[28] ) );
INV_X4 _u0_U15247  ( .A(1'b1), .ZN(_u0_ch16_adr0[27] ) );
INV_X4 _u0_U15245  ( .A(1'b1), .ZN(_u0_ch16_adr0[26] ) );
INV_X4 _u0_U15243  ( .A(1'b1), .ZN(_u0_ch16_adr0[25] ) );
INV_X4 _u0_U15241  ( .A(1'b1), .ZN(_u0_ch16_adr0[24] ) );
INV_X4 _u0_U15239  ( .A(1'b1), .ZN(_u0_ch16_adr0[23] ) );
INV_X4 _u0_U15237  ( .A(1'b1), .ZN(_u0_ch16_adr0[22] ) );
INV_X4 _u0_U15235  ( .A(1'b1), .ZN(_u0_ch16_adr0[21] ) );
INV_X4 _u0_U15233  ( .A(1'b1), .ZN(_u0_ch16_adr0[20] ) );
INV_X4 _u0_U15231  ( .A(1'b1), .ZN(_u0_ch16_adr0[19] ) );
INV_X4 _u0_U15229  ( .A(1'b1), .ZN(_u0_ch16_adr0[18] ) );
INV_X4 _u0_U15227  ( .A(1'b1), .ZN(_u0_ch16_adr0[17] ) );
INV_X4 _u0_U15225  ( .A(1'b1), .ZN(_u0_ch16_adr0[16] ) );
INV_X4 _u0_U15223  ( .A(1'b1), .ZN(_u0_ch16_adr0[15] ) );
INV_X4 _u0_U15221  ( .A(1'b1), .ZN(_u0_ch16_adr0[14] ) );
INV_X4 _u0_U15219  ( .A(1'b1), .ZN(_u0_ch16_adr0[13] ) );
INV_X4 _u0_U15217  ( .A(1'b1), .ZN(_u0_ch16_adr0[12] ) );
INV_X4 _u0_U15215  ( .A(1'b1), .ZN(_u0_ch16_adr0[11] ) );
INV_X4 _u0_U15213  ( .A(1'b1), .ZN(_u0_ch16_adr0[10] ) );
INV_X4 _u0_U15211  ( .A(1'b1), .ZN(_u0_ch16_adr0[9] ) );
INV_X4 _u0_U15209  ( .A(1'b1), .ZN(_u0_ch16_adr0[8] ) );
INV_X4 _u0_U15207  ( .A(1'b1), .ZN(_u0_ch16_adr0[7] ) );
INV_X4 _u0_U15205  ( .A(1'b1), .ZN(_u0_ch16_adr0[6] ) );
INV_X4 _u0_U15203  ( .A(1'b1), .ZN(_u0_ch16_adr0[5] ) );
INV_X4 _u0_U15201  ( .A(1'b1), .ZN(_u0_ch16_adr0[4] ) );
INV_X4 _u0_U15199  ( .A(1'b1), .ZN(_u0_ch16_adr0[3] ) );
INV_X4 _u0_U15197  ( .A(1'b1), .ZN(_u0_ch16_adr0[2] ) );
INV_X4 _u0_U15195  ( .A(1'b1), .ZN(_u0_ch16_adr0[1] ) );
INV_X4 _u0_U15193  ( .A(1'b1), .ZN(_u0_ch16_adr0[0] ) );
INV_X4 _u0_U15191  ( .A(1'b1), .ZN(_u0_ch16_adr1[31] ) );
INV_X4 _u0_U15189  ( .A(1'b1), .ZN(_u0_ch16_adr1[30] ) );
INV_X4 _u0_U15187  ( .A(1'b1), .ZN(_u0_ch16_adr1[29] ) );
INV_X4 _u0_U15185  ( .A(1'b1), .ZN(_u0_ch16_adr1[28] ) );
INV_X4 _u0_U15183  ( .A(1'b1), .ZN(_u0_ch16_adr1[27] ) );
INV_X4 _u0_U15181  ( .A(1'b1), .ZN(_u0_ch16_adr1[26] ) );
INV_X4 _u0_U15179  ( .A(1'b1), .ZN(_u0_ch16_adr1[25] ) );
INV_X4 _u0_U15177  ( .A(1'b1), .ZN(_u0_ch16_adr1[24] ) );
INV_X4 _u0_U15175  ( .A(1'b1), .ZN(_u0_ch16_adr1[23] ) );
INV_X4 _u0_U15173  ( .A(1'b1), .ZN(_u0_ch16_adr1[22] ) );
INV_X4 _u0_U15171  ( .A(1'b1), .ZN(_u0_ch16_adr1[21] ) );
INV_X4 _u0_U15169  ( .A(1'b1), .ZN(_u0_ch16_adr1[20] ) );
INV_X4 _u0_U15167  ( .A(1'b1), .ZN(_u0_ch16_adr1[19] ) );
INV_X4 _u0_U15165  ( .A(1'b1), .ZN(_u0_ch16_adr1[18] ) );
INV_X4 _u0_U15163  ( .A(1'b1), .ZN(_u0_ch16_adr1[17] ) );
INV_X4 _u0_U15161  ( .A(1'b1), .ZN(_u0_ch16_adr1[16] ) );
INV_X4 _u0_U15159  ( .A(1'b1), .ZN(_u0_ch16_adr1[15] ) );
INV_X4 _u0_U15157  ( .A(1'b1), .ZN(_u0_ch16_adr1[14] ) );
INV_X4 _u0_U15155  ( .A(1'b1), .ZN(_u0_ch16_adr1[13] ) );
INV_X4 _u0_U15153  ( .A(1'b1), .ZN(_u0_ch16_adr1[12] ) );
INV_X4 _u0_U15151  ( .A(1'b1), .ZN(_u0_ch16_adr1[11] ) );
INV_X4 _u0_U15149  ( .A(1'b1), .ZN(_u0_ch16_adr1[10] ) );
INV_X4 _u0_U15147  ( .A(1'b1), .ZN(_u0_ch16_adr1[9] ) );
INV_X4 _u0_U15145  ( .A(1'b1), .ZN(_u0_ch16_adr1[8] ) );
INV_X4 _u0_U15143  ( .A(1'b1), .ZN(_u0_ch16_adr1[7] ) );
INV_X4 _u0_U15141  ( .A(1'b1), .ZN(_u0_ch16_adr1[6] ) );
INV_X4 _u0_U15139  ( .A(1'b1), .ZN(_u0_ch16_adr1[5] ) );
INV_X4 _u0_U15137  ( .A(1'b1), .ZN(_u0_ch16_adr1[4] ) );
INV_X4 _u0_U15135  ( .A(1'b1), .ZN(_u0_ch16_adr1[3] ) );
INV_X4 _u0_U15133  ( .A(1'b1), .ZN(_u0_ch16_adr1[2] ) );
INV_X4 _u0_U15131  ( .A(1'b1), .ZN(_u0_ch16_adr1[1] ) );
INV_X4 _u0_U15129  ( .A(1'b1), .ZN(_u0_ch16_adr1[0] ) );
INV_X4 _u0_U15127  ( .A(1'b0), .ZN(_u0_ch16_am0[31] ) );
INV_X4 _u0_U15125  ( .A(1'b0), .ZN(_u0_ch16_am0[30] ) );
INV_X4 _u0_U15123  ( .A(1'b0), .ZN(_u0_ch16_am0[29] ) );
INV_X4 _u0_U15121  ( .A(1'b0), .ZN(_u0_ch16_am0[28] ) );
INV_X4 _u0_U15119  ( .A(1'b0), .ZN(_u0_ch16_am0[27] ) );
INV_X4 _u0_U15117  ( .A(1'b0), .ZN(_u0_ch16_am0[26] ) );
INV_X4 _u0_U15115  ( .A(1'b0), .ZN(_u0_ch16_am0[25] ) );
INV_X4 _u0_U15113  ( .A(1'b0), .ZN(_u0_ch16_am0[24] ) );
INV_X4 _u0_U15111  ( .A(1'b0), .ZN(_u0_ch16_am0[23] ) );
INV_X4 _u0_U15109  ( .A(1'b0), .ZN(_u0_ch16_am0[22] ) );
INV_X4 _u0_U15107  ( .A(1'b0), .ZN(_u0_ch16_am0[21] ) );
INV_X4 _u0_U15105  ( .A(1'b0), .ZN(_u0_ch16_am0[20] ) );
INV_X4 _u0_U15103  ( .A(1'b0), .ZN(_u0_ch16_am0[19] ) );
INV_X4 _u0_U15101  ( .A(1'b0), .ZN(_u0_ch16_am0[18] ) );
INV_X4 _u0_U15099  ( .A(1'b0), .ZN(_u0_ch16_am0[17] ) );
INV_X4 _u0_U15097  ( .A(1'b0), .ZN(_u0_ch16_am0[16] ) );
INV_X4 _u0_U15095  ( .A(1'b0), .ZN(_u0_ch16_am0[15] ) );
INV_X4 _u0_U15093  ( .A(1'b0), .ZN(_u0_ch16_am0[14] ) );
INV_X4 _u0_U15091  ( .A(1'b0), .ZN(_u0_ch16_am0[13] ) );
INV_X4 _u0_U15089  ( .A(1'b0), .ZN(_u0_ch16_am0[12] ) );
INV_X4 _u0_U15087  ( .A(1'b0), .ZN(_u0_ch16_am0[11] ) );
INV_X4 _u0_U15085  ( .A(1'b0), .ZN(_u0_ch16_am0[10] ) );
INV_X4 _u0_U15083  ( .A(1'b0), .ZN(_u0_ch16_am0[9] ) );
INV_X4 _u0_U15081  ( .A(1'b0), .ZN(_u0_ch16_am0[8] ) );
INV_X4 _u0_U15079  ( .A(1'b0), .ZN(_u0_ch16_am0[7] ) );
INV_X4 _u0_U15077  ( .A(1'b0), .ZN(_u0_ch16_am0[6] ) );
INV_X4 _u0_U15075  ( .A(1'b0), .ZN(_u0_ch16_am0[5] ) );
INV_X4 _u0_U15073  ( .A(1'b0), .ZN(_u0_ch16_am0[4] ) );
INV_X4 _u0_U15071  ( .A(1'b1), .ZN(_u0_ch16_am0[3] ) );
INV_X4 _u0_U15069  ( .A(1'b1), .ZN(_u0_ch16_am0[2] ) );
INV_X4 _u0_U15067  ( .A(1'b1), .ZN(_u0_ch16_am0[1] ) );
INV_X4 _u0_U15065  ( .A(1'b1), .ZN(_u0_ch16_am0[0] ) );
INV_X4 _u0_U15063  ( .A(1'b0), .ZN(_u0_ch16_am1[31] ) );
INV_X4 _u0_U15061  ( .A(1'b0), .ZN(_u0_ch16_am1[30] ) );
INV_X4 _u0_U15059  ( .A(1'b0), .ZN(_u0_ch16_am1[29] ) );
INV_X4 _u0_U15057  ( .A(1'b0), .ZN(_u0_ch16_am1[28] ) );
INV_X4 _u0_U15055  ( .A(1'b0), .ZN(_u0_ch16_am1[27] ) );
INV_X4 _u0_U15053  ( .A(1'b0), .ZN(_u0_ch16_am1[26] ) );
INV_X4 _u0_U15051  ( .A(1'b0), .ZN(_u0_ch16_am1[25] ) );
INV_X4 _u0_U15049  ( .A(1'b0), .ZN(_u0_ch16_am1[24] ) );
INV_X4 _u0_U15047  ( .A(1'b0), .ZN(_u0_ch16_am1[23] ) );
INV_X4 _u0_U15045  ( .A(1'b0), .ZN(_u0_ch16_am1[22] ) );
INV_X4 _u0_U15043  ( .A(1'b0), .ZN(_u0_ch16_am1[21] ) );
INV_X4 _u0_U15041  ( .A(1'b0), .ZN(_u0_ch16_am1[20] ) );
INV_X4 _u0_U15039  ( .A(1'b0), .ZN(_u0_ch16_am1[19] ) );
INV_X4 _u0_U15037  ( .A(1'b0), .ZN(_u0_ch16_am1[18] ) );
INV_X4 _u0_U15035  ( .A(1'b0), .ZN(_u0_ch16_am1[17] ) );
INV_X4 _u0_U15033  ( .A(1'b0), .ZN(_u0_ch16_am1[16] ) );
INV_X4 _u0_U15031  ( .A(1'b0), .ZN(_u0_ch16_am1[15] ) );
INV_X4 _u0_U15029  ( .A(1'b0), .ZN(_u0_ch16_am1[14] ) );
INV_X4 _u0_U15027  ( .A(1'b0), .ZN(_u0_ch16_am1[13] ) );
INV_X4 _u0_U15025  ( .A(1'b0), .ZN(_u0_ch16_am1[12] ) );
INV_X4 _u0_U15023  ( .A(1'b0), .ZN(_u0_ch16_am1[11] ) );
INV_X4 _u0_U15021  ( .A(1'b0), .ZN(_u0_ch16_am1[10] ) );
INV_X4 _u0_U15019  ( .A(1'b0), .ZN(_u0_ch16_am1[9] ) );
INV_X4 _u0_U15017  ( .A(1'b0), .ZN(_u0_ch16_am1[8] ) );
INV_X4 _u0_U15015  ( .A(1'b0), .ZN(_u0_ch16_am1[7] ) );
INV_X4 _u0_U15013  ( .A(1'b0), .ZN(_u0_ch16_am1[6] ) );
INV_X4 _u0_U15011  ( .A(1'b0), .ZN(_u0_ch16_am1[5] ) );
INV_X4 _u0_U15009  ( .A(1'b0), .ZN(_u0_ch16_am1[4] ) );
INV_X4 _u0_U15007  ( .A(1'b1), .ZN(_u0_ch16_am1[3] ) );
INV_X4 _u0_U15005  ( .A(1'b1), .ZN(_u0_ch16_am1[2] ) );
INV_X4 _u0_U15003  ( .A(1'b1), .ZN(_u0_ch16_am1[1] ) );
INV_X4 _u0_U15001  ( .A(1'b1), .ZN(_u0_ch16_am1[0] ) );
INV_X4 _u0_U14999  ( .A(1'b1), .ZN(_u0_pointer17[31] ) );
INV_X4 _u0_U14997  ( .A(1'b1), .ZN(_u0_pointer17[30] ) );
INV_X4 _u0_U14995  ( .A(1'b1), .ZN(_u0_pointer17[29] ) );
INV_X4 _u0_U14993  ( .A(1'b1), .ZN(_u0_pointer17[28] ) );
INV_X4 _u0_U14991  ( .A(1'b1), .ZN(_u0_pointer17[27] ) );
INV_X4 _u0_U14989  ( .A(1'b1), .ZN(_u0_pointer17[26] ) );
INV_X4 _u0_U14987  ( .A(1'b1), .ZN(_u0_pointer17[25] ) );
INV_X4 _u0_U14985  ( .A(1'b1), .ZN(_u0_pointer17[24] ) );
INV_X4 _u0_U14983  ( .A(1'b1), .ZN(_u0_pointer17[23] ) );
INV_X4 _u0_U14981  ( .A(1'b1), .ZN(_u0_pointer17[22] ) );
INV_X4 _u0_U14979  ( .A(1'b1), .ZN(_u0_pointer17[21] ) );
INV_X4 _u0_U14977  ( .A(1'b1), .ZN(_u0_pointer17[20] ) );
INV_X4 _u0_U14975  ( .A(1'b1), .ZN(_u0_pointer17[19] ) );
INV_X4 _u0_U14973  ( .A(1'b1), .ZN(_u0_pointer17[18] ) );
INV_X4 _u0_U14971  ( .A(1'b1), .ZN(_u0_pointer17[17] ) );
INV_X4 _u0_U14969  ( .A(1'b1), .ZN(_u0_pointer17[16] ) );
INV_X4 _u0_U14967  ( .A(1'b1), .ZN(_u0_pointer17[15] ) );
INV_X4 _u0_U14965  ( .A(1'b1), .ZN(_u0_pointer17[14] ) );
INV_X4 _u0_U14963  ( .A(1'b1), .ZN(_u0_pointer17[13] ) );
INV_X4 _u0_U14961  ( .A(1'b1), .ZN(_u0_pointer17[12] ) );
INV_X4 _u0_U14959  ( .A(1'b1), .ZN(_u0_pointer17[11] ) );
INV_X4 _u0_U14957  ( .A(1'b1), .ZN(_u0_pointer17[10] ) );
INV_X4 _u0_U14955  ( .A(1'b1), .ZN(_u0_pointer17[9] ) );
INV_X4 _u0_U14953  ( .A(1'b1), .ZN(_u0_pointer17[8] ) );
INV_X4 _u0_U14951  ( .A(1'b1), .ZN(_u0_pointer17[7] ) );
INV_X4 _u0_U14949  ( .A(1'b1), .ZN(_u0_pointer17[6] ) );
INV_X4 _u0_U14947  ( .A(1'b1), .ZN(_u0_pointer17[5] ) );
INV_X4 _u0_U14945  ( .A(1'b1), .ZN(_u0_pointer17[4] ) );
INV_X4 _u0_U14943  ( .A(1'b1), .ZN(_u0_pointer17[3] ) );
INV_X4 _u0_U14941  ( .A(1'b1), .ZN(_u0_pointer17[2] ) );
INV_X4 _u0_U14939  ( .A(1'b1), .ZN(_u0_pointer17[1] ) );
INV_X4 _u0_U14937  ( .A(1'b1), .ZN(_u0_pointer17[0] ) );
INV_X4 _u0_U14935  ( .A(1'b1), .ZN(_u0_pointer17_s[31] ) );
INV_X4 _u0_U14933  ( .A(1'b1), .ZN(_u0_pointer17_s[30] ) );
INV_X4 _u0_U14931  ( .A(1'b1), .ZN(_u0_pointer17_s[29] ) );
INV_X4 _u0_U14929  ( .A(1'b1), .ZN(_u0_pointer17_s[28] ) );
INV_X4 _u0_U14927  ( .A(1'b1), .ZN(_u0_pointer17_s[27] ) );
INV_X4 _u0_U14925  ( .A(1'b1), .ZN(_u0_pointer17_s[26] ) );
INV_X4 _u0_U14923  ( .A(1'b1), .ZN(_u0_pointer17_s[25] ) );
INV_X4 _u0_U14921  ( .A(1'b1), .ZN(_u0_pointer17_s[24] ) );
INV_X4 _u0_U14919  ( .A(1'b1), .ZN(_u0_pointer17_s[23] ) );
INV_X4 _u0_U14917  ( .A(1'b1), .ZN(_u0_pointer17_s[22] ) );
INV_X4 _u0_U14915  ( .A(1'b1), .ZN(_u0_pointer17_s[21] ) );
INV_X4 _u0_U14913  ( .A(1'b1), .ZN(_u0_pointer17_s[20] ) );
INV_X4 _u0_U14911  ( .A(1'b1), .ZN(_u0_pointer17_s[19] ) );
INV_X4 _u0_U14909  ( .A(1'b1), .ZN(_u0_pointer17_s[18] ) );
INV_X4 _u0_U14907  ( .A(1'b1), .ZN(_u0_pointer17_s[17] ) );
INV_X4 _u0_U14905  ( .A(1'b1), .ZN(_u0_pointer17_s[16] ) );
INV_X4 _u0_U14903  ( .A(1'b1), .ZN(_u0_pointer17_s[15] ) );
INV_X4 _u0_U14901  ( .A(1'b1), .ZN(_u0_pointer17_s[14] ) );
INV_X4 _u0_U14899  ( .A(1'b1), .ZN(_u0_pointer17_s[13] ) );
INV_X4 _u0_U14897  ( .A(1'b1), .ZN(_u0_pointer17_s[12] ) );
INV_X4 _u0_U14895  ( .A(1'b1), .ZN(_u0_pointer17_s[11] ) );
INV_X4 _u0_U14893  ( .A(1'b1), .ZN(_u0_pointer17_s[10] ) );
INV_X4 _u0_U14891  ( .A(1'b1), .ZN(_u0_pointer17_s[9] ) );
INV_X4 _u0_U14889  ( .A(1'b1), .ZN(_u0_pointer17_s[8] ) );
INV_X4 _u0_U14887  ( .A(1'b1), .ZN(_u0_pointer17_s[7] ) );
INV_X4 _u0_U14885  ( .A(1'b1), .ZN(_u0_pointer17_s[6] ) );
INV_X4 _u0_U14883  ( .A(1'b1), .ZN(_u0_pointer17_s[5] ) );
INV_X4 _u0_U14881  ( .A(1'b1), .ZN(_u0_pointer17_s[4] ) );
INV_X4 _u0_U14879  ( .A(1'b1), .ZN(_u0_pointer17_s[3] ) );
INV_X4 _u0_U14877  ( .A(1'b1), .ZN(_u0_pointer17_s[2] ) );
INV_X4 _u0_U14875  ( .A(1'b1), .ZN(_u0_pointer17_s[1] ) );
INV_X4 _u0_U14873  ( .A(1'b1), .ZN(_u0_pointer17_s[0] ) );
INV_X4 _u0_U14871  ( .A(1'b1), .ZN(_u0_ch17_csr[31] ) );
INV_X4 _u0_U14869  ( .A(1'b1), .ZN(_u0_ch17_csr[30] ) );
INV_X4 _u0_U14867  ( .A(1'b1), .ZN(_u0_ch17_csr[29] ) );
INV_X4 _u0_U14865  ( .A(1'b1), .ZN(_u0_ch17_csr[28] ) );
INV_X4 _u0_U14863  ( .A(1'b1), .ZN(_u0_ch17_csr[27] ) );
INV_X4 _u0_U14861  ( .A(1'b1), .ZN(_u0_ch17_csr[26] ) );
INV_X4 _u0_U14859  ( .A(1'b1), .ZN(_u0_ch17_csr[25] ) );
INV_X4 _u0_U14857  ( .A(1'b1), .ZN(_u0_ch17_csr[24] ) );
INV_X4 _u0_U14855  ( .A(1'b1), .ZN(_u0_ch17_csr[23] ) );
INV_X4 _u0_U14853  ( .A(1'b1), .ZN(_u0_ch17_csr[22] ) );
INV_X4 _u0_U14851  ( .A(1'b1), .ZN(_u0_ch17_csr[21] ) );
INV_X4 _u0_U14849  ( .A(1'b1), .ZN(_u0_ch17_csr[20] ) );
INV_X4 _u0_U14847  ( .A(1'b1), .ZN(_u0_ch17_csr[19] ) );
INV_X4 _u0_U14845  ( .A(1'b1), .ZN(_u0_ch17_csr[18] ) );
INV_X4 _u0_U14843  ( .A(1'b1), .ZN(_u0_ch17_csr[17] ) );
INV_X4 _u0_U14841  ( .A(1'b1), .ZN(_u0_ch17_csr[16] ) );
INV_X4 _u0_U14839  ( .A(1'b1), .ZN(_u0_ch17_csr[15] ) );
INV_X4 _u0_U14837  ( .A(1'b1), .ZN(_u0_ch17_csr[14] ) );
INV_X4 _u0_U14835  ( .A(1'b1), .ZN(_u0_ch17_csr[13] ) );
INV_X4 _u0_U14833  ( .A(1'b1), .ZN(_u0_ch17_csr[12] ) );
INV_X4 _u0_U14831  ( .A(1'b1), .ZN(_u0_ch17_csr[11] ) );
INV_X4 _u0_U14829  ( .A(1'b1), .ZN(_u0_ch17_csr[10] ) );
INV_X4 _u0_U14827  ( .A(1'b1), .ZN(_u0_ch17_csr[9] ) );
INV_X4 _u0_U14825  ( .A(1'b1), .ZN(_u0_ch17_csr[8] ) );
INV_X4 _u0_U14823  ( .A(1'b1), .ZN(_u0_ch17_csr[7] ) );
INV_X4 _u0_U14821  ( .A(1'b1), .ZN(_u0_ch17_csr[6] ) );
INV_X4 _u0_U14819  ( .A(1'b1), .ZN(_u0_ch17_csr[5] ) );
INV_X4 _u0_U14817  ( .A(1'b1), .ZN(_u0_ch17_csr[4] ) );
INV_X4 _u0_U14815  ( .A(1'b1), .ZN(_u0_ch17_csr[3] ) );
INV_X4 _u0_U14813  ( .A(1'b1), .ZN(_u0_ch17_csr[2] ) );
INV_X4 _u0_U14811  ( .A(1'b1), .ZN(_u0_ch17_csr[1] ) );
INV_X4 _u0_U14809  ( .A(1'b1), .ZN(_u0_ch17_csr[0] ) );
INV_X4 _u0_U14807  ( .A(1'b1), .ZN(_u0_ch17_txsz[31] ) );
INV_X4 _u0_U14805  ( .A(1'b1), .ZN(_u0_ch17_txsz[30] ) );
INV_X4 _u0_U14803  ( .A(1'b1), .ZN(_u0_ch17_txsz[29] ) );
INV_X4 _u0_U14801  ( .A(1'b1), .ZN(_u0_ch17_txsz[28] ) );
INV_X4 _u0_U14799  ( .A(1'b1), .ZN(_u0_ch17_txsz[27] ) );
INV_X4 _u0_U14797  ( .A(1'b1), .ZN(_u0_ch17_txsz[26] ) );
INV_X4 _u0_U14795  ( .A(1'b1), .ZN(_u0_ch17_txsz[25] ) );
INV_X4 _u0_U14793  ( .A(1'b1), .ZN(_u0_ch17_txsz[24] ) );
INV_X4 _u0_U14791  ( .A(1'b1), .ZN(_u0_ch17_txsz[23] ) );
INV_X4 _u0_U14789  ( .A(1'b1), .ZN(_u0_ch17_txsz[22] ) );
INV_X4 _u0_U14787  ( .A(1'b1), .ZN(_u0_ch17_txsz[21] ) );
INV_X4 _u0_U14785  ( .A(1'b1), .ZN(_u0_ch17_txsz[20] ) );
INV_X4 _u0_U14783  ( .A(1'b1), .ZN(_u0_ch17_txsz[19] ) );
INV_X4 _u0_U14781  ( .A(1'b1), .ZN(_u0_ch17_txsz[18] ) );
INV_X4 _u0_U14779  ( .A(1'b1), .ZN(_u0_ch17_txsz[17] ) );
INV_X4 _u0_U14777  ( .A(1'b1), .ZN(_u0_ch17_txsz[16] ) );
INV_X4 _u0_U14775  ( .A(1'b1), .ZN(_u0_ch17_txsz[15] ) );
INV_X4 _u0_U14773  ( .A(1'b1), .ZN(_u0_ch17_txsz[14] ) );
INV_X4 _u0_U14771  ( .A(1'b1), .ZN(_u0_ch17_txsz[13] ) );
INV_X4 _u0_U14769  ( .A(1'b1), .ZN(_u0_ch17_txsz[12] ) );
INV_X4 _u0_U14767  ( .A(1'b1), .ZN(_u0_ch17_txsz[11] ) );
INV_X4 _u0_U14765  ( .A(1'b1), .ZN(_u0_ch17_txsz[10] ) );
INV_X4 _u0_U14763  ( .A(1'b1), .ZN(_u0_ch17_txsz[9] ) );
INV_X4 _u0_U14761  ( .A(1'b1), .ZN(_u0_ch17_txsz[8] ) );
INV_X4 _u0_U14759  ( .A(1'b1), .ZN(_u0_ch17_txsz[7] ) );
INV_X4 _u0_U14757  ( .A(1'b1), .ZN(_u0_ch17_txsz[6] ) );
INV_X4 _u0_U14755  ( .A(1'b1), .ZN(_u0_ch17_txsz[5] ) );
INV_X4 _u0_U14753  ( .A(1'b1), .ZN(_u0_ch17_txsz[4] ) );
INV_X4 _u0_U14751  ( .A(1'b1), .ZN(_u0_ch17_txsz[3] ) );
INV_X4 _u0_U14749  ( .A(1'b1), .ZN(_u0_ch17_txsz[2] ) );
INV_X4 _u0_U14747  ( .A(1'b1), .ZN(_u0_ch17_txsz[1] ) );
INV_X4 _u0_U14745  ( .A(1'b1), .ZN(_u0_ch17_txsz[0] ) );
INV_X4 _u0_U14743  ( .A(1'b1), .ZN(_u0_ch17_adr0[31] ) );
INV_X4 _u0_U14741  ( .A(1'b1), .ZN(_u0_ch17_adr0[30] ) );
INV_X4 _u0_U14739  ( .A(1'b1), .ZN(_u0_ch17_adr0[29] ) );
INV_X4 _u0_U14737  ( .A(1'b1), .ZN(_u0_ch17_adr0[28] ) );
INV_X4 _u0_U14735  ( .A(1'b1), .ZN(_u0_ch17_adr0[27] ) );
INV_X4 _u0_U14733  ( .A(1'b1), .ZN(_u0_ch17_adr0[26] ) );
INV_X4 _u0_U14731  ( .A(1'b1), .ZN(_u0_ch17_adr0[25] ) );
INV_X4 _u0_U14729  ( .A(1'b1), .ZN(_u0_ch17_adr0[24] ) );
INV_X4 _u0_U14727  ( .A(1'b1), .ZN(_u0_ch17_adr0[23] ) );
INV_X4 _u0_U14725  ( .A(1'b1), .ZN(_u0_ch17_adr0[22] ) );
INV_X4 _u0_U14723  ( .A(1'b1), .ZN(_u0_ch17_adr0[21] ) );
INV_X4 _u0_U14721  ( .A(1'b1), .ZN(_u0_ch17_adr0[20] ) );
INV_X4 _u0_U14719  ( .A(1'b1), .ZN(_u0_ch17_adr0[19] ) );
INV_X4 _u0_U14717  ( .A(1'b1), .ZN(_u0_ch17_adr0[18] ) );
INV_X4 _u0_U14715  ( .A(1'b1), .ZN(_u0_ch17_adr0[17] ) );
INV_X4 _u0_U14713  ( .A(1'b1), .ZN(_u0_ch17_adr0[16] ) );
INV_X4 _u0_U14711  ( .A(1'b1), .ZN(_u0_ch17_adr0[15] ) );
INV_X4 _u0_U14709  ( .A(1'b1), .ZN(_u0_ch17_adr0[14] ) );
INV_X4 _u0_U14707  ( .A(1'b1), .ZN(_u0_ch17_adr0[13] ) );
INV_X4 _u0_U14705  ( .A(1'b1), .ZN(_u0_ch17_adr0[12] ) );
INV_X4 _u0_U14703  ( .A(1'b1), .ZN(_u0_ch17_adr0[11] ) );
INV_X4 _u0_U14701  ( .A(1'b1), .ZN(_u0_ch17_adr0[10] ) );
INV_X4 _u0_U14699  ( .A(1'b1), .ZN(_u0_ch17_adr0[9] ) );
INV_X4 _u0_U14697  ( .A(1'b1), .ZN(_u0_ch17_adr0[8] ) );
INV_X4 _u0_U14695  ( .A(1'b1), .ZN(_u0_ch17_adr0[7] ) );
INV_X4 _u0_U14693  ( .A(1'b1), .ZN(_u0_ch17_adr0[6] ) );
INV_X4 _u0_U14691  ( .A(1'b1), .ZN(_u0_ch17_adr0[5] ) );
INV_X4 _u0_U14689  ( .A(1'b1), .ZN(_u0_ch17_adr0[4] ) );
INV_X4 _u0_U14687  ( .A(1'b1), .ZN(_u0_ch17_adr0[3] ) );
INV_X4 _u0_U14685  ( .A(1'b1), .ZN(_u0_ch17_adr0[2] ) );
INV_X4 _u0_U14683  ( .A(1'b1), .ZN(_u0_ch17_adr0[1] ) );
INV_X4 _u0_U14681  ( .A(1'b1), .ZN(_u0_ch17_adr0[0] ) );
INV_X4 _u0_U14679  ( .A(1'b1), .ZN(_u0_ch17_adr1[31] ) );
INV_X4 _u0_U14677  ( .A(1'b1), .ZN(_u0_ch17_adr1[30] ) );
INV_X4 _u0_U14675  ( .A(1'b1), .ZN(_u0_ch17_adr1[29] ) );
INV_X4 _u0_U14673  ( .A(1'b1), .ZN(_u0_ch17_adr1[28] ) );
INV_X4 _u0_U14671  ( .A(1'b1), .ZN(_u0_ch17_adr1[27] ) );
INV_X4 _u0_U14669  ( .A(1'b1), .ZN(_u0_ch17_adr1[26] ) );
INV_X4 _u0_U14667  ( .A(1'b1), .ZN(_u0_ch17_adr1[25] ) );
INV_X4 _u0_U14665  ( .A(1'b1), .ZN(_u0_ch17_adr1[24] ) );
INV_X4 _u0_U14663  ( .A(1'b1), .ZN(_u0_ch17_adr1[23] ) );
INV_X4 _u0_U14661  ( .A(1'b1), .ZN(_u0_ch17_adr1[22] ) );
INV_X4 _u0_U14659  ( .A(1'b1), .ZN(_u0_ch17_adr1[21] ) );
INV_X4 _u0_U14657  ( .A(1'b1), .ZN(_u0_ch17_adr1[20] ) );
INV_X4 _u0_U14655  ( .A(1'b1), .ZN(_u0_ch17_adr1[19] ) );
INV_X4 _u0_U14653  ( .A(1'b1), .ZN(_u0_ch17_adr1[18] ) );
INV_X4 _u0_U14651  ( .A(1'b1), .ZN(_u0_ch17_adr1[17] ) );
INV_X4 _u0_U14649  ( .A(1'b1), .ZN(_u0_ch17_adr1[16] ) );
INV_X4 _u0_U14647  ( .A(1'b1), .ZN(_u0_ch17_adr1[15] ) );
INV_X4 _u0_U14645  ( .A(1'b1), .ZN(_u0_ch17_adr1[14] ) );
INV_X4 _u0_U14643  ( .A(1'b1), .ZN(_u0_ch17_adr1[13] ) );
INV_X4 _u0_U14641  ( .A(1'b1), .ZN(_u0_ch17_adr1[12] ) );
INV_X4 _u0_U14639  ( .A(1'b1), .ZN(_u0_ch17_adr1[11] ) );
INV_X4 _u0_U14637  ( .A(1'b1), .ZN(_u0_ch17_adr1[10] ) );
INV_X4 _u0_U14635  ( .A(1'b1), .ZN(_u0_ch17_adr1[9] ) );
INV_X4 _u0_U14633  ( .A(1'b1), .ZN(_u0_ch17_adr1[8] ) );
INV_X4 _u0_U14631  ( .A(1'b1), .ZN(_u0_ch17_adr1[7] ) );
INV_X4 _u0_U14629  ( .A(1'b1), .ZN(_u0_ch17_adr1[6] ) );
INV_X4 _u0_U14627  ( .A(1'b1), .ZN(_u0_ch17_adr1[5] ) );
INV_X4 _u0_U14625  ( .A(1'b1), .ZN(_u0_ch17_adr1[4] ) );
INV_X4 _u0_U14623  ( .A(1'b1), .ZN(_u0_ch17_adr1[3] ) );
INV_X4 _u0_U14621  ( .A(1'b1), .ZN(_u0_ch17_adr1[2] ) );
INV_X4 _u0_U14619  ( .A(1'b1), .ZN(_u0_ch17_adr1[1] ) );
INV_X4 _u0_U14617  ( .A(1'b1), .ZN(_u0_ch17_adr1[0] ) );
INV_X4 _u0_U14615  ( .A(1'b0), .ZN(_u0_ch17_am0[31] ) );
INV_X4 _u0_U14613  ( .A(1'b0), .ZN(_u0_ch17_am0[30] ) );
INV_X4 _u0_U14611  ( .A(1'b0), .ZN(_u0_ch17_am0[29] ) );
INV_X4 _u0_U14609  ( .A(1'b0), .ZN(_u0_ch17_am0[28] ) );
INV_X4 _u0_U14607  ( .A(1'b0), .ZN(_u0_ch17_am0[27] ) );
INV_X4 _u0_U14605  ( .A(1'b0), .ZN(_u0_ch17_am0[26] ) );
INV_X4 _u0_U14603  ( .A(1'b0), .ZN(_u0_ch17_am0[25] ) );
INV_X4 _u0_U14601  ( .A(1'b0), .ZN(_u0_ch17_am0[24] ) );
INV_X4 _u0_U14599  ( .A(1'b0), .ZN(_u0_ch17_am0[23] ) );
INV_X4 _u0_U14597  ( .A(1'b0), .ZN(_u0_ch17_am0[22] ) );
INV_X4 _u0_U14595  ( .A(1'b0), .ZN(_u0_ch17_am0[21] ) );
INV_X4 _u0_U14593  ( .A(1'b0), .ZN(_u0_ch17_am0[20] ) );
INV_X4 _u0_U14591  ( .A(1'b0), .ZN(_u0_ch17_am0[19] ) );
INV_X4 _u0_U14589  ( .A(1'b0), .ZN(_u0_ch17_am0[18] ) );
INV_X4 _u0_U14587  ( .A(1'b0), .ZN(_u0_ch17_am0[17] ) );
INV_X4 _u0_U14585  ( .A(1'b0), .ZN(_u0_ch17_am0[16] ) );
INV_X4 _u0_U14583  ( .A(1'b0), .ZN(_u0_ch17_am0[15] ) );
INV_X4 _u0_U14581  ( .A(1'b0), .ZN(_u0_ch17_am0[14] ) );
INV_X4 _u0_U14579  ( .A(1'b0), .ZN(_u0_ch17_am0[13] ) );
INV_X4 _u0_U14577  ( .A(1'b0), .ZN(_u0_ch17_am0[12] ) );
INV_X4 _u0_U14575  ( .A(1'b0), .ZN(_u0_ch17_am0[11] ) );
INV_X4 _u0_U14573  ( .A(1'b0), .ZN(_u0_ch17_am0[10] ) );
INV_X4 _u0_U14571  ( .A(1'b0), .ZN(_u0_ch17_am0[9] ) );
INV_X4 _u0_U14569  ( .A(1'b0), .ZN(_u0_ch17_am0[8] ) );
INV_X4 _u0_U14567  ( .A(1'b0), .ZN(_u0_ch17_am0[7] ) );
INV_X4 _u0_U14565  ( .A(1'b0), .ZN(_u0_ch17_am0[6] ) );
INV_X4 _u0_U14563  ( .A(1'b0), .ZN(_u0_ch17_am0[5] ) );
INV_X4 _u0_U14561  ( .A(1'b0), .ZN(_u0_ch17_am0[4] ) );
INV_X4 _u0_U14559  ( .A(1'b1), .ZN(_u0_ch17_am0[3] ) );
INV_X4 _u0_U14557  ( .A(1'b1), .ZN(_u0_ch17_am0[2] ) );
INV_X4 _u0_U14555  ( .A(1'b1), .ZN(_u0_ch17_am0[1] ) );
INV_X4 _u0_U14553  ( .A(1'b1), .ZN(_u0_ch17_am0[0] ) );
INV_X4 _u0_U14551  ( .A(1'b0), .ZN(_u0_ch17_am1[31] ) );
INV_X4 _u0_U14549  ( .A(1'b0), .ZN(_u0_ch17_am1[30] ) );
INV_X4 _u0_U14547  ( .A(1'b0), .ZN(_u0_ch17_am1[29] ) );
INV_X4 _u0_U14545  ( .A(1'b0), .ZN(_u0_ch17_am1[28] ) );
INV_X4 _u0_U14543  ( .A(1'b0), .ZN(_u0_ch17_am1[27] ) );
INV_X4 _u0_U14541  ( .A(1'b0), .ZN(_u0_ch17_am1[26] ) );
INV_X4 _u0_U14539  ( .A(1'b0), .ZN(_u0_ch17_am1[25] ) );
INV_X4 _u0_U14537  ( .A(1'b0), .ZN(_u0_ch17_am1[24] ) );
INV_X4 _u0_U14535  ( .A(1'b0), .ZN(_u0_ch17_am1[23] ) );
INV_X4 _u0_U14533  ( .A(1'b0), .ZN(_u0_ch17_am1[22] ) );
INV_X4 _u0_U14531  ( .A(1'b0), .ZN(_u0_ch17_am1[21] ) );
INV_X4 _u0_U14529  ( .A(1'b0), .ZN(_u0_ch17_am1[20] ) );
INV_X4 _u0_U14527  ( .A(1'b0), .ZN(_u0_ch17_am1[19] ) );
INV_X4 _u0_U14525  ( .A(1'b0), .ZN(_u0_ch17_am1[18] ) );
INV_X4 _u0_U14523  ( .A(1'b0), .ZN(_u0_ch17_am1[17] ) );
INV_X4 _u0_U14521  ( .A(1'b0), .ZN(_u0_ch17_am1[16] ) );
INV_X4 _u0_U14519  ( .A(1'b0), .ZN(_u0_ch17_am1[15] ) );
INV_X4 _u0_U14517  ( .A(1'b0), .ZN(_u0_ch17_am1[14] ) );
INV_X4 _u0_U14515  ( .A(1'b0), .ZN(_u0_ch17_am1[13] ) );
INV_X4 _u0_U14513  ( .A(1'b0), .ZN(_u0_ch17_am1[12] ) );
INV_X4 _u0_U14511  ( .A(1'b0), .ZN(_u0_ch17_am1[11] ) );
INV_X4 _u0_U14509  ( .A(1'b0), .ZN(_u0_ch17_am1[10] ) );
INV_X4 _u0_U14507  ( .A(1'b0), .ZN(_u0_ch17_am1[9] ) );
INV_X4 _u0_U14505  ( .A(1'b0), .ZN(_u0_ch17_am1[8] ) );
INV_X4 _u0_U14503  ( .A(1'b0), .ZN(_u0_ch17_am1[7] ) );
INV_X4 _u0_U14501  ( .A(1'b0), .ZN(_u0_ch17_am1[6] ) );
INV_X4 _u0_U14499  ( .A(1'b0), .ZN(_u0_ch17_am1[5] ) );
INV_X4 _u0_U14497  ( .A(1'b0), .ZN(_u0_ch17_am1[4] ) );
INV_X4 _u0_U14495  ( .A(1'b1), .ZN(_u0_ch17_am1[3] ) );
INV_X4 _u0_U14493  ( .A(1'b1), .ZN(_u0_ch17_am1[2] ) );
INV_X4 _u0_U14491  ( .A(1'b1), .ZN(_u0_ch17_am1[1] ) );
INV_X4 _u0_U14489  ( .A(1'b1), .ZN(_u0_ch17_am1[0] ) );
INV_X4 _u0_U14487  ( .A(1'b1), .ZN(_u0_pointer18[31] ) );
INV_X4 _u0_U14485  ( .A(1'b1), .ZN(_u0_pointer18[30] ) );
INV_X4 _u0_U14483  ( .A(1'b1), .ZN(_u0_pointer18[29] ) );
INV_X4 _u0_U14481  ( .A(1'b1), .ZN(_u0_pointer18[28] ) );
INV_X4 _u0_U14479  ( .A(1'b1), .ZN(_u0_pointer18[27] ) );
INV_X4 _u0_U14477  ( .A(1'b1), .ZN(_u0_pointer18[26] ) );
INV_X4 _u0_U14475  ( .A(1'b1), .ZN(_u0_pointer18[25] ) );
INV_X4 _u0_U14473  ( .A(1'b1), .ZN(_u0_pointer18[24] ) );
INV_X4 _u0_U14471  ( .A(1'b1), .ZN(_u0_pointer18[23] ) );
INV_X4 _u0_U14469  ( .A(1'b1), .ZN(_u0_pointer18[22] ) );
INV_X4 _u0_U14467  ( .A(1'b1), .ZN(_u0_pointer18[21] ) );
INV_X4 _u0_U14465  ( .A(1'b1), .ZN(_u0_pointer18[20] ) );
INV_X4 _u0_U14463  ( .A(1'b1), .ZN(_u0_pointer18[19] ) );
INV_X4 _u0_U14461  ( .A(1'b1), .ZN(_u0_pointer18[18] ) );
INV_X4 _u0_U14459  ( .A(1'b1), .ZN(_u0_pointer18[17] ) );
INV_X4 _u0_U14457  ( .A(1'b1), .ZN(_u0_pointer18[16] ) );
INV_X4 _u0_U14455  ( .A(1'b1), .ZN(_u0_pointer18[15] ) );
INV_X4 _u0_U14453  ( .A(1'b1), .ZN(_u0_pointer18[14] ) );
INV_X4 _u0_U14451  ( .A(1'b1), .ZN(_u0_pointer18[13] ) );
INV_X4 _u0_U14449  ( .A(1'b1), .ZN(_u0_pointer18[12] ) );
INV_X4 _u0_U14447  ( .A(1'b1), .ZN(_u0_pointer18[11] ) );
INV_X4 _u0_U14445  ( .A(1'b1), .ZN(_u0_pointer18[10] ) );
INV_X4 _u0_U14443  ( .A(1'b1), .ZN(_u0_pointer18[9] ) );
INV_X4 _u0_U14441  ( .A(1'b1), .ZN(_u0_pointer18[8] ) );
INV_X4 _u0_U14439  ( .A(1'b1), .ZN(_u0_pointer18[7] ) );
INV_X4 _u0_U14437  ( .A(1'b1), .ZN(_u0_pointer18[6] ) );
INV_X4 _u0_U14435  ( .A(1'b1), .ZN(_u0_pointer18[5] ) );
INV_X4 _u0_U14433  ( .A(1'b1), .ZN(_u0_pointer18[4] ) );
INV_X4 _u0_U14431  ( .A(1'b1), .ZN(_u0_pointer18[3] ) );
INV_X4 _u0_U14429  ( .A(1'b1), .ZN(_u0_pointer18[2] ) );
INV_X4 _u0_U14427  ( .A(1'b1), .ZN(_u0_pointer18[1] ) );
INV_X4 _u0_U14425  ( .A(1'b1), .ZN(_u0_pointer18[0] ) );
INV_X4 _u0_U14423  ( .A(1'b1), .ZN(_u0_pointer18_s[31] ) );
INV_X4 _u0_U14421  ( .A(1'b1), .ZN(_u0_pointer18_s[30] ) );
INV_X4 _u0_U14419  ( .A(1'b1), .ZN(_u0_pointer18_s[29] ) );
INV_X4 _u0_U14417  ( .A(1'b1), .ZN(_u0_pointer18_s[28] ) );
INV_X4 _u0_U14415  ( .A(1'b1), .ZN(_u0_pointer18_s[27] ) );
INV_X4 _u0_U14413  ( .A(1'b1), .ZN(_u0_pointer18_s[26] ) );
INV_X4 _u0_U14411  ( .A(1'b1), .ZN(_u0_pointer18_s[25] ) );
INV_X4 _u0_U14409  ( .A(1'b1), .ZN(_u0_pointer18_s[24] ) );
INV_X4 _u0_U14407  ( .A(1'b1), .ZN(_u0_pointer18_s[23] ) );
INV_X4 _u0_U14405  ( .A(1'b1), .ZN(_u0_pointer18_s[22] ) );
INV_X4 _u0_U14403  ( .A(1'b1), .ZN(_u0_pointer18_s[21] ) );
INV_X4 _u0_U14401  ( .A(1'b1), .ZN(_u0_pointer18_s[20] ) );
INV_X4 _u0_U14399  ( .A(1'b1), .ZN(_u0_pointer18_s[19] ) );
INV_X4 _u0_U14397  ( .A(1'b1), .ZN(_u0_pointer18_s[18] ) );
INV_X4 _u0_U14395  ( .A(1'b1), .ZN(_u0_pointer18_s[17] ) );
INV_X4 _u0_U14393  ( .A(1'b1), .ZN(_u0_pointer18_s[16] ) );
INV_X4 _u0_U14391  ( .A(1'b1), .ZN(_u0_pointer18_s[15] ) );
INV_X4 _u0_U14389  ( .A(1'b1), .ZN(_u0_pointer18_s[14] ) );
INV_X4 _u0_U14387  ( .A(1'b1), .ZN(_u0_pointer18_s[13] ) );
INV_X4 _u0_U14385  ( .A(1'b1), .ZN(_u0_pointer18_s[12] ) );
INV_X4 _u0_U14383  ( .A(1'b1), .ZN(_u0_pointer18_s[11] ) );
INV_X4 _u0_U14381  ( .A(1'b1), .ZN(_u0_pointer18_s[10] ) );
INV_X4 _u0_U14379  ( .A(1'b1), .ZN(_u0_pointer18_s[9] ) );
INV_X4 _u0_U14377  ( .A(1'b1), .ZN(_u0_pointer18_s[8] ) );
INV_X4 _u0_U14375  ( .A(1'b1), .ZN(_u0_pointer18_s[7] ) );
INV_X4 _u0_U14373  ( .A(1'b1), .ZN(_u0_pointer18_s[6] ) );
INV_X4 _u0_U14371  ( .A(1'b1), .ZN(_u0_pointer18_s[5] ) );
INV_X4 _u0_U14369  ( .A(1'b1), .ZN(_u0_pointer18_s[4] ) );
INV_X4 _u0_U14367  ( .A(1'b1), .ZN(_u0_pointer18_s[3] ) );
INV_X4 _u0_U14365  ( .A(1'b1), .ZN(_u0_pointer18_s[2] ) );
INV_X4 _u0_U14363  ( .A(1'b1), .ZN(_u0_pointer18_s[1] ) );
INV_X4 _u0_U14361  ( .A(1'b1), .ZN(_u0_pointer18_s[0] ) );
INV_X4 _u0_U14359  ( .A(1'b1), .ZN(_u0_ch18_csr[31] ) );
INV_X4 _u0_U14357  ( .A(1'b1), .ZN(_u0_ch18_csr[30] ) );
INV_X4 _u0_U14355  ( .A(1'b1), .ZN(_u0_ch18_csr[29] ) );
INV_X4 _u0_U14353  ( .A(1'b1), .ZN(_u0_ch18_csr[28] ) );
INV_X4 _u0_U14351  ( .A(1'b1), .ZN(_u0_ch18_csr[27] ) );
INV_X4 _u0_U14349  ( .A(1'b1), .ZN(_u0_ch18_csr[26] ) );
INV_X4 _u0_U14347  ( .A(1'b1), .ZN(_u0_ch18_csr[25] ) );
INV_X4 _u0_U14345  ( .A(1'b1), .ZN(_u0_ch18_csr[24] ) );
INV_X4 _u0_U14343  ( .A(1'b1), .ZN(_u0_ch18_csr[23] ) );
INV_X4 _u0_U14341  ( .A(1'b1), .ZN(_u0_ch18_csr[22] ) );
INV_X4 _u0_U14339  ( .A(1'b1), .ZN(_u0_ch18_csr[21] ) );
INV_X4 _u0_U14337  ( .A(1'b1), .ZN(_u0_ch18_csr[20] ) );
INV_X4 _u0_U14335  ( .A(1'b1), .ZN(_u0_ch18_csr[19] ) );
INV_X4 _u0_U14333  ( .A(1'b1), .ZN(_u0_ch18_csr[18] ) );
INV_X4 _u0_U14331  ( .A(1'b1), .ZN(_u0_ch18_csr[17] ) );
INV_X4 _u0_U14329  ( .A(1'b1), .ZN(_u0_ch18_csr[16] ) );
INV_X4 _u0_U14327  ( .A(1'b1), .ZN(_u0_ch18_csr[15] ) );
INV_X4 _u0_U14325  ( .A(1'b1), .ZN(_u0_ch18_csr[14] ) );
INV_X4 _u0_U14323  ( .A(1'b1), .ZN(_u0_ch18_csr[13] ) );
INV_X4 _u0_U14321  ( .A(1'b1), .ZN(_u0_ch18_csr[12] ) );
INV_X4 _u0_U14319  ( .A(1'b1), .ZN(_u0_ch18_csr[11] ) );
INV_X4 _u0_U14317  ( .A(1'b1), .ZN(_u0_ch18_csr[10] ) );
INV_X4 _u0_U14315  ( .A(1'b1), .ZN(_u0_ch18_csr[9] ) );
INV_X4 _u0_U14313  ( .A(1'b1), .ZN(_u0_ch18_csr[8] ) );
INV_X4 _u0_U14311  ( .A(1'b1), .ZN(_u0_ch18_csr[7] ) );
INV_X4 _u0_U14309  ( .A(1'b1), .ZN(_u0_ch18_csr[6] ) );
INV_X4 _u0_U14307  ( .A(1'b1), .ZN(_u0_ch18_csr[5] ) );
INV_X4 _u0_U14305  ( .A(1'b1), .ZN(_u0_ch18_csr[4] ) );
INV_X4 _u0_U14303  ( .A(1'b1), .ZN(_u0_ch18_csr[3] ) );
INV_X4 _u0_U14301  ( .A(1'b1), .ZN(_u0_ch18_csr[2] ) );
INV_X4 _u0_U14299  ( .A(1'b1), .ZN(_u0_ch18_csr[1] ) );
INV_X4 _u0_U14297  ( .A(1'b1), .ZN(_u0_ch18_csr[0] ) );
INV_X4 _u0_U14295  ( .A(1'b1), .ZN(_u0_ch18_txsz[31] ) );
INV_X4 _u0_U14293  ( .A(1'b1), .ZN(_u0_ch18_txsz[30] ) );
INV_X4 _u0_U14291  ( .A(1'b1), .ZN(_u0_ch18_txsz[29] ) );
INV_X4 _u0_U14289  ( .A(1'b1), .ZN(_u0_ch18_txsz[28] ) );
INV_X4 _u0_U14287  ( .A(1'b1), .ZN(_u0_ch18_txsz[27] ) );
INV_X4 _u0_U14285  ( .A(1'b1), .ZN(_u0_ch18_txsz[26] ) );
INV_X4 _u0_U14283  ( .A(1'b1), .ZN(_u0_ch18_txsz[25] ) );
INV_X4 _u0_U14281  ( .A(1'b1), .ZN(_u0_ch18_txsz[24] ) );
INV_X4 _u0_U14279  ( .A(1'b1), .ZN(_u0_ch18_txsz[23] ) );
INV_X4 _u0_U14277  ( .A(1'b1), .ZN(_u0_ch18_txsz[22] ) );
INV_X4 _u0_U14275  ( .A(1'b1), .ZN(_u0_ch18_txsz[21] ) );
INV_X4 _u0_U14273  ( .A(1'b1), .ZN(_u0_ch18_txsz[20] ) );
INV_X4 _u0_U14271  ( .A(1'b1), .ZN(_u0_ch18_txsz[19] ) );
INV_X4 _u0_U14269  ( .A(1'b1), .ZN(_u0_ch18_txsz[18] ) );
INV_X4 _u0_U14267  ( .A(1'b1), .ZN(_u0_ch18_txsz[17] ) );
INV_X4 _u0_U14265  ( .A(1'b1), .ZN(_u0_ch18_txsz[16] ) );
INV_X4 _u0_U14263  ( .A(1'b1), .ZN(_u0_ch18_txsz[15] ) );
INV_X4 _u0_U14261  ( .A(1'b1), .ZN(_u0_ch18_txsz[14] ) );
INV_X4 _u0_U14259  ( .A(1'b1), .ZN(_u0_ch18_txsz[13] ) );
INV_X4 _u0_U14257  ( .A(1'b1), .ZN(_u0_ch18_txsz[12] ) );
INV_X4 _u0_U14255  ( .A(1'b1), .ZN(_u0_ch18_txsz[11] ) );
INV_X4 _u0_U14253  ( .A(1'b1), .ZN(_u0_ch18_txsz[10] ) );
INV_X4 _u0_U14251  ( .A(1'b1), .ZN(_u0_ch18_txsz[9] ) );
INV_X4 _u0_U14249  ( .A(1'b1), .ZN(_u0_ch18_txsz[8] ) );
INV_X4 _u0_U14247  ( .A(1'b1), .ZN(_u0_ch18_txsz[7] ) );
INV_X4 _u0_U14245  ( .A(1'b1), .ZN(_u0_ch18_txsz[6] ) );
INV_X4 _u0_U14243  ( .A(1'b1), .ZN(_u0_ch18_txsz[5] ) );
INV_X4 _u0_U14241  ( .A(1'b1), .ZN(_u0_ch18_txsz[4] ) );
INV_X4 _u0_U14239  ( .A(1'b1), .ZN(_u0_ch18_txsz[3] ) );
INV_X4 _u0_U14237  ( .A(1'b1), .ZN(_u0_ch18_txsz[2] ) );
INV_X4 _u0_U14235  ( .A(1'b1), .ZN(_u0_ch18_txsz[1] ) );
INV_X4 _u0_U14233  ( .A(1'b1), .ZN(_u0_ch18_txsz[0] ) );
INV_X4 _u0_U14231  ( .A(1'b1), .ZN(_u0_ch18_adr0[31] ) );
INV_X4 _u0_U14229  ( .A(1'b1), .ZN(_u0_ch18_adr0[30] ) );
INV_X4 _u0_U14227  ( .A(1'b1), .ZN(_u0_ch18_adr0[29] ) );
INV_X4 _u0_U14225  ( .A(1'b1), .ZN(_u0_ch18_adr0[28] ) );
INV_X4 _u0_U14223  ( .A(1'b1), .ZN(_u0_ch18_adr0[27] ) );
INV_X4 _u0_U14221  ( .A(1'b1), .ZN(_u0_ch18_adr0[26] ) );
INV_X4 _u0_U14219  ( .A(1'b1), .ZN(_u0_ch18_adr0[25] ) );
INV_X4 _u0_U14217  ( .A(1'b1), .ZN(_u0_ch18_adr0[24] ) );
INV_X4 _u0_U14215  ( .A(1'b1), .ZN(_u0_ch18_adr0[23] ) );
INV_X4 _u0_U14213  ( .A(1'b1), .ZN(_u0_ch18_adr0[22] ) );
INV_X4 _u0_U14211  ( .A(1'b1), .ZN(_u0_ch18_adr0[21] ) );
INV_X4 _u0_U14209  ( .A(1'b1), .ZN(_u0_ch18_adr0[20] ) );
INV_X4 _u0_U14207  ( .A(1'b1), .ZN(_u0_ch18_adr0[19] ) );
INV_X4 _u0_U14205  ( .A(1'b1), .ZN(_u0_ch18_adr0[18] ) );
INV_X4 _u0_U14203  ( .A(1'b1), .ZN(_u0_ch18_adr0[17] ) );
INV_X4 _u0_U14201  ( .A(1'b1), .ZN(_u0_ch18_adr0[16] ) );
INV_X4 _u0_U14199  ( .A(1'b1), .ZN(_u0_ch18_adr0[15] ) );
INV_X4 _u0_U14197  ( .A(1'b1), .ZN(_u0_ch18_adr0[14] ) );
INV_X4 _u0_U14195  ( .A(1'b1), .ZN(_u0_ch18_adr0[13] ) );
INV_X4 _u0_U14193  ( .A(1'b1), .ZN(_u0_ch18_adr0[12] ) );
INV_X4 _u0_U14191  ( .A(1'b1), .ZN(_u0_ch18_adr0[11] ) );
INV_X4 _u0_U14189  ( .A(1'b1), .ZN(_u0_ch18_adr0[10] ) );
INV_X4 _u0_U14187  ( .A(1'b1), .ZN(_u0_ch18_adr0[9] ) );
INV_X4 _u0_U14185  ( .A(1'b1), .ZN(_u0_ch18_adr0[8] ) );
INV_X4 _u0_U14183  ( .A(1'b1), .ZN(_u0_ch18_adr0[7] ) );
INV_X4 _u0_U14181  ( .A(1'b1), .ZN(_u0_ch18_adr0[6] ) );
INV_X4 _u0_U14179  ( .A(1'b1), .ZN(_u0_ch18_adr0[5] ) );
INV_X4 _u0_U14177  ( .A(1'b1), .ZN(_u0_ch18_adr0[4] ) );
INV_X4 _u0_U14175  ( .A(1'b1), .ZN(_u0_ch18_adr0[3] ) );
INV_X4 _u0_U14173  ( .A(1'b1), .ZN(_u0_ch18_adr0[2] ) );
INV_X4 _u0_U14171  ( .A(1'b1), .ZN(_u0_ch18_adr0[1] ) );
INV_X4 _u0_U14169  ( .A(1'b1), .ZN(_u0_ch18_adr0[0] ) );
INV_X4 _u0_U14167  ( .A(1'b1), .ZN(_u0_ch18_adr1[31] ) );
INV_X4 _u0_U14165  ( .A(1'b1), .ZN(_u0_ch18_adr1[30] ) );
INV_X4 _u0_U14163  ( .A(1'b1), .ZN(_u0_ch18_adr1[29] ) );
INV_X4 _u0_U14161  ( .A(1'b1), .ZN(_u0_ch18_adr1[28] ) );
INV_X4 _u0_U14159  ( .A(1'b1), .ZN(_u0_ch18_adr1[27] ) );
INV_X4 _u0_U14157  ( .A(1'b1), .ZN(_u0_ch18_adr1[26] ) );
INV_X4 _u0_U14155  ( .A(1'b1), .ZN(_u0_ch18_adr1[25] ) );
INV_X4 _u0_U14153  ( .A(1'b1), .ZN(_u0_ch18_adr1[24] ) );
INV_X4 _u0_U14151  ( .A(1'b1), .ZN(_u0_ch18_adr1[23] ) );
INV_X4 _u0_U14149  ( .A(1'b1), .ZN(_u0_ch18_adr1[22] ) );
INV_X4 _u0_U14147  ( .A(1'b1), .ZN(_u0_ch18_adr1[21] ) );
INV_X4 _u0_U14145  ( .A(1'b1), .ZN(_u0_ch18_adr1[20] ) );
INV_X4 _u0_U14143  ( .A(1'b1), .ZN(_u0_ch18_adr1[19] ) );
INV_X4 _u0_U14141  ( .A(1'b1), .ZN(_u0_ch18_adr1[18] ) );
INV_X4 _u0_U14139  ( .A(1'b1), .ZN(_u0_ch18_adr1[17] ) );
INV_X4 _u0_U14137  ( .A(1'b1), .ZN(_u0_ch18_adr1[16] ) );
INV_X4 _u0_U14135  ( .A(1'b1), .ZN(_u0_ch18_adr1[15] ) );
INV_X4 _u0_U14133  ( .A(1'b1), .ZN(_u0_ch18_adr1[14] ) );
INV_X4 _u0_U14131  ( .A(1'b1), .ZN(_u0_ch18_adr1[13] ) );
INV_X4 _u0_U14129  ( .A(1'b1), .ZN(_u0_ch18_adr1[12] ) );
INV_X4 _u0_U14127  ( .A(1'b1), .ZN(_u0_ch18_adr1[11] ) );
INV_X4 _u0_U14125  ( .A(1'b1), .ZN(_u0_ch18_adr1[10] ) );
INV_X4 _u0_U14123  ( .A(1'b1), .ZN(_u0_ch18_adr1[9] ) );
INV_X4 _u0_U14121  ( .A(1'b1), .ZN(_u0_ch18_adr1[8] ) );
INV_X4 _u0_U14119  ( .A(1'b1), .ZN(_u0_ch18_adr1[7] ) );
INV_X4 _u0_U14117  ( .A(1'b1), .ZN(_u0_ch18_adr1[6] ) );
INV_X4 _u0_U14115  ( .A(1'b1), .ZN(_u0_ch18_adr1[5] ) );
INV_X4 _u0_U14113  ( .A(1'b1), .ZN(_u0_ch18_adr1[4] ) );
INV_X4 _u0_U14111  ( .A(1'b1), .ZN(_u0_ch18_adr1[3] ) );
INV_X4 _u0_U14109  ( .A(1'b1), .ZN(_u0_ch18_adr1[2] ) );
INV_X4 _u0_U14107  ( .A(1'b1), .ZN(_u0_ch18_adr1[1] ) );
INV_X4 _u0_U14105  ( .A(1'b1), .ZN(_u0_ch18_adr1[0] ) );
INV_X4 _u0_U14103  ( .A(1'b0), .ZN(_u0_ch18_am0[31] ) );
INV_X4 _u0_U14101  ( .A(1'b0), .ZN(_u0_ch18_am0[30] ) );
INV_X4 _u0_U14099  ( .A(1'b0), .ZN(_u0_ch18_am0[29] ) );
INV_X4 _u0_U14097  ( .A(1'b0), .ZN(_u0_ch18_am0[28] ) );
INV_X4 _u0_U14095  ( .A(1'b0), .ZN(_u0_ch18_am0[27] ) );
INV_X4 _u0_U14093  ( .A(1'b0), .ZN(_u0_ch18_am0[26] ) );
INV_X4 _u0_U14091  ( .A(1'b0), .ZN(_u0_ch18_am0[25] ) );
INV_X4 _u0_U14089  ( .A(1'b0), .ZN(_u0_ch18_am0[24] ) );
INV_X4 _u0_U14087  ( .A(1'b0), .ZN(_u0_ch18_am0[23] ) );
INV_X4 _u0_U14085  ( .A(1'b0), .ZN(_u0_ch18_am0[22] ) );
INV_X4 _u0_U14083  ( .A(1'b0), .ZN(_u0_ch18_am0[21] ) );
INV_X4 _u0_U14081  ( .A(1'b0), .ZN(_u0_ch18_am0[20] ) );
INV_X4 _u0_U14079  ( .A(1'b0), .ZN(_u0_ch18_am0[19] ) );
INV_X4 _u0_U14077  ( .A(1'b0), .ZN(_u0_ch18_am0[18] ) );
INV_X4 _u0_U14075  ( .A(1'b0), .ZN(_u0_ch18_am0[17] ) );
INV_X4 _u0_U14073  ( .A(1'b0), .ZN(_u0_ch18_am0[16] ) );
INV_X4 _u0_U14071  ( .A(1'b0), .ZN(_u0_ch18_am0[15] ) );
INV_X4 _u0_U14069  ( .A(1'b0), .ZN(_u0_ch18_am0[14] ) );
INV_X4 _u0_U14067  ( .A(1'b0), .ZN(_u0_ch18_am0[13] ) );
INV_X4 _u0_U14065  ( .A(1'b0), .ZN(_u0_ch18_am0[12] ) );
INV_X4 _u0_U14063  ( .A(1'b0), .ZN(_u0_ch18_am0[11] ) );
INV_X4 _u0_U14061  ( .A(1'b0), .ZN(_u0_ch18_am0[10] ) );
INV_X4 _u0_U14059  ( .A(1'b0), .ZN(_u0_ch18_am0[9] ) );
INV_X4 _u0_U14057  ( .A(1'b0), .ZN(_u0_ch18_am0[8] ) );
INV_X4 _u0_U14055  ( .A(1'b0), .ZN(_u0_ch18_am0[7] ) );
INV_X4 _u0_U14053  ( .A(1'b0), .ZN(_u0_ch18_am0[6] ) );
INV_X4 _u0_U14051  ( .A(1'b0), .ZN(_u0_ch18_am0[5] ) );
INV_X4 _u0_U14049  ( .A(1'b0), .ZN(_u0_ch18_am0[4] ) );
INV_X4 _u0_U14047  ( .A(1'b1), .ZN(_u0_ch18_am0[3] ) );
INV_X4 _u0_U14045  ( .A(1'b1), .ZN(_u0_ch18_am0[2] ) );
INV_X4 _u0_U14043  ( .A(1'b1), .ZN(_u0_ch18_am0[1] ) );
INV_X4 _u0_U14041  ( .A(1'b1), .ZN(_u0_ch18_am0[0] ) );
INV_X4 _u0_U14039  ( .A(1'b0), .ZN(_u0_ch18_am1[31] ) );
INV_X4 _u0_U14037  ( .A(1'b0), .ZN(_u0_ch18_am1[30] ) );
INV_X4 _u0_U14035  ( .A(1'b0), .ZN(_u0_ch18_am1[29] ) );
INV_X4 _u0_U14033  ( .A(1'b0), .ZN(_u0_ch18_am1[28] ) );
INV_X4 _u0_U14031  ( .A(1'b0), .ZN(_u0_ch18_am1[27] ) );
INV_X4 _u0_U14029  ( .A(1'b0), .ZN(_u0_ch18_am1[26] ) );
INV_X4 _u0_U14027  ( .A(1'b0), .ZN(_u0_ch18_am1[25] ) );
INV_X4 _u0_U14025  ( .A(1'b0), .ZN(_u0_ch18_am1[24] ) );
INV_X4 _u0_U14023  ( .A(1'b0), .ZN(_u0_ch18_am1[23] ) );
INV_X4 _u0_U14021  ( .A(1'b0), .ZN(_u0_ch18_am1[22] ) );
INV_X4 _u0_U14019  ( .A(1'b0), .ZN(_u0_ch18_am1[21] ) );
INV_X4 _u0_U14017  ( .A(1'b0), .ZN(_u0_ch18_am1[20] ) );
INV_X4 _u0_U14015  ( .A(1'b0), .ZN(_u0_ch18_am1[19] ) );
INV_X4 _u0_U14013  ( .A(1'b0), .ZN(_u0_ch18_am1[18] ) );
INV_X4 _u0_U14011  ( .A(1'b0), .ZN(_u0_ch18_am1[17] ) );
INV_X4 _u0_U14009  ( .A(1'b0), .ZN(_u0_ch18_am1[16] ) );
INV_X4 _u0_U14007  ( .A(1'b0), .ZN(_u0_ch18_am1[15] ) );
INV_X4 _u0_U14005  ( .A(1'b0), .ZN(_u0_ch18_am1[14] ) );
INV_X4 _u0_U14003  ( .A(1'b0), .ZN(_u0_ch18_am1[13] ) );
INV_X4 _u0_U14001  ( .A(1'b0), .ZN(_u0_ch18_am1[12] ) );
INV_X4 _u0_U13999  ( .A(1'b0), .ZN(_u0_ch18_am1[11] ) );
INV_X4 _u0_U13997  ( .A(1'b0), .ZN(_u0_ch18_am1[10] ) );
INV_X4 _u0_U13995  ( .A(1'b0), .ZN(_u0_ch18_am1[9] ) );
INV_X4 _u0_U13993  ( .A(1'b0), .ZN(_u0_ch18_am1[8] ) );
INV_X4 _u0_U13991  ( .A(1'b0), .ZN(_u0_ch18_am1[7] ) );
INV_X4 _u0_U13989  ( .A(1'b0), .ZN(_u0_ch18_am1[6] ) );
INV_X4 _u0_U13987  ( .A(1'b0), .ZN(_u0_ch18_am1[5] ) );
INV_X4 _u0_U13985  ( .A(1'b0), .ZN(_u0_ch18_am1[4] ) );
INV_X4 _u0_U13983  ( .A(1'b1), .ZN(_u0_ch18_am1[3] ) );
INV_X4 _u0_U13981  ( .A(1'b1), .ZN(_u0_ch18_am1[2] ) );
INV_X4 _u0_U13979  ( .A(1'b1), .ZN(_u0_ch18_am1[1] ) );
INV_X4 _u0_U13977  ( .A(1'b1), .ZN(_u0_ch18_am1[0] ) );
INV_X4 _u0_U13975  ( .A(1'b1), .ZN(_u0_pointer19[31] ) );
INV_X4 _u0_U13973  ( .A(1'b1), .ZN(_u0_pointer19[30] ) );
INV_X4 _u0_U13971  ( .A(1'b1), .ZN(_u0_pointer19[29] ) );
INV_X4 _u0_U13969  ( .A(1'b1), .ZN(_u0_pointer19[28] ) );
INV_X4 _u0_U13967  ( .A(1'b1), .ZN(_u0_pointer19[27] ) );
INV_X4 _u0_U13965  ( .A(1'b1), .ZN(_u0_pointer19[26] ) );
INV_X4 _u0_U13963  ( .A(1'b1), .ZN(_u0_pointer19[25] ) );
INV_X4 _u0_U13961  ( .A(1'b1), .ZN(_u0_pointer19[24] ) );
INV_X4 _u0_U13959  ( .A(1'b1), .ZN(_u0_pointer19[23] ) );
INV_X4 _u0_U13957  ( .A(1'b1), .ZN(_u0_pointer19[22] ) );
INV_X4 _u0_U13955  ( .A(1'b1), .ZN(_u0_pointer19[21] ) );
INV_X4 _u0_U13953  ( .A(1'b1), .ZN(_u0_pointer19[20] ) );
INV_X4 _u0_U13951  ( .A(1'b1), .ZN(_u0_pointer19[19] ) );
INV_X4 _u0_U13949  ( .A(1'b1), .ZN(_u0_pointer19[18] ) );
INV_X4 _u0_U13947  ( .A(1'b1), .ZN(_u0_pointer19[17] ) );
INV_X4 _u0_U13945  ( .A(1'b1), .ZN(_u0_pointer19[16] ) );
INV_X4 _u0_U13943  ( .A(1'b1), .ZN(_u0_pointer19[15] ) );
INV_X4 _u0_U13941  ( .A(1'b1), .ZN(_u0_pointer19[14] ) );
INV_X4 _u0_U13939  ( .A(1'b1), .ZN(_u0_pointer19[13] ) );
INV_X4 _u0_U13937  ( .A(1'b1), .ZN(_u0_pointer19[12] ) );
INV_X4 _u0_U13935  ( .A(1'b1), .ZN(_u0_pointer19[11] ) );
INV_X4 _u0_U13933  ( .A(1'b1), .ZN(_u0_pointer19[10] ) );
INV_X4 _u0_U13931  ( .A(1'b1), .ZN(_u0_pointer19[9] ) );
INV_X4 _u0_U13929  ( .A(1'b1), .ZN(_u0_pointer19[8] ) );
INV_X4 _u0_U13927  ( .A(1'b1), .ZN(_u0_pointer19[7] ) );
INV_X4 _u0_U13925  ( .A(1'b1), .ZN(_u0_pointer19[6] ) );
INV_X4 _u0_U13923  ( .A(1'b1), .ZN(_u0_pointer19[5] ) );
INV_X4 _u0_U13921  ( .A(1'b1), .ZN(_u0_pointer19[4] ) );
INV_X4 _u0_U13919  ( .A(1'b1), .ZN(_u0_pointer19[3] ) );
INV_X4 _u0_U13917  ( .A(1'b1), .ZN(_u0_pointer19[2] ) );
INV_X4 _u0_U13915  ( .A(1'b1), .ZN(_u0_pointer19[1] ) );
INV_X4 _u0_U13913  ( .A(1'b1), .ZN(_u0_pointer19[0] ) );
INV_X4 _u0_U13911  ( .A(1'b1), .ZN(_u0_pointer19_s[31] ) );
INV_X4 _u0_U13909  ( .A(1'b1), .ZN(_u0_pointer19_s[30] ) );
INV_X4 _u0_U13907  ( .A(1'b1), .ZN(_u0_pointer19_s[29] ) );
INV_X4 _u0_U13905  ( .A(1'b1), .ZN(_u0_pointer19_s[28] ) );
INV_X4 _u0_U13903  ( .A(1'b1), .ZN(_u0_pointer19_s[27] ) );
INV_X4 _u0_U13901  ( .A(1'b1), .ZN(_u0_pointer19_s[26] ) );
INV_X4 _u0_U13899  ( .A(1'b1), .ZN(_u0_pointer19_s[25] ) );
INV_X4 _u0_U13897  ( .A(1'b1), .ZN(_u0_pointer19_s[24] ) );
INV_X4 _u0_U13895  ( .A(1'b1), .ZN(_u0_pointer19_s[23] ) );
INV_X4 _u0_U13893  ( .A(1'b1), .ZN(_u0_pointer19_s[22] ) );
INV_X4 _u0_U13891  ( .A(1'b1), .ZN(_u0_pointer19_s[21] ) );
INV_X4 _u0_U13889  ( .A(1'b1), .ZN(_u0_pointer19_s[20] ) );
INV_X4 _u0_U13887  ( .A(1'b1), .ZN(_u0_pointer19_s[19] ) );
INV_X4 _u0_U13885  ( .A(1'b1), .ZN(_u0_pointer19_s[18] ) );
INV_X4 _u0_U13883  ( .A(1'b1), .ZN(_u0_pointer19_s[17] ) );
INV_X4 _u0_U13881  ( .A(1'b1), .ZN(_u0_pointer19_s[16] ) );
INV_X4 _u0_U13879  ( .A(1'b1), .ZN(_u0_pointer19_s[15] ) );
INV_X4 _u0_U13877  ( .A(1'b1), .ZN(_u0_pointer19_s[14] ) );
INV_X4 _u0_U13875  ( .A(1'b1), .ZN(_u0_pointer19_s[13] ) );
INV_X4 _u0_U13873  ( .A(1'b1), .ZN(_u0_pointer19_s[12] ) );
INV_X4 _u0_U13871  ( .A(1'b1), .ZN(_u0_pointer19_s[11] ) );
INV_X4 _u0_U13869  ( .A(1'b1), .ZN(_u0_pointer19_s[10] ) );
INV_X4 _u0_U13867  ( .A(1'b1), .ZN(_u0_pointer19_s[9] ) );
INV_X4 _u0_U13865  ( .A(1'b1), .ZN(_u0_pointer19_s[8] ) );
INV_X4 _u0_U13863  ( .A(1'b1), .ZN(_u0_pointer19_s[7] ) );
INV_X4 _u0_U13861  ( .A(1'b1), .ZN(_u0_pointer19_s[6] ) );
INV_X4 _u0_U13859  ( .A(1'b1), .ZN(_u0_pointer19_s[5] ) );
INV_X4 _u0_U13857  ( .A(1'b1), .ZN(_u0_pointer19_s[4] ) );
INV_X4 _u0_U13855  ( .A(1'b1), .ZN(_u0_pointer19_s[3] ) );
INV_X4 _u0_U13853  ( .A(1'b1), .ZN(_u0_pointer19_s[2] ) );
INV_X4 _u0_U13851  ( .A(1'b1), .ZN(_u0_pointer19_s[1] ) );
INV_X4 _u0_U13849  ( .A(1'b1), .ZN(_u0_pointer19_s[0] ) );
INV_X4 _u0_U13847  ( .A(1'b1), .ZN(_u0_ch19_csr[31] ) );
INV_X4 _u0_U13845  ( .A(1'b1), .ZN(_u0_ch19_csr[30] ) );
INV_X4 _u0_U13843  ( .A(1'b1), .ZN(_u0_ch19_csr[29] ) );
INV_X4 _u0_U13841  ( .A(1'b1), .ZN(_u0_ch19_csr[28] ) );
INV_X4 _u0_U13839  ( .A(1'b1), .ZN(_u0_ch19_csr[27] ) );
INV_X4 _u0_U13837  ( .A(1'b1), .ZN(_u0_ch19_csr[26] ) );
INV_X4 _u0_U13835  ( .A(1'b1), .ZN(_u0_ch19_csr[25] ) );
INV_X4 _u0_U13833  ( .A(1'b1), .ZN(_u0_ch19_csr[24] ) );
INV_X4 _u0_U13831  ( .A(1'b1), .ZN(_u0_ch19_csr[23] ) );
INV_X4 _u0_U13829  ( .A(1'b1), .ZN(_u0_ch19_csr[22] ) );
INV_X4 _u0_U13827  ( .A(1'b1), .ZN(_u0_ch19_csr[21] ) );
INV_X4 _u0_U13825  ( .A(1'b1), .ZN(_u0_ch19_csr[20] ) );
INV_X4 _u0_U13823  ( .A(1'b1), .ZN(_u0_ch19_csr[19] ) );
INV_X4 _u0_U13821  ( .A(1'b1), .ZN(_u0_ch19_csr[18] ) );
INV_X4 _u0_U13819  ( .A(1'b1), .ZN(_u0_ch19_csr[17] ) );
INV_X4 _u0_U13817  ( .A(1'b1), .ZN(_u0_ch19_csr[16] ) );
INV_X4 _u0_U13815  ( .A(1'b1), .ZN(_u0_ch19_csr[15] ) );
INV_X4 _u0_U13813  ( .A(1'b1), .ZN(_u0_ch19_csr[14] ) );
INV_X4 _u0_U13811  ( .A(1'b1), .ZN(_u0_ch19_csr[13] ) );
INV_X4 _u0_U13809  ( .A(1'b1), .ZN(_u0_ch19_csr[12] ) );
INV_X4 _u0_U13807  ( .A(1'b1), .ZN(_u0_ch19_csr[11] ) );
INV_X4 _u0_U13805  ( .A(1'b1), .ZN(_u0_ch19_csr[10] ) );
INV_X4 _u0_U13803  ( .A(1'b1), .ZN(_u0_ch19_csr[9] ) );
INV_X4 _u0_U13801  ( .A(1'b1), .ZN(_u0_ch19_csr[8] ) );
INV_X4 _u0_U13799  ( .A(1'b1), .ZN(_u0_ch19_csr[7] ) );
INV_X4 _u0_U13797  ( .A(1'b1), .ZN(_u0_ch19_csr[6] ) );
INV_X4 _u0_U13795  ( .A(1'b1), .ZN(_u0_ch19_csr[5] ) );
INV_X4 _u0_U13793  ( .A(1'b1), .ZN(_u0_ch19_csr[4] ) );
INV_X4 _u0_U13791  ( .A(1'b1), .ZN(_u0_ch19_csr[3] ) );
INV_X4 _u0_U13789  ( .A(1'b1), .ZN(_u0_ch19_csr[2] ) );
INV_X4 _u0_U13787  ( .A(1'b1), .ZN(_u0_ch19_csr[1] ) );
INV_X4 _u0_U13785  ( .A(1'b1), .ZN(_u0_ch19_csr[0] ) );
INV_X4 _u0_U13783  ( .A(1'b1), .ZN(_u0_ch19_txsz[31] ) );
INV_X4 _u0_U13781  ( .A(1'b1), .ZN(_u0_ch19_txsz[30] ) );
INV_X4 _u0_U13779  ( .A(1'b1), .ZN(_u0_ch19_txsz[29] ) );
INV_X4 _u0_U13777  ( .A(1'b1), .ZN(_u0_ch19_txsz[28] ) );
INV_X4 _u0_U13775  ( .A(1'b1), .ZN(_u0_ch19_txsz[27] ) );
INV_X4 _u0_U13773  ( .A(1'b1), .ZN(_u0_ch19_txsz[26] ) );
INV_X4 _u0_U13771  ( .A(1'b1), .ZN(_u0_ch19_txsz[25] ) );
INV_X4 _u0_U13769  ( .A(1'b1), .ZN(_u0_ch19_txsz[24] ) );
INV_X4 _u0_U13767  ( .A(1'b1), .ZN(_u0_ch19_txsz[23] ) );
INV_X4 _u0_U13765  ( .A(1'b1), .ZN(_u0_ch19_txsz[22] ) );
INV_X4 _u0_U13763  ( .A(1'b1), .ZN(_u0_ch19_txsz[21] ) );
INV_X4 _u0_U13761  ( .A(1'b1), .ZN(_u0_ch19_txsz[20] ) );
INV_X4 _u0_U13759  ( .A(1'b1), .ZN(_u0_ch19_txsz[19] ) );
INV_X4 _u0_U13757  ( .A(1'b1), .ZN(_u0_ch19_txsz[18] ) );
INV_X4 _u0_U13755  ( .A(1'b1), .ZN(_u0_ch19_txsz[17] ) );
INV_X4 _u0_U13753  ( .A(1'b1), .ZN(_u0_ch19_txsz[16] ) );
INV_X4 _u0_U13751  ( .A(1'b1), .ZN(_u0_ch19_txsz[15] ) );
INV_X4 _u0_U13749  ( .A(1'b1), .ZN(_u0_ch19_txsz[14] ) );
INV_X4 _u0_U13747  ( .A(1'b1), .ZN(_u0_ch19_txsz[13] ) );
INV_X4 _u0_U13745  ( .A(1'b1), .ZN(_u0_ch19_txsz[12] ) );
INV_X4 _u0_U13743  ( .A(1'b1), .ZN(_u0_ch19_txsz[11] ) );
INV_X4 _u0_U13741  ( .A(1'b1), .ZN(_u0_ch19_txsz[10] ) );
INV_X4 _u0_U13739  ( .A(1'b1), .ZN(_u0_ch19_txsz[9] ) );
INV_X4 _u0_U13737  ( .A(1'b1), .ZN(_u0_ch19_txsz[8] ) );
INV_X4 _u0_U13735  ( .A(1'b1), .ZN(_u0_ch19_txsz[7] ) );
INV_X4 _u0_U13733  ( .A(1'b1), .ZN(_u0_ch19_txsz[6] ) );
INV_X4 _u0_U13731  ( .A(1'b1), .ZN(_u0_ch19_txsz[5] ) );
INV_X4 _u0_U13729  ( .A(1'b1), .ZN(_u0_ch19_txsz[4] ) );
INV_X4 _u0_U13727  ( .A(1'b1), .ZN(_u0_ch19_txsz[3] ) );
INV_X4 _u0_U13725  ( .A(1'b1), .ZN(_u0_ch19_txsz[2] ) );
INV_X4 _u0_U13723  ( .A(1'b1), .ZN(_u0_ch19_txsz[1] ) );
INV_X4 _u0_U13721  ( .A(1'b1), .ZN(_u0_ch19_txsz[0] ) );
INV_X4 _u0_U13719  ( .A(1'b1), .ZN(_u0_ch19_adr0[31] ) );
INV_X4 _u0_U13717  ( .A(1'b1), .ZN(_u0_ch19_adr0[30] ) );
INV_X4 _u0_U13715  ( .A(1'b1), .ZN(_u0_ch19_adr0[29] ) );
INV_X4 _u0_U13713  ( .A(1'b1), .ZN(_u0_ch19_adr0[28] ) );
INV_X4 _u0_U13711  ( .A(1'b1), .ZN(_u0_ch19_adr0[27] ) );
INV_X4 _u0_U13709  ( .A(1'b1), .ZN(_u0_ch19_adr0[26] ) );
INV_X4 _u0_U13707  ( .A(1'b1), .ZN(_u0_ch19_adr0[25] ) );
INV_X4 _u0_U13705  ( .A(1'b1), .ZN(_u0_ch19_adr0[24] ) );
INV_X4 _u0_U13703  ( .A(1'b1), .ZN(_u0_ch19_adr0[23] ) );
INV_X4 _u0_U13701  ( .A(1'b1), .ZN(_u0_ch19_adr0[22] ) );
INV_X4 _u0_U13699  ( .A(1'b1), .ZN(_u0_ch19_adr0[21] ) );
INV_X4 _u0_U13697  ( .A(1'b1), .ZN(_u0_ch19_adr0[20] ) );
INV_X4 _u0_U13695  ( .A(1'b1), .ZN(_u0_ch19_adr0[19] ) );
INV_X4 _u0_U13693  ( .A(1'b1), .ZN(_u0_ch19_adr0[18] ) );
INV_X4 _u0_U13691  ( .A(1'b1), .ZN(_u0_ch19_adr0[17] ) );
INV_X4 _u0_U13689  ( .A(1'b1), .ZN(_u0_ch19_adr0[16] ) );
INV_X4 _u0_U13687  ( .A(1'b1), .ZN(_u0_ch19_adr0[15] ) );
INV_X4 _u0_U13685  ( .A(1'b1), .ZN(_u0_ch19_adr0[14] ) );
INV_X4 _u0_U13683  ( .A(1'b1), .ZN(_u0_ch19_adr0[13] ) );
INV_X4 _u0_U13681  ( .A(1'b1), .ZN(_u0_ch19_adr0[12] ) );
INV_X4 _u0_U13679  ( .A(1'b1), .ZN(_u0_ch19_adr0[11] ) );
INV_X4 _u0_U13677  ( .A(1'b1), .ZN(_u0_ch19_adr0[10] ) );
INV_X4 _u0_U13675  ( .A(1'b1), .ZN(_u0_ch19_adr0[9] ) );
INV_X4 _u0_U13673  ( .A(1'b1), .ZN(_u0_ch19_adr0[8] ) );
INV_X4 _u0_U13671  ( .A(1'b1), .ZN(_u0_ch19_adr0[7] ) );
INV_X4 _u0_U13669  ( .A(1'b1), .ZN(_u0_ch19_adr0[6] ) );
INV_X4 _u0_U13667  ( .A(1'b1), .ZN(_u0_ch19_adr0[5] ) );
INV_X4 _u0_U13665  ( .A(1'b1), .ZN(_u0_ch19_adr0[4] ) );
INV_X4 _u0_U13663  ( .A(1'b1), .ZN(_u0_ch19_adr0[3] ) );
INV_X4 _u0_U13661  ( .A(1'b1), .ZN(_u0_ch19_adr0[2] ) );
INV_X4 _u0_U13659  ( .A(1'b1), .ZN(_u0_ch19_adr0[1] ) );
INV_X4 _u0_U13657  ( .A(1'b1), .ZN(_u0_ch19_adr0[0] ) );
INV_X4 _u0_U13655  ( .A(1'b1), .ZN(_u0_ch19_adr1[31] ) );
INV_X4 _u0_U13653  ( .A(1'b1), .ZN(_u0_ch19_adr1[30] ) );
INV_X4 _u0_U13651  ( .A(1'b1), .ZN(_u0_ch19_adr1[29] ) );
INV_X4 _u0_U13649  ( .A(1'b1), .ZN(_u0_ch19_adr1[28] ) );
INV_X4 _u0_U13647  ( .A(1'b1), .ZN(_u0_ch19_adr1[27] ) );
INV_X4 _u0_U13645  ( .A(1'b1), .ZN(_u0_ch19_adr1[26] ) );
INV_X4 _u0_U13643  ( .A(1'b1), .ZN(_u0_ch19_adr1[25] ) );
INV_X4 _u0_U13641  ( .A(1'b1), .ZN(_u0_ch19_adr1[24] ) );
INV_X4 _u0_U13639  ( .A(1'b1), .ZN(_u0_ch19_adr1[23] ) );
INV_X4 _u0_U13637  ( .A(1'b1), .ZN(_u0_ch19_adr1[22] ) );
INV_X4 _u0_U13635  ( .A(1'b1), .ZN(_u0_ch19_adr1[21] ) );
INV_X4 _u0_U13633  ( .A(1'b1), .ZN(_u0_ch19_adr1[20] ) );
INV_X4 _u0_U13631  ( .A(1'b1), .ZN(_u0_ch19_adr1[19] ) );
INV_X4 _u0_U13629  ( .A(1'b1), .ZN(_u0_ch19_adr1[18] ) );
INV_X4 _u0_U13627  ( .A(1'b1), .ZN(_u0_ch19_adr1[17] ) );
INV_X4 _u0_U13625  ( .A(1'b1), .ZN(_u0_ch19_adr1[16] ) );
INV_X4 _u0_U13623  ( .A(1'b1), .ZN(_u0_ch19_adr1[15] ) );
INV_X4 _u0_U13621  ( .A(1'b1), .ZN(_u0_ch19_adr1[14] ) );
INV_X4 _u0_U13619  ( .A(1'b1), .ZN(_u0_ch19_adr1[13] ) );
INV_X4 _u0_U13617  ( .A(1'b1), .ZN(_u0_ch19_adr1[12] ) );
INV_X4 _u0_U13615  ( .A(1'b1), .ZN(_u0_ch19_adr1[11] ) );
INV_X4 _u0_U13613  ( .A(1'b1), .ZN(_u0_ch19_adr1[10] ) );
INV_X4 _u0_U13611  ( .A(1'b1), .ZN(_u0_ch19_adr1[9] ) );
INV_X4 _u0_U13609  ( .A(1'b1), .ZN(_u0_ch19_adr1[8] ) );
INV_X4 _u0_U13607  ( .A(1'b1), .ZN(_u0_ch19_adr1[7] ) );
INV_X4 _u0_U13605  ( .A(1'b1), .ZN(_u0_ch19_adr1[6] ) );
INV_X4 _u0_U13603  ( .A(1'b1), .ZN(_u0_ch19_adr1[5] ) );
INV_X4 _u0_U13601  ( .A(1'b1), .ZN(_u0_ch19_adr1[4] ) );
INV_X4 _u0_U13599  ( .A(1'b1), .ZN(_u0_ch19_adr1[3] ) );
INV_X4 _u0_U13597  ( .A(1'b1), .ZN(_u0_ch19_adr1[2] ) );
INV_X4 _u0_U13595  ( .A(1'b1), .ZN(_u0_ch19_adr1[1] ) );
INV_X4 _u0_U13593  ( .A(1'b1), .ZN(_u0_ch19_adr1[0] ) );
INV_X4 _u0_U13591  ( .A(1'b0), .ZN(_u0_ch19_am0[31] ) );
INV_X4 _u0_U13589  ( .A(1'b0), .ZN(_u0_ch19_am0[30] ) );
INV_X4 _u0_U13587  ( .A(1'b0), .ZN(_u0_ch19_am0[29] ) );
INV_X4 _u0_U13585  ( .A(1'b0), .ZN(_u0_ch19_am0[28] ) );
INV_X4 _u0_U13583  ( .A(1'b0), .ZN(_u0_ch19_am0[27] ) );
INV_X4 _u0_U13581  ( .A(1'b0), .ZN(_u0_ch19_am0[26] ) );
INV_X4 _u0_U13579  ( .A(1'b0), .ZN(_u0_ch19_am0[25] ) );
INV_X4 _u0_U13577  ( .A(1'b0), .ZN(_u0_ch19_am0[24] ) );
INV_X4 _u0_U13575  ( .A(1'b0), .ZN(_u0_ch19_am0[23] ) );
INV_X4 _u0_U13573  ( .A(1'b0), .ZN(_u0_ch19_am0[22] ) );
INV_X4 _u0_U13571  ( .A(1'b0), .ZN(_u0_ch19_am0[21] ) );
INV_X4 _u0_U13569  ( .A(1'b0), .ZN(_u0_ch19_am0[20] ) );
INV_X4 _u0_U13567  ( .A(1'b0), .ZN(_u0_ch19_am0[19] ) );
INV_X4 _u0_U13565  ( .A(1'b0), .ZN(_u0_ch19_am0[18] ) );
INV_X4 _u0_U13563  ( .A(1'b0), .ZN(_u0_ch19_am0[17] ) );
INV_X4 _u0_U13561  ( .A(1'b0), .ZN(_u0_ch19_am0[16] ) );
INV_X4 _u0_U13559  ( .A(1'b0), .ZN(_u0_ch19_am0[15] ) );
INV_X4 _u0_U13557  ( .A(1'b0), .ZN(_u0_ch19_am0[14] ) );
INV_X4 _u0_U13555  ( .A(1'b0), .ZN(_u0_ch19_am0[13] ) );
INV_X4 _u0_U13553  ( .A(1'b0), .ZN(_u0_ch19_am0[12] ) );
INV_X4 _u0_U13551  ( .A(1'b0), .ZN(_u0_ch19_am0[11] ) );
INV_X4 _u0_U13549  ( .A(1'b0), .ZN(_u0_ch19_am0[10] ) );
INV_X4 _u0_U13547  ( .A(1'b0), .ZN(_u0_ch19_am0[9] ) );
INV_X4 _u0_U13545  ( .A(1'b0), .ZN(_u0_ch19_am0[8] ) );
INV_X4 _u0_U13543  ( .A(1'b0), .ZN(_u0_ch19_am0[7] ) );
INV_X4 _u0_U13541  ( .A(1'b0), .ZN(_u0_ch19_am0[6] ) );
INV_X4 _u0_U13539  ( .A(1'b0), .ZN(_u0_ch19_am0[5] ) );
INV_X4 _u0_U13537  ( .A(1'b0), .ZN(_u0_ch19_am0[4] ) );
INV_X4 _u0_U13535  ( .A(1'b1), .ZN(_u0_ch19_am0[3] ) );
INV_X4 _u0_U13533  ( .A(1'b1), .ZN(_u0_ch19_am0[2] ) );
INV_X4 _u0_U13531  ( .A(1'b1), .ZN(_u0_ch19_am0[1] ) );
INV_X4 _u0_U13529  ( .A(1'b1), .ZN(_u0_ch19_am0[0] ) );
INV_X4 _u0_U13527  ( .A(1'b0), .ZN(_u0_ch19_am1[31] ) );
INV_X4 _u0_U13525  ( .A(1'b0), .ZN(_u0_ch19_am1[30] ) );
INV_X4 _u0_U13523  ( .A(1'b0), .ZN(_u0_ch19_am1[29] ) );
INV_X4 _u0_U13521  ( .A(1'b0), .ZN(_u0_ch19_am1[28] ) );
INV_X4 _u0_U13519  ( .A(1'b0), .ZN(_u0_ch19_am1[27] ) );
INV_X4 _u0_U13517  ( .A(1'b0), .ZN(_u0_ch19_am1[26] ) );
INV_X4 _u0_U13515  ( .A(1'b0), .ZN(_u0_ch19_am1[25] ) );
INV_X4 _u0_U13513  ( .A(1'b0), .ZN(_u0_ch19_am1[24] ) );
INV_X4 _u0_U13511  ( .A(1'b0), .ZN(_u0_ch19_am1[23] ) );
INV_X4 _u0_U13509  ( .A(1'b0), .ZN(_u0_ch19_am1[22] ) );
INV_X4 _u0_U13507  ( .A(1'b0), .ZN(_u0_ch19_am1[21] ) );
INV_X4 _u0_U13505  ( .A(1'b0), .ZN(_u0_ch19_am1[20] ) );
INV_X4 _u0_U13503  ( .A(1'b0), .ZN(_u0_ch19_am1[19] ) );
INV_X4 _u0_U13501  ( .A(1'b0), .ZN(_u0_ch19_am1[18] ) );
INV_X4 _u0_U13499  ( .A(1'b0), .ZN(_u0_ch19_am1[17] ) );
INV_X4 _u0_U13497  ( .A(1'b0), .ZN(_u0_ch19_am1[16] ) );
INV_X4 _u0_U13495  ( .A(1'b0), .ZN(_u0_ch19_am1[15] ) );
INV_X4 _u0_U13493  ( .A(1'b0), .ZN(_u0_ch19_am1[14] ) );
INV_X4 _u0_U13491  ( .A(1'b0), .ZN(_u0_ch19_am1[13] ) );
INV_X4 _u0_U13489  ( .A(1'b0), .ZN(_u0_ch19_am1[12] ) );
INV_X4 _u0_U13487  ( .A(1'b0), .ZN(_u0_ch19_am1[11] ) );
INV_X4 _u0_U13485  ( .A(1'b0), .ZN(_u0_ch19_am1[10] ) );
INV_X4 _u0_U13483  ( .A(1'b0), .ZN(_u0_ch19_am1[9] ) );
INV_X4 _u0_U13481  ( .A(1'b0), .ZN(_u0_ch19_am1[8] ) );
INV_X4 _u0_U13479  ( .A(1'b0), .ZN(_u0_ch19_am1[7] ) );
INV_X4 _u0_U13477  ( .A(1'b0), .ZN(_u0_ch19_am1[6] ) );
INV_X4 _u0_U13475  ( .A(1'b0), .ZN(_u0_ch19_am1[5] ) );
INV_X4 _u0_U13473  ( .A(1'b0), .ZN(_u0_ch19_am1[4] ) );
INV_X4 _u0_U13471  ( .A(1'b1), .ZN(_u0_ch19_am1[3] ) );
INV_X4 _u0_U13469  ( .A(1'b1), .ZN(_u0_ch19_am1[2] ) );
INV_X4 _u0_U13467  ( .A(1'b1), .ZN(_u0_ch19_am1[1] ) );
INV_X4 _u0_U13465  ( .A(1'b1), .ZN(_u0_ch19_am1[0] ) );
INV_X4 _u0_U13463  ( .A(1'b1), .ZN(_u0_pointer20[31] ) );
INV_X4 _u0_U13461  ( .A(1'b1), .ZN(_u0_pointer20[30] ) );
INV_X4 _u0_U13459  ( .A(1'b1), .ZN(_u0_pointer20[29] ) );
INV_X4 _u0_U13457  ( .A(1'b1), .ZN(_u0_pointer20[28] ) );
INV_X4 _u0_U13455  ( .A(1'b1), .ZN(_u0_pointer20[27] ) );
INV_X4 _u0_U13453  ( .A(1'b1), .ZN(_u0_pointer20[26] ) );
INV_X4 _u0_U13451  ( .A(1'b1), .ZN(_u0_pointer20[25] ) );
INV_X4 _u0_U13449  ( .A(1'b1), .ZN(_u0_pointer20[24] ) );
INV_X4 _u0_U13447  ( .A(1'b1), .ZN(_u0_pointer20[23] ) );
INV_X4 _u0_U13445  ( .A(1'b1), .ZN(_u0_pointer20[22] ) );
INV_X4 _u0_U13443  ( .A(1'b1), .ZN(_u0_pointer20[21] ) );
INV_X4 _u0_U13441  ( .A(1'b1), .ZN(_u0_pointer20[20] ) );
INV_X4 _u0_U13439  ( .A(1'b1), .ZN(_u0_pointer20[19] ) );
INV_X4 _u0_U13437  ( .A(1'b1), .ZN(_u0_pointer20[18] ) );
INV_X4 _u0_U13435  ( .A(1'b1), .ZN(_u0_pointer20[17] ) );
INV_X4 _u0_U13433  ( .A(1'b1), .ZN(_u0_pointer20[16] ) );
INV_X4 _u0_U13431  ( .A(1'b1), .ZN(_u0_pointer20[15] ) );
INV_X4 _u0_U13429  ( .A(1'b1), .ZN(_u0_pointer20[14] ) );
INV_X4 _u0_U13427  ( .A(1'b1), .ZN(_u0_pointer20[13] ) );
INV_X4 _u0_U13425  ( .A(1'b1), .ZN(_u0_pointer20[12] ) );
INV_X4 _u0_U13423  ( .A(1'b1), .ZN(_u0_pointer20[11] ) );
INV_X4 _u0_U13421  ( .A(1'b1), .ZN(_u0_pointer20[10] ) );
INV_X4 _u0_U13419  ( .A(1'b1), .ZN(_u0_pointer20[9] ) );
INV_X4 _u0_U13417  ( .A(1'b1), .ZN(_u0_pointer20[8] ) );
INV_X4 _u0_U13415  ( .A(1'b1), .ZN(_u0_pointer20[7] ) );
INV_X4 _u0_U13413  ( .A(1'b1), .ZN(_u0_pointer20[6] ) );
INV_X4 _u0_U13411  ( .A(1'b1), .ZN(_u0_pointer20[5] ) );
INV_X4 _u0_U13409  ( .A(1'b1), .ZN(_u0_pointer20[4] ) );
INV_X4 _u0_U13407  ( .A(1'b1), .ZN(_u0_pointer20[3] ) );
INV_X4 _u0_U13405  ( .A(1'b1), .ZN(_u0_pointer20[2] ) );
INV_X4 _u0_U13403  ( .A(1'b1), .ZN(_u0_pointer20[1] ) );
INV_X4 _u0_U13401  ( .A(1'b1), .ZN(_u0_pointer20[0] ) );
INV_X4 _u0_U13399  ( .A(1'b1), .ZN(_u0_pointer20_s[31] ) );
INV_X4 _u0_U13397  ( .A(1'b1), .ZN(_u0_pointer20_s[30] ) );
INV_X4 _u0_U13395  ( .A(1'b1), .ZN(_u0_pointer20_s[29] ) );
INV_X4 _u0_U13393  ( .A(1'b1), .ZN(_u0_pointer20_s[28] ) );
INV_X4 _u0_U13391  ( .A(1'b1), .ZN(_u0_pointer20_s[27] ) );
INV_X4 _u0_U13389  ( .A(1'b1), .ZN(_u0_pointer20_s[26] ) );
INV_X4 _u0_U13387  ( .A(1'b1), .ZN(_u0_pointer20_s[25] ) );
INV_X4 _u0_U13385  ( .A(1'b1), .ZN(_u0_pointer20_s[24] ) );
INV_X4 _u0_U13383  ( .A(1'b1), .ZN(_u0_pointer20_s[23] ) );
INV_X4 _u0_U13381  ( .A(1'b1), .ZN(_u0_pointer20_s[22] ) );
INV_X4 _u0_U13379  ( .A(1'b1), .ZN(_u0_pointer20_s[21] ) );
INV_X4 _u0_U13377  ( .A(1'b1), .ZN(_u0_pointer20_s[20] ) );
INV_X4 _u0_U13375  ( .A(1'b1), .ZN(_u0_pointer20_s[19] ) );
INV_X4 _u0_U13373  ( .A(1'b1), .ZN(_u0_pointer20_s[18] ) );
INV_X4 _u0_U13371  ( .A(1'b1), .ZN(_u0_pointer20_s[17] ) );
INV_X4 _u0_U13369  ( .A(1'b1), .ZN(_u0_pointer20_s[16] ) );
INV_X4 _u0_U13367  ( .A(1'b1), .ZN(_u0_pointer20_s[15] ) );
INV_X4 _u0_U13365  ( .A(1'b1), .ZN(_u0_pointer20_s[14] ) );
INV_X4 _u0_U13363  ( .A(1'b1), .ZN(_u0_pointer20_s[13] ) );
INV_X4 _u0_U13361  ( .A(1'b1), .ZN(_u0_pointer20_s[12] ) );
INV_X4 _u0_U13359  ( .A(1'b1), .ZN(_u0_pointer20_s[11] ) );
INV_X4 _u0_U13357  ( .A(1'b1), .ZN(_u0_pointer20_s[10] ) );
INV_X4 _u0_U13355  ( .A(1'b1), .ZN(_u0_pointer20_s[9] ) );
INV_X4 _u0_U13353  ( .A(1'b1), .ZN(_u0_pointer20_s[8] ) );
INV_X4 _u0_U13351  ( .A(1'b1), .ZN(_u0_pointer20_s[7] ) );
INV_X4 _u0_U13349  ( .A(1'b1), .ZN(_u0_pointer20_s[6] ) );
INV_X4 _u0_U13347  ( .A(1'b1), .ZN(_u0_pointer20_s[5] ) );
INV_X4 _u0_U13345  ( .A(1'b1), .ZN(_u0_pointer20_s[4] ) );
INV_X4 _u0_U13343  ( .A(1'b1), .ZN(_u0_pointer20_s[3] ) );
INV_X4 _u0_U13341  ( .A(1'b1), .ZN(_u0_pointer20_s[2] ) );
INV_X4 _u0_U13339  ( .A(1'b1), .ZN(_u0_pointer20_s[1] ) );
INV_X4 _u0_U13337  ( .A(1'b1), .ZN(_u0_pointer20_s[0] ) );
INV_X4 _u0_U13335  ( .A(1'b1), .ZN(_u0_ch20_csr[31] ) );
INV_X4 _u0_U13333  ( .A(1'b1), .ZN(_u0_ch20_csr[30] ) );
INV_X4 _u0_U13331  ( .A(1'b1), .ZN(_u0_ch20_csr[29] ) );
INV_X4 _u0_U13329  ( .A(1'b1), .ZN(_u0_ch20_csr[28] ) );
INV_X4 _u0_U13327  ( .A(1'b1), .ZN(_u0_ch20_csr[27] ) );
INV_X4 _u0_U13325  ( .A(1'b1), .ZN(_u0_ch20_csr[26] ) );
INV_X4 _u0_U13323  ( .A(1'b1), .ZN(_u0_ch20_csr[25] ) );
INV_X4 _u0_U13321  ( .A(1'b1), .ZN(_u0_ch20_csr[24] ) );
INV_X4 _u0_U13319  ( .A(1'b1), .ZN(_u0_ch20_csr[23] ) );
INV_X4 _u0_U13317  ( .A(1'b1), .ZN(_u0_ch20_csr[22] ) );
INV_X4 _u0_U13315  ( .A(1'b1), .ZN(_u0_ch20_csr[21] ) );
INV_X4 _u0_U13313  ( .A(1'b1), .ZN(_u0_ch20_csr[20] ) );
INV_X4 _u0_U13311  ( .A(1'b1), .ZN(_u0_ch20_csr[19] ) );
INV_X4 _u0_U13309  ( .A(1'b1), .ZN(_u0_ch20_csr[18] ) );
INV_X4 _u0_U13307  ( .A(1'b1), .ZN(_u0_ch20_csr[17] ) );
INV_X4 _u0_U13305  ( .A(1'b1), .ZN(_u0_ch20_csr[16] ) );
INV_X4 _u0_U13303  ( .A(1'b1), .ZN(_u0_ch20_csr[15] ) );
INV_X4 _u0_U13301  ( .A(1'b1), .ZN(_u0_ch20_csr[14] ) );
INV_X4 _u0_U13299  ( .A(1'b1), .ZN(_u0_ch20_csr[13] ) );
INV_X4 _u0_U13297  ( .A(1'b1), .ZN(_u0_ch20_csr[12] ) );
INV_X4 _u0_U13295  ( .A(1'b1), .ZN(_u0_ch20_csr[11] ) );
INV_X4 _u0_U13293  ( .A(1'b1), .ZN(_u0_ch20_csr[10] ) );
INV_X4 _u0_U13291  ( .A(1'b1), .ZN(_u0_ch20_csr[9] ) );
INV_X4 _u0_U13289  ( .A(1'b1), .ZN(_u0_ch20_csr[8] ) );
INV_X4 _u0_U13287  ( .A(1'b1), .ZN(_u0_ch20_csr[7] ) );
INV_X4 _u0_U13285  ( .A(1'b1), .ZN(_u0_ch20_csr[6] ) );
INV_X4 _u0_U13283  ( .A(1'b1), .ZN(_u0_ch20_csr[5] ) );
INV_X4 _u0_U13281  ( .A(1'b1), .ZN(_u0_ch20_csr[4] ) );
INV_X4 _u0_U13279  ( .A(1'b1), .ZN(_u0_ch20_csr[3] ) );
INV_X4 _u0_U13277  ( .A(1'b1), .ZN(_u0_ch20_csr[2] ) );
INV_X4 _u0_U13275  ( .A(1'b1), .ZN(_u0_ch20_csr[1] ) );
INV_X4 _u0_U13273  ( .A(1'b1), .ZN(_u0_ch20_csr[0] ) );
INV_X4 _u0_U13271  ( .A(1'b1), .ZN(_u0_ch20_txsz[31] ) );
INV_X4 _u0_U13269  ( .A(1'b1), .ZN(_u0_ch20_txsz[30] ) );
INV_X4 _u0_U13267  ( .A(1'b1), .ZN(_u0_ch20_txsz[29] ) );
INV_X4 _u0_U13265  ( .A(1'b1), .ZN(_u0_ch20_txsz[28] ) );
INV_X4 _u0_U13263  ( .A(1'b1), .ZN(_u0_ch20_txsz[27] ) );
INV_X4 _u0_U13261  ( .A(1'b1), .ZN(_u0_ch20_txsz[26] ) );
INV_X4 _u0_U13259  ( .A(1'b1), .ZN(_u0_ch20_txsz[25] ) );
INV_X4 _u0_U13257  ( .A(1'b1), .ZN(_u0_ch20_txsz[24] ) );
INV_X4 _u0_U13255  ( .A(1'b1), .ZN(_u0_ch20_txsz[23] ) );
INV_X4 _u0_U13253  ( .A(1'b1), .ZN(_u0_ch20_txsz[22] ) );
INV_X4 _u0_U13251  ( .A(1'b1), .ZN(_u0_ch20_txsz[21] ) );
INV_X4 _u0_U13249  ( .A(1'b1), .ZN(_u0_ch20_txsz[20] ) );
INV_X4 _u0_U13247  ( .A(1'b1), .ZN(_u0_ch20_txsz[19] ) );
INV_X4 _u0_U13245  ( .A(1'b1), .ZN(_u0_ch20_txsz[18] ) );
INV_X4 _u0_U13243  ( .A(1'b1), .ZN(_u0_ch20_txsz[17] ) );
INV_X4 _u0_U13241  ( .A(1'b1), .ZN(_u0_ch20_txsz[16] ) );
INV_X4 _u0_U13239  ( .A(1'b1), .ZN(_u0_ch20_txsz[15] ) );
INV_X4 _u0_U13237  ( .A(1'b1), .ZN(_u0_ch20_txsz[14] ) );
INV_X4 _u0_U13235  ( .A(1'b1), .ZN(_u0_ch20_txsz[13] ) );
INV_X4 _u0_U13233  ( .A(1'b1), .ZN(_u0_ch20_txsz[12] ) );
INV_X4 _u0_U13231  ( .A(1'b1), .ZN(_u0_ch20_txsz[11] ) );
INV_X4 _u0_U13229  ( .A(1'b1), .ZN(_u0_ch20_txsz[10] ) );
INV_X4 _u0_U13227  ( .A(1'b1), .ZN(_u0_ch20_txsz[9] ) );
INV_X4 _u0_U13225  ( .A(1'b1), .ZN(_u0_ch20_txsz[8] ) );
INV_X4 _u0_U13223  ( .A(1'b1), .ZN(_u0_ch20_txsz[7] ) );
INV_X4 _u0_U13221  ( .A(1'b1), .ZN(_u0_ch20_txsz[6] ) );
INV_X4 _u0_U13219  ( .A(1'b1), .ZN(_u0_ch20_txsz[5] ) );
INV_X4 _u0_U13217  ( .A(1'b1), .ZN(_u0_ch20_txsz[4] ) );
INV_X4 _u0_U13215  ( .A(1'b1), .ZN(_u0_ch20_txsz[3] ) );
INV_X4 _u0_U13213  ( .A(1'b1), .ZN(_u0_ch20_txsz[2] ) );
INV_X4 _u0_U13211  ( .A(1'b1), .ZN(_u0_ch20_txsz[1] ) );
INV_X4 _u0_U13209  ( .A(1'b1), .ZN(_u0_ch20_txsz[0] ) );
INV_X4 _u0_U13207  ( .A(1'b1), .ZN(_u0_ch20_adr0[31] ) );
INV_X4 _u0_U13205  ( .A(1'b1), .ZN(_u0_ch20_adr0[30] ) );
INV_X4 _u0_U13203  ( .A(1'b1), .ZN(_u0_ch20_adr0[29] ) );
INV_X4 _u0_U13201  ( .A(1'b1), .ZN(_u0_ch20_adr0[28] ) );
INV_X4 _u0_U13199  ( .A(1'b1), .ZN(_u0_ch20_adr0[27] ) );
INV_X4 _u0_U13197  ( .A(1'b1), .ZN(_u0_ch20_adr0[26] ) );
INV_X4 _u0_U13195  ( .A(1'b1), .ZN(_u0_ch20_adr0[25] ) );
INV_X4 _u0_U13193  ( .A(1'b1), .ZN(_u0_ch20_adr0[24] ) );
INV_X4 _u0_U13191  ( .A(1'b1), .ZN(_u0_ch20_adr0[23] ) );
INV_X4 _u0_U13189  ( .A(1'b1), .ZN(_u0_ch20_adr0[22] ) );
INV_X4 _u0_U13187  ( .A(1'b1), .ZN(_u0_ch20_adr0[21] ) );
INV_X4 _u0_U13185  ( .A(1'b1), .ZN(_u0_ch20_adr0[20] ) );
INV_X4 _u0_U13183  ( .A(1'b1), .ZN(_u0_ch20_adr0[19] ) );
INV_X4 _u0_U13181  ( .A(1'b1), .ZN(_u0_ch20_adr0[18] ) );
INV_X4 _u0_U13179  ( .A(1'b1), .ZN(_u0_ch20_adr0[17] ) );
INV_X4 _u0_U13177  ( .A(1'b1), .ZN(_u0_ch20_adr0[16] ) );
INV_X4 _u0_U13175  ( .A(1'b1), .ZN(_u0_ch20_adr0[15] ) );
INV_X4 _u0_U13173  ( .A(1'b1), .ZN(_u0_ch20_adr0[14] ) );
INV_X4 _u0_U13171  ( .A(1'b1), .ZN(_u0_ch20_adr0[13] ) );
INV_X4 _u0_U13169  ( .A(1'b1), .ZN(_u0_ch20_adr0[12] ) );
INV_X4 _u0_U13167  ( .A(1'b1), .ZN(_u0_ch20_adr0[11] ) );
INV_X4 _u0_U13165  ( .A(1'b1), .ZN(_u0_ch20_adr0[10] ) );
INV_X4 _u0_U13163  ( .A(1'b1), .ZN(_u0_ch20_adr0[9] ) );
INV_X4 _u0_U13161  ( .A(1'b1), .ZN(_u0_ch20_adr0[8] ) );
INV_X4 _u0_U13159  ( .A(1'b1), .ZN(_u0_ch20_adr0[7] ) );
INV_X4 _u0_U13157  ( .A(1'b1), .ZN(_u0_ch20_adr0[6] ) );
INV_X4 _u0_U13155  ( .A(1'b1), .ZN(_u0_ch20_adr0[5] ) );
INV_X4 _u0_U13153  ( .A(1'b1), .ZN(_u0_ch20_adr0[4] ) );
INV_X4 _u0_U13151  ( .A(1'b1), .ZN(_u0_ch20_adr0[3] ) );
INV_X4 _u0_U13149  ( .A(1'b1), .ZN(_u0_ch20_adr0[2] ) );
INV_X4 _u0_U13147  ( .A(1'b1), .ZN(_u0_ch20_adr0[1] ) );
INV_X4 _u0_U13145  ( .A(1'b1), .ZN(_u0_ch20_adr0[0] ) );
INV_X4 _u0_U13143  ( .A(1'b1), .ZN(_u0_ch20_adr1[31] ) );
INV_X4 _u0_U13141  ( .A(1'b1), .ZN(_u0_ch20_adr1[30] ) );
INV_X4 _u0_U13139  ( .A(1'b1), .ZN(_u0_ch20_adr1[29] ) );
INV_X4 _u0_U13137  ( .A(1'b1), .ZN(_u0_ch20_adr1[28] ) );
INV_X4 _u0_U13135  ( .A(1'b1), .ZN(_u0_ch20_adr1[27] ) );
INV_X4 _u0_U13133  ( .A(1'b1), .ZN(_u0_ch20_adr1[26] ) );
INV_X4 _u0_U13131  ( .A(1'b1), .ZN(_u0_ch20_adr1[25] ) );
INV_X4 _u0_U13129  ( .A(1'b1), .ZN(_u0_ch20_adr1[24] ) );
INV_X4 _u0_U13127  ( .A(1'b1), .ZN(_u0_ch20_adr1[23] ) );
INV_X4 _u0_U13125  ( .A(1'b1), .ZN(_u0_ch20_adr1[22] ) );
INV_X4 _u0_U13123  ( .A(1'b1), .ZN(_u0_ch20_adr1[21] ) );
INV_X4 _u0_U13121  ( .A(1'b1), .ZN(_u0_ch20_adr1[20] ) );
INV_X4 _u0_U13119  ( .A(1'b1), .ZN(_u0_ch20_adr1[19] ) );
INV_X4 _u0_U13117  ( .A(1'b1), .ZN(_u0_ch20_adr1[18] ) );
INV_X4 _u0_U13115  ( .A(1'b1), .ZN(_u0_ch20_adr1[17] ) );
INV_X4 _u0_U13113  ( .A(1'b1), .ZN(_u0_ch20_adr1[16] ) );
INV_X4 _u0_U13111  ( .A(1'b1), .ZN(_u0_ch20_adr1[15] ) );
INV_X4 _u0_U13109  ( .A(1'b1), .ZN(_u0_ch20_adr1[14] ) );
INV_X4 _u0_U13107  ( .A(1'b1), .ZN(_u0_ch20_adr1[13] ) );
INV_X4 _u0_U13105  ( .A(1'b1), .ZN(_u0_ch20_adr1[12] ) );
INV_X4 _u0_U13103  ( .A(1'b1), .ZN(_u0_ch20_adr1[11] ) );
INV_X4 _u0_U13101  ( .A(1'b1), .ZN(_u0_ch20_adr1[10] ) );
INV_X4 _u0_U13099  ( .A(1'b1), .ZN(_u0_ch20_adr1[9] ) );
INV_X4 _u0_U13097  ( .A(1'b1), .ZN(_u0_ch20_adr1[8] ) );
INV_X4 _u0_U13095  ( .A(1'b1), .ZN(_u0_ch20_adr1[7] ) );
INV_X4 _u0_U13093  ( .A(1'b1), .ZN(_u0_ch20_adr1[6] ) );
INV_X4 _u0_U13091  ( .A(1'b1), .ZN(_u0_ch20_adr1[5] ) );
INV_X4 _u0_U13089  ( .A(1'b1), .ZN(_u0_ch20_adr1[4] ) );
INV_X4 _u0_U13087  ( .A(1'b1), .ZN(_u0_ch20_adr1[3] ) );
INV_X4 _u0_U13085  ( .A(1'b1), .ZN(_u0_ch20_adr1[2] ) );
INV_X4 _u0_U13083  ( .A(1'b1), .ZN(_u0_ch20_adr1[1] ) );
INV_X4 _u0_U13081  ( .A(1'b1), .ZN(_u0_ch20_adr1[0] ) );
INV_X4 _u0_U13079  ( .A(1'b0), .ZN(_u0_ch20_am0[31] ) );
INV_X4 _u0_U13077  ( .A(1'b0), .ZN(_u0_ch20_am0[30] ) );
INV_X4 _u0_U13075  ( .A(1'b0), .ZN(_u0_ch20_am0[29] ) );
INV_X4 _u0_U13073  ( .A(1'b0), .ZN(_u0_ch20_am0[28] ) );
INV_X4 _u0_U13071  ( .A(1'b0), .ZN(_u0_ch20_am0[27] ) );
INV_X4 _u0_U13069  ( .A(1'b0), .ZN(_u0_ch20_am0[26] ) );
INV_X4 _u0_U13067  ( .A(1'b0), .ZN(_u0_ch20_am0[25] ) );
INV_X4 _u0_U13065  ( .A(1'b0), .ZN(_u0_ch20_am0[24] ) );
INV_X4 _u0_U13063  ( .A(1'b0), .ZN(_u0_ch20_am0[23] ) );
INV_X4 _u0_U13061  ( .A(1'b0), .ZN(_u0_ch20_am0[22] ) );
INV_X4 _u0_U13059  ( .A(1'b0), .ZN(_u0_ch20_am0[21] ) );
INV_X4 _u0_U13057  ( .A(1'b0), .ZN(_u0_ch20_am0[20] ) );
INV_X4 _u0_U13055  ( .A(1'b0), .ZN(_u0_ch20_am0[19] ) );
INV_X4 _u0_U13053  ( .A(1'b0), .ZN(_u0_ch20_am0[18] ) );
INV_X4 _u0_U13051  ( .A(1'b0), .ZN(_u0_ch20_am0[17] ) );
INV_X4 _u0_U13049  ( .A(1'b0), .ZN(_u0_ch20_am0[16] ) );
INV_X4 _u0_U13047  ( .A(1'b0), .ZN(_u0_ch20_am0[15] ) );
INV_X4 _u0_U13045  ( .A(1'b0), .ZN(_u0_ch20_am0[14] ) );
INV_X4 _u0_U13043  ( .A(1'b0), .ZN(_u0_ch20_am0[13] ) );
INV_X4 _u0_U13041  ( .A(1'b0), .ZN(_u0_ch20_am0[12] ) );
INV_X4 _u0_U13039  ( .A(1'b0), .ZN(_u0_ch20_am0[11] ) );
INV_X4 _u0_U13037  ( .A(1'b0), .ZN(_u0_ch20_am0[10] ) );
INV_X4 _u0_U13035  ( .A(1'b0), .ZN(_u0_ch20_am0[9] ) );
INV_X4 _u0_U13033  ( .A(1'b0), .ZN(_u0_ch20_am0[8] ) );
INV_X4 _u0_U13031  ( .A(1'b0), .ZN(_u0_ch20_am0[7] ) );
INV_X4 _u0_U13029  ( .A(1'b0), .ZN(_u0_ch20_am0[6] ) );
INV_X4 _u0_U13027  ( .A(1'b0), .ZN(_u0_ch20_am0[5] ) );
INV_X4 _u0_U13025  ( .A(1'b0), .ZN(_u0_ch20_am0[4] ) );
INV_X4 _u0_U13023  ( .A(1'b1), .ZN(_u0_ch20_am0[3] ) );
INV_X4 _u0_U13021  ( .A(1'b1), .ZN(_u0_ch20_am0[2] ) );
INV_X4 _u0_U13019  ( .A(1'b1), .ZN(_u0_ch20_am0[1] ) );
INV_X4 _u0_U13017  ( .A(1'b1), .ZN(_u0_ch20_am0[0] ) );
INV_X4 _u0_U13015  ( .A(1'b0), .ZN(_u0_ch20_am1[31] ) );
INV_X4 _u0_U13013  ( .A(1'b0), .ZN(_u0_ch20_am1[30] ) );
INV_X4 _u0_U13011  ( .A(1'b0), .ZN(_u0_ch20_am1[29] ) );
INV_X4 _u0_U13009  ( .A(1'b0), .ZN(_u0_ch20_am1[28] ) );
INV_X4 _u0_U13007  ( .A(1'b0), .ZN(_u0_ch20_am1[27] ) );
INV_X4 _u0_U13005  ( .A(1'b0), .ZN(_u0_ch20_am1[26] ) );
INV_X4 _u0_U13003  ( .A(1'b0), .ZN(_u0_ch20_am1[25] ) );
INV_X4 _u0_U13001  ( .A(1'b0), .ZN(_u0_ch20_am1[24] ) );
INV_X4 _u0_U12999  ( .A(1'b0), .ZN(_u0_ch20_am1[23] ) );
INV_X4 _u0_U12997  ( .A(1'b0), .ZN(_u0_ch20_am1[22] ) );
INV_X4 _u0_U12995  ( .A(1'b0), .ZN(_u0_ch20_am1[21] ) );
INV_X4 _u0_U12993  ( .A(1'b0), .ZN(_u0_ch20_am1[20] ) );
INV_X4 _u0_U12991  ( .A(1'b0), .ZN(_u0_ch20_am1[19] ) );
INV_X4 _u0_U12989  ( .A(1'b0), .ZN(_u0_ch20_am1[18] ) );
INV_X4 _u0_U12987  ( .A(1'b0), .ZN(_u0_ch20_am1[17] ) );
INV_X4 _u0_U12985  ( .A(1'b0), .ZN(_u0_ch20_am1[16] ) );
INV_X4 _u0_U12983  ( .A(1'b0), .ZN(_u0_ch20_am1[15] ) );
INV_X4 _u0_U12981  ( .A(1'b0), .ZN(_u0_ch20_am1[14] ) );
INV_X4 _u0_U12979  ( .A(1'b0), .ZN(_u0_ch20_am1[13] ) );
INV_X4 _u0_U12977  ( .A(1'b0), .ZN(_u0_ch20_am1[12] ) );
INV_X4 _u0_U12975  ( .A(1'b0), .ZN(_u0_ch20_am1[11] ) );
INV_X4 _u0_U12973  ( .A(1'b0), .ZN(_u0_ch20_am1[10] ) );
INV_X4 _u0_U12971  ( .A(1'b0), .ZN(_u0_ch20_am1[9] ) );
INV_X4 _u0_U12969  ( .A(1'b0), .ZN(_u0_ch20_am1[8] ) );
INV_X4 _u0_U12967  ( .A(1'b0), .ZN(_u0_ch20_am1[7] ) );
INV_X4 _u0_U12965  ( .A(1'b0), .ZN(_u0_ch20_am1[6] ) );
INV_X4 _u0_U12963  ( .A(1'b0), .ZN(_u0_ch20_am1[5] ) );
INV_X4 _u0_U12961  ( .A(1'b0), .ZN(_u0_ch20_am1[4] ) );
INV_X4 _u0_U12959  ( .A(1'b1), .ZN(_u0_ch20_am1[3] ) );
INV_X4 _u0_U12957  ( .A(1'b1), .ZN(_u0_ch20_am1[2] ) );
INV_X4 _u0_U12955  ( .A(1'b1), .ZN(_u0_ch20_am1[1] ) );
INV_X4 _u0_U12953  ( .A(1'b1), .ZN(_u0_ch20_am1[0] ) );
INV_X4 _u0_U12951  ( .A(1'b1), .ZN(_u0_pointer21[31] ) );
INV_X4 _u0_U12949  ( .A(1'b1), .ZN(_u0_pointer21[30] ) );
INV_X4 _u0_U12947  ( .A(1'b1), .ZN(_u0_pointer21[29] ) );
INV_X4 _u0_U12945  ( .A(1'b1), .ZN(_u0_pointer21[28] ) );
INV_X4 _u0_U12943  ( .A(1'b1), .ZN(_u0_pointer21[27] ) );
INV_X4 _u0_U12941  ( .A(1'b1), .ZN(_u0_pointer21[26] ) );
INV_X4 _u0_U12939  ( .A(1'b1), .ZN(_u0_pointer21[25] ) );
INV_X4 _u0_U12937  ( .A(1'b1), .ZN(_u0_pointer21[24] ) );
INV_X4 _u0_U12935  ( .A(1'b1), .ZN(_u0_pointer21[23] ) );
INV_X4 _u0_U12933  ( .A(1'b1), .ZN(_u0_pointer21[22] ) );
INV_X4 _u0_U12931  ( .A(1'b1), .ZN(_u0_pointer21[21] ) );
INV_X4 _u0_U12929  ( .A(1'b1), .ZN(_u0_pointer21[20] ) );
INV_X4 _u0_U12927  ( .A(1'b1), .ZN(_u0_pointer21[19] ) );
INV_X4 _u0_U12925  ( .A(1'b1), .ZN(_u0_pointer21[18] ) );
INV_X4 _u0_U12923  ( .A(1'b1), .ZN(_u0_pointer21[17] ) );
INV_X4 _u0_U12921  ( .A(1'b1), .ZN(_u0_pointer21[16] ) );
INV_X4 _u0_U12919  ( .A(1'b1), .ZN(_u0_pointer21[15] ) );
INV_X4 _u0_U12917  ( .A(1'b1), .ZN(_u0_pointer21[14] ) );
INV_X4 _u0_U12915  ( .A(1'b1), .ZN(_u0_pointer21[13] ) );
INV_X4 _u0_U12913  ( .A(1'b1), .ZN(_u0_pointer21[12] ) );
INV_X4 _u0_U12911  ( .A(1'b1), .ZN(_u0_pointer21[11] ) );
INV_X4 _u0_U12909  ( .A(1'b1), .ZN(_u0_pointer21[10] ) );
INV_X4 _u0_U12907  ( .A(1'b1), .ZN(_u0_pointer21[9] ) );
INV_X4 _u0_U12905  ( .A(1'b1), .ZN(_u0_pointer21[8] ) );
INV_X4 _u0_U12903  ( .A(1'b1), .ZN(_u0_pointer21[7] ) );
INV_X4 _u0_U12901  ( .A(1'b1), .ZN(_u0_pointer21[6] ) );
INV_X4 _u0_U12899  ( .A(1'b1), .ZN(_u0_pointer21[5] ) );
INV_X4 _u0_U12897  ( .A(1'b1), .ZN(_u0_pointer21[4] ) );
INV_X4 _u0_U12895  ( .A(1'b1), .ZN(_u0_pointer21[3] ) );
INV_X4 _u0_U12893  ( .A(1'b1), .ZN(_u0_pointer21[2] ) );
INV_X4 _u0_U12891  ( .A(1'b1), .ZN(_u0_pointer21[1] ) );
INV_X4 _u0_U12889  ( .A(1'b1), .ZN(_u0_pointer21[0] ) );
INV_X4 _u0_U12887  ( .A(1'b1), .ZN(_u0_pointer21_s[31] ) );
INV_X4 _u0_U12885  ( .A(1'b1), .ZN(_u0_pointer21_s[30] ) );
INV_X4 _u0_U12883  ( .A(1'b1), .ZN(_u0_pointer21_s[29] ) );
INV_X4 _u0_U12881  ( .A(1'b1), .ZN(_u0_pointer21_s[28] ) );
INV_X4 _u0_U12879  ( .A(1'b1), .ZN(_u0_pointer21_s[27] ) );
INV_X4 _u0_U12877  ( .A(1'b1), .ZN(_u0_pointer21_s[26] ) );
INV_X4 _u0_U12875  ( .A(1'b1), .ZN(_u0_pointer21_s[25] ) );
INV_X4 _u0_U12873  ( .A(1'b1), .ZN(_u0_pointer21_s[24] ) );
INV_X4 _u0_U12871  ( .A(1'b1), .ZN(_u0_pointer21_s[23] ) );
INV_X4 _u0_U12869  ( .A(1'b1), .ZN(_u0_pointer21_s[22] ) );
INV_X4 _u0_U12867  ( .A(1'b1), .ZN(_u0_pointer21_s[21] ) );
INV_X4 _u0_U12865  ( .A(1'b1), .ZN(_u0_pointer21_s[20] ) );
INV_X4 _u0_U12863  ( .A(1'b1), .ZN(_u0_pointer21_s[19] ) );
INV_X4 _u0_U12861  ( .A(1'b1), .ZN(_u0_pointer21_s[18] ) );
INV_X4 _u0_U12859  ( .A(1'b1), .ZN(_u0_pointer21_s[17] ) );
INV_X4 _u0_U12857  ( .A(1'b1), .ZN(_u0_pointer21_s[16] ) );
INV_X4 _u0_U12855  ( .A(1'b1), .ZN(_u0_pointer21_s[15] ) );
INV_X4 _u0_U12853  ( .A(1'b1), .ZN(_u0_pointer21_s[14] ) );
INV_X4 _u0_U12851  ( .A(1'b1), .ZN(_u0_pointer21_s[13] ) );
INV_X4 _u0_U12849  ( .A(1'b1), .ZN(_u0_pointer21_s[12] ) );
INV_X4 _u0_U12847  ( .A(1'b1), .ZN(_u0_pointer21_s[11] ) );
INV_X4 _u0_U12845  ( .A(1'b1), .ZN(_u0_pointer21_s[10] ) );
INV_X4 _u0_U12843  ( .A(1'b1), .ZN(_u0_pointer21_s[9] ) );
INV_X4 _u0_U12841  ( .A(1'b1), .ZN(_u0_pointer21_s[8] ) );
INV_X4 _u0_U12839  ( .A(1'b1), .ZN(_u0_pointer21_s[7] ) );
INV_X4 _u0_U12837  ( .A(1'b1), .ZN(_u0_pointer21_s[6] ) );
INV_X4 _u0_U12835  ( .A(1'b1), .ZN(_u0_pointer21_s[5] ) );
INV_X4 _u0_U12833  ( .A(1'b1), .ZN(_u0_pointer21_s[4] ) );
INV_X4 _u0_U12831  ( .A(1'b1), .ZN(_u0_pointer21_s[3] ) );
INV_X4 _u0_U12829  ( .A(1'b1), .ZN(_u0_pointer21_s[2] ) );
INV_X4 _u0_U12827  ( .A(1'b1), .ZN(_u0_pointer21_s[1] ) );
INV_X4 _u0_U12825  ( .A(1'b1), .ZN(_u0_pointer21_s[0] ) );
INV_X4 _u0_U12823  ( .A(1'b1), .ZN(_u0_ch21_csr[31] ) );
INV_X4 _u0_U12821  ( .A(1'b1), .ZN(_u0_ch21_csr[30] ) );
INV_X4 _u0_U12819  ( .A(1'b1), .ZN(_u0_ch21_csr[29] ) );
INV_X4 _u0_U12817  ( .A(1'b1), .ZN(_u0_ch21_csr[28] ) );
INV_X4 _u0_U12815  ( .A(1'b1), .ZN(_u0_ch21_csr[27] ) );
INV_X4 _u0_U12813  ( .A(1'b1), .ZN(_u0_ch21_csr[26] ) );
INV_X4 _u0_U12811  ( .A(1'b1), .ZN(_u0_ch21_csr[25] ) );
INV_X4 _u0_U12809  ( .A(1'b1), .ZN(_u0_ch21_csr[24] ) );
INV_X4 _u0_U12807  ( .A(1'b1), .ZN(_u0_ch21_csr[23] ) );
INV_X4 _u0_U12805  ( .A(1'b1), .ZN(_u0_ch21_csr[22] ) );
INV_X4 _u0_U12803  ( .A(1'b1), .ZN(_u0_ch21_csr[21] ) );
INV_X4 _u0_U12801  ( .A(1'b1), .ZN(_u0_ch21_csr[20] ) );
INV_X4 _u0_U12799  ( .A(1'b1), .ZN(_u0_ch21_csr[19] ) );
INV_X4 _u0_U12797  ( .A(1'b1), .ZN(_u0_ch21_csr[18] ) );
INV_X4 _u0_U12795  ( .A(1'b1), .ZN(_u0_ch21_csr[17] ) );
INV_X4 _u0_U12793  ( .A(1'b1), .ZN(_u0_ch21_csr[16] ) );
INV_X4 _u0_U12791  ( .A(1'b1), .ZN(_u0_ch21_csr[15] ) );
INV_X4 _u0_U12789  ( .A(1'b1), .ZN(_u0_ch21_csr[14] ) );
INV_X4 _u0_U12787  ( .A(1'b1), .ZN(_u0_ch21_csr[13] ) );
INV_X4 _u0_U12785  ( .A(1'b1), .ZN(_u0_ch21_csr[12] ) );
INV_X4 _u0_U12783  ( .A(1'b1), .ZN(_u0_ch21_csr[11] ) );
INV_X4 _u0_U12781  ( .A(1'b1), .ZN(_u0_ch21_csr[10] ) );
INV_X4 _u0_U12779  ( .A(1'b1), .ZN(_u0_ch21_csr[9] ) );
INV_X4 _u0_U12777  ( .A(1'b1), .ZN(_u0_ch21_csr[8] ) );
INV_X4 _u0_U12775  ( .A(1'b1), .ZN(_u0_ch21_csr[7] ) );
INV_X4 _u0_U12773  ( .A(1'b1), .ZN(_u0_ch21_csr[6] ) );
INV_X4 _u0_U12771  ( .A(1'b1), .ZN(_u0_ch21_csr[5] ) );
INV_X4 _u0_U12769  ( .A(1'b1), .ZN(_u0_ch21_csr[4] ) );
INV_X4 _u0_U12767  ( .A(1'b1), .ZN(_u0_ch21_csr[3] ) );
INV_X4 _u0_U12765  ( .A(1'b1), .ZN(_u0_ch21_csr[2] ) );
INV_X4 _u0_U12763  ( .A(1'b1), .ZN(_u0_ch21_csr[1] ) );
INV_X4 _u0_U12761  ( .A(1'b1), .ZN(_u0_ch21_csr[0] ) );
INV_X4 _u0_U12759  ( .A(1'b1), .ZN(_u0_ch21_txsz[31] ) );
INV_X4 _u0_U12757  ( .A(1'b1), .ZN(_u0_ch21_txsz[30] ) );
INV_X4 _u0_U12755  ( .A(1'b1), .ZN(_u0_ch21_txsz[29] ) );
INV_X4 _u0_U12753  ( .A(1'b1), .ZN(_u0_ch21_txsz[28] ) );
INV_X4 _u0_U12751  ( .A(1'b1), .ZN(_u0_ch21_txsz[27] ) );
INV_X4 _u0_U12749  ( .A(1'b1), .ZN(_u0_ch21_txsz[26] ) );
INV_X4 _u0_U12747  ( .A(1'b1), .ZN(_u0_ch21_txsz[25] ) );
INV_X4 _u0_U12745  ( .A(1'b1), .ZN(_u0_ch21_txsz[24] ) );
INV_X4 _u0_U12743  ( .A(1'b1), .ZN(_u0_ch21_txsz[23] ) );
INV_X4 _u0_U12741  ( .A(1'b1), .ZN(_u0_ch21_txsz[22] ) );
INV_X4 _u0_U12739  ( .A(1'b1), .ZN(_u0_ch21_txsz[21] ) );
INV_X4 _u0_U12737  ( .A(1'b1), .ZN(_u0_ch21_txsz[20] ) );
INV_X4 _u0_U12735  ( .A(1'b1), .ZN(_u0_ch21_txsz[19] ) );
INV_X4 _u0_U12733  ( .A(1'b1), .ZN(_u0_ch21_txsz[18] ) );
INV_X4 _u0_U12731  ( .A(1'b1), .ZN(_u0_ch21_txsz[17] ) );
INV_X4 _u0_U12729  ( .A(1'b1), .ZN(_u0_ch21_txsz[16] ) );
INV_X4 _u0_U12727  ( .A(1'b1), .ZN(_u0_ch21_txsz[15] ) );
INV_X4 _u0_U12725  ( .A(1'b1), .ZN(_u0_ch21_txsz[14] ) );
INV_X4 _u0_U12723  ( .A(1'b1), .ZN(_u0_ch21_txsz[13] ) );
INV_X4 _u0_U12721  ( .A(1'b1), .ZN(_u0_ch21_txsz[12] ) );
INV_X4 _u0_U12719  ( .A(1'b1), .ZN(_u0_ch21_txsz[11] ) );
INV_X4 _u0_U12717  ( .A(1'b1), .ZN(_u0_ch21_txsz[10] ) );
INV_X4 _u0_U12715  ( .A(1'b1), .ZN(_u0_ch21_txsz[9] ) );
INV_X4 _u0_U12713  ( .A(1'b1), .ZN(_u0_ch21_txsz[8] ) );
INV_X4 _u0_U12711  ( .A(1'b1), .ZN(_u0_ch21_txsz[7] ) );
INV_X4 _u0_U12709  ( .A(1'b1), .ZN(_u0_ch21_txsz[6] ) );
INV_X4 _u0_U12707  ( .A(1'b1), .ZN(_u0_ch21_txsz[5] ) );
INV_X4 _u0_U12705  ( .A(1'b1), .ZN(_u0_ch21_txsz[4] ) );
INV_X4 _u0_U12703  ( .A(1'b1), .ZN(_u0_ch21_txsz[3] ) );
INV_X4 _u0_U12701  ( .A(1'b1), .ZN(_u0_ch21_txsz[2] ) );
INV_X4 _u0_U12699  ( .A(1'b1), .ZN(_u0_ch21_txsz[1] ) );
INV_X4 _u0_U12697  ( .A(1'b1), .ZN(_u0_ch21_txsz[0] ) );
INV_X4 _u0_U12695  ( .A(1'b1), .ZN(_u0_ch21_adr0[31] ) );
INV_X4 _u0_U12693  ( .A(1'b1), .ZN(_u0_ch21_adr0[30] ) );
INV_X4 _u0_U12691  ( .A(1'b1), .ZN(_u0_ch21_adr0[29] ) );
INV_X4 _u0_U12689  ( .A(1'b1), .ZN(_u0_ch21_adr0[28] ) );
INV_X4 _u0_U12687  ( .A(1'b1), .ZN(_u0_ch21_adr0[27] ) );
INV_X4 _u0_U12685  ( .A(1'b1), .ZN(_u0_ch21_adr0[26] ) );
INV_X4 _u0_U12683  ( .A(1'b1), .ZN(_u0_ch21_adr0[25] ) );
INV_X4 _u0_U12681  ( .A(1'b1), .ZN(_u0_ch21_adr0[24] ) );
INV_X4 _u0_U12679  ( .A(1'b1), .ZN(_u0_ch21_adr0[23] ) );
INV_X4 _u0_U12677  ( .A(1'b1), .ZN(_u0_ch21_adr0[22] ) );
INV_X4 _u0_U12675  ( .A(1'b1), .ZN(_u0_ch21_adr0[21] ) );
INV_X4 _u0_U12673  ( .A(1'b1), .ZN(_u0_ch21_adr0[20] ) );
INV_X4 _u0_U12671  ( .A(1'b1), .ZN(_u0_ch21_adr0[19] ) );
INV_X4 _u0_U12669  ( .A(1'b1), .ZN(_u0_ch21_adr0[18] ) );
INV_X4 _u0_U12667  ( .A(1'b1), .ZN(_u0_ch21_adr0[17] ) );
INV_X4 _u0_U12665  ( .A(1'b1), .ZN(_u0_ch21_adr0[16] ) );
INV_X4 _u0_U12663  ( .A(1'b1), .ZN(_u0_ch21_adr0[15] ) );
INV_X4 _u0_U12661  ( .A(1'b1), .ZN(_u0_ch21_adr0[14] ) );
INV_X4 _u0_U12659  ( .A(1'b1), .ZN(_u0_ch21_adr0[13] ) );
INV_X4 _u0_U12657  ( .A(1'b1), .ZN(_u0_ch21_adr0[12] ) );
INV_X4 _u0_U12655  ( .A(1'b1), .ZN(_u0_ch21_adr0[11] ) );
INV_X4 _u0_U12653  ( .A(1'b1), .ZN(_u0_ch21_adr0[10] ) );
INV_X4 _u0_U12651  ( .A(1'b1), .ZN(_u0_ch21_adr0[9] ) );
INV_X4 _u0_U12649  ( .A(1'b1), .ZN(_u0_ch21_adr0[8] ) );
INV_X4 _u0_U12647  ( .A(1'b1), .ZN(_u0_ch21_adr0[7] ) );
INV_X4 _u0_U12645  ( .A(1'b1), .ZN(_u0_ch21_adr0[6] ) );
INV_X4 _u0_U12643  ( .A(1'b1), .ZN(_u0_ch21_adr0[5] ) );
INV_X4 _u0_U12641  ( .A(1'b1), .ZN(_u0_ch21_adr0[4] ) );
INV_X4 _u0_U12639  ( .A(1'b1), .ZN(_u0_ch21_adr0[3] ) );
INV_X4 _u0_U12637  ( .A(1'b1), .ZN(_u0_ch21_adr0[2] ) );
INV_X4 _u0_U12635  ( .A(1'b1), .ZN(_u0_ch21_adr0[1] ) );
INV_X4 _u0_U12633  ( .A(1'b1), .ZN(_u0_ch21_adr0[0] ) );
INV_X4 _u0_U12631  ( .A(1'b1), .ZN(_u0_ch21_adr1[31] ) );
INV_X4 _u0_U12629  ( .A(1'b1), .ZN(_u0_ch21_adr1[30] ) );
INV_X4 _u0_U12627  ( .A(1'b1), .ZN(_u0_ch21_adr1[29] ) );
INV_X4 _u0_U12625  ( .A(1'b1), .ZN(_u0_ch21_adr1[28] ) );
INV_X4 _u0_U12623  ( .A(1'b1), .ZN(_u0_ch21_adr1[27] ) );
INV_X4 _u0_U12621  ( .A(1'b1), .ZN(_u0_ch21_adr1[26] ) );
INV_X4 _u0_U12619  ( .A(1'b1), .ZN(_u0_ch21_adr1[25] ) );
INV_X4 _u0_U12617  ( .A(1'b1), .ZN(_u0_ch21_adr1[24] ) );
INV_X4 _u0_U12615  ( .A(1'b1), .ZN(_u0_ch21_adr1[23] ) );
INV_X4 _u0_U12613  ( .A(1'b1), .ZN(_u0_ch21_adr1[22] ) );
INV_X4 _u0_U12611  ( .A(1'b1), .ZN(_u0_ch21_adr1[21] ) );
INV_X4 _u0_U12609  ( .A(1'b1), .ZN(_u0_ch21_adr1[20] ) );
INV_X4 _u0_U12607  ( .A(1'b1), .ZN(_u0_ch21_adr1[19] ) );
INV_X4 _u0_U12605  ( .A(1'b1), .ZN(_u0_ch21_adr1[18] ) );
INV_X4 _u0_U12603  ( .A(1'b1), .ZN(_u0_ch21_adr1[17] ) );
INV_X4 _u0_U12601  ( .A(1'b1), .ZN(_u0_ch21_adr1[16] ) );
INV_X4 _u0_U12599  ( .A(1'b1), .ZN(_u0_ch21_adr1[15] ) );
INV_X4 _u0_U12597  ( .A(1'b1), .ZN(_u0_ch21_adr1[14] ) );
INV_X4 _u0_U12595  ( .A(1'b1), .ZN(_u0_ch21_adr1[13] ) );
INV_X4 _u0_U12593  ( .A(1'b1), .ZN(_u0_ch21_adr1[12] ) );
INV_X4 _u0_U12591  ( .A(1'b1), .ZN(_u0_ch21_adr1[11] ) );
INV_X4 _u0_U12589  ( .A(1'b1), .ZN(_u0_ch21_adr1[10] ) );
INV_X4 _u0_U12587  ( .A(1'b1), .ZN(_u0_ch21_adr1[9] ) );
INV_X4 _u0_U12585  ( .A(1'b1), .ZN(_u0_ch21_adr1[8] ) );
INV_X4 _u0_U12583  ( .A(1'b1), .ZN(_u0_ch21_adr1[7] ) );
INV_X4 _u0_U12581  ( .A(1'b1), .ZN(_u0_ch21_adr1[6] ) );
INV_X4 _u0_U12579  ( .A(1'b1), .ZN(_u0_ch21_adr1[5] ) );
INV_X4 _u0_U12577  ( .A(1'b1), .ZN(_u0_ch21_adr1[4] ) );
INV_X4 _u0_U12575  ( .A(1'b1), .ZN(_u0_ch21_adr1[3] ) );
INV_X4 _u0_U12573  ( .A(1'b1), .ZN(_u0_ch21_adr1[2] ) );
INV_X4 _u0_U12571  ( .A(1'b1), .ZN(_u0_ch21_adr1[1] ) );
INV_X4 _u0_U12569  ( .A(1'b1), .ZN(_u0_ch21_adr1[0] ) );
INV_X4 _u0_U12567  ( .A(1'b0), .ZN(_u0_ch21_am0[31] ) );
INV_X4 _u0_U12565  ( .A(1'b0), .ZN(_u0_ch21_am0[30] ) );
INV_X4 _u0_U12563  ( .A(1'b0), .ZN(_u0_ch21_am0[29] ) );
INV_X4 _u0_U12561  ( .A(1'b0), .ZN(_u0_ch21_am0[28] ) );
INV_X4 _u0_U12559  ( .A(1'b0), .ZN(_u0_ch21_am0[27] ) );
INV_X4 _u0_U12557  ( .A(1'b0), .ZN(_u0_ch21_am0[26] ) );
INV_X4 _u0_U12555  ( .A(1'b0), .ZN(_u0_ch21_am0[25] ) );
INV_X4 _u0_U12553  ( .A(1'b0), .ZN(_u0_ch21_am0[24] ) );
INV_X4 _u0_U12551  ( .A(1'b0), .ZN(_u0_ch21_am0[23] ) );
INV_X4 _u0_U12549  ( .A(1'b0), .ZN(_u0_ch21_am0[22] ) );
INV_X4 _u0_U12547  ( .A(1'b0), .ZN(_u0_ch21_am0[21] ) );
INV_X4 _u0_U12545  ( .A(1'b0), .ZN(_u0_ch21_am0[20] ) );
INV_X4 _u0_U12543  ( .A(1'b0), .ZN(_u0_ch21_am0[19] ) );
INV_X4 _u0_U12541  ( .A(1'b0), .ZN(_u0_ch21_am0[18] ) );
INV_X4 _u0_U12539  ( .A(1'b0), .ZN(_u0_ch21_am0[17] ) );
INV_X4 _u0_U12537  ( .A(1'b0), .ZN(_u0_ch21_am0[16] ) );
INV_X4 _u0_U12535  ( .A(1'b0), .ZN(_u0_ch21_am0[15] ) );
INV_X4 _u0_U12533  ( .A(1'b0), .ZN(_u0_ch21_am0[14] ) );
INV_X4 _u0_U12531  ( .A(1'b0), .ZN(_u0_ch21_am0[13] ) );
INV_X4 _u0_U12529  ( .A(1'b0), .ZN(_u0_ch21_am0[12] ) );
INV_X4 _u0_U12527  ( .A(1'b0), .ZN(_u0_ch21_am0[11] ) );
INV_X4 _u0_U12525  ( .A(1'b0), .ZN(_u0_ch21_am0[10] ) );
INV_X4 _u0_U12523  ( .A(1'b0), .ZN(_u0_ch21_am0[9] ) );
INV_X4 _u0_U12521  ( .A(1'b0), .ZN(_u0_ch21_am0[8] ) );
INV_X4 _u0_U12519  ( .A(1'b0), .ZN(_u0_ch21_am0[7] ) );
INV_X4 _u0_U12517  ( .A(1'b0), .ZN(_u0_ch21_am0[6] ) );
INV_X4 _u0_U12515  ( .A(1'b0), .ZN(_u0_ch21_am0[5] ) );
INV_X4 _u0_U12513  ( .A(1'b0), .ZN(_u0_ch21_am0[4] ) );
INV_X4 _u0_U12511  ( .A(1'b1), .ZN(_u0_ch21_am0[3] ) );
INV_X4 _u0_U12509  ( .A(1'b1), .ZN(_u0_ch21_am0[2] ) );
INV_X4 _u0_U12507  ( .A(1'b1), .ZN(_u0_ch21_am0[1] ) );
INV_X4 _u0_U12505  ( .A(1'b1), .ZN(_u0_ch21_am0[0] ) );
INV_X4 _u0_U12503  ( .A(1'b0), .ZN(_u0_ch21_am1[31] ) );
INV_X4 _u0_U12501  ( .A(1'b0), .ZN(_u0_ch21_am1[30] ) );
INV_X4 _u0_U12499  ( .A(1'b0), .ZN(_u0_ch21_am1[29] ) );
INV_X4 _u0_U12497  ( .A(1'b0), .ZN(_u0_ch21_am1[28] ) );
INV_X4 _u0_U12495  ( .A(1'b0), .ZN(_u0_ch21_am1[27] ) );
INV_X4 _u0_U12493  ( .A(1'b0), .ZN(_u0_ch21_am1[26] ) );
INV_X4 _u0_U12491  ( .A(1'b0), .ZN(_u0_ch21_am1[25] ) );
INV_X4 _u0_U12489  ( .A(1'b0), .ZN(_u0_ch21_am1[24] ) );
INV_X4 _u0_U12487  ( .A(1'b0), .ZN(_u0_ch21_am1[23] ) );
INV_X4 _u0_U12485  ( .A(1'b0), .ZN(_u0_ch21_am1[22] ) );
INV_X4 _u0_U12483  ( .A(1'b0), .ZN(_u0_ch21_am1[21] ) );
INV_X4 _u0_U12481  ( .A(1'b0), .ZN(_u0_ch21_am1[20] ) );
INV_X4 _u0_U12479  ( .A(1'b0), .ZN(_u0_ch21_am1[19] ) );
INV_X4 _u0_U12477  ( .A(1'b0), .ZN(_u0_ch21_am1[18] ) );
INV_X4 _u0_U12475  ( .A(1'b0), .ZN(_u0_ch21_am1[17] ) );
INV_X4 _u0_U12473  ( .A(1'b0), .ZN(_u0_ch21_am1[16] ) );
INV_X4 _u0_U12471  ( .A(1'b0), .ZN(_u0_ch21_am1[15] ) );
INV_X4 _u0_U12469  ( .A(1'b0), .ZN(_u0_ch21_am1[14] ) );
INV_X4 _u0_U12467  ( .A(1'b0), .ZN(_u0_ch21_am1[13] ) );
INV_X4 _u0_U12465  ( .A(1'b0), .ZN(_u0_ch21_am1[12] ) );
INV_X4 _u0_U12463  ( .A(1'b0), .ZN(_u0_ch21_am1[11] ) );
INV_X4 _u0_U12461  ( .A(1'b0), .ZN(_u0_ch21_am1[10] ) );
INV_X4 _u0_U12459  ( .A(1'b0), .ZN(_u0_ch21_am1[9] ) );
INV_X4 _u0_U12457  ( .A(1'b0), .ZN(_u0_ch21_am1[8] ) );
INV_X4 _u0_U12455  ( .A(1'b0), .ZN(_u0_ch21_am1[7] ) );
INV_X4 _u0_U12453  ( .A(1'b0), .ZN(_u0_ch21_am1[6] ) );
INV_X4 _u0_U12451  ( .A(1'b0), .ZN(_u0_ch21_am1[5] ) );
INV_X4 _u0_U12449  ( .A(1'b0), .ZN(_u0_ch21_am1[4] ) );
INV_X4 _u0_U12447  ( .A(1'b1), .ZN(_u0_ch21_am1[3] ) );
INV_X4 _u0_U12445  ( .A(1'b1), .ZN(_u0_ch21_am1[2] ) );
INV_X4 _u0_U12443  ( .A(1'b1), .ZN(_u0_ch21_am1[1] ) );
INV_X4 _u0_U12441  ( .A(1'b1), .ZN(_u0_ch21_am1[0] ) );
INV_X4 _u0_U12439  ( .A(1'b1), .ZN(_u0_pointer22[31] ) );
INV_X4 _u0_U12437  ( .A(1'b1), .ZN(_u0_pointer22[30] ) );
INV_X4 _u0_U12435  ( .A(1'b1), .ZN(_u0_pointer22[29] ) );
INV_X4 _u0_U12433  ( .A(1'b1), .ZN(_u0_pointer22[28] ) );
INV_X4 _u0_U12431  ( .A(1'b1), .ZN(_u0_pointer22[27] ) );
INV_X4 _u0_U12429  ( .A(1'b1), .ZN(_u0_pointer22[26] ) );
INV_X4 _u0_U12427  ( .A(1'b1), .ZN(_u0_pointer22[25] ) );
INV_X4 _u0_U12425  ( .A(1'b1), .ZN(_u0_pointer22[24] ) );
INV_X4 _u0_U12423  ( .A(1'b1), .ZN(_u0_pointer22[23] ) );
INV_X4 _u0_U12421  ( .A(1'b1), .ZN(_u0_pointer22[22] ) );
INV_X4 _u0_U12419  ( .A(1'b1), .ZN(_u0_pointer22[21] ) );
INV_X4 _u0_U12417  ( .A(1'b1), .ZN(_u0_pointer22[20] ) );
INV_X4 _u0_U12415  ( .A(1'b1), .ZN(_u0_pointer22[19] ) );
INV_X4 _u0_U12413  ( .A(1'b1), .ZN(_u0_pointer22[18] ) );
INV_X4 _u0_U12411  ( .A(1'b1), .ZN(_u0_pointer22[17] ) );
INV_X4 _u0_U12409  ( .A(1'b1), .ZN(_u0_pointer22[16] ) );
INV_X4 _u0_U12407  ( .A(1'b1), .ZN(_u0_pointer22[15] ) );
INV_X4 _u0_U12405  ( .A(1'b1), .ZN(_u0_pointer22[14] ) );
INV_X4 _u0_U12403  ( .A(1'b1), .ZN(_u0_pointer22[13] ) );
INV_X4 _u0_U12401  ( .A(1'b1), .ZN(_u0_pointer22[12] ) );
INV_X4 _u0_U12399  ( .A(1'b1), .ZN(_u0_pointer22[11] ) );
INV_X4 _u0_U12397  ( .A(1'b1), .ZN(_u0_pointer22[10] ) );
INV_X4 _u0_U12395  ( .A(1'b1), .ZN(_u0_pointer22[9] ) );
INV_X4 _u0_U12393  ( .A(1'b1), .ZN(_u0_pointer22[8] ) );
INV_X4 _u0_U12391  ( .A(1'b1), .ZN(_u0_pointer22[7] ) );
INV_X4 _u0_U12389  ( .A(1'b1), .ZN(_u0_pointer22[6] ) );
INV_X4 _u0_U12387  ( .A(1'b1), .ZN(_u0_pointer22[5] ) );
INV_X4 _u0_U12385  ( .A(1'b1), .ZN(_u0_pointer22[4] ) );
INV_X4 _u0_U12383  ( .A(1'b1), .ZN(_u0_pointer22[3] ) );
INV_X4 _u0_U12381  ( .A(1'b1), .ZN(_u0_pointer22[2] ) );
INV_X4 _u0_U12379  ( .A(1'b1), .ZN(_u0_pointer22[1] ) );
INV_X4 _u0_U12377  ( .A(1'b1), .ZN(_u0_pointer22[0] ) );
INV_X4 _u0_U12375  ( .A(1'b1), .ZN(_u0_pointer22_s[31] ) );
INV_X4 _u0_U12373  ( .A(1'b1), .ZN(_u0_pointer22_s[30] ) );
INV_X4 _u0_U12371  ( .A(1'b1), .ZN(_u0_pointer22_s[29] ) );
INV_X4 _u0_U12369  ( .A(1'b1), .ZN(_u0_pointer22_s[28] ) );
INV_X4 _u0_U12367  ( .A(1'b1), .ZN(_u0_pointer22_s[27] ) );
INV_X4 _u0_U12365  ( .A(1'b1), .ZN(_u0_pointer22_s[26] ) );
INV_X4 _u0_U12363  ( .A(1'b1), .ZN(_u0_pointer22_s[25] ) );
INV_X4 _u0_U12361  ( .A(1'b1), .ZN(_u0_pointer22_s[24] ) );
INV_X4 _u0_U12359  ( .A(1'b1), .ZN(_u0_pointer22_s[23] ) );
INV_X4 _u0_U12357  ( .A(1'b1), .ZN(_u0_pointer22_s[22] ) );
INV_X4 _u0_U12355  ( .A(1'b1), .ZN(_u0_pointer22_s[21] ) );
INV_X4 _u0_U12353  ( .A(1'b1), .ZN(_u0_pointer22_s[20] ) );
INV_X4 _u0_U12351  ( .A(1'b1), .ZN(_u0_pointer22_s[19] ) );
INV_X4 _u0_U12349  ( .A(1'b1), .ZN(_u0_pointer22_s[18] ) );
INV_X4 _u0_U12347  ( .A(1'b1), .ZN(_u0_pointer22_s[17] ) );
INV_X4 _u0_U12345  ( .A(1'b1), .ZN(_u0_pointer22_s[16] ) );
INV_X4 _u0_U12343  ( .A(1'b1), .ZN(_u0_pointer22_s[15] ) );
INV_X4 _u0_U12341  ( .A(1'b1), .ZN(_u0_pointer22_s[14] ) );
INV_X4 _u0_U12339  ( .A(1'b1), .ZN(_u0_pointer22_s[13] ) );
INV_X4 _u0_U12337  ( .A(1'b1), .ZN(_u0_pointer22_s[12] ) );
INV_X4 _u0_U12335  ( .A(1'b1), .ZN(_u0_pointer22_s[11] ) );
INV_X4 _u0_U12333  ( .A(1'b1), .ZN(_u0_pointer22_s[10] ) );
INV_X4 _u0_U12331  ( .A(1'b1), .ZN(_u0_pointer22_s[9] ) );
INV_X4 _u0_U12329  ( .A(1'b1), .ZN(_u0_pointer22_s[8] ) );
INV_X4 _u0_U12327  ( .A(1'b1), .ZN(_u0_pointer22_s[7] ) );
INV_X4 _u0_U12325  ( .A(1'b1), .ZN(_u0_pointer22_s[6] ) );
INV_X4 _u0_U12323  ( .A(1'b1), .ZN(_u0_pointer22_s[5] ) );
INV_X4 _u0_U12321  ( .A(1'b1), .ZN(_u0_pointer22_s[4] ) );
INV_X4 _u0_U12319  ( .A(1'b1), .ZN(_u0_pointer22_s[3] ) );
INV_X4 _u0_U12317  ( .A(1'b1), .ZN(_u0_pointer22_s[2] ) );
INV_X4 _u0_U12315  ( .A(1'b1), .ZN(_u0_pointer22_s[1] ) );
INV_X4 _u0_U12313  ( .A(1'b1), .ZN(_u0_pointer22_s[0] ) );
INV_X4 _u0_U12311  ( .A(1'b1), .ZN(_u0_ch22_csr[31] ) );
INV_X4 _u0_U12309  ( .A(1'b1), .ZN(_u0_ch22_csr[30] ) );
INV_X4 _u0_U12307  ( .A(1'b1), .ZN(_u0_ch22_csr[29] ) );
INV_X4 _u0_U12305  ( .A(1'b1), .ZN(_u0_ch22_csr[28] ) );
INV_X4 _u0_U12303  ( .A(1'b1), .ZN(_u0_ch22_csr[27] ) );
INV_X4 _u0_U12301  ( .A(1'b1), .ZN(_u0_ch22_csr[26] ) );
INV_X4 _u0_U12299  ( .A(1'b1), .ZN(_u0_ch22_csr[25] ) );
INV_X4 _u0_U12297  ( .A(1'b1), .ZN(_u0_ch22_csr[24] ) );
INV_X4 _u0_U12295  ( .A(1'b1), .ZN(_u0_ch22_csr[23] ) );
INV_X4 _u0_U12293  ( .A(1'b1), .ZN(_u0_ch22_csr[22] ) );
INV_X4 _u0_U12291  ( .A(1'b1), .ZN(_u0_ch22_csr[21] ) );
INV_X4 _u0_U12289  ( .A(1'b1), .ZN(_u0_ch22_csr[20] ) );
INV_X4 _u0_U12287  ( .A(1'b1), .ZN(_u0_ch22_csr[19] ) );
INV_X4 _u0_U12285  ( .A(1'b1), .ZN(_u0_ch22_csr[18] ) );
INV_X4 _u0_U12283  ( .A(1'b1), .ZN(_u0_ch22_csr[17] ) );
INV_X4 _u0_U12281  ( .A(1'b1), .ZN(_u0_ch22_csr[16] ) );
INV_X4 _u0_U12279  ( .A(1'b1), .ZN(_u0_ch22_csr[15] ) );
INV_X4 _u0_U12277  ( .A(1'b1), .ZN(_u0_ch22_csr[14] ) );
INV_X4 _u0_U12275  ( .A(1'b1), .ZN(_u0_ch22_csr[13] ) );
INV_X4 _u0_U12273  ( .A(1'b1), .ZN(_u0_ch22_csr[12] ) );
INV_X4 _u0_U12271  ( .A(1'b1), .ZN(_u0_ch22_csr[11] ) );
INV_X4 _u0_U12269  ( .A(1'b1), .ZN(_u0_ch22_csr[10] ) );
INV_X4 _u0_U12267  ( .A(1'b1), .ZN(_u0_ch22_csr[9] ) );
INV_X4 _u0_U12265  ( .A(1'b1), .ZN(_u0_ch22_csr[8] ) );
INV_X4 _u0_U12263  ( .A(1'b1), .ZN(_u0_ch22_csr[7] ) );
INV_X4 _u0_U12261  ( .A(1'b1), .ZN(_u0_ch22_csr[6] ) );
INV_X4 _u0_U12259  ( .A(1'b1), .ZN(_u0_ch22_csr[5] ) );
INV_X4 _u0_U12257  ( .A(1'b1), .ZN(_u0_ch22_csr[4] ) );
INV_X4 _u0_U12255  ( .A(1'b1), .ZN(_u0_ch22_csr[3] ) );
INV_X4 _u0_U12253  ( .A(1'b1), .ZN(_u0_ch22_csr[2] ) );
INV_X4 _u0_U12251  ( .A(1'b1), .ZN(_u0_ch22_csr[1] ) );
INV_X4 _u0_U12249  ( .A(1'b1), .ZN(_u0_ch22_csr[0] ) );
INV_X4 _u0_U12247  ( .A(1'b1), .ZN(_u0_ch22_txsz[31] ) );
INV_X4 _u0_U12245  ( .A(1'b1), .ZN(_u0_ch22_txsz[30] ) );
INV_X4 _u0_U12243  ( .A(1'b1), .ZN(_u0_ch22_txsz[29] ) );
INV_X4 _u0_U12241  ( .A(1'b1), .ZN(_u0_ch22_txsz[28] ) );
INV_X4 _u0_U12239  ( .A(1'b1), .ZN(_u0_ch22_txsz[27] ) );
INV_X4 _u0_U12237  ( .A(1'b1), .ZN(_u0_ch22_txsz[26] ) );
INV_X4 _u0_U12235  ( .A(1'b1), .ZN(_u0_ch22_txsz[25] ) );
INV_X4 _u0_U12233  ( .A(1'b1), .ZN(_u0_ch22_txsz[24] ) );
INV_X4 _u0_U12231  ( .A(1'b1), .ZN(_u0_ch22_txsz[23] ) );
INV_X4 _u0_U12229  ( .A(1'b1), .ZN(_u0_ch22_txsz[22] ) );
INV_X4 _u0_U12227  ( .A(1'b1), .ZN(_u0_ch22_txsz[21] ) );
INV_X4 _u0_U12225  ( .A(1'b1), .ZN(_u0_ch22_txsz[20] ) );
INV_X4 _u0_U12223  ( .A(1'b1), .ZN(_u0_ch22_txsz[19] ) );
INV_X4 _u0_U12221  ( .A(1'b1), .ZN(_u0_ch22_txsz[18] ) );
INV_X4 _u0_U12219  ( .A(1'b1), .ZN(_u0_ch22_txsz[17] ) );
INV_X4 _u0_U12217  ( .A(1'b1), .ZN(_u0_ch22_txsz[16] ) );
INV_X4 _u0_U12215  ( .A(1'b1), .ZN(_u0_ch22_txsz[15] ) );
INV_X4 _u0_U12213  ( .A(1'b1), .ZN(_u0_ch22_txsz[14] ) );
INV_X4 _u0_U12211  ( .A(1'b1), .ZN(_u0_ch22_txsz[13] ) );
INV_X4 _u0_U12209  ( .A(1'b1), .ZN(_u0_ch22_txsz[12] ) );
INV_X4 _u0_U12207  ( .A(1'b1), .ZN(_u0_ch22_txsz[11] ) );
INV_X4 _u0_U12205  ( .A(1'b1), .ZN(_u0_ch22_txsz[10] ) );
INV_X4 _u0_U12203  ( .A(1'b1), .ZN(_u0_ch22_txsz[9] ) );
INV_X4 _u0_U12201  ( .A(1'b1), .ZN(_u0_ch22_txsz[8] ) );
INV_X4 _u0_U12199  ( .A(1'b1), .ZN(_u0_ch22_txsz[7] ) );
INV_X4 _u0_U12197  ( .A(1'b1), .ZN(_u0_ch22_txsz[6] ) );
INV_X4 _u0_U12195  ( .A(1'b1), .ZN(_u0_ch22_txsz[5] ) );
INV_X4 _u0_U12193  ( .A(1'b1), .ZN(_u0_ch22_txsz[4] ) );
INV_X4 _u0_U12191  ( .A(1'b1), .ZN(_u0_ch22_txsz[3] ) );
INV_X4 _u0_U12189  ( .A(1'b1), .ZN(_u0_ch22_txsz[2] ) );
INV_X4 _u0_U12187  ( .A(1'b1), .ZN(_u0_ch22_txsz[1] ) );
INV_X4 _u0_U12185  ( .A(1'b1), .ZN(_u0_ch22_txsz[0] ) );
INV_X4 _u0_U12183  ( .A(1'b1), .ZN(_u0_ch22_adr0[31] ) );
INV_X4 _u0_U12181  ( .A(1'b1), .ZN(_u0_ch22_adr0[30] ) );
INV_X4 _u0_U12179  ( .A(1'b1), .ZN(_u0_ch22_adr0[29] ) );
INV_X4 _u0_U12177  ( .A(1'b1), .ZN(_u0_ch22_adr0[28] ) );
INV_X4 _u0_U12175  ( .A(1'b1), .ZN(_u0_ch22_adr0[27] ) );
INV_X4 _u0_U12173  ( .A(1'b1), .ZN(_u0_ch22_adr0[26] ) );
INV_X4 _u0_U12171  ( .A(1'b1), .ZN(_u0_ch22_adr0[25] ) );
INV_X4 _u0_U12169  ( .A(1'b1), .ZN(_u0_ch22_adr0[24] ) );
INV_X4 _u0_U12167  ( .A(1'b1), .ZN(_u0_ch22_adr0[23] ) );
INV_X4 _u0_U12165  ( .A(1'b1), .ZN(_u0_ch22_adr0[22] ) );
INV_X4 _u0_U12163  ( .A(1'b1), .ZN(_u0_ch22_adr0[21] ) );
INV_X4 _u0_U12161  ( .A(1'b1), .ZN(_u0_ch22_adr0[20] ) );
INV_X4 _u0_U12159  ( .A(1'b1), .ZN(_u0_ch22_adr0[19] ) );
INV_X4 _u0_U12157  ( .A(1'b1), .ZN(_u0_ch22_adr0[18] ) );
INV_X4 _u0_U12155  ( .A(1'b1), .ZN(_u0_ch22_adr0[17] ) );
INV_X4 _u0_U12153  ( .A(1'b1), .ZN(_u0_ch22_adr0[16] ) );
INV_X4 _u0_U12151  ( .A(1'b1), .ZN(_u0_ch22_adr0[15] ) );
INV_X4 _u0_U12149  ( .A(1'b1), .ZN(_u0_ch22_adr0[14] ) );
INV_X4 _u0_U12147  ( .A(1'b1), .ZN(_u0_ch22_adr0[13] ) );
INV_X4 _u0_U12145  ( .A(1'b1), .ZN(_u0_ch22_adr0[12] ) );
INV_X4 _u0_U12143  ( .A(1'b1), .ZN(_u0_ch22_adr0[11] ) );
INV_X4 _u0_U12141  ( .A(1'b1), .ZN(_u0_ch22_adr0[10] ) );
INV_X4 _u0_U12139  ( .A(1'b1), .ZN(_u0_ch22_adr0[9] ) );
INV_X4 _u0_U12137  ( .A(1'b1), .ZN(_u0_ch22_adr0[8] ) );
INV_X4 _u0_U12135  ( .A(1'b1), .ZN(_u0_ch22_adr0[7] ) );
INV_X4 _u0_U12133  ( .A(1'b1), .ZN(_u0_ch22_adr0[6] ) );
INV_X4 _u0_U12131  ( .A(1'b1), .ZN(_u0_ch22_adr0[5] ) );
INV_X4 _u0_U12129  ( .A(1'b1), .ZN(_u0_ch22_adr0[4] ) );
INV_X4 _u0_U12127  ( .A(1'b1), .ZN(_u0_ch22_adr0[3] ) );
INV_X4 _u0_U12125  ( .A(1'b1), .ZN(_u0_ch22_adr0[2] ) );
INV_X4 _u0_U12123  ( .A(1'b1), .ZN(_u0_ch22_adr0[1] ) );
INV_X4 _u0_U12121  ( .A(1'b1), .ZN(_u0_ch22_adr0[0] ) );
INV_X4 _u0_U12119  ( .A(1'b1), .ZN(_u0_ch22_adr1[31] ) );
INV_X4 _u0_U12117  ( .A(1'b1), .ZN(_u0_ch22_adr1[30] ) );
INV_X4 _u0_U12115  ( .A(1'b1), .ZN(_u0_ch22_adr1[29] ) );
INV_X4 _u0_U12113  ( .A(1'b1), .ZN(_u0_ch22_adr1[28] ) );
INV_X4 _u0_U12111  ( .A(1'b1), .ZN(_u0_ch22_adr1[27] ) );
INV_X4 _u0_U12109  ( .A(1'b1), .ZN(_u0_ch22_adr1[26] ) );
INV_X4 _u0_U12107  ( .A(1'b1), .ZN(_u0_ch22_adr1[25] ) );
INV_X4 _u0_U12105  ( .A(1'b1), .ZN(_u0_ch22_adr1[24] ) );
INV_X4 _u0_U12103  ( .A(1'b1), .ZN(_u0_ch22_adr1[23] ) );
INV_X4 _u0_U12101  ( .A(1'b1), .ZN(_u0_ch22_adr1[22] ) );
INV_X4 _u0_U12099  ( .A(1'b1), .ZN(_u0_ch22_adr1[21] ) );
INV_X4 _u0_U12097  ( .A(1'b1), .ZN(_u0_ch22_adr1[20] ) );
INV_X4 _u0_U12095  ( .A(1'b1), .ZN(_u0_ch22_adr1[19] ) );
INV_X4 _u0_U12093  ( .A(1'b1), .ZN(_u0_ch22_adr1[18] ) );
INV_X4 _u0_U12091  ( .A(1'b1), .ZN(_u0_ch22_adr1[17] ) );
INV_X4 _u0_U12089  ( .A(1'b1), .ZN(_u0_ch22_adr1[16] ) );
INV_X4 _u0_U12087  ( .A(1'b1), .ZN(_u0_ch22_adr1[15] ) );
INV_X4 _u0_U12085  ( .A(1'b1), .ZN(_u0_ch22_adr1[14] ) );
INV_X4 _u0_U12083  ( .A(1'b1), .ZN(_u0_ch22_adr1[13] ) );
INV_X4 _u0_U12081  ( .A(1'b1), .ZN(_u0_ch22_adr1[12] ) );
INV_X4 _u0_U12079  ( .A(1'b1), .ZN(_u0_ch22_adr1[11] ) );
INV_X4 _u0_U12077  ( .A(1'b1), .ZN(_u0_ch22_adr1[10] ) );
INV_X4 _u0_U12075  ( .A(1'b1), .ZN(_u0_ch22_adr1[9] ) );
INV_X4 _u0_U12073  ( .A(1'b1), .ZN(_u0_ch22_adr1[8] ) );
INV_X4 _u0_U12071  ( .A(1'b1), .ZN(_u0_ch22_adr1[7] ) );
INV_X4 _u0_U12069  ( .A(1'b1), .ZN(_u0_ch22_adr1[6] ) );
INV_X4 _u0_U12067  ( .A(1'b1), .ZN(_u0_ch22_adr1[5] ) );
INV_X4 _u0_U12065  ( .A(1'b1), .ZN(_u0_ch22_adr1[4] ) );
INV_X4 _u0_U12063  ( .A(1'b1), .ZN(_u0_ch22_adr1[3] ) );
INV_X4 _u0_U12061  ( .A(1'b1), .ZN(_u0_ch22_adr1[2] ) );
INV_X4 _u0_U12059  ( .A(1'b1), .ZN(_u0_ch22_adr1[1] ) );
INV_X4 _u0_U12057  ( .A(1'b1), .ZN(_u0_ch22_adr1[0] ) );
INV_X4 _u0_U12055  ( .A(1'b0), .ZN(_u0_ch22_am0[31] ) );
INV_X4 _u0_U12053  ( .A(1'b0), .ZN(_u0_ch22_am0[30] ) );
INV_X4 _u0_U12051  ( .A(1'b0), .ZN(_u0_ch22_am0[29] ) );
INV_X4 _u0_U12049  ( .A(1'b0), .ZN(_u0_ch22_am0[28] ) );
INV_X4 _u0_U12047  ( .A(1'b0), .ZN(_u0_ch22_am0[27] ) );
INV_X4 _u0_U12045  ( .A(1'b0), .ZN(_u0_ch22_am0[26] ) );
INV_X4 _u0_U12043  ( .A(1'b0), .ZN(_u0_ch22_am0[25] ) );
INV_X4 _u0_U12041  ( .A(1'b0), .ZN(_u0_ch22_am0[24] ) );
INV_X4 _u0_U12039  ( .A(1'b0), .ZN(_u0_ch22_am0[23] ) );
INV_X4 _u0_U12037  ( .A(1'b0), .ZN(_u0_ch22_am0[22] ) );
INV_X4 _u0_U12035  ( .A(1'b0), .ZN(_u0_ch22_am0[21] ) );
INV_X4 _u0_U12033  ( .A(1'b0), .ZN(_u0_ch22_am0[20] ) );
INV_X4 _u0_U12031  ( .A(1'b0), .ZN(_u0_ch22_am0[19] ) );
INV_X4 _u0_U12029  ( .A(1'b0), .ZN(_u0_ch22_am0[18] ) );
INV_X4 _u0_U12027  ( .A(1'b0), .ZN(_u0_ch22_am0[17] ) );
INV_X4 _u0_U12025  ( .A(1'b0), .ZN(_u0_ch22_am0[16] ) );
INV_X4 _u0_U12023  ( .A(1'b0), .ZN(_u0_ch22_am0[15] ) );
INV_X4 _u0_U12021  ( .A(1'b0), .ZN(_u0_ch22_am0[14] ) );
INV_X4 _u0_U12019  ( .A(1'b0), .ZN(_u0_ch22_am0[13] ) );
INV_X4 _u0_U12017  ( .A(1'b0), .ZN(_u0_ch22_am0[12] ) );
INV_X4 _u0_U12015  ( .A(1'b0), .ZN(_u0_ch22_am0[11] ) );
INV_X4 _u0_U12013  ( .A(1'b0), .ZN(_u0_ch22_am0[10] ) );
INV_X4 _u0_U12011  ( .A(1'b0), .ZN(_u0_ch22_am0[9] ) );
INV_X4 _u0_U12009  ( .A(1'b0), .ZN(_u0_ch22_am0[8] ) );
INV_X4 _u0_U12007  ( .A(1'b0), .ZN(_u0_ch22_am0[7] ) );
INV_X4 _u0_U12005  ( .A(1'b0), .ZN(_u0_ch22_am0[6] ) );
INV_X4 _u0_U12003  ( .A(1'b0), .ZN(_u0_ch22_am0[5] ) );
INV_X4 _u0_U12001  ( .A(1'b0), .ZN(_u0_ch22_am0[4] ) );
INV_X4 _u0_U11999  ( .A(1'b1), .ZN(_u0_ch22_am0[3] ) );
INV_X4 _u0_U11997  ( .A(1'b1), .ZN(_u0_ch22_am0[2] ) );
INV_X4 _u0_U11995  ( .A(1'b1), .ZN(_u0_ch22_am0[1] ) );
INV_X4 _u0_U11993  ( .A(1'b1), .ZN(_u0_ch22_am0[0] ) );
INV_X4 _u0_U11991  ( .A(1'b0), .ZN(_u0_ch22_am1[31] ) );
INV_X4 _u0_U11989  ( .A(1'b0), .ZN(_u0_ch22_am1[30] ) );
INV_X4 _u0_U11987  ( .A(1'b0), .ZN(_u0_ch22_am1[29] ) );
INV_X4 _u0_U11985  ( .A(1'b0), .ZN(_u0_ch22_am1[28] ) );
INV_X4 _u0_U11983  ( .A(1'b0), .ZN(_u0_ch22_am1[27] ) );
INV_X4 _u0_U11981  ( .A(1'b0), .ZN(_u0_ch22_am1[26] ) );
INV_X4 _u0_U11979  ( .A(1'b0), .ZN(_u0_ch22_am1[25] ) );
INV_X4 _u0_U11977  ( .A(1'b0), .ZN(_u0_ch22_am1[24] ) );
INV_X4 _u0_U11975  ( .A(1'b0), .ZN(_u0_ch22_am1[23] ) );
INV_X4 _u0_U11973  ( .A(1'b0), .ZN(_u0_ch22_am1[22] ) );
INV_X4 _u0_U11971  ( .A(1'b0), .ZN(_u0_ch22_am1[21] ) );
INV_X4 _u0_U11969  ( .A(1'b0), .ZN(_u0_ch22_am1[20] ) );
INV_X4 _u0_U11967  ( .A(1'b0), .ZN(_u0_ch22_am1[19] ) );
INV_X4 _u0_U11965  ( .A(1'b0), .ZN(_u0_ch22_am1[18] ) );
INV_X4 _u0_U11963  ( .A(1'b0), .ZN(_u0_ch22_am1[17] ) );
INV_X4 _u0_U11961  ( .A(1'b0), .ZN(_u0_ch22_am1[16] ) );
INV_X4 _u0_U11959  ( .A(1'b0), .ZN(_u0_ch22_am1[15] ) );
INV_X4 _u0_U11957  ( .A(1'b0), .ZN(_u0_ch22_am1[14] ) );
INV_X4 _u0_U11955  ( .A(1'b0), .ZN(_u0_ch22_am1[13] ) );
INV_X4 _u0_U11953  ( .A(1'b0), .ZN(_u0_ch22_am1[12] ) );
INV_X4 _u0_U11951  ( .A(1'b0), .ZN(_u0_ch22_am1[11] ) );
INV_X4 _u0_U11949  ( .A(1'b0), .ZN(_u0_ch22_am1[10] ) );
INV_X4 _u0_U11947  ( .A(1'b0), .ZN(_u0_ch22_am1[9] ) );
INV_X4 _u0_U11945  ( .A(1'b0), .ZN(_u0_ch22_am1[8] ) );
INV_X4 _u0_U11943  ( .A(1'b0), .ZN(_u0_ch22_am1[7] ) );
INV_X4 _u0_U11941  ( .A(1'b0), .ZN(_u0_ch22_am1[6] ) );
INV_X4 _u0_U11939  ( .A(1'b0), .ZN(_u0_ch22_am1[5] ) );
INV_X4 _u0_U11937  ( .A(1'b0), .ZN(_u0_ch22_am1[4] ) );
INV_X4 _u0_U11935  ( .A(1'b1), .ZN(_u0_ch22_am1[3] ) );
INV_X4 _u0_U11933  ( .A(1'b1), .ZN(_u0_ch22_am1[2] ) );
INV_X4 _u0_U11931  ( .A(1'b1), .ZN(_u0_ch22_am1[1] ) );
INV_X4 _u0_U11929  ( .A(1'b1), .ZN(_u0_ch22_am1[0] ) );
INV_X4 _u0_U11927  ( .A(1'b1), .ZN(_u0_pointer23[31] ) );
INV_X4 _u0_U11925  ( .A(1'b1), .ZN(_u0_pointer23[30] ) );
INV_X4 _u0_U11923  ( .A(1'b1), .ZN(_u0_pointer23[29] ) );
INV_X4 _u0_U11921  ( .A(1'b1), .ZN(_u0_pointer23[28] ) );
INV_X4 _u0_U11919  ( .A(1'b1), .ZN(_u0_pointer23[27] ) );
INV_X4 _u0_U11917  ( .A(1'b1), .ZN(_u0_pointer23[26] ) );
INV_X4 _u0_U11915  ( .A(1'b1), .ZN(_u0_pointer23[25] ) );
INV_X4 _u0_U11913  ( .A(1'b1), .ZN(_u0_pointer23[24] ) );
INV_X4 _u0_U11911  ( .A(1'b1), .ZN(_u0_pointer23[23] ) );
INV_X4 _u0_U11909  ( .A(1'b1), .ZN(_u0_pointer23[22] ) );
INV_X4 _u0_U11907  ( .A(1'b1), .ZN(_u0_pointer23[21] ) );
INV_X4 _u0_U11905  ( .A(1'b1), .ZN(_u0_pointer23[20] ) );
INV_X4 _u0_U11903  ( .A(1'b1), .ZN(_u0_pointer23[19] ) );
INV_X4 _u0_U11901  ( .A(1'b1), .ZN(_u0_pointer23[18] ) );
INV_X4 _u0_U11899  ( .A(1'b1), .ZN(_u0_pointer23[17] ) );
INV_X4 _u0_U11897  ( .A(1'b1), .ZN(_u0_pointer23[16] ) );
INV_X4 _u0_U11895  ( .A(1'b1), .ZN(_u0_pointer23[15] ) );
INV_X4 _u0_U11893  ( .A(1'b1), .ZN(_u0_pointer23[14] ) );
INV_X4 _u0_U11891  ( .A(1'b1), .ZN(_u0_pointer23[13] ) );
INV_X4 _u0_U11889  ( .A(1'b1), .ZN(_u0_pointer23[12] ) );
INV_X4 _u0_U11887  ( .A(1'b1), .ZN(_u0_pointer23[11] ) );
INV_X4 _u0_U11885  ( .A(1'b1), .ZN(_u0_pointer23[10] ) );
INV_X4 _u0_U11883  ( .A(1'b1), .ZN(_u0_pointer23[9] ) );
INV_X4 _u0_U11881  ( .A(1'b1), .ZN(_u0_pointer23[8] ) );
INV_X4 _u0_U11879  ( .A(1'b1), .ZN(_u0_pointer23[7] ) );
INV_X4 _u0_U11877  ( .A(1'b1), .ZN(_u0_pointer23[6] ) );
INV_X4 _u0_U11875  ( .A(1'b1), .ZN(_u0_pointer23[5] ) );
INV_X4 _u0_U11873  ( .A(1'b1), .ZN(_u0_pointer23[4] ) );
INV_X4 _u0_U11871  ( .A(1'b1), .ZN(_u0_pointer23[3] ) );
INV_X4 _u0_U11869  ( .A(1'b1), .ZN(_u0_pointer23[2] ) );
INV_X4 _u0_U11867  ( .A(1'b1), .ZN(_u0_pointer23[1] ) );
INV_X4 _u0_U11865  ( .A(1'b1), .ZN(_u0_pointer23[0] ) );
INV_X4 _u0_U11863  ( .A(1'b1), .ZN(_u0_pointer23_s[31] ) );
INV_X4 _u0_U11861  ( .A(1'b1), .ZN(_u0_pointer23_s[30] ) );
INV_X4 _u0_U11859  ( .A(1'b1), .ZN(_u0_pointer23_s[29] ) );
INV_X4 _u0_U11857  ( .A(1'b1), .ZN(_u0_pointer23_s[28] ) );
INV_X4 _u0_U11855  ( .A(1'b1), .ZN(_u0_pointer23_s[27] ) );
INV_X4 _u0_U11853  ( .A(1'b1), .ZN(_u0_pointer23_s[26] ) );
INV_X4 _u0_U11851  ( .A(1'b1), .ZN(_u0_pointer23_s[25] ) );
INV_X4 _u0_U11849  ( .A(1'b1), .ZN(_u0_pointer23_s[24] ) );
INV_X4 _u0_U11847  ( .A(1'b1), .ZN(_u0_pointer23_s[23] ) );
INV_X4 _u0_U11845  ( .A(1'b1), .ZN(_u0_pointer23_s[22] ) );
INV_X4 _u0_U11843  ( .A(1'b1), .ZN(_u0_pointer23_s[21] ) );
INV_X4 _u0_U11841  ( .A(1'b1), .ZN(_u0_pointer23_s[20] ) );
INV_X4 _u0_U11839  ( .A(1'b1), .ZN(_u0_pointer23_s[19] ) );
INV_X4 _u0_U11837  ( .A(1'b1), .ZN(_u0_pointer23_s[18] ) );
INV_X4 _u0_U11835  ( .A(1'b1), .ZN(_u0_pointer23_s[17] ) );
INV_X4 _u0_U11833  ( .A(1'b1), .ZN(_u0_pointer23_s[16] ) );
INV_X4 _u0_U11831  ( .A(1'b1), .ZN(_u0_pointer23_s[15] ) );
INV_X4 _u0_U11829  ( .A(1'b1), .ZN(_u0_pointer23_s[14] ) );
INV_X4 _u0_U11827  ( .A(1'b1), .ZN(_u0_pointer23_s[13] ) );
INV_X4 _u0_U11825  ( .A(1'b1), .ZN(_u0_pointer23_s[12] ) );
INV_X4 _u0_U11823  ( .A(1'b1), .ZN(_u0_pointer23_s[11] ) );
INV_X4 _u0_U11821  ( .A(1'b1), .ZN(_u0_pointer23_s[10] ) );
INV_X4 _u0_U11819  ( .A(1'b1), .ZN(_u0_pointer23_s[9] ) );
INV_X4 _u0_U11817  ( .A(1'b1), .ZN(_u0_pointer23_s[8] ) );
INV_X4 _u0_U11815  ( .A(1'b1), .ZN(_u0_pointer23_s[7] ) );
INV_X4 _u0_U11813  ( .A(1'b1), .ZN(_u0_pointer23_s[6] ) );
INV_X4 _u0_U11811  ( .A(1'b1), .ZN(_u0_pointer23_s[5] ) );
INV_X4 _u0_U11809  ( .A(1'b1), .ZN(_u0_pointer23_s[4] ) );
INV_X4 _u0_U11807  ( .A(1'b1), .ZN(_u0_pointer23_s[3] ) );
INV_X4 _u0_U11805  ( .A(1'b1), .ZN(_u0_pointer23_s[2] ) );
INV_X4 _u0_U11803  ( .A(1'b1), .ZN(_u0_pointer23_s[1] ) );
INV_X4 _u0_U11801  ( .A(1'b1), .ZN(_u0_pointer23_s[0] ) );
INV_X4 _u0_U11799  ( .A(1'b1), .ZN(_u0_ch23_csr[31] ) );
INV_X4 _u0_U11797  ( .A(1'b1), .ZN(_u0_ch23_csr[30] ) );
INV_X4 _u0_U11795  ( .A(1'b1), .ZN(_u0_ch23_csr[29] ) );
INV_X4 _u0_U11793  ( .A(1'b1), .ZN(_u0_ch23_csr[28] ) );
INV_X4 _u0_U11791  ( .A(1'b1), .ZN(_u0_ch23_csr[27] ) );
INV_X4 _u0_U11789  ( .A(1'b1), .ZN(_u0_ch23_csr[26] ) );
INV_X4 _u0_U11787  ( .A(1'b1), .ZN(_u0_ch23_csr[25] ) );
INV_X4 _u0_U11785  ( .A(1'b1), .ZN(_u0_ch23_csr[24] ) );
INV_X4 _u0_U11783  ( .A(1'b1), .ZN(_u0_ch23_csr[23] ) );
INV_X4 _u0_U11781  ( .A(1'b1), .ZN(_u0_ch23_csr[22] ) );
INV_X4 _u0_U11779  ( .A(1'b1), .ZN(_u0_ch23_csr[21] ) );
INV_X4 _u0_U11777  ( .A(1'b1), .ZN(_u0_ch23_csr[20] ) );
INV_X4 _u0_U11775  ( .A(1'b1), .ZN(_u0_ch23_csr[19] ) );
INV_X4 _u0_U11773  ( .A(1'b1), .ZN(_u0_ch23_csr[18] ) );
INV_X4 _u0_U11771  ( .A(1'b1), .ZN(_u0_ch23_csr[17] ) );
INV_X4 _u0_U11769  ( .A(1'b1), .ZN(_u0_ch23_csr[16] ) );
INV_X4 _u0_U11767  ( .A(1'b1), .ZN(_u0_ch23_csr[15] ) );
INV_X4 _u0_U11765  ( .A(1'b1), .ZN(_u0_ch23_csr[14] ) );
INV_X4 _u0_U11763  ( .A(1'b1), .ZN(_u0_ch23_csr[13] ) );
INV_X4 _u0_U11761  ( .A(1'b1), .ZN(_u0_ch23_csr[12] ) );
INV_X4 _u0_U11759  ( .A(1'b1), .ZN(_u0_ch23_csr[11] ) );
INV_X4 _u0_U11757  ( .A(1'b1), .ZN(_u0_ch23_csr[10] ) );
INV_X4 _u0_U11755  ( .A(1'b1), .ZN(_u0_ch23_csr[9] ) );
INV_X4 _u0_U11753  ( .A(1'b1), .ZN(_u0_ch23_csr[8] ) );
INV_X4 _u0_U11751  ( .A(1'b1), .ZN(_u0_ch23_csr[7] ) );
INV_X4 _u0_U11749  ( .A(1'b1), .ZN(_u0_ch23_csr[6] ) );
INV_X4 _u0_U11747  ( .A(1'b1), .ZN(_u0_ch23_csr[5] ) );
INV_X4 _u0_U11745  ( .A(1'b1), .ZN(_u0_ch23_csr[4] ) );
INV_X4 _u0_U11743  ( .A(1'b1), .ZN(_u0_ch23_csr[3] ) );
INV_X4 _u0_U11741  ( .A(1'b1), .ZN(_u0_ch23_csr[2] ) );
INV_X4 _u0_U11739  ( .A(1'b1), .ZN(_u0_ch23_csr[1] ) );
INV_X4 _u0_U11737  ( .A(1'b1), .ZN(_u0_ch23_csr[0] ) );
INV_X4 _u0_U11735  ( .A(1'b1), .ZN(_u0_ch23_txsz[31] ) );
INV_X4 _u0_U11733  ( .A(1'b1), .ZN(_u0_ch23_txsz[30] ) );
INV_X4 _u0_U11731  ( .A(1'b1), .ZN(_u0_ch23_txsz[29] ) );
INV_X4 _u0_U11729  ( .A(1'b1), .ZN(_u0_ch23_txsz[28] ) );
INV_X4 _u0_U11727  ( .A(1'b1), .ZN(_u0_ch23_txsz[27] ) );
INV_X4 _u0_U11725  ( .A(1'b1), .ZN(_u0_ch23_txsz[26] ) );
INV_X4 _u0_U11723  ( .A(1'b1), .ZN(_u0_ch23_txsz[25] ) );
INV_X4 _u0_U11721  ( .A(1'b1), .ZN(_u0_ch23_txsz[24] ) );
INV_X4 _u0_U11719  ( .A(1'b1), .ZN(_u0_ch23_txsz[23] ) );
INV_X4 _u0_U11717  ( .A(1'b1), .ZN(_u0_ch23_txsz[22] ) );
INV_X4 _u0_U11715  ( .A(1'b1), .ZN(_u0_ch23_txsz[21] ) );
INV_X4 _u0_U11713  ( .A(1'b1), .ZN(_u0_ch23_txsz[20] ) );
INV_X4 _u0_U11711  ( .A(1'b1), .ZN(_u0_ch23_txsz[19] ) );
INV_X4 _u0_U11709  ( .A(1'b1), .ZN(_u0_ch23_txsz[18] ) );
INV_X4 _u0_U11707  ( .A(1'b1), .ZN(_u0_ch23_txsz[17] ) );
INV_X4 _u0_U11705  ( .A(1'b1), .ZN(_u0_ch23_txsz[16] ) );
INV_X4 _u0_U11703  ( .A(1'b1), .ZN(_u0_ch23_txsz[15] ) );
INV_X4 _u0_U11701  ( .A(1'b1), .ZN(_u0_ch23_txsz[14] ) );
INV_X4 _u0_U11699  ( .A(1'b1), .ZN(_u0_ch23_txsz[13] ) );
INV_X4 _u0_U11697  ( .A(1'b1), .ZN(_u0_ch23_txsz[12] ) );
INV_X4 _u0_U11695  ( .A(1'b1), .ZN(_u0_ch23_txsz[11] ) );
INV_X4 _u0_U11693  ( .A(1'b1), .ZN(_u0_ch23_txsz[10] ) );
INV_X4 _u0_U11691  ( .A(1'b1), .ZN(_u0_ch23_txsz[9] ) );
INV_X4 _u0_U11689  ( .A(1'b1), .ZN(_u0_ch23_txsz[8] ) );
INV_X4 _u0_U11687  ( .A(1'b1), .ZN(_u0_ch23_txsz[7] ) );
INV_X4 _u0_U11685  ( .A(1'b1), .ZN(_u0_ch23_txsz[6] ) );
INV_X4 _u0_U11683  ( .A(1'b1), .ZN(_u0_ch23_txsz[5] ) );
INV_X4 _u0_U11681  ( .A(1'b1), .ZN(_u0_ch23_txsz[4] ) );
INV_X4 _u0_U11679  ( .A(1'b1), .ZN(_u0_ch23_txsz[3] ) );
INV_X4 _u0_U11677  ( .A(1'b1), .ZN(_u0_ch23_txsz[2] ) );
INV_X4 _u0_U11675  ( .A(1'b1), .ZN(_u0_ch23_txsz[1] ) );
INV_X4 _u0_U11673  ( .A(1'b1), .ZN(_u0_ch23_txsz[0] ) );
INV_X4 _u0_U11671  ( .A(1'b1), .ZN(_u0_ch23_adr0[31] ) );
INV_X4 _u0_U11669  ( .A(1'b1), .ZN(_u0_ch23_adr0[30] ) );
INV_X4 _u0_U11667  ( .A(1'b1), .ZN(_u0_ch23_adr0[29] ) );
INV_X4 _u0_U11665  ( .A(1'b1), .ZN(_u0_ch23_adr0[28] ) );
INV_X4 _u0_U11663  ( .A(1'b1), .ZN(_u0_ch23_adr0[27] ) );
INV_X4 _u0_U11661  ( .A(1'b1), .ZN(_u0_ch23_adr0[26] ) );
INV_X4 _u0_U11659  ( .A(1'b1), .ZN(_u0_ch23_adr0[25] ) );
INV_X4 _u0_U11657  ( .A(1'b1), .ZN(_u0_ch23_adr0[24] ) );
INV_X4 _u0_U11655  ( .A(1'b1), .ZN(_u0_ch23_adr0[23] ) );
INV_X4 _u0_U11653  ( .A(1'b1), .ZN(_u0_ch23_adr0[22] ) );
INV_X4 _u0_U11651  ( .A(1'b1), .ZN(_u0_ch23_adr0[21] ) );
INV_X4 _u0_U11649  ( .A(1'b1), .ZN(_u0_ch23_adr0[20] ) );
INV_X4 _u0_U11647  ( .A(1'b1), .ZN(_u0_ch23_adr0[19] ) );
INV_X4 _u0_U11645  ( .A(1'b1), .ZN(_u0_ch23_adr0[18] ) );
INV_X4 _u0_U11643  ( .A(1'b1), .ZN(_u0_ch23_adr0[17] ) );
INV_X4 _u0_U11641  ( .A(1'b1), .ZN(_u0_ch23_adr0[16] ) );
INV_X4 _u0_U11639  ( .A(1'b1), .ZN(_u0_ch23_adr0[15] ) );
INV_X4 _u0_U11637  ( .A(1'b1), .ZN(_u0_ch23_adr0[14] ) );
INV_X4 _u0_U11635  ( .A(1'b1), .ZN(_u0_ch23_adr0[13] ) );
INV_X4 _u0_U11633  ( .A(1'b1), .ZN(_u0_ch23_adr0[12] ) );
INV_X4 _u0_U11631  ( .A(1'b1), .ZN(_u0_ch23_adr0[11] ) );
INV_X4 _u0_U11629  ( .A(1'b1), .ZN(_u0_ch23_adr0[10] ) );
INV_X4 _u0_U11627  ( .A(1'b1), .ZN(_u0_ch23_adr0[9] ) );
INV_X4 _u0_U11625  ( .A(1'b1), .ZN(_u0_ch23_adr0[8] ) );
INV_X4 _u0_U11623  ( .A(1'b1), .ZN(_u0_ch23_adr0[7] ) );
INV_X4 _u0_U11621  ( .A(1'b1), .ZN(_u0_ch23_adr0[6] ) );
INV_X4 _u0_U11619  ( .A(1'b1), .ZN(_u0_ch23_adr0[5] ) );
INV_X4 _u0_U11617  ( .A(1'b1), .ZN(_u0_ch23_adr0[4] ) );
INV_X4 _u0_U11615  ( .A(1'b1), .ZN(_u0_ch23_adr0[3] ) );
INV_X4 _u0_U11613  ( .A(1'b1), .ZN(_u0_ch23_adr0[2] ) );
INV_X4 _u0_U11611  ( .A(1'b1), .ZN(_u0_ch23_adr0[1] ) );
INV_X4 _u0_U11609  ( .A(1'b1), .ZN(_u0_ch23_adr0[0] ) );
INV_X4 _u0_U11607  ( .A(1'b1), .ZN(_u0_ch23_adr1[31] ) );
INV_X4 _u0_U11605  ( .A(1'b1), .ZN(_u0_ch23_adr1[30] ) );
INV_X4 _u0_U11603  ( .A(1'b1), .ZN(_u0_ch23_adr1[29] ) );
INV_X4 _u0_U11601  ( .A(1'b1), .ZN(_u0_ch23_adr1[28] ) );
INV_X4 _u0_U11599  ( .A(1'b1), .ZN(_u0_ch23_adr1[27] ) );
INV_X4 _u0_U11597  ( .A(1'b1), .ZN(_u0_ch23_adr1[26] ) );
INV_X4 _u0_U11595  ( .A(1'b1), .ZN(_u0_ch23_adr1[25] ) );
INV_X4 _u0_U11593  ( .A(1'b1), .ZN(_u0_ch23_adr1[24] ) );
INV_X4 _u0_U11591  ( .A(1'b1), .ZN(_u0_ch23_adr1[23] ) );
INV_X4 _u0_U11589  ( .A(1'b1), .ZN(_u0_ch23_adr1[22] ) );
INV_X4 _u0_U11587  ( .A(1'b1), .ZN(_u0_ch23_adr1[21] ) );
INV_X4 _u0_U11585  ( .A(1'b1), .ZN(_u0_ch23_adr1[20] ) );
INV_X4 _u0_U11583  ( .A(1'b1), .ZN(_u0_ch23_adr1[19] ) );
INV_X4 _u0_U11581  ( .A(1'b1), .ZN(_u0_ch23_adr1[18] ) );
INV_X4 _u0_U11579  ( .A(1'b1), .ZN(_u0_ch23_adr1[17] ) );
INV_X4 _u0_U11577  ( .A(1'b1), .ZN(_u0_ch23_adr1[16] ) );
INV_X4 _u0_U11575  ( .A(1'b1), .ZN(_u0_ch23_adr1[15] ) );
INV_X4 _u0_U11573  ( .A(1'b1), .ZN(_u0_ch23_adr1[14] ) );
INV_X4 _u0_U11571  ( .A(1'b1), .ZN(_u0_ch23_adr1[13] ) );
INV_X4 _u0_U11569  ( .A(1'b1), .ZN(_u0_ch23_adr1[12] ) );
INV_X4 _u0_U11567  ( .A(1'b1), .ZN(_u0_ch23_adr1[11] ) );
INV_X4 _u0_U11565  ( .A(1'b1), .ZN(_u0_ch23_adr1[10] ) );
INV_X4 _u0_U11563  ( .A(1'b1), .ZN(_u0_ch23_adr1[9] ) );
INV_X4 _u0_U11561  ( .A(1'b1), .ZN(_u0_ch23_adr1[8] ) );
INV_X4 _u0_U11559  ( .A(1'b1), .ZN(_u0_ch23_adr1[7] ) );
INV_X4 _u0_U11557  ( .A(1'b1), .ZN(_u0_ch23_adr1[6] ) );
INV_X4 _u0_U11555  ( .A(1'b1), .ZN(_u0_ch23_adr1[5] ) );
INV_X4 _u0_U11553  ( .A(1'b1), .ZN(_u0_ch23_adr1[4] ) );
INV_X4 _u0_U11551  ( .A(1'b1), .ZN(_u0_ch23_adr1[3] ) );
INV_X4 _u0_U11549  ( .A(1'b1), .ZN(_u0_ch23_adr1[2] ) );
INV_X4 _u0_U11547  ( .A(1'b1), .ZN(_u0_ch23_adr1[1] ) );
INV_X4 _u0_U11545  ( .A(1'b1), .ZN(_u0_ch23_adr1[0] ) );
INV_X4 _u0_U11543  ( .A(1'b0), .ZN(_u0_ch23_am0[31] ) );
INV_X4 _u0_U11541  ( .A(1'b0), .ZN(_u0_ch23_am0[30] ) );
INV_X4 _u0_U11539  ( .A(1'b0), .ZN(_u0_ch23_am0[29] ) );
INV_X4 _u0_U11537  ( .A(1'b0), .ZN(_u0_ch23_am0[28] ) );
INV_X4 _u0_U11535  ( .A(1'b0), .ZN(_u0_ch23_am0[27] ) );
INV_X4 _u0_U11533  ( .A(1'b0), .ZN(_u0_ch23_am0[26] ) );
INV_X4 _u0_U11531  ( .A(1'b0), .ZN(_u0_ch23_am0[25] ) );
INV_X4 _u0_U11529  ( .A(1'b0), .ZN(_u0_ch23_am0[24] ) );
INV_X4 _u0_U11527  ( .A(1'b0), .ZN(_u0_ch23_am0[23] ) );
INV_X4 _u0_U11525  ( .A(1'b0), .ZN(_u0_ch23_am0[22] ) );
INV_X4 _u0_U11523  ( .A(1'b0), .ZN(_u0_ch23_am0[21] ) );
INV_X4 _u0_U11521  ( .A(1'b0), .ZN(_u0_ch23_am0[20] ) );
INV_X4 _u0_U11519  ( .A(1'b0), .ZN(_u0_ch23_am0[19] ) );
INV_X4 _u0_U11517  ( .A(1'b0), .ZN(_u0_ch23_am0[18] ) );
INV_X4 _u0_U11515  ( .A(1'b0), .ZN(_u0_ch23_am0[17] ) );
INV_X4 _u0_U11513  ( .A(1'b0), .ZN(_u0_ch23_am0[16] ) );
INV_X4 _u0_U11511  ( .A(1'b0), .ZN(_u0_ch23_am0[15] ) );
INV_X4 _u0_U11509  ( .A(1'b0), .ZN(_u0_ch23_am0[14] ) );
INV_X4 _u0_U11507  ( .A(1'b0), .ZN(_u0_ch23_am0[13] ) );
INV_X4 _u0_U11505  ( .A(1'b0), .ZN(_u0_ch23_am0[12] ) );
INV_X4 _u0_U11503  ( .A(1'b0), .ZN(_u0_ch23_am0[11] ) );
INV_X4 _u0_U11501  ( .A(1'b0), .ZN(_u0_ch23_am0[10] ) );
INV_X4 _u0_U11499  ( .A(1'b0), .ZN(_u0_ch23_am0[9] ) );
INV_X4 _u0_U11497  ( .A(1'b0), .ZN(_u0_ch23_am0[8] ) );
INV_X4 _u0_U11495  ( .A(1'b0), .ZN(_u0_ch23_am0[7] ) );
INV_X4 _u0_U11493  ( .A(1'b0), .ZN(_u0_ch23_am0[6] ) );
INV_X4 _u0_U11491  ( .A(1'b0), .ZN(_u0_ch23_am0[5] ) );
INV_X4 _u0_U11489  ( .A(1'b0), .ZN(_u0_ch23_am0[4] ) );
INV_X4 _u0_U11487  ( .A(1'b1), .ZN(_u0_ch23_am0[3] ) );
INV_X4 _u0_U11485  ( .A(1'b1), .ZN(_u0_ch23_am0[2] ) );
INV_X4 _u0_U11483  ( .A(1'b1), .ZN(_u0_ch23_am0[1] ) );
INV_X4 _u0_U11481  ( .A(1'b1), .ZN(_u0_ch23_am0[0] ) );
INV_X4 _u0_U11479  ( .A(1'b0), .ZN(_u0_ch23_am1[31] ) );
INV_X4 _u0_U11477  ( .A(1'b0), .ZN(_u0_ch23_am1[30] ) );
INV_X4 _u0_U11475  ( .A(1'b0), .ZN(_u0_ch23_am1[29] ) );
INV_X4 _u0_U11473  ( .A(1'b0), .ZN(_u0_ch23_am1[28] ) );
INV_X4 _u0_U11471  ( .A(1'b0), .ZN(_u0_ch23_am1[27] ) );
INV_X4 _u0_U11469  ( .A(1'b0), .ZN(_u0_ch23_am1[26] ) );
INV_X4 _u0_U11467  ( .A(1'b0), .ZN(_u0_ch23_am1[25] ) );
INV_X4 _u0_U11465  ( .A(1'b0), .ZN(_u0_ch23_am1[24] ) );
INV_X4 _u0_U11463  ( .A(1'b0), .ZN(_u0_ch23_am1[23] ) );
INV_X4 _u0_U11461  ( .A(1'b0), .ZN(_u0_ch23_am1[22] ) );
INV_X4 _u0_U11459  ( .A(1'b0), .ZN(_u0_ch23_am1[21] ) );
INV_X4 _u0_U11457  ( .A(1'b0), .ZN(_u0_ch23_am1[20] ) );
INV_X4 _u0_U11455  ( .A(1'b0), .ZN(_u0_ch23_am1[19] ) );
INV_X4 _u0_U11453  ( .A(1'b0), .ZN(_u0_ch23_am1[18] ) );
INV_X4 _u0_U11451  ( .A(1'b0), .ZN(_u0_ch23_am1[17] ) );
INV_X4 _u0_U11449  ( .A(1'b0), .ZN(_u0_ch23_am1[16] ) );
INV_X4 _u0_U11447  ( .A(1'b0), .ZN(_u0_ch23_am1[15] ) );
INV_X4 _u0_U11445  ( .A(1'b0), .ZN(_u0_ch23_am1[14] ) );
INV_X4 _u0_U11443  ( .A(1'b0), .ZN(_u0_ch23_am1[13] ) );
INV_X4 _u0_U11441  ( .A(1'b0), .ZN(_u0_ch23_am1[12] ) );
INV_X4 _u0_U11439  ( .A(1'b0), .ZN(_u0_ch23_am1[11] ) );
INV_X4 _u0_U11437  ( .A(1'b0), .ZN(_u0_ch23_am1[10] ) );
INV_X4 _u0_U11435  ( .A(1'b0), .ZN(_u0_ch23_am1[9] ) );
INV_X4 _u0_U11433  ( .A(1'b0), .ZN(_u0_ch23_am1[8] ) );
INV_X4 _u0_U11431  ( .A(1'b0), .ZN(_u0_ch23_am1[7] ) );
INV_X4 _u0_U11429  ( .A(1'b0), .ZN(_u0_ch23_am1[6] ) );
INV_X4 _u0_U11427  ( .A(1'b0), .ZN(_u0_ch23_am1[5] ) );
INV_X4 _u0_U11425  ( .A(1'b0), .ZN(_u0_ch23_am1[4] ) );
INV_X4 _u0_U11423  ( .A(1'b1), .ZN(_u0_ch23_am1[3] ) );
INV_X4 _u0_U11421  ( .A(1'b1), .ZN(_u0_ch23_am1[2] ) );
INV_X4 _u0_U11419  ( .A(1'b1), .ZN(_u0_ch23_am1[1] ) );
INV_X4 _u0_U11417  ( .A(1'b1), .ZN(_u0_ch23_am1[0] ) );
INV_X4 _u0_U11415  ( .A(1'b1), .ZN(_u0_pointer24[31] ) );
INV_X4 _u0_U11413  ( .A(1'b1), .ZN(_u0_pointer24[30] ) );
INV_X4 _u0_U11411  ( .A(1'b1), .ZN(_u0_pointer24[29] ) );
INV_X4 _u0_U11409  ( .A(1'b1), .ZN(_u0_pointer24[28] ) );
INV_X4 _u0_U11407  ( .A(1'b1), .ZN(_u0_pointer24[27] ) );
INV_X4 _u0_U11405  ( .A(1'b1), .ZN(_u0_pointer24[26] ) );
INV_X4 _u0_U11403  ( .A(1'b1), .ZN(_u0_pointer24[25] ) );
INV_X4 _u0_U11401  ( .A(1'b1), .ZN(_u0_pointer24[24] ) );
INV_X4 _u0_U11399  ( .A(1'b1), .ZN(_u0_pointer24[23] ) );
INV_X4 _u0_U11397  ( .A(1'b1), .ZN(_u0_pointer24[22] ) );
INV_X4 _u0_U11395  ( .A(1'b1), .ZN(_u0_pointer24[21] ) );
INV_X4 _u0_U11393  ( .A(1'b1), .ZN(_u0_pointer24[20] ) );
INV_X4 _u0_U11391  ( .A(1'b1), .ZN(_u0_pointer24[19] ) );
INV_X4 _u0_U11389  ( .A(1'b1), .ZN(_u0_pointer24[18] ) );
INV_X4 _u0_U11387  ( .A(1'b1), .ZN(_u0_pointer24[17] ) );
INV_X4 _u0_U11385  ( .A(1'b1), .ZN(_u0_pointer24[16] ) );
INV_X4 _u0_U11383  ( .A(1'b1), .ZN(_u0_pointer24[15] ) );
INV_X4 _u0_U11381  ( .A(1'b1), .ZN(_u0_pointer24[14] ) );
INV_X4 _u0_U11379  ( .A(1'b1), .ZN(_u0_pointer24[13] ) );
INV_X4 _u0_U11377  ( .A(1'b1), .ZN(_u0_pointer24[12] ) );
INV_X4 _u0_U11375  ( .A(1'b1), .ZN(_u0_pointer24[11] ) );
INV_X4 _u0_U11373  ( .A(1'b1), .ZN(_u0_pointer24[10] ) );
INV_X4 _u0_U11371  ( .A(1'b1), .ZN(_u0_pointer24[9] ) );
INV_X4 _u0_U11369  ( .A(1'b1), .ZN(_u0_pointer24[8] ) );
INV_X4 _u0_U11367  ( .A(1'b1), .ZN(_u0_pointer24[7] ) );
INV_X4 _u0_U11365  ( .A(1'b1), .ZN(_u0_pointer24[6] ) );
INV_X4 _u0_U11363  ( .A(1'b1), .ZN(_u0_pointer24[5] ) );
INV_X4 _u0_U11361  ( .A(1'b1), .ZN(_u0_pointer24[4] ) );
INV_X4 _u0_U11359  ( .A(1'b1), .ZN(_u0_pointer24[3] ) );
INV_X4 _u0_U11357  ( .A(1'b1), .ZN(_u0_pointer24[2] ) );
INV_X4 _u0_U11355  ( .A(1'b1), .ZN(_u0_pointer24[1] ) );
INV_X4 _u0_U11353  ( .A(1'b1), .ZN(_u0_pointer24[0] ) );
INV_X4 _u0_U11351  ( .A(1'b1), .ZN(_u0_pointer24_s[31] ) );
INV_X4 _u0_U11349  ( .A(1'b1), .ZN(_u0_pointer24_s[30] ) );
INV_X4 _u0_U11347  ( .A(1'b1), .ZN(_u0_pointer24_s[29] ) );
INV_X4 _u0_U11345  ( .A(1'b1), .ZN(_u0_pointer24_s[28] ) );
INV_X4 _u0_U11343  ( .A(1'b1), .ZN(_u0_pointer24_s[27] ) );
INV_X4 _u0_U11341  ( .A(1'b1), .ZN(_u0_pointer24_s[26] ) );
INV_X4 _u0_U11339  ( .A(1'b1), .ZN(_u0_pointer24_s[25] ) );
INV_X4 _u0_U11337  ( .A(1'b1), .ZN(_u0_pointer24_s[24] ) );
INV_X4 _u0_U11335  ( .A(1'b1), .ZN(_u0_pointer24_s[23] ) );
INV_X4 _u0_U11333  ( .A(1'b1), .ZN(_u0_pointer24_s[22] ) );
INV_X4 _u0_U11331  ( .A(1'b1), .ZN(_u0_pointer24_s[21] ) );
INV_X4 _u0_U11329  ( .A(1'b1), .ZN(_u0_pointer24_s[20] ) );
INV_X4 _u0_U11327  ( .A(1'b1), .ZN(_u0_pointer24_s[19] ) );
INV_X4 _u0_U11325  ( .A(1'b1), .ZN(_u0_pointer24_s[18] ) );
INV_X4 _u0_U11323  ( .A(1'b1), .ZN(_u0_pointer24_s[17] ) );
INV_X4 _u0_U11321  ( .A(1'b1), .ZN(_u0_pointer24_s[16] ) );
INV_X4 _u0_U11319  ( .A(1'b1), .ZN(_u0_pointer24_s[15] ) );
INV_X4 _u0_U11317  ( .A(1'b1), .ZN(_u0_pointer24_s[14] ) );
INV_X4 _u0_U11315  ( .A(1'b1), .ZN(_u0_pointer24_s[13] ) );
INV_X4 _u0_U11313  ( .A(1'b1), .ZN(_u0_pointer24_s[12] ) );
INV_X4 _u0_U11311  ( .A(1'b1), .ZN(_u0_pointer24_s[11] ) );
INV_X4 _u0_U11309  ( .A(1'b1), .ZN(_u0_pointer24_s[10] ) );
INV_X4 _u0_U11307  ( .A(1'b1), .ZN(_u0_pointer24_s[9] ) );
INV_X4 _u0_U11305  ( .A(1'b1), .ZN(_u0_pointer24_s[8] ) );
INV_X4 _u0_U11303  ( .A(1'b1), .ZN(_u0_pointer24_s[7] ) );
INV_X4 _u0_U11301  ( .A(1'b1), .ZN(_u0_pointer24_s[6] ) );
INV_X4 _u0_U11299  ( .A(1'b1), .ZN(_u0_pointer24_s[5] ) );
INV_X4 _u0_U11297  ( .A(1'b1), .ZN(_u0_pointer24_s[4] ) );
INV_X4 _u0_U11295  ( .A(1'b1), .ZN(_u0_pointer24_s[3] ) );
INV_X4 _u0_U11293  ( .A(1'b1), .ZN(_u0_pointer24_s[2] ) );
INV_X4 _u0_U11291  ( .A(1'b1), .ZN(_u0_pointer24_s[1] ) );
INV_X4 _u0_U11289  ( .A(1'b1), .ZN(_u0_pointer24_s[0] ) );
INV_X4 _u0_U11287  ( .A(1'b1), .ZN(_u0_ch24_csr[31] ) );
INV_X4 _u0_U11285  ( .A(1'b1), .ZN(_u0_ch24_csr[30] ) );
INV_X4 _u0_U11283  ( .A(1'b1), .ZN(_u0_ch24_csr[29] ) );
INV_X4 _u0_U11281  ( .A(1'b1), .ZN(_u0_ch24_csr[28] ) );
INV_X4 _u0_U11279  ( .A(1'b1), .ZN(_u0_ch24_csr[27] ) );
INV_X4 _u0_U11277  ( .A(1'b1), .ZN(_u0_ch24_csr[26] ) );
INV_X4 _u0_U11275  ( .A(1'b1), .ZN(_u0_ch24_csr[25] ) );
INV_X4 _u0_U11273  ( .A(1'b1), .ZN(_u0_ch24_csr[24] ) );
INV_X4 _u0_U11271  ( .A(1'b1), .ZN(_u0_ch24_csr[23] ) );
INV_X4 _u0_U11269  ( .A(1'b1), .ZN(_u0_ch24_csr[22] ) );
INV_X4 _u0_U11267  ( .A(1'b1), .ZN(_u0_ch24_csr[21] ) );
INV_X4 _u0_U11265  ( .A(1'b1), .ZN(_u0_ch24_csr[20] ) );
INV_X4 _u0_U11263  ( .A(1'b1), .ZN(_u0_ch24_csr[19] ) );
INV_X4 _u0_U11261  ( .A(1'b1), .ZN(_u0_ch24_csr[18] ) );
INV_X4 _u0_U11259  ( .A(1'b1), .ZN(_u0_ch24_csr[17] ) );
INV_X4 _u0_U11257  ( .A(1'b1), .ZN(_u0_ch24_csr[16] ) );
INV_X4 _u0_U11255  ( .A(1'b1), .ZN(_u0_ch24_csr[15] ) );
INV_X4 _u0_U11253  ( .A(1'b1), .ZN(_u0_ch24_csr[14] ) );
INV_X4 _u0_U11251  ( .A(1'b1), .ZN(_u0_ch24_csr[13] ) );
INV_X4 _u0_U11249  ( .A(1'b1), .ZN(_u0_ch24_csr[12] ) );
INV_X4 _u0_U11247  ( .A(1'b1), .ZN(_u0_ch24_csr[11] ) );
INV_X4 _u0_U11245  ( .A(1'b1), .ZN(_u0_ch24_csr[10] ) );
INV_X4 _u0_U11243  ( .A(1'b1), .ZN(_u0_ch24_csr[9] ) );
INV_X4 _u0_U11241  ( .A(1'b1), .ZN(_u0_ch24_csr[8] ) );
INV_X4 _u0_U11239  ( .A(1'b1), .ZN(_u0_ch24_csr[7] ) );
INV_X4 _u0_U11237  ( .A(1'b1), .ZN(_u0_ch24_csr[6] ) );
INV_X4 _u0_U11235  ( .A(1'b1), .ZN(_u0_ch24_csr[5] ) );
INV_X4 _u0_U11233  ( .A(1'b1), .ZN(_u0_ch24_csr[4] ) );
INV_X4 _u0_U11231  ( .A(1'b1), .ZN(_u0_ch24_csr[3] ) );
INV_X4 _u0_U11229  ( .A(1'b1), .ZN(_u0_ch24_csr[2] ) );
INV_X4 _u0_U11227  ( .A(1'b1), .ZN(_u0_ch24_csr[1] ) );
INV_X4 _u0_U11225  ( .A(1'b1), .ZN(_u0_ch24_csr[0] ) );
INV_X4 _u0_U11223  ( .A(1'b1), .ZN(_u0_ch24_txsz[31] ) );
INV_X4 _u0_U11221  ( .A(1'b1), .ZN(_u0_ch24_txsz[30] ) );
INV_X4 _u0_U11219  ( .A(1'b1), .ZN(_u0_ch24_txsz[29] ) );
INV_X4 _u0_U11217  ( .A(1'b1), .ZN(_u0_ch24_txsz[28] ) );
INV_X4 _u0_U11215  ( .A(1'b1), .ZN(_u0_ch24_txsz[27] ) );
INV_X4 _u0_U11213  ( .A(1'b1), .ZN(_u0_ch24_txsz[26] ) );
INV_X4 _u0_U11211  ( .A(1'b1), .ZN(_u0_ch24_txsz[25] ) );
INV_X4 _u0_U11209  ( .A(1'b1), .ZN(_u0_ch24_txsz[24] ) );
INV_X4 _u0_U11207  ( .A(1'b1), .ZN(_u0_ch24_txsz[23] ) );
INV_X4 _u0_U11205  ( .A(1'b1), .ZN(_u0_ch24_txsz[22] ) );
INV_X4 _u0_U11203  ( .A(1'b1), .ZN(_u0_ch24_txsz[21] ) );
INV_X4 _u0_U11201  ( .A(1'b1), .ZN(_u0_ch24_txsz[20] ) );
INV_X4 _u0_U11199  ( .A(1'b1), .ZN(_u0_ch24_txsz[19] ) );
INV_X4 _u0_U11197  ( .A(1'b1), .ZN(_u0_ch24_txsz[18] ) );
INV_X4 _u0_U11195  ( .A(1'b1), .ZN(_u0_ch24_txsz[17] ) );
INV_X4 _u0_U11193  ( .A(1'b1), .ZN(_u0_ch24_txsz[16] ) );
INV_X4 _u0_U11191  ( .A(1'b1), .ZN(_u0_ch24_txsz[15] ) );
INV_X4 _u0_U11189  ( .A(1'b1), .ZN(_u0_ch24_txsz[14] ) );
INV_X4 _u0_U11187  ( .A(1'b1), .ZN(_u0_ch24_txsz[13] ) );
INV_X4 _u0_U11185  ( .A(1'b1), .ZN(_u0_ch24_txsz[12] ) );
INV_X4 _u0_U11183  ( .A(1'b1), .ZN(_u0_ch24_txsz[11] ) );
INV_X4 _u0_U11181  ( .A(1'b1), .ZN(_u0_ch24_txsz[10] ) );
INV_X4 _u0_U11179  ( .A(1'b1), .ZN(_u0_ch24_txsz[9] ) );
INV_X4 _u0_U11177  ( .A(1'b1), .ZN(_u0_ch24_txsz[8] ) );
INV_X4 _u0_U11175  ( .A(1'b1), .ZN(_u0_ch24_txsz[7] ) );
INV_X4 _u0_U11173  ( .A(1'b1), .ZN(_u0_ch24_txsz[6] ) );
INV_X4 _u0_U11171  ( .A(1'b1), .ZN(_u0_ch24_txsz[5] ) );
INV_X4 _u0_U11169  ( .A(1'b1), .ZN(_u0_ch24_txsz[4] ) );
INV_X4 _u0_U11167  ( .A(1'b1), .ZN(_u0_ch24_txsz[3] ) );
INV_X4 _u0_U11165  ( .A(1'b1), .ZN(_u0_ch24_txsz[2] ) );
INV_X4 _u0_U11163  ( .A(1'b1), .ZN(_u0_ch24_txsz[1] ) );
INV_X4 _u0_U11161  ( .A(1'b1), .ZN(_u0_ch24_txsz[0] ) );
INV_X4 _u0_U11159  ( .A(1'b1), .ZN(_u0_ch24_adr0[31] ) );
INV_X4 _u0_U11157  ( .A(1'b1), .ZN(_u0_ch24_adr0[30] ) );
INV_X4 _u0_U11155  ( .A(1'b1), .ZN(_u0_ch24_adr0[29] ) );
INV_X4 _u0_U11153  ( .A(1'b1), .ZN(_u0_ch24_adr0[28] ) );
INV_X4 _u0_U11151  ( .A(1'b1), .ZN(_u0_ch24_adr0[27] ) );
INV_X4 _u0_U11149  ( .A(1'b1), .ZN(_u0_ch24_adr0[26] ) );
INV_X4 _u0_U11147  ( .A(1'b1), .ZN(_u0_ch24_adr0[25] ) );
INV_X4 _u0_U11145  ( .A(1'b1), .ZN(_u0_ch24_adr0[24] ) );
INV_X4 _u0_U11143  ( .A(1'b1), .ZN(_u0_ch24_adr0[23] ) );
INV_X4 _u0_U11141  ( .A(1'b1), .ZN(_u0_ch24_adr0[22] ) );
INV_X4 _u0_U11139  ( .A(1'b1), .ZN(_u0_ch24_adr0[21] ) );
INV_X4 _u0_U11137  ( .A(1'b1), .ZN(_u0_ch24_adr0[20] ) );
INV_X4 _u0_U11135  ( .A(1'b1), .ZN(_u0_ch24_adr0[19] ) );
INV_X4 _u0_U11133  ( .A(1'b1), .ZN(_u0_ch24_adr0[18] ) );
INV_X4 _u0_U11131  ( .A(1'b1), .ZN(_u0_ch24_adr0[17] ) );
INV_X4 _u0_U11129  ( .A(1'b1), .ZN(_u0_ch24_adr0[16] ) );
INV_X4 _u0_U11127  ( .A(1'b1), .ZN(_u0_ch24_adr0[15] ) );
INV_X4 _u0_U11125  ( .A(1'b1), .ZN(_u0_ch24_adr0[14] ) );
INV_X4 _u0_U11123  ( .A(1'b1), .ZN(_u0_ch24_adr0[13] ) );
INV_X4 _u0_U11121  ( .A(1'b1), .ZN(_u0_ch24_adr0[12] ) );
INV_X4 _u0_U11119  ( .A(1'b1), .ZN(_u0_ch24_adr0[11] ) );
INV_X4 _u0_U11117  ( .A(1'b1), .ZN(_u0_ch24_adr0[10] ) );
INV_X4 _u0_U11115  ( .A(1'b1), .ZN(_u0_ch24_adr0[9] ) );
INV_X4 _u0_U11113  ( .A(1'b1), .ZN(_u0_ch24_adr0[8] ) );
INV_X4 _u0_U11111  ( .A(1'b1), .ZN(_u0_ch24_adr0[7] ) );
INV_X4 _u0_U11109  ( .A(1'b1), .ZN(_u0_ch24_adr0[6] ) );
INV_X4 _u0_U11107  ( .A(1'b1), .ZN(_u0_ch24_adr0[5] ) );
INV_X4 _u0_U11105  ( .A(1'b1), .ZN(_u0_ch24_adr0[4] ) );
INV_X4 _u0_U11103  ( .A(1'b1), .ZN(_u0_ch24_adr0[3] ) );
INV_X4 _u0_U11101  ( .A(1'b1), .ZN(_u0_ch24_adr0[2] ) );
INV_X4 _u0_U11099  ( .A(1'b1), .ZN(_u0_ch24_adr0[1] ) );
INV_X4 _u0_U11097  ( .A(1'b1), .ZN(_u0_ch24_adr0[0] ) );
INV_X4 _u0_U11095  ( .A(1'b1), .ZN(_u0_ch24_adr1[31] ) );
INV_X4 _u0_U11093  ( .A(1'b1), .ZN(_u0_ch24_adr1[30] ) );
INV_X4 _u0_U11091  ( .A(1'b1), .ZN(_u0_ch24_adr1[29] ) );
INV_X4 _u0_U11089  ( .A(1'b1), .ZN(_u0_ch24_adr1[28] ) );
INV_X4 _u0_U11087  ( .A(1'b1), .ZN(_u0_ch24_adr1[27] ) );
INV_X4 _u0_U11085  ( .A(1'b1), .ZN(_u0_ch24_adr1[26] ) );
INV_X4 _u0_U11083  ( .A(1'b1), .ZN(_u0_ch24_adr1[25] ) );
INV_X4 _u0_U11081  ( .A(1'b1), .ZN(_u0_ch24_adr1[24] ) );
INV_X4 _u0_U11079  ( .A(1'b1), .ZN(_u0_ch24_adr1[23] ) );
INV_X4 _u0_U11077  ( .A(1'b1), .ZN(_u0_ch24_adr1[22] ) );
INV_X4 _u0_U11075  ( .A(1'b1), .ZN(_u0_ch24_adr1[21] ) );
INV_X4 _u0_U11073  ( .A(1'b1), .ZN(_u0_ch24_adr1[20] ) );
INV_X4 _u0_U11071  ( .A(1'b1), .ZN(_u0_ch24_adr1[19] ) );
INV_X4 _u0_U11069  ( .A(1'b1), .ZN(_u0_ch24_adr1[18] ) );
INV_X4 _u0_U11067  ( .A(1'b1), .ZN(_u0_ch24_adr1[17] ) );
INV_X4 _u0_U11065  ( .A(1'b1), .ZN(_u0_ch24_adr1[16] ) );
INV_X4 _u0_U11063  ( .A(1'b1), .ZN(_u0_ch24_adr1[15] ) );
INV_X4 _u0_U11061  ( .A(1'b1), .ZN(_u0_ch24_adr1[14] ) );
INV_X4 _u0_U11059  ( .A(1'b1), .ZN(_u0_ch24_adr1[13] ) );
INV_X4 _u0_U11057  ( .A(1'b1), .ZN(_u0_ch24_adr1[12] ) );
INV_X4 _u0_U11055  ( .A(1'b1), .ZN(_u0_ch24_adr1[11] ) );
INV_X4 _u0_U11053  ( .A(1'b1), .ZN(_u0_ch24_adr1[10] ) );
INV_X4 _u0_U11051  ( .A(1'b1), .ZN(_u0_ch24_adr1[9] ) );
INV_X4 _u0_U11049  ( .A(1'b1), .ZN(_u0_ch24_adr1[8] ) );
INV_X4 _u0_U11047  ( .A(1'b1), .ZN(_u0_ch24_adr1[7] ) );
INV_X4 _u0_U11045  ( .A(1'b1), .ZN(_u0_ch24_adr1[6] ) );
INV_X4 _u0_U11043  ( .A(1'b1), .ZN(_u0_ch24_adr1[5] ) );
INV_X4 _u0_U11041  ( .A(1'b1), .ZN(_u0_ch24_adr1[4] ) );
INV_X4 _u0_U11039  ( .A(1'b1), .ZN(_u0_ch24_adr1[3] ) );
INV_X4 _u0_U11037  ( .A(1'b1), .ZN(_u0_ch24_adr1[2] ) );
INV_X4 _u0_U11035  ( .A(1'b1), .ZN(_u0_ch24_adr1[1] ) );
INV_X4 _u0_U11033  ( .A(1'b1), .ZN(_u0_ch24_adr1[0] ) );
INV_X4 _u0_U11031  ( .A(1'b0), .ZN(_u0_ch24_am0[31] ) );
INV_X4 _u0_U11029  ( .A(1'b0), .ZN(_u0_ch24_am0[30] ) );
INV_X4 _u0_U11027  ( .A(1'b0), .ZN(_u0_ch24_am0[29] ) );
INV_X4 _u0_U11025  ( .A(1'b0), .ZN(_u0_ch24_am0[28] ) );
INV_X4 _u0_U11023  ( .A(1'b0), .ZN(_u0_ch24_am0[27] ) );
INV_X4 _u0_U11021  ( .A(1'b0), .ZN(_u0_ch24_am0[26] ) );
INV_X4 _u0_U11019  ( .A(1'b0), .ZN(_u0_ch24_am0[25] ) );
INV_X4 _u0_U11017  ( .A(1'b0), .ZN(_u0_ch24_am0[24] ) );
INV_X4 _u0_U11015  ( .A(1'b0), .ZN(_u0_ch24_am0[23] ) );
INV_X4 _u0_U11013  ( .A(1'b0), .ZN(_u0_ch24_am0[22] ) );
INV_X4 _u0_U11011  ( .A(1'b0), .ZN(_u0_ch24_am0[21] ) );
INV_X4 _u0_U11009  ( .A(1'b0), .ZN(_u0_ch24_am0[20] ) );
INV_X4 _u0_U11007  ( .A(1'b0), .ZN(_u0_ch24_am0[19] ) );
INV_X4 _u0_U11005  ( .A(1'b0), .ZN(_u0_ch24_am0[18] ) );
INV_X4 _u0_U11003  ( .A(1'b0), .ZN(_u0_ch24_am0[17] ) );
INV_X4 _u0_U11001  ( .A(1'b0), .ZN(_u0_ch24_am0[16] ) );
INV_X4 _u0_U10999  ( .A(1'b0), .ZN(_u0_ch24_am0[15] ) );
INV_X4 _u0_U10997  ( .A(1'b0), .ZN(_u0_ch24_am0[14] ) );
INV_X4 _u0_U10995  ( .A(1'b0), .ZN(_u0_ch24_am0[13] ) );
INV_X4 _u0_U10993  ( .A(1'b0), .ZN(_u0_ch24_am0[12] ) );
INV_X4 _u0_U10991  ( .A(1'b0), .ZN(_u0_ch24_am0[11] ) );
INV_X4 _u0_U10989  ( .A(1'b0), .ZN(_u0_ch24_am0[10] ) );
INV_X4 _u0_U10987  ( .A(1'b0), .ZN(_u0_ch24_am0[9] ) );
INV_X4 _u0_U10985  ( .A(1'b0), .ZN(_u0_ch24_am0[8] ) );
INV_X4 _u0_U10983  ( .A(1'b0), .ZN(_u0_ch24_am0[7] ) );
INV_X4 _u0_U10981  ( .A(1'b0), .ZN(_u0_ch24_am0[6] ) );
INV_X4 _u0_U10979  ( .A(1'b0), .ZN(_u0_ch24_am0[5] ) );
INV_X4 _u0_U10977  ( .A(1'b0), .ZN(_u0_ch24_am0[4] ) );
INV_X4 _u0_U10975  ( .A(1'b1), .ZN(_u0_ch24_am0[3] ) );
INV_X4 _u0_U10973  ( .A(1'b1), .ZN(_u0_ch24_am0[2] ) );
INV_X4 _u0_U10971  ( .A(1'b1), .ZN(_u0_ch24_am0[1] ) );
INV_X4 _u0_U10969  ( .A(1'b1), .ZN(_u0_ch24_am0[0] ) );
INV_X4 _u0_U10967  ( .A(1'b0), .ZN(_u0_ch24_am1[31] ) );
INV_X4 _u0_U10965  ( .A(1'b0), .ZN(_u0_ch24_am1[30] ) );
INV_X4 _u0_U10963  ( .A(1'b0), .ZN(_u0_ch24_am1[29] ) );
INV_X4 _u0_U10961  ( .A(1'b0), .ZN(_u0_ch24_am1[28] ) );
INV_X4 _u0_U10959  ( .A(1'b0), .ZN(_u0_ch24_am1[27] ) );
INV_X4 _u0_U10957  ( .A(1'b0), .ZN(_u0_ch24_am1[26] ) );
INV_X4 _u0_U10955  ( .A(1'b0), .ZN(_u0_ch24_am1[25] ) );
INV_X4 _u0_U10953  ( .A(1'b0), .ZN(_u0_ch24_am1[24] ) );
INV_X4 _u0_U10951  ( .A(1'b0), .ZN(_u0_ch24_am1[23] ) );
INV_X4 _u0_U10949  ( .A(1'b0), .ZN(_u0_ch24_am1[22] ) );
INV_X4 _u0_U10947  ( .A(1'b0), .ZN(_u0_ch24_am1[21] ) );
INV_X4 _u0_U10945  ( .A(1'b0), .ZN(_u0_ch24_am1[20] ) );
INV_X4 _u0_U10943  ( .A(1'b0), .ZN(_u0_ch24_am1[19] ) );
INV_X4 _u0_U10941  ( .A(1'b0), .ZN(_u0_ch24_am1[18] ) );
INV_X4 _u0_U10939  ( .A(1'b0), .ZN(_u0_ch24_am1[17] ) );
INV_X4 _u0_U10937  ( .A(1'b0), .ZN(_u0_ch24_am1[16] ) );
INV_X4 _u0_U10935  ( .A(1'b0), .ZN(_u0_ch24_am1[15] ) );
INV_X4 _u0_U10933  ( .A(1'b0), .ZN(_u0_ch24_am1[14] ) );
INV_X4 _u0_U10931  ( .A(1'b0), .ZN(_u0_ch24_am1[13] ) );
INV_X4 _u0_U10929  ( .A(1'b0), .ZN(_u0_ch24_am1[12] ) );
INV_X4 _u0_U10927  ( .A(1'b0), .ZN(_u0_ch24_am1[11] ) );
INV_X4 _u0_U10925  ( .A(1'b0), .ZN(_u0_ch24_am1[10] ) );
INV_X4 _u0_U10923  ( .A(1'b0), .ZN(_u0_ch24_am1[9] ) );
INV_X4 _u0_U10921  ( .A(1'b0), .ZN(_u0_ch24_am1[8] ) );
INV_X4 _u0_U10919  ( .A(1'b0), .ZN(_u0_ch24_am1[7] ) );
INV_X4 _u0_U10917  ( .A(1'b0), .ZN(_u0_ch24_am1[6] ) );
INV_X4 _u0_U10915  ( .A(1'b0), .ZN(_u0_ch24_am1[5] ) );
INV_X4 _u0_U10913  ( .A(1'b0), .ZN(_u0_ch24_am1[4] ) );
INV_X4 _u0_U10911  ( .A(1'b1), .ZN(_u0_ch24_am1[3] ) );
INV_X4 _u0_U10909  ( .A(1'b1), .ZN(_u0_ch24_am1[2] ) );
INV_X4 _u0_U10907  ( .A(1'b1), .ZN(_u0_ch24_am1[1] ) );
INV_X4 _u0_U10905  ( .A(1'b1), .ZN(_u0_ch24_am1[0] ) );
INV_X4 _u0_U10903  ( .A(1'b1), .ZN(_u0_pointer25[31] ) );
INV_X4 _u0_U10901  ( .A(1'b1), .ZN(_u0_pointer25[30] ) );
INV_X4 _u0_U10899  ( .A(1'b1), .ZN(_u0_pointer25[29] ) );
INV_X4 _u0_U10897  ( .A(1'b1), .ZN(_u0_pointer25[28] ) );
INV_X4 _u0_U10895  ( .A(1'b1), .ZN(_u0_pointer25[27] ) );
INV_X4 _u0_U10893  ( .A(1'b1), .ZN(_u0_pointer25[26] ) );
INV_X4 _u0_U10891  ( .A(1'b1), .ZN(_u0_pointer25[25] ) );
INV_X4 _u0_U10889  ( .A(1'b1), .ZN(_u0_pointer25[24] ) );
INV_X4 _u0_U10887  ( .A(1'b1), .ZN(_u0_pointer25[23] ) );
INV_X4 _u0_U10885  ( .A(1'b1), .ZN(_u0_pointer25[22] ) );
INV_X4 _u0_U10883  ( .A(1'b1), .ZN(_u0_pointer25[21] ) );
INV_X4 _u0_U10881  ( .A(1'b1), .ZN(_u0_pointer25[20] ) );
INV_X4 _u0_U10879  ( .A(1'b1), .ZN(_u0_pointer25[19] ) );
INV_X4 _u0_U10877  ( .A(1'b1), .ZN(_u0_pointer25[18] ) );
INV_X4 _u0_U10875  ( .A(1'b1), .ZN(_u0_pointer25[17] ) );
INV_X4 _u0_U10873  ( .A(1'b1), .ZN(_u0_pointer25[16] ) );
INV_X4 _u0_U10871  ( .A(1'b1), .ZN(_u0_pointer25[15] ) );
INV_X4 _u0_U10869  ( .A(1'b1), .ZN(_u0_pointer25[14] ) );
INV_X4 _u0_U10867  ( .A(1'b1), .ZN(_u0_pointer25[13] ) );
INV_X4 _u0_U10865  ( .A(1'b1), .ZN(_u0_pointer25[12] ) );
INV_X4 _u0_U10863  ( .A(1'b1), .ZN(_u0_pointer25[11] ) );
INV_X4 _u0_U10861  ( .A(1'b1), .ZN(_u0_pointer25[10] ) );
INV_X4 _u0_U10859  ( .A(1'b1), .ZN(_u0_pointer25[9] ) );
INV_X4 _u0_U10857  ( .A(1'b1), .ZN(_u0_pointer25[8] ) );
INV_X4 _u0_U10855  ( .A(1'b1), .ZN(_u0_pointer25[7] ) );
INV_X4 _u0_U10853  ( .A(1'b1), .ZN(_u0_pointer25[6] ) );
INV_X4 _u0_U10851  ( .A(1'b1), .ZN(_u0_pointer25[5] ) );
INV_X4 _u0_U10849  ( .A(1'b1), .ZN(_u0_pointer25[4] ) );
INV_X4 _u0_U10847  ( .A(1'b1), .ZN(_u0_pointer25[3] ) );
INV_X4 _u0_U10845  ( .A(1'b1), .ZN(_u0_pointer25[2] ) );
INV_X4 _u0_U10843  ( .A(1'b1), .ZN(_u0_pointer25[1] ) );
INV_X4 _u0_U10841  ( .A(1'b1), .ZN(_u0_pointer25[0] ) );
INV_X4 _u0_U10839  ( .A(1'b1), .ZN(_u0_pointer25_s[31] ) );
INV_X4 _u0_U10837  ( .A(1'b1), .ZN(_u0_pointer25_s[30] ) );
INV_X4 _u0_U10835  ( .A(1'b1), .ZN(_u0_pointer25_s[29] ) );
INV_X4 _u0_U10833  ( .A(1'b1), .ZN(_u0_pointer25_s[28] ) );
INV_X4 _u0_U10831  ( .A(1'b1), .ZN(_u0_pointer25_s[27] ) );
INV_X4 _u0_U10829  ( .A(1'b1), .ZN(_u0_pointer25_s[26] ) );
INV_X4 _u0_U10827  ( .A(1'b1), .ZN(_u0_pointer25_s[25] ) );
INV_X4 _u0_U10825  ( .A(1'b1), .ZN(_u0_pointer25_s[24] ) );
INV_X4 _u0_U10823  ( .A(1'b1), .ZN(_u0_pointer25_s[23] ) );
INV_X4 _u0_U10821  ( .A(1'b1), .ZN(_u0_pointer25_s[22] ) );
INV_X4 _u0_U10819  ( .A(1'b1), .ZN(_u0_pointer25_s[21] ) );
INV_X4 _u0_U10817  ( .A(1'b1), .ZN(_u0_pointer25_s[20] ) );
INV_X4 _u0_U10815  ( .A(1'b1), .ZN(_u0_pointer25_s[19] ) );
INV_X4 _u0_U10813  ( .A(1'b1), .ZN(_u0_pointer25_s[18] ) );
INV_X4 _u0_U10811  ( .A(1'b1), .ZN(_u0_pointer25_s[17] ) );
INV_X4 _u0_U10809  ( .A(1'b1), .ZN(_u0_pointer25_s[16] ) );
INV_X4 _u0_U10807  ( .A(1'b1), .ZN(_u0_pointer25_s[15] ) );
INV_X4 _u0_U10805  ( .A(1'b1), .ZN(_u0_pointer25_s[14] ) );
INV_X4 _u0_U10803  ( .A(1'b1), .ZN(_u0_pointer25_s[13] ) );
INV_X4 _u0_U10801  ( .A(1'b1), .ZN(_u0_pointer25_s[12] ) );
INV_X4 _u0_U10799  ( .A(1'b1), .ZN(_u0_pointer25_s[11] ) );
INV_X4 _u0_U10797  ( .A(1'b1), .ZN(_u0_pointer25_s[10] ) );
INV_X4 _u0_U10795  ( .A(1'b1), .ZN(_u0_pointer25_s[9] ) );
INV_X4 _u0_U10793  ( .A(1'b1), .ZN(_u0_pointer25_s[8] ) );
INV_X4 _u0_U10791  ( .A(1'b1), .ZN(_u0_pointer25_s[7] ) );
INV_X4 _u0_U10789  ( .A(1'b1), .ZN(_u0_pointer25_s[6] ) );
INV_X4 _u0_U10787  ( .A(1'b1), .ZN(_u0_pointer25_s[5] ) );
INV_X4 _u0_U10785  ( .A(1'b1), .ZN(_u0_pointer25_s[4] ) );
INV_X4 _u0_U10783  ( .A(1'b1), .ZN(_u0_pointer25_s[3] ) );
INV_X4 _u0_U10781  ( .A(1'b1), .ZN(_u0_pointer25_s[2] ) );
INV_X4 _u0_U10779  ( .A(1'b1), .ZN(_u0_pointer25_s[1] ) );
INV_X4 _u0_U10777  ( .A(1'b1), .ZN(_u0_pointer25_s[0] ) );
INV_X4 _u0_U10775  ( .A(1'b1), .ZN(_u0_ch25_csr[31] ) );
INV_X4 _u0_U10773  ( .A(1'b1), .ZN(_u0_ch25_csr[30] ) );
INV_X4 _u0_U10771  ( .A(1'b1), .ZN(_u0_ch25_csr[29] ) );
INV_X4 _u0_U10769  ( .A(1'b1), .ZN(_u0_ch25_csr[28] ) );
INV_X4 _u0_U10767  ( .A(1'b1), .ZN(_u0_ch25_csr[27] ) );
INV_X4 _u0_U10765  ( .A(1'b1), .ZN(_u0_ch25_csr[26] ) );
INV_X4 _u0_U10763  ( .A(1'b1), .ZN(_u0_ch25_csr[25] ) );
INV_X4 _u0_U10761  ( .A(1'b1), .ZN(_u0_ch25_csr[24] ) );
INV_X4 _u0_U10759  ( .A(1'b1), .ZN(_u0_ch25_csr[23] ) );
INV_X4 _u0_U10757  ( .A(1'b1), .ZN(_u0_ch25_csr[22] ) );
INV_X4 _u0_U10755  ( .A(1'b1), .ZN(_u0_ch25_csr[21] ) );
INV_X4 _u0_U10753  ( .A(1'b1), .ZN(_u0_ch25_csr[20] ) );
INV_X4 _u0_U10751  ( .A(1'b1), .ZN(_u0_ch25_csr[19] ) );
INV_X4 _u0_U10749  ( .A(1'b1), .ZN(_u0_ch25_csr[18] ) );
INV_X4 _u0_U10747  ( .A(1'b1), .ZN(_u0_ch25_csr[17] ) );
INV_X4 _u0_U10745  ( .A(1'b1), .ZN(_u0_ch25_csr[16] ) );
INV_X4 _u0_U10743  ( .A(1'b1), .ZN(_u0_ch25_csr[15] ) );
INV_X4 _u0_U10741  ( .A(1'b1), .ZN(_u0_ch25_csr[14] ) );
INV_X4 _u0_U10739  ( .A(1'b1), .ZN(_u0_ch25_csr[13] ) );
INV_X4 _u0_U10737  ( .A(1'b1), .ZN(_u0_ch25_csr[12] ) );
INV_X4 _u0_U10735  ( .A(1'b1), .ZN(_u0_ch25_csr[11] ) );
INV_X4 _u0_U10733  ( .A(1'b1), .ZN(_u0_ch25_csr[10] ) );
INV_X4 _u0_U10731  ( .A(1'b1), .ZN(_u0_ch25_csr[9] ) );
INV_X4 _u0_U10729  ( .A(1'b1), .ZN(_u0_ch25_csr[8] ) );
INV_X4 _u0_U10727  ( .A(1'b1), .ZN(_u0_ch25_csr[7] ) );
INV_X4 _u0_U10725  ( .A(1'b1), .ZN(_u0_ch25_csr[6] ) );
INV_X4 _u0_U10723  ( .A(1'b1), .ZN(_u0_ch25_csr[5] ) );
INV_X4 _u0_U10721  ( .A(1'b1), .ZN(_u0_ch25_csr[4] ) );
INV_X4 _u0_U10719  ( .A(1'b1), .ZN(_u0_ch25_csr[3] ) );
INV_X4 _u0_U10717  ( .A(1'b1), .ZN(_u0_ch25_csr[2] ) );
INV_X4 _u0_U10715  ( .A(1'b1), .ZN(_u0_ch25_csr[1] ) );
INV_X4 _u0_U10713  ( .A(1'b1), .ZN(_u0_ch25_csr[0] ) );
INV_X4 _u0_U10711  ( .A(1'b1), .ZN(_u0_ch25_txsz[31] ) );
INV_X4 _u0_U10709  ( .A(1'b1), .ZN(_u0_ch25_txsz[30] ) );
INV_X4 _u0_U10707  ( .A(1'b1), .ZN(_u0_ch25_txsz[29] ) );
INV_X4 _u0_U10705  ( .A(1'b1), .ZN(_u0_ch25_txsz[28] ) );
INV_X4 _u0_U10703  ( .A(1'b1), .ZN(_u0_ch25_txsz[27] ) );
INV_X4 _u0_U10701  ( .A(1'b1), .ZN(_u0_ch25_txsz[26] ) );
INV_X4 _u0_U10699  ( .A(1'b1), .ZN(_u0_ch25_txsz[25] ) );
INV_X4 _u0_U10697  ( .A(1'b1), .ZN(_u0_ch25_txsz[24] ) );
INV_X4 _u0_U10695  ( .A(1'b1), .ZN(_u0_ch25_txsz[23] ) );
INV_X4 _u0_U10693  ( .A(1'b1), .ZN(_u0_ch25_txsz[22] ) );
INV_X4 _u0_U10691  ( .A(1'b1), .ZN(_u0_ch25_txsz[21] ) );
INV_X4 _u0_U10689  ( .A(1'b1), .ZN(_u0_ch25_txsz[20] ) );
INV_X4 _u0_U10687  ( .A(1'b1), .ZN(_u0_ch25_txsz[19] ) );
INV_X4 _u0_U10685  ( .A(1'b1), .ZN(_u0_ch25_txsz[18] ) );
INV_X4 _u0_U10683  ( .A(1'b1), .ZN(_u0_ch25_txsz[17] ) );
INV_X4 _u0_U10681  ( .A(1'b1), .ZN(_u0_ch25_txsz[16] ) );
INV_X4 _u0_U10679  ( .A(1'b1), .ZN(_u0_ch25_txsz[15] ) );
INV_X4 _u0_U10677  ( .A(1'b1), .ZN(_u0_ch25_txsz[14] ) );
INV_X4 _u0_U10675  ( .A(1'b1), .ZN(_u0_ch25_txsz[13] ) );
INV_X4 _u0_U10673  ( .A(1'b1), .ZN(_u0_ch25_txsz[12] ) );
INV_X4 _u0_U10671  ( .A(1'b1), .ZN(_u0_ch25_txsz[11] ) );
INV_X4 _u0_U10669  ( .A(1'b1), .ZN(_u0_ch25_txsz[10] ) );
INV_X4 _u0_U10667  ( .A(1'b1), .ZN(_u0_ch25_txsz[9] ) );
INV_X4 _u0_U10665  ( .A(1'b1), .ZN(_u0_ch25_txsz[8] ) );
INV_X4 _u0_U10663  ( .A(1'b1), .ZN(_u0_ch25_txsz[7] ) );
INV_X4 _u0_U10661  ( .A(1'b1), .ZN(_u0_ch25_txsz[6] ) );
INV_X4 _u0_U10659  ( .A(1'b1), .ZN(_u0_ch25_txsz[5] ) );
INV_X4 _u0_U10657  ( .A(1'b1), .ZN(_u0_ch25_txsz[4] ) );
INV_X4 _u0_U10655  ( .A(1'b1), .ZN(_u0_ch25_txsz[3] ) );
INV_X4 _u0_U10653  ( .A(1'b1), .ZN(_u0_ch25_txsz[2] ) );
INV_X4 _u0_U10651  ( .A(1'b1), .ZN(_u0_ch25_txsz[1] ) );
INV_X4 _u0_U10649  ( .A(1'b1), .ZN(_u0_ch25_txsz[0] ) );
INV_X4 _u0_U10647  ( .A(1'b1), .ZN(_u0_ch25_adr0[31] ) );
INV_X4 _u0_U10645  ( .A(1'b1), .ZN(_u0_ch25_adr0[30] ) );
INV_X4 _u0_U10643  ( .A(1'b1), .ZN(_u0_ch25_adr0[29] ) );
INV_X4 _u0_U10641  ( .A(1'b1), .ZN(_u0_ch25_adr0[28] ) );
INV_X4 _u0_U10639  ( .A(1'b1), .ZN(_u0_ch25_adr0[27] ) );
INV_X4 _u0_U10637  ( .A(1'b1), .ZN(_u0_ch25_adr0[26] ) );
INV_X4 _u0_U10635  ( .A(1'b1), .ZN(_u0_ch25_adr0[25] ) );
INV_X4 _u0_U10633  ( .A(1'b1), .ZN(_u0_ch25_adr0[24] ) );
INV_X4 _u0_U10631  ( .A(1'b1), .ZN(_u0_ch25_adr0[23] ) );
INV_X4 _u0_U10629  ( .A(1'b1), .ZN(_u0_ch25_adr0[22] ) );
INV_X4 _u0_U10627  ( .A(1'b1), .ZN(_u0_ch25_adr0[21] ) );
INV_X4 _u0_U10625  ( .A(1'b1), .ZN(_u0_ch25_adr0[20] ) );
INV_X4 _u0_U10623  ( .A(1'b1), .ZN(_u0_ch25_adr0[19] ) );
INV_X4 _u0_U10621  ( .A(1'b1), .ZN(_u0_ch25_adr0[18] ) );
INV_X4 _u0_U10619  ( .A(1'b1), .ZN(_u0_ch25_adr0[17] ) );
INV_X4 _u0_U10617  ( .A(1'b1), .ZN(_u0_ch25_adr0[16] ) );
INV_X4 _u0_U10615  ( .A(1'b1), .ZN(_u0_ch25_adr0[15] ) );
INV_X4 _u0_U10613  ( .A(1'b1), .ZN(_u0_ch25_adr0[14] ) );
INV_X4 _u0_U10611  ( .A(1'b1), .ZN(_u0_ch25_adr0[13] ) );
INV_X4 _u0_U10609  ( .A(1'b1), .ZN(_u0_ch25_adr0[12] ) );
INV_X4 _u0_U10607  ( .A(1'b1), .ZN(_u0_ch25_adr0[11] ) );
INV_X4 _u0_U10605  ( .A(1'b1), .ZN(_u0_ch25_adr0[10] ) );
INV_X4 _u0_U10603  ( .A(1'b1), .ZN(_u0_ch25_adr0[9] ) );
INV_X4 _u0_U10601  ( .A(1'b1), .ZN(_u0_ch25_adr0[8] ) );
INV_X4 _u0_U10599  ( .A(1'b1), .ZN(_u0_ch25_adr0[7] ) );
INV_X4 _u0_U10597  ( .A(1'b1), .ZN(_u0_ch25_adr0[6] ) );
INV_X4 _u0_U10595  ( .A(1'b1), .ZN(_u0_ch25_adr0[5] ) );
INV_X4 _u0_U10593  ( .A(1'b1), .ZN(_u0_ch25_adr0[4] ) );
INV_X4 _u0_U10591  ( .A(1'b1), .ZN(_u0_ch25_adr0[3] ) );
INV_X4 _u0_U10589  ( .A(1'b1), .ZN(_u0_ch25_adr0[2] ) );
INV_X4 _u0_U10587  ( .A(1'b1), .ZN(_u0_ch25_adr0[1] ) );
INV_X4 _u0_U10585  ( .A(1'b1), .ZN(_u0_ch25_adr0[0] ) );
INV_X4 _u0_U10583  ( .A(1'b1), .ZN(_u0_ch25_adr1[31] ) );
INV_X4 _u0_U10581  ( .A(1'b1), .ZN(_u0_ch25_adr1[30] ) );
INV_X4 _u0_U10579  ( .A(1'b1), .ZN(_u0_ch25_adr1[29] ) );
INV_X4 _u0_U10577  ( .A(1'b1), .ZN(_u0_ch25_adr1[28] ) );
INV_X4 _u0_U10575  ( .A(1'b1), .ZN(_u0_ch25_adr1[27] ) );
INV_X4 _u0_U10573  ( .A(1'b1), .ZN(_u0_ch25_adr1[26] ) );
INV_X4 _u0_U10571  ( .A(1'b1), .ZN(_u0_ch25_adr1[25] ) );
INV_X4 _u0_U10569  ( .A(1'b1), .ZN(_u0_ch25_adr1[24] ) );
INV_X4 _u0_U10567  ( .A(1'b1), .ZN(_u0_ch25_adr1[23] ) );
INV_X4 _u0_U10565  ( .A(1'b1), .ZN(_u0_ch25_adr1[22] ) );
INV_X4 _u0_U10563  ( .A(1'b1), .ZN(_u0_ch25_adr1[21] ) );
INV_X4 _u0_U10561  ( .A(1'b1), .ZN(_u0_ch25_adr1[20] ) );
INV_X4 _u0_U10559  ( .A(1'b1), .ZN(_u0_ch25_adr1[19] ) );
INV_X4 _u0_U10557  ( .A(1'b1), .ZN(_u0_ch25_adr1[18] ) );
INV_X4 _u0_U10555  ( .A(1'b1), .ZN(_u0_ch25_adr1[17] ) );
INV_X4 _u0_U10553  ( .A(1'b1), .ZN(_u0_ch25_adr1[16] ) );
INV_X4 _u0_U10551  ( .A(1'b1), .ZN(_u0_ch25_adr1[15] ) );
INV_X4 _u0_U10549  ( .A(1'b1), .ZN(_u0_ch25_adr1[14] ) );
INV_X4 _u0_U10547  ( .A(1'b1), .ZN(_u0_ch25_adr1[13] ) );
INV_X4 _u0_U10545  ( .A(1'b1), .ZN(_u0_ch25_adr1[12] ) );
INV_X4 _u0_U10543  ( .A(1'b1), .ZN(_u0_ch25_adr1[11] ) );
INV_X4 _u0_U10541  ( .A(1'b1), .ZN(_u0_ch25_adr1[10] ) );
INV_X4 _u0_U10539  ( .A(1'b1), .ZN(_u0_ch25_adr1[9] ) );
INV_X4 _u0_U10537  ( .A(1'b1), .ZN(_u0_ch25_adr1[8] ) );
INV_X4 _u0_U10535  ( .A(1'b1), .ZN(_u0_ch25_adr1[7] ) );
INV_X4 _u0_U10533  ( .A(1'b1), .ZN(_u0_ch25_adr1[6] ) );
INV_X4 _u0_U10531  ( .A(1'b1), .ZN(_u0_ch25_adr1[5] ) );
INV_X4 _u0_U10529  ( .A(1'b1), .ZN(_u0_ch25_adr1[4] ) );
INV_X4 _u0_U10527  ( .A(1'b1), .ZN(_u0_ch25_adr1[3] ) );
INV_X4 _u0_U10525  ( .A(1'b1), .ZN(_u0_ch25_adr1[2] ) );
INV_X4 _u0_U10523  ( .A(1'b1), .ZN(_u0_ch25_adr1[1] ) );
INV_X4 _u0_U10521  ( .A(1'b1), .ZN(_u0_ch25_adr1[0] ) );
INV_X4 _u0_U10519  ( .A(1'b0), .ZN(_u0_ch25_am0[31] ) );
INV_X4 _u0_U10517  ( .A(1'b0), .ZN(_u0_ch25_am0[30] ) );
INV_X4 _u0_U10515  ( .A(1'b0), .ZN(_u0_ch25_am0[29] ) );
INV_X4 _u0_U10513  ( .A(1'b0), .ZN(_u0_ch25_am0[28] ) );
INV_X4 _u0_U10511  ( .A(1'b0), .ZN(_u0_ch25_am0[27] ) );
INV_X4 _u0_U10509  ( .A(1'b0), .ZN(_u0_ch25_am0[26] ) );
INV_X4 _u0_U10507  ( .A(1'b0), .ZN(_u0_ch25_am0[25] ) );
INV_X4 _u0_U10505  ( .A(1'b0), .ZN(_u0_ch25_am0[24] ) );
INV_X4 _u0_U10503  ( .A(1'b0), .ZN(_u0_ch25_am0[23] ) );
INV_X4 _u0_U10501  ( .A(1'b0), .ZN(_u0_ch25_am0[22] ) );
INV_X4 _u0_U10499  ( .A(1'b0), .ZN(_u0_ch25_am0[21] ) );
INV_X4 _u0_U10497  ( .A(1'b0), .ZN(_u0_ch25_am0[20] ) );
INV_X4 _u0_U10495  ( .A(1'b0), .ZN(_u0_ch25_am0[19] ) );
INV_X4 _u0_U10493  ( .A(1'b0), .ZN(_u0_ch25_am0[18] ) );
INV_X4 _u0_U10491  ( .A(1'b0), .ZN(_u0_ch25_am0[17] ) );
INV_X4 _u0_U10489  ( .A(1'b0), .ZN(_u0_ch25_am0[16] ) );
INV_X4 _u0_U10487  ( .A(1'b0), .ZN(_u0_ch25_am0[15] ) );
INV_X4 _u0_U10485  ( .A(1'b0), .ZN(_u0_ch25_am0[14] ) );
INV_X4 _u0_U10483  ( .A(1'b0), .ZN(_u0_ch25_am0[13] ) );
INV_X4 _u0_U10481  ( .A(1'b0), .ZN(_u0_ch25_am0[12] ) );
INV_X4 _u0_U10479  ( .A(1'b0), .ZN(_u0_ch25_am0[11] ) );
INV_X4 _u0_U10477  ( .A(1'b0), .ZN(_u0_ch25_am0[10] ) );
INV_X4 _u0_U10475  ( .A(1'b0), .ZN(_u0_ch25_am0[9] ) );
INV_X4 _u0_U10473  ( .A(1'b0), .ZN(_u0_ch25_am0[8] ) );
INV_X4 _u0_U10471  ( .A(1'b0), .ZN(_u0_ch25_am0[7] ) );
INV_X4 _u0_U10469  ( .A(1'b0), .ZN(_u0_ch25_am0[6] ) );
INV_X4 _u0_U10467  ( .A(1'b0), .ZN(_u0_ch25_am0[5] ) );
INV_X4 _u0_U10465  ( .A(1'b0), .ZN(_u0_ch25_am0[4] ) );
INV_X4 _u0_U10463  ( .A(1'b1), .ZN(_u0_ch25_am0[3] ) );
INV_X4 _u0_U10461  ( .A(1'b1), .ZN(_u0_ch25_am0[2] ) );
INV_X4 _u0_U10459  ( .A(1'b1), .ZN(_u0_ch25_am0[1] ) );
INV_X4 _u0_U10457  ( .A(1'b1), .ZN(_u0_ch25_am0[0] ) );
INV_X4 _u0_U10455  ( .A(1'b0), .ZN(_u0_ch25_am1[31] ) );
INV_X4 _u0_U10453  ( .A(1'b0), .ZN(_u0_ch25_am1[30] ) );
INV_X4 _u0_U10451  ( .A(1'b0), .ZN(_u0_ch25_am1[29] ) );
INV_X4 _u0_U10449  ( .A(1'b0), .ZN(_u0_ch25_am1[28] ) );
INV_X4 _u0_U10447  ( .A(1'b0), .ZN(_u0_ch25_am1[27] ) );
INV_X4 _u0_U10445  ( .A(1'b0), .ZN(_u0_ch25_am1[26] ) );
INV_X4 _u0_U10443  ( .A(1'b0), .ZN(_u0_ch25_am1[25] ) );
INV_X4 _u0_U10441  ( .A(1'b0), .ZN(_u0_ch25_am1[24] ) );
INV_X4 _u0_U10439  ( .A(1'b0), .ZN(_u0_ch25_am1[23] ) );
INV_X4 _u0_U10437  ( .A(1'b0), .ZN(_u0_ch25_am1[22] ) );
INV_X4 _u0_U10435  ( .A(1'b0), .ZN(_u0_ch25_am1[21] ) );
INV_X4 _u0_U10433  ( .A(1'b0), .ZN(_u0_ch25_am1[20] ) );
INV_X4 _u0_U10431  ( .A(1'b0), .ZN(_u0_ch25_am1[19] ) );
INV_X4 _u0_U10429  ( .A(1'b0), .ZN(_u0_ch25_am1[18] ) );
INV_X4 _u0_U10427  ( .A(1'b0), .ZN(_u0_ch25_am1[17] ) );
INV_X4 _u0_U10425  ( .A(1'b0), .ZN(_u0_ch25_am1[16] ) );
INV_X4 _u0_U10423  ( .A(1'b0), .ZN(_u0_ch25_am1[15] ) );
INV_X4 _u0_U10421  ( .A(1'b0), .ZN(_u0_ch25_am1[14] ) );
INV_X4 _u0_U10419  ( .A(1'b0), .ZN(_u0_ch25_am1[13] ) );
INV_X4 _u0_U10417  ( .A(1'b0), .ZN(_u0_ch25_am1[12] ) );
INV_X4 _u0_U10415  ( .A(1'b0), .ZN(_u0_ch25_am1[11] ) );
INV_X4 _u0_U10413  ( .A(1'b0), .ZN(_u0_ch25_am1[10] ) );
INV_X4 _u0_U10411  ( .A(1'b0), .ZN(_u0_ch25_am1[9] ) );
INV_X4 _u0_U10409  ( .A(1'b0), .ZN(_u0_ch25_am1[8] ) );
INV_X4 _u0_U10407  ( .A(1'b0), .ZN(_u0_ch25_am1[7] ) );
INV_X4 _u0_U10405  ( .A(1'b0), .ZN(_u0_ch25_am1[6] ) );
INV_X4 _u0_U10403  ( .A(1'b0), .ZN(_u0_ch25_am1[5] ) );
INV_X4 _u0_U10401  ( .A(1'b0), .ZN(_u0_ch25_am1[4] ) );
INV_X4 _u0_U10399  ( .A(1'b1), .ZN(_u0_ch25_am1[3] ) );
INV_X4 _u0_U10397  ( .A(1'b1), .ZN(_u0_ch25_am1[2] ) );
INV_X4 _u0_U10395  ( .A(1'b1), .ZN(_u0_ch25_am1[1] ) );
INV_X4 _u0_U10393  ( .A(1'b1), .ZN(_u0_ch25_am1[0] ) );
INV_X4 _u0_U10391  ( .A(1'b1), .ZN(_u0_pointer26[31] ) );
INV_X4 _u0_U10389  ( .A(1'b1), .ZN(_u0_pointer26[30] ) );
INV_X4 _u0_U10387  ( .A(1'b1), .ZN(_u0_pointer26[29] ) );
INV_X4 _u0_U10385  ( .A(1'b1), .ZN(_u0_pointer26[28] ) );
INV_X4 _u0_U10383  ( .A(1'b1), .ZN(_u0_pointer26[27] ) );
INV_X4 _u0_U10381  ( .A(1'b1), .ZN(_u0_pointer26[26] ) );
INV_X4 _u0_U10379  ( .A(1'b1), .ZN(_u0_pointer26[25] ) );
INV_X4 _u0_U10377  ( .A(1'b1), .ZN(_u0_pointer26[24] ) );
INV_X4 _u0_U10375  ( .A(1'b1), .ZN(_u0_pointer26[23] ) );
INV_X4 _u0_U10373  ( .A(1'b1), .ZN(_u0_pointer26[22] ) );
INV_X4 _u0_U10371  ( .A(1'b1), .ZN(_u0_pointer26[21] ) );
INV_X4 _u0_U10369  ( .A(1'b1), .ZN(_u0_pointer26[20] ) );
INV_X4 _u0_U10367  ( .A(1'b1), .ZN(_u0_pointer26[19] ) );
INV_X4 _u0_U10365  ( .A(1'b1), .ZN(_u0_pointer26[18] ) );
INV_X4 _u0_U10363  ( .A(1'b1), .ZN(_u0_pointer26[17] ) );
INV_X4 _u0_U10361  ( .A(1'b1), .ZN(_u0_pointer26[16] ) );
INV_X4 _u0_U10359  ( .A(1'b1), .ZN(_u0_pointer26[15] ) );
INV_X4 _u0_U10357  ( .A(1'b1), .ZN(_u0_pointer26[14] ) );
INV_X4 _u0_U10355  ( .A(1'b1), .ZN(_u0_pointer26[13] ) );
INV_X4 _u0_U10353  ( .A(1'b1), .ZN(_u0_pointer26[12] ) );
INV_X4 _u0_U10351  ( .A(1'b1), .ZN(_u0_pointer26[11] ) );
INV_X4 _u0_U10349  ( .A(1'b1), .ZN(_u0_pointer26[10] ) );
INV_X4 _u0_U10347  ( .A(1'b1), .ZN(_u0_pointer26[9] ) );
INV_X4 _u0_U10345  ( .A(1'b1), .ZN(_u0_pointer26[8] ) );
INV_X4 _u0_U10343  ( .A(1'b1), .ZN(_u0_pointer26[7] ) );
INV_X4 _u0_U10341  ( .A(1'b1), .ZN(_u0_pointer26[6] ) );
INV_X4 _u0_U10339  ( .A(1'b1), .ZN(_u0_pointer26[5] ) );
INV_X4 _u0_U10337  ( .A(1'b1), .ZN(_u0_pointer26[4] ) );
INV_X4 _u0_U10335  ( .A(1'b1), .ZN(_u0_pointer26[3] ) );
INV_X4 _u0_U10333  ( .A(1'b1), .ZN(_u0_pointer26[2] ) );
INV_X4 _u0_U10331  ( .A(1'b1), .ZN(_u0_pointer26[1] ) );
INV_X4 _u0_U10329  ( .A(1'b1), .ZN(_u0_pointer26[0] ) );
INV_X4 _u0_U10327  ( .A(1'b1), .ZN(_u0_pointer26_s[31] ) );
INV_X4 _u0_U10325  ( .A(1'b1), .ZN(_u0_pointer26_s[30] ) );
INV_X4 _u0_U10323  ( .A(1'b1), .ZN(_u0_pointer26_s[29] ) );
INV_X4 _u0_U10321  ( .A(1'b1), .ZN(_u0_pointer26_s[28] ) );
INV_X4 _u0_U10319  ( .A(1'b1), .ZN(_u0_pointer26_s[27] ) );
INV_X4 _u0_U10317  ( .A(1'b1), .ZN(_u0_pointer26_s[26] ) );
INV_X4 _u0_U10315  ( .A(1'b1), .ZN(_u0_pointer26_s[25] ) );
INV_X4 _u0_U10313  ( .A(1'b1), .ZN(_u0_pointer26_s[24] ) );
INV_X4 _u0_U10311  ( .A(1'b1), .ZN(_u0_pointer26_s[23] ) );
INV_X4 _u0_U10309  ( .A(1'b1), .ZN(_u0_pointer26_s[22] ) );
INV_X4 _u0_U10307  ( .A(1'b1), .ZN(_u0_pointer26_s[21] ) );
INV_X4 _u0_U10305  ( .A(1'b1), .ZN(_u0_pointer26_s[20] ) );
INV_X4 _u0_U10303  ( .A(1'b1), .ZN(_u0_pointer26_s[19] ) );
INV_X4 _u0_U10301  ( .A(1'b1), .ZN(_u0_pointer26_s[18] ) );
INV_X4 _u0_U10299  ( .A(1'b1), .ZN(_u0_pointer26_s[17] ) );
INV_X4 _u0_U10297  ( .A(1'b1), .ZN(_u0_pointer26_s[16] ) );
INV_X4 _u0_U10295  ( .A(1'b1), .ZN(_u0_pointer26_s[15] ) );
INV_X4 _u0_U10293  ( .A(1'b1), .ZN(_u0_pointer26_s[14] ) );
INV_X4 _u0_U10291  ( .A(1'b1), .ZN(_u0_pointer26_s[13] ) );
INV_X4 _u0_U10289  ( .A(1'b1), .ZN(_u0_pointer26_s[12] ) );
INV_X4 _u0_U10287  ( .A(1'b1), .ZN(_u0_pointer26_s[11] ) );
INV_X4 _u0_U10285  ( .A(1'b1), .ZN(_u0_pointer26_s[10] ) );
INV_X4 _u0_U10283  ( .A(1'b1), .ZN(_u0_pointer26_s[9] ) );
INV_X4 _u0_U10281  ( .A(1'b1), .ZN(_u0_pointer26_s[8] ) );
INV_X4 _u0_U10279  ( .A(1'b1), .ZN(_u0_pointer26_s[7] ) );
INV_X4 _u0_U10277  ( .A(1'b1), .ZN(_u0_pointer26_s[6] ) );
INV_X4 _u0_U10275  ( .A(1'b1), .ZN(_u0_pointer26_s[5] ) );
INV_X4 _u0_U10273  ( .A(1'b1), .ZN(_u0_pointer26_s[4] ) );
INV_X4 _u0_U10271  ( .A(1'b1), .ZN(_u0_pointer26_s[3] ) );
INV_X4 _u0_U10269  ( .A(1'b1), .ZN(_u0_pointer26_s[2] ) );
INV_X4 _u0_U10267  ( .A(1'b1), .ZN(_u0_pointer26_s[1] ) );
INV_X4 _u0_U10265  ( .A(1'b1), .ZN(_u0_pointer26_s[0] ) );
INV_X4 _u0_U10263  ( .A(1'b1), .ZN(_u0_ch26_csr[31] ) );
INV_X4 _u0_U10261  ( .A(1'b1), .ZN(_u0_ch26_csr[30] ) );
INV_X4 _u0_U10259  ( .A(1'b1), .ZN(_u0_ch26_csr[29] ) );
INV_X4 _u0_U10257  ( .A(1'b1), .ZN(_u0_ch26_csr[28] ) );
INV_X4 _u0_U10255  ( .A(1'b1), .ZN(_u0_ch26_csr[27] ) );
INV_X4 _u0_U10253  ( .A(1'b1), .ZN(_u0_ch26_csr[26] ) );
INV_X4 _u0_U10251  ( .A(1'b1), .ZN(_u0_ch26_csr[25] ) );
INV_X4 _u0_U10249  ( .A(1'b1), .ZN(_u0_ch26_csr[24] ) );
INV_X4 _u0_U10247  ( .A(1'b1), .ZN(_u0_ch26_csr[23] ) );
INV_X4 _u0_U10245  ( .A(1'b1), .ZN(_u0_ch26_csr[22] ) );
INV_X4 _u0_U10243  ( .A(1'b1), .ZN(_u0_ch26_csr[21] ) );
INV_X4 _u0_U10241  ( .A(1'b1), .ZN(_u0_ch26_csr[20] ) );
INV_X4 _u0_U10239  ( .A(1'b1), .ZN(_u0_ch26_csr[19] ) );
INV_X4 _u0_U10237  ( .A(1'b1), .ZN(_u0_ch26_csr[18] ) );
INV_X4 _u0_U10235  ( .A(1'b1), .ZN(_u0_ch26_csr[17] ) );
INV_X4 _u0_U10233  ( .A(1'b1), .ZN(_u0_ch26_csr[16] ) );
INV_X4 _u0_U10231  ( .A(1'b1), .ZN(_u0_ch26_csr[15] ) );
INV_X4 _u0_U10229  ( .A(1'b1), .ZN(_u0_ch26_csr[14] ) );
INV_X4 _u0_U10227  ( .A(1'b1), .ZN(_u0_ch26_csr[13] ) );
INV_X4 _u0_U10225  ( .A(1'b1), .ZN(_u0_ch26_csr[12] ) );
INV_X4 _u0_U10223  ( .A(1'b1), .ZN(_u0_ch26_csr[11] ) );
INV_X4 _u0_U10221  ( .A(1'b1), .ZN(_u0_ch26_csr[10] ) );
INV_X4 _u0_U10219  ( .A(1'b1), .ZN(_u0_ch26_csr[9] ) );
INV_X4 _u0_U10217  ( .A(1'b1), .ZN(_u0_ch26_csr[8] ) );
INV_X4 _u0_U10215  ( .A(1'b1), .ZN(_u0_ch26_csr[7] ) );
INV_X4 _u0_U10213  ( .A(1'b1), .ZN(_u0_ch26_csr[6] ) );
INV_X4 _u0_U10211  ( .A(1'b1), .ZN(_u0_ch26_csr[5] ) );
INV_X4 _u0_U10209  ( .A(1'b1), .ZN(_u0_ch26_csr[4] ) );
INV_X4 _u0_U10207  ( .A(1'b1), .ZN(_u0_ch26_csr[3] ) );
INV_X4 _u0_U10205  ( .A(1'b1), .ZN(_u0_ch26_csr[2] ) );
INV_X4 _u0_U10203  ( .A(1'b1), .ZN(_u0_ch26_csr[1] ) );
INV_X4 _u0_U10201  ( .A(1'b1), .ZN(_u0_ch26_csr[0] ) );
INV_X4 _u0_U10199  ( .A(1'b1), .ZN(_u0_ch26_txsz[31] ) );
INV_X4 _u0_U10197  ( .A(1'b1), .ZN(_u0_ch26_txsz[30] ) );
INV_X4 _u0_U10195  ( .A(1'b1), .ZN(_u0_ch26_txsz[29] ) );
INV_X4 _u0_U10193  ( .A(1'b1), .ZN(_u0_ch26_txsz[28] ) );
INV_X4 _u0_U10191  ( .A(1'b1), .ZN(_u0_ch26_txsz[27] ) );
INV_X4 _u0_U10189  ( .A(1'b1), .ZN(_u0_ch26_txsz[26] ) );
INV_X4 _u0_U10187  ( .A(1'b1), .ZN(_u0_ch26_txsz[25] ) );
INV_X4 _u0_U10185  ( .A(1'b1), .ZN(_u0_ch26_txsz[24] ) );
INV_X4 _u0_U10183  ( .A(1'b1), .ZN(_u0_ch26_txsz[23] ) );
INV_X4 _u0_U10181  ( .A(1'b1), .ZN(_u0_ch26_txsz[22] ) );
INV_X4 _u0_U10179  ( .A(1'b1), .ZN(_u0_ch26_txsz[21] ) );
INV_X4 _u0_U10177  ( .A(1'b1), .ZN(_u0_ch26_txsz[20] ) );
INV_X4 _u0_U10175  ( .A(1'b1), .ZN(_u0_ch26_txsz[19] ) );
INV_X4 _u0_U10173  ( .A(1'b1), .ZN(_u0_ch26_txsz[18] ) );
INV_X4 _u0_U10171  ( .A(1'b1), .ZN(_u0_ch26_txsz[17] ) );
INV_X4 _u0_U10169  ( .A(1'b1), .ZN(_u0_ch26_txsz[16] ) );
INV_X4 _u0_U10167  ( .A(1'b1), .ZN(_u0_ch26_txsz[15] ) );
INV_X4 _u0_U10165  ( .A(1'b1), .ZN(_u0_ch26_txsz[14] ) );
INV_X4 _u0_U10163  ( .A(1'b1), .ZN(_u0_ch26_txsz[13] ) );
INV_X4 _u0_U10161  ( .A(1'b1), .ZN(_u0_ch26_txsz[12] ) );
INV_X4 _u0_U10159  ( .A(1'b1), .ZN(_u0_ch26_txsz[11] ) );
INV_X4 _u0_U10157  ( .A(1'b1), .ZN(_u0_ch26_txsz[10] ) );
INV_X4 _u0_U10155  ( .A(1'b1), .ZN(_u0_ch26_txsz[9] ) );
INV_X4 _u0_U10153  ( .A(1'b1), .ZN(_u0_ch26_txsz[8] ) );
INV_X4 _u0_U10151  ( .A(1'b1), .ZN(_u0_ch26_txsz[7] ) );
INV_X4 _u0_U10149  ( .A(1'b1), .ZN(_u0_ch26_txsz[6] ) );
INV_X4 _u0_U10147  ( .A(1'b1), .ZN(_u0_ch26_txsz[5] ) );
INV_X4 _u0_U10145  ( .A(1'b1), .ZN(_u0_ch26_txsz[4] ) );
INV_X4 _u0_U10143  ( .A(1'b1), .ZN(_u0_ch26_txsz[3] ) );
INV_X4 _u0_U10141  ( .A(1'b1), .ZN(_u0_ch26_txsz[2] ) );
INV_X4 _u0_U10139  ( .A(1'b1), .ZN(_u0_ch26_txsz[1] ) );
INV_X4 _u0_U10137  ( .A(1'b1), .ZN(_u0_ch26_txsz[0] ) );
INV_X4 _u0_U10135  ( .A(1'b1), .ZN(_u0_ch26_adr0[31] ) );
INV_X4 _u0_U10133  ( .A(1'b1), .ZN(_u0_ch26_adr0[30] ) );
INV_X4 _u0_U10131  ( .A(1'b1), .ZN(_u0_ch26_adr0[29] ) );
INV_X4 _u0_U10129  ( .A(1'b1), .ZN(_u0_ch26_adr0[28] ) );
INV_X4 _u0_U10127  ( .A(1'b1), .ZN(_u0_ch26_adr0[27] ) );
INV_X4 _u0_U10125  ( .A(1'b1), .ZN(_u0_ch26_adr0[26] ) );
INV_X4 _u0_U10123  ( .A(1'b1), .ZN(_u0_ch26_adr0[25] ) );
INV_X4 _u0_U10121  ( .A(1'b1), .ZN(_u0_ch26_adr0[24] ) );
INV_X4 _u0_U10119  ( .A(1'b1), .ZN(_u0_ch26_adr0[23] ) );
INV_X4 _u0_U10117  ( .A(1'b1), .ZN(_u0_ch26_adr0[22] ) );
INV_X4 _u0_U10115  ( .A(1'b1), .ZN(_u0_ch26_adr0[21] ) );
INV_X4 _u0_U10113  ( .A(1'b1), .ZN(_u0_ch26_adr0[20] ) );
INV_X4 _u0_U10111  ( .A(1'b1), .ZN(_u0_ch26_adr0[19] ) );
INV_X4 _u0_U10109  ( .A(1'b1), .ZN(_u0_ch26_adr0[18] ) );
INV_X4 _u0_U10107  ( .A(1'b1), .ZN(_u0_ch26_adr0[17] ) );
INV_X4 _u0_U10105  ( .A(1'b1), .ZN(_u0_ch26_adr0[16] ) );
INV_X4 _u0_U10103  ( .A(1'b1), .ZN(_u0_ch26_adr0[15] ) );
INV_X4 _u0_U10101  ( .A(1'b1), .ZN(_u0_ch26_adr0[14] ) );
INV_X4 _u0_U10099  ( .A(1'b1), .ZN(_u0_ch26_adr0[13] ) );
INV_X4 _u0_U10097  ( .A(1'b1), .ZN(_u0_ch26_adr0[12] ) );
INV_X4 _u0_U10095  ( .A(1'b1), .ZN(_u0_ch26_adr0[11] ) );
INV_X4 _u0_U10093  ( .A(1'b1), .ZN(_u0_ch26_adr0[10] ) );
INV_X4 _u0_U10091  ( .A(1'b1), .ZN(_u0_ch26_adr0[9] ) );
INV_X4 _u0_U10089  ( .A(1'b1), .ZN(_u0_ch26_adr0[8] ) );
INV_X4 _u0_U10087  ( .A(1'b1), .ZN(_u0_ch26_adr0[7] ) );
INV_X4 _u0_U10085  ( .A(1'b1), .ZN(_u0_ch26_adr0[6] ) );
INV_X4 _u0_U10083  ( .A(1'b1), .ZN(_u0_ch26_adr0[5] ) );
INV_X4 _u0_U10081  ( .A(1'b1), .ZN(_u0_ch26_adr0[4] ) );
INV_X4 _u0_U10079  ( .A(1'b1), .ZN(_u0_ch26_adr0[3] ) );
INV_X4 _u0_U10077  ( .A(1'b1), .ZN(_u0_ch26_adr0[2] ) );
INV_X4 _u0_U10075  ( .A(1'b1), .ZN(_u0_ch26_adr0[1] ) );
INV_X4 _u0_U10073  ( .A(1'b1), .ZN(_u0_ch26_adr0[0] ) );
INV_X4 _u0_U10071  ( .A(1'b1), .ZN(_u0_ch26_adr1[31] ) );
INV_X4 _u0_U10069  ( .A(1'b1), .ZN(_u0_ch26_adr1[30] ) );
INV_X4 _u0_U10067  ( .A(1'b1), .ZN(_u0_ch26_adr1[29] ) );
INV_X4 _u0_U10065  ( .A(1'b1), .ZN(_u0_ch26_adr1[28] ) );
INV_X4 _u0_U10063  ( .A(1'b1), .ZN(_u0_ch26_adr1[27] ) );
INV_X4 _u0_U10061  ( .A(1'b1), .ZN(_u0_ch26_adr1[26] ) );
INV_X4 _u0_U10059  ( .A(1'b1), .ZN(_u0_ch26_adr1[25] ) );
INV_X4 _u0_U10057  ( .A(1'b1), .ZN(_u0_ch26_adr1[24] ) );
INV_X4 _u0_U10055  ( .A(1'b1), .ZN(_u0_ch26_adr1[23] ) );
INV_X4 _u0_U10053  ( .A(1'b1), .ZN(_u0_ch26_adr1[22] ) );
INV_X4 _u0_U10051  ( .A(1'b1), .ZN(_u0_ch26_adr1[21] ) );
INV_X4 _u0_U10049  ( .A(1'b1), .ZN(_u0_ch26_adr1[20] ) );
INV_X4 _u0_U10047  ( .A(1'b1), .ZN(_u0_ch26_adr1[19] ) );
INV_X4 _u0_U10045  ( .A(1'b1), .ZN(_u0_ch26_adr1[18] ) );
INV_X4 _u0_U10043  ( .A(1'b1), .ZN(_u0_ch26_adr1[17] ) );
INV_X4 _u0_U10041  ( .A(1'b1), .ZN(_u0_ch26_adr1[16] ) );
INV_X4 _u0_U10039  ( .A(1'b1), .ZN(_u0_ch26_adr1[15] ) );
INV_X4 _u0_U10037  ( .A(1'b1), .ZN(_u0_ch26_adr1[14] ) );
INV_X4 _u0_U10035  ( .A(1'b1), .ZN(_u0_ch26_adr1[13] ) );
INV_X4 _u0_U10033  ( .A(1'b1), .ZN(_u0_ch26_adr1[12] ) );
INV_X4 _u0_U10031  ( .A(1'b1), .ZN(_u0_ch26_adr1[11] ) );
INV_X4 _u0_U10029  ( .A(1'b1), .ZN(_u0_ch26_adr1[10] ) );
INV_X4 _u0_U10027  ( .A(1'b1), .ZN(_u0_ch26_adr1[9] ) );
INV_X4 _u0_U10025  ( .A(1'b1), .ZN(_u0_ch26_adr1[8] ) );
INV_X4 _u0_U10023  ( .A(1'b1), .ZN(_u0_ch26_adr1[7] ) );
INV_X4 _u0_U10021  ( .A(1'b1), .ZN(_u0_ch26_adr1[6] ) );
INV_X4 _u0_U10019  ( .A(1'b1), .ZN(_u0_ch26_adr1[5] ) );
INV_X4 _u0_U10017  ( .A(1'b1), .ZN(_u0_ch26_adr1[4] ) );
INV_X4 _u0_U10015  ( .A(1'b1), .ZN(_u0_ch26_adr1[3] ) );
INV_X4 _u0_U10013  ( .A(1'b1), .ZN(_u0_ch26_adr1[2] ) );
INV_X4 _u0_U10011  ( .A(1'b1), .ZN(_u0_ch26_adr1[1] ) );
INV_X4 _u0_U10009  ( .A(1'b1), .ZN(_u0_ch26_adr1[0] ) );
INV_X4 _u0_U10007  ( .A(1'b0), .ZN(_u0_ch26_am0[31] ) );
INV_X4 _u0_U10005  ( .A(1'b0), .ZN(_u0_ch26_am0[30] ) );
INV_X4 _u0_U10003  ( .A(1'b0), .ZN(_u0_ch26_am0[29] ) );
INV_X4 _u0_U10001  ( .A(1'b0), .ZN(_u0_ch26_am0[28] ) );
INV_X4 _u0_U9999  ( .A(1'b0), .ZN(_u0_ch26_am0[27] ) );
INV_X4 _u0_U9997  ( .A(1'b0), .ZN(_u0_ch26_am0[26] ) );
INV_X4 _u0_U9995  ( .A(1'b0), .ZN(_u0_ch26_am0[25] ) );
INV_X4 _u0_U9993  ( .A(1'b0), .ZN(_u0_ch26_am0[24] ) );
INV_X4 _u0_U9991  ( .A(1'b0), .ZN(_u0_ch26_am0[23] ) );
INV_X4 _u0_U9989  ( .A(1'b0), .ZN(_u0_ch26_am0[22] ) );
INV_X4 _u0_U9987  ( .A(1'b0), .ZN(_u0_ch26_am0[21] ) );
INV_X4 _u0_U9985  ( .A(1'b0), .ZN(_u0_ch26_am0[20] ) );
INV_X4 _u0_U9983  ( .A(1'b0), .ZN(_u0_ch26_am0[19] ) );
INV_X4 _u0_U9981  ( .A(1'b0), .ZN(_u0_ch26_am0[18] ) );
INV_X4 _u0_U9979  ( .A(1'b0), .ZN(_u0_ch26_am0[17] ) );
INV_X4 _u0_U9977  ( .A(1'b0), .ZN(_u0_ch26_am0[16] ) );
INV_X4 _u0_U9975  ( .A(1'b0), .ZN(_u0_ch26_am0[15] ) );
INV_X4 _u0_U9973  ( .A(1'b0), .ZN(_u0_ch26_am0[14] ) );
INV_X4 _u0_U9971  ( .A(1'b0), .ZN(_u0_ch26_am0[13] ) );
INV_X4 _u0_U9969  ( .A(1'b0), .ZN(_u0_ch26_am0[12] ) );
INV_X4 _u0_U9967  ( .A(1'b0), .ZN(_u0_ch26_am0[11] ) );
INV_X4 _u0_U9965  ( .A(1'b0), .ZN(_u0_ch26_am0[10] ) );
INV_X4 _u0_U9963  ( .A(1'b0), .ZN(_u0_ch26_am0[9] ) );
INV_X4 _u0_U9961  ( .A(1'b0), .ZN(_u0_ch26_am0[8] ) );
INV_X4 _u0_U9959  ( .A(1'b0), .ZN(_u0_ch26_am0[7] ) );
INV_X4 _u0_U9957  ( .A(1'b0), .ZN(_u0_ch26_am0[6] ) );
INV_X4 _u0_U9955  ( .A(1'b0), .ZN(_u0_ch26_am0[5] ) );
INV_X4 _u0_U9953  ( .A(1'b0), .ZN(_u0_ch26_am0[4] ) );
INV_X4 _u0_U9951  ( .A(1'b1), .ZN(_u0_ch26_am0[3] ) );
INV_X4 _u0_U9949  ( .A(1'b1), .ZN(_u0_ch26_am0[2] ) );
INV_X4 _u0_U9947  ( .A(1'b1), .ZN(_u0_ch26_am0[1] ) );
INV_X4 _u0_U9945  ( .A(1'b1), .ZN(_u0_ch26_am0[0] ) );
INV_X4 _u0_U9943  ( .A(1'b0), .ZN(_u0_ch26_am1[31] ) );
INV_X4 _u0_U9941  ( .A(1'b0), .ZN(_u0_ch26_am1[30] ) );
INV_X4 _u0_U9939  ( .A(1'b0), .ZN(_u0_ch26_am1[29] ) );
INV_X4 _u0_U9937  ( .A(1'b0), .ZN(_u0_ch26_am1[28] ) );
INV_X4 _u0_U9935  ( .A(1'b0), .ZN(_u0_ch26_am1[27] ) );
INV_X4 _u0_U9933  ( .A(1'b0), .ZN(_u0_ch26_am1[26] ) );
INV_X4 _u0_U9931  ( .A(1'b0), .ZN(_u0_ch26_am1[25] ) );
INV_X4 _u0_U9929  ( .A(1'b0), .ZN(_u0_ch26_am1[24] ) );
INV_X4 _u0_U9927  ( .A(1'b0), .ZN(_u0_ch26_am1[23] ) );
INV_X4 _u0_U9925  ( .A(1'b0), .ZN(_u0_ch26_am1[22] ) );
INV_X4 _u0_U9923  ( .A(1'b0), .ZN(_u0_ch26_am1[21] ) );
INV_X4 _u0_U9921  ( .A(1'b0), .ZN(_u0_ch26_am1[20] ) );
INV_X4 _u0_U9919  ( .A(1'b0), .ZN(_u0_ch26_am1[19] ) );
INV_X4 _u0_U9917  ( .A(1'b0), .ZN(_u0_ch26_am1[18] ) );
INV_X4 _u0_U9915  ( .A(1'b0), .ZN(_u0_ch26_am1[17] ) );
INV_X4 _u0_U9913  ( .A(1'b0), .ZN(_u0_ch26_am1[16] ) );
INV_X4 _u0_U9911  ( .A(1'b0), .ZN(_u0_ch26_am1[15] ) );
INV_X4 _u0_U9909  ( .A(1'b0), .ZN(_u0_ch26_am1[14] ) );
INV_X4 _u0_U9907  ( .A(1'b0), .ZN(_u0_ch26_am1[13] ) );
INV_X4 _u0_U9905  ( .A(1'b0), .ZN(_u0_ch26_am1[12] ) );
INV_X4 _u0_U9903  ( .A(1'b0), .ZN(_u0_ch26_am1[11] ) );
INV_X4 _u0_U9901  ( .A(1'b0), .ZN(_u0_ch26_am1[10] ) );
INV_X4 _u0_U9899  ( .A(1'b0), .ZN(_u0_ch26_am1[9] ) );
INV_X4 _u0_U9897  ( .A(1'b0), .ZN(_u0_ch26_am1[8] ) );
INV_X4 _u0_U9895  ( .A(1'b0), .ZN(_u0_ch26_am1[7] ) );
INV_X4 _u0_U9893  ( .A(1'b0), .ZN(_u0_ch26_am1[6] ) );
INV_X4 _u0_U9891  ( .A(1'b0), .ZN(_u0_ch26_am1[5] ) );
INV_X4 _u0_U9889  ( .A(1'b0), .ZN(_u0_ch26_am1[4] ) );
INV_X4 _u0_U9887  ( .A(1'b1), .ZN(_u0_ch26_am1[3] ) );
INV_X4 _u0_U9885  ( .A(1'b1), .ZN(_u0_ch26_am1[2] ) );
INV_X4 _u0_U9883  ( .A(1'b1), .ZN(_u0_ch26_am1[1] ) );
INV_X4 _u0_U9881  ( .A(1'b1), .ZN(_u0_ch26_am1[0] ) );
INV_X4 _u0_U9879  ( .A(1'b1), .ZN(_u0_pointer27[31] ) );
INV_X4 _u0_U9877  ( .A(1'b1), .ZN(_u0_pointer27[30] ) );
INV_X4 _u0_U9875  ( .A(1'b1), .ZN(_u0_pointer27[29] ) );
INV_X4 _u0_U9873  ( .A(1'b1), .ZN(_u0_pointer27[28] ) );
INV_X4 _u0_U9871  ( .A(1'b1), .ZN(_u0_pointer27[27] ) );
INV_X4 _u0_U9869  ( .A(1'b1), .ZN(_u0_pointer27[26] ) );
INV_X4 _u0_U9867  ( .A(1'b1), .ZN(_u0_pointer27[25] ) );
INV_X4 _u0_U9865  ( .A(1'b1), .ZN(_u0_pointer27[24] ) );
INV_X4 _u0_U9863  ( .A(1'b1), .ZN(_u0_pointer27[23] ) );
INV_X4 _u0_U9861  ( .A(1'b1), .ZN(_u0_pointer27[22] ) );
INV_X4 _u0_U9859  ( .A(1'b1), .ZN(_u0_pointer27[21] ) );
INV_X4 _u0_U9857  ( .A(1'b1), .ZN(_u0_pointer27[20] ) );
INV_X4 _u0_U9855  ( .A(1'b1), .ZN(_u0_pointer27[19] ) );
INV_X4 _u0_U9853  ( .A(1'b1), .ZN(_u0_pointer27[18] ) );
INV_X4 _u0_U9851  ( .A(1'b1), .ZN(_u0_pointer27[17] ) );
INV_X4 _u0_U9849  ( .A(1'b1), .ZN(_u0_pointer27[16] ) );
INV_X4 _u0_U9847  ( .A(1'b1), .ZN(_u0_pointer27[15] ) );
INV_X4 _u0_U9845  ( .A(1'b1), .ZN(_u0_pointer27[14] ) );
INV_X4 _u0_U9843  ( .A(1'b1), .ZN(_u0_pointer27[13] ) );
INV_X4 _u0_U9841  ( .A(1'b1), .ZN(_u0_pointer27[12] ) );
INV_X4 _u0_U9839  ( .A(1'b1), .ZN(_u0_pointer27[11] ) );
INV_X4 _u0_U9837  ( .A(1'b1), .ZN(_u0_pointer27[10] ) );
INV_X4 _u0_U9835  ( .A(1'b1), .ZN(_u0_pointer27[9] ) );
INV_X4 _u0_U9833  ( .A(1'b1), .ZN(_u0_pointer27[8] ) );
INV_X4 _u0_U9831  ( .A(1'b1), .ZN(_u0_pointer27[7] ) );
INV_X4 _u0_U9829  ( .A(1'b1), .ZN(_u0_pointer27[6] ) );
INV_X4 _u0_U9827  ( .A(1'b1), .ZN(_u0_pointer27[5] ) );
INV_X4 _u0_U9825  ( .A(1'b1), .ZN(_u0_pointer27[4] ) );
INV_X4 _u0_U9823  ( .A(1'b1), .ZN(_u0_pointer27[3] ) );
INV_X4 _u0_U9821  ( .A(1'b1), .ZN(_u0_pointer27[2] ) );
INV_X4 _u0_U9819  ( .A(1'b1), .ZN(_u0_pointer27[1] ) );
INV_X4 _u0_U9817  ( .A(1'b1), .ZN(_u0_pointer27[0] ) );
INV_X4 _u0_U9815  ( .A(1'b1), .ZN(_u0_pointer27_s[31] ) );
INV_X4 _u0_U9813  ( .A(1'b1), .ZN(_u0_pointer27_s[30] ) );
INV_X4 _u0_U9811  ( .A(1'b1), .ZN(_u0_pointer27_s[29] ) );
INV_X4 _u0_U9809  ( .A(1'b1), .ZN(_u0_pointer27_s[28] ) );
INV_X4 _u0_U9807  ( .A(1'b1), .ZN(_u0_pointer27_s[27] ) );
INV_X4 _u0_U9805  ( .A(1'b1), .ZN(_u0_pointer27_s[26] ) );
INV_X4 _u0_U9803  ( .A(1'b1), .ZN(_u0_pointer27_s[25] ) );
INV_X4 _u0_U9801  ( .A(1'b1), .ZN(_u0_pointer27_s[24] ) );
INV_X4 _u0_U9799  ( .A(1'b1), .ZN(_u0_pointer27_s[23] ) );
INV_X4 _u0_U9797  ( .A(1'b1), .ZN(_u0_pointer27_s[22] ) );
INV_X4 _u0_U9795  ( .A(1'b1), .ZN(_u0_pointer27_s[21] ) );
INV_X4 _u0_U9793  ( .A(1'b1), .ZN(_u0_pointer27_s[20] ) );
INV_X4 _u0_U9791  ( .A(1'b1), .ZN(_u0_pointer27_s[19] ) );
INV_X4 _u0_U9789  ( .A(1'b1), .ZN(_u0_pointer27_s[18] ) );
INV_X4 _u0_U9787  ( .A(1'b1), .ZN(_u0_pointer27_s[17] ) );
INV_X4 _u0_U9785  ( .A(1'b1), .ZN(_u0_pointer27_s[16] ) );
INV_X4 _u0_U9783  ( .A(1'b1), .ZN(_u0_pointer27_s[15] ) );
INV_X4 _u0_U9781  ( .A(1'b1), .ZN(_u0_pointer27_s[14] ) );
INV_X4 _u0_U9779  ( .A(1'b1), .ZN(_u0_pointer27_s[13] ) );
INV_X4 _u0_U9777  ( .A(1'b1), .ZN(_u0_pointer27_s[12] ) );
INV_X4 _u0_U9775  ( .A(1'b1), .ZN(_u0_pointer27_s[11] ) );
INV_X4 _u0_U9773  ( .A(1'b1), .ZN(_u0_pointer27_s[10] ) );
INV_X4 _u0_U9771  ( .A(1'b1), .ZN(_u0_pointer27_s[9] ) );
INV_X4 _u0_U9769  ( .A(1'b1), .ZN(_u0_pointer27_s[8] ) );
INV_X4 _u0_U9767  ( .A(1'b1), .ZN(_u0_pointer27_s[7] ) );
INV_X4 _u0_U9765  ( .A(1'b1), .ZN(_u0_pointer27_s[6] ) );
INV_X4 _u0_U9763  ( .A(1'b1), .ZN(_u0_pointer27_s[5] ) );
INV_X4 _u0_U9761  ( .A(1'b1), .ZN(_u0_pointer27_s[4] ) );
INV_X4 _u0_U9759  ( .A(1'b1), .ZN(_u0_pointer27_s[3] ) );
INV_X4 _u0_U9757  ( .A(1'b1), .ZN(_u0_pointer27_s[2] ) );
INV_X4 _u0_U9755  ( .A(1'b1), .ZN(_u0_pointer27_s[1] ) );
INV_X4 _u0_U9753  ( .A(1'b1), .ZN(_u0_pointer27_s[0] ) );
INV_X4 _u0_U9751  ( .A(1'b1), .ZN(_u0_ch27_csr[31] ) );
INV_X4 _u0_U9749  ( .A(1'b1), .ZN(_u0_ch27_csr[30] ) );
INV_X4 _u0_U9747  ( .A(1'b1), .ZN(_u0_ch27_csr[29] ) );
INV_X4 _u0_U9745  ( .A(1'b1), .ZN(_u0_ch27_csr[28] ) );
INV_X4 _u0_U9743  ( .A(1'b1), .ZN(_u0_ch27_csr[27] ) );
INV_X4 _u0_U9741  ( .A(1'b1), .ZN(_u0_ch27_csr[26] ) );
INV_X4 _u0_U9739  ( .A(1'b1), .ZN(_u0_ch27_csr[25] ) );
INV_X4 _u0_U9737  ( .A(1'b1), .ZN(_u0_ch27_csr[24] ) );
INV_X4 _u0_U9735  ( .A(1'b1), .ZN(_u0_ch27_csr[23] ) );
INV_X4 _u0_U9733  ( .A(1'b1), .ZN(_u0_ch27_csr[22] ) );
INV_X4 _u0_U9731  ( .A(1'b1), .ZN(_u0_ch27_csr[21] ) );
INV_X4 _u0_U9729  ( .A(1'b1), .ZN(_u0_ch27_csr[20] ) );
INV_X4 _u0_U9727  ( .A(1'b1), .ZN(_u0_ch27_csr[19] ) );
INV_X4 _u0_U9725  ( .A(1'b1), .ZN(_u0_ch27_csr[18] ) );
INV_X4 _u0_U9723  ( .A(1'b1), .ZN(_u0_ch27_csr[17] ) );
INV_X4 _u0_U9721  ( .A(1'b1), .ZN(_u0_ch27_csr[16] ) );
INV_X4 _u0_U9719  ( .A(1'b1), .ZN(_u0_ch27_csr[15] ) );
INV_X4 _u0_U9717  ( .A(1'b1), .ZN(_u0_ch27_csr[14] ) );
INV_X4 _u0_U9715  ( .A(1'b1), .ZN(_u0_ch27_csr[13] ) );
INV_X4 _u0_U9713  ( .A(1'b1), .ZN(_u0_ch27_csr[12] ) );
INV_X4 _u0_U9711  ( .A(1'b1), .ZN(_u0_ch27_csr[11] ) );
INV_X4 _u0_U9709  ( .A(1'b1), .ZN(_u0_ch27_csr[10] ) );
INV_X4 _u0_U9707  ( .A(1'b1), .ZN(_u0_ch27_csr[9] ) );
INV_X4 _u0_U9705  ( .A(1'b1), .ZN(_u0_ch27_csr[8] ) );
INV_X4 _u0_U9703  ( .A(1'b1), .ZN(_u0_ch27_csr[7] ) );
INV_X4 _u0_U9701  ( .A(1'b1), .ZN(_u0_ch27_csr[6] ) );
INV_X4 _u0_U9699  ( .A(1'b1), .ZN(_u0_ch27_csr[5] ) );
INV_X4 _u0_U9697  ( .A(1'b1), .ZN(_u0_ch27_csr[4] ) );
INV_X4 _u0_U9695  ( .A(1'b1), .ZN(_u0_ch27_csr[3] ) );
INV_X4 _u0_U9693  ( .A(1'b1), .ZN(_u0_ch27_csr[2] ) );
INV_X4 _u0_U9691  ( .A(1'b1), .ZN(_u0_ch27_csr[1] ) );
INV_X4 _u0_U9689  ( .A(1'b1), .ZN(_u0_ch27_csr[0] ) );
INV_X4 _u0_U9687  ( .A(1'b1), .ZN(_u0_ch27_txsz[31] ) );
INV_X4 _u0_U9685  ( .A(1'b1), .ZN(_u0_ch27_txsz[30] ) );
INV_X4 _u0_U9683  ( .A(1'b1), .ZN(_u0_ch27_txsz[29] ) );
INV_X4 _u0_U9681  ( .A(1'b1), .ZN(_u0_ch27_txsz[28] ) );
INV_X4 _u0_U9679  ( .A(1'b1), .ZN(_u0_ch27_txsz[27] ) );
INV_X4 _u0_U9677  ( .A(1'b1), .ZN(_u0_ch27_txsz[26] ) );
INV_X4 _u0_U9675  ( .A(1'b1), .ZN(_u0_ch27_txsz[25] ) );
INV_X4 _u0_U9673  ( .A(1'b1), .ZN(_u0_ch27_txsz[24] ) );
INV_X4 _u0_U9671  ( .A(1'b1), .ZN(_u0_ch27_txsz[23] ) );
INV_X4 _u0_U9669  ( .A(1'b1), .ZN(_u0_ch27_txsz[22] ) );
INV_X4 _u0_U9667  ( .A(1'b1), .ZN(_u0_ch27_txsz[21] ) );
INV_X4 _u0_U9665  ( .A(1'b1), .ZN(_u0_ch27_txsz[20] ) );
INV_X4 _u0_U9663  ( .A(1'b1), .ZN(_u0_ch27_txsz[19] ) );
INV_X4 _u0_U9661  ( .A(1'b1), .ZN(_u0_ch27_txsz[18] ) );
INV_X4 _u0_U9659  ( .A(1'b1), .ZN(_u0_ch27_txsz[17] ) );
INV_X4 _u0_U9657  ( .A(1'b1), .ZN(_u0_ch27_txsz[16] ) );
INV_X4 _u0_U9655  ( .A(1'b1), .ZN(_u0_ch27_txsz[15] ) );
INV_X4 _u0_U9653  ( .A(1'b1), .ZN(_u0_ch27_txsz[14] ) );
INV_X4 _u0_U9651  ( .A(1'b1), .ZN(_u0_ch27_txsz[13] ) );
INV_X4 _u0_U9649  ( .A(1'b1), .ZN(_u0_ch27_txsz[12] ) );
INV_X4 _u0_U9647  ( .A(1'b1), .ZN(_u0_ch27_txsz[11] ) );
INV_X4 _u0_U9645  ( .A(1'b1), .ZN(_u0_ch27_txsz[10] ) );
INV_X4 _u0_U9643  ( .A(1'b1), .ZN(_u0_ch27_txsz[9] ) );
INV_X4 _u0_U9641  ( .A(1'b1), .ZN(_u0_ch27_txsz[8] ) );
INV_X4 _u0_U9639  ( .A(1'b1), .ZN(_u0_ch27_txsz[7] ) );
INV_X4 _u0_U9637  ( .A(1'b1), .ZN(_u0_ch27_txsz[6] ) );
INV_X4 _u0_U9635  ( .A(1'b1), .ZN(_u0_ch27_txsz[5] ) );
INV_X4 _u0_U9633  ( .A(1'b1), .ZN(_u0_ch27_txsz[4] ) );
INV_X4 _u0_U9631  ( .A(1'b1), .ZN(_u0_ch27_txsz[3] ) );
INV_X4 _u0_U9629  ( .A(1'b1), .ZN(_u0_ch27_txsz[2] ) );
INV_X4 _u0_U9627  ( .A(1'b1), .ZN(_u0_ch27_txsz[1] ) );
INV_X4 _u0_U9625  ( .A(1'b1), .ZN(_u0_ch27_txsz[0] ) );
INV_X4 _u0_U9623  ( .A(1'b1), .ZN(_u0_ch27_adr0[31] ) );
INV_X4 _u0_U9621  ( .A(1'b1), .ZN(_u0_ch27_adr0[30] ) );
INV_X4 _u0_U9619  ( .A(1'b1), .ZN(_u0_ch27_adr0[29] ) );
INV_X4 _u0_U9617  ( .A(1'b1), .ZN(_u0_ch27_adr0[28] ) );
INV_X4 _u0_U9615  ( .A(1'b1), .ZN(_u0_ch27_adr0[27] ) );
INV_X4 _u0_U9613  ( .A(1'b1), .ZN(_u0_ch27_adr0[26] ) );
INV_X4 _u0_U9611  ( .A(1'b1), .ZN(_u0_ch27_adr0[25] ) );
INV_X4 _u0_U9609  ( .A(1'b1), .ZN(_u0_ch27_adr0[24] ) );
INV_X4 _u0_U9607  ( .A(1'b1), .ZN(_u0_ch27_adr0[23] ) );
INV_X4 _u0_U9605  ( .A(1'b1), .ZN(_u0_ch27_adr0[22] ) );
INV_X4 _u0_U9603  ( .A(1'b1), .ZN(_u0_ch27_adr0[21] ) );
INV_X4 _u0_U9601  ( .A(1'b1), .ZN(_u0_ch27_adr0[20] ) );
INV_X4 _u0_U9599  ( .A(1'b1), .ZN(_u0_ch27_adr0[19] ) );
INV_X4 _u0_U9597  ( .A(1'b1), .ZN(_u0_ch27_adr0[18] ) );
INV_X4 _u0_U9595  ( .A(1'b1), .ZN(_u0_ch27_adr0[17] ) );
INV_X4 _u0_U9593  ( .A(1'b1), .ZN(_u0_ch27_adr0[16] ) );
INV_X4 _u0_U9591  ( .A(1'b1), .ZN(_u0_ch27_adr0[15] ) );
INV_X4 _u0_U9589  ( .A(1'b1), .ZN(_u0_ch27_adr0[14] ) );
INV_X4 _u0_U9587  ( .A(1'b1), .ZN(_u0_ch27_adr0[13] ) );
INV_X4 _u0_U9585  ( .A(1'b1), .ZN(_u0_ch27_adr0[12] ) );
INV_X4 _u0_U9583  ( .A(1'b1), .ZN(_u0_ch27_adr0[11] ) );
INV_X4 _u0_U9581  ( .A(1'b1), .ZN(_u0_ch27_adr0[10] ) );
INV_X4 _u0_U9579  ( .A(1'b1), .ZN(_u0_ch27_adr0[9] ) );
INV_X4 _u0_U9577  ( .A(1'b1), .ZN(_u0_ch27_adr0[8] ) );
INV_X4 _u0_U9575  ( .A(1'b1), .ZN(_u0_ch27_adr0[7] ) );
INV_X4 _u0_U9573  ( .A(1'b1), .ZN(_u0_ch27_adr0[6] ) );
INV_X4 _u0_U9571  ( .A(1'b1), .ZN(_u0_ch27_adr0[5] ) );
INV_X4 _u0_U9569  ( .A(1'b1), .ZN(_u0_ch27_adr0[4] ) );
INV_X4 _u0_U9567  ( .A(1'b1), .ZN(_u0_ch27_adr0[3] ) );
INV_X4 _u0_U9565  ( .A(1'b1), .ZN(_u0_ch27_adr0[2] ) );
INV_X4 _u0_U9563  ( .A(1'b1), .ZN(_u0_ch27_adr0[1] ) );
INV_X4 _u0_U9561  ( .A(1'b1), .ZN(_u0_ch27_adr0[0] ) );
INV_X4 _u0_U9559  ( .A(1'b1), .ZN(_u0_ch27_adr1[31] ) );
INV_X4 _u0_U9557  ( .A(1'b1), .ZN(_u0_ch27_adr1[30] ) );
INV_X4 _u0_U9555  ( .A(1'b1), .ZN(_u0_ch27_adr1[29] ) );
INV_X4 _u0_U9553  ( .A(1'b1), .ZN(_u0_ch27_adr1[28] ) );
INV_X4 _u0_U9551  ( .A(1'b1), .ZN(_u0_ch27_adr1[27] ) );
INV_X4 _u0_U9549  ( .A(1'b1), .ZN(_u0_ch27_adr1[26] ) );
INV_X4 _u0_U9547  ( .A(1'b1), .ZN(_u0_ch27_adr1[25] ) );
INV_X4 _u0_U9545  ( .A(1'b1), .ZN(_u0_ch27_adr1[24] ) );
INV_X4 _u0_U9543  ( .A(1'b1), .ZN(_u0_ch27_adr1[23] ) );
INV_X4 _u0_U9541  ( .A(1'b1), .ZN(_u0_ch27_adr1[22] ) );
INV_X4 _u0_U9539  ( .A(1'b1), .ZN(_u0_ch27_adr1[21] ) );
INV_X4 _u0_U9537  ( .A(1'b1), .ZN(_u0_ch27_adr1[20] ) );
INV_X4 _u0_U9535  ( .A(1'b1), .ZN(_u0_ch27_adr1[19] ) );
INV_X4 _u0_U9533  ( .A(1'b1), .ZN(_u0_ch27_adr1[18] ) );
INV_X4 _u0_U9531  ( .A(1'b1), .ZN(_u0_ch27_adr1[17] ) );
INV_X4 _u0_U9529  ( .A(1'b1), .ZN(_u0_ch27_adr1[16] ) );
INV_X4 _u0_U9527  ( .A(1'b1), .ZN(_u0_ch27_adr1[15] ) );
INV_X4 _u0_U9525  ( .A(1'b1), .ZN(_u0_ch27_adr1[14] ) );
INV_X4 _u0_U9523  ( .A(1'b1), .ZN(_u0_ch27_adr1[13] ) );
INV_X4 _u0_U9521  ( .A(1'b1), .ZN(_u0_ch27_adr1[12] ) );
INV_X4 _u0_U9519  ( .A(1'b1), .ZN(_u0_ch27_adr1[11] ) );
INV_X4 _u0_U9517  ( .A(1'b1), .ZN(_u0_ch27_adr1[10] ) );
INV_X4 _u0_U9515  ( .A(1'b1), .ZN(_u0_ch27_adr1[9] ) );
INV_X4 _u0_U9513  ( .A(1'b1), .ZN(_u0_ch27_adr1[8] ) );
INV_X4 _u0_U9511  ( .A(1'b1), .ZN(_u0_ch27_adr1[7] ) );
INV_X4 _u0_U9509  ( .A(1'b1), .ZN(_u0_ch27_adr1[6] ) );
INV_X4 _u0_U9507  ( .A(1'b1), .ZN(_u0_ch27_adr1[5] ) );
INV_X4 _u0_U9505  ( .A(1'b1), .ZN(_u0_ch27_adr1[4] ) );
INV_X4 _u0_U9503  ( .A(1'b1), .ZN(_u0_ch27_adr1[3] ) );
INV_X4 _u0_U9501  ( .A(1'b1), .ZN(_u0_ch27_adr1[2] ) );
INV_X4 _u0_U9499  ( .A(1'b1), .ZN(_u0_ch27_adr1[1] ) );
INV_X4 _u0_U9497  ( .A(1'b1), .ZN(_u0_ch27_adr1[0] ) );
INV_X4 _u0_U9495  ( .A(1'b0), .ZN(_u0_ch27_am0[31] ) );
INV_X4 _u0_U9493  ( .A(1'b0), .ZN(_u0_ch27_am0[30] ) );
INV_X4 _u0_U9491  ( .A(1'b0), .ZN(_u0_ch27_am0[29] ) );
INV_X4 _u0_U9489  ( .A(1'b0), .ZN(_u0_ch27_am0[28] ) );
INV_X4 _u0_U9487  ( .A(1'b0), .ZN(_u0_ch27_am0[27] ) );
INV_X4 _u0_U9485  ( .A(1'b0), .ZN(_u0_ch27_am0[26] ) );
INV_X4 _u0_U9483  ( .A(1'b0), .ZN(_u0_ch27_am0[25] ) );
INV_X4 _u0_U9481  ( .A(1'b0), .ZN(_u0_ch27_am0[24] ) );
INV_X4 _u0_U9479  ( .A(1'b0), .ZN(_u0_ch27_am0[23] ) );
INV_X4 _u0_U9477  ( .A(1'b0), .ZN(_u0_ch27_am0[22] ) );
INV_X4 _u0_U9475  ( .A(1'b0), .ZN(_u0_ch27_am0[21] ) );
INV_X4 _u0_U9473  ( .A(1'b0), .ZN(_u0_ch27_am0[20] ) );
INV_X4 _u0_U9471  ( .A(1'b0), .ZN(_u0_ch27_am0[19] ) );
INV_X4 _u0_U9469  ( .A(1'b0), .ZN(_u0_ch27_am0[18] ) );
INV_X4 _u0_U9467  ( .A(1'b0), .ZN(_u0_ch27_am0[17] ) );
INV_X4 _u0_U9465  ( .A(1'b0), .ZN(_u0_ch27_am0[16] ) );
INV_X4 _u0_U9463  ( .A(1'b0), .ZN(_u0_ch27_am0[15] ) );
INV_X4 _u0_U9461  ( .A(1'b0), .ZN(_u0_ch27_am0[14] ) );
INV_X4 _u0_U9459  ( .A(1'b0), .ZN(_u0_ch27_am0[13] ) );
INV_X4 _u0_U9457  ( .A(1'b0), .ZN(_u0_ch27_am0[12] ) );
INV_X4 _u0_U9455  ( .A(1'b0), .ZN(_u0_ch27_am0[11] ) );
INV_X4 _u0_U9453  ( .A(1'b0), .ZN(_u0_ch27_am0[10] ) );
INV_X4 _u0_U9451  ( .A(1'b0), .ZN(_u0_ch27_am0[9] ) );
INV_X4 _u0_U9449  ( .A(1'b0), .ZN(_u0_ch27_am0[8] ) );
INV_X4 _u0_U9447  ( .A(1'b0), .ZN(_u0_ch27_am0[7] ) );
INV_X4 _u0_U9445  ( .A(1'b0), .ZN(_u0_ch27_am0[6] ) );
INV_X4 _u0_U9443  ( .A(1'b0), .ZN(_u0_ch27_am0[5] ) );
INV_X4 _u0_U9441  ( .A(1'b0), .ZN(_u0_ch27_am0[4] ) );
INV_X4 _u0_U9439  ( .A(1'b1), .ZN(_u0_ch27_am0[3] ) );
INV_X4 _u0_U9437  ( .A(1'b1), .ZN(_u0_ch27_am0[2] ) );
INV_X4 _u0_U9435  ( .A(1'b1), .ZN(_u0_ch27_am0[1] ) );
INV_X4 _u0_U9433  ( .A(1'b1), .ZN(_u0_ch27_am0[0] ) );
INV_X4 _u0_U9431  ( .A(1'b0), .ZN(_u0_ch27_am1[31] ) );
INV_X4 _u0_U9429  ( .A(1'b0), .ZN(_u0_ch27_am1[30] ) );
INV_X4 _u0_U9427  ( .A(1'b0), .ZN(_u0_ch27_am1[29] ) );
INV_X4 _u0_U9425  ( .A(1'b0), .ZN(_u0_ch27_am1[28] ) );
INV_X4 _u0_U9423  ( .A(1'b0), .ZN(_u0_ch27_am1[27] ) );
INV_X4 _u0_U9421  ( .A(1'b0), .ZN(_u0_ch27_am1[26] ) );
INV_X4 _u0_U9419  ( .A(1'b0), .ZN(_u0_ch27_am1[25] ) );
INV_X4 _u0_U9417  ( .A(1'b0), .ZN(_u0_ch27_am1[24] ) );
INV_X4 _u0_U9415  ( .A(1'b0), .ZN(_u0_ch27_am1[23] ) );
INV_X4 _u0_U9413  ( .A(1'b0), .ZN(_u0_ch27_am1[22] ) );
INV_X4 _u0_U9411  ( .A(1'b0), .ZN(_u0_ch27_am1[21] ) );
INV_X4 _u0_U9409  ( .A(1'b0), .ZN(_u0_ch27_am1[20] ) );
INV_X4 _u0_U9407  ( .A(1'b0), .ZN(_u0_ch27_am1[19] ) );
INV_X4 _u0_U9405  ( .A(1'b0), .ZN(_u0_ch27_am1[18] ) );
INV_X4 _u0_U9403  ( .A(1'b0), .ZN(_u0_ch27_am1[17] ) );
INV_X4 _u0_U9401  ( .A(1'b0), .ZN(_u0_ch27_am1[16] ) );
INV_X4 _u0_U9399  ( .A(1'b0), .ZN(_u0_ch27_am1[15] ) );
INV_X4 _u0_U9397  ( .A(1'b0), .ZN(_u0_ch27_am1[14] ) );
INV_X4 _u0_U9395  ( .A(1'b0), .ZN(_u0_ch27_am1[13] ) );
INV_X4 _u0_U9393  ( .A(1'b0), .ZN(_u0_ch27_am1[12] ) );
INV_X4 _u0_U9391  ( .A(1'b0), .ZN(_u0_ch27_am1[11] ) );
INV_X4 _u0_U9389  ( .A(1'b0), .ZN(_u0_ch27_am1[10] ) );
INV_X4 _u0_U9387  ( .A(1'b0), .ZN(_u0_ch27_am1[9] ) );
INV_X4 _u0_U9385  ( .A(1'b0), .ZN(_u0_ch27_am1[8] ) );
INV_X4 _u0_U9383  ( .A(1'b0), .ZN(_u0_ch27_am1[7] ) );
INV_X4 _u0_U9381  ( .A(1'b0), .ZN(_u0_ch27_am1[6] ) );
INV_X4 _u0_U9379  ( .A(1'b0), .ZN(_u0_ch27_am1[5] ) );
INV_X4 _u0_U9377  ( .A(1'b0), .ZN(_u0_ch27_am1[4] ) );
INV_X4 _u0_U9375  ( .A(1'b1), .ZN(_u0_ch27_am1[3] ) );
INV_X4 _u0_U9373  ( .A(1'b1), .ZN(_u0_ch27_am1[2] ) );
INV_X4 _u0_U9371  ( .A(1'b1), .ZN(_u0_ch27_am1[1] ) );
INV_X4 _u0_U9369  ( .A(1'b1), .ZN(_u0_ch27_am1[0] ) );
INV_X4 _u0_U9367  ( .A(1'b1), .ZN(_u0_pointer28[31] ) );
INV_X4 _u0_U9365  ( .A(1'b1), .ZN(_u0_pointer28[30] ) );
INV_X4 _u0_U9363  ( .A(1'b1), .ZN(_u0_pointer28[29] ) );
INV_X4 _u0_U9361  ( .A(1'b1), .ZN(_u0_pointer28[28] ) );
INV_X4 _u0_U9359  ( .A(1'b1), .ZN(_u0_pointer28[27] ) );
INV_X4 _u0_U9357  ( .A(1'b1), .ZN(_u0_pointer28[26] ) );
INV_X4 _u0_U9355  ( .A(1'b1), .ZN(_u0_pointer28[25] ) );
INV_X4 _u0_U9353  ( .A(1'b1), .ZN(_u0_pointer28[24] ) );
INV_X4 _u0_U9351  ( .A(1'b1), .ZN(_u0_pointer28[23] ) );
INV_X4 _u0_U9349  ( .A(1'b1), .ZN(_u0_pointer28[22] ) );
INV_X4 _u0_U9347  ( .A(1'b1), .ZN(_u0_pointer28[21] ) );
INV_X4 _u0_U9345  ( .A(1'b1), .ZN(_u0_pointer28[20] ) );
INV_X4 _u0_U9343  ( .A(1'b1), .ZN(_u0_pointer28[19] ) );
INV_X4 _u0_U9341  ( .A(1'b1), .ZN(_u0_pointer28[18] ) );
INV_X4 _u0_U9339  ( .A(1'b1), .ZN(_u0_pointer28[17] ) );
INV_X4 _u0_U9337  ( .A(1'b1), .ZN(_u0_pointer28[16] ) );
INV_X4 _u0_U9335  ( .A(1'b1), .ZN(_u0_pointer28[15] ) );
INV_X4 _u0_U9333  ( .A(1'b1), .ZN(_u0_pointer28[14] ) );
INV_X4 _u0_U9331  ( .A(1'b1), .ZN(_u0_pointer28[13] ) );
INV_X4 _u0_U9329  ( .A(1'b1), .ZN(_u0_pointer28[12] ) );
INV_X4 _u0_U9327  ( .A(1'b1), .ZN(_u0_pointer28[11] ) );
INV_X4 _u0_U9325  ( .A(1'b1), .ZN(_u0_pointer28[10] ) );
INV_X4 _u0_U9323  ( .A(1'b1), .ZN(_u0_pointer28[9] ) );
INV_X4 _u0_U9321  ( .A(1'b1), .ZN(_u0_pointer28[8] ) );
INV_X4 _u0_U9319  ( .A(1'b1), .ZN(_u0_pointer28[7] ) );
INV_X4 _u0_U9317  ( .A(1'b1), .ZN(_u0_pointer28[6] ) );
INV_X4 _u0_U9315  ( .A(1'b1), .ZN(_u0_pointer28[5] ) );
INV_X4 _u0_U9313  ( .A(1'b1), .ZN(_u0_pointer28[4] ) );
INV_X4 _u0_U9311  ( .A(1'b1), .ZN(_u0_pointer28[3] ) );
INV_X4 _u0_U9309  ( .A(1'b1), .ZN(_u0_pointer28[2] ) );
INV_X4 _u0_U9307  ( .A(1'b1), .ZN(_u0_pointer28[1] ) );
INV_X4 _u0_U9305  ( .A(1'b1), .ZN(_u0_pointer28[0] ) );
INV_X4 _u0_U9303  ( .A(1'b1), .ZN(_u0_pointer28_s[31] ) );
INV_X4 _u0_U9301  ( .A(1'b1), .ZN(_u0_pointer28_s[30] ) );
INV_X4 _u0_U9299  ( .A(1'b1), .ZN(_u0_pointer28_s[29] ) );
INV_X4 _u0_U9297  ( .A(1'b1), .ZN(_u0_pointer28_s[28] ) );
INV_X4 _u0_U9295  ( .A(1'b1), .ZN(_u0_pointer28_s[27] ) );
INV_X4 _u0_U9293  ( .A(1'b1), .ZN(_u0_pointer28_s[26] ) );
INV_X4 _u0_U9291  ( .A(1'b1), .ZN(_u0_pointer28_s[25] ) );
INV_X4 _u0_U9289  ( .A(1'b1), .ZN(_u0_pointer28_s[24] ) );
INV_X4 _u0_U9287  ( .A(1'b1), .ZN(_u0_pointer28_s[23] ) );
INV_X4 _u0_U9285  ( .A(1'b1), .ZN(_u0_pointer28_s[22] ) );
INV_X4 _u0_U9283  ( .A(1'b1), .ZN(_u0_pointer28_s[21] ) );
INV_X4 _u0_U9281  ( .A(1'b1), .ZN(_u0_pointer28_s[20] ) );
INV_X4 _u0_U9279  ( .A(1'b1), .ZN(_u0_pointer28_s[19] ) );
INV_X4 _u0_U9277  ( .A(1'b1), .ZN(_u0_pointer28_s[18] ) );
INV_X4 _u0_U9275  ( .A(1'b1), .ZN(_u0_pointer28_s[17] ) );
INV_X4 _u0_U9273  ( .A(1'b1), .ZN(_u0_pointer28_s[16] ) );
INV_X4 _u0_U9271  ( .A(1'b1), .ZN(_u0_pointer28_s[15] ) );
INV_X4 _u0_U9269  ( .A(1'b1), .ZN(_u0_pointer28_s[14] ) );
INV_X4 _u0_U9267  ( .A(1'b1), .ZN(_u0_pointer28_s[13] ) );
INV_X4 _u0_U9265  ( .A(1'b1), .ZN(_u0_pointer28_s[12] ) );
INV_X4 _u0_U9263  ( .A(1'b1), .ZN(_u0_pointer28_s[11] ) );
INV_X4 _u0_U9261  ( .A(1'b1), .ZN(_u0_pointer28_s[10] ) );
INV_X4 _u0_U9259  ( .A(1'b1), .ZN(_u0_pointer28_s[9] ) );
INV_X4 _u0_U9257  ( .A(1'b1), .ZN(_u0_pointer28_s[8] ) );
INV_X4 _u0_U9255  ( .A(1'b1), .ZN(_u0_pointer28_s[7] ) );
INV_X4 _u0_U9253  ( .A(1'b1), .ZN(_u0_pointer28_s[6] ) );
INV_X4 _u0_U9251  ( .A(1'b1), .ZN(_u0_pointer28_s[5] ) );
INV_X4 _u0_U9249  ( .A(1'b1), .ZN(_u0_pointer28_s[4] ) );
INV_X4 _u0_U9247  ( .A(1'b1), .ZN(_u0_pointer28_s[3] ) );
INV_X4 _u0_U9245  ( .A(1'b1), .ZN(_u0_pointer28_s[2] ) );
INV_X4 _u0_U9243  ( .A(1'b1), .ZN(_u0_pointer28_s[1] ) );
INV_X4 _u0_U9241  ( .A(1'b1), .ZN(_u0_pointer28_s[0] ) );
INV_X4 _u0_U9239  ( .A(1'b1), .ZN(_u0_ch28_csr[31] ) );
INV_X4 _u0_U9237  ( .A(1'b1), .ZN(_u0_ch28_csr[30] ) );
INV_X4 _u0_U9235  ( .A(1'b1), .ZN(_u0_ch28_csr[29] ) );
INV_X4 _u0_U9233  ( .A(1'b1), .ZN(_u0_ch28_csr[28] ) );
INV_X4 _u0_U9231  ( .A(1'b1), .ZN(_u0_ch28_csr[27] ) );
INV_X4 _u0_U9229  ( .A(1'b1), .ZN(_u0_ch28_csr[26] ) );
INV_X4 _u0_U9227  ( .A(1'b1), .ZN(_u0_ch28_csr[25] ) );
INV_X4 _u0_U9225  ( .A(1'b1), .ZN(_u0_ch28_csr[24] ) );
INV_X4 _u0_U9223  ( .A(1'b1), .ZN(_u0_ch28_csr[23] ) );
INV_X4 _u0_U9221  ( .A(1'b1), .ZN(_u0_ch28_csr[22] ) );
INV_X4 _u0_U9219  ( .A(1'b1), .ZN(_u0_ch28_csr[21] ) );
INV_X4 _u0_U9217  ( .A(1'b1), .ZN(_u0_ch28_csr[20] ) );
INV_X4 _u0_U9215  ( .A(1'b1), .ZN(_u0_ch28_csr[19] ) );
INV_X4 _u0_U9213  ( .A(1'b1), .ZN(_u0_ch28_csr[18] ) );
INV_X4 _u0_U9211  ( .A(1'b1), .ZN(_u0_ch28_csr[17] ) );
INV_X4 _u0_U9209  ( .A(1'b1), .ZN(_u0_ch28_csr[16] ) );
INV_X4 _u0_U9207  ( .A(1'b1), .ZN(_u0_ch28_csr[15] ) );
INV_X4 _u0_U9205  ( .A(1'b1), .ZN(_u0_ch28_csr[14] ) );
INV_X4 _u0_U9203  ( .A(1'b1), .ZN(_u0_ch28_csr[13] ) );
INV_X4 _u0_U9201  ( .A(1'b1), .ZN(_u0_ch28_csr[12] ) );
INV_X4 _u0_U9199  ( .A(1'b1), .ZN(_u0_ch28_csr[11] ) );
INV_X4 _u0_U9197  ( .A(1'b1), .ZN(_u0_ch28_csr[10] ) );
INV_X4 _u0_U9195  ( .A(1'b1), .ZN(_u0_ch28_csr[9] ) );
INV_X4 _u0_U9193  ( .A(1'b1), .ZN(_u0_ch28_csr[8] ) );
INV_X4 _u0_U9191  ( .A(1'b1), .ZN(_u0_ch28_csr[7] ) );
INV_X4 _u0_U9189  ( .A(1'b1), .ZN(_u0_ch28_csr[6] ) );
INV_X4 _u0_U9187  ( .A(1'b1), .ZN(_u0_ch28_csr[5] ) );
INV_X4 _u0_U9185  ( .A(1'b1), .ZN(_u0_ch28_csr[4] ) );
INV_X4 _u0_U9183  ( .A(1'b1), .ZN(_u0_ch28_csr[3] ) );
INV_X4 _u0_U9181  ( .A(1'b1), .ZN(_u0_ch28_csr[2] ) );
INV_X4 _u0_U9179  ( .A(1'b1), .ZN(_u0_ch28_csr[1] ) );
INV_X4 _u0_U9177  ( .A(1'b1), .ZN(_u0_ch28_csr[0] ) );
INV_X4 _u0_U9175  ( .A(1'b1), .ZN(_u0_ch28_txsz[31] ) );
INV_X4 _u0_U9173  ( .A(1'b1), .ZN(_u0_ch28_txsz[30] ) );
INV_X4 _u0_U9171  ( .A(1'b1), .ZN(_u0_ch28_txsz[29] ) );
INV_X4 _u0_U9169  ( .A(1'b1), .ZN(_u0_ch28_txsz[28] ) );
INV_X4 _u0_U9167  ( .A(1'b1), .ZN(_u0_ch28_txsz[27] ) );
INV_X4 _u0_U9165  ( .A(1'b1), .ZN(_u0_ch28_txsz[26] ) );
INV_X4 _u0_U9163  ( .A(1'b1), .ZN(_u0_ch28_txsz[25] ) );
INV_X4 _u0_U9161  ( .A(1'b1), .ZN(_u0_ch28_txsz[24] ) );
INV_X4 _u0_U9159  ( .A(1'b1), .ZN(_u0_ch28_txsz[23] ) );
INV_X4 _u0_U9157  ( .A(1'b1), .ZN(_u0_ch28_txsz[22] ) );
INV_X4 _u0_U9155  ( .A(1'b1), .ZN(_u0_ch28_txsz[21] ) );
INV_X4 _u0_U9153  ( .A(1'b1), .ZN(_u0_ch28_txsz[20] ) );
INV_X4 _u0_U9151  ( .A(1'b1), .ZN(_u0_ch28_txsz[19] ) );
INV_X4 _u0_U9149  ( .A(1'b1), .ZN(_u0_ch28_txsz[18] ) );
INV_X4 _u0_U9147  ( .A(1'b1), .ZN(_u0_ch28_txsz[17] ) );
INV_X4 _u0_U9145  ( .A(1'b1), .ZN(_u0_ch28_txsz[16] ) );
INV_X4 _u0_U9143  ( .A(1'b1), .ZN(_u0_ch28_txsz[15] ) );
INV_X4 _u0_U9141  ( .A(1'b1), .ZN(_u0_ch28_txsz[14] ) );
INV_X4 _u0_U9139  ( .A(1'b1), .ZN(_u0_ch28_txsz[13] ) );
INV_X4 _u0_U9137  ( .A(1'b1), .ZN(_u0_ch28_txsz[12] ) );
INV_X4 _u0_U9135  ( .A(1'b1), .ZN(_u0_ch28_txsz[11] ) );
INV_X4 _u0_U9133  ( .A(1'b1), .ZN(_u0_ch28_txsz[10] ) );
INV_X4 _u0_U9131  ( .A(1'b1), .ZN(_u0_ch28_txsz[9] ) );
INV_X4 _u0_U9129  ( .A(1'b1), .ZN(_u0_ch28_txsz[8] ) );
INV_X4 _u0_U9127  ( .A(1'b1), .ZN(_u0_ch28_txsz[7] ) );
INV_X4 _u0_U9125  ( .A(1'b1), .ZN(_u0_ch28_txsz[6] ) );
INV_X4 _u0_U9123  ( .A(1'b1), .ZN(_u0_ch28_txsz[5] ) );
INV_X4 _u0_U9121  ( .A(1'b1), .ZN(_u0_ch28_txsz[4] ) );
INV_X4 _u0_U9119  ( .A(1'b1), .ZN(_u0_ch28_txsz[3] ) );
INV_X4 _u0_U9117  ( .A(1'b1), .ZN(_u0_ch28_txsz[2] ) );
INV_X4 _u0_U9115  ( .A(1'b1), .ZN(_u0_ch28_txsz[1] ) );
INV_X4 _u0_U9113  ( .A(1'b1), .ZN(_u0_ch28_txsz[0] ) );
INV_X4 _u0_U9111  ( .A(1'b1), .ZN(_u0_ch28_adr0[31] ) );
INV_X4 _u0_U9109  ( .A(1'b1), .ZN(_u0_ch28_adr0[30] ) );
INV_X4 _u0_U9107  ( .A(1'b1), .ZN(_u0_ch28_adr0[29] ) );
INV_X4 _u0_U9105  ( .A(1'b1), .ZN(_u0_ch28_adr0[28] ) );
INV_X4 _u0_U9103  ( .A(1'b1), .ZN(_u0_ch28_adr0[27] ) );
INV_X4 _u0_U9101  ( .A(1'b1), .ZN(_u0_ch28_adr0[26] ) );
INV_X4 _u0_U9099  ( .A(1'b1), .ZN(_u0_ch28_adr0[25] ) );
INV_X4 _u0_U9097  ( .A(1'b1), .ZN(_u0_ch28_adr0[24] ) );
INV_X4 _u0_U9095  ( .A(1'b1), .ZN(_u0_ch28_adr0[23] ) );
INV_X4 _u0_U9093  ( .A(1'b1), .ZN(_u0_ch28_adr0[22] ) );
INV_X4 _u0_U9091  ( .A(1'b1), .ZN(_u0_ch28_adr0[21] ) );
INV_X4 _u0_U9089  ( .A(1'b1), .ZN(_u0_ch28_adr0[20] ) );
INV_X4 _u0_U9087  ( .A(1'b1), .ZN(_u0_ch28_adr0[19] ) );
INV_X4 _u0_U9085  ( .A(1'b1), .ZN(_u0_ch28_adr0[18] ) );
INV_X4 _u0_U9083  ( .A(1'b1), .ZN(_u0_ch28_adr0[17] ) );
INV_X4 _u0_U9081  ( .A(1'b1), .ZN(_u0_ch28_adr0[16] ) );
INV_X4 _u0_U9079  ( .A(1'b1), .ZN(_u0_ch28_adr0[15] ) );
INV_X4 _u0_U9077  ( .A(1'b1), .ZN(_u0_ch28_adr0[14] ) );
INV_X4 _u0_U9075  ( .A(1'b1), .ZN(_u0_ch28_adr0[13] ) );
INV_X4 _u0_U9073  ( .A(1'b1), .ZN(_u0_ch28_adr0[12] ) );
INV_X4 _u0_U9071  ( .A(1'b1), .ZN(_u0_ch28_adr0[11] ) );
INV_X4 _u0_U9069  ( .A(1'b1), .ZN(_u0_ch28_adr0[10] ) );
INV_X4 _u0_U9067  ( .A(1'b1), .ZN(_u0_ch28_adr0[9] ) );
INV_X4 _u0_U9065  ( .A(1'b1), .ZN(_u0_ch28_adr0[8] ) );
INV_X4 _u0_U9063  ( .A(1'b1), .ZN(_u0_ch28_adr0[7] ) );
INV_X4 _u0_U9061  ( .A(1'b1), .ZN(_u0_ch28_adr0[6] ) );
INV_X4 _u0_U9059  ( .A(1'b1), .ZN(_u0_ch28_adr0[5] ) );
INV_X4 _u0_U9057  ( .A(1'b1), .ZN(_u0_ch28_adr0[4] ) );
INV_X4 _u0_U9055  ( .A(1'b1), .ZN(_u0_ch28_adr0[3] ) );
INV_X4 _u0_U9053  ( .A(1'b1), .ZN(_u0_ch28_adr0[2] ) );
INV_X4 _u0_U9051  ( .A(1'b1), .ZN(_u0_ch28_adr0[1] ) );
INV_X4 _u0_U9049  ( .A(1'b1), .ZN(_u0_ch28_adr0[0] ) );
INV_X4 _u0_U9047  ( .A(1'b1), .ZN(_u0_ch28_adr1[31] ) );
INV_X4 _u0_U9045  ( .A(1'b1), .ZN(_u0_ch28_adr1[30] ) );
INV_X4 _u0_U9043  ( .A(1'b1), .ZN(_u0_ch28_adr1[29] ) );
INV_X4 _u0_U9041  ( .A(1'b1), .ZN(_u0_ch28_adr1[28] ) );
INV_X4 _u0_U9039  ( .A(1'b1), .ZN(_u0_ch28_adr1[27] ) );
INV_X4 _u0_U9037  ( .A(1'b1), .ZN(_u0_ch28_adr1[26] ) );
INV_X4 _u0_U9035  ( .A(1'b1), .ZN(_u0_ch28_adr1[25] ) );
INV_X4 _u0_U9033  ( .A(1'b1), .ZN(_u0_ch28_adr1[24] ) );
INV_X4 _u0_U9031  ( .A(1'b1), .ZN(_u0_ch28_adr1[23] ) );
INV_X4 _u0_U9029  ( .A(1'b1), .ZN(_u0_ch28_adr1[22] ) );
INV_X4 _u0_U9027  ( .A(1'b1), .ZN(_u0_ch28_adr1[21] ) );
INV_X4 _u0_U9025  ( .A(1'b1), .ZN(_u0_ch28_adr1[20] ) );
INV_X4 _u0_U9023  ( .A(1'b1), .ZN(_u0_ch28_adr1[19] ) );
INV_X4 _u0_U9021  ( .A(1'b1), .ZN(_u0_ch28_adr1[18] ) );
INV_X4 _u0_U9019  ( .A(1'b1), .ZN(_u0_ch28_adr1[17] ) );
INV_X4 _u0_U9017  ( .A(1'b1), .ZN(_u0_ch28_adr1[16] ) );
INV_X4 _u0_U9015  ( .A(1'b1), .ZN(_u0_ch28_adr1[15] ) );
INV_X4 _u0_U9013  ( .A(1'b1), .ZN(_u0_ch28_adr1[14] ) );
INV_X4 _u0_U9011  ( .A(1'b1), .ZN(_u0_ch28_adr1[13] ) );
INV_X4 _u0_U9009  ( .A(1'b1), .ZN(_u0_ch28_adr1[12] ) );
INV_X4 _u0_U9007  ( .A(1'b1), .ZN(_u0_ch28_adr1[11] ) );
INV_X4 _u0_U9005  ( .A(1'b1), .ZN(_u0_ch28_adr1[10] ) );
INV_X4 _u0_U9003  ( .A(1'b1), .ZN(_u0_ch28_adr1[9] ) );
INV_X4 _u0_U9001  ( .A(1'b1), .ZN(_u0_ch28_adr1[8] ) );
INV_X4 _u0_U8999  ( .A(1'b1), .ZN(_u0_ch28_adr1[7] ) );
INV_X4 _u0_U8997  ( .A(1'b1), .ZN(_u0_ch28_adr1[6] ) );
INV_X4 _u0_U8995  ( .A(1'b1), .ZN(_u0_ch28_adr1[5] ) );
INV_X4 _u0_U8993  ( .A(1'b1), .ZN(_u0_ch28_adr1[4] ) );
INV_X4 _u0_U8991  ( .A(1'b1), .ZN(_u0_ch28_adr1[3] ) );
INV_X4 _u0_U8989  ( .A(1'b1), .ZN(_u0_ch28_adr1[2] ) );
INV_X4 _u0_U8987  ( .A(1'b1), .ZN(_u0_ch28_adr1[1] ) );
INV_X4 _u0_U8985  ( .A(1'b1), .ZN(_u0_ch28_adr1[0] ) );
INV_X4 _u0_U8983  ( .A(1'b0), .ZN(_u0_ch28_am0[31] ) );
INV_X4 _u0_U8981  ( .A(1'b0), .ZN(_u0_ch28_am0[30] ) );
INV_X4 _u0_U8979  ( .A(1'b0), .ZN(_u0_ch28_am0[29] ) );
INV_X4 _u0_U8977  ( .A(1'b0), .ZN(_u0_ch28_am0[28] ) );
INV_X4 _u0_U8975  ( .A(1'b0), .ZN(_u0_ch28_am0[27] ) );
INV_X4 _u0_U8973  ( .A(1'b0), .ZN(_u0_ch28_am0[26] ) );
INV_X4 _u0_U8971  ( .A(1'b0), .ZN(_u0_ch28_am0[25] ) );
INV_X4 _u0_U8969  ( .A(1'b0), .ZN(_u0_ch28_am0[24] ) );
INV_X4 _u0_U8967  ( .A(1'b0), .ZN(_u0_ch28_am0[23] ) );
INV_X4 _u0_U8965  ( .A(1'b0), .ZN(_u0_ch28_am0[22] ) );
INV_X4 _u0_U8963  ( .A(1'b0), .ZN(_u0_ch28_am0[21] ) );
INV_X4 _u0_U8961  ( .A(1'b0), .ZN(_u0_ch28_am0[20] ) );
INV_X4 _u0_U8959  ( .A(1'b0), .ZN(_u0_ch28_am0[19] ) );
INV_X4 _u0_U8957  ( .A(1'b0), .ZN(_u0_ch28_am0[18] ) );
INV_X4 _u0_U8955  ( .A(1'b0), .ZN(_u0_ch28_am0[17] ) );
INV_X4 _u0_U8953  ( .A(1'b0), .ZN(_u0_ch28_am0[16] ) );
INV_X4 _u0_U8951  ( .A(1'b0), .ZN(_u0_ch28_am0[15] ) );
INV_X4 _u0_U8949  ( .A(1'b0), .ZN(_u0_ch28_am0[14] ) );
INV_X4 _u0_U8947  ( .A(1'b0), .ZN(_u0_ch28_am0[13] ) );
INV_X4 _u0_U8945  ( .A(1'b0), .ZN(_u0_ch28_am0[12] ) );
INV_X4 _u0_U8943  ( .A(1'b0), .ZN(_u0_ch28_am0[11] ) );
INV_X4 _u0_U8941  ( .A(1'b0), .ZN(_u0_ch28_am0[10] ) );
INV_X4 _u0_U8939  ( .A(1'b0), .ZN(_u0_ch28_am0[9] ) );
INV_X4 _u0_U8937  ( .A(1'b0), .ZN(_u0_ch28_am0[8] ) );
INV_X4 _u0_U8935  ( .A(1'b0), .ZN(_u0_ch28_am0[7] ) );
INV_X4 _u0_U8933  ( .A(1'b0), .ZN(_u0_ch28_am0[6] ) );
INV_X4 _u0_U8931  ( .A(1'b0), .ZN(_u0_ch28_am0[5] ) );
INV_X4 _u0_U8929  ( .A(1'b0), .ZN(_u0_ch28_am0[4] ) );
INV_X4 _u0_U8927  ( .A(1'b1), .ZN(_u0_ch28_am0[3] ) );
INV_X4 _u0_U8925  ( .A(1'b1), .ZN(_u0_ch28_am0[2] ) );
INV_X4 _u0_U8923  ( .A(1'b1), .ZN(_u0_ch28_am0[1] ) );
INV_X4 _u0_U8921  ( .A(1'b1), .ZN(_u0_ch28_am0[0] ) );
INV_X4 _u0_U8919  ( .A(1'b0), .ZN(_u0_ch28_am1[31] ) );
INV_X4 _u0_U8917  ( .A(1'b0), .ZN(_u0_ch28_am1[30] ) );
INV_X4 _u0_U8915  ( .A(1'b0), .ZN(_u0_ch28_am1[29] ) );
INV_X4 _u0_U8913  ( .A(1'b0), .ZN(_u0_ch28_am1[28] ) );
INV_X4 _u0_U8911  ( .A(1'b0), .ZN(_u0_ch28_am1[27] ) );
INV_X4 _u0_U8909  ( .A(1'b0), .ZN(_u0_ch28_am1[26] ) );
INV_X4 _u0_U8907  ( .A(1'b0), .ZN(_u0_ch28_am1[25] ) );
INV_X4 _u0_U8905  ( .A(1'b0), .ZN(_u0_ch28_am1[24] ) );
INV_X4 _u0_U8903  ( .A(1'b0), .ZN(_u0_ch28_am1[23] ) );
INV_X4 _u0_U8901  ( .A(1'b0), .ZN(_u0_ch28_am1[22] ) );
INV_X4 _u0_U8899  ( .A(1'b0), .ZN(_u0_ch28_am1[21] ) );
INV_X4 _u0_U8897  ( .A(1'b0), .ZN(_u0_ch28_am1[20] ) );
INV_X4 _u0_U8895  ( .A(1'b0), .ZN(_u0_ch28_am1[19] ) );
INV_X4 _u0_U8893  ( .A(1'b0), .ZN(_u0_ch28_am1[18] ) );
INV_X4 _u0_U8891  ( .A(1'b0), .ZN(_u0_ch28_am1[17] ) );
INV_X4 _u0_U8889  ( .A(1'b0), .ZN(_u0_ch28_am1[16] ) );
INV_X4 _u0_U8887  ( .A(1'b0), .ZN(_u0_ch28_am1[15] ) );
INV_X4 _u0_U8885  ( .A(1'b0), .ZN(_u0_ch28_am1[14] ) );
INV_X4 _u0_U8883  ( .A(1'b0), .ZN(_u0_ch28_am1[13] ) );
INV_X4 _u0_U8881  ( .A(1'b0), .ZN(_u0_ch28_am1[12] ) );
INV_X4 _u0_U8879  ( .A(1'b0), .ZN(_u0_ch28_am1[11] ) );
INV_X4 _u0_U8877  ( .A(1'b0), .ZN(_u0_ch28_am1[10] ) );
INV_X4 _u0_U8875  ( .A(1'b0), .ZN(_u0_ch28_am1[9] ) );
INV_X4 _u0_U8873  ( .A(1'b0), .ZN(_u0_ch28_am1[8] ) );
INV_X4 _u0_U8871  ( .A(1'b0), .ZN(_u0_ch28_am1[7] ) );
INV_X4 _u0_U8869  ( .A(1'b0), .ZN(_u0_ch28_am1[6] ) );
INV_X4 _u0_U8867  ( .A(1'b0), .ZN(_u0_ch28_am1[5] ) );
INV_X4 _u0_U8865  ( .A(1'b0), .ZN(_u0_ch28_am1[4] ) );
INV_X4 _u0_U8863  ( .A(1'b1), .ZN(_u0_ch28_am1[3] ) );
INV_X4 _u0_U8861  ( .A(1'b1), .ZN(_u0_ch28_am1[2] ) );
INV_X4 _u0_U8859  ( .A(1'b1), .ZN(_u0_ch28_am1[1] ) );
INV_X4 _u0_U8857  ( .A(1'b1), .ZN(_u0_ch28_am1[0] ) );
INV_X4 _u0_U8855  ( .A(1'b1), .ZN(_u0_pointer29[31] ) );
INV_X4 _u0_U8853  ( .A(1'b1), .ZN(_u0_pointer29[30] ) );
INV_X4 _u0_U8851  ( .A(1'b1), .ZN(_u0_pointer29[29] ) );
INV_X4 _u0_U8849  ( .A(1'b1), .ZN(_u0_pointer29[28] ) );
INV_X4 _u0_U8847  ( .A(1'b1), .ZN(_u0_pointer29[27] ) );
INV_X4 _u0_U8845  ( .A(1'b1), .ZN(_u0_pointer29[26] ) );
INV_X4 _u0_U8843  ( .A(1'b1), .ZN(_u0_pointer29[25] ) );
INV_X4 _u0_U8841  ( .A(1'b1), .ZN(_u0_pointer29[24] ) );
INV_X4 _u0_U8839  ( .A(1'b1), .ZN(_u0_pointer29[23] ) );
INV_X4 _u0_U8837  ( .A(1'b1), .ZN(_u0_pointer29[22] ) );
INV_X4 _u0_U8835  ( .A(1'b1), .ZN(_u0_pointer29[21] ) );
INV_X4 _u0_U8833  ( .A(1'b1), .ZN(_u0_pointer29[20] ) );
INV_X4 _u0_U8831  ( .A(1'b1), .ZN(_u0_pointer29[19] ) );
INV_X4 _u0_U8829  ( .A(1'b1), .ZN(_u0_pointer29[18] ) );
INV_X4 _u0_U8827  ( .A(1'b1), .ZN(_u0_pointer29[17] ) );
INV_X4 _u0_U8825  ( .A(1'b1), .ZN(_u0_pointer29[16] ) );
INV_X4 _u0_U8823  ( .A(1'b1), .ZN(_u0_pointer29[15] ) );
INV_X4 _u0_U8821  ( .A(1'b1), .ZN(_u0_pointer29[14] ) );
INV_X4 _u0_U8819  ( .A(1'b1), .ZN(_u0_pointer29[13] ) );
INV_X4 _u0_U8817  ( .A(1'b1), .ZN(_u0_pointer29[12] ) );
INV_X4 _u0_U8815  ( .A(1'b1), .ZN(_u0_pointer29[11] ) );
INV_X4 _u0_U8813  ( .A(1'b1), .ZN(_u0_pointer29[10] ) );
INV_X4 _u0_U8811  ( .A(1'b1), .ZN(_u0_pointer29[9] ) );
INV_X4 _u0_U8809  ( .A(1'b1), .ZN(_u0_pointer29[8] ) );
INV_X4 _u0_U8807  ( .A(1'b1), .ZN(_u0_pointer29[7] ) );
INV_X4 _u0_U8805  ( .A(1'b1), .ZN(_u0_pointer29[6] ) );
INV_X4 _u0_U8803  ( .A(1'b1), .ZN(_u0_pointer29[5] ) );
INV_X4 _u0_U8801  ( .A(1'b1), .ZN(_u0_pointer29[4] ) );
INV_X4 _u0_U8799  ( .A(1'b1), .ZN(_u0_pointer29[3] ) );
INV_X4 _u0_U8797  ( .A(1'b1), .ZN(_u0_pointer29[2] ) );
INV_X4 _u0_U8795  ( .A(1'b1), .ZN(_u0_pointer29[1] ) );
INV_X4 _u0_U8793  ( .A(1'b1), .ZN(_u0_pointer29[0] ) );
INV_X4 _u0_U8791  ( .A(1'b1), .ZN(_u0_pointer29_s[31] ) );
INV_X4 _u0_U8789  ( .A(1'b1), .ZN(_u0_pointer29_s[30] ) );
INV_X4 _u0_U8787  ( .A(1'b1), .ZN(_u0_pointer29_s[29] ) );
INV_X4 _u0_U8785  ( .A(1'b1), .ZN(_u0_pointer29_s[28] ) );
INV_X4 _u0_U8783  ( .A(1'b1), .ZN(_u0_pointer29_s[27] ) );
INV_X4 _u0_U8781  ( .A(1'b1), .ZN(_u0_pointer29_s[26] ) );
INV_X4 _u0_U8779  ( .A(1'b1), .ZN(_u0_pointer29_s[25] ) );
INV_X4 _u0_U8777  ( .A(1'b1), .ZN(_u0_pointer29_s[24] ) );
INV_X4 _u0_U8775  ( .A(1'b1), .ZN(_u0_pointer29_s[23] ) );
INV_X4 _u0_U8773  ( .A(1'b1), .ZN(_u0_pointer29_s[22] ) );
INV_X4 _u0_U8771  ( .A(1'b1), .ZN(_u0_pointer29_s[21] ) );
INV_X4 _u0_U8769  ( .A(1'b1), .ZN(_u0_pointer29_s[20] ) );
INV_X4 _u0_U8767  ( .A(1'b1), .ZN(_u0_pointer29_s[19] ) );
INV_X4 _u0_U8765  ( .A(1'b1), .ZN(_u0_pointer29_s[18] ) );
INV_X4 _u0_U8763  ( .A(1'b1), .ZN(_u0_pointer29_s[17] ) );
INV_X4 _u0_U8761  ( .A(1'b1), .ZN(_u0_pointer29_s[16] ) );
INV_X4 _u0_U8759  ( .A(1'b1), .ZN(_u0_pointer29_s[15] ) );
INV_X4 _u0_U8757  ( .A(1'b1), .ZN(_u0_pointer29_s[14] ) );
INV_X4 _u0_U8755  ( .A(1'b1), .ZN(_u0_pointer29_s[13] ) );
INV_X4 _u0_U8753  ( .A(1'b1), .ZN(_u0_pointer29_s[12] ) );
INV_X4 _u0_U8751  ( .A(1'b1), .ZN(_u0_pointer29_s[11] ) );
INV_X4 _u0_U8749  ( .A(1'b1), .ZN(_u0_pointer29_s[10] ) );
INV_X4 _u0_U8747  ( .A(1'b1), .ZN(_u0_pointer29_s[9] ) );
INV_X4 _u0_U8745  ( .A(1'b1), .ZN(_u0_pointer29_s[8] ) );
INV_X4 _u0_U8743  ( .A(1'b1), .ZN(_u0_pointer29_s[7] ) );
INV_X4 _u0_U8741  ( .A(1'b1), .ZN(_u0_pointer29_s[6] ) );
INV_X4 _u0_U8739  ( .A(1'b1), .ZN(_u0_pointer29_s[5] ) );
INV_X4 _u0_U8737  ( .A(1'b1), .ZN(_u0_pointer29_s[4] ) );
INV_X4 _u0_U8735  ( .A(1'b1), .ZN(_u0_pointer29_s[3] ) );
INV_X4 _u0_U8733  ( .A(1'b1), .ZN(_u0_pointer29_s[2] ) );
INV_X4 _u0_U8731  ( .A(1'b1), .ZN(_u0_pointer29_s[1] ) );
INV_X4 _u0_U8729  ( .A(1'b1), .ZN(_u0_pointer29_s[0] ) );
INV_X4 _u0_U8727  ( .A(1'b1), .ZN(_u0_ch29_csr[31] ) );
INV_X4 _u0_U8725  ( .A(1'b1), .ZN(_u0_ch29_csr[30] ) );
INV_X4 _u0_U8723  ( .A(1'b1), .ZN(_u0_ch29_csr[29] ) );
INV_X4 _u0_U8721  ( .A(1'b1), .ZN(_u0_ch29_csr[28] ) );
INV_X4 _u0_U8719  ( .A(1'b1), .ZN(_u0_ch29_csr[27] ) );
INV_X4 _u0_U8717  ( .A(1'b1), .ZN(_u0_ch29_csr[26] ) );
INV_X4 _u0_U8715  ( .A(1'b1), .ZN(_u0_ch29_csr[25] ) );
INV_X4 _u0_U8713  ( .A(1'b1), .ZN(_u0_ch29_csr[24] ) );
INV_X4 _u0_U8711  ( .A(1'b1), .ZN(_u0_ch29_csr[23] ) );
INV_X4 _u0_U8709  ( .A(1'b1), .ZN(_u0_ch29_csr[22] ) );
INV_X4 _u0_U8707  ( .A(1'b1), .ZN(_u0_ch29_csr[21] ) );
INV_X4 _u0_U8705  ( .A(1'b1), .ZN(_u0_ch29_csr[20] ) );
INV_X4 _u0_U8703  ( .A(1'b1), .ZN(_u0_ch29_csr[19] ) );
INV_X4 _u0_U8701  ( .A(1'b1), .ZN(_u0_ch29_csr[18] ) );
INV_X4 _u0_U8699  ( .A(1'b1), .ZN(_u0_ch29_csr[17] ) );
INV_X4 _u0_U8697  ( .A(1'b1), .ZN(_u0_ch29_csr[16] ) );
INV_X4 _u0_U8695  ( .A(1'b1), .ZN(_u0_ch29_csr[15] ) );
INV_X4 _u0_U8693  ( .A(1'b1), .ZN(_u0_ch29_csr[14] ) );
INV_X4 _u0_U8691  ( .A(1'b1), .ZN(_u0_ch29_csr[13] ) );
INV_X4 _u0_U8689  ( .A(1'b1), .ZN(_u0_ch29_csr[12] ) );
INV_X4 _u0_U8687  ( .A(1'b1), .ZN(_u0_ch29_csr[11] ) );
INV_X4 _u0_U8685  ( .A(1'b1), .ZN(_u0_ch29_csr[10] ) );
INV_X4 _u0_U8683  ( .A(1'b1), .ZN(_u0_ch29_csr[9] ) );
INV_X4 _u0_U8681  ( .A(1'b1), .ZN(_u0_ch29_csr[8] ) );
INV_X4 _u0_U8679  ( .A(1'b1), .ZN(_u0_ch29_csr[7] ) );
INV_X4 _u0_U8677  ( .A(1'b1), .ZN(_u0_ch29_csr[6] ) );
INV_X4 _u0_U8675  ( .A(1'b1), .ZN(_u0_ch29_csr[5] ) );
INV_X4 _u0_U8673  ( .A(1'b1), .ZN(_u0_ch29_csr[4] ) );
INV_X4 _u0_U8671  ( .A(1'b1), .ZN(_u0_ch29_csr[3] ) );
INV_X4 _u0_U8669  ( .A(1'b1), .ZN(_u0_ch29_csr[2] ) );
INV_X4 _u0_U8667  ( .A(1'b1), .ZN(_u0_ch29_csr[1] ) );
INV_X4 _u0_U8665  ( .A(1'b1), .ZN(_u0_ch29_csr[0] ) );
INV_X4 _u0_U8663  ( .A(1'b1), .ZN(_u0_ch29_txsz[31] ) );
INV_X4 _u0_U8661  ( .A(1'b1), .ZN(_u0_ch29_txsz[30] ) );
INV_X4 _u0_U8659  ( .A(1'b1), .ZN(_u0_ch29_txsz[29] ) );
INV_X4 _u0_U8657  ( .A(1'b1), .ZN(_u0_ch29_txsz[28] ) );
INV_X4 _u0_U8655  ( .A(1'b1), .ZN(_u0_ch29_txsz[27] ) );
INV_X4 _u0_U8653  ( .A(1'b1), .ZN(_u0_ch29_txsz[26] ) );
INV_X4 _u0_U8651  ( .A(1'b1), .ZN(_u0_ch29_txsz[25] ) );
INV_X4 _u0_U8649  ( .A(1'b1), .ZN(_u0_ch29_txsz[24] ) );
INV_X4 _u0_U8647  ( .A(1'b1), .ZN(_u0_ch29_txsz[23] ) );
INV_X4 _u0_U8645  ( .A(1'b1), .ZN(_u0_ch29_txsz[22] ) );
INV_X4 _u0_U8643  ( .A(1'b1), .ZN(_u0_ch29_txsz[21] ) );
INV_X4 _u0_U8641  ( .A(1'b1), .ZN(_u0_ch29_txsz[20] ) );
INV_X4 _u0_U8639  ( .A(1'b1), .ZN(_u0_ch29_txsz[19] ) );
INV_X4 _u0_U8637  ( .A(1'b1), .ZN(_u0_ch29_txsz[18] ) );
INV_X4 _u0_U8635  ( .A(1'b1), .ZN(_u0_ch29_txsz[17] ) );
INV_X4 _u0_U8633  ( .A(1'b1), .ZN(_u0_ch29_txsz[16] ) );
INV_X4 _u0_U8631  ( .A(1'b1), .ZN(_u0_ch29_txsz[15] ) );
INV_X4 _u0_U8629  ( .A(1'b1), .ZN(_u0_ch29_txsz[14] ) );
INV_X4 _u0_U8627  ( .A(1'b1), .ZN(_u0_ch29_txsz[13] ) );
INV_X4 _u0_U8625  ( .A(1'b1), .ZN(_u0_ch29_txsz[12] ) );
INV_X4 _u0_U8623  ( .A(1'b1), .ZN(_u0_ch29_txsz[11] ) );
INV_X4 _u0_U8621  ( .A(1'b1), .ZN(_u0_ch29_txsz[10] ) );
INV_X4 _u0_U8619  ( .A(1'b1), .ZN(_u0_ch29_txsz[9] ) );
INV_X4 _u0_U8617  ( .A(1'b1), .ZN(_u0_ch29_txsz[8] ) );
INV_X4 _u0_U8615  ( .A(1'b1), .ZN(_u0_ch29_txsz[7] ) );
INV_X4 _u0_U8613  ( .A(1'b1), .ZN(_u0_ch29_txsz[6] ) );
INV_X4 _u0_U8611  ( .A(1'b1), .ZN(_u0_ch29_txsz[5] ) );
INV_X4 _u0_U8609  ( .A(1'b1), .ZN(_u0_ch29_txsz[4] ) );
INV_X4 _u0_U8607  ( .A(1'b1), .ZN(_u0_ch29_txsz[3] ) );
INV_X4 _u0_U8605  ( .A(1'b1), .ZN(_u0_ch29_txsz[2] ) );
INV_X4 _u0_U8603  ( .A(1'b1), .ZN(_u0_ch29_txsz[1] ) );
INV_X4 _u0_U8601  ( .A(1'b1), .ZN(_u0_ch29_txsz[0] ) );
INV_X4 _u0_U8599  ( .A(1'b1), .ZN(_u0_ch29_adr0[31] ) );
INV_X4 _u0_U8597  ( .A(1'b1), .ZN(_u0_ch29_adr0[30] ) );
INV_X4 _u0_U8595  ( .A(1'b1), .ZN(_u0_ch29_adr0[29] ) );
INV_X4 _u0_U8593  ( .A(1'b1), .ZN(_u0_ch29_adr0[28] ) );
INV_X4 _u0_U8591  ( .A(1'b1), .ZN(_u0_ch29_adr0[27] ) );
INV_X4 _u0_U8589  ( .A(1'b1), .ZN(_u0_ch29_adr0[26] ) );
INV_X4 _u0_U8587  ( .A(1'b1), .ZN(_u0_ch29_adr0[25] ) );
INV_X4 _u0_U8585  ( .A(1'b1), .ZN(_u0_ch29_adr0[24] ) );
INV_X4 _u0_U8583  ( .A(1'b1), .ZN(_u0_ch29_adr0[23] ) );
INV_X4 _u0_U8581  ( .A(1'b1), .ZN(_u0_ch29_adr0[22] ) );
INV_X4 _u0_U8579  ( .A(1'b1), .ZN(_u0_ch29_adr0[21] ) );
INV_X4 _u0_U8577  ( .A(1'b1), .ZN(_u0_ch29_adr0[20] ) );
INV_X4 _u0_U8575  ( .A(1'b1), .ZN(_u0_ch29_adr0[19] ) );
INV_X4 _u0_U8573  ( .A(1'b1), .ZN(_u0_ch29_adr0[18] ) );
INV_X4 _u0_U8571  ( .A(1'b1), .ZN(_u0_ch29_adr0[17] ) );
INV_X4 _u0_U8569  ( .A(1'b1), .ZN(_u0_ch29_adr0[16] ) );
INV_X4 _u0_U8567  ( .A(1'b1), .ZN(_u0_ch29_adr0[15] ) );
INV_X4 _u0_U8565  ( .A(1'b1), .ZN(_u0_ch29_adr0[14] ) );
INV_X4 _u0_U8563  ( .A(1'b1), .ZN(_u0_ch29_adr0[13] ) );
INV_X4 _u0_U8561  ( .A(1'b1), .ZN(_u0_ch29_adr0[12] ) );
INV_X4 _u0_U8559  ( .A(1'b1), .ZN(_u0_ch29_adr0[11] ) );
INV_X4 _u0_U8557  ( .A(1'b1), .ZN(_u0_ch29_adr0[10] ) );
INV_X4 _u0_U8555  ( .A(1'b1), .ZN(_u0_ch29_adr0[9] ) );
INV_X4 _u0_U8553  ( .A(1'b1), .ZN(_u0_ch29_adr0[8] ) );
INV_X4 _u0_U8551  ( .A(1'b1), .ZN(_u0_ch29_adr0[7] ) );
INV_X4 _u0_U8549  ( .A(1'b1), .ZN(_u0_ch29_adr0[6] ) );
INV_X4 _u0_U8547  ( .A(1'b1), .ZN(_u0_ch29_adr0[5] ) );
INV_X4 _u0_U8545  ( .A(1'b1), .ZN(_u0_ch29_adr0[4] ) );
INV_X4 _u0_U8543  ( .A(1'b1), .ZN(_u0_ch29_adr0[3] ) );
INV_X4 _u0_U8541  ( .A(1'b1), .ZN(_u0_ch29_adr0[2] ) );
INV_X4 _u0_U8539  ( .A(1'b1), .ZN(_u0_ch29_adr0[1] ) );
INV_X4 _u0_U8537  ( .A(1'b1), .ZN(_u0_ch29_adr0[0] ) );
INV_X4 _u0_U8535  ( .A(1'b1), .ZN(_u0_ch29_adr1[31] ) );
INV_X4 _u0_U8533  ( .A(1'b1), .ZN(_u0_ch29_adr1[30] ) );
INV_X4 _u0_U8531  ( .A(1'b1), .ZN(_u0_ch29_adr1[29] ) );
INV_X4 _u0_U8529  ( .A(1'b1), .ZN(_u0_ch29_adr1[28] ) );
INV_X4 _u0_U8527  ( .A(1'b1), .ZN(_u0_ch29_adr1[27] ) );
INV_X4 _u0_U8525  ( .A(1'b1), .ZN(_u0_ch29_adr1[26] ) );
INV_X4 _u0_U8523  ( .A(1'b1), .ZN(_u0_ch29_adr1[25] ) );
INV_X4 _u0_U8521  ( .A(1'b1), .ZN(_u0_ch29_adr1[24] ) );
INV_X4 _u0_U8519  ( .A(1'b1), .ZN(_u0_ch29_adr1[23] ) );
INV_X4 _u0_U8517  ( .A(1'b1), .ZN(_u0_ch29_adr1[22] ) );
INV_X4 _u0_U8515  ( .A(1'b1), .ZN(_u0_ch29_adr1[21] ) );
INV_X4 _u0_U8513  ( .A(1'b1), .ZN(_u0_ch29_adr1[20] ) );
INV_X4 _u0_U8511  ( .A(1'b1), .ZN(_u0_ch29_adr1[19] ) );
INV_X4 _u0_U8509  ( .A(1'b1), .ZN(_u0_ch29_adr1[18] ) );
INV_X4 _u0_U8507  ( .A(1'b1), .ZN(_u0_ch29_adr1[17] ) );
INV_X4 _u0_U8505  ( .A(1'b1), .ZN(_u0_ch29_adr1[16] ) );
INV_X4 _u0_U8503  ( .A(1'b1), .ZN(_u0_ch29_adr1[15] ) );
INV_X4 _u0_U8501  ( .A(1'b1), .ZN(_u0_ch29_adr1[14] ) );
INV_X4 _u0_U8499  ( .A(1'b1), .ZN(_u0_ch29_adr1[13] ) );
INV_X4 _u0_U8497  ( .A(1'b1), .ZN(_u0_ch29_adr1[12] ) );
INV_X4 _u0_U8495  ( .A(1'b1), .ZN(_u0_ch29_adr1[11] ) );
INV_X4 _u0_U8493  ( .A(1'b1), .ZN(_u0_ch29_adr1[10] ) );
INV_X4 _u0_U8491  ( .A(1'b1), .ZN(_u0_ch29_adr1[9] ) );
INV_X4 _u0_U8489  ( .A(1'b1), .ZN(_u0_ch29_adr1[8] ) );
INV_X4 _u0_U8487  ( .A(1'b1), .ZN(_u0_ch29_adr1[7] ) );
INV_X4 _u0_U8485  ( .A(1'b1), .ZN(_u0_ch29_adr1[6] ) );
INV_X4 _u0_U8483  ( .A(1'b1), .ZN(_u0_ch29_adr1[5] ) );
INV_X4 _u0_U8481  ( .A(1'b1), .ZN(_u0_ch29_adr1[4] ) );
INV_X4 _u0_U8479  ( .A(1'b1), .ZN(_u0_ch29_adr1[3] ) );
INV_X4 _u0_U8477  ( .A(1'b1), .ZN(_u0_ch29_adr1[2] ) );
INV_X4 _u0_U8475  ( .A(1'b1), .ZN(_u0_ch29_adr1[1] ) );
INV_X4 _u0_U8473  ( .A(1'b1), .ZN(_u0_ch29_adr1[0] ) );
INV_X4 _u0_U8471  ( .A(1'b0), .ZN(_u0_ch29_am0[31] ) );
INV_X4 _u0_U8469  ( .A(1'b0), .ZN(_u0_ch29_am0[30] ) );
INV_X4 _u0_U8467  ( .A(1'b0), .ZN(_u0_ch29_am0[29] ) );
INV_X4 _u0_U8465  ( .A(1'b0), .ZN(_u0_ch29_am0[28] ) );
INV_X4 _u0_U8463  ( .A(1'b0), .ZN(_u0_ch29_am0[27] ) );
INV_X4 _u0_U8461  ( .A(1'b0), .ZN(_u0_ch29_am0[26] ) );
INV_X4 _u0_U8459  ( .A(1'b0), .ZN(_u0_ch29_am0[25] ) );
INV_X4 _u0_U8457  ( .A(1'b0), .ZN(_u0_ch29_am0[24] ) );
INV_X4 _u0_U8455  ( .A(1'b0), .ZN(_u0_ch29_am0[23] ) );
INV_X4 _u0_U8453  ( .A(1'b0), .ZN(_u0_ch29_am0[22] ) );
INV_X4 _u0_U8451  ( .A(1'b0), .ZN(_u0_ch29_am0[21] ) );
INV_X4 _u0_U8449  ( .A(1'b0), .ZN(_u0_ch29_am0[20] ) );
INV_X4 _u0_U8447  ( .A(1'b0), .ZN(_u0_ch29_am0[19] ) );
INV_X4 _u0_U8445  ( .A(1'b0), .ZN(_u0_ch29_am0[18] ) );
INV_X4 _u0_U8443  ( .A(1'b0), .ZN(_u0_ch29_am0[17] ) );
INV_X4 _u0_U8441  ( .A(1'b0), .ZN(_u0_ch29_am0[16] ) );
INV_X4 _u0_U8439  ( .A(1'b0), .ZN(_u0_ch29_am0[15] ) );
INV_X4 _u0_U8437  ( .A(1'b0), .ZN(_u0_ch29_am0[14] ) );
INV_X4 _u0_U8435  ( .A(1'b0), .ZN(_u0_ch29_am0[13] ) );
INV_X4 _u0_U8433  ( .A(1'b0), .ZN(_u0_ch29_am0[12] ) );
INV_X4 _u0_U8431  ( .A(1'b0), .ZN(_u0_ch29_am0[11] ) );
INV_X4 _u0_U8429  ( .A(1'b0), .ZN(_u0_ch29_am0[10] ) );
INV_X4 _u0_U8427  ( .A(1'b0), .ZN(_u0_ch29_am0[9] ) );
INV_X4 _u0_U8425  ( .A(1'b0), .ZN(_u0_ch29_am0[8] ) );
INV_X4 _u0_U8423  ( .A(1'b0), .ZN(_u0_ch29_am0[7] ) );
INV_X4 _u0_U8421  ( .A(1'b0), .ZN(_u0_ch29_am0[6] ) );
INV_X4 _u0_U8419  ( .A(1'b0), .ZN(_u0_ch29_am0[5] ) );
INV_X4 _u0_U8417  ( .A(1'b0), .ZN(_u0_ch29_am0[4] ) );
INV_X4 _u0_U8415  ( .A(1'b1), .ZN(_u0_ch29_am0[3] ) );
INV_X4 _u0_U8413  ( .A(1'b1), .ZN(_u0_ch29_am0[2] ) );
INV_X4 _u0_U8411  ( .A(1'b1), .ZN(_u0_ch29_am0[1] ) );
INV_X4 _u0_U8409  ( .A(1'b1), .ZN(_u0_ch29_am0[0] ) );
INV_X4 _u0_U8407  ( .A(1'b0), .ZN(_u0_ch29_am1[31] ) );
INV_X4 _u0_U8405  ( .A(1'b0), .ZN(_u0_ch29_am1[30] ) );
INV_X4 _u0_U8403  ( .A(1'b0), .ZN(_u0_ch29_am1[29] ) );
INV_X4 _u0_U8401  ( .A(1'b0), .ZN(_u0_ch29_am1[28] ) );
INV_X4 _u0_U8399  ( .A(1'b0), .ZN(_u0_ch29_am1[27] ) );
INV_X4 _u0_U8397  ( .A(1'b0), .ZN(_u0_ch29_am1[26] ) );
INV_X4 _u0_U8395  ( .A(1'b0), .ZN(_u0_ch29_am1[25] ) );
INV_X4 _u0_U8393  ( .A(1'b0), .ZN(_u0_ch29_am1[24] ) );
INV_X4 _u0_U8391  ( .A(1'b0), .ZN(_u0_ch29_am1[23] ) );
INV_X4 _u0_U8389  ( .A(1'b0), .ZN(_u0_ch29_am1[22] ) );
INV_X4 _u0_U8387  ( .A(1'b0), .ZN(_u0_ch29_am1[21] ) );
INV_X4 _u0_U8385  ( .A(1'b0), .ZN(_u0_ch29_am1[20] ) );
INV_X4 _u0_U8383  ( .A(1'b0), .ZN(_u0_ch29_am1[19] ) );
INV_X4 _u0_U8381  ( .A(1'b0), .ZN(_u0_ch29_am1[18] ) );
INV_X4 _u0_U8379  ( .A(1'b0), .ZN(_u0_ch29_am1[17] ) );
INV_X4 _u0_U8377  ( .A(1'b0), .ZN(_u0_ch29_am1[16] ) );
INV_X4 _u0_U8375  ( .A(1'b0), .ZN(_u0_ch29_am1[15] ) );
INV_X4 _u0_U8373  ( .A(1'b0), .ZN(_u0_ch29_am1[14] ) );
INV_X4 _u0_U8371  ( .A(1'b0), .ZN(_u0_ch29_am1[13] ) );
INV_X4 _u0_U8369  ( .A(1'b0), .ZN(_u0_ch29_am1[12] ) );
INV_X4 _u0_U8367  ( .A(1'b0), .ZN(_u0_ch29_am1[11] ) );
INV_X4 _u0_U8365  ( .A(1'b0), .ZN(_u0_ch29_am1[10] ) );
INV_X4 _u0_U8363  ( .A(1'b0), .ZN(_u0_ch29_am1[9] ) );
INV_X4 _u0_U8361  ( .A(1'b0), .ZN(_u0_ch29_am1[8] ) );
INV_X4 _u0_U8359  ( .A(1'b0), .ZN(_u0_ch29_am1[7] ) );
INV_X4 _u0_U8357  ( .A(1'b0), .ZN(_u0_ch29_am1[6] ) );
INV_X4 _u0_U8355  ( .A(1'b0), .ZN(_u0_ch29_am1[5] ) );
INV_X4 _u0_U8353  ( .A(1'b0), .ZN(_u0_ch29_am1[4] ) );
INV_X4 _u0_U8351  ( .A(1'b1), .ZN(_u0_ch29_am1[3] ) );
INV_X4 _u0_U8349  ( .A(1'b1), .ZN(_u0_ch29_am1[2] ) );
INV_X4 _u0_U8347  ( .A(1'b1), .ZN(_u0_ch29_am1[1] ) );
INV_X4 _u0_U8345  ( .A(1'b1), .ZN(_u0_ch29_am1[0] ) );
INV_X4 _u0_U8343  ( .A(1'b1), .ZN(_u0_pointer30[31] ) );
INV_X4 _u0_U8341  ( .A(1'b1), .ZN(_u0_pointer30[30] ) );
INV_X4 _u0_U8339  ( .A(1'b1), .ZN(_u0_pointer30[29] ) );
INV_X4 _u0_U8337  ( .A(1'b1), .ZN(_u0_pointer30[28] ) );
INV_X4 _u0_U8335  ( .A(1'b1), .ZN(_u0_pointer30[27] ) );
INV_X4 _u0_U8333  ( .A(1'b1), .ZN(_u0_pointer30[26] ) );
INV_X4 _u0_U8331  ( .A(1'b1), .ZN(_u0_pointer30[25] ) );
INV_X4 _u0_U8329  ( .A(1'b1), .ZN(_u0_pointer30[24] ) );
INV_X4 _u0_U8327  ( .A(1'b1), .ZN(_u0_pointer30[23] ) );
INV_X4 _u0_U8325  ( .A(1'b1), .ZN(_u0_pointer30[22] ) );
INV_X4 _u0_U8323  ( .A(1'b1), .ZN(_u0_pointer30[21] ) );
INV_X4 _u0_U8321  ( .A(1'b1), .ZN(_u0_pointer30[20] ) );
INV_X4 _u0_U8319  ( .A(1'b1), .ZN(_u0_pointer30[19] ) );
INV_X4 _u0_U8317  ( .A(1'b1), .ZN(_u0_pointer30[18] ) );
INV_X4 _u0_U8315  ( .A(1'b1), .ZN(_u0_pointer30[17] ) );
INV_X4 _u0_U8313  ( .A(1'b1), .ZN(_u0_pointer30[16] ) );
INV_X4 _u0_U8311  ( .A(1'b1), .ZN(_u0_pointer30[15] ) );
INV_X4 _u0_U8309  ( .A(1'b1), .ZN(_u0_pointer30[14] ) );
INV_X4 _u0_U8307  ( .A(1'b1), .ZN(_u0_pointer30[13] ) );
INV_X4 _u0_U8305  ( .A(1'b1), .ZN(_u0_pointer30[12] ) );
INV_X4 _u0_U8303  ( .A(1'b1), .ZN(_u0_pointer30[11] ) );
INV_X4 _u0_U8301  ( .A(1'b1), .ZN(_u0_pointer30[10] ) );
INV_X4 _u0_U8299  ( .A(1'b1), .ZN(_u0_pointer30[9] ) );
INV_X4 _u0_U8297  ( .A(1'b1), .ZN(_u0_pointer30[8] ) );
INV_X4 _u0_U8295  ( .A(1'b1), .ZN(_u0_pointer30[7] ) );
INV_X4 _u0_U8293  ( .A(1'b1), .ZN(_u0_pointer30[6] ) );
INV_X4 _u0_U8291  ( .A(1'b1), .ZN(_u0_pointer30[5] ) );
INV_X4 _u0_U8289  ( .A(1'b1), .ZN(_u0_pointer30[4] ) );
INV_X4 _u0_U8287  ( .A(1'b1), .ZN(_u0_pointer30[3] ) );
INV_X4 _u0_U8285  ( .A(1'b1), .ZN(_u0_pointer30[2] ) );
INV_X4 _u0_U8283  ( .A(1'b1), .ZN(_u0_pointer30[1] ) );
INV_X4 _u0_U8281  ( .A(1'b1), .ZN(_u0_pointer30[0] ) );
INV_X4 _u0_U8279  ( .A(1'b1), .ZN(_u0_pointer30_s[31] ) );
INV_X4 _u0_U8277  ( .A(1'b1), .ZN(_u0_pointer30_s[30] ) );
INV_X4 _u0_U8275  ( .A(1'b1), .ZN(_u0_pointer30_s[29] ) );
INV_X4 _u0_U8273  ( .A(1'b1), .ZN(_u0_pointer30_s[28] ) );
INV_X4 _u0_U8271  ( .A(1'b1), .ZN(_u0_pointer30_s[27] ) );
INV_X4 _u0_U8269  ( .A(1'b1), .ZN(_u0_pointer30_s[26] ) );
INV_X4 _u0_U8267  ( .A(1'b1), .ZN(_u0_pointer30_s[25] ) );
INV_X4 _u0_U8265  ( .A(1'b1), .ZN(_u0_pointer30_s[24] ) );
INV_X4 _u0_U8263  ( .A(1'b1), .ZN(_u0_pointer30_s[23] ) );
INV_X4 _u0_U8261  ( .A(1'b1), .ZN(_u0_pointer30_s[22] ) );
INV_X4 _u0_U8259  ( .A(1'b1), .ZN(_u0_pointer30_s[21] ) );
INV_X4 _u0_U8257  ( .A(1'b1), .ZN(_u0_pointer30_s[20] ) );
INV_X4 _u0_U8255  ( .A(1'b1), .ZN(_u0_pointer30_s[19] ) );
INV_X4 _u0_U8253  ( .A(1'b1), .ZN(_u0_pointer30_s[18] ) );
INV_X4 _u0_U8251  ( .A(1'b1), .ZN(_u0_pointer30_s[17] ) );
INV_X4 _u0_U8249  ( .A(1'b1), .ZN(_u0_pointer30_s[16] ) );
INV_X4 _u0_U8247  ( .A(1'b1), .ZN(_u0_pointer30_s[15] ) );
INV_X4 _u0_U8245  ( .A(1'b1), .ZN(_u0_pointer30_s[14] ) );
INV_X4 _u0_U8243  ( .A(1'b1), .ZN(_u0_pointer30_s[13] ) );
INV_X4 _u0_U8241  ( .A(1'b1), .ZN(_u0_pointer30_s[12] ) );
INV_X4 _u0_U8239  ( .A(1'b1), .ZN(_u0_pointer30_s[11] ) );
INV_X4 _u0_U8237  ( .A(1'b1), .ZN(_u0_pointer30_s[10] ) );
INV_X4 _u0_U8235  ( .A(1'b1), .ZN(_u0_pointer30_s[9] ) );
INV_X4 _u0_U8233  ( .A(1'b1), .ZN(_u0_pointer30_s[8] ) );
INV_X4 _u0_U8231  ( .A(1'b1), .ZN(_u0_pointer30_s[7] ) );
INV_X4 _u0_U8229  ( .A(1'b1), .ZN(_u0_pointer30_s[6] ) );
INV_X4 _u0_U8227  ( .A(1'b1), .ZN(_u0_pointer30_s[5] ) );
INV_X4 _u0_U8225  ( .A(1'b1), .ZN(_u0_pointer30_s[4] ) );
INV_X4 _u0_U8223  ( .A(1'b1), .ZN(_u0_pointer30_s[3] ) );
INV_X4 _u0_U8221  ( .A(1'b1), .ZN(_u0_pointer30_s[2] ) );
INV_X4 _u0_U8219  ( .A(1'b1), .ZN(_u0_pointer30_s[1] ) );
INV_X4 _u0_U8217  ( .A(1'b1), .ZN(_u0_pointer30_s[0] ) );
INV_X4 _u0_U8215  ( .A(1'b1), .ZN(_u0_ch30_csr[31] ) );
INV_X4 _u0_U8213  ( .A(1'b1), .ZN(_u0_ch30_csr[30] ) );
INV_X4 _u0_U8211  ( .A(1'b1), .ZN(_u0_ch30_csr[29] ) );
INV_X4 _u0_U8209  ( .A(1'b1), .ZN(_u0_ch30_csr[28] ) );
INV_X4 _u0_U8207  ( .A(1'b1), .ZN(_u0_ch30_csr[27] ) );
INV_X4 _u0_U8205  ( .A(1'b1), .ZN(_u0_ch30_csr[26] ) );
INV_X4 _u0_U8203  ( .A(1'b1), .ZN(_u0_ch30_csr[25] ) );
INV_X4 _u0_U8201  ( .A(1'b1), .ZN(_u0_ch30_csr[24] ) );
INV_X4 _u0_U8199  ( .A(1'b1), .ZN(_u0_ch30_csr[23] ) );
INV_X4 _u0_U8197  ( .A(1'b1), .ZN(_u0_ch30_csr[22] ) );
INV_X4 _u0_U8195  ( .A(1'b1), .ZN(_u0_ch30_csr[21] ) );
INV_X4 _u0_U8193  ( .A(1'b1), .ZN(_u0_ch30_csr[20] ) );
INV_X4 _u0_U8191  ( .A(1'b1), .ZN(_u0_ch30_csr[19] ) );
INV_X4 _u0_U8189  ( .A(1'b1), .ZN(_u0_ch30_csr[18] ) );
INV_X4 _u0_U8187  ( .A(1'b1), .ZN(_u0_ch30_csr[17] ) );
INV_X4 _u0_U8185  ( .A(1'b1), .ZN(_u0_ch30_csr[16] ) );
INV_X4 _u0_U8183  ( .A(1'b1), .ZN(_u0_ch30_csr[15] ) );
INV_X4 _u0_U8181  ( .A(1'b1), .ZN(_u0_ch30_csr[14] ) );
INV_X4 _u0_U8179  ( .A(1'b1), .ZN(_u0_ch30_csr[13] ) );
INV_X4 _u0_U8177  ( .A(1'b1), .ZN(_u0_ch30_csr[12] ) );
INV_X4 _u0_U8175  ( .A(1'b1), .ZN(_u0_ch30_csr[11] ) );
INV_X4 _u0_U8173  ( .A(1'b1), .ZN(_u0_ch30_csr[10] ) );
INV_X4 _u0_U8171  ( .A(1'b1), .ZN(_u0_ch30_csr[9] ) );
INV_X4 _u0_U8169  ( .A(1'b1), .ZN(_u0_ch30_csr[8] ) );
INV_X4 _u0_U8167  ( .A(1'b1), .ZN(_u0_ch30_csr[7] ) );
INV_X4 _u0_U8165  ( .A(1'b1), .ZN(_u0_ch30_csr[6] ) );
INV_X4 _u0_U8163  ( .A(1'b1), .ZN(_u0_ch30_csr[5] ) );
INV_X4 _u0_U8161  ( .A(1'b1), .ZN(_u0_ch30_csr[4] ) );
INV_X4 _u0_U329  ( .A(1'b1), .ZN(_u0_ch30_csr[3] ) );
INV_X4 _u0_U327  ( .A(1'b1), .ZN(_u0_ch30_csr[2] ) );
INV_X4 _u0_U325  ( .A(1'b1), .ZN(_u0_ch30_csr[1] ) );
INV_X4 _u0_U323  ( .A(1'b1), .ZN(_u0_ch30_csr[0] ) );
INV_X4 _u0_U321  ( .A(1'b1), .ZN(_u0_ch30_txsz[31] ) );
INV_X4 _u0_U319  ( .A(1'b1), .ZN(_u0_ch30_txsz[30] ) );
INV_X4 _u0_U317  ( .A(1'b1), .ZN(_u0_ch30_txsz[29] ) );
INV_X4 _u0_U315  ( .A(1'b1), .ZN(_u0_ch30_txsz[28] ) );
INV_X4 _u0_U313  ( .A(1'b1), .ZN(_u0_ch30_txsz[27] ) );
INV_X4 _u0_U311  ( .A(1'b1), .ZN(_u0_ch30_txsz[26] ) );
INV_X4 _u0_U309  ( .A(1'b1), .ZN(_u0_ch30_txsz[25] ) );
INV_X4 _u0_U307  ( .A(1'b1), .ZN(_u0_ch30_txsz[24] ) );
INV_X4 _u0_U305  ( .A(1'b1), .ZN(_u0_ch30_txsz[23] ) );
INV_X4 _u0_U303  ( .A(1'b1), .ZN(_u0_ch30_txsz[22] ) );
INV_X4 _u0_U301  ( .A(1'b1), .ZN(_u0_ch30_txsz[21] ) );
INV_X4 _u0_U299  ( .A(1'b1), .ZN(_u0_ch30_txsz[20] ) );
INV_X4 _u0_U297  ( .A(1'b1), .ZN(_u0_ch30_txsz[19] ) );
INV_X4 _u0_U295  ( .A(1'b1), .ZN(_u0_ch30_txsz[18] ) );
INV_X4 _u0_U293  ( .A(1'b1), .ZN(_u0_ch30_txsz[17] ) );
INV_X4 _u0_U291  ( .A(1'b1), .ZN(_u0_ch30_txsz[16] ) );
INV_X4 _u0_U289  ( .A(1'b1), .ZN(_u0_ch30_txsz[15] ) );
INV_X4 _u0_U287  ( .A(1'b1), .ZN(_u0_ch30_txsz[14] ) );
INV_X4 _u0_U285  ( .A(1'b1), .ZN(_u0_ch30_txsz[13] ) );
INV_X4 _u0_U283  ( .A(1'b1), .ZN(_u0_ch30_txsz[12] ) );
INV_X4 _u0_U281  ( .A(1'b1), .ZN(_u0_ch30_txsz[11] ) );
INV_X4 _u0_U279  ( .A(1'b1), .ZN(_u0_ch30_txsz[10] ) );
INV_X4 _u0_U277  ( .A(1'b1), .ZN(_u0_ch30_txsz[9] ) );
INV_X4 _u0_U275  ( .A(1'b1), .ZN(_u0_ch30_txsz[8] ) );
INV_X4 _u0_U273  ( .A(1'b1), .ZN(_u0_ch30_txsz[7] ) );
INV_X4 _u0_U271  ( .A(1'b1), .ZN(_u0_ch30_txsz[6] ) );
INV_X4 _u0_U269  ( .A(1'b1), .ZN(_u0_ch30_txsz[5] ) );
INV_X4 _u0_U267  ( .A(1'b1), .ZN(_u0_ch30_txsz[4] ) );
INV_X4 _u0_U265  ( .A(1'b1), .ZN(_u0_ch30_txsz[3] ) );
INV_X4 _u0_U263  ( .A(1'b1), .ZN(_u0_ch30_txsz[2] ) );
INV_X4 _u0_U261  ( .A(1'b1), .ZN(_u0_ch30_txsz[1] ) );
INV_X4 _u0_U259  ( .A(1'b1), .ZN(_u0_ch30_txsz[0] ) );
INV_X4 _u0_U257  ( .A(1'b1), .ZN(_u0_ch30_adr0[31] ) );
INV_X4 _u0_U255  ( .A(1'b1), .ZN(_u0_ch30_adr0[30] ) );
INV_X4 _u0_U253  ( .A(1'b1), .ZN(_u0_ch30_adr0[29] ) );
INV_X4 _u0_U251  ( .A(1'b1), .ZN(_u0_ch30_adr0[28] ) );
INV_X4 _u0_U249  ( .A(1'b1), .ZN(_u0_ch30_adr0[27] ) );
INV_X4 _u0_U247  ( .A(1'b1), .ZN(_u0_ch30_adr0[26] ) );
INV_X4 _u0_U245  ( .A(1'b1), .ZN(_u0_ch30_adr0[25] ) );
INV_X4 _u0_U243  ( .A(1'b1), .ZN(_u0_ch30_adr0[24] ) );
INV_X4 _u0_U241  ( .A(1'b1), .ZN(_u0_ch30_adr0[23] ) );
INV_X4 _u0_U239  ( .A(1'b1), .ZN(_u0_ch30_adr0[22] ) );
INV_X4 _u0_U237  ( .A(1'b1), .ZN(_u0_ch30_adr0[21] ) );
INV_X4 _u0_U235  ( .A(1'b1), .ZN(_u0_ch30_adr0[20] ) );
INV_X4 _u0_U233  ( .A(1'b1), .ZN(_u0_ch30_adr0[19] ) );
INV_X4 _u0_U231  ( .A(1'b1), .ZN(_u0_ch30_adr0[18] ) );
INV_X4 _u0_U229  ( .A(1'b1), .ZN(_u0_ch30_adr0[17] ) );
INV_X4 _u0_U227  ( .A(1'b1), .ZN(_u0_ch30_adr0[16] ) );
INV_X4 _u0_U225  ( .A(1'b1), .ZN(_u0_ch30_adr0[15] ) );
INV_X4 _u0_U223  ( .A(1'b1), .ZN(_u0_ch30_adr0[14] ) );
INV_X4 _u0_U221  ( .A(1'b1), .ZN(_u0_ch30_adr0[13] ) );
INV_X4 _u0_U219  ( .A(1'b1), .ZN(_u0_ch30_adr0[12] ) );
INV_X4 _u0_U217  ( .A(1'b1), .ZN(_u0_ch30_adr0[11] ) );
INV_X4 _u0_U215  ( .A(1'b1), .ZN(_u0_ch30_adr0[10] ) );
INV_X4 _u0_U213  ( .A(1'b1), .ZN(_u0_ch30_adr0[9] ) );
INV_X4 _u0_U211  ( .A(1'b1), .ZN(_u0_ch30_adr0[8] ) );
INV_X4 _u0_U209  ( .A(1'b1), .ZN(_u0_ch30_adr0[7] ) );
INV_X4 _u0_U207  ( .A(1'b1), .ZN(_u0_ch30_adr0[6] ) );
INV_X4 _u0_U205  ( .A(1'b1), .ZN(_u0_ch30_adr0[5] ) );
INV_X4 _u0_U203  ( .A(1'b1), .ZN(_u0_ch30_adr0[4] ) );
INV_X4 _u0_U201  ( .A(1'b1), .ZN(_u0_ch30_adr0[3] ) );
INV_X4 _u0_U199  ( .A(1'b1), .ZN(_u0_ch30_adr0[2] ) );
INV_X4 _u0_U197  ( .A(1'b1), .ZN(_u0_ch30_adr0[1] ) );
INV_X4 _u0_U195  ( .A(1'b1), .ZN(_u0_ch30_adr0[0] ) );
INV_X4 _u0_U193  ( .A(1'b1), .ZN(_u0_ch30_adr1[31] ) );
INV_X4 _u0_U191  ( .A(1'b1), .ZN(_u0_ch30_adr1[30] ) );
INV_X4 _u0_U189  ( .A(1'b1), .ZN(_u0_ch30_adr1[29] ) );
INV_X4 _u0_U187  ( .A(1'b1), .ZN(_u0_ch30_adr1[28] ) );
INV_X4 _u0_U185  ( .A(1'b1), .ZN(_u0_ch30_adr1[27] ) );
INV_X4 _u0_U183  ( .A(1'b1), .ZN(_u0_ch30_adr1[26] ) );
INV_X4 _u0_U181  ( .A(1'b1), .ZN(_u0_ch30_adr1[25] ) );
INV_X4 _u0_U179  ( .A(1'b1), .ZN(_u0_ch30_adr1[24] ) );
INV_X4 _u0_U177  ( .A(1'b1), .ZN(_u0_ch30_adr1[23] ) );
INV_X4 _u0_U175  ( .A(1'b1), .ZN(_u0_ch30_adr1[22] ) );
INV_X4 _u0_U173  ( .A(1'b1), .ZN(_u0_ch30_adr1[21] ) );
INV_X4 _u0_U171  ( .A(1'b1), .ZN(_u0_ch30_adr1[20] ) );
INV_X4 _u0_U169  ( .A(1'b1), .ZN(_u0_ch30_adr1[19] ) );
INV_X4 _u0_U167  ( .A(1'b1), .ZN(_u0_ch30_adr1[18] ) );
INV_X4 _u0_U165  ( .A(1'b1), .ZN(_u0_ch30_adr1[17] ) );
INV_X4 _u0_U163  ( .A(1'b1), .ZN(_u0_ch30_adr1[16] ) );
INV_X4 _u0_U161  ( .A(1'b1), .ZN(_u0_ch30_adr1[15] ) );
INV_X4 _u0_U159  ( .A(1'b1), .ZN(_u0_ch30_adr1[14] ) );
INV_X4 _u0_U157  ( .A(1'b1), .ZN(_u0_ch30_adr1[13] ) );
INV_X4 _u0_U155  ( .A(1'b1), .ZN(_u0_ch30_adr1[12] ) );
INV_X4 _u0_U153  ( .A(1'b1), .ZN(_u0_ch30_adr1[11] ) );
INV_X4 _u0_U151  ( .A(1'b1), .ZN(_u0_ch30_adr1[10] ) );
INV_X4 _u0_U149  ( .A(1'b1), .ZN(_u0_ch30_adr1[9] ) );
INV_X4 _u0_U147  ( .A(1'b1), .ZN(_u0_ch30_adr1[8] ) );
INV_X4 _u0_U145  ( .A(1'b1), .ZN(_u0_ch30_adr1[7] ) );
INV_X4 _u0_U143  ( .A(1'b1), .ZN(_u0_ch30_adr1[6] ) );
INV_X4 _u0_U141  ( .A(1'b1), .ZN(_u0_ch30_adr1[5] ) );
INV_X4 _u0_U139  ( .A(1'b1), .ZN(_u0_ch30_adr1[4] ) );
INV_X4 _u0_U137  ( .A(1'b1), .ZN(_u0_ch30_adr1[3] ) );
INV_X4 _u0_U135  ( .A(1'b1), .ZN(_u0_ch30_adr1[2] ) );
INV_X4 _u0_U133  ( .A(1'b1), .ZN(_u0_ch30_adr1[1] ) );
INV_X4 _u0_U131  ( .A(1'b1), .ZN(_u0_ch30_adr1[0] ) );
INV_X4 _u0_U129  ( .A(1'b0), .ZN(_u0_ch30_am0[31] ) );
INV_X4 _u0_U127  ( .A(1'b0), .ZN(_u0_ch30_am0[30] ) );
INV_X4 _u0_U125  ( .A(1'b0), .ZN(_u0_ch30_am0[29] ) );
INV_X4 _u0_U123  ( .A(1'b0), .ZN(_u0_ch30_am0[28] ) );
INV_X4 _u0_U121  ( .A(1'b0), .ZN(_u0_ch30_am0[27] ) );
INV_X4 _u0_U119  ( .A(1'b0), .ZN(_u0_ch30_am0[26] ) );
INV_X4 _u0_U117  ( .A(1'b0), .ZN(_u0_ch30_am0[25] ) );
INV_X4 _u0_U115  ( .A(1'b0), .ZN(_u0_ch30_am0[24] ) );
INV_X4 _u0_U113  ( .A(1'b0), .ZN(_u0_ch30_am0[23] ) );
INV_X4 _u0_U111  ( .A(1'b0), .ZN(_u0_ch30_am0[22] ) );
INV_X4 _u0_U109  ( .A(1'b0), .ZN(_u0_ch30_am0[21] ) );
INV_X4 _u0_U107  ( .A(1'b0), .ZN(_u0_ch30_am0[20] ) );
INV_X4 _u0_U105  ( .A(1'b0), .ZN(_u0_ch30_am0[19] ) );
INV_X4 _u0_U103  ( .A(1'b0), .ZN(_u0_ch30_am0[18] ) );
INV_X4 _u0_U101  ( .A(1'b0), .ZN(_u0_ch30_am0[17] ) );
INV_X4 _u0_U99  ( .A(1'b0), .ZN(_u0_ch30_am0[16] ) );
INV_X4 _u0_U97  ( .A(1'b0), .ZN(_u0_ch30_am0[15] ) );
INV_X4 _u0_U95  ( .A(1'b0), .ZN(_u0_ch30_am0[14] ) );
INV_X4 _u0_U93  ( .A(1'b0), .ZN(_u0_ch30_am0[13] ) );
INV_X4 _u0_U91  ( .A(1'b0), .ZN(_u0_ch30_am0[12] ) );
INV_X4 _u0_U89  ( .A(1'b0), .ZN(_u0_ch30_am0[11] ) );
INV_X4 _u0_U87  ( .A(1'b0), .ZN(_u0_ch30_am0[10] ) );
INV_X4 _u0_U85  ( .A(1'b0), .ZN(_u0_ch30_am0[9] ) );
INV_X4 _u0_U83  ( .A(1'b0), .ZN(_u0_ch30_am0[8] ) );
INV_X4 _u0_U81  ( .A(1'b0), .ZN(_u0_ch30_am0[7] ) );
INV_X4 _u0_U79  ( .A(1'b0), .ZN(_u0_ch30_am0[6] ) );
INV_X4 _u0_U77  ( .A(1'b0), .ZN(_u0_ch30_am0[5] ) );
INV_X4 _u0_U75  ( .A(1'b0), .ZN(_u0_ch30_am0[4] ) );
INV_X4 _u0_U73  ( .A(1'b1), .ZN(_u0_ch30_am0[3] ) );
INV_X4 _u0_U71  ( .A(1'b1), .ZN(_u0_ch30_am0[2] ) );
INV_X4 _u0_U69  ( .A(1'b1), .ZN(_u0_ch30_am0[1] ) );
INV_X4 _u0_U67  ( .A(1'b1), .ZN(_u0_ch30_am0[0] ) );
INV_X4 _u0_U65  ( .A(1'b0), .ZN(_u0_ch30_am1[31] ) );
INV_X4 _u0_U63  ( .A(1'b0), .ZN(_u0_ch30_am1[30] ) );
INV_X4 _u0_U61  ( .A(1'b0), .ZN(_u0_ch30_am1[29] ) );
INV_X4 _u0_U59  ( .A(1'b0), .ZN(_u0_ch30_am1[28] ) );
INV_X4 _u0_U57  ( .A(1'b0), .ZN(_u0_ch30_am1[27] ) );
INV_X4 _u0_U55  ( .A(1'b0), .ZN(_u0_ch30_am1[26] ) );
INV_X4 _u0_U53  ( .A(1'b0), .ZN(_u0_ch30_am1[25] ) );
INV_X4 _u0_U51  ( .A(1'b0), .ZN(_u0_ch30_am1[24] ) );
INV_X4 _u0_U49  ( .A(1'b0), .ZN(_u0_ch30_am1[23] ) );
INV_X4 _u0_U47  ( .A(1'b0), .ZN(_u0_ch30_am1[22] ) );
INV_X4 _u0_U45  ( .A(1'b0), .ZN(_u0_ch30_am1[21] ) );
INV_X4 _u0_U43  ( .A(1'b0), .ZN(_u0_ch30_am1[20] ) );
INV_X4 _u0_U41  ( .A(1'b0), .ZN(_u0_ch30_am1[19] ) );
INV_X4 _u0_U39  ( .A(1'b0), .ZN(_u0_ch30_am1[18] ) );
INV_X4 _u0_U37  ( .A(1'b0), .ZN(_u0_ch30_am1[17] ) );
INV_X4 _u0_U35  ( .A(1'b0), .ZN(_u0_ch30_am1[16] ) );
INV_X4 _u0_U33  ( .A(1'b0), .ZN(_u0_ch30_am1[15] ) );
INV_X4 _u0_U3100  ( .A(1'b0), .ZN(_u0_ch30_am1[14] ) );
INV_X4 _u0_U2900  ( .A(1'b0), .ZN(_u0_ch30_am1[13] ) );
INV_X4 _u0_U2700  ( .A(1'b0), .ZN(_u0_ch30_am1[12] ) );
INV_X4 _u0_U2500  ( .A(1'b0), .ZN(_u0_ch30_am1[11] ) );
INV_X4 _u0_U2300  ( .A(1'b0), .ZN(_u0_ch30_am1[10] ) );
INV_X4 _u0_U2100  ( .A(1'b0), .ZN(_u0_ch30_am1[9] ) );
INV_X4 _u0_U1900  ( .A(1'b0), .ZN(_u0_ch30_am1[8] ) );
INV_X4 _u0_U1700  ( .A(1'b0), .ZN(_u0_ch30_am1[7] ) );
INV_X4 _u0_U1500  ( .A(1'b0), .ZN(_u0_ch30_am1[6] ) );
INV_X4 _u0_U1300  ( .A(1'b0), .ZN(_u0_ch30_am1[5] ) );
INV_X4 _u0_U1100  ( .A(1'b0), .ZN(_u0_ch30_am1[4] ) );
INV_X4 _u0_U900  ( .A(1'b1), .ZN(_u0_ch30_am1[3] ) );
INV_X4 _u0_U700  ( .A(1'b1), .ZN(_u0_ch30_am1[2] ) );
INV_X4 _u0_U500  ( .A(1'b1), .ZN(_u0_ch30_am1[1] ) );
INV_X4 _u0_U3110  ( .A(1'b1), .ZN(_u0_ch30_am1[0] ) );
DFF_X2 _u0_intb_o_reg  ( .D(_u0_n453 ), .CK(clk_i), .Q(intb_o), .QN() );
DFF_X2 _u0_inta_o_reg  ( .D(_u0_N3078 ), .CK(clk_i), .Q(inta_o), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_0_  ( .D(_u0_N3043 ), .CK(clk_i), .Q(slv0_din[0]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_1_  ( .D(_u0_N3044 ), .CK(clk_i), .Q(slv0_din[1]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_2_  ( .D(_u0_N3045 ), .CK(clk_i), .Q(slv0_din[2]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_3_  ( .D(_u0_N3046 ), .CK(clk_i), .Q(slv0_din[3]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_4_  ( .D(_u0_N3047 ), .CK(clk_i), .Q(slv0_din[4]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_5_  ( .D(_u0_N3048 ), .CK(clk_i), .Q(slv0_din[5]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_6_  ( .D(_u0_N3049 ), .CK(clk_i), .Q(slv0_din[6]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_7_  ( .D(_u0_N3050 ), .CK(clk_i), .Q(slv0_din[7]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_8_  ( .D(_u0_N3051 ), .CK(clk_i), .Q(slv0_din[8]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_9_  ( .D(_u0_N3052 ), .CK(clk_i), .Q(slv0_din[9]),.QN() );
DFF_X2 _u0_wb_rf_dout_reg_10_  ( .D(_u0_N3053 ), .CK(clk_i), .Q(slv0_din[10]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_11_  ( .D(_u0_N3054 ), .CK(clk_i), .Q(slv0_din[11]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_12_  ( .D(_u0_N3055 ), .CK(clk_i), .Q(slv0_din[12]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_13_  ( .D(_u0_N3056 ), .CK(clk_i), .Q(slv0_din[13]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_14_  ( .D(_u0_N3057 ), .CK(clk_i), .Q(slv0_din[14]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_15_  ( .D(_u0_N3058 ), .CK(clk_i), .Q(slv0_din[15]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_16_  ( .D(_u0_N3059 ), .CK(clk_i), .Q(slv0_din[16]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_17_  ( .D(_u0_N3060 ), .CK(clk_i), .Q(slv0_din[17]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_18_  ( .D(_u0_N3061 ), .CK(clk_i), .Q(slv0_din[18]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_19_  ( .D(_u0_N3062 ), .CK(clk_i), .Q(slv0_din[19]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_20_  ( .D(_u0_N3063 ), .CK(clk_i), .Q(slv0_din[20]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_21_  ( .D(_u0_N3064 ), .CK(clk_i), .Q(slv0_din[21]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_22_  ( .D(_u0_N3065 ), .CK(clk_i), .Q(slv0_din[22]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_23_  ( .D(_u0_N3066 ), .CK(clk_i), .Q(slv0_din[23]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_24_  ( .D(_u0_N3067 ), .CK(clk_i), .Q(slv0_din[24]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_25_  ( .D(_u0_N3068 ), .CK(clk_i), .Q(slv0_din[25]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_26_  ( .D(_u0_N3069 ), .CK(clk_i), .Q(slv0_din[26]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_27_  ( .D(_u0_N3070 ), .CK(clk_i), .Q(slv0_din[27]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_28_  ( .D(_u0_N3071 ), .CK(clk_i), .Q(slv0_din[28]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_29_  ( .D(_u0_N3072 ), .CK(clk_i), .Q(slv0_din[29]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_30_  ( .D(_u0_N3073 ), .CK(clk_i), .Q(slv0_din[30]), .QN() );
DFF_X2 _u0_wb_rf_dout_reg_31_  ( .D(_u0_N3074 ), .CK(clk_i), .Q(slv0_din[31]), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_0_  ( .D(_u0_n853 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16276 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_1_  ( .D(_u0_n854 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16277 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_2_  ( .D(_u0_n855 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16275 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_3_  ( .D(_u0_n856 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16273 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_4_  ( .D(_u0_n857 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16278 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_5_  ( .D(_u0_n858 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16279 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_6_  ( .D(_u0_n859 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16280 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_7_  ( .D(_u0_n860 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16281 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_8_  ( .D(_u0_n861 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16282 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_9_  ( .D(_u0_n862 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16270 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_10_  ( .D(_u0_n863 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16283 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_11_  ( .D(_u0_n864 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16284 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_12_  ( .D(_u0_n865 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16269 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_13_  ( .D(_u0_n866 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16267 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_14_  ( .D(_u0_n867 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16265 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_15_  ( .D(_u0_n868 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16285 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_16_  ( .D(_u0_n869 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16286 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_17_  ( .D(_u0_n870 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16287 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_18_  ( .D(_u0_n871 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16288 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_19_  ( .D(_u0_n872 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16289 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_20_  ( .D(_u0_n873 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16290 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_21_  ( .D(_u0_n874 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16291 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_22_  ( .D(_u0_n875 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16292 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_23_  ( .D(_u0_n876 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16262 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_24_  ( .D(_u0_n877 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16260 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_25_  ( .D(_u0_n878 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16258 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_26_  ( .D(_u0_n879 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16256 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_27_  ( .D(_u0_n880 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16255 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_28_  ( .D(_u0_n881 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16253 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_29_  ( .D(_u0_n882 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16251 ), .QN() );
DFFR_X1 _u0_int_maskb_r_reg_30_  ( .D(_u0_n883 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16249 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_0_  ( .D(_u0_n884 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16293 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_1_  ( .D(_u0_n885 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16294 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_2_  ( .D(_u0_n886 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16274 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_3_  ( .D(_u0_n887 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16272 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_4_  ( .D(_u0_n888 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16295 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_5_  ( .D(_u0_n889 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16296 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_6_  ( .D(_u0_n890 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16297 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_7_  ( .D(_u0_n891 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16298 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_8_  ( .D(_u0_n892 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16299 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_9_  ( .D(_u0_n893 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16271 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_10_  ( .D(_u0_n894 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16300 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_11_  ( .D(_u0_n895 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16301 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_12_  ( .D(_u0_n896 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16268 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_13_  ( .D(_u0_n897 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16266 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_14_  ( .D(_u0_n898 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16264 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_15_  ( .D(_u0_n899 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16302 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_16_  ( .D(_u0_n900 ), .CK(clk_i), .RN(_u0_n16018 ), .Q(_u0_n16303 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_17_  ( .D(_u0_n901 ), .CK(clk_i), .RN(n5), .Q(_u0_n16304 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_18_  ( .D(_u0_n902 ), .CK(clk_i), .RN(n5), .Q(_u0_n16305 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_19_  ( .D(_u0_n903 ), .CK(clk_i), .RN(n5), .Q(_u0_n16306 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_20_  ( .D(_u0_n904 ), .CK(clk_i), .RN(n5), .Q(_u0_n16307 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_21_  ( .D(_u0_n905 ), .CK(clk_i), .RN(n5), .Q(_u0_n16308 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_22_  ( .D(_u0_n906 ), .CK(clk_i), .RN(n5), .Q(_u0_n16309 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_23_  ( .D(_u0_n907 ), .CK(clk_i), .RN(n5), .Q(_u0_n16263 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_24_  ( .D(_u0_n908 ), .CK(clk_i), .RN(n5), .Q(_u0_n16261 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_25_  ( .D(_u0_n909 ), .CK(clk_i), .RN(n5), .Q(_u0_n16259 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_26_  ( .D(_u0_n910 ), .CK(clk_i), .RN(n5), .Q(_u0_n16257 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_27_  ( .D(_u0_n911 ), .CK(clk_i), .RN(n5), .Q(_u0_n16254 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_28_  ( .D(_u0_n912 ), .CK(clk_i), .RN(n5), .Q(_u0_n16252 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_29_  ( .D(_u0_n913 ), .CK(clk_i), .RN(n5), .Q(_u0_n16250 ), .QN() );
DFFR_X1 _u0_int_maska_r_reg_30_  ( .D(_u0_n914 ), .CK(clk_i), .RN(n5), .Q(_u0_n16248 ), .QN() );
DFFR_X1 _u0_csr_r_reg_0_  ( .D(_u0_n915 ), .CK(clk_i), .RN(n5), .Q(pause_req), .QN() );
OR3_X1 _u0_u0_U809  ( .A1(ch_sel[4]), .A2(ch_sel[3]), .A3(ch_sel[2]), .ZN(_u0_u0_n1025 ) );
NOR3_X1 _u0_u0_U808  ( .A1(ch_sel[1]), .A2(ch_sel[0]), .A3(_u0_u0_n1025 ),.ZN(_u0_u0_n771 ) );
AND2_X1 _u0_u0_U807  ( .A1(dma_busy), .A2(_u0_u0_n771 ), .ZN(_u0_u0_N23 ) );
INV_X1 _u0_u0_U806  ( .A(slv0_adr[6]), .ZN(_u0_u0_n1023 ) );
NOR3_X1 _u0_u0_U805  ( .A1(slv0_adr[7]), .A2(slv0_adr[9]), .A3(slv0_adr[8]),.ZN(_u0_u0_n1024 ) );
AND3_X1 _u0_u0_U804  ( .A1(slv0_adr[5]), .A2(_u0_u0_n1023 ), .A3(_u0_u0_n1024 ), .ZN(_u0_u0_n787 ) );
INV_X1 _u0_u0_U803  ( .A(slv0_adr[4]), .ZN(_u0_u0_n788 ) );
NAND3_X1 _u0_u0_U802  ( .A1(_u0_u0_n787 ), .A2(_u0_u0_n788 ), .A3(slv0_we),.ZN(_u0_u0_n1019 ) );
INV_X1 _u0_u0_U801  ( .A(_u0_u0_n1019 ), .ZN(_u0_u0_n923 ) );
NOR2_X1 _u0_u0_U800  ( .A1(slv0_adr[3]), .A2(slv0_adr[2]), .ZN(_u0_u0_n786 ));
NAND2_X1 _u0_u0_U799  ( .A1(_u0_u0_n923 ), .A2(_u0_u0_n786 ), .ZN(_u0_u0_n770 ) );
AND2_X1 _u0_u0_U798  ( .A1(_u0_u0_n757 ), .A2(slv0_dout[9]), .ZN(_u0_u0_N24 ) );
NAND2_X1 _u0_u0_U797  ( .A1(ch0_csr[19]), .A2(ch0_csr[22]), .ZN(_u0_u0_n1020 ) );
NAND2_X1 _u0_u0_U796  ( .A1(ch0_csr[17]), .A2(ch0_csr[20]), .ZN(_u0_u0_n1021 ) );
NAND2_X1 _u0_u0_U795  ( .A1(ch0_csr[18]), .A2(ch0_csr[21]), .ZN(_u0_u0_n1022 ) );
NAND3_X1 _u0_u0_U794  ( .A1(_u0_u0_n1020 ), .A2(_u0_u0_n1021 ), .A3(_u0_u0_n1022 ), .ZN(_u0_ch_int_0_ ) );
INV_X1 _u0_u0_U793  ( .A(slv0_adr[2]), .ZN(_u0_u0_n924 ) );
MUX2_X1 _u0_u0_U792  ( .A(ch0_txsz[15]), .B(slv0_dout[15]), .S(_u0_u0_n792 ),.Z(_u0_u0_n335 ) );
MUX2_X1 _u0_u0_U791  ( .A(ch0_csr[17]), .B(slv0_dout[17]), .S(_u0_u0_n757 ),.Z(_u0_u0_n336 ) );
MUX2_X1 _u0_u0_U790  ( .A(ch0_csr[18]), .B(slv0_dout[18]), .S(_u0_u0_n757 ),.Z(_u0_u0_n337 ) );
MUX2_X1 _u0_u0_U789  ( .A(ch0_csr[19]), .B(slv0_dout[19]), .S(_u0_u0_n757 ),.Z(_u0_u0_n338 ) );
MUX2_X1 _u0_u0_U788  ( .A(ch0_csr[16]), .B(slv0_dout[16]), .S(_u0_u0_n757 ),.Z(_u0_u0_n339 ) );
MUX2_X1 _u0_u0_U787  ( .A(ch0_csr[13]), .B(slv0_dout[13]), .S(_u0_u0_n757 ),.Z(_u0_u0_n340 ) );
MUX2_X1 _u0_u0_U786  ( .A(ch0_csr[14]), .B(slv0_dout[14]), .S(_u0_u0_n757 ),.Z(_u0_u0_n341 ) );
MUX2_X1 _u0_u0_U785  ( .A(ch0_csr[15]), .B(slv0_dout[15]), .S(_u0_u0_n757 ),.Z(_u0_u0_n342 ) );
MUX2_X1 _u0_u0_U784  ( .A(ch0_csr[5]), .B(slv0_dout[5]), .S(_u0_u0_n757 ),.Z(_u0_u0_n343 ) );
MUX2_X1 _u0_u0_U783  ( .A(ch0_csr[6]), .B(slv0_dout[6]), .S(_u0_u0_n757 ),.Z(_u0_u0_n344 ) );
MUX2_X1 _u0_u0_U782  ( .A(ch0_csr[7]), .B(slv0_dout[7]), .S(_u0_u0_n757 ),.Z(_u0_u0_n345 ) );
MUX2_X1 _u0_u0_U781  ( .A(ch0_csr[8]), .B(slv0_dout[8]), .S(_u0_u0_n757 ),.Z(_u0_u0_n346 ) );
NAND4_X1 _u0_u0_U780  ( .A1(slv0_adr[4]), .A2(_u0_u0_n786 ), .A3(slv0_we),.A4(_u0_u0_n787 ), .ZN(_u0_u0_n1018 ) );
NAND2_X1 _u0_u0_U779  ( .A1(de_adr1[2]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n1015 ) );
NAND2_X1 _u0_u0_U778  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[2]), .ZN(_u0_u0_n1016 ) );
NAND2_X1 _u0_u0_U777  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[2]), .ZN(_u0_u0_n1017 ) );
NAND3_X1 _u0_u0_U776  ( .A1(_u0_u0_n1015 ), .A2(_u0_u0_n1016 ), .A3(_u0_u0_n1017 ), .ZN(_u0_u0_n347 ) );
NAND2_X1 _u0_u0_U775  ( .A1(de_adr1[3]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n1012 ) );
NAND2_X1 _u0_u0_U774  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[3]), .ZN(_u0_u0_n1013 ) );
NAND2_X1 _u0_u0_U773  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[3]), .ZN(_u0_u0_n1014 ) );
NAND3_X1 _u0_u0_U772  ( .A1(_u0_u0_n1012 ), .A2(_u0_u0_n1013 ), .A3(_u0_u0_n1014 ), .ZN(_u0_u0_n348 ) );
NAND2_X1 _u0_u0_U771  ( .A1(de_adr1[4]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n1009 ) );
NAND2_X1 _u0_u0_U770  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[4]), .ZN(_u0_u0_n1010 ) );
NAND2_X1 _u0_u0_U769  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[4]), .ZN(_u0_u0_n1011 ) );
NAND3_X1 _u0_u0_U768  ( .A1(_u0_u0_n1009 ), .A2(_u0_u0_n1010 ), .A3(_u0_u0_n1011 ), .ZN(_u0_u0_n349 ) );
NAND2_X1 _u0_u0_U767  ( .A1(de_adr1[5]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n1006 ) );
NAND2_X1 _u0_u0_U766  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[5]), .ZN(_u0_u0_n1007 ) );
NAND2_X1 _u0_u0_U765  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[5]), .ZN(_u0_u0_n1008 ) );
NAND3_X1 _u0_u0_U764  ( .A1(_u0_u0_n1006 ), .A2(_u0_u0_n1007 ), .A3(_u0_u0_n1008 ), .ZN(_u0_u0_n350 ) );
NAND2_X1 _u0_u0_U763  ( .A1(de_adr1[6]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n1003 ) );
NAND2_X1 _u0_u0_U762  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[6]), .ZN(_u0_u0_n1004 ) );
NAND2_X1 _u0_u0_U761  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[6]), .ZN(_u0_u0_n1005 ) );
NAND3_X1 _u0_u0_U760  ( .A1(_u0_u0_n1003 ), .A2(_u0_u0_n1004 ), .A3(_u0_u0_n1005 ), .ZN(_u0_u0_n351 ) );
NAND2_X1 _u0_u0_U759  ( .A1(de_adr1[7]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n1000 ) );
NAND2_X1 _u0_u0_U758  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[7]), .ZN(_u0_u0_n1001 ) );
NAND2_X1 _u0_u0_U757  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[7]), .ZN(_u0_u0_n1002 ) );
NAND3_X1 _u0_u0_U756  ( .A1(_u0_u0_n1000 ), .A2(_u0_u0_n1001 ), .A3(_u0_u0_n1002 ), .ZN(_u0_u0_n352 ) );
NAND2_X1 _u0_u0_U755  ( .A1(de_adr1[8]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n997 ) );
NAND2_X1 _u0_u0_U754  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[8]), .ZN(_u0_u0_n998 ) );
NAND2_X1 _u0_u0_U753  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[8]), .ZN(_u0_u0_n999 ) );
NAND3_X1 _u0_u0_U752  ( .A1(_u0_u0_n997 ), .A2(_u0_u0_n998 ), .A3(_u0_u0_n999 ), .ZN(_u0_u0_n353 ) );
NAND2_X1 _u0_u0_U751  ( .A1(de_adr1[9]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n994 ) );
NAND2_X1 _u0_u0_U750  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[9]), .ZN(_u0_u0_n995 ) );
NAND2_X1 _u0_u0_U749  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[9]), .ZN(_u0_u0_n996 ) );
NAND3_X1 _u0_u0_U748  ( .A1(_u0_u0_n994 ), .A2(_u0_u0_n995 ), .A3(_u0_u0_n996 ), .ZN(_u0_u0_n354 ) );
NAND2_X1 _u0_u0_U747  ( .A1(de_adr1[10]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n991 ) );
NAND2_X1 _u0_u0_U746  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[10]), .ZN(_u0_u0_n992 ) );
NAND2_X1 _u0_u0_U745  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[10]), .ZN(_u0_u0_n993 ) );
NAND3_X1 _u0_u0_U744  ( .A1(_u0_u0_n991 ), .A2(_u0_u0_n992 ), .A3(_u0_u0_n993 ), .ZN(_u0_u0_n355 ) );
NAND2_X1 _u0_u0_U743  ( .A1(de_adr1[11]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n988 ) );
NAND2_X1 _u0_u0_U742  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[11]), .ZN(_u0_u0_n989 ) );
NAND2_X1 _u0_u0_U741  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[11]), .ZN(_u0_u0_n990 ) );
NAND3_X1 _u0_u0_U740  ( .A1(_u0_u0_n988 ), .A2(_u0_u0_n989 ), .A3(_u0_u0_n990 ), .ZN(_u0_u0_n356 ) );
NAND2_X1 _u0_u0_U739  ( .A1(de_adr1[12]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n985 ) );
NAND2_X1 _u0_u0_U738  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[12]), .ZN(_u0_u0_n986 ) );
NAND2_X1 _u0_u0_U737  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[12]), .ZN(_u0_u0_n987 ) );
NAND3_X1 _u0_u0_U736  ( .A1(_u0_u0_n985 ), .A2(_u0_u0_n986 ), .A3(_u0_u0_n987 ), .ZN(_u0_u0_n357 ) );
NAND2_X1 _u0_u0_U735  ( .A1(de_adr1[13]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n982 ) );
NAND2_X1 _u0_u0_U734  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[13]), .ZN(_u0_u0_n983 ) );
NAND2_X1 _u0_u0_U733  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[13]), .ZN(_u0_u0_n984 ) );
NAND3_X1 _u0_u0_U732  ( .A1(_u0_u0_n982 ), .A2(_u0_u0_n983 ), .A3(_u0_u0_n984 ), .ZN(_u0_u0_n358 ) );
NAND2_X1 _u0_u0_U731  ( .A1(de_adr1[14]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n979 ) );
NAND2_X1 _u0_u0_U730  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[14]), .ZN(_u0_u0_n980 ) );
NAND2_X1 _u0_u0_U729  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[14]), .ZN(_u0_u0_n981 ) );
NAND3_X1 _u0_u0_U728  ( .A1(_u0_u0_n979 ), .A2(_u0_u0_n980 ), .A3(_u0_u0_n981 ), .ZN(_u0_u0_n359 ) );
NAND2_X1 _u0_u0_U727  ( .A1(de_adr1[15]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n976 ) );
NAND2_X1 _u0_u0_U726  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[15]), .ZN(_u0_u0_n977 ) );
NAND2_X1 _u0_u0_U725  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[15]), .ZN(_u0_u0_n978 ) );
NAND3_X1 _u0_u0_U724  ( .A1(_u0_u0_n976 ), .A2(_u0_u0_n977 ), .A3(_u0_u0_n978 ), .ZN(_u0_u0_n360 ) );
NAND2_X1 _u0_u0_U723  ( .A1(de_adr1[16]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n973 ) );
NAND2_X1 _u0_u0_U722  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[16]), .ZN(_u0_u0_n974 ) );
NAND2_X1 _u0_u0_U721  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[16]), .ZN(_u0_u0_n975 ) );
NAND3_X1 _u0_u0_U720  ( .A1(_u0_u0_n973 ), .A2(_u0_u0_n974 ), .A3(_u0_u0_n975 ), .ZN(_u0_u0_n361 ) );
NAND2_X1 _u0_u0_U719  ( .A1(de_adr1[17]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n970 ) );
NAND2_X1 _u0_u0_U718  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[17]), .ZN(_u0_u0_n971 ) );
NAND2_X1 _u0_u0_U717  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[17]), .ZN(_u0_u0_n972 ) );
NAND3_X1 _u0_u0_U716  ( .A1(_u0_u0_n970 ), .A2(_u0_u0_n971 ), .A3(_u0_u0_n972 ), .ZN(_u0_u0_n362 ) );
NAND2_X1 _u0_u0_U715  ( .A1(de_adr1[18]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n967 ) );
NAND2_X1 _u0_u0_U714  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[18]), .ZN(_u0_u0_n968 ) );
NAND2_X1 _u0_u0_U713  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[18]), .ZN(_u0_u0_n969 ) );
NAND3_X1 _u0_u0_U712  ( .A1(_u0_u0_n967 ), .A2(_u0_u0_n968 ), .A3(_u0_u0_n969 ), .ZN(_u0_u0_n363 ) );
NAND2_X1 _u0_u0_U711  ( .A1(de_adr1[19]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n964 ) );
NAND2_X1 _u0_u0_U710  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[19]), .ZN(_u0_u0_n965 ) );
NAND2_X1 _u0_u0_U709  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[19]), .ZN(_u0_u0_n966 ) );
NAND3_X1 _u0_u0_U708  ( .A1(_u0_u0_n964 ), .A2(_u0_u0_n965 ), .A3(_u0_u0_n966 ), .ZN(_u0_u0_n364 ) );
NAND2_X1 _u0_u0_U707  ( .A1(de_adr1[20]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n961 ) );
NAND2_X1 _u0_u0_U706  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[20]), .ZN(_u0_u0_n962 ) );
NAND2_X1 _u0_u0_U705  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[20]), .ZN(_u0_u0_n963 ) );
NAND3_X1 _u0_u0_U704  ( .A1(_u0_u0_n961 ), .A2(_u0_u0_n962 ), .A3(_u0_u0_n963 ), .ZN(_u0_u0_n365 ) );
NAND2_X1 _u0_u0_U703  ( .A1(de_adr1[21]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n958 ) );
NAND2_X1 _u0_u0_U702  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[21]), .ZN(_u0_u0_n959 ) );
NAND2_X1 _u0_u0_U701  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[21]), .ZN(_u0_u0_n960 ) );
NAND3_X1 _u0_u0_U700  ( .A1(_u0_u0_n958 ), .A2(_u0_u0_n959 ), .A3(_u0_u0_n960 ), .ZN(_u0_u0_n366 ) );
NAND2_X1 _u0_u0_U699  ( .A1(de_adr1[22]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n955 ) );
NAND2_X1 _u0_u0_U698  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[22]), .ZN(_u0_u0_n956 ) );
NAND2_X1 _u0_u0_U697  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[22]), .ZN(_u0_u0_n957 ) );
NAND3_X1 _u0_u0_U696  ( .A1(_u0_u0_n955 ), .A2(_u0_u0_n956 ), .A3(_u0_u0_n957 ), .ZN(_u0_u0_n367 ) );
NAND2_X1 _u0_u0_U695  ( .A1(de_adr1[23]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n952 ) );
NAND2_X1 _u0_u0_U694  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[23]), .ZN(_u0_u0_n953 ) );
NAND2_X1 _u0_u0_U693  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[23]), .ZN(_u0_u0_n954 ) );
NAND3_X1 _u0_u0_U692  ( .A1(_u0_u0_n952 ), .A2(_u0_u0_n953 ), .A3(_u0_u0_n954 ), .ZN(_u0_u0_n368 ) );
NAND2_X1 _u0_u0_U691  ( .A1(de_adr1[24]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n949 ) );
NAND2_X1 _u0_u0_U690  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[24]), .ZN(_u0_u0_n950 ) );
NAND2_X1 _u0_u0_U689  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[24]), .ZN(_u0_u0_n951 ) );
NAND3_X1 _u0_u0_U688  ( .A1(_u0_u0_n949 ), .A2(_u0_u0_n950 ), .A3(_u0_u0_n951 ), .ZN(_u0_u0_n369 ) );
NAND2_X1 _u0_u0_U687  ( .A1(de_adr1[25]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n946 ) );
NAND2_X1 _u0_u0_U686  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[25]), .ZN(_u0_u0_n947 ) );
NAND2_X1 _u0_u0_U685  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[25]), .ZN(_u0_u0_n948 ) );
NAND3_X1 _u0_u0_U684  ( .A1(_u0_u0_n946 ), .A2(_u0_u0_n947 ), .A3(_u0_u0_n948 ), .ZN(_u0_u0_n370 ) );
NAND2_X1 _u0_u0_U683  ( .A1(de_adr1[26]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n943 ) );
NAND2_X1 _u0_u0_U682  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[26]), .ZN(_u0_u0_n944 ) );
NAND2_X1 _u0_u0_U681  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[26]), .ZN(_u0_u0_n945 ) );
NAND3_X1 _u0_u0_U680  ( .A1(_u0_u0_n943 ), .A2(_u0_u0_n944 ), .A3(_u0_u0_n945 ), .ZN(_u0_u0_n371 ) );
NAND2_X1 _u0_u0_U679  ( .A1(de_adr1[27]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n940 ) );
NAND2_X1 _u0_u0_U678  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[27]), .ZN(_u0_u0_n941 ) );
NAND2_X1 _u0_u0_U677  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[27]), .ZN(_u0_u0_n942 ) );
NAND3_X1 _u0_u0_U676  ( .A1(_u0_u0_n940 ), .A2(_u0_u0_n941 ), .A3(_u0_u0_n942 ), .ZN(_u0_u0_n372 ) );
NAND2_X1 _u0_u0_U675  ( .A1(de_adr1[28]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n937 ) );
NAND2_X1 _u0_u0_U674  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[28]), .ZN(_u0_u0_n938 ) );
NAND2_X1 _u0_u0_U673  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[28]), .ZN(_u0_u0_n939 ) );
NAND3_X1 _u0_u0_U672  ( .A1(_u0_u0_n937 ), .A2(_u0_u0_n938 ), .A3(_u0_u0_n939 ), .ZN(_u0_u0_n373 ) );
NAND2_X1 _u0_u0_U671  ( .A1(de_adr1[29]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n934 ) );
NAND2_X1 _u0_u0_U670  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[29]), .ZN(_u0_u0_n935 ) );
NAND2_X1 _u0_u0_U669  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[29]), .ZN(_u0_u0_n936 ) );
NAND3_X1 _u0_u0_U668  ( .A1(_u0_u0_n934 ), .A2(_u0_u0_n935 ), .A3(_u0_u0_n936 ), .ZN(_u0_u0_n374 ) );
NAND2_X1 _u0_u0_U667  ( .A1(de_adr1[30]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n931 ) );
NAND2_X1 _u0_u0_U666  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[30]), .ZN(_u0_u0_n932 ) );
NAND2_X1 _u0_u0_U665  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[30]), .ZN(_u0_u0_n933 ) );
NAND3_X1 _u0_u0_U664  ( .A1(_u0_u0_n931 ), .A2(_u0_u0_n932 ), .A3(_u0_u0_n933 ), .ZN(_u0_u0_n375 ) );
NAND2_X1 _u0_u0_U663  ( .A1(de_adr1[31]), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n925 ) );
NAND2_X1 _u0_u0_U662  ( .A1(_u0_u0_n929 ), .A2(ch0_adr1[31]), .ZN(_u0_u0_n926 ) );
NAND2_X1 _u0_u0_U661  ( .A1(_u0_u0_n928 ), .A2(slv0_dout[31]), .ZN(_u0_u0_n927 ) );
NAND3_X1 _u0_u0_U660  ( .A1(_u0_u0_n925 ), .A2(_u0_u0_n926 ), .A3(_u0_u0_n927 ), .ZN(_u0_u0_n376 ) );
NAND3_X1 _u0_u0_U659  ( .A1(_u0_u0_n923 ), .A2(_u0_u0_n924 ), .A3(slv0_adr[3]), .ZN(_u0_u0_n922 ) );
NAND2_X1 _u0_u0_U658  ( .A1(de_adr0[2]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n919 ) );
NAND2_X1 _u0_u0_U657  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[2]), .ZN(_u0_u0_n920 ) );
NAND2_X1 _u0_u0_U656  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[2]), .ZN(_u0_u0_n921 ) );
NAND3_X1 _u0_u0_U655  ( .A1(_u0_u0_n919 ), .A2(_u0_u0_n920 ), .A3(_u0_u0_n921 ), .ZN(_u0_u0_n377 ) );
NAND2_X1 _u0_u0_U654  ( .A1(de_adr0[3]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n916 ) );
NAND2_X1 _u0_u0_U653  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[3]), .ZN(_u0_u0_n917 ) );
NAND2_X1 _u0_u0_U652  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[3]), .ZN(_u0_u0_n918 ) );
NAND3_X1 _u0_u0_U651  ( .A1(_u0_u0_n916 ), .A2(_u0_u0_n917 ), .A3(_u0_u0_n918 ), .ZN(_u0_u0_n378 ) );
NAND2_X1 _u0_u0_U650  ( .A1(de_adr0[4]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n913 ) );
NAND2_X1 _u0_u0_U649  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[4]), .ZN(_u0_u0_n914 ) );
NAND2_X1 _u0_u0_U648  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[4]), .ZN(_u0_u0_n915 ) );
NAND3_X1 _u0_u0_U647  ( .A1(_u0_u0_n913 ), .A2(_u0_u0_n914 ), .A3(_u0_u0_n915 ), .ZN(_u0_u0_n379 ) );
NAND2_X1 _u0_u0_U646  ( .A1(de_adr0[5]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n910 ) );
NAND2_X1 _u0_u0_U645  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[5]), .ZN(_u0_u0_n911 ) );
NAND2_X1 _u0_u0_U644  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[5]), .ZN(_u0_u0_n912 ) );
NAND3_X1 _u0_u0_U643  ( .A1(_u0_u0_n910 ), .A2(_u0_u0_n911 ), .A3(_u0_u0_n912 ), .ZN(_u0_u0_n380 ) );
NAND2_X1 _u0_u0_U642  ( .A1(de_adr0[6]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n907 ) );
NAND2_X1 _u0_u0_U641  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[6]), .ZN(_u0_u0_n908 ) );
NAND2_X1 _u0_u0_U640  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[6]), .ZN(_u0_u0_n909 ) );
NAND3_X1 _u0_u0_U639  ( .A1(_u0_u0_n907 ), .A2(_u0_u0_n908 ), .A3(_u0_u0_n909 ), .ZN(_u0_u0_n381 ) );
NAND2_X1 _u0_u0_U638  ( .A1(de_adr0[7]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n904 ) );
NAND2_X1 _u0_u0_U637  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[7]), .ZN(_u0_u0_n905 ) );
NAND2_X1 _u0_u0_U636  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[7]), .ZN(_u0_u0_n906 ) );
NAND3_X1 _u0_u0_U635  ( .A1(_u0_u0_n904 ), .A2(_u0_u0_n905 ), .A3(_u0_u0_n906 ), .ZN(_u0_u0_n382 ) );
NAND2_X1 _u0_u0_U634  ( .A1(de_adr0[8]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n901 ) );
NAND2_X1 _u0_u0_U633  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[8]), .ZN(_u0_u0_n902 ) );
NAND2_X1 _u0_u0_U632  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[8]), .ZN(_u0_u0_n903 ) );
NAND3_X1 _u0_u0_U631  ( .A1(_u0_u0_n901 ), .A2(_u0_u0_n902 ), .A3(_u0_u0_n903 ), .ZN(_u0_u0_n383 ) );
NAND2_X1 _u0_u0_U630  ( .A1(de_adr0[9]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n898 ) );
NAND2_X1 _u0_u0_U629  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[9]), .ZN(_u0_u0_n899 ) );
NAND2_X1 _u0_u0_U628  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[9]), .ZN(_u0_u0_n900 ) );
NAND3_X1 _u0_u0_U627  ( .A1(_u0_u0_n898 ), .A2(_u0_u0_n899 ), .A3(_u0_u0_n900 ), .ZN(_u0_u0_n384 ) );
NAND2_X1 _u0_u0_U626  ( .A1(de_adr0[10]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n895 ) );
NAND2_X1 _u0_u0_U625  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[10]), .ZN(_u0_u0_n896 ) );
NAND2_X1 _u0_u0_U624  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[10]), .ZN(_u0_u0_n897 ) );
NAND3_X1 _u0_u0_U623  ( .A1(_u0_u0_n895 ), .A2(_u0_u0_n896 ), .A3(_u0_u0_n897 ), .ZN(_u0_u0_n385 ) );
NAND2_X1 _u0_u0_U622  ( .A1(de_adr0[11]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n892 ) );
NAND2_X1 _u0_u0_U621  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[11]), .ZN(_u0_u0_n893 ) );
NAND2_X1 _u0_u0_U620  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[11]), .ZN(_u0_u0_n894 ) );
NAND3_X1 _u0_u0_U619  ( .A1(_u0_u0_n892 ), .A2(_u0_u0_n893 ), .A3(_u0_u0_n894 ), .ZN(_u0_u0_n386 ) );
NAND2_X1 _u0_u0_U618  ( .A1(de_adr0[12]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n889 ) );
NAND2_X1 _u0_u0_U617  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[12]), .ZN(_u0_u0_n890 ) );
NAND2_X1 _u0_u0_U616  ( .A1(slv0_dout[12]), .A2(_u0_u0_n832 ), .ZN(_u0_u0_n891 ) );
NAND3_X1 _u0_u0_U615  ( .A1(_u0_u0_n889 ), .A2(_u0_u0_n890 ), .A3(_u0_u0_n891 ), .ZN(_u0_u0_n387 ) );
NAND2_X1 _u0_u0_U614  ( .A1(de_adr0[13]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n886 ) );
NAND2_X1 _u0_u0_U613  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[13]), .ZN(_u0_u0_n887 ) );
NAND2_X1 _u0_u0_U612  ( .A1(slv0_dout[13]), .A2(_u0_u0_n832 ), .ZN(_u0_u0_n888 ) );
NAND3_X1 _u0_u0_U611  ( .A1(_u0_u0_n886 ), .A2(_u0_u0_n887 ), .A3(_u0_u0_n888 ), .ZN(_u0_u0_n388 ) );
NAND2_X1 _u0_u0_U610  ( .A1(de_adr0[14]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n883 ) );
NAND2_X1 _u0_u0_U609  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[14]), .ZN(_u0_u0_n884 ) );
NAND2_X1 _u0_u0_U608  ( .A1(slv0_dout[14]), .A2(_u0_u0_n832 ), .ZN(_u0_u0_n885 ) );
NAND3_X1 _u0_u0_U607  ( .A1(_u0_u0_n883 ), .A2(_u0_u0_n884 ), .A3(_u0_u0_n885 ), .ZN(_u0_u0_n389 ) );
NAND2_X1 _u0_u0_U606  ( .A1(de_adr0[15]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n880 ) );
NAND2_X1 _u0_u0_U605  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[15]), .ZN(_u0_u0_n881 ) );
NAND2_X1 _u0_u0_U604  ( .A1(slv0_dout[15]), .A2(_u0_u0_n832 ), .ZN(_u0_u0_n882 ) );
NAND3_X1 _u0_u0_U603  ( .A1(_u0_u0_n880 ), .A2(_u0_u0_n881 ), .A3(_u0_u0_n882 ), .ZN(_u0_u0_n390 ) );
NAND2_X1 _u0_u0_U602  ( .A1(de_adr0[16]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n877 ) );
NAND2_X1 _u0_u0_U601  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[16]), .ZN(_u0_u0_n878 ) );
NAND2_X1 _u0_u0_U600  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[16]), .ZN(_u0_u0_n879 ) );
NAND3_X1 _u0_u0_U599  ( .A1(_u0_u0_n877 ), .A2(_u0_u0_n878 ), .A3(_u0_u0_n879 ), .ZN(_u0_u0_n391 ) );
NAND2_X1 _u0_u0_U598  ( .A1(de_adr0[17]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n874 ) );
NAND2_X1 _u0_u0_U597  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[17]), .ZN(_u0_u0_n875 ) );
NAND2_X1 _u0_u0_U596  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[17]), .ZN(_u0_u0_n876 ) );
NAND3_X1 _u0_u0_U595  ( .A1(_u0_u0_n874 ), .A2(_u0_u0_n875 ), .A3(_u0_u0_n876 ), .ZN(_u0_u0_n392 ) );
NAND2_X1 _u0_u0_U594  ( .A1(de_adr0[18]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n871 ) );
NAND2_X1 _u0_u0_U593  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[18]), .ZN(_u0_u0_n872 ) );
NAND2_X1 _u0_u0_U592  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[18]), .ZN(_u0_u0_n873 ) );
NAND3_X1 _u0_u0_U591  ( .A1(_u0_u0_n871 ), .A2(_u0_u0_n872 ), .A3(_u0_u0_n873 ), .ZN(_u0_u0_n393 ) );
NAND2_X1 _u0_u0_U590  ( .A1(de_adr0[19]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n868 ) );
NAND2_X1 _u0_u0_U589  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[19]), .ZN(_u0_u0_n869 ) );
NAND2_X1 _u0_u0_U588  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[19]), .ZN(_u0_u0_n870 ) );
NAND3_X1 _u0_u0_U587  ( .A1(_u0_u0_n868 ), .A2(_u0_u0_n869 ), .A3(_u0_u0_n870 ), .ZN(_u0_u0_n394 ) );
NAND2_X1 _u0_u0_U586  ( .A1(de_adr0[20]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n865 ) );
NAND2_X1 _u0_u0_U585  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[20]), .ZN(_u0_u0_n866 ) );
NAND2_X1 _u0_u0_U584  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[20]), .ZN(_u0_u0_n867 ) );
NAND3_X1 _u0_u0_U583  ( .A1(_u0_u0_n865 ), .A2(_u0_u0_n866 ), .A3(_u0_u0_n867 ), .ZN(_u0_u0_n395 ) );
NAND2_X1 _u0_u0_U582  ( .A1(de_adr0[21]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n862 ) );
NAND2_X1 _u0_u0_U581  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[21]), .ZN(_u0_u0_n863 ) );
NAND2_X1 _u0_u0_U580  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[21]), .ZN(_u0_u0_n864 ) );
NAND3_X1 _u0_u0_U579  ( .A1(_u0_u0_n862 ), .A2(_u0_u0_n863 ), .A3(_u0_u0_n864 ), .ZN(_u0_u0_n396 ) );
NAND2_X1 _u0_u0_U578  ( .A1(de_adr0[22]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n859 ) );
NAND2_X1 _u0_u0_U577  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[22]), .ZN(_u0_u0_n860 ) );
NAND2_X1 _u0_u0_U576  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[22]), .ZN(_u0_u0_n861 ) );
NAND3_X1 _u0_u0_U575  ( .A1(_u0_u0_n859 ), .A2(_u0_u0_n860 ), .A3(_u0_u0_n861 ), .ZN(_u0_u0_n397 ) );
NAND2_X1 _u0_u0_U574  ( .A1(de_adr0[23]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n856 ) );
NAND2_X1 _u0_u0_U573  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[23]), .ZN(_u0_u0_n857 ) );
NAND2_X1 _u0_u0_U572  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[23]), .ZN(_u0_u0_n858 ) );
NAND3_X1 _u0_u0_U571  ( .A1(_u0_u0_n856 ), .A2(_u0_u0_n857 ), .A3(_u0_u0_n858 ), .ZN(_u0_u0_n398 ) );
NAND2_X1 _u0_u0_U570  ( .A1(de_adr0[24]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n853 ) );
NAND2_X1 _u0_u0_U569  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[24]), .ZN(_u0_u0_n854 ) );
NAND2_X1 _u0_u0_U568  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[24]), .ZN(_u0_u0_n855 ) );
NAND3_X1 _u0_u0_U567  ( .A1(_u0_u0_n853 ), .A2(_u0_u0_n854 ), .A3(_u0_u0_n855 ), .ZN(_u0_u0_n399 ) );
NAND2_X1 _u0_u0_U566  ( .A1(de_adr0[25]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n850 ) );
NAND2_X1 _u0_u0_U565  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[25]), .ZN(_u0_u0_n851 ) );
NAND2_X1 _u0_u0_U564  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[25]), .ZN(_u0_u0_n852 ) );
NAND3_X1 _u0_u0_U563  ( .A1(_u0_u0_n850 ), .A2(_u0_u0_n851 ), .A3(_u0_u0_n852 ), .ZN(_u0_u0_n400 ) );
NAND2_X1 _u0_u0_U562  ( .A1(de_adr0[26]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n847 ) );
NAND2_X1 _u0_u0_U561  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[26]), .ZN(_u0_u0_n848 ) );
NAND2_X1 _u0_u0_U560  ( .A1(_u0_u0_n832 ), .A2(slv0_dout[26]), .ZN(_u0_u0_n849 ) );
NAND3_X1 _u0_u0_U559  ( .A1(_u0_u0_n847 ), .A2(_u0_u0_n848 ), .A3(_u0_u0_n849 ), .ZN(_u0_u0_n401 ) );
NAND2_X1 _u0_u0_U558  ( .A1(de_adr0[27]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n844 ) );
NAND2_X1 _u0_u0_U557  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[27]), .ZN(_u0_u0_n845 ) );
NAND2_X1 _u0_u0_U556  ( .A1(slv0_dout[27]), .A2(_u0_u0_n832 ), .ZN(_u0_u0_n846 ) );
NAND3_X1 _u0_u0_U555  ( .A1(_u0_u0_n844 ), .A2(_u0_u0_n845 ), .A3(_u0_u0_n846 ), .ZN(_u0_u0_n402 ) );
NAND2_X1 _u0_u0_U554  ( .A1(de_adr0[28]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n841 ) );
NAND2_X1 _u0_u0_U553  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[28]), .ZN(_u0_u0_n842 ) );
NAND2_X1 _u0_u0_U552  ( .A1(slv0_dout[28]), .A2(_u0_u0_n832 ), .ZN(_u0_u0_n843 ) );
NAND3_X1 _u0_u0_U551  ( .A1(_u0_u0_n841 ), .A2(_u0_u0_n842 ), .A3(_u0_u0_n843 ), .ZN(_u0_u0_n403 ) );
NAND2_X1 _u0_u0_U550  ( .A1(de_adr0[29]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n838 ) );
NAND2_X1 _u0_u0_U549  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[29]), .ZN(_u0_u0_n839 ) );
NAND2_X1 _u0_u0_U548  ( .A1(slv0_dout[29]), .A2(_u0_u0_n832 ), .ZN(_u0_u0_n840 ) );
NAND3_X1 _u0_u0_U547  ( .A1(_u0_u0_n838 ), .A2(_u0_u0_n839 ), .A3(_u0_u0_n840 ), .ZN(_u0_u0_n404 ) );
NAND2_X1 _u0_u0_U546  ( .A1(de_adr0[30]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n835 ) );
NAND2_X1 _u0_u0_U545  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[30]), .ZN(_u0_u0_n836 ) );
NAND2_X1 _u0_u0_U544  ( .A1(slv0_dout[30]), .A2(_u0_u0_n832 ), .ZN(_u0_u0_n837 ) );
NAND3_X1 _u0_u0_U543  ( .A1(_u0_u0_n835 ), .A2(_u0_u0_n836 ), .A3(_u0_u0_n837 ), .ZN(_u0_u0_n405 ) );
NAND2_X1 _u0_u0_U542  ( .A1(de_adr0[31]), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n829 ) );
NAND2_X1 _u0_u0_U541  ( .A1(_u0_u0_n833 ), .A2(ch0_adr0[31]), .ZN(_u0_u0_n830 ) );
NAND2_X1 _u0_u0_U540  ( .A1(slv0_dout[31]), .A2(_u0_u0_n832 ), .ZN(_u0_u0_n831 ) );
NAND3_X1 _u0_u0_U539  ( .A1(_u0_u0_n829 ), .A2(_u0_u0_n830 ), .A3(_u0_u0_n831 ), .ZN(_u0_u0_n406 ) );
MUX2_X1 _u0_u0_U538  ( .A(ch0_txsz[16]), .B(slv0_dout[16]), .S(_u0_u0_n792 ),.Z(_u0_u0_n407 ) );
MUX2_X1 _u0_u0_U537  ( .A(ch0_txsz[17]), .B(slv0_dout[17]), .S(_u0_u0_n792 ),.Z(_u0_u0_n408 ) );
MUX2_X1 _u0_u0_U536  ( .A(ch0_txsz[18]), .B(slv0_dout[18]), .S(_u0_u0_n792 ),.Z(_u0_u0_n409 ) );
MUX2_X1 _u0_u0_U535  ( .A(ch0_txsz[19]), .B(slv0_dout[19]), .S(_u0_u0_n792 ),.Z(_u0_u0_n410 ) );
MUX2_X1 _u0_u0_U534  ( .A(ch0_txsz[20]), .B(slv0_dout[20]), .S(_u0_u0_n792 ),.Z(_u0_u0_n411 ) );
MUX2_X1 _u0_u0_U533  ( .A(ch0_txsz[21]), .B(slv0_dout[21]), .S(_u0_u0_n792 ),.Z(_u0_u0_n412 ) );
MUX2_X1 _u0_u0_U532  ( .A(ch0_txsz[22]), .B(slv0_dout[22]), .S(_u0_u0_n792 ),.Z(_u0_u0_n413 ) );
MUX2_X1 _u0_u0_U531  ( .A(ch0_txsz[23]), .B(slv0_dout[23]), .S(_u0_u0_n792 ),.Z(_u0_u0_n414 ) );
MUX2_X1 _u0_u0_U530  ( .A(ch0_txsz[24]), .B(slv0_dout[24]), .S(_u0_u0_n792 ),.Z(_u0_u0_n415 ) );
MUX2_X1 _u0_u0_U529  ( .A(ch0_txsz[25]), .B(slv0_dout[25]), .S(_u0_u0_n792 ),.Z(_u0_u0_n416 ) );
MUX2_X1 _u0_u0_U528  ( .A(ch0_txsz[26]), .B(slv0_dout[26]), .S(_u0_u0_n792 ),.Z(_u0_u0_n417 ) );
INV_X1 _u0_u0_U527  ( .A(_u0_u0_n792 ), .ZN(_u0_u0_n828 ) );
AND3_X1 _u0_u0_U526  ( .A1(_u0_u0_n771 ), .A2(_u0_u0_n828 ), .A3(de_txsz_we),.ZN(_u0_u0_n794 ) );
NAND2_X1 _u0_u0_U525  ( .A1(de_txsz[0]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n825 ) );
NOR2_X1 _u0_u0_U524  ( .A1(_u0_u0_n792 ), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n793 ) );
NAND2_X1 _u0_u0_U523  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[0]), .ZN(_u0_u0_n826 ) );
NAND2_X1 _u0_u0_U522  ( .A1(_u0_u0_n792 ), .A2(slv0_dout[0]), .ZN(_u0_u0_n827 ) );
NAND3_X1 _u0_u0_U521  ( .A1(_u0_u0_n825 ), .A2(_u0_u0_n826 ), .A3(_u0_u0_n827 ), .ZN(_u0_u0_n418 ) );
NAND2_X1 _u0_u0_U520  ( .A1(de_txsz[1]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n822 ) );
NAND2_X1 _u0_u0_U519  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[1]), .ZN(_u0_u0_n823 ) );
NAND2_X1 _u0_u0_U518  ( .A1(_u0_u0_n792 ), .A2(slv0_dout[1]), .ZN(_u0_u0_n824 ) );
NAND3_X1 _u0_u0_U517  ( .A1(_u0_u0_n822 ), .A2(_u0_u0_n823 ), .A3(_u0_u0_n824 ), .ZN(_u0_u0_n419 ) );
NAND2_X1 _u0_u0_U516  ( .A1(de_txsz[2]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n819 ) );
NAND2_X1 _u0_u0_U515  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[2]), .ZN(_u0_u0_n820 ) );
NAND2_X1 _u0_u0_U514  ( .A1(_u0_u0_n792 ), .A2(slv0_dout[2]), .ZN(_u0_u0_n821 ) );
NAND3_X1 _u0_u0_U513  ( .A1(_u0_u0_n819 ), .A2(_u0_u0_n820 ), .A3(_u0_u0_n821 ), .ZN(_u0_u0_n420 ) );
NAND2_X1 _u0_u0_U512  ( .A1(de_txsz[3]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n816 ) );
NAND2_X1 _u0_u0_U511  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[3]), .ZN(_u0_u0_n817 ) );
NAND2_X1 _u0_u0_U510  ( .A1(_u0_u0_n792 ), .A2(slv0_dout[3]), .ZN(_u0_u0_n818 ) );
NAND3_X1 _u0_u0_U509  ( .A1(_u0_u0_n816 ), .A2(_u0_u0_n817 ), .A3(_u0_u0_n818 ), .ZN(_u0_u0_n421 ) );
NAND2_X1 _u0_u0_U508  ( .A1(de_txsz[4]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n813 ) );
NAND2_X1 _u0_u0_U507  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[4]), .ZN(_u0_u0_n814 ) );
NAND2_X1 _u0_u0_U506  ( .A1(_u0_u0_n792 ), .A2(slv0_dout[4]), .ZN(_u0_u0_n815 ) );
NAND3_X1 _u0_u0_U505  ( .A1(_u0_u0_n813 ), .A2(_u0_u0_n814 ), .A3(_u0_u0_n815 ), .ZN(_u0_u0_n422 ) );
NAND2_X1 _u0_u0_U504  ( .A1(de_txsz[5]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n810 ) );
NAND2_X1 _u0_u0_U503  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[5]), .ZN(_u0_u0_n811 ) );
NAND2_X1 _u0_u0_U502  ( .A1(slv0_dout[5]), .A2(_u0_u0_n792 ), .ZN(_u0_u0_n812 ) );
NAND3_X1 _u0_u0_U501  ( .A1(_u0_u0_n810 ), .A2(_u0_u0_n811 ), .A3(_u0_u0_n812 ), .ZN(_u0_u0_n423 ) );
NAND2_X1 _u0_u0_U500  ( .A1(de_txsz[6]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n807 ) );
NAND2_X1 _u0_u0_U499  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[6]), .ZN(_u0_u0_n808 ) );
NAND2_X1 _u0_u0_U498  ( .A1(slv0_dout[6]), .A2(_u0_u0_n792 ), .ZN(_u0_u0_n809 ) );
NAND3_X1 _u0_u0_U497  ( .A1(_u0_u0_n807 ), .A2(_u0_u0_n808 ), .A3(_u0_u0_n809 ), .ZN(_u0_u0_n424 ) );
NAND2_X1 _u0_u0_U496  ( .A1(de_txsz[7]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n804 ) );
NAND2_X1 _u0_u0_U495  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[7]), .ZN(_u0_u0_n805 ) );
NAND2_X1 _u0_u0_U494  ( .A1(slv0_dout[7]), .A2(_u0_u0_n792 ), .ZN(_u0_u0_n806 ) );
NAND3_X1 _u0_u0_U435  ( .A1(_u0_u0_n804 ), .A2(_u0_u0_n805 ), .A3(_u0_u0_n806 ), .ZN(_u0_u0_n425 ) );
NAND2_X1 _u0_u0_U434  ( .A1(de_txsz[8]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n801 ) );
NAND2_X1 _u0_u0_U433  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[8]), .ZN(_u0_u0_n802 ) );
NAND2_X1 _u0_u0_U432  ( .A1(slv0_dout[8]), .A2(_u0_u0_n792 ), .ZN(_u0_u0_n803 ) );
NAND3_X1 _u0_u0_U431  ( .A1(_u0_u0_n801 ), .A2(_u0_u0_n802 ), .A3(_u0_u0_n803 ), .ZN(_u0_u0_n426 ) );
NAND2_X1 _u0_u0_U430  ( .A1(de_txsz[9]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n798 ) );
NAND2_X1 _u0_u0_U429  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[9]), .ZN(_u0_u0_n799 ) );
NAND2_X1 _u0_u0_U428  ( .A1(slv0_dout[9]), .A2(_u0_u0_n792 ), .ZN(_u0_u0_n800 ) );
NAND3_X1 _u0_u0_U427  ( .A1(_u0_u0_n798 ), .A2(_u0_u0_n799 ), .A3(_u0_u0_n800 ), .ZN(_u0_u0_n427 ) );
NAND2_X1 _u0_u0_U426  ( .A1(de_txsz[10]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n795 ) );
NAND2_X1 _u0_u0_U425  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[10]), .ZN(_u0_u0_n796 ) );
NAND2_X1 _u0_u0_U424  ( .A1(slv0_dout[10]), .A2(_u0_u0_n792 ), .ZN(_u0_u0_n797 ) );
NAND3_X1 _u0_u0_U423  ( .A1(_u0_u0_n795 ), .A2(_u0_u0_n796 ), .A3(_u0_u0_n797 ), .ZN(_u0_u0_n428 ) );
NAND2_X1 _u0_u0_U422  ( .A1(de_txsz[11]), .A2(_u0_u0_n794 ), .ZN(_u0_u0_n789 ) );
NAND2_X1 _u0_u0_U421  ( .A1(_u0_u0_n793 ), .A2(ch0_txsz[11]), .ZN(_u0_u0_n790 ) );
NAND2_X1 _u0_u0_U420  ( .A1(slv0_dout[11]), .A2(_u0_u0_n792 ), .ZN(_u0_u0_n791 ) );
NAND3_X1 _u0_u0_U419  ( .A1(_u0_u0_n789 ), .A2(_u0_u0_n790 ), .A3(_u0_u0_n791 ), .ZN(_u0_u0_n429 ) );
NAND2_X1 _u0_u0_U418  ( .A1(dma_err), .A2(_u0_u0_n771 ), .ZN(_u0_u0_n777 ));
NAND4_X1 _u0_u0_U417  ( .A1(slv0_re), .A2(_u0_u0_n786 ), .A3(_u0_u0_n787 ),.A4(_u0_u0_n788 ), .ZN(_u0_u0_n779 ) );
NAND2_X1 _u0_u0_U416  ( .A1(_u0_u0_n779 ), .A2(ch0_csr[20]), .ZN(_u0_u0_n785 ) );
NAND2_X1 _u0_u0_U415  ( .A1(_u0_u0_n777 ), .A2(_u0_u0_n785 ), .ZN(_u0_u0_n430 ) );
AND2_X1 _u0_u0_U414  ( .A1(dma_done_all), .A2(_u0_u0_n771 ), .ZN(_u0_u0_n784 ) );
OR2_X1 _u0_u0_U413  ( .A1(ndnr[0]), .A2(_u0_u0_n784 ), .ZN(_u0_u0_n783 ) );
NAND3_X1 _u0_u0_U412  ( .A1(_u0_u0_n333 ), .A2(_u0_u0_n783 ), .A3(_u0_u0_n334 ), .ZN(_u0_u0_n774 ) );
NAND2_X1 _u0_u0_U411  ( .A1(_u0_u0_n779 ), .A2(ch0_csr[21]), .ZN(_u0_u0_n782 ) );
NAND2_X1 _u0_u0_U410  ( .A1(_u0_u0_n774 ), .A2(_u0_u0_n782 ), .ZN(_u0_u0_n431 ) );
NAND2_X1 _u0_u0_U409  ( .A1(dma_done), .A2(_u0_u0_n771 ), .ZN(_u0_u0_n780 ));
NAND2_X1 _u0_u0_U408  ( .A1(_u0_u0_n779 ), .A2(ch0_csr[22]), .ZN(_u0_u0_n781 ) );
NAND2_X1 _u0_u0_U407  ( .A1(_u0_u0_n780 ), .A2(_u0_u0_n781 ), .ZN(_u0_u0_n432 ) );
NAND2_X1 _u0_u0_U406  ( .A1(_u0_u0_n779 ), .A2(ch0_csr[12]), .ZN(_u0_u0_n778 ) );
NAND2_X1 _u0_u0_U405  ( .A1(_u0_u0_n777 ), .A2(_u0_u0_n778 ), .ZN(_u0_u0_n433 ) );
NAND2_X1 _u0_u0_U404  ( .A1(_u0_u0_n326 ), .A2(_u0_u0_n774 ), .ZN(_u0_u0_n775 ) );
INV_X1 _u0_u0_U403  ( .A(slv0_dout[0]), .ZN(_u0_u0_n776 ) );
MUX2_X1 _u0_u0_U402  ( .A(_u0_u0_n775 ), .B(_u0_u0_n776 ), .S(_u0_u0_n757 ),.Z(_u0_u0_n434 ) );
INV_X1 _u0_u0_U401  ( .A(_u0_u0_n774 ), .ZN(_u0_u0_n773 ) );
NOR2_X1 _u0_u0_U400  ( .A1(_u0_u0_n1026 ), .A2(_u0_u0_n773 ), .ZN(_u0_u0_n772 ) );
MUX2_X1 _u0_u0_U399  ( .A(_u0_u0_n772 ), .B(slv0_dout[0]), .S(_u0_u0_n757 ),.Z(_u0_u0_n435 ) );
NAND2_X1 _u0_u0_U398  ( .A1(de_csr_we), .A2(_u0_u0_n771 ), .ZN(_u0_u0_n769 ));
AND2_X1 _u0_u0_U397  ( .A1(_u0_u0_n769 ), .A2(_u0_u0_n770 ), .ZN(_u0_u0_n759 ) );
NAND2_X1 _u0_u0_U396  ( .A1(_u0_u0_n759 ), .A2(ch0_csr[1]), .ZN(_u0_u0_n766 ) );
NOR2_X1 _u0_u0_U395  ( .A1(_u0_u0_n757 ), .A2(_u0_u0_n759 ), .ZN(_u0_u0_n758 ) );
NAND2_X1 _u0_u0_U394  ( .A1(de_csr[16]), .A2(_u0_u0_n758 ), .ZN(_u0_u0_n767 ) );
NAND2_X1 _u0_u0_U393  ( .A1(slv0_dout[1]), .A2(_u0_u0_n757 ), .ZN(_u0_u0_n768 ) );
NAND3_X1 _u0_u0_U392  ( .A1(_u0_u0_n766 ), .A2(_u0_u0_n767 ), .A3(_u0_u0_n768 ), .ZN(_u0_u0_n436 ) );
NAND2_X1 _u0_u0_U391  ( .A1(_u0_u0_n759 ), .A2(ch0_csr[2]), .ZN(_u0_u0_n763 ) );
NAND2_X1 _u0_u0_U390  ( .A1(de_csr[17]), .A2(_u0_u0_n758 ), .ZN(_u0_u0_n764 ) );
NAND2_X1 _u0_u0_U389  ( .A1(slv0_dout[2]), .A2(_u0_u0_n757 ), .ZN(_u0_u0_n765 ) );
NAND3_X1 _u0_u0_U388  ( .A1(_u0_u0_n763 ), .A2(_u0_u0_n764 ), .A3(_u0_u0_n765 ), .ZN(_u0_u0_n437 ) );
NAND2_X1 _u0_u0_U387  ( .A1(_u0_u0_n759 ), .A2(ch0_csr[3]), .ZN(_u0_u0_n760 ) );
NAND2_X1 _u0_u0_U386  ( .A1(de_csr[18]), .A2(_u0_u0_n758 ), .ZN(_u0_u0_n761 ) );
NAND2_X1 _u0_u0_U385  ( .A1(slv0_dout[3]), .A2(_u0_u0_n757 ), .ZN(_u0_u0_n762 ) );
NAND3_X1 _u0_u0_U384  ( .A1(_u0_u0_n760 ), .A2(_u0_u0_n761 ), .A3(_u0_u0_n762 ), .ZN(_u0_u0_n438 ) );
NAND2_X1 _u0_u0_U383  ( .A1(_u0_u0_n759 ), .A2(ch0_csr[4]), .ZN(_u0_u0_n754 ) );
NAND2_X1 _u0_u0_U382  ( .A1(de_csr[19]), .A2(_u0_u0_n758 ), .ZN(_u0_u0_n755 ) );
NAND2_X1 _u0_u0_U381  ( .A1(slv0_dout[4]), .A2(_u0_u0_n757 ), .ZN(_u0_u0_n756 ) );
NAND3_X1 _u0_u0_U380  ( .A1(_u0_u0_n754 ), .A2(_u0_u0_n755 ), .A3(_u0_u0_n756 ), .ZN(_u0_u0_n439 ) );
INV_X4 _u0_u0_U379  ( .A(_u0_n16018 ), .ZN(_u0_u0_n753 ) );
INV_X4 _u0_u0_U378  ( .A(_u0_u0_n753 ), .ZN(_u0_u0_n752 ) );
INV_X4 _u0_u0_U377  ( .A(_u0_u0_n753 ), .ZN(_u0_u0_n751 ) );
NOR3_X2 _u0_u0_U376  ( .A1(_u0_u0_n1019 ), .A2(slv0_adr[3]), .A3(_u0_u0_n924 ), .ZN(_u0_u0_n792 ) );
NOR2_X2 _u0_u0_U375  ( .A1(_u0_u0_n928 ), .A2(_u0_u0_n930 ), .ZN(_u0_u0_n929 ) );
NOR2_X2 _u0_u0_U374  ( .A1(_u0_u0_n832 ), .A2(_u0_u0_n834 ), .ZN(_u0_u0_n833 ) );
INV_X4 _u0_u0_U373  ( .A(_u0_u0_n1018 ), .ZN(_u0_u0_n928 ) );
INV_X4 _u0_u0_U372  ( .A(_u0_u0_n922 ), .ZN(_u0_u0_n832 ) );
INV_X4 _u0_u0_U371  ( .A(_u0_u0_n770 ), .ZN(_u0_u0_n757 ) );
AND3_X4 _u0_u0_U370  ( .A1(_u0_u0_n771 ), .A2(_u0_u0_n1018 ), .A3(de_adr1_we), .ZN(_u0_u0_n930 ) );
AND3_X4 _u0_u0_U369  ( .A1(_u0_u0_n771 ), .A2(_u0_u0_n922 ), .A3(de_adr0_we),.ZN(_u0_u0_n834 ) );
INV_X4 _u0_u0_U367  ( .A(1'b1), .ZN(_u0_u0_pointer[31] ) );
INV_X4 _u0_u0_U365  ( .A(1'b1), .ZN(_u0_u0_pointer[30] ) );
INV_X4 _u0_u0_U363  ( .A(1'b1), .ZN(_u0_u0_pointer[29] ) );
INV_X4 _u0_u0_U361  ( .A(1'b1), .ZN(_u0_u0_pointer[28] ) );
INV_X4 _u0_u0_U359  ( .A(1'b1), .ZN(_u0_u0_pointer[27] ) );
INV_X4 _u0_u0_U357  ( .A(1'b1), .ZN(_u0_u0_pointer[26] ) );
INV_X4 _u0_u0_U355  ( .A(1'b1), .ZN(_u0_u0_pointer[25] ) );
INV_X4 _u0_u0_U353  ( .A(1'b1), .ZN(_u0_u0_pointer[24] ) );
INV_X4 _u0_u0_U351  ( .A(1'b1), .ZN(_u0_u0_pointer[23] ) );
INV_X4 _u0_u0_U349  ( .A(1'b1), .ZN(_u0_u0_pointer[22] ) );
INV_X4 _u0_u0_U347  ( .A(1'b1), .ZN(_u0_u0_pointer[21] ) );
INV_X4 _u0_u0_U345  ( .A(1'b1), .ZN(_u0_u0_pointer[20] ) );
INV_X4 _u0_u0_U343  ( .A(1'b1), .ZN(_u0_u0_pointer[19] ) );
INV_X4 _u0_u0_U341  ( .A(1'b1), .ZN(_u0_u0_pointer[18] ) );
INV_X4 _u0_u0_U339  ( .A(1'b1), .ZN(_u0_u0_pointer[17] ) );
INV_X4 _u0_u0_U337  ( .A(1'b1), .ZN(_u0_u0_pointer[16] ) );
INV_X4 _u0_u0_U335  ( .A(1'b1), .ZN(_u0_u0_pointer[15] ) );
INV_X4 _u0_u0_U333  ( .A(1'b1), .ZN(_u0_u0_pointer[14] ) );
INV_X4 _u0_u0_U331  ( .A(1'b1), .ZN(_u0_u0_pointer[13] ) );
INV_X4 _u0_u0_U329  ( .A(1'b1), .ZN(_u0_u0_pointer[12] ) );
INV_X4 _u0_u0_U327  ( .A(1'b1), .ZN(_u0_u0_pointer[11] ) );
INV_X4 _u0_u0_U325  ( .A(1'b1), .ZN(_u0_u0_pointer[10] ) );
INV_X4 _u0_u0_U323  ( .A(1'b1), .ZN(_u0_u0_pointer[9] ) );
INV_X4 _u0_u0_U321  ( .A(1'b1), .ZN(_u0_u0_pointer[8] ) );
INV_X4 _u0_u0_U319  ( .A(1'b1), .ZN(_u0_u0_pointer[7] ) );
INV_X4 _u0_u0_U317  ( .A(1'b1), .ZN(_u0_u0_pointer[6] ) );
INV_X4 _u0_u0_U315  ( .A(1'b1), .ZN(_u0_u0_pointer[5] ) );
INV_X4 _u0_u0_U313  ( .A(1'b1), .ZN(_u0_u0_pointer[4] ) );
INV_X4 _u0_u0_U311  ( .A(1'b1), .ZN(_u0_u0_pointer[3] ) );
INV_X4 _u0_u0_U309  ( .A(1'b1), .ZN(_u0_u0_pointer[2] ) );
INV_X4 _u0_u0_U307  ( .A(1'b1), .ZN(_u0_u0_pointer[1] ) );
INV_X4 _u0_u0_U305  ( .A(1'b1), .ZN(_u0_u0_pointer[0] ) );
INV_X4 _u0_u0_U303  ( .A(1'b1), .ZN(_u0_u0_pointer_s[31] ) );
INV_X4 _u0_u0_U301  ( .A(1'b1), .ZN(_u0_u0_pointer_s[30] ) );
INV_X4 _u0_u0_U299  ( .A(1'b1), .ZN(_u0_u0_pointer_s[29] ) );
INV_X4 _u0_u0_U297  ( .A(1'b1), .ZN(_u0_u0_pointer_s[28] ) );
INV_X4 _u0_u0_U295  ( .A(1'b1), .ZN(_u0_u0_pointer_s[27] ) );
INV_X4 _u0_u0_U293  ( .A(1'b1), .ZN(_u0_u0_pointer_s[26] ) );
INV_X4 _u0_u0_U291  ( .A(1'b1), .ZN(_u0_u0_pointer_s[25] ) );
INV_X4 _u0_u0_U289  ( .A(1'b1), .ZN(_u0_u0_pointer_s[24] ) );
INV_X4 _u0_u0_U287  ( .A(1'b1), .ZN(_u0_u0_pointer_s[23] ) );
INV_X4 _u0_u0_U285  ( .A(1'b1), .ZN(_u0_u0_pointer_s[22] ) );
INV_X4 _u0_u0_U283  ( .A(1'b1), .ZN(_u0_u0_pointer_s[21] ) );
INV_X4 _u0_u0_U281  ( .A(1'b1), .ZN(_u0_u0_pointer_s[20] ) );
INV_X4 _u0_u0_U279  ( .A(1'b1), .ZN(_u0_u0_pointer_s[19] ) );
INV_X4 _u0_u0_U277  ( .A(1'b1), .ZN(_u0_u0_pointer_s[18] ) );
INV_X4 _u0_u0_U275  ( .A(1'b1), .ZN(_u0_u0_pointer_s[17] ) );
INV_X4 _u0_u0_U273  ( .A(1'b1), .ZN(_u0_u0_pointer_s[16] ) );
INV_X4 _u0_u0_U271  ( .A(1'b1), .ZN(_u0_u0_pointer_s[15] ) );
INV_X4 _u0_u0_U269  ( .A(1'b1), .ZN(_u0_u0_pointer_s[14] ) );
INV_X4 _u0_u0_U267  ( .A(1'b1), .ZN(_u0_u0_pointer_s[13] ) );
INV_X4 _u0_u0_U265  ( .A(1'b1), .ZN(_u0_u0_pointer_s[12] ) );
INV_X4 _u0_u0_U263  ( .A(1'b1), .ZN(_u0_u0_pointer_s[11] ) );
INV_X4 _u0_u0_U261  ( .A(1'b1), .ZN(_u0_u0_pointer_s[10] ) );
INV_X4 _u0_u0_U259  ( .A(1'b1), .ZN(_u0_u0_pointer_s[9] ) );
INV_X4 _u0_u0_U257  ( .A(1'b1), .ZN(_u0_u0_pointer_s[8] ) );
INV_X4 _u0_u0_U255  ( .A(1'b1), .ZN(_u0_u0_pointer_s[7] ) );
INV_X4 _u0_u0_U253  ( .A(1'b1), .ZN(_u0_u0_pointer_s[6] ) );
INV_X4 _u0_u0_U251  ( .A(1'b1), .ZN(_u0_u0_pointer_s[5] ) );
INV_X4 _u0_u0_U249  ( .A(1'b1), .ZN(_u0_u0_pointer_s[4] ) );
INV_X4 _u0_u0_U247  ( .A(1'b1), .ZN(_u0_u0_pointer_s[3] ) );
INV_X4 _u0_u0_U245  ( .A(1'b1), .ZN(_u0_u0_pointer_s[2] ) );
INV_X4 _u0_u0_U243  ( .A(1'b1), .ZN(_u0_u0_pointer_s[1] ) );
INV_X4 _u0_u0_U241  ( .A(1'b1), .ZN(_u0_u0_pointer_s[0] ) );
INV_X4 _u0_u0_U239  ( .A(1'b1), .ZN(_u0_u0_ch_csr[31] ) );
INV_X4 _u0_u0_U237  ( .A(1'b1), .ZN(_u0_u0_ch_csr[30] ) );
INV_X4 _u0_u0_U235  ( .A(1'b1), .ZN(_u0_u0_ch_csr[29] ) );
INV_X4 _u0_u0_U233  ( .A(1'b1), .ZN(_u0_u0_ch_csr[28] ) );
INV_X4 _u0_u0_U231  ( .A(1'b1), .ZN(_u0_u0_ch_csr[27] ) );
INV_X4 _u0_u0_U229  ( .A(1'b1), .ZN(_u0_u0_ch_csr[26] ) );
INV_X4 _u0_u0_U227  ( .A(1'b1), .ZN(_u0_u0_ch_csr[25] ) );
INV_X4 _u0_u0_U225  ( .A(1'b1), .ZN(_u0_u0_ch_csr[24] ) );
INV_X4 _u0_u0_U223  ( .A(1'b1), .ZN(_u0_u0_ch_csr[23] ) );
INV_X4 _u0_u0_U221  ( .A(1'b1), .ZN(_u0_u0_ch_csr[9] ) );
INV_X4 _u0_u0_U219  ( .A(1'b1), .ZN(_u0_u0_ch_txsz[31] ) );
INV_X4 _u0_u0_U217  ( .A(1'b1), .ZN(_u0_u0_ch_txsz[30] ) );
INV_X4 _u0_u0_U215  ( .A(1'b1), .ZN(_u0_u0_ch_txsz[29] ) );
INV_X4 _u0_u0_U213  ( .A(1'b1), .ZN(_u0_u0_ch_txsz[28] ) );
INV_X4 _u0_u0_U211  ( .A(1'b1), .ZN(_u0_u0_ch_txsz[27] ) );
INV_X4 _u0_u0_U209  ( .A(1'b1), .ZN(_u0_u0_ch_txsz[14] ) );
INV_X4 _u0_u0_U207  ( .A(1'b1), .ZN(_u0_u0_ch_txsz[13] ) );
INV_X4 _u0_u0_U205  ( .A(1'b1), .ZN(_u0_u0_ch_txsz[12] ) );
INV_X4 _u0_u0_U203  ( .A(1'b1), .ZN(_u0_u0_ch_adr0[1] ) );
INV_X4 _u0_u0_U201  ( .A(1'b1), .ZN(_u0_u0_ch_adr0[0] ) );
INV_X4 _u0_u0_U199  ( .A(1'b1), .ZN(_u0_u0_ch_adr1[1] ) );
INV_X4 _u0_u0_U197  ( .A(1'b1), .ZN(_u0_u0_ch_adr1[0] ) );
INV_X4 _u0_u0_U195  ( .A(1'b0), .ZN(_u0_u0_ch_am0[31] ) );
INV_X4 _u0_u0_U193  ( .A(1'b0), .ZN(_u0_u0_ch_am0[30] ) );
INV_X4 _u0_u0_U191  ( .A(1'b0), .ZN(_u0_u0_ch_am0[29] ) );
INV_X4 _u0_u0_U189  ( .A(1'b0), .ZN(_u0_u0_ch_am0[28] ) );
INV_X4 _u0_u0_U187  ( .A(1'b0), .ZN(_u0_u0_ch_am0[27] ) );
INV_X4 _u0_u0_U185  ( .A(1'b0), .ZN(_u0_u0_ch_am0[26] ) );
INV_X4 _u0_u0_U183  ( .A(1'b0), .ZN(_u0_u0_ch_am0[25] ) );
INV_X4 _u0_u0_U181  ( .A(1'b0), .ZN(_u0_u0_ch_am0[24] ) );
INV_X4 _u0_u0_U179  ( .A(1'b0), .ZN(_u0_u0_ch_am0[23] ) );
INV_X4 _u0_u0_U177  ( .A(1'b0), .ZN(_u0_u0_ch_am0[22] ) );
INV_X4 _u0_u0_U175  ( .A(1'b0), .ZN(_u0_u0_ch_am0[21] ) );
INV_X4 _u0_u0_U173  ( .A(1'b0), .ZN(_u0_u0_ch_am0[20] ) );
INV_X4 _u0_u0_U171  ( .A(1'b0), .ZN(_u0_u0_ch_am0[19] ) );
INV_X4 _u0_u0_U169  ( .A(1'b0), .ZN(_u0_u0_ch_am0[18] ) );
INV_X4 _u0_u0_U167  ( .A(1'b0), .ZN(_u0_u0_ch_am0[17] ) );
INV_X4 _u0_u0_U165  ( .A(1'b0), .ZN(_u0_u0_ch_am0[16] ) );
INV_X4 _u0_u0_U163  ( .A(1'b0), .ZN(_u0_u0_ch_am0[15] ) );
INV_X4 _u0_u0_U161  ( .A(1'b0), .ZN(_u0_u0_ch_am0[14] ) );
INV_X4 _u0_u0_U159  ( .A(1'b0), .ZN(_u0_u0_ch_am0[13] ) );
INV_X4 _u0_u0_U157  ( .A(1'b0), .ZN(_u0_u0_ch_am0[12] ) );
INV_X4 _u0_u0_U155  ( .A(1'b0), .ZN(_u0_u0_ch_am0[11] ) );
INV_X4 _u0_u0_U153  ( .A(1'b0), .ZN(_u0_u0_ch_am0[10] ) );
INV_X4 _u0_u0_U151  ( .A(1'b0), .ZN(_u0_u0_ch_am0[9] ) );
INV_X4 _u0_u0_U149  ( .A(1'b0), .ZN(_u0_u0_ch_am0[8] ) );
INV_X4 _u0_u0_U147  ( .A(1'b0), .ZN(_u0_u0_ch_am0[7] ) );
INV_X4 _u0_u0_U145  ( .A(1'b0), .ZN(_u0_u0_ch_am0[6] ) );
INV_X4 _u0_u0_U143  ( .A(1'b0), .ZN(_u0_u0_ch_am0[5] ) );
INV_X4 _u0_u0_U141  ( .A(1'b0), .ZN(_u0_u0_ch_am0[4] ) );
INV_X4 _u0_u0_U139  ( .A(1'b1), .ZN(_u0_u0_ch_am0[3] ) );
INV_X4 _u0_u0_U137  ( .A(1'b1), .ZN(_u0_u0_ch_am0[2] ) );
INV_X4 _u0_u0_U135  ( .A(1'b1), .ZN(_u0_u0_ch_am0[1] ) );
INV_X4 _u0_u0_U133  ( .A(1'b1), .ZN(_u0_u0_ch_am0[0] ) );
INV_X4 _u0_u0_U131  ( .A(1'b0), .ZN(_u0_u0_ch_am1[31] ) );
INV_X4 _u0_u0_U129  ( .A(1'b0), .ZN(_u0_u0_ch_am1[30] ) );
INV_X4 _u0_u0_U127  ( .A(1'b0), .ZN(_u0_u0_ch_am1[29] ) );
INV_X4 _u0_u0_U125  ( .A(1'b0), .ZN(_u0_u0_ch_am1[28] ) );
INV_X4 _u0_u0_U123  ( .A(1'b0), .ZN(_u0_u0_ch_am1[27] ) );
INV_X4 _u0_u0_U121  ( .A(1'b0), .ZN(_u0_u0_ch_am1[26] ) );
INV_X4 _u0_u0_U119  ( .A(1'b0), .ZN(_u0_u0_ch_am1[25] ) );
INV_X4 _u0_u0_U117  ( .A(1'b0), .ZN(_u0_u0_ch_am1[24] ) );
INV_X4 _u0_u0_U115  ( .A(1'b0), .ZN(_u0_u0_ch_am1[23] ) );
INV_X4 _u0_u0_U113  ( .A(1'b0), .ZN(_u0_u0_ch_am1[22] ) );
INV_X4 _u0_u0_U111  ( .A(1'b0), .ZN(_u0_u0_ch_am1[21] ) );
INV_X4 _u0_u0_U109  ( .A(1'b0), .ZN(_u0_u0_ch_am1[20] ) );
INV_X4 _u0_u0_U107  ( .A(1'b0), .ZN(_u0_u0_ch_am1[19] ) );
INV_X4 _u0_u0_U105  ( .A(1'b0), .ZN(_u0_u0_ch_am1[18] ) );
INV_X4 _u0_u0_U103  ( .A(1'b0), .ZN(_u0_u0_ch_am1[17] ) );
INV_X4 _u0_u0_U101  ( .A(1'b0), .ZN(_u0_u0_ch_am1[16] ) );
INV_X4 _u0_u0_U99  ( .A(1'b0), .ZN(_u0_u0_ch_am1[15] ) );
INV_X4 _u0_u0_U97  ( .A(1'b0), .ZN(_u0_u0_ch_am1[14] ) );
INV_X4 _u0_u0_U95  ( .A(1'b0), .ZN(_u0_u0_ch_am1[13] ) );
INV_X4 _u0_u0_U93  ( .A(1'b0), .ZN(_u0_u0_ch_am1[12] ) );
INV_X4 _u0_u0_U91  ( .A(1'b0), .ZN(_u0_u0_ch_am1[11] ) );
INV_X4 _u0_u0_U89  ( .A(1'b0), .ZN(_u0_u0_ch_am1[10] ) );
INV_X4 _u0_u0_U87  ( .A(1'b0), .ZN(_u0_u0_ch_am1[9] ) );
INV_X4 _u0_u0_U85  ( .A(1'b0), .ZN(_u0_u0_ch_am1[8] ) );
INV_X4 _u0_u0_U83  ( .A(1'b0), .ZN(_u0_u0_ch_am1[7] ) );
INV_X4 _u0_u0_U81  ( .A(1'b0), .ZN(_u0_u0_ch_am1[6] ) );
INV_X4 _u0_u0_U79  ( .A(1'b0), .ZN(_u0_u0_ch_am1[5] ) );
INV_X4 _u0_u0_U77  ( .A(1'b0), .ZN(_u0_u0_ch_am1[4] ) );
INV_X4 _u0_u0_U75  ( .A(1'b1), .ZN(_u0_u0_ch_am1[3] ) );
INV_X4 _u0_u0_U73  ( .A(1'b1), .ZN(_u0_u0_ch_am1[2] ) );
INV_X4 _u0_u0_U71  ( .A(1'b1), .ZN(_u0_u0_ch_am1[1] ) );
INV_X4 _u0_u0_U69  ( .A(1'b1), .ZN(_u0_u0_ch_am1[0] ) );
INV_X4 _u0_u0_U67  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[31] ) );
INV_X4 _u0_u0_U65  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[30] ) );
INV_X4 _u0_u0_U63  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[29] ) );
INV_X4 _u0_u0_U61  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[28] ) );
INV_X4 _u0_u0_U59  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[27] ) );
INV_X4 _u0_u0_U57  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[26] ) );
INV_X4 _u0_u0_U55  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[25] ) );
INV_X4 _u0_u0_U53  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[24] ) );
INV_X4 _u0_u0_U51  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[23] ) );
INV_X4 _u0_u0_U49  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[22] ) );
INV_X4 _u0_u0_U47  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[21] ) );
INV_X4 _u0_u0_U45  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[20] ) );
INV_X4 _u0_u0_U43  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[19] ) );
INV_X4 _u0_u0_U41  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[18] ) );
INV_X4 _u0_u0_U39  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[17] ) );
INV_X4 _u0_u0_U37  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[16] ) );
INV_X4 _u0_u0_U35  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[15] ) );
INV_X4 _u0_u0_U33  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[14] ) );
INV_X4 _u0_u0_U31  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[13] ) );
INV_X4 _u0_u0_U29  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[12] ) );
INV_X4 _u0_u0_U27  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[11] ) );
INV_X4 _u0_u0_U25  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[10] ) );
INV_X4 _u0_u0_U23  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[9] ) );
INV_X4 _u0_u0_U21  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[8] ) );
INV_X4 _u0_u0_U19  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[7] ) );
INV_X4 _u0_u0_U17  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[6] ) );
INV_X4 _u0_u0_U15  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[5] ) );
INV_X4 _u0_u0_U13  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[4] ) );
INV_X4 _u0_u0_U11  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[3] ) );
INV_X4 _u0_u0_U9  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[2] ) );
INV_X4 _u0_u0_U7  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[1] ) );
INV_X4 _u0_u0_U5  ( .A(1'b1), .ZN(_u0_u0_sw_pointer[0] ) );
INV_X4 _u0_u0_U3  ( .A(1'b1), .ZN(_u0_u0_ch_dis ) );
DFF_X2 _u0_u0_ch_adr1_r_reg_0_  ( .D(_u0_u0_n347 ), .CK(clk_i), .Q(ch0_adr1[2]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_1_  ( .D(_u0_u0_n348 ), .CK(clk_i), .Q(ch0_adr1[3]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_2_  ( .D(_u0_u0_n349 ), .CK(clk_i), .Q(ch0_adr1[4]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_3_  ( .D(_u0_u0_n350 ), .CK(clk_i), .Q(ch0_adr1[5]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_4_  ( .D(_u0_u0_n351 ), .CK(clk_i), .Q(ch0_adr1[6]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_5_  ( .D(_u0_u0_n352 ), .CK(clk_i), .Q(ch0_adr1[7]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_6_  ( .D(_u0_u0_n353 ), .CK(clk_i), .Q(ch0_adr1[8]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_7_  ( .D(_u0_u0_n354 ), .CK(clk_i), .Q(ch0_adr1[9]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_8_  ( .D(_u0_u0_n355 ), .CK(clk_i), .Q(ch0_adr1[10]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_9_  ( .D(_u0_u0_n356 ), .CK(clk_i), .Q(ch0_adr1[11]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_10_  ( .D(_u0_u0_n357 ), .CK(clk_i), .Q(ch0_adr1[12]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_11_  ( .D(_u0_u0_n358 ), .CK(clk_i), .Q(ch0_adr1[13]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_12_  ( .D(_u0_u0_n359 ), .CK(clk_i), .Q(ch0_adr1[14]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_13_  ( .D(_u0_u0_n360 ), .CK(clk_i), .Q(ch0_adr1[15]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_14_  ( .D(_u0_u0_n361 ), .CK(clk_i), .Q(ch0_adr1[16]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_15_  ( .D(_u0_u0_n362 ), .CK(clk_i), .Q(ch0_adr1[17]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_16_  ( .D(_u0_u0_n363 ), .CK(clk_i), .Q(ch0_adr1[18]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_17_  ( .D(_u0_u0_n364 ), .CK(clk_i), .Q(ch0_adr1[19]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_18_  ( .D(_u0_u0_n365 ), .CK(clk_i), .Q(ch0_adr1[20]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_19_  ( .D(_u0_u0_n366 ), .CK(clk_i), .Q(ch0_adr1[21]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_20_  ( .D(_u0_u0_n367 ), .CK(clk_i), .Q(ch0_adr1[22]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_21_  ( .D(_u0_u0_n368 ), .CK(clk_i), .Q(ch0_adr1[23]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_22_  ( .D(_u0_u0_n369 ), .CK(clk_i), .Q(ch0_adr1[24]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_23_  ( .D(_u0_u0_n370 ), .CK(clk_i), .Q(ch0_adr1[25]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_24_  ( .D(_u0_u0_n371 ), .CK(clk_i), .Q(ch0_adr1[26]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_25_  ( .D(_u0_u0_n372 ), .CK(clk_i), .Q(ch0_adr1[27]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_26_  ( .D(_u0_u0_n373 ), .CK(clk_i), .Q(ch0_adr1[28]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_27_  ( .D(_u0_u0_n374 ), .CK(clk_i), .Q(ch0_adr1[29]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_28_  ( .D(_u0_u0_n375 ), .CK(clk_i), .Q(ch0_adr1[30]), .QN() );
DFF_X2 _u0_u0_ch_adr1_r_reg_29_  ( .D(_u0_u0_n376 ), .CK(clk_i), .Q(ch0_adr1[31]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_0_  ( .D(_u0_u0_n377 ), .CK(clk_i), .Q(ch0_adr0[2]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_1_  ( .D(_u0_u0_n378 ), .CK(clk_i), .Q(ch0_adr0[3]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_2_  ( .D(_u0_u0_n379 ), .CK(clk_i), .Q(ch0_adr0[4]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_3_  ( .D(_u0_u0_n380 ), .CK(clk_i), .Q(ch0_adr0[5]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_4_  ( .D(_u0_u0_n381 ), .CK(clk_i), .Q(ch0_adr0[6]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_5_  ( .D(_u0_u0_n382 ), .CK(clk_i), .Q(ch0_adr0[7]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_6_  ( .D(_u0_u0_n383 ), .CK(clk_i), .Q(ch0_adr0[8]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_7_  ( .D(_u0_u0_n384 ), .CK(clk_i), .Q(ch0_adr0[9]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_8_  ( .D(_u0_u0_n385 ), .CK(clk_i), .Q(ch0_adr0[10]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_9_  ( .D(_u0_u0_n386 ), .CK(clk_i), .Q(ch0_adr0[11]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_10_  ( .D(_u0_u0_n387 ), .CK(clk_i), .Q(ch0_adr0[12]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_11_  ( .D(_u0_u0_n388 ), .CK(clk_i), .Q(ch0_adr0[13]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_12_  ( .D(_u0_u0_n389 ), .CK(clk_i), .Q(ch0_adr0[14]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_13_  ( .D(_u0_u0_n390 ), .CK(clk_i), .Q(ch0_adr0[15]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_14_  ( .D(_u0_u0_n391 ), .CK(clk_i), .Q(ch0_adr0[16]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_15_  ( .D(_u0_u0_n392 ), .CK(clk_i), .Q(ch0_adr0[17]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_16_  ( .D(_u0_u0_n393 ), .CK(clk_i), .Q(ch0_adr0[18]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_17_  ( .D(_u0_u0_n394 ), .CK(clk_i), .Q(ch0_adr0[19]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_18_  ( .D(_u0_u0_n395 ), .CK(clk_i), .Q(ch0_adr0[20]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_19_  ( .D(_u0_u0_n396 ), .CK(clk_i), .Q(ch0_adr0[21]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_20_  ( .D(_u0_u0_n397 ), .CK(clk_i), .Q(ch0_adr0[22]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_21_  ( .D(_u0_u0_n398 ), .CK(clk_i), .Q(ch0_adr0[23]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_22_  ( .D(_u0_u0_n399 ), .CK(clk_i), .Q(ch0_adr0[24]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_23_  ( .D(_u0_u0_n400 ), .CK(clk_i), .Q(ch0_adr0[25]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_24_  ( .D(_u0_u0_n401 ), .CK(clk_i), .Q(ch0_adr0[26]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_25_  ( .D(_u0_u0_n402 ), .CK(clk_i), .Q(ch0_adr0[27]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_26_  ( .D(_u0_u0_n403 ), .CK(clk_i), .Q(ch0_adr0[28]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_27_  ( .D(_u0_u0_n404 ), .CK(clk_i), .Q(ch0_adr0[29]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_28_  ( .D(_u0_u0_n405 ), .CK(clk_i), .Q(ch0_adr0[30]), .QN() );
DFF_X2 _u0_u0_ch_adr0_r_reg_29_  ( .D(_u0_u0_n406 ), .CK(clk_i), .Q(ch0_adr0[31]), .QN() );
DFF_X2 _u0_u0_ch_sz_inf_reg  ( .D(_u0_u0_n335 ), .CK(clk_i), .Q(ch0_txsz[15]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_0_  ( .D(_u0_u0_n407 ), .CK(clk_i), .Q(ch0_txsz[16]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_1_  ( .D(_u0_u0_n408 ), .CK(clk_i), .Q(ch0_txsz[17]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_2_  ( .D(_u0_u0_n409 ), .CK(clk_i), .Q(ch0_txsz[18]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_3_  ( .D(_u0_u0_n410 ), .CK(clk_i), .Q(ch0_txsz[19]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_4_  ( .D(_u0_u0_n411 ), .CK(clk_i), .Q(ch0_txsz[20]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_5_  ( .D(_u0_u0_n412 ), .CK(clk_i), .Q(ch0_txsz[21]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_6_  ( .D(_u0_u0_n413 ), .CK(clk_i), .Q(ch0_txsz[22]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_7_  ( .D(_u0_u0_n414 ), .CK(clk_i), .Q(ch0_txsz[23]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_8_  ( .D(_u0_u0_n415 ), .CK(clk_i), .Q(ch0_txsz[24]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_9_  ( .D(_u0_u0_n416 ), .CK(clk_i), .Q(ch0_txsz[25]), .QN() );
DFF_X2 _u0_u0_ch_chk_sz_r_reg_10_  ( .D(_u0_u0_n417 ), .CK(clk_i), .Q(ch0_txsz[26]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_0_  ( .D(_u0_u0_n418 ), .CK(clk_i), .Q(ch0_txsz[0]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_1_  ( .D(_u0_u0_n419 ), .CK(clk_i), .Q(ch0_txsz[1]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_2_  ( .D(_u0_u0_n420 ), .CK(clk_i), .Q(ch0_txsz[2]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_3_  ( .D(_u0_u0_n421 ), .CK(clk_i), .Q(ch0_txsz[3]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_4_  ( .D(_u0_u0_n422 ), .CK(clk_i), .Q(ch0_txsz[4]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_5_  ( .D(_u0_u0_n423 ), .CK(clk_i), .Q(ch0_txsz[5]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_6_  ( .D(_u0_u0_n424 ), .CK(clk_i), .Q(ch0_txsz[6]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_7_  ( .D(_u0_u0_n425 ), .CK(clk_i), .Q(ch0_txsz[7]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_8_  ( .D(_u0_u0_n426 ), .CK(clk_i), .Q(ch0_txsz[8]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_9_  ( .D(_u0_u0_n427 ), .CK(clk_i), .Q(ch0_txsz[9]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_10_  ( .D(_u0_u0_n428 ), .CK(clk_i), .Q(ch0_txsz[10]), .QN() );
DFF_X2 _u0_u0_ch_tot_sz_r_reg_11_  ( .D(_u0_u0_n429 ), .CK(clk_i), .Q(ch0_txsz[11]), .QN() );
DFF_X2 _u0_u0_ch_stop_reg  ( .D(_u0_u0_N24 ), .CK(clk_i), .Q(dma_abort),.QN() );
DFF_X2 _u0_u0_ch_busy_reg  ( .D(_u0_u0_N23 ), .CK(clk_i), .Q(ch0_csr[10]),.QN() );
DFFR_X1 _u0_u0_int_src_r_reg_0_  ( .D(_u0_u0_n430 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[20]), .QN() );
DFFR_X1 _u0_u0_int_src_r_reg_1_  ( .D(_u0_u0_n431 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[21]), .QN() );
DFFR_X1 _u0_u0_int_src_r_reg_2_  ( .D(_u0_u0_n432 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[22]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r3_reg_0_  ( .D(_u0_u0_n336 ), .CK(clk_i), .RN(_u0_u0_n752 ), .Q(ch0_csr[17]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r3_reg_1_  ( .D(_u0_u0_n337 ), .CK(clk_i), .RN(_u0_u0_n752 ), .Q(ch0_csr[18]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r3_reg_2_  ( .D(_u0_u0_n338 ), .CK(clk_i), .RN(_u0_u0_n752 ), .Q(ch0_csr[19]), .QN() );
DFFR_X1 _u0_u0_rest_en_reg  ( .D(_u0_u0_n339 ), .CK(clk_i), .RN(_u0_u0_n752 ), .Q(ch0_csr[16]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r2_reg_0_  ( .D(_u0_u0_n340 ), .CK(clk_i), .RN(_u0_u0_n752 ), .Q(ch0_csr[13]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r2_reg_1_  ( .D(_u0_u0_n341 ), .CK(clk_i), .RN(_u0_u0_n752 ), .Q(ch0_csr[14]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r2_reg_2_  ( .D(_u0_u0_n342 ), .CK(clk_i), .RN(_u0_u0_n752 ), .Q(ch0_csr[15]), .QN() );
DFFR_X1 _u0_u0_ch_err_reg  ( .D(_u0_u0_n433 ), .CK(clk_i), .RN(_u0_u0_n751 ),.Q(ch0_csr[12]), .QN() );
DFFR_X1 _u0_u0_ch_done_reg  ( .D(_u0_u0_n434 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[11]), .QN(_u0_u0_n326 ) );
DFFR_X1 _u0_u0_ch_csr_r_reg_0_  ( .D(_u0_u0_n435 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[0]), .QN(_u0_u0_n1026 ) );
DFFR_X1 _u0_u0_ch_csr_r_reg_1_  ( .D(_u0_u0_n436 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[1]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r_reg_2_  ( .D(_u0_u0_n437 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[2]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r_reg_3_  ( .D(_u0_u0_n438 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[3]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r_reg_4_  ( .D(_u0_u0_n439 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[4]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r_reg_5_  ( .D(_u0_u0_n343 ), .CK(clk_i), .RN(_u0_u0_n752 ), .Q(ch0_csr[5]), .QN() );
DFFR_X1 _u0_u0_ch_csr_r_reg_6_  ( .D(_u0_u0_n344 ), .CK(clk_i), .RN(_u0_u0_n752 ), .Q(ch0_csr[6]), .QN(_u0_u0_n333 ) );
DFFR_X1 _u0_u0_ch_csr_r_reg_7_  ( .D(_u0_u0_n345 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[7]), .QN(_u0_u0_n334 ) );
DFFR_X1 _u0_u0_ch_csr_r_reg_8_  ( .D(_u0_u0_n346 ), .CK(clk_i), .RN(_u0_u0_n751 ), .Q(ch0_csr[8]), .QN() );
INV_X4 _u0_u1_U585  ( .A(1'b1), .ZN(_u0_u1_pointer[31] ) );
INV_X4 _u0_u1_U583  ( .A(1'b1), .ZN(_u0_u1_pointer[30] ) );
INV_X4 _u0_u1_U581  ( .A(1'b1), .ZN(_u0_u1_pointer[29] ) );
INV_X4 _u0_u1_U579  ( .A(1'b1), .ZN(_u0_u1_pointer[28] ) );
INV_X4 _u0_u1_U577  ( .A(1'b1), .ZN(_u0_u1_pointer[27] ) );
INV_X4 _u0_u1_U575  ( .A(1'b1), .ZN(_u0_u1_pointer[26] ) );
INV_X4 _u0_u1_U573  ( .A(1'b1), .ZN(_u0_u1_pointer[25] ) );
INV_X4 _u0_u1_U571  ( .A(1'b1), .ZN(_u0_u1_pointer[24] ) );
INV_X4 _u0_u1_U569  ( .A(1'b1), .ZN(_u0_u1_pointer[23] ) );
INV_X4 _u0_u1_U567  ( .A(1'b1), .ZN(_u0_u1_pointer[22] ) );
INV_X4 _u0_u1_U565  ( .A(1'b1), .ZN(_u0_u1_pointer[21] ) );
INV_X4 _u0_u1_U563  ( .A(1'b1), .ZN(_u0_u1_pointer[20] ) );
INV_X4 _u0_u1_U561  ( .A(1'b1), .ZN(_u0_u1_pointer[19] ) );
INV_X4 _u0_u1_U559  ( .A(1'b1), .ZN(_u0_u1_pointer[18] ) );
INV_X4 _u0_u1_U557  ( .A(1'b1), .ZN(_u0_u1_pointer[17] ) );
INV_X4 _u0_u1_U555  ( .A(1'b1), .ZN(_u0_u1_pointer[16] ) );
INV_X4 _u0_u1_U553  ( .A(1'b1), .ZN(_u0_u1_pointer[15] ) );
INV_X4 _u0_u1_U551  ( .A(1'b1), .ZN(_u0_u1_pointer[14] ) );
INV_X4 _u0_u1_U549  ( .A(1'b1), .ZN(_u0_u1_pointer[13] ) );
INV_X4 _u0_u1_U547  ( .A(1'b1), .ZN(_u0_u1_pointer[12] ) );
INV_X4 _u0_u1_U545  ( .A(1'b1), .ZN(_u0_u1_pointer[11] ) );
INV_X4 _u0_u1_U543  ( .A(1'b1), .ZN(_u0_u1_pointer[10] ) );
INV_X4 _u0_u1_U541  ( .A(1'b1), .ZN(_u0_u1_pointer[9] ) );
INV_X4 _u0_u1_U539  ( .A(1'b1), .ZN(_u0_u1_pointer[8] ) );
INV_X4 _u0_u1_U537  ( .A(1'b1), .ZN(_u0_u1_pointer[7] ) );
INV_X4 _u0_u1_U535  ( .A(1'b1), .ZN(_u0_u1_pointer[6] ) );
INV_X4 _u0_u1_U533  ( .A(1'b1), .ZN(_u0_u1_pointer[5] ) );
INV_X4 _u0_u1_U531  ( .A(1'b1), .ZN(_u0_u1_pointer[4] ) );
INV_X4 _u0_u1_U529  ( .A(1'b1), .ZN(_u0_u1_pointer[3] ) );
INV_X4 _u0_u1_U527  ( .A(1'b1), .ZN(_u0_u1_pointer[2] ) );
INV_X4 _u0_u1_U525  ( .A(1'b1), .ZN(_u0_u1_pointer[1] ) );
INV_X4 _u0_u1_U523  ( .A(1'b1), .ZN(_u0_u1_pointer[0] ) );
INV_X4 _u0_u1_U521  ( .A(1'b1), .ZN(_u0_u1_pointer_s[31] ) );
INV_X4 _u0_u1_U519  ( .A(1'b1), .ZN(_u0_u1_pointer_s[30] ) );
INV_X4 _u0_u1_U517  ( .A(1'b1), .ZN(_u0_u1_pointer_s[29] ) );
INV_X4 _u0_u1_U515  ( .A(1'b1), .ZN(_u0_u1_pointer_s[28] ) );
INV_X4 _u0_u1_U513  ( .A(1'b1), .ZN(_u0_u1_pointer_s[27] ) );
INV_X4 _u0_u1_U511  ( .A(1'b1), .ZN(_u0_u1_pointer_s[26] ) );
INV_X4 _u0_u1_U509  ( .A(1'b1), .ZN(_u0_u1_pointer_s[25] ) );
INV_X4 _u0_u1_U507  ( .A(1'b1), .ZN(_u0_u1_pointer_s[24] ) );
INV_X4 _u0_u1_U505  ( .A(1'b1), .ZN(_u0_u1_pointer_s[23] ) );
INV_X4 _u0_u1_U503  ( .A(1'b1), .ZN(_u0_u1_pointer_s[22] ) );
INV_X4 _u0_u1_U501  ( .A(1'b1), .ZN(_u0_u1_pointer_s[21] ) );
INV_X4 _u0_u1_U499  ( .A(1'b1), .ZN(_u0_u1_pointer_s[20] ) );
INV_X4 _u0_u1_U497  ( .A(1'b1), .ZN(_u0_u1_pointer_s[19] ) );
INV_X4 _u0_u1_U495  ( .A(1'b1), .ZN(_u0_u1_pointer_s[18] ) );
INV_X4 _u0_u1_U493  ( .A(1'b1), .ZN(_u0_u1_pointer_s[17] ) );
INV_X4 _u0_u1_U491  ( .A(1'b1), .ZN(_u0_u1_pointer_s[16] ) );
INV_X4 _u0_u1_U489  ( .A(1'b1), .ZN(_u0_u1_pointer_s[15] ) );
INV_X4 _u0_u1_U487  ( .A(1'b1), .ZN(_u0_u1_pointer_s[14] ) );
INV_X4 _u0_u1_U485  ( .A(1'b1), .ZN(_u0_u1_pointer_s[13] ) );
INV_X4 _u0_u1_U483  ( .A(1'b1), .ZN(_u0_u1_pointer_s[12] ) );
INV_X4 _u0_u1_U481  ( .A(1'b1), .ZN(_u0_u1_pointer_s[11] ) );
INV_X4 _u0_u1_U479  ( .A(1'b1), .ZN(_u0_u1_pointer_s[10] ) );
INV_X4 _u0_u1_U477  ( .A(1'b1), .ZN(_u0_u1_pointer_s[9] ) );
INV_X4 _u0_u1_U475  ( .A(1'b1), .ZN(_u0_u1_pointer_s[8] ) );
INV_X4 _u0_u1_U473  ( .A(1'b1), .ZN(_u0_u1_pointer_s[7] ) );
INV_X4 _u0_u1_U471  ( .A(1'b1), .ZN(_u0_u1_pointer_s[6] ) );
INV_X4 _u0_u1_U469  ( .A(1'b1), .ZN(_u0_u1_pointer_s[5] ) );
INV_X4 _u0_u1_U467  ( .A(1'b1), .ZN(_u0_u1_pointer_s[4] ) );
INV_X4 _u0_u1_U465  ( .A(1'b1), .ZN(_u0_u1_pointer_s[3] ) );
INV_X4 _u0_u1_U463  ( .A(1'b1), .ZN(_u0_u1_pointer_s[2] ) );
INV_X4 _u0_u1_U461  ( .A(1'b1), .ZN(_u0_u1_pointer_s[1] ) );
INV_X4 _u0_u1_U459  ( .A(1'b1), .ZN(_u0_u1_pointer_s[0] ) );
INV_X4 _u0_u1_U457  ( .A(1'b1), .ZN(_u0_u1_ch_csr[31] ) );
INV_X4 _u0_u1_U455  ( .A(1'b1), .ZN(_u0_u1_ch_csr[30] ) );
INV_X4 _u0_u1_U453  ( .A(1'b1), .ZN(_u0_u1_ch_csr[29] ) );
INV_X4 _u0_u1_U451  ( .A(1'b1), .ZN(_u0_u1_ch_csr[28] ) );
INV_X4 _u0_u1_U449  ( .A(1'b1), .ZN(_u0_u1_ch_csr[27] ) );
INV_X4 _u0_u1_U447  ( .A(1'b1), .ZN(_u0_u1_ch_csr[26] ) );
INV_X4 _u0_u1_U445  ( .A(1'b1), .ZN(_u0_u1_ch_csr[25] ) );
INV_X4 _u0_u1_U443  ( .A(1'b1), .ZN(_u0_u1_ch_csr[24] ) );
INV_X4 _u0_u1_U441  ( .A(1'b1), .ZN(_u0_u1_ch_csr[23] ) );
INV_X4 _u0_u1_U439  ( .A(1'b1), .ZN(_u0_u1_ch_csr[22] ) );
INV_X4 _u0_u1_U437  ( .A(1'b1), .ZN(_u0_u1_ch_csr[21] ) );
INV_X4 _u0_u1_U435  ( .A(1'b1), .ZN(_u0_u1_ch_csr[20] ) );
INV_X4 _u0_u1_U433  ( .A(1'b1), .ZN(_u0_u1_ch_csr[19] ) );
INV_X4 _u0_u1_U431  ( .A(1'b1), .ZN(_u0_u1_ch_csr[18] ) );
INV_X4 _u0_u1_U429  ( .A(1'b1), .ZN(_u0_u1_ch_csr[17] ) );
INV_X4 _u0_u1_U427  ( .A(1'b1), .ZN(_u0_u1_ch_csr[16] ) );
INV_X4 _u0_u1_U425  ( .A(1'b1), .ZN(_u0_u1_ch_csr[15] ) );
INV_X4 _u0_u1_U423  ( .A(1'b1), .ZN(_u0_u1_ch_csr[14] ) );
INV_X4 _u0_u1_U421  ( .A(1'b1), .ZN(_u0_u1_ch_csr[13] ) );
INV_X4 _u0_u1_U419  ( .A(1'b1), .ZN(_u0_u1_ch_csr[12] ) );
INV_X4 _u0_u1_U417  ( .A(1'b1), .ZN(_u0_u1_ch_csr[11] ) );
INV_X4 _u0_u1_U415  ( .A(1'b1), .ZN(_u0_u1_ch_csr[10] ) );
INV_X4 _u0_u1_U413  ( .A(1'b1), .ZN(_u0_u1_ch_csr[9] ) );
INV_X4 _u0_u1_U411  ( .A(1'b1), .ZN(_u0_u1_ch_csr[8] ) );
INV_X4 _u0_u1_U409  ( .A(1'b1), .ZN(_u0_u1_ch_csr[7] ) );
INV_X4 _u0_u1_U407  ( .A(1'b1), .ZN(_u0_u1_ch_csr[6] ) );
INV_X4 _u0_u1_U405  ( .A(1'b1), .ZN(_u0_u1_ch_csr[5] ) );
INV_X4 _u0_u1_U403  ( .A(1'b1), .ZN(_u0_u1_ch_csr[4] ) );
INV_X4 _u0_u1_U401  ( .A(1'b1), .ZN(_u0_u1_ch_csr[3] ) );
INV_X4 _u0_u1_U399  ( .A(1'b1), .ZN(_u0_u1_ch_csr[2] ) );
INV_X4 _u0_u1_U397  ( .A(1'b1), .ZN(_u0_u1_ch_csr[1] ) );
INV_X4 _u0_u1_U395  ( .A(1'b1), .ZN(_u0_u1_ch_csr[0] ) );
INV_X4 _u0_u1_U393  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[31] ) );
INV_X4 _u0_u1_U391  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[30] ) );
INV_X4 _u0_u1_U389  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[29] ) );
INV_X4 _u0_u1_U387  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[28] ) );
INV_X4 _u0_u1_U385  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[27] ) );
INV_X4 _u0_u1_U383  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[26] ) );
INV_X4 _u0_u1_U381  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[25] ) );
INV_X4 _u0_u1_U379  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[24] ) );
INV_X4 _u0_u1_U377  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[23] ) );
INV_X4 _u0_u1_U375  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[22] ) );
INV_X4 _u0_u1_U373  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[21] ) );
INV_X4 _u0_u1_U371  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[20] ) );
INV_X4 _u0_u1_U369  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[19] ) );
INV_X4 _u0_u1_U367  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[18] ) );
INV_X4 _u0_u1_U365  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[17] ) );
INV_X4 _u0_u1_U363  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[16] ) );
INV_X4 _u0_u1_U361  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[15] ) );
INV_X4 _u0_u1_U359  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[14] ) );
INV_X4 _u0_u1_U357  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[13] ) );
INV_X4 _u0_u1_U355  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[12] ) );
INV_X4 _u0_u1_U353  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[11] ) );
INV_X4 _u0_u1_U351  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[10] ) );
INV_X4 _u0_u1_U349  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[9] ) );
INV_X4 _u0_u1_U347  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[8] ) );
INV_X4 _u0_u1_U345  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[7] ) );
INV_X4 _u0_u1_U343  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[6] ) );
INV_X4 _u0_u1_U341  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[5] ) );
INV_X4 _u0_u1_U339  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[4] ) );
INV_X4 _u0_u1_U337  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[3] ) );
INV_X4 _u0_u1_U335  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[2] ) );
INV_X4 _u0_u1_U333  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[1] ) );
INV_X4 _u0_u1_U331  ( .A(1'b1), .ZN(_u0_u1_ch_txsz[0] ) );
INV_X4 _u0_u1_U329  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[31] ) );
INV_X4 _u0_u1_U327  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[30] ) );
INV_X4 _u0_u1_U325  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[29] ) );
INV_X4 _u0_u1_U323  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[28] ) );
INV_X4 _u0_u1_U321  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[27] ) );
INV_X4 _u0_u1_U319  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[26] ) );
INV_X4 _u0_u1_U317  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[25] ) );
INV_X4 _u0_u1_U315  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[24] ) );
INV_X4 _u0_u1_U313  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[23] ) );
INV_X4 _u0_u1_U311  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[22] ) );
INV_X4 _u0_u1_U309  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[21] ) );
INV_X4 _u0_u1_U307  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[20] ) );
INV_X4 _u0_u1_U305  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[19] ) );
INV_X4 _u0_u1_U303  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[18] ) );
INV_X4 _u0_u1_U301  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[17] ) );
INV_X4 _u0_u1_U299  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[16] ) );
INV_X4 _u0_u1_U297  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[15] ) );
INV_X4 _u0_u1_U295  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[14] ) );
INV_X4 _u0_u1_U293  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[13] ) );
INV_X4 _u0_u1_U291  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[12] ) );
INV_X4 _u0_u1_U289  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[11] ) );
INV_X4 _u0_u1_U287  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[10] ) );
INV_X4 _u0_u1_U285  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[9] ) );
INV_X4 _u0_u1_U283  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[8] ) );
INV_X4 _u0_u1_U281  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[7] ) );
INV_X4 _u0_u1_U279  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[6] ) );
INV_X4 _u0_u1_U277  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[5] ) );
INV_X4 _u0_u1_U275  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[4] ) );
INV_X4 _u0_u1_U273  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[3] ) );
INV_X4 _u0_u1_U271  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[2] ) );
INV_X4 _u0_u1_U269  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[1] ) );
INV_X4 _u0_u1_U267  ( .A(1'b1), .ZN(_u0_u1_ch_adr0[0] ) );
INV_X4 _u0_u1_U265  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[31] ) );
INV_X4 _u0_u1_U263  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[30] ) );
INV_X4 _u0_u1_U261  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[29] ) );
INV_X4 _u0_u1_U259  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[28] ) );
INV_X4 _u0_u1_U257  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[27] ) );
INV_X4 _u0_u1_U255  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[26] ) );
INV_X4 _u0_u1_U253  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[25] ) );
INV_X4 _u0_u1_U251  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[24] ) );
INV_X4 _u0_u1_U249  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[23] ) );
INV_X4 _u0_u1_U247  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[22] ) );
INV_X4 _u0_u1_U245  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[21] ) );
INV_X4 _u0_u1_U243  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[20] ) );
INV_X4 _u0_u1_U241  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[19] ) );
INV_X4 _u0_u1_U239  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[18] ) );
INV_X4 _u0_u1_U237  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[17] ) );
INV_X4 _u0_u1_U235  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[16] ) );
INV_X4 _u0_u1_U233  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[15] ) );
INV_X4 _u0_u1_U231  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[14] ) );
INV_X4 _u0_u1_U229  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[13] ) );
INV_X4 _u0_u1_U227  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[12] ) );
INV_X4 _u0_u1_U225  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[11] ) );
INV_X4 _u0_u1_U223  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[10] ) );
INV_X4 _u0_u1_U221  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[9] ) );
INV_X4 _u0_u1_U219  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[8] ) );
INV_X4 _u0_u1_U217  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[7] ) );
INV_X4 _u0_u1_U215  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[6] ) );
INV_X4 _u0_u1_U213  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[5] ) );
INV_X4 _u0_u1_U211  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[4] ) );
INV_X4 _u0_u1_U209  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[3] ) );
INV_X4 _u0_u1_U207  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[2] ) );
INV_X4 _u0_u1_U205  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[1] ) );
INV_X4 _u0_u1_U203  ( .A(1'b1), .ZN(_u0_u1_ch_adr1[0] ) );
INV_X4 _u0_u1_U201  ( .A(1'b0), .ZN(_u0_u1_ch_am0[31] ) );
INV_X4 _u0_u1_U199  ( .A(1'b0), .ZN(_u0_u1_ch_am0[30] ) );
INV_X4 _u0_u1_U197  ( .A(1'b0), .ZN(_u0_u1_ch_am0[29] ) );
INV_X4 _u0_u1_U195  ( .A(1'b0), .ZN(_u0_u1_ch_am0[28] ) );
INV_X4 _u0_u1_U193  ( .A(1'b0), .ZN(_u0_u1_ch_am0[27] ) );
INV_X4 _u0_u1_U191  ( .A(1'b0), .ZN(_u0_u1_ch_am0[26] ) );
INV_X4 _u0_u1_U189  ( .A(1'b0), .ZN(_u0_u1_ch_am0[25] ) );
INV_X4 _u0_u1_U187  ( .A(1'b0), .ZN(_u0_u1_ch_am0[24] ) );
INV_X4 _u0_u1_U185  ( .A(1'b0), .ZN(_u0_u1_ch_am0[23] ) );
INV_X4 _u0_u1_U183  ( .A(1'b0), .ZN(_u0_u1_ch_am0[22] ) );
INV_X4 _u0_u1_U181  ( .A(1'b0), .ZN(_u0_u1_ch_am0[21] ) );
INV_X4 _u0_u1_U179  ( .A(1'b0), .ZN(_u0_u1_ch_am0[20] ) );
INV_X4 _u0_u1_U177  ( .A(1'b0), .ZN(_u0_u1_ch_am0[19] ) );
INV_X4 _u0_u1_U175  ( .A(1'b0), .ZN(_u0_u1_ch_am0[18] ) );
INV_X4 _u0_u1_U173  ( .A(1'b0), .ZN(_u0_u1_ch_am0[17] ) );
INV_X4 _u0_u1_U171  ( .A(1'b0), .ZN(_u0_u1_ch_am0[16] ) );
INV_X4 _u0_u1_U169  ( .A(1'b0), .ZN(_u0_u1_ch_am0[15] ) );
INV_X4 _u0_u1_U167  ( .A(1'b0), .ZN(_u0_u1_ch_am0[14] ) );
INV_X4 _u0_u1_U165  ( .A(1'b0), .ZN(_u0_u1_ch_am0[13] ) );
INV_X4 _u0_u1_U163  ( .A(1'b0), .ZN(_u0_u1_ch_am0[12] ) );
INV_X4 _u0_u1_U161  ( .A(1'b0), .ZN(_u0_u1_ch_am0[11] ) );
INV_X4 _u0_u1_U159  ( .A(1'b0), .ZN(_u0_u1_ch_am0[10] ) );
INV_X4 _u0_u1_U157  ( .A(1'b0), .ZN(_u0_u1_ch_am0[9] ) );
INV_X4 _u0_u1_U155  ( .A(1'b0), .ZN(_u0_u1_ch_am0[8] ) );
INV_X4 _u0_u1_U153  ( .A(1'b0), .ZN(_u0_u1_ch_am0[7] ) );
INV_X4 _u0_u1_U151  ( .A(1'b0), .ZN(_u0_u1_ch_am0[6] ) );
INV_X4 _u0_u1_U149  ( .A(1'b0), .ZN(_u0_u1_ch_am0[5] ) );
INV_X4 _u0_u1_U147  ( .A(1'b0), .ZN(_u0_u1_ch_am0[4] ) );
INV_X4 _u0_u1_U145  ( .A(1'b1), .ZN(_u0_u1_ch_am0[3] ) );
INV_X4 _u0_u1_U143  ( .A(1'b1), .ZN(_u0_u1_ch_am0[2] ) );
INV_X4 _u0_u1_U141  ( .A(1'b1), .ZN(_u0_u1_ch_am0[1] ) );
INV_X4 _u0_u1_U139  ( .A(1'b1), .ZN(_u0_u1_ch_am0[0] ) );
INV_X4 _u0_u1_U137  ( .A(1'b0), .ZN(_u0_u1_ch_am1[31] ) );
INV_X4 _u0_u1_U135  ( .A(1'b0), .ZN(_u0_u1_ch_am1[30] ) );
INV_X4 _u0_u1_U133  ( .A(1'b0), .ZN(_u0_u1_ch_am1[29] ) );
INV_X4 _u0_u1_U131  ( .A(1'b0), .ZN(_u0_u1_ch_am1[28] ) );
INV_X4 _u0_u1_U129  ( .A(1'b0), .ZN(_u0_u1_ch_am1[27] ) );
INV_X4 _u0_u1_U127  ( .A(1'b0), .ZN(_u0_u1_ch_am1[26] ) );
INV_X4 _u0_u1_U125  ( .A(1'b0), .ZN(_u0_u1_ch_am1[25] ) );
INV_X4 _u0_u1_U123  ( .A(1'b0), .ZN(_u0_u1_ch_am1[24] ) );
INV_X4 _u0_u1_U121  ( .A(1'b0), .ZN(_u0_u1_ch_am1[23] ) );
INV_X4 _u0_u1_U119  ( .A(1'b0), .ZN(_u0_u1_ch_am1[22] ) );
INV_X4 _u0_u1_U117  ( .A(1'b0), .ZN(_u0_u1_ch_am1[21] ) );
INV_X4 _u0_u1_U115  ( .A(1'b0), .ZN(_u0_u1_ch_am1[20] ) );
INV_X4 _u0_u1_U113  ( .A(1'b0), .ZN(_u0_u1_ch_am1[19] ) );
INV_X4 _u0_u1_U111  ( .A(1'b0), .ZN(_u0_u1_ch_am1[18] ) );
INV_X4 _u0_u1_U109  ( .A(1'b0), .ZN(_u0_u1_ch_am1[17] ) );
INV_X4 _u0_u1_U107  ( .A(1'b0), .ZN(_u0_u1_ch_am1[16] ) );
INV_X4 _u0_u1_U105  ( .A(1'b0), .ZN(_u0_u1_ch_am1[15] ) );
INV_X4 _u0_u1_U103  ( .A(1'b0), .ZN(_u0_u1_ch_am1[14] ) );
INV_X4 _u0_u1_U101  ( .A(1'b0), .ZN(_u0_u1_ch_am1[13] ) );
INV_X4 _u0_u1_U99  ( .A(1'b0), .ZN(_u0_u1_ch_am1[12] ) );
INV_X4 _u0_u1_U97  ( .A(1'b0), .ZN(_u0_u1_ch_am1[11] ) );
INV_X4 _u0_u1_U95  ( .A(1'b0), .ZN(_u0_u1_ch_am1[10] ) );
INV_X4 _u0_u1_U93  ( .A(1'b0), .ZN(_u0_u1_ch_am1[9] ) );
INV_X4 _u0_u1_U91  ( .A(1'b0), .ZN(_u0_u1_ch_am1[8] ) );
INV_X4 _u0_u1_U89  ( .A(1'b0), .ZN(_u0_u1_ch_am1[7] ) );
INV_X4 _u0_u1_U87  ( .A(1'b0), .ZN(_u0_u1_ch_am1[6] ) );
INV_X4 _u0_u1_U85  ( .A(1'b0), .ZN(_u0_u1_ch_am1[5] ) );
INV_X4 _u0_u1_U83  ( .A(1'b0), .ZN(_u0_u1_ch_am1[4] ) );
INV_X4 _u0_u1_U81  ( .A(1'b1), .ZN(_u0_u1_ch_am1[3] ) );
INV_X4 _u0_u1_U79  ( .A(1'b1), .ZN(_u0_u1_ch_am1[2] ) );
INV_X4 _u0_u1_U77  ( .A(1'b1), .ZN(_u0_u1_ch_am1[1] ) );
INV_X4 _u0_u1_U75  ( .A(1'b1), .ZN(_u0_u1_ch_am1[0] ) );
INV_X4 _u0_u1_U73  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[31] ) );
INV_X4 _u0_u1_U71  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[30] ) );
INV_X4 _u0_u1_U69  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[29] ) );
INV_X4 _u0_u1_U67  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[28] ) );
INV_X4 _u0_u1_U65  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[27] ) );
INV_X4 _u0_u1_U63  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[26] ) );
INV_X4 _u0_u1_U61  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[25] ) );
INV_X4 _u0_u1_U59  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[24] ) );
INV_X4 _u0_u1_U57  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[23] ) );
INV_X4 _u0_u1_U55  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[22] ) );
INV_X4 _u0_u1_U53  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[21] ) );
INV_X4 _u0_u1_U51  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[20] ) );
INV_X4 _u0_u1_U49  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[19] ) );
INV_X4 _u0_u1_U47  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[18] ) );
INV_X4 _u0_u1_U45  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[17] ) );
INV_X4 _u0_u1_U43  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[16] ) );
INV_X4 _u0_u1_U41  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[15] ) );
INV_X4 _u0_u1_U39  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[14] ) );
INV_X4 _u0_u1_U37  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[13] ) );
INV_X4 _u0_u1_U35  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[12] ) );
INV_X4 _u0_u1_U33  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[11] ) );
INV_X4 _u0_u1_U31  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[10] ) );
INV_X4 _u0_u1_U29  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[9] ) );
INV_X4 _u0_u1_U27  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[8] ) );
INV_X4 _u0_u1_U25  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[7] ) );
INV_X4 _u0_u1_U23  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[6] ) );
INV_X4 _u0_u1_U21  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[5] ) );
INV_X4 _u0_u1_U19  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[4] ) );
INV_X4 _u0_u1_U17  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[3] ) );
INV_X4 _u0_u1_U15  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[2] ) );
INV_X4 _u0_u1_U13  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[1] ) );
INV_X4 _u0_u1_U11  ( .A(1'b1), .ZN(_u0_u1_sw_pointer[0] ) );
INV_X4 _u0_u1_U9  ( .A(1'b1), .ZN(_u0_u1_ch_stop ) );
INV_X4 _u0_u1_U7  ( .A(1'b1), .ZN(_u0_u1_ch_dis ) );
INV_X4 _u0_u1_U5  ( .A(1'b1), .ZN(_u0_u1_int ) );
INV_X4 _u0_u2_U585  ( .A(1'b1), .ZN(_u0_u2_pointer[31] ) );
INV_X4 _u0_u2_U583  ( .A(1'b1), .ZN(_u0_u2_pointer[30] ) );
INV_X4 _u0_u2_U581  ( .A(1'b1), .ZN(_u0_u2_pointer[29] ) );
INV_X4 _u0_u2_U579  ( .A(1'b1), .ZN(_u0_u2_pointer[28] ) );
INV_X4 _u0_u2_U577  ( .A(1'b1), .ZN(_u0_u2_pointer[27] ) );
INV_X4 _u0_u2_U575  ( .A(1'b1), .ZN(_u0_u2_pointer[26] ) );
INV_X4 _u0_u2_U573  ( .A(1'b1), .ZN(_u0_u2_pointer[25] ) );
INV_X4 _u0_u2_U571  ( .A(1'b1), .ZN(_u0_u2_pointer[24] ) );
INV_X4 _u0_u2_U569  ( .A(1'b1), .ZN(_u0_u2_pointer[23] ) );
INV_X4 _u0_u2_U567  ( .A(1'b1), .ZN(_u0_u2_pointer[22] ) );
INV_X4 _u0_u2_U565  ( .A(1'b1), .ZN(_u0_u2_pointer[21] ) );
INV_X4 _u0_u2_U563  ( .A(1'b1), .ZN(_u0_u2_pointer[20] ) );
INV_X4 _u0_u2_U561  ( .A(1'b1), .ZN(_u0_u2_pointer[19] ) );
INV_X4 _u0_u2_U559  ( .A(1'b1), .ZN(_u0_u2_pointer[18] ) );
INV_X4 _u0_u2_U557  ( .A(1'b1), .ZN(_u0_u2_pointer[17] ) );
INV_X4 _u0_u2_U555  ( .A(1'b1), .ZN(_u0_u2_pointer[16] ) );
INV_X4 _u0_u2_U553  ( .A(1'b1), .ZN(_u0_u2_pointer[15] ) );
INV_X4 _u0_u2_U551  ( .A(1'b1), .ZN(_u0_u2_pointer[14] ) );
INV_X4 _u0_u2_U549  ( .A(1'b1), .ZN(_u0_u2_pointer[13] ) );
INV_X4 _u0_u2_U547  ( .A(1'b1), .ZN(_u0_u2_pointer[12] ) );
INV_X4 _u0_u2_U545  ( .A(1'b1), .ZN(_u0_u2_pointer[11] ) );
INV_X4 _u0_u2_U543  ( .A(1'b1), .ZN(_u0_u2_pointer[10] ) );
INV_X4 _u0_u2_U541  ( .A(1'b1), .ZN(_u0_u2_pointer[9] ) );
INV_X4 _u0_u2_U539  ( .A(1'b1), .ZN(_u0_u2_pointer[8] ) );
INV_X4 _u0_u2_U537  ( .A(1'b1), .ZN(_u0_u2_pointer[7] ) );
INV_X4 _u0_u2_U535  ( .A(1'b1), .ZN(_u0_u2_pointer[6] ) );
INV_X4 _u0_u2_U533  ( .A(1'b1), .ZN(_u0_u2_pointer[5] ) );
INV_X4 _u0_u2_U531  ( .A(1'b1), .ZN(_u0_u2_pointer[4] ) );
INV_X4 _u0_u2_U529  ( .A(1'b1), .ZN(_u0_u2_pointer[3] ) );
INV_X4 _u0_u2_U527  ( .A(1'b1), .ZN(_u0_u2_pointer[2] ) );
INV_X4 _u0_u2_U525  ( .A(1'b1), .ZN(_u0_u2_pointer[1] ) );
INV_X4 _u0_u2_U523  ( .A(1'b1), .ZN(_u0_u2_pointer[0] ) );
INV_X4 _u0_u2_U521  ( .A(1'b1), .ZN(_u0_u2_pointer_s[31] ) );
INV_X4 _u0_u2_U519  ( .A(1'b1), .ZN(_u0_u2_pointer_s[30] ) );
INV_X4 _u0_u2_U517  ( .A(1'b1), .ZN(_u0_u2_pointer_s[29] ) );
INV_X4 _u0_u2_U515  ( .A(1'b1), .ZN(_u0_u2_pointer_s[28] ) );
INV_X4 _u0_u2_U513  ( .A(1'b1), .ZN(_u0_u2_pointer_s[27] ) );
INV_X4 _u0_u2_U511  ( .A(1'b1), .ZN(_u0_u2_pointer_s[26] ) );
INV_X4 _u0_u2_U509  ( .A(1'b1), .ZN(_u0_u2_pointer_s[25] ) );
INV_X4 _u0_u2_U507  ( .A(1'b1), .ZN(_u0_u2_pointer_s[24] ) );
INV_X4 _u0_u2_U505  ( .A(1'b1), .ZN(_u0_u2_pointer_s[23] ) );
INV_X4 _u0_u2_U503  ( .A(1'b1), .ZN(_u0_u2_pointer_s[22] ) );
INV_X4 _u0_u2_U501  ( .A(1'b1), .ZN(_u0_u2_pointer_s[21] ) );
INV_X4 _u0_u2_U499  ( .A(1'b1), .ZN(_u0_u2_pointer_s[20] ) );
INV_X4 _u0_u2_U497  ( .A(1'b1), .ZN(_u0_u2_pointer_s[19] ) );
INV_X4 _u0_u2_U495  ( .A(1'b1), .ZN(_u0_u2_pointer_s[18] ) );
INV_X4 _u0_u2_U493  ( .A(1'b1), .ZN(_u0_u2_pointer_s[17] ) );
INV_X4 _u0_u2_U491  ( .A(1'b1), .ZN(_u0_u2_pointer_s[16] ) );
INV_X4 _u0_u2_U489  ( .A(1'b1), .ZN(_u0_u2_pointer_s[15] ) );
INV_X4 _u0_u2_U487  ( .A(1'b1), .ZN(_u0_u2_pointer_s[14] ) );
INV_X4 _u0_u2_U485  ( .A(1'b1), .ZN(_u0_u2_pointer_s[13] ) );
INV_X4 _u0_u2_U483  ( .A(1'b1), .ZN(_u0_u2_pointer_s[12] ) );
INV_X4 _u0_u2_U481  ( .A(1'b1), .ZN(_u0_u2_pointer_s[11] ) );
INV_X4 _u0_u2_U479  ( .A(1'b1), .ZN(_u0_u2_pointer_s[10] ) );
INV_X4 _u0_u2_U477  ( .A(1'b1), .ZN(_u0_u2_pointer_s[9] ) );
INV_X4 _u0_u2_U475  ( .A(1'b1), .ZN(_u0_u2_pointer_s[8] ) );
INV_X4 _u0_u2_U473  ( .A(1'b1), .ZN(_u0_u2_pointer_s[7] ) );
INV_X4 _u0_u2_U471  ( .A(1'b1), .ZN(_u0_u2_pointer_s[6] ) );
INV_X4 _u0_u2_U469  ( .A(1'b1), .ZN(_u0_u2_pointer_s[5] ) );
INV_X4 _u0_u2_U467  ( .A(1'b1), .ZN(_u0_u2_pointer_s[4] ) );
INV_X4 _u0_u2_U465  ( .A(1'b1), .ZN(_u0_u2_pointer_s[3] ) );
INV_X4 _u0_u2_U463  ( .A(1'b1), .ZN(_u0_u2_pointer_s[2] ) );
INV_X4 _u0_u2_U461  ( .A(1'b1), .ZN(_u0_u2_pointer_s[1] ) );
INV_X4 _u0_u2_U459  ( .A(1'b1), .ZN(_u0_u2_pointer_s[0] ) );
INV_X4 _u0_u2_U457  ( .A(1'b1), .ZN(_u0_u2_ch_csr[31] ) );
INV_X4 _u0_u2_U455  ( .A(1'b1), .ZN(_u0_u2_ch_csr[30] ) );
INV_X4 _u0_u2_U453  ( .A(1'b1), .ZN(_u0_u2_ch_csr[29] ) );
INV_X4 _u0_u2_U451  ( .A(1'b1), .ZN(_u0_u2_ch_csr[28] ) );
INV_X4 _u0_u2_U449  ( .A(1'b1), .ZN(_u0_u2_ch_csr[27] ) );
INV_X4 _u0_u2_U447  ( .A(1'b1), .ZN(_u0_u2_ch_csr[26] ) );
INV_X4 _u0_u2_U445  ( .A(1'b1), .ZN(_u0_u2_ch_csr[25] ) );
INV_X4 _u0_u2_U443  ( .A(1'b1), .ZN(_u0_u2_ch_csr[24] ) );
INV_X4 _u0_u2_U441  ( .A(1'b1), .ZN(_u0_u2_ch_csr[23] ) );
INV_X4 _u0_u2_U439  ( .A(1'b1), .ZN(_u0_u2_ch_csr[22] ) );
INV_X4 _u0_u2_U437  ( .A(1'b1), .ZN(_u0_u2_ch_csr[21] ) );
INV_X4 _u0_u2_U435  ( .A(1'b1), .ZN(_u0_u2_ch_csr[20] ) );
INV_X4 _u0_u2_U433  ( .A(1'b1), .ZN(_u0_u2_ch_csr[19] ) );
INV_X4 _u0_u2_U431  ( .A(1'b1), .ZN(_u0_u2_ch_csr[18] ) );
INV_X4 _u0_u2_U429  ( .A(1'b1), .ZN(_u0_u2_ch_csr[17] ) );
INV_X4 _u0_u2_U427  ( .A(1'b1), .ZN(_u0_u2_ch_csr[16] ) );
INV_X4 _u0_u2_U425  ( .A(1'b1), .ZN(_u0_u2_ch_csr[15] ) );
INV_X4 _u0_u2_U423  ( .A(1'b1), .ZN(_u0_u2_ch_csr[14] ) );
INV_X4 _u0_u2_U421  ( .A(1'b1), .ZN(_u0_u2_ch_csr[13] ) );
INV_X4 _u0_u2_U419  ( .A(1'b1), .ZN(_u0_u2_ch_csr[12] ) );
INV_X4 _u0_u2_U417  ( .A(1'b1), .ZN(_u0_u2_ch_csr[11] ) );
INV_X4 _u0_u2_U415  ( .A(1'b1), .ZN(_u0_u2_ch_csr[10] ) );
INV_X4 _u0_u2_U413  ( .A(1'b1), .ZN(_u0_u2_ch_csr[9] ) );
INV_X4 _u0_u2_U411  ( .A(1'b1), .ZN(_u0_u2_ch_csr[8] ) );
INV_X4 _u0_u2_U409  ( .A(1'b1), .ZN(_u0_u2_ch_csr[7] ) );
INV_X4 _u0_u2_U407  ( .A(1'b1), .ZN(_u0_u2_ch_csr[6] ) );
INV_X4 _u0_u2_U405  ( .A(1'b1), .ZN(_u0_u2_ch_csr[5] ) );
INV_X4 _u0_u2_U403  ( .A(1'b1), .ZN(_u0_u2_ch_csr[4] ) );
INV_X4 _u0_u2_U401  ( .A(1'b1), .ZN(_u0_u2_ch_csr[3] ) );
INV_X4 _u0_u2_U399  ( .A(1'b1), .ZN(_u0_u2_ch_csr[2] ) );
INV_X4 _u0_u2_U397  ( .A(1'b1), .ZN(_u0_u2_ch_csr[1] ) );
INV_X4 _u0_u2_U395  ( .A(1'b1), .ZN(_u0_u2_ch_csr[0] ) );
INV_X4 _u0_u2_U393  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[31] ) );
INV_X4 _u0_u2_U391  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[30] ) );
INV_X4 _u0_u2_U389  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[29] ) );
INV_X4 _u0_u2_U387  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[28] ) );
INV_X4 _u0_u2_U385  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[27] ) );
INV_X4 _u0_u2_U383  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[26] ) );
INV_X4 _u0_u2_U381  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[25] ) );
INV_X4 _u0_u2_U379  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[24] ) );
INV_X4 _u0_u2_U377  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[23] ) );
INV_X4 _u0_u2_U375  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[22] ) );
INV_X4 _u0_u2_U373  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[21] ) );
INV_X4 _u0_u2_U371  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[20] ) );
INV_X4 _u0_u2_U369  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[19] ) );
INV_X4 _u0_u2_U367  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[18] ) );
INV_X4 _u0_u2_U365  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[17] ) );
INV_X4 _u0_u2_U363  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[16] ) );
INV_X4 _u0_u2_U361  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[15] ) );
INV_X4 _u0_u2_U359  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[14] ) );
INV_X4 _u0_u2_U357  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[13] ) );
INV_X4 _u0_u2_U355  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[12] ) );
INV_X4 _u0_u2_U353  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[11] ) );
INV_X4 _u0_u2_U351  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[10] ) );
INV_X4 _u0_u2_U349  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[9] ) );
INV_X4 _u0_u2_U347  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[8] ) );
INV_X4 _u0_u2_U345  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[7] ) );
INV_X4 _u0_u2_U343  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[6] ) );
INV_X4 _u0_u2_U341  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[5] ) );
INV_X4 _u0_u2_U339  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[4] ) );
INV_X4 _u0_u2_U337  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[3] ) );
INV_X4 _u0_u2_U335  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[2] ) );
INV_X4 _u0_u2_U333  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[1] ) );
INV_X4 _u0_u2_U331  ( .A(1'b1), .ZN(_u0_u2_ch_txsz[0] ) );
INV_X4 _u0_u2_U329  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[31] ) );
INV_X4 _u0_u2_U327  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[30] ) );
INV_X4 _u0_u2_U325  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[29] ) );
INV_X4 _u0_u2_U323  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[28] ) );
INV_X4 _u0_u2_U321  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[27] ) );
INV_X4 _u0_u2_U319  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[26] ) );
INV_X4 _u0_u2_U317  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[25] ) );
INV_X4 _u0_u2_U315  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[24] ) );
INV_X4 _u0_u2_U313  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[23] ) );
INV_X4 _u0_u2_U311  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[22] ) );
INV_X4 _u0_u2_U309  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[21] ) );
INV_X4 _u0_u2_U307  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[20] ) );
INV_X4 _u0_u2_U305  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[19] ) );
INV_X4 _u0_u2_U303  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[18] ) );
INV_X4 _u0_u2_U301  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[17] ) );
INV_X4 _u0_u2_U299  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[16] ) );
INV_X4 _u0_u2_U297  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[15] ) );
INV_X4 _u0_u2_U295  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[14] ) );
INV_X4 _u0_u2_U293  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[13] ) );
INV_X4 _u0_u2_U291  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[12] ) );
INV_X4 _u0_u2_U289  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[11] ) );
INV_X4 _u0_u2_U287  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[10] ) );
INV_X4 _u0_u2_U285  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[9] ) );
INV_X4 _u0_u2_U283  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[8] ) );
INV_X4 _u0_u2_U281  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[7] ) );
INV_X4 _u0_u2_U279  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[6] ) );
INV_X4 _u0_u2_U277  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[5] ) );
INV_X4 _u0_u2_U275  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[4] ) );
INV_X4 _u0_u2_U273  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[3] ) );
INV_X4 _u0_u2_U271  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[2] ) );
INV_X4 _u0_u2_U269  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[1] ) );
INV_X4 _u0_u2_U267  ( .A(1'b1), .ZN(_u0_u2_ch_adr0[0] ) );
INV_X4 _u0_u2_U265  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[31] ) );
INV_X4 _u0_u2_U263  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[30] ) );
INV_X4 _u0_u2_U261  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[29] ) );
INV_X4 _u0_u2_U259  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[28] ) );
INV_X4 _u0_u2_U257  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[27] ) );
INV_X4 _u0_u2_U255  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[26] ) );
INV_X4 _u0_u2_U253  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[25] ) );
INV_X4 _u0_u2_U251  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[24] ) );
INV_X4 _u0_u2_U249  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[23] ) );
INV_X4 _u0_u2_U247  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[22] ) );
INV_X4 _u0_u2_U245  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[21] ) );
INV_X4 _u0_u2_U243  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[20] ) );
INV_X4 _u0_u2_U241  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[19] ) );
INV_X4 _u0_u2_U239  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[18] ) );
INV_X4 _u0_u2_U237  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[17] ) );
INV_X4 _u0_u2_U235  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[16] ) );
INV_X4 _u0_u2_U233  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[15] ) );
INV_X4 _u0_u2_U231  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[14] ) );
INV_X4 _u0_u2_U229  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[13] ) );
INV_X4 _u0_u2_U227  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[12] ) );
INV_X4 _u0_u2_U225  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[11] ) );
INV_X4 _u0_u2_U223  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[10] ) );
INV_X4 _u0_u2_U221  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[9] ) );
INV_X4 _u0_u2_U219  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[8] ) );
INV_X4 _u0_u2_U217  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[7] ) );
INV_X4 _u0_u2_U215  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[6] ) );
INV_X4 _u0_u2_U213  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[5] ) );
INV_X4 _u0_u2_U211  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[4] ) );
INV_X4 _u0_u2_U209  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[3] ) );
INV_X4 _u0_u2_U207  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[2] ) );
INV_X4 _u0_u2_U205  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[1] ) );
INV_X4 _u0_u2_U203  ( .A(1'b1), .ZN(_u0_u2_ch_adr1[0] ) );
INV_X4 _u0_u2_U201  ( .A(1'b0), .ZN(_u0_u2_ch_am0[31] ) );
INV_X4 _u0_u2_U199  ( .A(1'b0), .ZN(_u0_u2_ch_am0[30] ) );
INV_X4 _u0_u2_U197  ( .A(1'b0), .ZN(_u0_u2_ch_am0[29] ) );
INV_X4 _u0_u2_U195  ( .A(1'b0), .ZN(_u0_u2_ch_am0[28] ) );
INV_X4 _u0_u2_U193  ( .A(1'b0), .ZN(_u0_u2_ch_am0[27] ) );
INV_X4 _u0_u2_U191  ( .A(1'b0), .ZN(_u0_u2_ch_am0[26] ) );
INV_X4 _u0_u2_U189  ( .A(1'b0), .ZN(_u0_u2_ch_am0[25] ) );
INV_X4 _u0_u2_U187  ( .A(1'b0), .ZN(_u0_u2_ch_am0[24] ) );
INV_X4 _u0_u2_U185  ( .A(1'b0), .ZN(_u0_u2_ch_am0[23] ) );
INV_X4 _u0_u2_U183  ( .A(1'b0), .ZN(_u0_u2_ch_am0[22] ) );
INV_X4 _u0_u2_U181  ( .A(1'b0), .ZN(_u0_u2_ch_am0[21] ) );
INV_X4 _u0_u2_U179  ( .A(1'b0), .ZN(_u0_u2_ch_am0[20] ) );
INV_X4 _u0_u2_U177  ( .A(1'b0), .ZN(_u0_u2_ch_am0[19] ) );
INV_X4 _u0_u2_U175  ( .A(1'b0), .ZN(_u0_u2_ch_am0[18] ) );
INV_X4 _u0_u2_U173  ( .A(1'b0), .ZN(_u0_u2_ch_am0[17] ) );
INV_X4 _u0_u2_U171  ( .A(1'b0), .ZN(_u0_u2_ch_am0[16] ) );
INV_X4 _u0_u2_U169  ( .A(1'b0), .ZN(_u0_u2_ch_am0[15] ) );
INV_X4 _u0_u2_U167  ( .A(1'b0), .ZN(_u0_u2_ch_am0[14] ) );
INV_X4 _u0_u2_U165  ( .A(1'b0), .ZN(_u0_u2_ch_am0[13] ) );
INV_X4 _u0_u2_U163  ( .A(1'b0), .ZN(_u0_u2_ch_am0[12] ) );
INV_X4 _u0_u2_U161  ( .A(1'b0), .ZN(_u0_u2_ch_am0[11] ) );
INV_X4 _u0_u2_U159  ( .A(1'b0), .ZN(_u0_u2_ch_am0[10] ) );
INV_X4 _u0_u2_U157  ( .A(1'b0), .ZN(_u0_u2_ch_am0[9] ) );
INV_X4 _u0_u2_U155  ( .A(1'b0), .ZN(_u0_u2_ch_am0[8] ) );
INV_X4 _u0_u2_U153  ( .A(1'b0), .ZN(_u0_u2_ch_am0[7] ) );
INV_X4 _u0_u2_U151  ( .A(1'b0), .ZN(_u0_u2_ch_am0[6] ) );
INV_X4 _u0_u2_U149  ( .A(1'b0), .ZN(_u0_u2_ch_am0[5] ) );
INV_X4 _u0_u2_U147  ( .A(1'b0), .ZN(_u0_u2_ch_am0[4] ) );
INV_X4 _u0_u2_U145  ( .A(1'b1), .ZN(_u0_u2_ch_am0[3] ) );
INV_X4 _u0_u2_U143  ( .A(1'b1), .ZN(_u0_u2_ch_am0[2] ) );
INV_X4 _u0_u2_U141  ( .A(1'b1), .ZN(_u0_u2_ch_am0[1] ) );
INV_X4 _u0_u2_U139  ( .A(1'b1), .ZN(_u0_u2_ch_am0[0] ) );
INV_X4 _u0_u2_U137  ( .A(1'b0), .ZN(_u0_u2_ch_am1[31] ) );
INV_X4 _u0_u2_U135  ( .A(1'b0), .ZN(_u0_u2_ch_am1[30] ) );
INV_X4 _u0_u2_U133  ( .A(1'b0), .ZN(_u0_u2_ch_am1[29] ) );
INV_X4 _u0_u2_U131  ( .A(1'b0), .ZN(_u0_u2_ch_am1[28] ) );
INV_X4 _u0_u2_U129  ( .A(1'b0), .ZN(_u0_u2_ch_am1[27] ) );
INV_X4 _u0_u2_U127  ( .A(1'b0), .ZN(_u0_u2_ch_am1[26] ) );
INV_X4 _u0_u2_U125  ( .A(1'b0), .ZN(_u0_u2_ch_am1[25] ) );
INV_X4 _u0_u2_U123  ( .A(1'b0), .ZN(_u0_u2_ch_am1[24] ) );
INV_X4 _u0_u2_U121  ( .A(1'b0), .ZN(_u0_u2_ch_am1[23] ) );
INV_X4 _u0_u2_U119  ( .A(1'b0), .ZN(_u0_u2_ch_am1[22] ) );
INV_X4 _u0_u2_U117  ( .A(1'b0), .ZN(_u0_u2_ch_am1[21] ) );
INV_X4 _u0_u2_U115  ( .A(1'b0), .ZN(_u0_u2_ch_am1[20] ) );
INV_X4 _u0_u2_U113  ( .A(1'b0), .ZN(_u0_u2_ch_am1[19] ) );
INV_X4 _u0_u2_U111  ( .A(1'b0), .ZN(_u0_u2_ch_am1[18] ) );
INV_X4 _u0_u2_U109  ( .A(1'b0), .ZN(_u0_u2_ch_am1[17] ) );
INV_X4 _u0_u2_U107  ( .A(1'b0), .ZN(_u0_u2_ch_am1[16] ) );
INV_X4 _u0_u2_U105  ( .A(1'b0), .ZN(_u0_u2_ch_am1[15] ) );
INV_X4 _u0_u2_U103  ( .A(1'b0), .ZN(_u0_u2_ch_am1[14] ) );
INV_X4 _u0_u2_U101  ( .A(1'b0), .ZN(_u0_u2_ch_am1[13] ) );
INV_X4 _u0_u2_U99  ( .A(1'b0), .ZN(_u0_u2_ch_am1[12] ) );
INV_X4 _u0_u2_U97  ( .A(1'b0), .ZN(_u0_u2_ch_am1[11] ) );
INV_X4 _u0_u2_U95  ( .A(1'b0), .ZN(_u0_u2_ch_am1[10] ) );
INV_X4 _u0_u2_U93  ( .A(1'b0), .ZN(_u0_u2_ch_am1[9] ) );
INV_X4 _u0_u2_U91  ( .A(1'b0), .ZN(_u0_u2_ch_am1[8] ) );
INV_X4 _u0_u2_U89  ( .A(1'b0), .ZN(_u0_u2_ch_am1[7] ) );
INV_X4 _u0_u2_U87  ( .A(1'b0), .ZN(_u0_u2_ch_am1[6] ) );
INV_X4 _u0_u2_U85  ( .A(1'b0), .ZN(_u0_u2_ch_am1[5] ) );
INV_X4 _u0_u2_U83  ( .A(1'b0), .ZN(_u0_u2_ch_am1[4] ) );
INV_X4 _u0_u2_U81  ( .A(1'b1), .ZN(_u0_u2_ch_am1[3] ) );
INV_X4 _u0_u2_U79  ( .A(1'b1), .ZN(_u0_u2_ch_am1[2] ) );
INV_X4 _u0_u2_U77  ( .A(1'b1), .ZN(_u0_u2_ch_am1[1] ) );
INV_X4 _u0_u2_U75  ( .A(1'b1), .ZN(_u0_u2_ch_am1[0] ) );
INV_X4 _u0_u2_U73  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[31] ) );
INV_X4 _u0_u2_U71  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[30] ) );
INV_X4 _u0_u2_U69  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[29] ) );
INV_X4 _u0_u2_U67  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[28] ) );
INV_X4 _u0_u2_U65  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[27] ) );
INV_X4 _u0_u2_U63  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[26] ) );
INV_X4 _u0_u2_U61  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[25] ) );
INV_X4 _u0_u2_U59  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[24] ) );
INV_X4 _u0_u2_U57  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[23] ) );
INV_X4 _u0_u2_U55  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[22] ) );
INV_X4 _u0_u2_U53  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[21] ) );
INV_X4 _u0_u2_U51  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[20] ) );
INV_X4 _u0_u2_U49  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[19] ) );
INV_X4 _u0_u2_U47  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[18] ) );
INV_X4 _u0_u2_U45  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[17] ) );
INV_X4 _u0_u2_U43  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[16] ) );
INV_X4 _u0_u2_U41  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[15] ) );
INV_X4 _u0_u2_U39  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[14] ) );
INV_X4 _u0_u2_U37  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[13] ) );
INV_X4 _u0_u2_U35  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[12] ) );
INV_X4 _u0_u2_U33  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[11] ) );
INV_X4 _u0_u2_U31  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[10] ) );
INV_X4 _u0_u2_U29  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[9] ) );
INV_X4 _u0_u2_U27  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[8] ) );
INV_X4 _u0_u2_U25  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[7] ) );
INV_X4 _u0_u2_U23  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[6] ) );
INV_X4 _u0_u2_U21  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[5] ) );
INV_X4 _u0_u2_U19  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[4] ) );
INV_X4 _u0_u2_U17  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[3] ) );
INV_X4 _u0_u2_U15  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[2] ) );
INV_X4 _u0_u2_U13  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[1] ) );
INV_X4 _u0_u2_U11  ( .A(1'b1), .ZN(_u0_u2_sw_pointer[0] ) );
INV_X4 _u0_u2_U9  ( .A(1'b1), .ZN(_u0_u2_ch_stop ) );
INV_X4 _u0_u2_U7  ( .A(1'b1), .ZN(_u0_u2_ch_dis ) );
INV_X4 _u0_u2_U5  ( .A(1'b1), .ZN(_u0_u2_int ) );
INV_X4 _u0_u3_U585  ( .A(1'b1), .ZN(_u0_u3_pointer[31] ) );
INV_X4 _u0_u3_U583  ( .A(1'b1), .ZN(_u0_u3_pointer[30] ) );
INV_X4 _u0_u3_U581  ( .A(1'b1), .ZN(_u0_u3_pointer[29] ) );
INV_X4 _u0_u3_U579  ( .A(1'b1), .ZN(_u0_u3_pointer[28] ) );
INV_X4 _u0_u3_U577  ( .A(1'b1), .ZN(_u0_u3_pointer[27] ) );
INV_X4 _u0_u3_U575  ( .A(1'b1), .ZN(_u0_u3_pointer[26] ) );
INV_X4 _u0_u3_U573  ( .A(1'b1), .ZN(_u0_u3_pointer[25] ) );
INV_X4 _u0_u3_U571  ( .A(1'b1), .ZN(_u0_u3_pointer[24] ) );
INV_X4 _u0_u3_U569  ( .A(1'b1), .ZN(_u0_u3_pointer[23] ) );
INV_X4 _u0_u3_U567  ( .A(1'b1), .ZN(_u0_u3_pointer[22] ) );
INV_X4 _u0_u3_U565  ( .A(1'b1), .ZN(_u0_u3_pointer[21] ) );
INV_X4 _u0_u3_U563  ( .A(1'b1), .ZN(_u0_u3_pointer[20] ) );
INV_X4 _u0_u3_U561  ( .A(1'b1), .ZN(_u0_u3_pointer[19] ) );
INV_X4 _u0_u3_U559  ( .A(1'b1), .ZN(_u0_u3_pointer[18] ) );
INV_X4 _u0_u3_U557  ( .A(1'b1), .ZN(_u0_u3_pointer[17] ) );
INV_X4 _u0_u3_U555  ( .A(1'b1), .ZN(_u0_u3_pointer[16] ) );
INV_X4 _u0_u3_U553  ( .A(1'b1), .ZN(_u0_u3_pointer[15] ) );
INV_X4 _u0_u3_U551  ( .A(1'b1), .ZN(_u0_u3_pointer[14] ) );
INV_X4 _u0_u3_U549  ( .A(1'b1), .ZN(_u0_u3_pointer[13] ) );
INV_X4 _u0_u3_U547  ( .A(1'b1), .ZN(_u0_u3_pointer[12] ) );
INV_X4 _u0_u3_U545  ( .A(1'b1), .ZN(_u0_u3_pointer[11] ) );
INV_X4 _u0_u3_U543  ( .A(1'b1), .ZN(_u0_u3_pointer[10] ) );
INV_X4 _u0_u3_U541  ( .A(1'b1), .ZN(_u0_u3_pointer[9] ) );
INV_X4 _u0_u3_U539  ( .A(1'b1), .ZN(_u0_u3_pointer[8] ) );
INV_X4 _u0_u3_U537  ( .A(1'b1), .ZN(_u0_u3_pointer[7] ) );
INV_X4 _u0_u3_U535  ( .A(1'b1), .ZN(_u0_u3_pointer[6] ) );
INV_X4 _u0_u3_U533  ( .A(1'b1), .ZN(_u0_u3_pointer[5] ) );
INV_X4 _u0_u3_U531  ( .A(1'b1), .ZN(_u0_u3_pointer[4] ) );
INV_X4 _u0_u3_U529  ( .A(1'b1), .ZN(_u0_u3_pointer[3] ) );
INV_X4 _u0_u3_U527  ( .A(1'b1), .ZN(_u0_u3_pointer[2] ) );
INV_X4 _u0_u3_U525  ( .A(1'b1), .ZN(_u0_u3_pointer[1] ) );
INV_X4 _u0_u3_U523  ( .A(1'b1), .ZN(_u0_u3_pointer[0] ) );
INV_X4 _u0_u3_U521  ( .A(1'b1), .ZN(_u0_u3_pointer_s[31] ) );
INV_X4 _u0_u3_U519  ( .A(1'b1), .ZN(_u0_u3_pointer_s[30] ) );
INV_X4 _u0_u3_U517  ( .A(1'b1), .ZN(_u0_u3_pointer_s[29] ) );
INV_X4 _u0_u3_U515  ( .A(1'b1), .ZN(_u0_u3_pointer_s[28] ) );
INV_X4 _u0_u3_U513  ( .A(1'b1), .ZN(_u0_u3_pointer_s[27] ) );
INV_X4 _u0_u3_U511  ( .A(1'b1), .ZN(_u0_u3_pointer_s[26] ) );
INV_X4 _u0_u3_U509  ( .A(1'b1), .ZN(_u0_u3_pointer_s[25] ) );
INV_X4 _u0_u3_U507  ( .A(1'b1), .ZN(_u0_u3_pointer_s[24] ) );
INV_X4 _u0_u3_U505  ( .A(1'b1), .ZN(_u0_u3_pointer_s[23] ) );
INV_X4 _u0_u3_U503  ( .A(1'b1), .ZN(_u0_u3_pointer_s[22] ) );
INV_X4 _u0_u3_U501  ( .A(1'b1), .ZN(_u0_u3_pointer_s[21] ) );
INV_X4 _u0_u3_U499  ( .A(1'b1), .ZN(_u0_u3_pointer_s[20] ) );
INV_X4 _u0_u3_U497  ( .A(1'b1), .ZN(_u0_u3_pointer_s[19] ) );
INV_X4 _u0_u3_U495  ( .A(1'b1), .ZN(_u0_u3_pointer_s[18] ) );
INV_X4 _u0_u3_U493  ( .A(1'b1), .ZN(_u0_u3_pointer_s[17] ) );
INV_X4 _u0_u3_U491  ( .A(1'b1), .ZN(_u0_u3_pointer_s[16] ) );
INV_X4 _u0_u3_U489  ( .A(1'b1), .ZN(_u0_u3_pointer_s[15] ) );
INV_X4 _u0_u3_U487  ( .A(1'b1), .ZN(_u0_u3_pointer_s[14] ) );
INV_X4 _u0_u3_U485  ( .A(1'b1), .ZN(_u0_u3_pointer_s[13] ) );
INV_X4 _u0_u3_U483  ( .A(1'b1), .ZN(_u0_u3_pointer_s[12] ) );
INV_X4 _u0_u3_U481  ( .A(1'b1), .ZN(_u0_u3_pointer_s[11] ) );
INV_X4 _u0_u3_U479  ( .A(1'b1), .ZN(_u0_u3_pointer_s[10] ) );
INV_X4 _u0_u3_U477  ( .A(1'b1), .ZN(_u0_u3_pointer_s[9] ) );
INV_X4 _u0_u3_U475  ( .A(1'b1), .ZN(_u0_u3_pointer_s[8] ) );
INV_X4 _u0_u3_U473  ( .A(1'b1), .ZN(_u0_u3_pointer_s[7] ) );
INV_X4 _u0_u3_U471  ( .A(1'b1), .ZN(_u0_u3_pointer_s[6] ) );
INV_X4 _u0_u3_U469  ( .A(1'b1), .ZN(_u0_u3_pointer_s[5] ) );
INV_X4 _u0_u3_U467  ( .A(1'b1), .ZN(_u0_u3_pointer_s[4] ) );
INV_X4 _u0_u3_U465  ( .A(1'b1), .ZN(_u0_u3_pointer_s[3] ) );
INV_X4 _u0_u3_U463  ( .A(1'b1), .ZN(_u0_u3_pointer_s[2] ) );
INV_X4 _u0_u3_U461  ( .A(1'b1), .ZN(_u0_u3_pointer_s[1] ) );
INV_X4 _u0_u3_U459  ( .A(1'b1), .ZN(_u0_u3_pointer_s[0] ) );
INV_X4 _u0_u3_U457  ( .A(1'b1), .ZN(_u0_u3_ch_csr[31] ) );
INV_X4 _u0_u3_U455  ( .A(1'b1), .ZN(_u0_u3_ch_csr[30] ) );
INV_X4 _u0_u3_U453  ( .A(1'b1), .ZN(_u0_u3_ch_csr[29] ) );
INV_X4 _u0_u3_U451  ( .A(1'b1), .ZN(_u0_u3_ch_csr[28] ) );
INV_X4 _u0_u3_U449  ( .A(1'b1), .ZN(_u0_u3_ch_csr[27] ) );
INV_X4 _u0_u3_U447  ( .A(1'b1), .ZN(_u0_u3_ch_csr[26] ) );
INV_X4 _u0_u3_U445  ( .A(1'b1), .ZN(_u0_u3_ch_csr[25] ) );
INV_X4 _u0_u3_U443  ( .A(1'b1), .ZN(_u0_u3_ch_csr[24] ) );
INV_X4 _u0_u3_U441  ( .A(1'b1), .ZN(_u0_u3_ch_csr[23] ) );
INV_X4 _u0_u3_U439  ( .A(1'b1), .ZN(_u0_u3_ch_csr[22] ) );
INV_X4 _u0_u3_U437  ( .A(1'b1), .ZN(_u0_u3_ch_csr[21] ) );
INV_X4 _u0_u3_U435  ( .A(1'b1), .ZN(_u0_u3_ch_csr[20] ) );
INV_X4 _u0_u3_U433  ( .A(1'b1), .ZN(_u0_u3_ch_csr[19] ) );
INV_X4 _u0_u3_U431  ( .A(1'b1), .ZN(_u0_u3_ch_csr[18] ) );
INV_X4 _u0_u3_U429  ( .A(1'b1), .ZN(_u0_u3_ch_csr[17] ) );
INV_X4 _u0_u3_U427  ( .A(1'b1), .ZN(_u0_u3_ch_csr[16] ) );
INV_X4 _u0_u3_U425  ( .A(1'b1), .ZN(_u0_u3_ch_csr[15] ) );
INV_X4 _u0_u3_U423  ( .A(1'b1), .ZN(_u0_u3_ch_csr[14] ) );
INV_X4 _u0_u3_U421  ( .A(1'b1), .ZN(_u0_u3_ch_csr[13] ) );
INV_X4 _u0_u3_U419  ( .A(1'b1), .ZN(_u0_u3_ch_csr[12] ) );
INV_X4 _u0_u3_U417  ( .A(1'b1), .ZN(_u0_u3_ch_csr[11] ) );
INV_X4 _u0_u3_U415  ( .A(1'b1), .ZN(_u0_u3_ch_csr[10] ) );
INV_X4 _u0_u3_U413  ( .A(1'b1), .ZN(_u0_u3_ch_csr[9] ) );
INV_X4 _u0_u3_U411  ( .A(1'b1), .ZN(_u0_u3_ch_csr[8] ) );
INV_X4 _u0_u3_U409  ( .A(1'b1), .ZN(_u0_u3_ch_csr[7] ) );
INV_X4 _u0_u3_U407  ( .A(1'b1), .ZN(_u0_u3_ch_csr[6] ) );
INV_X4 _u0_u3_U405  ( .A(1'b1), .ZN(_u0_u3_ch_csr[5] ) );
INV_X4 _u0_u3_U403  ( .A(1'b1), .ZN(_u0_u3_ch_csr[4] ) );
INV_X4 _u0_u3_U401  ( .A(1'b1), .ZN(_u0_u3_ch_csr[3] ) );
INV_X4 _u0_u3_U399  ( .A(1'b1), .ZN(_u0_u3_ch_csr[2] ) );
INV_X4 _u0_u3_U397  ( .A(1'b1), .ZN(_u0_u3_ch_csr[1] ) );
INV_X4 _u0_u3_U395  ( .A(1'b1), .ZN(_u0_u3_ch_csr[0] ) );
INV_X4 _u0_u3_U393  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[31] ) );
INV_X4 _u0_u3_U391  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[30] ) );
INV_X4 _u0_u3_U389  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[29] ) );
INV_X4 _u0_u3_U387  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[28] ) );
INV_X4 _u0_u3_U385  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[27] ) );
INV_X4 _u0_u3_U383  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[26] ) );
INV_X4 _u0_u3_U381  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[25] ) );
INV_X4 _u0_u3_U379  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[24] ) );
INV_X4 _u0_u3_U377  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[23] ) );
INV_X4 _u0_u3_U375  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[22] ) );
INV_X4 _u0_u3_U373  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[21] ) );
INV_X4 _u0_u3_U371  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[20] ) );
INV_X4 _u0_u3_U369  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[19] ) );
INV_X4 _u0_u3_U367  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[18] ) );
INV_X4 _u0_u3_U365  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[17] ) );
INV_X4 _u0_u3_U363  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[16] ) );
INV_X4 _u0_u3_U361  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[15] ) );
INV_X4 _u0_u3_U359  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[14] ) );
INV_X4 _u0_u3_U357  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[13] ) );
INV_X4 _u0_u3_U355  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[12] ) );
INV_X4 _u0_u3_U353  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[11] ) );
INV_X4 _u0_u3_U351  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[10] ) );
INV_X4 _u0_u3_U349  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[9] ) );
INV_X4 _u0_u3_U347  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[8] ) );
INV_X4 _u0_u3_U345  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[7] ) );
INV_X4 _u0_u3_U343  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[6] ) );
INV_X4 _u0_u3_U341  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[5] ) );
INV_X4 _u0_u3_U339  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[4] ) );
INV_X4 _u0_u3_U337  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[3] ) );
INV_X4 _u0_u3_U335  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[2] ) );
INV_X4 _u0_u3_U333  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[1] ) );
INV_X4 _u0_u3_U331  ( .A(1'b1), .ZN(_u0_u3_ch_txsz[0] ) );
INV_X4 _u0_u3_U329  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[31] ) );
INV_X4 _u0_u3_U327  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[30] ) );
INV_X4 _u0_u3_U325  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[29] ) );
INV_X4 _u0_u3_U323  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[28] ) );
INV_X4 _u0_u3_U321  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[27] ) );
INV_X4 _u0_u3_U319  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[26] ) );
INV_X4 _u0_u3_U317  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[25] ) );
INV_X4 _u0_u3_U315  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[24] ) );
INV_X4 _u0_u3_U313  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[23] ) );
INV_X4 _u0_u3_U311  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[22] ) );
INV_X4 _u0_u3_U309  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[21] ) );
INV_X4 _u0_u3_U307  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[20] ) );
INV_X4 _u0_u3_U305  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[19] ) );
INV_X4 _u0_u3_U303  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[18] ) );
INV_X4 _u0_u3_U301  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[17] ) );
INV_X4 _u0_u3_U299  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[16] ) );
INV_X4 _u0_u3_U297  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[15] ) );
INV_X4 _u0_u3_U295  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[14] ) );
INV_X4 _u0_u3_U293  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[13] ) );
INV_X4 _u0_u3_U291  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[12] ) );
INV_X4 _u0_u3_U289  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[11] ) );
INV_X4 _u0_u3_U287  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[10] ) );
INV_X4 _u0_u3_U285  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[9] ) );
INV_X4 _u0_u3_U283  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[8] ) );
INV_X4 _u0_u3_U281  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[7] ) );
INV_X4 _u0_u3_U279  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[6] ) );
INV_X4 _u0_u3_U277  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[5] ) );
INV_X4 _u0_u3_U275  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[4] ) );
INV_X4 _u0_u3_U273  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[3] ) );
INV_X4 _u0_u3_U271  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[2] ) );
INV_X4 _u0_u3_U269  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[1] ) );
INV_X4 _u0_u3_U267  ( .A(1'b1), .ZN(_u0_u3_ch_adr0[0] ) );
INV_X4 _u0_u3_U265  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[31] ) );
INV_X4 _u0_u3_U263  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[30] ) );
INV_X4 _u0_u3_U261  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[29] ) );
INV_X4 _u0_u3_U259  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[28] ) );
INV_X4 _u0_u3_U257  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[27] ) );
INV_X4 _u0_u3_U255  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[26] ) );
INV_X4 _u0_u3_U253  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[25] ) );
INV_X4 _u0_u3_U251  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[24] ) );
INV_X4 _u0_u3_U249  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[23] ) );
INV_X4 _u0_u3_U247  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[22] ) );
INV_X4 _u0_u3_U245  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[21] ) );
INV_X4 _u0_u3_U243  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[20] ) );
INV_X4 _u0_u3_U241  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[19] ) );
INV_X4 _u0_u3_U239  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[18] ) );
INV_X4 _u0_u3_U237  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[17] ) );
INV_X4 _u0_u3_U235  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[16] ) );
INV_X4 _u0_u3_U233  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[15] ) );
INV_X4 _u0_u3_U231  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[14] ) );
INV_X4 _u0_u3_U229  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[13] ) );
INV_X4 _u0_u3_U227  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[12] ) );
INV_X4 _u0_u3_U225  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[11] ) );
INV_X4 _u0_u3_U223  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[10] ) );
INV_X4 _u0_u3_U221  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[9] ) );
INV_X4 _u0_u3_U219  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[8] ) );
INV_X4 _u0_u3_U217  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[7] ) );
INV_X4 _u0_u3_U215  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[6] ) );
INV_X4 _u0_u3_U213  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[5] ) );
INV_X4 _u0_u3_U211  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[4] ) );
INV_X4 _u0_u3_U209  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[3] ) );
INV_X4 _u0_u3_U207  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[2] ) );
INV_X4 _u0_u3_U205  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[1] ) );
INV_X4 _u0_u3_U203  ( .A(1'b1), .ZN(_u0_u3_ch_adr1[0] ) );
INV_X4 _u0_u3_U201  ( .A(1'b0), .ZN(_u0_u3_ch_am0[31] ) );
INV_X4 _u0_u3_U199  ( .A(1'b0), .ZN(_u0_u3_ch_am0[30] ) );
INV_X4 _u0_u3_U197  ( .A(1'b0), .ZN(_u0_u3_ch_am0[29] ) );
INV_X4 _u0_u3_U195  ( .A(1'b0), .ZN(_u0_u3_ch_am0[28] ) );
INV_X4 _u0_u3_U193  ( .A(1'b0), .ZN(_u0_u3_ch_am0[27] ) );
INV_X4 _u0_u3_U191  ( .A(1'b0), .ZN(_u0_u3_ch_am0[26] ) );
INV_X4 _u0_u3_U189  ( .A(1'b0), .ZN(_u0_u3_ch_am0[25] ) );
INV_X4 _u0_u3_U187  ( .A(1'b0), .ZN(_u0_u3_ch_am0[24] ) );
INV_X4 _u0_u3_U185  ( .A(1'b0), .ZN(_u0_u3_ch_am0[23] ) );
INV_X4 _u0_u3_U183  ( .A(1'b0), .ZN(_u0_u3_ch_am0[22] ) );
INV_X4 _u0_u3_U181  ( .A(1'b0), .ZN(_u0_u3_ch_am0[21] ) );
INV_X4 _u0_u3_U179  ( .A(1'b0), .ZN(_u0_u3_ch_am0[20] ) );
INV_X4 _u0_u3_U177  ( .A(1'b0), .ZN(_u0_u3_ch_am0[19] ) );
INV_X4 _u0_u3_U175  ( .A(1'b0), .ZN(_u0_u3_ch_am0[18] ) );
INV_X4 _u0_u3_U173  ( .A(1'b0), .ZN(_u0_u3_ch_am0[17] ) );
INV_X4 _u0_u3_U171  ( .A(1'b0), .ZN(_u0_u3_ch_am0[16] ) );
INV_X4 _u0_u3_U169  ( .A(1'b0), .ZN(_u0_u3_ch_am0[15] ) );
INV_X4 _u0_u3_U167  ( .A(1'b0), .ZN(_u0_u3_ch_am0[14] ) );
INV_X4 _u0_u3_U165  ( .A(1'b0), .ZN(_u0_u3_ch_am0[13] ) );
INV_X4 _u0_u3_U163  ( .A(1'b0), .ZN(_u0_u3_ch_am0[12] ) );
INV_X4 _u0_u3_U161  ( .A(1'b0), .ZN(_u0_u3_ch_am0[11] ) );
INV_X4 _u0_u3_U159  ( .A(1'b0), .ZN(_u0_u3_ch_am0[10] ) );
INV_X4 _u0_u3_U157  ( .A(1'b0), .ZN(_u0_u3_ch_am0[9] ) );
INV_X4 _u0_u3_U155  ( .A(1'b0), .ZN(_u0_u3_ch_am0[8] ) );
INV_X4 _u0_u3_U153  ( .A(1'b0), .ZN(_u0_u3_ch_am0[7] ) );
INV_X4 _u0_u3_U151  ( .A(1'b0), .ZN(_u0_u3_ch_am0[6] ) );
INV_X4 _u0_u3_U149  ( .A(1'b0), .ZN(_u0_u3_ch_am0[5] ) );
INV_X4 _u0_u3_U147  ( .A(1'b0), .ZN(_u0_u3_ch_am0[4] ) );
INV_X4 _u0_u3_U145  ( .A(1'b1), .ZN(_u0_u3_ch_am0[3] ) );
INV_X4 _u0_u3_U143  ( .A(1'b1), .ZN(_u0_u3_ch_am0[2] ) );
INV_X4 _u0_u3_U141  ( .A(1'b1), .ZN(_u0_u3_ch_am0[1] ) );
INV_X4 _u0_u3_U139  ( .A(1'b1), .ZN(_u0_u3_ch_am0[0] ) );
INV_X4 _u0_u3_U137  ( .A(1'b0), .ZN(_u0_u3_ch_am1[31] ) );
INV_X4 _u0_u3_U135  ( .A(1'b0), .ZN(_u0_u3_ch_am1[30] ) );
INV_X4 _u0_u3_U133  ( .A(1'b0), .ZN(_u0_u3_ch_am1[29] ) );
INV_X4 _u0_u3_U131  ( .A(1'b0), .ZN(_u0_u3_ch_am1[28] ) );
INV_X4 _u0_u3_U129  ( .A(1'b0), .ZN(_u0_u3_ch_am1[27] ) );
INV_X4 _u0_u3_U127  ( .A(1'b0), .ZN(_u0_u3_ch_am1[26] ) );
INV_X4 _u0_u3_U125  ( .A(1'b0), .ZN(_u0_u3_ch_am1[25] ) );
INV_X4 _u0_u3_U123  ( .A(1'b0), .ZN(_u0_u3_ch_am1[24] ) );
INV_X4 _u0_u3_U121  ( .A(1'b0), .ZN(_u0_u3_ch_am1[23] ) );
INV_X4 _u0_u3_U119  ( .A(1'b0), .ZN(_u0_u3_ch_am1[22] ) );
INV_X4 _u0_u3_U117  ( .A(1'b0), .ZN(_u0_u3_ch_am1[21] ) );
INV_X4 _u0_u3_U115  ( .A(1'b0), .ZN(_u0_u3_ch_am1[20] ) );
INV_X4 _u0_u3_U113  ( .A(1'b0), .ZN(_u0_u3_ch_am1[19] ) );
INV_X4 _u0_u3_U111  ( .A(1'b0), .ZN(_u0_u3_ch_am1[18] ) );
INV_X4 _u0_u3_U109  ( .A(1'b0), .ZN(_u0_u3_ch_am1[17] ) );
INV_X4 _u0_u3_U107  ( .A(1'b0), .ZN(_u0_u3_ch_am1[16] ) );
INV_X4 _u0_u3_U105  ( .A(1'b0), .ZN(_u0_u3_ch_am1[15] ) );
INV_X4 _u0_u3_U103  ( .A(1'b0), .ZN(_u0_u3_ch_am1[14] ) );
INV_X4 _u0_u3_U101  ( .A(1'b0), .ZN(_u0_u3_ch_am1[13] ) );
INV_X4 _u0_u3_U99  ( .A(1'b0), .ZN(_u0_u3_ch_am1[12] ) );
INV_X4 _u0_u3_U97  ( .A(1'b0), .ZN(_u0_u3_ch_am1[11] ) );
INV_X4 _u0_u3_U95  ( .A(1'b0), .ZN(_u0_u3_ch_am1[10] ) );
INV_X4 _u0_u3_U93  ( .A(1'b0), .ZN(_u0_u3_ch_am1[9] ) );
INV_X4 _u0_u3_U91  ( .A(1'b0), .ZN(_u0_u3_ch_am1[8] ) );
INV_X4 _u0_u3_U89  ( .A(1'b0), .ZN(_u0_u3_ch_am1[7] ) );
INV_X4 _u0_u3_U87  ( .A(1'b0), .ZN(_u0_u3_ch_am1[6] ) );
INV_X4 _u0_u3_U85  ( .A(1'b0), .ZN(_u0_u3_ch_am1[5] ) );
INV_X4 _u0_u3_U83  ( .A(1'b0), .ZN(_u0_u3_ch_am1[4] ) );
INV_X4 _u0_u3_U81  ( .A(1'b1), .ZN(_u0_u3_ch_am1[3] ) );
INV_X4 _u0_u3_U79  ( .A(1'b1), .ZN(_u0_u3_ch_am1[2] ) );
INV_X4 _u0_u3_U77  ( .A(1'b1), .ZN(_u0_u3_ch_am1[1] ) );
INV_X4 _u0_u3_U75  ( .A(1'b1), .ZN(_u0_u3_ch_am1[0] ) );
INV_X4 _u0_u3_U73  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[31] ) );
INV_X4 _u0_u3_U71  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[30] ) );
INV_X4 _u0_u3_U69  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[29] ) );
INV_X4 _u0_u3_U67  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[28] ) );
INV_X4 _u0_u3_U65  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[27] ) );
INV_X4 _u0_u3_U63  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[26] ) );
INV_X4 _u0_u3_U61  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[25] ) );
INV_X4 _u0_u3_U59  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[24] ) );
INV_X4 _u0_u3_U57  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[23] ) );
INV_X4 _u0_u3_U55  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[22] ) );
INV_X4 _u0_u3_U53  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[21] ) );
INV_X4 _u0_u3_U51  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[20] ) );
INV_X4 _u0_u3_U49  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[19] ) );
INV_X4 _u0_u3_U47  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[18] ) );
INV_X4 _u0_u3_U45  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[17] ) );
INV_X4 _u0_u3_U43  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[16] ) );
INV_X4 _u0_u3_U41  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[15] ) );
INV_X4 _u0_u3_U39  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[14] ) );
INV_X4 _u0_u3_U37  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[13] ) );
INV_X4 _u0_u3_U35  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[12] ) );
INV_X4 _u0_u3_U33  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[11] ) );
INV_X4 _u0_u3_U31  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[10] ) );
INV_X4 _u0_u3_U29  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[9] ) );
INV_X4 _u0_u3_U27  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[8] ) );
INV_X4 _u0_u3_U25  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[7] ) );
INV_X4 _u0_u3_U23  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[6] ) );
INV_X4 _u0_u3_U21  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[5] ) );
INV_X4 _u0_u3_U19  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[4] ) );
INV_X4 _u0_u3_U17  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[3] ) );
INV_X4 _u0_u3_U15  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[2] ) );
INV_X4 _u0_u3_U13  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[1] ) );
INV_X4 _u0_u3_U11  ( .A(1'b1), .ZN(_u0_u3_sw_pointer[0] ) );
INV_X4 _u0_u3_U9  ( .A(1'b1), .ZN(_u0_u3_ch_stop ) );
INV_X4 _u0_u3_U7  ( .A(1'b1), .ZN(_u0_u3_ch_dis ) );
INV_X4 _u0_u3_U5  ( .A(1'b1), .ZN(_u0_u3_int ) );
INV_X4 _u0_u4_U585  ( .A(1'b1), .ZN(_u0_u4_pointer[31] ) );
INV_X4 _u0_u4_U583  ( .A(1'b1), .ZN(_u0_u4_pointer[30] ) );
INV_X4 _u0_u4_U581  ( .A(1'b1), .ZN(_u0_u4_pointer[29] ) );
INV_X4 _u0_u4_U579  ( .A(1'b1), .ZN(_u0_u4_pointer[28] ) );
INV_X4 _u0_u4_U577  ( .A(1'b1), .ZN(_u0_u4_pointer[27] ) );
INV_X4 _u0_u4_U575  ( .A(1'b1), .ZN(_u0_u4_pointer[26] ) );
INV_X4 _u0_u4_U573  ( .A(1'b1), .ZN(_u0_u4_pointer[25] ) );
INV_X4 _u0_u4_U571  ( .A(1'b1), .ZN(_u0_u4_pointer[24] ) );
INV_X4 _u0_u4_U569  ( .A(1'b1), .ZN(_u0_u4_pointer[23] ) );
INV_X4 _u0_u4_U567  ( .A(1'b1), .ZN(_u0_u4_pointer[22] ) );
INV_X4 _u0_u4_U565  ( .A(1'b1), .ZN(_u0_u4_pointer[21] ) );
INV_X4 _u0_u4_U563  ( .A(1'b1), .ZN(_u0_u4_pointer[20] ) );
INV_X4 _u0_u4_U561  ( .A(1'b1), .ZN(_u0_u4_pointer[19] ) );
INV_X4 _u0_u4_U559  ( .A(1'b1), .ZN(_u0_u4_pointer[18] ) );
INV_X4 _u0_u4_U557  ( .A(1'b1), .ZN(_u0_u4_pointer[17] ) );
INV_X4 _u0_u4_U555  ( .A(1'b1), .ZN(_u0_u4_pointer[16] ) );
INV_X4 _u0_u4_U553  ( .A(1'b1), .ZN(_u0_u4_pointer[15] ) );
INV_X4 _u0_u4_U551  ( .A(1'b1), .ZN(_u0_u4_pointer[14] ) );
INV_X4 _u0_u4_U549  ( .A(1'b1), .ZN(_u0_u4_pointer[13] ) );
INV_X4 _u0_u4_U547  ( .A(1'b1), .ZN(_u0_u4_pointer[12] ) );
INV_X4 _u0_u4_U545  ( .A(1'b1), .ZN(_u0_u4_pointer[11] ) );
INV_X4 _u0_u4_U543  ( .A(1'b1), .ZN(_u0_u4_pointer[10] ) );
INV_X4 _u0_u4_U541  ( .A(1'b1), .ZN(_u0_u4_pointer[9] ) );
INV_X4 _u0_u4_U539  ( .A(1'b1), .ZN(_u0_u4_pointer[8] ) );
INV_X4 _u0_u4_U537  ( .A(1'b1), .ZN(_u0_u4_pointer[7] ) );
INV_X4 _u0_u4_U535  ( .A(1'b1), .ZN(_u0_u4_pointer[6] ) );
INV_X4 _u0_u4_U533  ( .A(1'b1), .ZN(_u0_u4_pointer[5] ) );
INV_X4 _u0_u4_U531  ( .A(1'b1), .ZN(_u0_u4_pointer[4] ) );
INV_X4 _u0_u4_U529  ( .A(1'b1), .ZN(_u0_u4_pointer[3] ) );
INV_X4 _u0_u4_U527  ( .A(1'b1), .ZN(_u0_u4_pointer[2] ) );
INV_X4 _u0_u4_U525  ( .A(1'b1), .ZN(_u0_u4_pointer[1] ) );
INV_X4 _u0_u4_U523  ( .A(1'b1), .ZN(_u0_u4_pointer[0] ) );
INV_X4 _u0_u4_U521  ( .A(1'b1), .ZN(_u0_u4_pointer_s[31] ) );
INV_X4 _u0_u4_U519  ( .A(1'b1), .ZN(_u0_u4_pointer_s[30] ) );
INV_X4 _u0_u4_U517  ( .A(1'b1), .ZN(_u0_u4_pointer_s[29] ) );
INV_X4 _u0_u4_U515  ( .A(1'b1), .ZN(_u0_u4_pointer_s[28] ) );
INV_X4 _u0_u4_U513  ( .A(1'b1), .ZN(_u0_u4_pointer_s[27] ) );
INV_X4 _u0_u4_U511  ( .A(1'b1), .ZN(_u0_u4_pointer_s[26] ) );
INV_X4 _u0_u4_U509  ( .A(1'b1), .ZN(_u0_u4_pointer_s[25] ) );
INV_X4 _u0_u4_U507  ( .A(1'b1), .ZN(_u0_u4_pointer_s[24] ) );
INV_X4 _u0_u4_U505  ( .A(1'b1), .ZN(_u0_u4_pointer_s[23] ) );
INV_X4 _u0_u4_U503  ( .A(1'b1), .ZN(_u0_u4_pointer_s[22] ) );
INV_X4 _u0_u4_U501  ( .A(1'b1), .ZN(_u0_u4_pointer_s[21] ) );
INV_X4 _u0_u4_U499  ( .A(1'b1), .ZN(_u0_u4_pointer_s[20] ) );
INV_X4 _u0_u4_U497  ( .A(1'b1), .ZN(_u0_u4_pointer_s[19] ) );
INV_X4 _u0_u4_U495  ( .A(1'b1), .ZN(_u0_u4_pointer_s[18] ) );
INV_X4 _u0_u4_U493  ( .A(1'b1), .ZN(_u0_u4_pointer_s[17] ) );
INV_X4 _u0_u4_U491  ( .A(1'b1), .ZN(_u0_u4_pointer_s[16] ) );
INV_X4 _u0_u4_U489  ( .A(1'b1), .ZN(_u0_u4_pointer_s[15] ) );
INV_X4 _u0_u4_U487  ( .A(1'b1), .ZN(_u0_u4_pointer_s[14] ) );
INV_X4 _u0_u4_U485  ( .A(1'b1), .ZN(_u0_u4_pointer_s[13] ) );
INV_X4 _u0_u4_U483  ( .A(1'b1), .ZN(_u0_u4_pointer_s[12] ) );
INV_X4 _u0_u4_U481  ( .A(1'b1), .ZN(_u0_u4_pointer_s[11] ) );
INV_X4 _u0_u4_U479  ( .A(1'b1), .ZN(_u0_u4_pointer_s[10] ) );
INV_X4 _u0_u4_U477  ( .A(1'b1), .ZN(_u0_u4_pointer_s[9] ) );
INV_X4 _u0_u4_U475  ( .A(1'b1), .ZN(_u0_u4_pointer_s[8] ) );
INV_X4 _u0_u4_U473  ( .A(1'b1), .ZN(_u0_u4_pointer_s[7] ) );
INV_X4 _u0_u4_U471  ( .A(1'b1), .ZN(_u0_u4_pointer_s[6] ) );
INV_X4 _u0_u4_U469  ( .A(1'b1), .ZN(_u0_u4_pointer_s[5] ) );
INV_X4 _u0_u4_U467  ( .A(1'b1), .ZN(_u0_u4_pointer_s[4] ) );
INV_X4 _u0_u4_U465  ( .A(1'b1), .ZN(_u0_u4_pointer_s[3] ) );
INV_X4 _u0_u4_U463  ( .A(1'b1), .ZN(_u0_u4_pointer_s[2] ) );
INV_X4 _u0_u4_U461  ( .A(1'b1), .ZN(_u0_u4_pointer_s[1] ) );
INV_X4 _u0_u4_U459  ( .A(1'b1), .ZN(_u0_u4_pointer_s[0] ) );
INV_X4 _u0_u4_U457  ( .A(1'b1), .ZN(_u0_u4_ch_csr[31] ) );
INV_X4 _u0_u4_U455  ( .A(1'b1), .ZN(_u0_u4_ch_csr[30] ) );
INV_X4 _u0_u4_U453  ( .A(1'b1), .ZN(_u0_u4_ch_csr[29] ) );
INV_X4 _u0_u4_U451  ( .A(1'b1), .ZN(_u0_u4_ch_csr[28] ) );
INV_X4 _u0_u4_U449  ( .A(1'b1), .ZN(_u0_u4_ch_csr[27] ) );
INV_X4 _u0_u4_U447  ( .A(1'b1), .ZN(_u0_u4_ch_csr[26] ) );
INV_X4 _u0_u4_U445  ( .A(1'b1), .ZN(_u0_u4_ch_csr[25] ) );
INV_X4 _u0_u4_U443  ( .A(1'b1), .ZN(_u0_u4_ch_csr[24] ) );
INV_X4 _u0_u4_U441  ( .A(1'b1), .ZN(_u0_u4_ch_csr[23] ) );
INV_X4 _u0_u4_U439  ( .A(1'b1), .ZN(_u0_u4_ch_csr[22] ) );
INV_X4 _u0_u4_U437  ( .A(1'b1), .ZN(_u0_u4_ch_csr[21] ) );
INV_X4 _u0_u4_U435  ( .A(1'b1), .ZN(_u0_u4_ch_csr[20] ) );
INV_X4 _u0_u4_U433  ( .A(1'b1), .ZN(_u0_u4_ch_csr[19] ) );
INV_X4 _u0_u4_U431  ( .A(1'b1), .ZN(_u0_u4_ch_csr[18] ) );
INV_X4 _u0_u4_U429  ( .A(1'b1), .ZN(_u0_u4_ch_csr[17] ) );
INV_X4 _u0_u4_U427  ( .A(1'b1), .ZN(_u0_u4_ch_csr[16] ) );
INV_X4 _u0_u4_U425  ( .A(1'b1), .ZN(_u0_u4_ch_csr[15] ) );
INV_X4 _u0_u4_U423  ( .A(1'b1), .ZN(_u0_u4_ch_csr[14] ) );
INV_X4 _u0_u4_U421  ( .A(1'b1), .ZN(_u0_u4_ch_csr[13] ) );
INV_X4 _u0_u4_U419  ( .A(1'b1), .ZN(_u0_u4_ch_csr[12] ) );
INV_X4 _u0_u4_U417  ( .A(1'b1), .ZN(_u0_u4_ch_csr[11] ) );
INV_X4 _u0_u4_U415  ( .A(1'b1), .ZN(_u0_u4_ch_csr[10] ) );
INV_X4 _u0_u4_U413  ( .A(1'b1), .ZN(_u0_u4_ch_csr[9] ) );
INV_X4 _u0_u4_U411  ( .A(1'b1), .ZN(_u0_u4_ch_csr[8] ) );
INV_X4 _u0_u4_U409  ( .A(1'b1), .ZN(_u0_u4_ch_csr[7] ) );
INV_X4 _u0_u4_U407  ( .A(1'b1), .ZN(_u0_u4_ch_csr[6] ) );
INV_X4 _u0_u4_U405  ( .A(1'b1), .ZN(_u0_u4_ch_csr[5] ) );
INV_X4 _u0_u4_U403  ( .A(1'b1), .ZN(_u0_u4_ch_csr[4] ) );
INV_X4 _u0_u4_U401  ( .A(1'b1), .ZN(_u0_u4_ch_csr[3] ) );
INV_X4 _u0_u4_U399  ( .A(1'b1), .ZN(_u0_u4_ch_csr[2] ) );
INV_X4 _u0_u4_U397  ( .A(1'b1), .ZN(_u0_u4_ch_csr[1] ) );
INV_X4 _u0_u4_U395  ( .A(1'b1), .ZN(_u0_u4_ch_csr[0] ) );
INV_X4 _u0_u4_U393  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[31] ) );
INV_X4 _u0_u4_U391  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[30] ) );
INV_X4 _u0_u4_U389  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[29] ) );
INV_X4 _u0_u4_U387  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[28] ) );
INV_X4 _u0_u4_U385  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[27] ) );
INV_X4 _u0_u4_U383  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[26] ) );
INV_X4 _u0_u4_U381  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[25] ) );
INV_X4 _u0_u4_U379  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[24] ) );
INV_X4 _u0_u4_U377  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[23] ) );
INV_X4 _u0_u4_U375  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[22] ) );
INV_X4 _u0_u4_U373  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[21] ) );
INV_X4 _u0_u4_U371  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[20] ) );
INV_X4 _u0_u4_U369  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[19] ) );
INV_X4 _u0_u4_U367  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[18] ) );
INV_X4 _u0_u4_U365  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[17] ) );
INV_X4 _u0_u4_U363  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[16] ) );
INV_X4 _u0_u4_U361  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[15] ) );
INV_X4 _u0_u4_U359  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[14] ) );
INV_X4 _u0_u4_U357  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[13] ) );
INV_X4 _u0_u4_U355  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[12] ) );
INV_X4 _u0_u4_U353  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[11] ) );
INV_X4 _u0_u4_U351  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[10] ) );
INV_X4 _u0_u4_U349  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[9] ) );
INV_X4 _u0_u4_U347  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[8] ) );
INV_X4 _u0_u4_U345  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[7] ) );
INV_X4 _u0_u4_U343  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[6] ) );
INV_X4 _u0_u4_U341  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[5] ) );
INV_X4 _u0_u4_U339  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[4] ) );
INV_X4 _u0_u4_U337  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[3] ) );
INV_X4 _u0_u4_U335  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[2] ) );
INV_X4 _u0_u4_U333  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[1] ) );
INV_X4 _u0_u4_U331  ( .A(1'b1), .ZN(_u0_u4_ch_txsz[0] ) );
INV_X4 _u0_u4_U329  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[31] ) );
INV_X4 _u0_u4_U327  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[30] ) );
INV_X4 _u0_u4_U325  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[29] ) );
INV_X4 _u0_u4_U323  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[28] ) );
INV_X4 _u0_u4_U321  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[27] ) );
INV_X4 _u0_u4_U319  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[26] ) );
INV_X4 _u0_u4_U317  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[25] ) );
INV_X4 _u0_u4_U315  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[24] ) );
INV_X4 _u0_u4_U313  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[23] ) );
INV_X4 _u0_u4_U311  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[22] ) );
INV_X4 _u0_u4_U309  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[21] ) );
INV_X4 _u0_u4_U307  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[20] ) );
INV_X4 _u0_u4_U305  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[19] ) );
INV_X4 _u0_u4_U303  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[18] ) );
INV_X4 _u0_u4_U301  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[17] ) );
INV_X4 _u0_u4_U299  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[16] ) );
INV_X4 _u0_u4_U297  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[15] ) );
INV_X4 _u0_u4_U295  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[14] ) );
INV_X4 _u0_u4_U293  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[13] ) );
INV_X4 _u0_u4_U291  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[12] ) );
INV_X4 _u0_u4_U289  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[11] ) );
INV_X4 _u0_u4_U287  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[10] ) );
INV_X4 _u0_u4_U285  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[9] ) );
INV_X4 _u0_u4_U283  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[8] ) );
INV_X4 _u0_u4_U281  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[7] ) );
INV_X4 _u0_u4_U279  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[6] ) );
INV_X4 _u0_u4_U277  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[5] ) );
INV_X4 _u0_u4_U275  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[4] ) );
INV_X4 _u0_u4_U273  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[3] ) );
INV_X4 _u0_u4_U271  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[2] ) );
INV_X4 _u0_u4_U269  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[1] ) );
INV_X4 _u0_u4_U267  ( .A(1'b1), .ZN(_u0_u4_ch_adr0[0] ) );
INV_X4 _u0_u4_U265  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[31] ) );
INV_X4 _u0_u4_U263  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[30] ) );
INV_X4 _u0_u4_U261  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[29] ) );
INV_X4 _u0_u4_U259  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[28] ) );
INV_X4 _u0_u4_U257  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[27] ) );
INV_X4 _u0_u4_U255  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[26] ) );
INV_X4 _u0_u4_U253  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[25] ) );
INV_X4 _u0_u4_U251  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[24] ) );
INV_X4 _u0_u4_U249  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[23] ) );
INV_X4 _u0_u4_U247  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[22] ) );
INV_X4 _u0_u4_U245  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[21] ) );
INV_X4 _u0_u4_U243  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[20] ) );
INV_X4 _u0_u4_U241  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[19] ) );
INV_X4 _u0_u4_U239  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[18] ) );
INV_X4 _u0_u4_U237  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[17] ) );
INV_X4 _u0_u4_U235  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[16] ) );
INV_X4 _u0_u4_U233  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[15] ) );
INV_X4 _u0_u4_U231  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[14] ) );
INV_X4 _u0_u4_U229  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[13] ) );
INV_X4 _u0_u4_U227  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[12] ) );
INV_X4 _u0_u4_U225  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[11] ) );
INV_X4 _u0_u4_U223  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[10] ) );
INV_X4 _u0_u4_U221  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[9] ) );
INV_X4 _u0_u4_U219  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[8] ) );
INV_X4 _u0_u4_U217  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[7] ) );
INV_X4 _u0_u4_U215  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[6] ) );
INV_X4 _u0_u4_U213  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[5] ) );
INV_X4 _u0_u4_U211  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[4] ) );
INV_X4 _u0_u4_U209  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[3] ) );
INV_X4 _u0_u4_U207  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[2] ) );
INV_X4 _u0_u4_U205  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[1] ) );
INV_X4 _u0_u4_U203  ( .A(1'b1), .ZN(_u0_u4_ch_adr1[0] ) );
INV_X4 _u0_u4_U201  ( .A(1'b0), .ZN(_u0_u4_ch_am0[31] ) );
INV_X4 _u0_u4_U199  ( .A(1'b0), .ZN(_u0_u4_ch_am0[30] ) );
INV_X4 _u0_u4_U197  ( .A(1'b0), .ZN(_u0_u4_ch_am0[29] ) );
INV_X4 _u0_u4_U195  ( .A(1'b0), .ZN(_u0_u4_ch_am0[28] ) );
INV_X4 _u0_u4_U193  ( .A(1'b0), .ZN(_u0_u4_ch_am0[27] ) );
INV_X4 _u0_u4_U191  ( .A(1'b0), .ZN(_u0_u4_ch_am0[26] ) );
INV_X4 _u0_u4_U189  ( .A(1'b0), .ZN(_u0_u4_ch_am0[25] ) );
INV_X4 _u0_u4_U187  ( .A(1'b0), .ZN(_u0_u4_ch_am0[24] ) );
INV_X4 _u0_u4_U185  ( .A(1'b0), .ZN(_u0_u4_ch_am0[23] ) );
INV_X4 _u0_u4_U183  ( .A(1'b0), .ZN(_u0_u4_ch_am0[22] ) );
INV_X4 _u0_u4_U181  ( .A(1'b0), .ZN(_u0_u4_ch_am0[21] ) );
INV_X4 _u0_u4_U179  ( .A(1'b0), .ZN(_u0_u4_ch_am0[20] ) );
INV_X4 _u0_u4_U177  ( .A(1'b0), .ZN(_u0_u4_ch_am0[19] ) );
INV_X4 _u0_u4_U175  ( .A(1'b0), .ZN(_u0_u4_ch_am0[18] ) );
INV_X4 _u0_u4_U173  ( .A(1'b0), .ZN(_u0_u4_ch_am0[17] ) );
INV_X4 _u0_u4_U171  ( .A(1'b0), .ZN(_u0_u4_ch_am0[16] ) );
INV_X4 _u0_u4_U169  ( .A(1'b0), .ZN(_u0_u4_ch_am0[15] ) );
INV_X4 _u0_u4_U167  ( .A(1'b0), .ZN(_u0_u4_ch_am0[14] ) );
INV_X4 _u0_u4_U165  ( .A(1'b0), .ZN(_u0_u4_ch_am0[13] ) );
INV_X4 _u0_u4_U163  ( .A(1'b0), .ZN(_u0_u4_ch_am0[12] ) );
INV_X4 _u0_u4_U161  ( .A(1'b0), .ZN(_u0_u4_ch_am0[11] ) );
INV_X4 _u0_u4_U159  ( .A(1'b0), .ZN(_u0_u4_ch_am0[10] ) );
INV_X4 _u0_u4_U157  ( .A(1'b0), .ZN(_u0_u4_ch_am0[9] ) );
INV_X4 _u0_u4_U155  ( .A(1'b0), .ZN(_u0_u4_ch_am0[8] ) );
INV_X4 _u0_u4_U153  ( .A(1'b0), .ZN(_u0_u4_ch_am0[7] ) );
INV_X4 _u0_u4_U151  ( .A(1'b0), .ZN(_u0_u4_ch_am0[6] ) );
INV_X4 _u0_u4_U149  ( .A(1'b0), .ZN(_u0_u4_ch_am0[5] ) );
INV_X4 _u0_u4_U147  ( .A(1'b0), .ZN(_u0_u4_ch_am0[4] ) );
INV_X4 _u0_u4_U145  ( .A(1'b1), .ZN(_u0_u4_ch_am0[3] ) );
INV_X4 _u0_u4_U143  ( .A(1'b1), .ZN(_u0_u4_ch_am0[2] ) );
INV_X4 _u0_u4_U141  ( .A(1'b1), .ZN(_u0_u4_ch_am0[1] ) );
INV_X4 _u0_u4_U139  ( .A(1'b1), .ZN(_u0_u4_ch_am0[0] ) );
INV_X4 _u0_u4_U137  ( .A(1'b0), .ZN(_u0_u4_ch_am1[31] ) );
INV_X4 _u0_u4_U135  ( .A(1'b0), .ZN(_u0_u4_ch_am1[30] ) );
INV_X4 _u0_u4_U133  ( .A(1'b0), .ZN(_u0_u4_ch_am1[29] ) );
INV_X4 _u0_u4_U131  ( .A(1'b0), .ZN(_u0_u4_ch_am1[28] ) );
INV_X4 _u0_u4_U129  ( .A(1'b0), .ZN(_u0_u4_ch_am1[27] ) );
INV_X4 _u0_u4_U127  ( .A(1'b0), .ZN(_u0_u4_ch_am1[26] ) );
INV_X4 _u0_u4_U125  ( .A(1'b0), .ZN(_u0_u4_ch_am1[25] ) );
INV_X4 _u0_u4_U123  ( .A(1'b0), .ZN(_u0_u4_ch_am1[24] ) );
INV_X4 _u0_u4_U121  ( .A(1'b0), .ZN(_u0_u4_ch_am1[23] ) );
INV_X4 _u0_u4_U119  ( .A(1'b0), .ZN(_u0_u4_ch_am1[22] ) );
INV_X4 _u0_u4_U117  ( .A(1'b0), .ZN(_u0_u4_ch_am1[21] ) );
INV_X4 _u0_u4_U115  ( .A(1'b0), .ZN(_u0_u4_ch_am1[20] ) );
INV_X4 _u0_u4_U113  ( .A(1'b0), .ZN(_u0_u4_ch_am1[19] ) );
INV_X4 _u0_u4_U111  ( .A(1'b0), .ZN(_u0_u4_ch_am1[18] ) );
INV_X4 _u0_u4_U109  ( .A(1'b0), .ZN(_u0_u4_ch_am1[17] ) );
INV_X4 _u0_u4_U107  ( .A(1'b0), .ZN(_u0_u4_ch_am1[16] ) );
INV_X4 _u0_u4_U105  ( .A(1'b0), .ZN(_u0_u4_ch_am1[15] ) );
INV_X4 _u0_u4_U103  ( .A(1'b0), .ZN(_u0_u4_ch_am1[14] ) );
INV_X4 _u0_u4_U101  ( .A(1'b0), .ZN(_u0_u4_ch_am1[13] ) );
INV_X4 _u0_u4_U99  ( .A(1'b0), .ZN(_u0_u4_ch_am1[12] ) );
INV_X4 _u0_u4_U97  ( .A(1'b0), .ZN(_u0_u4_ch_am1[11] ) );
INV_X4 _u0_u4_U95  ( .A(1'b0), .ZN(_u0_u4_ch_am1[10] ) );
INV_X4 _u0_u4_U93  ( .A(1'b0), .ZN(_u0_u4_ch_am1[9] ) );
INV_X4 _u0_u4_U91  ( .A(1'b0), .ZN(_u0_u4_ch_am1[8] ) );
INV_X4 _u0_u4_U89  ( .A(1'b0), .ZN(_u0_u4_ch_am1[7] ) );
INV_X4 _u0_u4_U87  ( .A(1'b0), .ZN(_u0_u4_ch_am1[6] ) );
INV_X4 _u0_u4_U85  ( .A(1'b0), .ZN(_u0_u4_ch_am1[5] ) );
INV_X4 _u0_u4_U83  ( .A(1'b0), .ZN(_u0_u4_ch_am1[4] ) );
INV_X4 _u0_u4_U81  ( .A(1'b1), .ZN(_u0_u4_ch_am1[3] ) );
INV_X4 _u0_u4_U79  ( .A(1'b1), .ZN(_u0_u4_ch_am1[2] ) );
INV_X4 _u0_u4_U77  ( .A(1'b1), .ZN(_u0_u4_ch_am1[1] ) );
INV_X4 _u0_u4_U75  ( .A(1'b1), .ZN(_u0_u4_ch_am1[0] ) );
INV_X4 _u0_u4_U73  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[31] ) );
INV_X4 _u0_u4_U71  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[30] ) );
INV_X4 _u0_u4_U69  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[29] ) );
INV_X4 _u0_u4_U67  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[28] ) );
INV_X4 _u0_u4_U65  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[27] ) );
INV_X4 _u0_u4_U63  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[26] ) );
INV_X4 _u0_u4_U61  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[25] ) );
INV_X4 _u0_u4_U59  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[24] ) );
INV_X4 _u0_u4_U57  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[23] ) );
INV_X4 _u0_u4_U55  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[22] ) );
INV_X4 _u0_u4_U53  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[21] ) );
INV_X4 _u0_u4_U51  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[20] ) );
INV_X4 _u0_u4_U49  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[19] ) );
INV_X4 _u0_u4_U47  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[18] ) );
INV_X4 _u0_u4_U45  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[17] ) );
INV_X4 _u0_u4_U43  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[16] ) );
INV_X4 _u0_u4_U41  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[15] ) );
INV_X4 _u0_u4_U39  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[14] ) );
INV_X4 _u0_u4_U37  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[13] ) );
INV_X4 _u0_u4_U35  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[12] ) );
INV_X4 _u0_u4_U33  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[11] ) );
INV_X4 _u0_u4_U31  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[10] ) );
INV_X4 _u0_u4_U29  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[9] ) );
INV_X4 _u0_u4_U27  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[8] ) );
INV_X4 _u0_u4_U25  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[7] ) );
INV_X4 _u0_u4_U23  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[6] ) );
INV_X4 _u0_u4_U21  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[5] ) );
INV_X4 _u0_u4_U19  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[4] ) );
INV_X4 _u0_u4_U17  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[3] ) );
INV_X4 _u0_u4_U15  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[2] ) );
INV_X4 _u0_u4_U13  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[1] ) );
INV_X4 _u0_u4_U11  ( .A(1'b1), .ZN(_u0_u4_sw_pointer[0] ) );
INV_X4 _u0_u4_U9  ( .A(1'b1), .ZN(_u0_u4_ch_stop ) );
INV_X4 _u0_u4_U7  ( .A(1'b1), .ZN(_u0_u4_ch_dis ) );
INV_X4 _u0_u4_U5  ( .A(1'b1), .ZN(_u0_u4_int ) );
INV_X4 _u0_u5_U585  ( .A(1'b1), .ZN(_u0_u5_pointer[31] ) );
INV_X4 _u0_u5_U583  ( .A(1'b1), .ZN(_u0_u5_pointer[30] ) );
INV_X4 _u0_u5_U581  ( .A(1'b1), .ZN(_u0_u5_pointer[29] ) );
INV_X4 _u0_u5_U579  ( .A(1'b1), .ZN(_u0_u5_pointer[28] ) );
INV_X4 _u0_u5_U577  ( .A(1'b1), .ZN(_u0_u5_pointer[27] ) );
INV_X4 _u0_u5_U575  ( .A(1'b1), .ZN(_u0_u5_pointer[26] ) );
INV_X4 _u0_u5_U573  ( .A(1'b1), .ZN(_u0_u5_pointer[25] ) );
INV_X4 _u0_u5_U571  ( .A(1'b1), .ZN(_u0_u5_pointer[24] ) );
INV_X4 _u0_u5_U569  ( .A(1'b1), .ZN(_u0_u5_pointer[23] ) );
INV_X4 _u0_u5_U567  ( .A(1'b1), .ZN(_u0_u5_pointer[22] ) );
INV_X4 _u0_u5_U565  ( .A(1'b1), .ZN(_u0_u5_pointer[21] ) );
INV_X4 _u0_u5_U563  ( .A(1'b1), .ZN(_u0_u5_pointer[20] ) );
INV_X4 _u0_u5_U561  ( .A(1'b1), .ZN(_u0_u5_pointer[19] ) );
INV_X4 _u0_u5_U559  ( .A(1'b1), .ZN(_u0_u5_pointer[18] ) );
INV_X4 _u0_u5_U557  ( .A(1'b1), .ZN(_u0_u5_pointer[17] ) );
INV_X4 _u0_u5_U555  ( .A(1'b1), .ZN(_u0_u5_pointer[16] ) );
INV_X4 _u0_u5_U553  ( .A(1'b1), .ZN(_u0_u5_pointer[15] ) );
INV_X4 _u0_u5_U551  ( .A(1'b1), .ZN(_u0_u5_pointer[14] ) );
INV_X4 _u0_u5_U549  ( .A(1'b1), .ZN(_u0_u5_pointer[13] ) );
INV_X4 _u0_u5_U547  ( .A(1'b1), .ZN(_u0_u5_pointer[12] ) );
INV_X4 _u0_u5_U545  ( .A(1'b1), .ZN(_u0_u5_pointer[11] ) );
INV_X4 _u0_u5_U543  ( .A(1'b1), .ZN(_u0_u5_pointer[10] ) );
INV_X4 _u0_u5_U541  ( .A(1'b1), .ZN(_u0_u5_pointer[9] ) );
INV_X4 _u0_u5_U539  ( .A(1'b1), .ZN(_u0_u5_pointer[8] ) );
INV_X4 _u0_u5_U537  ( .A(1'b1), .ZN(_u0_u5_pointer[7] ) );
INV_X4 _u0_u5_U535  ( .A(1'b1), .ZN(_u0_u5_pointer[6] ) );
INV_X4 _u0_u5_U533  ( .A(1'b1), .ZN(_u0_u5_pointer[5] ) );
INV_X4 _u0_u5_U531  ( .A(1'b1), .ZN(_u0_u5_pointer[4] ) );
INV_X4 _u0_u5_U529  ( .A(1'b1), .ZN(_u0_u5_pointer[3] ) );
INV_X4 _u0_u5_U527  ( .A(1'b1), .ZN(_u0_u5_pointer[2] ) );
INV_X4 _u0_u5_U525  ( .A(1'b1), .ZN(_u0_u5_pointer[1] ) );
INV_X4 _u0_u5_U523  ( .A(1'b1), .ZN(_u0_u5_pointer[0] ) );
INV_X4 _u0_u5_U521  ( .A(1'b1), .ZN(_u0_u5_pointer_s[31] ) );
INV_X4 _u0_u5_U519  ( .A(1'b1), .ZN(_u0_u5_pointer_s[30] ) );
INV_X4 _u0_u5_U517  ( .A(1'b1), .ZN(_u0_u5_pointer_s[29] ) );
INV_X4 _u0_u5_U515  ( .A(1'b1), .ZN(_u0_u5_pointer_s[28] ) );
INV_X4 _u0_u5_U513  ( .A(1'b1), .ZN(_u0_u5_pointer_s[27] ) );
INV_X4 _u0_u5_U511  ( .A(1'b1), .ZN(_u0_u5_pointer_s[26] ) );
INV_X4 _u0_u5_U509  ( .A(1'b1), .ZN(_u0_u5_pointer_s[25] ) );
INV_X4 _u0_u5_U507  ( .A(1'b1), .ZN(_u0_u5_pointer_s[24] ) );
INV_X4 _u0_u5_U505  ( .A(1'b1), .ZN(_u0_u5_pointer_s[23] ) );
INV_X4 _u0_u5_U503  ( .A(1'b1), .ZN(_u0_u5_pointer_s[22] ) );
INV_X4 _u0_u5_U501  ( .A(1'b1), .ZN(_u0_u5_pointer_s[21] ) );
INV_X4 _u0_u5_U499  ( .A(1'b1), .ZN(_u0_u5_pointer_s[20] ) );
INV_X4 _u0_u5_U497  ( .A(1'b1), .ZN(_u0_u5_pointer_s[19] ) );
INV_X4 _u0_u5_U495  ( .A(1'b1), .ZN(_u0_u5_pointer_s[18] ) );
INV_X4 _u0_u5_U493  ( .A(1'b1), .ZN(_u0_u5_pointer_s[17] ) );
INV_X4 _u0_u5_U491  ( .A(1'b1), .ZN(_u0_u5_pointer_s[16] ) );
INV_X4 _u0_u5_U489  ( .A(1'b1), .ZN(_u0_u5_pointer_s[15] ) );
INV_X4 _u0_u5_U487  ( .A(1'b1), .ZN(_u0_u5_pointer_s[14] ) );
INV_X4 _u0_u5_U485  ( .A(1'b1), .ZN(_u0_u5_pointer_s[13] ) );
INV_X4 _u0_u5_U483  ( .A(1'b1), .ZN(_u0_u5_pointer_s[12] ) );
INV_X4 _u0_u5_U481  ( .A(1'b1), .ZN(_u0_u5_pointer_s[11] ) );
INV_X4 _u0_u5_U479  ( .A(1'b1), .ZN(_u0_u5_pointer_s[10] ) );
INV_X4 _u0_u5_U477  ( .A(1'b1), .ZN(_u0_u5_pointer_s[9] ) );
INV_X4 _u0_u5_U475  ( .A(1'b1), .ZN(_u0_u5_pointer_s[8] ) );
INV_X4 _u0_u5_U473  ( .A(1'b1), .ZN(_u0_u5_pointer_s[7] ) );
INV_X4 _u0_u5_U471  ( .A(1'b1), .ZN(_u0_u5_pointer_s[6] ) );
INV_X4 _u0_u5_U469  ( .A(1'b1), .ZN(_u0_u5_pointer_s[5] ) );
INV_X4 _u0_u5_U467  ( .A(1'b1), .ZN(_u0_u5_pointer_s[4] ) );
INV_X4 _u0_u5_U465  ( .A(1'b1), .ZN(_u0_u5_pointer_s[3] ) );
INV_X4 _u0_u5_U463  ( .A(1'b1), .ZN(_u0_u5_pointer_s[2] ) );
INV_X4 _u0_u5_U461  ( .A(1'b1), .ZN(_u0_u5_pointer_s[1] ) );
INV_X4 _u0_u5_U459  ( .A(1'b1), .ZN(_u0_u5_pointer_s[0] ) );
INV_X4 _u0_u5_U457  ( .A(1'b1), .ZN(_u0_u5_ch_csr[31] ) );
INV_X4 _u0_u5_U455  ( .A(1'b1), .ZN(_u0_u5_ch_csr[30] ) );
INV_X4 _u0_u5_U453  ( .A(1'b1), .ZN(_u0_u5_ch_csr[29] ) );
INV_X4 _u0_u5_U451  ( .A(1'b1), .ZN(_u0_u5_ch_csr[28] ) );
INV_X4 _u0_u5_U449  ( .A(1'b1), .ZN(_u0_u5_ch_csr[27] ) );
INV_X4 _u0_u5_U447  ( .A(1'b1), .ZN(_u0_u5_ch_csr[26] ) );
INV_X4 _u0_u5_U445  ( .A(1'b1), .ZN(_u0_u5_ch_csr[25] ) );
INV_X4 _u0_u5_U443  ( .A(1'b1), .ZN(_u0_u5_ch_csr[24] ) );
INV_X4 _u0_u5_U441  ( .A(1'b1), .ZN(_u0_u5_ch_csr[23] ) );
INV_X4 _u0_u5_U439  ( .A(1'b1), .ZN(_u0_u5_ch_csr[22] ) );
INV_X4 _u0_u5_U437  ( .A(1'b1), .ZN(_u0_u5_ch_csr[21] ) );
INV_X4 _u0_u5_U435  ( .A(1'b1), .ZN(_u0_u5_ch_csr[20] ) );
INV_X4 _u0_u5_U433  ( .A(1'b1), .ZN(_u0_u5_ch_csr[19] ) );
INV_X4 _u0_u5_U431  ( .A(1'b1), .ZN(_u0_u5_ch_csr[18] ) );
INV_X4 _u0_u5_U429  ( .A(1'b1), .ZN(_u0_u5_ch_csr[17] ) );
INV_X4 _u0_u5_U427  ( .A(1'b1), .ZN(_u0_u5_ch_csr[16] ) );
INV_X4 _u0_u5_U425  ( .A(1'b1), .ZN(_u0_u5_ch_csr[15] ) );
INV_X4 _u0_u5_U423  ( .A(1'b1), .ZN(_u0_u5_ch_csr[14] ) );
INV_X4 _u0_u5_U421  ( .A(1'b1), .ZN(_u0_u5_ch_csr[13] ) );
INV_X4 _u0_u5_U419  ( .A(1'b1), .ZN(_u0_u5_ch_csr[12] ) );
INV_X4 _u0_u5_U417  ( .A(1'b1), .ZN(_u0_u5_ch_csr[11] ) );
INV_X4 _u0_u5_U415  ( .A(1'b1), .ZN(_u0_u5_ch_csr[10] ) );
INV_X4 _u0_u5_U413  ( .A(1'b1), .ZN(_u0_u5_ch_csr[9] ) );
INV_X4 _u0_u5_U411  ( .A(1'b1), .ZN(_u0_u5_ch_csr[8] ) );
INV_X4 _u0_u5_U409  ( .A(1'b1), .ZN(_u0_u5_ch_csr[7] ) );
INV_X4 _u0_u5_U407  ( .A(1'b1), .ZN(_u0_u5_ch_csr[6] ) );
INV_X4 _u0_u5_U405  ( .A(1'b1), .ZN(_u0_u5_ch_csr[5] ) );
INV_X4 _u0_u5_U403  ( .A(1'b1), .ZN(_u0_u5_ch_csr[4] ) );
INV_X4 _u0_u5_U401  ( .A(1'b1), .ZN(_u0_u5_ch_csr[3] ) );
INV_X4 _u0_u5_U399  ( .A(1'b1), .ZN(_u0_u5_ch_csr[2] ) );
INV_X4 _u0_u5_U397  ( .A(1'b1), .ZN(_u0_u5_ch_csr[1] ) );
INV_X4 _u0_u5_U395  ( .A(1'b1), .ZN(_u0_u5_ch_csr[0] ) );
INV_X4 _u0_u5_U393  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[31] ) );
INV_X4 _u0_u5_U391  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[30] ) );
INV_X4 _u0_u5_U389  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[29] ) );
INV_X4 _u0_u5_U387  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[28] ) );
INV_X4 _u0_u5_U385  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[27] ) );
INV_X4 _u0_u5_U383  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[26] ) );
INV_X4 _u0_u5_U381  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[25] ) );
INV_X4 _u0_u5_U379  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[24] ) );
INV_X4 _u0_u5_U377  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[23] ) );
INV_X4 _u0_u5_U375  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[22] ) );
INV_X4 _u0_u5_U373  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[21] ) );
INV_X4 _u0_u5_U371  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[20] ) );
INV_X4 _u0_u5_U369  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[19] ) );
INV_X4 _u0_u5_U367  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[18] ) );
INV_X4 _u0_u5_U365  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[17] ) );
INV_X4 _u0_u5_U363  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[16] ) );
INV_X4 _u0_u5_U361  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[15] ) );
INV_X4 _u0_u5_U359  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[14] ) );
INV_X4 _u0_u5_U357  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[13] ) );
INV_X4 _u0_u5_U355  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[12] ) );
INV_X4 _u0_u5_U353  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[11] ) );
INV_X4 _u0_u5_U351  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[10] ) );
INV_X4 _u0_u5_U349  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[9] ) );
INV_X4 _u0_u5_U347  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[8] ) );
INV_X4 _u0_u5_U345  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[7] ) );
INV_X4 _u0_u5_U343  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[6] ) );
INV_X4 _u0_u5_U341  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[5] ) );
INV_X4 _u0_u5_U339  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[4] ) );
INV_X4 _u0_u5_U337  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[3] ) );
INV_X4 _u0_u5_U335  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[2] ) );
INV_X4 _u0_u5_U333  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[1] ) );
INV_X4 _u0_u5_U331  ( .A(1'b1), .ZN(_u0_u5_ch_txsz[0] ) );
INV_X4 _u0_u5_U329  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[31] ) );
INV_X4 _u0_u5_U327  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[30] ) );
INV_X4 _u0_u5_U325  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[29] ) );
INV_X4 _u0_u5_U323  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[28] ) );
INV_X4 _u0_u5_U321  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[27] ) );
INV_X4 _u0_u5_U319  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[26] ) );
INV_X4 _u0_u5_U317  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[25] ) );
INV_X4 _u0_u5_U315  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[24] ) );
INV_X4 _u0_u5_U313  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[23] ) );
INV_X4 _u0_u5_U311  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[22] ) );
INV_X4 _u0_u5_U309  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[21] ) );
INV_X4 _u0_u5_U307  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[20] ) );
INV_X4 _u0_u5_U305  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[19] ) );
INV_X4 _u0_u5_U303  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[18] ) );
INV_X4 _u0_u5_U301  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[17] ) );
INV_X4 _u0_u5_U299  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[16] ) );
INV_X4 _u0_u5_U297  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[15] ) );
INV_X4 _u0_u5_U295  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[14] ) );
INV_X4 _u0_u5_U293  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[13] ) );
INV_X4 _u0_u5_U291  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[12] ) );
INV_X4 _u0_u5_U289  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[11] ) );
INV_X4 _u0_u5_U287  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[10] ) );
INV_X4 _u0_u5_U285  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[9] ) );
INV_X4 _u0_u5_U283  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[8] ) );
INV_X4 _u0_u5_U281  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[7] ) );
INV_X4 _u0_u5_U279  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[6] ) );
INV_X4 _u0_u5_U277  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[5] ) );
INV_X4 _u0_u5_U275  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[4] ) );
INV_X4 _u0_u5_U273  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[3] ) );
INV_X4 _u0_u5_U271  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[2] ) );
INV_X4 _u0_u5_U269  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[1] ) );
INV_X4 _u0_u5_U267  ( .A(1'b1), .ZN(_u0_u5_ch_adr0[0] ) );
INV_X4 _u0_u5_U265  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[31] ) );
INV_X4 _u0_u5_U263  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[30] ) );
INV_X4 _u0_u5_U261  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[29] ) );
INV_X4 _u0_u5_U259  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[28] ) );
INV_X4 _u0_u5_U257  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[27] ) );
INV_X4 _u0_u5_U255  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[26] ) );
INV_X4 _u0_u5_U253  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[25] ) );
INV_X4 _u0_u5_U251  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[24] ) );
INV_X4 _u0_u5_U249  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[23] ) );
INV_X4 _u0_u5_U247  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[22] ) );
INV_X4 _u0_u5_U245  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[21] ) );
INV_X4 _u0_u5_U243  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[20] ) );
INV_X4 _u0_u5_U241  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[19] ) );
INV_X4 _u0_u5_U239  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[18] ) );
INV_X4 _u0_u5_U237  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[17] ) );
INV_X4 _u0_u5_U235  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[16] ) );
INV_X4 _u0_u5_U233  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[15] ) );
INV_X4 _u0_u5_U231  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[14] ) );
INV_X4 _u0_u5_U229  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[13] ) );
INV_X4 _u0_u5_U227  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[12] ) );
INV_X4 _u0_u5_U225  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[11] ) );
INV_X4 _u0_u5_U223  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[10] ) );
INV_X4 _u0_u5_U221  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[9] ) );
INV_X4 _u0_u5_U219  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[8] ) );
INV_X4 _u0_u5_U217  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[7] ) );
INV_X4 _u0_u5_U215  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[6] ) );
INV_X4 _u0_u5_U213  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[5] ) );
INV_X4 _u0_u5_U211  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[4] ) );
INV_X4 _u0_u5_U209  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[3] ) );
INV_X4 _u0_u5_U207  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[2] ) );
INV_X4 _u0_u5_U205  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[1] ) );
INV_X4 _u0_u5_U203  ( .A(1'b1), .ZN(_u0_u5_ch_adr1[0] ) );
INV_X4 _u0_u5_U201  ( .A(1'b0), .ZN(_u0_u5_ch_am0[31] ) );
INV_X4 _u0_u5_U199  ( .A(1'b0), .ZN(_u0_u5_ch_am0[30] ) );
INV_X4 _u0_u5_U197  ( .A(1'b0), .ZN(_u0_u5_ch_am0[29] ) );
INV_X4 _u0_u5_U195  ( .A(1'b0), .ZN(_u0_u5_ch_am0[28] ) );
INV_X4 _u0_u5_U193  ( .A(1'b0), .ZN(_u0_u5_ch_am0[27] ) );
INV_X4 _u0_u5_U191  ( .A(1'b0), .ZN(_u0_u5_ch_am0[26] ) );
INV_X4 _u0_u5_U189  ( .A(1'b0), .ZN(_u0_u5_ch_am0[25] ) );
INV_X4 _u0_u5_U187  ( .A(1'b0), .ZN(_u0_u5_ch_am0[24] ) );
INV_X4 _u0_u5_U185  ( .A(1'b0), .ZN(_u0_u5_ch_am0[23] ) );
INV_X4 _u0_u5_U183  ( .A(1'b0), .ZN(_u0_u5_ch_am0[22] ) );
INV_X4 _u0_u5_U181  ( .A(1'b0), .ZN(_u0_u5_ch_am0[21] ) );
INV_X4 _u0_u5_U179  ( .A(1'b0), .ZN(_u0_u5_ch_am0[20] ) );
INV_X4 _u0_u5_U177  ( .A(1'b0), .ZN(_u0_u5_ch_am0[19] ) );
INV_X4 _u0_u5_U175  ( .A(1'b0), .ZN(_u0_u5_ch_am0[18] ) );
INV_X4 _u0_u5_U173  ( .A(1'b0), .ZN(_u0_u5_ch_am0[17] ) );
INV_X4 _u0_u5_U171  ( .A(1'b0), .ZN(_u0_u5_ch_am0[16] ) );
INV_X4 _u0_u5_U169  ( .A(1'b0), .ZN(_u0_u5_ch_am0[15] ) );
INV_X4 _u0_u5_U167  ( .A(1'b0), .ZN(_u0_u5_ch_am0[14] ) );
INV_X4 _u0_u5_U165  ( .A(1'b0), .ZN(_u0_u5_ch_am0[13] ) );
INV_X4 _u0_u5_U163  ( .A(1'b0), .ZN(_u0_u5_ch_am0[12] ) );
INV_X4 _u0_u5_U161  ( .A(1'b0), .ZN(_u0_u5_ch_am0[11] ) );
INV_X4 _u0_u5_U159  ( .A(1'b0), .ZN(_u0_u5_ch_am0[10] ) );
INV_X4 _u0_u5_U157  ( .A(1'b0), .ZN(_u0_u5_ch_am0[9] ) );
INV_X4 _u0_u5_U155  ( .A(1'b0), .ZN(_u0_u5_ch_am0[8] ) );
INV_X4 _u0_u5_U153  ( .A(1'b0), .ZN(_u0_u5_ch_am0[7] ) );
INV_X4 _u0_u5_U151  ( .A(1'b0), .ZN(_u0_u5_ch_am0[6] ) );
INV_X4 _u0_u5_U149  ( .A(1'b0), .ZN(_u0_u5_ch_am0[5] ) );
INV_X4 _u0_u5_U147  ( .A(1'b0), .ZN(_u0_u5_ch_am0[4] ) );
INV_X4 _u0_u5_U145  ( .A(1'b1), .ZN(_u0_u5_ch_am0[3] ) );
INV_X4 _u0_u5_U143  ( .A(1'b1), .ZN(_u0_u5_ch_am0[2] ) );
INV_X4 _u0_u5_U141  ( .A(1'b1), .ZN(_u0_u5_ch_am0[1] ) );
INV_X4 _u0_u5_U139  ( .A(1'b1), .ZN(_u0_u5_ch_am0[0] ) );
INV_X4 _u0_u5_U137  ( .A(1'b0), .ZN(_u0_u5_ch_am1[31] ) );
INV_X4 _u0_u5_U135  ( .A(1'b0), .ZN(_u0_u5_ch_am1[30] ) );
INV_X4 _u0_u5_U133  ( .A(1'b0), .ZN(_u0_u5_ch_am1[29] ) );
INV_X4 _u0_u5_U131  ( .A(1'b0), .ZN(_u0_u5_ch_am1[28] ) );
INV_X4 _u0_u5_U129  ( .A(1'b0), .ZN(_u0_u5_ch_am1[27] ) );
INV_X4 _u0_u5_U127  ( .A(1'b0), .ZN(_u0_u5_ch_am1[26] ) );
INV_X4 _u0_u5_U125  ( .A(1'b0), .ZN(_u0_u5_ch_am1[25] ) );
INV_X4 _u0_u5_U123  ( .A(1'b0), .ZN(_u0_u5_ch_am1[24] ) );
INV_X4 _u0_u5_U121  ( .A(1'b0), .ZN(_u0_u5_ch_am1[23] ) );
INV_X4 _u0_u5_U119  ( .A(1'b0), .ZN(_u0_u5_ch_am1[22] ) );
INV_X4 _u0_u5_U117  ( .A(1'b0), .ZN(_u0_u5_ch_am1[21] ) );
INV_X4 _u0_u5_U115  ( .A(1'b0), .ZN(_u0_u5_ch_am1[20] ) );
INV_X4 _u0_u5_U113  ( .A(1'b0), .ZN(_u0_u5_ch_am1[19] ) );
INV_X4 _u0_u5_U111  ( .A(1'b0), .ZN(_u0_u5_ch_am1[18] ) );
INV_X4 _u0_u5_U109  ( .A(1'b0), .ZN(_u0_u5_ch_am1[17] ) );
INV_X4 _u0_u5_U107  ( .A(1'b0), .ZN(_u0_u5_ch_am1[16] ) );
INV_X4 _u0_u5_U105  ( .A(1'b0), .ZN(_u0_u5_ch_am1[15] ) );
INV_X4 _u0_u5_U103  ( .A(1'b0), .ZN(_u0_u5_ch_am1[14] ) );
INV_X4 _u0_u5_U101  ( .A(1'b0), .ZN(_u0_u5_ch_am1[13] ) );
INV_X4 _u0_u5_U99  ( .A(1'b0), .ZN(_u0_u5_ch_am1[12] ) );
INV_X4 _u0_u5_U97  ( .A(1'b0), .ZN(_u0_u5_ch_am1[11] ) );
INV_X4 _u0_u5_U95  ( .A(1'b0), .ZN(_u0_u5_ch_am1[10] ) );
INV_X4 _u0_u5_U93  ( .A(1'b0), .ZN(_u0_u5_ch_am1[9] ) );
INV_X4 _u0_u5_U91  ( .A(1'b0), .ZN(_u0_u5_ch_am1[8] ) );
INV_X4 _u0_u5_U89  ( .A(1'b0), .ZN(_u0_u5_ch_am1[7] ) );
INV_X4 _u0_u5_U87  ( .A(1'b0), .ZN(_u0_u5_ch_am1[6] ) );
INV_X4 _u0_u5_U85  ( .A(1'b0), .ZN(_u0_u5_ch_am1[5] ) );
INV_X4 _u0_u5_U83  ( .A(1'b0), .ZN(_u0_u5_ch_am1[4] ) );
INV_X4 _u0_u5_U81  ( .A(1'b1), .ZN(_u0_u5_ch_am1[3] ) );
INV_X4 _u0_u5_U79  ( .A(1'b1), .ZN(_u0_u5_ch_am1[2] ) );
INV_X4 _u0_u5_U77  ( .A(1'b1), .ZN(_u0_u5_ch_am1[1] ) );
INV_X4 _u0_u5_U75  ( .A(1'b1), .ZN(_u0_u5_ch_am1[0] ) );
INV_X4 _u0_u5_U73  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[31] ) );
INV_X4 _u0_u5_U71  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[30] ) );
INV_X4 _u0_u5_U69  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[29] ) );
INV_X4 _u0_u5_U67  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[28] ) );
INV_X4 _u0_u5_U65  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[27] ) );
INV_X4 _u0_u5_U63  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[26] ) );
INV_X4 _u0_u5_U61  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[25] ) );
INV_X4 _u0_u5_U59  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[24] ) );
INV_X4 _u0_u5_U57  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[23] ) );
INV_X4 _u0_u5_U55  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[22] ) );
INV_X4 _u0_u5_U53  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[21] ) );
INV_X4 _u0_u5_U51  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[20] ) );
INV_X4 _u0_u5_U49  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[19] ) );
INV_X4 _u0_u5_U47  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[18] ) );
INV_X4 _u0_u5_U45  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[17] ) );
INV_X4 _u0_u5_U43  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[16] ) );
INV_X4 _u0_u5_U41  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[15] ) );
INV_X4 _u0_u5_U39  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[14] ) );
INV_X4 _u0_u5_U37  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[13] ) );
INV_X4 _u0_u5_U35  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[12] ) );
INV_X4 _u0_u5_U33  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[11] ) );
INV_X4 _u0_u5_U31  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[10] ) );
INV_X4 _u0_u5_U29  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[9] ) );
INV_X4 _u0_u5_U27  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[8] ) );
INV_X4 _u0_u5_U25  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[7] ) );
INV_X4 _u0_u5_U23  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[6] ) );
INV_X4 _u0_u5_U21  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[5] ) );
INV_X4 _u0_u5_U19  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[4] ) );
INV_X4 _u0_u5_U17  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[3] ) );
INV_X4 _u0_u5_U15  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[2] ) );
INV_X4 _u0_u5_U13  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[1] ) );
INV_X4 _u0_u5_U11  ( .A(1'b1), .ZN(_u0_u5_sw_pointer[0] ) );
INV_X4 _u0_u5_U9  ( .A(1'b1), .ZN(_u0_u5_ch_stop ) );
INV_X4 _u0_u5_U7  ( .A(1'b1), .ZN(_u0_u5_ch_dis ) );
INV_X4 _u0_u5_U5  ( .A(1'b1), .ZN(_u0_u5_int ) );
INV_X4 _u0_u6_U585  ( .A(1'b1), .ZN(_u0_u6_pointer[31] ) );
INV_X4 _u0_u6_U583  ( .A(1'b1), .ZN(_u0_u6_pointer[30] ) );
INV_X4 _u0_u6_U581  ( .A(1'b1), .ZN(_u0_u6_pointer[29] ) );
INV_X4 _u0_u6_U579  ( .A(1'b1), .ZN(_u0_u6_pointer[28] ) );
INV_X4 _u0_u6_U577  ( .A(1'b1), .ZN(_u0_u6_pointer[27] ) );
INV_X4 _u0_u6_U575  ( .A(1'b1), .ZN(_u0_u6_pointer[26] ) );
INV_X4 _u0_u6_U573  ( .A(1'b1), .ZN(_u0_u6_pointer[25] ) );
INV_X4 _u0_u6_U571  ( .A(1'b1), .ZN(_u0_u6_pointer[24] ) );
INV_X4 _u0_u6_U569  ( .A(1'b1), .ZN(_u0_u6_pointer[23] ) );
INV_X4 _u0_u6_U567  ( .A(1'b1), .ZN(_u0_u6_pointer[22] ) );
INV_X4 _u0_u6_U565  ( .A(1'b1), .ZN(_u0_u6_pointer[21] ) );
INV_X4 _u0_u6_U563  ( .A(1'b1), .ZN(_u0_u6_pointer[20] ) );
INV_X4 _u0_u6_U561  ( .A(1'b1), .ZN(_u0_u6_pointer[19] ) );
INV_X4 _u0_u6_U559  ( .A(1'b1), .ZN(_u0_u6_pointer[18] ) );
INV_X4 _u0_u6_U557  ( .A(1'b1), .ZN(_u0_u6_pointer[17] ) );
INV_X4 _u0_u6_U555  ( .A(1'b1), .ZN(_u0_u6_pointer[16] ) );
INV_X4 _u0_u6_U553  ( .A(1'b1), .ZN(_u0_u6_pointer[15] ) );
INV_X4 _u0_u6_U551  ( .A(1'b1), .ZN(_u0_u6_pointer[14] ) );
INV_X4 _u0_u6_U549  ( .A(1'b1), .ZN(_u0_u6_pointer[13] ) );
INV_X4 _u0_u6_U547  ( .A(1'b1), .ZN(_u0_u6_pointer[12] ) );
INV_X4 _u0_u6_U545  ( .A(1'b1), .ZN(_u0_u6_pointer[11] ) );
INV_X4 _u0_u6_U543  ( .A(1'b1), .ZN(_u0_u6_pointer[10] ) );
INV_X4 _u0_u6_U541  ( .A(1'b1), .ZN(_u0_u6_pointer[9] ) );
INV_X4 _u0_u6_U539  ( .A(1'b1), .ZN(_u0_u6_pointer[8] ) );
INV_X4 _u0_u6_U537  ( .A(1'b1), .ZN(_u0_u6_pointer[7] ) );
INV_X4 _u0_u6_U535  ( .A(1'b1), .ZN(_u0_u6_pointer[6] ) );
INV_X4 _u0_u6_U533  ( .A(1'b1), .ZN(_u0_u6_pointer[5] ) );
INV_X4 _u0_u6_U531  ( .A(1'b1), .ZN(_u0_u6_pointer[4] ) );
INV_X4 _u0_u6_U529  ( .A(1'b1), .ZN(_u0_u6_pointer[3] ) );
INV_X4 _u0_u6_U527  ( .A(1'b1), .ZN(_u0_u6_pointer[2] ) );
INV_X4 _u0_u6_U525  ( .A(1'b1), .ZN(_u0_u6_pointer[1] ) );
INV_X4 _u0_u6_U523  ( .A(1'b1), .ZN(_u0_u6_pointer[0] ) );
INV_X4 _u0_u6_U521  ( .A(1'b1), .ZN(_u0_u6_pointer_s[31] ) );
INV_X4 _u0_u6_U519  ( .A(1'b1), .ZN(_u0_u6_pointer_s[30] ) );
INV_X4 _u0_u6_U517  ( .A(1'b1), .ZN(_u0_u6_pointer_s[29] ) );
INV_X4 _u0_u6_U515  ( .A(1'b1), .ZN(_u0_u6_pointer_s[28] ) );
INV_X4 _u0_u6_U513  ( .A(1'b1), .ZN(_u0_u6_pointer_s[27] ) );
INV_X4 _u0_u6_U511  ( .A(1'b1), .ZN(_u0_u6_pointer_s[26] ) );
INV_X4 _u0_u6_U509  ( .A(1'b1), .ZN(_u0_u6_pointer_s[25] ) );
INV_X4 _u0_u6_U507  ( .A(1'b1), .ZN(_u0_u6_pointer_s[24] ) );
INV_X4 _u0_u6_U505  ( .A(1'b1), .ZN(_u0_u6_pointer_s[23] ) );
INV_X4 _u0_u6_U503  ( .A(1'b1), .ZN(_u0_u6_pointer_s[22] ) );
INV_X4 _u0_u6_U501  ( .A(1'b1), .ZN(_u0_u6_pointer_s[21] ) );
INV_X4 _u0_u6_U499  ( .A(1'b1), .ZN(_u0_u6_pointer_s[20] ) );
INV_X4 _u0_u6_U497  ( .A(1'b1), .ZN(_u0_u6_pointer_s[19] ) );
INV_X4 _u0_u6_U495  ( .A(1'b1), .ZN(_u0_u6_pointer_s[18] ) );
INV_X4 _u0_u6_U493  ( .A(1'b1), .ZN(_u0_u6_pointer_s[17] ) );
INV_X4 _u0_u6_U491  ( .A(1'b1), .ZN(_u0_u6_pointer_s[16] ) );
INV_X4 _u0_u6_U489  ( .A(1'b1), .ZN(_u0_u6_pointer_s[15] ) );
INV_X4 _u0_u6_U487  ( .A(1'b1), .ZN(_u0_u6_pointer_s[14] ) );
INV_X4 _u0_u6_U485  ( .A(1'b1), .ZN(_u0_u6_pointer_s[13] ) );
INV_X4 _u0_u6_U483  ( .A(1'b1), .ZN(_u0_u6_pointer_s[12] ) );
INV_X4 _u0_u6_U481  ( .A(1'b1), .ZN(_u0_u6_pointer_s[11] ) );
INV_X4 _u0_u6_U479  ( .A(1'b1), .ZN(_u0_u6_pointer_s[10] ) );
INV_X4 _u0_u6_U477  ( .A(1'b1), .ZN(_u0_u6_pointer_s[9] ) );
INV_X4 _u0_u6_U475  ( .A(1'b1), .ZN(_u0_u6_pointer_s[8] ) );
INV_X4 _u0_u6_U473  ( .A(1'b1), .ZN(_u0_u6_pointer_s[7] ) );
INV_X4 _u0_u6_U471  ( .A(1'b1), .ZN(_u0_u6_pointer_s[6] ) );
INV_X4 _u0_u6_U469  ( .A(1'b1), .ZN(_u0_u6_pointer_s[5] ) );
INV_X4 _u0_u6_U467  ( .A(1'b1), .ZN(_u0_u6_pointer_s[4] ) );
INV_X4 _u0_u6_U465  ( .A(1'b1), .ZN(_u0_u6_pointer_s[3] ) );
INV_X4 _u0_u6_U463  ( .A(1'b1), .ZN(_u0_u6_pointer_s[2] ) );
INV_X4 _u0_u6_U461  ( .A(1'b1), .ZN(_u0_u6_pointer_s[1] ) );
INV_X4 _u0_u6_U459  ( .A(1'b1), .ZN(_u0_u6_pointer_s[0] ) );
INV_X4 _u0_u6_U457  ( .A(1'b1), .ZN(_u0_u6_ch_csr[31] ) );
INV_X4 _u0_u6_U455  ( .A(1'b1), .ZN(_u0_u6_ch_csr[30] ) );
INV_X4 _u0_u6_U453  ( .A(1'b1), .ZN(_u0_u6_ch_csr[29] ) );
INV_X4 _u0_u6_U451  ( .A(1'b1), .ZN(_u0_u6_ch_csr[28] ) );
INV_X4 _u0_u6_U449  ( .A(1'b1), .ZN(_u0_u6_ch_csr[27] ) );
INV_X4 _u0_u6_U447  ( .A(1'b1), .ZN(_u0_u6_ch_csr[26] ) );
INV_X4 _u0_u6_U445  ( .A(1'b1), .ZN(_u0_u6_ch_csr[25] ) );
INV_X4 _u0_u6_U443  ( .A(1'b1), .ZN(_u0_u6_ch_csr[24] ) );
INV_X4 _u0_u6_U441  ( .A(1'b1), .ZN(_u0_u6_ch_csr[23] ) );
INV_X4 _u0_u6_U439  ( .A(1'b1), .ZN(_u0_u6_ch_csr[22] ) );
INV_X4 _u0_u6_U437  ( .A(1'b1), .ZN(_u0_u6_ch_csr[21] ) );
INV_X4 _u0_u6_U435  ( .A(1'b1), .ZN(_u0_u6_ch_csr[20] ) );
INV_X4 _u0_u6_U433  ( .A(1'b1), .ZN(_u0_u6_ch_csr[19] ) );
INV_X4 _u0_u6_U431  ( .A(1'b1), .ZN(_u0_u6_ch_csr[18] ) );
INV_X4 _u0_u6_U429  ( .A(1'b1), .ZN(_u0_u6_ch_csr[17] ) );
INV_X4 _u0_u6_U427  ( .A(1'b1), .ZN(_u0_u6_ch_csr[16] ) );
INV_X4 _u0_u6_U425  ( .A(1'b1), .ZN(_u0_u6_ch_csr[15] ) );
INV_X4 _u0_u6_U423  ( .A(1'b1), .ZN(_u0_u6_ch_csr[14] ) );
INV_X4 _u0_u6_U421  ( .A(1'b1), .ZN(_u0_u6_ch_csr[13] ) );
INV_X4 _u0_u6_U419  ( .A(1'b1), .ZN(_u0_u6_ch_csr[12] ) );
INV_X4 _u0_u6_U417  ( .A(1'b1), .ZN(_u0_u6_ch_csr[11] ) );
INV_X4 _u0_u6_U415  ( .A(1'b1), .ZN(_u0_u6_ch_csr[10] ) );
INV_X4 _u0_u6_U413  ( .A(1'b1), .ZN(_u0_u6_ch_csr[9] ) );
INV_X4 _u0_u6_U411  ( .A(1'b1), .ZN(_u0_u6_ch_csr[8] ) );
INV_X4 _u0_u6_U409  ( .A(1'b1), .ZN(_u0_u6_ch_csr[7] ) );
INV_X4 _u0_u6_U407  ( .A(1'b1), .ZN(_u0_u6_ch_csr[6] ) );
INV_X4 _u0_u6_U405  ( .A(1'b1), .ZN(_u0_u6_ch_csr[5] ) );
INV_X4 _u0_u6_U403  ( .A(1'b1), .ZN(_u0_u6_ch_csr[4] ) );
INV_X4 _u0_u6_U401  ( .A(1'b1), .ZN(_u0_u6_ch_csr[3] ) );
INV_X4 _u0_u6_U399  ( .A(1'b1), .ZN(_u0_u6_ch_csr[2] ) );
INV_X4 _u0_u6_U397  ( .A(1'b1), .ZN(_u0_u6_ch_csr[1] ) );
INV_X4 _u0_u6_U395  ( .A(1'b1), .ZN(_u0_u6_ch_csr[0] ) );
INV_X4 _u0_u6_U393  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[31] ) );
INV_X4 _u0_u6_U391  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[30] ) );
INV_X4 _u0_u6_U389  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[29] ) );
INV_X4 _u0_u6_U387  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[28] ) );
INV_X4 _u0_u6_U385  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[27] ) );
INV_X4 _u0_u6_U383  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[26] ) );
INV_X4 _u0_u6_U381  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[25] ) );
INV_X4 _u0_u6_U379  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[24] ) );
INV_X4 _u0_u6_U377  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[23] ) );
INV_X4 _u0_u6_U375  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[22] ) );
INV_X4 _u0_u6_U373  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[21] ) );
INV_X4 _u0_u6_U371  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[20] ) );
INV_X4 _u0_u6_U369  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[19] ) );
INV_X4 _u0_u6_U367  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[18] ) );
INV_X4 _u0_u6_U365  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[17] ) );
INV_X4 _u0_u6_U363  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[16] ) );
INV_X4 _u0_u6_U361  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[15] ) );
INV_X4 _u0_u6_U359  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[14] ) );
INV_X4 _u0_u6_U357  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[13] ) );
INV_X4 _u0_u6_U355  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[12] ) );
INV_X4 _u0_u6_U353  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[11] ) );
INV_X4 _u0_u6_U351  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[10] ) );
INV_X4 _u0_u6_U349  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[9] ) );
INV_X4 _u0_u6_U347  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[8] ) );
INV_X4 _u0_u6_U345  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[7] ) );
INV_X4 _u0_u6_U343  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[6] ) );
INV_X4 _u0_u6_U341  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[5] ) );
INV_X4 _u0_u6_U339  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[4] ) );
INV_X4 _u0_u6_U337  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[3] ) );
INV_X4 _u0_u6_U335  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[2] ) );
INV_X4 _u0_u6_U333  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[1] ) );
INV_X4 _u0_u6_U331  ( .A(1'b1), .ZN(_u0_u6_ch_txsz[0] ) );
INV_X4 _u0_u6_U329  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[31] ) );
INV_X4 _u0_u6_U327  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[30] ) );
INV_X4 _u0_u6_U325  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[29] ) );
INV_X4 _u0_u6_U323  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[28] ) );
INV_X4 _u0_u6_U321  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[27] ) );
INV_X4 _u0_u6_U319  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[26] ) );
INV_X4 _u0_u6_U317  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[25] ) );
INV_X4 _u0_u6_U315  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[24] ) );
INV_X4 _u0_u6_U313  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[23] ) );
INV_X4 _u0_u6_U311  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[22] ) );
INV_X4 _u0_u6_U309  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[21] ) );
INV_X4 _u0_u6_U307  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[20] ) );
INV_X4 _u0_u6_U305  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[19] ) );
INV_X4 _u0_u6_U303  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[18] ) );
INV_X4 _u0_u6_U301  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[17] ) );
INV_X4 _u0_u6_U299  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[16] ) );
INV_X4 _u0_u6_U297  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[15] ) );
INV_X4 _u0_u6_U295  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[14] ) );
INV_X4 _u0_u6_U293  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[13] ) );
INV_X4 _u0_u6_U291  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[12] ) );
INV_X4 _u0_u6_U289  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[11] ) );
INV_X4 _u0_u6_U287  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[10] ) );
INV_X4 _u0_u6_U285  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[9] ) );
INV_X4 _u0_u6_U283  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[8] ) );
INV_X4 _u0_u6_U281  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[7] ) );
INV_X4 _u0_u6_U279  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[6] ) );
INV_X4 _u0_u6_U277  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[5] ) );
INV_X4 _u0_u6_U275  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[4] ) );
INV_X4 _u0_u6_U273  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[3] ) );
INV_X4 _u0_u6_U271  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[2] ) );
INV_X4 _u0_u6_U269  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[1] ) );
INV_X4 _u0_u6_U267  ( .A(1'b1), .ZN(_u0_u6_ch_adr0[0] ) );
INV_X4 _u0_u6_U265  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[31] ) );
INV_X4 _u0_u6_U263  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[30] ) );
INV_X4 _u0_u6_U261  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[29] ) );
INV_X4 _u0_u6_U259  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[28] ) );
INV_X4 _u0_u6_U257  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[27] ) );
INV_X4 _u0_u6_U255  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[26] ) );
INV_X4 _u0_u6_U253  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[25] ) );
INV_X4 _u0_u6_U251  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[24] ) );
INV_X4 _u0_u6_U249  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[23] ) );
INV_X4 _u0_u6_U247  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[22] ) );
INV_X4 _u0_u6_U245  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[21] ) );
INV_X4 _u0_u6_U243  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[20] ) );
INV_X4 _u0_u6_U241  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[19] ) );
INV_X4 _u0_u6_U239  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[18] ) );
INV_X4 _u0_u6_U237  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[17] ) );
INV_X4 _u0_u6_U235  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[16] ) );
INV_X4 _u0_u6_U233  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[15] ) );
INV_X4 _u0_u6_U231  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[14] ) );
INV_X4 _u0_u6_U229  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[13] ) );
INV_X4 _u0_u6_U227  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[12] ) );
INV_X4 _u0_u6_U225  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[11] ) );
INV_X4 _u0_u6_U223  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[10] ) );
INV_X4 _u0_u6_U221  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[9] ) );
INV_X4 _u0_u6_U219  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[8] ) );
INV_X4 _u0_u6_U217  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[7] ) );
INV_X4 _u0_u6_U215  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[6] ) );
INV_X4 _u0_u6_U213  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[5] ) );
INV_X4 _u0_u6_U211  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[4] ) );
INV_X4 _u0_u6_U209  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[3] ) );
INV_X4 _u0_u6_U207  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[2] ) );
INV_X4 _u0_u6_U205  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[1] ) );
INV_X4 _u0_u6_U203  ( .A(1'b1), .ZN(_u0_u6_ch_adr1[0] ) );
INV_X4 _u0_u6_U201  ( .A(1'b0), .ZN(_u0_u6_ch_am0[31] ) );
INV_X4 _u0_u6_U199  ( .A(1'b0), .ZN(_u0_u6_ch_am0[30] ) );
INV_X4 _u0_u6_U197  ( .A(1'b0), .ZN(_u0_u6_ch_am0[29] ) );
INV_X4 _u0_u6_U195  ( .A(1'b0), .ZN(_u0_u6_ch_am0[28] ) );
INV_X4 _u0_u6_U193  ( .A(1'b0), .ZN(_u0_u6_ch_am0[27] ) );
INV_X4 _u0_u6_U191  ( .A(1'b0), .ZN(_u0_u6_ch_am0[26] ) );
INV_X4 _u0_u6_U189  ( .A(1'b0), .ZN(_u0_u6_ch_am0[25] ) );
INV_X4 _u0_u6_U187  ( .A(1'b0), .ZN(_u0_u6_ch_am0[24] ) );
INV_X4 _u0_u6_U185  ( .A(1'b0), .ZN(_u0_u6_ch_am0[23] ) );
INV_X4 _u0_u6_U183  ( .A(1'b0), .ZN(_u0_u6_ch_am0[22] ) );
INV_X4 _u0_u6_U181  ( .A(1'b0), .ZN(_u0_u6_ch_am0[21] ) );
INV_X4 _u0_u6_U179  ( .A(1'b0), .ZN(_u0_u6_ch_am0[20] ) );
INV_X4 _u0_u6_U177  ( .A(1'b0), .ZN(_u0_u6_ch_am0[19] ) );
INV_X4 _u0_u6_U175  ( .A(1'b0), .ZN(_u0_u6_ch_am0[18] ) );
INV_X4 _u0_u6_U173  ( .A(1'b0), .ZN(_u0_u6_ch_am0[17] ) );
INV_X4 _u0_u6_U171  ( .A(1'b0), .ZN(_u0_u6_ch_am0[16] ) );
INV_X4 _u0_u6_U169  ( .A(1'b0), .ZN(_u0_u6_ch_am0[15] ) );
INV_X4 _u0_u6_U167  ( .A(1'b0), .ZN(_u0_u6_ch_am0[14] ) );
INV_X4 _u0_u6_U165  ( .A(1'b0), .ZN(_u0_u6_ch_am0[13] ) );
INV_X4 _u0_u6_U163  ( .A(1'b0), .ZN(_u0_u6_ch_am0[12] ) );
INV_X4 _u0_u6_U161  ( .A(1'b0), .ZN(_u0_u6_ch_am0[11] ) );
INV_X4 _u0_u6_U159  ( .A(1'b0), .ZN(_u0_u6_ch_am0[10] ) );
INV_X4 _u0_u6_U157  ( .A(1'b0), .ZN(_u0_u6_ch_am0[9] ) );
INV_X4 _u0_u6_U155  ( .A(1'b0), .ZN(_u0_u6_ch_am0[8] ) );
INV_X4 _u0_u6_U153  ( .A(1'b0), .ZN(_u0_u6_ch_am0[7] ) );
INV_X4 _u0_u6_U151  ( .A(1'b0), .ZN(_u0_u6_ch_am0[6] ) );
INV_X4 _u0_u6_U149  ( .A(1'b0), .ZN(_u0_u6_ch_am0[5] ) );
INV_X4 _u0_u6_U147  ( .A(1'b0), .ZN(_u0_u6_ch_am0[4] ) );
INV_X4 _u0_u6_U145  ( .A(1'b1), .ZN(_u0_u6_ch_am0[3] ) );
INV_X4 _u0_u6_U143  ( .A(1'b1), .ZN(_u0_u6_ch_am0[2] ) );
INV_X4 _u0_u6_U141  ( .A(1'b1), .ZN(_u0_u6_ch_am0[1] ) );
INV_X4 _u0_u6_U139  ( .A(1'b1), .ZN(_u0_u6_ch_am0[0] ) );
INV_X4 _u0_u6_U137  ( .A(1'b0), .ZN(_u0_u6_ch_am1[31] ) );
INV_X4 _u0_u6_U135  ( .A(1'b0), .ZN(_u0_u6_ch_am1[30] ) );
INV_X4 _u0_u6_U133  ( .A(1'b0), .ZN(_u0_u6_ch_am1[29] ) );
INV_X4 _u0_u6_U131  ( .A(1'b0), .ZN(_u0_u6_ch_am1[28] ) );
INV_X4 _u0_u6_U129  ( .A(1'b0), .ZN(_u0_u6_ch_am1[27] ) );
INV_X4 _u0_u6_U127  ( .A(1'b0), .ZN(_u0_u6_ch_am1[26] ) );
INV_X4 _u0_u6_U125  ( .A(1'b0), .ZN(_u0_u6_ch_am1[25] ) );
INV_X4 _u0_u6_U123  ( .A(1'b0), .ZN(_u0_u6_ch_am1[24] ) );
INV_X4 _u0_u6_U121  ( .A(1'b0), .ZN(_u0_u6_ch_am1[23] ) );
INV_X4 _u0_u6_U119  ( .A(1'b0), .ZN(_u0_u6_ch_am1[22] ) );
INV_X4 _u0_u6_U117  ( .A(1'b0), .ZN(_u0_u6_ch_am1[21] ) );
INV_X4 _u0_u6_U115  ( .A(1'b0), .ZN(_u0_u6_ch_am1[20] ) );
INV_X4 _u0_u6_U113  ( .A(1'b0), .ZN(_u0_u6_ch_am1[19] ) );
INV_X4 _u0_u6_U111  ( .A(1'b0), .ZN(_u0_u6_ch_am1[18] ) );
INV_X4 _u0_u6_U109  ( .A(1'b0), .ZN(_u0_u6_ch_am1[17] ) );
INV_X4 _u0_u6_U107  ( .A(1'b0), .ZN(_u0_u6_ch_am1[16] ) );
INV_X4 _u0_u6_U105  ( .A(1'b0), .ZN(_u0_u6_ch_am1[15] ) );
INV_X4 _u0_u6_U103  ( .A(1'b0), .ZN(_u0_u6_ch_am1[14] ) );
INV_X4 _u0_u6_U101  ( .A(1'b0), .ZN(_u0_u6_ch_am1[13] ) );
INV_X4 _u0_u6_U99  ( .A(1'b0), .ZN(_u0_u6_ch_am1[12] ) );
INV_X4 _u0_u6_U97  ( .A(1'b0), .ZN(_u0_u6_ch_am1[11] ) );
INV_X4 _u0_u6_U95  ( .A(1'b0), .ZN(_u0_u6_ch_am1[10] ) );
INV_X4 _u0_u6_U93  ( .A(1'b0), .ZN(_u0_u6_ch_am1[9] ) );
INV_X4 _u0_u6_U91  ( .A(1'b0), .ZN(_u0_u6_ch_am1[8] ) );
INV_X4 _u0_u6_U89  ( .A(1'b0), .ZN(_u0_u6_ch_am1[7] ) );
INV_X4 _u0_u6_U87  ( .A(1'b0), .ZN(_u0_u6_ch_am1[6] ) );
INV_X4 _u0_u6_U85  ( .A(1'b0), .ZN(_u0_u6_ch_am1[5] ) );
INV_X4 _u0_u6_U83  ( .A(1'b0), .ZN(_u0_u6_ch_am1[4] ) );
INV_X4 _u0_u6_U81  ( .A(1'b1), .ZN(_u0_u6_ch_am1[3] ) );
INV_X4 _u0_u6_U79  ( .A(1'b1), .ZN(_u0_u6_ch_am1[2] ) );
INV_X4 _u0_u6_U77  ( .A(1'b1), .ZN(_u0_u6_ch_am1[1] ) );
INV_X4 _u0_u6_U75  ( .A(1'b1), .ZN(_u0_u6_ch_am1[0] ) );
INV_X4 _u0_u6_U73  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[31] ) );
INV_X4 _u0_u6_U71  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[30] ) );
INV_X4 _u0_u6_U69  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[29] ) );
INV_X4 _u0_u6_U67  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[28] ) );
INV_X4 _u0_u6_U65  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[27] ) );
INV_X4 _u0_u6_U63  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[26] ) );
INV_X4 _u0_u6_U61  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[25] ) );
INV_X4 _u0_u6_U59  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[24] ) );
INV_X4 _u0_u6_U57  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[23] ) );
INV_X4 _u0_u6_U55  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[22] ) );
INV_X4 _u0_u6_U53  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[21] ) );
INV_X4 _u0_u6_U51  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[20] ) );
INV_X4 _u0_u6_U49  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[19] ) );
INV_X4 _u0_u6_U47  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[18] ) );
INV_X4 _u0_u6_U45  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[17] ) );
INV_X4 _u0_u6_U43  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[16] ) );
INV_X4 _u0_u6_U41  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[15] ) );
INV_X4 _u0_u6_U39  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[14] ) );
INV_X4 _u0_u6_U37  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[13] ) );
INV_X4 _u0_u6_U35  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[12] ) );
INV_X4 _u0_u6_U33  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[11] ) );
INV_X4 _u0_u6_U31  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[10] ) );
INV_X4 _u0_u6_U29  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[9] ) );
INV_X4 _u0_u6_U27  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[8] ) );
INV_X4 _u0_u6_U25  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[7] ) );
INV_X4 _u0_u6_U23  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[6] ) );
INV_X4 _u0_u6_U21  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[5] ) );
INV_X4 _u0_u6_U19  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[4] ) );
INV_X4 _u0_u6_U17  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[3] ) );
INV_X4 _u0_u6_U15  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[2] ) );
INV_X4 _u0_u6_U13  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[1] ) );
INV_X4 _u0_u6_U11  ( .A(1'b1), .ZN(_u0_u6_sw_pointer[0] ) );
INV_X4 _u0_u6_U9  ( .A(1'b1), .ZN(_u0_u6_ch_stop ) );
INV_X4 _u0_u6_U7  ( .A(1'b1), .ZN(_u0_u6_ch_dis ) );
INV_X4 _u0_u6_U5  ( .A(1'b1), .ZN(_u0_u6_int ) );
INV_X4 _u0_u7_U585  ( .A(1'b1), .ZN(_u0_u7_pointer[31] ) );
INV_X4 _u0_u7_U583  ( .A(1'b1), .ZN(_u0_u7_pointer[30] ) );
INV_X4 _u0_u7_U581  ( .A(1'b1), .ZN(_u0_u7_pointer[29] ) );
INV_X4 _u0_u7_U579  ( .A(1'b1), .ZN(_u0_u7_pointer[28] ) );
INV_X4 _u0_u7_U577  ( .A(1'b1), .ZN(_u0_u7_pointer[27] ) );
INV_X4 _u0_u7_U575  ( .A(1'b1), .ZN(_u0_u7_pointer[26] ) );
INV_X4 _u0_u7_U573  ( .A(1'b1), .ZN(_u0_u7_pointer[25] ) );
INV_X4 _u0_u7_U571  ( .A(1'b1), .ZN(_u0_u7_pointer[24] ) );
INV_X4 _u0_u7_U569  ( .A(1'b1), .ZN(_u0_u7_pointer[23] ) );
INV_X4 _u0_u7_U567  ( .A(1'b1), .ZN(_u0_u7_pointer[22] ) );
INV_X4 _u0_u7_U565  ( .A(1'b1), .ZN(_u0_u7_pointer[21] ) );
INV_X4 _u0_u7_U563  ( .A(1'b1), .ZN(_u0_u7_pointer[20] ) );
INV_X4 _u0_u7_U561  ( .A(1'b1), .ZN(_u0_u7_pointer[19] ) );
INV_X4 _u0_u7_U559  ( .A(1'b1), .ZN(_u0_u7_pointer[18] ) );
INV_X4 _u0_u7_U557  ( .A(1'b1), .ZN(_u0_u7_pointer[17] ) );
INV_X4 _u0_u7_U555  ( .A(1'b1), .ZN(_u0_u7_pointer[16] ) );
INV_X4 _u0_u7_U553  ( .A(1'b1), .ZN(_u0_u7_pointer[15] ) );
INV_X4 _u0_u7_U551  ( .A(1'b1), .ZN(_u0_u7_pointer[14] ) );
INV_X4 _u0_u7_U549  ( .A(1'b1), .ZN(_u0_u7_pointer[13] ) );
INV_X4 _u0_u7_U547  ( .A(1'b1), .ZN(_u0_u7_pointer[12] ) );
INV_X4 _u0_u7_U545  ( .A(1'b1), .ZN(_u0_u7_pointer[11] ) );
INV_X4 _u0_u7_U543  ( .A(1'b1), .ZN(_u0_u7_pointer[10] ) );
INV_X4 _u0_u7_U541  ( .A(1'b1), .ZN(_u0_u7_pointer[9] ) );
INV_X4 _u0_u7_U539  ( .A(1'b1), .ZN(_u0_u7_pointer[8] ) );
INV_X4 _u0_u7_U537  ( .A(1'b1), .ZN(_u0_u7_pointer[7] ) );
INV_X4 _u0_u7_U535  ( .A(1'b1), .ZN(_u0_u7_pointer[6] ) );
INV_X4 _u0_u7_U533  ( .A(1'b1), .ZN(_u0_u7_pointer[5] ) );
INV_X4 _u0_u7_U531  ( .A(1'b1), .ZN(_u0_u7_pointer[4] ) );
INV_X4 _u0_u7_U529  ( .A(1'b1), .ZN(_u0_u7_pointer[3] ) );
INV_X4 _u0_u7_U527  ( .A(1'b1), .ZN(_u0_u7_pointer[2] ) );
INV_X4 _u0_u7_U525  ( .A(1'b1), .ZN(_u0_u7_pointer[1] ) );
INV_X4 _u0_u7_U523  ( .A(1'b1), .ZN(_u0_u7_pointer[0] ) );
INV_X4 _u0_u7_U521  ( .A(1'b1), .ZN(_u0_u7_pointer_s[31] ) );
INV_X4 _u0_u7_U519  ( .A(1'b1), .ZN(_u0_u7_pointer_s[30] ) );
INV_X4 _u0_u7_U517  ( .A(1'b1), .ZN(_u0_u7_pointer_s[29] ) );
INV_X4 _u0_u7_U515  ( .A(1'b1), .ZN(_u0_u7_pointer_s[28] ) );
INV_X4 _u0_u7_U513  ( .A(1'b1), .ZN(_u0_u7_pointer_s[27] ) );
INV_X4 _u0_u7_U511  ( .A(1'b1), .ZN(_u0_u7_pointer_s[26] ) );
INV_X4 _u0_u7_U509  ( .A(1'b1), .ZN(_u0_u7_pointer_s[25] ) );
INV_X4 _u0_u7_U507  ( .A(1'b1), .ZN(_u0_u7_pointer_s[24] ) );
INV_X4 _u0_u7_U505  ( .A(1'b1), .ZN(_u0_u7_pointer_s[23] ) );
INV_X4 _u0_u7_U503  ( .A(1'b1), .ZN(_u0_u7_pointer_s[22] ) );
INV_X4 _u0_u7_U501  ( .A(1'b1), .ZN(_u0_u7_pointer_s[21] ) );
INV_X4 _u0_u7_U499  ( .A(1'b1), .ZN(_u0_u7_pointer_s[20] ) );
INV_X4 _u0_u7_U497  ( .A(1'b1), .ZN(_u0_u7_pointer_s[19] ) );
INV_X4 _u0_u7_U495  ( .A(1'b1), .ZN(_u0_u7_pointer_s[18] ) );
INV_X4 _u0_u7_U493  ( .A(1'b1), .ZN(_u0_u7_pointer_s[17] ) );
INV_X4 _u0_u7_U491  ( .A(1'b1), .ZN(_u0_u7_pointer_s[16] ) );
INV_X4 _u0_u7_U489  ( .A(1'b1), .ZN(_u0_u7_pointer_s[15] ) );
INV_X4 _u0_u7_U487  ( .A(1'b1), .ZN(_u0_u7_pointer_s[14] ) );
INV_X4 _u0_u7_U485  ( .A(1'b1), .ZN(_u0_u7_pointer_s[13] ) );
INV_X4 _u0_u7_U483  ( .A(1'b1), .ZN(_u0_u7_pointer_s[12] ) );
INV_X4 _u0_u7_U481  ( .A(1'b1), .ZN(_u0_u7_pointer_s[11] ) );
INV_X4 _u0_u7_U479  ( .A(1'b1), .ZN(_u0_u7_pointer_s[10] ) );
INV_X4 _u0_u7_U477  ( .A(1'b1), .ZN(_u0_u7_pointer_s[9] ) );
INV_X4 _u0_u7_U475  ( .A(1'b1), .ZN(_u0_u7_pointer_s[8] ) );
INV_X4 _u0_u7_U473  ( .A(1'b1), .ZN(_u0_u7_pointer_s[7] ) );
INV_X4 _u0_u7_U471  ( .A(1'b1), .ZN(_u0_u7_pointer_s[6] ) );
INV_X4 _u0_u7_U469  ( .A(1'b1), .ZN(_u0_u7_pointer_s[5] ) );
INV_X4 _u0_u7_U467  ( .A(1'b1), .ZN(_u0_u7_pointer_s[4] ) );
INV_X4 _u0_u7_U465  ( .A(1'b1), .ZN(_u0_u7_pointer_s[3] ) );
INV_X4 _u0_u7_U463  ( .A(1'b1), .ZN(_u0_u7_pointer_s[2] ) );
INV_X4 _u0_u7_U461  ( .A(1'b1), .ZN(_u0_u7_pointer_s[1] ) );
INV_X4 _u0_u7_U459  ( .A(1'b1), .ZN(_u0_u7_pointer_s[0] ) );
INV_X4 _u0_u7_U457  ( .A(1'b1), .ZN(_u0_u7_ch_csr[31] ) );
INV_X4 _u0_u7_U455  ( .A(1'b1), .ZN(_u0_u7_ch_csr[30] ) );
INV_X4 _u0_u7_U453  ( .A(1'b1), .ZN(_u0_u7_ch_csr[29] ) );
INV_X4 _u0_u7_U451  ( .A(1'b1), .ZN(_u0_u7_ch_csr[28] ) );
INV_X4 _u0_u7_U449  ( .A(1'b1), .ZN(_u0_u7_ch_csr[27] ) );
INV_X4 _u0_u7_U447  ( .A(1'b1), .ZN(_u0_u7_ch_csr[26] ) );
INV_X4 _u0_u7_U445  ( .A(1'b1), .ZN(_u0_u7_ch_csr[25] ) );
INV_X4 _u0_u7_U443  ( .A(1'b1), .ZN(_u0_u7_ch_csr[24] ) );
INV_X4 _u0_u7_U441  ( .A(1'b1), .ZN(_u0_u7_ch_csr[23] ) );
INV_X4 _u0_u7_U439  ( .A(1'b1), .ZN(_u0_u7_ch_csr[22] ) );
INV_X4 _u0_u7_U437  ( .A(1'b1), .ZN(_u0_u7_ch_csr[21] ) );
INV_X4 _u0_u7_U435  ( .A(1'b1), .ZN(_u0_u7_ch_csr[20] ) );
INV_X4 _u0_u7_U433  ( .A(1'b1), .ZN(_u0_u7_ch_csr[19] ) );
INV_X4 _u0_u7_U431  ( .A(1'b1), .ZN(_u0_u7_ch_csr[18] ) );
INV_X4 _u0_u7_U429  ( .A(1'b1), .ZN(_u0_u7_ch_csr[17] ) );
INV_X4 _u0_u7_U427  ( .A(1'b1), .ZN(_u0_u7_ch_csr[16] ) );
INV_X4 _u0_u7_U425  ( .A(1'b1), .ZN(_u0_u7_ch_csr[15] ) );
INV_X4 _u0_u7_U423  ( .A(1'b1), .ZN(_u0_u7_ch_csr[14] ) );
INV_X4 _u0_u7_U421  ( .A(1'b1), .ZN(_u0_u7_ch_csr[13] ) );
INV_X4 _u0_u7_U419  ( .A(1'b1), .ZN(_u0_u7_ch_csr[12] ) );
INV_X4 _u0_u7_U417  ( .A(1'b1), .ZN(_u0_u7_ch_csr[11] ) );
INV_X4 _u0_u7_U415  ( .A(1'b1), .ZN(_u0_u7_ch_csr[10] ) );
INV_X4 _u0_u7_U413  ( .A(1'b1), .ZN(_u0_u7_ch_csr[9] ) );
INV_X4 _u0_u7_U411  ( .A(1'b1), .ZN(_u0_u7_ch_csr[8] ) );
INV_X4 _u0_u7_U409  ( .A(1'b1), .ZN(_u0_u7_ch_csr[7] ) );
INV_X4 _u0_u7_U407  ( .A(1'b1), .ZN(_u0_u7_ch_csr[6] ) );
INV_X4 _u0_u7_U405  ( .A(1'b1), .ZN(_u0_u7_ch_csr[5] ) );
INV_X4 _u0_u7_U403  ( .A(1'b1), .ZN(_u0_u7_ch_csr[4] ) );
INV_X4 _u0_u7_U401  ( .A(1'b1), .ZN(_u0_u7_ch_csr[3] ) );
INV_X4 _u0_u7_U399  ( .A(1'b1), .ZN(_u0_u7_ch_csr[2] ) );
INV_X4 _u0_u7_U397  ( .A(1'b1), .ZN(_u0_u7_ch_csr[1] ) );
INV_X4 _u0_u7_U395  ( .A(1'b1), .ZN(_u0_u7_ch_csr[0] ) );
INV_X4 _u0_u7_U393  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[31] ) );
INV_X4 _u0_u7_U391  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[30] ) );
INV_X4 _u0_u7_U389  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[29] ) );
INV_X4 _u0_u7_U387  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[28] ) );
INV_X4 _u0_u7_U385  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[27] ) );
INV_X4 _u0_u7_U383  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[26] ) );
INV_X4 _u0_u7_U381  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[25] ) );
INV_X4 _u0_u7_U379  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[24] ) );
INV_X4 _u0_u7_U377  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[23] ) );
INV_X4 _u0_u7_U375  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[22] ) );
INV_X4 _u0_u7_U373  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[21] ) );
INV_X4 _u0_u7_U371  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[20] ) );
INV_X4 _u0_u7_U369  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[19] ) );
INV_X4 _u0_u7_U367  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[18] ) );
INV_X4 _u0_u7_U365  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[17] ) );
INV_X4 _u0_u7_U363  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[16] ) );
INV_X4 _u0_u7_U361  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[15] ) );
INV_X4 _u0_u7_U359  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[14] ) );
INV_X4 _u0_u7_U357  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[13] ) );
INV_X4 _u0_u7_U355  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[12] ) );
INV_X4 _u0_u7_U353  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[11] ) );
INV_X4 _u0_u7_U351  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[10] ) );
INV_X4 _u0_u7_U349  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[9] ) );
INV_X4 _u0_u7_U347  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[8] ) );
INV_X4 _u0_u7_U345  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[7] ) );
INV_X4 _u0_u7_U343  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[6] ) );
INV_X4 _u0_u7_U341  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[5] ) );
INV_X4 _u0_u7_U339  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[4] ) );
INV_X4 _u0_u7_U337  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[3] ) );
INV_X4 _u0_u7_U335  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[2] ) );
INV_X4 _u0_u7_U333  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[1] ) );
INV_X4 _u0_u7_U331  ( .A(1'b1), .ZN(_u0_u7_ch_txsz[0] ) );
INV_X4 _u0_u7_U329  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[31] ) );
INV_X4 _u0_u7_U327  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[30] ) );
INV_X4 _u0_u7_U325  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[29] ) );
INV_X4 _u0_u7_U323  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[28] ) );
INV_X4 _u0_u7_U321  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[27] ) );
INV_X4 _u0_u7_U319  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[26] ) );
INV_X4 _u0_u7_U317  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[25] ) );
INV_X4 _u0_u7_U315  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[24] ) );
INV_X4 _u0_u7_U313  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[23] ) );
INV_X4 _u0_u7_U311  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[22] ) );
INV_X4 _u0_u7_U309  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[21] ) );
INV_X4 _u0_u7_U307  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[20] ) );
INV_X4 _u0_u7_U305  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[19] ) );
INV_X4 _u0_u7_U303  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[18] ) );
INV_X4 _u0_u7_U301  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[17] ) );
INV_X4 _u0_u7_U299  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[16] ) );
INV_X4 _u0_u7_U297  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[15] ) );
INV_X4 _u0_u7_U295  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[14] ) );
INV_X4 _u0_u7_U293  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[13] ) );
INV_X4 _u0_u7_U291  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[12] ) );
INV_X4 _u0_u7_U289  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[11] ) );
INV_X4 _u0_u7_U287  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[10] ) );
INV_X4 _u0_u7_U285  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[9] ) );
INV_X4 _u0_u7_U283  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[8] ) );
INV_X4 _u0_u7_U281  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[7] ) );
INV_X4 _u0_u7_U279  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[6] ) );
INV_X4 _u0_u7_U277  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[5] ) );
INV_X4 _u0_u7_U275  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[4] ) );
INV_X4 _u0_u7_U273  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[3] ) );
INV_X4 _u0_u7_U271  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[2] ) );
INV_X4 _u0_u7_U269  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[1] ) );
INV_X4 _u0_u7_U267  ( .A(1'b1), .ZN(_u0_u7_ch_adr0[0] ) );
INV_X4 _u0_u7_U265  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[31] ) );
INV_X4 _u0_u7_U263  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[30] ) );
INV_X4 _u0_u7_U261  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[29] ) );
INV_X4 _u0_u7_U259  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[28] ) );
INV_X4 _u0_u7_U257  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[27] ) );
INV_X4 _u0_u7_U255  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[26] ) );
INV_X4 _u0_u7_U253  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[25] ) );
INV_X4 _u0_u7_U251  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[24] ) );
INV_X4 _u0_u7_U249  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[23] ) );
INV_X4 _u0_u7_U247  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[22] ) );
INV_X4 _u0_u7_U245  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[21] ) );
INV_X4 _u0_u7_U243  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[20] ) );
INV_X4 _u0_u7_U241  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[19] ) );
INV_X4 _u0_u7_U239  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[18] ) );
INV_X4 _u0_u7_U237  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[17] ) );
INV_X4 _u0_u7_U235  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[16] ) );
INV_X4 _u0_u7_U233  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[15] ) );
INV_X4 _u0_u7_U231  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[14] ) );
INV_X4 _u0_u7_U229  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[13] ) );
INV_X4 _u0_u7_U227  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[12] ) );
INV_X4 _u0_u7_U225  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[11] ) );
INV_X4 _u0_u7_U223  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[10] ) );
INV_X4 _u0_u7_U221  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[9] ) );
INV_X4 _u0_u7_U219  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[8] ) );
INV_X4 _u0_u7_U217  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[7] ) );
INV_X4 _u0_u7_U215  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[6] ) );
INV_X4 _u0_u7_U213  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[5] ) );
INV_X4 _u0_u7_U211  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[4] ) );
INV_X4 _u0_u7_U209  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[3] ) );
INV_X4 _u0_u7_U207  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[2] ) );
INV_X4 _u0_u7_U205  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[1] ) );
INV_X4 _u0_u7_U203  ( .A(1'b1), .ZN(_u0_u7_ch_adr1[0] ) );
INV_X4 _u0_u7_U201  ( .A(1'b0), .ZN(_u0_u7_ch_am0[31] ) );
INV_X4 _u0_u7_U199  ( .A(1'b0), .ZN(_u0_u7_ch_am0[30] ) );
INV_X4 _u0_u7_U197  ( .A(1'b0), .ZN(_u0_u7_ch_am0[29] ) );
INV_X4 _u0_u7_U195  ( .A(1'b0), .ZN(_u0_u7_ch_am0[28] ) );
INV_X4 _u0_u7_U193  ( .A(1'b0), .ZN(_u0_u7_ch_am0[27] ) );
INV_X4 _u0_u7_U191  ( .A(1'b0), .ZN(_u0_u7_ch_am0[26] ) );
INV_X4 _u0_u7_U189  ( .A(1'b0), .ZN(_u0_u7_ch_am0[25] ) );
INV_X4 _u0_u7_U187  ( .A(1'b0), .ZN(_u0_u7_ch_am0[24] ) );
INV_X4 _u0_u7_U185  ( .A(1'b0), .ZN(_u0_u7_ch_am0[23] ) );
INV_X4 _u0_u7_U183  ( .A(1'b0), .ZN(_u0_u7_ch_am0[22] ) );
INV_X4 _u0_u7_U181  ( .A(1'b0), .ZN(_u0_u7_ch_am0[21] ) );
INV_X4 _u0_u7_U179  ( .A(1'b0), .ZN(_u0_u7_ch_am0[20] ) );
INV_X4 _u0_u7_U177  ( .A(1'b0), .ZN(_u0_u7_ch_am0[19] ) );
INV_X4 _u0_u7_U175  ( .A(1'b0), .ZN(_u0_u7_ch_am0[18] ) );
INV_X4 _u0_u7_U173  ( .A(1'b0), .ZN(_u0_u7_ch_am0[17] ) );
INV_X4 _u0_u7_U171  ( .A(1'b0), .ZN(_u0_u7_ch_am0[16] ) );
INV_X4 _u0_u7_U169  ( .A(1'b0), .ZN(_u0_u7_ch_am0[15] ) );
INV_X4 _u0_u7_U167  ( .A(1'b0), .ZN(_u0_u7_ch_am0[14] ) );
INV_X4 _u0_u7_U165  ( .A(1'b0), .ZN(_u0_u7_ch_am0[13] ) );
INV_X4 _u0_u7_U163  ( .A(1'b0), .ZN(_u0_u7_ch_am0[12] ) );
INV_X4 _u0_u7_U161  ( .A(1'b0), .ZN(_u0_u7_ch_am0[11] ) );
INV_X4 _u0_u7_U159  ( .A(1'b0), .ZN(_u0_u7_ch_am0[10] ) );
INV_X4 _u0_u7_U157  ( .A(1'b0), .ZN(_u0_u7_ch_am0[9] ) );
INV_X4 _u0_u7_U155  ( .A(1'b0), .ZN(_u0_u7_ch_am0[8] ) );
INV_X4 _u0_u7_U153  ( .A(1'b0), .ZN(_u0_u7_ch_am0[7] ) );
INV_X4 _u0_u7_U151  ( .A(1'b0), .ZN(_u0_u7_ch_am0[6] ) );
INV_X4 _u0_u7_U149  ( .A(1'b0), .ZN(_u0_u7_ch_am0[5] ) );
INV_X4 _u0_u7_U147  ( .A(1'b0), .ZN(_u0_u7_ch_am0[4] ) );
INV_X4 _u0_u7_U145  ( .A(1'b1), .ZN(_u0_u7_ch_am0[3] ) );
INV_X4 _u0_u7_U143  ( .A(1'b1), .ZN(_u0_u7_ch_am0[2] ) );
INV_X4 _u0_u7_U141  ( .A(1'b1), .ZN(_u0_u7_ch_am0[1] ) );
INV_X4 _u0_u7_U139  ( .A(1'b1), .ZN(_u0_u7_ch_am0[0] ) );
INV_X4 _u0_u7_U137  ( .A(1'b0), .ZN(_u0_u7_ch_am1[31] ) );
INV_X4 _u0_u7_U135  ( .A(1'b0), .ZN(_u0_u7_ch_am1[30] ) );
INV_X4 _u0_u7_U133  ( .A(1'b0), .ZN(_u0_u7_ch_am1[29] ) );
INV_X4 _u0_u7_U131  ( .A(1'b0), .ZN(_u0_u7_ch_am1[28] ) );
INV_X4 _u0_u7_U129  ( .A(1'b0), .ZN(_u0_u7_ch_am1[27] ) );
INV_X4 _u0_u7_U127  ( .A(1'b0), .ZN(_u0_u7_ch_am1[26] ) );
INV_X4 _u0_u7_U125  ( .A(1'b0), .ZN(_u0_u7_ch_am1[25] ) );
INV_X4 _u0_u7_U123  ( .A(1'b0), .ZN(_u0_u7_ch_am1[24] ) );
INV_X4 _u0_u7_U121  ( .A(1'b0), .ZN(_u0_u7_ch_am1[23] ) );
INV_X4 _u0_u7_U119  ( .A(1'b0), .ZN(_u0_u7_ch_am1[22] ) );
INV_X4 _u0_u7_U117  ( .A(1'b0), .ZN(_u0_u7_ch_am1[21] ) );
INV_X4 _u0_u7_U115  ( .A(1'b0), .ZN(_u0_u7_ch_am1[20] ) );
INV_X4 _u0_u7_U113  ( .A(1'b0), .ZN(_u0_u7_ch_am1[19] ) );
INV_X4 _u0_u7_U111  ( .A(1'b0), .ZN(_u0_u7_ch_am1[18] ) );
INV_X4 _u0_u7_U109  ( .A(1'b0), .ZN(_u0_u7_ch_am1[17] ) );
INV_X4 _u0_u7_U107  ( .A(1'b0), .ZN(_u0_u7_ch_am1[16] ) );
INV_X4 _u0_u7_U105  ( .A(1'b0), .ZN(_u0_u7_ch_am1[15] ) );
INV_X4 _u0_u7_U103  ( .A(1'b0), .ZN(_u0_u7_ch_am1[14] ) );
INV_X4 _u0_u7_U101  ( .A(1'b0), .ZN(_u0_u7_ch_am1[13] ) );
INV_X4 _u0_u7_U99  ( .A(1'b0), .ZN(_u0_u7_ch_am1[12] ) );
INV_X4 _u0_u7_U97  ( .A(1'b0), .ZN(_u0_u7_ch_am1[11] ) );
INV_X4 _u0_u7_U95  ( .A(1'b0), .ZN(_u0_u7_ch_am1[10] ) );
INV_X4 _u0_u7_U93  ( .A(1'b0), .ZN(_u0_u7_ch_am1[9] ) );
INV_X4 _u0_u7_U91  ( .A(1'b0), .ZN(_u0_u7_ch_am1[8] ) );
INV_X4 _u0_u7_U89  ( .A(1'b0), .ZN(_u0_u7_ch_am1[7] ) );
INV_X4 _u0_u7_U87  ( .A(1'b0), .ZN(_u0_u7_ch_am1[6] ) );
INV_X4 _u0_u7_U85  ( .A(1'b0), .ZN(_u0_u7_ch_am1[5] ) );
INV_X4 _u0_u7_U83  ( .A(1'b0), .ZN(_u0_u7_ch_am1[4] ) );
INV_X4 _u0_u7_U81  ( .A(1'b1), .ZN(_u0_u7_ch_am1[3] ) );
INV_X4 _u0_u7_U79  ( .A(1'b1), .ZN(_u0_u7_ch_am1[2] ) );
INV_X4 _u0_u7_U77  ( .A(1'b1), .ZN(_u0_u7_ch_am1[1] ) );
INV_X4 _u0_u7_U75  ( .A(1'b1), .ZN(_u0_u7_ch_am1[0] ) );
INV_X4 _u0_u7_U73  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[31] ) );
INV_X4 _u0_u7_U71  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[30] ) );
INV_X4 _u0_u7_U69  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[29] ) );
INV_X4 _u0_u7_U67  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[28] ) );
INV_X4 _u0_u7_U65  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[27] ) );
INV_X4 _u0_u7_U63  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[26] ) );
INV_X4 _u0_u7_U61  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[25] ) );
INV_X4 _u0_u7_U59  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[24] ) );
INV_X4 _u0_u7_U57  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[23] ) );
INV_X4 _u0_u7_U55  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[22] ) );
INV_X4 _u0_u7_U53  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[21] ) );
INV_X4 _u0_u7_U51  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[20] ) );
INV_X4 _u0_u7_U49  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[19] ) );
INV_X4 _u0_u7_U47  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[18] ) );
INV_X4 _u0_u7_U45  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[17] ) );
INV_X4 _u0_u7_U43  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[16] ) );
INV_X4 _u0_u7_U41  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[15] ) );
INV_X4 _u0_u7_U39  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[14] ) );
INV_X4 _u0_u7_U37  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[13] ) );
INV_X4 _u0_u7_U35  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[12] ) );
INV_X4 _u0_u7_U33  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[11] ) );
INV_X4 _u0_u7_U31  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[10] ) );
INV_X4 _u0_u7_U29  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[9] ) );
INV_X4 _u0_u7_U27  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[8] ) );
INV_X4 _u0_u7_U25  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[7] ) );
INV_X4 _u0_u7_U23  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[6] ) );
INV_X4 _u0_u7_U21  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[5] ) );
INV_X4 _u0_u7_U19  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[4] ) );
INV_X4 _u0_u7_U17  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[3] ) );
INV_X4 _u0_u7_U15  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[2] ) );
INV_X4 _u0_u7_U13  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[1] ) );
INV_X4 _u0_u7_U11  ( .A(1'b1), .ZN(_u0_u7_sw_pointer[0] ) );
INV_X4 _u0_u7_U9  ( .A(1'b1), .ZN(_u0_u7_ch_stop ) );
INV_X4 _u0_u7_U7  ( .A(1'b1), .ZN(_u0_u7_ch_dis ) );
INV_X4 _u0_u7_U5  ( .A(1'b1), .ZN(_u0_u7_int ) );
INV_X4 _u0_u8_U585  ( .A(1'b1), .ZN(_u0_u8_pointer[31] ) );
INV_X4 _u0_u8_U583  ( .A(1'b1), .ZN(_u0_u8_pointer[30] ) );
INV_X4 _u0_u8_U581  ( .A(1'b1), .ZN(_u0_u8_pointer[29] ) );
INV_X4 _u0_u8_U579  ( .A(1'b1), .ZN(_u0_u8_pointer[28] ) );
INV_X4 _u0_u8_U577  ( .A(1'b1), .ZN(_u0_u8_pointer[27] ) );
INV_X4 _u0_u8_U575  ( .A(1'b1), .ZN(_u0_u8_pointer[26] ) );
INV_X4 _u0_u8_U573  ( .A(1'b1), .ZN(_u0_u8_pointer[25] ) );
INV_X4 _u0_u8_U571  ( .A(1'b1), .ZN(_u0_u8_pointer[24] ) );
INV_X4 _u0_u8_U569  ( .A(1'b1), .ZN(_u0_u8_pointer[23] ) );
INV_X4 _u0_u8_U567  ( .A(1'b1), .ZN(_u0_u8_pointer[22] ) );
INV_X4 _u0_u8_U565  ( .A(1'b1), .ZN(_u0_u8_pointer[21] ) );
INV_X4 _u0_u8_U563  ( .A(1'b1), .ZN(_u0_u8_pointer[20] ) );
INV_X4 _u0_u8_U561  ( .A(1'b1), .ZN(_u0_u8_pointer[19] ) );
INV_X4 _u0_u8_U559  ( .A(1'b1), .ZN(_u0_u8_pointer[18] ) );
INV_X4 _u0_u8_U557  ( .A(1'b1), .ZN(_u0_u8_pointer[17] ) );
INV_X4 _u0_u8_U555  ( .A(1'b1), .ZN(_u0_u8_pointer[16] ) );
INV_X4 _u0_u8_U553  ( .A(1'b1), .ZN(_u0_u8_pointer[15] ) );
INV_X4 _u0_u8_U551  ( .A(1'b1), .ZN(_u0_u8_pointer[14] ) );
INV_X4 _u0_u8_U549  ( .A(1'b1), .ZN(_u0_u8_pointer[13] ) );
INV_X4 _u0_u8_U547  ( .A(1'b1), .ZN(_u0_u8_pointer[12] ) );
INV_X4 _u0_u8_U545  ( .A(1'b1), .ZN(_u0_u8_pointer[11] ) );
INV_X4 _u0_u8_U543  ( .A(1'b1), .ZN(_u0_u8_pointer[10] ) );
INV_X4 _u0_u8_U541  ( .A(1'b1), .ZN(_u0_u8_pointer[9] ) );
INV_X4 _u0_u8_U539  ( .A(1'b1), .ZN(_u0_u8_pointer[8] ) );
INV_X4 _u0_u8_U537  ( .A(1'b1), .ZN(_u0_u8_pointer[7] ) );
INV_X4 _u0_u8_U535  ( .A(1'b1), .ZN(_u0_u8_pointer[6] ) );
INV_X4 _u0_u8_U533  ( .A(1'b1), .ZN(_u0_u8_pointer[5] ) );
INV_X4 _u0_u8_U531  ( .A(1'b1), .ZN(_u0_u8_pointer[4] ) );
INV_X4 _u0_u8_U529  ( .A(1'b1), .ZN(_u0_u8_pointer[3] ) );
INV_X4 _u0_u8_U527  ( .A(1'b1), .ZN(_u0_u8_pointer[2] ) );
INV_X4 _u0_u8_U525  ( .A(1'b1), .ZN(_u0_u8_pointer[1] ) );
INV_X4 _u0_u8_U523  ( .A(1'b1), .ZN(_u0_u8_pointer[0] ) );
INV_X4 _u0_u8_U521  ( .A(1'b1), .ZN(_u0_u8_pointer_s[31] ) );
INV_X4 _u0_u8_U519  ( .A(1'b1), .ZN(_u0_u8_pointer_s[30] ) );
INV_X4 _u0_u8_U517  ( .A(1'b1), .ZN(_u0_u8_pointer_s[29] ) );
INV_X4 _u0_u8_U515  ( .A(1'b1), .ZN(_u0_u8_pointer_s[28] ) );
INV_X4 _u0_u8_U513  ( .A(1'b1), .ZN(_u0_u8_pointer_s[27] ) );
INV_X4 _u0_u8_U511  ( .A(1'b1), .ZN(_u0_u8_pointer_s[26] ) );
INV_X4 _u0_u8_U509  ( .A(1'b1), .ZN(_u0_u8_pointer_s[25] ) );
INV_X4 _u0_u8_U507  ( .A(1'b1), .ZN(_u0_u8_pointer_s[24] ) );
INV_X4 _u0_u8_U505  ( .A(1'b1), .ZN(_u0_u8_pointer_s[23] ) );
INV_X4 _u0_u8_U503  ( .A(1'b1), .ZN(_u0_u8_pointer_s[22] ) );
INV_X4 _u0_u8_U501  ( .A(1'b1), .ZN(_u0_u8_pointer_s[21] ) );
INV_X4 _u0_u8_U499  ( .A(1'b1), .ZN(_u0_u8_pointer_s[20] ) );
INV_X4 _u0_u8_U497  ( .A(1'b1), .ZN(_u0_u8_pointer_s[19] ) );
INV_X4 _u0_u8_U495  ( .A(1'b1), .ZN(_u0_u8_pointer_s[18] ) );
INV_X4 _u0_u8_U493  ( .A(1'b1), .ZN(_u0_u8_pointer_s[17] ) );
INV_X4 _u0_u8_U491  ( .A(1'b1), .ZN(_u0_u8_pointer_s[16] ) );
INV_X4 _u0_u8_U489  ( .A(1'b1), .ZN(_u0_u8_pointer_s[15] ) );
INV_X4 _u0_u8_U487  ( .A(1'b1), .ZN(_u0_u8_pointer_s[14] ) );
INV_X4 _u0_u8_U485  ( .A(1'b1), .ZN(_u0_u8_pointer_s[13] ) );
INV_X4 _u0_u8_U483  ( .A(1'b1), .ZN(_u0_u8_pointer_s[12] ) );
INV_X4 _u0_u8_U481  ( .A(1'b1), .ZN(_u0_u8_pointer_s[11] ) );
INV_X4 _u0_u8_U479  ( .A(1'b1), .ZN(_u0_u8_pointer_s[10] ) );
INV_X4 _u0_u8_U477  ( .A(1'b1), .ZN(_u0_u8_pointer_s[9] ) );
INV_X4 _u0_u8_U475  ( .A(1'b1), .ZN(_u0_u8_pointer_s[8] ) );
INV_X4 _u0_u8_U473  ( .A(1'b1), .ZN(_u0_u8_pointer_s[7] ) );
INV_X4 _u0_u8_U471  ( .A(1'b1), .ZN(_u0_u8_pointer_s[6] ) );
INV_X4 _u0_u8_U469  ( .A(1'b1), .ZN(_u0_u8_pointer_s[5] ) );
INV_X4 _u0_u8_U467  ( .A(1'b1), .ZN(_u0_u8_pointer_s[4] ) );
INV_X4 _u0_u8_U465  ( .A(1'b1), .ZN(_u0_u8_pointer_s[3] ) );
INV_X4 _u0_u8_U463  ( .A(1'b1), .ZN(_u0_u8_pointer_s[2] ) );
INV_X4 _u0_u8_U461  ( .A(1'b1), .ZN(_u0_u8_pointer_s[1] ) );
INV_X4 _u0_u8_U459  ( .A(1'b1), .ZN(_u0_u8_pointer_s[0] ) );
INV_X4 _u0_u8_U457  ( .A(1'b1), .ZN(_u0_u8_ch_csr[31] ) );
INV_X4 _u0_u8_U455  ( .A(1'b1), .ZN(_u0_u8_ch_csr[30] ) );
INV_X4 _u0_u8_U453  ( .A(1'b1), .ZN(_u0_u8_ch_csr[29] ) );
INV_X4 _u0_u8_U451  ( .A(1'b1), .ZN(_u0_u8_ch_csr[28] ) );
INV_X4 _u0_u8_U449  ( .A(1'b1), .ZN(_u0_u8_ch_csr[27] ) );
INV_X4 _u0_u8_U447  ( .A(1'b1), .ZN(_u0_u8_ch_csr[26] ) );
INV_X4 _u0_u8_U445  ( .A(1'b1), .ZN(_u0_u8_ch_csr[25] ) );
INV_X4 _u0_u8_U443  ( .A(1'b1), .ZN(_u0_u8_ch_csr[24] ) );
INV_X4 _u0_u8_U441  ( .A(1'b1), .ZN(_u0_u8_ch_csr[23] ) );
INV_X4 _u0_u8_U439  ( .A(1'b1), .ZN(_u0_u8_ch_csr[22] ) );
INV_X4 _u0_u8_U437  ( .A(1'b1), .ZN(_u0_u8_ch_csr[21] ) );
INV_X4 _u0_u8_U435  ( .A(1'b1), .ZN(_u0_u8_ch_csr[20] ) );
INV_X4 _u0_u8_U433  ( .A(1'b1), .ZN(_u0_u8_ch_csr[19] ) );
INV_X4 _u0_u8_U431  ( .A(1'b1), .ZN(_u0_u8_ch_csr[18] ) );
INV_X4 _u0_u8_U429  ( .A(1'b1), .ZN(_u0_u8_ch_csr[17] ) );
INV_X4 _u0_u8_U427  ( .A(1'b1), .ZN(_u0_u8_ch_csr[16] ) );
INV_X4 _u0_u8_U425  ( .A(1'b1), .ZN(_u0_u8_ch_csr[15] ) );
INV_X4 _u0_u8_U423  ( .A(1'b1), .ZN(_u0_u8_ch_csr[14] ) );
INV_X4 _u0_u8_U421  ( .A(1'b1), .ZN(_u0_u8_ch_csr[13] ) );
INV_X4 _u0_u8_U419  ( .A(1'b1), .ZN(_u0_u8_ch_csr[12] ) );
INV_X4 _u0_u8_U417  ( .A(1'b1), .ZN(_u0_u8_ch_csr[11] ) );
INV_X4 _u0_u8_U415  ( .A(1'b1), .ZN(_u0_u8_ch_csr[10] ) );
INV_X4 _u0_u8_U413  ( .A(1'b1), .ZN(_u0_u8_ch_csr[9] ) );
INV_X4 _u0_u8_U411  ( .A(1'b1), .ZN(_u0_u8_ch_csr[8] ) );
INV_X4 _u0_u8_U409  ( .A(1'b1), .ZN(_u0_u8_ch_csr[7] ) );
INV_X4 _u0_u8_U407  ( .A(1'b1), .ZN(_u0_u8_ch_csr[6] ) );
INV_X4 _u0_u8_U405  ( .A(1'b1), .ZN(_u0_u8_ch_csr[5] ) );
INV_X4 _u0_u8_U403  ( .A(1'b1), .ZN(_u0_u8_ch_csr[4] ) );
INV_X4 _u0_u8_U401  ( .A(1'b1), .ZN(_u0_u8_ch_csr[3] ) );
INV_X4 _u0_u8_U399  ( .A(1'b1), .ZN(_u0_u8_ch_csr[2] ) );
INV_X4 _u0_u8_U397  ( .A(1'b1), .ZN(_u0_u8_ch_csr[1] ) );
INV_X4 _u0_u8_U395  ( .A(1'b1), .ZN(_u0_u8_ch_csr[0] ) );
INV_X4 _u0_u8_U393  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[31] ) );
INV_X4 _u0_u8_U391  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[30] ) );
INV_X4 _u0_u8_U389  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[29] ) );
INV_X4 _u0_u8_U387  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[28] ) );
INV_X4 _u0_u8_U385  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[27] ) );
INV_X4 _u0_u8_U383  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[26] ) );
INV_X4 _u0_u8_U381  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[25] ) );
INV_X4 _u0_u8_U379  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[24] ) );
INV_X4 _u0_u8_U377  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[23] ) );
INV_X4 _u0_u8_U375  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[22] ) );
INV_X4 _u0_u8_U373  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[21] ) );
INV_X4 _u0_u8_U371  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[20] ) );
INV_X4 _u0_u8_U369  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[19] ) );
INV_X4 _u0_u8_U367  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[18] ) );
INV_X4 _u0_u8_U365  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[17] ) );
INV_X4 _u0_u8_U363  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[16] ) );
INV_X4 _u0_u8_U361  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[15] ) );
INV_X4 _u0_u8_U359  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[14] ) );
INV_X4 _u0_u8_U357  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[13] ) );
INV_X4 _u0_u8_U355  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[12] ) );
INV_X4 _u0_u8_U353  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[11] ) );
INV_X4 _u0_u8_U351  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[10] ) );
INV_X4 _u0_u8_U349  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[9] ) );
INV_X4 _u0_u8_U347  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[8] ) );
INV_X4 _u0_u8_U345  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[7] ) );
INV_X4 _u0_u8_U343  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[6] ) );
INV_X4 _u0_u8_U341  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[5] ) );
INV_X4 _u0_u8_U339  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[4] ) );
INV_X4 _u0_u8_U337  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[3] ) );
INV_X4 _u0_u8_U335  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[2] ) );
INV_X4 _u0_u8_U333  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[1] ) );
INV_X4 _u0_u8_U331  ( .A(1'b1), .ZN(_u0_u8_ch_txsz[0] ) );
INV_X4 _u0_u8_U329  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[31] ) );
INV_X4 _u0_u8_U327  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[30] ) );
INV_X4 _u0_u8_U325  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[29] ) );
INV_X4 _u0_u8_U323  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[28] ) );
INV_X4 _u0_u8_U321  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[27] ) );
INV_X4 _u0_u8_U319  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[26] ) );
INV_X4 _u0_u8_U317  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[25] ) );
INV_X4 _u0_u8_U315  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[24] ) );
INV_X4 _u0_u8_U313  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[23] ) );
INV_X4 _u0_u8_U311  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[22] ) );
INV_X4 _u0_u8_U309  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[21] ) );
INV_X4 _u0_u8_U307  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[20] ) );
INV_X4 _u0_u8_U305  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[19] ) );
INV_X4 _u0_u8_U303  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[18] ) );
INV_X4 _u0_u8_U301  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[17] ) );
INV_X4 _u0_u8_U299  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[16] ) );
INV_X4 _u0_u8_U297  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[15] ) );
INV_X4 _u0_u8_U295  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[14] ) );
INV_X4 _u0_u8_U293  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[13] ) );
INV_X4 _u0_u8_U291  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[12] ) );
INV_X4 _u0_u8_U289  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[11] ) );
INV_X4 _u0_u8_U287  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[10] ) );
INV_X4 _u0_u8_U285  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[9] ) );
INV_X4 _u0_u8_U283  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[8] ) );
INV_X4 _u0_u8_U281  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[7] ) );
INV_X4 _u0_u8_U279  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[6] ) );
INV_X4 _u0_u8_U277  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[5] ) );
INV_X4 _u0_u8_U275  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[4] ) );
INV_X4 _u0_u8_U273  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[3] ) );
INV_X4 _u0_u8_U271  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[2] ) );
INV_X4 _u0_u8_U269  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[1] ) );
INV_X4 _u0_u8_U267  ( .A(1'b1), .ZN(_u0_u8_ch_adr0[0] ) );
INV_X4 _u0_u8_U265  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[31] ) );
INV_X4 _u0_u8_U263  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[30] ) );
INV_X4 _u0_u8_U261  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[29] ) );
INV_X4 _u0_u8_U259  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[28] ) );
INV_X4 _u0_u8_U257  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[27] ) );
INV_X4 _u0_u8_U255  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[26] ) );
INV_X4 _u0_u8_U253  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[25] ) );
INV_X4 _u0_u8_U251  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[24] ) );
INV_X4 _u0_u8_U249  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[23] ) );
INV_X4 _u0_u8_U247  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[22] ) );
INV_X4 _u0_u8_U245  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[21] ) );
INV_X4 _u0_u8_U243  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[20] ) );
INV_X4 _u0_u8_U241  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[19] ) );
INV_X4 _u0_u8_U239  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[18] ) );
INV_X4 _u0_u8_U237  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[17] ) );
INV_X4 _u0_u8_U235  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[16] ) );
INV_X4 _u0_u8_U233  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[15] ) );
INV_X4 _u0_u8_U231  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[14] ) );
INV_X4 _u0_u8_U229  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[13] ) );
INV_X4 _u0_u8_U227  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[12] ) );
INV_X4 _u0_u8_U225  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[11] ) );
INV_X4 _u0_u8_U223  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[10] ) );
INV_X4 _u0_u8_U221  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[9] ) );
INV_X4 _u0_u8_U219  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[8] ) );
INV_X4 _u0_u8_U217  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[7] ) );
INV_X4 _u0_u8_U215  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[6] ) );
INV_X4 _u0_u8_U213  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[5] ) );
INV_X4 _u0_u8_U211  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[4] ) );
INV_X4 _u0_u8_U209  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[3] ) );
INV_X4 _u0_u8_U207  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[2] ) );
INV_X4 _u0_u8_U205  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[1] ) );
INV_X4 _u0_u8_U203  ( .A(1'b1), .ZN(_u0_u8_ch_adr1[0] ) );
INV_X4 _u0_u8_U201  ( .A(1'b0), .ZN(_u0_u8_ch_am0[31] ) );
INV_X4 _u0_u8_U199  ( .A(1'b0), .ZN(_u0_u8_ch_am0[30] ) );
INV_X4 _u0_u8_U197  ( .A(1'b0), .ZN(_u0_u8_ch_am0[29] ) );
INV_X4 _u0_u8_U195  ( .A(1'b0), .ZN(_u0_u8_ch_am0[28] ) );
INV_X4 _u0_u8_U193  ( .A(1'b0), .ZN(_u0_u8_ch_am0[27] ) );
INV_X4 _u0_u8_U191  ( .A(1'b0), .ZN(_u0_u8_ch_am0[26] ) );
INV_X4 _u0_u8_U189  ( .A(1'b0), .ZN(_u0_u8_ch_am0[25] ) );
INV_X4 _u0_u8_U187  ( .A(1'b0), .ZN(_u0_u8_ch_am0[24] ) );
INV_X4 _u0_u8_U185  ( .A(1'b0), .ZN(_u0_u8_ch_am0[23] ) );
INV_X4 _u0_u8_U183  ( .A(1'b0), .ZN(_u0_u8_ch_am0[22] ) );
INV_X4 _u0_u8_U181  ( .A(1'b0), .ZN(_u0_u8_ch_am0[21] ) );
INV_X4 _u0_u8_U179  ( .A(1'b0), .ZN(_u0_u8_ch_am0[20] ) );
INV_X4 _u0_u8_U177  ( .A(1'b0), .ZN(_u0_u8_ch_am0[19] ) );
INV_X4 _u0_u8_U175  ( .A(1'b0), .ZN(_u0_u8_ch_am0[18] ) );
INV_X4 _u0_u8_U173  ( .A(1'b0), .ZN(_u0_u8_ch_am0[17] ) );
INV_X4 _u0_u8_U171  ( .A(1'b0), .ZN(_u0_u8_ch_am0[16] ) );
INV_X4 _u0_u8_U169  ( .A(1'b0), .ZN(_u0_u8_ch_am0[15] ) );
INV_X4 _u0_u8_U167  ( .A(1'b0), .ZN(_u0_u8_ch_am0[14] ) );
INV_X4 _u0_u8_U165  ( .A(1'b0), .ZN(_u0_u8_ch_am0[13] ) );
INV_X4 _u0_u8_U163  ( .A(1'b0), .ZN(_u0_u8_ch_am0[12] ) );
INV_X4 _u0_u8_U161  ( .A(1'b0), .ZN(_u0_u8_ch_am0[11] ) );
INV_X4 _u0_u8_U159  ( .A(1'b0), .ZN(_u0_u8_ch_am0[10] ) );
INV_X4 _u0_u8_U157  ( .A(1'b0), .ZN(_u0_u8_ch_am0[9] ) );
INV_X4 _u0_u8_U155  ( .A(1'b0), .ZN(_u0_u8_ch_am0[8] ) );
INV_X4 _u0_u8_U153  ( .A(1'b0), .ZN(_u0_u8_ch_am0[7] ) );
INV_X4 _u0_u8_U151  ( .A(1'b0), .ZN(_u0_u8_ch_am0[6] ) );
INV_X4 _u0_u8_U149  ( .A(1'b0), .ZN(_u0_u8_ch_am0[5] ) );
INV_X4 _u0_u8_U147  ( .A(1'b0), .ZN(_u0_u8_ch_am0[4] ) );
INV_X4 _u0_u8_U145  ( .A(1'b1), .ZN(_u0_u8_ch_am0[3] ) );
INV_X4 _u0_u8_U143  ( .A(1'b1), .ZN(_u0_u8_ch_am0[2] ) );
INV_X4 _u0_u8_U141  ( .A(1'b1), .ZN(_u0_u8_ch_am0[1] ) );
INV_X4 _u0_u8_U139  ( .A(1'b1), .ZN(_u0_u8_ch_am0[0] ) );
INV_X4 _u0_u8_U137  ( .A(1'b0), .ZN(_u0_u8_ch_am1[31] ) );
INV_X4 _u0_u8_U135  ( .A(1'b0), .ZN(_u0_u8_ch_am1[30] ) );
INV_X4 _u0_u8_U133  ( .A(1'b0), .ZN(_u0_u8_ch_am1[29] ) );
INV_X4 _u0_u8_U131  ( .A(1'b0), .ZN(_u0_u8_ch_am1[28] ) );
INV_X4 _u0_u8_U129  ( .A(1'b0), .ZN(_u0_u8_ch_am1[27] ) );
INV_X4 _u0_u8_U127  ( .A(1'b0), .ZN(_u0_u8_ch_am1[26] ) );
INV_X4 _u0_u8_U125  ( .A(1'b0), .ZN(_u0_u8_ch_am1[25] ) );
INV_X4 _u0_u8_U123  ( .A(1'b0), .ZN(_u0_u8_ch_am1[24] ) );
INV_X4 _u0_u8_U121  ( .A(1'b0), .ZN(_u0_u8_ch_am1[23] ) );
INV_X4 _u0_u8_U119  ( .A(1'b0), .ZN(_u0_u8_ch_am1[22] ) );
INV_X4 _u0_u8_U117  ( .A(1'b0), .ZN(_u0_u8_ch_am1[21] ) );
INV_X4 _u0_u8_U115  ( .A(1'b0), .ZN(_u0_u8_ch_am1[20] ) );
INV_X4 _u0_u8_U113  ( .A(1'b0), .ZN(_u0_u8_ch_am1[19] ) );
INV_X4 _u0_u8_U111  ( .A(1'b0), .ZN(_u0_u8_ch_am1[18] ) );
INV_X4 _u0_u8_U109  ( .A(1'b0), .ZN(_u0_u8_ch_am1[17] ) );
INV_X4 _u0_u8_U107  ( .A(1'b0), .ZN(_u0_u8_ch_am1[16] ) );
INV_X4 _u0_u8_U105  ( .A(1'b0), .ZN(_u0_u8_ch_am1[15] ) );
INV_X4 _u0_u8_U103  ( .A(1'b0), .ZN(_u0_u8_ch_am1[14] ) );
INV_X4 _u0_u8_U101  ( .A(1'b0), .ZN(_u0_u8_ch_am1[13] ) );
INV_X4 _u0_u8_U99  ( .A(1'b0), .ZN(_u0_u8_ch_am1[12] ) );
INV_X4 _u0_u8_U97  ( .A(1'b0), .ZN(_u0_u8_ch_am1[11] ) );
INV_X4 _u0_u8_U95  ( .A(1'b0), .ZN(_u0_u8_ch_am1[10] ) );
INV_X4 _u0_u8_U93  ( .A(1'b0), .ZN(_u0_u8_ch_am1[9] ) );
INV_X4 _u0_u8_U91  ( .A(1'b0), .ZN(_u0_u8_ch_am1[8] ) );
INV_X4 _u0_u8_U89  ( .A(1'b0), .ZN(_u0_u8_ch_am1[7] ) );
INV_X4 _u0_u8_U87  ( .A(1'b0), .ZN(_u0_u8_ch_am1[6] ) );
INV_X4 _u0_u8_U85  ( .A(1'b0), .ZN(_u0_u8_ch_am1[5] ) );
INV_X4 _u0_u8_U83  ( .A(1'b0), .ZN(_u0_u8_ch_am1[4] ) );
INV_X4 _u0_u8_U81  ( .A(1'b1), .ZN(_u0_u8_ch_am1[3] ) );
INV_X4 _u0_u8_U79  ( .A(1'b1), .ZN(_u0_u8_ch_am1[2] ) );
INV_X4 _u0_u8_U77  ( .A(1'b1), .ZN(_u0_u8_ch_am1[1] ) );
INV_X4 _u0_u8_U75  ( .A(1'b1), .ZN(_u0_u8_ch_am1[0] ) );
INV_X4 _u0_u8_U73  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[31] ) );
INV_X4 _u0_u8_U71  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[30] ) );
INV_X4 _u0_u8_U69  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[29] ) );
INV_X4 _u0_u8_U67  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[28] ) );
INV_X4 _u0_u8_U65  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[27] ) );
INV_X4 _u0_u8_U63  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[26] ) );
INV_X4 _u0_u8_U61  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[25] ) );
INV_X4 _u0_u8_U59  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[24] ) );
INV_X4 _u0_u8_U57  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[23] ) );
INV_X4 _u0_u8_U55  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[22] ) );
INV_X4 _u0_u8_U53  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[21] ) );
INV_X4 _u0_u8_U51  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[20] ) );
INV_X4 _u0_u8_U49  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[19] ) );
INV_X4 _u0_u8_U47  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[18] ) );
INV_X4 _u0_u8_U45  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[17] ) );
INV_X4 _u0_u8_U43  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[16] ) );
INV_X4 _u0_u8_U41  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[15] ) );
INV_X4 _u0_u8_U39  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[14] ) );
INV_X4 _u0_u8_U37  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[13] ) );
INV_X4 _u0_u8_U35  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[12] ) );
INV_X4 _u0_u8_U33  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[11] ) );
INV_X4 _u0_u8_U31  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[10] ) );
INV_X4 _u0_u8_U29  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[9] ) );
INV_X4 _u0_u8_U27  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[8] ) );
INV_X4 _u0_u8_U25  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[7] ) );
INV_X4 _u0_u8_U23  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[6] ) );
INV_X4 _u0_u8_U21  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[5] ) );
INV_X4 _u0_u8_U19  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[4] ) );
INV_X4 _u0_u8_U17  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[3] ) );
INV_X4 _u0_u8_U15  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[2] ) );
INV_X4 _u0_u8_U13  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[1] ) );
INV_X4 _u0_u8_U11  ( .A(1'b1), .ZN(_u0_u8_sw_pointer[0] ) );
INV_X4 _u0_u8_U9  ( .A(1'b1), .ZN(_u0_u8_ch_stop ) );
INV_X4 _u0_u8_U7  ( .A(1'b1), .ZN(_u0_u8_ch_dis ) );
INV_X4 _u0_u8_U5  ( .A(1'b1), .ZN(_u0_u8_int ) );
INV_X4 _u0_u9_U585  ( .A(1'b1), .ZN(_u0_u9_pointer[31] ) );
INV_X4 _u0_u9_U583  ( .A(1'b1), .ZN(_u0_u9_pointer[30] ) );
INV_X4 _u0_u9_U581  ( .A(1'b1), .ZN(_u0_u9_pointer[29] ) );
INV_X4 _u0_u9_U579  ( .A(1'b1), .ZN(_u0_u9_pointer[28] ) );
INV_X4 _u0_u9_U577  ( .A(1'b1), .ZN(_u0_u9_pointer[27] ) );
INV_X4 _u0_u9_U575  ( .A(1'b1), .ZN(_u0_u9_pointer[26] ) );
INV_X4 _u0_u9_U573  ( .A(1'b1), .ZN(_u0_u9_pointer[25] ) );
INV_X4 _u0_u9_U571  ( .A(1'b1), .ZN(_u0_u9_pointer[24] ) );
INV_X4 _u0_u9_U569  ( .A(1'b1), .ZN(_u0_u9_pointer[23] ) );
INV_X4 _u0_u9_U567  ( .A(1'b1), .ZN(_u0_u9_pointer[22] ) );
INV_X4 _u0_u9_U565  ( .A(1'b1), .ZN(_u0_u9_pointer[21] ) );
INV_X4 _u0_u9_U563  ( .A(1'b1), .ZN(_u0_u9_pointer[20] ) );
INV_X4 _u0_u9_U561  ( .A(1'b1), .ZN(_u0_u9_pointer[19] ) );
INV_X4 _u0_u9_U559  ( .A(1'b1), .ZN(_u0_u9_pointer[18] ) );
INV_X4 _u0_u9_U557  ( .A(1'b1), .ZN(_u0_u9_pointer[17] ) );
INV_X4 _u0_u9_U555  ( .A(1'b1), .ZN(_u0_u9_pointer[16] ) );
INV_X4 _u0_u9_U553  ( .A(1'b1), .ZN(_u0_u9_pointer[15] ) );
INV_X4 _u0_u9_U551  ( .A(1'b1), .ZN(_u0_u9_pointer[14] ) );
INV_X4 _u0_u9_U549  ( .A(1'b1), .ZN(_u0_u9_pointer[13] ) );
INV_X4 _u0_u9_U547  ( .A(1'b1), .ZN(_u0_u9_pointer[12] ) );
INV_X4 _u0_u9_U545  ( .A(1'b1), .ZN(_u0_u9_pointer[11] ) );
INV_X4 _u0_u9_U543  ( .A(1'b1), .ZN(_u0_u9_pointer[10] ) );
INV_X4 _u0_u9_U541  ( .A(1'b1), .ZN(_u0_u9_pointer[9] ) );
INV_X4 _u0_u9_U539  ( .A(1'b1), .ZN(_u0_u9_pointer[8] ) );
INV_X4 _u0_u9_U537  ( .A(1'b1), .ZN(_u0_u9_pointer[7] ) );
INV_X4 _u0_u9_U535  ( .A(1'b1), .ZN(_u0_u9_pointer[6] ) );
INV_X4 _u0_u9_U533  ( .A(1'b1), .ZN(_u0_u9_pointer[5] ) );
INV_X4 _u0_u9_U531  ( .A(1'b1), .ZN(_u0_u9_pointer[4] ) );
INV_X4 _u0_u9_U529  ( .A(1'b1), .ZN(_u0_u9_pointer[3] ) );
INV_X4 _u0_u9_U527  ( .A(1'b1), .ZN(_u0_u9_pointer[2] ) );
INV_X4 _u0_u9_U525  ( .A(1'b1), .ZN(_u0_u9_pointer[1] ) );
INV_X4 _u0_u9_U523  ( .A(1'b1), .ZN(_u0_u9_pointer[0] ) );
INV_X4 _u0_u9_U521  ( .A(1'b1), .ZN(_u0_u9_pointer_s[31] ) );
INV_X4 _u0_u9_U519  ( .A(1'b1), .ZN(_u0_u9_pointer_s[30] ) );
INV_X4 _u0_u9_U517  ( .A(1'b1), .ZN(_u0_u9_pointer_s[29] ) );
INV_X4 _u0_u9_U515  ( .A(1'b1), .ZN(_u0_u9_pointer_s[28] ) );
INV_X4 _u0_u9_U513  ( .A(1'b1), .ZN(_u0_u9_pointer_s[27] ) );
INV_X4 _u0_u9_U511  ( .A(1'b1), .ZN(_u0_u9_pointer_s[26] ) );
INV_X4 _u0_u9_U509  ( .A(1'b1), .ZN(_u0_u9_pointer_s[25] ) );
INV_X4 _u0_u9_U507  ( .A(1'b1), .ZN(_u0_u9_pointer_s[24] ) );
INV_X4 _u0_u9_U505  ( .A(1'b1), .ZN(_u0_u9_pointer_s[23] ) );
INV_X4 _u0_u9_U503  ( .A(1'b1), .ZN(_u0_u9_pointer_s[22] ) );
INV_X4 _u0_u9_U501  ( .A(1'b1), .ZN(_u0_u9_pointer_s[21] ) );
INV_X4 _u0_u9_U499  ( .A(1'b1), .ZN(_u0_u9_pointer_s[20] ) );
INV_X4 _u0_u9_U497  ( .A(1'b1), .ZN(_u0_u9_pointer_s[19] ) );
INV_X4 _u0_u9_U495  ( .A(1'b1), .ZN(_u0_u9_pointer_s[18] ) );
INV_X4 _u0_u9_U493  ( .A(1'b1), .ZN(_u0_u9_pointer_s[17] ) );
INV_X4 _u0_u9_U491  ( .A(1'b1), .ZN(_u0_u9_pointer_s[16] ) );
INV_X4 _u0_u9_U489  ( .A(1'b1), .ZN(_u0_u9_pointer_s[15] ) );
INV_X4 _u0_u9_U487  ( .A(1'b1), .ZN(_u0_u9_pointer_s[14] ) );
INV_X4 _u0_u9_U485  ( .A(1'b1), .ZN(_u0_u9_pointer_s[13] ) );
INV_X4 _u0_u9_U483  ( .A(1'b1), .ZN(_u0_u9_pointer_s[12] ) );
INV_X4 _u0_u9_U481  ( .A(1'b1), .ZN(_u0_u9_pointer_s[11] ) );
INV_X4 _u0_u9_U479  ( .A(1'b1), .ZN(_u0_u9_pointer_s[10] ) );
INV_X4 _u0_u9_U477  ( .A(1'b1), .ZN(_u0_u9_pointer_s[9] ) );
INV_X4 _u0_u9_U475  ( .A(1'b1), .ZN(_u0_u9_pointer_s[8] ) );
INV_X4 _u0_u9_U473  ( .A(1'b1), .ZN(_u0_u9_pointer_s[7] ) );
INV_X4 _u0_u9_U471  ( .A(1'b1), .ZN(_u0_u9_pointer_s[6] ) );
INV_X4 _u0_u9_U469  ( .A(1'b1), .ZN(_u0_u9_pointer_s[5] ) );
INV_X4 _u0_u9_U467  ( .A(1'b1), .ZN(_u0_u9_pointer_s[4] ) );
INV_X4 _u0_u9_U465  ( .A(1'b1), .ZN(_u0_u9_pointer_s[3] ) );
INV_X4 _u0_u9_U463  ( .A(1'b1), .ZN(_u0_u9_pointer_s[2] ) );
INV_X4 _u0_u9_U461  ( .A(1'b1), .ZN(_u0_u9_pointer_s[1] ) );
INV_X4 _u0_u9_U459  ( .A(1'b1), .ZN(_u0_u9_pointer_s[0] ) );
INV_X4 _u0_u9_U457  ( .A(1'b1), .ZN(_u0_u9_ch_csr[31] ) );
INV_X4 _u0_u9_U455  ( .A(1'b1), .ZN(_u0_u9_ch_csr[30] ) );
INV_X4 _u0_u9_U453  ( .A(1'b1), .ZN(_u0_u9_ch_csr[29] ) );
INV_X4 _u0_u9_U451  ( .A(1'b1), .ZN(_u0_u9_ch_csr[28] ) );
INV_X4 _u0_u9_U449  ( .A(1'b1), .ZN(_u0_u9_ch_csr[27] ) );
INV_X4 _u0_u9_U447  ( .A(1'b1), .ZN(_u0_u9_ch_csr[26] ) );
INV_X4 _u0_u9_U445  ( .A(1'b1), .ZN(_u0_u9_ch_csr[25] ) );
INV_X4 _u0_u9_U443  ( .A(1'b1), .ZN(_u0_u9_ch_csr[24] ) );
INV_X4 _u0_u9_U441  ( .A(1'b1), .ZN(_u0_u9_ch_csr[23] ) );
INV_X4 _u0_u9_U439  ( .A(1'b1), .ZN(_u0_u9_ch_csr[22] ) );
INV_X4 _u0_u9_U437  ( .A(1'b1), .ZN(_u0_u9_ch_csr[21] ) );
INV_X4 _u0_u9_U435  ( .A(1'b1), .ZN(_u0_u9_ch_csr[20] ) );
INV_X4 _u0_u9_U433  ( .A(1'b1), .ZN(_u0_u9_ch_csr[19] ) );
INV_X4 _u0_u9_U431  ( .A(1'b1), .ZN(_u0_u9_ch_csr[18] ) );
INV_X4 _u0_u9_U429  ( .A(1'b1), .ZN(_u0_u9_ch_csr[17] ) );
INV_X4 _u0_u9_U427  ( .A(1'b1), .ZN(_u0_u9_ch_csr[16] ) );
INV_X4 _u0_u9_U425  ( .A(1'b1), .ZN(_u0_u9_ch_csr[15] ) );
INV_X4 _u0_u9_U423  ( .A(1'b1), .ZN(_u0_u9_ch_csr[14] ) );
INV_X4 _u0_u9_U421  ( .A(1'b1), .ZN(_u0_u9_ch_csr[13] ) );
INV_X4 _u0_u9_U419  ( .A(1'b1), .ZN(_u0_u9_ch_csr[12] ) );
INV_X4 _u0_u9_U417  ( .A(1'b1), .ZN(_u0_u9_ch_csr[11] ) );
INV_X4 _u0_u9_U415  ( .A(1'b1), .ZN(_u0_u9_ch_csr[10] ) );
INV_X4 _u0_u9_U413  ( .A(1'b1), .ZN(_u0_u9_ch_csr[9] ) );
INV_X4 _u0_u9_U411  ( .A(1'b1), .ZN(_u0_u9_ch_csr[8] ) );
INV_X4 _u0_u9_U409  ( .A(1'b1), .ZN(_u0_u9_ch_csr[7] ) );
INV_X4 _u0_u9_U407  ( .A(1'b1), .ZN(_u0_u9_ch_csr[6] ) );
INV_X4 _u0_u9_U405  ( .A(1'b1), .ZN(_u0_u9_ch_csr[5] ) );
INV_X4 _u0_u9_U403  ( .A(1'b1), .ZN(_u0_u9_ch_csr[4] ) );
INV_X4 _u0_u9_U401  ( .A(1'b1), .ZN(_u0_u9_ch_csr[3] ) );
INV_X4 _u0_u9_U399  ( .A(1'b1), .ZN(_u0_u9_ch_csr[2] ) );
INV_X4 _u0_u9_U397  ( .A(1'b1), .ZN(_u0_u9_ch_csr[1] ) );
INV_X4 _u0_u9_U395  ( .A(1'b1), .ZN(_u0_u9_ch_csr[0] ) );
INV_X4 _u0_u9_U393  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[31] ) );
INV_X4 _u0_u9_U391  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[30] ) );
INV_X4 _u0_u9_U389  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[29] ) );
INV_X4 _u0_u9_U387  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[28] ) );
INV_X4 _u0_u9_U385  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[27] ) );
INV_X4 _u0_u9_U383  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[26] ) );
INV_X4 _u0_u9_U381  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[25] ) );
INV_X4 _u0_u9_U379  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[24] ) );
INV_X4 _u0_u9_U377  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[23] ) );
INV_X4 _u0_u9_U375  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[22] ) );
INV_X4 _u0_u9_U373  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[21] ) );
INV_X4 _u0_u9_U371  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[20] ) );
INV_X4 _u0_u9_U369  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[19] ) );
INV_X4 _u0_u9_U367  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[18] ) );
INV_X4 _u0_u9_U365  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[17] ) );
INV_X4 _u0_u9_U363  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[16] ) );
INV_X4 _u0_u9_U361  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[15] ) );
INV_X4 _u0_u9_U359  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[14] ) );
INV_X4 _u0_u9_U357  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[13] ) );
INV_X4 _u0_u9_U355  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[12] ) );
INV_X4 _u0_u9_U353  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[11] ) );
INV_X4 _u0_u9_U351  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[10] ) );
INV_X4 _u0_u9_U349  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[9] ) );
INV_X4 _u0_u9_U347  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[8] ) );
INV_X4 _u0_u9_U345  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[7] ) );
INV_X4 _u0_u9_U343  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[6] ) );
INV_X4 _u0_u9_U341  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[5] ) );
INV_X4 _u0_u9_U339  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[4] ) );
INV_X4 _u0_u9_U337  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[3] ) );
INV_X4 _u0_u9_U335  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[2] ) );
INV_X4 _u0_u9_U333  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[1] ) );
INV_X4 _u0_u9_U331  ( .A(1'b1), .ZN(_u0_u9_ch_txsz[0] ) );
INV_X4 _u0_u9_U329  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[31] ) );
INV_X4 _u0_u9_U327  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[30] ) );
INV_X4 _u0_u9_U325  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[29] ) );
INV_X4 _u0_u9_U323  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[28] ) );
INV_X4 _u0_u9_U321  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[27] ) );
INV_X4 _u0_u9_U319  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[26] ) );
INV_X4 _u0_u9_U317  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[25] ) );
INV_X4 _u0_u9_U315  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[24] ) );
INV_X4 _u0_u9_U313  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[23] ) );
INV_X4 _u0_u9_U311  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[22] ) );
INV_X4 _u0_u9_U309  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[21] ) );
INV_X4 _u0_u9_U307  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[20] ) );
INV_X4 _u0_u9_U305  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[19] ) );
INV_X4 _u0_u9_U303  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[18] ) );
INV_X4 _u0_u9_U301  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[17] ) );
INV_X4 _u0_u9_U299  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[16] ) );
INV_X4 _u0_u9_U297  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[15] ) );
INV_X4 _u0_u9_U295  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[14] ) );
INV_X4 _u0_u9_U293  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[13] ) );
INV_X4 _u0_u9_U291  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[12] ) );
INV_X4 _u0_u9_U289  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[11] ) );
INV_X4 _u0_u9_U287  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[10] ) );
INV_X4 _u0_u9_U285  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[9] ) );
INV_X4 _u0_u9_U283  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[8] ) );
INV_X4 _u0_u9_U281  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[7] ) );
INV_X4 _u0_u9_U279  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[6] ) );
INV_X4 _u0_u9_U277  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[5] ) );
INV_X4 _u0_u9_U275  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[4] ) );
INV_X4 _u0_u9_U273  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[3] ) );
INV_X4 _u0_u9_U271  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[2] ) );
INV_X4 _u0_u9_U269  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[1] ) );
INV_X4 _u0_u9_U267  ( .A(1'b1), .ZN(_u0_u9_ch_adr0[0] ) );
INV_X4 _u0_u9_U265  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[31] ) );
INV_X4 _u0_u9_U263  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[30] ) );
INV_X4 _u0_u9_U261  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[29] ) );
INV_X4 _u0_u9_U259  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[28] ) );
INV_X4 _u0_u9_U257  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[27] ) );
INV_X4 _u0_u9_U255  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[26] ) );
INV_X4 _u0_u9_U253  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[25] ) );
INV_X4 _u0_u9_U251  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[24] ) );
INV_X4 _u0_u9_U249  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[23] ) );
INV_X4 _u0_u9_U247  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[22] ) );
INV_X4 _u0_u9_U245  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[21] ) );
INV_X4 _u0_u9_U243  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[20] ) );
INV_X4 _u0_u9_U241  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[19] ) );
INV_X4 _u0_u9_U239  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[18] ) );
INV_X4 _u0_u9_U237  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[17] ) );
INV_X4 _u0_u9_U235  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[16] ) );
INV_X4 _u0_u9_U233  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[15] ) );
INV_X4 _u0_u9_U231  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[14] ) );
INV_X4 _u0_u9_U229  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[13] ) );
INV_X4 _u0_u9_U227  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[12] ) );
INV_X4 _u0_u9_U225  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[11] ) );
INV_X4 _u0_u9_U223  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[10] ) );
INV_X4 _u0_u9_U221  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[9] ) );
INV_X4 _u0_u9_U219  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[8] ) );
INV_X4 _u0_u9_U217  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[7] ) );
INV_X4 _u0_u9_U215  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[6] ) );
INV_X4 _u0_u9_U213  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[5] ) );
INV_X4 _u0_u9_U211  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[4] ) );
INV_X4 _u0_u9_U209  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[3] ) );
INV_X4 _u0_u9_U207  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[2] ) );
INV_X4 _u0_u9_U205  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[1] ) );
INV_X4 _u0_u9_U203  ( .A(1'b1), .ZN(_u0_u9_ch_adr1[0] ) );
INV_X4 _u0_u9_U201  ( .A(1'b0), .ZN(_u0_u9_ch_am0[31] ) );
INV_X4 _u0_u9_U199  ( .A(1'b0), .ZN(_u0_u9_ch_am0[30] ) );
INV_X4 _u0_u9_U197  ( .A(1'b0), .ZN(_u0_u9_ch_am0[29] ) );
INV_X4 _u0_u9_U195  ( .A(1'b0), .ZN(_u0_u9_ch_am0[28] ) );
INV_X4 _u0_u9_U193  ( .A(1'b0), .ZN(_u0_u9_ch_am0[27] ) );
INV_X4 _u0_u9_U191  ( .A(1'b0), .ZN(_u0_u9_ch_am0[26] ) );
INV_X4 _u0_u9_U189  ( .A(1'b0), .ZN(_u0_u9_ch_am0[25] ) );
INV_X4 _u0_u9_U187  ( .A(1'b0), .ZN(_u0_u9_ch_am0[24] ) );
INV_X4 _u0_u9_U185  ( .A(1'b0), .ZN(_u0_u9_ch_am0[23] ) );
INV_X4 _u0_u9_U183  ( .A(1'b0), .ZN(_u0_u9_ch_am0[22] ) );
INV_X4 _u0_u9_U181  ( .A(1'b0), .ZN(_u0_u9_ch_am0[21] ) );
INV_X4 _u0_u9_U179  ( .A(1'b0), .ZN(_u0_u9_ch_am0[20] ) );
INV_X4 _u0_u9_U177  ( .A(1'b0), .ZN(_u0_u9_ch_am0[19] ) );
INV_X4 _u0_u9_U175  ( .A(1'b0), .ZN(_u0_u9_ch_am0[18] ) );
INV_X4 _u0_u9_U173  ( .A(1'b0), .ZN(_u0_u9_ch_am0[17] ) );
INV_X4 _u0_u9_U171  ( .A(1'b0), .ZN(_u0_u9_ch_am0[16] ) );
INV_X4 _u0_u9_U169  ( .A(1'b0), .ZN(_u0_u9_ch_am0[15] ) );
INV_X4 _u0_u9_U167  ( .A(1'b0), .ZN(_u0_u9_ch_am0[14] ) );
INV_X4 _u0_u9_U165  ( .A(1'b0), .ZN(_u0_u9_ch_am0[13] ) );
INV_X4 _u0_u9_U163  ( .A(1'b0), .ZN(_u0_u9_ch_am0[12] ) );
INV_X4 _u0_u9_U161  ( .A(1'b0), .ZN(_u0_u9_ch_am0[11] ) );
INV_X4 _u0_u9_U159  ( .A(1'b0), .ZN(_u0_u9_ch_am0[10] ) );
INV_X4 _u0_u9_U157  ( .A(1'b0), .ZN(_u0_u9_ch_am0[9] ) );
INV_X4 _u0_u9_U155  ( .A(1'b0), .ZN(_u0_u9_ch_am0[8] ) );
INV_X4 _u0_u9_U153  ( .A(1'b0), .ZN(_u0_u9_ch_am0[7] ) );
INV_X4 _u0_u9_U151  ( .A(1'b0), .ZN(_u0_u9_ch_am0[6] ) );
INV_X4 _u0_u9_U149  ( .A(1'b0), .ZN(_u0_u9_ch_am0[5] ) );
INV_X4 _u0_u9_U147  ( .A(1'b0), .ZN(_u0_u9_ch_am0[4] ) );
INV_X4 _u0_u9_U145  ( .A(1'b1), .ZN(_u0_u9_ch_am0[3] ) );
INV_X4 _u0_u9_U143  ( .A(1'b1), .ZN(_u0_u9_ch_am0[2] ) );
INV_X4 _u0_u9_U141  ( .A(1'b1), .ZN(_u0_u9_ch_am0[1] ) );
INV_X4 _u0_u9_U139  ( .A(1'b1), .ZN(_u0_u9_ch_am0[0] ) );
INV_X4 _u0_u9_U137  ( .A(1'b0), .ZN(_u0_u9_ch_am1[31] ) );
INV_X4 _u0_u9_U135  ( .A(1'b0), .ZN(_u0_u9_ch_am1[30] ) );
INV_X4 _u0_u9_U133  ( .A(1'b0), .ZN(_u0_u9_ch_am1[29] ) );
INV_X4 _u0_u9_U131  ( .A(1'b0), .ZN(_u0_u9_ch_am1[28] ) );
INV_X4 _u0_u9_U129  ( .A(1'b0), .ZN(_u0_u9_ch_am1[27] ) );
INV_X4 _u0_u9_U127  ( .A(1'b0), .ZN(_u0_u9_ch_am1[26] ) );
INV_X4 _u0_u9_U125  ( .A(1'b0), .ZN(_u0_u9_ch_am1[25] ) );
INV_X4 _u0_u9_U123  ( .A(1'b0), .ZN(_u0_u9_ch_am1[24] ) );
INV_X4 _u0_u9_U121  ( .A(1'b0), .ZN(_u0_u9_ch_am1[23] ) );
INV_X4 _u0_u9_U119  ( .A(1'b0), .ZN(_u0_u9_ch_am1[22] ) );
INV_X4 _u0_u9_U117  ( .A(1'b0), .ZN(_u0_u9_ch_am1[21] ) );
INV_X4 _u0_u9_U115  ( .A(1'b0), .ZN(_u0_u9_ch_am1[20] ) );
INV_X4 _u0_u9_U113  ( .A(1'b0), .ZN(_u0_u9_ch_am1[19] ) );
INV_X4 _u0_u9_U111  ( .A(1'b0), .ZN(_u0_u9_ch_am1[18] ) );
INV_X4 _u0_u9_U109  ( .A(1'b0), .ZN(_u0_u9_ch_am1[17] ) );
INV_X4 _u0_u9_U107  ( .A(1'b0), .ZN(_u0_u9_ch_am1[16] ) );
INV_X4 _u0_u9_U105  ( .A(1'b0), .ZN(_u0_u9_ch_am1[15] ) );
INV_X4 _u0_u9_U103  ( .A(1'b0), .ZN(_u0_u9_ch_am1[14] ) );
INV_X4 _u0_u9_U101  ( .A(1'b0), .ZN(_u0_u9_ch_am1[13] ) );
INV_X4 _u0_u9_U99  ( .A(1'b0), .ZN(_u0_u9_ch_am1[12] ) );
INV_X4 _u0_u9_U97  ( .A(1'b0), .ZN(_u0_u9_ch_am1[11] ) );
INV_X4 _u0_u9_U95  ( .A(1'b0), .ZN(_u0_u9_ch_am1[10] ) );
INV_X4 _u0_u9_U93  ( .A(1'b0), .ZN(_u0_u9_ch_am1[9] ) );
INV_X4 _u0_u9_U91  ( .A(1'b0), .ZN(_u0_u9_ch_am1[8] ) );
INV_X4 _u0_u9_U89  ( .A(1'b0), .ZN(_u0_u9_ch_am1[7] ) );
INV_X4 _u0_u9_U87  ( .A(1'b0), .ZN(_u0_u9_ch_am1[6] ) );
INV_X4 _u0_u9_U85  ( .A(1'b0), .ZN(_u0_u9_ch_am1[5] ) );
INV_X4 _u0_u9_U83  ( .A(1'b0), .ZN(_u0_u9_ch_am1[4] ) );
INV_X4 _u0_u9_U81  ( .A(1'b1), .ZN(_u0_u9_ch_am1[3] ) );
INV_X4 _u0_u9_U79  ( .A(1'b1), .ZN(_u0_u9_ch_am1[2] ) );
INV_X4 _u0_u9_U77  ( .A(1'b1), .ZN(_u0_u9_ch_am1[1] ) );
INV_X4 _u0_u9_U75  ( .A(1'b1), .ZN(_u0_u9_ch_am1[0] ) );
INV_X4 _u0_u9_U73  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[31] ) );
INV_X4 _u0_u9_U71  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[30] ) );
INV_X4 _u0_u9_U69  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[29] ) );
INV_X4 _u0_u9_U67  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[28] ) );
INV_X4 _u0_u9_U65  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[27] ) );
INV_X4 _u0_u9_U63  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[26] ) );
INV_X4 _u0_u9_U61  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[25] ) );
INV_X4 _u0_u9_U59  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[24] ) );
INV_X4 _u0_u9_U57  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[23] ) );
INV_X4 _u0_u9_U55  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[22] ) );
INV_X4 _u0_u9_U53  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[21] ) );
INV_X4 _u0_u9_U51  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[20] ) );
INV_X4 _u0_u9_U49  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[19] ) );
INV_X4 _u0_u9_U47  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[18] ) );
INV_X4 _u0_u9_U45  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[17] ) );
INV_X4 _u0_u9_U43  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[16] ) );
INV_X4 _u0_u9_U41  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[15] ) );
INV_X4 _u0_u9_U39  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[14] ) );
INV_X4 _u0_u9_U37  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[13] ) );
INV_X4 _u0_u9_U35  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[12] ) );
INV_X4 _u0_u9_U33  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[11] ) );
INV_X4 _u0_u9_U31  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[10] ) );
INV_X4 _u0_u9_U29  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[9] ) );
INV_X4 _u0_u9_U27  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[8] ) );
INV_X4 _u0_u9_U25  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[7] ) );
INV_X4 _u0_u9_U23  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[6] ) );
INV_X4 _u0_u9_U21  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[5] ) );
INV_X4 _u0_u9_U19  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[4] ) );
INV_X4 _u0_u9_U17  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[3] ) );
INV_X4 _u0_u9_U15  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[2] ) );
INV_X4 _u0_u9_U13  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[1] ) );
INV_X4 _u0_u9_U11  ( .A(1'b1), .ZN(_u0_u9_sw_pointer[0] ) );
INV_X4 _u0_u9_U9  ( .A(1'b1), .ZN(_u0_u9_ch_stop ) );
INV_X4 _u0_u9_U7  ( .A(1'b1), .ZN(_u0_u9_ch_dis ) );
INV_X4 _u0_u9_U5  ( .A(1'b1), .ZN(_u0_u9_int ) );
INV_X4 _u0_u10_U585  ( .A(1'b1), .ZN(_u0_u10_pointer[31] ) );
INV_X4 _u0_u10_U583  ( .A(1'b1), .ZN(_u0_u10_pointer[30] ) );
INV_X4 _u0_u10_U581  ( .A(1'b1), .ZN(_u0_u10_pointer[29] ) );
INV_X4 _u0_u10_U579  ( .A(1'b1), .ZN(_u0_u10_pointer[28] ) );
INV_X4 _u0_u10_U577  ( .A(1'b1), .ZN(_u0_u10_pointer[27] ) );
INV_X4 _u0_u10_U575  ( .A(1'b1), .ZN(_u0_u10_pointer[26] ) );
INV_X4 _u0_u10_U573  ( .A(1'b1), .ZN(_u0_u10_pointer[25] ) );
INV_X4 _u0_u10_U571  ( .A(1'b1), .ZN(_u0_u10_pointer[24] ) );
INV_X4 _u0_u10_U569  ( .A(1'b1), .ZN(_u0_u10_pointer[23] ) );
INV_X4 _u0_u10_U567  ( .A(1'b1), .ZN(_u0_u10_pointer[22] ) );
INV_X4 _u0_u10_U565  ( .A(1'b1), .ZN(_u0_u10_pointer[21] ) );
INV_X4 _u0_u10_U563  ( .A(1'b1), .ZN(_u0_u10_pointer[20] ) );
INV_X4 _u0_u10_U561  ( .A(1'b1), .ZN(_u0_u10_pointer[19] ) );
INV_X4 _u0_u10_U559  ( .A(1'b1), .ZN(_u0_u10_pointer[18] ) );
INV_X4 _u0_u10_U557  ( .A(1'b1), .ZN(_u0_u10_pointer[17] ) );
INV_X4 _u0_u10_U555  ( .A(1'b1), .ZN(_u0_u10_pointer[16] ) );
INV_X4 _u0_u10_U553  ( .A(1'b1), .ZN(_u0_u10_pointer[15] ) );
INV_X4 _u0_u10_U551  ( .A(1'b1), .ZN(_u0_u10_pointer[14] ) );
INV_X4 _u0_u10_U549  ( .A(1'b1), .ZN(_u0_u10_pointer[13] ) );
INV_X4 _u0_u10_U547  ( .A(1'b1), .ZN(_u0_u10_pointer[12] ) );
INV_X4 _u0_u10_U545  ( .A(1'b1), .ZN(_u0_u10_pointer[11] ) );
INV_X4 _u0_u10_U543  ( .A(1'b1), .ZN(_u0_u10_pointer[10] ) );
INV_X4 _u0_u10_U541  ( .A(1'b1), .ZN(_u0_u10_pointer[9] ) );
INV_X4 _u0_u10_U539  ( .A(1'b1), .ZN(_u0_u10_pointer[8] ) );
INV_X4 _u0_u10_U537  ( .A(1'b1), .ZN(_u0_u10_pointer[7] ) );
INV_X4 _u0_u10_U535  ( .A(1'b1), .ZN(_u0_u10_pointer[6] ) );
INV_X4 _u0_u10_U533  ( .A(1'b1), .ZN(_u0_u10_pointer[5] ) );
INV_X4 _u0_u10_U531  ( .A(1'b1), .ZN(_u0_u10_pointer[4] ) );
INV_X4 _u0_u10_U529  ( .A(1'b1), .ZN(_u0_u10_pointer[3] ) );
INV_X4 _u0_u10_U527  ( .A(1'b1), .ZN(_u0_u10_pointer[2] ) );
INV_X4 _u0_u10_U525  ( .A(1'b1), .ZN(_u0_u10_pointer[1] ) );
INV_X4 _u0_u10_U523  ( .A(1'b1), .ZN(_u0_u10_pointer[0] ) );
INV_X4 _u0_u10_U521  ( .A(1'b1), .ZN(_u0_u10_pointer_s[31] ) );
INV_X4 _u0_u10_U519  ( .A(1'b1), .ZN(_u0_u10_pointer_s[30] ) );
INV_X4 _u0_u10_U517  ( .A(1'b1), .ZN(_u0_u10_pointer_s[29] ) );
INV_X4 _u0_u10_U515  ( .A(1'b1), .ZN(_u0_u10_pointer_s[28] ) );
INV_X4 _u0_u10_U513  ( .A(1'b1), .ZN(_u0_u10_pointer_s[27] ) );
INV_X4 _u0_u10_U511  ( .A(1'b1), .ZN(_u0_u10_pointer_s[26] ) );
INV_X4 _u0_u10_U509  ( .A(1'b1), .ZN(_u0_u10_pointer_s[25] ) );
INV_X4 _u0_u10_U507  ( .A(1'b1), .ZN(_u0_u10_pointer_s[24] ) );
INV_X4 _u0_u10_U505  ( .A(1'b1), .ZN(_u0_u10_pointer_s[23] ) );
INV_X4 _u0_u10_U503  ( .A(1'b1), .ZN(_u0_u10_pointer_s[22] ) );
INV_X4 _u0_u10_U501  ( .A(1'b1), .ZN(_u0_u10_pointer_s[21] ) );
INV_X4 _u0_u10_U499  ( .A(1'b1), .ZN(_u0_u10_pointer_s[20] ) );
INV_X4 _u0_u10_U497  ( .A(1'b1), .ZN(_u0_u10_pointer_s[19] ) );
INV_X4 _u0_u10_U495  ( .A(1'b1), .ZN(_u0_u10_pointer_s[18] ) );
INV_X4 _u0_u10_U493  ( .A(1'b1), .ZN(_u0_u10_pointer_s[17] ) );
INV_X4 _u0_u10_U491  ( .A(1'b1), .ZN(_u0_u10_pointer_s[16] ) );
INV_X4 _u0_u10_U489  ( .A(1'b1), .ZN(_u0_u10_pointer_s[15] ) );
INV_X4 _u0_u10_U487  ( .A(1'b1), .ZN(_u0_u10_pointer_s[14] ) );
INV_X4 _u0_u10_U485  ( .A(1'b1), .ZN(_u0_u10_pointer_s[13] ) );
INV_X4 _u0_u10_U483  ( .A(1'b1), .ZN(_u0_u10_pointer_s[12] ) );
INV_X4 _u0_u10_U481  ( .A(1'b1), .ZN(_u0_u10_pointer_s[11] ) );
INV_X4 _u0_u10_U479  ( .A(1'b1), .ZN(_u0_u10_pointer_s[10] ) );
INV_X4 _u0_u10_U477  ( .A(1'b1), .ZN(_u0_u10_pointer_s[9] ) );
INV_X4 _u0_u10_U475  ( .A(1'b1), .ZN(_u0_u10_pointer_s[8] ) );
INV_X4 _u0_u10_U473  ( .A(1'b1), .ZN(_u0_u10_pointer_s[7] ) );
INV_X4 _u0_u10_U471  ( .A(1'b1), .ZN(_u0_u10_pointer_s[6] ) );
INV_X4 _u0_u10_U469  ( .A(1'b1), .ZN(_u0_u10_pointer_s[5] ) );
INV_X4 _u0_u10_U467  ( .A(1'b1), .ZN(_u0_u10_pointer_s[4] ) );
INV_X4 _u0_u10_U465  ( .A(1'b1), .ZN(_u0_u10_pointer_s[3] ) );
INV_X4 _u0_u10_U463  ( .A(1'b1), .ZN(_u0_u10_pointer_s[2] ) );
INV_X4 _u0_u10_U461  ( .A(1'b1), .ZN(_u0_u10_pointer_s[1] ) );
INV_X4 _u0_u10_U459  ( .A(1'b1), .ZN(_u0_u10_pointer_s[0] ) );
INV_X4 _u0_u10_U457  ( .A(1'b1), .ZN(_u0_u10_ch_csr[31] ) );
INV_X4 _u0_u10_U455  ( .A(1'b1), .ZN(_u0_u10_ch_csr[30] ) );
INV_X4 _u0_u10_U453  ( .A(1'b1), .ZN(_u0_u10_ch_csr[29] ) );
INV_X4 _u0_u10_U451  ( .A(1'b1), .ZN(_u0_u10_ch_csr[28] ) );
INV_X4 _u0_u10_U449  ( .A(1'b1), .ZN(_u0_u10_ch_csr[27] ) );
INV_X4 _u0_u10_U447  ( .A(1'b1), .ZN(_u0_u10_ch_csr[26] ) );
INV_X4 _u0_u10_U445  ( .A(1'b1), .ZN(_u0_u10_ch_csr[25] ) );
INV_X4 _u0_u10_U443  ( .A(1'b1), .ZN(_u0_u10_ch_csr[24] ) );
INV_X4 _u0_u10_U441  ( .A(1'b1), .ZN(_u0_u10_ch_csr[23] ) );
INV_X4 _u0_u10_U439  ( .A(1'b1), .ZN(_u0_u10_ch_csr[22] ) );
INV_X4 _u0_u10_U437  ( .A(1'b1), .ZN(_u0_u10_ch_csr[21] ) );
INV_X4 _u0_u10_U435  ( .A(1'b1), .ZN(_u0_u10_ch_csr[20] ) );
INV_X4 _u0_u10_U433  ( .A(1'b1), .ZN(_u0_u10_ch_csr[19] ) );
INV_X4 _u0_u10_U431  ( .A(1'b1), .ZN(_u0_u10_ch_csr[18] ) );
INV_X4 _u0_u10_U429  ( .A(1'b1), .ZN(_u0_u10_ch_csr[17] ) );
INV_X4 _u0_u10_U427  ( .A(1'b1), .ZN(_u0_u10_ch_csr[16] ) );
INV_X4 _u0_u10_U425  ( .A(1'b1), .ZN(_u0_u10_ch_csr[15] ) );
INV_X4 _u0_u10_U423  ( .A(1'b1), .ZN(_u0_u10_ch_csr[14] ) );
INV_X4 _u0_u10_U421  ( .A(1'b1), .ZN(_u0_u10_ch_csr[13] ) );
INV_X4 _u0_u10_U419  ( .A(1'b1), .ZN(_u0_u10_ch_csr[12] ) );
INV_X4 _u0_u10_U417  ( .A(1'b1), .ZN(_u0_u10_ch_csr[11] ) );
INV_X4 _u0_u10_U415  ( .A(1'b1), .ZN(_u0_u10_ch_csr[10] ) );
INV_X4 _u0_u10_U413  ( .A(1'b1), .ZN(_u0_u10_ch_csr[9] ) );
INV_X4 _u0_u10_U411  ( .A(1'b1), .ZN(_u0_u10_ch_csr[8] ) );
INV_X4 _u0_u10_U409  ( .A(1'b1), .ZN(_u0_u10_ch_csr[7] ) );
INV_X4 _u0_u10_U407  ( .A(1'b1), .ZN(_u0_u10_ch_csr[6] ) );
INV_X4 _u0_u10_U405  ( .A(1'b1), .ZN(_u0_u10_ch_csr[5] ) );
INV_X4 _u0_u10_U403  ( .A(1'b1), .ZN(_u0_u10_ch_csr[4] ) );
INV_X4 _u0_u10_U401  ( .A(1'b1), .ZN(_u0_u10_ch_csr[3] ) );
INV_X4 _u0_u10_U399  ( .A(1'b1), .ZN(_u0_u10_ch_csr[2] ) );
INV_X4 _u0_u10_U397  ( .A(1'b1), .ZN(_u0_u10_ch_csr[1] ) );
INV_X4 _u0_u10_U395  ( .A(1'b1), .ZN(_u0_u10_ch_csr[0] ) );
INV_X4 _u0_u10_U393  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[31] ) );
INV_X4 _u0_u10_U391  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[30] ) );
INV_X4 _u0_u10_U389  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[29] ) );
INV_X4 _u0_u10_U387  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[28] ) );
INV_X4 _u0_u10_U385  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[27] ) );
INV_X4 _u0_u10_U383  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[26] ) );
INV_X4 _u0_u10_U381  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[25] ) );
INV_X4 _u0_u10_U379  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[24] ) );
INV_X4 _u0_u10_U377  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[23] ) );
INV_X4 _u0_u10_U375  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[22] ) );
INV_X4 _u0_u10_U373  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[21] ) );
INV_X4 _u0_u10_U371  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[20] ) );
INV_X4 _u0_u10_U369  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[19] ) );
INV_X4 _u0_u10_U367  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[18] ) );
INV_X4 _u0_u10_U365  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[17] ) );
INV_X4 _u0_u10_U363  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[16] ) );
INV_X4 _u0_u10_U361  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[15] ) );
INV_X4 _u0_u10_U359  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[14] ) );
INV_X4 _u0_u10_U357  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[13] ) );
INV_X4 _u0_u10_U355  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[12] ) );
INV_X4 _u0_u10_U353  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[11] ) );
INV_X4 _u0_u10_U351  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[10] ) );
INV_X4 _u0_u10_U349  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[9] ) );
INV_X4 _u0_u10_U347  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[8] ) );
INV_X4 _u0_u10_U345  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[7] ) );
INV_X4 _u0_u10_U343  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[6] ) );
INV_X4 _u0_u10_U341  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[5] ) );
INV_X4 _u0_u10_U339  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[4] ) );
INV_X4 _u0_u10_U337  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[3] ) );
INV_X4 _u0_u10_U335  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[2] ) );
INV_X4 _u0_u10_U333  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[1] ) );
INV_X4 _u0_u10_U331  ( .A(1'b1), .ZN(_u0_u10_ch_txsz[0] ) );
INV_X4 _u0_u10_U329  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[31] ) );
INV_X4 _u0_u10_U327  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[30] ) );
INV_X4 _u0_u10_U325  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[29] ) );
INV_X4 _u0_u10_U323  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[28] ) );
INV_X4 _u0_u10_U321  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[27] ) );
INV_X4 _u0_u10_U319  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[26] ) );
INV_X4 _u0_u10_U317  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[25] ) );
INV_X4 _u0_u10_U315  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[24] ) );
INV_X4 _u0_u10_U313  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[23] ) );
INV_X4 _u0_u10_U311  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[22] ) );
INV_X4 _u0_u10_U309  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[21] ) );
INV_X4 _u0_u10_U307  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[20] ) );
INV_X4 _u0_u10_U305  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[19] ) );
INV_X4 _u0_u10_U303  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[18] ) );
INV_X4 _u0_u10_U301  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[17] ) );
INV_X4 _u0_u10_U299  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[16] ) );
INV_X4 _u0_u10_U297  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[15] ) );
INV_X4 _u0_u10_U295  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[14] ) );
INV_X4 _u0_u10_U293  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[13] ) );
INV_X4 _u0_u10_U291  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[12] ) );
INV_X4 _u0_u10_U289  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[11] ) );
INV_X4 _u0_u10_U287  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[10] ) );
INV_X4 _u0_u10_U285  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[9] ) );
INV_X4 _u0_u10_U283  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[8] ) );
INV_X4 _u0_u10_U281  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[7] ) );
INV_X4 _u0_u10_U279  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[6] ) );
INV_X4 _u0_u10_U277  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[5] ) );
INV_X4 _u0_u10_U275  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[4] ) );
INV_X4 _u0_u10_U273  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[3] ) );
INV_X4 _u0_u10_U271  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[2] ) );
INV_X4 _u0_u10_U269  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[1] ) );
INV_X4 _u0_u10_U267  ( .A(1'b1), .ZN(_u0_u10_ch_adr0[0] ) );
INV_X4 _u0_u10_U265  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[31] ) );
INV_X4 _u0_u10_U263  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[30] ) );
INV_X4 _u0_u10_U261  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[29] ) );
INV_X4 _u0_u10_U259  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[28] ) );
INV_X4 _u0_u10_U257  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[27] ) );
INV_X4 _u0_u10_U255  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[26] ) );
INV_X4 _u0_u10_U253  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[25] ) );
INV_X4 _u0_u10_U251  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[24] ) );
INV_X4 _u0_u10_U249  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[23] ) );
INV_X4 _u0_u10_U247  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[22] ) );
INV_X4 _u0_u10_U245  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[21] ) );
INV_X4 _u0_u10_U243  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[20] ) );
INV_X4 _u0_u10_U241  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[19] ) );
INV_X4 _u0_u10_U239  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[18] ) );
INV_X4 _u0_u10_U237  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[17] ) );
INV_X4 _u0_u10_U235  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[16] ) );
INV_X4 _u0_u10_U233  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[15] ) );
INV_X4 _u0_u10_U231  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[14] ) );
INV_X4 _u0_u10_U229  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[13] ) );
INV_X4 _u0_u10_U227  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[12] ) );
INV_X4 _u0_u10_U225  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[11] ) );
INV_X4 _u0_u10_U223  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[10] ) );
INV_X4 _u0_u10_U221  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[9] ) );
INV_X4 _u0_u10_U219  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[8] ) );
INV_X4 _u0_u10_U217  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[7] ) );
INV_X4 _u0_u10_U215  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[6] ) );
INV_X4 _u0_u10_U213  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[5] ) );
INV_X4 _u0_u10_U211  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[4] ) );
INV_X4 _u0_u10_U209  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[3] ) );
INV_X4 _u0_u10_U207  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[2] ) );
INV_X4 _u0_u10_U205  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[1] ) );
INV_X4 _u0_u10_U203  ( .A(1'b1), .ZN(_u0_u10_ch_adr1[0] ) );
INV_X4 _u0_u10_U201  ( .A(1'b0), .ZN(_u0_u10_ch_am0[31] ) );
INV_X4 _u0_u10_U199  ( .A(1'b0), .ZN(_u0_u10_ch_am0[30] ) );
INV_X4 _u0_u10_U197  ( .A(1'b0), .ZN(_u0_u10_ch_am0[29] ) );
INV_X4 _u0_u10_U195  ( .A(1'b0), .ZN(_u0_u10_ch_am0[28] ) );
INV_X4 _u0_u10_U193  ( .A(1'b0), .ZN(_u0_u10_ch_am0[27] ) );
INV_X4 _u0_u10_U191  ( .A(1'b0), .ZN(_u0_u10_ch_am0[26] ) );
INV_X4 _u0_u10_U189  ( .A(1'b0), .ZN(_u0_u10_ch_am0[25] ) );
INV_X4 _u0_u10_U187  ( .A(1'b0), .ZN(_u0_u10_ch_am0[24] ) );
INV_X4 _u0_u10_U185  ( .A(1'b0), .ZN(_u0_u10_ch_am0[23] ) );
INV_X4 _u0_u10_U183  ( .A(1'b0), .ZN(_u0_u10_ch_am0[22] ) );
INV_X4 _u0_u10_U181  ( .A(1'b0), .ZN(_u0_u10_ch_am0[21] ) );
INV_X4 _u0_u10_U179  ( .A(1'b0), .ZN(_u0_u10_ch_am0[20] ) );
INV_X4 _u0_u10_U177  ( .A(1'b0), .ZN(_u0_u10_ch_am0[19] ) );
INV_X4 _u0_u10_U175  ( .A(1'b0), .ZN(_u0_u10_ch_am0[18] ) );
INV_X4 _u0_u10_U173  ( .A(1'b0), .ZN(_u0_u10_ch_am0[17] ) );
INV_X4 _u0_u10_U171  ( .A(1'b0), .ZN(_u0_u10_ch_am0[16] ) );
INV_X4 _u0_u10_U169  ( .A(1'b0), .ZN(_u0_u10_ch_am0[15] ) );
INV_X4 _u0_u10_U167  ( .A(1'b0), .ZN(_u0_u10_ch_am0[14] ) );
INV_X4 _u0_u10_U165  ( .A(1'b0), .ZN(_u0_u10_ch_am0[13] ) );
INV_X4 _u0_u10_U163  ( .A(1'b0), .ZN(_u0_u10_ch_am0[12] ) );
INV_X4 _u0_u10_U161  ( .A(1'b0), .ZN(_u0_u10_ch_am0[11] ) );
INV_X4 _u0_u10_U159  ( .A(1'b0), .ZN(_u0_u10_ch_am0[10] ) );
INV_X4 _u0_u10_U157  ( .A(1'b0), .ZN(_u0_u10_ch_am0[9] ) );
INV_X4 _u0_u10_U155  ( .A(1'b0), .ZN(_u0_u10_ch_am0[8] ) );
INV_X4 _u0_u10_U153  ( .A(1'b0), .ZN(_u0_u10_ch_am0[7] ) );
INV_X4 _u0_u10_U151  ( .A(1'b0), .ZN(_u0_u10_ch_am0[6] ) );
INV_X4 _u0_u10_U149  ( .A(1'b0), .ZN(_u0_u10_ch_am0[5] ) );
INV_X4 _u0_u10_U147  ( .A(1'b0), .ZN(_u0_u10_ch_am0[4] ) );
INV_X4 _u0_u10_U145  ( .A(1'b1), .ZN(_u0_u10_ch_am0[3] ) );
INV_X4 _u0_u10_U143  ( .A(1'b1), .ZN(_u0_u10_ch_am0[2] ) );
INV_X4 _u0_u10_U141  ( .A(1'b1), .ZN(_u0_u10_ch_am0[1] ) );
INV_X4 _u0_u10_U139  ( .A(1'b1), .ZN(_u0_u10_ch_am0[0] ) );
INV_X4 _u0_u10_U137  ( .A(1'b0), .ZN(_u0_u10_ch_am1[31] ) );
INV_X4 _u0_u10_U135  ( .A(1'b0), .ZN(_u0_u10_ch_am1[30] ) );
INV_X4 _u0_u10_U133  ( .A(1'b0), .ZN(_u0_u10_ch_am1[29] ) );
INV_X4 _u0_u10_U131  ( .A(1'b0), .ZN(_u0_u10_ch_am1[28] ) );
INV_X4 _u0_u10_U129  ( .A(1'b0), .ZN(_u0_u10_ch_am1[27] ) );
INV_X4 _u0_u10_U127  ( .A(1'b0), .ZN(_u0_u10_ch_am1[26] ) );
INV_X4 _u0_u10_U125  ( .A(1'b0), .ZN(_u0_u10_ch_am1[25] ) );
INV_X4 _u0_u10_U123  ( .A(1'b0), .ZN(_u0_u10_ch_am1[24] ) );
INV_X4 _u0_u10_U121  ( .A(1'b0), .ZN(_u0_u10_ch_am1[23] ) );
INV_X4 _u0_u10_U119  ( .A(1'b0), .ZN(_u0_u10_ch_am1[22] ) );
INV_X4 _u0_u10_U117  ( .A(1'b0), .ZN(_u0_u10_ch_am1[21] ) );
INV_X4 _u0_u10_U115  ( .A(1'b0), .ZN(_u0_u10_ch_am1[20] ) );
INV_X4 _u0_u10_U113  ( .A(1'b0), .ZN(_u0_u10_ch_am1[19] ) );
INV_X4 _u0_u10_U111  ( .A(1'b0), .ZN(_u0_u10_ch_am1[18] ) );
INV_X4 _u0_u10_U109  ( .A(1'b0), .ZN(_u0_u10_ch_am1[17] ) );
INV_X4 _u0_u10_U107  ( .A(1'b0), .ZN(_u0_u10_ch_am1[16] ) );
INV_X4 _u0_u10_U105  ( .A(1'b0), .ZN(_u0_u10_ch_am1[15] ) );
INV_X4 _u0_u10_U103  ( .A(1'b0), .ZN(_u0_u10_ch_am1[14] ) );
INV_X4 _u0_u10_U101  ( .A(1'b0), .ZN(_u0_u10_ch_am1[13] ) );
INV_X4 _u0_u10_U99  ( .A(1'b0), .ZN(_u0_u10_ch_am1[12] ) );
INV_X4 _u0_u10_U97  ( .A(1'b0), .ZN(_u0_u10_ch_am1[11] ) );
INV_X4 _u0_u10_U95  ( .A(1'b0), .ZN(_u0_u10_ch_am1[10] ) );
INV_X4 _u0_u10_U93  ( .A(1'b0), .ZN(_u0_u10_ch_am1[9] ) );
INV_X4 _u0_u10_U91  ( .A(1'b0), .ZN(_u0_u10_ch_am1[8] ) );
INV_X4 _u0_u10_U89  ( .A(1'b0), .ZN(_u0_u10_ch_am1[7] ) );
INV_X4 _u0_u10_U87  ( .A(1'b0), .ZN(_u0_u10_ch_am1[6] ) );
INV_X4 _u0_u10_U85  ( .A(1'b0), .ZN(_u0_u10_ch_am1[5] ) );
INV_X4 _u0_u10_U83  ( .A(1'b0), .ZN(_u0_u10_ch_am1[4] ) );
INV_X4 _u0_u10_U81  ( .A(1'b1), .ZN(_u0_u10_ch_am1[3] ) );
INV_X4 _u0_u10_U79  ( .A(1'b1), .ZN(_u0_u10_ch_am1[2] ) );
INV_X4 _u0_u10_U77  ( .A(1'b1), .ZN(_u0_u10_ch_am1[1] ) );
INV_X4 _u0_u10_U75  ( .A(1'b1), .ZN(_u0_u10_ch_am1[0] ) );
INV_X4 _u0_u10_U73  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[31] ) );
INV_X4 _u0_u10_U71  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[30] ) );
INV_X4 _u0_u10_U69  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[29] ) );
INV_X4 _u0_u10_U67  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[28] ) );
INV_X4 _u0_u10_U65  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[27] ) );
INV_X4 _u0_u10_U63  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[26] ) );
INV_X4 _u0_u10_U61  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[25] ) );
INV_X4 _u0_u10_U59  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[24] ) );
INV_X4 _u0_u10_U57  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[23] ) );
INV_X4 _u0_u10_U55  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[22] ) );
INV_X4 _u0_u10_U53  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[21] ) );
INV_X4 _u0_u10_U51  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[20] ) );
INV_X4 _u0_u10_U49  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[19] ) );
INV_X4 _u0_u10_U47  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[18] ) );
INV_X4 _u0_u10_U45  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[17] ) );
INV_X4 _u0_u10_U43  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[16] ) );
INV_X4 _u0_u10_U41  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[15] ) );
INV_X4 _u0_u10_U39  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[14] ) );
INV_X4 _u0_u10_U37  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[13] ) );
INV_X4 _u0_u10_U35  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[12] ) );
INV_X4 _u0_u10_U33  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[11] ) );
INV_X4 _u0_u10_U31  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[10] ) );
INV_X4 _u0_u10_U29  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[9] ) );
INV_X4 _u0_u10_U27  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[8] ) );
INV_X4 _u0_u10_U25  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[7] ) );
INV_X4 _u0_u10_U23  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[6] ) );
INV_X4 _u0_u10_U21  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[5] ) );
INV_X4 _u0_u10_U19  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[4] ) );
INV_X4 _u0_u10_U17  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[3] ) );
INV_X4 _u0_u10_U15  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[2] ) );
INV_X4 _u0_u10_U13  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[1] ) );
INV_X4 _u0_u10_U11  ( .A(1'b1), .ZN(_u0_u10_sw_pointer[0] ) );
INV_X4 _u0_u10_U9  ( .A(1'b1), .ZN(_u0_u10_ch_stop ) );
INV_X4 _u0_u10_U7  ( .A(1'b1), .ZN(_u0_u10_ch_dis ) );
INV_X4 _u0_u10_U5  ( .A(1'b1), .ZN(_u0_u10_int ) );
INV_X4 _u0_u11_U585  ( .A(1'b1), .ZN(_u0_u11_pointer[31] ) );
INV_X4 _u0_u11_U583  ( .A(1'b1), .ZN(_u0_u11_pointer[30] ) );
INV_X4 _u0_u11_U581  ( .A(1'b1), .ZN(_u0_u11_pointer[29] ) );
INV_X4 _u0_u11_U579  ( .A(1'b1), .ZN(_u0_u11_pointer[28] ) );
INV_X4 _u0_u11_U577  ( .A(1'b1), .ZN(_u0_u11_pointer[27] ) );
INV_X4 _u0_u11_U575  ( .A(1'b1), .ZN(_u0_u11_pointer[26] ) );
INV_X4 _u0_u11_U573  ( .A(1'b1), .ZN(_u0_u11_pointer[25] ) );
INV_X4 _u0_u11_U571  ( .A(1'b1), .ZN(_u0_u11_pointer[24] ) );
INV_X4 _u0_u11_U569  ( .A(1'b1), .ZN(_u0_u11_pointer[23] ) );
INV_X4 _u0_u11_U567  ( .A(1'b1), .ZN(_u0_u11_pointer[22] ) );
INV_X4 _u0_u11_U565  ( .A(1'b1), .ZN(_u0_u11_pointer[21] ) );
INV_X4 _u0_u11_U563  ( .A(1'b1), .ZN(_u0_u11_pointer[20] ) );
INV_X4 _u0_u11_U561  ( .A(1'b1), .ZN(_u0_u11_pointer[19] ) );
INV_X4 _u0_u11_U559  ( .A(1'b1), .ZN(_u0_u11_pointer[18] ) );
INV_X4 _u0_u11_U557  ( .A(1'b1), .ZN(_u0_u11_pointer[17] ) );
INV_X4 _u0_u11_U555  ( .A(1'b1), .ZN(_u0_u11_pointer[16] ) );
INV_X4 _u0_u11_U553  ( .A(1'b1), .ZN(_u0_u11_pointer[15] ) );
INV_X4 _u0_u11_U551  ( .A(1'b1), .ZN(_u0_u11_pointer[14] ) );
INV_X4 _u0_u11_U549  ( .A(1'b1), .ZN(_u0_u11_pointer[13] ) );
INV_X4 _u0_u11_U547  ( .A(1'b1), .ZN(_u0_u11_pointer[12] ) );
INV_X4 _u0_u11_U545  ( .A(1'b1), .ZN(_u0_u11_pointer[11] ) );
INV_X4 _u0_u11_U543  ( .A(1'b1), .ZN(_u0_u11_pointer[10] ) );
INV_X4 _u0_u11_U541  ( .A(1'b1), .ZN(_u0_u11_pointer[9] ) );
INV_X4 _u0_u11_U539  ( .A(1'b1), .ZN(_u0_u11_pointer[8] ) );
INV_X4 _u0_u11_U537  ( .A(1'b1), .ZN(_u0_u11_pointer[7] ) );
INV_X4 _u0_u11_U535  ( .A(1'b1), .ZN(_u0_u11_pointer[6] ) );
INV_X4 _u0_u11_U533  ( .A(1'b1), .ZN(_u0_u11_pointer[5] ) );
INV_X4 _u0_u11_U531  ( .A(1'b1), .ZN(_u0_u11_pointer[4] ) );
INV_X4 _u0_u11_U529  ( .A(1'b1), .ZN(_u0_u11_pointer[3] ) );
INV_X4 _u0_u11_U527  ( .A(1'b1), .ZN(_u0_u11_pointer[2] ) );
INV_X4 _u0_u11_U525  ( .A(1'b1), .ZN(_u0_u11_pointer[1] ) );
INV_X4 _u0_u11_U523  ( .A(1'b1), .ZN(_u0_u11_pointer[0] ) );
INV_X4 _u0_u11_U521  ( .A(1'b1), .ZN(_u0_u11_pointer_s[31] ) );
INV_X4 _u0_u11_U519  ( .A(1'b1), .ZN(_u0_u11_pointer_s[30] ) );
INV_X4 _u0_u11_U517  ( .A(1'b1), .ZN(_u0_u11_pointer_s[29] ) );
INV_X4 _u0_u11_U515  ( .A(1'b1), .ZN(_u0_u11_pointer_s[28] ) );
INV_X4 _u0_u11_U513  ( .A(1'b1), .ZN(_u0_u11_pointer_s[27] ) );
INV_X4 _u0_u11_U511  ( .A(1'b1), .ZN(_u0_u11_pointer_s[26] ) );
INV_X4 _u0_u11_U509  ( .A(1'b1), .ZN(_u0_u11_pointer_s[25] ) );
INV_X4 _u0_u11_U507  ( .A(1'b1), .ZN(_u0_u11_pointer_s[24] ) );
INV_X4 _u0_u11_U505  ( .A(1'b1), .ZN(_u0_u11_pointer_s[23] ) );
INV_X4 _u0_u11_U503  ( .A(1'b1), .ZN(_u0_u11_pointer_s[22] ) );
INV_X4 _u0_u11_U501  ( .A(1'b1), .ZN(_u0_u11_pointer_s[21] ) );
INV_X4 _u0_u11_U499  ( .A(1'b1), .ZN(_u0_u11_pointer_s[20] ) );
INV_X4 _u0_u11_U497  ( .A(1'b1), .ZN(_u0_u11_pointer_s[19] ) );
INV_X4 _u0_u11_U495  ( .A(1'b1), .ZN(_u0_u11_pointer_s[18] ) );
INV_X4 _u0_u11_U493  ( .A(1'b1), .ZN(_u0_u11_pointer_s[17] ) );
INV_X4 _u0_u11_U491  ( .A(1'b1), .ZN(_u0_u11_pointer_s[16] ) );
INV_X4 _u0_u11_U489  ( .A(1'b1), .ZN(_u0_u11_pointer_s[15] ) );
INV_X4 _u0_u11_U487  ( .A(1'b1), .ZN(_u0_u11_pointer_s[14] ) );
INV_X4 _u0_u11_U485  ( .A(1'b1), .ZN(_u0_u11_pointer_s[13] ) );
INV_X4 _u0_u11_U483  ( .A(1'b1), .ZN(_u0_u11_pointer_s[12] ) );
INV_X4 _u0_u11_U481  ( .A(1'b1), .ZN(_u0_u11_pointer_s[11] ) );
INV_X4 _u0_u11_U479  ( .A(1'b1), .ZN(_u0_u11_pointer_s[10] ) );
INV_X4 _u0_u11_U477  ( .A(1'b1), .ZN(_u0_u11_pointer_s[9] ) );
INV_X4 _u0_u11_U475  ( .A(1'b1), .ZN(_u0_u11_pointer_s[8] ) );
INV_X4 _u0_u11_U473  ( .A(1'b1), .ZN(_u0_u11_pointer_s[7] ) );
INV_X4 _u0_u11_U471  ( .A(1'b1), .ZN(_u0_u11_pointer_s[6] ) );
INV_X4 _u0_u11_U469  ( .A(1'b1), .ZN(_u0_u11_pointer_s[5] ) );
INV_X4 _u0_u11_U467  ( .A(1'b1), .ZN(_u0_u11_pointer_s[4] ) );
INV_X4 _u0_u11_U465  ( .A(1'b1), .ZN(_u0_u11_pointer_s[3] ) );
INV_X4 _u0_u11_U463  ( .A(1'b1), .ZN(_u0_u11_pointer_s[2] ) );
INV_X4 _u0_u11_U461  ( .A(1'b1), .ZN(_u0_u11_pointer_s[1] ) );
INV_X4 _u0_u11_U459  ( .A(1'b1), .ZN(_u0_u11_pointer_s[0] ) );
INV_X4 _u0_u11_U457  ( .A(1'b1), .ZN(_u0_u11_ch_csr[31] ) );
INV_X4 _u0_u11_U455  ( .A(1'b1), .ZN(_u0_u11_ch_csr[30] ) );
INV_X4 _u0_u11_U453  ( .A(1'b1), .ZN(_u0_u11_ch_csr[29] ) );
INV_X4 _u0_u11_U451  ( .A(1'b1), .ZN(_u0_u11_ch_csr[28] ) );
INV_X4 _u0_u11_U449  ( .A(1'b1), .ZN(_u0_u11_ch_csr[27] ) );
INV_X4 _u0_u11_U447  ( .A(1'b1), .ZN(_u0_u11_ch_csr[26] ) );
INV_X4 _u0_u11_U445  ( .A(1'b1), .ZN(_u0_u11_ch_csr[25] ) );
INV_X4 _u0_u11_U443  ( .A(1'b1), .ZN(_u0_u11_ch_csr[24] ) );
INV_X4 _u0_u11_U441  ( .A(1'b1), .ZN(_u0_u11_ch_csr[23] ) );
INV_X4 _u0_u11_U439  ( .A(1'b1), .ZN(_u0_u11_ch_csr[22] ) );
INV_X4 _u0_u11_U437  ( .A(1'b1), .ZN(_u0_u11_ch_csr[21] ) );
INV_X4 _u0_u11_U435  ( .A(1'b1), .ZN(_u0_u11_ch_csr[20] ) );
INV_X4 _u0_u11_U433  ( .A(1'b1), .ZN(_u0_u11_ch_csr[19] ) );
INV_X4 _u0_u11_U431  ( .A(1'b1), .ZN(_u0_u11_ch_csr[18] ) );
INV_X4 _u0_u11_U429  ( .A(1'b1), .ZN(_u0_u11_ch_csr[17] ) );
INV_X4 _u0_u11_U427  ( .A(1'b1), .ZN(_u0_u11_ch_csr[16] ) );
INV_X4 _u0_u11_U425  ( .A(1'b1), .ZN(_u0_u11_ch_csr[15] ) );
INV_X4 _u0_u11_U423  ( .A(1'b1), .ZN(_u0_u11_ch_csr[14] ) );
INV_X4 _u0_u11_U421  ( .A(1'b1), .ZN(_u0_u11_ch_csr[13] ) );
INV_X4 _u0_u11_U419  ( .A(1'b1), .ZN(_u0_u11_ch_csr[12] ) );
INV_X4 _u0_u11_U417  ( .A(1'b1), .ZN(_u0_u11_ch_csr[11] ) );
INV_X4 _u0_u11_U415  ( .A(1'b1), .ZN(_u0_u11_ch_csr[10] ) );
INV_X4 _u0_u11_U413  ( .A(1'b1), .ZN(_u0_u11_ch_csr[9] ) );
INV_X4 _u0_u11_U411  ( .A(1'b1), .ZN(_u0_u11_ch_csr[8] ) );
INV_X4 _u0_u11_U409  ( .A(1'b1), .ZN(_u0_u11_ch_csr[7] ) );
INV_X4 _u0_u11_U407  ( .A(1'b1), .ZN(_u0_u11_ch_csr[6] ) );
INV_X4 _u0_u11_U405  ( .A(1'b1), .ZN(_u0_u11_ch_csr[5] ) );
INV_X4 _u0_u11_U403  ( .A(1'b1), .ZN(_u0_u11_ch_csr[4] ) );
INV_X4 _u0_u11_U401  ( .A(1'b1), .ZN(_u0_u11_ch_csr[3] ) );
INV_X4 _u0_u11_U399  ( .A(1'b1), .ZN(_u0_u11_ch_csr[2] ) );
INV_X4 _u0_u11_U397  ( .A(1'b1), .ZN(_u0_u11_ch_csr[1] ) );
INV_X4 _u0_u11_U395  ( .A(1'b1), .ZN(_u0_u11_ch_csr[0] ) );
INV_X4 _u0_u11_U393  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[31] ) );
INV_X4 _u0_u11_U391  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[30] ) );
INV_X4 _u0_u11_U389  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[29] ) );
INV_X4 _u0_u11_U387  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[28] ) );
INV_X4 _u0_u11_U385  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[27] ) );
INV_X4 _u0_u11_U383  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[26] ) );
INV_X4 _u0_u11_U381  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[25] ) );
INV_X4 _u0_u11_U379  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[24] ) );
INV_X4 _u0_u11_U377  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[23] ) );
INV_X4 _u0_u11_U375  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[22] ) );
INV_X4 _u0_u11_U373  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[21] ) );
INV_X4 _u0_u11_U371  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[20] ) );
INV_X4 _u0_u11_U369  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[19] ) );
INV_X4 _u0_u11_U367  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[18] ) );
INV_X4 _u0_u11_U365  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[17] ) );
INV_X4 _u0_u11_U363  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[16] ) );
INV_X4 _u0_u11_U361  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[15] ) );
INV_X4 _u0_u11_U359  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[14] ) );
INV_X4 _u0_u11_U357  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[13] ) );
INV_X4 _u0_u11_U355  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[12] ) );
INV_X4 _u0_u11_U353  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[11] ) );
INV_X4 _u0_u11_U351  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[10] ) );
INV_X4 _u0_u11_U349  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[9] ) );
INV_X4 _u0_u11_U347  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[8] ) );
INV_X4 _u0_u11_U345  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[7] ) );
INV_X4 _u0_u11_U343  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[6] ) );
INV_X4 _u0_u11_U341  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[5] ) );
INV_X4 _u0_u11_U339  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[4] ) );
INV_X4 _u0_u11_U337  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[3] ) );
INV_X4 _u0_u11_U335  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[2] ) );
INV_X4 _u0_u11_U333  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[1] ) );
INV_X4 _u0_u11_U331  ( .A(1'b1), .ZN(_u0_u11_ch_txsz[0] ) );
INV_X4 _u0_u11_U329  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[31] ) );
INV_X4 _u0_u11_U327  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[30] ) );
INV_X4 _u0_u11_U325  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[29] ) );
INV_X4 _u0_u11_U323  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[28] ) );
INV_X4 _u0_u11_U321  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[27] ) );
INV_X4 _u0_u11_U319  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[26] ) );
INV_X4 _u0_u11_U317  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[25] ) );
INV_X4 _u0_u11_U315  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[24] ) );
INV_X4 _u0_u11_U313  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[23] ) );
INV_X4 _u0_u11_U311  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[22] ) );
INV_X4 _u0_u11_U309  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[21] ) );
INV_X4 _u0_u11_U307  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[20] ) );
INV_X4 _u0_u11_U305  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[19] ) );
INV_X4 _u0_u11_U303  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[18] ) );
INV_X4 _u0_u11_U301  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[17] ) );
INV_X4 _u0_u11_U299  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[16] ) );
INV_X4 _u0_u11_U297  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[15] ) );
INV_X4 _u0_u11_U295  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[14] ) );
INV_X4 _u0_u11_U293  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[13] ) );
INV_X4 _u0_u11_U291  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[12] ) );
INV_X4 _u0_u11_U289  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[11] ) );
INV_X4 _u0_u11_U287  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[10] ) );
INV_X4 _u0_u11_U285  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[9] ) );
INV_X4 _u0_u11_U283  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[8] ) );
INV_X4 _u0_u11_U281  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[7] ) );
INV_X4 _u0_u11_U279  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[6] ) );
INV_X4 _u0_u11_U277  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[5] ) );
INV_X4 _u0_u11_U275  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[4] ) );
INV_X4 _u0_u11_U273  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[3] ) );
INV_X4 _u0_u11_U271  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[2] ) );
INV_X4 _u0_u11_U269  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[1] ) );
INV_X4 _u0_u11_U267  ( .A(1'b1), .ZN(_u0_u11_ch_adr0[0] ) );
INV_X4 _u0_u11_U265  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[31] ) );
INV_X4 _u0_u11_U263  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[30] ) );
INV_X4 _u0_u11_U261  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[29] ) );
INV_X4 _u0_u11_U259  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[28] ) );
INV_X4 _u0_u11_U257  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[27] ) );
INV_X4 _u0_u11_U255  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[26] ) );
INV_X4 _u0_u11_U253  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[25] ) );
INV_X4 _u0_u11_U251  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[24] ) );
INV_X4 _u0_u11_U249  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[23] ) );
INV_X4 _u0_u11_U247  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[22] ) );
INV_X4 _u0_u11_U245  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[21] ) );
INV_X4 _u0_u11_U243  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[20] ) );
INV_X4 _u0_u11_U241  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[19] ) );
INV_X4 _u0_u11_U239  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[18] ) );
INV_X4 _u0_u11_U237  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[17] ) );
INV_X4 _u0_u11_U235  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[16] ) );
INV_X4 _u0_u11_U233  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[15] ) );
INV_X4 _u0_u11_U231  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[14] ) );
INV_X4 _u0_u11_U229  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[13] ) );
INV_X4 _u0_u11_U227  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[12] ) );
INV_X4 _u0_u11_U225  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[11] ) );
INV_X4 _u0_u11_U223  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[10] ) );
INV_X4 _u0_u11_U221  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[9] ) );
INV_X4 _u0_u11_U219  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[8] ) );
INV_X4 _u0_u11_U217  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[7] ) );
INV_X4 _u0_u11_U215  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[6] ) );
INV_X4 _u0_u11_U213  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[5] ) );
INV_X4 _u0_u11_U211  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[4] ) );
INV_X4 _u0_u11_U209  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[3] ) );
INV_X4 _u0_u11_U207  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[2] ) );
INV_X4 _u0_u11_U205  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[1] ) );
INV_X4 _u0_u11_U203  ( .A(1'b1), .ZN(_u0_u11_ch_adr1[0] ) );
INV_X4 _u0_u11_U201  ( .A(1'b0), .ZN(_u0_u11_ch_am0[31] ) );
INV_X4 _u0_u11_U199  ( .A(1'b0), .ZN(_u0_u11_ch_am0[30] ) );
INV_X4 _u0_u11_U197  ( .A(1'b0), .ZN(_u0_u11_ch_am0[29] ) );
INV_X4 _u0_u11_U195  ( .A(1'b0), .ZN(_u0_u11_ch_am0[28] ) );
INV_X4 _u0_u11_U193  ( .A(1'b0), .ZN(_u0_u11_ch_am0[27] ) );
INV_X4 _u0_u11_U191  ( .A(1'b0), .ZN(_u0_u11_ch_am0[26] ) );
INV_X4 _u0_u11_U189  ( .A(1'b0), .ZN(_u0_u11_ch_am0[25] ) );
INV_X4 _u0_u11_U187  ( .A(1'b0), .ZN(_u0_u11_ch_am0[24] ) );
INV_X4 _u0_u11_U185  ( .A(1'b0), .ZN(_u0_u11_ch_am0[23] ) );
INV_X4 _u0_u11_U183  ( .A(1'b0), .ZN(_u0_u11_ch_am0[22] ) );
INV_X4 _u0_u11_U181  ( .A(1'b0), .ZN(_u0_u11_ch_am0[21] ) );
INV_X4 _u0_u11_U179  ( .A(1'b0), .ZN(_u0_u11_ch_am0[20] ) );
INV_X4 _u0_u11_U177  ( .A(1'b0), .ZN(_u0_u11_ch_am0[19] ) );
INV_X4 _u0_u11_U175  ( .A(1'b0), .ZN(_u0_u11_ch_am0[18] ) );
INV_X4 _u0_u11_U173  ( .A(1'b0), .ZN(_u0_u11_ch_am0[17] ) );
INV_X4 _u0_u11_U171  ( .A(1'b0), .ZN(_u0_u11_ch_am0[16] ) );
INV_X4 _u0_u11_U169  ( .A(1'b0), .ZN(_u0_u11_ch_am0[15] ) );
INV_X4 _u0_u11_U167  ( .A(1'b0), .ZN(_u0_u11_ch_am0[14] ) );
INV_X4 _u0_u11_U165  ( .A(1'b0), .ZN(_u0_u11_ch_am0[13] ) );
INV_X4 _u0_u11_U163  ( .A(1'b0), .ZN(_u0_u11_ch_am0[12] ) );
INV_X4 _u0_u11_U161  ( .A(1'b0), .ZN(_u0_u11_ch_am0[11] ) );
INV_X4 _u0_u11_U159  ( .A(1'b0), .ZN(_u0_u11_ch_am0[10] ) );
INV_X4 _u0_u11_U157  ( .A(1'b0), .ZN(_u0_u11_ch_am0[9] ) );
INV_X4 _u0_u11_U155  ( .A(1'b0), .ZN(_u0_u11_ch_am0[8] ) );
INV_X4 _u0_u11_U153  ( .A(1'b0), .ZN(_u0_u11_ch_am0[7] ) );
INV_X4 _u0_u11_U151  ( .A(1'b0), .ZN(_u0_u11_ch_am0[6] ) );
INV_X4 _u0_u11_U149  ( .A(1'b0), .ZN(_u0_u11_ch_am0[5] ) );
INV_X4 _u0_u11_U147  ( .A(1'b0), .ZN(_u0_u11_ch_am0[4] ) );
INV_X4 _u0_u11_U145  ( .A(1'b1), .ZN(_u0_u11_ch_am0[3] ) );
INV_X4 _u0_u11_U143  ( .A(1'b1), .ZN(_u0_u11_ch_am0[2] ) );
INV_X4 _u0_u11_U141  ( .A(1'b1), .ZN(_u0_u11_ch_am0[1] ) );
INV_X4 _u0_u11_U139  ( .A(1'b1), .ZN(_u0_u11_ch_am0[0] ) );
INV_X4 _u0_u11_U137  ( .A(1'b0), .ZN(_u0_u11_ch_am1[31] ) );
INV_X4 _u0_u11_U135  ( .A(1'b0), .ZN(_u0_u11_ch_am1[30] ) );
INV_X4 _u0_u11_U133  ( .A(1'b0), .ZN(_u0_u11_ch_am1[29] ) );
INV_X4 _u0_u11_U131  ( .A(1'b0), .ZN(_u0_u11_ch_am1[28] ) );
INV_X4 _u0_u11_U129  ( .A(1'b0), .ZN(_u0_u11_ch_am1[27] ) );
INV_X4 _u0_u11_U127  ( .A(1'b0), .ZN(_u0_u11_ch_am1[26] ) );
INV_X4 _u0_u11_U125  ( .A(1'b0), .ZN(_u0_u11_ch_am1[25] ) );
INV_X4 _u0_u11_U123  ( .A(1'b0), .ZN(_u0_u11_ch_am1[24] ) );
INV_X4 _u0_u11_U121  ( .A(1'b0), .ZN(_u0_u11_ch_am1[23] ) );
INV_X4 _u0_u11_U119  ( .A(1'b0), .ZN(_u0_u11_ch_am1[22] ) );
INV_X4 _u0_u11_U117  ( .A(1'b0), .ZN(_u0_u11_ch_am1[21] ) );
INV_X4 _u0_u11_U115  ( .A(1'b0), .ZN(_u0_u11_ch_am1[20] ) );
INV_X4 _u0_u11_U113  ( .A(1'b0), .ZN(_u0_u11_ch_am1[19] ) );
INV_X4 _u0_u11_U111  ( .A(1'b0), .ZN(_u0_u11_ch_am1[18] ) );
INV_X4 _u0_u11_U109  ( .A(1'b0), .ZN(_u0_u11_ch_am1[17] ) );
INV_X4 _u0_u11_U107  ( .A(1'b0), .ZN(_u0_u11_ch_am1[16] ) );
INV_X4 _u0_u11_U105  ( .A(1'b0), .ZN(_u0_u11_ch_am1[15] ) );
INV_X4 _u0_u11_U103  ( .A(1'b0), .ZN(_u0_u11_ch_am1[14] ) );
INV_X4 _u0_u11_U101  ( .A(1'b0), .ZN(_u0_u11_ch_am1[13] ) );
INV_X4 _u0_u11_U99  ( .A(1'b0), .ZN(_u0_u11_ch_am1[12] ) );
INV_X4 _u0_u11_U97  ( .A(1'b0), .ZN(_u0_u11_ch_am1[11] ) );
INV_X4 _u0_u11_U95  ( .A(1'b0), .ZN(_u0_u11_ch_am1[10] ) );
INV_X4 _u0_u11_U93  ( .A(1'b0), .ZN(_u0_u11_ch_am1[9] ) );
INV_X4 _u0_u11_U91  ( .A(1'b0), .ZN(_u0_u11_ch_am1[8] ) );
INV_X4 _u0_u11_U89  ( .A(1'b0), .ZN(_u0_u11_ch_am1[7] ) );
INV_X4 _u0_u11_U87  ( .A(1'b0), .ZN(_u0_u11_ch_am1[6] ) );
INV_X4 _u0_u11_U85  ( .A(1'b0), .ZN(_u0_u11_ch_am1[5] ) );
INV_X4 _u0_u11_U83  ( .A(1'b0), .ZN(_u0_u11_ch_am1[4] ) );
INV_X4 _u0_u11_U81  ( .A(1'b1), .ZN(_u0_u11_ch_am1[3] ) );
INV_X4 _u0_u11_U79  ( .A(1'b1), .ZN(_u0_u11_ch_am1[2] ) );
INV_X4 _u0_u11_U77  ( .A(1'b1), .ZN(_u0_u11_ch_am1[1] ) );
INV_X4 _u0_u11_U75  ( .A(1'b1), .ZN(_u0_u11_ch_am1[0] ) );
INV_X4 _u0_u11_U73  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[31] ) );
INV_X4 _u0_u11_U71  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[30] ) );
INV_X4 _u0_u11_U69  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[29] ) );
INV_X4 _u0_u11_U67  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[28] ) );
INV_X4 _u0_u11_U65  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[27] ) );
INV_X4 _u0_u11_U63  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[26] ) );
INV_X4 _u0_u11_U61  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[25] ) );
INV_X4 _u0_u11_U59  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[24] ) );
INV_X4 _u0_u11_U57  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[23] ) );
INV_X4 _u0_u11_U55  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[22] ) );
INV_X4 _u0_u11_U53  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[21] ) );
INV_X4 _u0_u11_U51  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[20] ) );
INV_X4 _u0_u11_U49  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[19] ) );
INV_X4 _u0_u11_U47  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[18] ) );
INV_X4 _u0_u11_U45  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[17] ) );
INV_X4 _u0_u11_U43  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[16] ) );
INV_X4 _u0_u11_U41  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[15] ) );
INV_X4 _u0_u11_U39  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[14] ) );
INV_X4 _u0_u11_U37  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[13] ) );
INV_X4 _u0_u11_U35  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[12] ) );
INV_X4 _u0_u11_U33  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[11] ) );
INV_X4 _u0_u11_U31  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[10] ) );
INV_X4 _u0_u11_U29  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[9] ) );
INV_X4 _u0_u11_U27  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[8] ) );
INV_X4 _u0_u11_U25  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[7] ) );
INV_X4 _u0_u11_U23  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[6] ) );
INV_X4 _u0_u11_U21  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[5] ) );
INV_X4 _u0_u11_U19  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[4] ) );
INV_X4 _u0_u11_U17  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[3] ) );
INV_X4 _u0_u11_U15  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[2] ) );
INV_X4 _u0_u11_U13  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[1] ) );
INV_X4 _u0_u11_U11  ( .A(1'b1), .ZN(_u0_u11_sw_pointer[0] ) );
INV_X4 _u0_u11_U9  ( .A(1'b1), .ZN(_u0_u11_ch_stop ) );
INV_X4 _u0_u11_U7  ( .A(1'b1), .ZN(_u0_u11_ch_dis ) );
INV_X4 _u0_u11_U5  ( .A(1'b1), .ZN(_u0_u11_int ) );
INV_X4 _u0_u12_U585  ( .A(1'b1), .ZN(_u0_u12_pointer[31] ) );
INV_X4 _u0_u12_U583  ( .A(1'b1), .ZN(_u0_u12_pointer[30] ) );
INV_X4 _u0_u12_U581  ( .A(1'b1), .ZN(_u0_u12_pointer[29] ) );
INV_X4 _u0_u12_U579  ( .A(1'b1), .ZN(_u0_u12_pointer[28] ) );
INV_X4 _u0_u12_U577  ( .A(1'b1), .ZN(_u0_u12_pointer[27] ) );
INV_X4 _u0_u12_U575  ( .A(1'b1), .ZN(_u0_u12_pointer[26] ) );
INV_X4 _u0_u12_U573  ( .A(1'b1), .ZN(_u0_u12_pointer[25] ) );
INV_X4 _u0_u12_U571  ( .A(1'b1), .ZN(_u0_u12_pointer[24] ) );
INV_X4 _u0_u12_U569  ( .A(1'b1), .ZN(_u0_u12_pointer[23] ) );
INV_X4 _u0_u12_U567  ( .A(1'b1), .ZN(_u0_u12_pointer[22] ) );
INV_X4 _u0_u12_U565  ( .A(1'b1), .ZN(_u0_u12_pointer[21] ) );
INV_X4 _u0_u12_U563  ( .A(1'b1), .ZN(_u0_u12_pointer[20] ) );
INV_X4 _u0_u12_U561  ( .A(1'b1), .ZN(_u0_u12_pointer[19] ) );
INV_X4 _u0_u12_U559  ( .A(1'b1), .ZN(_u0_u12_pointer[18] ) );
INV_X4 _u0_u12_U557  ( .A(1'b1), .ZN(_u0_u12_pointer[17] ) );
INV_X4 _u0_u12_U555  ( .A(1'b1), .ZN(_u0_u12_pointer[16] ) );
INV_X4 _u0_u12_U553  ( .A(1'b1), .ZN(_u0_u12_pointer[15] ) );
INV_X4 _u0_u12_U551  ( .A(1'b1), .ZN(_u0_u12_pointer[14] ) );
INV_X4 _u0_u12_U549  ( .A(1'b1), .ZN(_u0_u12_pointer[13] ) );
INV_X4 _u0_u12_U547  ( .A(1'b1), .ZN(_u0_u12_pointer[12] ) );
INV_X4 _u0_u12_U545  ( .A(1'b1), .ZN(_u0_u12_pointer[11] ) );
INV_X4 _u0_u12_U543  ( .A(1'b1), .ZN(_u0_u12_pointer[10] ) );
INV_X4 _u0_u12_U541  ( .A(1'b1), .ZN(_u0_u12_pointer[9] ) );
INV_X4 _u0_u12_U539  ( .A(1'b1), .ZN(_u0_u12_pointer[8] ) );
INV_X4 _u0_u12_U537  ( .A(1'b1), .ZN(_u0_u12_pointer[7] ) );
INV_X4 _u0_u12_U535  ( .A(1'b1), .ZN(_u0_u12_pointer[6] ) );
INV_X4 _u0_u12_U533  ( .A(1'b1), .ZN(_u0_u12_pointer[5] ) );
INV_X4 _u0_u12_U531  ( .A(1'b1), .ZN(_u0_u12_pointer[4] ) );
INV_X4 _u0_u12_U529  ( .A(1'b1), .ZN(_u0_u12_pointer[3] ) );
INV_X4 _u0_u12_U527  ( .A(1'b1), .ZN(_u0_u12_pointer[2] ) );
INV_X4 _u0_u12_U525  ( .A(1'b1), .ZN(_u0_u12_pointer[1] ) );
INV_X4 _u0_u12_U523  ( .A(1'b1), .ZN(_u0_u12_pointer[0] ) );
INV_X4 _u0_u12_U521  ( .A(1'b1), .ZN(_u0_u12_pointer_s[31] ) );
INV_X4 _u0_u12_U519  ( .A(1'b1), .ZN(_u0_u12_pointer_s[30] ) );
INV_X4 _u0_u12_U517  ( .A(1'b1), .ZN(_u0_u12_pointer_s[29] ) );
INV_X4 _u0_u12_U515  ( .A(1'b1), .ZN(_u0_u12_pointer_s[28] ) );
INV_X4 _u0_u12_U513  ( .A(1'b1), .ZN(_u0_u12_pointer_s[27] ) );
INV_X4 _u0_u12_U511  ( .A(1'b1), .ZN(_u0_u12_pointer_s[26] ) );
INV_X4 _u0_u12_U509  ( .A(1'b1), .ZN(_u0_u12_pointer_s[25] ) );
INV_X4 _u0_u12_U507  ( .A(1'b1), .ZN(_u0_u12_pointer_s[24] ) );
INV_X4 _u0_u12_U505  ( .A(1'b1), .ZN(_u0_u12_pointer_s[23] ) );
INV_X4 _u0_u12_U503  ( .A(1'b1), .ZN(_u0_u12_pointer_s[22] ) );
INV_X4 _u0_u12_U501  ( .A(1'b1), .ZN(_u0_u12_pointer_s[21] ) );
INV_X4 _u0_u12_U499  ( .A(1'b1), .ZN(_u0_u12_pointer_s[20] ) );
INV_X4 _u0_u12_U497  ( .A(1'b1), .ZN(_u0_u12_pointer_s[19] ) );
INV_X4 _u0_u12_U495  ( .A(1'b1), .ZN(_u0_u12_pointer_s[18] ) );
INV_X4 _u0_u12_U493  ( .A(1'b1), .ZN(_u0_u12_pointer_s[17] ) );
INV_X4 _u0_u12_U491  ( .A(1'b1), .ZN(_u0_u12_pointer_s[16] ) );
INV_X4 _u0_u12_U489  ( .A(1'b1), .ZN(_u0_u12_pointer_s[15] ) );
INV_X4 _u0_u12_U487  ( .A(1'b1), .ZN(_u0_u12_pointer_s[14] ) );
INV_X4 _u0_u12_U485  ( .A(1'b1), .ZN(_u0_u12_pointer_s[13] ) );
INV_X4 _u0_u12_U483  ( .A(1'b1), .ZN(_u0_u12_pointer_s[12] ) );
INV_X4 _u0_u12_U481  ( .A(1'b1), .ZN(_u0_u12_pointer_s[11] ) );
INV_X4 _u0_u12_U479  ( .A(1'b1), .ZN(_u0_u12_pointer_s[10] ) );
INV_X4 _u0_u12_U477  ( .A(1'b1), .ZN(_u0_u12_pointer_s[9] ) );
INV_X4 _u0_u12_U475  ( .A(1'b1), .ZN(_u0_u12_pointer_s[8] ) );
INV_X4 _u0_u12_U473  ( .A(1'b1), .ZN(_u0_u12_pointer_s[7] ) );
INV_X4 _u0_u12_U471  ( .A(1'b1), .ZN(_u0_u12_pointer_s[6] ) );
INV_X4 _u0_u12_U469  ( .A(1'b1), .ZN(_u0_u12_pointer_s[5] ) );
INV_X4 _u0_u12_U467  ( .A(1'b1), .ZN(_u0_u12_pointer_s[4] ) );
INV_X4 _u0_u12_U465  ( .A(1'b1), .ZN(_u0_u12_pointer_s[3] ) );
INV_X4 _u0_u12_U463  ( .A(1'b1), .ZN(_u0_u12_pointer_s[2] ) );
INV_X4 _u0_u12_U461  ( .A(1'b1), .ZN(_u0_u12_pointer_s[1] ) );
INV_X4 _u0_u12_U459  ( .A(1'b1), .ZN(_u0_u12_pointer_s[0] ) );
INV_X4 _u0_u12_U457  ( .A(1'b1), .ZN(_u0_u12_ch_csr[31] ) );
INV_X4 _u0_u12_U455  ( .A(1'b1), .ZN(_u0_u12_ch_csr[30] ) );
INV_X4 _u0_u12_U453  ( .A(1'b1), .ZN(_u0_u12_ch_csr[29] ) );
INV_X4 _u0_u12_U451  ( .A(1'b1), .ZN(_u0_u12_ch_csr[28] ) );
INV_X4 _u0_u12_U449  ( .A(1'b1), .ZN(_u0_u12_ch_csr[27] ) );
INV_X4 _u0_u12_U447  ( .A(1'b1), .ZN(_u0_u12_ch_csr[26] ) );
INV_X4 _u0_u12_U445  ( .A(1'b1), .ZN(_u0_u12_ch_csr[25] ) );
INV_X4 _u0_u12_U443  ( .A(1'b1), .ZN(_u0_u12_ch_csr[24] ) );
INV_X4 _u0_u12_U441  ( .A(1'b1), .ZN(_u0_u12_ch_csr[23] ) );
INV_X4 _u0_u12_U439  ( .A(1'b1), .ZN(_u0_u12_ch_csr[22] ) );
INV_X4 _u0_u12_U437  ( .A(1'b1), .ZN(_u0_u12_ch_csr[21] ) );
INV_X4 _u0_u12_U435  ( .A(1'b1), .ZN(_u0_u12_ch_csr[20] ) );
INV_X4 _u0_u12_U433  ( .A(1'b1), .ZN(_u0_u12_ch_csr[19] ) );
INV_X4 _u0_u12_U431  ( .A(1'b1), .ZN(_u0_u12_ch_csr[18] ) );
INV_X4 _u0_u12_U429  ( .A(1'b1), .ZN(_u0_u12_ch_csr[17] ) );
INV_X4 _u0_u12_U427  ( .A(1'b1), .ZN(_u0_u12_ch_csr[16] ) );
INV_X4 _u0_u12_U425  ( .A(1'b1), .ZN(_u0_u12_ch_csr[15] ) );
INV_X4 _u0_u12_U423  ( .A(1'b1), .ZN(_u0_u12_ch_csr[14] ) );
INV_X4 _u0_u12_U421  ( .A(1'b1), .ZN(_u0_u12_ch_csr[13] ) );
INV_X4 _u0_u12_U419  ( .A(1'b1), .ZN(_u0_u12_ch_csr[12] ) );
INV_X4 _u0_u12_U417  ( .A(1'b1), .ZN(_u0_u12_ch_csr[11] ) );
INV_X4 _u0_u12_U415  ( .A(1'b1), .ZN(_u0_u12_ch_csr[10] ) );
INV_X4 _u0_u12_U413  ( .A(1'b1), .ZN(_u0_u12_ch_csr[9] ) );
INV_X4 _u0_u12_U411  ( .A(1'b1), .ZN(_u0_u12_ch_csr[8] ) );
INV_X4 _u0_u12_U409  ( .A(1'b1), .ZN(_u0_u12_ch_csr[7] ) );
INV_X4 _u0_u12_U407  ( .A(1'b1), .ZN(_u0_u12_ch_csr[6] ) );
INV_X4 _u0_u12_U405  ( .A(1'b1), .ZN(_u0_u12_ch_csr[5] ) );
INV_X4 _u0_u12_U403  ( .A(1'b1), .ZN(_u0_u12_ch_csr[4] ) );
INV_X4 _u0_u12_U401  ( .A(1'b1), .ZN(_u0_u12_ch_csr[3] ) );
INV_X4 _u0_u12_U399  ( .A(1'b1), .ZN(_u0_u12_ch_csr[2] ) );
INV_X4 _u0_u12_U397  ( .A(1'b1), .ZN(_u0_u12_ch_csr[1] ) );
INV_X4 _u0_u12_U395  ( .A(1'b1), .ZN(_u0_u12_ch_csr[0] ) );
INV_X4 _u0_u12_U393  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[31] ) );
INV_X4 _u0_u12_U391  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[30] ) );
INV_X4 _u0_u12_U389  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[29] ) );
INV_X4 _u0_u12_U387  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[28] ) );
INV_X4 _u0_u12_U385  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[27] ) );
INV_X4 _u0_u12_U383  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[26] ) );
INV_X4 _u0_u12_U381  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[25] ) );
INV_X4 _u0_u12_U379  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[24] ) );
INV_X4 _u0_u12_U377  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[23] ) );
INV_X4 _u0_u12_U375  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[22] ) );
INV_X4 _u0_u12_U373  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[21] ) );
INV_X4 _u0_u12_U371  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[20] ) );
INV_X4 _u0_u12_U369  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[19] ) );
INV_X4 _u0_u12_U367  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[18] ) );
INV_X4 _u0_u12_U365  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[17] ) );
INV_X4 _u0_u12_U363  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[16] ) );
INV_X4 _u0_u12_U361  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[15] ) );
INV_X4 _u0_u12_U359  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[14] ) );
INV_X4 _u0_u12_U357  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[13] ) );
INV_X4 _u0_u12_U355  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[12] ) );
INV_X4 _u0_u12_U353  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[11] ) );
INV_X4 _u0_u12_U351  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[10] ) );
INV_X4 _u0_u12_U349  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[9] ) );
INV_X4 _u0_u12_U347  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[8] ) );
INV_X4 _u0_u12_U345  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[7] ) );
INV_X4 _u0_u12_U343  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[6] ) );
INV_X4 _u0_u12_U341  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[5] ) );
INV_X4 _u0_u12_U339  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[4] ) );
INV_X4 _u0_u12_U337  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[3] ) );
INV_X4 _u0_u12_U335  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[2] ) );
INV_X4 _u0_u12_U333  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[1] ) );
INV_X4 _u0_u12_U331  ( .A(1'b1), .ZN(_u0_u12_ch_txsz[0] ) );
INV_X4 _u0_u12_U329  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[31] ) );
INV_X4 _u0_u12_U327  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[30] ) );
INV_X4 _u0_u12_U325  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[29] ) );
INV_X4 _u0_u12_U323  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[28] ) );
INV_X4 _u0_u12_U321  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[27] ) );
INV_X4 _u0_u12_U319  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[26] ) );
INV_X4 _u0_u12_U317  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[25] ) );
INV_X4 _u0_u12_U315  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[24] ) );
INV_X4 _u0_u12_U313  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[23] ) );
INV_X4 _u0_u12_U311  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[22] ) );
INV_X4 _u0_u12_U309  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[21] ) );
INV_X4 _u0_u12_U307  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[20] ) );
INV_X4 _u0_u12_U305  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[19] ) );
INV_X4 _u0_u12_U303  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[18] ) );
INV_X4 _u0_u12_U301  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[17] ) );
INV_X4 _u0_u12_U299  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[16] ) );
INV_X4 _u0_u12_U297  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[15] ) );
INV_X4 _u0_u12_U295  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[14] ) );
INV_X4 _u0_u12_U293  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[13] ) );
INV_X4 _u0_u12_U291  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[12] ) );
INV_X4 _u0_u12_U289  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[11] ) );
INV_X4 _u0_u12_U287  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[10] ) );
INV_X4 _u0_u12_U285  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[9] ) );
INV_X4 _u0_u12_U283  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[8] ) );
INV_X4 _u0_u12_U281  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[7] ) );
INV_X4 _u0_u12_U279  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[6] ) );
INV_X4 _u0_u12_U277  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[5] ) );
INV_X4 _u0_u12_U275  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[4] ) );
INV_X4 _u0_u12_U273  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[3] ) );
INV_X4 _u0_u12_U271  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[2] ) );
INV_X4 _u0_u12_U269  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[1] ) );
INV_X4 _u0_u12_U267  ( .A(1'b1), .ZN(_u0_u12_ch_adr0[0] ) );
INV_X4 _u0_u12_U265  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[31] ) );
INV_X4 _u0_u12_U263  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[30] ) );
INV_X4 _u0_u12_U261  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[29] ) );
INV_X4 _u0_u12_U259  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[28] ) );
INV_X4 _u0_u12_U257  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[27] ) );
INV_X4 _u0_u12_U255  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[26] ) );
INV_X4 _u0_u12_U253  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[25] ) );
INV_X4 _u0_u12_U251  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[24] ) );
INV_X4 _u0_u12_U249  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[23] ) );
INV_X4 _u0_u12_U247  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[22] ) );
INV_X4 _u0_u12_U245  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[21] ) );
INV_X4 _u0_u12_U243  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[20] ) );
INV_X4 _u0_u12_U241  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[19] ) );
INV_X4 _u0_u12_U239  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[18] ) );
INV_X4 _u0_u12_U237  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[17] ) );
INV_X4 _u0_u12_U235  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[16] ) );
INV_X4 _u0_u12_U233  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[15] ) );
INV_X4 _u0_u12_U231  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[14] ) );
INV_X4 _u0_u12_U229  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[13] ) );
INV_X4 _u0_u12_U227  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[12] ) );
INV_X4 _u0_u12_U225  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[11] ) );
INV_X4 _u0_u12_U223  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[10] ) );
INV_X4 _u0_u12_U221  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[9] ) );
INV_X4 _u0_u12_U219  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[8] ) );
INV_X4 _u0_u12_U217  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[7] ) );
INV_X4 _u0_u12_U215  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[6] ) );
INV_X4 _u0_u12_U213  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[5] ) );
INV_X4 _u0_u12_U211  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[4] ) );
INV_X4 _u0_u12_U209  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[3] ) );
INV_X4 _u0_u12_U207  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[2] ) );
INV_X4 _u0_u12_U205  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[1] ) );
INV_X4 _u0_u12_U203  ( .A(1'b1), .ZN(_u0_u12_ch_adr1[0] ) );
INV_X4 _u0_u12_U201  ( .A(1'b0), .ZN(_u0_u12_ch_am0[31] ) );
INV_X4 _u0_u12_U199  ( .A(1'b0), .ZN(_u0_u12_ch_am0[30] ) );
INV_X4 _u0_u12_U197  ( .A(1'b0), .ZN(_u0_u12_ch_am0[29] ) );
INV_X4 _u0_u12_U195  ( .A(1'b0), .ZN(_u0_u12_ch_am0[28] ) );
INV_X4 _u0_u12_U193  ( .A(1'b0), .ZN(_u0_u12_ch_am0[27] ) );
INV_X4 _u0_u12_U191  ( .A(1'b0), .ZN(_u0_u12_ch_am0[26] ) );
INV_X4 _u0_u12_U189  ( .A(1'b0), .ZN(_u0_u12_ch_am0[25] ) );
INV_X4 _u0_u12_U187  ( .A(1'b0), .ZN(_u0_u12_ch_am0[24] ) );
INV_X4 _u0_u12_U185  ( .A(1'b0), .ZN(_u0_u12_ch_am0[23] ) );
INV_X4 _u0_u12_U183  ( .A(1'b0), .ZN(_u0_u12_ch_am0[22] ) );
INV_X4 _u0_u12_U181  ( .A(1'b0), .ZN(_u0_u12_ch_am0[21] ) );
INV_X4 _u0_u12_U179  ( .A(1'b0), .ZN(_u0_u12_ch_am0[20] ) );
INV_X4 _u0_u12_U177  ( .A(1'b0), .ZN(_u0_u12_ch_am0[19] ) );
INV_X4 _u0_u12_U175  ( .A(1'b0), .ZN(_u0_u12_ch_am0[18] ) );
INV_X4 _u0_u12_U173  ( .A(1'b0), .ZN(_u0_u12_ch_am0[17] ) );
INV_X4 _u0_u12_U171  ( .A(1'b0), .ZN(_u0_u12_ch_am0[16] ) );
INV_X4 _u0_u12_U169  ( .A(1'b0), .ZN(_u0_u12_ch_am0[15] ) );
INV_X4 _u0_u12_U167  ( .A(1'b0), .ZN(_u0_u12_ch_am0[14] ) );
INV_X4 _u0_u12_U165  ( .A(1'b0), .ZN(_u0_u12_ch_am0[13] ) );
INV_X4 _u0_u12_U163  ( .A(1'b0), .ZN(_u0_u12_ch_am0[12] ) );
INV_X4 _u0_u12_U161  ( .A(1'b0), .ZN(_u0_u12_ch_am0[11] ) );
INV_X4 _u0_u12_U159  ( .A(1'b0), .ZN(_u0_u12_ch_am0[10] ) );
INV_X4 _u0_u12_U157  ( .A(1'b0), .ZN(_u0_u12_ch_am0[9] ) );
INV_X4 _u0_u12_U155  ( .A(1'b0), .ZN(_u0_u12_ch_am0[8] ) );
INV_X4 _u0_u12_U153  ( .A(1'b0), .ZN(_u0_u12_ch_am0[7] ) );
INV_X4 _u0_u12_U151  ( .A(1'b0), .ZN(_u0_u12_ch_am0[6] ) );
INV_X4 _u0_u12_U149  ( .A(1'b0), .ZN(_u0_u12_ch_am0[5] ) );
INV_X4 _u0_u12_U147  ( .A(1'b0), .ZN(_u0_u12_ch_am0[4] ) );
INV_X4 _u0_u12_U145  ( .A(1'b1), .ZN(_u0_u12_ch_am0[3] ) );
INV_X4 _u0_u12_U143  ( .A(1'b1), .ZN(_u0_u12_ch_am0[2] ) );
INV_X4 _u0_u12_U141  ( .A(1'b1), .ZN(_u0_u12_ch_am0[1] ) );
INV_X4 _u0_u12_U139  ( .A(1'b1), .ZN(_u0_u12_ch_am0[0] ) );
INV_X4 _u0_u12_U137  ( .A(1'b0), .ZN(_u0_u12_ch_am1[31] ) );
INV_X4 _u0_u12_U135  ( .A(1'b0), .ZN(_u0_u12_ch_am1[30] ) );
INV_X4 _u0_u12_U133  ( .A(1'b0), .ZN(_u0_u12_ch_am1[29] ) );
INV_X4 _u0_u12_U131  ( .A(1'b0), .ZN(_u0_u12_ch_am1[28] ) );
INV_X4 _u0_u12_U129  ( .A(1'b0), .ZN(_u0_u12_ch_am1[27] ) );
INV_X4 _u0_u12_U127  ( .A(1'b0), .ZN(_u0_u12_ch_am1[26] ) );
INV_X4 _u0_u12_U125  ( .A(1'b0), .ZN(_u0_u12_ch_am1[25] ) );
INV_X4 _u0_u12_U123  ( .A(1'b0), .ZN(_u0_u12_ch_am1[24] ) );
INV_X4 _u0_u12_U121  ( .A(1'b0), .ZN(_u0_u12_ch_am1[23] ) );
INV_X4 _u0_u12_U119  ( .A(1'b0), .ZN(_u0_u12_ch_am1[22] ) );
INV_X4 _u0_u12_U117  ( .A(1'b0), .ZN(_u0_u12_ch_am1[21] ) );
INV_X4 _u0_u12_U115  ( .A(1'b0), .ZN(_u0_u12_ch_am1[20] ) );
INV_X4 _u0_u12_U113  ( .A(1'b0), .ZN(_u0_u12_ch_am1[19] ) );
INV_X4 _u0_u12_U111  ( .A(1'b0), .ZN(_u0_u12_ch_am1[18] ) );
INV_X4 _u0_u12_U109  ( .A(1'b0), .ZN(_u0_u12_ch_am1[17] ) );
INV_X4 _u0_u12_U107  ( .A(1'b0), .ZN(_u0_u12_ch_am1[16] ) );
INV_X4 _u0_u12_U105  ( .A(1'b0), .ZN(_u0_u12_ch_am1[15] ) );
INV_X4 _u0_u12_U103  ( .A(1'b0), .ZN(_u0_u12_ch_am1[14] ) );
INV_X4 _u0_u12_U101  ( .A(1'b0), .ZN(_u0_u12_ch_am1[13] ) );
INV_X4 _u0_u12_U99  ( .A(1'b0), .ZN(_u0_u12_ch_am1[12] ) );
INV_X4 _u0_u12_U97  ( .A(1'b0), .ZN(_u0_u12_ch_am1[11] ) );
INV_X4 _u0_u12_U95  ( .A(1'b0), .ZN(_u0_u12_ch_am1[10] ) );
INV_X4 _u0_u12_U93  ( .A(1'b0), .ZN(_u0_u12_ch_am1[9] ) );
INV_X4 _u0_u12_U91  ( .A(1'b0), .ZN(_u0_u12_ch_am1[8] ) );
INV_X4 _u0_u12_U89  ( .A(1'b0), .ZN(_u0_u12_ch_am1[7] ) );
INV_X4 _u0_u12_U87  ( .A(1'b0), .ZN(_u0_u12_ch_am1[6] ) );
INV_X4 _u0_u12_U85  ( .A(1'b0), .ZN(_u0_u12_ch_am1[5] ) );
INV_X4 _u0_u12_U83  ( .A(1'b0), .ZN(_u0_u12_ch_am1[4] ) );
INV_X4 _u0_u12_U81  ( .A(1'b1), .ZN(_u0_u12_ch_am1[3] ) );
INV_X4 _u0_u12_U79  ( .A(1'b1), .ZN(_u0_u12_ch_am1[2] ) );
INV_X4 _u0_u12_U77  ( .A(1'b1), .ZN(_u0_u12_ch_am1[1] ) );
INV_X4 _u0_u12_U75  ( .A(1'b1), .ZN(_u0_u12_ch_am1[0] ) );
INV_X4 _u0_u12_U73  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[31] ) );
INV_X4 _u0_u12_U71  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[30] ) );
INV_X4 _u0_u12_U69  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[29] ) );
INV_X4 _u0_u12_U67  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[28] ) );
INV_X4 _u0_u12_U65  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[27] ) );
INV_X4 _u0_u12_U63  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[26] ) );
INV_X4 _u0_u12_U61  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[25] ) );
INV_X4 _u0_u12_U59  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[24] ) );
INV_X4 _u0_u12_U57  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[23] ) );
INV_X4 _u0_u12_U55  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[22] ) );
INV_X4 _u0_u12_U53  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[21] ) );
INV_X4 _u0_u12_U51  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[20] ) );
INV_X4 _u0_u12_U49  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[19] ) );
INV_X4 _u0_u12_U47  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[18] ) );
INV_X4 _u0_u12_U45  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[17] ) );
INV_X4 _u0_u12_U43  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[16] ) );
INV_X4 _u0_u12_U41  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[15] ) );
INV_X4 _u0_u12_U39  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[14] ) );
INV_X4 _u0_u12_U37  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[13] ) );
INV_X4 _u0_u12_U35  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[12] ) );
INV_X4 _u0_u12_U33  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[11] ) );
INV_X4 _u0_u12_U31  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[10] ) );
INV_X4 _u0_u12_U29  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[9] ) );
INV_X4 _u0_u12_U27  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[8] ) );
INV_X4 _u0_u12_U25  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[7] ) );
INV_X4 _u0_u12_U23  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[6] ) );
INV_X4 _u0_u12_U21  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[5] ) );
INV_X4 _u0_u12_U19  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[4] ) );
INV_X4 _u0_u12_U17  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[3] ) );
INV_X4 _u0_u12_U15  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[2] ) );
INV_X4 _u0_u12_U13  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[1] ) );
INV_X4 _u0_u12_U11  ( .A(1'b1), .ZN(_u0_u12_sw_pointer[0] ) );
INV_X4 _u0_u12_U9  ( .A(1'b1), .ZN(_u0_u12_ch_stop ) );
INV_X4 _u0_u12_U7  ( .A(1'b1), .ZN(_u0_u12_ch_dis ) );
INV_X4 _u0_u12_U5  ( .A(1'b1), .ZN(_u0_u12_int ) );
INV_X4 _u0_u13_U585  ( .A(1'b1), .ZN(_u0_u13_pointer[31] ) );
INV_X4 _u0_u13_U583  ( .A(1'b1), .ZN(_u0_u13_pointer[30] ) );
INV_X4 _u0_u13_U581  ( .A(1'b1), .ZN(_u0_u13_pointer[29] ) );
INV_X4 _u0_u13_U579  ( .A(1'b1), .ZN(_u0_u13_pointer[28] ) );
INV_X4 _u0_u13_U577  ( .A(1'b1), .ZN(_u0_u13_pointer[27] ) );
INV_X4 _u0_u13_U575  ( .A(1'b1), .ZN(_u0_u13_pointer[26] ) );
INV_X4 _u0_u13_U573  ( .A(1'b1), .ZN(_u0_u13_pointer[25] ) );
INV_X4 _u0_u13_U571  ( .A(1'b1), .ZN(_u0_u13_pointer[24] ) );
INV_X4 _u0_u13_U569  ( .A(1'b1), .ZN(_u0_u13_pointer[23] ) );
INV_X4 _u0_u13_U567  ( .A(1'b1), .ZN(_u0_u13_pointer[22] ) );
INV_X4 _u0_u13_U565  ( .A(1'b1), .ZN(_u0_u13_pointer[21] ) );
INV_X4 _u0_u13_U563  ( .A(1'b1), .ZN(_u0_u13_pointer[20] ) );
INV_X4 _u0_u13_U561  ( .A(1'b1), .ZN(_u0_u13_pointer[19] ) );
INV_X4 _u0_u13_U559  ( .A(1'b1), .ZN(_u0_u13_pointer[18] ) );
INV_X4 _u0_u13_U557  ( .A(1'b1), .ZN(_u0_u13_pointer[17] ) );
INV_X4 _u0_u13_U555  ( .A(1'b1), .ZN(_u0_u13_pointer[16] ) );
INV_X4 _u0_u13_U553  ( .A(1'b1), .ZN(_u0_u13_pointer[15] ) );
INV_X4 _u0_u13_U551  ( .A(1'b1), .ZN(_u0_u13_pointer[14] ) );
INV_X4 _u0_u13_U549  ( .A(1'b1), .ZN(_u0_u13_pointer[13] ) );
INV_X4 _u0_u13_U547  ( .A(1'b1), .ZN(_u0_u13_pointer[12] ) );
INV_X4 _u0_u13_U545  ( .A(1'b1), .ZN(_u0_u13_pointer[11] ) );
INV_X4 _u0_u13_U543  ( .A(1'b1), .ZN(_u0_u13_pointer[10] ) );
INV_X4 _u0_u13_U541  ( .A(1'b1), .ZN(_u0_u13_pointer[9] ) );
INV_X4 _u0_u13_U539  ( .A(1'b1), .ZN(_u0_u13_pointer[8] ) );
INV_X4 _u0_u13_U537  ( .A(1'b1), .ZN(_u0_u13_pointer[7] ) );
INV_X4 _u0_u13_U535  ( .A(1'b1), .ZN(_u0_u13_pointer[6] ) );
INV_X4 _u0_u13_U533  ( .A(1'b1), .ZN(_u0_u13_pointer[5] ) );
INV_X4 _u0_u13_U531  ( .A(1'b1), .ZN(_u0_u13_pointer[4] ) );
INV_X4 _u0_u13_U529  ( .A(1'b1), .ZN(_u0_u13_pointer[3] ) );
INV_X4 _u0_u13_U527  ( .A(1'b1), .ZN(_u0_u13_pointer[2] ) );
INV_X4 _u0_u13_U525  ( .A(1'b1), .ZN(_u0_u13_pointer[1] ) );
INV_X4 _u0_u13_U523  ( .A(1'b1), .ZN(_u0_u13_pointer[0] ) );
INV_X4 _u0_u13_U521  ( .A(1'b1), .ZN(_u0_u13_pointer_s[31] ) );
INV_X4 _u0_u13_U519  ( .A(1'b1), .ZN(_u0_u13_pointer_s[30] ) );
INV_X4 _u0_u13_U517  ( .A(1'b1), .ZN(_u0_u13_pointer_s[29] ) );
INV_X4 _u0_u13_U515  ( .A(1'b1), .ZN(_u0_u13_pointer_s[28] ) );
INV_X4 _u0_u13_U513  ( .A(1'b1), .ZN(_u0_u13_pointer_s[27] ) );
INV_X4 _u0_u13_U511  ( .A(1'b1), .ZN(_u0_u13_pointer_s[26] ) );
INV_X4 _u0_u13_U509  ( .A(1'b1), .ZN(_u0_u13_pointer_s[25] ) );
INV_X4 _u0_u13_U507  ( .A(1'b1), .ZN(_u0_u13_pointer_s[24] ) );
INV_X4 _u0_u13_U505  ( .A(1'b1), .ZN(_u0_u13_pointer_s[23] ) );
INV_X4 _u0_u13_U503  ( .A(1'b1), .ZN(_u0_u13_pointer_s[22] ) );
INV_X4 _u0_u13_U501  ( .A(1'b1), .ZN(_u0_u13_pointer_s[21] ) );
INV_X4 _u0_u13_U499  ( .A(1'b1), .ZN(_u0_u13_pointer_s[20] ) );
INV_X4 _u0_u13_U497  ( .A(1'b1), .ZN(_u0_u13_pointer_s[19] ) );
INV_X4 _u0_u13_U495  ( .A(1'b1), .ZN(_u0_u13_pointer_s[18] ) );
INV_X4 _u0_u13_U493  ( .A(1'b1), .ZN(_u0_u13_pointer_s[17] ) );
INV_X4 _u0_u13_U491  ( .A(1'b1), .ZN(_u0_u13_pointer_s[16] ) );
INV_X4 _u0_u13_U489  ( .A(1'b1), .ZN(_u0_u13_pointer_s[15] ) );
INV_X4 _u0_u13_U487  ( .A(1'b1), .ZN(_u0_u13_pointer_s[14] ) );
INV_X4 _u0_u13_U485  ( .A(1'b1), .ZN(_u0_u13_pointer_s[13] ) );
INV_X4 _u0_u13_U483  ( .A(1'b1), .ZN(_u0_u13_pointer_s[12] ) );
INV_X4 _u0_u13_U481  ( .A(1'b1), .ZN(_u0_u13_pointer_s[11] ) );
INV_X4 _u0_u13_U479  ( .A(1'b1), .ZN(_u0_u13_pointer_s[10] ) );
INV_X4 _u0_u13_U477  ( .A(1'b1), .ZN(_u0_u13_pointer_s[9] ) );
INV_X4 _u0_u13_U475  ( .A(1'b1), .ZN(_u0_u13_pointer_s[8] ) );
INV_X4 _u0_u13_U473  ( .A(1'b1), .ZN(_u0_u13_pointer_s[7] ) );
INV_X4 _u0_u13_U471  ( .A(1'b1), .ZN(_u0_u13_pointer_s[6] ) );
INV_X4 _u0_u13_U469  ( .A(1'b1), .ZN(_u0_u13_pointer_s[5] ) );
INV_X4 _u0_u13_U467  ( .A(1'b1), .ZN(_u0_u13_pointer_s[4] ) );
INV_X4 _u0_u13_U465  ( .A(1'b1), .ZN(_u0_u13_pointer_s[3] ) );
INV_X4 _u0_u13_U463  ( .A(1'b1), .ZN(_u0_u13_pointer_s[2] ) );
INV_X4 _u0_u13_U461  ( .A(1'b1), .ZN(_u0_u13_pointer_s[1] ) );
INV_X4 _u0_u13_U459  ( .A(1'b1), .ZN(_u0_u13_pointer_s[0] ) );
INV_X4 _u0_u13_U457  ( .A(1'b1), .ZN(_u0_u13_ch_csr[31] ) );
INV_X4 _u0_u13_U455  ( .A(1'b1), .ZN(_u0_u13_ch_csr[30] ) );
INV_X4 _u0_u13_U453  ( .A(1'b1), .ZN(_u0_u13_ch_csr[29] ) );
INV_X4 _u0_u13_U451  ( .A(1'b1), .ZN(_u0_u13_ch_csr[28] ) );
INV_X4 _u0_u13_U449  ( .A(1'b1), .ZN(_u0_u13_ch_csr[27] ) );
INV_X4 _u0_u13_U447  ( .A(1'b1), .ZN(_u0_u13_ch_csr[26] ) );
INV_X4 _u0_u13_U445  ( .A(1'b1), .ZN(_u0_u13_ch_csr[25] ) );
INV_X4 _u0_u13_U443  ( .A(1'b1), .ZN(_u0_u13_ch_csr[24] ) );
INV_X4 _u0_u13_U441  ( .A(1'b1), .ZN(_u0_u13_ch_csr[23] ) );
INV_X4 _u0_u13_U439  ( .A(1'b1), .ZN(_u0_u13_ch_csr[22] ) );
INV_X4 _u0_u13_U437  ( .A(1'b1), .ZN(_u0_u13_ch_csr[21] ) );
INV_X4 _u0_u13_U435  ( .A(1'b1), .ZN(_u0_u13_ch_csr[20] ) );
INV_X4 _u0_u13_U433  ( .A(1'b1), .ZN(_u0_u13_ch_csr[19] ) );
INV_X4 _u0_u13_U431  ( .A(1'b1), .ZN(_u0_u13_ch_csr[18] ) );
INV_X4 _u0_u13_U429  ( .A(1'b1), .ZN(_u0_u13_ch_csr[17] ) );
INV_X4 _u0_u13_U427  ( .A(1'b1), .ZN(_u0_u13_ch_csr[16] ) );
INV_X4 _u0_u13_U425  ( .A(1'b1), .ZN(_u0_u13_ch_csr[15] ) );
INV_X4 _u0_u13_U423  ( .A(1'b1), .ZN(_u0_u13_ch_csr[14] ) );
INV_X4 _u0_u13_U421  ( .A(1'b1), .ZN(_u0_u13_ch_csr[13] ) );
INV_X4 _u0_u13_U419  ( .A(1'b1), .ZN(_u0_u13_ch_csr[12] ) );
INV_X4 _u0_u13_U417  ( .A(1'b1), .ZN(_u0_u13_ch_csr[11] ) );
INV_X4 _u0_u13_U415  ( .A(1'b1), .ZN(_u0_u13_ch_csr[10] ) );
INV_X4 _u0_u13_U413  ( .A(1'b1), .ZN(_u0_u13_ch_csr[9] ) );
INV_X4 _u0_u13_U411  ( .A(1'b1), .ZN(_u0_u13_ch_csr[8] ) );
INV_X4 _u0_u13_U409  ( .A(1'b1), .ZN(_u0_u13_ch_csr[7] ) );
INV_X4 _u0_u13_U407  ( .A(1'b1), .ZN(_u0_u13_ch_csr[6] ) );
INV_X4 _u0_u13_U405  ( .A(1'b1), .ZN(_u0_u13_ch_csr[5] ) );
INV_X4 _u0_u13_U403  ( .A(1'b1), .ZN(_u0_u13_ch_csr[4] ) );
INV_X4 _u0_u13_U401  ( .A(1'b1), .ZN(_u0_u13_ch_csr[3] ) );
INV_X4 _u0_u13_U399  ( .A(1'b1), .ZN(_u0_u13_ch_csr[2] ) );
INV_X4 _u0_u13_U397  ( .A(1'b1), .ZN(_u0_u13_ch_csr[1] ) );
INV_X4 _u0_u13_U395  ( .A(1'b1), .ZN(_u0_u13_ch_csr[0] ) );
INV_X4 _u0_u13_U393  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[31] ) );
INV_X4 _u0_u13_U391  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[30] ) );
INV_X4 _u0_u13_U389  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[29] ) );
INV_X4 _u0_u13_U387  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[28] ) );
INV_X4 _u0_u13_U385  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[27] ) );
INV_X4 _u0_u13_U383  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[26] ) );
INV_X4 _u0_u13_U381  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[25] ) );
INV_X4 _u0_u13_U379  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[24] ) );
INV_X4 _u0_u13_U377  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[23] ) );
INV_X4 _u0_u13_U375  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[22] ) );
INV_X4 _u0_u13_U373  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[21] ) );
INV_X4 _u0_u13_U371  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[20] ) );
INV_X4 _u0_u13_U369  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[19] ) );
INV_X4 _u0_u13_U367  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[18] ) );
INV_X4 _u0_u13_U365  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[17] ) );
INV_X4 _u0_u13_U363  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[16] ) );
INV_X4 _u0_u13_U361  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[15] ) );
INV_X4 _u0_u13_U359  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[14] ) );
INV_X4 _u0_u13_U357  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[13] ) );
INV_X4 _u0_u13_U355  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[12] ) );
INV_X4 _u0_u13_U353  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[11] ) );
INV_X4 _u0_u13_U351  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[10] ) );
INV_X4 _u0_u13_U349  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[9] ) );
INV_X4 _u0_u13_U347  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[8] ) );
INV_X4 _u0_u13_U345  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[7] ) );
INV_X4 _u0_u13_U343  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[6] ) );
INV_X4 _u0_u13_U341  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[5] ) );
INV_X4 _u0_u13_U339  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[4] ) );
INV_X4 _u0_u13_U337  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[3] ) );
INV_X4 _u0_u13_U335  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[2] ) );
INV_X4 _u0_u13_U333  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[1] ) );
INV_X4 _u0_u13_U331  ( .A(1'b1), .ZN(_u0_u13_ch_txsz[0] ) );
INV_X4 _u0_u13_U329  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[31] ) );
INV_X4 _u0_u13_U327  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[30] ) );
INV_X4 _u0_u13_U325  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[29] ) );
INV_X4 _u0_u13_U323  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[28] ) );
INV_X4 _u0_u13_U321  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[27] ) );
INV_X4 _u0_u13_U319  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[26] ) );
INV_X4 _u0_u13_U317  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[25] ) );
INV_X4 _u0_u13_U315  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[24] ) );
INV_X4 _u0_u13_U313  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[23] ) );
INV_X4 _u0_u13_U311  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[22] ) );
INV_X4 _u0_u13_U309  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[21] ) );
INV_X4 _u0_u13_U307  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[20] ) );
INV_X4 _u0_u13_U305  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[19] ) );
INV_X4 _u0_u13_U303  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[18] ) );
INV_X4 _u0_u13_U301  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[17] ) );
INV_X4 _u0_u13_U299  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[16] ) );
INV_X4 _u0_u13_U297  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[15] ) );
INV_X4 _u0_u13_U295  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[14] ) );
INV_X4 _u0_u13_U293  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[13] ) );
INV_X4 _u0_u13_U291  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[12] ) );
INV_X4 _u0_u13_U289  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[11] ) );
INV_X4 _u0_u13_U287  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[10] ) );
INV_X4 _u0_u13_U285  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[9] ) );
INV_X4 _u0_u13_U283  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[8] ) );
INV_X4 _u0_u13_U281  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[7] ) );
INV_X4 _u0_u13_U279  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[6] ) );
INV_X4 _u0_u13_U277  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[5] ) );
INV_X4 _u0_u13_U275  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[4] ) );
INV_X4 _u0_u13_U273  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[3] ) );
INV_X4 _u0_u13_U271  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[2] ) );
INV_X4 _u0_u13_U269  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[1] ) );
INV_X4 _u0_u13_U267  ( .A(1'b1), .ZN(_u0_u13_ch_adr0[0] ) );
INV_X4 _u0_u13_U265  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[31] ) );
INV_X4 _u0_u13_U263  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[30] ) );
INV_X4 _u0_u13_U261  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[29] ) );
INV_X4 _u0_u13_U259  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[28] ) );
INV_X4 _u0_u13_U257  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[27] ) );
INV_X4 _u0_u13_U255  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[26] ) );
INV_X4 _u0_u13_U253  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[25] ) );
INV_X4 _u0_u13_U251  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[24] ) );
INV_X4 _u0_u13_U249  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[23] ) );
INV_X4 _u0_u13_U247  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[22] ) );
INV_X4 _u0_u13_U245  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[21] ) );
INV_X4 _u0_u13_U243  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[20] ) );
INV_X4 _u0_u13_U241  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[19] ) );
INV_X4 _u0_u13_U239  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[18] ) );
INV_X4 _u0_u13_U237  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[17] ) );
INV_X4 _u0_u13_U235  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[16] ) );
INV_X4 _u0_u13_U233  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[15] ) );
INV_X4 _u0_u13_U231  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[14] ) );
INV_X4 _u0_u13_U229  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[13] ) );
INV_X4 _u0_u13_U227  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[12] ) );
INV_X4 _u0_u13_U225  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[11] ) );
INV_X4 _u0_u13_U223  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[10] ) );
INV_X4 _u0_u13_U221  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[9] ) );
INV_X4 _u0_u13_U219  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[8] ) );
INV_X4 _u0_u13_U217  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[7] ) );
INV_X4 _u0_u13_U215  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[6] ) );
INV_X4 _u0_u13_U213  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[5] ) );
INV_X4 _u0_u13_U211  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[4] ) );
INV_X4 _u0_u13_U209  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[3] ) );
INV_X4 _u0_u13_U207  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[2] ) );
INV_X4 _u0_u13_U205  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[1] ) );
INV_X4 _u0_u13_U203  ( .A(1'b1), .ZN(_u0_u13_ch_adr1[0] ) );
INV_X4 _u0_u13_U201  ( .A(1'b0), .ZN(_u0_u13_ch_am0[31] ) );
INV_X4 _u0_u13_U199  ( .A(1'b0), .ZN(_u0_u13_ch_am0[30] ) );
INV_X4 _u0_u13_U197  ( .A(1'b0), .ZN(_u0_u13_ch_am0[29] ) );
INV_X4 _u0_u13_U195  ( .A(1'b0), .ZN(_u0_u13_ch_am0[28] ) );
INV_X4 _u0_u13_U193  ( .A(1'b0), .ZN(_u0_u13_ch_am0[27] ) );
INV_X4 _u0_u13_U191  ( .A(1'b0), .ZN(_u0_u13_ch_am0[26] ) );
INV_X4 _u0_u13_U189  ( .A(1'b0), .ZN(_u0_u13_ch_am0[25] ) );
INV_X4 _u0_u13_U187  ( .A(1'b0), .ZN(_u0_u13_ch_am0[24] ) );
INV_X4 _u0_u13_U185  ( .A(1'b0), .ZN(_u0_u13_ch_am0[23] ) );
INV_X4 _u0_u13_U183  ( .A(1'b0), .ZN(_u0_u13_ch_am0[22] ) );
INV_X4 _u0_u13_U181  ( .A(1'b0), .ZN(_u0_u13_ch_am0[21] ) );
INV_X4 _u0_u13_U179  ( .A(1'b0), .ZN(_u0_u13_ch_am0[20] ) );
INV_X4 _u0_u13_U177  ( .A(1'b0), .ZN(_u0_u13_ch_am0[19] ) );
INV_X4 _u0_u13_U175  ( .A(1'b0), .ZN(_u0_u13_ch_am0[18] ) );
INV_X4 _u0_u13_U173  ( .A(1'b0), .ZN(_u0_u13_ch_am0[17] ) );
INV_X4 _u0_u13_U171  ( .A(1'b0), .ZN(_u0_u13_ch_am0[16] ) );
INV_X4 _u0_u13_U169  ( .A(1'b0), .ZN(_u0_u13_ch_am0[15] ) );
INV_X4 _u0_u13_U167  ( .A(1'b0), .ZN(_u0_u13_ch_am0[14] ) );
INV_X4 _u0_u13_U165  ( .A(1'b0), .ZN(_u0_u13_ch_am0[13] ) );
INV_X4 _u0_u13_U163  ( .A(1'b0), .ZN(_u0_u13_ch_am0[12] ) );
INV_X4 _u0_u13_U161  ( .A(1'b0), .ZN(_u0_u13_ch_am0[11] ) );
INV_X4 _u0_u13_U159  ( .A(1'b0), .ZN(_u0_u13_ch_am0[10] ) );
INV_X4 _u0_u13_U157  ( .A(1'b0), .ZN(_u0_u13_ch_am0[9] ) );
INV_X4 _u0_u13_U155  ( .A(1'b0), .ZN(_u0_u13_ch_am0[8] ) );
INV_X4 _u0_u13_U153  ( .A(1'b0), .ZN(_u0_u13_ch_am0[7] ) );
INV_X4 _u0_u13_U151  ( .A(1'b0), .ZN(_u0_u13_ch_am0[6] ) );
INV_X4 _u0_u13_U149  ( .A(1'b0), .ZN(_u0_u13_ch_am0[5] ) );
INV_X4 _u0_u13_U147  ( .A(1'b0), .ZN(_u0_u13_ch_am0[4] ) );
INV_X4 _u0_u13_U145  ( .A(1'b1), .ZN(_u0_u13_ch_am0[3] ) );
INV_X4 _u0_u13_U143  ( .A(1'b1), .ZN(_u0_u13_ch_am0[2] ) );
INV_X4 _u0_u13_U141  ( .A(1'b1), .ZN(_u0_u13_ch_am0[1] ) );
INV_X4 _u0_u13_U139  ( .A(1'b1), .ZN(_u0_u13_ch_am0[0] ) );
INV_X4 _u0_u13_U137  ( .A(1'b0), .ZN(_u0_u13_ch_am1[31] ) );
INV_X4 _u0_u13_U135  ( .A(1'b0), .ZN(_u0_u13_ch_am1[30] ) );
INV_X4 _u0_u13_U133  ( .A(1'b0), .ZN(_u0_u13_ch_am1[29] ) );
INV_X4 _u0_u13_U131  ( .A(1'b0), .ZN(_u0_u13_ch_am1[28] ) );
INV_X4 _u0_u13_U129  ( .A(1'b0), .ZN(_u0_u13_ch_am1[27] ) );
INV_X4 _u0_u13_U127  ( .A(1'b0), .ZN(_u0_u13_ch_am1[26] ) );
INV_X4 _u0_u13_U125  ( .A(1'b0), .ZN(_u0_u13_ch_am1[25] ) );
INV_X4 _u0_u13_U123  ( .A(1'b0), .ZN(_u0_u13_ch_am1[24] ) );
INV_X4 _u0_u13_U121  ( .A(1'b0), .ZN(_u0_u13_ch_am1[23] ) );
INV_X4 _u0_u13_U119  ( .A(1'b0), .ZN(_u0_u13_ch_am1[22] ) );
INV_X4 _u0_u13_U117  ( .A(1'b0), .ZN(_u0_u13_ch_am1[21] ) );
INV_X4 _u0_u13_U115  ( .A(1'b0), .ZN(_u0_u13_ch_am1[20] ) );
INV_X4 _u0_u13_U113  ( .A(1'b0), .ZN(_u0_u13_ch_am1[19] ) );
INV_X4 _u0_u13_U111  ( .A(1'b0), .ZN(_u0_u13_ch_am1[18] ) );
INV_X4 _u0_u13_U109  ( .A(1'b0), .ZN(_u0_u13_ch_am1[17] ) );
INV_X4 _u0_u13_U107  ( .A(1'b0), .ZN(_u0_u13_ch_am1[16] ) );
INV_X4 _u0_u13_U105  ( .A(1'b0), .ZN(_u0_u13_ch_am1[15] ) );
INV_X4 _u0_u13_U103  ( .A(1'b0), .ZN(_u0_u13_ch_am1[14] ) );
INV_X4 _u0_u13_U101  ( .A(1'b0), .ZN(_u0_u13_ch_am1[13] ) );
INV_X4 _u0_u13_U99  ( .A(1'b0), .ZN(_u0_u13_ch_am1[12] ) );
INV_X4 _u0_u13_U97  ( .A(1'b0), .ZN(_u0_u13_ch_am1[11] ) );
INV_X4 _u0_u13_U95  ( .A(1'b0), .ZN(_u0_u13_ch_am1[10] ) );
INV_X4 _u0_u13_U93  ( .A(1'b0), .ZN(_u0_u13_ch_am1[9] ) );
INV_X4 _u0_u13_U91  ( .A(1'b0), .ZN(_u0_u13_ch_am1[8] ) );
INV_X4 _u0_u13_U89  ( .A(1'b0), .ZN(_u0_u13_ch_am1[7] ) );
INV_X4 _u0_u13_U87  ( .A(1'b0), .ZN(_u0_u13_ch_am1[6] ) );
INV_X4 _u0_u13_U85  ( .A(1'b0), .ZN(_u0_u13_ch_am1[5] ) );
INV_X4 _u0_u13_U83  ( .A(1'b0), .ZN(_u0_u13_ch_am1[4] ) );
INV_X4 _u0_u13_U81  ( .A(1'b1), .ZN(_u0_u13_ch_am1[3] ) );
INV_X4 _u0_u13_U79  ( .A(1'b1), .ZN(_u0_u13_ch_am1[2] ) );
INV_X4 _u0_u13_U77  ( .A(1'b1), .ZN(_u0_u13_ch_am1[1] ) );
INV_X4 _u0_u13_U75  ( .A(1'b1), .ZN(_u0_u13_ch_am1[0] ) );
INV_X4 _u0_u13_U73  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[31] ) );
INV_X4 _u0_u13_U71  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[30] ) );
INV_X4 _u0_u13_U69  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[29] ) );
INV_X4 _u0_u13_U67  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[28] ) );
INV_X4 _u0_u13_U65  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[27] ) );
INV_X4 _u0_u13_U63  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[26] ) );
INV_X4 _u0_u13_U61  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[25] ) );
INV_X4 _u0_u13_U59  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[24] ) );
INV_X4 _u0_u13_U57  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[23] ) );
INV_X4 _u0_u13_U55  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[22] ) );
INV_X4 _u0_u13_U53  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[21] ) );
INV_X4 _u0_u13_U51  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[20] ) );
INV_X4 _u0_u13_U49  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[19] ) );
INV_X4 _u0_u13_U47  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[18] ) );
INV_X4 _u0_u13_U45  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[17] ) );
INV_X4 _u0_u13_U43  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[16] ) );
INV_X4 _u0_u13_U41  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[15] ) );
INV_X4 _u0_u13_U39  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[14] ) );
INV_X4 _u0_u13_U37  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[13] ) );
INV_X4 _u0_u13_U35  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[12] ) );
INV_X4 _u0_u13_U33  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[11] ) );
INV_X4 _u0_u13_U31  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[10] ) );
INV_X4 _u0_u13_U29  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[9] ) );
INV_X4 _u0_u13_U27  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[8] ) );
INV_X4 _u0_u13_U25  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[7] ) );
INV_X4 _u0_u13_U23  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[6] ) );
INV_X4 _u0_u13_U21  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[5] ) );
INV_X4 _u0_u13_U19  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[4] ) );
INV_X4 _u0_u13_U17  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[3] ) );
INV_X4 _u0_u13_U15  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[2] ) );
INV_X4 _u0_u13_U13  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[1] ) );
INV_X4 _u0_u13_U11  ( .A(1'b1), .ZN(_u0_u13_sw_pointer[0] ) );
INV_X4 _u0_u13_U9  ( .A(1'b1), .ZN(_u0_u13_ch_stop ) );
INV_X4 _u0_u13_U7  ( .A(1'b1), .ZN(_u0_u13_ch_dis ) );
INV_X4 _u0_u13_U5  ( .A(1'b1), .ZN(_u0_u13_int ) );
INV_X4 _u0_u14_U585  ( .A(1'b1), .ZN(_u0_u14_pointer[31] ) );
INV_X4 _u0_u14_U583  ( .A(1'b1), .ZN(_u0_u14_pointer[30] ) );
INV_X4 _u0_u14_U581  ( .A(1'b1), .ZN(_u0_u14_pointer[29] ) );
INV_X4 _u0_u14_U579  ( .A(1'b1), .ZN(_u0_u14_pointer[28] ) );
INV_X4 _u0_u14_U577  ( .A(1'b1), .ZN(_u0_u14_pointer[27] ) );
INV_X4 _u0_u14_U575  ( .A(1'b1), .ZN(_u0_u14_pointer[26] ) );
INV_X4 _u0_u14_U573  ( .A(1'b1), .ZN(_u0_u14_pointer[25] ) );
INV_X4 _u0_u14_U571  ( .A(1'b1), .ZN(_u0_u14_pointer[24] ) );
INV_X4 _u0_u14_U569  ( .A(1'b1), .ZN(_u0_u14_pointer[23] ) );
INV_X4 _u0_u14_U567  ( .A(1'b1), .ZN(_u0_u14_pointer[22] ) );
INV_X4 _u0_u14_U565  ( .A(1'b1), .ZN(_u0_u14_pointer[21] ) );
INV_X4 _u0_u14_U563  ( .A(1'b1), .ZN(_u0_u14_pointer[20] ) );
INV_X4 _u0_u14_U561  ( .A(1'b1), .ZN(_u0_u14_pointer[19] ) );
INV_X4 _u0_u14_U559  ( .A(1'b1), .ZN(_u0_u14_pointer[18] ) );
INV_X4 _u0_u14_U557  ( .A(1'b1), .ZN(_u0_u14_pointer[17] ) );
INV_X4 _u0_u14_U555  ( .A(1'b1), .ZN(_u0_u14_pointer[16] ) );
INV_X4 _u0_u14_U553  ( .A(1'b1), .ZN(_u0_u14_pointer[15] ) );
INV_X4 _u0_u14_U551  ( .A(1'b1), .ZN(_u0_u14_pointer[14] ) );
INV_X4 _u0_u14_U549  ( .A(1'b1), .ZN(_u0_u14_pointer[13] ) );
INV_X4 _u0_u14_U547  ( .A(1'b1), .ZN(_u0_u14_pointer[12] ) );
INV_X4 _u0_u14_U545  ( .A(1'b1), .ZN(_u0_u14_pointer[11] ) );
INV_X4 _u0_u14_U543  ( .A(1'b1), .ZN(_u0_u14_pointer[10] ) );
INV_X4 _u0_u14_U541  ( .A(1'b1), .ZN(_u0_u14_pointer[9] ) );
INV_X4 _u0_u14_U539  ( .A(1'b1), .ZN(_u0_u14_pointer[8] ) );
INV_X4 _u0_u14_U537  ( .A(1'b1), .ZN(_u0_u14_pointer[7] ) );
INV_X4 _u0_u14_U535  ( .A(1'b1), .ZN(_u0_u14_pointer[6] ) );
INV_X4 _u0_u14_U533  ( .A(1'b1), .ZN(_u0_u14_pointer[5] ) );
INV_X4 _u0_u14_U531  ( .A(1'b1), .ZN(_u0_u14_pointer[4] ) );
INV_X4 _u0_u14_U529  ( .A(1'b1), .ZN(_u0_u14_pointer[3] ) );
INV_X4 _u0_u14_U527  ( .A(1'b1), .ZN(_u0_u14_pointer[2] ) );
INV_X4 _u0_u14_U525  ( .A(1'b1), .ZN(_u0_u14_pointer[1] ) );
INV_X4 _u0_u14_U523  ( .A(1'b1), .ZN(_u0_u14_pointer[0] ) );
INV_X4 _u0_u14_U521  ( .A(1'b1), .ZN(_u0_u14_pointer_s[31] ) );
INV_X4 _u0_u14_U519  ( .A(1'b1), .ZN(_u0_u14_pointer_s[30] ) );
INV_X4 _u0_u14_U517  ( .A(1'b1), .ZN(_u0_u14_pointer_s[29] ) );
INV_X4 _u0_u14_U515  ( .A(1'b1), .ZN(_u0_u14_pointer_s[28] ) );
INV_X4 _u0_u14_U513  ( .A(1'b1), .ZN(_u0_u14_pointer_s[27] ) );
INV_X4 _u0_u14_U511  ( .A(1'b1), .ZN(_u0_u14_pointer_s[26] ) );
INV_X4 _u0_u14_U509  ( .A(1'b1), .ZN(_u0_u14_pointer_s[25] ) );
INV_X4 _u0_u14_U507  ( .A(1'b1), .ZN(_u0_u14_pointer_s[24] ) );
INV_X4 _u0_u14_U505  ( .A(1'b1), .ZN(_u0_u14_pointer_s[23] ) );
INV_X4 _u0_u14_U503  ( .A(1'b1), .ZN(_u0_u14_pointer_s[22] ) );
INV_X4 _u0_u14_U501  ( .A(1'b1), .ZN(_u0_u14_pointer_s[21] ) );
INV_X4 _u0_u14_U499  ( .A(1'b1), .ZN(_u0_u14_pointer_s[20] ) );
INV_X4 _u0_u14_U497  ( .A(1'b1), .ZN(_u0_u14_pointer_s[19] ) );
INV_X4 _u0_u14_U495  ( .A(1'b1), .ZN(_u0_u14_pointer_s[18] ) );
INV_X4 _u0_u14_U493  ( .A(1'b1), .ZN(_u0_u14_pointer_s[17] ) );
INV_X4 _u0_u14_U491  ( .A(1'b1), .ZN(_u0_u14_pointer_s[16] ) );
INV_X4 _u0_u14_U489  ( .A(1'b1), .ZN(_u0_u14_pointer_s[15] ) );
INV_X4 _u0_u14_U487  ( .A(1'b1), .ZN(_u0_u14_pointer_s[14] ) );
INV_X4 _u0_u14_U485  ( .A(1'b1), .ZN(_u0_u14_pointer_s[13] ) );
INV_X4 _u0_u14_U483  ( .A(1'b1), .ZN(_u0_u14_pointer_s[12] ) );
INV_X4 _u0_u14_U481  ( .A(1'b1), .ZN(_u0_u14_pointer_s[11] ) );
INV_X4 _u0_u14_U479  ( .A(1'b1), .ZN(_u0_u14_pointer_s[10] ) );
INV_X4 _u0_u14_U477  ( .A(1'b1), .ZN(_u0_u14_pointer_s[9] ) );
INV_X4 _u0_u14_U475  ( .A(1'b1), .ZN(_u0_u14_pointer_s[8] ) );
INV_X4 _u0_u14_U473  ( .A(1'b1), .ZN(_u0_u14_pointer_s[7] ) );
INV_X4 _u0_u14_U471  ( .A(1'b1), .ZN(_u0_u14_pointer_s[6] ) );
INV_X4 _u0_u14_U469  ( .A(1'b1), .ZN(_u0_u14_pointer_s[5] ) );
INV_X4 _u0_u14_U467  ( .A(1'b1), .ZN(_u0_u14_pointer_s[4] ) );
INV_X4 _u0_u14_U465  ( .A(1'b1), .ZN(_u0_u14_pointer_s[3] ) );
INV_X4 _u0_u14_U463  ( .A(1'b1), .ZN(_u0_u14_pointer_s[2] ) );
INV_X4 _u0_u14_U461  ( .A(1'b1), .ZN(_u0_u14_pointer_s[1] ) );
INV_X4 _u0_u14_U459  ( .A(1'b1), .ZN(_u0_u14_pointer_s[0] ) );
INV_X4 _u0_u14_U457  ( .A(1'b1), .ZN(_u0_u14_ch_csr[31] ) );
INV_X4 _u0_u14_U455  ( .A(1'b1), .ZN(_u0_u14_ch_csr[30] ) );
INV_X4 _u0_u14_U453  ( .A(1'b1), .ZN(_u0_u14_ch_csr[29] ) );
INV_X4 _u0_u14_U451  ( .A(1'b1), .ZN(_u0_u14_ch_csr[28] ) );
INV_X4 _u0_u14_U449  ( .A(1'b1), .ZN(_u0_u14_ch_csr[27] ) );
INV_X4 _u0_u14_U447  ( .A(1'b1), .ZN(_u0_u14_ch_csr[26] ) );
INV_X4 _u0_u14_U445  ( .A(1'b1), .ZN(_u0_u14_ch_csr[25] ) );
INV_X4 _u0_u14_U443  ( .A(1'b1), .ZN(_u0_u14_ch_csr[24] ) );
INV_X4 _u0_u14_U441  ( .A(1'b1), .ZN(_u0_u14_ch_csr[23] ) );
INV_X4 _u0_u14_U439  ( .A(1'b1), .ZN(_u0_u14_ch_csr[22] ) );
INV_X4 _u0_u14_U437  ( .A(1'b1), .ZN(_u0_u14_ch_csr[21] ) );
INV_X4 _u0_u14_U435  ( .A(1'b1), .ZN(_u0_u14_ch_csr[20] ) );
INV_X4 _u0_u14_U433  ( .A(1'b1), .ZN(_u0_u14_ch_csr[19] ) );
INV_X4 _u0_u14_U431  ( .A(1'b1), .ZN(_u0_u14_ch_csr[18] ) );
INV_X4 _u0_u14_U429  ( .A(1'b1), .ZN(_u0_u14_ch_csr[17] ) );
INV_X4 _u0_u14_U427  ( .A(1'b1), .ZN(_u0_u14_ch_csr[16] ) );
INV_X4 _u0_u14_U425  ( .A(1'b1), .ZN(_u0_u14_ch_csr[15] ) );
INV_X4 _u0_u14_U423  ( .A(1'b1), .ZN(_u0_u14_ch_csr[14] ) );
INV_X4 _u0_u14_U421  ( .A(1'b1), .ZN(_u0_u14_ch_csr[13] ) );
INV_X4 _u0_u14_U419  ( .A(1'b1), .ZN(_u0_u14_ch_csr[12] ) );
INV_X4 _u0_u14_U417  ( .A(1'b1), .ZN(_u0_u14_ch_csr[11] ) );
INV_X4 _u0_u14_U415  ( .A(1'b1), .ZN(_u0_u14_ch_csr[10] ) );
INV_X4 _u0_u14_U413  ( .A(1'b1), .ZN(_u0_u14_ch_csr[9] ) );
INV_X4 _u0_u14_U411  ( .A(1'b1), .ZN(_u0_u14_ch_csr[8] ) );
INV_X4 _u0_u14_U409  ( .A(1'b1), .ZN(_u0_u14_ch_csr[7] ) );
INV_X4 _u0_u14_U407  ( .A(1'b1), .ZN(_u0_u14_ch_csr[6] ) );
INV_X4 _u0_u14_U405  ( .A(1'b1), .ZN(_u0_u14_ch_csr[5] ) );
INV_X4 _u0_u14_U403  ( .A(1'b1), .ZN(_u0_u14_ch_csr[4] ) );
INV_X4 _u0_u14_U401  ( .A(1'b1), .ZN(_u0_u14_ch_csr[3] ) );
INV_X4 _u0_u14_U399  ( .A(1'b1), .ZN(_u0_u14_ch_csr[2] ) );
INV_X4 _u0_u14_U397  ( .A(1'b1), .ZN(_u0_u14_ch_csr[1] ) );
INV_X4 _u0_u14_U395  ( .A(1'b1), .ZN(_u0_u14_ch_csr[0] ) );
INV_X4 _u0_u14_U393  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[31] ) );
INV_X4 _u0_u14_U391  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[30] ) );
INV_X4 _u0_u14_U389  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[29] ) );
INV_X4 _u0_u14_U387  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[28] ) );
INV_X4 _u0_u14_U385  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[27] ) );
INV_X4 _u0_u14_U383  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[26] ) );
INV_X4 _u0_u14_U381  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[25] ) );
INV_X4 _u0_u14_U379  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[24] ) );
INV_X4 _u0_u14_U377  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[23] ) );
INV_X4 _u0_u14_U375  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[22] ) );
INV_X4 _u0_u14_U373  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[21] ) );
INV_X4 _u0_u14_U371  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[20] ) );
INV_X4 _u0_u14_U369  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[19] ) );
INV_X4 _u0_u14_U367  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[18] ) );
INV_X4 _u0_u14_U365  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[17] ) );
INV_X4 _u0_u14_U363  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[16] ) );
INV_X4 _u0_u14_U361  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[15] ) );
INV_X4 _u0_u14_U359  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[14] ) );
INV_X4 _u0_u14_U357  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[13] ) );
INV_X4 _u0_u14_U355  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[12] ) );
INV_X4 _u0_u14_U353  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[11] ) );
INV_X4 _u0_u14_U351  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[10] ) );
INV_X4 _u0_u14_U349  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[9] ) );
INV_X4 _u0_u14_U347  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[8] ) );
INV_X4 _u0_u14_U345  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[7] ) );
INV_X4 _u0_u14_U343  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[6] ) );
INV_X4 _u0_u14_U341  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[5] ) );
INV_X4 _u0_u14_U339  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[4] ) );
INV_X4 _u0_u14_U337  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[3] ) );
INV_X4 _u0_u14_U335  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[2] ) );
INV_X4 _u0_u14_U333  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[1] ) );
INV_X4 _u0_u14_U331  ( .A(1'b1), .ZN(_u0_u14_ch_txsz[0] ) );
INV_X4 _u0_u14_U329  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[31] ) );
INV_X4 _u0_u14_U327  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[30] ) );
INV_X4 _u0_u14_U325  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[29] ) );
INV_X4 _u0_u14_U323  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[28] ) );
INV_X4 _u0_u14_U321  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[27] ) );
INV_X4 _u0_u14_U319  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[26] ) );
INV_X4 _u0_u14_U317  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[25] ) );
INV_X4 _u0_u14_U315  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[24] ) );
INV_X4 _u0_u14_U313  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[23] ) );
INV_X4 _u0_u14_U311  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[22] ) );
INV_X4 _u0_u14_U309  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[21] ) );
INV_X4 _u0_u14_U307  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[20] ) );
INV_X4 _u0_u14_U305  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[19] ) );
INV_X4 _u0_u14_U303  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[18] ) );
INV_X4 _u0_u14_U301  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[17] ) );
INV_X4 _u0_u14_U299  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[16] ) );
INV_X4 _u0_u14_U297  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[15] ) );
INV_X4 _u0_u14_U295  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[14] ) );
INV_X4 _u0_u14_U293  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[13] ) );
INV_X4 _u0_u14_U291  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[12] ) );
INV_X4 _u0_u14_U289  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[11] ) );
INV_X4 _u0_u14_U287  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[10] ) );
INV_X4 _u0_u14_U285  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[9] ) );
INV_X4 _u0_u14_U283  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[8] ) );
INV_X4 _u0_u14_U281  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[7] ) );
INV_X4 _u0_u14_U279  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[6] ) );
INV_X4 _u0_u14_U277  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[5] ) );
INV_X4 _u0_u14_U275  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[4] ) );
INV_X4 _u0_u14_U273  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[3] ) );
INV_X4 _u0_u14_U271  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[2] ) );
INV_X4 _u0_u14_U269  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[1] ) );
INV_X4 _u0_u14_U267  ( .A(1'b1), .ZN(_u0_u14_ch_adr0[0] ) );
INV_X4 _u0_u14_U265  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[31] ) );
INV_X4 _u0_u14_U263  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[30] ) );
INV_X4 _u0_u14_U261  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[29] ) );
INV_X4 _u0_u14_U259  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[28] ) );
INV_X4 _u0_u14_U257  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[27] ) );
INV_X4 _u0_u14_U255  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[26] ) );
INV_X4 _u0_u14_U253  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[25] ) );
INV_X4 _u0_u14_U251  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[24] ) );
INV_X4 _u0_u14_U249  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[23] ) );
INV_X4 _u0_u14_U247  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[22] ) );
INV_X4 _u0_u14_U245  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[21] ) );
INV_X4 _u0_u14_U243  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[20] ) );
INV_X4 _u0_u14_U241  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[19] ) );
INV_X4 _u0_u14_U239  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[18] ) );
INV_X4 _u0_u14_U237  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[17] ) );
INV_X4 _u0_u14_U235  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[16] ) );
INV_X4 _u0_u14_U233  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[15] ) );
INV_X4 _u0_u14_U231  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[14] ) );
INV_X4 _u0_u14_U229  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[13] ) );
INV_X4 _u0_u14_U227  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[12] ) );
INV_X4 _u0_u14_U225  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[11] ) );
INV_X4 _u0_u14_U223  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[10] ) );
INV_X4 _u0_u14_U221  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[9] ) );
INV_X4 _u0_u14_U219  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[8] ) );
INV_X4 _u0_u14_U217  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[7] ) );
INV_X4 _u0_u14_U215  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[6] ) );
INV_X4 _u0_u14_U213  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[5] ) );
INV_X4 _u0_u14_U211  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[4] ) );
INV_X4 _u0_u14_U209  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[3] ) );
INV_X4 _u0_u14_U207  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[2] ) );
INV_X4 _u0_u14_U205  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[1] ) );
INV_X4 _u0_u14_U203  ( .A(1'b1), .ZN(_u0_u14_ch_adr1[0] ) );
INV_X4 _u0_u14_U201  ( .A(1'b0), .ZN(_u0_u14_ch_am0[31] ) );
INV_X4 _u0_u14_U199  ( .A(1'b0), .ZN(_u0_u14_ch_am0[30] ) );
INV_X4 _u0_u14_U197  ( .A(1'b0), .ZN(_u0_u14_ch_am0[29] ) );
INV_X4 _u0_u14_U195  ( .A(1'b0), .ZN(_u0_u14_ch_am0[28] ) );
INV_X4 _u0_u14_U193  ( .A(1'b0), .ZN(_u0_u14_ch_am0[27] ) );
INV_X4 _u0_u14_U191  ( .A(1'b0), .ZN(_u0_u14_ch_am0[26] ) );
INV_X4 _u0_u14_U189  ( .A(1'b0), .ZN(_u0_u14_ch_am0[25] ) );
INV_X4 _u0_u14_U187  ( .A(1'b0), .ZN(_u0_u14_ch_am0[24] ) );
INV_X4 _u0_u14_U185  ( .A(1'b0), .ZN(_u0_u14_ch_am0[23] ) );
INV_X4 _u0_u14_U183  ( .A(1'b0), .ZN(_u0_u14_ch_am0[22] ) );
INV_X4 _u0_u14_U181  ( .A(1'b0), .ZN(_u0_u14_ch_am0[21] ) );
INV_X4 _u0_u14_U179  ( .A(1'b0), .ZN(_u0_u14_ch_am0[20] ) );
INV_X4 _u0_u14_U177  ( .A(1'b0), .ZN(_u0_u14_ch_am0[19] ) );
INV_X4 _u0_u14_U175  ( .A(1'b0), .ZN(_u0_u14_ch_am0[18] ) );
INV_X4 _u0_u14_U173  ( .A(1'b0), .ZN(_u0_u14_ch_am0[17] ) );
INV_X4 _u0_u14_U171  ( .A(1'b0), .ZN(_u0_u14_ch_am0[16] ) );
INV_X4 _u0_u14_U169  ( .A(1'b0), .ZN(_u0_u14_ch_am0[15] ) );
INV_X4 _u0_u14_U167  ( .A(1'b0), .ZN(_u0_u14_ch_am0[14] ) );
INV_X4 _u0_u14_U165  ( .A(1'b0), .ZN(_u0_u14_ch_am0[13] ) );
INV_X4 _u0_u14_U163  ( .A(1'b0), .ZN(_u0_u14_ch_am0[12] ) );
INV_X4 _u0_u14_U161  ( .A(1'b0), .ZN(_u0_u14_ch_am0[11] ) );
INV_X4 _u0_u14_U159  ( .A(1'b0), .ZN(_u0_u14_ch_am0[10] ) );
INV_X4 _u0_u14_U157  ( .A(1'b0), .ZN(_u0_u14_ch_am0[9] ) );
INV_X4 _u0_u14_U155  ( .A(1'b0), .ZN(_u0_u14_ch_am0[8] ) );
INV_X4 _u0_u14_U153  ( .A(1'b0), .ZN(_u0_u14_ch_am0[7] ) );
INV_X4 _u0_u14_U151  ( .A(1'b0), .ZN(_u0_u14_ch_am0[6] ) );
INV_X4 _u0_u14_U149  ( .A(1'b0), .ZN(_u0_u14_ch_am0[5] ) );
INV_X4 _u0_u14_U147  ( .A(1'b0), .ZN(_u0_u14_ch_am0[4] ) );
INV_X4 _u0_u14_U145  ( .A(1'b1), .ZN(_u0_u14_ch_am0[3] ) );
INV_X4 _u0_u14_U143  ( .A(1'b1), .ZN(_u0_u14_ch_am0[2] ) );
INV_X4 _u0_u14_U141  ( .A(1'b1), .ZN(_u0_u14_ch_am0[1] ) );
INV_X4 _u0_u14_U139  ( .A(1'b1), .ZN(_u0_u14_ch_am0[0] ) );
INV_X4 _u0_u14_U137  ( .A(1'b0), .ZN(_u0_u14_ch_am1[31] ) );
INV_X4 _u0_u14_U135  ( .A(1'b0), .ZN(_u0_u14_ch_am1[30] ) );
INV_X4 _u0_u14_U133  ( .A(1'b0), .ZN(_u0_u14_ch_am1[29] ) );
INV_X4 _u0_u14_U131  ( .A(1'b0), .ZN(_u0_u14_ch_am1[28] ) );
INV_X4 _u0_u14_U129  ( .A(1'b0), .ZN(_u0_u14_ch_am1[27] ) );
INV_X4 _u0_u14_U127  ( .A(1'b0), .ZN(_u0_u14_ch_am1[26] ) );
INV_X4 _u0_u14_U125  ( .A(1'b0), .ZN(_u0_u14_ch_am1[25] ) );
INV_X4 _u0_u14_U123  ( .A(1'b0), .ZN(_u0_u14_ch_am1[24] ) );
INV_X4 _u0_u14_U121  ( .A(1'b0), .ZN(_u0_u14_ch_am1[23] ) );
INV_X4 _u0_u14_U119  ( .A(1'b0), .ZN(_u0_u14_ch_am1[22] ) );
INV_X4 _u0_u14_U117  ( .A(1'b0), .ZN(_u0_u14_ch_am1[21] ) );
INV_X4 _u0_u14_U115  ( .A(1'b0), .ZN(_u0_u14_ch_am1[20] ) );
INV_X4 _u0_u14_U113  ( .A(1'b0), .ZN(_u0_u14_ch_am1[19] ) );
INV_X4 _u0_u14_U111  ( .A(1'b0), .ZN(_u0_u14_ch_am1[18] ) );
INV_X4 _u0_u14_U109  ( .A(1'b0), .ZN(_u0_u14_ch_am1[17] ) );
INV_X4 _u0_u14_U107  ( .A(1'b0), .ZN(_u0_u14_ch_am1[16] ) );
INV_X4 _u0_u14_U105  ( .A(1'b0), .ZN(_u0_u14_ch_am1[15] ) );
INV_X4 _u0_u14_U103  ( .A(1'b0), .ZN(_u0_u14_ch_am1[14] ) );
INV_X4 _u0_u14_U101  ( .A(1'b0), .ZN(_u0_u14_ch_am1[13] ) );
INV_X4 _u0_u14_U99  ( .A(1'b0), .ZN(_u0_u14_ch_am1[12] ) );
INV_X4 _u0_u14_U97  ( .A(1'b0), .ZN(_u0_u14_ch_am1[11] ) );
INV_X4 _u0_u14_U95  ( .A(1'b0), .ZN(_u0_u14_ch_am1[10] ) );
INV_X4 _u0_u14_U93  ( .A(1'b0), .ZN(_u0_u14_ch_am1[9] ) );
INV_X4 _u0_u14_U91  ( .A(1'b0), .ZN(_u0_u14_ch_am1[8] ) );
INV_X4 _u0_u14_U89  ( .A(1'b0), .ZN(_u0_u14_ch_am1[7] ) );
INV_X4 _u0_u14_U87  ( .A(1'b0), .ZN(_u0_u14_ch_am1[6] ) );
INV_X4 _u0_u14_U85  ( .A(1'b0), .ZN(_u0_u14_ch_am1[5] ) );
INV_X4 _u0_u14_U83  ( .A(1'b0), .ZN(_u0_u14_ch_am1[4] ) );
INV_X4 _u0_u14_U81  ( .A(1'b1), .ZN(_u0_u14_ch_am1[3] ) );
INV_X4 _u0_u14_U79  ( .A(1'b1), .ZN(_u0_u14_ch_am1[2] ) );
INV_X4 _u0_u14_U77  ( .A(1'b1), .ZN(_u0_u14_ch_am1[1] ) );
INV_X4 _u0_u14_U75  ( .A(1'b1), .ZN(_u0_u14_ch_am1[0] ) );
INV_X4 _u0_u14_U73  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[31] ) );
INV_X4 _u0_u14_U71  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[30] ) );
INV_X4 _u0_u14_U69  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[29] ) );
INV_X4 _u0_u14_U67  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[28] ) );
INV_X4 _u0_u14_U65  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[27] ) );
INV_X4 _u0_u14_U63  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[26] ) );
INV_X4 _u0_u14_U61  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[25] ) );
INV_X4 _u0_u14_U59  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[24] ) );
INV_X4 _u0_u14_U57  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[23] ) );
INV_X4 _u0_u14_U55  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[22] ) );
INV_X4 _u0_u14_U53  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[21] ) );
INV_X4 _u0_u14_U51  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[20] ) );
INV_X4 _u0_u14_U49  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[19] ) );
INV_X4 _u0_u14_U47  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[18] ) );
INV_X4 _u0_u14_U45  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[17] ) );
INV_X4 _u0_u14_U43  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[16] ) );
INV_X4 _u0_u14_U41  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[15] ) );
INV_X4 _u0_u14_U39  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[14] ) );
INV_X4 _u0_u14_U37  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[13] ) );
INV_X4 _u0_u14_U35  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[12] ) );
INV_X4 _u0_u14_U33  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[11] ) );
INV_X4 _u0_u14_U31  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[10] ) );
INV_X4 _u0_u14_U29  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[9] ) );
INV_X4 _u0_u14_U27  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[8] ) );
INV_X4 _u0_u14_U25  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[7] ) );
INV_X4 _u0_u14_U23  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[6] ) );
INV_X4 _u0_u14_U21  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[5] ) );
INV_X4 _u0_u14_U19  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[4] ) );
INV_X4 _u0_u14_U17  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[3] ) );
INV_X4 _u0_u14_U15  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[2] ) );
INV_X4 _u0_u14_U13  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[1] ) );
INV_X4 _u0_u14_U11  ( .A(1'b1), .ZN(_u0_u14_sw_pointer[0] ) );
INV_X4 _u0_u14_U9  ( .A(1'b1), .ZN(_u0_u14_ch_stop ) );
INV_X4 _u0_u14_U7  ( .A(1'b1), .ZN(_u0_u14_ch_dis ) );
INV_X4 _u0_u14_U5  ( .A(1'b1), .ZN(_u0_u14_int ) );
INV_X4 _u0_u15_U585  ( .A(1'b1), .ZN(_u0_u15_pointer[31] ) );
INV_X4 _u0_u15_U583  ( .A(1'b1), .ZN(_u0_u15_pointer[30] ) );
INV_X4 _u0_u15_U581  ( .A(1'b1), .ZN(_u0_u15_pointer[29] ) );
INV_X4 _u0_u15_U579  ( .A(1'b1), .ZN(_u0_u15_pointer[28] ) );
INV_X4 _u0_u15_U577  ( .A(1'b1), .ZN(_u0_u15_pointer[27] ) );
INV_X4 _u0_u15_U575  ( .A(1'b1), .ZN(_u0_u15_pointer[26] ) );
INV_X4 _u0_u15_U573  ( .A(1'b1), .ZN(_u0_u15_pointer[25] ) );
INV_X4 _u0_u15_U571  ( .A(1'b1), .ZN(_u0_u15_pointer[24] ) );
INV_X4 _u0_u15_U569  ( .A(1'b1), .ZN(_u0_u15_pointer[23] ) );
INV_X4 _u0_u15_U567  ( .A(1'b1), .ZN(_u0_u15_pointer[22] ) );
INV_X4 _u0_u15_U565  ( .A(1'b1), .ZN(_u0_u15_pointer[21] ) );
INV_X4 _u0_u15_U563  ( .A(1'b1), .ZN(_u0_u15_pointer[20] ) );
INV_X4 _u0_u15_U561  ( .A(1'b1), .ZN(_u0_u15_pointer[19] ) );
INV_X4 _u0_u15_U559  ( .A(1'b1), .ZN(_u0_u15_pointer[18] ) );
INV_X4 _u0_u15_U557  ( .A(1'b1), .ZN(_u0_u15_pointer[17] ) );
INV_X4 _u0_u15_U555  ( .A(1'b1), .ZN(_u0_u15_pointer[16] ) );
INV_X4 _u0_u15_U553  ( .A(1'b1), .ZN(_u0_u15_pointer[15] ) );
INV_X4 _u0_u15_U551  ( .A(1'b1), .ZN(_u0_u15_pointer[14] ) );
INV_X4 _u0_u15_U549  ( .A(1'b1), .ZN(_u0_u15_pointer[13] ) );
INV_X4 _u0_u15_U547  ( .A(1'b1), .ZN(_u0_u15_pointer[12] ) );
INV_X4 _u0_u15_U545  ( .A(1'b1), .ZN(_u0_u15_pointer[11] ) );
INV_X4 _u0_u15_U543  ( .A(1'b1), .ZN(_u0_u15_pointer[10] ) );
INV_X4 _u0_u15_U541  ( .A(1'b1), .ZN(_u0_u15_pointer[9] ) );
INV_X4 _u0_u15_U539  ( .A(1'b1), .ZN(_u0_u15_pointer[8] ) );
INV_X4 _u0_u15_U537  ( .A(1'b1), .ZN(_u0_u15_pointer[7] ) );
INV_X4 _u0_u15_U535  ( .A(1'b1), .ZN(_u0_u15_pointer[6] ) );
INV_X4 _u0_u15_U533  ( .A(1'b1), .ZN(_u0_u15_pointer[5] ) );
INV_X4 _u0_u15_U531  ( .A(1'b1), .ZN(_u0_u15_pointer[4] ) );
INV_X4 _u0_u15_U529  ( .A(1'b1), .ZN(_u0_u15_pointer[3] ) );
INV_X4 _u0_u15_U527  ( .A(1'b1), .ZN(_u0_u15_pointer[2] ) );
INV_X4 _u0_u15_U525  ( .A(1'b1), .ZN(_u0_u15_pointer[1] ) );
INV_X4 _u0_u15_U523  ( .A(1'b1), .ZN(_u0_u15_pointer[0] ) );
INV_X4 _u0_u15_U521  ( .A(1'b1), .ZN(_u0_u15_pointer_s[31] ) );
INV_X4 _u0_u15_U519  ( .A(1'b1), .ZN(_u0_u15_pointer_s[30] ) );
INV_X4 _u0_u15_U517  ( .A(1'b1), .ZN(_u0_u15_pointer_s[29] ) );
INV_X4 _u0_u15_U515  ( .A(1'b1), .ZN(_u0_u15_pointer_s[28] ) );
INV_X4 _u0_u15_U513  ( .A(1'b1), .ZN(_u0_u15_pointer_s[27] ) );
INV_X4 _u0_u15_U511  ( .A(1'b1), .ZN(_u0_u15_pointer_s[26] ) );
INV_X4 _u0_u15_U509  ( .A(1'b1), .ZN(_u0_u15_pointer_s[25] ) );
INV_X4 _u0_u15_U507  ( .A(1'b1), .ZN(_u0_u15_pointer_s[24] ) );
INV_X4 _u0_u15_U505  ( .A(1'b1), .ZN(_u0_u15_pointer_s[23] ) );
INV_X4 _u0_u15_U503  ( .A(1'b1), .ZN(_u0_u15_pointer_s[22] ) );
INV_X4 _u0_u15_U501  ( .A(1'b1), .ZN(_u0_u15_pointer_s[21] ) );
INV_X4 _u0_u15_U499  ( .A(1'b1), .ZN(_u0_u15_pointer_s[20] ) );
INV_X4 _u0_u15_U497  ( .A(1'b1), .ZN(_u0_u15_pointer_s[19] ) );
INV_X4 _u0_u15_U495  ( .A(1'b1), .ZN(_u0_u15_pointer_s[18] ) );
INV_X4 _u0_u15_U493  ( .A(1'b1), .ZN(_u0_u15_pointer_s[17] ) );
INV_X4 _u0_u15_U491  ( .A(1'b1), .ZN(_u0_u15_pointer_s[16] ) );
INV_X4 _u0_u15_U489  ( .A(1'b1), .ZN(_u0_u15_pointer_s[15] ) );
INV_X4 _u0_u15_U487  ( .A(1'b1), .ZN(_u0_u15_pointer_s[14] ) );
INV_X4 _u0_u15_U485  ( .A(1'b1), .ZN(_u0_u15_pointer_s[13] ) );
INV_X4 _u0_u15_U483  ( .A(1'b1), .ZN(_u0_u15_pointer_s[12] ) );
INV_X4 _u0_u15_U481  ( .A(1'b1), .ZN(_u0_u15_pointer_s[11] ) );
INV_X4 _u0_u15_U479  ( .A(1'b1), .ZN(_u0_u15_pointer_s[10] ) );
INV_X4 _u0_u15_U477  ( .A(1'b1), .ZN(_u0_u15_pointer_s[9] ) );
INV_X4 _u0_u15_U475  ( .A(1'b1), .ZN(_u0_u15_pointer_s[8] ) );
INV_X4 _u0_u15_U473  ( .A(1'b1), .ZN(_u0_u15_pointer_s[7] ) );
INV_X4 _u0_u15_U471  ( .A(1'b1), .ZN(_u0_u15_pointer_s[6] ) );
INV_X4 _u0_u15_U469  ( .A(1'b1), .ZN(_u0_u15_pointer_s[5] ) );
INV_X4 _u0_u15_U467  ( .A(1'b1), .ZN(_u0_u15_pointer_s[4] ) );
INV_X4 _u0_u15_U465  ( .A(1'b1), .ZN(_u0_u15_pointer_s[3] ) );
INV_X4 _u0_u15_U463  ( .A(1'b1), .ZN(_u0_u15_pointer_s[2] ) );
INV_X4 _u0_u15_U461  ( .A(1'b1), .ZN(_u0_u15_pointer_s[1] ) );
INV_X4 _u0_u15_U459  ( .A(1'b1), .ZN(_u0_u15_pointer_s[0] ) );
INV_X4 _u0_u15_U457  ( .A(1'b1), .ZN(_u0_u15_ch_csr[31] ) );
INV_X4 _u0_u15_U455  ( .A(1'b1), .ZN(_u0_u15_ch_csr[30] ) );
INV_X4 _u0_u15_U453  ( .A(1'b1), .ZN(_u0_u15_ch_csr[29] ) );
INV_X4 _u0_u15_U451  ( .A(1'b1), .ZN(_u0_u15_ch_csr[28] ) );
INV_X4 _u0_u15_U449  ( .A(1'b1), .ZN(_u0_u15_ch_csr[27] ) );
INV_X4 _u0_u15_U447  ( .A(1'b1), .ZN(_u0_u15_ch_csr[26] ) );
INV_X4 _u0_u15_U445  ( .A(1'b1), .ZN(_u0_u15_ch_csr[25] ) );
INV_X4 _u0_u15_U443  ( .A(1'b1), .ZN(_u0_u15_ch_csr[24] ) );
INV_X4 _u0_u15_U441  ( .A(1'b1), .ZN(_u0_u15_ch_csr[23] ) );
INV_X4 _u0_u15_U439  ( .A(1'b1), .ZN(_u0_u15_ch_csr[22] ) );
INV_X4 _u0_u15_U437  ( .A(1'b1), .ZN(_u0_u15_ch_csr[21] ) );
INV_X4 _u0_u15_U435  ( .A(1'b1), .ZN(_u0_u15_ch_csr[20] ) );
INV_X4 _u0_u15_U433  ( .A(1'b1), .ZN(_u0_u15_ch_csr[19] ) );
INV_X4 _u0_u15_U431  ( .A(1'b1), .ZN(_u0_u15_ch_csr[18] ) );
INV_X4 _u0_u15_U429  ( .A(1'b1), .ZN(_u0_u15_ch_csr[17] ) );
INV_X4 _u0_u15_U427  ( .A(1'b1), .ZN(_u0_u15_ch_csr[16] ) );
INV_X4 _u0_u15_U425  ( .A(1'b1), .ZN(_u0_u15_ch_csr[15] ) );
INV_X4 _u0_u15_U423  ( .A(1'b1), .ZN(_u0_u15_ch_csr[14] ) );
INV_X4 _u0_u15_U421  ( .A(1'b1), .ZN(_u0_u15_ch_csr[13] ) );
INV_X4 _u0_u15_U419  ( .A(1'b1), .ZN(_u0_u15_ch_csr[12] ) );
INV_X4 _u0_u15_U417  ( .A(1'b1), .ZN(_u0_u15_ch_csr[11] ) );
INV_X4 _u0_u15_U415  ( .A(1'b1), .ZN(_u0_u15_ch_csr[10] ) );
INV_X4 _u0_u15_U413  ( .A(1'b1), .ZN(_u0_u15_ch_csr[9] ) );
INV_X4 _u0_u15_U411  ( .A(1'b1), .ZN(_u0_u15_ch_csr[8] ) );
INV_X4 _u0_u15_U409  ( .A(1'b1), .ZN(_u0_u15_ch_csr[7] ) );
INV_X4 _u0_u15_U407  ( .A(1'b1), .ZN(_u0_u15_ch_csr[6] ) );
INV_X4 _u0_u15_U405  ( .A(1'b1), .ZN(_u0_u15_ch_csr[5] ) );
INV_X4 _u0_u15_U403  ( .A(1'b1), .ZN(_u0_u15_ch_csr[4] ) );
INV_X4 _u0_u15_U401  ( .A(1'b1), .ZN(_u0_u15_ch_csr[3] ) );
INV_X4 _u0_u15_U399  ( .A(1'b1), .ZN(_u0_u15_ch_csr[2] ) );
INV_X4 _u0_u15_U397  ( .A(1'b1), .ZN(_u0_u15_ch_csr[1] ) );
INV_X4 _u0_u15_U395  ( .A(1'b1), .ZN(_u0_u15_ch_csr[0] ) );
INV_X4 _u0_u15_U393  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[31] ) );
INV_X4 _u0_u15_U391  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[30] ) );
INV_X4 _u0_u15_U389  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[29] ) );
INV_X4 _u0_u15_U387  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[28] ) );
INV_X4 _u0_u15_U385  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[27] ) );
INV_X4 _u0_u15_U383  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[26] ) );
INV_X4 _u0_u15_U381  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[25] ) );
INV_X4 _u0_u15_U379  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[24] ) );
INV_X4 _u0_u15_U377  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[23] ) );
INV_X4 _u0_u15_U375  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[22] ) );
INV_X4 _u0_u15_U373  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[21] ) );
INV_X4 _u0_u15_U371  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[20] ) );
INV_X4 _u0_u15_U369  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[19] ) );
INV_X4 _u0_u15_U367  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[18] ) );
INV_X4 _u0_u15_U365  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[17] ) );
INV_X4 _u0_u15_U363  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[16] ) );
INV_X4 _u0_u15_U361  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[15] ) );
INV_X4 _u0_u15_U359  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[14] ) );
INV_X4 _u0_u15_U357  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[13] ) );
INV_X4 _u0_u15_U355  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[12] ) );
INV_X4 _u0_u15_U353  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[11] ) );
INV_X4 _u0_u15_U351  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[10] ) );
INV_X4 _u0_u15_U349  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[9] ) );
INV_X4 _u0_u15_U347  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[8] ) );
INV_X4 _u0_u15_U345  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[7] ) );
INV_X4 _u0_u15_U343  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[6] ) );
INV_X4 _u0_u15_U341  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[5] ) );
INV_X4 _u0_u15_U339  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[4] ) );
INV_X4 _u0_u15_U337  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[3] ) );
INV_X4 _u0_u15_U335  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[2] ) );
INV_X4 _u0_u15_U333  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[1] ) );
INV_X4 _u0_u15_U331  ( .A(1'b1), .ZN(_u0_u15_ch_txsz[0] ) );
INV_X4 _u0_u15_U329  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[31] ) );
INV_X4 _u0_u15_U327  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[30] ) );
INV_X4 _u0_u15_U325  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[29] ) );
INV_X4 _u0_u15_U323  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[28] ) );
INV_X4 _u0_u15_U321  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[27] ) );
INV_X4 _u0_u15_U319  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[26] ) );
INV_X4 _u0_u15_U317  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[25] ) );
INV_X4 _u0_u15_U315  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[24] ) );
INV_X4 _u0_u15_U313  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[23] ) );
INV_X4 _u0_u15_U311  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[22] ) );
INV_X4 _u0_u15_U309  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[21] ) );
INV_X4 _u0_u15_U307  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[20] ) );
INV_X4 _u0_u15_U305  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[19] ) );
INV_X4 _u0_u15_U303  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[18] ) );
INV_X4 _u0_u15_U301  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[17] ) );
INV_X4 _u0_u15_U299  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[16] ) );
INV_X4 _u0_u15_U297  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[15] ) );
INV_X4 _u0_u15_U295  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[14] ) );
INV_X4 _u0_u15_U293  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[13] ) );
INV_X4 _u0_u15_U291  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[12] ) );
INV_X4 _u0_u15_U289  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[11] ) );
INV_X4 _u0_u15_U287  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[10] ) );
INV_X4 _u0_u15_U285  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[9] ) );
INV_X4 _u0_u15_U283  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[8] ) );
INV_X4 _u0_u15_U281  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[7] ) );
INV_X4 _u0_u15_U279  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[6] ) );
INV_X4 _u0_u15_U277  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[5] ) );
INV_X4 _u0_u15_U275  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[4] ) );
INV_X4 _u0_u15_U273  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[3] ) );
INV_X4 _u0_u15_U271  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[2] ) );
INV_X4 _u0_u15_U269  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[1] ) );
INV_X4 _u0_u15_U267  ( .A(1'b1), .ZN(_u0_u15_ch_adr0[0] ) );
INV_X4 _u0_u15_U265  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[31] ) );
INV_X4 _u0_u15_U263  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[30] ) );
INV_X4 _u0_u15_U261  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[29] ) );
INV_X4 _u0_u15_U259  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[28] ) );
INV_X4 _u0_u15_U257  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[27] ) );
INV_X4 _u0_u15_U255  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[26] ) );
INV_X4 _u0_u15_U253  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[25] ) );
INV_X4 _u0_u15_U251  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[24] ) );
INV_X4 _u0_u15_U249  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[23] ) );
INV_X4 _u0_u15_U247  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[22] ) );
INV_X4 _u0_u15_U245  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[21] ) );
INV_X4 _u0_u15_U243  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[20] ) );
INV_X4 _u0_u15_U241  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[19] ) );
INV_X4 _u0_u15_U239  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[18] ) );
INV_X4 _u0_u15_U237  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[17] ) );
INV_X4 _u0_u15_U235  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[16] ) );
INV_X4 _u0_u15_U233  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[15] ) );
INV_X4 _u0_u15_U231  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[14] ) );
INV_X4 _u0_u15_U229  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[13] ) );
INV_X4 _u0_u15_U227  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[12] ) );
INV_X4 _u0_u15_U225  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[11] ) );
INV_X4 _u0_u15_U223  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[10] ) );
INV_X4 _u0_u15_U221  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[9] ) );
INV_X4 _u0_u15_U219  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[8] ) );
INV_X4 _u0_u15_U217  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[7] ) );
INV_X4 _u0_u15_U215  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[6] ) );
INV_X4 _u0_u15_U213  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[5] ) );
INV_X4 _u0_u15_U211  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[4] ) );
INV_X4 _u0_u15_U209  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[3] ) );
INV_X4 _u0_u15_U207  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[2] ) );
INV_X4 _u0_u15_U205  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[1] ) );
INV_X4 _u0_u15_U203  ( .A(1'b1), .ZN(_u0_u15_ch_adr1[0] ) );
INV_X4 _u0_u15_U201  ( .A(1'b0), .ZN(_u0_u15_ch_am0[31] ) );
INV_X4 _u0_u15_U199  ( .A(1'b0), .ZN(_u0_u15_ch_am0[30] ) );
INV_X4 _u0_u15_U197  ( .A(1'b0), .ZN(_u0_u15_ch_am0[29] ) );
INV_X4 _u0_u15_U195  ( .A(1'b0), .ZN(_u0_u15_ch_am0[28] ) );
INV_X4 _u0_u15_U193  ( .A(1'b0), .ZN(_u0_u15_ch_am0[27] ) );
INV_X4 _u0_u15_U191  ( .A(1'b0), .ZN(_u0_u15_ch_am0[26] ) );
INV_X4 _u0_u15_U189  ( .A(1'b0), .ZN(_u0_u15_ch_am0[25] ) );
INV_X4 _u0_u15_U187  ( .A(1'b0), .ZN(_u0_u15_ch_am0[24] ) );
INV_X4 _u0_u15_U185  ( .A(1'b0), .ZN(_u0_u15_ch_am0[23] ) );
INV_X4 _u0_u15_U183  ( .A(1'b0), .ZN(_u0_u15_ch_am0[22] ) );
INV_X4 _u0_u15_U181  ( .A(1'b0), .ZN(_u0_u15_ch_am0[21] ) );
INV_X4 _u0_u15_U179  ( .A(1'b0), .ZN(_u0_u15_ch_am0[20] ) );
INV_X4 _u0_u15_U177  ( .A(1'b0), .ZN(_u0_u15_ch_am0[19] ) );
INV_X4 _u0_u15_U175  ( .A(1'b0), .ZN(_u0_u15_ch_am0[18] ) );
INV_X4 _u0_u15_U173  ( .A(1'b0), .ZN(_u0_u15_ch_am0[17] ) );
INV_X4 _u0_u15_U171  ( .A(1'b0), .ZN(_u0_u15_ch_am0[16] ) );
INV_X4 _u0_u15_U169  ( .A(1'b0), .ZN(_u0_u15_ch_am0[15] ) );
INV_X4 _u0_u15_U167  ( .A(1'b0), .ZN(_u0_u15_ch_am0[14] ) );
INV_X4 _u0_u15_U165  ( .A(1'b0), .ZN(_u0_u15_ch_am0[13] ) );
INV_X4 _u0_u15_U163  ( .A(1'b0), .ZN(_u0_u15_ch_am0[12] ) );
INV_X4 _u0_u15_U161  ( .A(1'b0), .ZN(_u0_u15_ch_am0[11] ) );
INV_X4 _u0_u15_U159  ( .A(1'b0), .ZN(_u0_u15_ch_am0[10] ) );
INV_X4 _u0_u15_U157  ( .A(1'b0), .ZN(_u0_u15_ch_am0[9] ) );
INV_X4 _u0_u15_U155  ( .A(1'b0), .ZN(_u0_u15_ch_am0[8] ) );
INV_X4 _u0_u15_U153  ( .A(1'b0), .ZN(_u0_u15_ch_am0[7] ) );
INV_X4 _u0_u15_U151  ( .A(1'b0), .ZN(_u0_u15_ch_am0[6] ) );
INV_X4 _u0_u15_U149  ( .A(1'b0), .ZN(_u0_u15_ch_am0[5] ) );
INV_X4 _u0_u15_U147  ( .A(1'b0), .ZN(_u0_u15_ch_am0[4] ) );
INV_X4 _u0_u15_U145  ( .A(1'b1), .ZN(_u0_u15_ch_am0[3] ) );
INV_X4 _u0_u15_U143  ( .A(1'b1), .ZN(_u0_u15_ch_am0[2] ) );
INV_X4 _u0_u15_U141  ( .A(1'b1), .ZN(_u0_u15_ch_am0[1] ) );
INV_X4 _u0_u15_U139  ( .A(1'b1), .ZN(_u0_u15_ch_am0[0] ) );
INV_X4 _u0_u15_U137  ( .A(1'b0), .ZN(_u0_u15_ch_am1[31] ) );
INV_X4 _u0_u15_U135  ( .A(1'b0), .ZN(_u0_u15_ch_am1[30] ) );
INV_X4 _u0_u15_U133  ( .A(1'b0), .ZN(_u0_u15_ch_am1[29] ) );
INV_X4 _u0_u15_U131  ( .A(1'b0), .ZN(_u0_u15_ch_am1[28] ) );
INV_X4 _u0_u15_U129  ( .A(1'b0), .ZN(_u0_u15_ch_am1[27] ) );
INV_X4 _u0_u15_U127  ( .A(1'b0), .ZN(_u0_u15_ch_am1[26] ) );
INV_X4 _u0_u15_U125  ( .A(1'b0), .ZN(_u0_u15_ch_am1[25] ) );
INV_X4 _u0_u15_U123  ( .A(1'b0), .ZN(_u0_u15_ch_am1[24] ) );
INV_X4 _u0_u15_U121  ( .A(1'b0), .ZN(_u0_u15_ch_am1[23] ) );
INV_X4 _u0_u15_U119  ( .A(1'b0), .ZN(_u0_u15_ch_am1[22] ) );
INV_X4 _u0_u15_U117  ( .A(1'b0), .ZN(_u0_u15_ch_am1[21] ) );
INV_X4 _u0_u15_U115  ( .A(1'b0), .ZN(_u0_u15_ch_am1[20] ) );
INV_X4 _u0_u15_U113  ( .A(1'b0), .ZN(_u0_u15_ch_am1[19] ) );
INV_X4 _u0_u15_U111  ( .A(1'b0), .ZN(_u0_u15_ch_am1[18] ) );
INV_X4 _u0_u15_U109  ( .A(1'b0), .ZN(_u0_u15_ch_am1[17] ) );
INV_X4 _u0_u15_U107  ( .A(1'b0), .ZN(_u0_u15_ch_am1[16] ) );
INV_X4 _u0_u15_U105  ( .A(1'b0), .ZN(_u0_u15_ch_am1[15] ) );
INV_X4 _u0_u15_U103  ( .A(1'b0), .ZN(_u0_u15_ch_am1[14] ) );
INV_X4 _u0_u15_U101  ( .A(1'b0), .ZN(_u0_u15_ch_am1[13] ) );
INV_X4 _u0_u15_U99  ( .A(1'b0), .ZN(_u0_u15_ch_am1[12] ) );
INV_X4 _u0_u15_U97  ( .A(1'b0), .ZN(_u0_u15_ch_am1[11] ) );
INV_X4 _u0_u15_U95  ( .A(1'b0), .ZN(_u0_u15_ch_am1[10] ) );
INV_X4 _u0_u15_U93  ( .A(1'b0), .ZN(_u0_u15_ch_am1[9] ) );
INV_X4 _u0_u15_U91  ( .A(1'b0), .ZN(_u0_u15_ch_am1[8] ) );
INV_X4 _u0_u15_U89  ( .A(1'b0), .ZN(_u0_u15_ch_am1[7] ) );
INV_X4 _u0_u15_U87  ( .A(1'b0), .ZN(_u0_u15_ch_am1[6] ) );
INV_X4 _u0_u15_U85  ( .A(1'b0), .ZN(_u0_u15_ch_am1[5] ) );
INV_X4 _u0_u15_U83  ( .A(1'b0), .ZN(_u0_u15_ch_am1[4] ) );
INV_X4 _u0_u15_U81  ( .A(1'b1), .ZN(_u0_u15_ch_am1[3] ) );
INV_X4 _u0_u15_U79  ( .A(1'b1), .ZN(_u0_u15_ch_am1[2] ) );
INV_X4 _u0_u15_U77  ( .A(1'b1), .ZN(_u0_u15_ch_am1[1] ) );
INV_X4 _u0_u15_U75  ( .A(1'b1), .ZN(_u0_u15_ch_am1[0] ) );
INV_X4 _u0_u15_U73  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[31] ) );
INV_X4 _u0_u15_U71  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[30] ) );
INV_X4 _u0_u15_U69  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[29] ) );
INV_X4 _u0_u15_U67  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[28] ) );
INV_X4 _u0_u15_U65  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[27] ) );
INV_X4 _u0_u15_U63  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[26] ) );
INV_X4 _u0_u15_U61  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[25] ) );
INV_X4 _u0_u15_U59  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[24] ) );
INV_X4 _u0_u15_U57  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[23] ) );
INV_X4 _u0_u15_U55  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[22] ) );
INV_X4 _u0_u15_U53  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[21] ) );
INV_X4 _u0_u15_U51  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[20] ) );
INV_X4 _u0_u15_U49  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[19] ) );
INV_X4 _u0_u15_U47  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[18] ) );
INV_X4 _u0_u15_U45  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[17] ) );
INV_X4 _u0_u15_U43  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[16] ) );
INV_X4 _u0_u15_U41  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[15] ) );
INV_X4 _u0_u15_U39  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[14] ) );
INV_X4 _u0_u15_U37  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[13] ) );
INV_X4 _u0_u15_U35  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[12] ) );
INV_X4 _u0_u15_U33  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[11] ) );
INV_X4 _u0_u15_U31  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[10] ) );
INV_X4 _u0_u15_U29  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[9] ) );
INV_X4 _u0_u15_U27  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[8] ) );
INV_X4 _u0_u15_U25  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[7] ) );
INV_X4 _u0_u15_U23  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[6] ) );
INV_X4 _u0_u15_U21  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[5] ) );
INV_X4 _u0_u15_U19  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[4] ) );
INV_X4 _u0_u15_U17  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[3] ) );
INV_X4 _u0_u15_U15  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[2] ) );
INV_X4 _u0_u15_U13  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[1] ) );
INV_X4 _u0_u15_U11  ( .A(1'b1), .ZN(_u0_u15_sw_pointer[0] ) );
INV_X4 _u0_u15_U9  ( .A(1'b1), .ZN(_u0_u15_ch_stop ) );
INV_X4 _u0_u15_U7  ( .A(1'b1), .ZN(_u0_u15_ch_dis ) );
INV_X4 _u0_u15_U5  ( .A(1'b1), .ZN(_u0_u15_int ) );
INV_X4 _u0_u16_U585  ( .A(1'b1), .ZN(_u0_u16_pointer[31] ) );
INV_X4 _u0_u16_U583  ( .A(1'b1), .ZN(_u0_u16_pointer[30] ) );
INV_X4 _u0_u16_U581  ( .A(1'b1), .ZN(_u0_u16_pointer[29] ) );
INV_X4 _u0_u16_U579  ( .A(1'b1), .ZN(_u0_u16_pointer[28] ) );
INV_X4 _u0_u16_U577  ( .A(1'b1), .ZN(_u0_u16_pointer[27] ) );
INV_X4 _u0_u16_U575  ( .A(1'b1), .ZN(_u0_u16_pointer[26] ) );
INV_X4 _u0_u16_U573  ( .A(1'b1), .ZN(_u0_u16_pointer[25] ) );
INV_X4 _u0_u16_U571  ( .A(1'b1), .ZN(_u0_u16_pointer[24] ) );
INV_X4 _u0_u16_U569  ( .A(1'b1), .ZN(_u0_u16_pointer[23] ) );
INV_X4 _u0_u16_U567  ( .A(1'b1), .ZN(_u0_u16_pointer[22] ) );
INV_X4 _u0_u16_U565  ( .A(1'b1), .ZN(_u0_u16_pointer[21] ) );
INV_X4 _u0_u16_U563  ( .A(1'b1), .ZN(_u0_u16_pointer[20] ) );
INV_X4 _u0_u16_U561  ( .A(1'b1), .ZN(_u0_u16_pointer[19] ) );
INV_X4 _u0_u16_U559  ( .A(1'b1), .ZN(_u0_u16_pointer[18] ) );
INV_X4 _u0_u16_U557  ( .A(1'b1), .ZN(_u0_u16_pointer[17] ) );
INV_X4 _u0_u16_U555  ( .A(1'b1), .ZN(_u0_u16_pointer[16] ) );
INV_X4 _u0_u16_U553  ( .A(1'b1), .ZN(_u0_u16_pointer[15] ) );
INV_X4 _u0_u16_U551  ( .A(1'b1), .ZN(_u0_u16_pointer[14] ) );
INV_X4 _u0_u16_U549  ( .A(1'b1), .ZN(_u0_u16_pointer[13] ) );
INV_X4 _u0_u16_U547  ( .A(1'b1), .ZN(_u0_u16_pointer[12] ) );
INV_X4 _u0_u16_U545  ( .A(1'b1), .ZN(_u0_u16_pointer[11] ) );
INV_X4 _u0_u16_U543  ( .A(1'b1), .ZN(_u0_u16_pointer[10] ) );
INV_X4 _u0_u16_U541  ( .A(1'b1), .ZN(_u0_u16_pointer[9] ) );
INV_X4 _u0_u16_U539  ( .A(1'b1), .ZN(_u0_u16_pointer[8] ) );
INV_X4 _u0_u16_U537  ( .A(1'b1), .ZN(_u0_u16_pointer[7] ) );
INV_X4 _u0_u16_U535  ( .A(1'b1), .ZN(_u0_u16_pointer[6] ) );
INV_X4 _u0_u16_U533  ( .A(1'b1), .ZN(_u0_u16_pointer[5] ) );
INV_X4 _u0_u16_U531  ( .A(1'b1), .ZN(_u0_u16_pointer[4] ) );
INV_X4 _u0_u16_U529  ( .A(1'b1), .ZN(_u0_u16_pointer[3] ) );
INV_X4 _u0_u16_U527  ( .A(1'b1), .ZN(_u0_u16_pointer[2] ) );
INV_X4 _u0_u16_U525  ( .A(1'b1), .ZN(_u0_u16_pointer[1] ) );
INV_X4 _u0_u16_U523  ( .A(1'b1), .ZN(_u0_u16_pointer[0] ) );
INV_X4 _u0_u16_U521  ( .A(1'b1), .ZN(_u0_u16_pointer_s[31] ) );
INV_X4 _u0_u16_U519  ( .A(1'b1), .ZN(_u0_u16_pointer_s[30] ) );
INV_X4 _u0_u16_U517  ( .A(1'b1), .ZN(_u0_u16_pointer_s[29] ) );
INV_X4 _u0_u16_U515  ( .A(1'b1), .ZN(_u0_u16_pointer_s[28] ) );
INV_X4 _u0_u16_U513  ( .A(1'b1), .ZN(_u0_u16_pointer_s[27] ) );
INV_X4 _u0_u16_U511  ( .A(1'b1), .ZN(_u0_u16_pointer_s[26] ) );
INV_X4 _u0_u16_U509  ( .A(1'b1), .ZN(_u0_u16_pointer_s[25] ) );
INV_X4 _u0_u16_U507  ( .A(1'b1), .ZN(_u0_u16_pointer_s[24] ) );
INV_X4 _u0_u16_U505  ( .A(1'b1), .ZN(_u0_u16_pointer_s[23] ) );
INV_X4 _u0_u16_U503  ( .A(1'b1), .ZN(_u0_u16_pointer_s[22] ) );
INV_X4 _u0_u16_U501  ( .A(1'b1), .ZN(_u0_u16_pointer_s[21] ) );
INV_X4 _u0_u16_U499  ( .A(1'b1), .ZN(_u0_u16_pointer_s[20] ) );
INV_X4 _u0_u16_U497  ( .A(1'b1), .ZN(_u0_u16_pointer_s[19] ) );
INV_X4 _u0_u16_U495  ( .A(1'b1), .ZN(_u0_u16_pointer_s[18] ) );
INV_X4 _u0_u16_U493  ( .A(1'b1), .ZN(_u0_u16_pointer_s[17] ) );
INV_X4 _u0_u16_U491  ( .A(1'b1), .ZN(_u0_u16_pointer_s[16] ) );
INV_X4 _u0_u16_U489  ( .A(1'b1), .ZN(_u0_u16_pointer_s[15] ) );
INV_X4 _u0_u16_U487  ( .A(1'b1), .ZN(_u0_u16_pointer_s[14] ) );
INV_X4 _u0_u16_U485  ( .A(1'b1), .ZN(_u0_u16_pointer_s[13] ) );
INV_X4 _u0_u16_U483  ( .A(1'b1), .ZN(_u0_u16_pointer_s[12] ) );
INV_X4 _u0_u16_U481  ( .A(1'b1), .ZN(_u0_u16_pointer_s[11] ) );
INV_X4 _u0_u16_U479  ( .A(1'b1), .ZN(_u0_u16_pointer_s[10] ) );
INV_X4 _u0_u16_U477  ( .A(1'b1), .ZN(_u0_u16_pointer_s[9] ) );
INV_X4 _u0_u16_U475  ( .A(1'b1), .ZN(_u0_u16_pointer_s[8] ) );
INV_X4 _u0_u16_U473  ( .A(1'b1), .ZN(_u0_u16_pointer_s[7] ) );
INV_X4 _u0_u16_U471  ( .A(1'b1), .ZN(_u0_u16_pointer_s[6] ) );
INV_X4 _u0_u16_U469  ( .A(1'b1), .ZN(_u0_u16_pointer_s[5] ) );
INV_X4 _u0_u16_U467  ( .A(1'b1), .ZN(_u0_u16_pointer_s[4] ) );
INV_X4 _u0_u16_U465  ( .A(1'b1), .ZN(_u0_u16_pointer_s[3] ) );
INV_X4 _u0_u16_U463  ( .A(1'b1), .ZN(_u0_u16_pointer_s[2] ) );
INV_X4 _u0_u16_U461  ( .A(1'b1), .ZN(_u0_u16_pointer_s[1] ) );
INV_X4 _u0_u16_U459  ( .A(1'b1), .ZN(_u0_u16_pointer_s[0] ) );
INV_X4 _u0_u16_U457  ( .A(1'b1), .ZN(_u0_u16_ch_csr[31] ) );
INV_X4 _u0_u16_U455  ( .A(1'b1), .ZN(_u0_u16_ch_csr[30] ) );
INV_X4 _u0_u16_U453  ( .A(1'b1), .ZN(_u0_u16_ch_csr[29] ) );
INV_X4 _u0_u16_U451  ( .A(1'b1), .ZN(_u0_u16_ch_csr[28] ) );
INV_X4 _u0_u16_U449  ( .A(1'b1), .ZN(_u0_u16_ch_csr[27] ) );
INV_X4 _u0_u16_U447  ( .A(1'b1), .ZN(_u0_u16_ch_csr[26] ) );
INV_X4 _u0_u16_U445  ( .A(1'b1), .ZN(_u0_u16_ch_csr[25] ) );
INV_X4 _u0_u16_U443  ( .A(1'b1), .ZN(_u0_u16_ch_csr[24] ) );
INV_X4 _u0_u16_U441  ( .A(1'b1), .ZN(_u0_u16_ch_csr[23] ) );
INV_X4 _u0_u16_U439  ( .A(1'b1), .ZN(_u0_u16_ch_csr[22] ) );
INV_X4 _u0_u16_U437  ( .A(1'b1), .ZN(_u0_u16_ch_csr[21] ) );
INV_X4 _u0_u16_U435  ( .A(1'b1), .ZN(_u0_u16_ch_csr[20] ) );
INV_X4 _u0_u16_U433  ( .A(1'b1), .ZN(_u0_u16_ch_csr[19] ) );
INV_X4 _u0_u16_U431  ( .A(1'b1), .ZN(_u0_u16_ch_csr[18] ) );
INV_X4 _u0_u16_U429  ( .A(1'b1), .ZN(_u0_u16_ch_csr[17] ) );
INV_X4 _u0_u16_U427  ( .A(1'b1), .ZN(_u0_u16_ch_csr[16] ) );
INV_X4 _u0_u16_U425  ( .A(1'b1), .ZN(_u0_u16_ch_csr[15] ) );
INV_X4 _u0_u16_U423  ( .A(1'b1), .ZN(_u0_u16_ch_csr[14] ) );
INV_X4 _u0_u16_U421  ( .A(1'b1), .ZN(_u0_u16_ch_csr[13] ) );
INV_X4 _u0_u16_U419  ( .A(1'b1), .ZN(_u0_u16_ch_csr[12] ) );
INV_X4 _u0_u16_U417  ( .A(1'b1), .ZN(_u0_u16_ch_csr[11] ) );
INV_X4 _u0_u16_U415  ( .A(1'b1), .ZN(_u0_u16_ch_csr[10] ) );
INV_X4 _u0_u16_U413  ( .A(1'b1), .ZN(_u0_u16_ch_csr[9] ) );
INV_X4 _u0_u16_U411  ( .A(1'b1), .ZN(_u0_u16_ch_csr[8] ) );
INV_X4 _u0_u16_U409  ( .A(1'b1), .ZN(_u0_u16_ch_csr[7] ) );
INV_X4 _u0_u16_U407  ( .A(1'b1), .ZN(_u0_u16_ch_csr[6] ) );
INV_X4 _u0_u16_U405  ( .A(1'b1), .ZN(_u0_u16_ch_csr[5] ) );
INV_X4 _u0_u16_U403  ( .A(1'b1), .ZN(_u0_u16_ch_csr[4] ) );
INV_X4 _u0_u16_U401  ( .A(1'b1), .ZN(_u0_u16_ch_csr[3] ) );
INV_X4 _u0_u16_U399  ( .A(1'b1), .ZN(_u0_u16_ch_csr[2] ) );
INV_X4 _u0_u16_U397  ( .A(1'b1), .ZN(_u0_u16_ch_csr[1] ) );
INV_X4 _u0_u16_U395  ( .A(1'b1), .ZN(_u0_u16_ch_csr[0] ) );
INV_X4 _u0_u16_U393  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[31] ) );
INV_X4 _u0_u16_U391  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[30] ) );
INV_X4 _u0_u16_U389  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[29] ) );
INV_X4 _u0_u16_U387  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[28] ) );
INV_X4 _u0_u16_U385  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[27] ) );
INV_X4 _u0_u16_U383  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[26] ) );
INV_X4 _u0_u16_U381  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[25] ) );
INV_X4 _u0_u16_U379  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[24] ) );
INV_X4 _u0_u16_U377  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[23] ) );
INV_X4 _u0_u16_U375  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[22] ) );
INV_X4 _u0_u16_U373  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[21] ) );
INV_X4 _u0_u16_U371  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[20] ) );
INV_X4 _u0_u16_U369  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[19] ) );
INV_X4 _u0_u16_U367  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[18] ) );
INV_X4 _u0_u16_U365  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[17] ) );
INV_X4 _u0_u16_U363  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[16] ) );
INV_X4 _u0_u16_U361  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[15] ) );
INV_X4 _u0_u16_U359  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[14] ) );
INV_X4 _u0_u16_U357  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[13] ) );
INV_X4 _u0_u16_U355  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[12] ) );
INV_X4 _u0_u16_U353  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[11] ) );
INV_X4 _u0_u16_U351  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[10] ) );
INV_X4 _u0_u16_U349  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[9] ) );
INV_X4 _u0_u16_U347  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[8] ) );
INV_X4 _u0_u16_U345  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[7] ) );
INV_X4 _u0_u16_U343  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[6] ) );
INV_X4 _u0_u16_U341  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[5] ) );
INV_X4 _u0_u16_U339  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[4] ) );
INV_X4 _u0_u16_U337  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[3] ) );
INV_X4 _u0_u16_U335  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[2] ) );
INV_X4 _u0_u16_U333  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[1] ) );
INV_X4 _u0_u16_U331  ( .A(1'b1), .ZN(_u0_u16_ch_txsz[0] ) );
INV_X4 _u0_u16_U329  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[31] ) );
INV_X4 _u0_u16_U327  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[30] ) );
INV_X4 _u0_u16_U325  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[29] ) );
INV_X4 _u0_u16_U323  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[28] ) );
INV_X4 _u0_u16_U321  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[27] ) );
INV_X4 _u0_u16_U319  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[26] ) );
INV_X4 _u0_u16_U317  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[25] ) );
INV_X4 _u0_u16_U315  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[24] ) );
INV_X4 _u0_u16_U313  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[23] ) );
INV_X4 _u0_u16_U311  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[22] ) );
INV_X4 _u0_u16_U309  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[21] ) );
INV_X4 _u0_u16_U307  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[20] ) );
INV_X4 _u0_u16_U305  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[19] ) );
INV_X4 _u0_u16_U303  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[18] ) );
INV_X4 _u0_u16_U301  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[17] ) );
INV_X4 _u0_u16_U299  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[16] ) );
INV_X4 _u0_u16_U297  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[15] ) );
INV_X4 _u0_u16_U295  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[14] ) );
INV_X4 _u0_u16_U293  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[13] ) );
INV_X4 _u0_u16_U291  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[12] ) );
INV_X4 _u0_u16_U289  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[11] ) );
INV_X4 _u0_u16_U287  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[10] ) );
INV_X4 _u0_u16_U285  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[9] ) );
INV_X4 _u0_u16_U283  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[8] ) );
INV_X4 _u0_u16_U281  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[7] ) );
INV_X4 _u0_u16_U279  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[6] ) );
INV_X4 _u0_u16_U277  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[5] ) );
INV_X4 _u0_u16_U275  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[4] ) );
INV_X4 _u0_u16_U273  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[3] ) );
INV_X4 _u0_u16_U271  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[2] ) );
INV_X4 _u0_u16_U269  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[1] ) );
INV_X4 _u0_u16_U267  ( .A(1'b1), .ZN(_u0_u16_ch_adr0[0] ) );
INV_X4 _u0_u16_U265  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[31] ) );
INV_X4 _u0_u16_U263  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[30] ) );
INV_X4 _u0_u16_U261  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[29] ) );
INV_X4 _u0_u16_U259  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[28] ) );
INV_X4 _u0_u16_U257  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[27] ) );
INV_X4 _u0_u16_U255  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[26] ) );
INV_X4 _u0_u16_U253  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[25] ) );
INV_X4 _u0_u16_U251  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[24] ) );
INV_X4 _u0_u16_U249  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[23] ) );
INV_X4 _u0_u16_U247  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[22] ) );
INV_X4 _u0_u16_U245  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[21] ) );
INV_X4 _u0_u16_U243  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[20] ) );
INV_X4 _u0_u16_U241  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[19] ) );
INV_X4 _u0_u16_U239  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[18] ) );
INV_X4 _u0_u16_U237  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[17] ) );
INV_X4 _u0_u16_U235  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[16] ) );
INV_X4 _u0_u16_U233  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[15] ) );
INV_X4 _u0_u16_U231  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[14] ) );
INV_X4 _u0_u16_U229  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[13] ) );
INV_X4 _u0_u16_U227  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[12] ) );
INV_X4 _u0_u16_U225  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[11] ) );
INV_X4 _u0_u16_U223  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[10] ) );
INV_X4 _u0_u16_U221  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[9] ) );
INV_X4 _u0_u16_U219  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[8] ) );
INV_X4 _u0_u16_U217  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[7] ) );
INV_X4 _u0_u16_U215  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[6] ) );
INV_X4 _u0_u16_U213  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[5] ) );
INV_X4 _u0_u16_U211  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[4] ) );
INV_X4 _u0_u16_U209  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[3] ) );
INV_X4 _u0_u16_U207  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[2] ) );
INV_X4 _u0_u16_U205  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[1] ) );
INV_X4 _u0_u16_U203  ( .A(1'b1), .ZN(_u0_u16_ch_adr1[0] ) );
INV_X4 _u0_u16_U201  ( .A(1'b0), .ZN(_u0_u16_ch_am0[31] ) );
INV_X4 _u0_u16_U199  ( .A(1'b0), .ZN(_u0_u16_ch_am0[30] ) );
INV_X4 _u0_u16_U197  ( .A(1'b0), .ZN(_u0_u16_ch_am0[29] ) );
INV_X4 _u0_u16_U195  ( .A(1'b0), .ZN(_u0_u16_ch_am0[28] ) );
INV_X4 _u0_u16_U193  ( .A(1'b0), .ZN(_u0_u16_ch_am0[27] ) );
INV_X4 _u0_u16_U191  ( .A(1'b0), .ZN(_u0_u16_ch_am0[26] ) );
INV_X4 _u0_u16_U189  ( .A(1'b0), .ZN(_u0_u16_ch_am0[25] ) );
INV_X4 _u0_u16_U187  ( .A(1'b0), .ZN(_u0_u16_ch_am0[24] ) );
INV_X4 _u0_u16_U185  ( .A(1'b0), .ZN(_u0_u16_ch_am0[23] ) );
INV_X4 _u0_u16_U183  ( .A(1'b0), .ZN(_u0_u16_ch_am0[22] ) );
INV_X4 _u0_u16_U181  ( .A(1'b0), .ZN(_u0_u16_ch_am0[21] ) );
INV_X4 _u0_u16_U179  ( .A(1'b0), .ZN(_u0_u16_ch_am0[20] ) );
INV_X4 _u0_u16_U177  ( .A(1'b0), .ZN(_u0_u16_ch_am0[19] ) );
INV_X4 _u0_u16_U175  ( .A(1'b0), .ZN(_u0_u16_ch_am0[18] ) );
INV_X4 _u0_u16_U173  ( .A(1'b0), .ZN(_u0_u16_ch_am0[17] ) );
INV_X4 _u0_u16_U171  ( .A(1'b0), .ZN(_u0_u16_ch_am0[16] ) );
INV_X4 _u0_u16_U169  ( .A(1'b0), .ZN(_u0_u16_ch_am0[15] ) );
INV_X4 _u0_u16_U167  ( .A(1'b0), .ZN(_u0_u16_ch_am0[14] ) );
INV_X4 _u0_u16_U165  ( .A(1'b0), .ZN(_u0_u16_ch_am0[13] ) );
INV_X4 _u0_u16_U163  ( .A(1'b0), .ZN(_u0_u16_ch_am0[12] ) );
INV_X4 _u0_u16_U161  ( .A(1'b0), .ZN(_u0_u16_ch_am0[11] ) );
INV_X4 _u0_u16_U159  ( .A(1'b0), .ZN(_u0_u16_ch_am0[10] ) );
INV_X4 _u0_u16_U157  ( .A(1'b0), .ZN(_u0_u16_ch_am0[9] ) );
INV_X4 _u0_u16_U155  ( .A(1'b0), .ZN(_u0_u16_ch_am0[8] ) );
INV_X4 _u0_u16_U153  ( .A(1'b0), .ZN(_u0_u16_ch_am0[7] ) );
INV_X4 _u0_u16_U151  ( .A(1'b0), .ZN(_u0_u16_ch_am0[6] ) );
INV_X4 _u0_u16_U149  ( .A(1'b0), .ZN(_u0_u16_ch_am0[5] ) );
INV_X4 _u0_u16_U147  ( .A(1'b0), .ZN(_u0_u16_ch_am0[4] ) );
INV_X4 _u0_u16_U145  ( .A(1'b1), .ZN(_u0_u16_ch_am0[3] ) );
INV_X4 _u0_u16_U143  ( .A(1'b1), .ZN(_u0_u16_ch_am0[2] ) );
INV_X4 _u0_u16_U141  ( .A(1'b1), .ZN(_u0_u16_ch_am0[1] ) );
INV_X4 _u0_u16_U139  ( .A(1'b1), .ZN(_u0_u16_ch_am0[0] ) );
INV_X4 _u0_u16_U137  ( .A(1'b0), .ZN(_u0_u16_ch_am1[31] ) );
INV_X4 _u0_u16_U135  ( .A(1'b0), .ZN(_u0_u16_ch_am1[30] ) );
INV_X4 _u0_u16_U133  ( .A(1'b0), .ZN(_u0_u16_ch_am1[29] ) );
INV_X4 _u0_u16_U131  ( .A(1'b0), .ZN(_u0_u16_ch_am1[28] ) );
INV_X4 _u0_u16_U129  ( .A(1'b0), .ZN(_u0_u16_ch_am1[27] ) );
INV_X4 _u0_u16_U127  ( .A(1'b0), .ZN(_u0_u16_ch_am1[26] ) );
INV_X4 _u0_u16_U125  ( .A(1'b0), .ZN(_u0_u16_ch_am1[25] ) );
INV_X4 _u0_u16_U123  ( .A(1'b0), .ZN(_u0_u16_ch_am1[24] ) );
INV_X4 _u0_u16_U121  ( .A(1'b0), .ZN(_u0_u16_ch_am1[23] ) );
INV_X4 _u0_u16_U119  ( .A(1'b0), .ZN(_u0_u16_ch_am1[22] ) );
INV_X4 _u0_u16_U117  ( .A(1'b0), .ZN(_u0_u16_ch_am1[21] ) );
INV_X4 _u0_u16_U115  ( .A(1'b0), .ZN(_u0_u16_ch_am1[20] ) );
INV_X4 _u0_u16_U113  ( .A(1'b0), .ZN(_u0_u16_ch_am1[19] ) );
INV_X4 _u0_u16_U111  ( .A(1'b0), .ZN(_u0_u16_ch_am1[18] ) );
INV_X4 _u0_u16_U109  ( .A(1'b0), .ZN(_u0_u16_ch_am1[17] ) );
INV_X4 _u0_u16_U107  ( .A(1'b0), .ZN(_u0_u16_ch_am1[16] ) );
INV_X4 _u0_u16_U105  ( .A(1'b0), .ZN(_u0_u16_ch_am1[15] ) );
INV_X4 _u0_u16_U103  ( .A(1'b0), .ZN(_u0_u16_ch_am1[14] ) );
INV_X4 _u0_u16_U101  ( .A(1'b0), .ZN(_u0_u16_ch_am1[13] ) );
INV_X4 _u0_u16_U99  ( .A(1'b0), .ZN(_u0_u16_ch_am1[12] ) );
INV_X4 _u0_u16_U97  ( .A(1'b0), .ZN(_u0_u16_ch_am1[11] ) );
INV_X4 _u0_u16_U95  ( .A(1'b0), .ZN(_u0_u16_ch_am1[10] ) );
INV_X4 _u0_u16_U93  ( .A(1'b0), .ZN(_u0_u16_ch_am1[9] ) );
INV_X4 _u0_u16_U91  ( .A(1'b0), .ZN(_u0_u16_ch_am1[8] ) );
INV_X4 _u0_u16_U89  ( .A(1'b0), .ZN(_u0_u16_ch_am1[7] ) );
INV_X4 _u0_u16_U87  ( .A(1'b0), .ZN(_u0_u16_ch_am1[6] ) );
INV_X4 _u0_u16_U85  ( .A(1'b0), .ZN(_u0_u16_ch_am1[5] ) );
INV_X4 _u0_u16_U83  ( .A(1'b0), .ZN(_u0_u16_ch_am1[4] ) );
INV_X4 _u0_u16_U81  ( .A(1'b1), .ZN(_u0_u16_ch_am1[3] ) );
INV_X4 _u0_u16_U79  ( .A(1'b1), .ZN(_u0_u16_ch_am1[2] ) );
INV_X4 _u0_u16_U77  ( .A(1'b1), .ZN(_u0_u16_ch_am1[1] ) );
INV_X4 _u0_u16_U75  ( .A(1'b1), .ZN(_u0_u16_ch_am1[0] ) );
INV_X4 _u0_u16_U73  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[31] ) );
INV_X4 _u0_u16_U71  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[30] ) );
INV_X4 _u0_u16_U69  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[29] ) );
INV_X4 _u0_u16_U67  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[28] ) );
INV_X4 _u0_u16_U65  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[27] ) );
INV_X4 _u0_u16_U63  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[26] ) );
INV_X4 _u0_u16_U61  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[25] ) );
INV_X4 _u0_u16_U59  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[24] ) );
INV_X4 _u0_u16_U57  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[23] ) );
INV_X4 _u0_u16_U55  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[22] ) );
INV_X4 _u0_u16_U53  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[21] ) );
INV_X4 _u0_u16_U51  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[20] ) );
INV_X4 _u0_u16_U49  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[19] ) );
INV_X4 _u0_u16_U47  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[18] ) );
INV_X4 _u0_u16_U45  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[17] ) );
INV_X4 _u0_u16_U43  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[16] ) );
INV_X4 _u0_u16_U41  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[15] ) );
INV_X4 _u0_u16_U39  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[14] ) );
INV_X4 _u0_u16_U37  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[13] ) );
INV_X4 _u0_u16_U35  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[12] ) );
INV_X4 _u0_u16_U33  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[11] ) );
INV_X4 _u0_u16_U31  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[10] ) );
INV_X4 _u0_u16_U29  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[9] ) );
INV_X4 _u0_u16_U27  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[8] ) );
INV_X4 _u0_u16_U25  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[7] ) );
INV_X4 _u0_u16_U23  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[6] ) );
INV_X4 _u0_u16_U21  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[5] ) );
INV_X4 _u0_u16_U19  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[4] ) );
INV_X4 _u0_u16_U17  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[3] ) );
INV_X4 _u0_u16_U15  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[2] ) );
INV_X4 _u0_u16_U13  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[1] ) );
INV_X4 _u0_u16_U11  ( .A(1'b1), .ZN(_u0_u16_sw_pointer[0] ) );
INV_X4 _u0_u16_U9  ( .A(1'b1), .ZN(_u0_u16_ch_stop ) );
INV_X4 _u0_u16_U7  ( .A(1'b1), .ZN(_u0_u16_ch_dis ) );
INV_X4 _u0_u16_U5  ( .A(1'b1), .ZN(_u0_u16_int ) );
INV_X4 _u0_u17_U585  ( .A(1'b1), .ZN(_u0_u17_pointer[31] ) );
INV_X4 _u0_u17_U583  ( .A(1'b1), .ZN(_u0_u17_pointer[30] ) );
INV_X4 _u0_u17_U581  ( .A(1'b1), .ZN(_u0_u17_pointer[29] ) );
INV_X4 _u0_u17_U579  ( .A(1'b1), .ZN(_u0_u17_pointer[28] ) );
INV_X4 _u0_u17_U577  ( .A(1'b1), .ZN(_u0_u17_pointer[27] ) );
INV_X4 _u0_u17_U575  ( .A(1'b1), .ZN(_u0_u17_pointer[26] ) );
INV_X4 _u0_u17_U573  ( .A(1'b1), .ZN(_u0_u17_pointer[25] ) );
INV_X4 _u0_u17_U571  ( .A(1'b1), .ZN(_u0_u17_pointer[24] ) );
INV_X4 _u0_u17_U569  ( .A(1'b1), .ZN(_u0_u17_pointer[23] ) );
INV_X4 _u0_u17_U567  ( .A(1'b1), .ZN(_u0_u17_pointer[22] ) );
INV_X4 _u0_u17_U565  ( .A(1'b1), .ZN(_u0_u17_pointer[21] ) );
INV_X4 _u0_u17_U563  ( .A(1'b1), .ZN(_u0_u17_pointer[20] ) );
INV_X4 _u0_u17_U561  ( .A(1'b1), .ZN(_u0_u17_pointer[19] ) );
INV_X4 _u0_u17_U559  ( .A(1'b1), .ZN(_u0_u17_pointer[18] ) );
INV_X4 _u0_u17_U557  ( .A(1'b1), .ZN(_u0_u17_pointer[17] ) );
INV_X4 _u0_u17_U555  ( .A(1'b1), .ZN(_u0_u17_pointer[16] ) );
INV_X4 _u0_u17_U553  ( .A(1'b1), .ZN(_u0_u17_pointer[15] ) );
INV_X4 _u0_u17_U551  ( .A(1'b1), .ZN(_u0_u17_pointer[14] ) );
INV_X4 _u0_u17_U549  ( .A(1'b1), .ZN(_u0_u17_pointer[13] ) );
INV_X4 _u0_u17_U547  ( .A(1'b1), .ZN(_u0_u17_pointer[12] ) );
INV_X4 _u0_u17_U545  ( .A(1'b1), .ZN(_u0_u17_pointer[11] ) );
INV_X4 _u0_u17_U543  ( .A(1'b1), .ZN(_u0_u17_pointer[10] ) );
INV_X4 _u0_u17_U541  ( .A(1'b1), .ZN(_u0_u17_pointer[9] ) );
INV_X4 _u0_u17_U539  ( .A(1'b1), .ZN(_u0_u17_pointer[8] ) );
INV_X4 _u0_u17_U537  ( .A(1'b1), .ZN(_u0_u17_pointer[7] ) );
INV_X4 _u0_u17_U535  ( .A(1'b1), .ZN(_u0_u17_pointer[6] ) );
INV_X4 _u0_u17_U533  ( .A(1'b1), .ZN(_u0_u17_pointer[5] ) );
INV_X4 _u0_u17_U531  ( .A(1'b1), .ZN(_u0_u17_pointer[4] ) );
INV_X4 _u0_u17_U529  ( .A(1'b1), .ZN(_u0_u17_pointer[3] ) );
INV_X4 _u0_u17_U527  ( .A(1'b1), .ZN(_u0_u17_pointer[2] ) );
INV_X4 _u0_u17_U525  ( .A(1'b1), .ZN(_u0_u17_pointer[1] ) );
INV_X4 _u0_u17_U523  ( .A(1'b1), .ZN(_u0_u17_pointer[0] ) );
INV_X4 _u0_u17_U521  ( .A(1'b1), .ZN(_u0_u17_pointer_s[31] ) );
INV_X4 _u0_u17_U519  ( .A(1'b1), .ZN(_u0_u17_pointer_s[30] ) );
INV_X4 _u0_u17_U517  ( .A(1'b1), .ZN(_u0_u17_pointer_s[29] ) );
INV_X4 _u0_u17_U515  ( .A(1'b1), .ZN(_u0_u17_pointer_s[28] ) );
INV_X4 _u0_u17_U513  ( .A(1'b1), .ZN(_u0_u17_pointer_s[27] ) );
INV_X4 _u0_u17_U511  ( .A(1'b1), .ZN(_u0_u17_pointer_s[26] ) );
INV_X4 _u0_u17_U509  ( .A(1'b1), .ZN(_u0_u17_pointer_s[25] ) );
INV_X4 _u0_u17_U507  ( .A(1'b1), .ZN(_u0_u17_pointer_s[24] ) );
INV_X4 _u0_u17_U505  ( .A(1'b1), .ZN(_u0_u17_pointer_s[23] ) );
INV_X4 _u0_u17_U503  ( .A(1'b1), .ZN(_u0_u17_pointer_s[22] ) );
INV_X4 _u0_u17_U501  ( .A(1'b1), .ZN(_u0_u17_pointer_s[21] ) );
INV_X4 _u0_u17_U499  ( .A(1'b1), .ZN(_u0_u17_pointer_s[20] ) );
INV_X4 _u0_u17_U497  ( .A(1'b1), .ZN(_u0_u17_pointer_s[19] ) );
INV_X4 _u0_u17_U495  ( .A(1'b1), .ZN(_u0_u17_pointer_s[18] ) );
INV_X4 _u0_u17_U493  ( .A(1'b1), .ZN(_u0_u17_pointer_s[17] ) );
INV_X4 _u0_u17_U491  ( .A(1'b1), .ZN(_u0_u17_pointer_s[16] ) );
INV_X4 _u0_u17_U489  ( .A(1'b1), .ZN(_u0_u17_pointer_s[15] ) );
INV_X4 _u0_u17_U487  ( .A(1'b1), .ZN(_u0_u17_pointer_s[14] ) );
INV_X4 _u0_u17_U485  ( .A(1'b1), .ZN(_u0_u17_pointer_s[13] ) );
INV_X4 _u0_u17_U483  ( .A(1'b1), .ZN(_u0_u17_pointer_s[12] ) );
INV_X4 _u0_u17_U481  ( .A(1'b1), .ZN(_u0_u17_pointer_s[11] ) );
INV_X4 _u0_u17_U479  ( .A(1'b1), .ZN(_u0_u17_pointer_s[10] ) );
INV_X4 _u0_u17_U477  ( .A(1'b1), .ZN(_u0_u17_pointer_s[9] ) );
INV_X4 _u0_u17_U475  ( .A(1'b1), .ZN(_u0_u17_pointer_s[8] ) );
INV_X4 _u0_u17_U473  ( .A(1'b1), .ZN(_u0_u17_pointer_s[7] ) );
INV_X4 _u0_u17_U471  ( .A(1'b1), .ZN(_u0_u17_pointer_s[6] ) );
INV_X4 _u0_u17_U469  ( .A(1'b1), .ZN(_u0_u17_pointer_s[5] ) );
INV_X4 _u0_u17_U467  ( .A(1'b1), .ZN(_u0_u17_pointer_s[4] ) );
INV_X4 _u0_u17_U465  ( .A(1'b1), .ZN(_u0_u17_pointer_s[3] ) );
INV_X4 _u0_u17_U463  ( .A(1'b1), .ZN(_u0_u17_pointer_s[2] ) );
INV_X4 _u0_u17_U461  ( .A(1'b1), .ZN(_u0_u17_pointer_s[1] ) );
INV_X4 _u0_u17_U459  ( .A(1'b1), .ZN(_u0_u17_pointer_s[0] ) );
INV_X4 _u0_u17_U457  ( .A(1'b1), .ZN(_u0_u17_ch_csr[31] ) );
INV_X4 _u0_u17_U455  ( .A(1'b1), .ZN(_u0_u17_ch_csr[30] ) );
INV_X4 _u0_u17_U453  ( .A(1'b1), .ZN(_u0_u17_ch_csr[29] ) );
INV_X4 _u0_u17_U451  ( .A(1'b1), .ZN(_u0_u17_ch_csr[28] ) );
INV_X4 _u0_u17_U449  ( .A(1'b1), .ZN(_u0_u17_ch_csr[27] ) );
INV_X4 _u0_u17_U447  ( .A(1'b1), .ZN(_u0_u17_ch_csr[26] ) );
INV_X4 _u0_u17_U445  ( .A(1'b1), .ZN(_u0_u17_ch_csr[25] ) );
INV_X4 _u0_u17_U443  ( .A(1'b1), .ZN(_u0_u17_ch_csr[24] ) );
INV_X4 _u0_u17_U441  ( .A(1'b1), .ZN(_u0_u17_ch_csr[23] ) );
INV_X4 _u0_u17_U439  ( .A(1'b1), .ZN(_u0_u17_ch_csr[22] ) );
INV_X4 _u0_u17_U437  ( .A(1'b1), .ZN(_u0_u17_ch_csr[21] ) );
INV_X4 _u0_u17_U435  ( .A(1'b1), .ZN(_u0_u17_ch_csr[20] ) );
INV_X4 _u0_u17_U433  ( .A(1'b1), .ZN(_u0_u17_ch_csr[19] ) );
INV_X4 _u0_u17_U431  ( .A(1'b1), .ZN(_u0_u17_ch_csr[18] ) );
INV_X4 _u0_u17_U429  ( .A(1'b1), .ZN(_u0_u17_ch_csr[17] ) );
INV_X4 _u0_u17_U427  ( .A(1'b1), .ZN(_u0_u17_ch_csr[16] ) );
INV_X4 _u0_u17_U425  ( .A(1'b1), .ZN(_u0_u17_ch_csr[15] ) );
INV_X4 _u0_u17_U423  ( .A(1'b1), .ZN(_u0_u17_ch_csr[14] ) );
INV_X4 _u0_u17_U421  ( .A(1'b1), .ZN(_u0_u17_ch_csr[13] ) );
INV_X4 _u0_u17_U419  ( .A(1'b1), .ZN(_u0_u17_ch_csr[12] ) );
INV_X4 _u0_u17_U417  ( .A(1'b1), .ZN(_u0_u17_ch_csr[11] ) );
INV_X4 _u0_u17_U415  ( .A(1'b1), .ZN(_u0_u17_ch_csr[10] ) );
INV_X4 _u0_u17_U413  ( .A(1'b1), .ZN(_u0_u17_ch_csr[9] ) );
INV_X4 _u0_u17_U411  ( .A(1'b1), .ZN(_u0_u17_ch_csr[8] ) );
INV_X4 _u0_u17_U409  ( .A(1'b1), .ZN(_u0_u17_ch_csr[7] ) );
INV_X4 _u0_u17_U407  ( .A(1'b1), .ZN(_u0_u17_ch_csr[6] ) );
INV_X4 _u0_u17_U405  ( .A(1'b1), .ZN(_u0_u17_ch_csr[5] ) );
INV_X4 _u0_u17_U403  ( .A(1'b1), .ZN(_u0_u17_ch_csr[4] ) );
INV_X4 _u0_u17_U401  ( .A(1'b1), .ZN(_u0_u17_ch_csr[3] ) );
INV_X4 _u0_u17_U399  ( .A(1'b1), .ZN(_u0_u17_ch_csr[2] ) );
INV_X4 _u0_u17_U397  ( .A(1'b1), .ZN(_u0_u17_ch_csr[1] ) );
INV_X4 _u0_u17_U395  ( .A(1'b1), .ZN(_u0_u17_ch_csr[0] ) );
INV_X4 _u0_u17_U393  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[31] ) );
INV_X4 _u0_u17_U391  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[30] ) );
INV_X4 _u0_u17_U389  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[29] ) );
INV_X4 _u0_u17_U387  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[28] ) );
INV_X4 _u0_u17_U385  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[27] ) );
INV_X4 _u0_u17_U383  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[26] ) );
INV_X4 _u0_u17_U381  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[25] ) );
INV_X4 _u0_u17_U379  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[24] ) );
INV_X4 _u0_u17_U377  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[23] ) );
INV_X4 _u0_u17_U375  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[22] ) );
INV_X4 _u0_u17_U373  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[21] ) );
INV_X4 _u0_u17_U371  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[20] ) );
INV_X4 _u0_u17_U369  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[19] ) );
INV_X4 _u0_u17_U367  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[18] ) );
INV_X4 _u0_u17_U365  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[17] ) );
INV_X4 _u0_u17_U363  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[16] ) );
INV_X4 _u0_u17_U361  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[15] ) );
INV_X4 _u0_u17_U359  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[14] ) );
INV_X4 _u0_u17_U357  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[13] ) );
INV_X4 _u0_u17_U355  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[12] ) );
INV_X4 _u0_u17_U353  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[11] ) );
INV_X4 _u0_u17_U351  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[10] ) );
INV_X4 _u0_u17_U349  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[9] ) );
INV_X4 _u0_u17_U347  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[8] ) );
INV_X4 _u0_u17_U345  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[7] ) );
INV_X4 _u0_u17_U343  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[6] ) );
INV_X4 _u0_u17_U341  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[5] ) );
INV_X4 _u0_u17_U339  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[4] ) );
INV_X4 _u0_u17_U337  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[3] ) );
INV_X4 _u0_u17_U335  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[2] ) );
INV_X4 _u0_u17_U333  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[1] ) );
INV_X4 _u0_u17_U331  ( .A(1'b1), .ZN(_u0_u17_ch_txsz[0] ) );
INV_X4 _u0_u17_U329  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[31] ) );
INV_X4 _u0_u17_U327  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[30] ) );
INV_X4 _u0_u17_U325  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[29] ) );
INV_X4 _u0_u17_U323  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[28] ) );
INV_X4 _u0_u17_U321  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[27] ) );
INV_X4 _u0_u17_U319  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[26] ) );
INV_X4 _u0_u17_U317  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[25] ) );
INV_X4 _u0_u17_U315  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[24] ) );
INV_X4 _u0_u17_U313  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[23] ) );
INV_X4 _u0_u17_U311  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[22] ) );
INV_X4 _u0_u17_U309  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[21] ) );
INV_X4 _u0_u17_U307  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[20] ) );
INV_X4 _u0_u17_U305  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[19] ) );
INV_X4 _u0_u17_U303  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[18] ) );
INV_X4 _u0_u17_U301  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[17] ) );
INV_X4 _u0_u17_U299  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[16] ) );
INV_X4 _u0_u17_U297  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[15] ) );
INV_X4 _u0_u17_U295  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[14] ) );
INV_X4 _u0_u17_U293  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[13] ) );
INV_X4 _u0_u17_U291  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[12] ) );
INV_X4 _u0_u17_U289  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[11] ) );
INV_X4 _u0_u17_U287  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[10] ) );
INV_X4 _u0_u17_U285  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[9] ) );
INV_X4 _u0_u17_U283  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[8] ) );
INV_X4 _u0_u17_U281  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[7] ) );
INV_X4 _u0_u17_U279  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[6] ) );
INV_X4 _u0_u17_U277  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[5] ) );
INV_X4 _u0_u17_U275  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[4] ) );
INV_X4 _u0_u17_U273  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[3] ) );
INV_X4 _u0_u17_U271  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[2] ) );
INV_X4 _u0_u17_U269  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[1] ) );
INV_X4 _u0_u17_U267  ( .A(1'b1), .ZN(_u0_u17_ch_adr0[0] ) );
INV_X4 _u0_u17_U265  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[31] ) );
INV_X4 _u0_u17_U263  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[30] ) );
INV_X4 _u0_u17_U261  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[29] ) );
INV_X4 _u0_u17_U259  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[28] ) );
INV_X4 _u0_u17_U257  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[27] ) );
INV_X4 _u0_u17_U255  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[26] ) );
INV_X4 _u0_u17_U253  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[25] ) );
INV_X4 _u0_u17_U251  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[24] ) );
INV_X4 _u0_u17_U249  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[23] ) );
INV_X4 _u0_u17_U247  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[22] ) );
INV_X4 _u0_u17_U245  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[21] ) );
INV_X4 _u0_u17_U243  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[20] ) );
INV_X4 _u0_u17_U241  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[19] ) );
INV_X4 _u0_u17_U239  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[18] ) );
INV_X4 _u0_u17_U237  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[17] ) );
INV_X4 _u0_u17_U235  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[16] ) );
INV_X4 _u0_u17_U233  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[15] ) );
INV_X4 _u0_u17_U231  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[14] ) );
INV_X4 _u0_u17_U229  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[13] ) );
INV_X4 _u0_u17_U227  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[12] ) );
INV_X4 _u0_u17_U225  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[11] ) );
INV_X4 _u0_u17_U223  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[10] ) );
INV_X4 _u0_u17_U221  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[9] ) );
INV_X4 _u0_u17_U219  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[8] ) );
INV_X4 _u0_u17_U217  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[7] ) );
INV_X4 _u0_u17_U215  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[6] ) );
INV_X4 _u0_u17_U213  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[5] ) );
INV_X4 _u0_u17_U211  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[4] ) );
INV_X4 _u0_u17_U209  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[3] ) );
INV_X4 _u0_u17_U207  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[2] ) );
INV_X4 _u0_u17_U205  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[1] ) );
INV_X4 _u0_u17_U203  ( .A(1'b1), .ZN(_u0_u17_ch_adr1[0] ) );
INV_X4 _u0_u17_U201  ( .A(1'b0), .ZN(_u0_u17_ch_am0[31] ) );
INV_X4 _u0_u17_U199  ( .A(1'b0), .ZN(_u0_u17_ch_am0[30] ) );
INV_X4 _u0_u17_U197  ( .A(1'b0), .ZN(_u0_u17_ch_am0[29] ) );
INV_X4 _u0_u17_U195  ( .A(1'b0), .ZN(_u0_u17_ch_am0[28] ) );
INV_X4 _u0_u17_U193  ( .A(1'b0), .ZN(_u0_u17_ch_am0[27] ) );
INV_X4 _u0_u17_U191  ( .A(1'b0), .ZN(_u0_u17_ch_am0[26] ) );
INV_X4 _u0_u17_U189  ( .A(1'b0), .ZN(_u0_u17_ch_am0[25] ) );
INV_X4 _u0_u17_U187  ( .A(1'b0), .ZN(_u0_u17_ch_am0[24] ) );
INV_X4 _u0_u17_U185  ( .A(1'b0), .ZN(_u0_u17_ch_am0[23] ) );
INV_X4 _u0_u17_U183  ( .A(1'b0), .ZN(_u0_u17_ch_am0[22] ) );
INV_X4 _u0_u17_U181  ( .A(1'b0), .ZN(_u0_u17_ch_am0[21] ) );
INV_X4 _u0_u17_U179  ( .A(1'b0), .ZN(_u0_u17_ch_am0[20] ) );
INV_X4 _u0_u17_U177  ( .A(1'b0), .ZN(_u0_u17_ch_am0[19] ) );
INV_X4 _u0_u17_U175  ( .A(1'b0), .ZN(_u0_u17_ch_am0[18] ) );
INV_X4 _u0_u17_U173  ( .A(1'b0), .ZN(_u0_u17_ch_am0[17] ) );
INV_X4 _u0_u17_U171  ( .A(1'b0), .ZN(_u0_u17_ch_am0[16] ) );
INV_X4 _u0_u17_U169  ( .A(1'b0), .ZN(_u0_u17_ch_am0[15] ) );
INV_X4 _u0_u17_U167  ( .A(1'b0), .ZN(_u0_u17_ch_am0[14] ) );
INV_X4 _u0_u17_U165  ( .A(1'b0), .ZN(_u0_u17_ch_am0[13] ) );
INV_X4 _u0_u17_U163  ( .A(1'b0), .ZN(_u0_u17_ch_am0[12] ) );
INV_X4 _u0_u17_U161  ( .A(1'b0), .ZN(_u0_u17_ch_am0[11] ) );
INV_X4 _u0_u17_U159  ( .A(1'b0), .ZN(_u0_u17_ch_am0[10] ) );
INV_X4 _u0_u17_U157  ( .A(1'b0), .ZN(_u0_u17_ch_am0[9] ) );
INV_X4 _u0_u17_U155  ( .A(1'b0), .ZN(_u0_u17_ch_am0[8] ) );
INV_X4 _u0_u17_U153  ( .A(1'b0), .ZN(_u0_u17_ch_am0[7] ) );
INV_X4 _u0_u17_U151  ( .A(1'b0), .ZN(_u0_u17_ch_am0[6] ) );
INV_X4 _u0_u17_U149  ( .A(1'b0), .ZN(_u0_u17_ch_am0[5] ) );
INV_X4 _u0_u17_U147  ( .A(1'b0), .ZN(_u0_u17_ch_am0[4] ) );
INV_X4 _u0_u17_U145  ( .A(1'b1), .ZN(_u0_u17_ch_am0[3] ) );
INV_X4 _u0_u17_U143  ( .A(1'b1), .ZN(_u0_u17_ch_am0[2] ) );
INV_X4 _u0_u17_U141  ( .A(1'b1), .ZN(_u0_u17_ch_am0[1] ) );
INV_X4 _u0_u17_U139  ( .A(1'b1), .ZN(_u0_u17_ch_am0[0] ) );
INV_X4 _u0_u17_U137  ( .A(1'b0), .ZN(_u0_u17_ch_am1[31] ) );
INV_X4 _u0_u17_U135  ( .A(1'b0), .ZN(_u0_u17_ch_am1[30] ) );
INV_X4 _u0_u17_U133  ( .A(1'b0), .ZN(_u0_u17_ch_am1[29] ) );
INV_X4 _u0_u17_U131  ( .A(1'b0), .ZN(_u0_u17_ch_am1[28] ) );
INV_X4 _u0_u17_U129  ( .A(1'b0), .ZN(_u0_u17_ch_am1[27] ) );
INV_X4 _u0_u17_U127  ( .A(1'b0), .ZN(_u0_u17_ch_am1[26] ) );
INV_X4 _u0_u17_U125  ( .A(1'b0), .ZN(_u0_u17_ch_am1[25] ) );
INV_X4 _u0_u17_U123  ( .A(1'b0), .ZN(_u0_u17_ch_am1[24] ) );
INV_X4 _u0_u17_U121  ( .A(1'b0), .ZN(_u0_u17_ch_am1[23] ) );
INV_X4 _u0_u17_U119  ( .A(1'b0), .ZN(_u0_u17_ch_am1[22] ) );
INV_X4 _u0_u17_U117  ( .A(1'b0), .ZN(_u0_u17_ch_am1[21] ) );
INV_X4 _u0_u17_U115  ( .A(1'b0), .ZN(_u0_u17_ch_am1[20] ) );
INV_X4 _u0_u17_U113  ( .A(1'b0), .ZN(_u0_u17_ch_am1[19] ) );
INV_X4 _u0_u17_U111  ( .A(1'b0), .ZN(_u0_u17_ch_am1[18] ) );
INV_X4 _u0_u17_U109  ( .A(1'b0), .ZN(_u0_u17_ch_am1[17] ) );
INV_X4 _u0_u17_U107  ( .A(1'b0), .ZN(_u0_u17_ch_am1[16] ) );
INV_X4 _u0_u17_U105  ( .A(1'b0), .ZN(_u0_u17_ch_am1[15] ) );
INV_X4 _u0_u17_U103  ( .A(1'b0), .ZN(_u0_u17_ch_am1[14] ) );
INV_X4 _u0_u17_U101  ( .A(1'b0), .ZN(_u0_u17_ch_am1[13] ) );
INV_X4 _u0_u17_U99  ( .A(1'b0), .ZN(_u0_u17_ch_am1[12] ) );
INV_X4 _u0_u17_U97  ( .A(1'b0), .ZN(_u0_u17_ch_am1[11] ) );
INV_X4 _u0_u17_U95  ( .A(1'b0), .ZN(_u0_u17_ch_am1[10] ) );
INV_X4 _u0_u17_U93  ( .A(1'b0), .ZN(_u0_u17_ch_am1[9] ) );
INV_X4 _u0_u17_U91  ( .A(1'b0), .ZN(_u0_u17_ch_am1[8] ) );
INV_X4 _u0_u17_U89  ( .A(1'b0), .ZN(_u0_u17_ch_am1[7] ) );
INV_X4 _u0_u17_U87  ( .A(1'b0), .ZN(_u0_u17_ch_am1[6] ) );
INV_X4 _u0_u17_U85  ( .A(1'b0), .ZN(_u0_u17_ch_am1[5] ) );
INV_X4 _u0_u17_U83  ( .A(1'b0), .ZN(_u0_u17_ch_am1[4] ) );
INV_X4 _u0_u17_U81  ( .A(1'b1), .ZN(_u0_u17_ch_am1[3] ) );
INV_X4 _u0_u17_U79  ( .A(1'b1), .ZN(_u0_u17_ch_am1[2] ) );
INV_X4 _u0_u17_U77  ( .A(1'b1), .ZN(_u0_u17_ch_am1[1] ) );
INV_X4 _u0_u17_U75  ( .A(1'b1), .ZN(_u0_u17_ch_am1[0] ) );
INV_X4 _u0_u17_U73  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[31] ) );
INV_X4 _u0_u17_U71  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[30] ) );
INV_X4 _u0_u17_U69  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[29] ) );
INV_X4 _u0_u17_U67  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[28] ) );
INV_X4 _u0_u17_U65  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[27] ) );
INV_X4 _u0_u17_U63  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[26] ) );
INV_X4 _u0_u17_U61  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[25] ) );
INV_X4 _u0_u17_U59  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[24] ) );
INV_X4 _u0_u17_U57  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[23] ) );
INV_X4 _u0_u17_U55  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[22] ) );
INV_X4 _u0_u17_U53  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[21] ) );
INV_X4 _u0_u17_U51  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[20] ) );
INV_X4 _u0_u17_U49  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[19] ) );
INV_X4 _u0_u17_U47  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[18] ) );
INV_X4 _u0_u17_U45  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[17] ) );
INV_X4 _u0_u17_U43  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[16] ) );
INV_X4 _u0_u17_U41  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[15] ) );
INV_X4 _u0_u17_U39  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[14] ) );
INV_X4 _u0_u17_U37  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[13] ) );
INV_X4 _u0_u17_U35  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[12] ) );
INV_X4 _u0_u17_U33  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[11] ) );
INV_X4 _u0_u17_U31  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[10] ) );
INV_X4 _u0_u17_U29  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[9] ) );
INV_X4 _u0_u17_U27  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[8] ) );
INV_X4 _u0_u17_U25  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[7] ) );
INV_X4 _u0_u17_U23  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[6] ) );
INV_X4 _u0_u17_U21  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[5] ) );
INV_X4 _u0_u17_U19  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[4] ) );
INV_X4 _u0_u17_U17  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[3] ) );
INV_X4 _u0_u17_U15  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[2] ) );
INV_X4 _u0_u17_U13  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[1] ) );
INV_X4 _u0_u17_U11  ( .A(1'b1), .ZN(_u0_u17_sw_pointer[0] ) );
INV_X4 _u0_u17_U9  ( .A(1'b1), .ZN(_u0_u17_ch_stop ) );
INV_X4 _u0_u17_U7  ( .A(1'b1), .ZN(_u0_u17_ch_dis ) );
INV_X4 _u0_u17_U5  ( .A(1'b1), .ZN(_u0_u17_int ) );
INV_X4 _u0_u18_U585  ( .A(1'b1), .ZN(_u0_u18_pointer[31] ) );
INV_X4 _u0_u18_U583  ( .A(1'b1), .ZN(_u0_u18_pointer[30] ) );
INV_X4 _u0_u18_U581  ( .A(1'b1), .ZN(_u0_u18_pointer[29] ) );
INV_X4 _u0_u18_U579  ( .A(1'b1), .ZN(_u0_u18_pointer[28] ) );
INV_X4 _u0_u18_U577  ( .A(1'b1), .ZN(_u0_u18_pointer[27] ) );
INV_X4 _u0_u18_U575  ( .A(1'b1), .ZN(_u0_u18_pointer[26] ) );
INV_X4 _u0_u18_U573  ( .A(1'b1), .ZN(_u0_u18_pointer[25] ) );
INV_X4 _u0_u18_U571  ( .A(1'b1), .ZN(_u0_u18_pointer[24] ) );
INV_X4 _u0_u18_U569  ( .A(1'b1), .ZN(_u0_u18_pointer[23] ) );
INV_X4 _u0_u18_U567  ( .A(1'b1), .ZN(_u0_u18_pointer[22] ) );
INV_X4 _u0_u18_U565  ( .A(1'b1), .ZN(_u0_u18_pointer[21] ) );
INV_X4 _u0_u18_U563  ( .A(1'b1), .ZN(_u0_u18_pointer[20] ) );
INV_X4 _u0_u18_U561  ( .A(1'b1), .ZN(_u0_u18_pointer[19] ) );
INV_X4 _u0_u18_U559  ( .A(1'b1), .ZN(_u0_u18_pointer[18] ) );
INV_X4 _u0_u18_U557  ( .A(1'b1), .ZN(_u0_u18_pointer[17] ) );
INV_X4 _u0_u18_U555  ( .A(1'b1), .ZN(_u0_u18_pointer[16] ) );
INV_X4 _u0_u18_U553  ( .A(1'b1), .ZN(_u0_u18_pointer[15] ) );
INV_X4 _u0_u18_U551  ( .A(1'b1), .ZN(_u0_u18_pointer[14] ) );
INV_X4 _u0_u18_U549  ( .A(1'b1), .ZN(_u0_u18_pointer[13] ) );
INV_X4 _u0_u18_U547  ( .A(1'b1), .ZN(_u0_u18_pointer[12] ) );
INV_X4 _u0_u18_U545  ( .A(1'b1), .ZN(_u0_u18_pointer[11] ) );
INV_X4 _u0_u18_U543  ( .A(1'b1), .ZN(_u0_u18_pointer[10] ) );
INV_X4 _u0_u18_U541  ( .A(1'b1), .ZN(_u0_u18_pointer[9] ) );
INV_X4 _u0_u18_U539  ( .A(1'b1), .ZN(_u0_u18_pointer[8] ) );
INV_X4 _u0_u18_U537  ( .A(1'b1), .ZN(_u0_u18_pointer[7] ) );
INV_X4 _u0_u18_U535  ( .A(1'b1), .ZN(_u0_u18_pointer[6] ) );
INV_X4 _u0_u18_U533  ( .A(1'b1), .ZN(_u0_u18_pointer[5] ) );
INV_X4 _u0_u18_U531  ( .A(1'b1), .ZN(_u0_u18_pointer[4] ) );
INV_X4 _u0_u18_U529  ( .A(1'b1), .ZN(_u0_u18_pointer[3] ) );
INV_X4 _u0_u18_U527  ( .A(1'b1), .ZN(_u0_u18_pointer[2] ) );
INV_X4 _u0_u18_U525  ( .A(1'b1), .ZN(_u0_u18_pointer[1] ) );
INV_X4 _u0_u18_U523  ( .A(1'b1), .ZN(_u0_u18_pointer[0] ) );
INV_X4 _u0_u18_U521  ( .A(1'b1), .ZN(_u0_u18_pointer_s[31] ) );
INV_X4 _u0_u18_U519  ( .A(1'b1), .ZN(_u0_u18_pointer_s[30] ) );
INV_X4 _u0_u18_U517  ( .A(1'b1), .ZN(_u0_u18_pointer_s[29] ) );
INV_X4 _u0_u18_U515  ( .A(1'b1), .ZN(_u0_u18_pointer_s[28] ) );
INV_X4 _u0_u18_U513  ( .A(1'b1), .ZN(_u0_u18_pointer_s[27] ) );
INV_X4 _u0_u18_U511  ( .A(1'b1), .ZN(_u0_u18_pointer_s[26] ) );
INV_X4 _u0_u18_U509  ( .A(1'b1), .ZN(_u0_u18_pointer_s[25] ) );
INV_X4 _u0_u18_U507  ( .A(1'b1), .ZN(_u0_u18_pointer_s[24] ) );
INV_X4 _u0_u18_U505  ( .A(1'b1), .ZN(_u0_u18_pointer_s[23] ) );
INV_X4 _u0_u18_U503  ( .A(1'b1), .ZN(_u0_u18_pointer_s[22] ) );
INV_X4 _u0_u18_U501  ( .A(1'b1), .ZN(_u0_u18_pointer_s[21] ) );
INV_X4 _u0_u18_U499  ( .A(1'b1), .ZN(_u0_u18_pointer_s[20] ) );
INV_X4 _u0_u18_U497  ( .A(1'b1), .ZN(_u0_u18_pointer_s[19] ) );
INV_X4 _u0_u18_U495  ( .A(1'b1), .ZN(_u0_u18_pointer_s[18] ) );
INV_X4 _u0_u18_U493  ( .A(1'b1), .ZN(_u0_u18_pointer_s[17] ) );
INV_X4 _u0_u18_U491  ( .A(1'b1), .ZN(_u0_u18_pointer_s[16] ) );
INV_X4 _u0_u18_U489  ( .A(1'b1), .ZN(_u0_u18_pointer_s[15] ) );
INV_X4 _u0_u18_U487  ( .A(1'b1), .ZN(_u0_u18_pointer_s[14] ) );
INV_X4 _u0_u18_U485  ( .A(1'b1), .ZN(_u0_u18_pointer_s[13] ) );
INV_X4 _u0_u18_U483  ( .A(1'b1), .ZN(_u0_u18_pointer_s[12] ) );
INV_X4 _u0_u18_U481  ( .A(1'b1), .ZN(_u0_u18_pointer_s[11] ) );
INV_X4 _u0_u18_U479  ( .A(1'b1), .ZN(_u0_u18_pointer_s[10] ) );
INV_X4 _u0_u18_U477  ( .A(1'b1), .ZN(_u0_u18_pointer_s[9] ) );
INV_X4 _u0_u18_U475  ( .A(1'b1), .ZN(_u0_u18_pointer_s[8] ) );
INV_X4 _u0_u18_U473  ( .A(1'b1), .ZN(_u0_u18_pointer_s[7] ) );
INV_X4 _u0_u18_U471  ( .A(1'b1), .ZN(_u0_u18_pointer_s[6] ) );
INV_X4 _u0_u18_U469  ( .A(1'b1), .ZN(_u0_u18_pointer_s[5] ) );
INV_X4 _u0_u18_U467  ( .A(1'b1), .ZN(_u0_u18_pointer_s[4] ) );
INV_X4 _u0_u18_U465  ( .A(1'b1), .ZN(_u0_u18_pointer_s[3] ) );
INV_X4 _u0_u18_U463  ( .A(1'b1), .ZN(_u0_u18_pointer_s[2] ) );
INV_X4 _u0_u18_U461  ( .A(1'b1), .ZN(_u0_u18_pointer_s[1] ) );
INV_X4 _u0_u18_U459  ( .A(1'b1), .ZN(_u0_u18_pointer_s[0] ) );
INV_X4 _u0_u18_U457  ( .A(1'b1), .ZN(_u0_u18_ch_csr[31] ) );
INV_X4 _u0_u18_U455  ( .A(1'b1), .ZN(_u0_u18_ch_csr[30] ) );
INV_X4 _u0_u18_U453  ( .A(1'b1), .ZN(_u0_u18_ch_csr[29] ) );
INV_X4 _u0_u18_U451  ( .A(1'b1), .ZN(_u0_u18_ch_csr[28] ) );
INV_X4 _u0_u18_U449  ( .A(1'b1), .ZN(_u0_u18_ch_csr[27] ) );
INV_X4 _u0_u18_U447  ( .A(1'b1), .ZN(_u0_u18_ch_csr[26] ) );
INV_X4 _u0_u18_U445  ( .A(1'b1), .ZN(_u0_u18_ch_csr[25] ) );
INV_X4 _u0_u18_U443  ( .A(1'b1), .ZN(_u0_u18_ch_csr[24] ) );
INV_X4 _u0_u18_U441  ( .A(1'b1), .ZN(_u0_u18_ch_csr[23] ) );
INV_X4 _u0_u18_U439  ( .A(1'b1), .ZN(_u0_u18_ch_csr[22] ) );
INV_X4 _u0_u18_U437  ( .A(1'b1), .ZN(_u0_u18_ch_csr[21] ) );
INV_X4 _u0_u18_U435  ( .A(1'b1), .ZN(_u0_u18_ch_csr[20] ) );
INV_X4 _u0_u18_U433  ( .A(1'b1), .ZN(_u0_u18_ch_csr[19] ) );
INV_X4 _u0_u18_U431  ( .A(1'b1), .ZN(_u0_u18_ch_csr[18] ) );
INV_X4 _u0_u18_U429  ( .A(1'b1), .ZN(_u0_u18_ch_csr[17] ) );
INV_X4 _u0_u18_U427  ( .A(1'b1), .ZN(_u0_u18_ch_csr[16] ) );
INV_X4 _u0_u18_U425  ( .A(1'b1), .ZN(_u0_u18_ch_csr[15] ) );
INV_X4 _u0_u18_U423  ( .A(1'b1), .ZN(_u0_u18_ch_csr[14] ) );
INV_X4 _u0_u18_U421  ( .A(1'b1), .ZN(_u0_u18_ch_csr[13] ) );
INV_X4 _u0_u18_U419  ( .A(1'b1), .ZN(_u0_u18_ch_csr[12] ) );
INV_X4 _u0_u18_U417  ( .A(1'b1), .ZN(_u0_u18_ch_csr[11] ) );
INV_X4 _u0_u18_U415  ( .A(1'b1), .ZN(_u0_u18_ch_csr[10] ) );
INV_X4 _u0_u18_U413  ( .A(1'b1), .ZN(_u0_u18_ch_csr[9] ) );
INV_X4 _u0_u18_U411  ( .A(1'b1), .ZN(_u0_u18_ch_csr[8] ) );
INV_X4 _u0_u18_U409  ( .A(1'b1), .ZN(_u0_u18_ch_csr[7] ) );
INV_X4 _u0_u18_U407  ( .A(1'b1), .ZN(_u0_u18_ch_csr[6] ) );
INV_X4 _u0_u18_U405  ( .A(1'b1), .ZN(_u0_u18_ch_csr[5] ) );
INV_X4 _u0_u18_U403  ( .A(1'b1), .ZN(_u0_u18_ch_csr[4] ) );
INV_X4 _u0_u18_U401  ( .A(1'b1), .ZN(_u0_u18_ch_csr[3] ) );
INV_X4 _u0_u18_U399  ( .A(1'b1), .ZN(_u0_u18_ch_csr[2] ) );
INV_X4 _u0_u18_U397  ( .A(1'b1), .ZN(_u0_u18_ch_csr[1] ) );
INV_X4 _u0_u18_U395  ( .A(1'b1), .ZN(_u0_u18_ch_csr[0] ) );
INV_X4 _u0_u18_U393  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[31] ) );
INV_X4 _u0_u18_U391  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[30] ) );
INV_X4 _u0_u18_U389  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[29] ) );
INV_X4 _u0_u18_U387  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[28] ) );
INV_X4 _u0_u18_U385  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[27] ) );
INV_X4 _u0_u18_U383  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[26] ) );
INV_X4 _u0_u18_U381  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[25] ) );
INV_X4 _u0_u18_U379  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[24] ) );
INV_X4 _u0_u18_U377  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[23] ) );
INV_X4 _u0_u18_U375  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[22] ) );
INV_X4 _u0_u18_U373  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[21] ) );
INV_X4 _u0_u18_U371  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[20] ) );
INV_X4 _u0_u18_U369  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[19] ) );
INV_X4 _u0_u18_U367  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[18] ) );
INV_X4 _u0_u18_U365  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[17] ) );
INV_X4 _u0_u18_U363  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[16] ) );
INV_X4 _u0_u18_U361  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[15] ) );
INV_X4 _u0_u18_U359  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[14] ) );
INV_X4 _u0_u18_U357  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[13] ) );
INV_X4 _u0_u18_U355  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[12] ) );
INV_X4 _u0_u18_U353  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[11] ) );
INV_X4 _u0_u18_U351  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[10] ) );
INV_X4 _u0_u18_U349  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[9] ) );
INV_X4 _u0_u18_U347  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[8] ) );
INV_X4 _u0_u18_U345  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[7] ) );
INV_X4 _u0_u18_U343  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[6] ) );
INV_X4 _u0_u18_U341  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[5] ) );
INV_X4 _u0_u18_U339  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[4] ) );
INV_X4 _u0_u18_U337  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[3] ) );
INV_X4 _u0_u18_U335  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[2] ) );
INV_X4 _u0_u18_U333  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[1] ) );
INV_X4 _u0_u18_U331  ( .A(1'b1), .ZN(_u0_u18_ch_txsz[0] ) );
INV_X4 _u0_u18_U329  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[31] ) );
INV_X4 _u0_u18_U327  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[30] ) );
INV_X4 _u0_u18_U325  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[29] ) );
INV_X4 _u0_u18_U323  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[28] ) );
INV_X4 _u0_u18_U321  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[27] ) );
INV_X4 _u0_u18_U319  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[26] ) );
INV_X4 _u0_u18_U317  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[25] ) );
INV_X4 _u0_u18_U315  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[24] ) );
INV_X4 _u0_u18_U313  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[23] ) );
INV_X4 _u0_u18_U311  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[22] ) );
INV_X4 _u0_u18_U309  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[21] ) );
INV_X4 _u0_u18_U307  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[20] ) );
INV_X4 _u0_u18_U305  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[19] ) );
INV_X4 _u0_u18_U303  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[18] ) );
INV_X4 _u0_u18_U301  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[17] ) );
INV_X4 _u0_u18_U299  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[16] ) );
INV_X4 _u0_u18_U297  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[15] ) );
INV_X4 _u0_u18_U295  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[14] ) );
INV_X4 _u0_u18_U293  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[13] ) );
INV_X4 _u0_u18_U291  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[12] ) );
INV_X4 _u0_u18_U289  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[11] ) );
INV_X4 _u0_u18_U287  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[10] ) );
INV_X4 _u0_u18_U285  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[9] ) );
INV_X4 _u0_u18_U283  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[8] ) );
INV_X4 _u0_u18_U281  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[7] ) );
INV_X4 _u0_u18_U279  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[6] ) );
INV_X4 _u0_u18_U277  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[5] ) );
INV_X4 _u0_u18_U275  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[4] ) );
INV_X4 _u0_u18_U273  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[3] ) );
INV_X4 _u0_u18_U271  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[2] ) );
INV_X4 _u0_u18_U269  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[1] ) );
INV_X4 _u0_u18_U267  ( .A(1'b1), .ZN(_u0_u18_ch_adr0[0] ) );
INV_X4 _u0_u18_U265  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[31] ) );
INV_X4 _u0_u18_U263  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[30] ) );
INV_X4 _u0_u18_U261  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[29] ) );
INV_X4 _u0_u18_U259  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[28] ) );
INV_X4 _u0_u18_U257  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[27] ) );
INV_X4 _u0_u18_U255  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[26] ) );
INV_X4 _u0_u18_U253  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[25] ) );
INV_X4 _u0_u18_U251  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[24] ) );
INV_X4 _u0_u18_U249  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[23] ) );
INV_X4 _u0_u18_U247  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[22] ) );
INV_X4 _u0_u18_U245  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[21] ) );
INV_X4 _u0_u18_U243  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[20] ) );
INV_X4 _u0_u18_U241  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[19] ) );
INV_X4 _u0_u18_U239  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[18] ) );
INV_X4 _u0_u18_U237  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[17] ) );
INV_X4 _u0_u18_U235  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[16] ) );
INV_X4 _u0_u18_U233  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[15] ) );
INV_X4 _u0_u18_U231  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[14] ) );
INV_X4 _u0_u18_U229  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[13] ) );
INV_X4 _u0_u18_U227  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[12] ) );
INV_X4 _u0_u18_U225  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[11] ) );
INV_X4 _u0_u18_U223  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[10] ) );
INV_X4 _u0_u18_U221  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[9] ) );
INV_X4 _u0_u18_U219  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[8] ) );
INV_X4 _u0_u18_U217  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[7] ) );
INV_X4 _u0_u18_U215  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[6] ) );
INV_X4 _u0_u18_U213  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[5] ) );
INV_X4 _u0_u18_U211  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[4] ) );
INV_X4 _u0_u18_U209  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[3] ) );
INV_X4 _u0_u18_U207  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[2] ) );
INV_X4 _u0_u18_U205  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[1] ) );
INV_X4 _u0_u18_U203  ( .A(1'b1), .ZN(_u0_u18_ch_adr1[0] ) );
INV_X4 _u0_u18_U201  ( .A(1'b0), .ZN(_u0_u18_ch_am0[31] ) );
INV_X4 _u0_u18_U199  ( .A(1'b0), .ZN(_u0_u18_ch_am0[30] ) );
INV_X4 _u0_u18_U197  ( .A(1'b0), .ZN(_u0_u18_ch_am0[29] ) );
INV_X4 _u0_u18_U195  ( .A(1'b0), .ZN(_u0_u18_ch_am0[28] ) );
INV_X4 _u0_u18_U193  ( .A(1'b0), .ZN(_u0_u18_ch_am0[27] ) );
INV_X4 _u0_u18_U191  ( .A(1'b0), .ZN(_u0_u18_ch_am0[26] ) );
INV_X4 _u0_u18_U189  ( .A(1'b0), .ZN(_u0_u18_ch_am0[25] ) );
INV_X4 _u0_u18_U187  ( .A(1'b0), .ZN(_u0_u18_ch_am0[24] ) );
INV_X4 _u0_u18_U185  ( .A(1'b0), .ZN(_u0_u18_ch_am0[23] ) );
INV_X4 _u0_u18_U183  ( .A(1'b0), .ZN(_u0_u18_ch_am0[22] ) );
INV_X4 _u0_u18_U181  ( .A(1'b0), .ZN(_u0_u18_ch_am0[21] ) );
INV_X4 _u0_u18_U179  ( .A(1'b0), .ZN(_u0_u18_ch_am0[20] ) );
INV_X4 _u0_u18_U177  ( .A(1'b0), .ZN(_u0_u18_ch_am0[19] ) );
INV_X4 _u0_u18_U175  ( .A(1'b0), .ZN(_u0_u18_ch_am0[18] ) );
INV_X4 _u0_u18_U173  ( .A(1'b0), .ZN(_u0_u18_ch_am0[17] ) );
INV_X4 _u0_u18_U171  ( .A(1'b0), .ZN(_u0_u18_ch_am0[16] ) );
INV_X4 _u0_u18_U169  ( .A(1'b0), .ZN(_u0_u18_ch_am0[15] ) );
INV_X4 _u0_u18_U167  ( .A(1'b0), .ZN(_u0_u18_ch_am0[14] ) );
INV_X4 _u0_u18_U165  ( .A(1'b0), .ZN(_u0_u18_ch_am0[13] ) );
INV_X4 _u0_u18_U163  ( .A(1'b0), .ZN(_u0_u18_ch_am0[12] ) );
INV_X4 _u0_u18_U161  ( .A(1'b0), .ZN(_u0_u18_ch_am0[11] ) );
INV_X4 _u0_u18_U159  ( .A(1'b0), .ZN(_u0_u18_ch_am0[10] ) );
INV_X4 _u0_u18_U157  ( .A(1'b0), .ZN(_u0_u18_ch_am0[9] ) );
INV_X4 _u0_u18_U155  ( .A(1'b0), .ZN(_u0_u18_ch_am0[8] ) );
INV_X4 _u0_u18_U153  ( .A(1'b0), .ZN(_u0_u18_ch_am0[7] ) );
INV_X4 _u0_u18_U151  ( .A(1'b0), .ZN(_u0_u18_ch_am0[6] ) );
INV_X4 _u0_u18_U149  ( .A(1'b0), .ZN(_u0_u18_ch_am0[5] ) );
INV_X4 _u0_u18_U147  ( .A(1'b0), .ZN(_u0_u18_ch_am0[4] ) );
INV_X4 _u0_u18_U145  ( .A(1'b1), .ZN(_u0_u18_ch_am0[3] ) );
INV_X4 _u0_u18_U143  ( .A(1'b1), .ZN(_u0_u18_ch_am0[2] ) );
INV_X4 _u0_u18_U141  ( .A(1'b1), .ZN(_u0_u18_ch_am0[1] ) );
INV_X4 _u0_u18_U139  ( .A(1'b1), .ZN(_u0_u18_ch_am0[0] ) );
INV_X4 _u0_u18_U137  ( .A(1'b0), .ZN(_u0_u18_ch_am1[31] ) );
INV_X4 _u0_u18_U135  ( .A(1'b0), .ZN(_u0_u18_ch_am1[30] ) );
INV_X4 _u0_u18_U133  ( .A(1'b0), .ZN(_u0_u18_ch_am1[29] ) );
INV_X4 _u0_u18_U131  ( .A(1'b0), .ZN(_u0_u18_ch_am1[28] ) );
INV_X4 _u0_u18_U129  ( .A(1'b0), .ZN(_u0_u18_ch_am1[27] ) );
INV_X4 _u0_u18_U127  ( .A(1'b0), .ZN(_u0_u18_ch_am1[26] ) );
INV_X4 _u0_u18_U125  ( .A(1'b0), .ZN(_u0_u18_ch_am1[25] ) );
INV_X4 _u0_u18_U123  ( .A(1'b0), .ZN(_u0_u18_ch_am1[24] ) );
INV_X4 _u0_u18_U121  ( .A(1'b0), .ZN(_u0_u18_ch_am1[23] ) );
INV_X4 _u0_u18_U119  ( .A(1'b0), .ZN(_u0_u18_ch_am1[22] ) );
INV_X4 _u0_u18_U117  ( .A(1'b0), .ZN(_u0_u18_ch_am1[21] ) );
INV_X4 _u0_u18_U115  ( .A(1'b0), .ZN(_u0_u18_ch_am1[20] ) );
INV_X4 _u0_u18_U113  ( .A(1'b0), .ZN(_u0_u18_ch_am1[19] ) );
INV_X4 _u0_u18_U111  ( .A(1'b0), .ZN(_u0_u18_ch_am1[18] ) );
INV_X4 _u0_u18_U109  ( .A(1'b0), .ZN(_u0_u18_ch_am1[17] ) );
INV_X4 _u0_u18_U107  ( .A(1'b0), .ZN(_u0_u18_ch_am1[16] ) );
INV_X4 _u0_u18_U105  ( .A(1'b0), .ZN(_u0_u18_ch_am1[15] ) );
INV_X4 _u0_u18_U103  ( .A(1'b0), .ZN(_u0_u18_ch_am1[14] ) );
INV_X4 _u0_u18_U101  ( .A(1'b0), .ZN(_u0_u18_ch_am1[13] ) );
INV_X4 _u0_u18_U99  ( .A(1'b0), .ZN(_u0_u18_ch_am1[12] ) );
INV_X4 _u0_u18_U97  ( .A(1'b0), .ZN(_u0_u18_ch_am1[11] ) );
INV_X4 _u0_u18_U95  ( .A(1'b0), .ZN(_u0_u18_ch_am1[10] ) );
INV_X4 _u0_u18_U93  ( .A(1'b0), .ZN(_u0_u18_ch_am1[9] ) );
INV_X4 _u0_u18_U91  ( .A(1'b0), .ZN(_u0_u18_ch_am1[8] ) );
INV_X4 _u0_u18_U89  ( .A(1'b0), .ZN(_u0_u18_ch_am1[7] ) );
INV_X4 _u0_u18_U87  ( .A(1'b0), .ZN(_u0_u18_ch_am1[6] ) );
INV_X4 _u0_u18_U85  ( .A(1'b0), .ZN(_u0_u18_ch_am1[5] ) );
INV_X4 _u0_u18_U83  ( .A(1'b0), .ZN(_u0_u18_ch_am1[4] ) );
INV_X4 _u0_u18_U81  ( .A(1'b1), .ZN(_u0_u18_ch_am1[3] ) );
INV_X4 _u0_u18_U79  ( .A(1'b1), .ZN(_u0_u18_ch_am1[2] ) );
INV_X4 _u0_u18_U77  ( .A(1'b1), .ZN(_u0_u18_ch_am1[1] ) );
INV_X4 _u0_u18_U75  ( .A(1'b1), .ZN(_u0_u18_ch_am1[0] ) );
INV_X4 _u0_u18_U73  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[31] ) );
INV_X4 _u0_u18_U71  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[30] ) );
INV_X4 _u0_u18_U69  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[29] ) );
INV_X4 _u0_u18_U67  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[28] ) );
INV_X4 _u0_u18_U65  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[27] ) );
INV_X4 _u0_u18_U63  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[26] ) );
INV_X4 _u0_u18_U61  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[25] ) );
INV_X4 _u0_u18_U59  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[24] ) );
INV_X4 _u0_u18_U57  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[23] ) );
INV_X4 _u0_u18_U55  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[22] ) );
INV_X4 _u0_u18_U53  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[21] ) );
INV_X4 _u0_u18_U51  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[20] ) );
INV_X4 _u0_u18_U49  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[19] ) );
INV_X4 _u0_u18_U47  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[18] ) );
INV_X4 _u0_u18_U45  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[17] ) );
INV_X4 _u0_u18_U43  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[16] ) );
INV_X4 _u0_u18_U41  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[15] ) );
INV_X4 _u0_u18_U39  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[14] ) );
INV_X4 _u0_u18_U37  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[13] ) );
INV_X4 _u0_u18_U35  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[12] ) );
INV_X4 _u0_u18_U33  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[11] ) );
INV_X4 _u0_u18_U31  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[10] ) );
INV_X4 _u0_u18_U29  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[9] ) );
INV_X4 _u0_u18_U27  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[8] ) );
INV_X4 _u0_u18_U25  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[7] ) );
INV_X4 _u0_u18_U23  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[6] ) );
INV_X4 _u0_u18_U21  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[5] ) );
INV_X4 _u0_u18_U19  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[4] ) );
INV_X4 _u0_u18_U17  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[3] ) );
INV_X4 _u0_u18_U15  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[2] ) );
INV_X4 _u0_u18_U13  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[1] ) );
INV_X4 _u0_u18_U11  ( .A(1'b1), .ZN(_u0_u18_sw_pointer[0] ) );
INV_X4 _u0_u18_U9  ( .A(1'b1), .ZN(_u0_u18_ch_stop ) );
INV_X4 _u0_u18_U7  ( .A(1'b1), .ZN(_u0_u18_ch_dis ) );
INV_X4 _u0_u18_U5  ( .A(1'b1), .ZN(_u0_u18_int ) );
INV_X4 _u0_u19_U585  ( .A(1'b1), .ZN(_u0_u19_pointer[31] ) );
INV_X4 _u0_u19_U583  ( .A(1'b1), .ZN(_u0_u19_pointer[30] ) );
INV_X4 _u0_u19_U581  ( .A(1'b1), .ZN(_u0_u19_pointer[29] ) );
INV_X4 _u0_u19_U579  ( .A(1'b1), .ZN(_u0_u19_pointer[28] ) );
INV_X4 _u0_u19_U577  ( .A(1'b1), .ZN(_u0_u19_pointer[27] ) );
INV_X4 _u0_u19_U575  ( .A(1'b1), .ZN(_u0_u19_pointer[26] ) );
INV_X4 _u0_u19_U573  ( .A(1'b1), .ZN(_u0_u19_pointer[25] ) );
INV_X4 _u0_u19_U571  ( .A(1'b1), .ZN(_u0_u19_pointer[24] ) );
INV_X4 _u0_u19_U569  ( .A(1'b1), .ZN(_u0_u19_pointer[23] ) );
INV_X4 _u0_u19_U567  ( .A(1'b1), .ZN(_u0_u19_pointer[22] ) );
INV_X4 _u0_u19_U565  ( .A(1'b1), .ZN(_u0_u19_pointer[21] ) );
INV_X4 _u0_u19_U563  ( .A(1'b1), .ZN(_u0_u19_pointer[20] ) );
INV_X4 _u0_u19_U561  ( .A(1'b1), .ZN(_u0_u19_pointer[19] ) );
INV_X4 _u0_u19_U559  ( .A(1'b1), .ZN(_u0_u19_pointer[18] ) );
INV_X4 _u0_u19_U557  ( .A(1'b1), .ZN(_u0_u19_pointer[17] ) );
INV_X4 _u0_u19_U555  ( .A(1'b1), .ZN(_u0_u19_pointer[16] ) );
INV_X4 _u0_u19_U553  ( .A(1'b1), .ZN(_u0_u19_pointer[15] ) );
INV_X4 _u0_u19_U551  ( .A(1'b1), .ZN(_u0_u19_pointer[14] ) );
INV_X4 _u0_u19_U549  ( .A(1'b1), .ZN(_u0_u19_pointer[13] ) );
INV_X4 _u0_u19_U547  ( .A(1'b1), .ZN(_u0_u19_pointer[12] ) );
INV_X4 _u0_u19_U545  ( .A(1'b1), .ZN(_u0_u19_pointer[11] ) );
INV_X4 _u0_u19_U543  ( .A(1'b1), .ZN(_u0_u19_pointer[10] ) );
INV_X4 _u0_u19_U541  ( .A(1'b1), .ZN(_u0_u19_pointer[9] ) );
INV_X4 _u0_u19_U539  ( .A(1'b1), .ZN(_u0_u19_pointer[8] ) );
INV_X4 _u0_u19_U537  ( .A(1'b1), .ZN(_u0_u19_pointer[7] ) );
INV_X4 _u0_u19_U535  ( .A(1'b1), .ZN(_u0_u19_pointer[6] ) );
INV_X4 _u0_u19_U533  ( .A(1'b1), .ZN(_u0_u19_pointer[5] ) );
INV_X4 _u0_u19_U531  ( .A(1'b1), .ZN(_u0_u19_pointer[4] ) );
INV_X4 _u0_u19_U529  ( .A(1'b1), .ZN(_u0_u19_pointer[3] ) );
INV_X4 _u0_u19_U527  ( .A(1'b1), .ZN(_u0_u19_pointer[2] ) );
INV_X4 _u0_u19_U525  ( .A(1'b1), .ZN(_u0_u19_pointer[1] ) );
INV_X4 _u0_u19_U523  ( .A(1'b1), .ZN(_u0_u19_pointer[0] ) );
INV_X4 _u0_u19_U521  ( .A(1'b1), .ZN(_u0_u19_pointer_s[31] ) );
INV_X4 _u0_u19_U519  ( .A(1'b1), .ZN(_u0_u19_pointer_s[30] ) );
INV_X4 _u0_u19_U517  ( .A(1'b1), .ZN(_u0_u19_pointer_s[29] ) );
INV_X4 _u0_u19_U515  ( .A(1'b1), .ZN(_u0_u19_pointer_s[28] ) );
INV_X4 _u0_u19_U513  ( .A(1'b1), .ZN(_u0_u19_pointer_s[27] ) );
INV_X4 _u0_u19_U511  ( .A(1'b1), .ZN(_u0_u19_pointer_s[26] ) );
INV_X4 _u0_u19_U509  ( .A(1'b1), .ZN(_u0_u19_pointer_s[25] ) );
INV_X4 _u0_u19_U507  ( .A(1'b1), .ZN(_u0_u19_pointer_s[24] ) );
INV_X4 _u0_u19_U505  ( .A(1'b1), .ZN(_u0_u19_pointer_s[23] ) );
INV_X4 _u0_u19_U503  ( .A(1'b1), .ZN(_u0_u19_pointer_s[22] ) );
INV_X4 _u0_u19_U501  ( .A(1'b1), .ZN(_u0_u19_pointer_s[21] ) );
INV_X4 _u0_u19_U499  ( .A(1'b1), .ZN(_u0_u19_pointer_s[20] ) );
INV_X4 _u0_u19_U497  ( .A(1'b1), .ZN(_u0_u19_pointer_s[19] ) );
INV_X4 _u0_u19_U495  ( .A(1'b1), .ZN(_u0_u19_pointer_s[18] ) );
INV_X4 _u0_u19_U493  ( .A(1'b1), .ZN(_u0_u19_pointer_s[17] ) );
INV_X4 _u0_u19_U491  ( .A(1'b1), .ZN(_u0_u19_pointer_s[16] ) );
INV_X4 _u0_u19_U489  ( .A(1'b1), .ZN(_u0_u19_pointer_s[15] ) );
INV_X4 _u0_u19_U487  ( .A(1'b1), .ZN(_u0_u19_pointer_s[14] ) );
INV_X4 _u0_u19_U485  ( .A(1'b1), .ZN(_u0_u19_pointer_s[13] ) );
INV_X4 _u0_u19_U483  ( .A(1'b1), .ZN(_u0_u19_pointer_s[12] ) );
INV_X4 _u0_u19_U481  ( .A(1'b1), .ZN(_u0_u19_pointer_s[11] ) );
INV_X4 _u0_u19_U479  ( .A(1'b1), .ZN(_u0_u19_pointer_s[10] ) );
INV_X4 _u0_u19_U477  ( .A(1'b1), .ZN(_u0_u19_pointer_s[9] ) );
INV_X4 _u0_u19_U475  ( .A(1'b1), .ZN(_u0_u19_pointer_s[8] ) );
INV_X4 _u0_u19_U473  ( .A(1'b1), .ZN(_u0_u19_pointer_s[7] ) );
INV_X4 _u0_u19_U471  ( .A(1'b1), .ZN(_u0_u19_pointer_s[6] ) );
INV_X4 _u0_u19_U469  ( .A(1'b1), .ZN(_u0_u19_pointer_s[5] ) );
INV_X4 _u0_u19_U467  ( .A(1'b1), .ZN(_u0_u19_pointer_s[4] ) );
INV_X4 _u0_u19_U465  ( .A(1'b1), .ZN(_u0_u19_pointer_s[3] ) );
INV_X4 _u0_u19_U463  ( .A(1'b1), .ZN(_u0_u19_pointer_s[2] ) );
INV_X4 _u0_u19_U461  ( .A(1'b1), .ZN(_u0_u19_pointer_s[1] ) );
INV_X4 _u0_u19_U459  ( .A(1'b1), .ZN(_u0_u19_pointer_s[0] ) );
INV_X4 _u0_u19_U457  ( .A(1'b1), .ZN(_u0_u19_ch_csr[31] ) );
INV_X4 _u0_u19_U455  ( .A(1'b1), .ZN(_u0_u19_ch_csr[30] ) );
INV_X4 _u0_u19_U453  ( .A(1'b1), .ZN(_u0_u19_ch_csr[29] ) );
INV_X4 _u0_u19_U451  ( .A(1'b1), .ZN(_u0_u19_ch_csr[28] ) );
INV_X4 _u0_u19_U449  ( .A(1'b1), .ZN(_u0_u19_ch_csr[27] ) );
INV_X4 _u0_u19_U447  ( .A(1'b1), .ZN(_u0_u19_ch_csr[26] ) );
INV_X4 _u0_u19_U445  ( .A(1'b1), .ZN(_u0_u19_ch_csr[25] ) );
INV_X4 _u0_u19_U443  ( .A(1'b1), .ZN(_u0_u19_ch_csr[24] ) );
INV_X4 _u0_u19_U441  ( .A(1'b1), .ZN(_u0_u19_ch_csr[23] ) );
INV_X4 _u0_u19_U439  ( .A(1'b1), .ZN(_u0_u19_ch_csr[22] ) );
INV_X4 _u0_u19_U437  ( .A(1'b1), .ZN(_u0_u19_ch_csr[21] ) );
INV_X4 _u0_u19_U435  ( .A(1'b1), .ZN(_u0_u19_ch_csr[20] ) );
INV_X4 _u0_u19_U433  ( .A(1'b1), .ZN(_u0_u19_ch_csr[19] ) );
INV_X4 _u0_u19_U431  ( .A(1'b1), .ZN(_u0_u19_ch_csr[18] ) );
INV_X4 _u0_u19_U429  ( .A(1'b1), .ZN(_u0_u19_ch_csr[17] ) );
INV_X4 _u0_u19_U427  ( .A(1'b1), .ZN(_u0_u19_ch_csr[16] ) );
INV_X4 _u0_u19_U425  ( .A(1'b1), .ZN(_u0_u19_ch_csr[15] ) );
INV_X4 _u0_u19_U423  ( .A(1'b1), .ZN(_u0_u19_ch_csr[14] ) );
INV_X4 _u0_u19_U421  ( .A(1'b1), .ZN(_u0_u19_ch_csr[13] ) );
INV_X4 _u0_u19_U419  ( .A(1'b1), .ZN(_u0_u19_ch_csr[12] ) );
INV_X4 _u0_u19_U417  ( .A(1'b1), .ZN(_u0_u19_ch_csr[11] ) );
INV_X4 _u0_u19_U415  ( .A(1'b1), .ZN(_u0_u19_ch_csr[10] ) );
INV_X4 _u0_u19_U413  ( .A(1'b1), .ZN(_u0_u19_ch_csr[9] ) );
INV_X4 _u0_u19_U411  ( .A(1'b1), .ZN(_u0_u19_ch_csr[8] ) );
INV_X4 _u0_u19_U409  ( .A(1'b1), .ZN(_u0_u19_ch_csr[7] ) );
INV_X4 _u0_u19_U407  ( .A(1'b1), .ZN(_u0_u19_ch_csr[6] ) );
INV_X4 _u0_u19_U405  ( .A(1'b1), .ZN(_u0_u19_ch_csr[5] ) );
INV_X4 _u0_u19_U403  ( .A(1'b1), .ZN(_u0_u19_ch_csr[4] ) );
INV_X4 _u0_u19_U401  ( .A(1'b1), .ZN(_u0_u19_ch_csr[3] ) );
INV_X4 _u0_u19_U399  ( .A(1'b1), .ZN(_u0_u19_ch_csr[2] ) );
INV_X4 _u0_u19_U397  ( .A(1'b1), .ZN(_u0_u19_ch_csr[1] ) );
INV_X4 _u0_u19_U395  ( .A(1'b1), .ZN(_u0_u19_ch_csr[0] ) );
INV_X4 _u0_u19_U393  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[31] ) );
INV_X4 _u0_u19_U391  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[30] ) );
INV_X4 _u0_u19_U389  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[29] ) );
INV_X4 _u0_u19_U387  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[28] ) );
INV_X4 _u0_u19_U385  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[27] ) );
INV_X4 _u0_u19_U383  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[26] ) );
INV_X4 _u0_u19_U381  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[25] ) );
INV_X4 _u0_u19_U379  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[24] ) );
INV_X4 _u0_u19_U377  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[23] ) );
INV_X4 _u0_u19_U375  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[22] ) );
INV_X4 _u0_u19_U373  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[21] ) );
INV_X4 _u0_u19_U371  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[20] ) );
INV_X4 _u0_u19_U369  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[19] ) );
INV_X4 _u0_u19_U367  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[18] ) );
INV_X4 _u0_u19_U365  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[17] ) );
INV_X4 _u0_u19_U363  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[16] ) );
INV_X4 _u0_u19_U361  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[15] ) );
INV_X4 _u0_u19_U359  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[14] ) );
INV_X4 _u0_u19_U357  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[13] ) );
INV_X4 _u0_u19_U355  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[12] ) );
INV_X4 _u0_u19_U353  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[11] ) );
INV_X4 _u0_u19_U351  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[10] ) );
INV_X4 _u0_u19_U349  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[9] ) );
INV_X4 _u0_u19_U347  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[8] ) );
INV_X4 _u0_u19_U345  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[7] ) );
INV_X4 _u0_u19_U343  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[6] ) );
INV_X4 _u0_u19_U341  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[5] ) );
INV_X4 _u0_u19_U339  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[4] ) );
INV_X4 _u0_u19_U337  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[3] ) );
INV_X4 _u0_u19_U335  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[2] ) );
INV_X4 _u0_u19_U333  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[1] ) );
INV_X4 _u0_u19_U331  ( .A(1'b1), .ZN(_u0_u19_ch_txsz[0] ) );
INV_X4 _u0_u19_U329  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[31] ) );
INV_X4 _u0_u19_U327  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[30] ) );
INV_X4 _u0_u19_U325  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[29] ) );
INV_X4 _u0_u19_U323  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[28] ) );
INV_X4 _u0_u19_U321  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[27] ) );
INV_X4 _u0_u19_U319  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[26] ) );
INV_X4 _u0_u19_U317  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[25] ) );
INV_X4 _u0_u19_U315  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[24] ) );
INV_X4 _u0_u19_U313  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[23] ) );
INV_X4 _u0_u19_U311  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[22] ) );
INV_X4 _u0_u19_U309  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[21] ) );
INV_X4 _u0_u19_U307  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[20] ) );
INV_X4 _u0_u19_U305  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[19] ) );
INV_X4 _u0_u19_U303  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[18] ) );
INV_X4 _u0_u19_U301  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[17] ) );
INV_X4 _u0_u19_U299  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[16] ) );
INV_X4 _u0_u19_U297  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[15] ) );
INV_X4 _u0_u19_U295  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[14] ) );
INV_X4 _u0_u19_U293  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[13] ) );
INV_X4 _u0_u19_U291  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[12] ) );
INV_X4 _u0_u19_U289  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[11] ) );
INV_X4 _u0_u19_U287  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[10] ) );
INV_X4 _u0_u19_U285  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[9] ) );
INV_X4 _u0_u19_U283  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[8] ) );
INV_X4 _u0_u19_U281  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[7] ) );
INV_X4 _u0_u19_U279  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[6] ) );
INV_X4 _u0_u19_U277  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[5] ) );
INV_X4 _u0_u19_U275  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[4] ) );
INV_X4 _u0_u19_U273  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[3] ) );
INV_X4 _u0_u19_U271  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[2] ) );
INV_X4 _u0_u19_U269  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[1] ) );
INV_X4 _u0_u19_U267  ( .A(1'b1), .ZN(_u0_u19_ch_adr0[0] ) );
INV_X4 _u0_u19_U265  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[31] ) );
INV_X4 _u0_u19_U263  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[30] ) );
INV_X4 _u0_u19_U261  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[29] ) );
INV_X4 _u0_u19_U259  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[28] ) );
INV_X4 _u0_u19_U257  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[27] ) );
INV_X4 _u0_u19_U255  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[26] ) );
INV_X4 _u0_u19_U253  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[25] ) );
INV_X4 _u0_u19_U251  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[24] ) );
INV_X4 _u0_u19_U249  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[23] ) );
INV_X4 _u0_u19_U247  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[22] ) );
INV_X4 _u0_u19_U245  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[21] ) );
INV_X4 _u0_u19_U243  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[20] ) );
INV_X4 _u0_u19_U241  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[19] ) );
INV_X4 _u0_u19_U239  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[18] ) );
INV_X4 _u0_u19_U237  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[17] ) );
INV_X4 _u0_u19_U235  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[16] ) );
INV_X4 _u0_u19_U233  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[15] ) );
INV_X4 _u0_u19_U231  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[14] ) );
INV_X4 _u0_u19_U229  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[13] ) );
INV_X4 _u0_u19_U227  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[12] ) );
INV_X4 _u0_u19_U225  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[11] ) );
INV_X4 _u0_u19_U223  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[10] ) );
INV_X4 _u0_u19_U221  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[9] ) );
INV_X4 _u0_u19_U219  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[8] ) );
INV_X4 _u0_u19_U217  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[7] ) );
INV_X4 _u0_u19_U215  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[6] ) );
INV_X4 _u0_u19_U213  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[5] ) );
INV_X4 _u0_u19_U211  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[4] ) );
INV_X4 _u0_u19_U209  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[3] ) );
INV_X4 _u0_u19_U207  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[2] ) );
INV_X4 _u0_u19_U205  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[1] ) );
INV_X4 _u0_u19_U203  ( .A(1'b1), .ZN(_u0_u19_ch_adr1[0] ) );
INV_X4 _u0_u19_U201  ( .A(1'b0), .ZN(_u0_u19_ch_am0[31] ) );
INV_X4 _u0_u19_U199  ( .A(1'b0), .ZN(_u0_u19_ch_am0[30] ) );
INV_X4 _u0_u19_U197  ( .A(1'b0), .ZN(_u0_u19_ch_am0[29] ) );
INV_X4 _u0_u19_U195  ( .A(1'b0), .ZN(_u0_u19_ch_am0[28] ) );
INV_X4 _u0_u19_U193  ( .A(1'b0), .ZN(_u0_u19_ch_am0[27] ) );
INV_X4 _u0_u19_U191  ( .A(1'b0), .ZN(_u0_u19_ch_am0[26] ) );
INV_X4 _u0_u19_U189  ( .A(1'b0), .ZN(_u0_u19_ch_am0[25] ) );
INV_X4 _u0_u19_U187  ( .A(1'b0), .ZN(_u0_u19_ch_am0[24] ) );
INV_X4 _u0_u19_U185  ( .A(1'b0), .ZN(_u0_u19_ch_am0[23] ) );
INV_X4 _u0_u19_U183  ( .A(1'b0), .ZN(_u0_u19_ch_am0[22] ) );
INV_X4 _u0_u19_U181  ( .A(1'b0), .ZN(_u0_u19_ch_am0[21] ) );
INV_X4 _u0_u19_U179  ( .A(1'b0), .ZN(_u0_u19_ch_am0[20] ) );
INV_X4 _u0_u19_U177  ( .A(1'b0), .ZN(_u0_u19_ch_am0[19] ) );
INV_X4 _u0_u19_U175  ( .A(1'b0), .ZN(_u0_u19_ch_am0[18] ) );
INV_X4 _u0_u19_U173  ( .A(1'b0), .ZN(_u0_u19_ch_am0[17] ) );
INV_X4 _u0_u19_U171  ( .A(1'b0), .ZN(_u0_u19_ch_am0[16] ) );
INV_X4 _u0_u19_U169  ( .A(1'b0), .ZN(_u0_u19_ch_am0[15] ) );
INV_X4 _u0_u19_U167  ( .A(1'b0), .ZN(_u0_u19_ch_am0[14] ) );
INV_X4 _u0_u19_U165  ( .A(1'b0), .ZN(_u0_u19_ch_am0[13] ) );
INV_X4 _u0_u19_U163  ( .A(1'b0), .ZN(_u0_u19_ch_am0[12] ) );
INV_X4 _u0_u19_U161  ( .A(1'b0), .ZN(_u0_u19_ch_am0[11] ) );
INV_X4 _u0_u19_U159  ( .A(1'b0), .ZN(_u0_u19_ch_am0[10] ) );
INV_X4 _u0_u19_U157  ( .A(1'b0), .ZN(_u0_u19_ch_am0[9] ) );
INV_X4 _u0_u19_U155  ( .A(1'b0), .ZN(_u0_u19_ch_am0[8] ) );
INV_X4 _u0_u19_U153  ( .A(1'b0), .ZN(_u0_u19_ch_am0[7] ) );
INV_X4 _u0_u19_U151  ( .A(1'b0), .ZN(_u0_u19_ch_am0[6] ) );
INV_X4 _u0_u19_U149  ( .A(1'b0), .ZN(_u0_u19_ch_am0[5] ) );
INV_X4 _u0_u19_U147  ( .A(1'b0), .ZN(_u0_u19_ch_am0[4] ) );
INV_X4 _u0_u19_U145  ( .A(1'b1), .ZN(_u0_u19_ch_am0[3] ) );
INV_X4 _u0_u19_U143  ( .A(1'b1), .ZN(_u0_u19_ch_am0[2] ) );
INV_X4 _u0_u19_U141  ( .A(1'b1), .ZN(_u0_u19_ch_am0[1] ) );
INV_X4 _u0_u19_U139  ( .A(1'b1), .ZN(_u0_u19_ch_am0[0] ) );
INV_X4 _u0_u19_U137  ( .A(1'b0), .ZN(_u0_u19_ch_am1[31] ) );
INV_X4 _u0_u19_U135  ( .A(1'b0), .ZN(_u0_u19_ch_am1[30] ) );
INV_X4 _u0_u19_U133  ( .A(1'b0), .ZN(_u0_u19_ch_am1[29] ) );
INV_X4 _u0_u19_U131  ( .A(1'b0), .ZN(_u0_u19_ch_am1[28] ) );
INV_X4 _u0_u19_U129  ( .A(1'b0), .ZN(_u0_u19_ch_am1[27] ) );
INV_X4 _u0_u19_U127  ( .A(1'b0), .ZN(_u0_u19_ch_am1[26] ) );
INV_X4 _u0_u19_U125  ( .A(1'b0), .ZN(_u0_u19_ch_am1[25] ) );
INV_X4 _u0_u19_U123  ( .A(1'b0), .ZN(_u0_u19_ch_am1[24] ) );
INV_X4 _u0_u19_U121  ( .A(1'b0), .ZN(_u0_u19_ch_am1[23] ) );
INV_X4 _u0_u19_U119  ( .A(1'b0), .ZN(_u0_u19_ch_am1[22] ) );
INV_X4 _u0_u19_U117  ( .A(1'b0), .ZN(_u0_u19_ch_am1[21] ) );
INV_X4 _u0_u19_U115  ( .A(1'b0), .ZN(_u0_u19_ch_am1[20] ) );
INV_X4 _u0_u19_U113  ( .A(1'b0), .ZN(_u0_u19_ch_am1[19] ) );
INV_X4 _u0_u19_U111  ( .A(1'b0), .ZN(_u0_u19_ch_am1[18] ) );
INV_X4 _u0_u19_U109  ( .A(1'b0), .ZN(_u0_u19_ch_am1[17] ) );
INV_X4 _u0_u19_U107  ( .A(1'b0), .ZN(_u0_u19_ch_am1[16] ) );
INV_X4 _u0_u19_U105  ( .A(1'b0), .ZN(_u0_u19_ch_am1[15] ) );
INV_X4 _u0_u19_U103  ( .A(1'b0), .ZN(_u0_u19_ch_am1[14] ) );
INV_X4 _u0_u19_U101  ( .A(1'b0), .ZN(_u0_u19_ch_am1[13] ) );
INV_X4 _u0_u19_U99  ( .A(1'b0), .ZN(_u0_u19_ch_am1[12] ) );
INV_X4 _u0_u19_U97  ( .A(1'b0), .ZN(_u0_u19_ch_am1[11] ) );
INV_X4 _u0_u19_U95  ( .A(1'b0), .ZN(_u0_u19_ch_am1[10] ) );
INV_X4 _u0_u19_U93  ( .A(1'b0), .ZN(_u0_u19_ch_am1[9] ) );
INV_X4 _u0_u19_U91  ( .A(1'b0), .ZN(_u0_u19_ch_am1[8] ) );
INV_X4 _u0_u19_U89  ( .A(1'b0), .ZN(_u0_u19_ch_am1[7] ) );
INV_X4 _u0_u19_U87  ( .A(1'b0), .ZN(_u0_u19_ch_am1[6] ) );
INV_X4 _u0_u19_U85  ( .A(1'b0), .ZN(_u0_u19_ch_am1[5] ) );
INV_X4 _u0_u19_U83  ( .A(1'b0), .ZN(_u0_u19_ch_am1[4] ) );
INV_X4 _u0_u19_U81  ( .A(1'b1), .ZN(_u0_u19_ch_am1[3] ) );
INV_X4 _u0_u19_U79  ( .A(1'b1), .ZN(_u0_u19_ch_am1[2] ) );
INV_X4 _u0_u19_U77  ( .A(1'b1), .ZN(_u0_u19_ch_am1[1] ) );
INV_X4 _u0_u19_U75  ( .A(1'b1), .ZN(_u0_u19_ch_am1[0] ) );
INV_X4 _u0_u19_U73  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[31] ) );
INV_X4 _u0_u19_U71  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[30] ) );
INV_X4 _u0_u19_U69  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[29] ) );
INV_X4 _u0_u19_U67  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[28] ) );
INV_X4 _u0_u19_U65  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[27] ) );
INV_X4 _u0_u19_U63  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[26] ) );
INV_X4 _u0_u19_U61  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[25] ) );
INV_X4 _u0_u19_U59  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[24] ) );
INV_X4 _u0_u19_U57  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[23] ) );
INV_X4 _u0_u19_U55  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[22] ) );
INV_X4 _u0_u19_U53  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[21] ) );
INV_X4 _u0_u19_U51  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[20] ) );
INV_X4 _u0_u19_U49  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[19] ) );
INV_X4 _u0_u19_U47  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[18] ) );
INV_X4 _u0_u19_U45  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[17] ) );
INV_X4 _u0_u19_U43  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[16] ) );
INV_X4 _u0_u19_U41  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[15] ) );
INV_X4 _u0_u19_U39  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[14] ) );
INV_X4 _u0_u19_U37  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[13] ) );
INV_X4 _u0_u19_U35  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[12] ) );
INV_X4 _u0_u19_U33  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[11] ) );
INV_X4 _u0_u19_U31  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[10] ) );
INV_X4 _u0_u19_U29  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[9] ) );
INV_X4 _u0_u19_U27  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[8] ) );
INV_X4 _u0_u19_U25  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[7] ) );
INV_X4 _u0_u19_U23  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[6] ) );
INV_X4 _u0_u19_U21  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[5] ) );
INV_X4 _u0_u19_U19  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[4] ) );
INV_X4 _u0_u19_U17  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[3] ) );
INV_X4 _u0_u19_U15  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[2] ) );
INV_X4 _u0_u19_U13  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[1] ) );
INV_X4 _u0_u19_U11  ( .A(1'b1), .ZN(_u0_u19_sw_pointer[0] ) );
INV_X4 _u0_u19_U9  ( .A(1'b1), .ZN(_u0_u19_ch_stop ) );
INV_X4 _u0_u19_U7  ( .A(1'b1), .ZN(_u0_u19_ch_dis ) );
INV_X4 _u0_u19_U5  ( .A(1'b1), .ZN(_u0_u19_int ) );
INV_X4 _u0_u20_U585  ( .A(1'b1), .ZN(_u0_u20_pointer[31] ) );
INV_X4 _u0_u20_U583  ( .A(1'b1), .ZN(_u0_u20_pointer[30] ) );
INV_X4 _u0_u20_U581  ( .A(1'b1), .ZN(_u0_u20_pointer[29] ) );
INV_X4 _u0_u20_U579  ( .A(1'b1), .ZN(_u0_u20_pointer[28] ) );
INV_X4 _u0_u20_U577  ( .A(1'b1), .ZN(_u0_u20_pointer[27] ) );
INV_X4 _u0_u20_U575  ( .A(1'b1), .ZN(_u0_u20_pointer[26] ) );
INV_X4 _u0_u20_U573  ( .A(1'b1), .ZN(_u0_u20_pointer[25] ) );
INV_X4 _u0_u20_U571  ( .A(1'b1), .ZN(_u0_u20_pointer[24] ) );
INV_X4 _u0_u20_U569  ( .A(1'b1), .ZN(_u0_u20_pointer[23] ) );
INV_X4 _u0_u20_U567  ( .A(1'b1), .ZN(_u0_u20_pointer[22] ) );
INV_X4 _u0_u20_U565  ( .A(1'b1), .ZN(_u0_u20_pointer[21] ) );
INV_X4 _u0_u20_U563  ( .A(1'b1), .ZN(_u0_u20_pointer[20] ) );
INV_X4 _u0_u20_U561  ( .A(1'b1), .ZN(_u0_u20_pointer[19] ) );
INV_X4 _u0_u20_U559  ( .A(1'b1), .ZN(_u0_u20_pointer[18] ) );
INV_X4 _u0_u20_U557  ( .A(1'b1), .ZN(_u0_u20_pointer[17] ) );
INV_X4 _u0_u20_U555  ( .A(1'b1), .ZN(_u0_u20_pointer[16] ) );
INV_X4 _u0_u20_U553  ( .A(1'b1), .ZN(_u0_u20_pointer[15] ) );
INV_X4 _u0_u20_U551  ( .A(1'b1), .ZN(_u0_u20_pointer[14] ) );
INV_X4 _u0_u20_U549  ( .A(1'b1), .ZN(_u0_u20_pointer[13] ) );
INV_X4 _u0_u20_U547  ( .A(1'b1), .ZN(_u0_u20_pointer[12] ) );
INV_X4 _u0_u20_U545  ( .A(1'b1), .ZN(_u0_u20_pointer[11] ) );
INV_X4 _u0_u20_U543  ( .A(1'b1), .ZN(_u0_u20_pointer[10] ) );
INV_X4 _u0_u20_U541  ( .A(1'b1), .ZN(_u0_u20_pointer[9] ) );
INV_X4 _u0_u20_U539  ( .A(1'b1), .ZN(_u0_u20_pointer[8] ) );
INV_X4 _u0_u20_U537  ( .A(1'b1), .ZN(_u0_u20_pointer[7] ) );
INV_X4 _u0_u20_U535  ( .A(1'b1), .ZN(_u0_u20_pointer[6] ) );
INV_X4 _u0_u20_U533  ( .A(1'b1), .ZN(_u0_u20_pointer[5] ) );
INV_X4 _u0_u20_U531  ( .A(1'b1), .ZN(_u0_u20_pointer[4] ) );
INV_X4 _u0_u20_U529  ( .A(1'b1), .ZN(_u0_u20_pointer[3] ) );
INV_X4 _u0_u20_U527  ( .A(1'b1), .ZN(_u0_u20_pointer[2] ) );
INV_X4 _u0_u20_U525  ( .A(1'b1), .ZN(_u0_u20_pointer[1] ) );
INV_X4 _u0_u20_U523  ( .A(1'b1), .ZN(_u0_u20_pointer[0] ) );
INV_X4 _u0_u20_U521  ( .A(1'b1), .ZN(_u0_u20_pointer_s[31] ) );
INV_X4 _u0_u20_U519  ( .A(1'b1), .ZN(_u0_u20_pointer_s[30] ) );
INV_X4 _u0_u20_U517  ( .A(1'b1), .ZN(_u0_u20_pointer_s[29] ) );
INV_X4 _u0_u20_U515  ( .A(1'b1), .ZN(_u0_u20_pointer_s[28] ) );
INV_X4 _u0_u20_U513  ( .A(1'b1), .ZN(_u0_u20_pointer_s[27] ) );
INV_X4 _u0_u20_U511  ( .A(1'b1), .ZN(_u0_u20_pointer_s[26] ) );
INV_X4 _u0_u20_U509  ( .A(1'b1), .ZN(_u0_u20_pointer_s[25] ) );
INV_X4 _u0_u20_U507  ( .A(1'b1), .ZN(_u0_u20_pointer_s[24] ) );
INV_X4 _u0_u20_U505  ( .A(1'b1), .ZN(_u0_u20_pointer_s[23] ) );
INV_X4 _u0_u20_U503  ( .A(1'b1), .ZN(_u0_u20_pointer_s[22] ) );
INV_X4 _u0_u20_U501  ( .A(1'b1), .ZN(_u0_u20_pointer_s[21] ) );
INV_X4 _u0_u20_U499  ( .A(1'b1), .ZN(_u0_u20_pointer_s[20] ) );
INV_X4 _u0_u20_U497  ( .A(1'b1), .ZN(_u0_u20_pointer_s[19] ) );
INV_X4 _u0_u20_U495  ( .A(1'b1), .ZN(_u0_u20_pointer_s[18] ) );
INV_X4 _u0_u20_U493  ( .A(1'b1), .ZN(_u0_u20_pointer_s[17] ) );
INV_X4 _u0_u20_U491  ( .A(1'b1), .ZN(_u0_u20_pointer_s[16] ) );
INV_X4 _u0_u20_U489  ( .A(1'b1), .ZN(_u0_u20_pointer_s[15] ) );
INV_X4 _u0_u20_U487  ( .A(1'b1), .ZN(_u0_u20_pointer_s[14] ) );
INV_X4 _u0_u20_U485  ( .A(1'b1), .ZN(_u0_u20_pointer_s[13] ) );
INV_X4 _u0_u20_U483  ( .A(1'b1), .ZN(_u0_u20_pointer_s[12] ) );
INV_X4 _u0_u20_U481  ( .A(1'b1), .ZN(_u0_u20_pointer_s[11] ) );
INV_X4 _u0_u20_U479  ( .A(1'b1), .ZN(_u0_u20_pointer_s[10] ) );
INV_X4 _u0_u20_U477  ( .A(1'b1), .ZN(_u0_u20_pointer_s[9] ) );
INV_X4 _u0_u20_U475  ( .A(1'b1), .ZN(_u0_u20_pointer_s[8] ) );
INV_X4 _u0_u20_U473  ( .A(1'b1), .ZN(_u0_u20_pointer_s[7] ) );
INV_X4 _u0_u20_U471  ( .A(1'b1), .ZN(_u0_u20_pointer_s[6] ) );
INV_X4 _u0_u20_U469  ( .A(1'b1), .ZN(_u0_u20_pointer_s[5] ) );
INV_X4 _u0_u20_U467  ( .A(1'b1), .ZN(_u0_u20_pointer_s[4] ) );
INV_X4 _u0_u20_U465  ( .A(1'b1), .ZN(_u0_u20_pointer_s[3] ) );
INV_X4 _u0_u20_U463  ( .A(1'b1), .ZN(_u0_u20_pointer_s[2] ) );
INV_X4 _u0_u20_U461  ( .A(1'b1), .ZN(_u0_u20_pointer_s[1] ) );
INV_X4 _u0_u20_U459  ( .A(1'b1), .ZN(_u0_u20_pointer_s[0] ) );
INV_X4 _u0_u20_U457  ( .A(1'b1), .ZN(_u0_u20_ch_csr[31] ) );
INV_X4 _u0_u20_U455  ( .A(1'b1), .ZN(_u0_u20_ch_csr[30] ) );
INV_X4 _u0_u20_U453  ( .A(1'b1), .ZN(_u0_u20_ch_csr[29] ) );
INV_X4 _u0_u20_U451  ( .A(1'b1), .ZN(_u0_u20_ch_csr[28] ) );
INV_X4 _u0_u20_U449  ( .A(1'b1), .ZN(_u0_u20_ch_csr[27] ) );
INV_X4 _u0_u20_U447  ( .A(1'b1), .ZN(_u0_u20_ch_csr[26] ) );
INV_X4 _u0_u20_U445  ( .A(1'b1), .ZN(_u0_u20_ch_csr[25] ) );
INV_X4 _u0_u20_U443  ( .A(1'b1), .ZN(_u0_u20_ch_csr[24] ) );
INV_X4 _u0_u20_U441  ( .A(1'b1), .ZN(_u0_u20_ch_csr[23] ) );
INV_X4 _u0_u20_U439  ( .A(1'b1), .ZN(_u0_u20_ch_csr[22] ) );
INV_X4 _u0_u20_U437  ( .A(1'b1), .ZN(_u0_u20_ch_csr[21] ) );
INV_X4 _u0_u20_U435  ( .A(1'b1), .ZN(_u0_u20_ch_csr[20] ) );
INV_X4 _u0_u20_U433  ( .A(1'b1), .ZN(_u0_u20_ch_csr[19] ) );
INV_X4 _u0_u20_U431  ( .A(1'b1), .ZN(_u0_u20_ch_csr[18] ) );
INV_X4 _u0_u20_U429  ( .A(1'b1), .ZN(_u0_u20_ch_csr[17] ) );
INV_X4 _u0_u20_U427  ( .A(1'b1), .ZN(_u0_u20_ch_csr[16] ) );
INV_X4 _u0_u20_U425  ( .A(1'b1), .ZN(_u0_u20_ch_csr[15] ) );
INV_X4 _u0_u20_U423  ( .A(1'b1), .ZN(_u0_u20_ch_csr[14] ) );
INV_X4 _u0_u20_U421  ( .A(1'b1), .ZN(_u0_u20_ch_csr[13] ) );
INV_X4 _u0_u20_U419  ( .A(1'b1), .ZN(_u0_u20_ch_csr[12] ) );
INV_X4 _u0_u20_U417  ( .A(1'b1), .ZN(_u0_u20_ch_csr[11] ) );
INV_X4 _u0_u20_U415  ( .A(1'b1), .ZN(_u0_u20_ch_csr[10] ) );
INV_X4 _u0_u20_U413  ( .A(1'b1), .ZN(_u0_u20_ch_csr[9] ) );
INV_X4 _u0_u20_U411  ( .A(1'b1), .ZN(_u0_u20_ch_csr[8] ) );
INV_X4 _u0_u20_U409  ( .A(1'b1), .ZN(_u0_u20_ch_csr[7] ) );
INV_X4 _u0_u20_U407  ( .A(1'b1), .ZN(_u0_u20_ch_csr[6] ) );
INV_X4 _u0_u20_U405  ( .A(1'b1), .ZN(_u0_u20_ch_csr[5] ) );
INV_X4 _u0_u20_U403  ( .A(1'b1), .ZN(_u0_u20_ch_csr[4] ) );
INV_X4 _u0_u20_U401  ( .A(1'b1), .ZN(_u0_u20_ch_csr[3] ) );
INV_X4 _u0_u20_U399  ( .A(1'b1), .ZN(_u0_u20_ch_csr[2] ) );
INV_X4 _u0_u20_U397  ( .A(1'b1), .ZN(_u0_u20_ch_csr[1] ) );
INV_X4 _u0_u20_U395  ( .A(1'b1), .ZN(_u0_u20_ch_csr[0] ) );
INV_X4 _u0_u20_U393  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[31] ) );
INV_X4 _u0_u20_U391  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[30] ) );
INV_X4 _u0_u20_U389  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[29] ) );
INV_X4 _u0_u20_U387  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[28] ) );
INV_X4 _u0_u20_U385  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[27] ) );
INV_X4 _u0_u20_U383  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[26] ) );
INV_X4 _u0_u20_U381  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[25] ) );
INV_X4 _u0_u20_U379  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[24] ) );
INV_X4 _u0_u20_U377  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[23] ) );
INV_X4 _u0_u20_U375  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[22] ) );
INV_X4 _u0_u20_U373  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[21] ) );
INV_X4 _u0_u20_U371  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[20] ) );
INV_X4 _u0_u20_U369  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[19] ) );
INV_X4 _u0_u20_U367  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[18] ) );
INV_X4 _u0_u20_U365  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[17] ) );
INV_X4 _u0_u20_U363  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[16] ) );
INV_X4 _u0_u20_U361  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[15] ) );
INV_X4 _u0_u20_U359  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[14] ) );
INV_X4 _u0_u20_U357  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[13] ) );
INV_X4 _u0_u20_U355  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[12] ) );
INV_X4 _u0_u20_U353  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[11] ) );
INV_X4 _u0_u20_U351  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[10] ) );
INV_X4 _u0_u20_U349  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[9] ) );
INV_X4 _u0_u20_U347  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[8] ) );
INV_X4 _u0_u20_U345  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[7] ) );
INV_X4 _u0_u20_U343  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[6] ) );
INV_X4 _u0_u20_U341  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[5] ) );
INV_X4 _u0_u20_U339  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[4] ) );
INV_X4 _u0_u20_U337  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[3] ) );
INV_X4 _u0_u20_U335  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[2] ) );
INV_X4 _u0_u20_U333  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[1] ) );
INV_X4 _u0_u20_U331  ( .A(1'b1), .ZN(_u0_u20_ch_txsz[0] ) );
INV_X4 _u0_u20_U329  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[31] ) );
INV_X4 _u0_u20_U327  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[30] ) );
INV_X4 _u0_u20_U325  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[29] ) );
INV_X4 _u0_u20_U323  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[28] ) );
INV_X4 _u0_u20_U321  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[27] ) );
INV_X4 _u0_u20_U319  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[26] ) );
INV_X4 _u0_u20_U317  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[25] ) );
INV_X4 _u0_u20_U315  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[24] ) );
INV_X4 _u0_u20_U313  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[23] ) );
INV_X4 _u0_u20_U311  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[22] ) );
INV_X4 _u0_u20_U309  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[21] ) );
INV_X4 _u0_u20_U307  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[20] ) );
INV_X4 _u0_u20_U305  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[19] ) );
INV_X4 _u0_u20_U303  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[18] ) );
INV_X4 _u0_u20_U301  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[17] ) );
INV_X4 _u0_u20_U299  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[16] ) );
INV_X4 _u0_u20_U297  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[15] ) );
INV_X4 _u0_u20_U295  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[14] ) );
INV_X4 _u0_u20_U293  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[13] ) );
INV_X4 _u0_u20_U291  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[12] ) );
INV_X4 _u0_u20_U289  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[11] ) );
INV_X4 _u0_u20_U287  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[10] ) );
INV_X4 _u0_u20_U285  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[9] ) );
INV_X4 _u0_u20_U283  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[8] ) );
INV_X4 _u0_u20_U281  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[7] ) );
INV_X4 _u0_u20_U279  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[6] ) );
INV_X4 _u0_u20_U277  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[5] ) );
INV_X4 _u0_u20_U275  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[4] ) );
INV_X4 _u0_u20_U273  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[3] ) );
INV_X4 _u0_u20_U271  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[2] ) );
INV_X4 _u0_u20_U269  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[1] ) );
INV_X4 _u0_u20_U267  ( .A(1'b1), .ZN(_u0_u20_ch_adr0[0] ) );
INV_X4 _u0_u20_U265  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[31] ) );
INV_X4 _u0_u20_U263  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[30] ) );
INV_X4 _u0_u20_U261  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[29] ) );
INV_X4 _u0_u20_U259  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[28] ) );
INV_X4 _u0_u20_U257  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[27] ) );
INV_X4 _u0_u20_U255  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[26] ) );
INV_X4 _u0_u20_U253  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[25] ) );
INV_X4 _u0_u20_U251  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[24] ) );
INV_X4 _u0_u20_U249  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[23] ) );
INV_X4 _u0_u20_U247  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[22] ) );
INV_X4 _u0_u20_U245  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[21] ) );
INV_X4 _u0_u20_U243  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[20] ) );
INV_X4 _u0_u20_U241  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[19] ) );
INV_X4 _u0_u20_U239  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[18] ) );
INV_X4 _u0_u20_U237  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[17] ) );
INV_X4 _u0_u20_U235  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[16] ) );
INV_X4 _u0_u20_U233  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[15] ) );
INV_X4 _u0_u20_U231  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[14] ) );
INV_X4 _u0_u20_U229  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[13] ) );
INV_X4 _u0_u20_U227  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[12] ) );
INV_X4 _u0_u20_U225  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[11] ) );
INV_X4 _u0_u20_U223  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[10] ) );
INV_X4 _u0_u20_U221  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[9] ) );
INV_X4 _u0_u20_U219  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[8] ) );
INV_X4 _u0_u20_U217  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[7] ) );
INV_X4 _u0_u20_U215  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[6] ) );
INV_X4 _u0_u20_U213  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[5] ) );
INV_X4 _u0_u20_U211  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[4] ) );
INV_X4 _u0_u20_U209  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[3] ) );
INV_X4 _u0_u20_U207  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[2] ) );
INV_X4 _u0_u20_U205  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[1] ) );
INV_X4 _u0_u20_U203  ( .A(1'b1), .ZN(_u0_u20_ch_adr1[0] ) );
INV_X4 _u0_u20_U201  ( .A(1'b0), .ZN(_u0_u20_ch_am0[31] ) );
INV_X4 _u0_u20_U199  ( .A(1'b0), .ZN(_u0_u20_ch_am0[30] ) );
INV_X4 _u0_u20_U197  ( .A(1'b0), .ZN(_u0_u20_ch_am0[29] ) );
INV_X4 _u0_u20_U195  ( .A(1'b0), .ZN(_u0_u20_ch_am0[28] ) );
INV_X4 _u0_u20_U193  ( .A(1'b0), .ZN(_u0_u20_ch_am0[27] ) );
INV_X4 _u0_u20_U191  ( .A(1'b0), .ZN(_u0_u20_ch_am0[26] ) );
INV_X4 _u0_u20_U189  ( .A(1'b0), .ZN(_u0_u20_ch_am0[25] ) );
INV_X4 _u0_u20_U187  ( .A(1'b0), .ZN(_u0_u20_ch_am0[24] ) );
INV_X4 _u0_u20_U185  ( .A(1'b0), .ZN(_u0_u20_ch_am0[23] ) );
INV_X4 _u0_u20_U183  ( .A(1'b0), .ZN(_u0_u20_ch_am0[22] ) );
INV_X4 _u0_u20_U181  ( .A(1'b0), .ZN(_u0_u20_ch_am0[21] ) );
INV_X4 _u0_u20_U179  ( .A(1'b0), .ZN(_u0_u20_ch_am0[20] ) );
INV_X4 _u0_u20_U177  ( .A(1'b0), .ZN(_u0_u20_ch_am0[19] ) );
INV_X4 _u0_u20_U175  ( .A(1'b0), .ZN(_u0_u20_ch_am0[18] ) );
INV_X4 _u0_u20_U173  ( .A(1'b0), .ZN(_u0_u20_ch_am0[17] ) );
INV_X4 _u0_u20_U171  ( .A(1'b0), .ZN(_u0_u20_ch_am0[16] ) );
INV_X4 _u0_u20_U169  ( .A(1'b0), .ZN(_u0_u20_ch_am0[15] ) );
INV_X4 _u0_u20_U167  ( .A(1'b0), .ZN(_u0_u20_ch_am0[14] ) );
INV_X4 _u0_u20_U165  ( .A(1'b0), .ZN(_u0_u20_ch_am0[13] ) );
INV_X4 _u0_u20_U163  ( .A(1'b0), .ZN(_u0_u20_ch_am0[12] ) );
INV_X4 _u0_u20_U161  ( .A(1'b0), .ZN(_u0_u20_ch_am0[11] ) );
INV_X4 _u0_u20_U159  ( .A(1'b0), .ZN(_u0_u20_ch_am0[10] ) );
INV_X4 _u0_u20_U157  ( .A(1'b0), .ZN(_u0_u20_ch_am0[9] ) );
INV_X4 _u0_u20_U155  ( .A(1'b0), .ZN(_u0_u20_ch_am0[8] ) );
INV_X4 _u0_u20_U153  ( .A(1'b0), .ZN(_u0_u20_ch_am0[7] ) );
INV_X4 _u0_u20_U151  ( .A(1'b0), .ZN(_u0_u20_ch_am0[6] ) );
INV_X4 _u0_u20_U149  ( .A(1'b0), .ZN(_u0_u20_ch_am0[5] ) );
INV_X4 _u0_u20_U147  ( .A(1'b0), .ZN(_u0_u20_ch_am0[4] ) );
INV_X4 _u0_u20_U145  ( .A(1'b1), .ZN(_u0_u20_ch_am0[3] ) );
INV_X4 _u0_u20_U143  ( .A(1'b1), .ZN(_u0_u20_ch_am0[2] ) );
INV_X4 _u0_u20_U141  ( .A(1'b1), .ZN(_u0_u20_ch_am0[1] ) );
INV_X4 _u0_u20_U139  ( .A(1'b1), .ZN(_u0_u20_ch_am0[0] ) );
INV_X4 _u0_u20_U137  ( .A(1'b0), .ZN(_u0_u20_ch_am1[31] ) );
INV_X4 _u0_u20_U135  ( .A(1'b0), .ZN(_u0_u20_ch_am1[30] ) );
INV_X4 _u0_u20_U133  ( .A(1'b0), .ZN(_u0_u20_ch_am1[29] ) );
INV_X4 _u0_u20_U131  ( .A(1'b0), .ZN(_u0_u20_ch_am1[28] ) );
INV_X4 _u0_u20_U129  ( .A(1'b0), .ZN(_u0_u20_ch_am1[27] ) );
INV_X4 _u0_u20_U127  ( .A(1'b0), .ZN(_u0_u20_ch_am1[26] ) );
INV_X4 _u0_u20_U125  ( .A(1'b0), .ZN(_u0_u20_ch_am1[25] ) );
INV_X4 _u0_u20_U123  ( .A(1'b0), .ZN(_u0_u20_ch_am1[24] ) );
INV_X4 _u0_u20_U121  ( .A(1'b0), .ZN(_u0_u20_ch_am1[23] ) );
INV_X4 _u0_u20_U119  ( .A(1'b0), .ZN(_u0_u20_ch_am1[22] ) );
INV_X4 _u0_u20_U117  ( .A(1'b0), .ZN(_u0_u20_ch_am1[21] ) );
INV_X4 _u0_u20_U115  ( .A(1'b0), .ZN(_u0_u20_ch_am1[20] ) );
INV_X4 _u0_u20_U113  ( .A(1'b0), .ZN(_u0_u20_ch_am1[19] ) );
INV_X4 _u0_u20_U111  ( .A(1'b0), .ZN(_u0_u20_ch_am1[18] ) );
INV_X4 _u0_u20_U109  ( .A(1'b0), .ZN(_u0_u20_ch_am1[17] ) );
INV_X4 _u0_u20_U107  ( .A(1'b0), .ZN(_u0_u20_ch_am1[16] ) );
INV_X4 _u0_u20_U105  ( .A(1'b0), .ZN(_u0_u20_ch_am1[15] ) );
INV_X4 _u0_u20_U103  ( .A(1'b0), .ZN(_u0_u20_ch_am1[14] ) );
INV_X4 _u0_u20_U101  ( .A(1'b0), .ZN(_u0_u20_ch_am1[13] ) );
INV_X4 _u0_u20_U99  ( .A(1'b0), .ZN(_u0_u20_ch_am1[12] ) );
INV_X4 _u0_u20_U97  ( .A(1'b0), .ZN(_u0_u20_ch_am1[11] ) );
INV_X4 _u0_u20_U95  ( .A(1'b0), .ZN(_u0_u20_ch_am1[10] ) );
INV_X4 _u0_u20_U93  ( .A(1'b0), .ZN(_u0_u20_ch_am1[9] ) );
INV_X4 _u0_u20_U91  ( .A(1'b0), .ZN(_u0_u20_ch_am1[8] ) );
INV_X4 _u0_u20_U89  ( .A(1'b0), .ZN(_u0_u20_ch_am1[7] ) );
INV_X4 _u0_u20_U87  ( .A(1'b0), .ZN(_u0_u20_ch_am1[6] ) );
INV_X4 _u0_u20_U85  ( .A(1'b0), .ZN(_u0_u20_ch_am1[5] ) );
INV_X4 _u0_u20_U83  ( .A(1'b0), .ZN(_u0_u20_ch_am1[4] ) );
INV_X4 _u0_u20_U81  ( .A(1'b1), .ZN(_u0_u20_ch_am1[3] ) );
INV_X4 _u0_u20_U79  ( .A(1'b1), .ZN(_u0_u20_ch_am1[2] ) );
INV_X4 _u0_u20_U77  ( .A(1'b1), .ZN(_u0_u20_ch_am1[1] ) );
INV_X4 _u0_u20_U75  ( .A(1'b1), .ZN(_u0_u20_ch_am1[0] ) );
INV_X4 _u0_u20_U73  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[31] ) );
INV_X4 _u0_u20_U71  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[30] ) );
INV_X4 _u0_u20_U69  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[29] ) );
INV_X4 _u0_u20_U67  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[28] ) );
INV_X4 _u0_u20_U65  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[27] ) );
INV_X4 _u0_u20_U63  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[26] ) );
INV_X4 _u0_u20_U61  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[25] ) );
INV_X4 _u0_u20_U59  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[24] ) );
INV_X4 _u0_u20_U57  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[23] ) );
INV_X4 _u0_u20_U55  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[22] ) );
INV_X4 _u0_u20_U53  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[21] ) );
INV_X4 _u0_u20_U51  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[20] ) );
INV_X4 _u0_u20_U49  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[19] ) );
INV_X4 _u0_u20_U47  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[18] ) );
INV_X4 _u0_u20_U45  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[17] ) );
INV_X4 _u0_u20_U43  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[16] ) );
INV_X4 _u0_u20_U41  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[15] ) );
INV_X4 _u0_u20_U39  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[14] ) );
INV_X4 _u0_u20_U37  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[13] ) );
INV_X4 _u0_u20_U35  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[12] ) );
INV_X4 _u0_u20_U33  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[11] ) );
INV_X4 _u0_u20_U31  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[10] ) );
INV_X4 _u0_u20_U29  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[9] ) );
INV_X4 _u0_u20_U27  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[8] ) );
INV_X4 _u0_u20_U25  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[7] ) );
INV_X4 _u0_u20_U23  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[6] ) );
INV_X4 _u0_u20_U21  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[5] ) );
INV_X4 _u0_u20_U19  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[4] ) );
INV_X4 _u0_u20_U17  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[3] ) );
INV_X4 _u0_u20_U15  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[2] ) );
INV_X4 _u0_u20_U13  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[1] ) );
INV_X4 _u0_u20_U11  ( .A(1'b1), .ZN(_u0_u20_sw_pointer[0] ) );
INV_X4 _u0_u20_U9  ( .A(1'b1), .ZN(_u0_u20_ch_stop ) );
INV_X4 _u0_u20_U7  ( .A(1'b1), .ZN(_u0_u20_ch_dis ) );
INV_X4 _u0_u20_U5  ( .A(1'b1), .ZN(_u0_u20_int ) );
INV_X4 _u0_u21_U585  ( .A(1'b1), .ZN(_u0_u21_pointer[31] ) );
INV_X4 _u0_u21_U583  ( .A(1'b1), .ZN(_u0_u21_pointer[30] ) );
INV_X4 _u0_u21_U581  ( .A(1'b1), .ZN(_u0_u21_pointer[29] ) );
INV_X4 _u0_u21_U579  ( .A(1'b1), .ZN(_u0_u21_pointer[28] ) );
INV_X4 _u0_u21_U577  ( .A(1'b1), .ZN(_u0_u21_pointer[27] ) );
INV_X4 _u0_u21_U575  ( .A(1'b1), .ZN(_u0_u21_pointer[26] ) );
INV_X4 _u0_u21_U573  ( .A(1'b1), .ZN(_u0_u21_pointer[25] ) );
INV_X4 _u0_u21_U571  ( .A(1'b1), .ZN(_u0_u21_pointer[24] ) );
INV_X4 _u0_u21_U569  ( .A(1'b1), .ZN(_u0_u21_pointer[23] ) );
INV_X4 _u0_u21_U567  ( .A(1'b1), .ZN(_u0_u21_pointer[22] ) );
INV_X4 _u0_u21_U565  ( .A(1'b1), .ZN(_u0_u21_pointer[21] ) );
INV_X4 _u0_u21_U563  ( .A(1'b1), .ZN(_u0_u21_pointer[20] ) );
INV_X4 _u0_u21_U561  ( .A(1'b1), .ZN(_u0_u21_pointer[19] ) );
INV_X4 _u0_u21_U559  ( .A(1'b1), .ZN(_u0_u21_pointer[18] ) );
INV_X4 _u0_u21_U557  ( .A(1'b1), .ZN(_u0_u21_pointer[17] ) );
INV_X4 _u0_u21_U555  ( .A(1'b1), .ZN(_u0_u21_pointer[16] ) );
INV_X4 _u0_u21_U553  ( .A(1'b1), .ZN(_u0_u21_pointer[15] ) );
INV_X4 _u0_u21_U551  ( .A(1'b1), .ZN(_u0_u21_pointer[14] ) );
INV_X4 _u0_u21_U549  ( .A(1'b1), .ZN(_u0_u21_pointer[13] ) );
INV_X4 _u0_u21_U547  ( .A(1'b1), .ZN(_u0_u21_pointer[12] ) );
INV_X4 _u0_u21_U545  ( .A(1'b1), .ZN(_u0_u21_pointer[11] ) );
INV_X4 _u0_u21_U543  ( .A(1'b1), .ZN(_u0_u21_pointer[10] ) );
INV_X4 _u0_u21_U541  ( .A(1'b1), .ZN(_u0_u21_pointer[9] ) );
INV_X4 _u0_u21_U539  ( .A(1'b1), .ZN(_u0_u21_pointer[8] ) );
INV_X4 _u0_u21_U537  ( .A(1'b1), .ZN(_u0_u21_pointer[7] ) );
INV_X4 _u0_u21_U535  ( .A(1'b1), .ZN(_u0_u21_pointer[6] ) );
INV_X4 _u0_u21_U533  ( .A(1'b1), .ZN(_u0_u21_pointer[5] ) );
INV_X4 _u0_u21_U531  ( .A(1'b1), .ZN(_u0_u21_pointer[4] ) );
INV_X4 _u0_u21_U529  ( .A(1'b1), .ZN(_u0_u21_pointer[3] ) );
INV_X4 _u0_u21_U527  ( .A(1'b1), .ZN(_u0_u21_pointer[2] ) );
INV_X4 _u0_u21_U525  ( .A(1'b1), .ZN(_u0_u21_pointer[1] ) );
INV_X4 _u0_u21_U523  ( .A(1'b1), .ZN(_u0_u21_pointer[0] ) );
INV_X4 _u0_u21_U521  ( .A(1'b1), .ZN(_u0_u21_pointer_s[31] ) );
INV_X4 _u0_u21_U519  ( .A(1'b1), .ZN(_u0_u21_pointer_s[30] ) );
INV_X4 _u0_u21_U517  ( .A(1'b1), .ZN(_u0_u21_pointer_s[29] ) );
INV_X4 _u0_u21_U515  ( .A(1'b1), .ZN(_u0_u21_pointer_s[28] ) );
INV_X4 _u0_u21_U513  ( .A(1'b1), .ZN(_u0_u21_pointer_s[27] ) );
INV_X4 _u0_u21_U511  ( .A(1'b1), .ZN(_u0_u21_pointer_s[26] ) );
INV_X4 _u0_u21_U509  ( .A(1'b1), .ZN(_u0_u21_pointer_s[25] ) );
INV_X4 _u0_u21_U507  ( .A(1'b1), .ZN(_u0_u21_pointer_s[24] ) );
INV_X4 _u0_u21_U505  ( .A(1'b1), .ZN(_u0_u21_pointer_s[23] ) );
INV_X4 _u0_u21_U503  ( .A(1'b1), .ZN(_u0_u21_pointer_s[22] ) );
INV_X4 _u0_u21_U501  ( .A(1'b1), .ZN(_u0_u21_pointer_s[21] ) );
INV_X4 _u0_u21_U499  ( .A(1'b1), .ZN(_u0_u21_pointer_s[20] ) );
INV_X4 _u0_u21_U497  ( .A(1'b1), .ZN(_u0_u21_pointer_s[19] ) );
INV_X4 _u0_u21_U495  ( .A(1'b1), .ZN(_u0_u21_pointer_s[18] ) );
INV_X4 _u0_u21_U493  ( .A(1'b1), .ZN(_u0_u21_pointer_s[17] ) );
INV_X4 _u0_u21_U491  ( .A(1'b1), .ZN(_u0_u21_pointer_s[16] ) );
INV_X4 _u0_u21_U489  ( .A(1'b1), .ZN(_u0_u21_pointer_s[15] ) );
INV_X4 _u0_u21_U487  ( .A(1'b1), .ZN(_u0_u21_pointer_s[14] ) );
INV_X4 _u0_u21_U485  ( .A(1'b1), .ZN(_u0_u21_pointer_s[13] ) );
INV_X4 _u0_u21_U483  ( .A(1'b1), .ZN(_u0_u21_pointer_s[12] ) );
INV_X4 _u0_u21_U481  ( .A(1'b1), .ZN(_u0_u21_pointer_s[11] ) );
INV_X4 _u0_u21_U479  ( .A(1'b1), .ZN(_u0_u21_pointer_s[10] ) );
INV_X4 _u0_u21_U477  ( .A(1'b1), .ZN(_u0_u21_pointer_s[9] ) );
INV_X4 _u0_u21_U475  ( .A(1'b1), .ZN(_u0_u21_pointer_s[8] ) );
INV_X4 _u0_u21_U473  ( .A(1'b1), .ZN(_u0_u21_pointer_s[7] ) );
INV_X4 _u0_u21_U471  ( .A(1'b1), .ZN(_u0_u21_pointer_s[6] ) );
INV_X4 _u0_u21_U469  ( .A(1'b1), .ZN(_u0_u21_pointer_s[5] ) );
INV_X4 _u0_u21_U467  ( .A(1'b1), .ZN(_u0_u21_pointer_s[4] ) );
INV_X4 _u0_u21_U465  ( .A(1'b1), .ZN(_u0_u21_pointer_s[3] ) );
INV_X4 _u0_u21_U463  ( .A(1'b1), .ZN(_u0_u21_pointer_s[2] ) );
INV_X4 _u0_u21_U461  ( .A(1'b1), .ZN(_u0_u21_pointer_s[1] ) );
INV_X4 _u0_u21_U459  ( .A(1'b1), .ZN(_u0_u21_pointer_s[0] ) );
INV_X4 _u0_u21_U457  ( .A(1'b1), .ZN(_u0_u21_ch_csr[31] ) );
INV_X4 _u0_u21_U455  ( .A(1'b1), .ZN(_u0_u21_ch_csr[30] ) );
INV_X4 _u0_u21_U453  ( .A(1'b1), .ZN(_u0_u21_ch_csr[29] ) );
INV_X4 _u0_u21_U451  ( .A(1'b1), .ZN(_u0_u21_ch_csr[28] ) );
INV_X4 _u0_u21_U449  ( .A(1'b1), .ZN(_u0_u21_ch_csr[27] ) );
INV_X4 _u0_u21_U447  ( .A(1'b1), .ZN(_u0_u21_ch_csr[26] ) );
INV_X4 _u0_u21_U445  ( .A(1'b1), .ZN(_u0_u21_ch_csr[25] ) );
INV_X4 _u0_u21_U443  ( .A(1'b1), .ZN(_u0_u21_ch_csr[24] ) );
INV_X4 _u0_u21_U441  ( .A(1'b1), .ZN(_u0_u21_ch_csr[23] ) );
INV_X4 _u0_u21_U439  ( .A(1'b1), .ZN(_u0_u21_ch_csr[22] ) );
INV_X4 _u0_u21_U437  ( .A(1'b1), .ZN(_u0_u21_ch_csr[21] ) );
INV_X4 _u0_u21_U435  ( .A(1'b1), .ZN(_u0_u21_ch_csr[20] ) );
INV_X4 _u0_u21_U433  ( .A(1'b1), .ZN(_u0_u21_ch_csr[19] ) );
INV_X4 _u0_u21_U431  ( .A(1'b1), .ZN(_u0_u21_ch_csr[18] ) );
INV_X4 _u0_u21_U429  ( .A(1'b1), .ZN(_u0_u21_ch_csr[17] ) );
INV_X4 _u0_u21_U427  ( .A(1'b1), .ZN(_u0_u21_ch_csr[16] ) );
INV_X4 _u0_u21_U425  ( .A(1'b1), .ZN(_u0_u21_ch_csr[15] ) );
INV_X4 _u0_u21_U423  ( .A(1'b1), .ZN(_u0_u21_ch_csr[14] ) );
INV_X4 _u0_u21_U421  ( .A(1'b1), .ZN(_u0_u21_ch_csr[13] ) );
INV_X4 _u0_u21_U419  ( .A(1'b1), .ZN(_u0_u21_ch_csr[12] ) );
INV_X4 _u0_u21_U417  ( .A(1'b1), .ZN(_u0_u21_ch_csr[11] ) );
INV_X4 _u0_u21_U415  ( .A(1'b1), .ZN(_u0_u21_ch_csr[10] ) );
INV_X4 _u0_u21_U413  ( .A(1'b1), .ZN(_u0_u21_ch_csr[9] ) );
INV_X4 _u0_u21_U411  ( .A(1'b1), .ZN(_u0_u21_ch_csr[8] ) );
INV_X4 _u0_u21_U409  ( .A(1'b1), .ZN(_u0_u21_ch_csr[7] ) );
INV_X4 _u0_u21_U407  ( .A(1'b1), .ZN(_u0_u21_ch_csr[6] ) );
INV_X4 _u0_u21_U405  ( .A(1'b1), .ZN(_u0_u21_ch_csr[5] ) );
INV_X4 _u0_u21_U403  ( .A(1'b1), .ZN(_u0_u21_ch_csr[4] ) );
INV_X4 _u0_u21_U401  ( .A(1'b1), .ZN(_u0_u21_ch_csr[3] ) );
INV_X4 _u0_u21_U399  ( .A(1'b1), .ZN(_u0_u21_ch_csr[2] ) );
INV_X4 _u0_u21_U397  ( .A(1'b1), .ZN(_u0_u21_ch_csr[1] ) );
INV_X4 _u0_u21_U395  ( .A(1'b1), .ZN(_u0_u21_ch_csr[0] ) );
INV_X4 _u0_u21_U393  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[31] ) );
INV_X4 _u0_u21_U391  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[30] ) );
INV_X4 _u0_u21_U389  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[29] ) );
INV_X4 _u0_u21_U387  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[28] ) );
INV_X4 _u0_u21_U385  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[27] ) );
INV_X4 _u0_u21_U383  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[26] ) );
INV_X4 _u0_u21_U381  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[25] ) );
INV_X4 _u0_u21_U379  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[24] ) );
INV_X4 _u0_u21_U377  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[23] ) );
INV_X4 _u0_u21_U375  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[22] ) );
INV_X4 _u0_u21_U373  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[21] ) );
INV_X4 _u0_u21_U371  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[20] ) );
INV_X4 _u0_u21_U369  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[19] ) );
INV_X4 _u0_u21_U367  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[18] ) );
INV_X4 _u0_u21_U365  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[17] ) );
INV_X4 _u0_u21_U363  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[16] ) );
INV_X4 _u0_u21_U361  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[15] ) );
INV_X4 _u0_u21_U359  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[14] ) );
INV_X4 _u0_u21_U357  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[13] ) );
INV_X4 _u0_u21_U355  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[12] ) );
INV_X4 _u0_u21_U353  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[11] ) );
INV_X4 _u0_u21_U351  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[10] ) );
INV_X4 _u0_u21_U349  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[9] ) );
INV_X4 _u0_u21_U347  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[8] ) );
INV_X4 _u0_u21_U345  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[7] ) );
INV_X4 _u0_u21_U343  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[6] ) );
INV_X4 _u0_u21_U341  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[5] ) );
INV_X4 _u0_u21_U339  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[4] ) );
INV_X4 _u0_u21_U337  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[3] ) );
INV_X4 _u0_u21_U335  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[2] ) );
INV_X4 _u0_u21_U333  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[1] ) );
INV_X4 _u0_u21_U331  ( .A(1'b1), .ZN(_u0_u21_ch_txsz[0] ) );
INV_X4 _u0_u21_U329  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[31] ) );
INV_X4 _u0_u21_U327  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[30] ) );
INV_X4 _u0_u21_U325  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[29] ) );
INV_X4 _u0_u21_U323  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[28] ) );
INV_X4 _u0_u21_U321  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[27] ) );
INV_X4 _u0_u21_U319  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[26] ) );
INV_X4 _u0_u21_U317  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[25] ) );
INV_X4 _u0_u21_U315  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[24] ) );
INV_X4 _u0_u21_U313  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[23] ) );
INV_X4 _u0_u21_U311  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[22] ) );
INV_X4 _u0_u21_U309  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[21] ) );
INV_X4 _u0_u21_U307  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[20] ) );
INV_X4 _u0_u21_U305  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[19] ) );
INV_X4 _u0_u21_U303  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[18] ) );
INV_X4 _u0_u21_U301  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[17] ) );
INV_X4 _u0_u21_U299  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[16] ) );
INV_X4 _u0_u21_U297  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[15] ) );
INV_X4 _u0_u21_U295  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[14] ) );
INV_X4 _u0_u21_U293  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[13] ) );
INV_X4 _u0_u21_U291  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[12] ) );
INV_X4 _u0_u21_U289  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[11] ) );
INV_X4 _u0_u21_U287  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[10] ) );
INV_X4 _u0_u21_U285  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[9] ) );
INV_X4 _u0_u21_U283  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[8] ) );
INV_X4 _u0_u21_U281  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[7] ) );
INV_X4 _u0_u21_U279  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[6] ) );
INV_X4 _u0_u21_U277  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[5] ) );
INV_X4 _u0_u21_U275  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[4] ) );
INV_X4 _u0_u21_U273  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[3] ) );
INV_X4 _u0_u21_U271  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[2] ) );
INV_X4 _u0_u21_U269  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[1] ) );
INV_X4 _u0_u21_U267  ( .A(1'b1), .ZN(_u0_u21_ch_adr0[0] ) );
INV_X4 _u0_u21_U265  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[31] ) );
INV_X4 _u0_u21_U263  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[30] ) );
INV_X4 _u0_u21_U261  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[29] ) );
INV_X4 _u0_u21_U259  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[28] ) );
INV_X4 _u0_u21_U257  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[27] ) );
INV_X4 _u0_u21_U255  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[26] ) );
INV_X4 _u0_u21_U253  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[25] ) );
INV_X4 _u0_u21_U251  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[24] ) );
INV_X4 _u0_u21_U249  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[23] ) );
INV_X4 _u0_u21_U247  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[22] ) );
INV_X4 _u0_u21_U245  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[21] ) );
INV_X4 _u0_u21_U243  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[20] ) );
INV_X4 _u0_u21_U241  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[19] ) );
INV_X4 _u0_u21_U239  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[18] ) );
INV_X4 _u0_u21_U237  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[17] ) );
INV_X4 _u0_u21_U235  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[16] ) );
INV_X4 _u0_u21_U233  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[15] ) );
INV_X4 _u0_u21_U231  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[14] ) );
INV_X4 _u0_u21_U229  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[13] ) );
INV_X4 _u0_u21_U227  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[12] ) );
INV_X4 _u0_u21_U225  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[11] ) );
INV_X4 _u0_u21_U223  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[10] ) );
INV_X4 _u0_u21_U221  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[9] ) );
INV_X4 _u0_u21_U219  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[8] ) );
INV_X4 _u0_u21_U217  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[7] ) );
INV_X4 _u0_u21_U215  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[6] ) );
INV_X4 _u0_u21_U213  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[5] ) );
INV_X4 _u0_u21_U211  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[4] ) );
INV_X4 _u0_u21_U209  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[3] ) );
INV_X4 _u0_u21_U207  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[2] ) );
INV_X4 _u0_u21_U205  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[1] ) );
INV_X4 _u0_u21_U203  ( .A(1'b1), .ZN(_u0_u21_ch_adr1[0] ) );
INV_X4 _u0_u21_U201  ( .A(1'b0), .ZN(_u0_u21_ch_am0[31] ) );
INV_X4 _u0_u21_U199  ( .A(1'b0), .ZN(_u0_u21_ch_am0[30] ) );
INV_X4 _u0_u21_U197  ( .A(1'b0), .ZN(_u0_u21_ch_am0[29] ) );
INV_X4 _u0_u21_U195  ( .A(1'b0), .ZN(_u0_u21_ch_am0[28] ) );
INV_X4 _u0_u21_U193  ( .A(1'b0), .ZN(_u0_u21_ch_am0[27] ) );
INV_X4 _u0_u21_U191  ( .A(1'b0), .ZN(_u0_u21_ch_am0[26] ) );
INV_X4 _u0_u21_U189  ( .A(1'b0), .ZN(_u0_u21_ch_am0[25] ) );
INV_X4 _u0_u21_U187  ( .A(1'b0), .ZN(_u0_u21_ch_am0[24] ) );
INV_X4 _u0_u21_U185  ( .A(1'b0), .ZN(_u0_u21_ch_am0[23] ) );
INV_X4 _u0_u21_U183  ( .A(1'b0), .ZN(_u0_u21_ch_am0[22] ) );
INV_X4 _u0_u21_U181  ( .A(1'b0), .ZN(_u0_u21_ch_am0[21] ) );
INV_X4 _u0_u21_U179  ( .A(1'b0), .ZN(_u0_u21_ch_am0[20] ) );
INV_X4 _u0_u21_U177  ( .A(1'b0), .ZN(_u0_u21_ch_am0[19] ) );
INV_X4 _u0_u21_U175  ( .A(1'b0), .ZN(_u0_u21_ch_am0[18] ) );
INV_X4 _u0_u21_U173  ( .A(1'b0), .ZN(_u0_u21_ch_am0[17] ) );
INV_X4 _u0_u21_U171  ( .A(1'b0), .ZN(_u0_u21_ch_am0[16] ) );
INV_X4 _u0_u21_U169  ( .A(1'b0), .ZN(_u0_u21_ch_am0[15] ) );
INV_X4 _u0_u21_U167  ( .A(1'b0), .ZN(_u0_u21_ch_am0[14] ) );
INV_X4 _u0_u21_U165  ( .A(1'b0), .ZN(_u0_u21_ch_am0[13] ) );
INV_X4 _u0_u21_U163  ( .A(1'b0), .ZN(_u0_u21_ch_am0[12] ) );
INV_X4 _u0_u21_U161  ( .A(1'b0), .ZN(_u0_u21_ch_am0[11] ) );
INV_X4 _u0_u21_U159  ( .A(1'b0), .ZN(_u0_u21_ch_am0[10] ) );
INV_X4 _u0_u21_U157  ( .A(1'b0), .ZN(_u0_u21_ch_am0[9] ) );
INV_X4 _u0_u21_U155  ( .A(1'b0), .ZN(_u0_u21_ch_am0[8] ) );
INV_X4 _u0_u21_U153  ( .A(1'b0), .ZN(_u0_u21_ch_am0[7] ) );
INV_X4 _u0_u21_U151  ( .A(1'b0), .ZN(_u0_u21_ch_am0[6] ) );
INV_X4 _u0_u21_U149  ( .A(1'b0), .ZN(_u0_u21_ch_am0[5] ) );
INV_X4 _u0_u21_U147  ( .A(1'b0), .ZN(_u0_u21_ch_am0[4] ) );
INV_X4 _u0_u21_U145  ( .A(1'b1), .ZN(_u0_u21_ch_am0[3] ) );
INV_X4 _u0_u21_U143  ( .A(1'b1), .ZN(_u0_u21_ch_am0[2] ) );
INV_X4 _u0_u21_U141  ( .A(1'b1), .ZN(_u0_u21_ch_am0[1] ) );
INV_X4 _u0_u21_U139  ( .A(1'b1), .ZN(_u0_u21_ch_am0[0] ) );
INV_X4 _u0_u21_U137  ( .A(1'b0), .ZN(_u0_u21_ch_am1[31] ) );
INV_X4 _u0_u21_U135  ( .A(1'b0), .ZN(_u0_u21_ch_am1[30] ) );
INV_X4 _u0_u21_U133  ( .A(1'b0), .ZN(_u0_u21_ch_am1[29] ) );
INV_X4 _u0_u21_U131  ( .A(1'b0), .ZN(_u0_u21_ch_am1[28] ) );
INV_X4 _u0_u21_U129  ( .A(1'b0), .ZN(_u0_u21_ch_am1[27] ) );
INV_X4 _u0_u21_U127  ( .A(1'b0), .ZN(_u0_u21_ch_am1[26] ) );
INV_X4 _u0_u21_U125  ( .A(1'b0), .ZN(_u0_u21_ch_am1[25] ) );
INV_X4 _u0_u21_U123  ( .A(1'b0), .ZN(_u0_u21_ch_am1[24] ) );
INV_X4 _u0_u21_U121  ( .A(1'b0), .ZN(_u0_u21_ch_am1[23] ) );
INV_X4 _u0_u21_U119  ( .A(1'b0), .ZN(_u0_u21_ch_am1[22] ) );
INV_X4 _u0_u21_U117  ( .A(1'b0), .ZN(_u0_u21_ch_am1[21] ) );
INV_X4 _u0_u21_U115  ( .A(1'b0), .ZN(_u0_u21_ch_am1[20] ) );
INV_X4 _u0_u21_U113  ( .A(1'b0), .ZN(_u0_u21_ch_am1[19] ) );
INV_X4 _u0_u21_U111  ( .A(1'b0), .ZN(_u0_u21_ch_am1[18] ) );
INV_X4 _u0_u21_U109  ( .A(1'b0), .ZN(_u0_u21_ch_am1[17] ) );
INV_X4 _u0_u21_U107  ( .A(1'b0), .ZN(_u0_u21_ch_am1[16] ) );
INV_X4 _u0_u21_U105  ( .A(1'b0), .ZN(_u0_u21_ch_am1[15] ) );
INV_X4 _u0_u21_U103  ( .A(1'b0), .ZN(_u0_u21_ch_am1[14] ) );
INV_X4 _u0_u21_U101  ( .A(1'b0), .ZN(_u0_u21_ch_am1[13] ) );
INV_X4 _u0_u21_U99  ( .A(1'b0), .ZN(_u0_u21_ch_am1[12] ) );
INV_X4 _u0_u21_U97  ( .A(1'b0), .ZN(_u0_u21_ch_am1[11] ) );
INV_X4 _u0_u21_U95  ( .A(1'b0), .ZN(_u0_u21_ch_am1[10] ) );
INV_X4 _u0_u21_U93  ( .A(1'b0), .ZN(_u0_u21_ch_am1[9] ) );
INV_X4 _u0_u21_U91  ( .A(1'b0), .ZN(_u0_u21_ch_am1[8] ) );
INV_X4 _u0_u21_U89  ( .A(1'b0), .ZN(_u0_u21_ch_am1[7] ) );
INV_X4 _u0_u21_U87  ( .A(1'b0), .ZN(_u0_u21_ch_am1[6] ) );
INV_X4 _u0_u21_U85  ( .A(1'b0), .ZN(_u0_u21_ch_am1[5] ) );
INV_X4 _u0_u21_U83  ( .A(1'b0), .ZN(_u0_u21_ch_am1[4] ) );
INV_X4 _u0_u21_U81  ( .A(1'b1), .ZN(_u0_u21_ch_am1[3] ) );
INV_X4 _u0_u21_U79  ( .A(1'b1), .ZN(_u0_u21_ch_am1[2] ) );
INV_X4 _u0_u21_U77  ( .A(1'b1), .ZN(_u0_u21_ch_am1[1] ) );
INV_X4 _u0_u21_U75  ( .A(1'b1), .ZN(_u0_u21_ch_am1[0] ) );
INV_X4 _u0_u21_U73  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[31] ) );
INV_X4 _u0_u21_U71  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[30] ) );
INV_X4 _u0_u21_U69  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[29] ) );
INV_X4 _u0_u21_U67  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[28] ) );
INV_X4 _u0_u21_U65  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[27] ) );
INV_X4 _u0_u21_U63  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[26] ) );
INV_X4 _u0_u21_U61  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[25] ) );
INV_X4 _u0_u21_U59  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[24] ) );
INV_X4 _u0_u21_U57  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[23] ) );
INV_X4 _u0_u21_U55  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[22] ) );
INV_X4 _u0_u21_U53  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[21] ) );
INV_X4 _u0_u21_U51  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[20] ) );
INV_X4 _u0_u21_U49  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[19] ) );
INV_X4 _u0_u21_U47  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[18] ) );
INV_X4 _u0_u21_U45  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[17] ) );
INV_X4 _u0_u21_U43  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[16] ) );
INV_X4 _u0_u21_U41  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[15] ) );
INV_X4 _u0_u21_U39  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[14] ) );
INV_X4 _u0_u21_U37  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[13] ) );
INV_X4 _u0_u21_U35  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[12] ) );
INV_X4 _u0_u21_U33  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[11] ) );
INV_X4 _u0_u21_U31  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[10] ) );
INV_X4 _u0_u21_U29  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[9] ) );
INV_X4 _u0_u21_U27  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[8] ) );
INV_X4 _u0_u21_U25  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[7] ) );
INV_X4 _u0_u21_U23  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[6] ) );
INV_X4 _u0_u21_U21  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[5] ) );
INV_X4 _u0_u21_U19  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[4] ) );
INV_X4 _u0_u21_U17  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[3] ) );
INV_X4 _u0_u21_U15  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[2] ) );
INV_X4 _u0_u21_U13  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[1] ) );
INV_X4 _u0_u21_U11  ( .A(1'b1), .ZN(_u0_u21_sw_pointer[0] ) );
INV_X4 _u0_u21_U9  ( .A(1'b1), .ZN(_u0_u21_ch_stop ) );
INV_X4 _u0_u21_U7  ( .A(1'b1), .ZN(_u0_u21_ch_dis ) );
INV_X4 _u0_u21_U5  ( .A(1'b1), .ZN(_u0_u21_int ) );
INV_X4 _u0_u22_U585  ( .A(1'b1), .ZN(_u0_u22_pointer[31] ) );
INV_X4 _u0_u22_U583  ( .A(1'b1), .ZN(_u0_u22_pointer[30] ) );
INV_X4 _u0_u22_U581  ( .A(1'b1), .ZN(_u0_u22_pointer[29] ) );
INV_X4 _u0_u22_U579  ( .A(1'b1), .ZN(_u0_u22_pointer[28] ) );
INV_X4 _u0_u22_U577  ( .A(1'b1), .ZN(_u0_u22_pointer[27] ) );
INV_X4 _u0_u22_U575  ( .A(1'b1), .ZN(_u0_u22_pointer[26] ) );
INV_X4 _u0_u22_U573  ( .A(1'b1), .ZN(_u0_u22_pointer[25] ) );
INV_X4 _u0_u22_U571  ( .A(1'b1), .ZN(_u0_u22_pointer[24] ) );
INV_X4 _u0_u22_U569  ( .A(1'b1), .ZN(_u0_u22_pointer[23] ) );
INV_X4 _u0_u22_U567  ( .A(1'b1), .ZN(_u0_u22_pointer[22] ) );
INV_X4 _u0_u22_U565  ( .A(1'b1), .ZN(_u0_u22_pointer[21] ) );
INV_X4 _u0_u22_U563  ( .A(1'b1), .ZN(_u0_u22_pointer[20] ) );
INV_X4 _u0_u22_U561  ( .A(1'b1), .ZN(_u0_u22_pointer[19] ) );
INV_X4 _u0_u22_U559  ( .A(1'b1), .ZN(_u0_u22_pointer[18] ) );
INV_X4 _u0_u22_U557  ( .A(1'b1), .ZN(_u0_u22_pointer[17] ) );
INV_X4 _u0_u22_U555  ( .A(1'b1), .ZN(_u0_u22_pointer[16] ) );
INV_X4 _u0_u22_U553  ( .A(1'b1), .ZN(_u0_u22_pointer[15] ) );
INV_X4 _u0_u22_U551  ( .A(1'b1), .ZN(_u0_u22_pointer[14] ) );
INV_X4 _u0_u22_U549  ( .A(1'b1), .ZN(_u0_u22_pointer[13] ) );
INV_X4 _u0_u22_U547  ( .A(1'b1), .ZN(_u0_u22_pointer[12] ) );
INV_X4 _u0_u22_U545  ( .A(1'b1), .ZN(_u0_u22_pointer[11] ) );
INV_X4 _u0_u22_U543  ( .A(1'b1), .ZN(_u0_u22_pointer[10] ) );
INV_X4 _u0_u22_U541  ( .A(1'b1), .ZN(_u0_u22_pointer[9] ) );
INV_X4 _u0_u22_U539  ( .A(1'b1), .ZN(_u0_u22_pointer[8] ) );
INV_X4 _u0_u22_U537  ( .A(1'b1), .ZN(_u0_u22_pointer[7] ) );
INV_X4 _u0_u22_U535  ( .A(1'b1), .ZN(_u0_u22_pointer[6] ) );
INV_X4 _u0_u22_U533  ( .A(1'b1), .ZN(_u0_u22_pointer[5] ) );
INV_X4 _u0_u22_U531  ( .A(1'b1), .ZN(_u0_u22_pointer[4] ) );
INV_X4 _u0_u22_U529  ( .A(1'b1), .ZN(_u0_u22_pointer[3] ) );
INV_X4 _u0_u22_U527  ( .A(1'b1), .ZN(_u0_u22_pointer[2] ) );
INV_X4 _u0_u22_U525  ( .A(1'b1), .ZN(_u0_u22_pointer[1] ) );
INV_X4 _u0_u22_U523  ( .A(1'b1), .ZN(_u0_u22_pointer[0] ) );
INV_X4 _u0_u22_U521  ( .A(1'b1), .ZN(_u0_u22_pointer_s[31] ) );
INV_X4 _u0_u22_U519  ( .A(1'b1), .ZN(_u0_u22_pointer_s[30] ) );
INV_X4 _u0_u22_U517  ( .A(1'b1), .ZN(_u0_u22_pointer_s[29] ) );
INV_X4 _u0_u22_U515  ( .A(1'b1), .ZN(_u0_u22_pointer_s[28] ) );
INV_X4 _u0_u22_U513  ( .A(1'b1), .ZN(_u0_u22_pointer_s[27] ) );
INV_X4 _u0_u22_U511  ( .A(1'b1), .ZN(_u0_u22_pointer_s[26] ) );
INV_X4 _u0_u22_U509  ( .A(1'b1), .ZN(_u0_u22_pointer_s[25] ) );
INV_X4 _u0_u22_U507  ( .A(1'b1), .ZN(_u0_u22_pointer_s[24] ) );
INV_X4 _u0_u22_U505  ( .A(1'b1), .ZN(_u0_u22_pointer_s[23] ) );
INV_X4 _u0_u22_U503  ( .A(1'b1), .ZN(_u0_u22_pointer_s[22] ) );
INV_X4 _u0_u22_U501  ( .A(1'b1), .ZN(_u0_u22_pointer_s[21] ) );
INV_X4 _u0_u22_U499  ( .A(1'b1), .ZN(_u0_u22_pointer_s[20] ) );
INV_X4 _u0_u22_U497  ( .A(1'b1), .ZN(_u0_u22_pointer_s[19] ) );
INV_X4 _u0_u22_U495  ( .A(1'b1), .ZN(_u0_u22_pointer_s[18] ) );
INV_X4 _u0_u22_U493  ( .A(1'b1), .ZN(_u0_u22_pointer_s[17] ) );
INV_X4 _u0_u22_U491  ( .A(1'b1), .ZN(_u0_u22_pointer_s[16] ) );
INV_X4 _u0_u22_U489  ( .A(1'b1), .ZN(_u0_u22_pointer_s[15] ) );
INV_X4 _u0_u22_U487  ( .A(1'b1), .ZN(_u0_u22_pointer_s[14] ) );
INV_X4 _u0_u22_U485  ( .A(1'b1), .ZN(_u0_u22_pointer_s[13] ) );
INV_X4 _u0_u22_U483  ( .A(1'b1), .ZN(_u0_u22_pointer_s[12] ) );
INV_X4 _u0_u22_U481  ( .A(1'b1), .ZN(_u0_u22_pointer_s[11] ) );
INV_X4 _u0_u22_U479  ( .A(1'b1), .ZN(_u0_u22_pointer_s[10] ) );
INV_X4 _u0_u22_U477  ( .A(1'b1), .ZN(_u0_u22_pointer_s[9] ) );
INV_X4 _u0_u22_U475  ( .A(1'b1), .ZN(_u0_u22_pointer_s[8] ) );
INV_X4 _u0_u22_U473  ( .A(1'b1), .ZN(_u0_u22_pointer_s[7] ) );
INV_X4 _u0_u22_U471  ( .A(1'b1), .ZN(_u0_u22_pointer_s[6] ) );
INV_X4 _u0_u22_U469  ( .A(1'b1), .ZN(_u0_u22_pointer_s[5] ) );
INV_X4 _u0_u22_U467  ( .A(1'b1), .ZN(_u0_u22_pointer_s[4] ) );
INV_X4 _u0_u22_U465  ( .A(1'b1), .ZN(_u0_u22_pointer_s[3] ) );
INV_X4 _u0_u22_U463  ( .A(1'b1), .ZN(_u0_u22_pointer_s[2] ) );
INV_X4 _u0_u22_U461  ( .A(1'b1), .ZN(_u0_u22_pointer_s[1] ) );
INV_X4 _u0_u22_U459  ( .A(1'b1), .ZN(_u0_u22_pointer_s[0] ) );
INV_X4 _u0_u22_U457  ( .A(1'b1), .ZN(_u0_u22_ch_csr[31] ) );
INV_X4 _u0_u22_U455  ( .A(1'b1), .ZN(_u0_u22_ch_csr[30] ) );
INV_X4 _u0_u22_U453  ( .A(1'b1), .ZN(_u0_u22_ch_csr[29] ) );
INV_X4 _u0_u22_U451  ( .A(1'b1), .ZN(_u0_u22_ch_csr[28] ) );
INV_X4 _u0_u22_U449  ( .A(1'b1), .ZN(_u0_u22_ch_csr[27] ) );
INV_X4 _u0_u22_U447  ( .A(1'b1), .ZN(_u0_u22_ch_csr[26] ) );
INV_X4 _u0_u22_U445  ( .A(1'b1), .ZN(_u0_u22_ch_csr[25] ) );
INV_X4 _u0_u22_U443  ( .A(1'b1), .ZN(_u0_u22_ch_csr[24] ) );
INV_X4 _u0_u22_U441  ( .A(1'b1), .ZN(_u0_u22_ch_csr[23] ) );
INV_X4 _u0_u22_U439  ( .A(1'b1), .ZN(_u0_u22_ch_csr[22] ) );
INV_X4 _u0_u22_U437  ( .A(1'b1), .ZN(_u0_u22_ch_csr[21] ) );
INV_X4 _u0_u22_U435  ( .A(1'b1), .ZN(_u0_u22_ch_csr[20] ) );
INV_X4 _u0_u22_U433  ( .A(1'b1), .ZN(_u0_u22_ch_csr[19] ) );
INV_X4 _u0_u22_U431  ( .A(1'b1), .ZN(_u0_u22_ch_csr[18] ) );
INV_X4 _u0_u22_U429  ( .A(1'b1), .ZN(_u0_u22_ch_csr[17] ) );
INV_X4 _u0_u22_U427  ( .A(1'b1), .ZN(_u0_u22_ch_csr[16] ) );
INV_X4 _u0_u22_U425  ( .A(1'b1), .ZN(_u0_u22_ch_csr[15] ) );
INV_X4 _u0_u22_U423  ( .A(1'b1), .ZN(_u0_u22_ch_csr[14] ) );
INV_X4 _u0_u22_U421  ( .A(1'b1), .ZN(_u0_u22_ch_csr[13] ) );
INV_X4 _u0_u22_U419  ( .A(1'b1), .ZN(_u0_u22_ch_csr[12] ) );
INV_X4 _u0_u22_U417  ( .A(1'b1), .ZN(_u0_u22_ch_csr[11] ) );
INV_X4 _u0_u22_U415  ( .A(1'b1), .ZN(_u0_u22_ch_csr[10] ) );
INV_X4 _u0_u22_U413  ( .A(1'b1), .ZN(_u0_u22_ch_csr[9] ) );
INV_X4 _u0_u22_U411  ( .A(1'b1), .ZN(_u0_u22_ch_csr[8] ) );
INV_X4 _u0_u22_U409  ( .A(1'b1), .ZN(_u0_u22_ch_csr[7] ) );
INV_X4 _u0_u22_U407  ( .A(1'b1), .ZN(_u0_u22_ch_csr[6] ) );
INV_X4 _u0_u22_U405  ( .A(1'b1), .ZN(_u0_u22_ch_csr[5] ) );
INV_X4 _u0_u22_U403  ( .A(1'b1), .ZN(_u0_u22_ch_csr[4] ) );
INV_X4 _u0_u22_U401  ( .A(1'b1), .ZN(_u0_u22_ch_csr[3] ) );
INV_X4 _u0_u22_U399  ( .A(1'b1), .ZN(_u0_u22_ch_csr[2] ) );
INV_X4 _u0_u22_U397  ( .A(1'b1), .ZN(_u0_u22_ch_csr[1] ) );
INV_X4 _u0_u22_U395  ( .A(1'b1), .ZN(_u0_u22_ch_csr[0] ) );
INV_X4 _u0_u22_U393  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[31] ) );
INV_X4 _u0_u22_U391  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[30] ) );
INV_X4 _u0_u22_U389  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[29] ) );
INV_X4 _u0_u22_U387  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[28] ) );
INV_X4 _u0_u22_U385  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[27] ) );
INV_X4 _u0_u22_U383  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[26] ) );
INV_X4 _u0_u22_U381  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[25] ) );
INV_X4 _u0_u22_U379  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[24] ) );
INV_X4 _u0_u22_U377  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[23] ) );
INV_X4 _u0_u22_U375  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[22] ) );
INV_X4 _u0_u22_U373  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[21] ) );
INV_X4 _u0_u22_U371  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[20] ) );
INV_X4 _u0_u22_U369  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[19] ) );
INV_X4 _u0_u22_U367  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[18] ) );
INV_X4 _u0_u22_U365  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[17] ) );
INV_X4 _u0_u22_U363  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[16] ) );
INV_X4 _u0_u22_U361  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[15] ) );
INV_X4 _u0_u22_U359  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[14] ) );
INV_X4 _u0_u22_U357  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[13] ) );
INV_X4 _u0_u22_U355  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[12] ) );
INV_X4 _u0_u22_U353  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[11] ) );
INV_X4 _u0_u22_U351  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[10] ) );
INV_X4 _u0_u22_U349  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[9] ) );
INV_X4 _u0_u22_U347  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[8] ) );
INV_X4 _u0_u22_U345  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[7] ) );
INV_X4 _u0_u22_U343  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[6] ) );
INV_X4 _u0_u22_U341  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[5] ) );
INV_X4 _u0_u22_U339  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[4] ) );
INV_X4 _u0_u22_U337  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[3] ) );
INV_X4 _u0_u22_U335  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[2] ) );
INV_X4 _u0_u22_U333  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[1] ) );
INV_X4 _u0_u22_U331  ( .A(1'b1), .ZN(_u0_u22_ch_txsz[0] ) );
INV_X4 _u0_u22_U329  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[31] ) );
INV_X4 _u0_u22_U327  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[30] ) );
INV_X4 _u0_u22_U325  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[29] ) );
INV_X4 _u0_u22_U323  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[28] ) );
INV_X4 _u0_u22_U321  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[27] ) );
INV_X4 _u0_u22_U319  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[26] ) );
INV_X4 _u0_u22_U317  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[25] ) );
INV_X4 _u0_u22_U315  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[24] ) );
INV_X4 _u0_u22_U313  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[23] ) );
INV_X4 _u0_u22_U311  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[22] ) );
INV_X4 _u0_u22_U309  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[21] ) );
INV_X4 _u0_u22_U307  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[20] ) );
INV_X4 _u0_u22_U305  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[19] ) );
INV_X4 _u0_u22_U303  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[18] ) );
INV_X4 _u0_u22_U301  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[17] ) );
INV_X4 _u0_u22_U299  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[16] ) );
INV_X4 _u0_u22_U297  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[15] ) );
INV_X4 _u0_u22_U295  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[14] ) );
INV_X4 _u0_u22_U293  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[13] ) );
INV_X4 _u0_u22_U291  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[12] ) );
INV_X4 _u0_u22_U289  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[11] ) );
INV_X4 _u0_u22_U287  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[10] ) );
INV_X4 _u0_u22_U285  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[9] ) );
INV_X4 _u0_u22_U283  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[8] ) );
INV_X4 _u0_u22_U281  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[7] ) );
INV_X4 _u0_u22_U279  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[6] ) );
INV_X4 _u0_u22_U277  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[5] ) );
INV_X4 _u0_u22_U275  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[4] ) );
INV_X4 _u0_u22_U273  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[3] ) );
INV_X4 _u0_u22_U271  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[2] ) );
INV_X4 _u0_u22_U269  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[1] ) );
INV_X4 _u0_u22_U267  ( .A(1'b1), .ZN(_u0_u22_ch_adr0[0] ) );
INV_X4 _u0_u22_U265  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[31] ) );
INV_X4 _u0_u22_U263  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[30] ) );
INV_X4 _u0_u22_U261  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[29] ) );
INV_X4 _u0_u22_U259  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[28] ) );
INV_X4 _u0_u22_U257  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[27] ) );
INV_X4 _u0_u22_U255  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[26] ) );
INV_X4 _u0_u22_U253  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[25] ) );
INV_X4 _u0_u22_U251  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[24] ) );
INV_X4 _u0_u22_U249  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[23] ) );
INV_X4 _u0_u22_U247  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[22] ) );
INV_X4 _u0_u22_U245  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[21] ) );
INV_X4 _u0_u22_U243  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[20] ) );
INV_X4 _u0_u22_U241  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[19] ) );
INV_X4 _u0_u22_U239  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[18] ) );
INV_X4 _u0_u22_U237  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[17] ) );
INV_X4 _u0_u22_U235  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[16] ) );
INV_X4 _u0_u22_U233  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[15] ) );
INV_X4 _u0_u22_U231  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[14] ) );
INV_X4 _u0_u22_U229  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[13] ) );
INV_X4 _u0_u22_U227  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[12] ) );
INV_X4 _u0_u22_U225  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[11] ) );
INV_X4 _u0_u22_U223  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[10] ) );
INV_X4 _u0_u22_U221  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[9] ) );
INV_X4 _u0_u22_U219  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[8] ) );
INV_X4 _u0_u22_U217  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[7] ) );
INV_X4 _u0_u22_U215  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[6] ) );
INV_X4 _u0_u22_U213  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[5] ) );
INV_X4 _u0_u22_U211  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[4] ) );
INV_X4 _u0_u22_U209  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[3] ) );
INV_X4 _u0_u22_U207  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[2] ) );
INV_X4 _u0_u22_U205  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[1] ) );
INV_X4 _u0_u22_U203  ( .A(1'b1), .ZN(_u0_u22_ch_adr1[0] ) );
INV_X4 _u0_u22_U201  ( .A(1'b0), .ZN(_u0_u22_ch_am0[31] ) );
INV_X4 _u0_u22_U199  ( .A(1'b0), .ZN(_u0_u22_ch_am0[30] ) );
INV_X4 _u0_u22_U197  ( .A(1'b0), .ZN(_u0_u22_ch_am0[29] ) );
INV_X4 _u0_u22_U195  ( .A(1'b0), .ZN(_u0_u22_ch_am0[28] ) );
INV_X4 _u0_u22_U193  ( .A(1'b0), .ZN(_u0_u22_ch_am0[27] ) );
INV_X4 _u0_u22_U191  ( .A(1'b0), .ZN(_u0_u22_ch_am0[26] ) );
INV_X4 _u0_u22_U189  ( .A(1'b0), .ZN(_u0_u22_ch_am0[25] ) );
INV_X4 _u0_u22_U187  ( .A(1'b0), .ZN(_u0_u22_ch_am0[24] ) );
INV_X4 _u0_u22_U185  ( .A(1'b0), .ZN(_u0_u22_ch_am0[23] ) );
INV_X4 _u0_u22_U183  ( .A(1'b0), .ZN(_u0_u22_ch_am0[22] ) );
INV_X4 _u0_u22_U181  ( .A(1'b0), .ZN(_u0_u22_ch_am0[21] ) );
INV_X4 _u0_u22_U179  ( .A(1'b0), .ZN(_u0_u22_ch_am0[20] ) );
INV_X4 _u0_u22_U177  ( .A(1'b0), .ZN(_u0_u22_ch_am0[19] ) );
INV_X4 _u0_u22_U175  ( .A(1'b0), .ZN(_u0_u22_ch_am0[18] ) );
INV_X4 _u0_u22_U173  ( .A(1'b0), .ZN(_u0_u22_ch_am0[17] ) );
INV_X4 _u0_u22_U171  ( .A(1'b0), .ZN(_u0_u22_ch_am0[16] ) );
INV_X4 _u0_u22_U169  ( .A(1'b0), .ZN(_u0_u22_ch_am0[15] ) );
INV_X4 _u0_u22_U167  ( .A(1'b0), .ZN(_u0_u22_ch_am0[14] ) );
INV_X4 _u0_u22_U165  ( .A(1'b0), .ZN(_u0_u22_ch_am0[13] ) );
INV_X4 _u0_u22_U163  ( .A(1'b0), .ZN(_u0_u22_ch_am0[12] ) );
INV_X4 _u0_u22_U161  ( .A(1'b0), .ZN(_u0_u22_ch_am0[11] ) );
INV_X4 _u0_u22_U159  ( .A(1'b0), .ZN(_u0_u22_ch_am0[10] ) );
INV_X4 _u0_u22_U157  ( .A(1'b0), .ZN(_u0_u22_ch_am0[9] ) );
INV_X4 _u0_u22_U155  ( .A(1'b0), .ZN(_u0_u22_ch_am0[8] ) );
INV_X4 _u0_u22_U153  ( .A(1'b0), .ZN(_u0_u22_ch_am0[7] ) );
INV_X4 _u0_u22_U151  ( .A(1'b0), .ZN(_u0_u22_ch_am0[6] ) );
INV_X4 _u0_u22_U149  ( .A(1'b0), .ZN(_u0_u22_ch_am0[5] ) );
INV_X4 _u0_u22_U147  ( .A(1'b0), .ZN(_u0_u22_ch_am0[4] ) );
INV_X4 _u0_u22_U145  ( .A(1'b1), .ZN(_u0_u22_ch_am0[3] ) );
INV_X4 _u0_u22_U143  ( .A(1'b1), .ZN(_u0_u22_ch_am0[2] ) );
INV_X4 _u0_u22_U141  ( .A(1'b1), .ZN(_u0_u22_ch_am0[1] ) );
INV_X4 _u0_u22_U139  ( .A(1'b1), .ZN(_u0_u22_ch_am0[0] ) );
INV_X4 _u0_u22_U137  ( .A(1'b0), .ZN(_u0_u22_ch_am1[31] ) );
INV_X4 _u0_u22_U135  ( .A(1'b0), .ZN(_u0_u22_ch_am1[30] ) );
INV_X4 _u0_u22_U133  ( .A(1'b0), .ZN(_u0_u22_ch_am1[29] ) );
INV_X4 _u0_u22_U131  ( .A(1'b0), .ZN(_u0_u22_ch_am1[28] ) );
INV_X4 _u0_u22_U129  ( .A(1'b0), .ZN(_u0_u22_ch_am1[27] ) );
INV_X4 _u0_u22_U127  ( .A(1'b0), .ZN(_u0_u22_ch_am1[26] ) );
INV_X4 _u0_u22_U125  ( .A(1'b0), .ZN(_u0_u22_ch_am1[25] ) );
INV_X4 _u0_u22_U123  ( .A(1'b0), .ZN(_u0_u22_ch_am1[24] ) );
INV_X4 _u0_u22_U121  ( .A(1'b0), .ZN(_u0_u22_ch_am1[23] ) );
INV_X4 _u0_u22_U119  ( .A(1'b0), .ZN(_u0_u22_ch_am1[22] ) );
INV_X4 _u0_u22_U117  ( .A(1'b0), .ZN(_u0_u22_ch_am1[21] ) );
INV_X4 _u0_u22_U115  ( .A(1'b0), .ZN(_u0_u22_ch_am1[20] ) );
INV_X4 _u0_u22_U113  ( .A(1'b0), .ZN(_u0_u22_ch_am1[19] ) );
INV_X4 _u0_u22_U111  ( .A(1'b0), .ZN(_u0_u22_ch_am1[18] ) );
INV_X4 _u0_u22_U109  ( .A(1'b0), .ZN(_u0_u22_ch_am1[17] ) );
INV_X4 _u0_u22_U107  ( .A(1'b0), .ZN(_u0_u22_ch_am1[16] ) );
INV_X4 _u0_u22_U105  ( .A(1'b0), .ZN(_u0_u22_ch_am1[15] ) );
INV_X4 _u0_u22_U103  ( .A(1'b0), .ZN(_u0_u22_ch_am1[14] ) );
INV_X4 _u0_u22_U101  ( .A(1'b0), .ZN(_u0_u22_ch_am1[13] ) );
INV_X4 _u0_u22_U99  ( .A(1'b0), .ZN(_u0_u22_ch_am1[12] ) );
INV_X4 _u0_u22_U97  ( .A(1'b0), .ZN(_u0_u22_ch_am1[11] ) );
INV_X4 _u0_u22_U95  ( .A(1'b0), .ZN(_u0_u22_ch_am1[10] ) );
INV_X4 _u0_u22_U93  ( .A(1'b0), .ZN(_u0_u22_ch_am1[9] ) );
INV_X4 _u0_u22_U91  ( .A(1'b0), .ZN(_u0_u22_ch_am1[8] ) );
INV_X4 _u0_u22_U89  ( .A(1'b0), .ZN(_u0_u22_ch_am1[7] ) );
INV_X4 _u0_u22_U87  ( .A(1'b0), .ZN(_u0_u22_ch_am1[6] ) );
INV_X4 _u0_u22_U85  ( .A(1'b0), .ZN(_u0_u22_ch_am1[5] ) );
INV_X4 _u0_u22_U83  ( .A(1'b0), .ZN(_u0_u22_ch_am1[4] ) );
INV_X4 _u0_u22_U81  ( .A(1'b1), .ZN(_u0_u22_ch_am1[3] ) );
INV_X4 _u0_u22_U79  ( .A(1'b1), .ZN(_u0_u22_ch_am1[2] ) );
INV_X4 _u0_u22_U77  ( .A(1'b1), .ZN(_u0_u22_ch_am1[1] ) );
INV_X4 _u0_u22_U75  ( .A(1'b1), .ZN(_u0_u22_ch_am1[0] ) );
INV_X4 _u0_u22_U73  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[31] ) );
INV_X4 _u0_u22_U71  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[30] ) );
INV_X4 _u0_u22_U69  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[29] ) );
INV_X4 _u0_u22_U67  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[28] ) );
INV_X4 _u0_u22_U65  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[27] ) );
INV_X4 _u0_u22_U63  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[26] ) );
INV_X4 _u0_u22_U61  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[25] ) );
INV_X4 _u0_u22_U59  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[24] ) );
INV_X4 _u0_u22_U57  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[23] ) );
INV_X4 _u0_u22_U55  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[22] ) );
INV_X4 _u0_u22_U53  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[21] ) );
INV_X4 _u0_u22_U51  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[20] ) );
INV_X4 _u0_u22_U49  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[19] ) );
INV_X4 _u0_u22_U47  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[18] ) );
INV_X4 _u0_u22_U45  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[17] ) );
INV_X4 _u0_u22_U43  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[16] ) );
INV_X4 _u0_u22_U41  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[15] ) );
INV_X4 _u0_u22_U39  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[14] ) );
INV_X4 _u0_u22_U37  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[13] ) );
INV_X4 _u0_u22_U35  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[12] ) );
INV_X4 _u0_u22_U33  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[11] ) );
INV_X4 _u0_u22_U31  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[10] ) );
INV_X4 _u0_u22_U29  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[9] ) );
INV_X4 _u0_u22_U27  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[8] ) );
INV_X4 _u0_u22_U25  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[7] ) );
INV_X4 _u0_u22_U23  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[6] ) );
INV_X4 _u0_u22_U21  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[5] ) );
INV_X4 _u0_u22_U19  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[4] ) );
INV_X4 _u0_u22_U17  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[3] ) );
INV_X4 _u0_u22_U15  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[2] ) );
INV_X4 _u0_u22_U13  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[1] ) );
INV_X4 _u0_u22_U11  ( .A(1'b1), .ZN(_u0_u22_sw_pointer[0] ) );
INV_X4 _u0_u22_U9  ( .A(1'b1), .ZN(_u0_u22_ch_stop ) );
INV_X4 _u0_u22_U7  ( .A(1'b1), .ZN(_u0_u22_ch_dis ) );
INV_X4 _u0_u22_U5  ( .A(1'b1), .ZN(_u0_u22_int ) );
INV_X4 _u0_u23_U585  ( .A(1'b1), .ZN(_u0_u23_pointer[31] ) );
INV_X4 _u0_u23_U583  ( .A(1'b1), .ZN(_u0_u23_pointer[30] ) );
INV_X4 _u0_u23_U581  ( .A(1'b1), .ZN(_u0_u23_pointer[29] ) );
INV_X4 _u0_u23_U579  ( .A(1'b1), .ZN(_u0_u23_pointer[28] ) );
INV_X4 _u0_u23_U577  ( .A(1'b1), .ZN(_u0_u23_pointer[27] ) );
INV_X4 _u0_u23_U575  ( .A(1'b1), .ZN(_u0_u23_pointer[26] ) );
INV_X4 _u0_u23_U573  ( .A(1'b1), .ZN(_u0_u23_pointer[25] ) );
INV_X4 _u0_u23_U571  ( .A(1'b1), .ZN(_u0_u23_pointer[24] ) );
INV_X4 _u0_u23_U569  ( .A(1'b1), .ZN(_u0_u23_pointer[23] ) );
INV_X4 _u0_u23_U567  ( .A(1'b1), .ZN(_u0_u23_pointer[22] ) );
INV_X4 _u0_u23_U565  ( .A(1'b1), .ZN(_u0_u23_pointer[21] ) );
INV_X4 _u0_u23_U563  ( .A(1'b1), .ZN(_u0_u23_pointer[20] ) );
INV_X4 _u0_u23_U561  ( .A(1'b1), .ZN(_u0_u23_pointer[19] ) );
INV_X4 _u0_u23_U559  ( .A(1'b1), .ZN(_u0_u23_pointer[18] ) );
INV_X4 _u0_u23_U557  ( .A(1'b1), .ZN(_u0_u23_pointer[17] ) );
INV_X4 _u0_u23_U555  ( .A(1'b1), .ZN(_u0_u23_pointer[16] ) );
INV_X4 _u0_u23_U553  ( .A(1'b1), .ZN(_u0_u23_pointer[15] ) );
INV_X4 _u0_u23_U551  ( .A(1'b1), .ZN(_u0_u23_pointer[14] ) );
INV_X4 _u0_u23_U549  ( .A(1'b1), .ZN(_u0_u23_pointer[13] ) );
INV_X4 _u0_u23_U547  ( .A(1'b1), .ZN(_u0_u23_pointer[12] ) );
INV_X4 _u0_u23_U545  ( .A(1'b1), .ZN(_u0_u23_pointer[11] ) );
INV_X4 _u0_u23_U543  ( .A(1'b1), .ZN(_u0_u23_pointer[10] ) );
INV_X4 _u0_u23_U541  ( .A(1'b1), .ZN(_u0_u23_pointer[9] ) );
INV_X4 _u0_u23_U539  ( .A(1'b1), .ZN(_u0_u23_pointer[8] ) );
INV_X4 _u0_u23_U537  ( .A(1'b1), .ZN(_u0_u23_pointer[7] ) );
INV_X4 _u0_u23_U535  ( .A(1'b1), .ZN(_u0_u23_pointer[6] ) );
INV_X4 _u0_u23_U533  ( .A(1'b1), .ZN(_u0_u23_pointer[5] ) );
INV_X4 _u0_u23_U531  ( .A(1'b1), .ZN(_u0_u23_pointer[4] ) );
INV_X4 _u0_u23_U529  ( .A(1'b1), .ZN(_u0_u23_pointer[3] ) );
INV_X4 _u0_u23_U527  ( .A(1'b1), .ZN(_u0_u23_pointer[2] ) );
INV_X4 _u0_u23_U525  ( .A(1'b1), .ZN(_u0_u23_pointer[1] ) );
INV_X4 _u0_u23_U523  ( .A(1'b1), .ZN(_u0_u23_pointer[0] ) );
INV_X4 _u0_u23_U521  ( .A(1'b1), .ZN(_u0_u23_pointer_s[31] ) );
INV_X4 _u0_u23_U519  ( .A(1'b1), .ZN(_u0_u23_pointer_s[30] ) );
INV_X4 _u0_u23_U517  ( .A(1'b1), .ZN(_u0_u23_pointer_s[29] ) );
INV_X4 _u0_u23_U515  ( .A(1'b1), .ZN(_u0_u23_pointer_s[28] ) );
INV_X4 _u0_u23_U513  ( .A(1'b1), .ZN(_u0_u23_pointer_s[27] ) );
INV_X4 _u0_u23_U511  ( .A(1'b1), .ZN(_u0_u23_pointer_s[26] ) );
INV_X4 _u0_u23_U509  ( .A(1'b1), .ZN(_u0_u23_pointer_s[25] ) );
INV_X4 _u0_u23_U507  ( .A(1'b1), .ZN(_u0_u23_pointer_s[24] ) );
INV_X4 _u0_u23_U505  ( .A(1'b1), .ZN(_u0_u23_pointer_s[23] ) );
INV_X4 _u0_u23_U503  ( .A(1'b1), .ZN(_u0_u23_pointer_s[22] ) );
INV_X4 _u0_u23_U501  ( .A(1'b1), .ZN(_u0_u23_pointer_s[21] ) );
INV_X4 _u0_u23_U499  ( .A(1'b1), .ZN(_u0_u23_pointer_s[20] ) );
INV_X4 _u0_u23_U497  ( .A(1'b1), .ZN(_u0_u23_pointer_s[19] ) );
INV_X4 _u0_u23_U495  ( .A(1'b1), .ZN(_u0_u23_pointer_s[18] ) );
INV_X4 _u0_u23_U493  ( .A(1'b1), .ZN(_u0_u23_pointer_s[17] ) );
INV_X4 _u0_u23_U491  ( .A(1'b1), .ZN(_u0_u23_pointer_s[16] ) );
INV_X4 _u0_u23_U489  ( .A(1'b1), .ZN(_u0_u23_pointer_s[15] ) );
INV_X4 _u0_u23_U487  ( .A(1'b1), .ZN(_u0_u23_pointer_s[14] ) );
INV_X4 _u0_u23_U485  ( .A(1'b1), .ZN(_u0_u23_pointer_s[13] ) );
INV_X4 _u0_u23_U483  ( .A(1'b1), .ZN(_u0_u23_pointer_s[12] ) );
INV_X4 _u0_u23_U481  ( .A(1'b1), .ZN(_u0_u23_pointer_s[11] ) );
INV_X4 _u0_u23_U479  ( .A(1'b1), .ZN(_u0_u23_pointer_s[10] ) );
INV_X4 _u0_u23_U477  ( .A(1'b1), .ZN(_u0_u23_pointer_s[9] ) );
INV_X4 _u0_u23_U475  ( .A(1'b1), .ZN(_u0_u23_pointer_s[8] ) );
INV_X4 _u0_u23_U473  ( .A(1'b1), .ZN(_u0_u23_pointer_s[7] ) );
INV_X4 _u0_u23_U471  ( .A(1'b1), .ZN(_u0_u23_pointer_s[6] ) );
INV_X4 _u0_u23_U469  ( .A(1'b1), .ZN(_u0_u23_pointer_s[5] ) );
INV_X4 _u0_u23_U467  ( .A(1'b1), .ZN(_u0_u23_pointer_s[4] ) );
INV_X4 _u0_u23_U465  ( .A(1'b1), .ZN(_u0_u23_pointer_s[3] ) );
INV_X4 _u0_u23_U463  ( .A(1'b1), .ZN(_u0_u23_pointer_s[2] ) );
INV_X4 _u0_u23_U461  ( .A(1'b1), .ZN(_u0_u23_pointer_s[1] ) );
INV_X4 _u0_u23_U459  ( .A(1'b1), .ZN(_u0_u23_pointer_s[0] ) );
INV_X4 _u0_u23_U457  ( .A(1'b1), .ZN(_u0_u23_ch_csr[31] ) );
INV_X4 _u0_u23_U455  ( .A(1'b1), .ZN(_u0_u23_ch_csr[30] ) );
INV_X4 _u0_u23_U453  ( .A(1'b1), .ZN(_u0_u23_ch_csr[29] ) );
INV_X4 _u0_u23_U451  ( .A(1'b1), .ZN(_u0_u23_ch_csr[28] ) );
INV_X4 _u0_u23_U449  ( .A(1'b1), .ZN(_u0_u23_ch_csr[27] ) );
INV_X4 _u0_u23_U447  ( .A(1'b1), .ZN(_u0_u23_ch_csr[26] ) );
INV_X4 _u0_u23_U445  ( .A(1'b1), .ZN(_u0_u23_ch_csr[25] ) );
INV_X4 _u0_u23_U443  ( .A(1'b1), .ZN(_u0_u23_ch_csr[24] ) );
INV_X4 _u0_u23_U441  ( .A(1'b1), .ZN(_u0_u23_ch_csr[23] ) );
INV_X4 _u0_u23_U439  ( .A(1'b1), .ZN(_u0_u23_ch_csr[22] ) );
INV_X4 _u0_u23_U437  ( .A(1'b1), .ZN(_u0_u23_ch_csr[21] ) );
INV_X4 _u0_u23_U435  ( .A(1'b1), .ZN(_u0_u23_ch_csr[20] ) );
INV_X4 _u0_u23_U433  ( .A(1'b1), .ZN(_u0_u23_ch_csr[19] ) );
INV_X4 _u0_u23_U431  ( .A(1'b1), .ZN(_u0_u23_ch_csr[18] ) );
INV_X4 _u0_u23_U429  ( .A(1'b1), .ZN(_u0_u23_ch_csr[17] ) );
INV_X4 _u0_u23_U427  ( .A(1'b1), .ZN(_u0_u23_ch_csr[16] ) );
INV_X4 _u0_u23_U425  ( .A(1'b1), .ZN(_u0_u23_ch_csr[15] ) );
INV_X4 _u0_u23_U423  ( .A(1'b1), .ZN(_u0_u23_ch_csr[14] ) );
INV_X4 _u0_u23_U421  ( .A(1'b1), .ZN(_u0_u23_ch_csr[13] ) );
INV_X4 _u0_u23_U419  ( .A(1'b1), .ZN(_u0_u23_ch_csr[12] ) );
INV_X4 _u0_u23_U417  ( .A(1'b1), .ZN(_u0_u23_ch_csr[11] ) );
INV_X4 _u0_u23_U415  ( .A(1'b1), .ZN(_u0_u23_ch_csr[10] ) );
INV_X4 _u0_u23_U413  ( .A(1'b1), .ZN(_u0_u23_ch_csr[9] ) );
INV_X4 _u0_u23_U411  ( .A(1'b1), .ZN(_u0_u23_ch_csr[8] ) );
INV_X4 _u0_u23_U409  ( .A(1'b1), .ZN(_u0_u23_ch_csr[7] ) );
INV_X4 _u0_u23_U407  ( .A(1'b1), .ZN(_u0_u23_ch_csr[6] ) );
INV_X4 _u0_u23_U405  ( .A(1'b1), .ZN(_u0_u23_ch_csr[5] ) );
INV_X4 _u0_u23_U403  ( .A(1'b1), .ZN(_u0_u23_ch_csr[4] ) );
INV_X4 _u0_u23_U401  ( .A(1'b1), .ZN(_u0_u23_ch_csr[3] ) );
INV_X4 _u0_u23_U399  ( .A(1'b1), .ZN(_u0_u23_ch_csr[2] ) );
INV_X4 _u0_u23_U397  ( .A(1'b1), .ZN(_u0_u23_ch_csr[1] ) );
INV_X4 _u0_u23_U395  ( .A(1'b1), .ZN(_u0_u23_ch_csr[0] ) );
INV_X4 _u0_u23_U393  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[31] ) );
INV_X4 _u0_u23_U391  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[30] ) );
INV_X4 _u0_u23_U389  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[29] ) );
INV_X4 _u0_u23_U387  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[28] ) );
INV_X4 _u0_u23_U385  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[27] ) );
INV_X4 _u0_u23_U383  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[26] ) );
INV_X4 _u0_u23_U381  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[25] ) );
INV_X4 _u0_u23_U379  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[24] ) );
INV_X4 _u0_u23_U377  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[23] ) );
INV_X4 _u0_u23_U375  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[22] ) );
INV_X4 _u0_u23_U373  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[21] ) );
INV_X4 _u0_u23_U371  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[20] ) );
INV_X4 _u0_u23_U369  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[19] ) );
INV_X4 _u0_u23_U367  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[18] ) );
INV_X4 _u0_u23_U365  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[17] ) );
INV_X4 _u0_u23_U363  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[16] ) );
INV_X4 _u0_u23_U361  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[15] ) );
INV_X4 _u0_u23_U359  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[14] ) );
INV_X4 _u0_u23_U357  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[13] ) );
INV_X4 _u0_u23_U355  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[12] ) );
INV_X4 _u0_u23_U353  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[11] ) );
INV_X4 _u0_u23_U351  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[10] ) );
INV_X4 _u0_u23_U349  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[9] ) );
INV_X4 _u0_u23_U347  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[8] ) );
INV_X4 _u0_u23_U345  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[7] ) );
INV_X4 _u0_u23_U343  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[6] ) );
INV_X4 _u0_u23_U341  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[5] ) );
INV_X4 _u0_u23_U339  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[4] ) );
INV_X4 _u0_u23_U337  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[3] ) );
INV_X4 _u0_u23_U335  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[2] ) );
INV_X4 _u0_u23_U333  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[1] ) );
INV_X4 _u0_u23_U331  ( .A(1'b1), .ZN(_u0_u23_ch_txsz[0] ) );
INV_X4 _u0_u23_U329  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[31] ) );
INV_X4 _u0_u23_U327  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[30] ) );
INV_X4 _u0_u23_U325  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[29] ) );
INV_X4 _u0_u23_U323  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[28] ) );
INV_X4 _u0_u23_U321  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[27] ) );
INV_X4 _u0_u23_U319  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[26] ) );
INV_X4 _u0_u23_U317  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[25] ) );
INV_X4 _u0_u23_U315  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[24] ) );
INV_X4 _u0_u23_U313  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[23] ) );
INV_X4 _u0_u23_U311  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[22] ) );
INV_X4 _u0_u23_U309  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[21] ) );
INV_X4 _u0_u23_U307  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[20] ) );
INV_X4 _u0_u23_U305  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[19] ) );
INV_X4 _u0_u23_U303  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[18] ) );
INV_X4 _u0_u23_U301  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[17] ) );
INV_X4 _u0_u23_U299  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[16] ) );
INV_X4 _u0_u23_U297  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[15] ) );
INV_X4 _u0_u23_U295  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[14] ) );
INV_X4 _u0_u23_U293  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[13] ) );
INV_X4 _u0_u23_U291  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[12] ) );
INV_X4 _u0_u23_U289  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[11] ) );
INV_X4 _u0_u23_U287  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[10] ) );
INV_X4 _u0_u23_U285  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[9] ) );
INV_X4 _u0_u23_U283  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[8] ) );
INV_X4 _u0_u23_U281  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[7] ) );
INV_X4 _u0_u23_U279  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[6] ) );
INV_X4 _u0_u23_U277  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[5] ) );
INV_X4 _u0_u23_U275  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[4] ) );
INV_X4 _u0_u23_U273  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[3] ) );
INV_X4 _u0_u23_U271  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[2] ) );
INV_X4 _u0_u23_U269  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[1] ) );
INV_X4 _u0_u23_U267  ( .A(1'b1), .ZN(_u0_u23_ch_adr0[0] ) );
INV_X4 _u0_u23_U265  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[31] ) );
INV_X4 _u0_u23_U263  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[30] ) );
INV_X4 _u0_u23_U261  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[29] ) );
INV_X4 _u0_u23_U259  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[28] ) );
INV_X4 _u0_u23_U257  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[27] ) );
INV_X4 _u0_u23_U255  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[26] ) );
INV_X4 _u0_u23_U253  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[25] ) );
INV_X4 _u0_u23_U251  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[24] ) );
INV_X4 _u0_u23_U249  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[23] ) );
INV_X4 _u0_u23_U247  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[22] ) );
INV_X4 _u0_u23_U245  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[21] ) );
INV_X4 _u0_u23_U243  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[20] ) );
INV_X4 _u0_u23_U241  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[19] ) );
INV_X4 _u0_u23_U239  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[18] ) );
INV_X4 _u0_u23_U237  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[17] ) );
INV_X4 _u0_u23_U235  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[16] ) );
INV_X4 _u0_u23_U233  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[15] ) );
INV_X4 _u0_u23_U231  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[14] ) );
INV_X4 _u0_u23_U229  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[13] ) );
INV_X4 _u0_u23_U227  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[12] ) );
INV_X4 _u0_u23_U225  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[11] ) );
INV_X4 _u0_u23_U223  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[10] ) );
INV_X4 _u0_u23_U221  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[9] ) );
INV_X4 _u0_u23_U219  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[8] ) );
INV_X4 _u0_u23_U217  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[7] ) );
INV_X4 _u0_u23_U215  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[6] ) );
INV_X4 _u0_u23_U213  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[5] ) );
INV_X4 _u0_u23_U211  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[4] ) );
INV_X4 _u0_u23_U209  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[3] ) );
INV_X4 _u0_u23_U207  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[2] ) );
INV_X4 _u0_u23_U205  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[1] ) );
INV_X4 _u0_u23_U203  ( .A(1'b1), .ZN(_u0_u23_ch_adr1[0] ) );
INV_X4 _u0_u23_U201  ( .A(1'b0), .ZN(_u0_u23_ch_am0[31] ) );
INV_X4 _u0_u23_U199  ( .A(1'b0), .ZN(_u0_u23_ch_am0[30] ) );
INV_X4 _u0_u23_U197  ( .A(1'b0), .ZN(_u0_u23_ch_am0[29] ) );
INV_X4 _u0_u23_U195  ( .A(1'b0), .ZN(_u0_u23_ch_am0[28] ) );
INV_X4 _u0_u23_U193  ( .A(1'b0), .ZN(_u0_u23_ch_am0[27] ) );
INV_X4 _u0_u23_U191  ( .A(1'b0), .ZN(_u0_u23_ch_am0[26] ) );
INV_X4 _u0_u23_U189  ( .A(1'b0), .ZN(_u0_u23_ch_am0[25] ) );
INV_X4 _u0_u23_U187  ( .A(1'b0), .ZN(_u0_u23_ch_am0[24] ) );
INV_X4 _u0_u23_U185  ( .A(1'b0), .ZN(_u0_u23_ch_am0[23] ) );
INV_X4 _u0_u23_U183  ( .A(1'b0), .ZN(_u0_u23_ch_am0[22] ) );
INV_X4 _u0_u23_U181  ( .A(1'b0), .ZN(_u0_u23_ch_am0[21] ) );
INV_X4 _u0_u23_U179  ( .A(1'b0), .ZN(_u0_u23_ch_am0[20] ) );
INV_X4 _u0_u23_U177  ( .A(1'b0), .ZN(_u0_u23_ch_am0[19] ) );
INV_X4 _u0_u23_U175  ( .A(1'b0), .ZN(_u0_u23_ch_am0[18] ) );
INV_X4 _u0_u23_U173  ( .A(1'b0), .ZN(_u0_u23_ch_am0[17] ) );
INV_X4 _u0_u23_U171  ( .A(1'b0), .ZN(_u0_u23_ch_am0[16] ) );
INV_X4 _u0_u23_U169  ( .A(1'b0), .ZN(_u0_u23_ch_am0[15] ) );
INV_X4 _u0_u23_U167  ( .A(1'b0), .ZN(_u0_u23_ch_am0[14] ) );
INV_X4 _u0_u23_U165  ( .A(1'b0), .ZN(_u0_u23_ch_am0[13] ) );
INV_X4 _u0_u23_U163  ( .A(1'b0), .ZN(_u0_u23_ch_am0[12] ) );
INV_X4 _u0_u23_U161  ( .A(1'b0), .ZN(_u0_u23_ch_am0[11] ) );
INV_X4 _u0_u23_U159  ( .A(1'b0), .ZN(_u0_u23_ch_am0[10] ) );
INV_X4 _u0_u23_U157  ( .A(1'b0), .ZN(_u0_u23_ch_am0[9] ) );
INV_X4 _u0_u23_U155  ( .A(1'b0), .ZN(_u0_u23_ch_am0[8] ) );
INV_X4 _u0_u23_U153  ( .A(1'b0), .ZN(_u0_u23_ch_am0[7] ) );
INV_X4 _u0_u23_U151  ( .A(1'b0), .ZN(_u0_u23_ch_am0[6] ) );
INV_X4 _u0_u23_U149  ( .A(1'b0), .ZN(_u0_u23_ch_am0[5] ) );
INV_X4 _u0_u23_U147  ( .A(1'b0), .ZN(_u0_u23_ch_am0[4] ) );
INV_X4 _u0_u23_U145  ( .A(1'b1), .ZN(_u0_u23_ch_am0[3] ) );
INV_X4 _u0_u23_U143  ( .A(1'b1), .ZN(_u0_u23_ch_am0[2] ) );
INV_X4 _u0_u23_U141  ( .A(1'b1), .ZN(_u0_u23_ch_am0[1] ) );
INV_X4 _u0_u23_U139  ( .A(1'b1), .ZN(_u0_u23_ch_am0[0] ) );
INV_X4 _u0_u23_U137  ( .A(1'b0), .ZN(_u0_u23_ch_am1[31] ) );
INV_X4 _u0_u23_U135  ( .A(1'b0), .ZN(_u0_u23_ch_am1[30] ) );
INV_X4 _u0_u23_U133  ( .A(1'b0), .ZN(_u0_u23_ch_am1[29] ) );
INV_X4 _u0_u23_U131  ( .A(1'b0), .ZN(_u0_u23_ch_am1[28] ) );
INV_X4 _u0_u23_U129  ( .A(1'b0), .ZN(_u0_u23_ch_am1[27] ) );
INV_X4 _u0_u23_U127  ( .A(1'b0), .ZN(_u0_u23_ch_am1[26] ) );
INV_X4 _u0_u23_U125  ( .A(1'b0), .ZN(_u0_u23_ch_am1[25] ) );
INV_X4 _u0_u23_U123  ( .A(1'b0), .ZN(_u0_u23_ch_am1[24] ) );
INV_X4 _u0_u23_U121  ( .A(1'b0), .ZN(_u0_u23_ch_am1[23] ) );
INV_X4 _u0_u23_U119  ( .A(1'b0), .ZN(_u0_u23_ch_am1[22] ) );
INV_X4 _u0_u23_U117  ( .A(1'b0), .ZN(_u0_u23_ch_am1[21] ) );
INV_X4 _u0_u23_U115  ( .A(1'b0), .ZN(_u0_u23_ch_am1[20] ) );
INV_X4 _u0_u23_U113  ( .A(1'b0), .ZN(_u0_u23_ch_am1[19] ) );
INV_X4 _u0_u23_U111  ( .A(1'b0), .ZN(_u0_u23_ch_am1[18] ) );
INV_X4 _u0_u23_U109  ( .A(1'b0), .ZN(_u0_u23_ch_am1[17] ) );
INV_X4 _u0_u23_U107  ( .A(1'b0), .ZN(_u0_u23_ch_am1[16] ) );
INV_X4 _u0_u23_U105  ( .A(1'b0), .ZN(_u0_u23_ch_am1[15] ) );
INV_X4 _u0_u23_U103  ( .A(1'b0), .ZN(_u0_u23_ch_am1[14] ) );
INV_X4 _u0_u23_U101  ( .A(1'b0), .ZN(_u0_u23_ch_am1[13] ) );
INV_X4 _u0_u23_U99  ( .A(1'b0), .ZN(_u0_u23_ch_am1[12] ) );
INV_X4 _u0_u23_U97  ( .A(1'b0), .ZN(_u0_u23_ch_am1[11] ) );
INV_X4 _u0_u23_U95  ( .A(1'b0), .ZN(_u0_u23_ch_am1[10] ) );
INV_X4 _u0_u23_U93  ( .A(1'b0), .ZN(_u0_u23_ch_am1[9] ) );
INV_X4 _u0_u23_U91  ( .A(1'b0), .ZN(_u0_u23_ch_am1[8] ) );
INV_X4 _u0_u23_U89  ( .A(1'b0), .ZN(_u0_u23_ch_am1[7] ) );
INV_X4 _u0_u23_U87  ( .A(1'b0), .ZN(_u0_u23_ch_am1[6] ) );
INV_X4 _u0_u23_U85  ( .A(1'b0), .ZN(_u0_u23_ch_am1[5] ) );
INV_X4 _u0_u23_U83  ( .A(1'b0), .ZN(_u0_u23_ch_am1[4] ) );
INV_X4 _u0_u23_U81  ( .A(1'b1), .ZN(_u0_u23_ch_am1[3] ) );
INV_X4 _u0_u23_U79  ( .A(1'b1), .ZN(_u0_u23_ch_am1[2] ) );
INV_X4 _u0_u23_U77  ( .A(1'b1), .ZN(_u0_u23_ch_am1[1] ) );
INV_X4 _u0_u23_U75  ( .A(1'b1), .ZN(_u0_u23_ch_am1[0] ) );
INV_X4 _u0_u23_U73  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[31] ) );
INV_X4 _u0_u23_U71  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[30] ) );
INV_X4 _u0_u23_U69  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[29] ) );
INV_X4 _u0_u23_U67  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[28] ) );
INV_X4 _u0_u23_U65  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[27] ) );
INV_X4 _u0_u23_U63  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[26] ) );
INV_X4 _u0_u23_U61  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[25] ) );
INV_X4 _u0_u23_U59  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[24] ) );
INV_X4 _u0_u23_U57  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[23] ) );
INV_X4 _u0_u23_U55  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[22] ) );
INV_X4 _u0_u23_U53  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[21] ) );
INV_X4 _u0_u23_U51  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[20] ) );
INV_X4 _u0_u23_U49  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[19] ) );
INV_X4 _u0_u23_U47  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[18] ) );
INV_X4 _u0_u23_U45  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[17] ) );
INV_X4 _u0_u23_U43  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[16] ) );
INV_X4 _u0_u23_U41  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[15] ) );
INV_X4 _u0_u23_U39  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[14] ) );
INV_X4 _u0_u23_U37  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[13] ) );
INV_X4 _u0_u23_U35  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[12] ) );
INV_X4 _u0_u23_U33  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[11] ) );
INV_X4 _u0_u23_U31  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[10] ) );
INV_X4 _u0_u23_U29  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[9] ) );
INV_X4 _u0_u23_U27  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[8] ) );
INV_X4 _u0_u23_U25  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[7] ) );
INV_X4 _u0_u23_U23  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[6] ) );
INV_X4 _u0_u23_U21  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[5] ) );
INV_X4 _u0_u23_U19  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[4] ) );
INV_X4 _u0_u23_U17  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[3] ) );
INV_X4 _u0_u23_U15  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[2] ) );
INV_X4 _u0_u23_U13  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[1] ) );
INV_X4 _u0_u23_U11  ( .A(1'b1), .ZN(_u0_u23_sw_pointer[0] ) );
INV_X4 _u0_u23_U9  ( .A(1'b1), .ZN(_u0_u23_ch_stop ) );
INV_X4 _u0_u23_U7  ( .A(1'b1), .ZN(_u0_u23_ch_dis ) );
INV_X4 _u0_u23_U5  ( .A(1'b1), .ZN(_u0_u23_int ) );
INV_X4 _u0_u24_U585  ( .A(1'b1), .ZN(_u0_u24_pointer[31] ) );
INV_X4 _u0_u24_U583  ( .A(1'b1), .ZN(_u0_u24_pointer[30] ) );
INV_X4 _u0_u24_U581  ( .A(1'b1), .ZN(_u0_u24_pointer[29] ) );
INV_X4 _u0_u24_U579  ( .A(1'b1), .ZN(_u0_u24_pointer[28] ) );
INV_X4 _u0_u24_U577  ( .A(1'b1), .ZN(_u0_u24_pointer[27] ) );
INV_X4 _u0_u24_U575  ( .A(1'b1), .ZN(_u0_u24_pointer[26] ) );
INV_X4 _u0_u24_U573  ( .A(1'b1), .ZN(_u0_u24_pointer[25] ) );
INV_X4 _u0_u24_U571  ( .A(1'b1), .ZN(_u0_u24_pointer[24] ) );
INV_X4 _u0_u24_U569  ( .A(1'b1), .ZN(_u0_u24_pointer[23] ) );
INV_X4 _u0_u24_U567  ( .A(1'b1), .ZN(_u0_u24_pointer[22] ) );
INV_X4 _u0_u24_U565  ( .A(1'b1), .ZN(_u0_u24_pointer[21] ) );
INV_X4 _u0_u24_U563  ( .A(1'b1), .ZN(_u0_u24_pointer[20] ) );
INV_X4 _u0_u24_U561  ( .A(1'b1), .ZN(_u0_u24_pointer[19] ) );
INV_X4 _u0_u24_U559  ( .A(1'b1), .ZN(_u0_u24_pointer[18] ) );
INV_X4 _u0_u24_U557  ( .A(1'b1), .ZN(_u0_u24_pointer[17] ) );
INV_X4 _u0_u24_U555  ( .A(1'b1), .ZN(_u0_u24_pointer[16] ) );
INV_X4 _u0_u24_U553  ( .A(1'b1), .ZN(_u0_u24_pointer[15] ) );
INV_X4 _u0_u24_U551  ( .A(1'b1), .ZN(_u0_u24_pointer[14] ) );
INV_X4 _u0_u24_U549  ( .A(1'b1), .ZN(_u0_u24_pointer[13] ) );
INV_X4 _u0_u24_U547  ( .A(1'b1), .ZN(_u0_u24_pointer[12] ) );
INV_X4 _u0_u24_U545  ( .A(1'b1), .ZN(_u0_u24_pointer[11] ) );
INV_X4 _u0_u24_U543  ( .A(1'b1), .ZN(_u0_u24_pointer[10] ) );
INV_X4 _u0_u24_U541  ( .A(1'b1), .ZN(_u0_u24_pointer[9] ) );
INV_X4 _u0_u24_U539  ( .A(1'b1), .ZN(_u0_u24_pointer[8] ) );
INV_X4 _u0_u24_U537  ( .A(1'b1), .ZN(_u0_u24_pointer[7] ) );
INV_X4 _u0_u24_U535  ( .A(1'b1), .ZN(_u0_u24_pointer[6] ) );
INV_X4 _u0_u24_U533  ( .A(1'b1), .ZN(_u0_u24_pointer[5] ) );
INV_X4 _u0_u24_U531  ( .A(1'b1), .ZN(_u0_u24_pointer[4] ) );
INV_X4 _u0_u24_U529  ( .A(1'b1), .ZN(_u0_u24_pointer[3] ) );
INV_X4 _u0_u24_U527  ( .A(1'b1), .ZN(_u0_u24_pointer[2] ) );
INV_X4 _u0_u24_U525  ( .A(1'b1), .ZN(_u0_u24_pointer[1] ) );
INV_X4 _u0_u24_U523  ( .A(1'b1), .ZN(_u0_u24_pointer[0] ) );
INV_X4 _u0_u24_U521  ( .A(1'b1), .ZN(_u0_u24_pointer_s[31] ) );
INV_X4 _u0_u24_U519  ( .A(1'b1), .ZN(_u0_u24_pointer_s[30] ) );
INV_X4 _u0_u24_U517  ( .A(1'b1), .ZN(_u0_u24_pointer_s[29] ) );
INV_X4 _u0_u24_U515  ( .A(1'b1), .ZN(_u0_u24_pointer_s[28] ) );
INV_X4 _u0_u24_U513  ( .A(1'b1), .ZN(_u0_u24_pointer_s[27] ) );
INV_X4 _u0_u24_U511  ( .A(1'b1), .ZN(_u0_u24_pointer_s[26] ) );
INV_X4 _u0_u24_U509  ( .A(1'b1), .ZN(_u0_u24_pointer_s[25] ) );
INV_X4 _u0_u24_U507  ( .A(1'b1), .ZN(_u0_u24_pointer_s[24] ) );
INV_X4 _u0_u24_U505  ( .A(1'b1), .ZN(_u0_u24_pointer_s[23] ) );
INV_X4 _u0_u24_U503  ( .A(1'b1), .ZN(_u0_u24_pointer_s[22] ) );
INV_X4 _u0_u24_U501  ( .A(1'b1), .ZN(_u0_u24_pointer_s[21] ) );
INV_X4 _u0_u24_U499  ( .A(1'b1), .ZN(_u0_u24_pointer_s[20] ) );
INV_X4 _u0_u24_U497  ( .A(1'b1), .ZN(_u0_u24_pointer_s[19] ) );
INV_X4 _u0_u24_U495  ( .A(1'b1), .ZN(_u0_u24_pointer_s[18] ) );
INV_X4 _u0_u24_U493  ( .A(1'b1), .ZN(_u0_u24_pointer_s[17] ) );
INV_X4 _u0_u24_U491  ( .A(1'b1), .ZN(_u0_u24_pointer_s[16] ) );
INV_X4 _u0_u24_U489  ( .A(1'b1), .ZN(_u0_u24_pointer_s[15] ) );
INV_X4 _u0_u24_U487  ( .A(1'b1), .ZN(_u0_u24_pointer_s[14] ) );
INV_X4 _u0_u24_U485  ( .A(1'b1), .ZN(_u0_u24_pointer_s[13] ) );
INV_X4 _u0_u24_U483  ( .A(1'b1), .ZN(_u0_u24_pointer_s[12] ) );
INV_X4 _u0_u24_U481  ( .A(1'b1), .ZN(_u0_u24_pointer_s[11] ) );
INV_X4 _u0_u24_U479  ( .A(1'b1), .ZN(_u0_u24_pointer_s[10] ) );
INV_X4 _u0_u24_U477  ( .A(1'b1), .ZN(_u0_u24_pointer_s[9] ) );
INV_X4 _u0_u24_U475  ( .A(1'b1), .ZN(_u0_u24_pointer_s[8] ) );
INV_X4 _u0_u24_U473  ( .A(1'b1), .ZN(_u0_u24_pointer_s[7] ) );
INV_X4 _u0_u24_U471  ( .A(1'b1), .ZN(_u0_u24_pointer_s[6] ) );
INV_X4 _u0_u24_U469  ( .A(1'b1), .ZN(_u0_u24_pointer_s[5] ) );
INV_X4 _u0_u24_U467  ( .A(1'b1), .ZN(_u0_u24_pointer_s[4] ) );
INV_X4 _u0_u24_U465  ( .A(1'b1), .ZN(_u0_u24_pointer_s[3] ) );
INV_X4 _u0_u24_U463  ( .A(1'b1), .ZN(_u0_u24_pointer_s[2] ) );
INV_X4 _u0_u24_U461  ( .A(1'b1), .ZN(_u0_u24_pointer_s[1] ) );
INV_X4 _u0_u24_U459  ( .A(1'b1), .ZN(_u0_u24_pointer_s[0] ) );
INV_X4 _u0_u24_U457  ( .A(1'b1), .ZN(_u0_u24_ch_csr[31] ) );
INV_X4 _u0_u24_U455  ( .A(1'b1), .ZN(_u0_u24_ch_csr[30] ) );
INV_X4 _u0_u24_U453  ( .A(1'b1), .ZN(_u0_u24_ch_csr[29] ) );
INV_X4 _u0_u24_U451  ( .A(1'b1), .ZN(_u0_u24_ch_csr[28] ) );
INV_X4 _u0_u24_U449  ( .A(1'b1), .ZN(_u0_u24_ch_csr[27] ) );
INV_X4 _u0_u24_U447  ( .A(1'b1), .ZN(_u0_u24_ch_csr[26] ) );
INV_X4 _u0_u24_U445  ( .A(1'b1), .ZN(_u0_u24_ch_csr[25] ) );
INV_X4 _u0_u24_U443  ( .A(1'b1), .ZN(_u0_u24_ch_csr[24] ) );
INV_X4 _u0_u24_U441  ( .A(1'b1), .ZN(_u0_u24_ch_csr[23] ) );
INV_X4 _u0_u24_U439  ( .A(1'b1), .ZN(_u0_u24_ch_csr[22] ) );
INV_X4 _u0_u24_U437  ( .A(1'b1), .ZN(_u0_u24_ch_csr[21] ) );
INV_X4 _u0_u24_U435  ( .A(1'b1), .ZN(_u0_u24_ch_csr[20] ) );
INV_X4 _u0_u24_U433  ( .A(1'b1), .ZN(_u0_u24_ch_csr[19] ) );
INV_X4 _u0_u24_U431  ( .A(1'b1), .ZN(_u0_u24_ch_csr[18] ) );
INV_X4 _u0_u24_U429  ( .A(1'b1), .ZN(_u0_u24_ch_csr[17] ) );
INV_X4 _u0_u24_U427  ( .A(1'b1), .ZN(_u0_u24_ch_csr[16] ) );
INV_X4 _u0_u24_U425  ( .A(1'b1), .ZN(_u0_u24_ch_csr[15] ) );
INV_X4 _u0_u24_U423  ( .A(1'b1), .ZN(_u0_u24_ch_csr[14] ) );
INV_X4 _u0_u24_U421  ( .A(1'b1), .ZN(_u0_u24_ch_csr[13] ) );
INV_X4 _u0_u24_U419  ( .A(1'b1), .ZN(_u0_u24_ch_csr[12] ) );
INV_X4 _u0_u24_U417  ( .A(1'b1), .ZN(_u0_u24_ch_csr[11] ) );
INV_X4 _u0_u24_U415  ( .A(1'b1), .ZN(_u0_u24_ch_csr[10] ) );
INV_X4 _u0_u24_U413  ( .A(1'b1), .ZN(_u0_u24_ch_csr[9] ) );
INV_X4 _u0_u24_U411  ( .A(1'b1), .ZN(_u0_u24_ch_csr[8] ) );
INV_X4 _u0_u24_U409  ( .A(1'b1), .ZN(_u0_u24_ch_csr[7] ) );
INV_X4 _u0_u24_U407  ( .A(1'b1), .ZN(_u0_u24_ch_csr[6] ) );
INV_X4 _u0_u24_U405  ( .A(1'b1), .ZN(_u0_u24_ch_csr[5] ) );
INV_X4 _u0_u24_U403  ( .A(1'b1), .ZN(_u0_u24_ch_csr[4] ) );
INV_X4 _u0_u24_U401  ( .A(1'b1), .ZN(_u0_u24_ch_csr[3] ) );
INV_X4 _u0_u24_U399  ( .A(1'b1), .ZN(_u0_u24_ch_csr[2] ) );
INV_X4 _u0_u24_U397  ( .A(1'b1), .ZN(_u0_u24_ch_csr[1] ) );
INV_X4 _u0_u24_U395  ( .A(1'b1), .ZN(_u0_u24_ch_csr[0] ) );
INV_X4 _u0_u24_U393  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[31] ) );
INV_X4 _u0_u24_U391  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[30] ) );
INV_X4 _u0_u24_U389  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[29] ) );
INV_X4 _u0_u24_U387  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[28] ) );
INV_X4 _u0_u24_U385  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[27] ) );
INV_X4 _u0_u24_U383  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[26] ) );
INV_X4 _u0_u24_U381  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[25] ) );
INV_X4 _u0_u24_U379  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[24] ) );
INV_X4 _u0_u24_U377  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[23] ) );
INV_X4 _u0_u24_U375  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[22] ) );
INV_X4 _u0_u24_U373  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[21] ) );
INV_X4 _u0_u24_U371  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[20] ) );
INV_X4 _u0_u24_U369  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[19] ) );
INV_X4 _u0_u24_U367  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[18] ) );
INV_X4 _u0_u24_U365  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[17] ) );
INV_X4 _u0_u24_U363  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[16] ) );
INV_X4 _u0_u24_U361  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[15] ) );
INV_X4 _u0_u24_U359  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[14] ) );
INV_X4 _u0_u24_U357  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[13] ) );
INV_X4 _u0_u24_U355  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[12] ) );
INV_X4 _u0_u24_U353  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[11] ) );
INV_X4 _u0_u24_U351  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[10] ) );
INV_X4 _u0_u24_U349  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[9] ) );
INV_X4 _u0_u24_U347  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[8] ) );
INV_X4 _u0_u24_U345  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[7] ) );
INV_X4 _u0_u24_U343  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[6] ) );
INV_X4 _u0_u24_U341  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[5] ) );
INV_X4 _u0_u24_U339  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[4] ) );
INV_X4 _u0_u24_U337  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[3] ) );
INV_X4 _u0_u24_U335  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[2] ) );
INV_X4 _u0_u24_U333  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[1] ) );
INV_X4 _u0_u24_U331  ( .A(1'b1), .ZN(_u0_u24_ch_txsz[0] ) );
INV_X4 _u0_u24_U329  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[31] ) );
INV_X4 _u0_u24_U327  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[30] ) );
INV_X4 _u0_u24_U325  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[29] ) );
INV_X4 _u0_u24_U323  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[28] ) );
INV_X4 _u0_u24_U321  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[27] ) );
INV_X4 _u0_u24_U319  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[26] ) );
INV_X4 _u0_u24_U317  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[25] ) );
INV_X4 _u0_u24_U315  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[24] ) );
INV_X4 _u0_u24_U313  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[23] ) );
INV_X4 _u0_u24_U311  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[22] ) );
INV_X4 _u0_u24_U309  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[21] ) );
INV_X4 _u0_u24_U307  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[20] ) );
INV_X4 _u0_u24_U305  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[19] ) );
INV_X4 _u0_u24_U303  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[18] ) );
INV_X4 _u0_u24_U301  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[17] ) );
INV_X4 _u0_u24_U299  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[16] ) );
INV_X4 _u0_u24_U297  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[15] ) );
INV_X4 _u0_u24_U295  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[14] ) );
INV_X4 _u0_u24_U293  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[13] ) );
INV_X4 _u0_u24_U291  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[12] ) );
INV_X4 _u0_u24_U289  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[11] ) );
INV_X4 _u0_u24_U287  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[10] ) );
INV_X4 _u0_u24_U285  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[9] ) );
INV_X4 _u0_u24_U283  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[8] ) );
INV_X4 _u0_u24_U281  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[7] ) );
INV_X4 _u0_u24_U279  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[6] ) );
INV_X4 _u0_u24_U277  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[5] ) );
INV_X4 _u0_u24_U275  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[4] ) );
INV_X4 _u0_u24_U273  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[3] ) );
INV_X4 _u0_u24_U271  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[2] ) );
INV_X4 _u0_u24_U269  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[1] ) );
INV_X4 _u0_u24_U267  ( .A(1'b1), .ZN(_u0_u24_ch_adr0[0] ) );
INV_X4 _u0_u24_U265  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[31] ) );
INV_X4 _u0_u24_U263  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[30] ) );
INV_X4 _u0_u24_U261  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[29] ) );
INV_X4 _u0_u24_U259  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[28] ) );
INV_X4 _u0_u24_U257  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[27] ) );
INV_X4 _u0_u24_U255  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[26] ) );
INV_X4 _u0_u24_U253  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[25] ) );
INV_X4 _u0_u24_U251  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[24] ) );
INV_X4 _u0_u24_U249  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[23] ) );
INV_X4 _u0_u24_U247  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[22] ) );
INV_X4 _u0_u24_U245  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[21] ) );
INV_X4 _u0_u24_U243  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[20] ) );
INV_X4 _u0_u24_U241  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[19] ) );
INV_X4 _u0_u24_U239  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[18] ) );
INV_X4 _u0_u24_U237  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[17] ) );
INV_X4 _u0_u24_U235  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[16] ) );
INV_X4 _u0_u24_U233  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[15] ) );
INV_X4 _u0_u24_U231  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[14] ) );
INV_X4 _u0_u24_U229  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[13] ) );
INV_X4 _u0_u24_U227  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[12] ) );
INV_X4 _u0_u24_U225  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[11] ) );
INV_X4 _u0_u24_U223  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[10] ) );
INV_X4 _u0_u24_U221  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[9] ) );
INV_X4 _u0_u24_U219  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[8] ) );
INV_X4 _u0_u24_U217  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[7] ) );
INV_X4 _u0_u24_U215  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[6] ) );
INV_X4 _u0_u24_U213  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[5] ) );
INV_X4 _u0_u24_U211  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[4] ) );
INV_X4 _u0_u24_U209  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[3] ) );
INV_X4 _u0_u24_U207  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[2] ) );
INV_X4 _u0_u24_U205  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[1] ) );
INV_X4 _u0_u24_U203  ( .A(1'b1), .ZN(_u0_u24_ch_adr1[0] ) );
INV_X4 _u0_u24_U201  ( .A(1'b0), .ZN(_u0_u24_ch_am0[31] ) );
INV_X4 _u0_u24_U199  ( .A(1'b0), .ZN(_u0_u24_ch_am0[30] ) );
INV_X4 _u0_u24_U197  ( .A(1'b0), .ZN(_u0_u24_ch_am0[29] ) );
INV_X4 _u0_u24_U195  ( .A(1'b0), .ZN(_u0_u24_ch_am0[28] ) );
INV_X4 _u0_u24_U193  ( .A(1'b0), .ZN(_u0_u24_ch_am0[27] ) );
INV_X4 _u0_u24_U191  ( .A(1'b0), .ZN(_u0_u24_ch_am0[26] ) );
INV_X4 _u0_u24_U189  ( .A(1'b0), .ZN(_u0_u24_ch_am0[25] ) );
INV_X4 _u0_u24_U187  ( .A(1'b0), .ZN(_u0_u24_ch_am0[24] ) );
INV_X4 _u0_u24_U185  ( .A(1'b0), .ZN(_u0_u24_ch_am0[23] ) );
INV_X4 _u0_u24_U183  ( .A(1'b0), .ZN(_u0_u24_ch_am0[22] ) );
INV_X4 _u0_u24_U181  ( .A(1'b0), .ZN(_u0_u24_ch_am0[21] ) );
INV_X4 _u0_u24_U179  ( .A(1'b0), .ZN(_u0_u24_ch_am0[20] ) );
INV_X4 _u0_u24_U177  ( .A(1'b0), .ZN(_u0_u24_ch_am0[19] ) );
INV_X4 _u0_u24_U175  ( .A(1'b0), .ZN(_u0_u24_ch_am0[18] ) );
INV_X4 _u0_u24_U173  ( .A(1'b0), .ZN(_u0_u24_ch_am0[17] ) );
INV_X4 _u0_u24_U171  ( .A(1'b0), .ZN(_u0_u24_ch_am0[16] ) );
INV_X4 _u0_u24_U169  ( .A(1'b0), .ZN(_u0_u24_ch_am0[15] ) );
INV_X4 _u0_u24_U167  ( .A(1'b0), .ZN(_u0_u24_ch_am0[14] ) );
INV_X4 _u0_u24_U165  ( .A(1'b0), .ZN(_u0_u24_ch_am0[13] ) );
INV_X4 _u0_u24_U163  ( .A(1'b0), .ZN(_u0_u24_ch_am0[12] ) );
INV_X4 _u0_u24_U161  ( .A(1'b0), .ZN(_u0_u24_ch_am0[11] ) );
INV_X4 _u0_u24_U159  ( .A(1'b0), .ZN(_u0_u24_ch_am0[10] ) );
INV_X4 _u0_u24_U157  ( .A(1'b0), .ZN(_u0_u24_ch_am0[9] ) );
INV_X4 _u0_u24_U155  ( .A(1'b0), .ZN(_u0_u24_ch_am0[8] ) );
INV_X4 _u0_u24_U153  ( .A(1'b0), .ZN(_u0_u24_ch_am0[7] ) );
INV_X4 _u0_u24_U151  ( .A(1'b0), .ZN(_u0_u24_ch_am0[6] ) );
INV_X4 _u0_u24_U149  ( .A(1'b0), .ZN(_u0_u24_ch_am0[5] ) );
INV_X4 _u0_u24_U147  ( .A(1'b0), .ZN(_u0_u24_ch_am0[4] ) );
INV_X4 _u0_u24_U145  ( .A(1'b1), .ZN(_u0_u24_ch_am0[3] ) );
INV_X4 _u0_u24_U143  ( .A(1'b1), .ZN(_u0_u24_ch_am0[2] ) );
INV_X4 _u0_u24_U141  ( .A(1'b1), .ZN(_u0_u24_ch_am0[1] ) );
INV_X4 _u0_u24_U139  ( .A(1'b1), .ZN(_u0_u24_ch_am0[0] ) );
INV_X4 _u0_u24_U137  ( .A(1'b0), .ZN(_u0_u24_ch_am1[31] ) );
INV_X4 _u0_u24_U135  ( .A(1'b0), .ZN(_u0_u24_ch_am1[30] ) );
INV_X4 _u0_u24_U133  ( .A(1'b0), .ZN(_u0_u24_ch_am1[29] ) );
INV_X4 _u0_u24_U131  ( .A(1'b0), .ZN(_u0_u24_ch_am1[28] ) );
INV_X4 _u0_u24_U129  ( .A(1'b0), .ZN(_u0_u24_ch_am1[27] ) );
INV_X4 _u0_u24_U127  ( .A(1'b0), .ZN(_u0_u24_ch_am1[26] ) );
INV_X4 _u0_u24_U125  ( .A(1'b0), .ZN(_u0_u24_ch_am1[25] ) );
INV_X4 _u0_u24_U123  ( .A(1'b0), .ZN(_u0_u24_ch_am1[24] ) );
INV_X4 _u0_u24_U121  ( .A(1'b0), .ZN(_u0_u24_ch_am1[23] ) );
INV_X4 _u0_u24_U119  ( .A(1'b0), .ZN(_u0_u24_ch_am1[22] ) );
INV_X4 _u0_u24_U117  ( .A(1'b0), .ZN(_u0_u24_ch_am1[21] ) );
INV_X4 _u0_u24_U115  ( .A(1'b0), .ZN(_u0_u24_ch_am1[20] ) );
INV_X4 _u0_u24_U113  ( .A(1'b0), .ZN(_u0_u24_ch_am1[19] ) );
INV_X4 _u0_u24_U111  ( .A(1'b0), .ZN(_u0_u24_ch_am1[18] ) );
INV_X4 _u0_u24_U109  ( .A(1'b0), .ZN(_u0_u24_ch_am1[17] ) );
INV_X4 _u0_u24_U107  ( .A(1'b0), .ZN(_u0_u24_ch_am1[16] ) );
INV_X4 _u0_u24_U105  ( .A(1'b0), .ZN(_u0_u24_ch_am1[15] ) );
INV_X4 _u0_u24_U103  ( .A(1'b0), .ZN(_u0_u24_ch_am1[14] ) );
INV_X4 _u0_u24_U101  ( .A(1'b0), .ZN(_u0_u24_ch_am1[13] ) );
INV_X4 _u0_u24_U99  ( .A(1'b0), .ZN(_u0_u24_ch_am1[12] ) );
INV_X4 _u0_u24_U97  ( .A(1'b0), .ZN(_u0_u24_ch_am1[11] ) );
INV_X4 _u0_u24_U95  ( .A(1'b0), .ZN(_u0_u24_ch_am1[10] ) );
INV_X4 _u0_u24_U93  ( .A(1'b0), .ZN(_u0_u24_ch_am1[9] ) );
INV_X4 _u0_u24_U91  ( .A(1'b0), .ZN(_u0_u24_ch_am1[8] ) );
INV_X4 _u0_u24_U89  ( .A(1'b0), .ZN(_u0_u24_ch_am1[7] ) );
INV_X4 _u0_u24_U87  ( .A(1'b0), .ZN(_u0_u24_ch_am1[6] ) );
INV_X4 _u0_u24_U85  ( .A(1'b0), .ZN(_u0_u24_ch_am1[5] ) );
INV_X4 _u0_u24_U83  ( .A(1'b0), .ZN(_u0_u24_ch_am1[4] ) );
INV_X4 _u0_u24_U81  ( .A(1'b1), .ZN(_u0_u24_ch_am1[3] ) );
INV_X4 _u0_u24_U79  ( .A(1'b1), .ZN(_u0_u24_ch_am1[2] ) );
INV_X4 _u0_u24_U77  ( .A(1'b1), .ZN(_u0_u24_ch_am1[1] ) );
INV_X4 _u0_u24_U75  ( .A(1'b1), .ZN(_u0_u24_ch_am1[0] ) );
INV_X4 _u0_u24_U73  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[31] ) );
INV_X4 _u0_u24_U71  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[30] ) );
INV_X4 _u0_u24_U69  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[29] ) );
INV_X4 _u0_u24_U67  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[28] ) );
INV_X4 _u0_u24_U65  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[27] ) );
INV_X4 _u0_u24_U63  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[26] ) );
INV_X4 _u0_u24_U61  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[25] ) );
INV_X4 _u0_u24_U59  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[24] ) );
INV_X4 _u0_u24_U57  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[23] ) );
INV_X4 _u0_u24_U55  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[22] ) );
INV_X4 _u0_u24_U53  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[21] ) );
INV_X4 _u0_u24_U51  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[20] ) );
INV_X4 _u0_u24_U49  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[19] ) );
INV_X4 _u0_u24_U47  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[18] ) );
INV_X4 _u0_u24_U45  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[17] ) );
INV_X4 _u0_u24_U43  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[16] ) );
INV_X4 _u0_u24_U41  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[15] ) );
INV_X4 _u0_u24_U39  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[14] ) );
INV_X4 _u0_u24_U37  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[13] ) );
INV_X4 _u0_u24_U35  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[12] ) );
INV_X4 _u0_u24_U33  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[11] ) );
INV_X4 _u0_u24_U31  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[10] ) );
INV_X4 _u0_u24_U29  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[9] ) );
INV_X4 _u0_u24_U27  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[8] ) );
INV_X4 _u0_u24_U25  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[7] ) );
INV_X4 _u0_u24_U23  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[6] ) );
INV_X4 _u0_u24_U21  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[5] ) );
INV_X4 _u0_u24_U19  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[4] ) );
INV_X4 _u0_u24_U17  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[3] ) );
INV_X4 _u0_u24_U15  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[2] ) );
INV_X4 _u0_u24_U13  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[1] ) );
INV_X4 _u0_u24_U11  ( .A(1'b1), .ZN(_u0_u24_sw_pointer[0] ) );
INV_X4 _u0_u24_U9  ( .A(1'b1), .ZN(_u0_u24_ch_stop ) );
INV_X4 _u0_u24_U7  ( .A(1'b1), .ZN(_u0_u24_ch_dis ) );
INV_X4 _u0_u24_U5  ( .A(1'b1), .ZN(_u0_u24_int ) );
INV_X4 _u0_u25_U585  ( .A(1'b1), .ZN(_u0_u25_pointer[31] ) );
INV_X4 _u0_u25_U583  ( .A(1'b1), .ZN(_u0_u25_pointer[30] ) );
INV_X4 _u0_u25_U581  ( .A(1'b1), .ZN(_u0_u25_pointer[29] ) );
INV_X4 _u0_u25_U579  ( .A(1'b1), .ZN(_u0_u25_pointer[28] ) );
INV_X4 _u0_u25_U577  ( .A(1'b1), .ZN(_u0_u25_pointer[27] ) );
INV_X4 _u0_u25_U575  ( .A(1'b1), .ZN(_u0_u25_pointer[26] ) );
INV_X4 _u0_u25_U573  ( .A(1'b1), .ZN(_u0_u25_pointer[25] ) );
INV_X4 _u0_u25_U571  ( .A(1'b1), .ZN(_u0_u25_pointer[24] ) );
INV_X4 _u0_u25_U569  ( .A(1'b1), .ZN(_u0_u25_pointer[23] ) );
INV_X4 _u0_u25_U567  ( .A(1'b1), .ZN(_u0_u25_pointer[22] ) );
INV_X4 _u0_u25_U565  ( .A(1'b1), .ZN(_u0_u25_pointer[21] ) );
INV_X4 _u0_u25_U563  ( .A(1'b1), .ZN(_u0_u25_pointer[20] ) );
INV_X4 _u0_u25_U561  ( .A(1'b1), .ZN(_u0_u25_pointer[19] ) );
INV_X4 _u0_u25_U559  ( .A(1'b1), .ZN(_u0_u25_pointer[18] ) );
INV_X4 _u0_u25_U557  ( .A(1'b1), .ZN(_u0_u25_pointer[17] ) );
INV_X4 _u0_u25_U555  ( .A(1'b1), .ZN(_u0_u25_pointer[16] ) );
INV_X4 _u0_u25_U553  ( .A(1'b1), .ZN(_u0_u25_pointer[15] ) );
INV_X4 _u0_u25_U551  ( .A(1'b1), .ZN(_u0_u25_pointer[14] ) );
INV_X4 _u0_u25_U549  ( .A(1'b1), .ZN(_u0_u25_pointer[13] ) );
INV_X4 _u0_u25_U547  ( .A(1'b1), .ZN(_u0_u25_pointer[12] ) );
INV_X4 _u0_u25_U545  ( .A(1'b1), .ZN(_u0_u25_pointer[11] ) );
INV_X4 _u0_u25_U543  ( .A(1'b1), .ZN(_u0_u25_pointer[10] ) );
INV_X4 _u0_u25_U541  ( .A(1'b1), .ZN(_u0_u25_pointer[9] ) );
INV_X4 _u0_u25_U539  ( .A(1'b1), .ZN(_u0_u25_pointer[8] ) );
INV_X4 _u0_u25_U537  ( .A(1'b1), .ZN(_u0_u25_pointer[7] ) );
INV_X4 _u0_u25_U535  ( .A(1'b1), .ZN(_u0_u25_pointer[6] ) );
INV_X4 _u0_u25_U533  ( .A(1'b1), .ZN(_u0_u25_pointer[5] ) );
INV_X4 _u0_u25_U531  ( .A(1'b1), .ZN(_u0_u25_pointer[4] ) );
INV_X4 _u0_u25_U529  ( .A(1'b1), .ZN(_u0_u25_pointer[3] ) );
INV_X4 _u0_u25_U527  ( .A(1'b1), .ZN(_u0_u25_pointer[2] ) );
INV_X4 _u0_u25_U525  ( .A(1'b1), .ZN(_u0_u25_pointer[1] ) );
INV_X4 _u0_u25_U523  ( .A(1'b1), .ZN(_u0_u25_pointer[0] ) );
INV_X4 _u0_u25_U521  ( .A(1'b1), .ZN(_u0_u25_pointer_s[31] ) );
INV_X4 _u0_u25_U519  ( .A(1'b1), .ZN(_u0_u25_pointer_s[30] ) );
INV_X4 _u0_u25_U517  ( .A(1'b1), .ZN(_u0_u25_pointer_s[29] ) );
INV_X4 _u0_u25_U515  ( .A(1'b1), .ZN(_u0_u25_pointer_s[28] ) );
INV_X4 _u0_u25_U513  ( .A(1'b1), .ZN(_u0_u25_pointer_s[27] ) );
INV_X4 _u0_u25_U511  ( .A(1'b1), .ZN(_u0_u25_pointer_s[26] ) );
INV_X4 _u0_u25_U509  ( .A(1'b1), .ZN(_u0_u25_pointer_s[25] ) );
INV_X4 _u0_u25_U507  ( .A(1'b1), .ZN(_u0_u25_pointer_s[24] ) );
INV_X4 _u0_u25_U505  ( .A(1'b1), .ZN(_u0_u25_pointer_s[23] ) );
INV_X4 _u0_u25_U503  ( .A(1'b1), .ZN(_u0_u25_pointer_s[22] ) );
INV_X4 _u0_u25_U501  ( .A(1'b1), .ZN(_u0_u25_pointer_s[21] ) );
INV_X4 _u0_u25_U499  ( .A(1'b1), .ZN(_u0_u25_pointer_s[20] ) );
INV_X4 _u0_u25_U497  ( .A(1'b1), .ZN(_u0_u25_pointer_s[19] ) );
INV_X4 _u0_u25_U495  ( .A(1'b1), .ZN(_u0_u25_pointer_s[18] ) );
INV_X4 _u0_u25_U493  ( .A(1'b1), .ZN(_u0_u25_pointer_s[17] ) );
INV_X4 _u0_u25_U491  ( .A(1'b1), .ZN(_u0_u25_pointer_s[16] ) );
INV_X4 _u0_u25_U489  ( .A(1'b1), .ZN(_u0_u25_pointer_s[15] ) );
INV_X4 _u0_u25_U487  ( .A(1'b1), .ZN(_u0_u25_pointer_s[14] ) );
INV_X4 _u0_u25_U485  ( .A(1'b1), .ZN(_u0_u25_pointer_s[13] ) );
INV_X4 _u0_u25_U483  ( .A(1'b1), .ZN(_u0_u25_pointer_s[12] ) );
INV_X4 _u0_u25_U481  ( .A(1'b1), .ZN(_u0_u25_pointer_s[11] ) );
INV_X4 _u0_u25_U479  ( .A(1'b1), .ZN(_u0_u25_pointer_s[10] ) );
INV_X4 _u0_u25_U477  ( .A(1'b1), .ZN(_u0_u25_pointer_s[9] ) );
INV_X4 _u0_u25_U475  ( .A(1'b1), .ZN(_u0_u25_pointer_s[8] ) );
INV_X4 _u0_u25_U473  ( .A(1'b1), .ZN(_u0_u25_pointer_s[7] ) );
INV_X4 _u0_u25_U471  ( .A(1'b1), .ZN(_u0_u25_pointer_s[6] ) );
INV_X4 _u0_u25_U469  ( .A(1'b1), .ZN(_u0_u25_pointer_s[5] ) );
INV_X4 _u0_u25_U467  ( .A(1'b1), .ZN(_u0_u25_pointer_s[4] ) );
INV_X4 _u0_u25_U465  ( .A(1'b1), .ZN(_u0_u25_pointer_s[3] ) );
INV_X4 _u0_u25_U463  ( .A(1'b1), .ZN(_u0_u25_pointer_s[2] ) );
INV_X4 _u0_u25_U461  ( .A(1'b1), .ZN(_u0_u25_pointer_s[1] ) );
INV_X4 _u0_u25_U459  ( .A(1'b1), .ZN(_u0_u25_pointer_s[0] ) );
INV_X4 _u0_u25_U457  ( .A(1'b1), .ZN(_u0_u25_ch_csr[31] ) );
INV_X4 _u0_u25_U455  ( .A(1'b1), .ZN(_u0_u25_ch_csr[30] ) );
INV_X4 _u0_u25_U453  ( .A(1'b1), .ZN(_u0_u25_ch_csr[29] ) );
INV_X4 _u0_u25_U451  ( .A(1'b1), .ZN(_u0_u25_ch_csr[28] ) );
INV_X4 _u0_u25_U449  ( .A(1'b1), .ZN(_u0_u25_ch_csr[27] ) );
INV_X4 _u0_u25_U447  ( .A(1'b1), .ZN(_u0_u25_ch_csr[26] ) );
INV_X4 _u0_u25_U445  ( .A(1'b1), .ZN(_u0_u25_ch_csr[25] ) );
INV_X4 _u0_u25_U443  ( .A(1'b1), .ZN(_u0_u25_ch_csr[24] ) );
INV_X4 _u0_u25_U441  ( .A(1'b1), .ZN(_u0_u25_ch_csr[23] ) );
INV_X4 _u0_u25_U439  ( .A(1'b1), .ZN(_u0_u25_ch_csr[22] ) );
INV_X4 _u0_u25_U437  ( .A(1'b1), .ZN(_u0_u25_ch_csr[21] ) );
INV_X4 _u0_u25_U435  ( .A(1'b1), .ZN(_u0_u25_ch_csr[20] ) );
INV_X4 _u0_u25_U433  ( .A(1'b1), .ZN(_u0_u25_ch_csr[19] ) );
INV_X4 _u0_u25_U431  ( .A(1'b1), .ZN(_u0_u25_ch_csr[18] ) );
INV_X4 _u0_u25_U429  ( .A(1'b1), .ZN(_u0_u25_ch_csr[17] ) );
INV_X4 _u0_u25_U427  ( .A(1'b1), .ZN(_u0_u25_ch_csr[16] ) );
INV_X4 _u0_u25_U425  ( .A(1'b1), .ZN(_u0_u25_ch_csr[15] ) );
INV_X4 _u0_u25_U423  ( .A(1'b1), .ZN(_u0_u25_ch_csr[14] ) );
INV_X4 _u0_u25_U421  ( .A(1'b1), .ZN(_u0_u25_ch_csr[13] ) );
INV_X4 _u0_u25_U419  ( .A(1'b1), .ZN(_u0_u25_ch_csr[12] ) );
INV_X4 _u0_u25_U417  ( .A(1'b1), .ZN(_u0_u25_ch_csr[11] ) );
INV_X4 _u0_u25_U415  ( .A(1'b1), .ZN(_u0_u25_ch_csr[10] ) );
INV_X4 _u0_u25_U413  ( .A(1'b1), .ZN(_u0_u25_ch_csr[9] ) );
INV_X4 _u0_u25_U411  ( .A(1'b1), .ZN(_u0_u25_ch_csr[8] ) );
INV_X4 _u0_u25_U409  ( .A(1'b1), .ZN(_u0_u25_ch_csr[7] ) );
INV_X4 _u0_u25_U407  ( .A(1'b1), .ZN(_u0_u25_ch_csr[6] ) );
INV_X4 _u0_u25_U405  ( .A(1'b1), .ZN(_u0_u25_ch_csr[5] ) );
INV_X4 _u0_u25_U403  ( .A(1'b1), .ZN(_u0_u25_ch_csr[4] ) );
INV_X4 _u0_u25_U401  ( .A(1'b1), .ZN(_u0_u25_ch_csr[3] ) );
INV_X4 _u0_u25_U399  ( .A(1'b1), .ZN(_u0_u25_ch_csr[2] ) );
INV_X4 _u0_u25_U397  ( .A(1'b1), .ZN(_u0_u25_ch_csr[1] ) );
INV_X4 _u0_u25_U395  ( .A(1'b1), .ZN(_u0_u25_ch_csr[0] ) );
INV_X4 _u0_u25_U393  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[31] ) );
INV_X4 _u0_u25_U391  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[30] ) );
INV_X4 _u0_u25_U389  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[29] ) );
INV_X4 _u0_u25_U387  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[28] ) );
INV_X4 _u0_u25_U385  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[27] ) );
INV_X4 _u0_u25_U383  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[26] ) );
INV_X4 _u0_u25_U381  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[25] ) );
INV_X4 _u0_u25_U379  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[24] ) );
INV_X4 _u0_u25_U377  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[23] ) );
INV_X4 _u0_u25_U375  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[22] ) );
INV_X4 _u0_u25_U373  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[21] ) );
INV_X4 _u0_u25_U371  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[20] ) );
INV_X4 _u0_u25_U369  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[19] ) );
INV_X4 _u0_u25_U367  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[18] ) );
INV_X4 _u0_u25_U365  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[17] ) );
INV_X4 _u0_u25_U363  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[16] ) );
INV_X4 _u0_u25_U361  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[15] ) );
INV_X4 _u0_u25_U359  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[14] ) );
INV_X4 _u0_u25_U357  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[13] ) );
INV_X4 _u0_u25_U355  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[12] ) );
INV_X4 _u0_u25_U353  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[11] ) );
INV_X4 _u0_u25_U351  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[10] ) );
INV_X4 _u0_u25_U349  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[9] ) );
INV_X4 _u0_u25_U347  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[8] ) );
INV_X4 _u0_u25_U345  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[7] ) );
INV_X4 _u0_u25_U343  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[6] ) );
INV_X4 _u0_u25_U341  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[5] ) );
INV_X4 _u0_u25_U339  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[4] ) );
INV_X4 _u0_u25_U337  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[3] ) );
INV_X4 _u0_u25_U335  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[2] ) );
INV_X4 _u0_u25_U333  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[1] ) );
INV_X4 _u0_u25_U331  ( .A(1'b1), .ZN(_u0_u25_ch_txsz[0] ) );
INV_X4 _u0_u25_U329  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[31] ) );
INV_X4 _u0_u25_U327  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[30] ) );
INV_X4 _u0_u25_U325  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[29] ) );
INV_X4 _u0_u25_U323  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[28] ) );
INV_X4 _u0_u25_U321  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[27] ) );
INV_X4 _u0_u25_U319  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[26] ) );
INV_X4 _u0_u25_U317  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[25] ) );
INV_X4 _u0_u25_U315  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[24] ) );
INV_X4 _u0_u25_U313  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[23] ) );
INV_X4 _u0_u25_U311  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[22] ) );
INV_X4 _u0_u25_U309  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[21] ) );
INV_X4 _u0_u25_U307  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[20] ) );
INV_X4 _u0_u25_U305  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[19] ) );
INV_X4 _u0_u25_U303  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[18] ) );
INV_X4 _u0_u25_U301  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[17] ) );
INV_X4 _u0_u25_U299  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[16] ) );
INV_X4 _u0_u25_U297  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[15] ) );
INV_X4 _u0_u25_U295  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[14] ) );
INV_X4 _u0_u25_U293  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[13] ) );
INV_X4 _u0_u25_U291  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[12] ) );
INV_X4 _u0_u25_U289  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[11] ) );
INV_X4 _u0_u25_U287  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[10] ) );
INV_X4 _u0_u25_U285  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[9] ) );
INV_X4 _u0_u25_U283  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[8] ) );
INV_X4 _u0_u25_U281  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[7] ) );
INV_X4 _u0_u25_U279  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[6] ) );
INV_X4 _u0_u25_U277  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[5] ) );
INV_X4 _u0_u25_U275  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[4] ) );
INV_X4 _u0_u25_U273  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[3] ) );
INV_X4 _u0_u25_U271  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[2] ) );
INV_X4 _u0_u25_U269  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[1] ) );
INV_X4 _u0_u25_U267  ( .A(1'b1), .ZN(_u0_u25_ch_adr0[0] ) );
INV_X4 _u0_u25_U265  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[31] ) );
INV_X4 _u0_u25_U263  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[30] ) );
INV_X4 _u0_u25_U261  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[29] ) );
INV_X4 _u0_u25_U259  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[28] ) );
INV_X4 _u0_u25_U257  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[27] ) );
INV_X4 _u0_u25_U255  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[26] ) );
INV_X4 _u0_u25_U253  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[25] ) );
INV_X4 _u0_u25_U251  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[24] ) );
INV_X4 _u0_u25_U249  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[23] ) );
INV_X4 _u0_u25_U247  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[22] ) );
INV_X4 _u0_u25_U245  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[21] ) );
INV_X4 _u0_u25_U243  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[20] ) );
INV_X4 _u0_u25_U241  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[19] ) );
INV_X4 _u0_u25_U239  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[18] ) );
INV_X4 _u0_u25_U237  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[17] ) );
INV_X4 _u0_u25_U235  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[16] ) );
INV_X4 _u0_u25_U233  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[15] ) );
INV_X4 _u0_u25_U231  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[14] ) );
INV_X4 _u0_u25_U229  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[13] ) );
INV_X4 _u0_u25_U227  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[12] ) );
INV_X4 _u0_u25_U225  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[11] ) );
INV_X4 _u0_u25_U223  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[10] ) );
INV_X4 _u0_u25_U221  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[9] ) );
INV_X4 _u0_u25_U219  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[8] ) );
INV_X4 _u0_u25_U217  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[7] ) );
INV_X4 _u0_u25_U215  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[6] ) );
INV_X4 _u0_u25_U213  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[5] ) );
INV_X4 _u0_u25_U211  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[4] ) );
INV_X4 _u0_u25_U209  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[3] ) );
INV_X4 _u0_u25_U207  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[2] ) );
INV_X4 _u0_u25_U205  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[1] ) );
INV_X4 _u0_u25_U203  ( .A(1'b1), .ZN(_u0_u25_ch_adr1[0] ) );
INV_X4 _u0_u25_U201  ( .A(1'b0), .ZN(_u0_u25_ch_am0[31] ) );
INV_X4 _u0_u25_U199  ( .A(1'b0), .ZN(_u0_u25_ch_am0[30] ) );
INV_X4 _u0_u25_U197  ( .A(1'b0), .ZN(_u0_u25_ch_am0[29] ) );
INV_X4 _u0_u25_U195  ( .A(1'b0), .ZN(_u0_u25_ch_am0[28] ) );
INV_X4 _u0_u25_U193  ( .A(1'b0), .ZN(_u0_u25_ch_am0[27] ) );
INV_X4 _u0_u25_U191  ( .A(1'b0), .ZN(_u0_u25_ch_am0[26] ) );
INV_X4 _u0_u25_U189  ( .A(1'b0), .ZN(_u0_u25_ch_am0[25] ) );
INV_X4 _u0_u25_U187  ( .A(1'b0), .ZN(_u0_u25_ch_am0[24] ) );
INV_X4 _u0_u25_U185  ( .A(1'b0), .ZN(_u0_u25_ch_am0[23] ) );
INV_X4 _u0_u25_U183  ( .A(1'b0), .ZN(_u0_u25_ch_am0[22] ) );
INV_X4 _u0_u25_U181  ( .A(1'b0), .ZN(_u0_u25_ch_am0[21] ) );
INV_X4 _u0_u25_U179  ( .A(1'b0), .ZN(_u0_u25_ch_am0[20] ) );
INV_X4 _u0_u25_U177  ( .A(1'b0), .ZN(_u0_u25_ch_am0[19] ) );
INV_X4 _u0_u25_U175  ( .A(1'b0), .ZN(_u0_u25_ch_am0[18] ) );
INV_X4 _u0_u25_U173  ( .A(1'b0), .ZN(_u0_u25_ch_am0[17] ) );
INV_X4 _u0_u25_U171  ( .A(1'b0), .ZN(_u0_u25_ch_am0[16] ) );
INV_X4 _u0_u25_U169  ( .A(1'b0), .ZN(_u0_u25_ch_am0[15] ) );
INV_X4 _u0_u25_U167  ( .A(1'b0), .ZN(_u0_u25_ch_am0[14] ) );
INV_X4 _u0_u25_U165  ( .A(1'b0), .ZN(_u0_u25_ch_am0[13] ) );
INV_X4 _u0_u25_U163  ( .A(1'b0), .ZN(_u0_u25_ch_am0[12] ) );
INV_X4 _u0_u25_U161  ( .A(1'b0), .ZN(_u0_u25_ch_am0[11] ) );
INV_X4 _u0_u25_U159  ( .A(1'b0), .ZN(_u0_u25_ch_am0[10] ) );
INV_X4 _u0_u25_U157  ( .A(1'b0), .ZN(_u0_u25_ch_am0[9] ) );
INV_X4 _u0_u25_U155  ( .A(1'b0), .ZN(_u0_u25_ch_am0[8] ) );
INV_X4 _u0_u25_U153  ( .A(1'b0), .ZN(_u0_u25_ch_am0[7] ) );
INV_X4 _u0_u25_U151  ( .A(1'b0), .ZN(_u0_u25_ch_am0[6] ) );
INV_X4 _u0_u25_U149  ( .A(1'b0), .ZN(_u0_u25_ch_am0[5] ) );
INV_X4 _u0_u25_U147  ( .A(1'b0), .ZN(_u0_u25_ch_am0[4] ) );
INV_X4 _u0_u25_U145  ( .A(1'b1), .ZN(_u0_u25_ch_am0[3] ) );
INV_X4 _u0_u25_U143  ( .A(1'b1), .ZN(_u0_u25_ch_am0[2] ) );
INV_X4 _u0_u25_U141  ( .A(1'b1), .ZN(_u0_u25_ch_am0[1] ) );
INV_X4 _u0_u25_U139  ( .A(1'b1), .ZN(_u0_u25_ch_am0[0] ) );
INV_X4 _u0_u25_U137  ( .A(1'b0), .ZN(_u0_u25_ch_am1[31] ) );
INV_X4 _u0_u25_U135  ( .A(1'b0), .ZN(_u0_u25_ch_am1[30] ) );
INV_X4 _u0_u25_U133  ( .A(1'b0), .ZN(_u0_u25_ch_am1[29] ) );
INV_X4 _u0_u25_U131  ( .A(1'b0), .ZN(_u0_u25_ch_am1[28] ) );
INV_X4 _u0_u25_U129  ( .A(1'b0), .ZN(_u0_u25_ch_am1[27] ) );
INV_X4 _u0_u25_U127  ( .A(1'b0), .ZN(_u0_u25_ch_am1[26] ) );
INV_X4 _u0_u25_U125  ( .A(1'b0), .ZN(_u0_u25_ch_am1[25] ) );
INV_X4 _u0_u25_U123  ( .A(1'b0), .ZN(_u0_u25_ch_am1[24] ) );
INV_X4 _u0_u25_U121  ( .A(1'b0), .ZN(_u0_u25_ch_am1[23] ) );
INV_X4 _u0_u25_U119  ( .A(1'b0), .ZN(_u0_u25_ch_am1[22] ) );
INV_X4 _u0_u25_U117  ( .A(1'b0), .ZN(_u0_u25_ch_am1[21] ) );
INV_X4 _u0_u25_U115  ( .A(1'b0), .ZN(_u0_u25_ch_am1[20] ) );
INV_X4 _u0_u25_U113  ( .A(1'b0), .ZN(_u0_u25_ch_am1[19] ) );
INV_X4 _u0_u25_U111  ( .A(1'b0), .ZN(_u0_u25_ch_am1[18] ) );
INV_X4 _u0_u25_U109  ( .A(1'b0), .ZN(_u0_u25_ch_am1[17] ) );
INV_X4 _u0_u25_U107  ( .A(1'b0), .ZN(_u0_u25_ch_am1[16] ) );
INV_X4 _u0_u25_U105  ( .A(1'b0), .ZN(_u0_u25_ch_am1[15] ) );
INV_X4 _u0_u25_U103  ( .A(1'b0), .ZN(_u0_u25_ch_am1[14] ) );
INV_X4 _u0_u25_U101  ( .A(1'b0), .ZN(_u0_u25_ch_am1[13] ) );
INV_X4 _u0_u25_U99  ( .A(1'b0), .ZN(_u0_u25_ch_am1[12] ) );
INV_X4 _u0_u25_U97  ( .A(1'b0), .ZN(_u0_u25_ch_am1[11] ) );
INV_X4 _u0_u25_U95  ( .A(1'b0), .ZN(_u0_u25_ch_am1[10] ) );
INV_X4 _u0_u25_U93  ( .A(1'b0), .ZN(_u0_u25_ch_am1[9] ) );
INV_X4 _u0_u25_U91  ( .A(1'b0), .ZN(_u0_u25_ch_am1[8] ) );
INV_X4 _u0_u25_U89  ( .A(1'b0), .ZN(_u0_u25_ch_am1[7] ) );
INV_X4 _u0_u25_U87  ( .A(1'b0), .ZN(_u0_u25_ch_am1[6] ) );
INV_X4 _u0_u25_U85  ( .A(1'b0), .ZN(_u0_u25_ch_am1[5] ) );
INV_X4 _u0_u25_U83  ( .A(1'b0), .ZN(_u0_u25_ch_am1[4] ) );
INV_X4 _u0_u25_U81  ( .A(1'b1), .ZN(_u0_u25_ch_am1[3] ) );
INV_X4 _u0_u25_U79  ( .A(1'b1), .ZN(_u0_u25_ch_am1[2] ) );
INV_X4 _u0_u25_U77  ( .A(1'b1), .ZN(_u0_u25_ch_am1[1] ) );
INV_X4 _u0_u25_U75  ( .A(1'b1), .ZN(_u0_u25_ch_am1[0] ) );
INV_X4 _u0_u25_U73  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[31] ) );
INV_X4 _u0_u25_U71  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[30] ) );
INV_X4 _u0_u25_U69  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[29] ) );
INV_X4 _u0_u25_U67  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[28] ) );
INV_X4 _u0_u25_U65  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[27] ) );
INV_X4 _u0_u25_U63  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[26] ) );
INV_X4 _u0_u25_U61  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[25] ) );
INV_X4 _u0_u25_U59  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[24] ) );
INV_X4 _u0_u25_U57  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[23] ) );
INV_X4 _u0_u25_U55  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[22] ) );
INV_X4 _u0_u25_U53  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[21] ) );
INV_X4 _u0_u25_U51  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[20] ) );
INV_X4 _u0_u25_U49  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[19] ) );
INV_X4 _u0_u25_U47  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[18] ) );
INV_X4 _u0_u25_U45  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[17] ) );
INV_X4 _u0_u25_U43  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[16] ) );
INV_X4 _u0_u25_U41  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[15] ) );
INV_X4 _u0_u25_U39  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[14] ) );
INV_X4 _u0_u25_U37  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[13] ) );
INV_X4 _u0_u25_U35  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[12] ) );
INV_X4 _u0_u25_U33  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[11] ) );
INV_X4 _u0_u25_U31  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[10] ) );
INV_X4 _u0_u25_U29  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[9] ) );
INV_X4 _u0_u25_U27  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[8] ) );
INV_X4 _u0_u25_U25  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[7] ) );
INV_X4 _u0_u25_U23  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[6] ) );
INV_X4 _u0_u25_U21  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[5] ) );
INV_X4 _u0_u25_U19  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[4] ) );
INV_X4 _u0_u25_U17  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[3] ) );
INV_X4 _u0_u25_U15  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[2] ) );
INV_X4 _u0_u25_U13  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[1] ) );
INV_X4 _u0_u25_U11  ( .A(1'b1), .ZN(_u0_u25_sw_pointer[0] ) );
INV_X4 _u0_u25_U9  ( .A(1'b1), .ZN(_u0_u25_ch_stop ) );
INV_X4 _u0_u25_U7  ( .A(1'b1), .ZN(_u0_u25_ch_dis ) );
INV_X4 _u0_u25_U5  ( .A(1'b1), .ZN(_u0_u25_int ) );
INV_X4 _u0_u26_U585  ( .A(1'b1), .ZN(_u0_u26_pointer[31] ) );
INV_X4 _u0_u26_U583  ( .A(1'b1), .ZN(_u0_u26_pointer[30] ) );
INV_X4 _u0_u26_U581  ( .A(1'b1), .ZN(_u0_u26_pointer[29] ) );
INV_X4 _u0_u26_U579  ( .A(1'b1), .ZN(_u0_u26_pointer[28] ) );
INV_X4 _u0_u26_U577  ( .A(1'b1), .ZN(_u0_u26_pointer[27] ) );
INV_X4 _u0_u26_U575  ( .A(1'b1), .ZN(_u0_u26_pointer[26] ) );
INV_X4 _u0_u26_U573  ( .A(1'b1), .ZN(_u0_u26_pointer[25] ) );
INV_X4 _u0_u26_U571  ( .A(1'b1), .ZN(_u0_u26_pointer[24] ) );
INV_X4 _u0_u26_U569  ( .A(1'b1), .ZN(_u0_u26_pointer[23] ) );
INV_X4 _u0_u26_U567  ( .A(1'b1), .ZN(_u0_u26_pointer[22] ) );
INV_X4 _u0_u26_U565  ( .A(1'b1), .ZN(_u0_u26_pointer[21] ) );
INV_X4 _u0_u26_U563  ( .A(1'b1), .ZN(_u0_u26_pointer[20] ) );
INV_X4 _u0_u26_U561  ( .A(1'b1), .ZN(_u0_u26_pointer[19] ) );
INV_X4 _u0_u26_U559  ( .A(1'b1), .ZN(_u0_u26_pointer[18] ) );
INV_X4 _u0_u26_U557  ( .A(1'b1), .ZN(_u0_u26_pointer[17] ) );
INV_X4 _u0_u26_U555  ( .A(1'b1), .ZN(_u0_u26_pointer[16] ) );
INV_X4 _u0_u26_U553  ( .A(1'b1), .ZN(_u0_u26_pointer[15] ) );
INV_X4 _u0_u26_U551  ( .A(1'b1), .ZN(_u0_u26_pointer[14] ) );
INV_X4 _u0_u26_U549  ( .A(1'b1), .ZN(_u0_u26_pointer[13] ) );
INV_X4 _u0_u26_U547  ( .A(1'b1), .ZN(_u0_u26_pointer[12] ) );
INV_X4 _u0_u26_U545  ( .A(1'b1), .ZN(_u0_u26_pointer[11] ) );
INV_X4 _u0_u26_U543  ( .A(1'b1), .ZN(_u0_u26_pointer[10] ) );
INV_X4 _u0_u26_U541  ( .A(1'b1), .ZN(_u0_u26_pointer[9] ) );
INV_X4 _u0_u26_U539  ( .A(1'b1), .ZN(_u0_u26_pointer[8] ) );
INV_X4 _u0_u26_U537  ( .A(1'b1), .ZN(_u0_u26_pointer[7] ) );
INV_X4 _u0_u26_U535  ( .A(1'b1), .ZN(_u0_u26_pointer[6] ) );
INV_X4 _u0_u26_U533  ( .A(1'b1), .ZN(_u0_u26_pointer[5] ) );
INV_X4 _u0_u26_U531  ( .A(1'b1), .ZN(_u0_u26_pointer[4] ) );
INV_X4 _u0_u26_U529  ( .A(1'b1), .ZN(_u0_u26_pointer[3] ) );
INV_X4 _u0_u26_U527  ( .A(1'b1), .ZN(_u0_u26_pointer[2] ) );
INV_X4 _u0_u26_U525  ( .A(1'b1), .ZN(_u0_u26_pointer[1] ) );
INV_X4 _u0_u26_U523  ( .A(1'b1), .ZN(_u0_u26_pointer[0] ) );
INV_X4 _u0_u26_U521  ( .A(1'b1), .ZN(_u0_u26_pointer_s[31] ) );
INV_X4 _u0_u26_U519  ( .A(1'b1), .ZN(_u0_u26_pointer_s[30] ) );
INV_X4 _u0_u26_U517  ( .A(1'b1), .ZN(_u0_u26_pointer_s[29] ) );
INV_X4 _u0_u26_U515  ( .A(1'b1), .ZN(_u0_u26_pointer_s[28] ) );
INV_X4 _u0_u26_U513  ( .A(1'b1), .ZN(_u0_u26_pointer_s[27] ) );
INV_X4 _u0_u26_U511  ( .A(1'b1), .ZN(_u0_u26_pointer_s[26] ) );
INV_X4 _u0_u26_U509  ( .A(1'b1), .ZN(_u0_u26_pointer_s[25] ) );
INV_X4 _u0_u26_U507  ( .A(1'b1), .ZN(_u0_u26_pointer_s[24] ) );
INV_X4 _u0_u26_U505  ( .A(1'b1), .ZN(_u0_u26_pointer_s[23] ) );
INV_X4 _u0_u26_U503  ( .A(1'b1), .ZN(_u0_u26_pointer_s[22] ) );
INV_X4 _u0_u26_U501  ( .A(1'b1), .ZN(_u0_u26_pointer_s[21] ) );
INV_X4 _u0_u26_U499  ( .A(1'b1), .ZN(_u0_u26_pointer_s[20] ) );
INV_X4 _u0_u26_U497  ( .A(1'b1), .ZN(_u0_u26_pointer_s[19] ) );
INV_X4 _u0_u26_U495  ( .A(1'b1), .ZN(_u0_u26_pointer_s[18] ) );
INV_X4 _u0_u26_U493  ( .A(1'b1), .ZN(_u0_u26_pointer_s[17] ) );
INV_X4 _u0_u26_U491  ( .A(1'b1), .ZN(_u0_u26_pointer_s[16] ) );
INV_X4 _u0_u26_U489  ( .A(1'b1), .ZN(_u0_u26_pointer_s[15] ) );
INV_X4 _u0_u26_U487  ( .A(1'b1), .ZN(_u0_u26_pointer_s[14] ) );
INV_X4 _u0_u26_U485  ( .A(1'b1), .ZN(_u0_u26_pointer_s[13] ) );
INV_X4 _u0_u26_U483  ( .A(1'b1), .ZN(_u0_u26_pointer_s[12] ) );
INV_X4 _u0_u26_U481  ( .A(1'b1), .ZN(_u0_u26_pointer_s[11] ) );
INV_X4 _u0_u26_U479  ( .A(1'b1), .ZN(_u0_u26_pointer_s[10] ) );
INV_X4 _u0_u26_U477  ( .A(1'b1), .ZN(_u0_u26_pointer_s[9] ) );
INV_X4 _u0_u26_U475  ( .A(1'b1), .ZN(_u0_u26_pointer_s[8] ) );
INV_X4 _u0_u26_U473  ( .A(1'b1), .ZN(_u0_u26_pointer_s[7] ) );
INV_X4 _u0_u26_U471  ( .A(1'b1), .ZN(_u0_u26_pointer_s[6] ) );
INV_X4 _u0_u26_U469  ( .A(1'b1), .ZN(_u0_u26_pointer_s[5] ) );
INV_X4 _u0_u26_U467  ( .A(1'b1), .ZN(_u0_u26_pointer_s[4] ) );
INV_X4 _u0_u26_U465  ( .A(1'b1), .ZN(_u0_u26_pointer_s[3] ) );
INV_X4 _u0_u26_U463  ( .A(1'b1), .ZN(_u0_u26_pointer_s[2] ) );
INV_X4 _u0_u26_U461  ( .A(1'b1), .ZN(_u0_u26_pointer_s[1] ) );
INV_X4 _u0_u26_U459  ( .A(1'b1), .ZN(_u0_u26_pointer_s[0] ) );
INV_X4 _u0_u26_U457  ( .A(1'b1), .ZN(_u0_u26_ch_csr[31] ) );
INV_X4 _u0_u26_U455  ( .A(1'b1), .ZN(_u0_u26_ch_csr[30] ) );
INV_X4 _u0_u26_U453  ( .A(1'b1), .ZN(_u0_u26_ch_csr[29] ) );
INV_X4 _u0_u26_U451  ( .A(1'b1), .ZN(_u0_u26_ch_csr[28] ) );
INV_X4 _u0_u26_U449  ( .A(1'b1), .ZN(_u0_u26_ch_csr[27] ) );
INV_X4 _u0_u26_U447  ( .A(1'b1), .ZN(_u0_u26_ch_csr[26] ) );
INV_X4 _u0_u26_U445  ( .A(1'b1), .ZN(_u0_u26_ch_csr[25] ) );
INV_X4 _u0_u26_U443  ( .A(1'b1), .ZN(_u0_u26_ch_csr[24] ) );
INV_X4 _u0_u26_U441  ( .A(1'b1), .ZN(_u0_u26_ch_csr[23] ) );
INV_X4 _u0_u26_U439  ( .A(1'b1), .ZN(_u0_u26_ch_csr[22] ) );
INV_X4 _u0_u26_U437  ( .A(1'b1), .ZN(_u0_u26_ch_csr[21] ) );
INV_X4 _u0_u26_U435  ( .A(1'b1), .ZN(_u0_u26_ch_csr[20] ) );
INV_X4 _u0_u26_U433  ( .A(1'b1), .ZN(_u0_u26_ch_csr[19] ) );
INV_X4 _u0_u26_U431  ( .A(1'b1), .ZN(_u0_u26_ch_csr[18] ) );
INV_X4 _u0_u26_U429  ( .A(1'b1), .ZN(_u0_u26_ch_csr[17] ) );
INV_X4 _u0_u26_U427  ( .A(1'b1), .ZN(_u0_u26_ch_csr[16] ) );
INV_X4 _u0_u26_U425  ( .A(1'b1), .ZN(_u0_u26_ch_csr[15] ) );
INV_X4 _u0_u26_U423  ( .A(1'b1), .ZN(_u0_u26_ch_csr[14] ) );
INV_X4 _u0_u26_U421  ( .A(1'b1), .ZN(_u0_u26_ch_csr[13] ) );
INV_X4 _u0_u26_U419  ( .A(1'b1), .ZN(_u0_u26_ch_csr[12] ) );
INV_X4 _u0_u26_U417  ( .A(1'b1), .ZN(_u0_u26_ch_csr[11] ) );
INV_X4 _u0_u26_U415  ( .A(1'b1), .ZN(_u0_u26_ch_csr[10] ) );
INV_X4 _u0_u26_U413  ( .A(1'b1), .ZN(_u0_u26_ch_csr[9] ) );
INV_X4 _u0_u26_U411  ( .A(1'b1), .ZN(_u0_u26_ch_csr[8] ) );
INV_X4 _u0_u26_U409  ( .A(1'b1), .ZN(_u0_u26_ch_csr[7] ) );
INV_X4 _u0_u26_U407  ( .A(1'b1), .ZN(_u0_u26_ch_csr[6] ) );
INV_X4 _u0_u26_U405  ( .A(1'b1), .ZN(_u0_u26_ch_csr[5] ) );
INV_X4 _u0_u26_U403  ( .A(1'b1), .ZN(_u0_u26_ch_csr[4] ) );
INV_X4 _u0_u26_U401  ( .A(1'b1), .ZN(_u0_u26_ch_csr[3] ) );
INV_X4 _u0_u26_U399  ( .A(1'b1), .ZN(_u0_u26_ch_csr[2] ) );
INV_X4 _u0_u26_U397  ( .A(1'b1), .ZN(_u0_u26_ch_csr[1] ) );
INV_X4 _u0_u26_U395  ( .A(1'b1), .ZN(_u0_u26_ch_csr[0] ) );
INV_X4 _u0_u26_U393  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[31] ) );
INV_X4 _u0_u26_U391  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[30] ) );
INV_X4 _u0_u26_U389  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[29] ) );
INV_X4 _u0_u26_U387  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[28] ) );
INV_X4 _u0_u26_U385  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[27] ) );
INV_X4 _u0_u26_U383  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[26] ) );
INV_X4 _u0_u26_U381  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[25] ) );
INV_X4 _u0_u26_U379  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[24] ) );
INV_X4 _u0_u26_U377  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[23] ) );
INV_X4 _u0_u26_U375  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[22] ) );
INV_X4 _u0_u26_U373  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[21] ) );
INV_X4 _u0_u26_U371  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[20] ) );
INV_X4 _u0_u26_U369  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[19] ) );
INV_X4 _u0_u26_U367  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[18] ) );
INV_X4 _u0_u26_U365  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[17] ) );
INV_X4 _u0_u26_U363  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[16] ) );
INV_X4 _u0_u26_U361  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[15] ) );
INV_X4 _u0_u26_U359  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[14] ) );
INV_X4 _u0_u26_U357  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[13] ) );
INV_X4 _u0_u26_U355  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[12] ) );
INV_X4 _u0_u26_U353  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[11] ) );
INV_X4 _u0_u26_U351  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[10] ) );
INV_X4 _u0_u26_U349  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[9] ) );
INV_X4 _u0_u26_U347  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[8] ) );
INV_X4 _u0_u26_U345  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[7] ) );
INV_X4 _u0_u26_U343  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[6] ) );
INV_X4 _u0_u26_U341  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[5] ) );
INV_X4 _u0_u26_U339  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[4] ) );
INV_X4 _u0_u26_U337  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[3] ) );
INV_X4 _u0_u26_U335  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[2] ) );
INV_X4 _u0_u26_U333  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[1] ) );
INV_X4 _u0_u26_U331  ( .A(1'b1), .ZN(_u0_u26_ch_txsz[0] ) );
INV_X4 _u0_u26_U329  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[31] ) );
INV_X4 _u0_u26_U327  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[30] ) );
INV_X4 _u0_u26_U325  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[29] ) );
INV_X4 _u0_u26_U323  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[28] ) );
INV_X4 _u0_u26_U321  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[27] ) );
INV_X4 _u0_u26_U319  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[26] ) );
INV_X4 _u0_u26_U317  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[25] ) );
INV_X4 _u0_u26_U315  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[24] ) );
INV_X4 _u0_u26_U313  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[23] ) );
INV_X4 _u0_u26_U311  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[22] ) );
INV_X4 _u0_u26_U309  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[21] ) );
INV_X4 _u0_u26_U307  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[20] ) );
INV_X4 _u0_u26_U305  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[19] ) );
INV_X4 _u0_u26_U303  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[18] ) );
INV_X4 _u0_u26_U301  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[17] ) );
INV_X4 _u0_u26_U299  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[16] ) );
INV_X4 _u0_u26_U297  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[15] ) );
INV_X4 _u0_u26_U295  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[14] ) );
INV_X4 _u0_u26_U293  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[13] ) );
INV_X4 _u0_u26_U291  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[12] ) );
INV_X4 _u0_u26_U289  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[11] ) );
INV_X4 _u0_u26_U287  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[10] ) );
INV_X4 _u0_u26_U285  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[9] ) );
INV_X4 _u0_u26_U283  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[8] ) );
INV_X4 _u0_u26_U281  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[7] ) );
INV_X4 _u0_u26_U279  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[6] ) );
INV_X4 _u0_u26_U277  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[5] ) );
INV_X4 _u0_u26_U275  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[4] ) );
INV_X4 _u0_u26_U273  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[3] ) );
INV_X4 _u0_u26_U271  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[2] ) );
INV_X4 _u0_u26_U269  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[1] ) );
INV_X4 _u0_u26_U267  ( .A(1'b1), .ZN(_u0_u26_ch_adr0[0] ) );
INV_X4 _u0_u26_U265  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[31] ) );
INV_X4 _u0_u26_U263  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[30] ) );
INV_X4 _u0_u26_U261  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[29] ) );
INV_X4 _u0_u26_U259  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[28] ) );
INV_X4 _u0_u26_U257  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[27] ) );
INV_X4 _u0_u26_U255  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[26] ) );
INV_X4 _u0_u26_U253  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[25] ) );
INV_X4 _u0_u26_U251  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[24] ) );
INV_X4 _u0_u26_U249  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[23] ) );
INV_X4 _u0_u26_U247  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[22] ) );
INV_X4 _u0_u26_U245  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[21] ) );
INV_X4 _u0_u26_U243  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[20] ) );
INV_X4 _u0_u26_U241  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[19] ) );
INV_X4 _u0_u26_U239  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[18] ) );
INV_X4 _u0_u26_U237  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[17] ) );
INV_X4 _u0_u26_U235  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[16] ) );
INV_X4 _u0_u26_U233  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[15] ) );
INV_X4 _u0_u26_U231  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[14] ) );
INV_X4 _u0_u26_U229  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[13] ) );
INV_X4 _u0_u26_U227  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[12] ) );
INV_X4 _u0_u26_U225  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[11] ) );
INV_X4 _u0_u26_U223  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[10] ) );
INV_X4 _u0_u26_U221  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[9] ) );
INV_X4 _u0_u26_U219  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[8] ) );
INV_X4 _u0_u26_U217  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[7] ) );
INV_X4 _u0_u26_U215  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[6] ) );
INV_X4 _u0_u26_U213  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[5] ) );
INV_X4 _u0_u26_U211  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[4] ) );
INV_X4 _u0_u26_U209  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[3] ) );
INV_X4 _u0_u26_U207  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[2] ) );
INV_X4 _u0_u26_U205  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[1] ) );
INV_X4 _u0_u26_U203  ( .A(1'b1), .ZN(_u0_u26_ch_adr1[0] ) );
INV_X4 _u0_u26_U201  ( .A(1'b0), .ZN(_u0_u26_ch_am0[31] ) );
INV_X4 _u0_u26_U199  ( .A(1'b0), .ZN(_u0_u26_ch_am0[30] ) );
INV_X4 _u0_u26_U197  ( .A(1'b0), .ZN(_u0_u26_ch_am0[29] ) );
INV_X4 _u0_u26_U195  ( .A(1'b0), .ZN(_u0_u26_ch_am0[28] ) );
INV_X4 _u0_u26_U193  ( .A(1'b0), .ZN(_u0_u26_ch_am0[27] ) );
INV_X4 _u0_u26_U191  ( .A(1'b0), .ZN(_u0_u26_ch_am0[26] ) );
INV_X4 _u0_u26_U189  ( .A(1'b0), .ZN(_u0_u26_ch_am0[25] ) );
INV_X4 _u0_u26_U187  ( .A(1'b0), .ZN(_u0_u26_ch_am0[24] ) );
INV_X4 _u0_u26_U185  ( .A(1'b0), .ZN(_u0_u26_ch_am0[23] ) );
INV_X4 _u0_u26_U183  ( .A(1'b0), .ZN(_u0_u26_ch_am0[22] ) );
INV_X4 _u0_u26_U181  ( .A(1'b0), .ZN(_u0_u26_ch_am0[21] ) );
INV_X4 _u0_u26_U179  ( .A(1'b0), .ZN(_u0_u26_ch_am0[20] ) );
INV_X4 _u0_u26_U177  ( .A(1'b0), .ZN(_u0_u26_ch_am0[19] ) );
INV_X4 _u0_u26_U175  ( .A(1'b0), .ZN(_u0_u26_ch_am0[18] ) );
INV_X4 _u0_u26_U173  ( .A(1'b0), .ZN(_u0_u26_ch_am0[17] ) );
INV_X4 _u0_u26_U171  ( .A(1'b0), .ZN(_u0_u26_ch_am0[16] ) );
INV_X4 _u0_u26_U169  ( .A(1'b0), .ZN(_u0_u26_ch_am0[15] ) );
INV_X4 _u0_u26_U167  ( .A(1'b0), .ZN(_u0_u26_ch_am0[14] ) );
INV_X4 _u0_u26_U165  ( .A(1'b0), .ZN(_u0_u26_ch_am0[13] ) );
INV_X4 _u0_u26_U163  ( .A(1'b0), .ZN(_u0_u26_ch_am0[12] ) );
INV_X4 _u0_u26_U161  ( .A(1'b0), .ZN(_u0_u26_ch_am0[11] ) );
INV_X4 _u0_u26_U159  ( .A(1'b0), .ZN(_u0_u26_ch_am0[10] ) );
INV_X4 _u0_u26_U157  ( .A(1'b0), .ZN(_u0_u26_ch_am0[9] ) );
INV_X4 _u0_u26_U155  ( .A(1'b0), .ZN(_u0_u26_ch_am0[8] ) );
INV_X4 _u0_u26_U153  ( .A(1'b0), .ZN(_u0_u26_ch_am0[7] ) );
INV_X4 _u0_u26_U151  ( .A(1'b0), .ZN(_u0_u26_ch_am0[6] ) );
INV_X4 _u0_u26_U149  ( .A(1'b0), .ZN(_u0_u26_ch_am0[5] ) );
INV_X4 _u0_u26_U147  ( .A(1'b0), .ZN(_u0_u26_ch_am0[4] ) );
INV_X4 _u0_u26_U145  ( .A(1'b1), .ZN(_u0_u26_ch_am0[3] ) );
INV_X4 _u0_u26_U143  ( .A(1'b1), .ZN(_u0_u26_ch_am0[2] ) );
INV_X4 _u0_u26_U141  ( .A(1'b1), .ZN(_u0_u26_ch_am0[1] ) );
INV_X4 _u0_u26_U139  ( .A(1'b1), .ZN(_u0_u26_ch_am0[0] ) );
INV_X4 _u0_u26_U137  ( .A(1'b0), .ZN(_u0_u26_ch_am1[31] ) );
INV_X4 _u0_u26_U135  ( .A(1'b0), .ZN(_u0_u26_ch_am1[30] ) );
INV_X4 _u0_u26_U133  ( .A(1'b0), .ZN(_u0_u26_ch_am1[29] ) );
INV_X4 _u0_u26_U131  ( .A(1'b0), .ZN(_u0_u26_ch_am1[28] ) );
INV_X4 _u0_u26_U129  ( .A(1'b0), .ZN(_u0_u26_ch_am1[27] ) );
INV_X4 _u0_u26_U127  ( .A(1'b0), .ZN(_u0_u26_ch_am1[26] ) );
INV_X4 _u0_u26_U125  ( .A(1'b0), .ZN(_u0_u26_ch_am1[25] ) );
INV_X4 _u0_u26_U123  ( .A(1'b0), .ZN(_u0_u26_ch_am1[24] ) );
INV_X4 _u0_u26_U121  ( .A(1'b0), .ZN(_u0_u26_ch_am1[23] ) );
INV_X4 _u0_u26_U119  ( .A(1'b0), .ZN(_u0_u26_ch_am1[22] ) );
INV_X4 _u0_u26_U117  ( .A(1'b0), .ZN(_u0_u26_ch_am1[21] ) );
INV_X4 _u0_u26_U115  ( .A(1'b0), .ZN(_u0_u26_ch_am1[20] ) );
INV_X4 _u0_u26_U113  ( .A(1'b0), .ZN(_u0_u26_ch_am1[19] ) );
INV_X4 _u0_u26_U111  ( .A(1'b0), .ZN(_u0_u26_ch_am1[18] ) );
INV_X4 _u0_u26_U109  ( .A(1'b0), .ZN(_u0_u26_ch_am1[17] ) );
INV_X4 _u0_u26_U107  ( .A(1'b0), .ZN(_u0_u26_ch_am1[16] ) );
INV_X4 _u0_u26_U105  ( .A(1'b0), .ZN(_u0_u26_ch_am1[15] ) );
INV_X4 _u0_u26_U103  ( .A(1'b0), .ZN(_u0_u26_ch_am1[14] ) );
INV_X4 _u0_u26_U101  ( .A(1'b0), .ZN(_u0_u26_ch_am1[13] ) );
INV_X4 _u0_u26_U99  ( .A(1'b0), .ZN(_u0_u26_ch_am1[12] ) );
INV_X4 _u0_u26_U97  ( .A(1'b0), .ZN(_u0_u26_ch_am1[11] ) );
INV_X4 _u0_u26_U95  ( .A(1'b0), .ZN(_u0_u26_ch_am1[10] ) );
INV_X4 _u0_u26_U93  ( .A(1'b0), .ZN(_u0_u26_ch_am1[9] ) );
INV_X4 _u0_u26_U91  ( .A(1'b0), .ZN(_u0_u26_ch_am1[8] ) );
INV_X4 _u0_u26_U89  ( .A(1'b0), .ZN(_u0_u26_ch_am1[7] ) );
INV_X4 _u0_u26_U87  ( .A(1'b0), .ZN(_u0_u26_ch_am1[6] ) );
INV_X4 _u0_u26_U85  ( .A(1'b0), .ZN(_u0_u26_ch_am1[5] ) );
INV_X4 _u0_u26_U83  ( .A(1'b0), .ZN(_u0_u26_ch_am1[4] ) );
INV_X4 _u0_u26_U81  ( .A(1'b1), .ZN(_u0_u26_ch_am1[3] ) );
INV_X4 _u0_u26_U79  ( .A(1'b1), .ZN(_u0_u26_ch_am1[2] ) );
INV_X4 _u0_u26_U77  ( .A(1'b1), .ZN(_u0_u26_ch_am1[1] ) );
INV_X4 _u0_u26_U75  ( .A(1'b1), .ZN(_u0_u26_ch_am1[0] ) );
INV_X4 _u0_u26_U73  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[31] ) );
INV_X4 _u0_u26_U71  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[30] ) );
INV_X4 _u0_u26_U69  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[29] ) );
INV_X4 _u0_u26_U67  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[28] ) );
INV_X4 _u0_u26_U65  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[27] ) );
INV_X4 _u0_u26_U63  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[26] ) );
INV_X4 _u0_u26_U61  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[25] ) );
INV_X4 _u0_u26_U59  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[24] ) );
INV_X4 _u0_u26_U57  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[23] ) );
INV_X4 _u0_u26_U55  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[22] ) );
INV_X4 _u0_u26_U53  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[21] ) );
INV_X4 _u0_u26_U51  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[20] ) );
INV_X4 _u0_u26_U49  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[19] ) );
INV_X4 _u0_u26_U47  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[18] ) );
INV_X4 _u0_u26_U45  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[17] ) );
INV_X4 _u0_u26_U43  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[16] ) );
INV_X4 _u0_u26_U41  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[15] ) );
INV_X4 _u0_u26_U39  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[14] ) );
INV_X4 _u0_u26_U37  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[13] ) );
INV_X4 _u0_u26_U35  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[12] ) );
INV_X4 _u0_u26_U33  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[11] ) );
INV_X4 _u0_u26_U31  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[10] ) );
INV_X4 _u0_u26_U29  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[9] ) );
INV_X4 _u0_u26_U27  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[8] ) );
INV_X4 _u0_u26_U25  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[7] ) );
INV_X4 _u0_u26_U23  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[6] ) );
INV_X4 _u0_u26_U21  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[5] ) );
INV_X4 _u0_u26_U19  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[4] ) );
INV_X4 _u0_u26_U17  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[3] ) );
INV_X4 _u0_u26_U15  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[2] ) );
INV_X4 _u0_u26_U13  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[1] ) );
INV_X4 _u0_u26_U11  ( .A(1'b1), .ZN(_u0_u26_sw_pointer[0] ) );
INV_X4 _u0_u26_U9  ( .A(1'b1), .ZN(_u0_u26_ch_stop ) );
INV_X4 _u0_u26_U7  ( .A(1'b1), .ZN(_u0_u26_ch_dis ) );
INV_X4 _u0_u26_U5  ( .A(1'b1), .ZN(_u0_u26_int ) );
INV_X4 _u0_u27_U585  ( .A(1'b1), .ZN(_u0_u27_pointer[31] ) );
INV_X4 _u0_u27_U583  ( .A(1'b1), .ZN(_u0_u27_pointer[30] ) );
INV_X4 _u0_u27_U581  ( .A(1'b1), .ZN(_u0_u27_pointer[29] ) );
INV_X4 _u0_u27_U579  ( .A(1'b1), .ZN(_u0_u27_pointer[28] ) );
INV_X4 _u0_u27_U577  ( .A(1'b1), .ZN(_u0_u27_pointer[27] ) );
INV_X4 _u0_u27_U575  ( .A(1'b1), .ZN(_u0_u27_pointer[26] ) );
INV_X4 _u0_u27_U573  ( .A(1'b1), .ZN(_u0_u27_pointer[25] ) );
INV_X4 _u0_u27_U571  ( .A(1'b1), .ZN(_u0_u27_pointer[24] ) );
INV_X4 _u0_u27_U569  ( .A(1'b1), .ZN(_u0_u27_pointer[23] ) );
INV_X4 _u0_u27_U567  ( .A(1'b1), .ZN(_u0_u27_pointer[22] ) );
INV_X4 _u0_u27_U565  ( .A(1'b1), .ZN(_u0_u27_pointer[21] ) );
INV_X4 _u0_u27_U563  ( .A(1'b1), .ZN(_u0_u27_pointer[20] ) );
INV_X4 _u0_u27_U561  ( .A(1'b1), .ZN(_u0_u27_pointer[19] ) );
INV_X4 _u0_u27_U559  ( .A(1'b1), .ZN(_u0_u27_pointer[18] ) );
INV_X4 _u0_u27_U557  ( .A(1'b1), .ZN(_u0_u27_pointer[17] ) );
INV_X4 _u0_u27_U555  ( .A(1'b1), .ZN(_u0_u27_pointer[16] ) );
INV_X4 _u0_u27_U553  ( .A(1'b1), .ZN(_u0_u27_pointer[15] ) );
INV_X4 _u0_u27_U551  ( .A(1'b1), .ZN(_u0_u27_pointer[14] ) );
INV_X4 _u0_u27_U549  ( .A(1'b1), .ZN(_u0_u27_pointer[13] ) );
INV_X4 _u0_u27_U547  ( .A(1'b1), .ZN(_u0_u27_pointer[12] ) );
INV_X4 _u0_u27_U545  ( .A(1'b1), .ZN(_u0_u27_pointer[11] ) );
INV_X4 _u0_u27_U543  ( .A(1'b1), .ZN(_u0_u27_pointer[10] ) );
INV_X4 _u0_u27_U541  ( .A(1'b1), .ZN(_u0_u27_pointer[9] ) );
INV_X4 _u0_u27_U539  ( .A(1'b1), .ZN(_u0_u27_pointer[8] ) );
INV_X4 _u0_u27_U537  ( .A(1'b1), .ZN(_u0_u27_pointer[7] ) );
INV_X4 _u0_u27_U535  ( .A(1'b1), .ZN(_u0_u27_pointer[6] ) );
INV_X4 _u0_u27_U533  ( .A(1'b1), .ZN(_u0_u27_pointer[5] ) );
INV_X4 _u0_u27_U531  ( .A(1'b1), .ZN(_u0_u27_pointer[4] ) );
INV_X4 _u0_u27_U529  ( .A(1'b1), .ZN(_u0_u27_pointer[3] ) );
INV_X4 _u0_u27_U527  ( .A(1'b1), .ZN(_u0_u27_pointer[2] ) );
INV_X4 _u0_u27_U525  ( .A(1'b1), .ZN(_u0_u27_pointer[1] ) );
INV_X4 _u0_u27_U523  ( .A(1'b1), .ZN(_u0_u27_pointer[0] ) );
INV_X4 _u0_u27_U521  ( .A(1'b1), .ZN(_u0_u27_pointer_s[31] ) );
INV_X4 _u0_u27_U519  ( .A(1'b1), .ZN(_u0_u27_pointer_s[30] ) );
INV_X4 _u0_u27_U517  ( .A(1'b1), .ZN(_u0_u27_pointer_s[29] ) );
INV_X4 _u0_u27_U515  ( .A(1'b1), .ZN(_u0_u27_pointer_s[28] ) );
INV_X4 _u0_u27_U513  ( .A(1'b1), .ZN(_u0_u27_pointer_s[27] ) );
INV_X4 _u0_u27_U511  ( .A(1'b1), .ZN(_u0_u27_pointer_s[26] ) );
INV_X4 _u0_u27_U509  ( .A(1'b1), .ZN(_u0_u27_pointer_s[25] ) );
INV_X4 _u0_u27_U507  ( .A(1'b1), .ZN(_u0_u27_pointer_s[24] ) );
INV_X4 _u0_u27_U505  ( .A(1'b1), .ZN(_u0_u27_pointer_s[23] ) );
INV_X4 _u0_u27_U503  ( .A(1'b1), .ZN(_u0_u27_pointer_s[22] ) );
INV_X4 _u0_u27_U501  ( .A(1'b1), .ZN(_u0_u27_pointer_s[21] ) );
INV_X4 _u0_u27_U499  ( .A(1'b1), .ZN(_u0_u27_pointer_s[20] ) );
INV_X4 _u0_u27_U497  ( .A(1'b1), .ZN(_u0_u27_pointer_s[19] ) );
INV_X4 _u0_u27_U495  ( .A(1'b1), .ZN(_u0_u27_pointer_s[18] ) );
INV_X4 _u0_u27_U493  ( .A(1'b1), .ZN(_u0_u27_pointer_s[17] ) );
INV_X4 _u0_u27_U491  ( .A(1'b1), .ZN(_u0_u27_pointer_s[16] ) );
INV_X4 _u0_u27_U489  ( .A(1'b1), .ZN(_u0_u27_pointer_s[15] ) );
INV_X4 _u0_u27_U487  ( .A(1'b1), .ZN(_u0_u27_pointer_s[14] ) );
INV_X4 _u0_u27_U485  ( .A(1'b1), .ZN(_u0_u27_pointer_s[13] ) );
INV_X4 _u0_u27_U483  ( .A(1'b1), .ZN(_u0_u27_pointer_s[12] ) );
INV_X4 _u0_u27_U481  ( .A(1'b1), .ZN(_u0_u27_pointer_s[11] ) );
INV_X4 _u0_u27_U479  ( .A(1'b1), .ZN(_u0_u27_pointer_s[10] ) );
INV_X4 _u0_u27_U477  ( .A(1'b1), .ZN(_u0_u27_pointer_s[9] ) );
INV_X4 _u0_u27_U475  ( .A(1'b1), .ZN(_u0_u27_pointer_s[8] ) );
INV_X4 _u0_u27_U473  ( .A(1'b1), .ZN(_u0_u27_pointer_s[7] ) );
INV_X4 _u0_u27_U471  ( .A(1'b1), .ZN(_u0_u27_pointer_s[6] ) );
INV_X4 _u0_u27_U469  ( .A(1'b1), .ZN(_u0_u27_pointer_s[5] ) );
INV_X4 _u0_u27_U467  ( .A(1'b1), .ZN(_u0_u27_pointer_s[4] ) );
INV_X4 _u0_u27_U465  ( .A(1'b1), .ZN(_u0_u27_pointer_s[3] ) );
INV_X4 _u0_u27_U463  ( .A(1'b1), .ZN(_u0_u27_pointer_s[2] ) );
INV_X4 _u0_u27_U461  ( .A(1'b1), .ZN(_u0_u27_pointer_s[1] ) );
INV_X4 _u0_u27_U459  ( .A(1'b1), .ZN(_u0_u27_pointer_s[0] ) );
INV_X4 _u0_u27_U457  ( .A(1'b1), .ZN(_u0_u27_ch_csr[31] ) );
INV_X4 _u0_u27_U455  ( .A(1'b1), .ZN(_u0_u27_ch_csr[30] ) );
INV_X4 _u0_u27_U453  ( .A(1'b1), .ZN(_u0_u27_ch_csr[29] ) );
INV_X4 _u0_u27_U451  ( .A(1'b1), .ZN(_u0_u27_ch_csr[28] ) );
INV_X4 _u0_u27_U449  ( .A(1'b1), .ZN(_u0_u27_ch_csr[27] ) );
INV_X4 _u0_u27_U447  ( .A(1'b1), .ZN(_u0_u27_ch_csr[26] ) );
INV_X4 _u0_u27_U445  ( .A(1'b1), .ZN(_u0_u27_ch_csr[25] ) );
INV_X4 _u0_u27_U443  ( .A(1'b1), .ZN(_u0_u27_ch_csr[24] ) );
INV_X4 _u0_u27_U441  ( .A(1'b1), .ZN(_u0_u27_ch_csr[23] ) );
INV_X4 _u0_u27_U439  ( .A(1'b1), .ZN(_u0_u27_ch_csr[22] ) );
INV_X4 _u0_u27_U437  ( .A(1'b1), .ZN(_u0_u27_ch_csr[21] ) );
INV_X4 _u0_u27_U435  ( .A(1'b1), .ZN(_u0_u27_ch_csr[20] ) );
INV_X4 _u0_u27_U433  ( .A(1'b1), .ZN(_u0_u27_ch_csr[19] ) );
INV_X4 _u0_u27_U431  ( .A(1'b1), .ZN(_u0_u27_ch_csr[18] ) );
INV_X4 _u0_u27_U429  ( .A(1'b1), .ZN(_u0_u27_ch_csr[17] ) );
INV_X4 _u0_u27_U427  ( .A(1'b1), .ZN(_u0_u27_ch_csr[16] ) );
INV_X4 _u0_u27_U425  ( .A(1'b1), .ZN(_u0_u27_ch_csr[15] ) );
INV_X4 _u0_u27_U423  ( .A(1'b1), .ZN(_u0_u27_ch_csr[14] ) );
INV_X4 _u0_u27_U421  ( .A(1'b1), .ZN(_u0_u27_ch_csr[13] ) );
INV_X4 _u0_u27_U419  ( .A(1'b1), .ZN(_u0_u27_ch_csr[12] ) );
INV_X4 _u0_u27_U417  ( .A(1'b1), .ZN(_u0_u27_ch_csr[11] ) );
INV_X4 _u0_u27_U415  ( .A(1'b1), .ZN(_u0_u27_ch_csr[10] ) );
INV_X4 _u0_u27_U413  ( .A(1'b1), .ZN(_u0_u27_ch_csr[9] ) );
INV_X4 _u0_u27_U411  ( .A(1'b1), .ZN(_u0_u27_ch_csr[8] ) );
INV_X4 _u0_u27_U409  ( .A(1'b1), .ZN(_u0_u27_ch_csr[7] ) );
INV_X4 _u0_u27_U407  ( .A(1'b1), .ZN(_u0_u27_ch_csr[6] ) );
INV_X4 _u0_u27_U405  ( .A(1'b1), .ZN(_u0_u27_ch_csr[5] ) );
INV_X4 _u0_u27_U403  ( .A(1'b1), .ZN(_u0_u27_ch_csr[4] ) );
INV_X4 _u0_u27_U401  ( .A(1'b1), .ZN(_u0_u27_ch_csr[3] ) );
INV_X4 _u0_u27_U399  ( .A(1'b1), .ZN(_u0_u27_ch_csr[2] ) );
INV_X4 _u0_u27_U397  ( .A(1'b1), .ZN(_u0_u27_ch_csr[1] ) );
INV_X4 _u0_u27_U395  ( .A(1'b1), .ZN(_u0_u27_ch_csr[0] ) );
INV_X4 _u0_u27_U393  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[31] ) );
INV_X4 _u0_u27_U391  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[30] ) );
INV_X4 _u0_u27_U389  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[29] ) );
INV_X4 _u0_u27_U387  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[28] ) );
INV_X4 _u0_u27_U385  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[27] ) );
INV_X4 _u0_u27_U383  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[26] ) );
INV_X4 _u0_u27_U381  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[25] ) );
INV_X4 _u0_u27_U379  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[24] ) );
INV_X4 _u0_u27_U377  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[23] ) );
INV_X4 _u0_u27_U375  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[22] ) );
INV_X4 _u0_u27_U373  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[21] ) );
INV_X4 _u0_u27_U371  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[20] ) );
INV_X4 _u0_u27_U369  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[19] ) );
INV_X4 _u0_u27_U367  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[18] ) );
INV_X4 _u0_u27_U365  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[17] ) );
INV_X4 _u0_u27_U363  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[16] ) );
INV_X4 _u0_u27_U361  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[15] ) );
INV_X4 _u0_u27_U359  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[14] ) );
INV_X4 _u0_u27_U357  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[13] ) );
INV_X4 _u0_u27_U355  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[12] ) );
INV_X4 _u0_u27_U353  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[11] ) );
INV_X4 _u0_u27_U351  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[10] ) );
INV_X4 _u0_u27_U349  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[9] ) );
INV_X4 _u0_u27_U347  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[8] ) );
INV_X4 _u0_u27_U345  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[7] ) );
INV_X4 _u0_u27_U343  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[6] ) );
INV_X4 _u0_u27_U341  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[5] ) );
INV_X4 _u0_u27_U339  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[4] ) );
INV_X4 _u0_u27_U337  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[3] ) );
INV_X4 _u0_u27_U335  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[2] ) );
INV_X4 _u0_u27_U333  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[1] ) );
INV_X4 _u0_u27_U331  ( .A(1'b1), .ZN(_u0_u27_ch_txsz[0] ) );
INV_X4 _u0_u27_U329  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[31] ) );
INV_X4 _u0_u27_U327  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[30] ) );
INV_X4 _u0_u27_U325  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[29] ) );
INV_X4 _u0_u27_U323  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[28] ) );
INV_X4 _u0_u27_U321  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[27] ) );
INV_X4 _u0_u27_U319  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[26] ) );
INV_X4 _u0_u27_U317  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[25] ) );
INV_X4 _u0_u27_U315  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[24] ) );
INV_X4 _u0_u27_U313  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[23] ) );
INV_X4 _u0_u27_U311  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[22] ) );
INV_X4 _u0_u27_U309  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[21] ) );
INV_X4 _u0_u27_U307  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[20] ) );
INV_X4 _u0_u27_U305  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[19] ) );
INV_X4 _u0_u27_U303  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[18] ) );
INV_X4 _u0_u27_U301  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[17] ) );
INV_X4 _u0_u27_U299  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[16] ) );
INV_X4 _u0_u27_U297  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[15] ) );
INV_X4 _u0_u27_U295  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[14] ) );
INV_X4 _u0_u27_U293  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[13] ) );
INV_X4 _u0_u27_U291  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[12] ) );
INV_X4 _u0_u27_U289  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[11] ) );
INV_X4 _u0_u27_U287  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[10] ) );
INV_X4 _u0_u27_U285  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[9] ) );
INV_X4 _u0_u27_U283  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[8] ) );
INV_X4 _u0_u27_U281  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[7] ) );
INV_X4 _u0_u27_U279  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[6] ) );
INV_X4 _u0_u27_U277  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[5] ) );
INV_X4 _u0_u27_U275  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[4] ) );
INV_X4 _u0_u27_U273  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[3] ) );
INV_X4 _u0_u27_U271  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[2] ) );
INV_X4 _u0_u27_U269  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[1] ) );
INV_X4 _u0_u27_U267  ( .A(1'b1), .ZN(_u0_u27_ch_adr0[0] ) );
INV_X4 _u0_u27_U265  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[31] ) );
INV_X4 _u0_u27_U263  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[30] ) );
INV_X4 _u0_u27_U261  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[29] ) );
INV_X4 _u0_u27_U259  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[28] ) );
INV_X4 _u0_u27_U257  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[27] ) );
INV_X4 _u0_u27_U255  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[26] ) );
INV_X4 _u0_u27_U253  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[25] ) );
INV_X4 _u0_u27_U251  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[24] ) );
INV_X4 _u0_u27_U249  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[23] ) );
INV_X4 _u0_u27_U247  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[22] ) );
INV_X4 _u0_u27_U245  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[21] ) );
INV_X4 _u0_u27_U243  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[20] ) );
INV_X4 _u0_u27_U241  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[19] ) );
INV_X4 _u0_u27_U239  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[18] ) );
INV_X4 _u0_u27_U237  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[17] ) );
INV_X4 _u0_u27_U235  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[16] ) );
INV_X4 _u0_u27_U233  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[15] ) );
INV_X4 _u0_u27_U231  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[14] ) );
INV_X4 _u0_u27_U229  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[13] ) );
INV_X4 _u0_u27_U227  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[12] ) );
INV_X4 _u0_u27_U225  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[11] ) );
INV_X4 _u0_u27_U223  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[10] ) );
INV_X4 _u0_u27_U221  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[9] ) );
INV_X4 _u0_u27_U219  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[8] ) );
INV_X4 _u0_u27_U217  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[7] ) );
INV_X4 _u0_u27_U215  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[6] ) );
INV_X4 _u0_u27_U213  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[5] ) );
INV_X4 _u0_u27_U211  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[4] ) );
INV_X4 _u0_u27_U209  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[3] ) );
INV_X4 _u0_u27_U207  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[2] ) );
INV_X4 _u0_u27_U205  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[1] ) );
INV_X4 _u0_u27_U203  ( .A(1'b1), .ZN(_u0_u27_ch_adr1[0] ) );
INV_X4 _u0_u27_U201  ( .A(1'b0), .ZN(_u0_u27_ch_am0[31] ) );
INV_X4 _u0_u27_U199  ( .A(1'b0), .ZN(_u0_u27_ch_am0[30] ) );
INV_X4 _u0_u27_U197  ( .A(1'b0), .ZN(_u0_u27_ch_am0[29] ) );
INV_X4 _u0_u27_U195  ( .A(1'b0), .ZN(_u0_u27_ch_am0[28] ) );
INV_X4 _u0_u27_U193  ( .A(1'b0), .ZN(_u0_u27_ch_am0[27] ) );
INV_X4 _u0_u27_U191  ( .A(1'b0), .ZN(_u0_u27_ch_am0[26] ) );
INV_X4 _u0_u27_U189  ( .A(1'b0), .ZN(_u0_u27_ch_am0[25] ) );
INV_X4 _u0_u27_U187  ( .A(1'b0), .ZN(_u0_u27_ch_am0[24] ) );
INV_X4 _u0_u27_U185  ( .A(1'b0), .ZN(_u0_u27_ch_am0[23] ) );
INV_X4 _u0_u27_U183  ( .A(1'b0), .ZN(_u0_u27_ch_am0[22] ) );
INV_X4 _u0_u27_U181  ( .A(1'b0), .ZN(_u0_u27_ch_am0[21] ) );
INV_X4 _u0_u27_U179  ( .A(1'b0), .ZN(_u0_u27_ch_am0[20] ) );
INV_X4 _u0_u27_U177  ( .A(1'b0), .ZN(_u0_u27_ch_am0[19] ) );
INV_X4 _u0_u27_U175  ( .A(1'b0), .ZN(_u0_u27_ch_am0[18] ) );
INV_X4 _u0_u27_U173  ( .A(1'b0), .ZN(_u0_u27_ch_am0[17] ) );
INV_X4 _u0_u27_U171  ( .A(1'b0), .ZN(_u0_u27_ch_am0[16] ) );
INV_X4 _u0_u27_U169  ( .A(1'b0), .ZN(_u0_u27_ch_am0[15] ) );
INV_X4 _u0_u27_U167  ( .A(1'b0), .ZN(_u0_u27_ch_am0[14] ) );
INV_X4 _u0_u27_U165  ( .A(1'b0), .ZN(_u0_u27_ch_am0[13] ) );
INV_X4 _u0_u27_U163  ( .A(1'b0), .ZN(_u0_u27_ch_am0[12] ) );
INV_X4 _u0_u27_U161  ( .A(1'b0), .ZN(_u0_u27_ch_am0[11] ) );
INV_X4 _u0_u27_U159  ( .A(1'b0), .ZN(_u0_u27_ch_am0[10] ) );
INV_X4 _u0_u27_U157  ( .A(1'b0), .ZN(_u0_u27_ch_am0[9] ) );
INV_X4 _u0_u27_U155  ( .A(1'b0), .ZN(_u0_u27_ch_am0[8] ) );
INV_X4 _u0_u27_U153  ( .A(1'b0), .ZN(_u0_u27_ch_am0[7] ) );
INV_X4 _u0_u27_U151  ( .A(1'b0), .ZN(_u0_u27_ch_am0[6] ) );
INV_X4 _u0_u27_U149  ( .A(1'b0), .ZN(_u0_u27_ch_am0[5] ) );
INV_X4 _u0_u27_U147  ( .A(1'b0), .ZN(_u0_u27_ch_am0[4] ) );
INV_X4 _u0_u27_U145  ( .A(1'b1), .ZN(_u0_u27_ch_am0[3] ) );
INV_X4 _u0_u27_U143  ( .A(1'b1), .ZN(_u0_u27_ch_am0[2] ) );
INV_X4 _u0_u27_U141  ( .A(1'b1), .ZN(_u0_u27_ch_am0[1] ) );
INV_X4 _u0_u27_U139  ( .A(1'b1), .ZN(_u0_u27_ch_am0[0] ) );
INV_X4 _u0_u27_U137  ( .A(1'b0), .ZN(_u0_u27_ch_am1[31] ) );
INV_X4 _u0_u27_U135  ( .A(1'b0), .ZN(_u0_u27_ch_am1[30] ) );
INV_X4 _u0_u27_U133  ( .A(1'b0), .ZN(_u0_u27_ch_am1[29] ) );
INV_X4 _u0_u27_U131  ( .A(1'b0), .ZN(_u0_u27_ch_am1[28] ) );
INV_X4 _u0_u27_U129  ( .A(1'b0), .ZN(_u0_u27_ch_am1[27] ) );
INV_X4 _u0_u27_U127  ( .A(1'b0), .ZN(_u0_u27_ch_am1[26] ) );
INV_X4 _u0_u27_U125  ( .A(1'b0), .ZN(_u0_u27_ch_am1[25] ) );
INV_X4 _u0_u27_U123  ( .A(1'b0), .ZN(_u0_u27_ch_am1[24] ) );
INV_X4 _u0_u27_U121  ( .A(1'b0), .ZN(_u0_u27_ch_am1[23] ) );
INV_X4 _u0_u27_U119  ( .A(1'b0), .ZN(_u0_u27_ch_am1[22] ) );
INV_X4 _u0_u27_U117  ( .A(1'b0), .ZN(_u0_u27_ch_am1[21] ) );
INV_X4 _u0_u27_U115  ( .A(1'b0), .ZN(_u0_u27_ch_am1[20] ) );
INV_X4 _u0_u27_U113  ( .A(1'b0), .ZN(_u0_u27_ch_am1[19] ) );
INV_X4 _u0_u27_U111  ( .A(1'b0), .ZN(_u0_u27_ch_am1[18] ) );
INV_X4 _u0_u27_U109  ( .A(1'b0), .ZN(_u0_u27_ch_am1[17] ) );
INV_X4 _u0_u27_U107  ( .A(1'b0), .ZN(_u0_u27_ch_am1[16] ) );
INV_X4 _u0_u27_U105  ( .A(1'b0), .ZN(_u0_u27_ch_am1[15] ) );
INV_X4 _u0_u27_U103  ( .A(1'b0), .ZN(_u0_u27_ch_am1[14] ) );
INV_X4 _u0_u27_U101  ( .A(1'b0), .ZN(_u0_u27_ch_am1[13] ) );
INV_X4 _u0_u27_U99  ( .A(1'b0), .ZN(_u0_u27_ch_am1[12] ) );
INV_X4 _u0_u27_U97  ( .A(1'b0), .ZN(_u0_u27_ch_am1[11] ) );
INV_X4 _u0_u27_U95  ( .A(1'b0), .ZN(_u0_u27_ch_am1[10] ) );
INV_X4 _u0_u27_U93  ( .A(1'b0), .ZN(_u0_u27_ch_am1[9] ) );
INV_X4 _u0_u27_U91  ( .A(1'b0), .ZN(_u0_u27_ch_am1[8] ) );
INV_X4 _u0_u27_U89  ( .A(1'b0), .ZN(_u0_u27_ch_am1[7] ) );
INV_X4 _u0_u27_U87  ( .A(1'b0), .ZN(_u0_u27_ch_am1[6] ) );
INV_X4 _u0_u27_U85  ( .A(1'b0), .ZN(_u0_u27_ch_am1[5] ) );
INV_X4 _u0_u27_U83  ( .A(1'b0), .ZN(_u0_u27_ch_am1[4] ) );
INV_X4 _u0_u27_U81  ( .A(1'b1), .ZN(_u0_u27_ch_am1[3] ) );
INV_X4 _u0_u27_U79  ( .A(1'b1), .ZN(_u0_u27_ch_am1[2] ) );
INV_X4 _u0_u27_U77  ( .A(1'b1), .ZN(_u0_u27_ch_am1[1] ) );
INV_X4 _u0_u27_U75  ( .A(1'b1), .ZN(_u0_u27_ch_am1[0] ) );
INV_X4 _u0_u27_U73  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[31] ) );
INV_X4 _u0_u27_U71  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[30] ) );
INV_X4 _u0_u27_U69  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[29] ) );
INV_X4 _u0_u27_U67  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[28] ) );
INV_X4 _u0_u27_U65  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[27] ) );
INV_X4 _u0_u27_U63  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[26] ) );
INV_X4 _u0_u27_U61  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[25] ) );
INV_X4 _u0_u27_U59  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[24] ) );
INV_X4 _u0_u27_U57  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[23] ) );
INV_X4 _u0_u27_U55  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[22] ) );
INV_X4 _u0_u27_U53  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[21] ) );
INV_X4 _u0_u27_U51  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[20] ) );
INV_X4 _u0_u27_U49  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[19] ) );
INV_X4 _u0_u27_U47  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[18] ) );
INV_X4 _u0_u27_U45  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[17] ) );
INV_X4 _u0_u27_U43  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[16] ) );
INV_X4 _u0_u27_U41  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[15] ) );
INV_X4 _u0_u27_U39  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[14] ) );
INV_X4 _u0_u27_U37  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[13] ) );
INV_X4 _u0_u27_U35  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[12] ) );
INV_X4 _u0_u27_U33  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[11] ) );
INV_X4 _u0_u27_U31  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[10] ) );
INV_X4 _u0_u27_U29  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[9] ) );
INV_X4 _u0_u27_U27  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[8] ) );
INV_X4 _u0_u27_U25  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[7] ) );
INV_X4 _u0_u27_U23  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[6] ) );
INV_X4 _u0_u27_U21  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[5] ) );
INV_X4 _u0_u27_U19  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[4] ) );
INV_X4 _u0_u27_U17  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[3] ) );
INV_X4 _u0_u27_U15  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[2] ) );
INV_X4 _u0_u27_U13  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[1] ) );
INV_X4 _u0_u27_U11  ( .A(1'b1), .ZN(_u0_u27_sw_pointer[0] ) );
INV_X4 _u0_u27_U9  ( .A(1'b1), .ZN(_u0_u27_ch_stop ) );
INV_X4 _u0_u27_U7  ( .A(1'b1), .ZN(_u0_u27_ch_dis ) );
INV_X4 _u0_u27_U5  ( .A(1'b1), .ZN(_u0_u27_int ) );
INV_X4 _u0_u28_U585  ( .A(1'b1), .ZN(_u0_u28_pointer[31] ) );
INV_X4 _u0_u28_U583  ( .A(1'b1), .ZN(_u0_u28_pointer[30] ) );
INV_X4 _u0_u28_U581  ( .A(1'b1), .ZN(_u0_u28_pointer[29] ) );
INV_X4 _u0_u28_U579  ( .A(1'b1), .ZN(_u0_u28_pointer[28] ) );
INV_X4 _u0_u28_U577  ( .A(1'b1), .ZN(_u0_u28_pointer[27] ) );
INV_X4 _u0_u28_U575  ( .A(1'b1), .ZN(_u0_u28_pointer[26] ) );
INV_X4 _u0_u28_U573  ( .A(1'b1), .ZN(_u0_u28_pointer[25] ) );
INV_X4 _u0_u28_U571  ( .A(1'b1), .ZN(_u0_u28_pointer[24] ) );
INV_X4 _u0_u28_U569  ( .A(1'b1), .ZN(_u0_u28_pointer[23] ) );
INV_X4 _u0_u28_U567  ( .A(1'b1), .ZN(_u0_u28_pointer[22] ) );
INV_X4 _u0_u28_U565  ( .A(1'b1), .ZN(_u0_u28_pointer[21] ) );
INV_X4 _u0_u28_U563  ( .A(1'b1), .ZN(_u0_u28_pointer[20] ) );
INV_X4 _u0_u28_U561  ( .A(1'b1), .ZN(_u0_u28_pointer[19] ) );
INV_X4 _u0_u28_U559  ( .A(1'b1), .ZN(_u0_u28_pointer[18] ) );
INV_X4 _u0_u28_U557  ( .A(1'b1), .ZN(_u0_u28_pointer[17] ) );
INV_X4 _u0_u28_U555  ( .A(1'b1), .ZN(_u0_u28_pointer[16] ) );
INV_X4 _u0_u28_U553  ( .A(1'b1), .ZN(_u0_u28_pointer[15] ) );
INV_X4 _u0_u28_U551  ( .A(1'b1), .ZN(_u0_u28_pointer[14] ) );
INV_X4 _u0_u28_U549  ( .A(1'b1), .ZN(_u0_u28_pointer[13] ) );
INV_X4 _u0_u28_U547  ( .A(1'b1), .ZN(_u0_u28_pointer[12] ) );
INV_X4 _u0_u28_U545  ( .A(1'b1), .ZN(_u0_u28_pointer[11] ) );
INV_X4 _u0_u28_U543  ( .A(1'b1), .ZN(_u0_u28_pointer[10] ) );
INV_X4 _u0_u28_U541  ( .A(1'b1), .ZN(_u0_u28_pointer[9] ) );
INV_X4 _u0_u28_U539  ( .A(1'b1), .ZN(_u0_u28_pointer[8] ) );
INV_X4 _u0_u28_U537  ( .A(1'b1), .ZN(_u0_u28_pointer[7] ) );
INV_X4 _u0_u28_U535  ( .A(1'b1), .ZN(_u0_u28_pointer[6] ) );
INV_X4 _u0_u28_U533  ( .A(1'b1), .ZN(_u0_u28_pointer[5] ) );
INV_X4 _u0_u28_U531  ( .A(1'b1), .ZN(_u0_u28_pointer[4] ) );
INV_X4 _u0_u28_U529  ( .A(1'b1), .ZN(_u0_u28_pointer[3] ) );
INV_X4 _u0_u28_U527  ( .A(1'b1), .ZN(_u0_u28_pointer[2] ) );
INV_X4 _u0_u28_U525  ( .A(1'b1), .ZN(_u0_u28_pointer[1] ) );
INV_X4 _u0_u28_U523  ( .A(1'b1), .ZN(_u0_u28_pointer[0] ) );
INV_X4 _u0_u28_U521  ( .A(1'b1), .ZN(_u0_u28_pointer_s[31] ) );
INV_X4 _u0_u28_U519  ( .A(1'b1), .ZN(_u0_u28_pointer_s[30] ) );
INV_X4 _u0_u28_U517  ( .A(1'b1), .ZN(_u0_u28_pointer_s[29] ) );
INV_X4 _u0_u28_U515  ( .A(1'b1), .ZN(_u0_u28_pointer_s[28] ) );
INV_X4 _u0_u28_U513  ( .A(1'b1), .ZN(_u0_u28_pointer_s[27] ) );
INV_X4 _u0_u28_U511  ( .A(1'b1), .ZN(_u0_u28_pointer_s[26] ) );
INV_X4 _u0_u28_U509  ( .A(1'b1), .ZN(_u0_u28_pointer_s[25] ) );
INV_X4 _u0_u28_U507  ( .A(1'b1), .ZN(_u0_u28_pointer_s[24] ) );
INV_X4 _u0_u28_U505  ( .A(1'b1), .ZN(_u0_u28_pointer_s[23] ) );
INV_X4 _u0_u28_U503  ( .A(1'b1), .ZN(_u0_u28_pointer_s[22] ) );
INV_X4 _u0_u28_U501  ( .A(1'b1), .ZN(_u0_u28_pointer_s[21] ) );
INV_X4 _u0_u28_U499  ( .A(1'b1), .ZN(_u0_u28_pointer_s[20] ) );
INV_X4 _u0_u28_U497  ( .A(1'b1), .ZN(_u0_u28_pointer_s[19] ) );
INV_X4 _u0_u28_U495  ( .A(1'b1), .ZN(_u0_u28_pointer_s[18] ) );
INV_X4 _u0_u28_U493  ( .A(1'b1), .ZN(_u0_u28_pointer_s[17] ) );
INV_X4 _u0_u28_U491  ( .A(1'b1), .ZN(_u0_u28_pointer_s[16] ) );
INV_X4 _u0_u28_U489  ( .A(1'b1), .ZN(_u0_u28_pointer_s[15] ) );
INV_X4 _u0_u28_U487  ( .A(1'b1), .ZN(_u0_u28_pointer_s[14] ) );
INV_X4 _u0_u28_U485  ( .A(1'b1), .ZN(_u0_u28_pointer_s[13] ) );
INV_X4 _u0_u28_U483  ( .A(1'b1), .ZN(_u0_u28_pointer_s[12] ) );
INV_X4 _u0_u28_U481  ( .A(1'b1), .ZN(_u0_u28_pointer_s[11] ) );
INV_X4 _u0_u28_U479  ( .A(1'b1), .ZN(_u0_u28_pointer_s[10] ) );
INV_X4 _u0_u28_U477  ( .A(1'b1), .ZN(_u0_u28_pointer_s[9] ) );
INV_X4 _u0_u28_U475  ( .A(1'b1), .ZN(_u0_u28_pointer_s[8] ) );
INV_X4 _u0_u28_U473  ( .A(1'b1), .ZN(_u0_u28_pointer_s[7] ) );
INV_X4 _u0_u28_U471  ( .A(1'b1), .ZN(_u0_u28_pointer_s[6] ) );
INV_X4 _u0_u28_U469  ( .A(1'b1), .ZN(_u0_u28_pointer_s[5] ) );
INV_X4 _u0_u28_U467  ( .A(1'b1), .ZN(_u0_u28_pointer_s[4] ) );
INV_X4 _u0_u28_U465  ( .A(1'b1), .ZN(_u0_u28_pointer_s[3] ) );
INV_X4 _u0_u28_U463  ( .A(1'b1), .ZN(_u0_u28_pointer_s[2] ) );
INV_X4 _u0_u28_U461  ( .A(1'b1), .ZN(_u0_u28_pointer_s[1] ) );
INV_X4 _u0_u28_U459  ( .A(1'b1), .ZN(_u0_u28_pointer_s[0] ) );
INV_X4 _u0_u28_U457  ( .A(1'b1), .ZN(_u0_u28_ch_csr[31] ) );
INV_X4 _u0_u28_U455  ( .A(1'b1), .ZN(_u0_u28_ch_csr[30] ) );
INV_X4 _u0_u28_U453  ( .A(1'b1), .ZN(_u0_u28_ch_csr[29] ) );
INV_X4 _u0_u28_U451  ( .A(1'b1), .ZN(_u0_u28_ch_csr[28] ) );
INV_X4 _u0_u28_U449  ( .A(1'b1), .ZN(_u0_u28_ch_csr[27] ) );
INV_X4 _u0_u28_U447  ( .A(1'b1), .ZN(_u0_u28_ch_csr[26] ) );
INV_X4 _u0_u28_U445  ( .A(1'b1), .ZN(_u0_u28_ch_csr[25] ) );
INV_X4 _u0_u28_U443  ( .A(1'b1), .ZN(_u0_u28_ch_csr[24] ) );
INV_X4 _u0_u28_U441  ( .A(1'b1), .ZN(_u0_u28_ch_csr[23] ) );
INV_X4 _u0_u28_U439  ( .A(1'b1), .ZN(_u0_u28_ch_csr[22] ) );
INV_X4 _u0_u28_U437  ( .A(1'b1), .ZN(_u0_u28_ch_csr[21] ) );
INV_X4 _u0_u28_U435  ( .A(1'b1), .ZN(_u0_u28_ch_csr[20] ) );
INV_X4 _u0_u28_U433  ( .A(1'b1), .ZN(_u0_u28_ch_csr[19] ) );
INV_X4 _u0_u28_U431  ( .A(1'b1), .ZN(_u0_u28_ch_csr[18] ) );
INV_X4 _u0_u28_U429  ( .A(1'b1), .ZN(_u0_u28_ch_csr[17] ) );
INV_X4 _u0_u28_U427  ( .A(1'b1), .ZN(_u0_u28_ch_csr[16] ) );
INV_X4 _u0_u28_U425  ( .A(1'b1), .ZN(_u0_u28_ch_csr[15] ) );
INV_X4 _u0_u28_U423  ( .A(1'b1), .ZN(_u0_u28_ch_csr[14] ) );
INV_X4 _u0_u28_U421  ( .A(1'b1), .ZN(_u0_u28_ch_csr[13] ) );
INV_X4 _u0_u28_U419  ( .A(1'b1), .ZN(_u0_u28_ch_csr[12] ) );
INV_X4 _u0_u28_U417  ( .A(1'b1), .ZN(_u0_u28_ch_csr[11] ) );
INV_X4 _u0_u28_U415  ( .A(1'b1), .ZN(_u0_u28_ch_csr[10] ) );
INV_X4 _u0_u28_U413  ( .A(1'b1), .ZN(_u0_u28_ch_csr[9] ) );
INV_X4 _u0_u28_U411  ( .A(1'b1), .ZN(_u0_u28_ch_csr[8] ) );
INV_X4 _u0_u28_U409  ( .A(1'b1), .ZN(_u0_u28_ch_csr[7] ) );
INV_X4 _u0_u28_U407  ( .A(1'b1), .ZN(_u0_u28_ch_csr[6] ) );
INV_X4 _u0_u28_U405  ( .A(1'b1), .ZN(_u0_u28_ch_csr[5] ) );
INV_X4 _u0_u28_U403  ( .A(1'b1), .ZN(_u0_u28_ch_csr[4] ) );
INV_X4 _u0_u28_U401  ( .A(1'b1), .ZN(_u0_u28_ch_csr[3] ) );
INV_X4 _u0_u28_U399  ( .A(1'b1), .ZN(_u0_u28_ch_csr[2] ) );
INV_X4 _u0_u28_U397  ( .A(1'b1), .ZN(_u0_u28_ch_csr[1] ) );
INV_X4 _u0_u28_U395  ( .A(1'b1), .ZN(_u0_u28_ch_csr[0] ) );
INV_X4 _u0_u28_U393  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[31] ) );
INV_X4 _u0_u28_U391  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[30] ) );
INV_X4 _u0_u28_U389  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[29] ) );
INV_X4 _u0_u28_U387  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[28] ) );
INV_X4 _u0_u28_U385  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[27] ) );
INV_X4 _u0_u28_U383  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[26] ) );
INV_X4 _u0_u28_U381  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[25] ) );
INV_X4 _u0_u28_U379  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[24] ) );
INV_X4 _u0_u28_U377  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[23] ) );
INV_X4 _u0_u28_U375  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[22] ) );
INV_X4 _u0_u28_U373  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[21] ) );
INV_X4 _u0_u28_U371  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[20] ) );
INV_X4 _u0_u28_U369  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[19] ) );
INV_X4 _u0_u28_U367  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[18] ) );
INV_X4 _u0_u28_U365  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[17] ) );
INV_X4 _u0_u28_U363  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[16] ) );
INV_X4 _u0_u28_U361  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[15] ) );
INV_X4 _u0_u28_U359  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[14] ) );
INV_X4 _u0_u28_U357  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[13] ) );
INV_X4 _u0_u28_U355  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[12] ) );
INV_X4 _u0_u28_U353  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[11] ) );
INV_X4 _u0_u28_U351  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[10] ) );
INV_X4 _u0_u28_U349  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[9] ) );
INV_X4 _u0_u28_U347  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[8] ) );
INV_X4 _u0_u28_U345  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[7] ) );
INV_X4 _u0_u28_U343  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[6] ) );
INV_X4 _u0_u28_U341  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[5] ) );
INV_X4 _u0_u28_U339  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[4] ) );
INV_X4 _u0_u28_U337  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[3] ) );
INV_X4 _u0_u28_U335  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[2] ) );
INV_X4 _u0_u28_U333  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[1] ) );
INV_X4 _u0_u28_U331  ( .A(1'b1), .ZN(_u0_u28_ch_txsz[0] ) );
INV_X4 _u0_u28_U329  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[31] ) );
INV_X4 _u0_u28_U327  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[30] ) );
INV_X4 _u0_u28_U325  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[29] ) );
INV_X4 _u0_u28_U323  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[28] ) );
INV_X4 _u0_u28_U321  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[27] ) );
INV_X4 _u0_u28_U319  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[26] ) );
INV_X4 _u0_u28_U317  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[25] ) );
INV_X4 _u0_u28_U315  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[24] ) );
INV_X4 _u0_u28_U313  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[23] ) );
INV_X4 _u0_u28_U311  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[22] ) );
INV_X4 _u0_u28_U309  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[21] ) );
INV_X4 _u0_u28_U307  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[20] ) );
INV_X4 _u0_u28_U305  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[19] ) );
INV_X4 _u0_u28_U303  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[18] ) );
INV_X4 _u0_u28_U301  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[17] ) );
INV_X4 _u0_u28_U299  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[16] ) );
INV_X4 _u0_u28_U297  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[15] ) );
INV_X4 _u0_u28_U295  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[14] ) );
INV_X4 _u0_u28_U293  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[13] ) );
INV_X4 _u0_u28_U291  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[12] ) );
INV_X4 _u0_u28_U289  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[11] ) );
INV_X4 _u0_u28_U287  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[10] ) );
INV_X4 _u0_u28_U285  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[9] ) );
INV_X4 _u0_u28_U283  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[8] ) );
INV_X4 _u0_u28_U281  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[7] ) );
INV_X4 _u0_u28_U279  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[6] ) );
INV_X4 _u0_u28_U277  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[5] ) );
INV_X4 _u0_u28_U275  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[4] ) );
INV_X4 _u0_u28_U273  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[3] ) );
INV_X4 _u0_u28_U271  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[2] ) );
INV_X4 _u0_u28_U269  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[1] ) );
INV_X4 _u0_u28_U267  ( .A(1'b1), .ZN(_u0_u28_ch_adr0[0] ) );
INV_X4 _u0_u28_U265  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[31] ) );
INV_X4 _u0_u28_U263  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[30] ) );
INV_X4 _u0_u28_U261  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[29] ) );
INV_X4 _u0_u28_U259  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[28] ) );
INV_X4 _u0_u28_U257  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[27] ) );
INV_X4 _u0_u28_U255  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[26] ) );
INV_X4 _u0_u28_U253  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[25] ) );
INV_X4 _u0_u28_U251  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[24] ) );
INV_X4 _u0_u28_U249  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[23] ) );
INV_X4 _u0_u28_U247  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[22] ) );
INV_X4 _u0_u28_U245  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[21] ) );
INV_X4 _u0_u28_U243  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[20] ) );
INV_X4 _u0_u28_U241  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[19] ) );
INV_X4 _u0_u28_U239  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[18] ) );
INV_X4 _u0_u28_U237  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[17] ) );
INV_X4 _u0_u28_U235  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[16] ) );
INV_X4 _u0_u28_U233  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[15] ) );
INV_X4 _u0_u28_U231  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[14] ) );
INV_X4 _u0_u28_U229  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[13] ) );
INV_X4 _u0_u28_U227  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[12] ) );
INV_X4 _u0_u28_U225  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[11] ) );
INV_X4 _u0_u28_U223  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[10] ) );
INV_X4 _u0_u28_U221  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[9] ) );
INV_X4 _u0_u28_U219  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[8] ) );
INV_X4 _u0_u28_U217  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[7] ) );
INV_X4 _u0_u28_U215  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[6] ) );
INV_X4 _u0_u28_U213  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[5] ) );
INV_X4 _u0_u28_U211  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[4] ) );
INV_X4 _u0_u28_U209  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[3] ) );
INV_X4 _u0_u28_U207  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[2] ) );
INV_X4 _u0_u28_U205  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[1] ) );
INV_X4 _u0_u28_U203  ( .A(1'b1), .ZN(_u0_u28_ch_adr1[0] ) );
INV_X4 _u0_u28_U201  ( .A(1'b0), .ZN(_u0_u28_ch_am0[31] ) );
INV_X4 _u0_u28_U199  ( .A(1'b0), .ZN(_u0_u28_ch_am0[30] ) );
INV_X4 _u0_u28_U197  ( .A(1'b0), .ZN(_u0_u28_ch_am0[29] ) );
INV_X4 _u0_u28_U195  ( .A(1'b0), .ZN(_u0_u28_ch_am0[28] ) );
INV_X4 _u0_u28_U193  ( .A(1'b0), .ZN(_u0_u28_ch_am0[27] ) );
INV_X4 _u0_u28_U191  ( .A(1'b0), .ZN(_u0_u28_ch_am0[26] ) );
INV_X4 _u0_u28_U189  ( .A(1'b0), .ZN(_u0_u28_ch_am0[25] ) );
INV_X4 _u0_u28_U187  ( .A(1'b0), .ZN(_u0_u28_ch_am0[24] ) );
INV_X4 _u0_u28_U185  ( .A(1'b0), .ZN(_u0_u28_ch_am0[23] ) );
INV_X4 _u0_u28_U183  ( .A(1'b0), .ZN(_u0_u28_ch_am0[22] ) );
INV_X4 _u0_u28_U181  ( .A(1'b0), .ZN(_u0_u28_ch_am0[21] ) );
INV_X4 _u0_u28_U179  ( .A(1'b0), .ZN(_u0_u28_ch_am0[20] ) );
INV_X4 _u0_u28_U177  ( .A(1'b0), .ZN(_u0_u28_ch_am0[19] ) );
INV_X4 _u0_u28_U175  ( .A(1'b0), .ZN(_u0_u28_ch_am0[18] ) );
INV_X4 _u0_u28_U173  ( .A(1'b0), .ZN(_u0_u28_ch_am0[17] ) );
INV_X4 _u0_u28_U171  ( .A(1'b0), .ZN(_u0_u28_ch_am0[16] ) );
INV_X4 _u0_u28_U169  ( .A(1'b0), .ZN(_u0_u28_ch_am0[15] ) );
INV_X4 _u0_u28_U167  ( .A(1'b0), .ZN(_u0_u28_ch_am0[14] ) );
INV_X4 _u0_u28_U165  ( .A(1'b0), .ZN(_u0_u28_ch_am0[13] ) );
INV_X4 _u0_u28_U163  ( .A(1'b0), .ZN(_u0_u28_ch_am0[12] ) );
INV_X4 _u0_u28_U161  ( .A(1'b0), .ZN(_u0_u28_ch_am0[11] ) );
INV_X4 _u0_u28_U159  ( .A(1'b0), .ZN(_u0_u28_ch_am0[10] ) );
INV_X4 _u0_u28_U157  ( .A(1'b0), .ZN(_u0_u28_ch_am0[9] ) );
INV_X4 _u0_u28_U155  ( .A(1'b0), .ZN(_u0_u28_ch_am0[8] ) );
INV_X4 _u0_u28_U153  ( .A(1'b0), .ZN(_u0_u28_ch_am0[7] ) );
INV_X4 _u0_u28_U151  ( .A(1'b0), .ZN(_u0_u28_ch_am0[6] ) );
INV_X4 _u0_u28_U149  ( .A(1'b0), .ZN(_u0_u28_ch_am0[5] ) );
INV_X4 _u0_u28_U147  ( .A(1'b0), .ZN(_u0_u28_ch_am0[4] ) );
INV_X4 _u0_u28_U145  ( .A(1'b1), .ZN(_u0_u28_ch_am0[3] ) );
INV_X4 _u0_u28_U143  ( .A(1'b1), .ZN(_u0_u28_ch_am0[2] ) );
INV_X4 _u0_u28_U141  ( .A(1'b1), .ZN(_u0_u28_ch_am0[1] ) );
INV_X4 _u0_u28_U139  ( .A(1'b1), .ZN(_u0_u28_ch_am0[0] ) );
INV_X4 _u0_u28_U137  ( .A(1'b0), .ZN(_u0_u28_ch_am1[31] ) );
INV_X4 _u0_u28_U135  ( .A(1'b0), .ZN(_u0_u28_ch_am1[30] ) );
INV_X4 _u0_u28_U133  ( .A(1'b0), .ZN(_u0_u28_ch_am1[29] ) );
INV_X4 _u0_u28_U131  ( .A(1'b0), .ZN(_u0_u28_ch_am1[28] ) );
INV_X4 _u0_u28_U129  ( .A(1'b0), .ZN(_u0_u28_ch_am1[27] ) );
INV_X4 _u0_u28_U127  ( .A(1'b0), .ZN(_u0_u28_ch_am1[26] ) );
INV_X4 _u0_u28_U125  ( .A(1'b0), .ZN(_u0_u28_ch_am1[25] ) );
INV_X4 _u0_u28_U123  ( .A(1'b0), .ZN(_u0_u28_ch_am1[24] ) );
INV_X4 _u0_u28_U121  ( .A(1'b0), .ZN(_u0_u28_ch_am1[23] ) );
INV_X4 _u0_u28_U119  ( .A(1'b0), .ZN(_u0_u28_ch_am1[22] ) );
INV_X4 _u0_u28_U117  ( .A(1'b0), .ZN(_u0_u28_ch_am1[21] ) );
INV_X4 _u0_u28_U115  ( .A(1'b0), .ZN(_u0_u28_ch_am1[20] ) );
INV_X4 _u0_u28_U113  ( .A(1'b0), .ZN(_u0_u28_ch_am1[19] ) );
INV_X4 _u0_u28_U111  ( .A(1'b0), .ZN(_u0_u28_ch_am1[18] ) );
INV_X4 _u0_u28_U109  ( .A(1'b0), .ZN(_u0_u28_ch_am1[17] ) );
INV_X4 _u0_u28_U107  ( .A(1'b0), .ZN(_u0_u28_ch_am1[16] ) );
INV_X4 _u0_u28_U105  ( .A(1'b0), .ZN(_u0_u28_ch_am1[15] ) );
INV_X4 _u0_u28_U103  ( .A(1'b0), .ZN(_u0_u28_ch_am1[14] ) );
INV_X4 _u0_u28_U101  ( .A(1'b0), .ZN(_u0_u28_ch_am1[13] ) );
INV_X4 _u0_u28_U99  ( .A(1'b0), .ZN(_u0_u28_ch_am1[12] ) );
INV_X4 _u0_u28_U97  ( .A(1'b0), .ZN(_u0_u28_ch_am1[11] ) );
INV_X4 _u0_u28_U95  ( .A(1'b0), .ZN(_u0_u28_ch_am1[10] ) );
INV_X4 _u0_u28_U93  ( .A(1'b0), .ZN(_u0_u28_ch_am1[9] ) );
INV_X4 _u0_u28_U91  ( .A(1'b0), .ZN(_u0_u28_ch_am1[8] ) );
INV_X4 _u0_u28_U89  ( .A(1'b0), .ZN(_u0_u28_ch_am1[7] ) );
INV_X4 _u0_u28_U87  ( .A(1'b0), .ZN(_u0_u28_ch_am1[6] ) );
INV_X4 _u0_u28_U85  ( .A(1'b0), .ZN(_u0_u28_ch_am1[5] ) );
INV_X4 _u0_u28_U83  ( .A(1'b0), .ZN(_u0_u28_ch_am1[4] ) );
INV_X4 _u0_u28_U81  ( .A(1'b1), .ZN(_u0_u28_ch_am1[3] ) );
INV_X4 _u0_u28_U79  ( .A(1'b1), .ZN(_u0_u28_ch_am1[2] ) );
INV_X4 _u0_u28_U77  ( .A(1'b1), .ZN(_u0_u28_ch_am1[1] ) );
INV_X4 _u0_u28_U75  ( .A(1'b1), .ZN(_u0_u28_ch_am1[0] ) );
INV_X4 _u0_u28_U73  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[31] ) );
INV_X4 _u0_u28_U71  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[30] ) );
INV_X4 _u0_u28_U69  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[29] ) );
INV_X4 _u0_u28_U67  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[28] ) );
INV_X4 _u0_u28_U65  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[27] ) );
INV_X4 _u0_u28_U63  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[26] ) );
INV_X4 _u0_u28_U61  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[25] ) );
INV_X4 _u0_u28_U59  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[24] ) );
INV_X4 _u0_u28_U57  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[23] ) );
INV_X4 _u0_u28_U55  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[22] ) );
INV_X4 _u0_u28_U53  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[21] ) );
INV_X4 _u0_u28_U51  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[20] ) );
INV_X4 _u0_u28_U49  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[19] ) );
INV_X4 _u0_u28_U47  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[18] ) );
INV_X4 _u0_u28_U45  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[17] ) );
INV_X4 _u0_u28_U43  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[16] ) );
INV_X4 _u0_u28_U41  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[15] ) );
INV_X4 _u0_u28_U39  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[14] ) );
INV_X4 _u0_u28_U37  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[13] ) );
INV_X4 _u0_u28_U35  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[12] ) );
INV_X4 _u0_u28_U33  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[11] ) );
INV_X4 _u0_u28_U31  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[10] ) );
INV_X4 _u0_u28_U29  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[9] ) );
INV_X4 _u0_u28_U27  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[8] ) );
INV_X4 _u0_u28_U25  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[7] ) );
INV_X4 _u0_u28_U23  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[6] ) );
INV_X4 _u0_u28_U21  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[5] ) );
INV_X4 _u0_u28_U19  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[4] ) );
INV_X4 _u0_u28_U17  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[3] ) );
INV_X4 _u0_u28_U15  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[2] ) );
INV_X4 _u0_u28_U13  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[1] ) );
INV_X4 _u0_u28_U11  ( .A(1'b1), .ZN(_u0_u28_sw_pointer[0] ) );
INV_X4 _u0_u28_U9  ( .A(1'b1), .ZN(_u0_u28_ch_stop ) );
INV_X4 _u0_u28_U7  ( .A(1'b1), .ZN(_u0_u28_ch_dis ) );
INV_X4 _u0_u28_U5  ( .A(1'b1), .ZN(_u0_u28_int ) );
INV_X4 _u0_u29_U585  ( .A(1'b1), .ZN(_u0_u29_pointer[31] ) );
INV_X4 _u0_u29_U583  ( .A(1'b1), .ZN(_u0_u29_pointer[30] ) );
INV_X4 _u0_u29_U581  ( .A(1'b1), .ZN(_u0_u29_pointer[29] ) );
INV_X4 _u0_u29_U579  ( .A(1'b1), .ZN(_u0_u29_pointer[28] ) );
INV_X4 _u0_u29_U577  ( .A(1'b1), .ZN(_u0_u29_pointer[27] ) );
INV_X4 _u0_u29_U575  ( .A(1'b1), .ZN(_u0_u29_pointer[26] ) );
INV_X4 _u0_u29_U573  ( .A(1'b1), .ZN(_u0_u29_pointer[25] ) );
INV_X4 _u0_u29_U571  ( .A(1'b1), .ZN(_u0_u29_pointer[24] ) );
INV_X4 _u0_u29_U569  ( .A(1'b1), .ZN(_u0_u29_pointer[23] ) );
INV_X4 _u0_u29_U567  ( .A(1'b1), .ZN(_u0_u29_pointer[22] ) );
INV_X4 _u0_u29_U565  ( .A(1'b1), .ZN(_u0_u29_pointer[21] ) );
INV_X4 _u0_u29_U563  ( .A(1'b1), .ZN(_u0_u29_pointer[20] ) );
INV_X4 _u0_u29_U561  ( .A(1'b1), .ZN(_u0_u29_pointer[19] ) );
INV_X4 _u0_u29_U559  ( .A(1'b1), .ZN(_u0_u29_pointer[18] ) );
INV_X4 _u0_u29_U557  ( .A(1'b1), .ZN(_u0_u29_pointer[17] ) );
INV_X4 _u0_u29_U555  ( .A(1'b1), .ZN(_u0_u29_pointer[16] ) );
INV_X4 _u0_u29_U553  ( .A(1'b1), .ZN(_u0_u29_pointer[15] ) );
INV_X4 _u0_u29_U551  ( .A(1'b1), .ZN(_u0_u29_pointer[14] ) );
INV_X4 _u0_u29_U549  ( .A(1'b1), .ZN(_u0_u29_pointer[13] ) );
INV_X4 _u0_u29_U547  ( .A(1'b1), .ZN(_u0_u29_pointer[12] ) );
INV_X4 _u0_u29_U545  ( .A(1'b1), .ZN(_u0_u29_pointer[11] ) );
INV_X4 _u0_u29_U543  ( .A(1'b1), .ZN(_u0_u29_pointer[10] ) );
INV_X4 _u0_u29_U541  ( .A(1'b1), .ZN(_u0_u29_pointer[9] ) );
INV_X4 _u0_u29_U539  ( .A(1'b1), .ZN(_u0_u29_pointer[8] ) );
INV_X4 _u0_u29_U537  ( .A(1'b1), .ZN(_u0_u29_pointer[7] ) );
INV_X4 _u0_u29_U535  ( .A(1'b1), .ZN(_u0_u29_pointer[6] ) );
INV_X4 _u0_u29_U533  ( .A(1'b1), .ZN(_u0_u29_pointer[5] ) );
INV_X4 _u0_u29_U531  ( .A(1'b1), .ZN(_u0_u29_pointer[4] ) );
INV_X4 _u0_u29_U529  ( .A(1'b1), .ZN(_u0_u29_pointer[3] ) );
INV_X4 _u0_u29_U527  ( .A(1'b1), .ZN(_u0_u29_pointer[2] ) );
INV_X4 _u0_u29_U525  ( .A(1'b1), .ZN(_u0_u29_pointer[1] ) );
INV_X4 _u0_u29_U523  ( .A(1'b1), .ZN(_u0_u29_pointer[0] ) );
INV_X4 _u0_u29_U521  ( .A(1'b1), .ZN(_u0_u29_pointer_s[31] ) );
INV_X4 _u0_u29_U519  ( .A(1'b1), .ZN(_u0_u29_pointer_s[30] ) );
INV_X4 _u0_u29_U517  ( .A(1'b1), .ZN(_u0_u29_pointer_s[29] ) );
INV_X4 _u0_u29_U515  ( .A(1'b1), .ZN(_u0_u29_pointer_s[28] ) );
INV_X4 _u0_u29_U513  ( .A(1'b1), .ZN(_u0_u29_pointer_s[27] ) );
INV_X4 _u0_u29_U511  ( .A(1'b1), .ZN(_u0_u29_pointer_s[26] ) );
INV_X4 _u0_u29_U509  ( .A(1'b1), .ZN(_u0_u29_pointer_s[25] ) );
INV_X4 _u0_u29_U507  ( .A(1'b1), .ZN(_u0_u29_pointer_s[24] ) );
INV_X4 _u0_u29_U505  ( .A(1'b1), .ZN(_u0_u29_pointer_s[23] ) );
INV_X4 _u0_u29_U503  ( .A(1'b1), .ZN(_u0_u29_pointer_s[22] ) );
INV_X4 _u0_u29_U501  ( .A(1'b1), .ZN(_u0_u29_pointer_s[21] ) );
INV_X4 _u0_u29_U499  ( .A(1'b1), .ZN(_u0_u29_pointer_s[20] ) );
INV_X4 _u0_u29_U497  ( .A(1'b1), .ZN(_u0_u29_pointer_s[19] ) );
INV_X4 _u0_u29_U495  ( .A(1'b1), .ZN(_u0_u29_pointer_s[18] ) );
INV_X4 _u0_u29_U493  ( .A(1'b1), .ZN(_u0_u29_pointer_s[17] ) );
INV_X4 _u0_u29_U491  ( .A(1'b1), .ZN(_u0_u29_pointer_s[16] ) );
INV_X4 _u0_u29_U489  ( .A(1'b1), .ZN(_u0_u29_pointer_s[15] ) );
INV_X4 _u0_u29_U487  ( .A(1'b1), .ZN(_u0_u29_pointer_s[14] ) );
INV_X4 _u0_u29_U485  ( .A(1'b1), .ZN(_u0_u29_pointer_s[13] ) );
INV_X4 _u0_u29_U483  ( .A(1'b1), .ZN(_u0_u29_pointer_s[12] ) );
INV_X4 _u0_u29_U481  ( .A(1'b1), .ZN(_u0_u29_pointer_s[11] ) );
INV_X4 _u0_u29_U479  ( .A(1'b1), .ZN(_u0_u29_pointer_s[10] ) );
INV_X4 _u0_u29_U477  ( .A(1'b1), .ZN(_u0_u29_pointer_s[9] ) );
INV_X4 _u0_u29_U475  ( .A(1'b1), .ZN(_u0_u29_pointer_s[8] ) );
INV_X4 _u0_u29_U473  ( .A(1'b1), .ZN(_u0_u29_pointer_s[7] ) );
INV_X4 _u0_u29_U471  ( .A(1'b1), .ZN(_u0_u29_pointer_s[6] ) );
INV_X4 _u0_u29_U469  ( .A(1'b1), .ZN(_u0_u29_pointer_s[5] ) );
INV_X4 _u0_u29_U467  ( .A(1'b1), .ZN(_u0_u29_pointer_s[4] ) );
INV_X4 _u0_u29_U465  ( .A(1'b1), .ZN(_u0_u29_pointer_s[3] ) );
INV_X4 _u0_u29_U463  ( .A(1'b1), .ZN(_u0_u29_pointer_s[2] ) );
INV_X4 _u0_u29_U461  ( .A(1'b1), .ZN(_u0_u29_pointer_s[1] ) );
INV_X4 _u0_u29_U459  ( .A(1'b1), .ZN(_u0_u29_pointer_s[0] ) );
INV_X4 _u0_u29_U457  ( .A(1'b1), .ZN(_u0_u29_ch_csr[31] ) );
INV_X4 _u0_u29_U455  ( .A(1'b1), .ZN(_u0_u29_ch_csr[30] ) );
INV_X4 _u0_u29_U453  ( .A(1'b1), .ZN(_u0_u29_ch_csr[29] ) );
INV_X4 _u0_u29_U451  ( .A(1'b1), .ZN(_u0_u29_ch_csr[28] ) );
INV_X4 _u0_u29_U449  ( .A(1'b1), .ZN(_u0_u29_ch_csr[27] ) );
INV_X4 _u0_u29_U447  ( .A(1'b1), .ZN(_u0_u29_ch_csr[26] ) );
INV_X4 _u0_u29_U445  ( .A(1'b1), .ZN(_u0_u29_ch_csr[25] ) );
INV_X4 _u0_u29_U443  ( .A(1'b1), .ZN(_u0_u29_ch_csr[24] ) );
INV_X4 _u0_u29_U441  ( .A(1'b1), .ZN(_u0_u29_ch_csr[23] ) );
INV_X4 _u0_u29_U439  ( .A(1'b1), .ZN(_u0_u29_ch_csr[22] ) );
INV_X4 _u0_u29_U437  ( .A(1'b1), .ZN(_u0_u29_ch_csr[21] ) );
INV_X4 _u0_u29_U435  ( .A(1'b1), .ZN(_u0_u29_ch_csr[20] ) );
INV_X4 _u0_u29_U433  ( .A(1'b1), .ZN(_u0_u29_ch_csr[19] ) );
INV_X4 _u0_u29_U431  ( .A(1'b1), .ZN(_u0_u29_ch_csr[18] ) );
INV_X4 _u0_u29_U429  ( .A(1'b1), .ZN(_u0_u29_ch_csr[17] ) );
INV_X4 _u0_u29_U427  ( .A(1'b1), .ZN(_u0_u29_ch_csr[16] ) );
INV_X4 _u0_u29_U425  ( .A(1'b1), .ZN(_u0_u29_ch_csr[15] ) );
INV_X4 _u0_u29_U423  ( .A(1'b1), .ZN(_u0_u29_ch_csr[14] ) );
INV_X4 _u0_u29_U421  ( .A(1'b1), .ZN(_u0_u29_ch_csr[13] ) );
INV_X4 _u0_u29_U419  ( .A(1'b1), .ZN(_u0_u29_ch_csr[12] ) );
INV_X4 _u0_u29_U417  ( .A(1'b1), .ZN(_u0_u29_ch_csr[11] ) );
INV_X4 _u0_u29_U415  ( .A(1'b1), .ZN(_u0_u29_ch_csr[10] ) );
INV_X4 _u0_u29_U413  ( .A(1'b1), .ZN(_u0_u29_ch_csr[9] ) );
INV_X4 _u0_u29_U411  ( .A(1'b1), .ZN(_u0_u29_ch_csr[8] ) );
INV_X4 _u0_u29_U409  ( .A(1'b1), .ZN(_u0_u29_ch_csr[7] ) );
INV_X4 _u0_u29_U407  ( .A(1'b1), .ZN(_u0_u29_ch_csr[6] ) );
INV_X4 _u0_u29_U405  ( .A(1'b1), .ZN(_u0_u29_ch_csr[5] ) );
INV_X4 _u0_u29_U403  ( .A(1'b1), .ZN(_u0_u29_ch_csr[4] ) );
INV_X4 _u0_u29_U401  ( .A(1'b1), .ZN(_u0_u29_ch_csr[3] ) );
INV_X4 _u0_u29_U399  ( .A(1'b1), .ZN(_u0_u29_ch_csr[2] ) );
INV_X4 _u0_u29_U397  ( .A(1'b1), .ZN(_u0_u29_ch_csr[1] ) );
INV_X4 _u0_u29_U395  ( .A(1'b1), .ZN(_u0_u29_ch_csr[0] ) );
INV_X4 _u0_u29_U393  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[31] ) );
INV_X4 _u0_u29_U391  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[30] ) );
INV_X4 _u0_u29_U389  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[29] ) );
INV_X4 _u0_u29_U387  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[28] ) );
INV_X4 _u0_u29_U385  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[27] ) );
INV_X4 _u0_u29_U383  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[26] ) );
INV_X4 _u0_u29_U381  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[25] ) );
INV_X4 _u0_u29_U379  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[24] ) );
INV_X4 _u0_u29_U377  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[23] ) );
INV_X4 _u0_u29_U375  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[22] ) );
INV_X4 _u0_u29_U373  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[21] ) );
INV_X4 _u0_u29_U371  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[20] ) );
INV_X4 _u0_u29_U369  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[19] ) );
INV_X4 _u0_u29_U367  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[18] ) );
INV_X4 _u0_u29_U365  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[17] ) );
INV_X4 _u0_u29_U363  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[16] ) );
INV_X4 _u0_u29_U361  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[15] ) );
INV_X4 _u0_u29_U359  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[14] ) );
INV_X4 _u0_u29_U357  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[13] ) );
INV_X4 _u0_u29_U355  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[12] ) );
INV_X4 _u0_u29_U353  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[11] ) );
INV_X4 _u0_u29_U351  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[10] ) );
INV_X4 _u0_u29_U349  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[9] ) );
INV_X4 _u0_u29_U347  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[8] ) );
INV_X4 _u0_u29_U345  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[7] ) );
INV_X4 _u0_u29_U343  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[6] ) );
INV_X4 _u0_u29_U341  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[5] ) );
INV_X4 _u0_u29_U339  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[4] ) );
INV_X4 _u0_u29_U337  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[3] ) );
INV_X4 _u0_u29_U335  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[2] ) );
INV_X4 _u0_u29_U333  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[1] ) );
INV_X4 _u0_u29_U331  ( .A(1'b1), .ZN(_u0_u29_ch_txsz[0] ) );
INV_X4 _u0_u29_U329  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[31] ) );
INV_X4 _u0_u29_U327  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[30] ) );
INV_X4 _u0_u29_U325  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[29] ) );
INV_X4 _u0_u29_U323  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[28] ) );
INV_X4 _u0_u29_U321  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[27] ) );
INV_X4 _u0_u29_U319  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[26] ) );
INV_X4 _u0_u29_U317  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[25] ) );
INV_X4 _u0_u29_U315  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[24] ) );
INV_X4 _u0_u29_U313  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[23] ) );
INV_X4 _u0_u29_U311  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[22] ) );
INV_X4 _u0_u29_U309  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[21] ) );
INV_X4 _u0_u29_U307  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[20] ) );
INV_X4 _u0_u29_U305  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[19] ) );
INV_X4 _u0_u29_U303  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[18] ) );
INV_X4 _u0_u29_U301  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[17] ) );
INV_X4 _u0_u29_U299  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[16] ) );
INV_X4 _u0_u29_U297  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[15] ) );
INV_X4 _u0_u29_U295  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[14] ) );
INV_X4 _u0_u29_U293  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[13] ) );
INV_X4 _u0_u29_U291  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[12] ) );
INV_X4 _u0_u29_U289  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[11] ) );
INV_X4 _u0_u29_U287  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[10] ) );
INV_X4 _u0_u29_U285  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[9] ) );
INV_X4 _u0_u29_U283  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[8] ) );
INV_X4 _u0_u29_U281  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[7] ) );
INV_X4 _u0_u29_U279  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[6] ) );
INV_X4 _u0_u29_U277  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[5] ) );
INV_X4 _u0_u29_U275  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[4] ) );
INV_X4 _u0_u29_U273  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[3] ) );
INV_X4 _u0_u29_U271  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[2] ) );
INV_X4 _u0_u29_U269  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[1] ) );
INV_X4 _u0_u29_U267  ( .A(1'b1), .ZN(_u0_u29_ch_adr0[0] ) );
INV_X4 _u0_u29_U265  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[31] ) );
INV_X4 _u0_u29_U263  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[30] ) );
INV_X4 _u0_u29_U261  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[29] ) );
INV_X4 _u0_u29_U259  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[28] ) );
INV_X4 _u0_u29_U257  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[27] ) );
INV_X4 _u0_u29_U255  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[26] ) );
INV_X4 _u0_u29_U253  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[25] ) );
INV_X4 _u0_u29_U251  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[24] ) );
INV_X4 _u0_u29_U249  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[23] ) );
INV_X4 _u0_u29_U247  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[22] ) );
INV_X4 _u0_u29_U245  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[21] ) );
INV_X4 _u0_u29_U243  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[20] ) );
INV_X4 _u0_u29_U241  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[19] ) );
INV_X4 _u0_u29_U239  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[18] ) );
INV_X4 _u0_u29_U237  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[17] ) );
INV_X4 _u0_u29_U235  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[16] ) );
INV_X4 _u0_u29_U233  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[15] ) );
INV_X4 _u0_u29_U231  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[14] ) );
INV_X4 _u0_u29_U229  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[13] ) );
INV_X4 _u0_u29_U227  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[12] ) );
INV_X4 _u0_u29_U225  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[11] ) );
INV_X4 _u0_u29_U223  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[10] ) );
INV_X4 _u0_u29_U221  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[9] ) );
INV_X4 _u0_u29_U219  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[8] ) );
INV_X4 _u0_u29_U217  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[7] ) );
INV_X4 _u0_u29_U215  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[6] ) );
INV_X4 _u0_u29_U213  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[5] ) );
INV_X4 _u0_u29_U211  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[4] ) );
INV_X4 _u0_u29_U209  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[3] ) );
INV_X4 _u0_u29_U207  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[2] ) );
INV_X4 _u0_u29_U205  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[1] ) );
INV_X4 _u0_u29_U203  ( .A(1'b1), .ZN(_u0_u29_ch_adr1[0] ) );
INV_X4 _u0_u29_U201  ( .A(1'b0), .ZN(_u0_u29_ch_am0[31] ) );
INV_X4 _u0_u29_U199  ( .A(1'b0), .ZN(_u0_u29_ch_am0[30] ) );
INV_X4 _u0_u29_U197  ( .A(1'b0), .ZN(_u0_u29_ch_am0[29] ) );
INV_X4 _u0_u29_U195  ( .A(1'b0), .ZN(_u0_u29_ch_am0[28] ) );
INV_X4 _u0_u29_U193  ( .A(1'b0), .ZN(_u0_u29_ch_am0[27] ) );
INV_X4 _u0_u29_U191  ( .A(1'b0), .ZN(_u0_u29_ch_am0[26] ) );
INV_X4 _u0_u29_U189  ( .A(1'b0), .ZN(_u0_u29_ch_am0[25] ) );
INV_X4 _u0_u29_U187  ( .A(1'b0), .ZN(_u0_u29_ch_am0[24] ) );
INV_X4 _u0_u29_U185  ( .A(1'b0), .ZN(_u0_u29_ch_am0[23] ) );
INV_X4 _u0_u29_U183  ( .A(1'b0), .ZN(_u0_u29_ch_am0[22] ) );
INV_X4 _u0_u29_U181  ( .A(1'b0), .ZN(_u0_u29_ch_am0[21] ) );
INV_X4 _u0_u29_U179  ( .A(1'b0), .ZN(_u0_u29_ch_am0[20] ) );
INV_X4 _u0_u29_U177  ( .A(1'b0), .ZN(_u0_u29_ch_am0[19] ) );
INV_X4 _u0_u29_U175  ( .A(1'b0), .ZN(_u0_u29_ch_am0[18] ) );
INV_X4 _u0_u29_U173  ( .A(1'b0), .ZN(_u0_u29_ch_am0[17] ) );
INV_X4 _u0_u29_U171  ( .A(1'b0), .ZN(_u0_u29_ch_am0[16] ) );
INV_X4 _u0_u29_U169  ( .A(1'b0), .ZN(_u0_u29_ch_am0[15] ) );
INV_X4 _u0_u29_U167  ( .A(1'b0), .ZN(_u0_u29_ch_am0[14] ) );
INV_X4 _u0_u29_U165  ( .A(1'b0), .ZN(_u0_u29_ch_am0[13] ) );
INV_X4 _u0_u29_U163  ( .A(1'b0), .ZN(_u0_u29_ch_am0[12] ) );
INV_X4 _u0_u29_U161  ( .A(1'b0), .ZN(_u0_u29_ch_am0[11] ) );
INV_X4 _u0_u29_U159  ( .A(1'b0), .ZN(_u0_u29_ch_am0[10] ) );
INV_X4 _u0_u29_U157  ( .A(1'b0), .ZN(_u0_u29_ch_am0[9] ) );
INV_X4 _u0_u29_U155  ( .A(1'b0), .ZN(_u0_u29_ch_am0[8] ) );
INV_X4 _u0_u29_U153  ( .A(1'b0), .ZN(_u0_u29_ch_am0[7] ) );
INV_X4 _u0_u29_U151  ( .A(1'b0), .ZN(_u0_u29_ch_am0[6] ) );
INV_X4 _u0_u29_U149  ( .A(1'b0), .ZN(_u0_u29_ch_am0[5] ) );
INV_X4 _u0_u29_U147  ( .A(1'b0), .ZN(_u0_u29_ch_am0[4] ) );
INV_X4 _u0_u29_U145  ( .A(1'b1), .ZN(_u0_u29_ch_am0[3] ) );
INV_X4 _u0_u29_U143  ( .A(1'b1), .ZN(_u0_u29_ch_am0[2] ) );
INV_X4 _u0_u29_U141  ( .A(1'b1), .ZN(_u0_u29_ch_am0[1] ) );
INV_X4 _u0_u29_U139  ( .A(1'b1), .ZN(_u0_u29_ch_am0[0] ) );
INV_X4 _u0_u29_U137  ( .A(1'b0), .ZN(_u0_u29_ch_am1[31] ) );
INV_X4 _u0_u29_U135  ( .A(1'b0), .ZN(_u0_u29_ch_am1[30] ) );
INV_X4 _u0_u29_U133  ( .A(1'b0), .ZN(_u0_u29_ch_am1[29] ) );
INV_X4 _u0_u29_U131  ( .A(1'b0), .ZN(_u0_u29_ch_am1[28] ) );
INV_X4 _u0_u29_U129  ( .A(1'b0), .ZN(_u0_u29_ch_am1[27] ) );
INV_X4 _u0_u29_U127  ( .A(1'b0), .ZN(_u0_u29_ch_am1[26] ) );
INV_X4 _u0_u29_U125  ( .A(1'b0), .ZN(_u0_u29_ch_am1[25] ) );
INV_X4 _u0_u29_U123  ( .A(1'b0), .ZN(_u0_u29_ch_am1[24] ) );
INV_X4 _u0_u29_U121  ( .A(1'b0), .ZN(_u0_u29_ch_am1[23] ) );
INV_X4 _u0_u29_U119  ( .A(1'b0), .ZN(_u0_u29_ch_am1[22] ) );
INV_X4 _u0_u29_U117  ( .A(1'b0), .ZN(_u0_u29_ch_am1[21] ) );
INV_X4 _u0_u29_U115  ( .A(1'b0), .ZN(_u0_u29_ch_am1[20] ) );
INV_X4 _u0_u29_U113  ( .A(1'b0), .ZN(_u0_u29_ch_am1[19] ) );
INV_X4 _u0_u29_U111  ( .A(1'b0), .ZN(_u0_u29_ch_am1[18] ) );
INV_X4 _u0_u29_U109  ( .A(1'b0), .ZN(_u0_u29_ch_am1[17] ) );
INV_X4 _u0_u29_U107  ( .A(1'b0), .ZN(_u0_u29_ch_am1[16] ) );
INV_X4 _u0_u29_U105  ( .A(1'b0), .ZN(_u0_u29_ch_am1[15] ) );
INV_X4 _u0_u29_U103  ( .A(1'b0), .ZN(_u0_u29_ch_am1[14] ) );
INV_X4 _u0_u29_U101  ( .A(1'b0), .ZN(_u0_u29_ch_am1[13] ) );
INV_X4 _u0_u29_U99  ( .A(1'b0), .ZN(_u0_u29_ch_am1[12] ) );
INV_X4 _u0_u29_U97  ( .A(1'b0), .ZN(_u0_u29_ch_am1[11] ) );
INV_X4 _u0_u29_U95  ( .A(1'b0), .ZN(_u0_u29_ch_am1[10] ) );
INV_X4 _u0_u29_U93  ( .A(1'b0), .ZN(_u0_u29_ch_am1[9] ) );
INV_X4 _u0_u29_U91  ( .A(1'b0), .ZN(_u0_u29_ch_am1[8] ) );
INV_X4 _u0_u29_U89  ( .A(1'b0), .ZN(_u0_u29_ch_am1[7] ) );
INV_X4 _u0_u29_U87  ( .A(1'b0), .ZN(_u0_u29_ch_am1[6] ) );
INV_X4 _u0_u29_U85  ( .A(1'b0), .ZN(_u0_u29_ch_am1[5] ) );
INV_X4 _u0_u29_U83  ( .A(1'b0), .ZN(_u0_u29_ch_am1[4] ) );
INV_X4 _u0_u29_U81  ( .A(1'b1), .ZN(_u0_u29_ch_am1[3] ) );
INV_X4 _u0_u29_U79  ( .A(1'b1), .ZN(_u0_u29_ch_am1[2] ) );
INV_X4 _u0_u29_U77  ( .A(1'b1), .ZN(_u0_u29_ch_am1[1] ) );
INV_X4 _u0_u29_U75  ( .A(1'b1), .ZN(_u0_u29_ch_am1[0] ) );
INV_X4 _u0_u29_U73  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[31] ) );
INV_X4 _u0_u29_U71  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[30] ) );
INV_X4 _u0_u29_U69  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[29] ) );
INV_X4 _u0_u29_U67  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[28] ) );
INV_X4 _u0_u29_U65  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[27] ) );
INV_X4 _u0_u29_U63  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[26] ) );
INV_X4 _u0_u29_U61  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[25] ) );
INV_X4 _u0_u29_U59  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[24] ) );
INV_X4 _u0_u29_U57  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[23] ) );
INV_X4 _u0_u29_U55  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[22] ) );
INV_X4 _u0_u29_U53  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[21] ) );
INV_X4 _u0_u29_U51  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[20] ) );
INV_X4 _u0_u29_U49  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[19] ) );
INV_X4 _u0_u29_U47  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[18] ) );
INV_X4 _u0_u29_U45  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[17] ) );
INV_X4 _u0_u29_U43  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[16] ) );
INV_X4 _u0_u29_U41  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[15] ) );
INV_X4 _u0_u29_U39  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[14] ) );
INV_X4 _u0_u29_U37  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[13] ) );
INV_X4 _u0_u29_U35  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[12] ) );
INV_X4 _u0_u29_U33  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[11] ) );
INV_X4 _u0_u29_U31  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[10] ) );
INV_X4 _u0_u29_U29  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[9] ) );
INV_X4 _u0_u29_U27  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[8] ) );
INV_X4 _u0_u29_U25  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[7] ) );
INV_X4 _u0_u29_U23  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[6] ) );
INV_X4 _u0_u29_U21  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[5] ) );
INV_X4 _u0_u29_U19  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[4] ) );
INV_X4 _u0_u29_U17  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[3] ) );
INV_X4 _u0_u29_U15  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[2] ) );
INV_X4 _u0_u29_U13  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[1] ) );
INV_X4 _u0_u29_U11  ( .A(1'b1), .ZN(_u0_u29_sw_pointer[0] ) );
INV_X4 _u0_u29_U9  ( .A(1'b1), .ZN(_u0_u29_ch_stop ) );
INV_X4 _u0_u29_U7  ( .A(1'b1), .ZN(_u0_u29_ch_dis ) );
INV_X4 _u0_u29_U5  ( .A(1'b1), .ZN(_u0_u29_int ) );
INV_X4 _u0_u30_U585  ( .A(1'b1), .ZN(_u0_u30_pointer[31] ) );
INV_X4 _u0_u30_U583  ( .A(1'b1), .ZN(_u0_u30_pointer[30] ) );
INV_X4 _u0_u30_U581  ( .A(1'b1), .ZN(_u0_u30_pointer[29] ) );
INV_X4 _u0_u30_U579  ( .A(1'b1), .ZN(_u0_u30_pointer[28] ) );
INV_X4 _u0_u30_U577  ( .A(1'b1), .ZN(_u0_u30_pointer[27] ) );
INV_X4 _u0_u30_U575  ( .A(1'b1), .ZN(_u0_u30_pointer[26] ) );
INV_X4 _u0_u30_U573  ( .A(1'b1), .ZN(_u0_u30_pointer[25] ) );
INV_X4 _u0_u30_U571  ( .A(1'b1), .ZN(_u0_u30_pointer[24] ) );
INV_X4 _u0_u30_U569  ( .A(1'b1), .ZN(_u0_u30_pointer[23] ) );
INV_X4 _u0_u30_U567  ( .A(1'b1), .ZN(_u0_u30_pointer[22] ) );
INV_X4 _u0_u30_U565  ( .A(1'b1), .ZN(_u0_u30_pointer[21] ) );
INV_X4 _u0_u30_U563  ( .A(1'b1), .ZN(_u0_u30_pointer[20] ) );
INV_X4 _u0_u30_U561  ( .A(1'b1), .ZN(_u0_u30_pointer[19] ) );
INV_X4 _u0_u30_U559  ( .A(1'b1), .ZN(_u0_u30_pointer[18] ) );
INV_X4 _u0_u30_U557  ( .A(1'b1), .ZN(_u0_u30_pointer[17] ) );
INV_X4 _u0_u30_U555  ( .A(1'b1), .ZN(_u0_u30_pointer[16] ) );
INV_X4 _u0_u30_U553  ( .A(1'b1), .ZN(_u0_u30_pointer[15] ) );
INV_X4 _u0_u30_U551  ( .A(1'b1), .ZN(_u0_u30_pointer[14] ) );
INV_X4 _u0_u30_U549  ( .A(1'b1), .ZN(_u0_u30_pointer[13] ) );
INV_X4 _u0_u30_U547  ( .A(1'b1), .ZN(_u0_u30_pointer[12] ) );
INV_X4 _u0_u30_U545  ( .A(1'b1), .ZN(_u0_u30_pointer[11] ) );
INV_X4 _u0_u30_U543  ( .A(1'b1), .ZN(_u0_u30_pointer[10] ) );
INV_X4 _u0_u30_U541  ( .A(1'b1), .ZN(_u0_u30_pointer[9] ) );
INV_X4 _u0_u30_U539  ( .A(1'b1), .ZN(_u0_u30_pointer[8] ) );
INV_X4 _u0_u30_U537  ( .A(1'b1), .ZN(_u0_u30_pointer[7] ) );
INV_X4 _u0_u30_U535  ( .A(1'b1), .ZN(_u0_u30_pointer[6] ) );
INV_X4 _u0_u30_U533  ( .A(1'b1), .ZN(_u0_u30_pointer[5] ) );
INV_X4 _u0_u30_U531  ( .A(1'b1), .ZN(_u0_u30_pointer[4] ) );
INV_X4 _u0_u30_U529  ( .A(1'b1), .ZN(_u0_u30_pointer[3] ) );
INV_X4 _u0_u30_U527  ( .A(1'b1), .ZN(_u0_u30_pointer[2] ) );
INV_X4 _u0_u30_U525  ( .A(1'b1), .ZN(_u0_u30_pointer[1] ) );
INV_X4 _u0_u30_U523  ( .A(1'b1), .ZN(_u0_u30_pointer[0] ) );
INV_X4 _u0_u30_U521  ( .A(1'b1), .ZN(_u0_u30_pointer_s[31] ) );
INV_X4 _u0_u30_U519  ( .A(1'b1), .ZN(_u0_u30_pointer_s[30] ) );
INV_X4 _u0_u30_U517  ( .A(1'b1), .ZN(_u0_u30_pointer_s[29] ) );
INV_X4 _u0_u30_U515  ( .A(1'b1), .ZN(_u0_u30_pointer_s[28] ) );
INV_X4 _u0_u30_U513  ( .A(1'b1), .ZN(_u0_u30_pointer_s[27] ) );
INV_X4 _u0_u30_U511  ( .A(1'b1), .ZN(_u0_u30_pointer_s[26] ) );
INV_X4 _u0_u30_U509  ( .A(1'b1), .ZN(_u0_u30_pointer_s[25] ) );
INV_X4 _u0_u30_U507  ( .A(1'b1), .ZN(_u0_u30_pointer_s[24] ) );
INV_X4 _u0_u30_U505  ( .A(1'b1), .ZN(_u0_u30_pointer_s[23] ) );
INV_X4 _u0_u30_U503  ( .A(1'b1), .ZN(_u0_u30_pointer_s[22] ) );
INV_X4 _u0_u30_U501  ( .A(1'b1), .ZN(_u0_u30_pointer_s[21] ) );
INV_X4 _u0_u30_U499  ( .A(1'b1), .ZN(_u0_u30_pointer_s[20] ) );
INV_X4 _u0_u30_U497  ( .A(1'b1), .ZN(_u0_u30_pointer_s[19] ) );
INV_X4 _u0_u30_U495  ( .A(1'b1), .ZN(_u0_u30_pointer_s[18] ) );
INV_X4 _u0_u30_U493  ( .A(1'b1), .ZN(_u0_u30_pointer_s[17] ) );
INV_X4 _u0_u30_U491  ( .A(1'b1), .ZN(_u0_u30_pointer_s[16] ) );
INV_X4 _u0_u30_U489  ( .A(1'b1), .ZN(_u0_u30_pointer_s[15] ) );
INV_X4 _u0_u30_U487  ( .A(1'b1), .ZN(_u0_u30_pointer_s[14] ) );
INV_X4 _u0_u30_U485  ( .A(1'b1), .ZN(_u0_u30_pointer_s[13] ) );
INV_X4 _u0_u30_U483  ( .A(1'b1), .ZN(_u0_u30_pointer_s[12] ) );
INV_X4 _u0_u30_U481  ( .A(1'b1), .ZN(_u0_u30_pointer_s[11] ) );
INV_X4 _u0_u30_U479  ( .A(1'b1), .ZN(_u0_u30_pointer_s[10] ) );
INV_X4 _u0_u30_U477  ( .A(1'b1), .ZN(_u0_u30_pointer_s[9] ) );
INV_X4 _u0_u30_U475  ( .A(1'b1), .ZN(_u0_u30_pointer_s[8] ) );
INV_X4 _u0_u30_U473  ( .A(1'b1), .ZN(_u0_u30_pointer_s[7] ) );
INV_X4 _u0_u30_U471  ( .A(1'b1), .ZN(_u0_u30_pointer_s[6] ) );
INV_X4 _u0_u30_U469  ( .A(1'b1), .ZN(_u0_u30_pointer_s[5] ) );
INV_X4 _u0_u30_U467  ( .A(1'b1), .ZN(_u0_u30_pointer_s[4] ) );
INV_X4 _u0_u30_U465  ( .A(1'b1), .ZN(_u0_u30_pointer_s[3] ) );
INV_X4 _u0_u30_U463  ( .A(1'b1), .ZN(_u0_u30_pointer_s[2] ) );
INV_X4 _u0_u30_U461  ( .A(1'b1), .ZN(_u0_u30_pointer_s[1] ) );
INV_X4 _u0_u30_U459  ( .A(1'b1), .ZN(_u0_u30_pointer_s[0] ) );
INV_X4 _u0_u30_U457  ( .A(1'b1), .ZN(_u0_u30_ch_csr[31] ) );
INV_X4 _u0_u30_U455  ( .A(1'b1), .ZN(_u0_u30_ch_csr[30] ) );
INV_X4 _u0_u30_U453  ( .A(1'b1), .ZN(_u0_u30_ch_csr[29] ) );
INV_X4 _u0_u30_U451  ( .A(1'b1), .ZN(_u0_u30_ch_csr[28] ) );
INV_X4 _u0_u30_U449  ( .A(1'b1), .ZN(_u0_u30_ch_csr[27] ) );
INV_X4 _u0_u30_U447  ( .A(1'b1), .ZN(_u0_u30_ch_csr[26] ) );
INV_X4 _u0_u30_U445  ( .A(1'b1), .ZN(_u0_u30_ch_csr[25] ) );
INV_X4 _u0_u30_U443  ( .A(1'b1), .ZN(_u0_u30_ch_csr[24] ) );
INV_X4 _u0_u30_U441  ( .A(1'b1), .ZN(_u0_u30_ch_csr[23] ) );
INV_X4 _u0_u30_U439  ( .A(1'b1), .ZN(_u0_u30_ch_csr[22] ) );
INV_X4 _u0_u30_U437  ( .A(1'b1), .ZN(_u0_u30_ch_csr[21] ) );
INV_X4 _u0_u30_U435  ( .A(1'b1), .ZN(_u0_u30_ch_csr[20] ) );
INV_X4 _u0_u30_U433  ( .A(1'b1), .ZN(_u0_u30_ch_csr[19] ) );
INV_X4 _u0_u30_U431  ( .A(1'b1), .ZN(_u0_u30_ch_csr[18] ) );
INV_X4 _u0_u30_U429  ( .A(1'b1), .ZN(_u0_u30_ch_csr[17] ) );
INV_X4 _u0_u30_U427  ( .A(1'b1), .ZN(_u0_u30_ch_csr[16] ) );
INV_X4 _u0_u30_U425  ( .A(1'b1), .ZN(_u0_u30_ch_csr[15] ) );
INV_X4 _u0_u30_U423  ( .A(1'b1), .ZN(_u0_u30_ch_csr[14] ) );
INV_X4 _u0_u30_U421  ( .A(1'b1), .ZN(_u0_u30_ch_csr[13] ) );
INV_X4 _u0_u30_U419  ( .A(1'b1), .ZN(_u0_u30_ch_csr[12] ) );
INV_X4 _u0_u30_U417  ( .A(1'b1), .ZN(_u0_u30_ch_csr[11] ) );
INV_X4 _u0_u30_U415  ( .A(1'b1), .ZN(_u0_u30_ch_csr[10] ) );
INV_X4 _u0_u30_U413  ( .A(1'b1), .ZN(_u0_u30_ch_csr[9] ) );
INV_X4 _u0_u30_U411  ( .A(1'b1), .ZN(_u0_u30_ch_csr[8] ) );
INV_X4 _u0_u30_U409  ( .A(1'b1), .ZN(_u0_u30_ch_csr[7] ) );
INV_X4 _u0_u30_U407  ( .A(1'b1), .ZN(_u0_u30_ch_csr[6] ) );
INV_X4 _u0_u30_U405  ( .A(1'b1), .ZN(_u0_u30_ch_csr[5] ) );
INV_X4 _u0_u30_U403  ( .A(1'b1), .ZN(_u0_u30_ch_csr[4] ) );
INV_X4 _u0_u30_U401  ( .A(1'b1), .ZN(_u0_u30_ch_csr[3] ) );
INV_X4 _u0_u30_U399  ( .A(1'b1), .ZN(_u0_u30_ch_csr[2] ) );
INV_X4 _u0_u30_U397  ( .A(1'b1), .ZN(_u0_u30_ch_csr[1] ) );
INV_X4 _u0_u30_U395  ( .A(1'b1), .ZN(_u0_u30_ch_csr[0] ) );
INV_X4 _u0_u30_U393  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[31] ) );
INV_X4 _u0_u30_U391  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[30] ) );
INV_X4 _u0_u30_U389  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[29] ) );
INV_X4 _u0_u30_U387  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[28] ) );
INV_X4 _u0_u30_U385  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[27] ) );
INV_X4 _u0_u30_U383  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[26] ) );
INV_X4 _u0_u30_U381  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[25] ) );
INV_X4 _u0_u30_U379  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[24] ) );
INV_X4 _u0_u30_U377  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[23] ) );
INV_X4 _u0_u30_U375  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[22] ) );
INV_X4 _u0_u30_U373  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[21] ) );
INV_X4 _u0_u30_U371  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[20] ) );
INV_X4 _u0_u30_U369  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[19] ) );
INV_X4 _u0_u30_U367  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[18] ) );
INV_X4 _u0_u30_U365  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[17] ) );
INV_X4 _u0_u30_U363  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[16] ) );
INV_X4 _u0_u30_U361  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[15] ) );
INV_X4 _u0_u30_U359  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[14] ) );
INV_X4 _u0_u30_U357  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[13] ) );
INV_X4 _u0_u30_U355  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[12] ) );
INV_X4 _u0_u30_U353  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[11] ) );
INV_X4 _u0_u30_U351  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[10] ) );
INV_X4 _u0_u30_U349  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[9] ) );
INV_X4 _u0_u30_U347  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[8] ) );
INV_X4 _u0_u30_U345  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[7] ) );
INV_X4 _u0_u30_U343  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[6] ) );
INV_X4 _u0_u30_U341  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[5] ) );
INV_X4 _u0_u30_U339  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[4] ) );
INV_X4 _u0_u30_U337  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[3] ) );
INV_X4 _u0_u30_U335  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[2] ) );
INV_X4 _u0_u30_U333  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[1] ) );
INV_X4 _u0_u30_U331  ( .A(1'b1), .ZN(_u0_u30_ch_txsz[0] ) );
INV_X4 _u0_u30_U329  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[31] ) );
INV_X4 _u0_u30_U327  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[30] ) );
INV_X4 _u0_u30_U325  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[29] ) );
INV_X4 _u0_u30_U323  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[28] ) );
INV_X4 _u0_u30_U321  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[27] ) );
INV_X4 _u0_u30_U319  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[26] ) );
INV_X4 _u0_u30_U317  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[25] ) );
INV_X4 _u0_u30_U315  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[24] ) );
INV_X4 _u0_u30_U313  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[23] ) );
INV_X4 _u0_u30_U311  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[22] ) );
INV_X4 _u0_u30_U309  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[21] ) );
INV_X4 _u0_u30_U307  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[20] ) );
INV_X4 _u0_u30_U305  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[19] ) );
INV_X4 _u0_u30_U303  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[18] ) );
INV_X4 _u0_u30_U301  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[17] ) );
INV_X4 _u0_u30_U299  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[16] ) );
INV_X4 _u0_u30_U297  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[15] ) );
INV_X4 _u0_u30_U295  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[14] ) );
INV_X4 _u0_u30_U293  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[13] ) );
INV_X4 _u0_u30_U291  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[12] ) );
INV_X4 _u0_u30_U289  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[11] ) );
INV_X4 _u0_u30_U287  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[10] ) );
INV_X4 _u0_u30_U285  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[9] ) );
INV_X4 _u0_u30_U283  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[8] ) );
INV_X4 _u0_u30_U281  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[7] ) );
INV_X4 _u0_u30_U279  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[6] ) );
INV_X4 _u0_u30_U277  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[5] ) );
INV_X4 _u0_u30_U275  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[4] ) );
INV_X4 _u0_u30_U273  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[3] ) );
INV_X4 _u0_u30_U271  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[2] ) );
INV_X4 _u0_u30_U269  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[1] ) );
INV_X4 _u0_u30_U267  ( .A(1'b1), .ZN(_u0_u30_ch_adr0[0] ) );
INV_X4 _u0_u30_U265  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[31] ) );
INV_X4 _u0_u30_U263  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[30] ) );
INV_X4 _u0_u30_U261  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[29] ) );
INV_X4 _u0_u30_U259  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[28] ) );
INV_X4 _u0_u30_U257  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[27] ) );
INV_X4 _u0_u30_U255  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[26] ) );
INV_X4 _u0_u30_U253  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[25] ) );
INV_X4 _u0_u30_U251  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[24] ) );
INV_X4 _u0_u30_U249  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[23] ) );
INV_X4 _u0_u30_U247  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[22] ) );
INV_X4 _u0_u30_U245  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[21] ) );
INV_X4 _u0_u30_U243  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[20] ) );
INV_X4 _u0_u30_U241  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[19] ) );
INV_X4 _u0_u30_U239  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[18] ) );
INV_X4 _u0_u30_U237  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[17] ) );
INV_X4 _u0_u30_U235  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[16] ) );
INV_X4 _u0_u30_U233  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[15] ) );
INV_X4 _u0_u30_U231  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[14] ) );
INV_X4 _u0_u30_U229  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[13] ) );
INV_X4 _u0_u30_U227  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[12] ) );
INV_X4 _u0_u30_U225  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[11] ) );
INV_X4 _u0_u30_U223  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[10] ) );
INV_X4 _u0_u30_U221  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[9] ) );
INV_X4 _u0_u30_U219  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[8] ) );
INV_X4 _u0_u30_U217  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[7] ) );
INV_X4 _u0_u30_U215  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[6] ) );
INV_X4 _u0_u30_U213  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[5] ) );
INV_X4 _u0_u30_U211  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[4] ) );
INV_X4 _u0_u30_U209  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[3] ) );
INV_X4 _u0_u30_U207  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[2] ) );
INV_X4 _u0_u30_U205  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[1] ) );
INV_X4 _u0_u30_U203  ( .A(1'b1), .ZN(_u0_u30_ch_adr1[0] ) );
INV_X4 _u0_u30_U201  ( .A(1'b0), .ZN(_u0_u30_ch_am0[31] ) );
INV_X4 _u0_u30_U199  ( .A(1'b0), .ZN(_u0_u30_ch_am0[30] ) );
INV_X4 _u0_u30_U197  ( .A(1'b0), .ZN(_u0_u30_ch_am0[29] ) );
INV_X4 _u0_u30_U195  ( .A(1'b0), .ZN(_u0_u30_ch_am0[28] ) );
INV_X4 _u0_u30_U193  ( .A(1'b0), .ZN(_u0_u30_ch_am0[27] ) );
INV_X4 _u0_u30_U191  ( .A(1'b0), .ZN(_u0_u30_ch_am0[26] ) );
INV_X4 _u0_u30_U189  ( .A(1'b0), .ZN(_u0_u30_ch_am0[25] ) );
INV_X4 _u0_u30_U187  ( .A(1'b0), .ZN(_u0_u30_ch_am0[24] ) );
INV_X4 _u0_u30_U185  ( .A(1'b0), .ZN(_u0_u30_ch_am0[23] ) );
INV_X4 _u0_u30_U183  ( .A(1'b0), .ZN(_u0_u30_ch_am0[22] ) );
INV_X4 _u0_u30_U181  ( .A(1'b0), .ZN(_u0_u30_ch_am0[21] ) );
INV_X4 _u0_u30_U179  ( .A(1'b0), .ZN(_u0_u30_ch_am0[20] ) );
INV_X4 _u0_u30_U177  ( .A(1'b0), .ZN(_u0_u30_ch_am0[19] ) );
INV_X4 _u0_u30_U175  ( .A(1'b0), .ZN(_u0_u30_ch_am0[18] ) );
INV_X4 _u0_u30_U173  ( .A(1'b0), .ZN(_u0_u30_ch_am0[17] ) );
INV_X4 _u0_u30_U171  ( .A(1'b0), .ZN(_u0_u30_ch_am0[16] ) );
INV_X4 _u0_u30_U169  ( .A(1'b0), .ZN(_u0_u30_ch_am0[15] ) );
INV_X4 _u0_u30_U167  ( .A(1'b0), .ZN(_u0_u30_ch_am0[14] ) );
INV_X4 _u0_u30_U165  ( .A(1'b0), .ZN(_u0_u30_ch_am0[13] ) );
INV_X4 _u0_u30_U163  ( .A(1'b0), .ZN(_u0_u30_ch_am0[12] ) );
INV_X4 _u0_u30_U161  ( .A(1'b0), .ZN(_u0_u30_ch_am0[11] ) );
INV_X4 _u0_u30_U159  ( .A(1'b0), .ZN(_u0_u30_ch_am0[10] ) );
INV_X4 _u0_u30_U157  ( .A(1'b0), .ZN(_u0_u30_ch_am0[9] ) );
INV_X4 _u0_u30_U155  ( .A(1'b0), .ZN(_u0_u30_ch_am0[8] ) );
INV_X4 _u0_u30_U153  ( .A(1'b0), .ZN(_u0_u30_ch_am0[7] ) );
INV_X4 _u0_u30_U151  ( .A(1'b0), .ZN(_u0_u30_ch_am0[6] ) );
INV_X4 _u0_u30_U149  ( .A(1'b0), .ZN(_u0_u30_ch_am0[5] ) );
INV_X4 _u0_u30_U147  ( .A(1'b0), .ZN(_u0_u30_ch_am0[4] ) );
INV_X4 _u0_u30_U145  ( .A(1'b1), .ZN(_u0_u30_ch_am0[3] ) );
INV_X4 _u0_u30_U143  ( .A(1'b1), .ZN(_u0_u30_ch_am0[2] ) );
INV_X4 _u0_u30_U141  ( .A(1'b1), .ZN(_u0_u30_ch_am0[1] ) );
INV_X4 _u0_u30_U139  ( .A(1'b1), .ZN(_u0_u30_ch_am0[0] ) );
INV_X4 _u0_u30_U137  ( .A(1'b0), .ZN(_u0_u30_ch_am1[31] ) );
INV_X4 _u0_u30_U135  ( .A(1'b0), .ZN(_u0_u30_ch_am1[30] ) );
INV_X4 _u0_u30_U133  ( .A(1'b0), .ZN(_u0_u30_ch_am1[29] ) );
INV_X4 _u0_u30_U131  ( .A(1'b0), .ZN(_u0_u30_ch_am1[28] ) );
INV_X4 _u0_u30_U129  ( .A(1'b0), .ZN(_u0_u30_ch_am1[27] ) );
INV_X4 _u0_u30_U127  ( .A(1'b0), .ZN(_u0_u30_ch_am1[26] ) );
INV_X4 _u0_u30_U125  ( .A(1'b0), .ZN(_u0_u30_ch_am1[25] ) );
INV_X4 _u0_u30_U123  ( .A(1'b0), .ZN(_u0_u30_ch_am1[24] ) );
INV_X4 _u0_u30_U121  ( .A(1'b0), .ZN(_u0_u30_ch_am1[23] ) );
INV_X4 _u0_u30_U119  ( .A(1'b0), .ZN(_u0_u30_ch_am1[22] ) );
INV_X4 _u0_u30_U117  ( .A(1'b0), .ZN(_u0_u30_ch_am1[21] ) );
INV_X4 _u0_u30_U115  ( .A(1'b0), .ZN(_u0_u30_ch_am1[20] ) );
INV_X4 _u0_u30_U113  ( .A(1'b0), .ZN(_u0_u30_ch_am1[19] ) );
INV_X4 _u0_u30_U111  ( .A(1'b0), .ZN(_u0_u30_ch_am1[18] ) );
INV_X4 _u0_u30_U109  ( .A(1'b0), .ZN(_u0_u30_ch_am1[17] ) );
INV_X4 _u0_u30_U107  ( .A(1'b0), .ZN(_u0_u30_ch_am1[16] ) );
INV_X4 _u0_u30_U105  ( .A(1'b0), .ZN(_u0_u30_ch_am1[15] ) );
INV_X4 _u0_u30_U103  ( .A(1'b0), .ZN(_u0_u30_ch_am1[14] ) );
INV_X4 _u0_u30_U101  ( .A(1'b0), .ZN(_u0_u30_ch_am1[13] ) );
INV_X4 _u0_u30_U99  ( .A(1'b0), .ZN(_u0_u30_ch_am1[12] ) );
INV_X4 _u0_u30_U97  ( .A(1'b0), .ZN(_u0_u30_ch_am1[11] ) );
INV_X4 _u0_u30_U95  ( .A(1'b0), .ZN(_u0_u30_ch_am1[10] ) );
INV_X4 _u0_u30_U93  ( .A(1'b0), .ZN(_u0_u30_ch_am1[9] ) );
INV_X4 _u0_u30_U91  ( .A(1'b0), .ZN(_u0_u30_ch_am1[8] ) );
INV_X4 _u0_u30_U89  ( .A(1'b0), .ZN(_u0_u30_ch_am1[7] ) );
INV_X4 _u0_u30_U87  ( .A(1'b0), .ZN(_u0_u30_ch_am1[6] ) );
INV_X4 _u0_u30_U85  ( .A(1'b0), .ZN(_u0_u30_ch_am1[5] ) );
INV_X4 _u0_u30_U83  ( .A(1'b0), .ZN(_u0_u30_ch_am1[4] ) );
INV_X4 _u0_u30_U81  ( .A(1'b1), .ZN(_u0_u30_ch_am1[3] ) );
INV_X4 _u0_u30_U79  ( .A(1'b1), .ZN(_u0_u30_ch_am1[2] ) );
INV_X4 _u0_u30_U77  ( .A(1'b1), .ZN(_u0_u30_ch_am1[1] ) );
INV_X4 _u0_u30_U75  ( .A(1'b1), .ZN(_u0_u30_ch_am1[0] ) );
INV_X4 _u0_u30_U73  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[31] ) );
INV_X4 _u0_u30_U71  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[30] ) );
INV_X4 _u0_u30_U69  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[29] ) );
INV_X4 _u0_u30_U67  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[28] ) );
INV_X4 _u0_u30_U65  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[27] ) );
INV_X4 _u0_u30_U63  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[26] ) );
INV_X4 _u0_u30_U61  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[25] ) );
INV_X4 _u0_u30_U59  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[24] ) );
INV_X4 _u0_u30_U57  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[23] ) );
INV_X4 _u0_u30_U55  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[22] ) );
INV_X4 _u0_u30_U53  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[21] ) );
INV_X4 _u0_u30_U51  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[20] ) );
INV_X4 _u0_u30_U49  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[19] ) );
INV_X4 _u0_u30_U47  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[18] ) );
INV_X4 _u0_u30_U45  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[17] ) );
INV_X4 _u0_u30_U43  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[16] ) );
INV_X4 _u0_u30_U41  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[15] ) );
INV_X4 _u0_u30_U39  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[14] ) );
INV_X4 _u0_u30_U37  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[13] ) );
INV_X4 _u0_u30_U35  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[12] ) );
INV_X4 _u0_u30_U33  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[11] ) );
INV_X4 _u0_u30_U31  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[10] ) );
INV_X4 _u0_u30_U29  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[9] ) );
INV_X4 _u0_u30_U27  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[8] ) );
INV_X4 _u0_u30_U25  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[7] ) );
INV_X4 _u0_u30_U23  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[6] ) );
INV_X4 _u0_u30_U21  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[5] ) );
INV_X4 _u0_u30_U19  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[4] ) );
INV_X4 _u0_u30_U17  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[3] ) );
INV_X4 _u0_u30_U15  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[2] ) );
INV_X4 _u0_u30_U13  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[1] ) );
INV_X4 _u0_u30_U11  ( .A(1'b1), .ZN(_u0_u30_sw_pointer[0] ) );
INV_X4 _u0_u30_U9  ( .A(1'b1), .ZN(_u0_u30_ch_stop ) );
INV_X4 _u0_u30_U7  ( .A(1'b1), .ZN(_u0_u30_ch_dis ) );
INV_X4 _u0_u30_U5  ( .A(1'b1), .ZN(_u0_u30_int ) );
AND2_X1 _u10_U11803  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N1000 ) );
INV_X1 _u10_U11802  ( .A(1'b0), .ZN(_u10_n22987 ) );
NOR2_X1 _u10_U11801  ( .A1(1'b0), .A2(_u10_n22987 ), .ZN(_u10_N1002 ) );
INV_X1 _u10_U11800  ( .A(1'b0), .ZN(_u10_n22986 ) );
NOR2_X1 _u10_U11799  ( .A1(1'b0), .A2(_u10_n22986 ), .ZN(_u10_N1003 ) );
INV_X1 _u10_U11798  ( .A(1'b0), .ZN(_u10_n22985 ) );
NOR2_X1 _u10_U11797  ( .A1(1'b0), .A2(_u10_n22985 ), .ZN(_u10_N1004 ) );
INV_X1 _u10_U11796  ( .A(1'b0), .ZN(_u10_n22984 ) );
NOR2_X1 _u10_U11795  ( .A1(1'b0), .A2(_u10_n22984 ), .ZN(_u10_N1005 ) );
INV_X1 _u10_U11794  ( .A(1'b0), .ZN(_u10_n22983 ) );
NOR2_X1 _u10_U11793  ( .A1(1'b0), .A2(_u10_n22983 ), .ZN(_u10_N1006 ) );
INV_X1 _u10_U11792  ( .A(1'b0), .ZN(_u10_n22982 ) );
NOR2_X1 _u10_U11791  ( .A1(1'b0), .A2(_u10_n22982 ), .ZN(_u10_N1007 ) );
INV_X1 _u10_U11790  ( .A(1'b0), .ZN(_u10_n22981 ) );
NOR2_X1 _u10_U11789  ( .A1(1'b0), .A2(_u10_n22981 ), .ZN(_u10_N1008 ) );
INV_X1 _u10_U11788  ( .A(1'b0), .ZN(_u10_n22980 ) );
NOR2_X1 _u10_U11787  ( .A1(1'b0), .A2(_u10_n22980 ), .ZN(_u10_N1009 ) );
INV_X1 _u10_U11786  ( .A(1'b0), .ZN(_u10_n22979 ) );
NOR2_X1 _u10_U11785  ( .A1(1'b0), .A2(_u10_n22979 ), .ZN(_u10_N1010 ) );
INV_X1 _u10_U11784  ( .A(1'b0), .ZN(_u10_n22978 ) );
NOR2_X1 _u10_U11783  ( .A1(1'b0), .A2(_u10_n22978 ), .ZN(_u10_N1011 ) );
INV_X1 _u10_U11782  ( .A(1'b0), .ZN(_u10_n22977 ) );
NOR2_X1 _u10_U11781  ( .A1(1'b0), .A2(_u10_n22977 ), .ZN(_u10_N1012 ) );
INV_X1 _u10_U11780  ( .A(1'b0), .ZN(_u10_n22976 ) );
NOR2_X1 _u10_U11779  ( .A1(1'b0), .A2(_u10_n22976 ), .ZN(_u10_N1013 ) );
INV_X1 _u10_U11778  ( .A(1'b0), .ZN(_u10_n22975 ) );
NOR2_X1 _u10_U11777  ( .A1(1'b0), .A2(_u10_n22975 ), .ZN(_u10_N1014 ) );
INV_X1 _u10_U11776  ( .A(1'b0), .ZN(_u10_n22974 ) );
NOR2_X1 _u10_U11775  ( .A1(1'b0), .A2(_u10_n22974 ), .ZN(_u10_N1015 ) );
INV_X1 _u10_U11774  ( .A(1'b0), .ZN(_u10_n22973 ) );
NOR2_X1 _u10_U11773  ( .A1(1'b0), .A2(_u10_n22973 ), .ZN(_u10_N1016 ) );
INV_X1 _u10_U11772  ( .A(1'b0), .ZN(_u10_n22972 ) );
NOR2_X1 _u10_U11771  ( .A1(1'b0), .A2(_u10_n22972 ), .ZN(_u10_N1017 ) );
INV_X1 _u10_U11770  ( .A(1'b0), .ZN(_u10_n22971 ) );
NOR2_X1 _u10_U11769  ( .A1(1'b0), .A2(_u10_n22971 ), .ZN(_u10_N1018 ) );
INV_X1 _u10_U11768  ( .A(1'b0), .ZN(_u10_n22970 ) );
NOR2_X1 _u10_U11767  ( .A1(1'b0), .A2(_u10_n22970 ), .ZN(_u10_N1019 ) );
INV_X1 _u10_U11766  ( .A(1'b0), .ZN(_u10_n22969 ) );
NOR2_X1 _u10_U11765  ( .A1(1'b0), .A2(_u10_n22969 ), .ZN(_u10_N1020 ) );
INV_X1 _u10_U11764  ( .A(1'b0), .ZN(_u10_n22968 ) );
NOR2_X1 _u10_U11763  ( .A1(1'b0), .A2(_u10_n22968 ), .ZN(_u10_N1021 ) );
INV_X1 _u10_U11762  ( .A(1'b0), .ZN(_u10_n22967 ) );
NOR2_X1 _u10_U11761  ( .A1(1'b0), .A2(_u10_n22967 ), .ZN(_u10_N1022 ) );
INV_X1 _u10_U11760  ( .A(1'b0), .ZN(_u10_n22966 ) );
NOR2_X1 _u10_U11759  ( .A1(1'b0), .A2(_u10_n22966 ), .ZN(_u10_N1023 ) );
INV_X1 _u10_U11758  ( .A(1'b0), .ZN(_u10_n22965 ) );
NOR2_X1 _u10_U11757  ( .A1(1'b0), .A2(_u10_n22965 ), .ZN(_u10_N1024 ) );
INV_X1 _u10_U11756  ( .A(1'b0), .ZN(_u10_n22964 ) );
NOR2_X1 _u10_U11755  ( .A1(1'b0), .A2(_u10_n22964 ), .ZN(_u10_N1025 ) );
INV_X1 _u10_U11754  ( .A(1'b0), .ZN(_u10_n22963 ) );
NOR2_X1 _u10_U11753  ( .A1(1'b0), .A2(_u10_n22963 ), .ZN(_u10_N1026 ) );
INV_X1 _u10_U11752  ( .A(1'b0), .ZN(_u10_n22962 ) );
NOR2_X1 _u10_U11751  ( .A1(1'b0), .A2(_u10_n22962 ), .ZN(_u10_N1027 ) );
INV_X1 _u10_U11750  ( .A(1'b0), .ZN(_u10_n22961 ) );
NOR2_X1 _u10_U11749  ( .A1(1'b0), .A2(_u10_n22961 ), .ZN(_u10_N1028 ) );
INV_X1 _u10_U11748  ( .A(1'b0), .ZN(_u10_n22960 ) );
NOR2_X1 _u10_U11747  ( .A1(1'b0), .A2(_u10_n22960 ), .ZN(_u10_N1029 ) );
INV_X1 _u10_U11746  ( .A(1'b0), .ZN(_u10_n22959 ) );
NOR2_X1 _u10_U11745  ( .A1(1'b0), .A2(_u10_n22959 ), .ZN(_u10_N1030 ) );
INV_X1 _u10_U11744  ( .A(1'b0), .ZN(_u10_n22958 ) );
NOR2_X1 _u10_U11743  ( .A1(1'b0), .A2(_u10_n22958 ), .ZN(_u10_N1031 ) );
INV_X1 _u10_U11742  ( .A(dma_req_i[0]), .ZN(_u10_n23001 ) );
AND2_X1 _u10_U11741  ( .A1(dma_nd_i[0]), .A2(_u10_n23001 ), .ZN(_u10_N1032 ));
NAND2_X1 _u10_U11740  ( .A1(_u10_req_r_0_ ), .A2(_u10_n5 ), .ZN(_u10_n22957 ) );
NAND2_X1 _u10_U11739  ( .A1(ch0_csr[5]), .A2(_u10_n22957 ), .ZN(_u10_n22956 ) );
NAND2_X1 _u10_U11738  ( .A1(ch0_csr[0]), .A2(_u10_n22956 ), .ZN(_u10_n13702 ) );
NOR3_X1 _u10_U11737  ( .A1(ch_sel[2]), .A2(ch_sel[3]), .A3(ch_sel[4]), .ZN(_u10_n22944 ) );
NOR2_X1 _u10_U11736  ( .A1(ch_sel[1]), .A2(ch_sel[0]), .ZN(_u10_n22909 ) );
NAND2_X1 _u10_U11735  ( .A1(_u10_n22944 ), .A2(_u10_n22909 ), .ZN(_u10_n16357 ) );
NOR2_X1 _u10_U11734  ( .A1(_u10_n13702 ), .A2(_u10_n16357 ), .ZN(_u10_n11552 ) );
AND2_X1 _u10_U11733  ( .A1(next_ch), .A2(_u10_n11552 ), .ZN(_u10_N1033 ) );
INV_X1 _u10_U11732  ( .A(_u10_n16357 ), .ZN(_u10_n12404 ) );
AND3_X1 _u10_U11731  ( .A1(ch0_csr[5]), .A2(_u10_n12000 ), .A3(de_ack), .ZN(_u10_N1034 ) );
AND2_X1 _u10_U11730  ( .A1(dma_req_i[0]), .A2(_u10_n5 ), .ZN(_u10_N967 ) );
AND2_X1 _u10_U11729  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N971 ) );
AND2_X1 _u10_U11728  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N972 ) );
AND2_X1 _u10_U11727  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N973 ) );
AND2_X1 _u10_U11726  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N974 ) );
AND2_X1 _u10_U11725  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N975 ) );
AND2_X1 _u10_U11724  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N976 ) );
AND2_X1 _u10_U11723  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N977 ) );
AND2_X1 _u10_U11722  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N978 ) );
AND2_X1 _u10_U11721  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N979 ) );
AND2_X1 _u10_U11720  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N980 ) );
AND2_X1 _u10_U11719  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N981 ) );
AND2_X1 _u10_U11718  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N982 ) );
AND2_X1 _u10_U11717  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N983 ) );
AND2_X1 _u10_U11716  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N984 ) );
AND2_X1 _u10_U11715  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N985 ) );
AND2_X1 _u10_U11714  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N986 ) );
AND2_X1 _u10_U11713  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N987 ) );
AND2_X1 _u10_U11712  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N988 ) );
AND2_X1 _u10_U11711  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N989 ) );
AND2_X1 _u10_U11710  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N990 ) );
AND2_X1 _u10_U11709  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N991 ) );
AND2_X1 _u10_U11708  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N992 ) );
AND2_X1 _u10_U11707  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N993 ) );
AND2_X1 _u10_U11706  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N994 ) );
AND2_X1 _u10_U11705  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N995 ) );
AND2_X1 _u10_U11704  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N996 ) );
AND2_X1 _u10_U11703  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N997 ) );
AND2_X1 _u10_U11702  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N998 ) );
AND2_X1 _u10_U11701  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_N999 ) );
INV_X1 _u10_U11700  ( .A(ch_sel[3]), .ZN(_u10_n22925 ) );
NOR3_X1 _u10_U11699  ( .A1(ch_sel[4]), .A2(ch_sel[2]), .A3(_u10_n22925 ),.ZN(_u10_n22938 ) );
INV_X1 _u10_U11698  ( .A(ch_sel[0]), .ZN(_u10_n22947 ) );
NOR2_X1 _u10_U11697  ( .A1(_u10_n22947 ), .A2(ch_sel[1]), .ZN(_u10_n22918 ));
NAND2_X1 _u10_U11696  ( .A1(_u10_n22938 ), .A2(_u10_n22918 ), .ZN(_u10_n16366 ) );
INV_X1 _u10_U11695  ( .A(_u10_n16366 ), .ZN(_u10_n12430 ) );
NAND2_X1 _u10_U11694  ( .A1(1'b0), .A2(_u10_n12353 ), .ZN(_u10_n22952 ) );
INV_X1 _u10_U11693  ( .A(ch_sel[1]), .ZN(_u10_n22946 ) );
NOR2_X1 _u10_U11692  ( .A1(_u10_n22946 ), .A2(ch_sel[0]), .ZN(_u10_n22917 ));
NAND2_X1 _u10_U11691  ( .A1(_u10_n22938 ), .A2(_u10_n22917 ), .ZN(_u10_n16367 ) );
INV_X1 _u10_U11690  ( .A(_u10_n16367 ), .ZN(_u10_n12429 ) );
NAND2_X1 _u10_U11689  ( .A1(1'b0), .A2(_u10_n12328 ), .ZN(_u10_n22953 ) );
INV_X1 _u10_U11688  ( .A(ch_sel[2]), .ZN(_u10_n22919 ) );
NOR3_X1 _u10_U11687  ( .A1(ch_sel[4]), .A2(ch_sel[3]), .A3(_u10_n22919 ),.ZN(_u10_n22939 ) );
NAND2_X1 _u10_U11686  ( .A1(_u10_n22939 ), .A2(_u10_n22918 ), .ZN(_u10_n16368 ) );
INV_X1 _u10_U11685  ( .A(_u10_n16368 ), .ZN(_u10_n12428 ) );
NAND2_X1 _u10_U11684  ( .A1(1'b0), .A2(_u10_n12303 ), .ZN(_u10_n22954 ) );
NAND2_X1 _u10_U11683  ( .A1(_u10_n22939 ), .A2(_u10_n22917 ), .ZN(_u10_n16369 ) );
INV_X1 _u10_U11682  ( .A(_u10_n16369 ), .ZN(_u10_n12427 ) );
NAND2_X1 _u10_U11681  ( .A1(1'b0), .A2(_u10_n12279 ), .ZN(_u10_n22955 ) );
NAND4_X1 _u10_U11680  ( .A1(_u10_n22952 ), .A2(_u10_n22953 ), .A3(_u10_n22954 ), .A4(_u10_n22955 ), .ZN(_u10_n22931 ) );
NOR3_X1 _u10_U11679  ( .A1(ch_sel[4]), .A2(_u10_n22925 ), .A3(_u10_n22919 ),.ZN(_u10_n22945 ) );
NAND2_X1 _u10_U11678  ( .A1(_u10_n22945 ), .A2(_u10_n22918 ), .ZN(_u10_n16374 ) );
INV_X1 _u10_U11677  ( .A(_u10_n16374 ), .ZN(_u10_n12422 ) );
NAND2_X1 _u10_U11676  ( .A1(1'b0), .A2(_u10_n12257 ), .ZN(_u10_n22948 ) );
NAND2_X1 _u10_U11675  ( .A1(_u10_n22945 ), .A2(_u10_n22917 ), .ZN(_u10_n16375 ) );
INV_X1 _u10_U11674  ( .A(_u10_n16375 ), .ZN(_u10_n12421 ) );
NAND2_X1 _u10_U11673  ( .A1(1'b0), .A2(_u10_n12233 ), .ZN(_u10_n22949 ) );
NAND2_X1 _u10_U11672  ( .A1(_u10_n22944 ), .A2(_u10_n22918 ), .ZN(_u10_n16376 ) );
INV_X1 _u10_U11671  ( .A(_u10_n16376 ), .ZN(_u10_n12420 ) );
NAND2_X1 _u10_U11670  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n22950 ) );
NAND2_X1 _u10_U11669  ( .A1(_u10_n22944 ), .A2(_u10_n22917 ), .ZN(_u10_n16377 ) );
INV_X1 _u10_U11668  ( .A(_u10_n16377 ), .ZN(_u10_n12419 ) );
NAND2_X1 _u10_U11667  ( .A1(1'b0), .A2(_u10_n12185 ), .ZN(_u10_n22951 ) );
NAND4_X1 _u10_U11666  ( .A1(_u10_n22948 ), .A2(_u10_n22949 ), .A3(_u10_n22950 ), .A4(_u10_n22951 ), .ZN(_u10_n22932 ) );
NOR2_X1 _u10_U11665  ( .A1(_u10_n22946 ), .A2(_u10_n22947 ), .ZN(_u10_n22911 ) );
AND2_X1 _u10_U11664  ( .A1(_u10_n22938 ), .A2(_u10_n22911 ), .ZN(_u10_n12414 ) );
NAND2_X1 _u10_U11663  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n22940 ) );
AND2_X1 _u10_U11662  ( .A1(_u10_n22945 ), .A2(_u10_n22909 ), .ZN(_u10_n12413 ) );
NAND2_X1 _u10_U11661  ( .A1(1'b0), .A2(_u10_n12136 ), .ZN(_u10_n22941 ) );
AND2_X1 _u10_U11660  ( .A1(_u10_n22944 ), .A2(_u10_n22911 ), .ZN(_u10_n12412 ) );
NAND2_X1 _u10_U11659  ( .A1(1'b0), .A2(_u10_n12112 ), .ZN(_u10_n22942 ) );
AND2_X1 _u10_U11658  ( .A1(_u10_n22939 ), .A2(_u10_n22909 ), .ZN(_u10_n12411 ) );
NAND2_X1 _u10_U11657  ( .A1(1'b0), .A2(_u10_n12088 ), .ZN(_u10_n22943 ) );
NAND4_X1 _u10_U11656  ( .A1(_u10_n22940 ), .A2(_u10_n22941 ), .A3(_u10_n22942 ), .A4(_u10_n22943 ), .ZN(_u10_n22933 ) );
NAND2_X1 _u10_U11655  ( .A1(_u10_n22939 ), .A2(_u10_n22911 ), .ZN(_u10_n16355 ) );
INV_X1 _u10_U11654  ( .A(_u10_n16355 ), .ZN(_u10_n12406 ) );
NAND2_X1 _u10_U11653  ( .A1(1'b0), .A2(_u10_n12065 ), .ZN(_u10_n22935 ) );
NAND2_X1 _u10_U11652  ( .A1(_u10_n22938 ), .A2(_u10_n22909 ), .ZN(_u10_n16356 ) );
INV_X1 _u10_U11651  ( .A(_u10_n16356 ), .ZN(_u10_n12405 ) );
NAND2_X1 _u10_U11650  ( .A1(1'b0), .A2(_u10_n12041 ), .ZN(_u10_n22936 ) );
NAND2_X1 _u10_U11649  ( .A1(1'b0), .A2(_u10_n12000 ), .ZN(_u10_n22937 ) );
NAND3_X1 _u10_U11648  ( .A1(_u10_n22935 ), .A2(_u10_n22936 ), .A3(_u10_n22937 ), .ZN(_u10_n22934 ) );
NOR4_X1 _u10_U11647  ( .A1(_u10_n22931 ), .A2(_u10_n22932 ), .A3(_u10_n22933 ), .A4(_u10_n22934 ), .ZN(_u10_n22898 ) );
NAND2_X1 _u10_U11646  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n22927 ) );
AND3_X1 _u10_U11645  ( .A1(_u10_n22919 ), .A2(_u10_n22925 ), .A3(ch_sel[4]),.ZN(_u10_n22926 ) );
AND2_X1 _u10_U11644  ( .A1(_u10_n22909 ), .A2(_u10_n22926 ), .ZN(_u10_n12395 ) );
NAND2_X1 _u10_U11643  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n22928 ) );
AND2_X1 _u10_U11642  ( .A1(_u10_n22918 ), .A2(_u10_n22926 ), .ZN(_u10_n12394 ) );
NAND2_X1 _u10_U11641  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n22929 ) );
AND2_X1 _u10_U11640  ( .A1(_u10_n22917 ), .A2(_u10_n22926 ), .ZN(_u10_n12393 ) );
NAND2_X1 _u10_U11639  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n22930 ) );
NAND4_X1 _u10_U11638  ( .A1(_u10_n22927 ), .A2(_u10_n22928 ), .A3(_u10_n22929 ), .A4(_u10_n22930 ), .ZN(_u10_n22900 ) );
AND2_X1 _u10_U11637  ( .A1(_u10_n22911 ), .A2(_u10_n22926 ), .ZN(_u10_n12388 ) );
NAND2_X1 _u10_U11636  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n22920 ) );
AND2_X1 _u10_U11635  ( .A1(_u10_n22924 ), .A2(_u10_n22909 ), .ZN(_u10_n12387 ) );
NAND2_X1 _u10_U11634  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n22921 ) );
AND2_X1 _u10_U11633  ( .A1(_u10_n22924 ), .A2(_u10_n22918 ), .ZN(_u10_n12386 ) );
NAND2_X1 _u10_U11632  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n22922 ) );
AND2_X1 _u10_U11631  ( .A1(_u10_n22924 ), .A2(_u10_n22917 ), .ZN(_u10_n12385 ) );
NAND2_X1 _u10_U11630  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n22923 ) );
NAND4_X1 _u10_U11629  ( .A1(_u10_n22920 ), .A2(_u10_n22921 ), .A3(_u10_n22922 ), .A4(_u10_n22923 ), .ZN(_u10_n22901 ) );
NAND2_X1 _u10_U11628  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n22912 ) );
AND2_X1 _u10_U11627  ( .A1(ch_sel[3]), .A2(ch_sel[4]), .ZN(_u10_n22910 ) );
AND2_X1 _u10_U11626  ( .A1(_u10_n22910 ), .A2(_u10_n22919 ), .ZN(_u10_n22916 ) );
AND2_X1 _u10_U11625  ( .A1(_u10_n22916 ), .A2(_u10_n22909 ), .ZN(_u10_n12379 ) );
NAND2_X1 _u10_U11624  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n22913 ) );
AND2_X1 _u10_U11623  ( .A1(_u10_n22916 ), .A2(_u10_n22918 ), .ZN(_u10_n12378 ) );
NAND2_X1 _u10_U11622  ( .A1(1'b0), .A2(_u10_n11758 ), .ZN(_u10_n22914 ) );
AND2_X1 _u10_U11621  ( .A1(_u10_n22916 ), .A2(_u10_n22917 ), .ZN(_u10_n12377 ) );
NAND2_X1 _u10_U11620  ( .A1(1'b0), .A2(_u10_n11733 ), .ZN(_u10_n22915 ) );
NAND4_X1 _u10_U11619  ( .A1(_u10_n22912 ), .A2(_u10_n22913 ), .A3(_u10_n22914 ), .A4(_u10_n22915 ), .ZN(_u10_n22902 ) );
AND2_X1 _u10_U11618  ( .A1(_u10_n22910 ), .A2(_u10_n22911 ), .ZN(_u10_n12372 ) );
NAND2_X1 _u10_U11617  ( .A1(1'b0), .A2(_u10_n11710 ), .ZN(_u10_n22904 ) );
AND2_X1 _u10_U11616  ( .A1(_u10_n22910 ), .A2(ch_sel[2]), .ZN(_u10_n22908 ));
AND2_X1 _u10_U11615  ( .A1(_u10_n22908 ), .A2(_u10_n22909 ), .ZN(_u10_n12371 ) );
NAND2_X1 _u10_U11614  ( .A1(1'b0), .A2(_u10_n11685 ), .ZN(_u10_n22905 ) );
AND2_X1 _u10_U11613  ( .A1(_u10_n22908 ), .A2(ch_sel[0]), .ZN(_u10_n12370 ));
NAND2_X1 _u10_U11612  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n22906 ) );
AND2_X1 _u10_U11611  ( .A1(_u10_n22908 ), .A2(ch_sel[1]), .ZN(_u10_n12369 ));
NAND2_X1 _u10_U11610  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n22907 ) );
NAND4_X1 _u10_U11609  ( .A1(_u10_n22904 ), .A2(_u10_n22905 ), .A3(_u10_n22906 ), .A4(_u10_n22907 ), .ZN(_u10_n22903 ) );
NOR4_X1 _u10_U11608  ( .A1(_u10_n22900 ), .A2(_u10_n22901 ), .A3(_u10_n22902 ), .A4(_u10_n22903 ), .ZN(_u10_n22899 ) );
NAND2_X1 _u10_U11607  ( .A1(_u10_n22898 ), .A2(_u10_n22899 ), .ZN(adr0[0]));
NAND2_X1 _u10_U11606  ( .A1(1'b0), .A2(_u10_n12352 ), .ZN(_u10_n22894 ) );
NAND2_X1 _u10_U11605  ( .A1(1'b0), .A2(_u10_n12330 ), .ZN(_u10_n22895 ) );
NAND2_X1 _u10_U11604  ( .A1(1'b0), .A2(_u10_n12304 ), .ZN(_u10_n22896 ) );
NAND2_X1 _u10_U11603  ( .A1(1'b0), .A2(_u10_n12280 ), .ZN(_u10_n22897 ) );
NAND4_X1 _u10_U11602  ( .A1(_u10_n22894 ), .A2(_u10_n22895 ), .A3(_u10_n22896 ), .A4(_u10_n22897 ), .ZN(_u10_n22879 ) );
NAND2_X1 _u10_U11601  ( .A1(1'b0), .A2(_u10_n12256 ), .ZN(_u10_n22890 ) );
NAND2_X1 _u10_U11600  ( .A1(1'b0), .A2(_u10_n12232 ), .ZN(_u10_n22891 ) );
NAND2_X1 _u10_U11599  ( .A1(1'b0), .A2(_u10_n12206 ), .ZN(_u10_n22892 ) );
NAND2_X1 _u10_U11598  ( .A1(1'b0), .A2(_u10_n12184 ), .ZN(_u10_n22893 ) );
NAND4_X1 _u10_U11597  ( .A1(_u10_n22890 ), .A2(_u10_n22891 ), .A3(_u10_n22892 ), .A4(_u10_n22893 ), .ZN(_u10_n22880 ) );
NAND2_X1 _u10_U11596  ( .A1(1'b0), .A2(_u10_n12160 ), .ZN(_u10_n22886 ) );
NAND2_X1 _u10_U11595  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n22887 ) );
NAND2_X1 _u10_U11594  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n22888 ) );
NAND2_X1 _u10_U11593  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n22889 ) );
NAND4_X1 _u10_U11592  ( .A1(_u10_n22886 ), .A2(_u10_n22887 ), .A3(_u10_n22888 ), .A4(_u10_n22889 ), .ZN(_u10_n22881 ) );
NAND2_X1 _u10_U11591  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n22883 ) );
NAND2_X1 _u10_U11590  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n22884 ) );
NAND2_X1 _u10_U11589  ( .A1(ch0_adr0[10]), .A2(_u10_n12000 ), .ZN(_u10_n22885 ) );
NAND3_X1 _u10_U11588  ( .A1(_u10_n22883 ), .A2(_u10_n22884 ), .A3(_u10_n22885 ), .ZN(_u10_n22882 ) );
NOR4_X1 _u10_U11587  ( .A1(_u10_n22879 ), .A2(_u10_n22880 ), .A3(_u10_n22881 ), .A4(_u10_n22882 ), .ZN(_u10_n22857 ) );
NAND2_X1 _u10_U11586  ( .A1(1'b0), .A2(_u10_n11997 ), .ZN(_u10_n22875 ) );
NAND2_X1 _u10_U11585  ( .A1(1'b0), .A2(_u10_n11971 ), .ZN(_u10_n22876 ) );
NAND2_X1 _u10_U11584  ( .A1(1'b0), .A2(_u10_n11947 ), .ZN(_u10_n22877 ) );
NAND2_X1 _u10_U11583  ( .A1(1'b0), .A2(_u10_n11923 ), .ZN(_u10_n22878 ) );
NAND4_X1 _u10_U11582  ( .A1(_u10_n22875 ), .A2(_u10_n22876 ), .A3(_u10_n22877 ), .A4(_u10_n22878 ), .ZN(_u10_n22859 ) );
NAND2_X1 _u10_U11581  ( .A1(1'b0), .A2(_u10_n11901 ), .ZN(_u10_n22871 ) );
NAND2_X1 _u10_U11580  ( .A1(1'b0), .A2(_u10_n11877 ), .ZN(_u10_n22872 ) );
NAND2_X1 _u10_U11579  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n22873 ) );
NAND2_X1 _u10_U11578  ( .A1(1'b0), .A2(_u10_n11829 ), .ZN(_u10_n22874 ) );
NAND4_X1 _u10_U11577  ( .A1(_u10_n22871 ), .A2(_u10_n22872 ), .A3(_u10_n22873 ), .A4(_u10_n22874 ), .ZN(_u10_n22860 ) );
NAND2_X1 _u10_U11576  ( .A1(1'b0), .A2(_u10_n11805 ), .ZN(_u10_n22867 ) );
NAND2_X1 _u10_U11575  ( .A1(1'b0), .A2(_u10_n11781 ), .ZN(_u10_n22868 ) );
NAND2_X1 _u10_U11574  ( .A1(1'b0), .A2(_u10_n11757 ), .ZN(_u10_n22869 ) );
NAND2_X1 _u10_U11573  ( .A1(1'b0), .A2(_u10_n11733 ), .ZN(_u10_n22870 ) );
NAND4_X1 _u10_U11572  ( .A1(_u10_n22867 ), .A2(_u10_n22868 ), .A3(_u10_n22869 ), .A4(_u10_n22870 ), .ZN(_u10_n22861 ) );
NAND2_X1 _u10_U11571  ( .A1(1'b0), .A2(_u10_n11709 ), .ZN(_u10_n22863 ) );
NAND2_X1 _u10_U11570  ( .A1(1'b0), .A2(_u10_n11685 ), .ZN(_u10_n22864 ) );
NAND2_X1 _u10_U11569  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n22865 ) );
NAND2_X1 _u10_U11568  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n22866 ) );
NAND4_X1 _u10_U11567  ( .A1(_u10_n22863 ), .A2(_u10_n22864 ), .A3(_u10_n22865 ), .A4(_u10_n22866 ), .ZN(_u10_n22862 ) );
NOR4_X1 _u10_U11566  ( .A1(_u10_n22859 ), .A2(_u10_n22860 ), .A3(_u10_n22861 ), .A4(_u10_n22862 ), .ZN(_u10_n22858 ) );
NAND2_X1 _u10_U11565  ( .A1(_u10_n22857 ), .A2(_u10_n22858 ), .ZN(adr0[10]));
NAND2_X1 _u10_U11564  ( .A1(1'b0), .A2(_u10_n12356 ), .ZN(_u10_n22853 ) );
NAND2_X1 _u10_U11563  ( .A1(1'b0), .A2(_u10_n12332 ), .ZN(_u10_n22854 ) );
NAND2_X1 _u10_U11562  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n22855 ) );
NAND2_X1 _u10_U11561  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n22856 ) );
NAND4_X1 _u10_U11560  ( .A1(_u10_n22853 ), .A2(_u10_n22854 ), .A3(_u10_n22855 ), .A4(_u10_n22856 ), .ZN(_u10_n22838 ) );
NAND2_X1 _u10_U11559  ( .A1(1'b0), .A2(_u10_n12260 ), .ZN(_u10_n22849 ) );
NAND2_X1 _u10_U11558  ( .A1(1'b0), .A2(_u10_n12236 ), .ZN(_u10_n22850 ) );
NAND2_X1 _u10_U11557  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n22851 ) );
NAND2_X1 _u10_U11556  ( .A1(1'b0), .A2(_u10_n12188 ), .ZN(_u10_n22852 ) );
NAND4_X1 _u10_U11555  ( .A1(_u10_n22849 ), .A2(_u10_n22850 ), .A3(_u10_n22851 ), .A4(_u10_n22852 ), .ZN(_u10_n22839 ) );
NAND2_X1 _u10_U11554  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n22845 ) );
NAND2_X1 _u10_U11553  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n22846 ) );
NAND2_X1 _u10_U11552  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n22847 ) );
NAND2_X1 _u10_U11551  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n22848 ) );
NAND4_X1 _u10_U11550  ( .A1(_u10_n22845 ), .A2(_u10_n22846 ), .A3(_u10_n22847 ), .A4(_u10_n22848 ), .ZN(_u10_n22840 ) );
NAND2_X1 _u10_U11549  ( .A1(1'b0), .A2(_u10_n12068 ), .ZN(_u10_n22842 ) );
NAND2_X1 _u10_U11548  ( .A1(1'b0), .A2(_u10_n12044 ), .ZN(_u10_n22843 ) );
NAND2_X1 _u10_U11547  ( .A1(ch0_adr0[11]), .A2(_u10_n12000 ), .ZN(_u10_n22844 ) );
NAND3_X1 _u10_U11546  ( .A1(_u10_n22842 ), .A2(_u10_n22843 ), .A3(_u10_n22844 ), .ZN(_u10_n22841 ) );
NOR4_X1 _u10_U11545  ( .A1(_u10_n22838 ), .A2(_u10_n22839 ), .A3(_u10_n22840 ), .A4(_u10_n22841 ), .ZN(_u10_n22816 ) );
NAND2_X1 _u10_U11544  ( .A1(1'b0), .A2(_u10_n11997 ), .ZN(_u10_n22834 ) );
NAND2_X1 _u10_U11543  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n22835 ) );
NAND2_X1 _u10_U11542  ( .A1(1'b0), .A2(_u10_n11948 ), .ZN(_u10_n22836 ) );
NAND2_X1 _u10_U11541  ( .A1(1'b0), .A2(_u10_n11924 ), .ZN(_u10_n22837 ) );
NAND4_X1 _u10_U11540  ( .A1(_u10_n22834 ), .A2(_u10_n22835 ), .A3(_u10_n22836 ), .A4(_u10_n22837 ), .ZN(_u10_n22818 ) );
NAND2_X1 _u10_U11539  ( .A1(1'b0), .A2(_u10_n11901 ), .ZN(_u10_n22830 ) );
NAND2_X1 _u10_U11538  ( .A1(1'b0), .A2(_u10_n11877 ), .ZN(_u10_n22831 ) );
NAND2_X1 _u10_U11537  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n22832 ) );
NAND2_X1 _u10_U11536  ( .A1(1'b0), .A2(_u10_n11829 ), .ZN(_u10_n22833 ) );
NAND4_X1 _u10_U11535  ( .A1(_u10_n22830 ), .A2(_u10_n22831 ), .A3(_u10_n22832 ), .A4(_u10_n22833 ), .ZN(_u10_n22819 ) );
NAND2_X1 _u10_U11534  ( .A1(1'b0), .A2(_u10_n11805 ), .ZN(_u10_n22826 ) );
NAND2_X1 _u10_U11533  ( .A1(1'b0), .A2(_u10_n11781 ), .ZN(_u10_n22827 ) );
NAND2_X1 _u10_U11532  ( .A1(1'b0), .A2(_u10_n11757 ), .ZN(_u10_n22828 ) );
NAND2_X1 _u10_U11531  ( .A1(1'b0), .A2(_u10_n11733 ), .ZN(_u10_n22829 ) );
NAND4_X1 _u10_U11530  ( .A1(_u10_n22826 ), .A2(_u10_n22827 ), .A3(_u10_n22828 ), .A4(_u10_n22829 ), .ZN(_u10_n22820 ) );
NAND2_X1 _u10_U11529  ( .A1(1'b0), .A2(_u10_n11709 ), .ZN(_u10_n22822 ) );
NAND2_X1 _u10_U11528  ( .A1(1'b0), .A2(_u10_n11685 ), .ZN(_u10_n22823 ) );
NAND2_X1 _u10_U11527  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n22824 ) );
NAND2_X1 _u10_U11526  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n22825 ) );
NAND4_X1 _u10_U11525  ( .A1(_u10_n22822 ), .A2(_u10_n22823 ), .A3(_u10_n22824 ), .A4(_u10_n22825 ), .ZN(_u10_n22821 ) );
NOR4_X1 _u10_U11524  ( .A1(_u10_n22818 ), .A2(_u10_n22819 ), .A3(_u10_n22820 ), .A4(_u10_n22821 ), .ZN(_u10_n22817 ) );
NAND2_X1 _u10_U11523  ( .A1(_u10_n22816 ), .A2(_u10_n22817 ), .ZN(adr0[11]));
NAND2_X1 _u10_U11522  ( .A1(1'b0), .A2(_u10_n12354 ), .ZN(_u10_n22812 ) );
NAND2_X1 _u10_U11521  ( .A1(1'b0), .A2(_u10_n12331 ), .ZN(_u10_n22813 ) );
NAND2_X1 _u10_U11520  ( .A1(1'b0), .A2(_u10_n12307 ), .ZN(_u10_n22814 ) );
NAND2_X1 _u10_U11519  ( .A1(1'b0), .A2(_u10_n12283 ), .ZN(_u10_n22815 ) );
NAND4_X1 _u10_U11518  ( .A1(_u10_n22812 ), .A2(_u10_n22813 ), .A3(_u10_n22814 ), .A4(_u10_n22815 ), .ZN(_u10_n22797 ) );
NAND2_X1 _u10_U11517  ( .A1(1'b0), .A2(_u10_n12258 ), .ZN(_u10_n22808 ) );
NAND2_X1 _u10_U11516  ( .A1(1'b0), .A2(_u10_n12234 ), .ZN(_u10_n22809 ) );
NAND2_X1 _u10_U11515  ( .A1(1'b0), .A2(_u10_n12209 ), .ZN(_u10_n22810 ) );
NAND2_X1 _u10_U11514  ( .A1(1'b0), .A2(_u10_n12186 ), .ZN(_u10_n22811 ) );
NAND4_X1 _u10_U11513  ( .A1(_u10_n22808 ), .A2(_u10_n22809 ), .A3(_u10_n22810 ), .A4(_u10_n22811 ), .ZN(_u10_n22798 ) );
NAND2_X1 _u10_U11512  ( .A1(1'b0), .A2(_u10_n12161 ), .ZN(_u10_n22804 ) );
NAND2_X1 _u10_U11511  ( .A1(1'b0), .A2(_u10_n12137 ), .ZN(_u10_n22805 ) );
NAND2_X1 _u10_U11510  ( .A1(1'b0), .A2(_u10_n12113 ), .ZN(_u10_n22806 ) );
NAND2_X1 _u10_U11509  ( .A1(1'b0), .A2(_u10_n12089 ), .ZN(_u10_n22807 ) );
NAND4_X1 _u10_U11508  ( .A1(_u10_n22804 ), .A2(_u10_n22805 ), .A3(_u10_n22806 ), .A4(_u10_n22807 ), .ZN(_u10_n22799 ) );
NAND2_X1 _u10_U11507  ( .A1(1'b0), .A2(_u10_n12065 ), .ZN(_u10_n22801 ) );
NAND2_X1 _u10_U11506  ( .A1(1'b0), .A2(_u10_n12041 ), .ZN(_u10_n22802 ) );
NAND2_X1 _u10_U11505  ( .A1(ch0_adr0[12]), .A2(_u10_n12000 ), .ZN(_u10_n22803 ) );
NAND3_X1 _u10_U11504  ( .A1(_u10_n22801 ), .A2(_u10_n22802 ), .A3(_u10_n22803 ), .ZN(_u10_n22800 ) );
NOR4_X1 _u10_U11503  ( .A1(_u10_n22797 ), .A2(_u10_n22798 ), .A3(_u10_n22799 ), .A4(_u10_n22800 ), .ZN(_u10_n22775 ) );
NAND2_X1 _u10_U11502  ( .A1(1'b0), .A2(_u10_n11998 ), .ZN(_u10_n22793 ) );
NAND2_X1 _u10_U11501  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n22794 ) );
NAND2_X1 _u10_U11500  ( .A1(1'b0), .A2(_u10_n11951 ), .ZN(_u10_n22795 ) );
NAND2_X1 _u10_U11499  ( .A1(1'b0), .A2(_u10_n11927 ), .ZN(_u10_n22796 ) );
NAND4_X1 _u10_U11498  ( .A1(_u10_n22793 ), .A2(_u10_n22794 ), .A3(_u10_n22795 ), .A4(_u10_n22796 ), .ZN(_u10_n22777 ) );
NAND2_X1 _u10_U11497  ( .A1(1'b0), .A2(_u10_n11902 ), .ZN(_u10_n22789 ) );
NAND2_X1 _u10_U11496  ( .A1(1'b0), .A2(_u10_n11878 ), .ZN(_u10_n22790 ) );
NAND2_X1 _u10_U11495  ( .A1(1'b0), .A2(_u10_n11854 ), .ZN(_u10_n22791 ) );
NAND2_X1 _u10_U11494  ( .A1(1'b0), .A2(_u10_n11830 ), .ZN(_u10_n22792 ) );
NAND4_X1 _u10_U11493  ( .A1(_u10_n22789 ), .A2(_u10_n22790 ), .A3(_u10_n22791 ), .A4(_u10_n22792 ), .ZN(_u10_n22778 ) );
NAND2_X1 _u10_U11492  ( .A1(1'b0), .A2(_u10_n11806 ), .ZN(_u10_n22785 ) );
NAND2_X1 _u10_U11491  ( .A1(1'b0), .A2(_u10_n11782 ), .ZN(_u10_n22786 ) );
NAND2_X1 _u10_U11490  ( .A1(1'b0), .A2(_u10_n11759 ), .ZN(_u10_n22787 ) );
NAND2_X1 _u10_U11489  ( .A1(1'b0), .A2(_u10_n11735 ), .ZN(_u10_n22788 ) );
NAND4_X1 _u10_U11488  ( .A1(_u10_n22785 ), .A2(_u10_n22786 ), .A3(_u10_n22787 ), .A4(_u10_n22788 ), .ZN(_u10_n22779 ) );
NAND2_X1 _u10_U11487  ( .A1(1'b0), .A2(_u10_n11711 ), .ZN(_u10_n22781 ) );
NAND2_X1 _u10_U11486  ( .A1(1'b0), .A2(_u10_n11687 ), .ZN(_u10_n22782 ) );
NAND2_X1 _u10_U11485  ( .A1(1'b0), .A2(_u10_n11662 ), .ZN(_u10_n22783 ) );
NAND2_X1 _u10_U11484  ( .A1(1'b0), .A2(_u10_n11638 ), .ZN(_u10_n22784 ) );
NAND4_X1 _u10_U11483  ( .A1(_u10_n22781 ), .A2(_u10_n22782 ), .A3(_u10_n22783 ), .A4(_u10_n22784 ), .ZN(_u10_n22780 ) );
NOR4_X1 _u10_U11482  ( .A1(_u10_n22777 ), .A2(_u10_n22778 ), .A3(_u10_n22779 ), .A4(_u10_n22780 ), .ZN(_u10_n22776 ) );
NAND2_X1 _u10_U11481  ( .A1(_u10_n22775 ), .A2(_u10_n22776 ), .ZN(adr0[12]));
NAND2_X1 _u10_U11480  ( .A1(1'b0), .A2(_u10_n12355 ), .ZN(_u10_n22771 ) );
NAND2_X1 _u10_U11479  ( .A1(1'b0), .A2(_u10_n12330 ), .ZN(_u10_n22772 ) );
NAND2_X1 _u10_U11478  ( .A1(1'b0), .A2(_u10_n12306 ), .ZN(_u10_n22773 ) );
NAND2_X1 _u10_U11477  ( .A1(1'b0), .A2(_u10_n12282 ), .ZN(_u10_n22774 ) );
NAND4_X1 _u10_U11476  ( .A1(_u10_n22771 ), .A2(_u10_n22772 ), .A3(_u10_n22773 ), .A4(_u10_n22774 ), .ZN(_u10_n22756 ) );
NAND2_X1 _u10_U11475  ( .A1(1'b0), .A2(_u10_n12259 ), .ZN(_u10_n22767 ) );
NAND2_X1 _u10_U11474  ( .A1(1'b0), .A2(_u10_n12235 ), .ZN(_u10_n22768 ) );
NAND2_X1 _u10_U11473  ( .A1(1'b0), .A2(_u10_n12211 ), .ZN(_u10_n22769 ) );
NAND2_X1 _u10_U11472  ( .A1(1'b0), .A2(_u10_n12187 ), .ZN(_u10_n22770 ) );
NAND4_X1 _u10_U11471  ( .A1(_u10_n22767 ), .A2(_u10_n22768 ), .A3(_u10_n22769 ), .A4(_u10_n22770 ), .ZN(_u10_n22757 ) );
NAND2_X1 _u10_U11470  ( .A1(1'b0), .A2(_u10_n12163 ), .ZN(_u10_n22763 ) );
NAND2_X1 _u10_U11469  ( .A1(1'b0), .A2(_u10_n12139 ), .ZN(_u10_n22764 ) );
NAND2_X1 _u10_U11468  ( .A1(1'b0), .A2(_u10_n12115 ), .ZN(_u10_n22765 ) );
NAND2_X1 _u10_U11467  ( .A1(1'b0), .A2(_u10_n12091 ), .ZN(_u10_n22766 ) );
NAND4_X1 _u10_U11466  ( .A1(_u10_n22763 ), .A2(_u10_n22764 ), .A3(_u10_n22765 ), .A4(_u10_n22766 ), .ZN(_u10_n22758 ) );
NAND2_X1 _u10_U11465  ( .A1(1'b0), .A2(_u10_n12067 ), .ZN(_u10_n22760 ) );
NAND2_X1 _u10_U11464  ( .A1(1'b0), .A2(_u10_n12043 ), .ZN(_u10_n22761 ) );
NAND2_X1 _u10_U11463  ( .A1(ch0_adr0[13]), .A2(_u10_n12000 ), .ZN(_u10_n22762 ) );
NAND3_X1 _u10_U11462  ( .A1(_u10_n22760 ), .A2(_u10_n22761 ), .A3(_u10_n22762 ), .ZN(_u10_n22759 ) );
NOR4_X1 _u10_U11461  ( .A1(_u10_n22756 ), .A2(_u10_n22757 ), .A3(_u10_n22758 ), .A4(_u10_n22759 ), .ZN(_u10_n22734 ) );
NAND2_X1 _u10_U11460  ( .A1(1'b0), .A2(_u10_n11998 ), .ZN(_u10_n22752 ) );
NAND2_X1 _u10_U11459  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n22753 ) );
NAND2_X1 _u10_U11458  ( .A1(1'b0), .A2(_u10_n12394 ), .ZN(_u10_n22754 ) );
NAND2_X1 _u10_U11457  ( .A1(1'b0), .A2(_u10_n12393 ), .ZN(_u10_n22755 ) );
NAND4_X1 _u10_U11456  ( .A1(_u10_n22752 ), .A2(_u10_n22753 ), .A3(_u10_n22754 ), .A4(_u10_n22755 ), .ZN(_u10_n22736 ) );
NAND2_X1 _u10_U11455  ( .A1(1'b0), .A2(_u10_n11902 ), .ZN(_u10_n22748 ) );
NAND2_X1 _u10_U11454  ( .A1(1'b0), .A2(_u10_n11878 ), .ZN(_u10_n22749 ) );
NAND2_X1 _u10_U11453  ( .A1(1'b0), .A2(_u10_n11854 ), .ZN(_u10_n22750 ) );
NAND2_X1 _u10_U11452  ( .A1(1'b0), .A2(_u10_n11830 ), .ZN(_u10_n22751 ) );
NAND4_X1 _u10_U11451  ( .A1(_u10_n22748 ), .A2(_u10_n22749 ), .A3(_u10_n22750 ), .A4(_u10_n22751 ), .ZN(_u10_n22737 ) );
NAND2_X1 _u10_U11450  ( .A1(1'b0), .A2(_u10_n11806 ), .ZN(_u10_n22744 ) );
NAND2_X1 _u10_U11449  ( .A1(1'b0), .A2(_u10_n11778 ), .ZN(_u10_n22745 ) );
NAND2_X1 _u10_U11448  ( .A1(1'b0), .A2(_u10_n11758 ), .ZN(_u10_n22746 ) );
NAND2_X1 _u10_U11447  ( .A1(1'b0), .A2(_u10_n11734 ), .ZN(_u10_n22747 ) );
NAND4_X1 _u10_U11446  ( .A1(_u10_n22744 ), .A2(_u10_n22745 ), .A3(_u10_n22746 ), .A4(_u10_n22747 ), .ZN(_u10_n22738 ) );
NAND2_X1 _u10_U11445  ( .A1(1'b0), .A2(_u10_n11710 ), .ZN(_u10_n22740 ) );
NAND2_X1 _u10_U11444  ( .A1(1'b0), .A2(_u10_n11686 ), .ZN(_u10_n22741 ) );
NAND2_X1 _u10_U11443  ( .A1(1'b0), .A2(_u10_n11662 ), .ZN(_u10_n22742 ) );
NAND2_X1 _u10_U11442  ( .A1(1'b0), .A2(_u10_n11638 ), .ZN(_u10_n22743 ) );
NAND4_X1 _u10_U11441  ( .A1(_u10_n22740 ), .A2(_u10_n22741 ), .A3(_u10_n22742 ), .A4(_u10_n22743 ), .ZN(_u10_n22739 ) );
NOR4_X1 _u10_U11440  ( .A1(_u10_n22736 ), .A2(_u10_n22737 ), .A3(_u10_n22738 ), .A4(_u10_n22739 ), .ZN(_u10_n22735 ) );
NAND2_X1 _u10_U11439  ( .A1(_u10_n22734 ), .A2(_u10_n22735 ), .ZN(adr0[13]));
NAND2_X1 _u10_U11438  ( .A1(1'b0), .A2(_u10_n12352 ), .ZN(_u10_n22730 ) );
NAND2_X1 _u10_U11437  ( .A1(1'b0), .A2(_u10_n12329 ), .ZN(_u10_n22731 ) );
NAND2_X1 _u10_U11436  ( .A1(1'b0), .A2(_u10_n12305 ), .ZN(_u10_n22732 ) );
NAND2_X1 _u10_U11435  ( .A1(1'b0), .A2(_u10_n12281 ), .ZN(_u10_n22733 ) );
NAND4_X1 _u10_U11434  ( .A1(_u10_n22730 ), .A2(_u10_n22731 ), .A3(_u10_n22732 ), .A4(_u10_n22733 ), .ZN(_u10_n22715 ) );
NAND2_X1 _u10_U11433  ( .A1(1'b0), .A2(_u10_n12256 ), .ZN(_u10_n22726 ) );
NAND2_X1 _u10_U11432  ( .A1(1'b0), .A2(_u10_n12232 ), .ZN(_u10_n22727 ) );
NAND2_X1 _u10_U11431  ( .A1(1'b0), .A2(_u10_n12210 ), .ZN(_u10_n22728 ) );
NAND2_X1 _u10_U11430  ( .A1(1'b0), .A2(_u10_n12184 ), .ZN(_u10_n22729 ) );
NAND4_X1 _u10_U11429  ( .A1(_u10_n22726 ), .A2(_u10_n22727 ), .A3(_u10_n22728 ), .A4(_u10_n22729 ), .ZN(_u10_n22716 ) );
NAND2_X1 _u10_U11428  ( .A1(1'b0), .A2(_u10_n12162 ), .ZN(_u10_n22722 ) );
NAND2_X1 _u10_U11427  ( .A1(1'b0), .A2(_u10_n12138 ), .ZN(_u10_n22723 ) );
NAND2_X1 _u10_U11426  ( .A1(1'b0), .A2(_u10_n12114 ), .ZN(_u10_n22724 ) );
NAND2_X1 _u10_U11425  ( .A1(1'b0), .A2(_u10_n12090 ), .ZN(_u10_n22725 ) );
NAND4_X1 _u10_U11424  ( .A1(_u10_n22722 ), .A2(_u10_n22723 ), .A3(_u10_n22724 ), .A4(_u10_n22725 ), .ZN(_u10_n22717 ) );
NAND2_X1 _u10_U11423  ( .A1(1'b0), .A2(_u10_n12066 ), .ZN(_u10_n22719 ) );
NAND2_X1 _u10_U11422  ( .A1(1'b0), .A2(_u10_n12042 ), .ZN(_u10_n22720 ) );
NAND2_X1 _u10_U11421  ( .A1(ch0_adr0[14]), .A2(_u10_n12000 ), .ZN(_u10_n22721 ) );
NAND3_X1 _u10_U11420  ( .A1(_u10_n22719 ), .A2(_u10_n22720 ), .A3(_u10_n22721 ), .ZN(_u10_n22718 ) );
NOR4_X1 _u10_U11419  ( .A1(_u10_n22715 ), .A2(_u10_n22716 ), .A3(_u10_n22717 ), .A4(_u10_n22718 ), .ZN(_u10_n22693 ) );
NAND2_X1 _u10_U11418  ( .A1(1'b0), .A2(_u10_n11995 ), .ZN(_u10_n22711 ) );
NAND2_X1 _u10_U11417  ( .A1(1'b0), .A2(_u10_n11969 ), .ZN(_u10_n22712 ) );
NAND2_X1 _u10_U11416  ( .A1(1'b0), .A2(_u10_n11948 ), .ZN(_u10_n22713 ) );
NAND2_X1 _u10_U11415  ( .A1(1'b0), .A2(_u10_n11924 ), .ZN(_u10_n22714 ) );
NAND4_X1 _u10_U11414  ( .A1(_u10_n22711 ), .A2(_u10_n22712 ), .A3(_u10_n22713 ), .A4(_u10_n22714 ), .ZN(_u10_n22695 ) );
NAND2_X1 _u10_U11413  ( .A1(1'b0), .A2(_u10_n11899 ), .ZN(_u10_n22707 ) );
NAND2_X1 _u10_U11412  ( .A1(1'b0), .A2(_u10_n11875 ), .ZN(_u10_n22708 ) );
NAND2_X1 _u10_U11411  ( .A1(1'b0), .A2(_u10_n11851 ), .ZN(_u10_n22709 ) );
NAND2_X1 _u10_U11410  ( .A1(1'b0), .A2(_u10_n11827 ), .ZN(_u10_n22710 ) );
NAND4_X1 _u10_U11409  ( .A1(_u10_n22707 ), .A2(_u10_n22708 ), .A3(_u10_n22709 ), .A4(_u10_n22710 ), .ZN(_u10_n22696 ) );
NAND2_X1 _u10_U11408  ( .A1(1'b0), .A2(_u10_n11803 ), .ZN(_u10_n22703 ) );
NAND2_X1 _u10_U11407  ( .A1(1'b0), .A2(_u10_n11779 ), .ZN(_u10_n22704 ) );
NAND2_X1 _u10_U11406  ( .A1(1'b0), .A2(_u10_n11755 ), .ZN(_u10_n22705 ) );
NAND2_X1 _u10_U11405  ( .A1(1'b0), .A2(_u10_n11731 ), .ZN(_u10_n22706 ) );
NAND4_X1 _u10_U11404  ( .A1(_u10_n22703 ), .A2(_u10_n22704 ), .A3(_u10_n22705 ), .A4(_u10_n22706 ), .ZN(_u10_n22697 ) );
NAND2_X1 _u10_U11403  ( .A1(1'b0), .A2(_u10_n11707 ), .ZN(_u10_n22699 ) );
NAND2_X1 _u10_U11402  ( .A1(1'b0), .A2(_u10_n11683 ), .ZN(_u10_n22700 ) );
NAND2_X1 _u10_U11401  ( .A1(1'b0), .A2(_u10_n11659 ), .ZN(_u10_n22701 ) );
NAND2_X1 _u10_U11400  ( .A1(1'b0), .A2(_u10_n11635 ), .ZN(_u10_n22702 ) );
NAND4_X1 _u10_U11399  ( .A1(_u10_n22699 ), .A2(_u10_n22700 ), .A3(_u10_n22701 ), .A4(_u10_n22702 ), .ZN(_u10_n22698 ) );
NOR4_X1 _u10_U11398  ( .A1(_u10_n22695 ), .A2(_u10_n22696 ), .A3(_u10_n22697 ), .A4(_u10_n22698 ), .ZN(_u10_n22694 ) );
NAND2_X1 _u10_U11397  ( .A1(_u10_n22693 ), .A2(_u10_n22694 ), .ZN(adr0[14]));
NAND2_X1 _u10_U11396  ( .A1(1'b0), .A2(_u10_n12353 ), .ZN(_u10_n22689 ) );
NAND2_X1 _u10_U11395  ( .A1(1'b0), .A2(_u10_n12328 ), .ZN(_u10_n22690 ) );
NAND2_X1 _u10_U11394  ( .A1(1'b0), .A2(_u10_n12304 ), .ZN(_u10_n22691 ) );
NAND2_X1 _u10_U11393  ( .A1(1'b0), .A2(_u10_n12280 ), .ZN(_u10_n22692 ) );
NAND4_X1 _u10_U11392  ( .A1(_u10_n22689 ), .A2(_u10_n22690 ), .A3(_u10_n22691 ), .A4(_u10_n22692 ), .ZN(_u10_n22674 ) );
NAND2_X1 _u10_U11391  ( .A1(1'b0), .A2(_u10_n12257 ), .ZN(_u10_n22685 ) );
NAND2_X1 _u10_U11390  ( .A1(1'b0), .A2(_u10_n12233 ), .ZN(_u10_n22686 ) );
NAND2_X1 _u10_U11389  ( .A1(1'b0), .A2(_u10_n12207 ), .ZN(_u10_n22687 ) );
NAND2_X1 _u10_U11388  ( .A1(1'b0), .A2(_u10_n12185 ), .ZN(_u10_n22688 ) );
NAND4_X1 _u10_U11387  ( .A1(_u10_n22685 ), .A2(_u10_n22686 ), .A3(_u10_n22687 ), .A4(_u10_n22688 ), .ZN(_u10_n22675 ) );
NAND2_X1 _u10_U11386  ( .A1(1'b0), .A2(_u10_n12159 ), .ZN(_u10_n22681 ) );
NAND2_X1 _u10_U11385  ( .A1(1'b0), .A2(_u10_n12135 ), .ZN(_u10_n22682 ) );
NAND2_X1 _u10_U11384  ( .A1(1'b0), .A2(_u10_n12111 ), .ZN(_u10_n22683 ) );
NAND2_X1 _u10_U11383  ( .A1(1'b0), .A2(_u10_n12087 ), .ZN(_u10_n22684 ) );
NAND4_X1 _u10_U11382  ( .A1(_u10_n22681 ), .A2(_u10_n22682 ), .A3(_u10_n22683 ), .A4(_u10_n22684 ), .ZN(_u10_n22676 ) );
NAND2_X1 _u10_U11381  ( .A1(1'b0), .A2(_u10_n12063 ), .ZN(_u10_n22678 ) );
NAND2_X1 _u10_U11380  ( .A1(1'b0), .A2(_u10_n12039 ), .ZN(_u10_n22679 ) );
NAND2_X1 _u10_U11379  ( .A1(ch0_adr0[15]), .A2(_u10_n12000 ), .ZN(_u10_n22680 ) );
NAND3_X1 _u10_U11378  ( .A1(_u10_n22678 ), .A2(_u10_n22679 ), .A3(_u10_n22680 ), .ZN(_u10_n22677 ) );
NOR4_X1 _u10_U11377  ( .A1(_u10_n22674 ), .A2(_u10_n22675 ), .A3(_u10_n22676 ), .A4(_u10_n22677 ), .ZN(_u10_n22652 ) );
NAND2_X1 _u10_U11376  ( .A1(1'b0), .A2(_u10_n11998 ), .ZN(_u10_n22670 ) );
NAND2_X1 _u10_U11375  ( .A1(1'b0), .A2(_u10_n11974 ), .ZN(_u10_n22671 ) );
NAND2_X1 _u10_U11374  ( .A1(1'b0), .A2(_u10_n11948 ), .ZN(_u10_n22672 ) );
NAND2_X1 _u10_U11373  ( .A1(1'b0), .A2(_u10_n11924 ), .ZN(_u10_n22673 ) );
NAND4_X1 _u10_U11372  ( .A1(_u10_n22670 ), .A2(_u10_n22671 ), .A3(_u10_n22672 ), .A4(_u10_n22673 ), .ZN(_u10_n22654 ) );
NAND2_X1 _u10_U11371  ( .A1(1'b0), .A2(_u10_n12388 ), .ZN(_u10_n22666 ) );
NAND2_X1 _u10_U11370  ( .A1(1'b0), .A2(_u10_n11878 ), .ZN(_u10_n22667 ) );
NAND2_X1 _u10_U11369  ( .A1(1'b0), .A2(_u10_n11850 ), .ZN(_u10_n22668 ) );
NAND2_X1 _u10_U11368  ( .A1(1'b0), .A2(_u10_n12385 ), .ZN(_u10_n22669 ) );
NAND4_X1 _u10_U11367  ( .A1(_u10_n22666 ), .A2(_u10_n22667 ), .A3(_u10_n22668 ), .A4(_u10_n22669 ), .ZN(_u10_n22655 ) );
NAND2_X1 _u10_U11366  ( .A1(1'b0), .A2(_u10_n11806 ), .ZN(_u10_n22662 ) );
NAND2_X1 _u10_U11365  ( .A1(1'b0), .A2(_u10_n11782 ), .ZN(_u10_n22663 ) );
NAND2_X1 _u10_U11364  ( .A1(1'b0), .A2(_u10_n11759 ), .ZN(_u10_n22664 ) );
NAND2_X1 _u10_U11363  ( .A1(1'b0), .A2(_u10_n11735 ), .ZN(_u10_n22665 ) );
NAND4_X1 _u10_U11362  ( .A1(_u10_n22662 ), .A2(_u10_n22663 ), .A3(_u10_n22664 ), .A4(_u10_n22665 ), .ZN(_u10_n22656 ) );
NAND2_X1 _u10_U11361  ( .A1(1'b0), .A2(_u10_n11711 ), .ZN(_u10_n22658 ) );
NAND2_X1 _u10_U11360  ( .A1(1'b0), .A2(_u10_n11687 ), .ZN(_u10_n22659 ) );
NAND2_X1 _u10_U11359  ( .A1(1'b0), .A2(_u10_n11658 ), .ZN(_u10_n22660 ) );
NAND2_X1 _u10_U11358  ( .A1(1'b0), .A2(_u10_n11634 ), .ZN(_u10_n22661 ) );
NAND4_X1 _u10_U11357  ( .A1(_u10_n22658 ), .A2(_u10_n22659 ), .A3(_u10_n22660 ), .A4(_u10_n22661 ), .ZN(_u10_n22657 ) );
NOR4_X1 _u10_U11356  ( .A1(_u10_n22654 ), .A2(_u10_n22655 ), .A3(_u10_n22656 ), .A4(_u10_n22657 ), .ZN(_u10_n22653 ) );
NAND2_X1 _u10_U11355  ( .A1(_u10_n22652 ), .A2(_u10_n22653 ), .ZN(adr0[15]));
NAND2_X1 _u10_U11354  ( .A1(1'b0), .A2(_u10_n12355 ), .ZN(_u10_n22648 ) );
NAND2_X1 _u10_U11353  ( .A1(1'b0), .A2(_u10_n12330 ), .ZN(_u10_n22649 ) );
NAND2_X1 _u10_U11352  ( .A1(1'b0), .A2(_u10_n12304 ), .ZN(_u10_n22650 ) );
NAND2_X1 _u10_U11351  ( .A1(1'b0), .A2(_u10_n12280 ), .ZN(_u10_n22651 ) );
NAND4_X1 _u10_U11350  ( .A1(_u10_n22648 ), .A2(_u10_n22649 ), .A3(_u10_n22650 ), .A4(_u10_n22651 ), .ZN(_u10_n22633 ) );
NAND2_X1 _u10_U11349  ( .A1(1'b0), .A2(_u10_n12259 ), .ZN(_u10_n22644 ) );
NAND2_X1 _u10_U11348  ( .A1(1'b0), .A2(_u10_n12235 ), .ZN(_u10_n22645 ) );
NAND2_X1 _u10_U11347  ( .A1(1'b0), .A2(_u10_n12207 ), .ZN(_u10_n22646 ) );
NAND2_X1 _u10_U11346  ( .A1(1'b0), .A2(_u10_n12187 ), .ZN(_u10_n22647 ) );
NAND4_X1 _u10_U11345  ( .A1(_u10_n22644 ), .A2(_u10_n22645 ), .A3(_u10_n22646 ), .A4(_u10_n22647 ), .ZN(_u10_n22634 ) );
NAND2_X1 _u10_U11344  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n22640 ) );
NAND2_X1 _u10_U11343  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n22641 ) );
NAND2_X1 _u10_U11342  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n22642 ) );
NAND2_X1 _u10_U11341  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n22643 ) );
NAND4_X1 _u10_U11340  ( .A1(_u10_n22640 ), .A2(_u10_n22641 ), .A3(_u10_n22642 ), .A4(_u10_n22643 ), .ZN(_u10_n22635 ) );
NAND2_X1 _u10_U11339  ( .A1(1'b0), .A2(_u10_n12067 ), .ZN(_u10_n22637 ) );
NAND2_X1 _u10_U11338  ( .A1(1'b0), .A2(_u10_n12043 ), .ZN(_u10_n22638 ) );
NAND2_X1 _u10_U11337  ( .A1(ch0_adr0[16]), .A2(_u10_n12000 ), .ZN(_u10_n22639 ) );
NAND3_X1 _u10_U11336  ( .A1(_u10_n22637 ), .A2(_u10_n22638 ), .A3(_u10_n22639 ), .ZN(_u10_n22636 ) );
NOR4_X1 _u10_U11335  ( .A1(_u10_n22633 ), .A2(_u10_n22634 ), .A3(_u10_n22635 ), .A4(_u10_n22636 ), .ZN(_u10_n22611 ) );
NAND2_X1 _u10_U11334  ( .A1(1'b0), .A2(_u10_n11999 ), .ZN(_u10_n22629 ) );
NAND2_X1 _u10_U11333  ( .A1(1'b0), .A2(_u10_n11971 ), .ZN(_u10_n22630 ) );
NAND2_X1 _u10_U11332  ( .A1(1'b0), .A2(_u10_n11950 ), .ZN(_u10_n22631 ) );
NAND2_X1 _u10_U11331  ( .A1(1'b0), .A2(_u10_n11926 ), .ZN(_u10_n22632 ) );
NAND4_X1 _u10_U11330  ( .A1(_u10_n22629 ), .A2(_u10_n22630 ), .A3(_u10_n22631 ), .A4(_u10_n22632 ), .ZN(_u10_n22613 ) );
NAND2_X1 _u10_U11329  ( .A1(1'b0), .A2(_u10_n11903 ), .ZN(_u10_n22625 ) );
NAND2_X1 _u10_U11328  ( .A1(1'b0), .A2(_u10_n11879 ), .ZN(_u10_n22626 ) );
NAND2_X1 _u10_U11327  ( .A1(1'b0), .A2(_u10_n12386 ), .ZN(_u10_n22627 ) );
NAND2_X1 _u10_U11326  ( .A1(1'b0), .A2(_u10_n11831 ), .ZN(_u10_n22628 ) );
NAND4_X1 _u10_U11325  ( .A1(_u10_n22625 ), .A2(_u10_n22626 ), .A3(_u10_n22627 ), .A4(_u10_n22628 ), .ZN(_u10_n22614 ) );
NAND2_X1 _u10_U11324  ( .A1(1'b0), .A2(_u10_n11807 ), .ZN(_u10_n22621 ) );
NAND2_X1 _u10_U11323  ( .A1(1'b0), .A2(_u10_n11783 ), .ZN(_u10_n22622 ) );
NAND2_X1 _u10_U11322  ( .A1(1'b0), .A2(_u10_n11754 ), .ZN(_u10_n22623 ) );
NAND2_X1 _u10_U11321  ( .A1(1'b0), .A2(_u10_n11730 ), .ZN(_u10_n22624 ) );
NAND4_X1 _u10_U11320  ( .A1(_u10_n22621 ), .A2(_u10_n22622 ), .A3(_u10_n22623 ), .A4(_u10_n22624 ), .ZN(_u10_n22615 ) );
NAND2_X1 _u10_U11319  ( .A1(1'b0), .A2(_u10_n11706 ), .ZN(_u10_n22617 ) );
NAND2_X1 _u10_U11318  ( .A1(1'b0), .A2(_u10_n11682 ), .ZN(_u10_n22618 ) );
NAND2_X1 _u10_U11317  ( .A1(1'b0), .A2(_u10_n12370 ), .ZN(_u10_n22619 ) );
NAND2_X1 _u10_U11316  ( .A1(1'b0), .A2(_u10_n12369 ), .ZN(_u10_n22620 ) );
NAND4_X1 _u10_U11315  ( .A1(_u10_n22617 ), .A2(_u10_n22618 ), .A3(_u10_n22619 ), .A4(_u10_n22620 ), .ZN(_u10_n22616 ) );
NOR4_X1 _u10_U11314  ( .A1(_u10_n22613 ), .A2(_u10_n22614 ), .A3(_u10_n22615 ), .A4(_u10_n22616 ), .ZN(_u10_n22612 ) );
NAND2_X1 _u10_U11313  ( .A1(_u10_n22611 ), .A2(_u10_n22612 ), .ZN(adr0[16]));
NAND2_X1 _u10_U11312  ( .A1(1'b0), .A2(_u10_n12355 ), .ZN(_u10_n22607 ) );
NAND2_X1 _u10_U11311  ( .A1(1'b0), .A2(_u10_n12329 ), .ZN(_u10_n22608 ) );
NAND2_X1 _u10_U11310  ( .A1(1'b0), .A2(_u10_n12304 ), .ZN(_u10_n22609 ) );
NAND2_X1 _u10_U11309  ( .A1(1'b0), .A2(_u10_n12280 ), .ZN(_u10_n22610 ) );
NAND4_X1 _u10_U11308  ( .A1(_u10_n22607 ), .A2(_u10_n22608 ), .A3(_u10_n22609 ), .A4(_u10_n22610 ), .ZN(_u10_n22592 ) );
NAND2_X1 _u10_U11307  ( .A1(1'b0), .A2(_u10_n12259 ), .ZN(_u10_n22603 ) );
NAND2_X1 _u10_U11306  ( .A1(1'b0), .A2(_u10_n12235 ), .ZN(_u10_n22604 ) );
NAND2_X1 _u10_U11305  ( .A1(1'b0), .A2(_u10_n12209 ), .ZN(_u10_n22605 ) );
NAND2_X1 _u10_U11304  ( .A1(1'b0), .A2(_u10_n12187 ), .ZN(_u10_n22606 ) );
NAND4_X1 _u10_U11303  ( .A1(_u10_n22603 ), .A2(_u10_n22604 ), .A3(_u10_n22605 ), .A4(_u10_n22606 ), .ZN(_u10_n22593 ) );
NAND2_X1 _u10_U11302  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n22599 ) );
NAND2_X1 _u10_U11301  ( .A1(1'b0), .A2(_u10_n12136 ), .ZN(_u10_n22600 ) );
NAND2_X1 _u10_U11300  ( .A1(1'b0), .A2(_u10_n12112 ), .ZN(_u10_n22601 ) );
NAND2_X1 _u10_U11299  ( .A1(1'b0), .A2(_u10_n12088 ), .ZN(_u10_n22602 ) );
NAND4_X1 _u10_U11298  ( .A1(_u10_n22599 ), .A2(_u10_n22600 ), .A3(_u10_n22601 ), .A4(_u10_n22602 ), .ZN(_u10_n22594 ) );
NAND2_X1 _u10_U11297  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n22596 ) );
NAND2_X1 _u10_U11296  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n22597 ) );
NAND2_X1 _u10_U11295  ( .A1(ch0_adr0[17]), .A2(_u10_n12000 ), .ZN(_u10_n22598 ) );
NAND3_X1 _u10_U11294  ( .A1(_u10_n22596 ), .A2(_u10_n22597 ), .A3(_u10_n22598 ), .ZN(_u10_n22595 ) );
NOR4_X1 _u10_U11293  ( .A1(_u10_n22592 ), .A2(_u10_n22593 ), .A3(_u10_n22594 ), .A4(_u10_n22595 ), .ZN(_u10_n22570 ) );
NAND2_X1 _u10_U11292  ( .A1(1'b0), .A2(_u10_n11994 ), .ZN(_u10_n22588 ) );
NAND2_X1 _u10_U11291  ( .A1(1'b0), .A2(_u10_n11969 ), .ZN(_u10_n22589 ) );
NAND2_X1 _u10_U11290  ( .A1(1'b0), .A2(_u10_n11945 ), .ZN(_u10_n22590 ) );
NAND2_X1 _u10_U11289  ( .A1(1'b0), .A2(_u10_n11921 ), .ZN(_u10_n22591 ) );
NAND4_X1 _u10_U11288  ( .A1(_u10_n22588 ), .A2(_u10_n22589 ), .A3(_u10_n22590 ), .A4(_u10_n22591 ), .ZN(_u10_n22572 ) );
NAND2_X1 _u10_U11287  ( .A1(1'b0), .A2(_u10_n11898 ), .ZN(_u10_n22584 ) );
NAND2_X1 _u10_U11286  ( .A1(1'b0), .A2(_u10_n11874 ), .ZN(_u10_n22585 ) );
NAND2_X1 _u10_U11285  ( .A1(1'b0), .A2(_u10_n11855 ), .ZN(_u10_n22586 ) );
NAND2_X1 _u10_U11284  ( .A1(1'b0), .A2(_u10_n11826 ), .ZN(_u10_n22587 ) );
NAND4_X1 _u10_U11283  ( .A1(_u10_n22584 ), .A2(_u10_n22585 ), .A3(_u10_n22586 ), .A4(_u10_n22587 ), .ZN(_u10_n22573 ) );
NAND2_X1 _u10_U11282  ( .A1(1'b0), .A2(_u10_n11802 ), .ZN(_u10_n22580 ) );
NAND2_X1 _u10_U11281  ( .A1(1'b0), .A2(_u10_n11778 ), .ZN(_u10_n22581 ) );
NAND2_X1 _u10_U11280  ( .A1(1'b0), .A2(_u10_n11757 ), .ZN(_u10_n22582 ) );
NAND2_X1 _u10_U11279  ( .A1(1'b0), .A2(_u10_n11734 ), .ZN(_u10_n22583 ) );
NAND4_X1 _u10_U11278  ( .A1(_u10_n22580 ), .A2(_u10_n22581 ), .A3(_u10_n22582 ), .A4(_u10_n22583 ), .ZN(_u10_n22574 ) );
NAND2_X1 _u10_U11277  ( .A1(1'b0), .A2(_u10_n11709 ), .ZN(_u10_n22576 ) );
NAND2_X1 _u10_U11276  ( .A1(1'b0), .A2(_u10_n11686 ), .ZN(_u10_n22577 ) );
NAND2_X1 _u10_U11275  ( .A1(1'b0), .A2(_u10_n11663 ), .ZN(_u10_n22578 ) );
NAND2_X1 _u10_U11274  ( .A1(1'b0), .A2(_u10_n11639 ), .ZN(_u10_n22579 ) );
NAND4_X1 _u10_U11273  ( .A1(_u10_n22576 ), .A2(_u10_n22577 ), .A3(_u10_n22578 ), .A4(_u10_n22579 ), .ZN(_u10_n22575 ) );
NOR4_X1 _u10_U11272  ( .A1(_u10_n22572 ), .A2(_u10_n22573 ), .A3(_u10_n22574 ), .A4(_u10_n22575 ), .ZN(_u10_n22571 ) );
NAND2_X1 _u10_U11271  ( .A1(_u10_n22570 ), .A2(_u10_n22571 ), .ZN(adr0[17]));
NAND2_X1 _u10_U11270  ( .A1(1'b0), .A2(_u10_n12430 ), .ZN(_u10_n22566 ) );
NAND2_X1 _u10_U11269  ( .A1(1'b0), .A2(_u10_n12429 ), .ZN(_u10_n22567 ) );
NAND2_X1 _u10_U11268  ( .A1(1'b0), .A2(_u10_n12303 ), .ZN(_u10_n22568 ) );
NAND2_X1 _u10_U11267  ( .A1(1'b0), .A2(_u10_n12279 ), .ZN(_u10_n22569 ) );
NAND4_X1 _u10_U11266  ( .A1(_u10_n22566 ), .A2(_u10_n22567 ), .A3(_u10_n22568 ), .A4(_u10_n22569 ), .ZN(_u10_n22551 ) );
NAND2_X1 _u10_U11265  ( .A1(1'b0), .A2(_u10_n12422 ), .ZN(_u10_n22562 ) );
NAND2_X1 _u10_U11264  ( .A1(1'b0), .A2(_u10_n12421 ), .ZN(_u10_n22563 ) );
NAND2_X1 _u10_U11263  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n22564 ) );
NAND2_X1 _u10_U11262  ( .A1(1'b0), .A2(_u10_n12419 ), .ZN(_u10_n22565 ) );
NAND4_X1 _u10_U11261  ( .A1(_u10_n22562 ), .A2(_u10_n22563 ), .A3(_u10_n22564 ), .A4(_u10_n22565 ), .ZN(_u10_n22552 ) );
NAND2_X1 _u10_U11260  ( .A1(1'b0), .A2(_u10_n12160 ), .ZN(_u10_n22558 ) );
NAND2_X1 _u10_U11259  ( .A1(1'b0), .A2(_u10_n12137 ), .ZN(_u10_n22559 ) );
NAND2_X1 _u10_U11258  ( .A1(1'b0), .A2(_u10_n12113 ), .ZN(_u10_n22560 ) );
NAND2_X1 _u10_U11257  ( .A1(1'b0), .A2(_u10_n12089 ), .ZN(_u10_n22561 ) );
NAND4_X1 _u10_U11256  ( .A1(_u10_n22558 ), .A2(_u10_n22559 ), .A3(_u10_n22560 ), .A4(_u10_n22561 ), .ZN(_u10_n22553 ) );
NAND2_X1 _u10_U11255  ( .A1(1'b0), .A2(_u10_n12067 ), .ZN(_u10_n22555 ) );
NAND2_X1 _u10_U11254  ( .A1(1'b0), .A2(_u10_n12043 ), .ZN(_u10_n22556 ) );
NAND2_X1 _u10_U11253  ( .A1(ch0_adr0[18]), .A2(_u10_n12000 ), .ZN(_u10_n22557 ) );
NAND3_X1 _u10_U11252  ( .A1(_u10_n22555 ), .A2(_u10_n22556 ), .A3(_u10_n22557 ), .ZN(_u10_n22554 ) );
NOR4_X1 _u10_U11251  ( .A1(_u10_n22551 ), .A2(_u10_n22552 ), .A3(_u10_n22553 ), .A4(_u10_n22554 ), .ZN(_u10_n22529 ) );
NAND2_X1 _u10_U11250  ( .A1(1'b0), .A2(_u10_n11993 ), .ZN(_u10_n22547 ) );
NAND2_X1 _u10_U11249  ( .A1(1'b0), .A2(_u10_n11973 ), .ZN(_u10_n22548 ) );
NAND2_X1 _u10_U11248  ( .A1(1'b0), .A2(_u10_n11949 ), .ZN(_u10_n22549 ) );
NAND2_X1 _u10_U11247  ( .A1(1'b0), .A2(_u10_n11925 ), .ZN(_u10_n22550 ) );
NAND4_X1 _u10_U11246  ( .A1(_u10_n22547 ), .A2(_u10_n22548 ), .A3(_u10_n22549 ), .A4(_u10_n22550 ), .ZN(_u10_n22531 ) );
NAND2_X1 _u10_U11245  ( .A1(1'b0), .A2(_u10_n11897 ), .ZN(_u10_n22543 ) );
NAND2_X1 _u10_U11244  ( .A1(1'b0), .A2(_u10_n11873 ), .ZN(_u10_n22544 ) );
NAND2_X1 _u10_U11243  ( .A1(1'b0), .A2(_u10_n11849 ), .ZN(_u10_n22545 ) );
NAND2_X1 _u10_U11242  ( .A1(1'b0), .A2(_u10_n11825 ), .ZN(_u10_n22546 ) );
NAND4_X1 _u10_U11241  ( .A1(_u10_n22543 ), .A2(_u10_n22544 ), .A3(_u10_n22545 ), .A4(_u10_n22546 ), .ZN(_u10_n22532 ) );
NAND2_X1 _u10_U11240  ( .A1(1'b0), .A2(_u10_n11801 ), .ZN(_u10_n22539 ) );
NAND2_X1 _u10_U11239  ( .A1(1'b0), .A2(_u10_n11777 ), .ZN(_u10_n22540 ) );
NAND2_X1 _u10_U11238  ( .A1(1'b0), .A2(_u10_n11753 ), .ZN(_u10_n22541 ) );
NAND2_X1 _u10_U11237  ( .A1(1'b0), .A2(_u10_n11729 ), .ZN(_u10_n22542 ) );
NAND4_X1 _u10_U11236  ( .A1(_u10_n22539 ), .A2(_u10_n22540 ), .A3(_u10_n22541 ), .A4(_u10_n22542 ), .ZN(_u10_n22533 ) );
NAND2_X1 _u10_U11235  ( .A1(1'b0), .A2(_u10_n11705 ), .ZN(_u10_n22535 ) );
NAND2_X1 _u10_U11234  ( .A1(1'b0), .A2(_u10_n11681 ), .ZN(_u10_n22536 ) );
NAND2_X1 _u10_U11233  ( .A1(1'b0), .A2(_u10_n11657 ), .ZN(_u10_n22537 ) );
NAND2_X1 _u10_U11232  ( .A1(1'b0), .A2(_u10_n11633 ), .ZN(_u10_n22538 ) );
NAND4_X1 _u10_U11231  ( .A1(_u10_n22535 ), .A2(_u10_n22536 ), .A3(_u10_n22537 ), .A4(_u10_n22538 ), .ZN(_u10_n22534 ) );
NOR4_X1 _u10_U11230  ( .A1(_u10_n22531 ), .A2(_u10_n22532 ), .A3(_u10_n22533 ), .A4(_u10_n22534 ), .ZN(_u10_n22530 ) );
NAND2_X1 _u10_U11229  ( .A1(_u10_n22529 ), .A2(_u10_n22530 ), .ZN(adr0[18]));
NAND2_X1 _u10_U11228  ( .A1(1'b0), .A2(_u10_n12356 ), .ZN(_u10_n22525 ) );
NAND2_X1 _u10_U11227  ( .A1(1'b0), .A2(_u10_n12332 ), .ZN(_u10_n22526 ) );
NAND2_X1 _u10_U11226  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n22527 ) );
NAND2_X1 _u10_U11225  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n22528 ) );
NAND4_X1 _u10_U11224  ( .A1(_u10_n22525 ), .A2(_u10_n22526 ), .A3(_u10_n22527 ), .A4(_u10_n22528 ), .ZN(_u10_n22510 ) );
NAND2_X1 _u10_U11223  ( .A1(1'b0), .A2(_u10_n12260 ), .ZN(_u10_n22521 ) );
NAND2_X1 _u10_U11222  ( .A1(1'b0), .A2(_u10_n12236 ), .ZN(_u10_n22522 ) );
NAND2_X1 _u10_U11221  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n22523 ) );
NAND2_X1 _u10_U11220  ( .A1(1'b0), .A2(_u10_n12188 ), .ZN(_u10_n22524 ) );
NAND4_X1 _u10_U11219  ( .A1(_u10_n22521 ), .A2(_u10_n22522 ), .A3(_u10_n22523 ), .A4(_u10_n22524 ), .ZN(_u10_n22511 ) );
NAND2_X1 _u10_U11218  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n22517 ) );
NAND2_X1 _u10_U11217  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n22518 ) );
NAND2_X1 _u10_U11216  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n22519 ) );
NAND2_X1 _u10_U11215  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n22520 ) );
NAND4_X1 _u10_U11214  ( .A1(_u10_n22517 ), .A2(_u10_n22518 ), .A3(_u10_n22519 ), .A4(_u10_n22520 ), .ZN(_u10_n22512 ) );
NAND2_X1 _u10_U11213  ( .A1(1'b0), .A2(_u10_n12068 ), .ZN(_u10_n22514 ) );
NAND2_X1 _u10_U11212  ( .A1(1'b0), .A2(_u10_n12044 ), .ZN(_u10_n22515 ) );
NAND2_X1 _u10_U11211  ( .A1(ch0_adr0[19]), .A2(_u10_n12000 ), .ZN(_u10_n22516 ) );
NAND3_X1 _u10_U11210  ( .A1(_u10_n22514 ), .A2(_u10_n22515 ), .A3(_u10_n22516 ), .ZN(_u10_n22513 ) );
NOR4_X1 _u10_U11209  ( .A1(_u10_n22510 ), .A2(_u10_n22511 ), .A3(_u10_n22512 ), .A4(_u10_n22513 ), .ZN(_u10_n22488 ) );
NAND2_X1 _u10_U11208  ( .A1(1'b0), .A2(_u10_n11997 ), .ZN(_u10_n22506 ) );
NAND2_X1 _u10_U11207  ( .A1(1'b0), .A2(_u10_n11972 ), .ZN(_u10_n22507 ) );
NAND2_X1 _u10_U11206  ( .A1(1'b0), .A2(_u10_n11948 ), .ZN(_u10_n22508 ) );
NAND2_X1 _u10_U11205  ( .A1(1'b0), .A2(_u10_n11924 ), .ZN(_u10_n22509 ) );
NAND4_X1 _u10_U11204  ( .A1(_u10_n22506 ), .A2(_u10_n22507 ), .A3(_u10_n22508 ), .A4(_u10_n22509 ), .ZN(_u10_n22490 ) );
NAND2_X1 _u10_U11203  ( .A1(1'b0), .A2(_u10_n11901 ), .ZN(_u10_n22502 ) );
NAND2_X1 _u10_U11202  ( .A1(1'b0), .A2(_u10_n11877 ), .ZN(_u10_n22503 ) );
NAND2_X1 _u10_U11201  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n22504 ) );
NAND2_X1 _u10_U11200  ( .A1(1'b0), .A2(_u10_n11829 ), .ZN(_u10_n22505 ) );
NAND4_X1 _u10_U11199  ( .A1(_u10_n22502 ), .A2(_u10_n22503 ), .A3(_u10_n22504 ), .A4(_u10_n22505 ), .ZN(_u10_n22491 ) );
NAND2_X1 _u10_U11198  ( .A1(1'b0), .A2(_u10_n11805 ), .ZN(_u10_n22498 ) );
NAND2_X1 _u10_U11197  ( .A1(1'b0), .A2(_u10_n11781 ), .ZN(_u10_n22499 ) );
NAND2_X1 _u10_U11196  ( .A1(1'b0), .A2(_u10_n11757 ), .ZN(_u10_n22500 ) );
NAND2_X1 _u10_U11195  ( .A1(1'b0), .A2(_u10_n11733 ), .ZN(_u10_n22501 ) );
NAND4_X1 _u10_U11194  ( .A1(_u10_n22498 ), .A2(_u10_n22499 ), .A3(_u10_n22500 ), .A4(_u10_n22501 ), .ZN(_u10_n22492 ) );
NAND2_X1 _u10_U11193  ( .A1(1'b0), .A2(_u10_n11709 ), .ZN(_u10_n22494 ) );
NAND2_X1 _u10_U11192  ( .A1(1'b0), .A2(_u10_n11685 ), .ZN(_u10_n22495 ) );
NAND2_X1 _u10_U11191  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n22496 ) );
NAND2_X1 _u10_U11190  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n22497 ) );
NAND4_X1 _u10_U11189  ( .A1(_u10_n22494 ), .A2(_u10_n22495 ), .A3(_u10_n22496 ), .A4(_u10_n22497 ), .ZN(_u10_n22493 ) );
NOR4_X1 _u10_U11188  ( .A1(_u10_n22490 ), .A2(_u10_n22491 ), .A3(_u10_n22492 ), .A4(_u10_n22493 ), .ZN(_u10_n22489 ) );
NAND2_X1 _u10_U11187  ( .A1(_u10_n22488 ), .A2(_u10_n22489 ), .ZN(adr0[19]));
NAND2_X1 _u10_U11186  ( .A1(1'b0), .A2(_u10_n12430 ), .ZN(_u10_n22484 ) );
NAND2_X1 _u10_U11185  ( .A1(1'b0), .A2(_u10_n12429 ), .ZN(_u10_n22485 ) );
NAND2_X1 _u10_U11184  ( .A1(1'b0), .A2(_u10_n12307 ), .ZN(_u10_n22486 ) );
NAND2_X1 _u10_U11183  ( .A1(1'b0), .A2(_u10_n12283 ), .ZN(_u10_n22487 ) );
NAND4_X1 _u10_U11182  ( .A1(_u10_n22484 ), .A2(_u10_n22485 ), .A3(_u10_n22486 ), .A4(_u10_n22487 ), .ZN(_u10_n22469 ) );
NAND2_X1 _u10_U11181  ( .A1(1'b0), .A2(_u10_n12422 ), .ZN(_u10_n22480 ) );
NAND2_X1 _u10_U11180  ( .A1(1'b0), .A2(_u10_n12421 ), .ZN(_u10_n22481 ) );
NAND2_X1 _u10_U11179  ( .A1(1'b0), .A2(_u10_n12211 ), .ZN(_u10_n22482 ) );
NAND2_X1 _u10_U11178  ( .A1(1'b0), .A2(_u10_n12419 ), .ZN(_u10_n22483 ) );
NAND4_X1 _u10_U11177  ( .A1(_u10_n22480 ), .A2(_u10_n22481 ), .A3(_u10_n22482 ), .A4(_u10_n22483 ), .ZN(_u10_n22470 ) );
NAND2_X1 _u10_U11176  ( .A1(1'b0), .A2(_u10_n12162 ), .ZN(_u10_n22476 ) );
NAND2_X1 _u10_U11175  ( .A1(1'b0), .A2(_u10_n12137 ), .ZN(_u10_n22477 ) );
NAND2_X1 _u10_U11174  ( .A1(1'b0), .A2(_u10_n12113 ), .ZN(_u10_n22478 ) );
NAND2_X1 _u10_U11173  ( .A1(1'b0), .A2(_u10_n12089 ), .ZN(_u10_n22479 ) );
NAND4_X1 _u10_U11172  ( .A1(_u10_n22476 ), .A2(_u10_n22477 ), .A3(_u10_n22478 ), .A4(_u10_n22479 ), .ZN(_u10_n22471 ) );
NAND2_X1 _u10_U11171  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n22473 ) );
NAND2_X1 _u10_U11170  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n22474 ) );
NAND2_X1 _u10_U11169  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n22475 ) );
NAND3_X1 _u10_U11168  ( .A1(_u10_n22473 ), .A2(_u10_n22474 ), .A3(_u10_n22475 ), .ZN(_u10_n22472 ) );
NOR4_X1 _u10_U11167  ( .A1(_u10_n22469 ), .A2(_u10_n22470 ), .A3(_u10_n22471 ), .A4(_u10_n22472 ), .ZN(_u10_n22447 ) );
NAND2_X1 _u10_U11166  ( .A1(1'b0), .A2(_u10_n11996 ), .ZN(_u10_n22465 ) );
NAND2_X1 _u10_U11165  ( .A1(1'b0), .A2(_u10_n11975 ), .ZN(_u10_n22466 ) );
NAND2_X1 _u10_U11164  ( .A1(1'b0), .A2(_u10_n11951 ), .ZN(_u10_n22467 ) );
NAND2_X1 _u10_U11163  ( .A1(1'b0), .A2(_u10_n11927 ), .ZN(_u10_n22468 ) );
NAND4_X1 _u10_U11162  ( .A1(_u10_n22465 ), .A2(_u10_n22466 ), .A3(_u10_n22467 ), .A4(_u10_n22468 ), .ZN(_u10_n22449 ) );
NAND2_X1 _u10_U11161  ( .A1(1'b0), .A2(_u10_n11900 ), .ZN(_u10_n22461 ) );
NAND2_X1 _u10_U11160  ( .A1(1'b0), .A2(_u10_n11876 ), .ZN(_u10_n22462 ) );
NAND2_X1 _u10_U11159  ( .A1(1'b0), .A2(_u10_n11852 ), .ZN(_u10_n22463 ) );
NAND2_X1 _u10_U11158  ( .A1(1'b0), .A2(_u10_n11828 ), .ZN(_u10_n22464 ) );
NAND4_X1 _u10_U11157  ( .A1(_u10_n22461 ), .A2(_u10_n22462 ), .A3(_u10_n22463 ), .A4(_u10_n22464 ), .ZN(_u10_n22450 ) );
NAND2_X1 _u10_U11156  ( .A1(1'b0), .A2(_u10_n11804 ), .ZN(_u10_n22457 ) );
NAND2_X1 _u10_U11155  ( .A1(1'b0), .A2(_u10_n11780 ), .ZN(_u10_n22458 ) );
NAND2_X1 _u10_U11154  ( .A1(1'b0), .A2(_u10_n11756 ), .ZN(_u10_n22459 ) );
NAND2_X1 _u10_U11153  ( .A1(1'b0), .A2(_u10_n11732 ), .ZN(_u10_n22460 ) );
NAND4_X1 _u10_U11152  ( .A1(_u10_n22457 ), .A2(_u10_n22458 ), .A3(_u10_n22459 ), .A4(_u10_n22460 ), .ZN(_u10_n22451 ) );
NAND2_X1 _u10_U11151  ( .A1(1'b0), .A2(_u10_n11708 ), .ZN(_u10_n22453 ) );
NAND2_X1 _u10_U11150  ( .A1(1'b0), .A2(_u10_n11684 ), .ZN(_u10_n22454 ) );
NAND2_X1 _u10_U11149  ( .A1(1'b0), .A2(_u10_n11660 ), .ZN(_u10_n22455 ) );
NAND2_X1 _u10_U11148  ( .A1(1'b0), .A2(_u10_n11636 ), .ZN(_u10_n22456 ) );
NAND4_X1 _u10_U11147  ( .A1(_u10_n22453 ), .A2(_u10_n22454 ), .A3(_u10_n22455 ), .A4(_u10_n22456 ), .ZN(_u10_n22452 ) );
NOR4_X1 _u10_U11146  ( .A1(_u10_n22449 ), .A2(_u10_n22450 ), .A3(_u10_n22451 ), .A4(_u10_n22452 ), .ZN(_u10_n22448 ) );
NAND2_X1 _u10_U11145  ( .A1(_u10_n22447 ), .A2(_u10_n22448 ), .ZN(adr0[1]));
NAND2_X1 _u10_U11144  ( .A1(1'b0), .A2(_u10_n12352 ), .ZN(_u10_n22443 ) );
NAND2_X1 _u10_U11143  ( .A1(1'b0), .A2(_u10_n12332 ), .ZN(_u10_n22444 ) );
NAND2_X1 _u10_U11142  ( .A1(1'b0), .A2(_u10_n12303 ), .ZN(_u10_n22445 ) );
NAND2_X1 _u10_U11141  ( .A1(1'b0), .A2(_u10_n12279 ), .ZN(_u10_n22446 ) );
NAND4_X1 _u10_U11140  ( .A1(_u10_n22443 ), .A2(_u10_n22444 ), .A3(_u10_n22445 ), .A4(_u10_n22446 ), .ZN(_u10_n22428 ) );
NAND2_X1 _u10_U11139  ( .A1(1'b0), .A2(_u10_n12256 ), .ZN(_u10_n22439 ) );
NAND2_X1 _u10_U11138  ( .A1(1'b0), .A2(_u10_n12232 ), .ZN(_u10_n22440 ) );
NAND2_X1 _u10_U11137  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n22441 ) );
NAND2_X1 _u10_U11136  ( .A1(1'b0), .A2(_u10_n12184 ), .ZN(_u10_n22442 ) );
NAND4_X1 _u10_U11135  ( .A1(_u10_n22439 ), .A2(_u10_n22440 ), .A3(_u10_n22441 ), .A4(_u10_n22442 ), .ZN(_u10_n22429 ) );
NAND2_X1 _u10_U11134  ( .A1(1'b0), .A2(_u10_n12161 ), .ZN(_u10_n22435 ) );
NAND2_X1 _u10_U11133  ( .A1(1'b0), .A2(_u10_n12136 ), .ZN(_u10_n22436 ) );
NAND2_X1 _u10_U11132  ( .A1(1'b0), .A2(_u10_n12112 ), .ZN(_u10_n22437 ) );
NAND2_X1 _u10_U11131  ( .A1(1'b0), .A2(_u10_n12088 ), .ZN(_u10_n22438 ) );
NAND4_X1 _u10_U11130  ( .A1(_u10_n22435 ), .A2(_u10_n22436 ), .A3(_u10_n22437 ), .A4(_u10_n22438 ), .ZN(_u10_n22430 ) );
NAND2_X1 _u10_U11129  ( .A1(1'b0), .A2(_u10_n12066 ), .ZN(_u10_n22432 ) );
NAND2_X1 _u10_U11128  ( .A1(1'b0), .A2(_u10_n12042 ), .ZN(_u10_n22433 ) );
NAND2_X1 _u10_U11127  ( .A1(ch0_adr0[20]), .A2(_u10_n12014 ), .ZN(_u10_n22434 ) );
NAND3_X1 _u10_U11126  ( .A1(_u10_n22432 ), .A2(_u10_n22433 ), .A3(_u10_n22434 ), .ZN(_u10_n22431 ) );
NOR4_X1 _u10_U11125  ( .A1(_u10_n22428 ), .A2(_u10_n22429 ), .A3(_u10_n22430 ), .A4(_u10_n22431 ), .ZN(_u10_n22406 ) );
NAND2_X1 _u10_U11124  ( .A1(1'b0), .A2(_u10_n12396 ), .ZN(_u10_n22424 ) );
NAND2_X1 _u10_U11123  ( .A1(1'b0), .A2(_u10_n11971 ), .ZN(_u10_n22425 ) );
NAND2_X1 _u10_U11122  ( .A1(1'b0), .A2(_u10_n11947 ), .ZN(_u10_n22426 ) );
NAND2_X1 _u10_U11121  ( .A1(1'b0), .A2(_u10_n11923 ), .ZN(_u10_n22427 ) );
NAND4_X1 _u10_U11120  ( .A1(_u10_n22424 ), .A2(_u10_n22425 ), .A3(_u10_n22426 ), .A4(_u10_n22427 ), .ZN(_u10_n22408 ) );
NAND2_X1 _u10_U11119  ( .A1(1'b0), .A2(_u10_n11902 ), .ZN(_u10_n22420 ) );
NAND2_X1 _u10_U11118  ( .A1(1'b0), .A2(_u10_n12387 ), .ZN(_u10_n22421 ) );
NAND2_X1 _u10_U11117  ( .A1(1'b0), .A2(_u10_n11854 ), .ZN(_u10_n22422 ) );
NAND2_X1 _u10_U11116  ( .A1(1'b0), .A2(_u10_n11830 ), .ZN(_u10_n22423 ) );
NAND4_X1 _u10_U11115  ( .A1(_u10_n22420 ), .A2(_u10_n22421 ), .A3(_u10_n22422 ), .A4(_u10_n22423 ), .ZN(_u10_n22409 ) );
NAND2_X1 _u10_U11114  ( .A1(1'b0), .A2(_u10_n12380 ), .ZN(_u10_n22416 ) );
NAND2_X1 _u10_U11113  ( .A1(1'b0), .A2(_u10_n11779 ), .ZN(_u10_n22417 ) );
NAND2_X1 _u10_U11112  ( .A1(1'b0), .A2(_u10_n11758 ), .ZN(_u10_n22418 ) );
NAND2_X1 _u10_U11111  ( .A1(1'b0), .A2(_u10_n11734 ), .ZN(_u10_n22419 ) );
NAND4_X1 _u10_U11110  ( .A1(_u10_n22416 ), .A2(_u10_n22417 ), .A3(_u10_n22418 ), .A4(_u10_n22419 ), .ZN(_u10_n22410 ) );
NAND2_X1 _u10_U11109  ( .A1(1'b0), .A2(_u10_n11710 ), .ZN(_u10_n22412 ) );
NAND2_X1 _u10_U11108  ( .A1(1'b0), .A2(_u10_n11686 ), .ZN(_u10_n22413 ) );
NAND2_X1 _u10_U11107  ( .A1(1'b0), .A2(_u10_n11662 ), .ZN(_u10_n22414 ) );
NAND2_X1 _u10_U11106  ( .A1(1'b0), .A2(_u10_n11638 ), .ZN(_u10_n22415 ) );
NAND4_X1 _u10_U11105  ( .A1(_u10_n22412 ), .A2(_u10_n22413 ), .A3(_u10_n22414 ), .A4(_u10_n22415 ), .ZN(_u10_n22411 ) );
NOR4_X1 _u10_U11104  ( .A1(_u10_n22408 ), .A2(_u10_n22409 ), .A3(_u10_n22410 ), .A4(_u10_n22411 ), .ZN(_u10_n22407 ) );
NAND2_X1 _u10_U11103  ( .A1(_u10_n22406 ), .A2(_u10_n22407 ), .ZN(adr0[20]));
NAND2_X1 _u10_U11102  ( .A1(1'b0), .A2(_u10_n12352 ), .ZN(_u10_n22402 ) );
NAND2_X1 _u10_U11101  ( .A1(1'b0), .A2(_u10_n12329 ), .ZN(_u10_n22403 ) );
NAND2_X1 _u10_U11100  ( .A1(1'b0), .A2(_u10_n12303 ), .ZN(_u10_n22404 ) );
NAND2_X1 _u10_U11099  ( .A1(1'b0), .A2(_u10_n12279 ), .ZN(_u10_n22405 ) );
NAND4_X1 _u10_U11098  ( .A1(_u10_n22402 ), .A2(_u10_n22403 ), .A3(_u10_n22404 ), .A4(_u10_n22405 ), .ZN(_u10_n22387 ) );
NAND2_X1 _u10_U11097  ( .A1(1'b0), .A2(_u10_n12256 ), .ZN(_u10_n22398 ) );
NAND2_X1 _u10_U11096  ( .A1(1'b0), .A2(_u10_n12232 ), .ZN(_u10_n22399 ) );
NAND2_X1 _u10_U11095  ( .A1(1'b0), .A2(_u10_n12206 ), .ZN(_u10_n22400 ) );
NAND2_X1 _u10_U11094  ( .A1(1'b0), .A2(_u10_n12184 ), .ZN(_u10_n22401 ) );
NAND4_X1 _u10_U11093  ( .A1(_u10_n22398 ), .A2(_u10_n22399 ), .A3(_u10_n22400 ), .A4(_u10_n22401 ), .ZN(_u10_n22388 ) );
NAND2_X1 _u10_U11092  ( .A1(1'b0), .A2(_u10_n12160 ), .ZN(_u10_n22394 ) );
NAND2_X1 _u10_U11091  ( .A1(1'b0), .A2(_u10_n12139 ), .ZN(_u10_n22395 ) );
NAND2_X1 _u10_U11090  ( .A1(1'b0), .A2(_u10_n12115 ), .ZN(_u10_n22396 ) );
NAND2_X1 _u10_U11089  ( .A1(1'b0), .A2(_u10_n12091 ), .ZN(_u10_n22397 ) );
NAND4_X1 _u10_U11088  ( .A1(_u10_n22394 ), .A2(_u10_n22395 ), .A3(_u10_n22396 ), .A4(_u10_n22397 ), .ZN(_u10_n22389 ) );
NAND2_X1 _u10_U11087  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n22391 ) );
NAND2_X1 _u10_U11086  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n22392 ) );
NAND2_X1 _u10_U11085  ( .A1(ch0_adr0[21]), .A2(_u10_n12013 ), .ZN(_u10_n22393 ) );
NAND3_X1 _u10_U11084  ( .A1(_u10_n22391 ), .A2(_u10_n22392 ), .A3(_u10_n22393 ), .ZN(_u10_n22390 ) );
NOR4_X1 _u10_U11083  ( .A1(_u10_n22387 ), .A2(_u10_n22388 ), .A3(_u10_n22389 ), .A4(_u10_n22390 ), .ZN(_u10_n22365 ) );
NAND2_X1 _u10_U11082  ( .A1(1'b0), .A2(_u10_n11994 ), .ZN(_u10_n22383 ) );
NAND2_X1 _u10_U11081  ( .A1(1'b0), .A2(_u10_n11970 ), .ZN(_u10_n22384 ) );
NAND2_X1 _u10_U11080  ( .A1(1'b0), .A2(_u10_n11946 ), .ZN(_u10_n22385 ) );
NAND2_X1 _u10_U11079  ( .A1(1'b0), .A2(_u10_n11922 ), .ZN(_u10_n22386 ) );
NAND4_X1 _u10_U11078  ( .A1(_u10_n22383 ), .A2(_u10_n22384 ), .A3(_u10_n22385 ), .A4(_u10_n22386 ), .ZN(_u10_n22367 ) );
NAND2_X1 _u10_U11077  ( .A1(1'b0), .A2(_u10_n11898 ), .ZN(_u10_n22379 ) );
NAND2_X1 _u10_U11076  ( .A1(1'b0), .A2(_u10_n11874 ), .ZN(_u10_n22380 ) );
NAND2_X1 _u10_U11075  ( .A1(1'b0), .A2(_u10_n11850 ), .ZN(_u10_n22381 ) );
NAND2_X1 _u10_U11074  ( .A1(1'b0), .A2(_u10_n11826 ), .ZN(_u10_n22382 ) );
NAND4_X1 _u10_U11073  ( .A1(_u10_n22379 ), .A2(_u10_n22380 ), .A3(_u10_n22381 ), .A4(_u10_n22382 ), .ZN(_u10_n22368 ) );
NAND2_X1 _u10_U11072  ( .A1(1'b0), .A2(_u10_n11802 ), .ZN(_u10_n22375 ) );
NAND2_X1 _u10_U11071  ( .A1(1'b0), .A2(_u10_n11778 ), .ZN(_u10_n22376 ) );
NAND2_X1 _u10_U11070  ( .A1(1'b0), .A2(_u10_n11754 ), .ZN(_u10_n22377 ) );
NAND2_X1 _u10_U11069  ( .A1(1'b0), .A2(_u10_n11730 ), .ZN(_u10_n22378 ) );
NAND4_X1 _u10_U11068  ( .A1(_u10_n22375 ), .A2(_u10_n22376 ), .A3(_u10_n22377 ), .A4(_u10_n22378 ), .ZN(_u10_n22369 ) );
NAND2_X1 _u10_U11067  ( .A1(1'b0), .A2(_u10_n11706 ), .ZN(_u10_n22371 ) );
NAND2_X1 _u10_U11066  ( .A1(1'b0), .A2(_u10_n11682 ), .ZN(_u10_n22372 ) );
NAND2_X1 _u10_U11065  ( .A1(1'b0), .A2(_u10_n11658 ), .ZN(_u10_n22373 ) );
NAND2_X1 _u10_U11064  ( .A1(1'b0), .A2(_u10_n11634 ), .ZN(_u10_n22374 ) );
NAND4_X1 _u10_U11063  ( .A1(_u10_n22371 ), .A2(_u10_n22372 ), .A3(_u10_n22373 ), .A4(_u10_n22374 ), .ZN(_u10_n22370 ) );
NOR4_X1 _u10_U11062  ( .A1(_u10_n22367 ), .A2(_u10_n22368 ), .A3(_u10_n22369 ), .A4(_u10_n22370 ), .ZN(_u10_n22366 ) );
NAND2_X1 _u10_U11061  ( .A1(_u10_n22365 ), .A2(_u10_n22366 ), .ZN(adr0[21]));
NAND2_X1 _u10_U11060  ( .A1(1'b0), .A2(_u10_n12356 ), .ZN(_u10_n22361 ) );
NAND2_X1 _u10_U11059  ( .A1(1'b0), .A2(_u10_n12332 ), .ZN(_u10_n22362 ) );
NAND2_X1 _u10_U11058  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n22363 ) );
NAND2_X1 _u10_U11057  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n22364 ) );
NAND4_X1 _u10_U11056  ( .A1(_u10_n22361 ), .A2(_u10_n22362 ), .A3(_u10_n22363 ), .A4(_u10_n22364 ), .ZN(_u10_n22346 ) );
NAND2_X1 _u10_U11055  ( .A1(1'b0), .A2(_u10_n12260 ), .ZN(_u10_n22357 ) );
NAND2_X1 _u10_U11054  ( .A1(1'b0), .A2(_u10_n12236 ), .ZN(_u10_n22358 ) );
NAND2_X1 _u10_U11053  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n22359 ) );
NAND2_X1 _u10_U11052  ( .A1(1'b0), .A2(_u10_n12188 ), .ZN(_u10_n22360 ) );
NAND4_X1 _u10_U11051  ( .A1(_u10_n22357 ), .A2(_u10_n22358 ), .A3(_u10_n22359 ), .A4(_u10_n22360 ), .ZN(_u10_n22347 ) );
NAND2_X1 _u10_U11050  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n22353 ) );
NAND2_X1 _u10_U11049  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n22354 ) );
NAND2_X1 _u10_U11048  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n22355 ) );
NAND2_X1 _u10_U11047  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n22356 ) );
NAND4_X1 _u10_U11046  ( .A1(_u10_n22353 ), .A2(_u10_n22354 ), .A3(_u10_n22355 ), .A4(_u10_n22356 ), .ZN(_u10_n22348 ) );
NAND2_X1 _u10_U11045  ( .A1(1'b0), .A2(_u10_n12068 ), .ZN(_u10_n22350 ) );
NAND2_X1 _u10_U11044  ( .A1(1'b0), .A2(_u10_n12044 ), .ZN(_u10_n22351 ) );
NAND2_X1 _u10_U11043  ( .A1(ch0_adr0[22]), .A2(_u10_n12012 ), .ZN(_u10_n22352 ) );
NAND3_X1 _u10_U11042  ( .A1(_u10_n22350 ), .A2(_u10_n22351 ), .A3(_u10_n22352 ), .ZN(_u10_n22349 ) );
NOR4_X1 _u10_U11041  ( .A1(_u10_n22346 ), .A2(_u10_n22347 ), .A3(_u10_n22348 ), .A4(_u10_n22349 ), .ZN(_u10_n22324 ) );
NAND2_X1 _u10_U11040  ( .A1(1'b0), .A2(_u10_n11995 ), .ZN(_u10_n22342 ) );
NAND2_X1 _u10_U11039  ( .A1(1'b0), .A2(_u10_n11972 ), .ZN(_u10_n22343 ) );
NAND2_X1 _u10_U11038  ( .A1(1'b0), .A2(_u10_n11947 ), .ZN(_u10_n22344 ) );
NAND2_X1 _u10_U11037  ( .A1(1'b0), .A2(_u10_n11923 ), .ZN(_u10_n22345 ) );
NAND4_X1 _u10_U11035  ( .A1(_u10_n22342 ), .A2(_u10_n22343 ), .A3(_u10_n22344 ), .A4(_u10_n22345 ), .ZN(_u10_n22326 ) );
NAND2_X1 _u10_U11034  ( .A1(1'b0), .A2(_u10_n11899 ), .ZN(_u10_n22338 ) );
NAND2_X1 _u10_U11033  ( .A1(1'b0), .A2(_u10_n11875 ), .ZN(_u10_n22339 ) );
NAND2_X1 _u10_U11032  ( .A1(1'b0), .A2(_u10_n11851 ), .ZN(_u10_n22340 ) );
NAND2_X1 _u10_U11031  ( .A1(1'b0), .A2(_u10_n11827 ), .ZN(_u10_n22341 ) );
NAND4_X1 _u10_U11030  ( .A1(_u10_n22338 ), .A2(_u10_n22339 ), .A3(_u10_n22340 ), .A4(_u10_n22341 ), .ZN(_u10_n22327 ) );
NAND2_X1 _u10_U11029  ( .A1(1'b0), .A2(_u10_n11803 ), .ZN(_u10_n22334 ) );
NAND2_X1 _u10_U11028  ( .A1(1'b0), .A2(_u10_n11779 ), .ZN(_u10_n22335 ) );
NAND2_X1 _u10_U11027  ( .A1(1'b0), .A2(_u10_n11755 ), .ZN(_u10_n22336 ) );
NAND2_X1 _u10_U11026  ( .A1(1'b0), .A2(_u10_n11731 ), .ZN(_u10_n22337 ) );
NAND4_X1 _u10_U11025  ( .A1(_u10_n22334 ), .A2(_u10_n22335 ), .A3(_u10_n22336 ), .A4(_u10_n22337 ), .ZN(_u10_n22328 ) );
NAND2_X1 _u10_U11024  ( .A1(1'b0), .A2(_u10_n11707 ), .ZN(_u10_n22330 ) );
NAND2_X1 _u10_U11023  ( .A1(1'b0), .A2(_u10_n11683 ), .ZN(_u10_n22331 ) );
NAND2_X1 _u10_U11022  ( .A1(1'b0), .A2(_u10_n11659 ), .ZN(_u10_n22332 ) );
NAND2_X1 _u10_U11021  ( .A1(1'b0), .A2(_u10_n11635 ), .ZN(_u10_n22333 ) );
NAND4_X1 _u10_U11020  ( .A1(_u10_n22330 ), .A2(_u10_n22331 ), .A3(_u10_n22332 ), .A4(_u10_n22333 ), .ZN(_u10_n22329 ) );
NOR4_X1 _u10_U11019  ( .A1(_u10_n22326 ), .A2(_u10_n22327 ), .A3(_u10_n22328 ), .A4(_u10_n22329 ), .ZN(_u10_n22325 ) );
NAND2_X1 _u10_U11018  ( .A1(_u10_n22324 ), .A2(_u10_n22325 ), .ZN(adr0[22]));
NAND2_X1 _u10_U11017  ( .A1(1'b0), .A2(_u10_n12354 ), .ZN(_u10_n22320 ) );
NAND2_X1 _u10_U11016  ( .A1(1'b0), .A2(_u10_n12331 ), .ZN(_u10_n22321 ) );
NAND2_X1 _u10_U11015  ( .A1(1'b0), .A2(_u10_n12307 ), .ZN(_u10_n22322 ) );
NAND2_X1 _u10_U11014  ( .A1(1'b0), .A2(_u10_n12283 ), .ZN(_u10_n22323 ) );
NAND4_X1 _u10_U11013  ( .A1(_u10_n22320 ), .A2(_u10_n22321 ), .A3(_u10_n22322 ), .A4(_u10_n22323 ), .ZN(_u10_n22305 ) );
NAND2_X1 _u10_U11012  ( .A1(1'b0), .A2(_u10_n12258 ), .ZN(_u10_n22316 ) );
NAND2_X1 _u10_U11011  ( .A1(1'b0), .A2(_u10_n12234 ), .ZN(_u10_n22317 ) );
NAND2_X1 _u10_U11010  ( .A1(1'b0), .A2(_u10_n12209 ), .ZN(_u10_n22318 ) );
NAND2_X1 _u10_U11009  ( .A1(1'b0), .A2(_u10_n12186 ), .ZN(_u10_n22319 ) );
NAND4_X1 _u10_U11008  ( .A1(_u10_n22316 ), .A2(_u10_n22317 ), .A3(_u10_n22318 ), .A4(_u10_n22319 ), .ZN(_u10_n22306 ) );
NAND2_X1 _u10_U11007  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n22312 ) );
NAND2_X1 _u10_U11006  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n22313 ) );
NAND2_X1 _u10_U11005  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n22314 ) );
NAND2_X1 _u10_U11004  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n22315 ) );
NAND4_X1 _u10_U11003  ( .A1(_u10_n22312 ), .A2(_u10_n22313 ), .A3(_u10_n22314 ), .A4(_u10_n22315 ), .ZN(_u10_n22307 ) );
NAND2_X1 _u10_U11002  ( .A1(1'b0), .A2(_u10_n12065 ), .ZN(_u10_n22309 ) );
NAND2_X1 _u10_U11001  ( .A1(1'b0), .A2(_u10_n12041 ), .ZN(_u10_n22310 ) );
NAND2_X1 _u10_U11000  ( .A1(ch0_adr0[23]), .A2(_u10_n12011 ), .ZN(_u10_n22311 ) );
NAND3_X1 _u10_U10999  ( .A1(_u10_n22309 ), .A2(_u10_n22310 ), .A3(_u10_n22311 ), .ZN(_u10_n22308 ) );
NOR4_X1 _u10_U10998  ( .A1(_u10_n22305 ), .A2(_u10_n22306 ), .A3(_u10_n22307 ), .A4(_u10_n22308 ), .ZN(_u10_n22283 ) );
NAND2_X1 _u10_U10997  ( .A1(1'b0), .A2(_u10_n11997 ), .ZN(_u10_n22301 ) );
NAND2_X1 _u10_U10996  ( .A1(1'b0), .A2(_u10_n11973 ), .ZN(_u10_n22302 ) );
NAND2_X1 _u10_U10995  ( .A1(1'b0), .A2(_u10_n11949 ), .ZN(_u10_n22303 ) );
NAND2_X1 _u10_U10994  ( .A1(1'b0), .A2(_u10_n11925 ), .ZN(_u10_n22304 ) );
NAND4_X1 _u10_U10993  ( .A1(_u10_n22301 ), .A2(_u10_n22302 ), .A3(_u10_n22303 ), .A4(_u10_n22304 ), .ZN(_u10_n22285 ) );
NAND2_X1 _u10_U10992  ( .A1(1'b0), .A2(_u10_n11901 ), .ZN(_u10_n22297 ) );
NAND2_X1 _u10_U10991  ( .A1(1'b0), .A2(_u10_n11877 ), .ZN(_u10_n22298 ) );
NAND2_X1 _u10_U10990  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n22299 ) );
NAND2_X1 _u10_U10989  ( .A1(1'b0), .A2(_u10_n11829 ), .ZN(_u10_n22300 ) );
NAND4_X1 _u10_U10988  ( .A1(_u10_n22297 ), .A2(_u10_n22298 ), .A3(_u10_n22299 ), .A4(_u10_n22300 ), .ZN(_u10_n22286 ) );
NAND2_X1 _u10_U10987  ( .A1(1'b0), .A2(_u10_n11805 ), .ZN(_u10_n22293 ) );
NAND2_X1 _u10_U10986  ( .A1(1'b0), .A2(_u10_n11781 ), .ZN(_u10_n22294 ) );
NAND2_X1 _u10_U10985  ( .A1(1'b0), .A2(_u10_n11757 ), .ZN(_u10_n22295 ) );
NAND2_X1 _u10_U10984  ( .A1(1'b0), .A2(_u10_n11733 ), .ZN(_u10_n22296 ) );
NAND4_X1 _u10_U10983  ( .A1(_u10_n22293 ), .A2(_u10_n22294 ), .A3(_u10_n22295 ), .A4(_u10_n22296 ), .ZN(_u10_n22287 ) );
NAND2_X1 _u10_U10982  ( .A1(1'b0), .A2(_u10_n11709 ), .ZN(_u10_n22289 ) );
NAND2_X1 _u10_U10981  ( .A1(1'b0), .A2(_u10_n11685 ), .ZN(_u10_n22290 ) );
NAND2_X1 _u10_U10980  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n22291 ) );
NAND2_X1 _u10_U10979  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n22292 ) );
NAND4_X1 _u10_U10978  ( .A1(_u10_n22289 ), .A2(_u10_n22290 ), .A3(_u10_n22291 ), .A4(_u10_n22292 ), .ZN(_u10_n22288 ) );
NOR4_X1 _u10_U10977  ( .A1(_u10_n22285 ), .A2(_u10_n22286 ), .A3(_u10_n22287 ), .A4(_u10_n22288 ), .ZN(_u10_n22284 ) );
NAND2_X1 _u10_U10976  ( .A1(_u10_n22283 ), .A2(_u10_n22284 ), .ZN(adr0[23]));
NAND2_X1 _u10_U10975  ( .A1(1'b0), .A2(_u10_n12355 ), .ZN(_u10_n22279 ) );
NAND2_X1 _u10_U10974  ( .A1(1'b0), .A2(_u10_n12330 ), .ZN(_u10_n22280 ) );
NAND2_X1 _u10_U10973  ( .A1(1'b0), .A2(_u10_n12306 ), .ZN(_u10_n22281 ) );
NAND2_X1 _u10_U10972  ( .A1(1'b0), .A2(_u10_n12282 ), .ZN(_u10_n22282 ) );
NAND4_X1 _u10_U10971  ( .A1(_u10_n22279 ), .A2(_u10_n22280 ), .A3(_u10_n22281 ), .A4(_u10_n22282 ), .ZN(_u10_n22264 ) );
NAND2_X1 _u10_U10970  ( .A1(1'b0), .A2(_u10_n12259 ), .ZN(_u10_n22275 ) );
NAND2_X1 _u10_U10969  ( .A1(1'b0), .A2(_u10_n12235 ), .ZN(_u10_n22276 ) );
NAND2_X1 _u10_U10968  ( .A1(1'b0), .A2(_u10_n12211 ), .ZN(_u10_n22277 ) );
NAND2_X1 _u10_U10967  ( .A1(1'b0), .A2(_u10_n12187 ), .ZN(_u10_n22278 ) );
NAND4_X1 _u10_U10966  ( .A1(_u10_n22275 ), .A2(_u10_n22276 ), .A3(_u10_n22277 ), .A4(_u10_n22278 ), .ZN(_u10_n22265 ) );
NAND2_X1 _u10_U10965  ( .A1(1'b0), .A2(_u10_n12161 ), .ZN(_u10_n22271 ) );
NAND2_X1 _u10_U10964  ( .A1(1'b0), .A2(_u10_n12137 ), .ZN(_u10_n22272 ) );
NAND2_X1 _u10_U10963  ( .A1(1'b0), .A2(_u10_n12113 ), .ZN(_u10_n22273 ) );
NAND2_X1 _u10_U10962  ( .A1(1'b0), .A2(_u10_n12089 ), .ZN(_u10_n22274 ) );
NAND4_X1 _u10_U10961  ( .A1(_u10_n22271 ), .A2(_u10_n22272 ), .A3(_u10_n22273 ), .A4(_u10_n22274 ), .ZN(_u10_n22266 ) );
NAND2_X1 _u10_U10960  ( .A1(1'b0), .A2(_u10_n12067 ), .ZN(_u10_n22268 ) );
NAND2_X1 _u10_U10959  ( .A1(1'b0), .A2(_u10_n12043 ), .ZN(_u10_n22269 ) );
NAND2_X1 _u10_U10958  ( .A1(ch0_adr0[24]), .A2(_u10_n12020 ), .ZN(_u10_n22270 ) );
NAND3_X1 _u10_U10957  ( .A1(_u10_n22268 ), .A2(_u10_n22269 ), .A3(_u10_n22270 ), .ZN(_u10_n22267 ) );
NOR4_X1 _u10_U10956  ( .A1(_u10_n22264 ), .A2(_u10_n22265 ), .A3(_u10_n22266 ), .A4(_u10_n22267 ), .ZN(_u10_n22242 ) );
NAND2_X1 _u10_U10955  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n22260 ) );
NAND2_X1 _u10_U10954  ( .A1(1'b0), .A2(_u10_n11970 ), .ZN(_u10_n22261 ) );
NAND2_X1 _u10_U10953  ( .A1(1'b0), .A2(_u10_n11946 ), .ZN(_u10_n22262 ) );
NAND2_X1 _u10_U10952  ( .A1(1'b0), .A2(_u10_n11922 ), .ZN(_u10_n22263 ) );
NAND4_X1 _u10_U10951  ( .A1(_u10_n22260 ), .A2(_u10_n22261 ), .A3(_u10_n22262 ), .A4(_u10_n22263 ), .ZN(_u10_n22244 ) );
NAND2_X1 _u10_U10950  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n22256 ) );
NAND2_X1 _u10_U10949  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n22257 ) );
NAND2_X1 _u10_U10948  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n22258 ) );
NAND2_X1 _u10_U10947  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n22259 ) );
NAND4_X1 _u10_U10946  ( .A1(_u10_n22256 ), .A2(_u10_n22257 ), .A3(_u10_n22258 ), .A4(_u10_n22259 ), .ZN(_u10_n22245 ) );
NAND2_X1 _u10_U10945  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n22252 ) );
NAND2_X1 _u10_U10944  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n22253 ) );
NAND2_X1 _u10_U10943  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n22254 ) );
NAND2_X1 _u10_U10942  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n22255 ) );
NAND4_X1 _u10_U10941  ( .A1(_u10_n22252 ), .A2(_u10_n22253 ), .A3(_u10_n22254 ), .A4(_u10_n22255 ), .ZN(_u10_n22246 ) );
NAND2_X1 _u10_U10940  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n22248 ) );
NAND2_X1 _u10_U10939  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n22249 ) );
NAND2_X1 _u10_U10938  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n22250 ) );
NAND2_X1 _u10_U10937  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n22251 ) );
NAND4_X1 _u10_U10936  ( .A1(_u10_n22248 ), .A2(_u10_n22249 ), .A3(_u10_n22250 ), .A4(_u10_n22251 ), .ZN(_u10_n22247 ) );
NOR4_X1 _u10_U10935  ( .A1(_u10_n22244 ), .A2(_u10_n22245 ), .A3(_u10_n22246 ), .A4(_u10_n22247 ), .ZN(_u10_n22243 ) );
NAND2_X1 _u10_U10934  ( .A1(_u10_n22242 ), .A2(_u10_n22243 ), .ZN(adr0[24]));
NAND2_X1 _u10_U10933  ( .A1(1'b0), .A2(_u10_n12356 ), .ZN(_u10_n22238 ) );
NAND2_X1 _u10_U10932  ( .A1(1'b0), .A2(_u10_n12329 ), .ZN(_u10_n22239 ) );
NAND2_X1 _u10_U10931  ( .A1(1'b0), .A2(_u10_n12305 ), .ZN(_u10_n22240 ) );
NAND2_X1 _u10_U10930  ( .A1(1'b0), .A2(_u10_n12281 ), .ZN(_u10_n22241 ) );
NAND4_X1 _u10_U10929  ( .A1(_u10_n22238 ), .A2(_u10_n22239 ), .A3(_u10_n22240 ), .A4(_u10_n22241 ), .ZN(_u10_n22223 ) );
NAND2_X1 _u10_U10928  ( .A1(1'b0), .A2(_u10_n12260 ), .ZN(_u10_n22234 ) );
NAND2_X1 _u10_U10927  ( .A1(1'b0), .A2(_u10_n12236 ), .ZN(_u10_n22235 ) );
NAND2_X1 _u10_U10926  ( .A1(1'b0), .A2(_u10_n12210 ), .ZN(_u10_n22236 ) );
NAND2_X1 _u10_U10925  ( .A1(1'b0), .A2(_u10_n12188 ), .ZN(_u10_n22237 ) );
NAND4_X1 _u10_U10924  ( .A1(_u10_n22234 ), .A2(_u10_n22235 ), .A3(_u10_n22236 ), .A4(_u10_n22237 ), .ZN(_u10_n22224 ) );
NAND2_X1 _u10_U10923  ( .A1(1'b0), .A2(_u10_n12163 ), .ZN(_u10_n22230 ) );
NAND2_X1 _u10_U10922  ( .A1(1'b0), .A2(_u10_n12139 ), .ZN(_u10_n22231 ) );
NAND2_X1 _u10_U10921  ( .A1(1'b0), .A2(_u10_n12115 ), .ZN(_u10_n22232 ) );
NAND2_X1 _u10_U10920  ( .A1(1'b0), .A2(_u10_n12091 ), .ZN(_u10_n22233 ) );
NAND4_X1 _u10_U10919  ( .A1(_u10_n22230 ), .A2(_u10_n22231 ), .A3(_u10_n22232 ), .A4(_u10_n22233 ), .ZN(_u10_n22225 ) );
NAND2_X1 _u10_U10918  ( .A1(1'b0), .A2(_u10_n12066 ), .ZN(_u10_n22227 ) );
NAND2_X1 _u10_U10917  ( .A1(1'b0), .A2(_u10_n12042 ), .ZN(_u10_n22228 ) );
NAND2_X1 _u10_U10916  ( .A1(ch0_adr0[25]), .A2(_u10_n12020 ), .ZN(_u10_n22229 ) );
NAND3_X1 _u10_U10915  ( .A1(_u10_n22227 ), .A2(_u10_n22228 ), .A3(_u10_n22229 ), .ZN(_u10_n22226 ) );
NOR4_X1 _u10_U10914  ( .A1(_u10_n22223 ), .A2(_u10_n22224 ), .A3(_u10_n22225 ), .A4(_u10_n22226 ), .ZN(_u10_n22201 ) );
NAND2_X1 _u10_U10913  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n22219 ) );
NAND2_X1 _u10_U10912  ( .A1(1'b0), .A2(_u10_n12395 ), .ZN(_u10_n22220 ) );
NAND2_X1 _u10_U10911  ( .A1(1'b0), .A2(_u10_n11951 ), .ZN(_u10_n22221 ) );
NAND2_X1 _u10_U10910  ( .A1(1'b0), .A2(_u10_n11927 ), .ZN(_u10_n22222 ) );
NAND4_X1 _u10_U10909  ( .A1(_u10_n22219 ), .A2(_u10_n22220 ), .A3(_u10_n22221 ), .A4(_u10_n22222 ), .ZN(_u10_n22203 ) );
NAND2_X1 _u10_U10908  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n22215 ) );
NAND2_X1 _u10_U10907  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n22216 ) );
NAND2_X1 _u10_U10906  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n22217 ) );
NAND2_X1 _u10_U10905  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n22218 ) );
NAND4_X1 _u10_U10904  ( .A1(_u10_n22215 ), .A2(_u10_n22216 ), .A3(_u10_n22217 ), .A4(_u10_n22218 ), .ZN(_u10_n22204 ) );
NAND2_X1 _u10_U10903  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n22211 ) );
NAND2_X1 _u10_U10902  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n22212 ) );
NAND2_X1 _u10_U10901  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n22213 ) );
NAND2_X1 _u10_U10900  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n22214 ) );
NAND4_X1 _u10_U10899  ( .A1(_u10_n22211 ), .A2(_u10_n22212 ), .A3(_u10_n22213 ), .A4(_u10_n22214 ), .ZN(_u10_n22205 ) );
NAND2_X1 _u10_U10898  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n22207 ) );
NAND2_X1 _u10_U10897  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n22208 ) );
NAND2_X1 _u10_U10896  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n22209 ) );
NAND2_X1 _u10_U10895  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n22210 ) );
NAND4_X1 _u10_U10894  ( .A1(_u10_n22207 ), .A2(_u10_n22208 ), .A3(_u10_n22209 ), .A4(_u10_n22210 ), .ZN(_u10_n22206 ) );
NOR4_X1 _u10_U10893  ( .A1(_u10_n22203 ), .A2(_u10_n22204 ), .A3(_u10_n22205 ), .A4(_u10_n22206 ), .ZN(_u10_n22202 ) );
NAND2_X1 _u10_U10892  ( .A1(_u10_n22201 ), .A2(_u10_n22202 ), .ZN(adr0[25]));
NAND2_X1 _u10_U10891  ( .A1(1'b0), .A2(_u10_n12353 ), .ZN(_u10_n22197 ) );
NAND2_X1 _u10_U10890  ( .A1(1'b0), .A2(_u10_n12328 ), .ZN(_u10_n22198 ) );
NAND2_X1 _u10_U10889  ( .A1(1'b0), .A2(_u10_n12304 ), .ZN(_u10_n22199 ) );
NAND2_X1 _u10_U10888  ( .A1(1'b0), .A2(_u10_n12280 ), .ZN(_u10_n22200 ) );
NAND4_X1 _u10_U10887  ( .A1(_u10_n22197 ), .A2(_u10_n22198 ), .A3(_u10_n22199 ), .A4(_u10_n22200 ), .ZN(_u10_n22182 ) );
NAND2_X1 _u10_U10886  ( .A1(1'b0), .A2(_u10_n12257 ), .ZN(_u10_n22193 ) );
NAND2_X1 _u10_U10885  ( .A1(1'b0), .A2(_u10_n12233 ), .ZN(_u10_n22194 ) );
NAND2_X1 _u10_U10884  ( .A1(1'b0), .A2(_u10_n12207 ), .ZN(_u10_n22195 ) );
NAND2_X1 _u10_U10883  ( .A1(1'b0), .A2(_u10_n12185 ), .ZN(_u10_n22196 ) );
NAND4_X1 _u10_U10882  ( .A1(_u10_n22193 ), .A2(_u10_n22194 ), .A3(_u10_n22195 ), .A4(_u10_n22196 ), .ZN(_u10_n22183 ) );
NAND2_X1 _u10_U10881  ( .A1(1'b0), .A2(_u10_n12162 ), .ZN(_u10_n22189 ) );
NAND2_X1 _u10_U10880  ( .A1(1'b0), .A2(_u10_n12138 ), .ZN(_u10_n22190 ) );
NAND2_X1 _u10_U10879  ( .A1(1'b0), .A2(_u10_n12114 ), .ZN(_u10_n22191 ) );
NAND2_X1 _u10_U10878  ( .A1(1'b0), .A2(_u10_n12090 ), .ZN(_u10_n22192 ) );
NAND4_X1 _u10_U10877  ( .A1(_u10_n22189 ), .A2(_u10_n22190 ), .A3(_u10_n22191 ), .A4(_u10_n22192 ), .ZN(_u10_n22184 ) );
NAND2_X1 _u10_U10876  ( .A1(1'b0), .A2(_u10_n12063 ), .ZN(_u10_n22186 ) );
NAND2_X1 _u10_U10875  ( .A1(1'b0), .A2(_u10_n12039 ), .ZN(_u10_n22187 ) );
NAND2_X1 _u10_U10874  ( .A1(ch0_adr0[26]), .A2(_u10_n12020 ), .ZN(_u10_n22188 ) );
NAND3_X1 _u10_U10873  ( .A1(_u10_n22186 ), .A2(_u10_n22187 ), .A3(_u10_n22188 ), .ZN(_u10_n22185 ) );
NOR4_X1 _u10_U10872  ( .A1(_u10_n22182 ), .A2(_u10_n22183 ), .A3(_u10_n22184 ), .A4(_u10_n22185 ), .ZN(_u10_n22160 ) );
NAND2_X1 _u10_U10871  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n22178 ) );
NAND2_X1 _u10_U10870  ( .A1(1'b0), .A2(_u10_n11974 ), .ZN(_u10_n22179 ) );
NAND2_X1 _u10_U10869  ( .A1(1'b0), .A2(_u10_n12394 ), .ZN(_u10_n22180 ) );
NAND2_X1 _u10_U10868  ( .A1(1'b0), .A2(_u10_n12393 ), .ZN(_u10_n22181 ) );
NAND4_X1 _u10_U10867  ( .A1(_u10_n22178 ), .A2(_u10_n22179 ), .A3(_u10_n22180 ), .A4(_u10_n22181 ), .ZN(_u10_n22162 ) );
NAND2_X1 _u10_U10866  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n22174 ) );
NAND2_X1 _u10_U10865  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n22175 ) );
NAND2_X1 _u10_U10864  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n22176 ) );
NAND2_X1 _u10_U10863  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n22177 ) );
NAND4_X1 _u10_U10862  ( .A1(_u10_n22174 ), .A2(_u10_n22175 ), .A3(_u10_n22176 ), .A4(_u10_n22177 ), .ZN(_u10_n22163 ) );
NAND2_X1 _u10_U10861  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n22170 ) );
NAND2_X1 _u10_U10860  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n22171 ) );
NAND2_X1 _u10_U10859  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n22172 ) );
NAND2_X1 _u10_U10858  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n22173 ) );
NAND4_X1 _u10_U10857  ( .A1(_u10_n22170 ), .A2(_u10_n22171 ), .A3(_u10_n22172 ), .A4(_u10_n22173 ), .ZN(_u10_n22164 ) );
NAND2_X1 _u10_U10856  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n22166 ) );
NAND2_X1 _u10_U10855  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n22167 ) );
NAND2_X1 _u10_U10854  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n22168 ) );
NAND2_X1 _u10_U10853  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n22169 ) );
NAND4_X1 _u10_U10852  ( .A1(_u10_n22166 ), .A2(_u10_n22167 ), .A3(_u10_n22168 ), .A4(_u10_n22169 ), .ZN(_u10_n22165 ) );
NOR4_X1 _u10_U10851  ( .A1(_u10_n22162 ), .A2(_u10_n22163 ), .A3(_u10_n22164 ), .A4(_u10_n22165 ), .ZN(_u10_n22161 ) );
NAND2_X1 _u10_U10850  ( .A1(_u10_n22160 ), .A2(_u10_n22161 ), .ZN(adr0[26]));
NAND2_X1 _u10_U10849  ( .A1(1'b0), .A2(_u10_n12353 ), .ZN(_u10_n22156 ) );
NAND2_X1 _u10_U10848  ( .A1(1'b0), .A2(_u10_n12329 ), .ZN(_u10_n22157 ) );
NAND2_X1 _u10_U10847  ( .A1(1'b0), .A2(_u10_n12307 ), .ZN(_u10_n22158 ) );
NAND2_X1 _u10_U10846  ( .A1(1'b0), .A2(_u10_n12283 ), .ZN(_u10_n22159 ) );
NAND4_X1 _u10_U10845  ( .A1(_u10_n22156 ), .A2(_u10_n22157 ), .A3(_u10_n22158 ), .A4(_u10_n22159 ), .ZN(_u10_n22141 ) );
NAND2_X1 _u10_U10844  ( .A1(1'b0), .A2(_u10_n12257 ), .ZN(_u10_n22152 ) );
NAND2_X1 _u10_U10843  ( .A1(1'b0), .A2(_u10_n12233 ), .ZN(_u10_n22153 ) );
NAND2_X1 _u10_U10842  ( .A1(1'b0), .A2(_u10_n12209 ), .ZN(_u10_n22154 ) );
NAND2_X1 _u10_U10841  ( .A1(1'b0), .A2(_u10_n12185 ), .ZN(_u10_n22155 ) );
NAND4_X1 _u10_U10840  ( .A1(_u10_n22152 ), .A2(_u10_n22153 ), .A3(_u10_n22154 ), .A4(_u10_n22155 ), .ZN(_u10_n22142 ) );
NAND2_X1 _u10_U10839  ( .A1(1'b0), .A2(_u10_n12159 ), .ZN(_u10_n22148 ) );
NAND2_X1 _u10_U10838  ( .A1(1'b0), .A2(_u10_n12135 ), .ZN(_u10_n22149 ) );
NAND2_X1 _u10_U10837  ( .A1(1'b0), .A2(_u10_n12111 ), .ZN(_u10_n22150 ) );
NAND2_X1 _u10_U10836  ( .A1(1'b0), .A2(_u10_n12087 ), .ZN(_u10_n22151 ) );
NAND4_X1 _u10_U10835  ( .A1(_u10_n22148 ), .A2(_u10_n22149 ), .A3(_u10_n22150 ), .A4(_u10_n22151 ), .ZN(_u10_n22143 ) );
NAND2_X1 _u10_U10834  ( .A1(1'b0), .A2(_u10_n12066 ), .ZN(_u10_n22145 ) );
NAND2_X1 _u10_U10833  ( .A1(1'b0), .A2(_u10_n12042 ), .ZN(_u10_n22146 ) );
NAND2_X1 _u10_U10832  ( .A1(ch0_adr0[27]), .A2(_u10_n12020 ), .ZN(_u10_n22147 ) );
NAND3_X1 _u10_U10831  ( .A1(_u10_n22145 ), .A2(_u10_n22146 ), .A3(_u10_n22147 ), .ZN(_u10_n22144 ) );
NOR4_X1 _u10_U10830  ( .A1(_u10_n22141 ), .A2(_u10_n22142 ), .A3(_u10_n22143 ), .A4(_u10_n22144 ), .ZN(_u10_n22119 ) );
NAND2_X1 _u10_U10829  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n22137 ) );
NAND2_X1 _u10_U10828  ( .A1(1'b0), .A2(_u10_n11975 ), .ZN(_u10_n22138 ) );
NAND2_X1 _u10_U10827  ( .A1(1'b0), .A2(_u10_n11950 ), .ZN(_u10_n22139 ) );
NAND2_X1 _u10_U10826  ( .A1(1'b0), .A2(_u10_n11926 ), .ZN(_u10_n22140 ) );
NAND4_X1 _u10_U10825  ( .A1(_u10_n22137 ), .A2(_u10_n22138 ), .A3(_u10_n22139 ), .A4(_u10_n22140 ), .ZN(_u10_n22121 ) );
NAND2_X1 _u10_U10824  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n22133 ) );
NAND2_X1 _u10_U10823  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n22134 ) );
NAND2_X1 _u10_U10822  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n22135 ) );
NAND2_X1 _u10_U10821  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n22136 ) );
NAND4_X1 _u10_U10820  ( .A1(_u10_n22133 ), .A2(_u10_n22134 ), .A3(_u10_n22135 ), .A4(_u10_n22136 ), .ZN(_u10_n22122 ) );
NAND2_X1 _u10_U10819  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n22129 ) );
NAND2_X1 _u10_U10818  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n22130 ) );
NAND2_X1 _u10_U10817  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n22131 ) );
NAND2_X1 _u10_U10816  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n22132 ) );
NAND4_X1 _u10_U10815  ( .A1(_u10_n22129 ), .A2(_u10_n22130 ), .A3(_u10_n22131 ), .A4(_u10_n22132 ), .ZN(_u10_n22123 ) );
NAND2_X1 _u10_U10814  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n22125 ) );
NAND2_X1 _u10_U10813  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n22126 ) );
NAND2_X1 _u10_U10812  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n22127 ) );
NAND2_X1 _u10_U10811  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n22128 ) );
NAND4_X1 _u10_U10810  ( .A1(_u10_n22125 ), .A2(_u10_n22126 ), .A3(_u10_n22127 ), .A4(_u10_n22128 ), .ZN(_u10_n22124 ) );
NOR4_X1 _u10_U10809  ( .A1(_u10_n22121 ), .A2(_u10_n22122 ), .A3(_u10_n22123 ), .A4(_u10_n22124 ), .ZN(_u10_n22120 ) );
NAND2_X1 _u10_U10808  ( .A1(_u10_n22119 ), .A2(_u10_n22120 ), .ZN(adr0[27]));
NAND2_X1 _u10_U10807  ( .A1(1'b0), .A2(_u10_n12354 ), .ZN(_u10_n22115 ) );
NAND2_X1 _u10_U10806  ( .A1(1'b0), .A2(_u10_n12332 ), .ZN(_u10_n22116 ) );
NAND2_X1 _u10_U10805  ( .A1(1'b0), .A2(_u10_n12306 ), .ZN(_u10_n22117 ) );
NAND2_X1 _u10_U10804  ( .A1(1'b0), .A2(_u10_n12282 ), .ZN(_u10_n22118 ) );
NAND4_X1 _u10_U10803  ( .A1(_u10_n22115 ), .A2(_u10_n22116 ), .A3(_u10_n22117 ), .A4(_u10_n22118 ), .ZN(_u10_n22100 ) );
NAND2_X1 _u10_U10802  ( .A1(1'b0), .A2(_u10_n12258 ), .ZN(_u10_n22111 ) );
NAND2_X1 _u10_U10801  ( .A1(1'b0), .A2(_u10_n12234 ), .ZN(_u10_n22112 ) );
NAND2_X1 _u10_U10800  ( .A1(1'b0), .A2(_u10_n12210 ), .ZN(_u10_n22113 ) );
NAND2_X1 _u10_U10799  ( .A1(1'b0), .A2(_u10_n12186 ), .ZN(_u10_n22114 ) );
NAND4_X1 _u10_U10798  ( .A1(_u10_n22111 ), .A2(_u10_n22112 ), .A3(_u10_n22113 ), .A4(_u10_n22114 ), .ZN(_u10_n22101 ) );
NAND2_X1 _u10_U10797  ( .A1(1'b0), .A2(_u10_n12161 ), .ZN(_u10_n22107 ) );
NAND2_X1 _u10_U10796  ( .A1(1'b0), .A2(_u10_n12139 ), .ZN(_u10_n22108 ) );
NAND2_X1 _u10_U10795  ( .A1(1'b0), .A2(_u10_n12115 ), .ZN(_u10_n22109 ) );
NAND2_X1 _u10_U10794  ( .A1(1'b0), .A2(_u10_n12091 ), .ZN(_u10_n22110 ) );
NAND4_X1 _u10_U10793  ( .A1(_u10_n22107 ), .A2(_u10_n22108 ), .A3(_u10_n22109 ), .A4(_u10_n22110 ), .ZN(_u10_n22102 ) );
NAND2_X1 _u10_U10792  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n22104 ) );
NAND2_X1 _u10_U10791  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n22105 ) );
NAND2_X1 _u10_U10790  ( .A1(ch0_adr0[28]), .A2(_u10_n12020 ), .ZN(_u10_n22106 ) );
NAND3_X1 _u10_U10789  ( .A1(_u10_n22104 ), .A2(_u10_n22105 ), .A3(_u10_n22106 ), .ZN(_u10_n22103 ) );
NOR4_X1 _u10_U10788  ( .A1(_u10_n22100 ), .A2(_u10_n22101 ), .A3(_u10_n22102 ), .A4(_u10_n22103 ), .ZN(_u10_n22078 ) );
NAND2_X1 _u10_U10787  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n22096 ) );
NAND2_X1 _u10_U10786  ( .A1(1'b0), .A2(_u10_n11969 ), .ZN(_u10_n22097 ) );
NAND2_X1 _u10_U10785  ( .A1(1'b0), .A2(_u10_n11945 ), .ZN(_u10_n22098 ) );
NAND2_X1 _u10_U10784  ( .A1(1'b0), .A2(_u10_n11921 ), .ZN(_u10_n22099 ) );
NAND4_X1 _u10_U10783  ( .A1(_u10_n22096 ), .A2(_u10_n22097 ), .A3(_u10_n22098 ), .A4(_u10_n22099 ), .ZN(_u10_n22080 ) );
NAND2_X1 _u10_U10782  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n22092 ) );
NAND2_X1 _u10_U10781  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n22093 ) );
NAND2_X1 _u10_U10780  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n22094 ) );
NAND2_X1 _u10_U10779  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n22095 ) );
NAND4_X1 _u10_U10778  ( .A1(_u10_n22092 ), .A2(_u10_n22093 ), .A3(_u10_n22094 ), .A4(_u10_n22095 ), .ZN(_u10_n22081 ) );
NAND2_X1 _u10_U10777  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n22088 ) );
NAND2_X1 _u10_U10776  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n22089 ) );
NAND2_X1 _u10_U10775  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n22090 ) );
NAND2_X1 _u10_U10774  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n22091 ) );
NAND4_X1 _u10_U10773  ( .A1(_u10_n22088 ), .A2(_u10_n22089 ), .A3(_u10_n22090 ), .A4(_u10_n22091 ), .ZN(_u10_n22082 ) );
NAND2_X1 _u10_U10772  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n22084 ) );
NAND2_X1 _u10_U10771  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n22085 ) );
NAND2_X1 _u10_U10770  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n22086 ) );
NAND2_X1 _u10_U10769  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n22087 ) );
NAND4_X1 _u10_U10768  ( .A1(_u10_n22084 ), .A2(_u10_n22085 ), .A3(_u10_n22086 ), .A4(_u10_n22087 ), .ZN(_u10_n22083 ) );
NOR4_X1 _u10_U10767  ( .A1(_u10_n22080 ), .A2(_u10_n22081 ), .A3(_u10_n22082 ), .A4(_u10_n22083 ), .ZN(_u10_n22079 ) );
NAND2_X1 _u10_U10766  ( .A1(_u10_n22078 ), .A2(_u10_n22079 ), .ZN(adr0[28]));
NAND2_X1 _u10_U10765  ( .A1(1'b0), .A2(_u10_n12356 ), .ZN(_u10_n22074 ) );
NAND2_X1 _u10_U10764  ( .A1(1'b0), .A2(_u10_n12332 ), .ZN(_u10_n22075 ) );
NAND2_X1 _u10_U10763  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n22076 ) );
NAND2_X1 _u10_U10762  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n22077 ) );
NAND4_X1 _u10_U10761  ( .A1(_u10_n22074 ), .A2(_u10_n22075 ), .A3(_u10_n22076 ), .A4(_u10_n22077 ), .ZN(_u10_n22059 ) );
NAND2_X1 _u10_U10760  ( .A1(1'b0), .A2(_u10_n12260 ), .ZN(_u10_n22070 ) );
NAND2_X1 _u10_U10759  ( .A1(1'b0), .A2(_u10_n12236 ), .ZN(_u10_n22071 ) );
NAND2_X1 _u10_U10758  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n22072 ) );
NAND2_X1 _u10_U10757  ( .A1(1'b0), .A2(_u10_n12188 ), .ZN(_u10_n22073 ) );
NAND4_X1 _u10_U10756  ( .A1(_u10_n22070 ), .A2(_u10_n22071 ), .A3(_u10_n22072 ), .A4(_u10_n22073 ), .ZN(_u10_n22060 ) );
NAND2_X1 _u10_U10755  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n22066 ) );
NAND2_X1 _u10_U10754  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n22067 ) );
NAND2_X1 _u10_U10753  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n22068 ) );
NAND2_X1 _u10_U10752  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n22069 ) );
NAND4_X1 _u10_U10751  ( .A1(_u10_n22066 ), .A2(_u10_n22067 ), .A3(_u10_n22068 ), .A4(_u10_n22069 ), .ZN(_u10_n22061 ) );
NAND2_X1 _u10_U10750  ( .A1(1'b0), .A2(_u10_n12068 ), .ZN(_u10_n22063 ) );
NAND2_X1 _u10_U10749  ( .A1(1'b0), .A2(_u10_n12044 ), .ZN(_u10_n22064 ) );
NAND2_X1 _u10_U10748  ( .A1(ch0_adr0[29]), .A2(_u10_n12020 ), .ZN(_u10_n22065 ) );
NAND3_X1 _u10_U10747  ( .A1(_u10_n22063 ), .A2(_u10_n22064 ), .A3(_u10_n22065 ), .ZN(_u10_n22062 ) );
NOR4_X1 _u10_U10746  ( .A1(_u10_n22059 ), .A2(_u10_n22060 ), .A3(_u10_n22061 ), .A4(_u10_n22062 ), .ZN(_u10_n22037 ) );
NAND2_X1 _u10_U10745  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n22055 ) );
NAND2_X1 _u10_U10744  ( .A1(1'b0), .A2(_u10_n11973 ), .ZN(_u10_n22056 ) );
NAND2_X1 _u10_U10743  ( .A1(1'b0), .A2(_u10_n11949 ), .ZN(_u10_n22057 ) );
NAND2_X1 _u10_U10742  ( .A1(1'b0), .A2(_u10_n11925 ), .ZN(_u10_n22058 ) );
NAND4_X1 _u10_U10741  ( .A1(_u10_n22055 ), .A2(_u10_n22056 ), .A3(_u10_n22057 ), .A4(_u10_n22058 ), .ZN(_u10_n22039 ) );
NAND2_X1 _u10_U10740  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n22051 ) );
NAND2_X1 _u10_U10739  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n22052 ) );
NAND2_X1 _u10_U10738  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n22053 ) );
NAND2_X1 _u10_U10737  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n22054 ) );
NAND4_X1 _u10_U10736  ( .A1(_u10_n22051 ), .A2(_u10_n22052 ), .A3(_u10_n22053 ), .A4(_u10_n22054 ), .ZN(_u10_n22040 ) );
NAND2_X1 _u10_U10735  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n22047 ) );
NAND2_X1 _u10_U10734  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n22048 ) );
NAND2_X1 _u10_U10733  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n22049 ) );
NAND2_X1 _u10_U10732  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n22050 ) );
NAND4_X1 _u10_U10731  ( .A1(_u10_n22047 ), .A2(_u10_n22048 ), .A3(_u10_n22049 ), .A4(_u10_n22050 ), .ZN(_u10_n22041 ) );
NAND2_X1 _u10_U10730  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n22043 ) );
NAND2_X1 _u10_U10729  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n22044 ) );
NAND2_X1 _u10_U10728  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n22045 ) );
NAND2_X1 _u10_U10727  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n22046 ) );
NAND4_X1 _u10_U10726  ( .A1(_u10_n22043 ), .A2(_u10_n22044 ), .A3(_u10_n22045 ), .A4(_u10_n22046 ), .ZN(_u10_n22042 ) );
NOR4_X1 _u10_U10725  ( .A1(_u10_n22039 ), .A2(_u10_n22040 ), .A3(_u10_n22041 ), .A4(_u10_n22042 ), .ZN(_u10_n22038 ) );
NAND2_X1 _u10_U10724  ( .A1(_u10_n22037 ), .A2(_u10_n22038 ), .ZN(adr0[29]));
NAND2_X1 _u10_U10723  ( .A1(1'b0), .A2(_u10_n12354 ), .ZN(_u10_n22033 ) );
NAND2_X1 _u10_U10722  ( .A1(1'b0), .A2(_u10_n12328 ), .ZN(_u10_n22034 ) );
NAND2_X1 _u10_U10721  ( .A1(1'b0), .A2(_u10_n12306 ), .ZN(_u10_n22035 ) );
NAND2_X1 _u10_U10720  ( .A1(1'b0), .A2(_u10_n12282 ), .ZN(_u10_n22036 ) );
NAND4_X1 _u10_U10719  ( .A1(_u10_n22033 ), .A2(_u10_n22034 ), .A3(_u10_n22035 ), .A4(_u10_n22036 ), .ZN(_u10_n22018 ) );
NAND2_X1 _u10_U10718  ( .A1(1'b0), .A2(_u10_n12258 ), .ZN(_u10_n22029 ) );
NAND2_X1 _u10_U10717  ( .A1(1'b0), .A2(_u10_n12234 ), .ZN(_u10_n22030 ) );
NAND2_X1 _u10_U10716  ( .A1(1'b0), .A2(_u10_n12211 ), .ZN(_u10_n22031 ) );
NAND2_X1 _u10_U10715  ( .A1(1'b0), .A2(_u10_n12186 ), .ZN(_u10_n22032 ) );
NAND4_X1 _u10_U10714  ( .A1(_u10_n22029 ), .A2(_u10_n22030 ), .A3(_u10_n22031 ), .A4(_u10_n22032 ), .ZN(_u10_n22019 ) );
NAND2_X1 _u10_U10713  ( .A1(1'b0), .A2(_u10_n12159 ), .ZN(_u10_n22025 ) );
NAND2_X1 _u10_U10712  ( .A1(1'b0), .A2(_u10_n12135 ), .ZN(_u10_n22026 ) );
NAND2_X1 _u10_U10711  ( .A1(1'b0), .A2(_u10_n12111 ), .ZN(_u10_n22027 ) );
NAND2_X1 _u10_U10710  ( .A1(1'b0), .A2(_u10_n12087 ), .ZN(_u10_n22028 ) );
NAND4_X1 _u10_U10709  ( .A1(_u10_n22025 ), .A2(_u10_n22026 ), .A3(_u10_n22027 ), .A4(_u10_n22028 ), .ZN(_u10_n22020 ) );
NAND2_X1 _u10_U10708  ( .A1(1'b0), .A2(_u10_n12063 ), .ZN(_u10_n22022 ) );
NAND2_X1 _u10_U10707  ( .A1(1'b0), .A2(_u10_n12039 ), .ZN(_u10_n22023 ) );
NAND2_X1 _u10_U10706  ( .A1(ch0_adr0[2]), .A2(_u10_n12020 ), .ZN(_u10_n22024 ) );
NAND3_X1 _u10_U10705  ( .A1(_u10_n22022 ), .A2(_u10_n22023 ), .A3(_u10_n22024 ), .ZN(_u10_n22021 ) );
NOR4_X1 _u10_U10704  ( .A1(_u10_n22018 ), .A2(_u10_n22019 ), .A3(_u10_n22020 ), .A4(_u10_n22021 ), .ZN(_u10_n21996 ) );
NAND2_X1 _u10_U10703  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n22014 ) );
NAND2_X1 _u10_U10702  ( .A1(1'b0), .A2(_u10_n11972 ), .ZN(_u10_n22015 ) );
NAND2_X1 _u10_U10701  ( .A1(1'b0), .A2(_u10_n11948 ), .ZN(_u10_n22016 ) );
NAND2_X1 _u10_U10700  ( .A1(1'b0), .A2(_u10_n11924 ), .ZN(_u10_n22017 ) );
NAND4_X1 _u10_U10699  ( .A1(_u10_n22014 ), .A2(_u10_n22015 ), .A3(_u10_n22016 ), .A4(_u10_n22017 ), .ZN(_u10_n21998 ) );
NAND2_X1 _u10_U10698  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n22010 ) );
NAND2_X1 _u10_U10697  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n22011 ) );
NAND2_X1 _u10_U10696  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n22012 ) );
NAND2_X1 _u10_U10695  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n22013 ) );
NAND4_X1 _u10_U10694  ( .A1(_u10_n22010 ), .A2(_u10_n22011 ), .A3(_u10_n22012 ), .A4(_u10_n22013 ), .ZN(_u10_n21999 ) );
NAND2_X1 _u10_U10693  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n22006 ) );
NAND2_X1 _u10_U10692  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n22007 ) );
NAND2_X1 _u10_U10691  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n22008 ) );
NAND2_X1 _u10_U10690  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n22009 ) );
NAND4_X1 _u10_U10689  ( .A1(_u10_n22006 ), .A2(_u10_n22007 ), .A3(_u10_n22008 ), .A4(_u10_n22009 ), .ZN(_u10_n22000 ) );
NAND2_X1 _u10_U10688  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n22002 ) );
NAND2_X1 _u10_U10687  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n22003 ) );
NAND2_X1 _u10_U10686  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n22004 ) );
NAND2_X1 _u10_U10685  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n22005 ) );
NAND4_X1 _u10_U10684  ( .A1(_u10_n22002 ), .A2(_u10_n22003 ), .A3(_u10_n22004 ), .A4(_u10_n22005 ), .ZN(_u10_n22001 ) );
NOR4_X1 _u10_U10683  ( .A1(_u10_n21998 ), .A2(_u10_n21999 ), .A3(_u10_n22000 ), .A4(_u10_n22001 ), .ZN(_u10_n21997 ) );
NAND2_X1 _u10_U10682  ( .A1(_u10_n21996 ), .A2(_u10_n21997 ), .ZN(adr0[2]));
NAND2_X1 _u10_U10681  ( .A1(1'b0), .A2(_u10_n12430 ), .ZN(_u10_n21992 ) );
NAND2_X1 _u10_U10680  ( .A1(1'b0), .A2(_u10_n12429 ), .ZN(_u10_n21993 ) );
NAND2_X1 _u10_U10679  ( .A1(1'b0), .A2(_u10_n12428 ), .ZN(_u10_n21994 ) );
NAND2_X1 _u10_U10678  ( .A1(1'b0), .A2(_u10_n12427 ), .ZN(_u10_n21995 ) );
NAND4_X1 _u10_U10677  ( .A1(_u10_n21992 ), .A2(_u10_n21993 ), .A3(_u10_n21994 ), .A4(_u10_n21995 ), .ZN(_u10_n21977 ) );
NAND2_X1 _u10_U10676  ( .A1(1'b0), .A2(_u10_n12422 ), .ZN(_u10_n21988 ) );
NAND2_X1 _u10_U10675  ( .A1(1'b0), .A2(_u10_n12421 ), .ZN(_u10_n21989 ) );
NAND2_X1 _u10_U10674  ( .A1(1'b0), .A2(_u10_n12420 ), .ZN(_u10_n21990 ) );
NAND2_X1 _u10_U10673  ( .A1(1'b0), .A2(_u10_n12419 ), .ZN(_u10_n21991 ) );
NAND4_X1 _u10_U10672  ( .A1(_u10_n21988 ), .A2(_u10_n21989 ), .A3(_u10_n21990 ), .A4(_u10_n21991 ), .ZN(_u10_n21978 ) );
NAND2_X1 _u10_U10671  ( .A1(1'b0), .A2(_u10_n12163 ), .ZN(_u10_n21984 ) );
NAND2_X1 _u10_U10670  ( .A1(1'b0), .A2(_u10_n12413 ), .ZN(_u10_n21985 ) );
NAND2_X1 _u10_U10669  ( .A1(1'b0), .A2(_u10_n12412 ), .ZN(_u10_n21986 ) );
NAND2_X1 _u10_U10668  ( .A1(1'b0), .A2(_u10_n12411 ), .ZN(_u10_n21987 ) );
NAND4_X1 _u10_U10667  ( .A1(_u10_n21984 ), .A2(_u10_n21985 ), .A3(_u10_n21986 ), .A4(_u10_n21987 ), .ZN(_u10_n21979 ) );
NAND2_X1 _u10_U10666  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n21981 ) );
NAND2_X1 _u10_U10665  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n21982 ) );
NAND2_X1 _u10_U10664  ( .A1(ch0_adr0[30]), .A2(_u10_n12001 ), .ZN(_u10_n21983 ) );
NAND3_X1 _u10_U10663  ( .A1(_u10_n21981 ), .A2(_u10_n21982 ), .A3(_u10_n21983 ), .ZN(_u10_n21980 ) );
NOR4_X1 _u10_U10662  ( .A1(_u10_n21977 ), .A2(_u10_n21978 ), .A3(_u10_n21979 ), .A4(_u10_n21980 ), .ZN(_u10_n21955 ) );
NAND2_X1 _u10_U10661  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n21973 ) );
NAND2_X1 _u10_U10660  ( .A1(1'b0), .A2(_u10_n11975 ), .ZN(_u10_n21974 ) );
NAND2_X1 _u10_U10659  ( .A1(1'b0), .A2(_u10_n11951 ), .ZN(_u10_n21975 ) );
NAND2_X1 _u10_U10658  ( .A1(1'b0), .A2(_u10_n11927 ), .ZN(_u10_n21976 ) );
NAND4_X1 _u10_U10657  ( .A1(_u10_n21973 ), .A2(_u10_n21974 ), .A3(_u10_n21975 ), .A4(_u10_n21976 ), .ZN(_u10_n21957 ) );
NAND2_X1 _u10_U10656  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n21969 ) );
NAND2_X1 _u10_U10655  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n21970 ) );
NAND2_X1 _u10_U10654  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n21971 ) );
NAND2_X1 _u10_U10653  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n21972 ) );
NAND4_X1 _u10_U10652  ( .A1(_u10_n21969 ), .A2(_u10_n21970 ), .A3(_u10_n21971 ), .A4(_u10_n21972 ), .ZN(_u10_n21958 ) );
NAND2_X1 _u10_U10651  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n21965 ) );
NAND2_X1 _u10_U10650  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n21966 ) );
NAND2_X1 _u10_U10649  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n21967 ) );
NAND2_X1 _u10_U10648  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n21968 ) );
NAND4_X1 _u10_U10647  ( .A1(_u10_n21965 ), .A2(_u10_n21966 ), .A3(_u10_n21967 ), .A4(_u10_n21968 ), .ZN(_u10_n21959 ) );
NAND2_X1 _u10_U10646  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n21961 ) );
NAND2_X1 _u10_U10645  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n21962 ) );
NAND2_X1 _u10_U10644  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n21963 ) );
NAND2_X1 _u10_U10643  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n21964 ) );
NAND4_X1 _u10_U10642  ( .A1(_u10_n21961 ), .A2(_u10_n21962 ), .A3(_u10_n21963 ), .A4(_u10_n21964 ), .ZN(_u10_n21960 ) );
NOR4_X1 _u10_U10641  ( .A1(_u10_n21957 ), .A2(_u10_n21958 ), .A3(_u10_n21959 ), .A4(_u10_n21960 ), .ZN(_u10_n21956 ) );
NAND2_X1 _u10_U10640  ( .A1(_u10_n21955 ), .A2(_u10_n21956 ), .ZN(adr0[30]));
NAND2_X1 _u10_U10639  ( .A1(1'b0), .A2(_u10_n12430 ), .ZN(_u10_n21951 ) );
NAND2_X1 _u10_U10638  ( .A1(1'b0), .A2(_u10_n12429 ), .ZN(_u10_n21952 ) );
NAND2_X1 _u10_U10637  ( .A1(1'b0), .A2(_u10_n12303 ), .ZN(_u10_n21953 ) );
NAND2_X1 _u10_U10636  ( .A1(1'b0), .A2(_u10_n12279 ), .ZN(_u10_n21954 ) );
NAND4_X1 _u10_U10635  ( .A1(_u10_n21951 ), .A2(_u10_n21952 ), .A3(_u10_n21953 ), .A4(_u10_n21954 ), .ZN(_u10_n21936 ) );
NAND2_X1 _u10_U10634  ( .A1(1'b0), .A2(_u10_n12422 ), .ZN(_u10_n21947 ) );
NAND2_X1 _u10_U10633  ( .A1(1'b0), .A2(_u10_n12421 ), .ZN(_u10_n21948 ) );
NAND2_X1 _u10_U10632  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n21949 ) );
NAND2_X1 _u10_U10631  ( .A1(1'b0), .A2(_u10_n12419 ), .ZN(_u10_n21950 ) );
NAND4_X1 _u10_U10630  ( .A1(_u10_n21947 ), .A2(_u10_n21948 ), .A3(_u10_n21949 ), .A4(_u10_n21950 ), .ZN(_u10_n21937 ) );
NAND2_X1 _u10_U10629  ( .A1(1'b0), .A2(_u10_n12414 ), .ZN(_u10_n21943 ) );
NAND2_X1 _u10_U10628  ( .A1(1'b0), .A2(_u10_n12136 ), .ZN(_u10_n21944 ) );
NAND2_X1 _u10_U10627  ( .A1(1'b0), .A2(_u10_n12112 ), .ZN(_u10_n21945 ) );
NAND2_X1 _u10_U10626  ( .A1(1'b0), .A2(_u10_n12088 ), .ZN(_u10_n21946 ) );
NAND4_X1 _u10_U10625  ( .A1(_u10_n21943 ), .A2(_u10_n21944 ), .A3(_u10_n21945 ), .A4(_u10_n21946 ), .ZN(_u10_n21938 ) );
NAND2_X1 _u10_U10624  ( .A1(1'b0), .A2(_u10_n12063 ), .ZN(_u10_n21940 ) );
NAND2_X1 _u10_U10623  ( .A1(1'b0), .A2(_u10_n12039 ), .ZN(_u10_n21941 ) );
NAND2_X1 _u10_U10622  ( .A1(ch0_adr0[31]), .A2(_u10_n12001 ), .ZN(_u10_n21942 ) );
NAND3_X1 _u10_U10621  ( .A1(_u10_n21940 ), .A2(_u10_n21941 ), .A3(_u10_n21942 ), .ZN(_u10_n21939 ) );
NOR4_X1 _u10_U10620  ( .A1(_u10_n21936 ), .A2(_u10_n21937 ), .A3(_u10_n21938 ), .A4(_u10_n21939 ), .ZN(_u10_n21914 ) );
NAND2_X1 _u10_U10619  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n21932 ) );
NAND2_X1 _u10_U10618  ( .A1(1'b0), .A2(_u10_n11971 ), .ZN(_u10_n21933 ) );
NAND2_X1 _u10_U10617  ( .A1(1'b0), .A2(_u10_n11947 ), .ZN(_u10_n21934 ) );
NAND2_X1 _u10_U10616  ( .A1(1'b0), .A2(_u10_n11923 ), .ZN(_u10_n21935 ) );
NAND4_X1 _u10_U10615  ( .A1(_u10_n21932 ), .A2(_u10_n21933 ), .A3(_u10_n21934 ), .A4(_u10_n21935 ), .ZN(_u10_n21916 ) );
NAND2_X1 _u10_U10614  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n21928 ) );
NAND2_X1 _u10_U10613  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n21929 ) );
NAND2_X1 _u10_U10612  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n21930 ) );
NAND2_X1 _u10_U10611  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n21931 ) );
NAND4_X1 _u10_U10610  ( .A1(_u10_n21928 ), .A2(_u10_n21929 ), .A3(_u10_n21930 ), .A4(_u10_n21931 ), .ZN(_u10_n21917 ) );
NAND2_X1 _u10_U10609  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n21924 ) );
NAND2_X1 _u10_U10608  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n21925 ) );
NAND2_X1 _u10_U10607  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n21926 ) );
NAND2_X1 _u10_U10606  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n21927 ) );
NAND4_X1 _u10_U10605  ( .A1(_u10_n21924 ), .A2(_u10_n21925 ), .A3(_u10_n21926 ), .A4(_u10_n21927 ), .ZN(_u10_n21918 ) );
NAND2_X1 _u10_U10604  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n21920 ) );
NAND2_X1 _u10_U10603  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n21921 ) );
NAND2_X1 _u10_U10602  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n21922 ) );
NAND2_X1 _u10_U10601  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n21923 ) );
NAND4_X1 _u10_U10600  ( .A1(_u10_n21920 ), .A2(_u10_n21921 ), .A3(_u10_n21922 ), .A4(_u10_n21923 ), .ZN(_u10_n21919 ) );
NOR4_X1 _u10_U10599  ( .A1(_u10_n21916 ), .A2(_u10_n21917 ), .A3(_u10_n21918 ), .A4(_u10_n21919 ), .ZN(_u10_n21915 ) );
NAND2_X1 _u10_U10598  ( .A1(_u10_n21914 ), .A2(_u10_n21915 ), .ZN(adr0[31]));
NAND2_X1 _u10_U10597  ( .A1(1'b0), .A2(_u10_n12352 ), .ZN(_u10_n21910 ) );
NAND2_X1 _u10_U10596  ( .A1(1'b0), .A2(_u10_n12328 ), .ZN(_u10_n21911 ) );
NAND2_X1 _u10_U10595  ( .A1(1'b0), .A2(_u10_n12306 ), .ZN(_u10_n21912 ) );
NAND2_X1 _u10_U10594  ( .A1(1'b0), .A2(_u10_n12282 ), .ZN(_u10_n21913 ) );
NAND4_X1 _u10_U10593  ( .A1(_u10_n21910 ), .A2(_u10_n21911 ), .A3(_u10_n21912 ), .A4(_u10_n21913 ), .ZN(_u10_n21895 ) );
NAND2_X1 _u10_U10592  ( .A1(1'b0), .A2(_u10_n12256 ), .ZN(_u10_n21906 ) );
NAND2_X1 _u10_U10591  ( .A1(1'b0), .A2(_u10_n12232 ), .ZN(_u10_n21907 ) );
NAND2_X1 _u10_U10590  ( .A1(1'b0), .A2(_u10_n12206 ), .ZN(_u10_n21908 ) );
NAND2_X1 _u10_U10589  ( .A1(1'b0), .A2(_u10_n12184 ), .ZN(_u10_n21909 ) );
NAND4_X1 _u10_U10588  ( .A1(_u10_n21906 ), .A2(_u10_n21907 ), .A3(_u10_n21908 ), .A4(_u10_n21909 ), .ZN(_u10_n21896 ) );
NAND2_X1 _u10_U10587  ( .A1(1'b0), .A2(_u10_n12160 ), .ZN(_u10_n21902 ) );
NAND2_X1 _u10_U10586  ( .A1(1'b0), .A2(_u10_n12138 ), .ZN(_u10_n21903 ) );
NAND2_X1 _u10_U10585  ( .A1(1'b0), .A2(_u10_n12114 ), .ZN(_u10_n21904 ) );
NAND2_X1 _u10_U10584  ( .A1(1'b0), .A2(_u10_n12090 ), .ZN(_u10_n21905 ) );
NAND4_X1 _u10_U10583  ( .A1(_u10_n21902 ), .A2(_u10_n21903 ), .A3(_u10_n21904 ), .A4(_u10_n21905 ), .ZN(_u10_n21897 ) );
NAND2_X1 _u10_U10582  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n21899 ) );
NAND2_X1 _u10_U10581  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n21900 ) );
NAND2_X1 _u10_U10580  ( .A1(ch0_adr0[3]), .A2(_u10_n12001 ), .ZN(_u10_n21901 ) );
NAND3_X1 _u10_U10579  ( .A1(_u10_n21899 ), .A2(_u10_n21900 ), .A3(_u10_n21901 ), .ZN(_u10_n21898 ) );
NOR4_X1 _u10_U10578  ( .A1(_u10_n21895 ), .A2(_u10_n21896 ), .A3(_u10_n21897 ), .A4(_u10_n21898 ), .ZN(_u10_n21873 ) );
NAND2_X1 _u10_U10577  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n21891 ) );
NAND2_X1 _u10_U10576  ( .A1(1'b0), .A2(_u10_n11970 ), .ZN(_u10_n21892 ) );
NAND2_X1 _u10_U10575  ( .A1(1'b0), .A2(_u10_n11946 ), .ZN(_u10_n21893 ) );
NAND2_X1 _u10_U10574  ( .A1(1'b0), .A2(_u10_n11922 ), .ZN(_u10_n21894 ) );
NAND4_X1 _u10_U10573  ( .A1(_u10_n21891 ), .A2(_u10_n21892 ), .A3(_u10_n21893 ), .A4(_u10_n21894 ), .ZN(_u10_n21875 ) );
NAND2_X1 _u10_U10572  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n21887 ) );
NAND2_X1 _u10_U10571  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n21888 ) );
NAND2_X1 _u10_U10570  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n21889 ) );
NAND2_X1 _u10_U10569  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n21890 ) );
NAND4_X1 _u10_U10568  ( .A1(_u10_n21887 ), .A2(_u10_n21888 ), .A3(_u10_n21889 ), .A4(_u10_n21890 ), .ZN(_u10_n21876 ) );
NAND2_X1 _u10_U10567  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n21883 ) );
NAND2_X1 _u10_U10566  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n21884 ) );
NAND2_X1 _u10_U10565  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n21885 ) );
NAND2_X1 _u10_U10564  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n21886 ) );
NAND4_X1 _u10_U10563  ( .A1(_u10_n21883 ), .A2(_u10_n21884 ), .A3(_u10_n21885 ), .A4(_u10_n21886 ), .ZN(_u10_n21877 ) );
NAND2_X1 _u10_U10562  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n21879 ) );
NAND2_X1 _u10_U10561  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n21880 ) );
NAND2_X1 _u10_U10560  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n21881 ) );
NAND2_X1 _u10_U10559  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n21882 ) );
NAND4_X1 _u10_U10558  ( .A1(_u10_n21879 ), .A2(_u10_n21880 ), .A3(_u10_n21881 ), .A4(_u10_n21882 ), .ZN(_u10_n21878 ) );
NOR4_X1 _u10_U10557  ( .A1(_u10_n21875 ), .A2(_u10_n21876 ), .A3(_u10_n21877 ), .A4(_u10_n21878 ), .ZN(_u10_n21874 ) );
NAND2_X1 _u10_U10556  ( .A1(_u10_n21873 ), .A2(_u10_n21874 ), .ZN(adr0[3]));
NAND2_X1 _u10_U10555  ( .A1(1'b0), .A2(_u10_n12356 ), .ZN(_u10_n21869 ) );
NAND2_X1 _u10_U10554  ( .A1(1'b0), .A2(_u10_n12332 ), .ZN(_u10_n21870 ) );
NAND2_X1 _u10_U10553  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n21871 ) );
NAND2_X1 _u10_U10552  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n21872 ) );
NAND4_X1 _u10_U10551  ( .A1(_u10_n21869 ), .A2(_u10_n21870 ), .A3(_u10_n21871 ), .A4(_u10_n21872 ), .ZN(_u10_n21854 ) );
NAND2_X1 _u10_U10550  ( .A1(1'b0), .A2(_u10_n12260 ), .ZN(_u10_n21865 ) );
NAND2_X1 _u10_U10549  ( .A1(1'b0), .A2(_u10_n12236 ), .ZN(_u10_n21866 ) );
NAND2_X1 _u10_U10548  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n21867 ) );
NAND2_X1 _u10_U10547  ( .A1(1'b0), .A2(_u10_n12188 ), .ZN(_u10_n21868 ) );
NAND4_X1 _u10_U10546  ( .A1(_u10_n21865 ), .A2(_u10_n21866 ), .A3(_u10_n21867 ), .A4(_u10_n21868 ), .ZN(_u10_n21855 ) );
NAND2_X1 _u10_U10545  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n21861 ) );
NAND2_X1 _u10_U10544  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n21862 ) );
NAND2_X1 _u10_U10543  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n21863 ) );
NAND2_X1 _u10_U10542  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n21864 ) );
NAND4_X1 _u10_U10541  ( .A1(_u10_n21861 ), .A2(_u10_n21862 ), .A3(_u10_n21863 ), .A4(_u10_n21864 ), .ZN(_u10_n21856 ) );
NAND2_X1 _u10_U10540  ( .A1(1'b0), .A2(_u10_n12068 ), .ZN(_u10_n21858 ) );
NAND2_X1 _u10_U10539  ( .A1(1'b0), .A2(_u10_n12044 ), .ZN(_u10_n21859 ) );
NAND2_X1 _u10_U10538  ( .A1(ch0_adr0[4]), .A2(_u10_n12001 ), .ZN(_u10_n21860 ) );
NAND3_X1 _u10_U10537  ( .A1(_u10_n21858 ), .A2(_u10_n21859 ), .A3(_u10_n21860 ), .ZN(_u10_n21857 ) );
NOR4_X1 _u10_U10536  ( .A1(_u10_n21854 ), .A2(_u10_n21855 ), .A3(_u10_n21856 ), .A4(_u10_n21857 ), .ZN(_u10_n21832 ) );
NAND2_X1 _u10_U10535  ( .A1(1'b0), .A2(_u10_n11984 ), .ZN(_u10_n21850 ) );
NAND2_X1 _u10_U10534  ( .A1(1'b0), .A2(_u10_n11973 ), .ZN(_u10_n21851 ) );
NAND2_X1 _u10_U10533  ( .A1(1'b0), .A2(_u10_n11949 ), .ZN(_u10_n21852 ) );
NAND2_X1 _u10_U10532  ( .A1(1'b0), .A2(_u10_n11925 ), .ZN(_u10_n21853 ) );
NAND4_X1 _u10_U10531  ( .A1(_u10_n21850 ), .A2(_u10_n21851 ), .A3(_u10_n21852 ), .A4(_u10_n21853 ), .ZN(_u10_n21834 ) );
NAND2_X1 _u10_U10530  ( .A1(1'b0), .A2(_u10_n11888 ), .ZN(_u10_n21846 ) );
NAND2_X1 _u10_U10529  ( .A1(1'b0), .A2(_u10_n11864 ), .ZN(_u10_n21847 ) );
NAND2_X1 _u10_U10528  ( .A1(1'b0), .A2(_u10_n11840 ), .ZN(_u10_n21848 ) );
NAND2_X1 _u10_U10527  ( .A1(1'b0), .A2(_u10_n11816 ), .ZN(_u10_n21849 ) );
NAND4_X1 _u10_U10526  ( .A1(_u10_n21846 ), .A2(_u10_n21847 ), .A3(_u10_n21848 ), .A4(_u10_n21849 ), .ZN(_u10_n21835 ) );
NAND2_X1 _u10_U10525  ( .A1(1'b0), .A2(_u10_n11792 ), .ZN(_u10_n21842 ) );
NAND2_X1 _u10_U10524  ( .A1(1'b0), .A2(_u10_n11768 ), .ZN(_u10_n21843 ) );
NAND2_X1 _u10_U10523  ( .A1(1'b0), .A2(_u10_n11744 ), .ZN(_u10_n21844 ) );
NAND2_X1 _u10_U10522  ( .A1(1'b0), .A2(_u10_n11720 ), .ZN(_u10_n21845 ) );
NAND4_X1 _u10_U10521  ( .A1(_u10_n21842 ), .A2(_u10_n21843 ), .A3(_u10_n21844 ), .A4(_u10_n21845 ), .ZN(_u10_n21836 ) );
NAND2_X1 _u10_U10520  ( .A1(1'b0), .A2(_u10_n11696 ), .ZN(_u10_n21838 ) );
NAND2_X1 _u10_U10519  ( .A1(1'b0), .A2(_u10_n11672 ), .ZN(_u10_n21839 ) );
NAND2_X1 _u10_U10518  ( .A1(1'b0), .A2(_u10_n11648 ), .ZN(_u10_n21840 ) );
NAND2_X1 _u10_U10517  ( .A1(1'b0), .A2(_u10_n11624 ), .ZN(_u10_n21841 ) );
NAND4_X1 _u10_U10516  ( .A1(_u10_n21838 ), .A2(_u10_n21839 ), .A3(_u10_n21840 ), .A4(_u10_n21841 ), .ZN(_u10_n21837 ) );
NOR4_X1 _u10_U10515  ( .A1(_u10_n21834 ), .A2(_u10_n21835 ), .A3(_u10_n21836 ), .A4(_u10_n21837 ), .ZN(_u10_n21833 ) );
NAND2_X1 _u10_U10514  ( .A1(_u10_n21832 ), .A2(_u10_n21833 ), .ZN(adr0[4]));
NAND2_X1 _u10_U10513  ( .A1(1'b0), .A2(_u10_n12354 ), .ZN(_u10_n21828 ) );
NAND2_X1 _u10_U10512  ( .A1(1'b0), .A2(_u10_n12331 ), .ZN(_u10_n21829 ) );
NAND2_X1 _u10_U10511  ( .A1(1'b0), .A2(_u10_n12307 ), .ZN(_u10_n21830 ) );
NAND2_X1 _u10_U10510  ( .A1(1'b0), .A2(_u10_n12283 ), .ZN(_u10_n21831 ) );
NAND4_X1 _u10_U10509  ( .A1(_u10_n21828 ), .A2(_u10_n21829 ), .A3(_u10_n21830 ), .A4(_u10_n21831 ), .ZN(_u10_n21813 ) );
NAND2_X1 _u10_U10508  ( .A1(1'b0), .A2(_u10_n12258 ), .ZN(_u10_n21824 ) );
NAND2_X1 _u10_U10507  ( .A1(1'b0), .A2(_u10_n12234 ), .ZN(_u10_n21825 ) );
NAND2_X1 _u10_U10506  ( .A1(1'b0), .A2(_u10_n12209 ), .ZN(_u10_n21826 ) );
NAND2_X1 _u10_U10505  ( .A1(1'b0), .A2(_u10_n12186 ), .ZN(_u10_n21827 ) );
NAND4_X1 _u10_U10504  ( .A1(_u10_n21824 ), .A2(_u10_n21825 ), .A3(_u10_n21826 ), .A4(_u10_n21827 ), .ZN(_u10_n21814 ) );
NAND2_X1 _u10_U10503  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n21820 ) );
NAND2_X1 _u10_U10502  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n21821 ) );
NAND2_X1 _u10_U10501  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n21822 ) );
NAND2_X1 _u10_U10500  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n21823 ) );
NAND4_X1 _u10_U10499  ( .A1(_u10_n21820 ), .A2(_u10_n21821 ), .A3(_u10_n21822 ), .A4(_u10_n21823 ), .ZN(_u10_n21815 ) );
NAND2_X1 _u10_U10498  ( .A1(1'b0), .A2(_u10_n12065 ), .ZN(_u10_n21817 ) );
NAND2_X1 _u10_U10497  ( .A1(1'b0), .A2(_u10_n12041 ), .ZN(_u10_n21818 ) );
NAND2_X1 _u10_U10496  ( .A1(ch0_adr0[5]), .A2(_u10_n12001 ), .ZN(_u10_n21819 ) );
NAND3_X1 _u10_U10495  ( .A1(_u10_n21817 ), .A2(_u10_n21818 ), .A3(_u10_n21819 ), .ZN(_u10_n21816 ) );
NOR4_X1 _u10_U10494  ( .A1(_u10_n21813 ), .A2(_u10_n21814 ), .A3(_u10_n21815 ), .A4(_u10_n21816 ), .ZN(_u10_n21791 ) );
NAND2_X1 _u10_U10493  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21809 ) );
NAND2_X1 _u10_U10492  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21810 ) );
NAND2_X1 _u10_U10491  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21811 ) );
NAND2_X1 _u10_U10490  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21812 ) );
NAND4_X1 _u10_U10489  ( .A1(_u10_n21809 ), .A2(_u10_n21810 ), .A3(_u10_n21811 ), .A4(_u10_n21812 ), .ZN(_u10_n21793 ) );
NAND2_X1 _u10_U10488  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21805 ) );
NAND2_X1 _u10_U10487  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21806 ) );
NAND2_X1 _u10_U10486  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21807 ) );
NAND2_X1 _u10_U10485  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21808 ) );
NAND4_X1 _u10_U10484  ( .A1(_u10_n21805 ), .A2(_u10_n21806 ), .A3(_u10_n21807 ), .A4(_u10_n21808 ), .ZN(_u10_n21794 ) );
NAND2_X1 _u10_U10483  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21801 ) );
NAND2_X1 _u10_U10482  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21802 ) );
NAND2_X1 _u10_U10481  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21803 ) );
NAND2_X1 _u10_U10480  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21804 ) );
NAND4_X1 _u10_U10479  ( .A1(_u10_n21801 ), .A2(_u10_n21802 ), .A3(_u10_n21803 ), .A4(_u10_n21804 ), .ZN(_u10_n21795 ) );
NAND2_X1 _u10_U10478  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21797 ) );
NAND2_X1 _u10_U10477  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21798 ) );
NAND2_X1 _u10_U10476  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21799 ) );
NAND2_X1 _u10_U10475  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21800 ) );
NAND4_X1 _u10_U10474  ( .A1(_u10_n21797 ), .A2(_u10_n21798 ), .A3(_u10_n21799 ), .A4(_u10_n21800 ), .ZN(_u10_n21796 ) );
NOR4_X1 _u10_U10473  ( .A1(_u10_n21793 ), .A2(_u10_n21794 ), .A3(_u10_n21795 ), .A4(_u10_n21796 ), .ZN(_u10_n21792 ) );
NAND2_X1 _u10_U10472  ( .A1(_u10_n21791 ), .A2(_u10_n21792 ), .ZN(adr0[5]));
NAND2_X1 _u10_U10471  ( .A1(1'b0), .A2(_u10_n12355 ), .ZN(_u10_n21787 ) );
NAND2_X1 _u10_U10470  ( .A1(1'b0), .A2(_u10_n12330 ), .ZN(_u10_n21788 ) );
NAND2_X1 _u10_U10469  ( .A1(1'b0), .A2(_u10_n12306 ), .ZN(_u10_n21789 ) );
NAND2_X1 _u10_U10468  ( .A1(1'b0), .A2(_u10_n12282 ), .ZN(_u10_n21790 ) );
NAND4_X1 _u10_U10467  ( .A1(_u10_n21787 ), .A2(_u10_n21788 ), .A3(_u10_n21789 ), .A4(_u10_n21790 ), .ZN(_u10_n21772 ) );
NAND2_X1 _u10_U10466  ( .A1(1'b0), .A2(_u10_n12259 ), .ZN(_u10_n21783 ) );
NAND2_X1 _u10_U10465  ( .A1(1'b0), .A2(_u10_n12235 ), .ZN(_u10_n21784 ) );
NAND2_X1 _u10_U10464  ( .A1(1'b0), .A2(_u10_n12211 ), .ZN(_u10_n21785 ) );
NAND2_X1 _u10_U10463  ( .A1(1'b0), .A2(_u10_n12187 ), .ZN(_u10_n21786 ) );
NAND4_X1 _u10_U10462  ( .A1(_u10_n21783 ), .A2(_u10_n21784 ), .A3(_u10_n21785 ), .A4(_u10_n21786 ), .ZN(_u10_n21773 ) );
NAND2_X1 _u10_U10461  ( .A1(1'b0), .A2(_u10_n12161 ), .ZN(_u10_n21779 ) );
NAND2_X1 _u10_U10460  ( .A1(1'b0), .A2(_u10_n12137 ), .ZN(_u10_n21780 ) );
NAND2_X1 _u10_U10459  ( .A1(1'b0), .A2(_u10_n12113 ), .ZN(_u10_n21781 ) );
NAND2_X1 _u10_U10458  ( .A1(1'b0), .A2(_u10_n12089 ), .ZN(_u10_n21782 ) );
NAND4_X1 _u10_U10457  ( .A1(_u10_n21779 ), .A2(_u10_n21780 ), .A3(_u10_n21781 ), .A4(_u10_n21782 ), .ZN(_u10_n21774 ) );
NAND2_X1 _u10_U10456  ( .A1(1'b0), .A2(_u10_n12067 ), .ZN(_u10_n21776 ) );
NAND2_X1 _u10_U10455  ( .A1(1'b0), .A2(_u10_n12043 ), .ZN(_u10_n21777 ) );
NAND2_X1 _u10_U10454  ( .A1(ch0_adr0[6]), .A2(_u10_n12001 ), .ZN(_u10_n21778 ) );
NAND3_X1 _u10_U10453  ( .A1(_u10_n21776 ), .A2(_u10_n21777 ), .A3(_u10_n21778 ), .ZN(_u10_n21775 ) );
NOR4_X1 _u10_U10452  ( .A1(_u10_n21772 ), .A2(_u10_n21773 ), .A3(_u10_n21774 ), .A4(_u10_n21775 ), .ZN(_u10_n21750 ) );
NAND2_X1 _u10_U10451  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21768 ) );
NAND2_X1 _u10_U10450  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21769 ) );
NAND2_X1 _u10_U10449  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21770 ) );
NAND2_X1 _u10_U10448  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21771 ) );
NAND4_X1 _u10_U10447  ( .A1(_u10_n21768 ), .A2(_u10_n21769 ), .A3(_u10_n21770 ), .A4(_u10_n21771 ), .ZN(_u10_n21752 ) );
NAND2_X1 _u10_U10446  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21764 ) );
NAND2_X1 _u10_U10445  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21765 ) );
NAND2_X1 _u10_U10444  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21766 ) );
NAND2_X1 _u10_U10443  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21767 ) );
NAND4_X1 _u10_U10442  ( .A1(_u10_n21764 ), .A2(_u10_n21765 ), .A3(_u10_n21766 ), .A4(_u10_n21767 ), .ZN(_u10_n21753 ) );
NAND2_X1 _u10_U10441  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21760 ) );
NAND2_X1 _u10_U10440  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21761 ) );
NAND2_X1 _u10_U10439  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21762 ) );
NAND2_X1 _u10_U10438  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21763 ) );
NAND4_X1 _u10_U10437  ( .A1(_u10_n21760 ), .A2(_u10_n21761 ), .A3(_u10_n21762 ), .A4(_u10_n21763 ), .ZN(_u10_n21754 ) );
NAND2_X1 _u10_U10436  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21756 ) );
NAND2_X1 _u10_U10435  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21757 ) );
NAND2_X1 _u10_U10434  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21758 ) );
NAND2_X1 _u10_U10433  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21759 ) );
NAND4_X1 _u10_U10432  ( .A1(_u10_n21756 ), .A2(_u10_n21757 ), .A3(_u10_n21758 ), .A4(_u10_n21759 ), .ZN(_u10_n21755 ) );
NOR4_X1 _u10_U10431  ( .A1(_u10_n21752 ), .A2(_u10_n21753 ), .A3(_u10_n21754 ), .A4(_u10_n21755 ), .ZN(_u10_n21751 ) );
NAND2_X1 _u10_U10430  ( .A1(_u10_n21750 ), .A2(_u10_n21751 ), .ZN(adr0[6]));
NAND2_X1 _u10_U10429  ( .A1(1'b0), .A2(_u10_n12354 ), .ZN(_u10_n21746 ) );
NAND2_X1 _u10_U10428  ( .A1(1'b0), .A2(_u10_n12329 ), .ZN(_u10_n21747 ) );
NAND2_X1 _u10_U10427  ( .A1(1'b0), .A2(_u10_n12305 ), .ZN(_u10_n21748 ) );
NAND2_X1 _u10_U10426  ( .A1(1'b0), .A2(_u10_n12281 ), .ZN(_u10_n21749 ) );
NAND4_X1 _u10_U10425  ( .A1(_u10_n21746 ), .A2(_u10_n21747 ), .A3(_u10_n21748 ), .A4(_u10_n21749 ), .ZN(_u10_n21731 ) );
NAND2_X1 _u10_U10424  ( .A1(1'b0), .A2(_u10_n12258 ), .ZN(_u10_n21742 ) );
NAND2_X1 _u10_U10423  ( .A1(1'b0), .A2(_u10_n12234 ), .ZN(_u10_n21743 ) );
NAND2_X1 _u10_U10422  ( .A1(1'b0), .A2(_u10_n12210 ), .ZN(_u10_n21744 ) );
NAND2_X1 _u10_U10421  ( .A1(1'b0), .A2(_u10_n12186 ), .ZN(_u10_n21745 ) );
NAND4_X1 _u10_U10420  ( .A1(_u10_n21742 ), .A2(_u10_n21743 ), .A3(_u10_n21744 ), .A4(_u10_n21745 ), .ZN(_u10_n21732 ) );
NAND2_X1 _u10_U10419  ( .A1(1'b0), .A2(_u10_n12163 ), .ZN(_u10_n21738 ) );
NAND2_X1 _u10_U10418  ( .A1(1'b0), .A2(_u10_n12139 ), .ZN(_u10_n21739 ) );
NAND2_X1 _u10_U10417  ( .A1(1'b0), .A2(_u10_n12115 ), .ZN(_u10_n21740 ) );
NAND2_X1 _u10_U10416  ( .A1(1'b0), .A2(_u10_n12091 ), .ZN(_u10_n21741 ) );
NAND4_X1 _u10_U10415  ( .A1(_u10_n21738 ), .A2(_u10_n21739 ), .A3(_u10_n21740 ), .A4(_u10_n21741 ), .ZN(_u10_n21733 ) );
NAND2_X1 _u10_U10414  ( .A1(1'b0), .A2(_u10_n12066 ), .ZN(_u10_n21735 ) );
NAND2_X1 _u10_U10413  ( .A1(1'b0), .A2(_u10_n12042 ), .ZN(_u10_n21736 ) );
NAND2_X1 _u10_U10412  ( .A1(ch0_adr0[7]), .A2(_u10_n12001 ), .ZN(_u10_n21737 ) );
NAND3_X1 _u10_U10411  ( .A1(_u10_n21735 ), .A2(_u10_n21736 ), .A3(_u10_n21737 ), .ZN(_u10_n21734 ) );
NOR4_X1 _u10_U10410  ( .A1(_u10_n21731 ), .A2(_u10_n21732 ), .A3(_u10_n21733 ), .A4(_u10_n21734 ), .ZN(_u10_n21709 ) );
NAND2_X1 _u10_U10409  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21727 ) );
NAND2_X1 _u10_U10408  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21728 ) );
NAND2_X1 _u10_U10407  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21729 ) );
NAND2_X1 _u10_U10406  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21730 ) );
NAND4_X1 _u10_U10405  ( .A1(_u10_n21727 ), .A2(_u10_n21728 ), .A3(_u10_n21729 ), .A4(_u10_n21730 ), .ZN(_u10_n21711 ) );
NAND2_X1 _u10_U10404  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21723 ) );
NAND2_X1 _u10_U10403  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21724 ) );
NAND2_X1 _u10_U10402  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21725 ) );
NAND2_X1 _u10_U10401  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21726 ) );
NAND4_X1 _u10_U10400  ( .A1(_u10_n21723 ), .A2(_u10_n21724 ), .A3(_u10_n21725 ), .A4(_u10_n21726 ), .ZN(_u10_n21712 ) );
NAND2_X1 _u10_U10399  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21719 ) );
NAND2_X1 _u10_U10398  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21720 ) );
NAND2_X1 _u10_U10397  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21721 ) );
NAND2_X1 _u10_U10396  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21722 ) );
NAND4_X1 _u10_U10395  ( .A1(_u10_n21719 ), .A2(_u10_n21720 ), .A3(_u10_n21721 ), .A4(_u10_n21722 ), .ZN(_u10_n21713 ) );
NAND2_X1 _u10_U10394  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21715 ) );
NAND2_X1 _u10_U10393  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21716 ) );
NAND2_X1 _u10_U10392  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21717 ) );
NAND2_X1 _u10_U10391  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21718 ) );
NAND4_X1 _u10_U10390  ( .A1(_u10_n21715 ), .A2(_u10_n21716 ), .A3(_u10_n21717 ), .A4(_u10_n21718 ), .ZN(_u10_n21714 ) );
NOR4_X1 _u10_U10389  ( .A1(_u10_n21711 ), .A2(_u10_n21712 ), .A3(_u10_n21713 ), .A4(_u10_n21714 ), .ZN(_u10_n21710 ) );
NAND2_X1 _u10_U10388  ( .A1(_u10_n21709 ), .A2(_u10_n21710 ), .ZN(adr0[7]));
NAND2_X1 _u10_U10387  ( .A1(1'b0), .A2(_u10_n12353 ), .ZN(_u10_n21705 ) );
NAND2_X1 _u10_U10386  ( .A1(1'b0), .A2(_u10_n12328 ), .ZN(_u10_n21706 ) );
NAND2_X1 _u10_U10385  ( .A1(1'b0), .A2(_u10_n12304 ), .ZN(_u10_n21707 ) );
NAND2_X1 _u10_U10384  ( .A1(1'b0), .A2(_u10_n12280 ), .ZN(_u10_n21708 ) );
NAND4_X1 _u10_U10383  ( .A1(_u10_n21705 ), .A2(_u10_n21706 ), .A3(_u10_n21707 ), .A4(_u10_n21708 ), .ZN(_u10_n21690 ) );
NAND2_X1 _u10_U10382  ( .A1(1'b0), .A2(_u10_n12257 ), .ZN(_u10_n21701 ) );
NAND2_X1 _u10_U10381  ( .A1(1'b0), .A2(_u10_n12233 ), .ZN(_u10_n21702 ) );
NAND2_X1 _u10_U10380  ( .A1(1'b0), .A2(_u10_n12207 ), .ZN(_u10_n21703 ) );
NAND2_X1 _u10_U10379  ( .A1(1'b0), .A2(_u10_n12185 ), .ZN(_u10_n21704 ) );
NAND4_X1 _u10_U10378  ( .A1(_u10_n21701 ), .A2(_u10_n21702 ), .A3(_u10_n21703 ), .A4(_u10_n21704 ), .ZN(_u10_n21691 ) );
NAND2_X1 _u10_U10377  ( .A1(1'b0), .A2(_u10_n12162 ), .ZN(_u10_n21697 ) );
NAND2_X1 _u10_U10376  ( .A1(1'b0), .A2(_u10_n12138 ), .ZN(_u10_n21698 ) );
NAND2_X1 _u10_U10375  ( .A1(1'b0), .A2(_u10_n12114 ), .ZN(_u10_n21699 ) );
NAND2_X1 _u10_U10374  ( .A1(1'b0), .A2(_u10_n12090 ), .ZN(_u10_n21700 ) );
NAND4_X1 _u10_U10373  ( .A1(_u10_n21697 ), .A2(_u10_n21698 ), .A3(_u10_n21699 ), .A4(_u10_n21700 ), .ZN(_u10_n21692 ) );
NAND2_X1 _u10_U10372  ( .A1(1'b0), .A2(_u10_n12063 ), .ZN(_u10_n21694 ) );
NAND2_X1 _u10_U10371  ( .A1(1'b0), .A2(_u10_n12039 ), .ZN(_u10_n21695 ) );
NAND2_X1 _u10_U10370  ( .A1(ch0_adr0[8]), .A2(_u10_n12001 ), .ZN(_u10_n21696 ) );
NAND3_X1 _u10_U10369  ( .A1(_u10_n21694 ), .A2(_u10_n21695 ), .A3(_u10_n21696 ), .ZN(_u10_n21693 ) );
NOR4_X1 _u10_U10368  ( .A1(_u10_n21690 ), .A2(_u10_n21691 ), .A3(_u10_n21692 ), .A4(_u10_n21693 ), .ZN(_u10_n21668 ) );
NAND2_X1 _u10_U10367  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21686 ) );
NAND2_X1 _u10_U10366  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21687 ) );
NAND2_X1 _u10_U10365  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21688 ) );
NAND2_X1 _u10_U10364  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21689 ) );
NAND4_X1 _u10_U10363  ( .A1(_u10_n21686 ), .A2(_u10_n21687 ), .A3(_u10_n21688 ), .A4(_u10_n21689 ), .ZN(_u10_n21670 ) );
NAND2_X1 _u10_U10362  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21682 ) );
NAND2_X1 _u10_U10361  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21683 ) );
NAND2_X1 _u10_U10360  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21684 ) );
NAND2_X1 _u10_U10359  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21685 ) );
NAND4_X1 _u10_U10358  ( .A1(_u10_n21682 ), .A2(_u10_n21683 ), .A3(_u10_n21684 ), .A4(_u10_n21685 ), .ZN(_u10_n21671 ) );
NAND2_X1 _u10_U10357  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21678 ) );
NAND2_X1 _u10_U10356  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21679 ) );
NAND2_X1 _u10_U10355  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21680 ) );
NAND2_X1 _u10_U10354  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21681 ) );
NAND4_X1 _u10_U10353  ( .A1(_u10_n21678 ), .A2(_u10_n21679 ), .A3(_u10_n21680 ), .A4(_u10_n21681 ), .ZN(_u10_n21672 ) );
NAND2_X1 _u10_U10352  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21674 ) );
NAND2_X1 _u10_U10351  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21675 ) );
NAND2_X1 _u10_U10350  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21676 ) );
NAND2_X1 _u10_U10349  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21677 ) );
NAND4_X1 _u10_U10348  ( .A1(_u10_n21674 ), .A2(_u10_n21675 ), .A3(_u10_n21676 ), .A4(_u10_n21677 ), .ZN(_u10_n21673 ) );
NOR4_X1 _u10_U10347  ( .A1(_u10_n21670 ), .A2(_u10_n21671 ), .A3(_u10_n21672 ), .A4(_u10_n21673 ), .ZN(_u10_n21669 ) );
NAND2_X1 _u10_U10346  ( .A1(_u10_n21668 ), .A2(_u10_n21669 ), .ZN(adr0[8]));
NAND2_X1 _u10_U10345  ( .A1(1'b0), .A2(_u10_n12355 ), .ZN(_u10_n21664 ) );
NAND2_X1 _u10_U10344  ( .A1(1'b0), .A2(_u10_n12429 ), .ZN(_u10_n21665 ) );
NAND2_X1 _u10_U10343  ( .A1(1'b0), .A2(_u10_n12305 ), .ZN(_u10_n21666 ) );
NAND2_X1 _u10_U10342  ( .A1(1'b0), .A2(_u10_n12281 ), .ZN(_u10_n21667 ) );
NAND4_X1 _u10_U10341  ( .A1(_u10_n21664 ), .A2(_u10_n21665 ), .A3(_u10_n21666 ), .A4(_u10_n21667 ), .ZN(_u10_n21649 ) );
NAND2_X1 _u10_U10340  ( .A1(1'b0), .A2(_u10_n12259 ), .ZN(_u10_n21660 ) );
NAND2_X1 _u10_U10339  ( .A1(1'b0), .A2(_u10_n12235 ), .ZN(_u10_n21661 ) );
NAND2_X1 _u10_U10338  ( .A1(1'b0), .A2(_u10_n12210 ), .ZN(_u10_n21662 ) );
NAND2_X1 _u10_U10337  ( .A1(1'b0), .A2(_u10_n12187 ), .ZN(_u10_n21663 ) );
NAND4_X1 _u10_U10336  ( .A1(_u10_n21660 ), .A2(_u10_n21661 ), .A3(_u10_n21662 ), .A4(_u10_n21663 ), .ZN(_u10_n21650 ) );
NAND2_X1 _u10_U10335  ( .A1(1'b0), .A2(_u10_n12159 ), .ZN(_u10_n21656 ) );
NAND2_X1 _u10_U10334  ( .A1(1'b0), .A2(_u10_n12135 ), .ZN(_u10_n21657 ) );
NAND2_X1 _u10_U10333  ( .A1(1'b0), .A2(_u10_n12111 ), .ZN(_u10_n21658 ) );
NAND2_X1 _u10_U10332  ( .A1(1'b0), .A2(_u10_n12087 ), .ZN(_u10_n21659 ) );
NAND4_X1 _u10_U10331  ( .A1(_u10_n21656 ), .A2(_u10_n21657 ), .A3(_u10_n21658 ), .A4(_u10_n21659 ), .ZN(_u10_n21651 ) );
NAND2_X1 _u10_U10330  ( .A1(1'b0), .A2(_u10_n12406 ), .ZN(_u10_n21653 ) );
NAND2_X1 _u10_U10329  ( .A1(1'b0), .A2(_u10_n12405 ), .ZN(_u10_n21654 ) );
NAND2_X1 _u10_U10328  ( .A1(ch0_adr0[9]), .A2(_u10_n12001 ), .ZN(_u10_n21655 ) );
NAND3_X1 _u10_U10327  ( .A1(_u10_n21653 ), .A2(_u10_n21654 ), .A3(_u10_n21655 ), .ZN(_u10_n21652 ) );
NOR4_X1 _u10_U10326  ( .A1(_u10_n21649 ), .A2(_u10_n21650 ), .A3(_u10_n21651 ), .A4(_u10_n21652 ), .ZN(_u10_n21627 ) );
NAND2_X1 _u10_U10325  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21645 ) );
NAND2_X1 _u10_U10324  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21646 ) );
NAND2_X1 _u10_U10323  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21647 ) );
NAND2_X1 _u10_U10322  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21648 ) );
NAND4_X1 _u10_U10321  ( .A1(_u10_n21645 ), .A2(_u10_n21646 ), .A3(_u10_n21647 ), .A4(_u10_n21648 ), .ZN(_u10_n21629 ) );
NAND2_X1 _u10_U10320  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21641 ) );
NAND2_X1 _u10_U10319  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21642 ) );
NAND2_X1 _u10_U10318  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21643 ) );
NAND2_X1 _u10_U10317  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21644 ) );
NAND4_X1 _u10_U10316  ( .A1(_u10_n21641 ), .A2(_u10_n21642 ), .A3(_u10_n21643 ), .A4(_u10_n21644 ), .ZN(_u10_n21630 ) );
NAND2_X1 _u10_U10315  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21637 ) );
NAND2_X1 _u10_U10314  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21638 ) );
NAND2_X1 _u10_U10313  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21639 ) );
NAND2_X1 _u10_U10312  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21640 ) );
NAND4_X1 _u10_U10311  ( .A1(_u10_n21637 ), .A2(_u10_n21638 ), .A3(_u10_n21639 ), .A4(_u10_n21640 ), .ZN(_u10_n21631 ) );
NAND2_X1 _u10_U10310  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21633 ) );
NAND2_X1 _u10_U10309  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21634 ) );
NAND2_X1 _u10_U10308  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21635 ) );
NAND2_X1 _u10_U10307  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21636 ) );
NAND4_X1 _u10_U10306  ( .A1(_u10_n21633 ), .A2(_u10_n21634 ), .A3(_u10_n21635 ), .A4(_u10_n21636 ), .ZN(_u10_n21632 ) );
NOR4_X1 _u10_U10305  ( .A1(_u10_n21629 ), .A2(_u10_n21630 ), .A3(_u10_n21631 ), .A4(_u10_n21632 ), .ZN(_u10_n21628 ) );
NAND2_X1 _u10_U10304  ( .A1(_u10_n21627 ), .A2(_u10_n21628 ), .ZN(adr0[9]));
NAND2_X1 _u10_U10303  ( .A1(1'b0), .A2(_u10_n12356 ), .ZN(_u10_n21623 ) );
NAND2_X1 _u10_U10302  ( .A1(1'b0), .A2(_u10_n12332 ), .ZN(_u10_n21624 ) );
NAND2_X1 _u10_U10301  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n21625 ) );
NAND2_X1 _u10_U10300  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n21626 ) );
NAND4_X1 _u10_U10299  ( .A1(_u10_n21623 ), .A2(_u10_n21624 ), .A3(_u10_n21625 ), .A4(_u10_n21626 ), .ZN(_u10_n21608 ) );
NAND2_X1 _u10_U10298  ( .A1(1'b0), .A2(_u10_n12260 ), .ZN(_u10_n21619 ) );
NAND2_X1 _u10_U10297  ( .A1(1'b0), .A2(_u10_n12236 ), .ZN(_u10_n21620 ) );
NAND2_X1 _u10_U10296  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n21621 ) );
NAND2_X1 _u10_U10295  ( .A1(1'b0), .A2(_u10_n12188 ), .ZN(_u10_n21622 ) );
NAND4_X1 _u10_U10294  ( .A1(_u10_n21619 ), .A2(_u10_n21620 ), .A3(_u10_n21621 ), .A4(_u10_n21622 ), .ZN(_u10_n21609 ) );
NAND2_X1 _u10_U10293  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n21615 ) );
NAND2_X1 _u10_U10292  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n21616 ) );
NAND2_X1 _u10_U10291  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n21617 ) );
NAND2_X1 _u10_U10290  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n21618 ) );
NAND4_X1 _u10_U10289  ( .A1(_u10_n21615 ), .A2(_u10_n21616 ), .A3(_u10_n21617 ), .A4(_u10_n21618 ), .ZN(_u10_n21610 ) );
NAND2_X1 _u10_U10288  ( .A1(1'b0), .A2(_u10_n12068 ), .ZN(_u10_n21612 ) );
NAND2_X1 _u10_U10287  ( .A1(1'b0), .A2(_u10_n12044 ), .ZN(_u10_n21613 ) );
NAND2_X1 _u10_U10286  ( .A1(1'b0), .A2(_u10_n12001 ), .ZN(_u10_n21614 ) );
NAND3_X1 _u10_U10285  ( .A1(_u10_n21612 ), .A2(_u10_n21613 ), .A3(_u10_n21614 ), .ZN(_u10_n21611 ) );
NOR4_X1 _u10_U10284  ( .A1(_u10_n21608 ), .A2(_u10_n21609 ), .A3(_u10_n21610 ), .A4(_u10_n21611 ), .ZN(_u10_n21586 ) );
NAND2_X1 _u10_U10283  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21604 ) );
NAND2_X1 _u10_U10282  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21605 ) );
NAND2_X1 _u10_U10281  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21606 ) );
NAND2_X1 _u10_U10280  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21607 ) );
NAND4_X1 _u10_U10279  ( .A1(_u10_n21604 ), .A2(_u10_n21605 ), .A3(_u10_n21606 ), .A4(_u10_n21607 ), .ZN(_u10_n21588 ) );
NAND2_X1 _u10_U10278  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21600 ) );
NAND2_X1 _u10_U10277  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21601 ) );
NAND2_X1 _u10_U10276  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21602 ) );
NAND2_X1 _u10_U10275  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21603 ) );
NAND4_X1 _u10_U10274  ( .A1(_u10_n21600 ), .A2(_u10_n21601 ), .A3(_u10_n21602 ), .A4(_u10_n21603 ), .ZN(_u10_n21589 ) );
NAND2_X1 _u10_U10273  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21596 ) );
NAND2_X1 _u10_U10272  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21597 ) );
NAND2_X1 _u10_U10271  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21598 ) );
NAND2_X1 _u10_U10270  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21599 ) );
NAND4_X1 _u10_U10269  ( .A1(_u10_n21596 ), .A2(_u10_n21597 ), .A3(_u10_n21598 ), .A4(_u10_n21599 ), .ZN(_u10_n21590 ) );
NAND2_X1 _u10_U10268  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21592 ) );
NAND2_X1 _u10_U10267  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21593 ) );
NAND2_X1 _u10_U10266  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21594 ) );
NAND2_X1 _u10_U10265  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21595 ) );
NAND4_X1 _u10_U10264  ( .A1(_u10_n21592 ), .A2(_u10_n21593 ), .A3(_u10_n21594 ), .A4(_u10_n21595 ), .ZN(_u10_n21591 ) );
NOR4_X1 _u10_U10263  ( .A1(_u10_n21588 ), .A2(_u10_n21589 ), .A3(_u10_n21590 ), .A4(_u10_n21591 ), .ZN(_u10_n21587 ) );
NAND2_X1 _u10_U10262  ( .A1(_u10_n21586 ), .A2(_u10_n21587 ), .ZN(adr1[0]));
NAND2_X1 _u10_U10261  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21582 ) );
NAND2_X1 _u10_U10260  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21583 ) );
NAND2_X1 _u10_U10259  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21584 ) );
NAND2_X1 _u10_U10258  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21585 ) );
NAND4_X1 _u10_U10257  ( .A1(_u10_n21582 ), .A2(_u10_n21583 ), .A3(_u10_n21584 ), .A4(_u10_n21585 ), .ZN(_u10_n21567 ) );
NAND2_X1 _u10_U10256  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21578 ) );
NAND2_X1 _u10_U10255  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21579 ) );
NAND2_X1 _u10_U10254  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21580 ) );
NAND2_X1 _u10_U10253  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21581 ) );
NAND4_X1 _u10_U10252  ( .A1(_u10_n21578 ), .A2(_u10_n21579 ), .A3(_u10_n21580 ), .A4(_u10_n21581 ), .ZN(_u10_n21568 ) );
NAND2_X1 _u10_U10251  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21574 ) );
NAND2_X1 _u10_U10250  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21575 ) );
NAND2_X1 _u10_U10249  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21576 ) );
NAND2_X1 _u10_U10248  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21577 ) );
NAND4_X1 _u10_U10247  ( .A1(_u10_n21574 ), .A2(_u10_n21575 ), .A3(_u10_n21576 ), .A4(_u10_n21577 ), .ZN(_u10_n21569 ) );
NAND2_X1 _u10_U10246  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21571 ) );
NAND2_X1 _u10_U10245  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21572 ) );
NAND2_X1 _u10_U10244  ( .A1(ch0_adr1[10]), .A2(_u10_n12001 ), .ZN(_u10_n21573 ) );
NAND3_X1 _u10_U10243  ( .A1(_u10_n21571 ), .A2(_u10_n21572 ), .A3(_u10_n21573 ), .ZN(_u10_n21570 ) );
NOR4_X1 _u10_U10242  ( .A1(_u10_n21567 ), .A2(_u10_n21568 ), .A3(_u10_n21569 ), .A4(_u10_n21570 ), .ZN(_u10_n21545 ) );
NAND2_X1 _u10_U10241  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21563 ) );
NAND2_X1 _u10_U10240  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21564 ) );
NAND2_X1 _u10_U10239  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21565 ) );
NAND2_X1 _u10_U10238  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21566 ) );
NAND4_X1 _u10_U10237  ( .A1(_u10_n21563 ), .A2(_u10_n21564 ), .A3(_u10_n21565 ), .A4(_u10_n21566 ), .ZN(_u10_n21547 ) );
NAND2_X1 _u10_U10236  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21559 ) );
NAND2_X1 _u10_U10235  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21560 ) );
NAND2_X1 _u10_U10234  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21561 ) );
NAND2_X1 _u10_U10233  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21562 ) );
NAND4_X1 _u10_U10232  ( .A1(_u10_n21559 ), .A2(_u10_n21560 ), .A3(_u10_n21561 ), .A4(_u10_n21562 ), .ZN(_u10_n21548 ) );
NAND2_X1 _u10_U10231  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21555 ) );
NAND2_X1 _u10_U10230  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21556 ) );
NAND2_X1 _u10_U10229  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21557 ) );
NAND2_X1 _u10_U10228  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21558 ) );
NAND4_X1 _u10_U10227  ( .A1(_u10_n21555 ), .A2(_u10_n21556 ), .A3(_u10_n21557 ), .A4(_u10_n21558 ), .ZN(_u10_n21549 ) );
NAND2_X1 _u10_U10226  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21551 ) );
NAND2_X1 _u10_U10225  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21552 ) );
NAND2_X1 _u10_U10224  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21553 ) );
NAND2_X1 _u10_U10223  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21554 ) );
NAND4_X1 _u10_U10222  ( .A1(_u10_n21551 ), .A2(_u10_n21552 ), .A3(_u10_n21553 ), .A4(_u10_n21554 ), .ZN(_u10_n21550 ) );
NOR4_X1 _u10_U10221  ( .A1(_u10_n21547 ), .A2(_u10_n21548 ), .A3(_u10_n21549 ), .A4(_u10_n21550 ), .ZN(_u10_n21546 ) );
NAND2_X1 _u10_U10220  ( .A1(_u10_n21545 ), .A2(_u10_n21546 ), .ZN(adr1[10]));
NAND2_X1 _u10_U10219  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21541 ) );
NAND2_X1 _u10_U10218  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21542 ) );
NAND2_X1 _u10_U10217  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21543 ) );
NAND2_X1 _u10_U10216  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21544 ) );
NAND4_X1 _u10_U10215  ( .A1(_u10_n21541 ), .A2(_u10_n21542 ), .A3(_u10_n21543 ), .A4(_u10_n21544 ), .ZN(_u10_n21526 ) );
NAND2_X1 _u10_U10214  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21537 ) );
NAND2_X1 _u10_U10213  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21538 ) );
NAND2_X1 _u10_U10212  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21539 ) );
NAND2_X1 _u10_U10211  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21540 ) );
NAND4_X1 _u10_U10210  ( .A1(_u10_n21537 ), .A2(_u10_n21538 ), .A3(_u10_n21539 ), .A4(_u10_n21540 ), .ZN(_u10_n21527 ) );
NAND2_X1 _u10_U10209  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21533 ) );
NAND2_X1 _u10_U10208  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21534 ) );
NAND2_X1 _u10_U10207  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21535 ) );
NAND2_X1 _u10_U10206  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21536 ) );
NAND4_X1 _u10_U10205  ( .A1(_u10_n21533 ), .A2(_u10_n21534 ), .A3(_u10_n21535 ), .A4(_u10_n21536 ), .ZN(_u10_n21528 ) );
NAND2_X1 _u10_U10204  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21530 ) );
NAND2_X1 _u10_U10203  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21531 ) );
NAND2_X1 _u10_U10202  ( .A1(ch0_adr1[11]), .A2(_u10_n12001 ), .ZN(_u10_n21532 ) );
NAND3_X1 _u10_U10201  ( .A1(_u10_n21530 ), .A2(_u10_n21531 ), .A3(_u10_n21532 ), .ZN(_u10_n21529 ) );
NOR4_X1 _u10_U10200  ( .A1(_u10_n21526 ), .A2(_u10_n21527 ), .A3(_u10_n21528 ), .A4(_u10_n21529 ), .ZN(_u10_n21504 ) );
NAND2_X1 _u10_U10199  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21522 ) );
NAND2_X1 _u10_U10198  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21523 ) );
NAND2_X1 _u10_U10197  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21524 ) );
NAND2_X1 _u10_U10196  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21525 ) );
NAND4_X1 _u10_U10195  ( .A1(_u10_n21522 ), .A2(_u10_n21523 ), .A3(_u10_n21524 ), .A4(_u10_n21525 ), .ZN(_u10_n21506 ) );
NAND2_X1 _u10_U10194  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21518 ) );
NAND2_X1 _u10_U10193  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21519 ) );
NAND2_X1 _u10_U10192  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21520 ) );
NAND2_X1 _u10_U10191  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21521 ) );
NAND4_X1 _u10_U10190  ( .A1(_u10_n21518 ), .A2(_u10_n21519 ), .A3(_u10_n21520 ), .A4(_u10_n21521 ), .ZN(_u10_n21507 ) );
NAND2_X1 _u10_U10189  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21514 ) );
NAND2_X1 _u10_U10188  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21515 ) );
NAND2_X1 _u10_U10187  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21516 ) );
NAND2_X1 _u10_U10186  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21517 ) );
NAND4_X1 _u10_U10185  ( .A1(_u10_n21514 ), .A2(_u10_n21515 ), .A3(_u10_n21516 ), .A4(_u10_n21517 ), .ZN(_u10_n21508 ) );
NAND2_X1 _u10_U10184  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21510 ) );
NAND2_X1 _u10_U10183  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21511 ) );
NAND2_X1 _u10_U10182  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21512 ) );
NAND2_X1 _u10_U10181  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21513 ) );
NAND4_X1 _u10_U10180  ( .A1(_u10_n21510 ), .A2(_u10_n21511 ), .A3(_u10_n21512 ), .A4(_u10_n21513 ), .ZN(_u10_n21509 ) );
NOR4_X1 _u10_U10179  ( .A1(_u10_n21506 ), .A2(_u10_n21507 ), .A3(_u10_n21508 ), .A4(_u10_n21509 ), .ZN(_u10_n21505 ) );
NAND2_X1 _u10_U10178  ( .A1(_u10_n21504 ), .A2(_u10_n21505 ), .ZN(adr1[11]));
NAND2_X1 _u10_U10177  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21500 ) );
NAND2_X1 _u10_U10176  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21501 ) );
NAND2_X1 _u10_U10175  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21502 ) );
NAND2_X1 _u10_U10174  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21503 ) );
NAND4_X1 _u10_U10173  ( .A1(_u10_n21500 ), .A2(_u10_n21501 ), .A3(_u10_n21502 ), .A4(_u10_n21503 ), .ZN(_u10_n21485 ) );
NAND2_X1 _u10_U10172  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21496 ) );
NAND2_X1 _u10_U10171  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21497 ) );
NAND2_X1 _u10_U10170  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21498 ) );
NAND2_X1 _u10_U10169  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21499 ) );
NAND4_X1 _u10_U10168  ( .A1(_u10_n21496 ), .A2(_u10_n21497 ), .A3(_u10_n21498 ), .A4(_u10_n21499 ), .ZN(_u10_n21486 ) );
NAND2_X1 _u10_U10167  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21492 ) );
NAND2_X1 _u10_U10166  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21493 ) );
NAND2_X1 _u10_U10165  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21494 ) );
NAND2_X1 _u10_U10164  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21495 ) );
NAND4_X1 _u10_U10163  ( .A1(_u10_n21492 ), .A2(_u10_n21493 ), .A3(_u10_n21494 ), .A4(_u10_n21495 ), .ZN(_u10_n21487 ) );
NAND2_X1 _u10_U10162  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21489 ) );
NAND2_X1 _u10_U10161  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21490 ) );
NAND2_X1 _u10_U10160  ( .A1(ch0_adr1[12]), .A2(_u10_n12002 ), .ZN(_u10_n21491 ) );
NAND3_X1 _u10_U10159  ( .A1(_u10_n21489 ), .A2(_u10_n21490 ), .A3(_u10_n21491 ), .ZN(_u10_n21488 ) );
NOR4_X1 _u10_U10158  ( .A1(_u10_n21485 ), .A2(_u10_n21486 ), .A3(_u10_n21487 ), .A4(_u10_n21488 ), .ZN(_u10_n21463 ) );
NAND2_X1 _u10_U10157  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21481 ) );
NAND2_X1 _u10_U10156  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21482 ) );
NAND2_X1 _u10_U10155  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21483 ) );
NAND2_X1 _u10_U10154  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21484 ) );
NAND4_X1 _u10_U10153  ( .A1(_u10_n21481 ), .A2(_u10_n21482 ), .A3(_u10_n21483 ), .A4(_u10_n21484 ), .ZN(_u10_n21465 ) );
NAND2_X1 _u10_U10152  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21477 ) );
NAND2_X1 _u10_U10151  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21478 ) );
NAND2_X1 _u10_U10150  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21479 ) );
NAND2_X1 _u10_U10149  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21480 ) );
NAND4_X1 _u10_U10148  ( .A1(_u10_n21477 ), .A2(_u10_n21478 ), .A3(_u10_n21479 ), .A4(_u10_n21480 ), .ZN(_u10_n21466 ) );
NAND2_X1 _u10_U10147  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21473 ) );
NAND2_X1 _u10_U10146  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21474 ) );
NAND2_X1 _u10_U10145  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21475 ) );
NAND2_X1 _u10_U10144  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21476 ) );
NAND4_X1 _u10_U10143  ( .A1(_u10_n21473 ), .A2(_u10_n21474 ), .A3(_u10_n21475 ), .A4(_u10_n21476 ), .ZN(_u10_n21467 ) );
NAND2_X1 _u10_U10142  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21469 ) );
NAND2_X1 _u10_U10141  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21470 ) );
NAND2_X1 _u10_U10140  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21471 ) );
NAND2_X1 _u10_U10139  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21472 ) );
NAND4_X1 _u10_U10138  ( .A1(_u10_n21469 ), .A2(_u10_n21470 ), .A3(_u10_n21471 ), .A4(_u10_n21472 ), .ZN(_u10_n21468 ) );
NOR4_X1 _u10_U10137  ( .A1(_u10_n21465 ), .A2(_u10_n21466 ), .A3(_u10_n21467 ), .A4(_u10_n21468 ), .ZN(_u10_n21464 ) );
NAND2_X1 _u10_U10136  ( .A1(_u10_n21463 ), .A2(_u10_n21464 ), .ZN(adr1[12]));
NAND2_X1 _u10_U10135  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21459 ) );
NAND2_X1 _u10_U10134  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21460 ) );
NAND2_X1 _u10_U10133  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21461 ) );
NAND2_X1 _u10_U10132  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21462 ) );
NAND4_X1 _u10_U10131  ( .A1(_u10_n21459 ), .A2(_u10_n21460 ), .A3(_u10_n21461 ), .A4(_u10_n21462 ), .ZN(_u10_n21444 ) );
NAND2_X1 _u10_U10130  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21455 ) );
NAND2_X1 _u10_U10129  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21456 ) );
NAND2_X1 _u10_U10128  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21457 ) );
NAND2_X1 _u10_U10127  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21458 ) );
NAND4_X1 _u10_U10126  ( .A1(_u10_n21455 ), .A2(_u10_n21456 ), .A3(_u10_n21457 ), .A4(_u10_n21458 ), .ZN(_u10_n21445 ) );
NAND2_X1 _u10_U10125  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21451 ) );
NAND2_X1 _u10_U10124  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21452 ) );
NAND2_X1 _u10_U10123  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21453 ) );
NAND2_X1 _u10_U10122  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21454 ) );
NAND4_X1 _u10_U10121  ( .A1(_u10_n21451 ), .A2(_u10_n21452 ), .A3(_u10_n21453 ), .A4(_u10_n21454 ), .ZN(_u10_n21446 ) );
NAND2_X1 _u10_U10120  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21448 ) );
NAND2_X1 _u10_U10119  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21449 ) );
NAND2_X1 _u10_U10118  ( .A1(ch0_adr1[13]), .A2(_u10_n12002 ), .ZN(_u10_n21450 ) );
NAND3_X1 _u10_U10117  ( .A1(_u10_n21448 ), .A2(_u10_n21449 ), .A3(_u10_n21450 ), .ZN(_u10_n21447 ) );
NOR4_X1 _u10_U10116  ( .A1(_u10_n21444 ), .A2(_u10_n21445 ), .A3(_u10_n21446 ), .A4(_u10_n21447 ), .ZN(_u10_n21422 ) );
NAND2_X1 _u10_U10115  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21440 ) );
NAND2_X1 _u10_U10114  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21441 ) );
NAND2_X1 _u10_U10113  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21442 ) );
NAND2_X1 _u10_U10112  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21443 ) );
NAND4_X1 _u10_U10111  ( .A1(_u10_n21440 ), .A2(_u10_n21441 ), .A3(_u10_n21442 ), .A4(_u10_n21443 ), .ZN(_u10_n21424 ) );
NAND2_X1 _u10_U10110  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21436 ) );
NAND2_X1 _u10_U10109  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21437 ) );
NAND2_X1 _u10_U10108  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21438 ) );
NAND2_X1 _u10_U10107  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21439 ) );
NAND4_X1 _u10_U10106  ( .A1(_u10_n21436 ), .A2(_u10_n21437 ), .A3(_u10_n21438 ), .A4(_u10_n21439 ), .ZN(_u10_n21425 ) );
NAND2_X1 _u10_U10105  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21432 ) );
NAND2_X1 _u10_U10104  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21433 ) );
NAND2_X1 _u10_U10103  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21434 ) );
NAND2_X1 _u10_U10102  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21435 ) );
NAND4_X1 _u10_U10101  ( .A1(_u10_n21432 ), .A2(_u10_n21433 ), .A3(_u10_n21434 ), .A4(_u10_n21435 ), .ZN(_u10_n21426 ) );
NAND2_X1 _u10_U10100  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21428 ) );
NAND2_X1 _u10_U10099  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21429 ) );
NAND2_X1 _u10_U10098  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21430 ) );
NAND2_X1 _u10_U10097  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21431 ) );
NAND4_X1 _u10_U10096  ( .A1(_u10_n21428 ), .A2(_u10_n21429 ), .A3(_u10_n21430 ), .A4(_u10_n21431 ), .ZN(_u10_n21427 ) );
NOR4_X1 _u10_U10095  ( .A1(_u10_n21424 ), .A2(_u10_n21425 ), .A3(_u10_n21426 ), .A4(_u10_n21427 ), .ZN(_u10_n21423 ) );
NAND2_X1 _u10_U10094  ( .A1(_u10_n21422 ), .A2(_u10_n21423 ), .ZN(adr1[13]));
NAND2_X1 _u10_U10093  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21418 ) );
NAND2_X1 _u10_U10092  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21419 ) );
NAND2_X1 _u10_U10091  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21420 ) );
NAND2_X1 _u10_U10090  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21421 ) );
NAND4_X1 _u10_U10089  ( .A1(_u10_n21418 ), .A2(_u10_n21419 ), .A3(_u10_n21420 ), .A4(_u10_n21421 ), .ZN(_u10_n21403 ) );
NAND2_X1 _u10_U10088  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21414 ) );
NAND2_X1 _u10_U10087  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21415 ) );
NAND2_X1 _u10_U10086  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21416 ) );
NAND2_X1 _u10_U10085  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21417 ) );
NAND4_X1 _u10_U10084  ( .A1(_u10_n21414 ), .A2(_u10_n21415 ), .A3(_u10_n21416 ), .A4(_u10_n21417 ), .ZN(_u10_n21404 ) );
NAND2_X1 _u10_U10083  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21410 ) );
NAND2_X1 _u10_U10082  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21411 ) );
NAND2_X1 _u10_U10081  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21412 ) );
NAND2_X1 _u10_U10080  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21413 ) );
NAND4_X1 _u10_U10079  ( .A1(_u10_n21410 ), .A2(_u10_n21411 ), .A3(_u10_n21412 ), .A4(_u10_n21413 ), .ZN(_u10_n21405 ) );
NAND2_X1 _u10_U10078  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21407 ) );
NAND2_X1 _u10_U10077  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21408 ) );
NAND2_X1 _u10_U10076  ( .A1(ch0_adr1[14]), .A2(_u10_n12002 ), .ZN(_u10_n21409 ) );
NAND3_X1 _u10_U10075  ( .A1(_u10_n21407 ), .A2(_u10_n21408 ), .A3(_u10_n21409 ), .ZN(_u10_n21406 ) );
NOR4_X1 _u10_U10074  ( .A1(_u10_n21403 ), .A2(_u10_n21404 ), .A3(_u10_n21405 ), .A4(_u10_n21406 ), .ZN(_u10_n21381 ) );
NAND2_X1 _u10_U10073  ( .A1(1'b0), .A2(_u10_n11985 ), .ZN(_u10_n21399 ) );
NAND2_X1 _u10_U10072  ( .A1(1'b0), .A2(_u10_n11961 ), .ZN(_u10_n21400 ) );
NAND2_X1 _u10_U10071  ( .A1(1'b0), .A2(_u10_n11937 ), .ZN(_u10_n21401 ) );
NAND2_X1 _u10_U10070  ( .A1(1'b0), .A2(_u10_n11913 ), .ZN(_u10_n21402 ) );
NAND4_X1 _u10_U10069  ( .A1(_u10_n21399 ), .A2(_u10_n21400 ), .A3(_u10_n21401 ), .A4(_u10_n21402 ), .ZN(_u10_n21383 ) );
NAND2_X1 _u10_U10068  ( .A1(1'b0), .A2(_u10_n11889 ), .ZN(_u10_n21395 ) );
NAND2_X1 _u10_U10067  ( .A1(1'b0), .A2(_u10_n11865 ), .ZN(_u10_n21396 ) );
NAND2_X1 _u10_U10066  ( .A1(1'b0), .A2(_u10_n11841 ), .ZN(_u10_n21397 ) );
NAND2_X1 _u10_U10065  ( .A1(1'b0), .A2(_u10_n11817 ), .ZN(_u10_n21398 ) );
NAND4_X1 _u10_U10064  ( .A1(_u10_n21395 ), .A2(_u10_n21396 ), .A3(_u10_n21397 ), .A4(_u10_n21398 ), .ZN(_u10_n21384 ) );
NAND2_X1 _u10_U10063  ( .A1(1'b0), .A2(_u10_n11793 ), .ZN(_u10_n21391 ) );
NAND2_X1 _u10_U10062  ( .A1(1'b0), .A2(_u10_n11769 ), .ZN(_u10_n21392 ) );
NAND2_X1 _u10_U10061  ( .A1(1'b0), .A2(_u10_n11745 ), .ZN(_u10_n21393 ) );
NAND2_X1 _u10_U10060  ( .A1(1'b0), .A2(_u10_n11721 ), .ZN(_u10_n21394 ) );
NAND4_X1 _u10_U10059  ( .A1(_u10_n21391 ), .A2(_u10_n21392 ), .A3(_u10_n21393 ), .A4(_u10_n21394 ), .ZN(_u10_n21385 ) );
NAND2_X1 _u10_U10058  ( .A1(1'b0), .A2(_u10_n11697 ), .ZN(_u10_n21387 ) );
NAND2_X1 _u10_U10057  ( .A1(1'b0), .A2(_u10_n11673 ), .ZN(_u10_n21388 ) );
NAND2_X1 _u10_U10056  ( .A1(1'b0), .A2(_u10_n11649 ), .ZN(_u10_n21389 ) );
NAND2_X1 _u10_U10055  ( .A1(1'b0), .A2(_u10_n11625 ), .ZN(_u10_n21390 ) );
NAND4_X1 _u10_U10054  ( .A1(_u10_n21387 ), .A2(_u10_n21388 ), .A3(_u10_n21389 ), .A4(_u10_n21390 ), .ZN(_u10_n21386 ) );
NOR4_X1 _u10_U10053  ( .A1(_u10_n21383 ), .A2(_u10_n21384 ), .A3(_u10_n21385 ), .A4(_u10_n21386 ), .ZN(_u10_n21382 ) );
NAND2_X1 _u10_U10052  ( .A1(_u10_n21381 ), .A2(_u10_n21382 ), .ZN(adr1[14]));
NAND2_X1 _u10_U10051  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21377 ) );
NAND2_X1 _u10_U10050  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21378 ) );
NAND2_X1 _u10_U10049  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21379 ) );
NAND2_X1 _u10_U10048  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21380 ) );
NAND4_X1 _u10_U10047  ( .A1(_u10_n21377 ), .A2(_u10_n21378 ), .A3(_u10_n21379 ), .A4(_u10_n21380 ), .ZN(_u10_n21362 ) );
NAND2_X1 _u10_U10046  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21373 ) );
NAND2_X1 _u10_U10045  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21374 ) );
NAND2_X1 _u10_U10044  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21375 ) );
NAND2_X1 _u10_U10043  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21376 ) );
NAND4_X1 _u10_U10042  ( .A1(_u10_n21373 ), .A2(_u10_n21374 ), .A3(_u10_n21375 ), .A4(_u10_n21376 ), .ZN(_u10_n21363 ) );
NAND2_X1 _u10_U10041  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21369 ) );
NAND2_X1 _u10_U10040  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21370 ) );
NAND2_X1 _u10_U10039  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21371 ) );
NAND2_X1 _u10_U10038  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21372 ) );
NAND4_X1 _u10_U10037  ( .A1(_u10_n21369 ), .A2(_u10_n21370 ), .A3(_u10_n21371 ), .A4(_u10_n21372 ), .ZN(_u10_n21364 ) );
NAND2_X1 _u10_U10036  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21366 ) );
NAND2_X1 _u10_U10035  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21367 ) );
NAND2_X1 _u10_U10034  ( .A1(ch0_adr1[15]), .A2(_u10_n12002 ), .ZN(_u10_n21368 ) );
NAND3_X1 _u10_U10033  ( .A1(_u10_n21366 ), .A2(_u10_n21367 ), .A3(_u10_n21368 ), .ZN(_u10_n21365 ) );
NOR4_X1 _u10_U10032  ( .A1(_u10_n21362 ), .A2(_u10_n21363 ), .A3(_u10_n21364 ), .A4(_u10_n21365 ), .ZN(_u10_n21340 ) );
NAND2_X1 _u10_U10031  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n21358 ) );
NAND2_X1 _u10_U10030  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n21359 ) );
NAND2_X1 _u10_U10029  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n21360 ) );
NAND2_X1 _u10_U10028  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n21361 ) );
NAND4_X1 _u10_U10027  ( .A1(_u10_n21358 ), .A2(_u10_n21359 ), .A3(_u10_n21360 ), .A4(_u10_n21361 ), .ZN(_u10_n21342 ) );
NAND2_X1 _u10_U10026  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n21354 ) );
NAND2_X1 _u10_U10025  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n21355 ) );
NAND2_X1 _u10_U10024  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n21356 ) );
NAND2_X1 _u10_U10023  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n21357 ) );
NAND4_X1 _u10_U10022  ( .A1(_u10_n21354 ), .A2(_u10_n21355 ), .A3(_u10_n21356 ), .A4(_u10_n21357 ), .ZN(_u10_n21343 ) );
NAND2_X1 _u10_U10021  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n21350 ) );
NAND2_X1 _u10_U10020  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n21351 ) );
NAND2_X1 _u10_U10019  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n21352 ) );
NAND2_X1 _u10_U10018  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n21353 ) );
NAND4_X1 _u10_U10017  ( .A1(_u10_n21350 ), .A2(_u10_n21351 ), .A3(_u10_n21352 ), .A4(_u10_n21353 ), .ZN(_u10_n21344 ) );
NAND2_X1 _u10_U10016  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n21346 ) );
NAND2_X1 _u10_U10015  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n21347 ) );
NAND2_X1 _u10_U10014  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n21348 ) );
NAND2_X1 _u10_U10013  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n21349 ) );
NAND4_X1 _u10_U10012  ( .A1(_u10_n21346 ), .A2(_u10_n21347 ), .A3(_u10_n21348 ), .A4(_u10_n21349 ), .ZN(_u10_n21345 ) );
NOR4_X1 _u10_U10011  ( .A1(_u10_n21342 ), .A2(_u10_n21343 ), .A3(_u10_n21344 ), .A4(_u10_n21345 ), .ZN(_u10_n21341 ) );
NAND2_X1 _u10_U10010  ( .A1(_u10_n21340 ), .A2(_u10_n21341 ), .ZN(adr1[15]));
NAND2_X1 _u10_U10009  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21336 ) );
NAND2_X1 _u10_U10008  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21337 ) );
NAND2_X1 _u10_U10007  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21338 ) );
NAND2_X1 _u10_U10006  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21339 ) );
NAND4_X1 _u10_U10005  ( .A1(_u10_n21336 ), .A2(_u10_n21337 ), .A3(_u10_n21338 ), .A4(_u10_n21339 ), .ZN(_u10_n21321 ) );
NAND2_X1 _u10_U10004  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21332 ) );
NAND2_X1 _u10_U10003  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21333 ) );
NAND2_X1 _u10_U10002  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21334 ) );
NAND2_X1 _u10_U10001  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21335 ) );
NAND4_X1 _u10_U10000  ( .A1(_u10_n21332 ), .A2(_u10_n21333 ), .A3(_u10_n21334 ), .A4(_u10_n21335 ), .ZN(_u10_n21322 ) );
NAND2_X1 _u10_U9999  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21328 ) );
NAND2_X1 _u10_U9998  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21329 ) );
NAND2_X1 _u10_U9997  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21330 ) );
NAND2_X1 _u10_U9996  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21331 ) );
NAND4_X1 _u10_U9995  ( .A1(_u10_n21328 ), .A2(_u10_n21329 ), .A3(_u10_n21330 ), .A4(_u10_n21331 ), .ZN(_u10_n21323 ) );
NAND2_X1 _u10_U9994  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21325 ) );
NAND2_X1 _u10_U9993  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21326 ) );
NAND2_X1 _u10_U9992  ( .A1(ch0_adr1[16]), .A2(_u10_n12002 ), .ZN(_u10_n21327 ) );
NAND3_X1 _u10_U9991  ( .A1(_u10_n21325 ), .A2(_u10_n21326 ), .A3(_u10_n21327 ), .ZN(_u10_n21324 ) );
NOR4_X1 _u10_U9990  ( .A1(_u10_n21321 ), .A2(_u10_n21322 ), .A3(_u10_n21323 ), .A4(_u10_n21324 ), .ZN(_u10_n21299 ) );
NAND2_X1 _u10_U9989  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n21317 ) );
NAND2_X1 _u10_U9988  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n21318 ) );
NAND2_X1 _u10_U9987  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n21319 ) );
NAND2_X1 _u10_U9986  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n21320 ) );
NAND4_X1 _u10_U9985  ( .A1(_u10_n21317 ), .A2(_u10_n21318 ), .A3(_u10_n21319 ), .A4(_u10_n21320 ), .ZN(_u10_n21301 ) );
NAND2_X1 _u10_U9984  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n21313 ) );
NAND2_X1 _u10_U9983  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n21314 ) );
NAND2_X1 _u10_U9982  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n21315 ) );
NAND2_X1 _u10_U9981  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n21316 ) );
NAND4_X1 _u10_U9980  ( .A1(_u10_n21313 ), .A2(_u10_n21314 ), .A3(_u10_n21315 ), .A4(_u10_n21316 ), .ZN(_u10_n21302 ) );
NAND2_X1 _u10_U9979  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n21309 ) );
NAND2_X1 _u10_U9978  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n21310 ) );
NAND2_X1 _u10_U9977  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n21311 ) );
NAND2_X1 _u10_U9976  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n21312 ) );
NAND4_X1 _u10_U9975  ( .A1(_u10_n21309 ), .A2(_u10_n21310 ), .A3(_u10_n21311 ), .A4(_u10_n21312 ), .ZN(_u10_n21303 ) );
NAND2_X1 _u10_U9974  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n21305 ) );
NAND2_X1 _u10_U9973  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n21306 ) );
NAND2_X1 _u10_U9972  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n21307 ) );
NAND2_X1 _u10_U9971  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n21308 ) );
NAND4_X1 _u10_U9970  ( .A1(_u10_n21305 ), .A2(_u10_n21306 ), .A3(_u10_n21307 ), .A4(_u10_n21308 ), .ZN(_u10_n21304 ) );
NOR4_X1 _u10_U9969  ( .A1(_u10_n21301 ), .A2(_u10_n21302 ), .A3(_u10_n21303 ), .A4(_u10_n21304 ), .ZN(_u10_n21300 ) );
NAND2_X1 _u10_U9968  ( .A1(_u10_n21299 ), .A2(_u10_n21300 ), .ZN(adr1[16]));
NAND2_X1 _u10_U9967  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21295 ) );
NAND2_X1 _u10_U9966  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21296 ) );
NAND2_X1 _u10_U9965  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21297 ) );
NAND2_X1 _u10_U9964  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21298 ) );
NAND4_X1 _u10_U9963  ( .A1(_u10_n21295 ), .A2(_u10_n21296 ), .A3(_u10_n21297 ), .A4(_u10_n21298 ), .ZN(_u10_n21280 ) );
NAND2_X1 _u10_U9962  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21291 ) );
NAND2_X1 _u10_U9961  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21292 ) );
NAND2_X1 _u10_U9960  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21293 ) );
NAND2_X1 _u10_U9959  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21294 ) );
NAND4_X1 _u10_U9958  ( .A1(_u10_n21291 ), .A2(_u10_n21292 ), .A3(_u10_n21293 ), .A4(_u10_n21294 ), .ZN(_u10_n21281 ) );
NAND2_X1 _u10_U9957  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21287 ) );
NAND2_X1 _u10_U9956  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21288 ) );
NAND2_X1 _u10_U9955  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21289 ) );
NAND2_X1 _u10_U9954  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21290 ) );
NAND4_X1 _u10_U9953  ( .A1(_u10_n21287 ), .A2(_u10_n21288 ), .A3(_u10_n21289 ), .A4(_u10_n21290 ), .ZN(_u10_n21282 ) );
NAND2_X1 _u10_U9952  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21284 ) );
NAND2_X1 _u10_U9951  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21285 ) );
NAND2_X1 _u10_U9950  ( .A1(ch0_adr1[17]), .A2(_u10_n12002 ), .ZN(_u10_n21286 ) );
NAND3_X1 _u10_U9949  ( .A1(_u10_n21284 ), .A2(_u10_n21285 ), .A3(_u10_n21286 ), .ZN(_u10_n21283 ) );
NOR4_X1 _u10_U9948  ( .A1(_u10_n21280 ), .A2(_u10_n21281 ), .A3(_u10_n21282 ), .A4(_u10_n21283 ), .ZN(_u10_n21258 ) );
NAND2_X1 _u10_U9947  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n21276 ) );
NAND2_X1 _u10_U9946  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n21277 ) );
NAND2_X1 _u10_U9945  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n21278 ) );
NAND2_X1 _u10_U9944  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n21279 ) );
NAND4_X1 _u10_U9943  ( .A1(_u10_n21276 ), .A2(_u10_n21277 ), .A3(_u10_n21278 ), .A4(_u10_n21279 ), .ZN(_u10_n21260 ) );
NAND2_X1 _u10_U9942  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n21272 ) );
NAND2_X1 _u10_U9941  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n21273 ) );
NAND2_X1 _u10_U9940  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n21274 ) );
NAND2_X1 _u10_U9939  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n21275 ) );
NAND4_X1 _u10_U9938  ( .A1(_u10_n21272 ), .A2(_u10_n21273 ), .A3(_u10_n21274 ), .A4(_u10_n21275 ), .ZN(_u10_n21261 ) );
NAND2_X1 _u10_U9937  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n21268 ) );
NAND2_X1 _u10_U9936  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n21269 ) );
NAND2_X1 _u10_U9935  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n21270 ) );
NAND2_X1 _u10_U9934  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n21271 ) );
NAND4_X1 _u10_U9933  ( .A1(_u10_n21268 ), .A2(_u10_n21269 ), .A3(_u10_n21270 ), .A4(_u10_n21271 ), .ZN(_u10_n21262 ) );
NAND2_X1 _u10_U9932  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n21264 ) );
NAND2_X1 _u10_U9931  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n21265 ) );
NAND2_X1 _u10_U9930  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n21266 ) );
NAND2_X1 _u10_U9929  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n21267 ) );
NAND4_X1 _u10_U9928  ( .A1(_u10_n21264 ), .A2(_u10_n21265 ), .A3(_u10_n21266 ), .A4(_u10_n21267 ), .ZN(_u10_n21263 ) );
NOR4_X1 _u10_U9927  ( .A1(_u10_n21260 ), .A2(_u10_n21261 ), .A3(_u10_n21262 ), .A4(_u10_n21263 ), .ZN(_u10_n21259 ) );
NAND2_X1 _u10_U9926  ( .A1(_u10_n21258 ), .A2(_u10_n21259 ), .ZN(adr1[17]));
NAND2_X1 _u10_U9925  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21254 ) );
NAND2_X1 _u10_U9924  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21255 ) );
NAND2_X1 _u10_U9923  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21256 ) );
NAND2_X1 _u10_U9922  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21257 ) );
NAND4_X1 _u10_U9921  ( .A1(_u10_n21254 ), .A2(_u10_n21255 ), .A3(_u10_n21256 ), .A4(_u10_n21257 ), .ZN(_u10_n21239 ) );
NAND2_X1 _u10_U9920  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21250 ) );
NAND2_X1 _u10_U9919  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21251 ) );
NAND2_X1 _u10_U9918  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21252 ) );
NAND2_X1 _u10_U9917  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21253 ) );
NAND4_X1 _u10_U9916  ( .A1(_u10_n21250 ), .A2(_u10_n21251 ), .A3(_u10_n21252 ), .A4(_u10_n21253 ), .ZN(_u10_n21240 ) );
NAND2_X1 _u10_U9915  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21246 ) );
NAND2_X1 _u10_U9914  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21247 ) );
NAND2_X1 _u10_U9913  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21248 ) );
NAND2_X1 _u10_U9912  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21249 ) );
NAND4_X1 _u10_U9911  ( .A1(_u10_n21246 ), .A2(_u10_n21247 ), .A3(_u10_n21248 ), .A4(_u10_n21249 ), .ZN(_u10_n21241 ) );
NAND2_X1 _u10_U9910  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21243 ) );
NAND2_X1 _u10_U9909  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21244 ) );
NAND2_X1 _u10_U9908  ( .A1(ch0_adr1[18]), .A2(_u10_n12002 ), .ZN(_u10_n21245 ) );
NAND3_X1 _u10_U9907  ( .A1(_u10_n21243 ), .A2(_u10_n21244 ), .A3(_u10_n21245 ), .ZN(_u10_n21242 ) );
NOR4_X1 _u10_U9906  ( .A1(_u10_n21239 ), .A2(_u10_n21240 ), .A3(_u10_n21241 ), .A4(_u10_n21242 ), .ZN(_u10_n21217 ) );
NAND2_X1 _u10_U9905  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n21235 ) );
NAND2_X1 _u10_U9904  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n21236 ) );
NAND2_X1 _u10_U9903  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n21237 ) );
NAND2_X1 _u10_U9902  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n21238 ) );
NAND4_X1 _u10_U9901  ( .A1(_u10_n21235 ), .A2(_u10_n21236 ), .A3(_u10_n21237 ), .A4(_u10_n21238 ), .ZN(_u10_n21219 ) );
NAND2_X1 _u10_U9900  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n21231 ) );
NAND2_X1 _u10_U9899  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n21232 ) );
NAND2_X1 _u10_U9898  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n21233 ) );
NAND2_X1 _u10_U9897  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n21234 ) );
NAND4_X1 _u10_U9896  ( .A1(_u10_n21231 ), .A2(_u10_n21232 ), .A3(_u10_n21233 ), .A4(_u10_n21234 ), .ZN(_u10_n21220 ) );
NAND2_X1 _u10_U9895  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n21227 ) );
NAND2_X1 _u10_U9894  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n21228 ) );
NAND2_X1 _u10_U9893  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n21229 ) );
NAND2_X1 _u10_U9892  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n21230 ) );
NAND4_X1 _u10_U9891  ( .A1(_u10_n21227 ), .A2(_u10_n21228 ), .A3(_u10_n21229 ), .A4(_u10_n21230 ), .ZN(_u10_n21221 ) );
NAND2_X1 _u10_U9890  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n21223 ) );
NAND2_X1 _u10_U9889  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n21224 ) );
NAND2_X1 _u10_U9888  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n21225 ) );
NAND2_X1 _u10_U9887  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n21226 ) );
NAND4_X1 _u10_U9886  ( .A1(_u10_n21223 ), .A2(_u10_n21224 ), .A3(_u10_n21225 ), .A4(_u10_n21226 ), .ZN(_u10_n21222 ) );
NOR4_X1 _u10_U9885  ( .A1(_u10_n21219 ), .A2(_u10_n21220 ), .A3(_u10_n21221 ), .A4(_u10_n21222 ), .ZN(_u10_n21218 ) );
NAND2_X1 _u10_U9884  ( .A1(_u10_n21217 ), .A2(_u10_n21218 ), .ZN(adr1[18]));
NAND2_X1 _u10_U9883  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21213 ) );
NAND2_X1 _u10_U9882  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21214 ) );
NAND2_X1 _u10_U9881  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21215 ) );
NAND2_X1 _u10_U9880  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21216 ) );
NAND4_X1 _u10_U9879  ( .A1(_u10_n21213 ), .A2(_u10_n21214 ), .A3(_u10_n21215 ), .A4(_u10_n21216 ), .ZN(_u10_n21198 ) );
NAND2_X1 _u10_U9878  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21209 ) );
NAND2_X1 _u10_U9877  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21210 ) );
NAND2_X1 _u10_U9876  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21211 ) );
NAND2_X1 _u10_U9875  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21212 ) );
NAND4_X1 _u10_U9874  ( .A1(_u10_n21209 ), .A2(_u10_n21210 ), .A3(_u10_n21211 ), .A4(_u10_n21212 ), .ZN(_u10_n21199 ) );
NAND2_X1 _u10_U9873  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21205 ) );
NAND2_X1 _u10_U9872  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21206 ) );
NAND2_X1 _u10_U9871  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21207 ) );
NAND2_X1 _u10_U9870  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21208 ) );
NAND4_X1 _u10_U9869  ( .A1(_u10_n21205 ), .A2(_u10_n21206 ), .A3(_u10_n21207 ), .A4(_u10_n21208 ), .ZN(_u10_n21200 ) );
NAND2_X1 _u10_U9868  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21202 ) );
NAND2_X1 _u10_U9867  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21203 ) );
NAND2_X1 _u10_U9866  ( .A1(ch0_adr1[19]), .A2(_u10_n12002 ), .ZN(_u10_n21204 ) );
NAND3_X1 _u10_U9865  ( .A1(_u10_n21202 ), .A2(_u10_n21203 ), .A3(_u10_n21204 ), .ZN(_u10_n21201 ) );
NOR4_X1 _u10_U9864  ( .A1(_u10_n21198 ), .A2(_u10_n21199 ), .A3(_u10_n21200 ), .A4(_u10_n21201 ), .ZN(_u10_n21176 ) );
NAND2_X1 _u10_U9863  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n21194 ) );
NAND2_X1 _u10_U9862  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n21195 ) );
NAND2_X1 _u10_U9861  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n21196 ) );
NAND2_X1 _u10_U9860  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n21197 ) );
NAND4_X1 _u10_U9859  ( .A1(_u10_n21194 ), .A2(_u10_n21195 ), .A3(_u10_n21196 ), .A4(_u10_n21197 ), .ZN(_u10_n21178 ) );
NAND2_X1 _u10_U9858  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n21190 ) );
NAND2_X1 _u10_U9857  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n21191 ) );
NAND2_X1 _u10_U9856  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n21192 ) );
NAND2_X1 _u10_U9855  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n21193 ) );
NAND4_X1 _u10_U9854  ( .A1(_u10_n21190 ), .A2(_u10_n21191 ), .A3(_u10_n21192 ), .A4(_u10_n21193 ), .ZN(_u10_n21179 ) );
NAND2_X1 _u10_U9853  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n21186 ) );
NAND2_X1 _u10_U9852  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n21187 ) );
NAND2_X1 _u10_U9851  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n21188 ) );
NAND2_X1 _u10_U9850  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n21189 ) );
NAND4_X1 _u10_U9849  ( .A1(_u10_n21186 ), .A2(_u10_n21187 ), .A3(_u10_n21188 ), .A4(_u10_n21189 ), .ZN(_u10_n21180 ) );
NAND2_X1 _u10_U9848  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n21182 ) );
NAND2_X1 _u10_U9847  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n21183 ) );
NAND2_X1 _u10_U9846  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n21184 ) );
NAND2_X1 _u10_U9845  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n21185 ) );
NAND4_X1 _u10_U9844  ( .A1(_u10_n21182 ), .A2(_u10_n21183 ), .A3(_u10_n21184 ), .A4(_u10_n21185 ), .ZN(_u10_n21181 ) );
NOR4_X1 _u10_U9843  ( .A1(_u10_n21178 ), .A2(_u10_n21179 ), .A3(_u10_n21180 ), .A4(_u10_n21181 ), .ZN(_u10_n21177 ) );
NAND2_X1 _u10_U9842  ( .A1(_u10_n21176 ), .A2(_u10_n21177 ), .ZN(adr1[19]));
NAND2_X1 _u10_U9841  ( .A1(1'b0), .A2(_u10_n12333 ), .ZN(_u10_n21172 ) );
NAND2_X1 _u10_U9840  ( .A1(1'b0), .A2(_u10_n12309 ), .ZN(_u10_n21173 ) );
NAND2_X1 _u10_U9839  ( .A1(1'b0), .A2(_u10_n12285 ), .ZN(_u10_n21174 ) );
NAND2_X1 _u10_U9838  ( .A1(1'b0), .A2(_u10_n12261 ), .ZN(_u10_n21175 ) );
NAND4_X1 _u10_U9837  ( .A1(_u10_n21172 ), .A2(_u10_n21173 ), .A3(_u10_n21174 ), .A4(_u10_n21175 ), .ZN(_u10_n21157 ) );
NAND2_X1 _u10_U9836  ( .A1(1'b0), .A2(_u10_n12237 ), .ZN(_u10_n21168 ) );
NAND2_X1 _u10_U9835  ( .A1(1'b0), .A2(_u10_n12213 ), .ZN(_u10_n21169 ) );
NAND2_X1 _u10_U9834  ( .A1(1'b0), .A2(_u10_n12189 ), .ZN(_u10_n21170 ) );
NAND2_X1 _u10_U9833  ( .A1(1'b0), .A2(_u10_n12165 ), .ZN(_u10_n21171 ) );
NAND4_X1 _u10_U9832  ( .A1(_u10_n21168 ), .A2(_u10_n21169 ), .A3(_u10_n21170 ), .A4(_u10_n21171 ), .ZN(_u10_n21158 ) );
NAND2_X1 _u10_U9831  ( .A1(1'b0), .A2(_u10_n12141 ), .ZN(_u10_n21164 ) );
NAND2_X1 _u10_U9830  ( .A1(1'b0), .A2(_u10_n12117 ), .ZN(_u10_n21165 ) );
NAND2_X1 _u10_U9829  ( .A1(1'b0), .A2(_u10_n12093 ), .ZN(_u10_n21166 ) );
NAND2_X1 _u10_U9828  ( .A1(1'b0), .A2(_u10_n12069 ), .ZN(_u10_n21167 ) );
NAND4_X1 _u10_U9827  ( .A1(_u10_n21164 ), .A2(_u10_n21165 ), .A3(_u10_n21166 ), .A4(_u10_n21167 ), .ZN(_u10_n21159 ) );
NAND2_X1 _u10_U9826  ( .A1(1'b0), .A2(_u10_n12045 ), .ZN(_u10_n21161 ) );
NAND2_X1 _u10_U9825  ( .A1(1'b0), .A2(_u10_n12021 ), .ZN(_u10_n21162 ) );
NAND2_X1 _u10_U9824  ( .A1(1'b0), .A2(_u10_n12002 ), .ZN(_u10_n21163 ) );
NAND3_X1 _u10_U9823  ( .A1(_u10_n21161 ), .A2(_u10_n21162 ), .A3(_u10_n21163 ), .ZN(_u10_n21160 ) );
NOR4_X1 _u10_U9822  ( .A1(_u10_n21157 ), .A2(_u10_n21158 ), .A3(_u10_n21159 ), .A4(_u10_n21160 ), .ZN(_u10_n21135 ) );
NAND2_X1 _u10_U9821  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n21153 ) );
NAND2_X1 _u10_U9820  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n21154 ) );
NAND2_X1 _u10_U9819  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n21155 ) );
NAND2_X1 _u10_U9818  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n21156 ) );
NAND4_X1 _u10_U9817  ( .A1(_u10_n21153 ), .A2(_u10_n21154 ), .A3(_u10_n21155 ), .A4(_u10_n21156 ), .ZN(_u10_n21137 ) );
NAND2_X1 _u10_U9816  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n21149 ) );
NAND2_X1 _u10_U9815  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n21150 ) );
NAND2_X1 _u10_U9814  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n21151 ) );
NAND2_X1 _u10_U9813  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n21152 ) );
NAND4_X1 _u10_U9812  ( .A1(_u10_n21149 ), .A2(_u10_n21150 ), .A3(_u10_n21151 ), .A4(_u10_n21152 ), .ZN(_u10_n21138 ) );
NAND2_X1 _u10_U9811  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n21145 ) );
NAND2_X1 _u10_U9810  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n21146 ) );
NAND2_X1 _u10_U9809  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n21147 ) );
NAND2_X1 _u10_U9808  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n21148 ) );
NAND4_X1 _u10_U9807  ( .A1(_u10_n21145 ), .A2(_u10_n21146 ), .A3(_u10_n21147 ), .A4(_u10_n21148 ), .ZN(_u10_n21139 ) );
NAND2_X1 _u10_U9806  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n21141 ) );
NAND2_X1 _u10_U9805  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n21142 ) );
NAND2_X1 _u10_U9804  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n21143 ) );
NAND2_X1 _u10_U9803  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n21144 ) );
NAND4_X1 _u10_U9802  ( .A1(_u10_n21141 ), .A2(_u10_n21142 ), .A3(_u10_n21143 ), .A4(_u10_n21144 ), .ZN(_u10_n21140 ) );
NOR4_X1 _u10_U9801  ( .A1(_u10_n21137 ), .A2(_u10_n21138 ), .A3(_u10_n21139 ), .A4(_u10_n21140 ), .ZN(_u10_n21136 ) );
NAND2_X1 _u10_U9800  ( .A1(_u10_n21135 ), .A2(_u10_n21136 ), .ZN(adr1[1]) );
NAND2_X1 _u10_U9799  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n21131 ) );
NAND2_X1 _u10_U9798  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n21132 ) );
NAND2_X1 _u10_U9797  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n21133 ) );
NAND2_X1 _u10_U9796  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n21134 ) );
NAND4_X1 _u10_U9795  ( .A1(_u10_n21131 ), .A2(_u10_n21132 ), .A3(_u10_n21133 ), .A4(_u10_n21134 ), .ZN(_u10_n21116 ) );
NAND2_X1 _u10_U9794  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n21127 ) );
NAND2_X1 _u10_U9793  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n21128 ) );
NAND2_X1 _u10_U9792  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n21129 ) );
NAND2_X1 _u10_U9791  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n21130 ) );
NAND4_X1 _u10_U9790  ( .A1(_u10_n21127 ), .A2(_u10_n21128 ), .A3(_u10_n21129 ), .A4(_u10_n21130 ), .ZN(_u10_n21117 ) );
NAND2_X1 _u10_U9789  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n21123 ) );
NAND2_X1 _u10_U9788  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n21124 ) );
NAND2_X1 _u10_U9787  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n21125 ) );
NAND2_X1 _u10_U9786  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n21126 ) );
NAND4_X1 _u10_U9785  ( .A1(_u10_n21123 ), .A2(_u10_n21124 ), .A3(_u10_n21125 ), .A4(_u10_n21126 ), .ZN(_u10_n21118 ) );
NAND2_X1 _u10_U9784  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n21120 ) );
NAND2_X1 _u10_U9783  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n21121 ) );
NAND2_X1 _u10_U9782  ( .A1(ch0_adr1[20]), .A2(_u10_n12002 ), .ZN(_u10_n21122 ) );
NAND3_X1 _u10_U9781  ( .A1(_u10_n21120 ), .A2(_u10_n21121 ), .A3(_u10_n21122 ), .ZN(_u10_n21119 ) );
NOR4_X1 _u10_U9780  ( .A1(_u10_n21116 ), .A2(_u10_n21117 ), .A3(_u10_n21118 ), .A4(_u10_n21119 ), .ZN(_u10_n21094 ) );
NAND2_X1 _u10_U9779  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n21112 ) );
NAND2_X1 _u10_U9778  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n21113 ) );
NAND2_X1 _u10_U9777  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n21114 ) );
NAND2_X1 _u10_U9776  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n21115 ) );
NAND4_X1 _u10_U9775  ( .A1(_u10_n21112 ), .A2(_u10_n21113 ), .A3(_u10_n21114 ), .A4(_u10_n21115 ), .ZN(_u10_n21096 ) );
NAND2_X1 _u10_U9774  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n21108 ) );
NAND2_X1 _u10_U9773  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n21109 ) );
NAND2_X1 _u10_U9772  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n21110 ) );
NAND2_X1 _u10_U9771  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n21111 ) );
NAND4_X1 _u10_U9770  ( .A1(_u10_n21108 ), .A2(_u10_n21109 ), .A3(_u10_n21110 ), .A4(_u10_n21111 ), .ZN(_u10_n21097 ) );
NAND2_X1 _u10_U9769  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n21104 ) );
NAND2_X1 _u10_U9768  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n21105 ) );
NAND2_X1 _u10_U9767  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n21106 ) );
NAND2_X1 _u10_U9766  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n21107 ) );
NAND4_X1 _u10_U9765  ( .A1(_u10_n21104 ), .A2(_u10_n21105 ), .A3(_u10_n21106 ), .A4(_u10_n21107 ), .ZN(_u10_n21098 ) );
NAND2_X1 _u10_U9764  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n21100 ) );
NAND2_X1 _u10_U9763  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n21101 ) );
NAND2_X1 _u10_U9762  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n21102 ) );
NAND2_X1 _u10_U9761  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n21103 ) );
NAND4_X1 _u10_U9760  ( .A1(_u10_n21100 ), .A2(_u10_n21101 ), .A3(_u10_n21102 ), .A4(_u10_n21103 ), .ZN(_u10_n21099 ) );
NOR4_X1 _u10_U9759  ( .A1(_u10_n21096 ), .A2(_u10_n21097 ), .A3(_u10_n21098 ), .A4(_u10_n21099 ), .ZN(_u10_n21095 ) );
NAND2_X1 _u10_U9758  ( .A1(_u10_n21094 ), .A2(_u10_n21095 ), .ZN(adr1[20]));
NAND2_X1 _u10_U9757  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n21090 ) );
NAND2_X1 _u10_U9756  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n21091 ) );
NAND2_X1 _u10_U9755  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n21092 ) );
NAND2_X1 _u10_U9754  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n21093 ) );
NAND4_X1 _u10_U9753  ( .A1(_u10_n21090 ), .A2(_u10_n21091 ), .A3(_u10_n21092 ), .A4(_u10_n21093 ), .ZN(_u10_n21075 ) );
NAND2_X1 _u10_U9752  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n21086 ) );
NAND2_X1 _u10_U9751  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n21087 ) );
NAND2_X1 _u10_U9750  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n21088 ) );
NAND2_X1 _u10_U9749  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n21089 ) );
NAND4_X1 _u10_U9748  ( .A1(_u10_n21086 ), .A2(_u10_n21087 ), .A3(_u10_n21088 ), .A4(_u10_n21089 ), .ZN(_u10_n21076 ) );
NAND2_X1 _u10_U9747  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n21082 ) );
NAND2_X1 _u10_U9746  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n21083 ) );
NAND2_X1 _u10_U9745  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n21084 ) );
NAND2_X1 _u10_U9744  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n21085 ) );
NAND4_X1 _u10_U9743  ( .A1(_u10_n21082 ), .A2(_u10_n21083 ), .A3(_u10_n21084 ), .A4(_u10_n21085 ), .ZN(_u10_n21077 ) );
NAND2_X1 _u10_U9742  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n21079 ) );
NAND2_X1 _u10_U9741  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n21080 ) );
NAND2_X1 _u10_U9740  ( .A1(ch0_adr1[21]), .A2(_u10_n12002 ), .ZN(_u10_n21081 ) );
NAND3_X1 _u10_U9739  ( .A1(_u10_n21079 ), .A2(_u10_n21080 ), .A3(_u10_n21081 ), .ZN(_u10_n21078 ) );
NOR4_X1 _u10_U9738  ( .A1(_u10_n21075 ), .A2(_u10_n21076 ), .A3(_u10_n21077 ), .A4(_u10_n21078 ), .ZN(_u10_n21053 ) );
NAND2_X1 _u10_U9737  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n21071 ) );
NAND2_X1 _u10_U9736  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n21072 ) );
NAND2_X1 _u10_U9735  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n21073 ) );
NAND2_X1 _u10_U9734  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n21074 ) );
NAND4_X1 _u10_U9733  ( .A1(_u10_n21071 ), .A2(_u10_n21072 ), .A3(_u10_n21073 ), .A4(_u10_n21074 ), .ZN(_u10_n21055 ) );
NAND2_X1 _u10_U9732  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n21067 ) );
NAND2_X1 _u10_U9731  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n21068 ) );
NAND2_X1 _u10_U9730  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n21069 ) );
NAND2_X1 _u10_U9729  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n21070 ) );
NAND4_X1 _u10_U9728  ( .A1(_u10_n21067 ), .A2(_u10_n21068 ), .A3(_u10_n21069 ), .A4(_u10_n21070 ), .ZN(_u10_n21056 ) );
NAND2_X1 _u10_U9727  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n21063 ) );
NAND2_X1 _u10_U9726  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n21064 ) );
NAND2_X1 _u10_U9725  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n21065 ) );
NAND2_X1 _u10_U9724  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n21066 ) );
NAND4_X1 _u10_U9723  ( .A1(_u10_n21063 ), .A2(_u10_n21064 ), .A3(_u10_n21065 ), .A4(_u10_n21066 ), .ZN(_u10_n21057 ) );
NAND2_X1 _u10_U9722  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n21059 ) );
NAND2_X1 _u10_U9721  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n21060 ) );
NAND2_X1 _u10_U9720  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n21061 ) );
NAND2_X1 _u10_U9719  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n21062 ) );
NAND4_X1 _u10_U9718  ( .A1(_u10_n21059 ), .A2(_u10_n21060 ), .A3(_u10_n21061 ), .A4(_u10_n21062 ), .ZN(_u10_n21058 ) );
NOR4_X1 _u10_U9717  ( .A1(_u10_n21055 ), .A2(_u10_n21056 ), .A3(_u10_n21057 ), .A4(_u10_n21058 ), .ZN(_u10_n21054 ) );
NAND2_X1 _u10_U9716  ( .A1(_u10_n21053 ), .A2(_u10_n21054 ), .ZN(adr1[21]));
NAND2_X1 _u10_U9715  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n21049 ) );
NAND2_X1 _u10_U9714  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n21050 ) );
NAND2_X1 _u10_U9713  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n21051 ) );
NAND2_X1 _u10_U9712  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n21052 ) );
NAND4_X1 _u10_U9711  ( .A1(_u10_n21049 ), .A2(_u10_n21050 ), .A3(_u10_n21051 ), .A4(_u10_n21052 ), .ZN(_u10_n21034 ) );
NAND2_X1 _u10_U9710  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n21045 ) );
NAND2_X1 _u10_U9709  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n21046 ) );
NAND2_X1 _u10_U9708  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n21047 ) );
NAND2_X1 _u10_U9707  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n21048 ) );
NAND4_X1 _u10_U9706  ( .A1(_u10_n21045 ), .A2(_u10_n21046 ), .A3(_u10_n21047 ), .A4(_u10_n21048 ), .ZN(_u10_n21035 ) );
NAND2_X1 _u10_U9705  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n21041 ) );
NAND2_X1 _u10_U9704  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n21042 ) );
NAND2_X1 _u10_U9703  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n21043 ) );
NAND2_X1 _u10_U9702  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n21044 ) );
NAND4_X1 _u10_U9701  ( .A1(_u10_n21041 ), .A2(_u10_n21042 ), .A3(_u10_n21043 ), .A4(_u10_n21044 ), .ZN(_u10_n21036 ) );
NAND2_X1 _u10_U9700  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n21038 ) );
NAND2_X1 _u10_U9699  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n21039 ) );
NAND2_X1 _u10_U9698  ( .A1(ch0_adr1[22]), .A2(_u10_n12002 ), .ZN(_u10_n21040 ) );
NAND3_X1 _u10_U9697  ( .A1(_u10_n21038 ), .A2(_u10_n21039 ), .A3(_u10_n21040 ), .ZN(_u10_n21037 ) );
NOR4_X1 _u10_U9696  ( .A1(_u10_n21034 ), .A2(_u10_n21035 ), .A3(_u10_n21036 ), .A4(_u10_n21037 ), .ZN(_u10_n21012 ) );
NAND2_X1 _u10_U9695  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n21030 ) );
NAND2_X1 _u10_U9694  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n21031 ) );
NAND2_X1 _u10_U9693  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n21032 ) );
NAND2_X1 _u10_U9692  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n21033 ) );
NAND4_X1 _u10_U9691  ( .A1(_u10_n21030 ), .A2(_u10_n21031 ), .A3(_u10_n21032 ), .A4(_u10_n21033 ), .ZN(_u10_n21014 ) );
NAND2_X1 _u10_U9690  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n21026 ) );
NAND2_X1 _u10_U9689  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n21027 ) );
NAND2_X1 _u10_U9688  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n21028 ) );
NAND2_X1 _u10_U9687  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n21029 ) );
NAND4_X1 _u10_U9686  ( .A1(_u10_n21026 ), .A2(_u10_n21027 ), .A3(_u10_n21028 ), .A4(_u10_n21029 ), .ZN(_u10_n21015 ) );
NAND2_X1 _u10_U9685  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n21022 ) );
NAND2_X1 _u10_U9684  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n21023 ) );
NAND2_X1 _u10_U9683  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n21024 ) );
NAND2_X1 _u10_U9682  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n21025 ) );
NAND4_X1 _u10_U9681  ( .A1(_u10_n21022 ), .A2(_u10_n21023 ), .A3(_u10_n21024 ), .A4(_u10_n21025 ), .ZN(_u10_n21016 ) );
NAND2_X1 _u10_U9680  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n21018 ) );
NAND2_X1 _u10_U9679  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n21019 ) );
NAND2_X1 _u10_U9678  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n21020 ) );
NAND2_X1 _u10_U9677  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n21021 ) );
NAND4_X1 _u10_U9676  ( .A1(_u10_n21018 ), .A2(_u10_n21019 ), .A3(_u10_n21020 ), .A4(_u10_n21021 ), .ZN(_u10_n21017 ) );
NOR4_X1 _u10_U9675  ( .A1(_u10_n21014 ), .A2(_u10_n21015 ), .A3(_u10_n21016 ), .A4(_u10_n21017 ), .ZN(_u10_n21013 ) );
NAND2_X1 _u10_U9674  ( .A1(_u10_n21012 ), .A2(_u10_n21013 ), .ZN(adr1[22]));
NAND2_X1 _u10_U9673  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n21008 ) );
NAND2_X1 _u10_U9672  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n21009 ) );
NAND2_X1 _u10_U9671  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n21010 ) );
NAND2_X1 _u10_U9670  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n21011 ) );
NAND4_X1 _u10_U9669  ( .A1(_u10_n21008 ), .A2(_u10_n21009 ), .A3(_u10_n21010 ), .A4(_u10_n21011 ), .ZN(_u10_n20993 ) );
NAND2_X1 _u10_U9668  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n21004 ) );
NAND2_X1 _u10_U9667  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n21005 ) );
NAND2_X1 _u10_U9666  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n21006 ) );
NAND2_X1 _u10_U9665  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n21007 ) );
NAND4_X1 _u10_U9664  ( .A1(_u10_n21004 ), .A2(_u10_n21005 ), .A3(_u10_n21006 ), .A4(_u10_n21007 ), .ZN(_u10_n20994 ) );
NAND2_X1 _u10_U9663  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n21000 ) );
NAND2_X1 _u10_U9662  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n21001 ) );
NAND2_X1 _u10_U9661  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n21002 ) );
NAND2_X1 _u10_U9660  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n21003 ) );
NAND4_X1 _u10_U9659  ( .A1(_u10_n21000 ), .A2(_u10_n21001 ), .A3(_u10_n21002 ), .A4(_u10_n21003 ), .ZN(_u10_n20995 ) );
NAND2_X1 _u10_U9658  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n20997 ) );
NAND2_X1 _u10_U9657  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n20998 ) );
NAND2_X1 _u10_U9656  ( .A1(ch0_adr1[23]), .A2(_u10_n12003 ), .ZN(_u10_n20999 ) );
NAND3_X1 _u10_U9655  ( .A1(_u10_n20997 ), .A2(_u10_n20998 ), .A3(_u10_n20999 ), .ZN(_u10_n20996 ) );
NOR4_X1 _u10_U9654  ( .A1(_u10_n20993 ), .A2(_u10_n20994 ), .A3(_u10_n20995 ), .A4(_u10_n20996 ), .ZN(_u10_n20971 ) );
NAND2_X1 _u10_U9653  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n20989 ) );
NAND2_X1 _u10_U9652  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n20990 ) );
NAND2_X1 _u10_U9651  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n20991 ) );
NAND2_X1 _u10_U9650  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n20992 ) );
NAND4_X1 _u10_U9649  ( .A1(_u10_n20989 ), .A2(_u10_n20990 ), .A3(_u10_n20991 ), .A4(_u10_n20992 ), .ZN(_u10_n20973 ) );
NAND2_X1 _u10_U9648  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n20985 ) );
NAND2_X1 _u10_U9647  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n20986 ) );
NAND2_X1 _u10_U9646  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n20987 ) );
NAND2_X1 _u10_U9645  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n20988 ) );
NAND4_X1 _u10_U9644  ( .A1(_u10_n20985 ), .A2(_u10_n20986 ), .A3(_u10_n20987 ), .A4(_u10_n20988 ), .ZN(_u10_n20974 ) );
NAND2_X1 _u10_U9643  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n20981 ) );
NAND2_X1 _u10_U9642  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n20982 ) );
NAND2_X1 _u10_U9641  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n20983 ) );
NAND2_X1 _u10_U9640  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n20984 ) );
NAND4_X1 _u10_U9639  ( .A1(_u10_n20981 ), .A2(_u10_n20982 ), .A3(_u10_n20983 ), .A4(_u10_n20984 ), .ZN(_u10_n20975 ) );
NAND2_X1 _u10_U9638  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n20977 ) );
NAND2_X1 _u10_U9637  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n20978 ) );
NAND2_X1 _u10_U9636  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n20979 ) );
NAND2_X1 _u10_U9635  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n20980 ) );
NAND4_X1 _u10_U9634  ( .A1(_u10_n20977 ), .A2(_u10_n20978 ), .A3(_u10_n20979 ), .A4(_u10_n20980 ), .ZN(_u10_n20976 ) );
NOR4_X1 _u10_U9633  ( .A1(_u10_n20973 ), .A2(_u10_n20974 ), .A3(_u10_n20975 ), .A4(_u10_n20976 ), .ZN(_u10_n20972 ) );
NAND2_X1 _u10_U9632  ( .A1(_u10_n20971 ), .A2(_u10_n20972 ), .ZN(adr1[23]));
NAND2_X1 _u10_U9631  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n20967 ) );
NAND2_X1 _u10_U9630  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n20968 ) );
NAND2_X1 _u10_U9629  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n20969 ) );
NAND2_X1 _u10_U9628  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n20970 ) );
NAND4_X1 _u10_U9627  ( .A1(_u10_n20967 ), .A2(_u10_n20968 ), .A3(_u10_n20969 ), .A4(_u10_n20970 ), .ZN(_u10_n20952 ) );
NAND2_X1 _u10_U9626  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n20963 ) );
NAND2_X1 _u10_U9625  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n20964 ) );
NAND2_X1 _u10_U9624  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n20965 ) );
NAND2_X1 _u10_U9623  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n20966 ) );
NAND4_X1 _u10_U9622  ( .A1(_u10_n20963 ), .A2(_u10_n20964 ), .A3(_u10_n20965 ), .A4(_u10_n20966 ), .ZN(_u10_n20953 ) );
NAND2_X1 _u10_U9621  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n20959 ) );
NAND2_X1 _u10_U9620  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n20960 ) );
NAND2_X1 _u10_U9619  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n20961 ) );
NAND2_X1 _u10_U9618  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n20962 ) );
NAND4_X1 _u10_U9617  ( .A1(_u10_n20959 ), .A2(_u10_n20960 ), .A3(_u10_n20961 ), .A4(_u10_n20962 ), .ZN(_u10_n20954 ) );
NAND2_X1 _u10_U9616  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n20956 ) );
NAND2_X1 _u10_U9615  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n20957 ) );
NAND2_X1 _u10_U9614  ( .A1(ch0_adr1[24]), .A2(_u10_n12003 ), .ZN(_u10_n20958 ) );
NAND3_X1 _u10_U9613  ( .A1(_u10_n20956 ), .A2(_u10_n20957 ), .A3(_u10_n20958 ), .ZN(_u10_n20955 ) );
NOR4_X1 _u10_U9612  ( .A1(_u10_n20952 ), .A2(_u10_n20953 ), .A3(_u10_n20954 ), .A4(_u10_n20955 ), .ZN(_u10_n20930 ) );
NAND2_X1 _u10_U9611  ( .A1(1'b0), .A2(_u10_n11986 ), .ZN(_u10_n20948 ) );
NAND2_X1 _u10_U9610  ( .A1(1'b0), .A2(_u10_n11962 ), .ZN(_u10_n20949 ) );
NAND2_X1 _u10_U9609  ( .A1(1'b0), .A2(_u10_n11938 ), .ZN(_u10_n20950 ) );
NAND2_X1 _u10_U9608  ( .A1(1'b0), .A2(_u10_n11914 ), .ZN(_u10_n20951 ) );
NAND4_X1 _u10_U9607  ( .A1(_u10_n20948 ), .A2(_u10_n20949 ), .A3(_u10_n20950 ), .A4(_u10_n20951 ), .ZN(_u10_n20932 ) );
NAND2_X1 _u10_U9606  ( .A1(1'b0), .A2(_u10_n11890 ), .ZN(_u10_n20944 ) );
NAND2_X1 _u10_U9605  ( .A1(1'b0), .A2(_u10_n11866 ), .ZN(_u10_n20945 ) );
NAND2_X1 _u10_U9604  ( .A1(1'b0), .A2(_u10_n11842 ), .ZN(_u10_n20946 ) );
NAND2_X1 _u10_U9603  ( .A1(1'b0), .A2(_u10_n11818 ), .ZN(_u10_n20947 ) );
NAND4_X1 _u10_U9602  ( .A1(_u10_n20944 ), .A2(_u10_n20945 ), .A3(_u10_n20946 ), .A4(_u10_n20947 ), .ZN(_u10_n20933 ) );
NAND2_X1 _u10_U9601  ( .A1(1'b0), .A2(_u10_n11794 ), .ZN(_u10_n20940 ) );
NAND2_X1 _u10_U9600  ( .A1(1'b0), .A2(_u10_n11770 ), .ZN(_u10_n20941 ) );
NAND2_X1 _u10_U9599  ( .A1(1'b0), .A2(_u10_n11746 ), .ZN(_u10_n20942 ) );
NAND2_X1 _u10_U9598  ( .A1(1'b0), .A2(_u10_n11722 ), .ZN(_u10_n20943 ) );
NAND4_X1 _u10_U9597  ( .A1(_u10_n20940 ), .A2(_u10_n20941 ), .A3(_u10_n20942 ), .A4(_u10_n20943 ), .ZN(_u10_n20934 ) );
NAND2_X1 _u10_U9596  ( .A1(1'b0), .A2(_u10_n11698 ), .ZN(_u10_n20936 ) );
NAND2_X1 _u10_U9595  ( .A1(1'b0), .A2(_u10_n11674 ), .ZN(_u10_n20937 ) );
NAND2_X1 _u10_U9594  ( .A1(1'b0), .A2(_u10_n11650 ), .ZN(_u10_n20938 ) );
NAND2_X1 _u10_U9593  ( .A1(1'b0), .A2(_u10_n11626 ), .ZN(_u10_n20939 ) );
NAND4_X1 _u10_U9592  ( .A1(_u10_n20936 ), .A2(_u10_n20937 ), .A3(_u10_n20938 ), .A4(_u10_n20939 ), .ZN(_u10_n20935 ) );
NOR4_X1 _u10_U9591  ( .A1(_u10_n20932 ), .A2(_u10_n20933 ), .A3(_u10_n20934 ), .A4(_u10_n20935 ), .ZN(_u10_n20931 ) );
NAND2_X1 _u10_U9590  ( .A1(_u10_n20930 ), .A2(_u10_n20931 ), .ZN(adr1[24]));
NAND2_X1 _u10_U9589  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n20926 ) );
NAND2_X1 _u10_U9588  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n20927 ) );
NAND2_X1 _u10_U9587  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n20928 ) );
NAND2_X1 _u10_U9586  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n20929 ) );
NAND4_X1 _u10_U9585  ( .A1(_u10_n20926 ), .A2(_u10_n20927 ), .A3(_u10_n20928 ), .A4(_u10_n20929 ), .ZN(_u10_n20911 ) );
NAND2_X1 _u10_U9584  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n20922 ) );
NAND2_X1 _u10_U9583  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n20923 ) );
NAND2_X1 _u10_U9582  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n20924 ) );
NAND2_X1 _u10_U9581  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n20925 ) );
NAND4_X1 _u10_U9580  ( .A1(_u10_n20922 ), .A2(_u10_n20923 ), .A3(_u10_n20924 ), .A4(_u10_n20925 ), .ZN(_u10_n20912 ) );
NAND2_X1 _u10_U9579  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n20918 ) );
NAND2_X1 _u10_U9578  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n20919 ) );
NAND2_X1 _u10_U9577  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n20920 ) );
NAND2_X1 _u10_U9576  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n20921 ) );
NAND4_X1 _u10_U9575  ( .A1(_u10_n20918 ), .A2(_u10_n20919 ), .A3(_u10_n20920 ), .A4(_u10_n20921 ), .ZN(_u10_n20913 ) );
NAND2_X1 _u10_U9574  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n20915 ) );
NAND2_X1 _u10_U9573  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n20916 ) );
NAND2_X1 _u10_U9572  ( .A1(ch0_adr1[25]), .A2(_u10_n12003 ), .ZN(_u10_n20917 ) );
NAND3_X1 _u10_U9571  ( .A1(_u10_n20915 ), .A2(_u10_n20916 ), .A3(_u10_n20917 ), .ZN(_u10_n20914 ) );
NOR4_X1 _u10_U9570  ( .A1(_u10_n20911 ), .A2(_u10_n20912 ), .A3(_u10_n20913 ), .A4(_u10_n20914 ), .ZN(_u10_n20889 ) );
NAND2_X1 _u10_U9569  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20907 ) );
NAND2_X1 _u10_U9568  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20908 ) );
NAND2_X1 _u10_U9567  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20909 ) );
NAND2_X1 _u10_U9566  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20910 ) );
NAND4_X1 _u10_U9565  ( .A1(_u10_n20907 ), .A2(_u10_n20908 ), .A3(_u10_n20909 ), .A4(_u10_n20910 ), .ZN(_u10_n20891 ) );
NAND2_X1 _u10_U9564  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20903 ) );
NAND2_X1 _u10_U9563  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20904 ) );
NAND2_X1 _u10_U9562  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20905 ) );
NAND2_X1 _u10_U9561  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20906 ) );
NAND4_X1 _u10_U9560  ( .A1(_u10_n20903 ), .A2(_u10_n20904 ), .A3(_u10_n20905 ), .A4(_u10_n20906 ), .ZN(_u10_n20892 ) );
NAND2_X1 _u10_U9559  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20899 ) );
NAND2_X1 _u10_U9558  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20900 ) );
NAND2_X1 _u10_U9557  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20901 ) );
NAND2_X1 _u10_U9556  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20902 ) );
NAND4_X1 _u10_U9555  ( .A1(_u10_n20899 ), .A2(_u10_n20900 ), .A3(_u10_n20901 ), .A4(_u10_n20902 ), .ZN(_u10_n20893 ) );
NAND2_X1 _u10_U9554  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20895 ) );
NAND2_X1 _u10_U9553  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20896 ) );
NAND2_X1 _u10_U9552  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20897 ) );
NAND2_X1 _u10_U9551  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20898 ) );
NAND4_X1 _u10_U9550  ( .A1(_u10_n20895 ), .A2(_u10_n20896 ), .A3(_u10_n20897 ), .A4(_u10_n20898 ), .ZN(_u10_n20894 ) );
NOR4_X1 _u10_U9549  ( .A1(_u10_n20891 ), .A2(_u10_n20892 ), .A3(_u10_n20893 ), .A4(_u10_n20894 ), .ZN(_u10_n20890 ) );
NAND2_X1 _u10_U9548  ( .A1(_u10_n20889 ), .A2(_u10_n20890 ), .ZN(adr1[25]));
NAND2_X1 _u10_U9547  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n20885 ) );
NAND2_X1 _u10_U9546  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n20886 ) );
NAND2_X1 _u10_U9545  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n20887 ) );
NAND2_X1 _u10_U9544  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n20888 ) );
NAND4_X1 _u10_U9543  ( .A1(_u10_n20885 ), .A2(_u10_n20886 ), .A3(_u10_n20887 ), .A4(_u10_n20888 ), .ZN(_u10_n20870 ) );
NAND2_X1 _u10_U9542  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n20881 ) );
NAND2_X1 _u10_U9541  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n20882 ) );
NAND2_X1 _u10_U9540  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n20883 ) );
NAND2_X1 _u10_U9539  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n20884 ) );
NAND4_X1 _u10_U9538  ( .A1(_u10_n20881 ), .A2(_u10_n20882 ), .A3(_u10_n20883 ), .A4(_u10_n20884 ), .ZN(_u10_n20871 ) );
NAND2_X1 _u10_U9537  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n20877 ) );
NAND2_X1 _u10_U9536  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n20878 ) );
NAND2_X1 _u10_U9535  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n20879 ) );
NAND2_X1 _u10_U9534  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n20880 ) );
NAND4_X1 _u10_U9533  ( .A1(_u10_n20877 ), .A2(_u10_n20878 ), .A3(_u10_n20879 ), .A4(_u10_n20880 ), .ZN(_u10_n20872 ) );
NAND2_X1 _u10_U9532  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n20874 ) );
NAND2_X1 _u10_U9531  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n20875 ) );
NAND2_X1 _u10_U9530  ( .A1(ch0_adr1[26]), .A2(_u10_n12003 ), .ZN(_u10_n20876 ) );
NAND3_X1 _u10_U9529  ( .A1(_u10_n20874 ), .A2(_u10_n20875 ), .A3(_u10_n20876 ), .ZN(_u10_n20873 ) );
NOR4_X1 _u10_U9528  ( .A1(_u10_n20870 ), .A2(_u10_n20871 ), .A3(_u10_n20872 ), .A4(_u10_n20873 ), .ZN(_u10_n20848 ) );
NAND2_X1 _u10_U9527  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20866 ) );
NAND2_X1 _u10_U9526  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20867 ) );
NAND2_X1 _u10_U9525  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20868 ) );
NAND2_X1 _u10_U9524  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20869 ) );
NAND4_X1 _u10_U9523  ( .A1(_u10_n20866 ), .A2(_u10_n20867 ), .A3(_u10_n20868 ), .A4(_u10_n20869 ), .ZN(_u10_n20850 ) );
NAND2_X1 _u10_U9522  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20862 ) );
NAND2_X1 _u10_U9521  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20863 ) );
NAND2_X1 _u10_U9520  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20864 ) );
NAND2_X1 _u10_U9519  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20865 ) );
NAND4_X1 _u10_U9518  ( .A1(_u10_n20862 ), .A2(_u10_n20863 ), .A3(_u10_n20864 ), .A4(_u10_n20865 ), .ZN(_u10_n20851 ) );
NAND2_X1 _u10_U9517  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20858 ) );
NAND2_X1 _u10_U9516  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20859 ) );
NAND2_X1 _u10_U9515  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20860 ) );
NAND2_X1 _u10_U9514  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20861 ) );
NAND4_X1 _u10_U9513  ( .A1(_u10_n20858 ), .A2(_u10_n20859 ), .A3(_u10_n20860 ), .A4(_u10_n20861 ), .ZN(_u10_n20852 ) );
NAND2_X1 _u10_U9512  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20854 ) );
NAND2_X1 _u10_U9511  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20855 ) );
NAND2_X1 _u10_U9510  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20856 ) );
NAND2_X1 _u10_U9509  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20857 ) );
NAND4_X1 _u10_U9508  ( .A1(_u10_n20854 ), .A2(_u10_n20855 ), .A3(_u10_n20856 ), .A4(_u10_n20857 ), .ZN(_u10_n20853 ) );
NOR4_X1 _u10_U9507  ( .A1(_u10_n20850 ), .A2(_u10_n20851 ), .A3(_u10_n20852 ), .A4(_u10_n20853 ), .ZN(_u10_n20849 ) );
NAND2_X1 _u10_U9506  ( .A1(_u10_n20848 ), .A2(_u10_n20849 ), .ZN(adr1[26]));
NAND2_X1 _u10_U9505  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n20844 ) );
NAND2_X1 _u10_U9504  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n20845 ) );
NAND2_X1 _u10_U9503  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n20846 ) );
NAND2_X1 _u10_U9502  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n20847 ) );
NAND4_X1 _u10_U9501  ( .A1(_u10_n20844 ), .A2(_u10_n20845 ), .A3(_u10_n20846 ), .A4(_u10_n20847 ), .ZN(_u10_n20829 ) );
NAND2_X1 _u10_U9500  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n20840 ) );
NAND2_X1 _u10_U9499  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n20841 ) );
NAND2_X1 _u10_U9498  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n20842 ) );
NAND2_X1 _u10_U9497  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n20843 ) );
NAND4_X1 _u10_U9496  ( .A1(_u10_n20840 ), .A2(_u10_n20841 ), .A3(_u10_n20842 ), .A4(_u10_n20843 ), .ZN(_u10_n20830 ) );
NAND2_X1 _u10_U9495  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n20836 ) );
NAND2_X1 _u10_U9494  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n20837 ) );
NAND2_X1 _u10_U9493  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n20838 ) );
NAND2_X1 _u10_U9492  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n20839 ) );
NAND4_X1 _u10_U9491  ( .A1(_u10_n20836 ), .A2(_u10_n20837 ), .A3(_u10_n20838 ), .A4(_u10_n20839 ), .ZN(_u10_n20831 ) );
NAND2_X1 _u10_U9490  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n20833 ) );
NAND2_X1 _u10_U9489  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n20834 ) );
NAND2_X1 _u10_U9488  ( .A1(ch0_adr1[27]), .A2(_u10_n12003 ), .ZN(_u10_n20835 ) );
NAND3_X1 _u10_U9487  ( .A1(_u10_n20833 ), .A2(_u10_n20834 ), .A3(_u10_n20835 ), .ZN(_u10_n20832 ) );
NOR4_X1 _u10_U9486  ( .A1(_u10_n20829 ), .A2(_u10_n20830 ), .A3(_u10_n20831 ), .A4(_u10_n20832 ), .ZN(_u10_n20807 ) );
NAND2_X1 _u10_U9485  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20825 ) );
NAND2_X1 _u10_U9484  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20826 ) );
NAND2_X1 _u10_U9483  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20827 ) );
NAND2_X1 _u10_U9482  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20828 ) );
NAND4_X1 _u10_U9481  ( .A1(_u10_n20825 ), .A2(_u10_n20826 ), .A3(_u10_n20827 ), .A4(_u10_n20828 ), .ZN(_u10_n20809 ) );
NAND2_X1 _u10_U9480  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20821 ) );
NAND2_X1 _u10_U9479  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20822 ) );
NAND2_X1 _u10_U9478  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20823 ) );
NAND2_X1 _u10_U9477  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20824 ) );
NAND4_X1 _u10_U9476  ( .A1(_u10_n20821 ), .A2(_u10_n20822 ), .A3(_u10_n20823 ), .A4(_u10_n20824 ), .ZN(_u10_n20810 ) );
NAND2_X1 _u10_U9475  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20817 ) );
NAND2_X1 _u10_U9474  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20818 ) );
NAND2_X1 _u10_U9473  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20819 ) );
NAND2_X1 _u10_U9472  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20820 ) );
NAND4_X1 _u10_U9471  ( .A1(_u10_n20817 ), .A2(_u10_n20818 ), .A3(_u10_n20819 ), .A4(_u10_n20820 ), .ZN(_u10_n20811 ) );
NAND2_X1 _u10_U9470  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20813 ) );
NAND2_X1 _u10_U9469  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20814 ) );
NAND2_X1 _u10_U9468  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20815 ) );
NAND2_X1 _u10_U9467  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20816 ) );
NAND4_X1 _u10_U9466  ( .A1(_u10_n20813 ), .A2(_u10_n20814 ), .A3(_u10_n20815 ), .A4(_u10_n20816 ), .ZN(_u10_n20812 ) );
NOR4_X1 _u10_U9465  ( .A1(_u10_n20809 ), .A2(_u10_n20810 ), .A3(_u10_n20811 ), .A4(_u10_n20812 ), .ZN(_u10_n20808 ) );
NAND2_X1 _u10_U9464  ( .A1(_u10_n20807 ), .A2(_u10_n20808 ), .ZN(adr1[27]));
NAND2_X1 _u10_U9463  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n20803 ) );
NAND2_X1 _u10_U9462  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n20804 ) );
NAND2_X1 _u10_U9461  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n20805 ) );
NAND2_X1 _u10_U9460  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n20806 ) );
NAND4_X1 _u10_U9459  ( .A1(_u10_n20803 ), .A2(_u10_n20804 ), .A3(_u10_n20805 ), .A4(_u10_n20806 ), .ZN(_u10_n20788 ) );
NAND2_X1 _u10_U9458  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n20799 ) );
NAND2_X1 _u10_U9457  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n20800 ) );
NAND2_X1 _u10_U9456  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n20801 ) );
NAND2_X1 _u10_U9455  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n20802 ) );
NAND4_X1 _u10_U9454  ( .A1(_u10_n20799 ), .A2(_u10_n20800 ), .A3(_u10_n20801 ), .A4(_u10_n20802 ), .ZN(_u10_n20789 ) );
NAND2_X1 _u10_U9453  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n20795 ) );
NAND2_X1 _u10_U9452  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n20796 ) );
NAND2_X1 _u10_U9451  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n20797 ) );
NAND2_X1 _u10_U9450  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n20798 ) );
NAND4_X1 _u10_U9449  ( .A1(_u10_n20795 ), .A2(_u10_n20796 ), .A3(_u10_n20797 ), .A4(_u10_n20798 ), .ZN(_u10_n20790 ) );
NAND2_X1 _u10_U9448  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n20792 ) );
NAND2_X1 _u10_U9447  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n20793 ) );
NAND2_X1 _u10_U9446  ( .A1(ch0_adr1[28]), .A2(_u10_n12003 ), .ZN(_u10_n20794 ) );
NAND3_X1 _u10_U9445  ( .A1(_u10_n20792 ), .A2(_u10_n20793 ), .A3(_u10_n20794 ), .ZN(_u10_n20791 ) );
NOR4_X1 _u10_U9444  ( .A1(_u10_n20788 ), .A2(_u10_n20789 ), .A3(_u10_n20790 ), .A4(_u10_n20791 ), .ZN(_u10_n20766 ) );
NAND2_X1 _u10_U9443  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20784 ) );
NAND2_X1 _u10_U9442  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20785 ) );
NAND2_X1 _u10_U9441  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20786 ) );
NAND2_X1 _u10_U9440  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20787 ) );
NAND4_X1 _u10_U9439  ( .A1(_u10_n20784 ), .A2(_u10_n20785 ), .A3(_u10_n20786 ), .A4(_u10_n20787 ), .ZN(_u10_n20768 ) );
NAND2_X1 _u10_U9438  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20780 ) );
NAND2_X1 _u10_U9437  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20781 ) );
NAND2_X1 _u10_U9436  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20782 ) );
NAND2_X1 _u10_U9435  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20783 ) );
NAND4_X1 _u10_U9434  ( .A1(_u10_n20780 ), .A2(_u10_n20781 ), .A3(_u10_n20782 ), .A4(_u10_n20783 ), .ZN(_u10_n20769 ) );
NAND2_X1 _u10_U9433  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20776 ) );
NAND2_X1 _u10_U9432  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20777 ) );
NAND2_X1 _u10_U9431  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20778 ) );
NAND2_X1 _u10_U9430  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20779 ) );
NAND4_X1 _u10_U9429  ( .A1(_u10_n20776 ), .A2(_u10_n20777 ), .A3(_u10_n20778 ), .A4(_u10_n20779 ), .ZN(_u10_n20770 ) );
NAND2_X1 _u10_U9428  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20772 ) );
NAND2_X1 _u10_U9427  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20773 ) );
NAND2_X1 _u10_U9426  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20774 ) );
NAND2_X1 _u10_U9425  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20775 ) );
NAND4_X1 _u10_U9424  ( .A1(_u10_n20772 ), .A2(_u10_n20773 ), .A3(_u10_n20774 ), .A4(_u10_n20775 ), .ZN(_u10_n20771 ) );
NOR4_X1 _u10_U9423  ( .A1(_u10_n20768 ), .A2(_u10_n20769 ), .A3(_u10_n20770 ), .A4(_u10_n20771 ), .ZN(_u10_n20767 ) );
NAND2_X1 _u10_U9422  ( .A1(_u10_n20766 ), .A2(_u10_n20767 ), .ZN(adr1[28]));
NAND2_X1 _u10_U9421  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n20762 ) );
NAND2_X1 _u10_U9420  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n20763 ) );
NAND2_X1 _u10_U9419  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n20764 ) );
NAND2_X1 _u10_U9418  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n20765 ) );
NAND4_X1 _u10_U9417  ( .A1(_u10_n20762 ), .A2(_u10_n20763 ), .A3(_u10_n20764 ), .A4(_u10_n20765 ), .ZN(_u10_n20747 ) );
NAND2_X1 _u10_U9416  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n20758 ) );
NAND2_X1 _u10_U9415  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n20759 ) );
NAND2_X1 _u10_U9414  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n20760 ) );
NAND2_X1 _u10_U9413  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n20761 ) );
NAND4_X1 _u10_U9412  ( .A1(_u10_n20758 ), .A2(_u10_n20759 ), .A3(_u10_n20760 ), .A4(_u10_n20761 ), .ZN(_u10_n20748 ) );
NAND2_X1 _u10_U9411  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n20754 ) );
NAND2_X1 _u10_U9410  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n20755 ) );
NAND2_X1 _u10_U9409  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n20756 ) );
NAND2_X1 _u10_U9408  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n20757 ) );
NAND4_X1 _u10_U9407  ( .A1(_u10_n20754 ), .A2(_u10_n20755 ), .A3(_u10_n20756 ), .A4(_u10_n20757 ), .ZN(_u10_n20749 ) );
NAND2_X1 _u10_U9406  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n20751 ) );
NAND2_X1 _u10_U9405  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n20752 ) );
NAND2_X1 _u10_U9404  ( .A1(ch0_adr1[29]), .A2(_u10_n12003 ), .ZN(_u10_n20753 ) );
NAND3_X1 _u10_U9403  ( .A1(_u10_n20751 ), .A2(_u10_n20752 ), .A3(_u10_n20753 ), .ZN(_u10_n20750 ) );
NOR4_X1 _u10_U9402  ( .A1(_u10_n20747 ), .A2(_u10_n20748 ), .A3(_u10_n20749 ), .A4(_u10_n20750 ), .ZN(_u10_n20725 ) );
NAND2_X1 _u10_U9401  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20743 ) );
NAND2_X1 _u10_U9400  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20744 ) );
NAND2_X1 _u10_U9399  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20745 ) );
NAND2_X1 _u10_U9398  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20746 ) );
NAND4_X1 _u10_U9397  ( .A1(_u10_n20743 ), .A2(_u10_n20744 ), .A3(_u10_n20745 ), .A4(_u10_n20746 ), .ZN(_u10_n20727 ) );
NAND2_X1 _u10_U9396  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20739 ) );
NAND2_X1 _u10_U9395  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20740 ) );
NAND2_X1 _u10_U9394  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20741 ) );
NAND2_X1 _u10_U9393  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20742 ) );
NAND4_X1 _u10_U9392  ( .A1(_u10_n20739 ), .A2(_u10_n20740 ), .A3(_u10_n20741 ), .A4(_u10_n20742 ), .ZN(_u10_n20728 ) );
NAND2_X1 _u10_U9391  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20735 ) );
NAND2_X1 _u10_U9390  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20736 ) );
NAND2_X1 _u10_U9389  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20737 ) );
NAND2_X1 _u10_U9388  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20738 ) );
NAND4_X1 _u10_U9387  ( .A1(_u10_n20735 ), .A2(_u10_n20736 ), .A3(_u10_n20737 ), .A4(_u10_n20738 ), .ZN(_u10_n20729 ) );
NAND2_X1 _u10_U9386  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20731 ) );
NAND2_X1 _u10_U9385  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20732 ) );
NAND2_X1 _u10_U9384  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20733 ) );
NAND2_X1 _u10_U9383  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20734 ) );
NAND4_X1 _u10_U9382  ( .A1(_u10_n20731 ), .A2(_u10_n20732 ), .A3(_u10_n20733 ), .A4(_u10_n20734 ), .ZN(_u10_n20730 ) );
NOR4_X1 _u10_U9381  ( .A1(_u10_n20727 ), .A2(_u10_n20728 ), .A3(_u10_n20729 ), .A4(_u10_n20730 ), .ZN(_u10_n20726 ) );
NAND2_X1 _u10_U9380  ( .A1(_u10_n20725 ), .A2(_u10_n20726 ), .ZN(adr1[29]));
NAND2_X1 _u10_U9379  ( .A1(1'b0), .A2(_u10_n12334 ), .ZN(_u10_n20721 ) );
NAND2_X1 _u10_U9378  ( .A1(1'b0), .A2(_u10_n12310 ), .ZN(_u10_n20722 ) );
NAND2_X1 _u10_U9377  ( .A1(1'b0), .A2(_u10_n12286 ), .ZN(_u10_n20723 ) );
NAND2_X1 _u10_U9376  ( .A1(1'b0), .A2(_u10_n12262 ), .ZN(_u10_n20724 ) );
NAND4_X1 _u10_U9375  ( .A1(_u10_n20721 ), .A2(_u10_n20722 ), .A3(_u10_n20723 ), .A4(_u10_n20724 ), .ZN(_u10_n20706 ) );
NAND2_X1 _u10_U9374  ( .A1(1'b0), .A2(_u10_n12238 ), .ZN(_u10_n20717 ) );
NAND2_X1 _u10_U9373  ( .A1(1'b0), .A2(_u10_n12214 ), .ZN(_u10_n20718 ) );
NAND2_X1 _u10_U9372  ( .A1(1'b0), .A2(_u10_n12190 ), .ZN(_u10_n20719 ) );
NAND2_X1 _u10_U9371  ( .A1(1'b0), .A2(_u10_n12166 ), .ZN(_u10_n20720 ) );
NAND4_X1 _u10_U9370  ( .A1(_u10_n20717 ), .A2(_u10_n20718 ), .A3(_u10_n20719 ), .A4(_u10_n20720 ), .ZN(_u10_n20707 ) );
NAND2_X1 _u10_U9369  ( .A1(1'b0), .A2(_u10_n12142 ), .ZN(_u10_n20713 ) );
NAND2_X1 _u10_U9368  ( .A1(1'b0), .A2(_u10_n12118 ), .ZN(_u10_n20714 ) );
NAND2_X1 _u10_U9367  ( .A1(1'b0), .A2(_u10_n12094 ), .ZN(_u10_n20715 ) );
NAND2_X1 _u10_U9366  ( .A1(1'b0), .A2(_u10_n12070 ), .ZN(_u10_n20716 ) );
NAND4_X1 _u10_U9365  ( .A1(_u10_n20713 ), .A2(_u10_n20714 ), .A3(_u10_n20715 ), .A4(_u10_n20716 ), .ZN(_u10_n20708 ) );
NAND2_X1 _u10_U9364  ( .A1(1'b0), .A2(_u10_n12046 ), .ZN(_u10_n20710 ) );
NAND2_X1 _u10_U9363  ( .A1(1'b0), .A2(_u10_n12022 ), .ZN(_u10_n20711 ) );
NAND2_X1 _u10_U9362  ( .A1(ch0_adr1[2]), .A2(_u10_n12003 ), .ZN(_u10_n20712 ) );
NAND3_X1 _u10_U9361  ( .A1(_u10_n20710 ), .A2(_u10_n20711 ), .A3(_u10_n20712 ), .ZN(_u10_n20709 ) );
NOR4_X1 _u10_U9360  ( .A1(_u10_n20706 ), .A2(_u10_n20707 ), .A3(_u10_n20708 ), .A4(_u10_n20709 ), .ZN(_u10_n20684 ) );
NAND2_X1 _u10_U9359  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20702 ) );
NAND2_X1 _u10_U9358  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20703 ) );
NAND2_X1 _u10_U9357  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20704 ) );
NAND2_X1 _u10_U9356  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20705 ) );
NAND4_X1 _u10_U9355  ( .A1(_u10_n20702 ), .A2(_u10_n20703 ), .A3(_u10_n20704 ), .A4(_u10_n20705 ), .ZN(_u10_n20686 ) );
NAND2_X1 _u10_U9354  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20698 ) );
NAND2_X1 _u10_U9353  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20699 ) );
NAND2_X1 _u10_U9352  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20700 ) );
NAND2_X1 _u10_U9351  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20701 ) );
NAND4_X1 _u10_U9350  ( .A1(_u10_n20698 ), .A2(_u10_n20699 ), .A3(_u10_n20700 ), .A4(_u10_n20701 ), .ZN(_u10_n20687 ) );
NAND2_X1 _u10_U9349  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20694 ) );
NAND2_X1 _u10_U9348  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20695 ) );
NAND2_X1 _u10_U9347  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20696 ) );
NAND2_X1 _u10_U9346  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20697 ) );
NAND4_X1 _u10_U9345  ( .A1(_u10_n20694 ), .A2(_u10_n20695 ), .A3(_u10_n20696 ), .A4(_u10_n20697 ), .ZN(_u10_n20688 ) );
NAND2_X1 _u10_U9344  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20690 ) );
NAND2_X1 _u10_U9343  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20691 ) );
NAND2_X1 _u10_U9342  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20692 ) );
NAND2_X1 _u10_U9341  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20693 ) );
NAND4_X1 _u10_U9340  ( .A1(_u10_n20690 ), .A2(_u10_n20691 ), .A3(_u10_n20692 ), .A4(_u10_n20693 ), .ZN(_u10_n20689 ) );
NOR4_X1 _u10_U9339  ( .A1(_u10_n20686 ), .A2(_u10_n20687 ), .A3(_u10_n20688 ), .A4(_u10_n20689 ), .ZN(_u10_n20685 ) );
NAND2_X1 _u10_U9338  ( .A1(_u10_n20684 ), .A2(_u10_n20685 ), .ZN(adr1[2]) );
NAND2_X1 _u10_U9337  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20680 ) );
NAND2_X1 _u10_U9336  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20681 ) );
NAND2_X1 _u10_U9335  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20682 ) );
NAND2_X1 _u10_U9334  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20683 ) );
NAND4_X1 _u10_U9333  ( .A1(_u10_n20680 ), .A2(_u10_n20681 ), .A3(_u10_n20682 ), .A4(_u10_n20683 ), .ZN(_u10_n20665 ) );
NAND2_X1 _u10_U9332  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20676 ) );
NAND2_X1 _u10_U9331  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20677 ) );
NAND2_X1 _u10_U9330  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20678 ) );
NAND2_X1 _u10_U9329  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20679 ) );
NAND4_X1 _u10_U9328  ( .A1(_u10_n20676 ), .A2(_u10_n20677 ), .A3(_u10_n20678 ), .A4(_u10_n20679 ), .ZN(_u10_n20666 ) );
NAND2_X1 _u10_U9327  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20672 ) );
NAND2_X1 _u10_U9326  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20673 ) );
NAND2_X1 _u10_U9325  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20674 ) );
NAND2_X1 _u10_U9324  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20675 ) );
NAND4_X1 _u10_U9323  ( .A1(_u10_n20672 ), .A2(_u10_n20673 ), .A3(_u10_n20674 ), .A4(_u10_n20675 ), .ZN(_u10_n20667 ) );
NAND2_X1 _u10_U9322  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20669 ) );
NAND2_X1 _u10_U9321  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20670 ) );
NAND2_X1 _u10_U9320  ( .A1(ch0_adr1[30]), .A2(_u10_n12003 ), .ZN(_u10_n20671 ) );
NAND3_X1 _u10_U9319  ( .A1(_u10_n20669 ), .A2(_u10_n20670 ), .A3(_u10_n20671 ), .ZN(_u10_n20668 ) );
NOR4_X1 _u10_U9318  ( .A1(_u10_n20665 ), .A2(_u10_n20666 ), .A3(_u10_n20667 ), .A4(_u10_n20668 ), .ZN(_u10_n20643 ) );
NAND2_X1 _u10_U9317  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20661 ) );
NAND2_X1 _u10_U9316  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20662 ) );
NAND2_X1 _u10_U9315  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20663 ) );
NAND2_X1 _u10_U9314  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20664 ) );
NAND4_X1 _u10_U9313  ( .A1(_u10_n20661 ), .A2(_u10_n20662 ), .A3(_u10_n20663 ), .A4(_u10_n20664 ), .ZN(_u10_n20645 ) );
NAND2_X1 _u10_U9312  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20657 ) );
NAND2_X1 _u10_U9311  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20658 ) );
NAND2_X1 _u10_U9310  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20659 ) );
NAND2_X1 _u10_U9309  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20660 ) );
NAND4_X1 _u10_U9308  ( .A1(_u10_n20657 ), .A2(_u10_n20658 ), .A3(_u10_n20659 ), .A4(_u10_n20660 ), .ZN(_u10_n20646 ) );
NAND2_X1 _u10_U9307  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20653 ) );
NAND2_X1 _u10_U9306  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20654 ) );
NAND2_X1 _u10_U9305  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20655 ) );
NAND2_X1 _u10_U9304  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20656 ) );
NAND4_X1 _u10_U9303  ( .A1(_u10_n20653 ), .A2(_u10_n20654 ), .A3(_u10_n20655 ), .A4(_u10_n20656 ), .ZN(_u10_n20647 ) );
NAND2_X1 _u10_U9302  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20649 ) );
NAND2_X1 _u10_U9301  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20650 ) );
NAND2_X1 _u10_U9300  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20651 ) );
NAND2_X1 _u10_U9299  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20652 ) );
NAND4_X1 _u10_U9298  ( .A1(_u10_n20649 ), .A2(_u10_n20650 ), .A3(_u10_n20651 ), .A4(_u10_n20652 ), .ZN(_u10_n20648 ) );
NOR4_X1 _u10_U9297  ( .A1(_u10_n20645 ), .A2(_u10_n20646 ), .A3(_u10_n20647 ), .A4(_u10_n20648 ), .ZN(_u10_n20644 ) );
NAND2_X1 _u10_U9296  ( .A1(_u10_n20643 ), .A2(_u10_n20644 ), .ZN(adr1[30]));
NAND2_X1 _u10_U9295  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20639 ) );
NAND2_X1 _u10_U9294  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20640 ) );
NAND2_X1 _u10_U9293  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20641 ) );
NAND2_X1 _u10_U9292  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20642 ) );
NAND4_X1 _u10_U9291  ( .A1(_u10_n20639 ), .A2(_u10_n20640 ), .A3(_u10_n20641 ), .A4(_u10_n20642 ), .ZN(_u10_n20624 ) );
NAND2_X1 _u10_U9290  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20635 ) );
NAND2_X1 _u10_U9289  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20636 ) );
NAND2_X1 _u10_U9288  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20637 ) );
NAND2_X1 _u10_U9287  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20638 ) );
NAND4_X1 _u10_U9286  ( .A1(_u10_n20635 ), .A2(_u10_n20636 ), .A3(_u10_n20637 ), .A4(_u10_n20638 ), .ZN(_u10_n20625 ) );
NAND2_X1 _u10_U9285  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20631 ) );
NAND2_X1 _u10_U9284  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20632 ) );
NAND2_X1 _u10_U9283  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20633 ) );
NAND2_X1 _u10_U9282  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20634 ) );
NAND4_X1 _u10_U9281  ( .A1(_u10_n20631 ), .A2(_u10_n20632 ), .A3(_u10_n20633 ), .A4(_u10_n20634 ), .ZN(_u10_n20626 ) );
NAND2_X1 _u10_U9280  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20628 ) );
NAND2_X1 _u10_U9279  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20629 ) );
NAND2_X1 _u10_U9278  ( .A1(ch0_adr1[31]), .A2(_u10_n12003 ), .ZN(_u10_n20630 ) );
NAND3_X1 _u10_U9277  ( .A1(_u10_n20628 ), .A2(_u10_n20629 ), .A3(_u10_n20630 ), .ZN(_u10_n20627 ) );
NOR4_X1 _u10_U9276  ( .A1(_u10_n20624 ), .A2(_u10_n20625 ), .A3(_u10_n20626 ), .A4(_u10_n20627 ), .ZN(_u10_n20602 ) );
NAND2_X1 _u10_U9275  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20620 ) );
NAND2_X1 _u10_U9274  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20621 ) );
NAND2_X1 _u10_U9273  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20622 ) );
NAND2_X1 _u10_U9272  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20623 ) );
NAND4_X1 _u10_U9271  ( .A1(_u10_n20620 ), .A2(_u10_n20621 ), .A3(_u10_n20622 ), .A4(_u10_n20623 ), .ZN(_u10_n20604 ) );
NAND2_X1 _u10_U9270  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20616 ) );
NAND2_X1 _u10_U9269  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20617 ) );
NAND2_X1 _u10_U9268  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20618 ) );
NAND2_X1 _u10_U9267  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20619 ) );
NAND4_X1 _u10_U9266  ( .A1(_u10_n20616 ), .A2(_u10_n20617 ), .A3(_u10_n20618 ), .A4(_u10_n20619 ), .ZN(_u10_n20605 ) );
NAND2_X1 _u10_U9265  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20612 ) );
NAND2_X1 _u10_U9264  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20613 ) );
NAND2_X1 _u10_U9263  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20614 ) );
NAND2_X1 _u10_U9262  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20615 ) );
NAND4_X1 _u10_U9261  ( .A1(_u10_n20612 ), .A2(_u10_n20613 ), .A3(_u10_n20614 ), .A4(_u10_n20615 ), .ZN(_u10_n20606 ) );
NAND2_X1 _u10_U9260  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20608 ) );
NAND2_X1 _u10_U9259  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20609 ) );
NAND2_X1 _u10_U9258  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20610 ) );
NAND2_X1 _u10_U9257  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20611 ) );
NAND4_X1 _u10_U9256  ( .A1(_u10_n20608 ), .A2(_u10_n20609 ), .A3(_u10_n20610 ), .A4(_u10_n20611 ), .ZN(_u10_n20607 ) );
NOR4_X1 _u10_U9255  ( .A1(_u10_n20604 ), .A2(_u10_n20605 ), .A3(_u10_n20606 ), .A4(_u10_n20607 ), .ZN(_u10_n20603 ) );
NAND2_X1 _u10_U9254  ( .A1(_u10_n20602 ), .A2(_u10_n20603 ), .ZN(adr1[31]));
NAND2_X1 _u10_U9253  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20598 ) );
NAND2_X1 _u10_U9252  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20599 ) );
NAND2_X1 _u10_U9251  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20600 ) );
NAND2_X1 _u10_U9250  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20601 ) );
NAND4_X1 _u10_U9249  ( .A1(_u10_n20598 ), .A2(_u10_n20599 ), .A3(_u10_n20600 ), .A4(_u10_n20601 ), .ZN(_u10_n20583 ) );
NAND2_X1 _u10_U9248  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20594 ) );
NAND2_X1 _u10_U9247  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20595 ) );
NAND2_X1 _u10_U9246  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20596 ) );
NAND2_X1 _u10_U9245  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20597 ) );
NAND4_X1 _u10_U9244  ( .A1(_u10_n20594 ), .A2(_u10_n20595 ), .A3(_u10_n20596 ), .A4(_u10_n20597 ), .ZN(_u10_n20584 ) );
NAND2_X1 _u10_U9243  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20590 ) );
NAND2_X1 _u10_U9242  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20591 ) );
NAND2_X1 _u10_U9241  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20592 ) );
NAND2_X1 _u10_U9240  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20593 ) );
NAND4_X1 _u10_U9239  ( .A1(_u10_n20590 ), .A2(_u10_n20591 ), .A3(_u10_n20592 ), .A4(_u10_n20593 ), .ZN(_u10_n20585 ) );
NAND2_X1 _u10_U9238  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20587 ) );
NAND2_X1 _u10_U9237  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20588 ) );
NAND2_X1 _u10_U9236  ( .A1(ch0_adr1[3]), .A2(_u10_n12003 ), .ZN(_u10_n20589 ) );
NAND3_X1 _u10_U9235  ( .A1(_u10_n20587 ), .A2(_u10_n20588 ), .A3(_u10_n20589 ), .ZN(_u10_n20586 ) );
NOR4_X1 _u10_U9234  ( .A1(_u10_n20583 ), .A2(_u10_n20584 ), .A3(_u10_n20585 ), .A4(_u10_n20586 ), .ZN(_u10_n20561 ) );
NAND2_X1 _u10_U9233  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20579 ) );
NAND2_X1 _u10_U9232  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20580 ) );
NAND2_X1 _u10_U9231  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20581 ) );
NAND2_X1 _u10_U9230  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20582 ) );
NAND4_X1 _u10_U9229  ( .A1(_u10_n20579 ), .A2(_u10_n20580 ), .A3(_u10_n20581 ), .A4(_u10_n20582 ), .ZN(_u10_n20563 ) );
NAND2_X1 _u10_U9228  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20575 ) );
NAND2_X1 _u10_U9227  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20576 ) );
NAND2_X1 _u10_U9226  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20577 ) );
NAND2_X1 _u10_U9225  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20578 ) );
NAND4_X1 _u10_U9224  ( .A1(_u10_n20575 ), .A2(_u10_n20576 ), .A3(_u10_n20577 ), .A4(_u10_n20578 ), .ZN(_u10_n20564 ) );
NAND2_X1 _u10_U9223  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20571 ) );
NAND2_X1 _u10_U9222  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20572 ) );
NAND2_X1 _u10_U9221  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20573 ) );
NAND2_X1 _u10_U9220  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20574 ) );
NAND4_X1 _u10_U9219  ( .A1(_u10_n20571 ), .A2(_u10_n20572 ), .A3(_u10_n20573 ), .A4(_u10_n20574 ), .ZN(_u10_n20565 ) );
NAND2_X1 _u10_U9218  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20567 ) );
NAND2_X1 _u10_U9217  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20568 ) );
NAND2_X1 _u10_U9216  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20569 ) );
NAND2_X1 _u10_U9215  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20570 ) );
NAND4_X1 _u10_U9214  ( .A1(_u10_n20567 ), .A2(_u10_n20568 ), .A3(_u10_n20569 ), .A4(_u10_n20570 ), .ZN(_u10_n20566 ) );
NOR4_X1 _u10_U9213  ( .A1(_u10_n20563 ), .A2(_u10_n20564 ), .A3(_u10_n20565 ), .A4(_u10_n20566 ), .ZN(_u10_n20562 ) );
NAND2_X1 _u10_U9212  ( .A1(_u10_n20561 ), .A2(_u10_n20562 ), .ZN(adr1[3]) );
NAND2_X1 _u10_U9211  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20557 ) );
NAND2_X1 _u10_U9210  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20558 ) );
NAND2_X1 _u10_U9209  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20559 ) );
NAND2_X1 _u10_U9208  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20560 ) );
NAND4_X1 _u10_U9207  ( .A1(_u10_n20557 ), .A2(_u10_n20558 ), .A3(_u10_n20559 ), .A4(_u10_n20560 ), .ZN(_u10_n20542 ) );
NAND2_X1 _u10_U9206  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20553 ) );
NAND2_X1 _u10_U9205  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20554 ) );
NAND2_X1 _u10_U9204  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20555 ) );
NAND2_X1 _u10_U9203  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20556 ) );
NAND4_X1 _u10_U9202  ( .A1(_u10_n20553 ), .A2(_u10_n20554 ), .A3(_u10_n20555 ), .A4(_u10_n20556 ), .ZN(_u10_n20543 ) );
NAND2_X1 _u10_U9201  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20549 ) );
NAND2_X1 _u10_U9200  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20550 ) );
NAND2_X1 _u10_U9199  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20551 ) );
NAND2_X1 _u10_U9198  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20552 ) );
NAND4_X1 _u10_U9197  ( .A1(_u10_n20549 ), .A2(_u10_n20550 ), .A3(_u10_n20551 ), .A4(_u10_n20552 ), .ZN(_u10_n20544 ) );
NAND2_X1 _u10_U9196  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20546 ) );
NAND2_X1 _u10_U9195  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20547 ) );
NAND2_X1 _u10_U9194  ( .A1(ch0_adr1[4]), .A2(_u10_n12003 ), .ZN(_u10_n20548 ) );
NAND3_X1 _u10_U9193  ( .A1(_u10_n20546 ), .A2(_u10_n20547 ), .A3(_u10_n20548 ), .ZN(_u10_n20545 ) );
NOR4_X1 _u10_U9192  ( .A1(_u10_n20542 ), .A2(_u10_n20543 ), .A3(_u10_n20544 ), .A4(_u10_n20545 ), .ZN(_u10_n20520 ) );
NAND2_X1 _u10_U9191  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20538 ) );
NAND2_X1 _u10_U9190  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20539 ) );
NAND2_X1 _u10_U9189  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20540 ) );
NAND2_X1 _u10_U9188  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20541 ) );
NAND4_X1 _u10_U9187  ( .A1(_u10_n20538 ), .A2(_u10_n20539 ), .A3(_u10_n20540 ), .A4(_u10_n20541 ), .ZN(_u10_n20522 ) );
NAND2_X1 _u10_U9186  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20534 ) );
NAND2_X1 _u10_U9185  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20535 ) );
NAND2_X1 _u10_U9184  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20536 ) );
NAND2_X1 _u10_U9183  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20537 ) );
NAND4_X1 _u10_U9182  ( .A1(_u10_n20534 ), .A2(_u10_n20535 ), .A3(_u10_n20536 ), .A4(_u10_n20537 ), .ZN(_u10_n20523 ) );
NAND2_X1 _u10_U9181  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20530 ) );
NAND2_X1 _u10_U9180  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20531 ) );
NAND2_X1 _u10_U9179  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20532 ) );
NAND2_X1 _u10_U9178  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20533 ) );
NAND4_X1 _u10_U9177  ( .A1(_u10_n20530 ), .A2(_u10_n20531 ), .A3(_u10_n20532 ), .A4(_u10_n20533 ), .ZN(_u10_n20524 ) );
NAND2_X1 _u10_U9176  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20526 ) );
NAND2_X1 _u10_U9175  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20527 ) );
NAND2_X1 _u10_U9174  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20528 ) );
NAND2_X1 _u10_U9173  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20529 ) );
NAND4_X1 _u10_U9172  ( .A1(_u10_n20526 ), .A2(_u10_n20527 ), .A3(_u10_n20528 ), .A4(_u10_n20529 ), .ZN(_u10_n20525 ) );
NOR4_X1 _u10_U9171  ( .A1(_u10_n20522 ), .A2(_u10_n20523 ), .A3(_u10_n20524 ), .A4(_u10_n20525 ), .ZN(_u10_n20521 ) );
NAND2_X1 _u10_U9170  ( .A1(_u10_n20520 ), .A2(_u10_n20521 ), .ZN(adr1[4]) );
NAND2_X1 _u10_U9169  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20516 ) );
NAND2_X1 _u10_U9168  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20517 ) );
NAND2_X1 _u10_U9167  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20518 ) );
NAND2_X1 _u10_U9166  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20519 ) );
NAND4_X1 _u10_U9165  ( .A1(_u10_n20516 ), .A2(_u10_n20517 ), .A3(_u10_n20518 ), .A4(_u10_n20519 ), .ZN(_u10_n20501 ) );
NAND2_X1 _u10_U9164  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20512 ) );
NAND2_X1 _u10_U9163  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20513 ) );
NAND2_X1 _u10_U9162  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20514 ) );
NAND2_X1 _u10_U9161  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20515 ) );
NAND4_X1 _u10_U9160  ( .A1(_u10_n20512 ), .A2(_u10_n20513 ), .A3(_u10_n20514 ), .A4(_u10_n20515 ), .ZN(_u10_n20502 ) );
NAND2_X1 _u10_U9159  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20508 ) );
NAND2_X1 _u10_U9158  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20509 ) );
NAND2_X1 _u10_U9157  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20510 ) );
NAND2_X1 _u10_U9156  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20511 ) );
NAND4_X1 _u10_U9155  ( .A1(_u10_n20508 ), .A2(_u10_n20509 ), .A3(_u10_n20510 ), .A4(_u10_n20511 ), .ZN(_u10_n20503 ) );
NAND2_X1 _u10_U9154  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20505 ) );
NAND2_X1 _u10_U9153  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20506 ) );
NAND2_X1 _u10_U9152  ( .A1(ch0_adr1[5]), .A2(_u10_n12004 ), .ZN(_u10_n20507 ) );
NAND3_X1 _u10_U9151  ( .A1(_u10_n20505 ), .A2(_u10_n20506 ), .A3(_u10_n20507 ), .ZN(_u10_n20504 ) );
NOR4_X1 _u10_U9150  ( .A1(_u10_n20501 ), .A2(_u10_n20502 ), .A3(_u10_n20503 ), .A4(_u10_n20504 ), .ZN(_u10_n20479 ) );
NAND2_X1 _u10_U9149  ( .A1(1'b0), .A2(_u10_n11987 ), .ZN(_u10_n20497 ) );
NAND2_X1 _u10_U9148  ( .A1(1'b0), .A2(_u10_n11963 ), .ZN(_u10_n20498 ) );
NAND2_X1 _u10_U9147  ( .A1(1'b0), .A2(_u10_n11939 ), .ZN(_u10_n20499 ) );
NAND2_X1 _u10_U9146  ( .A1(1'b0), .A2(_u10_n11915 ), .ZN(_u10_n20500 ) );
NAND4_X1 _u10_U9145  ( .A1(_u10_n20497 ), .A2(_u10_n20498 ), .A3(_u10_n20499 ), .A4(_u10_n20500 ), .ZN(_u10_n20481 ) );
NAND2_X1 _u10_U9144  ( .A1(1'b0), .A2(_u10_n11891 ), .ZN(_u10_n20493 ) );
NAND2_X1 _u10_U9143  ( .A1(1'b0), .A2(_u10_n11867 ), .ZN(_u10_n20494 ) );
NAND2_X1 _u10_U9142  ( .A1(1'b0), .A2(_u10_n11843 ), .ZN(_u10_n20495 ) );
NAND2_X1 _u10_U9141  ( .A1(1'b0), .A2(_u10_n11819 ), .ZN(_u10_n20496 ) );
NAND4_X1 _u10_U9140  ( .A1(_u10_n20493 ), .A2(_u10_n20494 ), .A3(_u10_n20495 ), .A4(_u10_n20496 ), .ZN(_u10_n20482 ) );
NAND2_X1 _u10_U9139  ( .A1(1'b0), .A2(_u10_n11795 ), .ZN(_u10_n20489 ) );
NAND2_X1 _u10_U9138  ( .A1(1'b0), .A2(_u10_n11771 ), .ZN(_u10_n20490 ) );
NAND2_X1 _u10_U9137  ( .A1(1'b0), .A2(_u10_n11747 ), .ZN(_u10_n20491 ) );
NAND2_X1 _u10_U9136  ( .A1(1'b0), .A2(_u10_n11723 ), .ZN(_u10_n20492 ) );
NAND4_X1 _u10_U9135  ( .A1(_u10_n20489 ), .A2(_u10_n20490 ), .A3(_u10_n20491 ), .A4(_u10_n20492 ), .ZN(_u10_n20483 ) );
NAND2_X1 _u10_U9134  ( .A1(1'b0), .A2(_u10_n11699 ), .ZN(_u10_n20485 ) );
NAND2_X1 _u10_U9133  ( .A1(1'b0), .A2(_u10_n11675 ), .ZN(_u10_n20486 ) );
NAND2_X1 _u10_U9132  ( .A1(1'b0), .A2(_u10_n11651 ), .ZN(_u10_n20487 ) );
NAND2_X1 _u10_U9131  ( .A1(1'b0), .A2(_u10_n11627 ), .ZN(_u10_n20488 ) );
NAND4_X1 _u10_U9130  ( .A1(_u10_n20485 ), .A2(_u10_n20486 ), .A3(_u10_n20487 ), .A4(_u10_n20488 ), .ZN(_u10_n20484 ) );
NOR4_X1 _u10_U9129  ( .A1(_u10_n20481 ), .A2(_u10_n20482 ), .A3(_u10_n20483 ), .A4(_u10_n20484 ), .ZN(_u10_n20480 ) );
NAND2_X1 _u10_U9128  ( .A1(_u10_n20479 ), .A2(_u10_n20480 ), .ZN(adr1[5]) );
NAND2_X1 _u10_U9127  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20475 ) );
NAND2_X1 _u10_U9126  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20476 ) );
NAND2_X1 _u10_U9125  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20477 ) );
NAND2_X1 _u10_U9124  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20478 ) );
NAND4_X1 _u10_U9123  ( .A1(_u10_n20475 ), .A2(_u10_n20476 ), .A3(_u10_n20477 ), .A4(_u10_n20478 ), .ZN(_u10_n20460 ) );
NAND2_X1 _u10_U9122  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20471 ) );
NAND2_X1 _u10_U9121  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20472 ) );
NAND2_X1 _u10_U9120  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20473 ) );
NAND2_X1 _u10_U9119  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20474 ) );
NAND4_X1 _u10_U9118  ( .A1(_u10_n20471 ), .A2(_u10_n20472 ), .A3(_u10_n20473 ), .A4(_u10_n20474 ), .ZN(_u10_n20461 ) );
NAND2_X1 _u10_U9117  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20467 ) );
NAND2_X1 _u10_U9116  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20468 ) );
NAND2_X1 _u10_U9115  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20469 ) );
NAND2_X1 _u10_U9114  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20470 ) );
NAND4_X1 _u10_U9113  ( .A1(_u10_n20467 ), .A2(_u10_n20468 ), .A3(_u10_n20469 ), .A4(_u10_n20470 ), .ZN(_u10_n20462 ) );
NAND2_X1 _u10_U9112  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20464 ) );
NAND2_X1 _u10_U9111  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20465 ) );
NAND2_X1 _u10_U9110  ( .A1(ch0_adr1[6]), .A2(_u10_n12004 ), .ZN(_u10_n20466 ) );
NAND3_X1 _u10_U9109  ( .A1(_u10_n20464 ), .A2(_u10_n20465 ), .A3(_u10_n20466 ), .ZN(_u10_n20463 ) );
NOR4_X1 _u10_U9108  ( .A1(_u10_n20460 ), .A2(_u10_n20461 ), .A3(_u10_n20462 ), .A4(_u10_n20463 ), .ZN(_u10_n20438 ) );
NAND2_X1 _u10_U9107  ( .A1(1'b0), .A2(_u10_n11999 ), .ZN(_u10_n20456 ) );
NAND2_X1 _u10_U9106  ( .A1(1'b0), .A2(_u10_n11974 ), .ZN(_u10_n20457 ) );
NAND2_X1 _u10_U9105  ( .A1(1'b0), .A2(_u10_n11949 ), .ZN(_u10_n20458 ) );
NAND2_X1 _u10_U9104  ( .A1(1'b0), .A2(_u10_n11925 ), .ZN(_u10_n20459 ) );
NAND4_X1 _u10_U9103  ( .A1(_u10_n20456 ), .A2(_u10_n20457 ), .A3(_u10_n20458 ), .A4(_u10_n20459 ), .ZN(_u10_n20440 ) );
NAND2_X1 _u10_U9102  ( .A1(1'b0), .A2(_u10_n11903 ), .ZN(_u10_n20452 ) );
NAND2_X1 _u10_U9101  ( .A1(1'b0), .A2(_u10_n11879 ), .ZN(_u10_n20453 ) );
NAND2_X1 _u10_U9100  ( .A1(1'b0), .A2(_u10_n11849 ), .ZN(_u10_n20454 ) );
NAND2_X1 _u10_U9099  ( .A1(1'b0), .A2(_u10_n11831 ), .ZN(_u10_n20455 ) );
NAND4_X1 _u10_U9098  ( .A1(_u10_n20452 ), .A2(_u10_n20453 ), .A3(_u10_n20454 ), .A4(_u10_n20455 ), .ZN(_u10_n20441 ) );
NAND2_X1 _u10_U9097  ( .A1(1'b0), .A2(_u10_n11807 ), .ZN(_u10_n20448 ) );
NAND2_X1 _u10_U9096  ( .A1(1'b0), .A2(_u10_n11783 ), .ZN(_u10_n20449 ) );
NAND2_X1 _u10_U9095  ( .A1(1'b0), .A2(_u10_n11756 ), .ZN(_u10_n20450 ) );
NAND2_X1 _u10_U9094  ( .A1(1'b0), .A2(_u10_n11732 ), .ZN(_u10_n20451 ) );
NAND4_X1 _u10_U9093  ( .A1(_u10_n20448 ), .A2(_u10_n20449 ), .A3(_u10_n20450 ), .A4(_u10_n20451 ), .ZN(_u10_n20442 ) );
NAND2_X1 _u10_U9092  ( .A1(1'b0), .A2(_u10_n11708 ), .ZN(_u10_n20444 ) );
NAND2_X1 _u10_U9091  ( .A1(1'b0), .A2(_u10_n11684 ), .ZN(_u10_n20445 ) );
NAND2_X1 _u10_U9090  ( .A1(1'b0), .A2(_u10_n11657 ), .ZN(_u10_n20446 ) );
NAND2_X1 _u10_U9089  ( .A1(1'b0), .A2(_u10_n11633 ), .ZN(_u10_n20447 ) );
NAND4_X1 _u10_U9088  ( .A1(_u10_n20444 ), .A2(_u10_n20445 ), .A3(_u10_n20446 ), .A4(_u10_n20447 ), .ZN(_u10_n20443 ) );
NOR4_X1 _u10_U9087  ( .A1(_u10_n20440 ), .A2(_u10_n20441 ), .A3(_u10_n20442 ), .A4(_u10_n20443 ), .ZN(_u10_n20439 ) );
NAND2_X1 _u10_U9086  ( .A1(_u10_n20438 ), .A2(_u10_n20439 ), .ZN(adr1[6]) );
NAND2_X1 _u10_U9085  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20434 ) );
NAND2_X1 _u10_U9084  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20435 ) );
NAND2_X1 _u10_U9083  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20436 ) );
NAND2_X1 _u10_U9082  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20437 ) );
NAND4_X1 _u10_U9081  ( .A1(_u10_n20434 ), .A2(_u10_n20435 ), .A3(_u10_n20436 ), .A4(_u10_n20437 ), .ZN(_u10_n20419 ) );
NAND2_X1 _u10_U9080  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20430 ) );
NAND2_X1 _u10_U9079  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20431 ) );
NAND2_X1 _u10_U9078  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20432 ) );
NAND2_X1 _u10_U9077  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20433 ) );
NAND4_X1 _u10_U9076  ( .A1(_u10_n20430 ), .A2(_u10_n20431 ), .A3(_u10_n20432 ), .A4(_u10_n20433 ), .ZN(_u10_n20420 ) );
NAND2_X1 _u10_U9075  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20426 ) );
NAND2_X1 _u10_U9074  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20427 ) );
NAND2_X1 _u10_U9073  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20428 ) );
NAND2_X1 _u10_U9072  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20429 ) );
NAND4_X1 _u10_U9071  ( .A1(_u10_n20426 ), .A2(_u10_n20427 ), .A3(_u10_n20428 ), .A4(_u10_n20429 ), .ZN(_u10_n20421 ) );
NAND2_X1 _u10_U9070  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20423 ) );
NAND2_X1 _u10_U9069  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20424 ) );
NAND2_X1 _u10_U9068  ( .A1(ch0_adr1[7]), .A2(_u10_n12004 ), .ZN(_u10_n20425 ) );
NAND3_X1 _u10_U9067  ( .A1(_u10_n20423 ), .A2(_u10_n20424 ), .A3(_u10_n20425 ), .ZN(_u10_n20422 ) );
NOR4_X1 _u10_U9066  ( .A1(_u10_n20419 ), .A2(_u10_n20420 ), .A3(_u10_n20421 ), .A4(_u10_n20422 ), .ZN(_u10_n20397 ) );
NAND2_X1 _u10_U9065  ( .A1(1'b0), .A2(_u10_n11996 ), .ZN(_u10_n20415 ) );
NAND2_X1 _u10_U9064  ( .A1(1'b0), .A2(_u10_n11973 ), .ZN(_u10_n20416 ) );
NAND2_X1 _u10_U9063  ( .A1(1'b0), .A2(_u10_n11950 ), .ZN(_u10_n20417 ) );
NAND2_X1 _u10_U9062  ( .A1(1'b0), .A2(_u10_n11926 ), .ZN(_u10_n20418 ) );
NAND4_X1 _u10_U9061  ( .A1(_u10_n20415 ), .A2(_u10_n20416 ), .A3(_u10_n20417 ), .A4(_u10_n20418 ), .ZN(_u10_n20399 ) );
NAND2_X1 _u10_U9060  ( .A1(1'b0), .A2(_u10_n11900 ), .ZN(_u10_n20411 ) );
NAND2_X1 _u10_U9059  ( .A1(1'b0), .A2(_u10_n11876 ), .ZN(_u10_n20412 ) );
NAND2_X1 _u10_U9058  ( .A1(1'b0), .A2(_u10_n11855 ), .ZN(_u10_n20413 ) );
NAND2_X1 _u10_U9057  ( .A1(1'b0), .A2(_u10_n11828 ), .ZN(_u10_n20414 ) );
NAND4_X1 _u10_U9056  ( .A1(_u10_n20411 ), .A2(_u10_n20412 ), .A3(_u10_n20413 ), .A4(_u10_n20414 ), .ZN(_u10_n20400 ) );
NAND2_X1 _u10_U9055  ( .A1(1'b0), .A2(_u10_n11804 ), .ZN(_u10_n20407 ) );
NAND2_X1 _u10_U9054  ( .A1(1'b0), .A2(_u10_n11780 ), .ZN(_u10_n20408 ) );
NAND2_X1 _u10_U9053  ( .A1(1'b0), .A2(_u10_n11759 ), .ZN(_u10_n20409 ) );
NAND2_X1 _u10_U9052  ( .A1(1'b0), .A2(_u10_n11735 ), .ZN(_u10_n20410 ) );
NAND4_X1 _u10_U9051  ( .A1(_u10_n20407 ), .A2(_u10_n20408 ), .A3(_u10_n20409 ), .A4(_u10_n20410 ), .ZN(_u10_n20401 ) );
NAND2_X1 _u10_U9050  ( .A1(1'b0), .A2(_u10_n11711 ), .ZN(_u10_n20403 ) );
NAND2_X1 _u10_U9049  ( .A1(1'b0), .A2(_u10_n11687 ), .ZN(_u10_n20404 ) );
NAND2_X1 _u10_U9048  ( .A1(1'b0), .A2(_u10_n11663 ), .ZN(_u10_n20405 ) );
NAND2_X1 _u10_U9047  ( .A1(1'b0), .A2(_u10_n11639 ), .ZN(_u10_n20406 ) );
NAND4_X1 _u10_U9046  ( .A1(_u10_n20403 ), .A2(_u10_n20404 ), .A3(_u10_n20405 ), .A4(_u10_n20406 ), .ZN(_u10_n20402 ) );
NOR4_X1 _u10_U9045  ( .A1(_u10_n20399 ), .A2(_u10_n20400 ), .A3(_u10_n20401 ), .A4(_u10_n20402 ), .ZN(_u10_n20398 ) );
NAND2_X1 _u10_U9044  ( .A1(_u10_n20397 ), .A2(_u10_n20398 ), .ZN(adr1[7]) );
NAND2_X1 _u10_U9043  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20393 ) );
NAND2_X1 _u10_U9042  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20394 ) );
NAND2_X1 _u10_U9041  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20395 ) );
NAND2_X1 _u10_U9040  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20396 ) );
NAND4_X1 _u10_U9039  ( .A1(_u10_n20393 ), .A2(_u10_n20394 ), .A3(_u10_n20395 ), .A4(_u10_n20396 ), .ZN(_u10_n20378 ) );
NAND2_X1 _u10_U9038  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20389 ) );
NAND2_X1 _u10_U9037  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20390 ) );
NAND2_X1 _u10_U9036  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20391 ) );
NAND2_X1 _u10_U9035  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20392 ) );
NAND4_X1 _u10_U9034  ( .A1(_u10_n20389 ), .A2(_u10_n20390 ), .A3(_u10_n20391 ), .A4(_u10_n20392 ), .ZN(_u10_n20379 ) );
NAND2_X1 _u10_U9033  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20385 ) );
NAND2_X1 _u10_U9032  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20386 ) );
NAND2_X1 _u10_U9031  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20387 ) );
NAND2_X1 _u10_U9030  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20388 ) );
NAND4_X1 _u10_U9029  ( .A1(_u10_n20385 ), .A2(_u10_n20386 ), .A3(_u10_n20387 ), .A4(_u10_n20388 ), .ZN(_u10_n20380 ) );
NAND2_X1 _u10_U9028  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20382 ) );
NAND2_X1 _u10_U9027  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20383 ) );
NAND2_X1 _u10_U9026  ( .A1(ch0_adr1[8]), .A2(_u10_n12004 ), .ZN(_u10_n20384 ) );
NAND3_X1 _u10_U9025  ( .A1(_u10_n20382 ), .A2(_u10_n20383 ), .A3(_u10_n20384 ), .ZN(_u10_n20381 ) );
NOR4_X1 _u10_U9024  ( .A1(_u10_n20378 ), .A2(_u10_n20379 ), .A3(_u10_n20380 ), .A4(_u10_n20381 ), .ZN(_u10_n20356 ) );
NAND2_X1 _u10_U9023  ( .A1(1'b0), .A2(_u10_n11996 ), .ZN(_u10_n20374 ) );
NAND2_X1 _u10_U9022  ( .A1(1'b0), .A2(_u10_n11972 ), .ZN(_u10_n20375 ) );
NAND2_X1 _u10_U9021  ( .A1(1'b0), .A2(_u10_n11948 ), .ZN(_u10_n20376 ) );
NAND2_X1 _u10_U9020  ( .A1(1'b0), .A2(_u10_n11924 ), .ZN(_u10_n20377 ) );
NAND4_X1 _u10_U9019  ( .A1(_u10_n20374 ), .A2(_u10_n20375 ), .A3(_u10_n20376 ), .A4(_u10_n20377 ), .ZN(_u10_n20358 ) );
NAND2_X1 _u10_U9018  ( .A1(1'b0), .A2(_u10_n11900 ), .ZN(_u10_n20370 ) );
NAND2_X1 _u10_U9017  ( .A1(1'b0), .A2(_u10_n11876 ), .ZN(_u10_n20371 ) );
NAND2_X1 _u10_U9016  ( .A1(1'b0), .A2(_u10_n11852 ), .ZN(_u10_n20372 ) );
NAND2_X1 _u10_U9015  ( .A1(1'b0), .A2(_u10_n11828 ), .ZN(_u10_n20373 ) );
NAND4_X1 _u10_U9014  ( .A1(_u10_n20370 ), .A2(_u10_n20371 ), .A3(_u10_n20372 ), .A4(_u10_n20373 ), .ZN(_u10_n20359 ) );
NAND2_X1 _u10_U9013  ( .A1(1'b0), .A2(_u10_n11804 ), .ZN(_u10_n20366 ) );
NAND2_X1 _u10_U9012  ( .A1(1'b0), .A2(_u10_n11780 ), .ZN(_u10_n20367 ) );
NAND2_X1 _u10_U9011  ( .A1(1'b0), .A2(_u10_n11756 ), .ZN(_u10_n20368 ) );
NAND2_X1 _u10_U9010  ( .A1(1'b0), .A2(_u10_n11732 ), .ZN(_u10_n20369 ) );
NAND4_X1 _u10_U9009  ( .A1(_u10_n20366 ), .A2(_u10_n20367 ), .A3(_u10_n20368 ), .A4(_u10_n20369 ), .ZN(_u10_n20360 ) );
NAND2_X1 _u10_U9008  ( .A1(1'b0), .A2(_u10_n11708 ), .ZN(_u10_n20362 ) );
NAND2_X1 _u10_U9007  ( .A1(1'b0), .A2(_u10_n11684 ), .ZN(_u10_n20363 ) );
NAND2_X1 _u10_U9006  ( .A1(1'b0), .A2(_u10_n11660 ), .ZN(_u10_n20364 ) );
NAND2_X1 _u10_U9005  ( .A1(1'b0), .A2(_u10_n11636 ), .ZN(_u10_n20365 ) );
NAND4_X1 _u10_U9004  ( .A1(_u10_n20362 ), .A2(_u10_n20363 ), .A3(_u10_n20364 ), .A4(_u10_n20365 ), .ZN(_u10_n20361 ) );
NOR4_X1 _u10_U9003  ( .A1(_u10_n20358 ), .A2(_u10_n20359 ), .A3(_u10_n20360 ), .A4(_u10_n20361 ), .ZN(_u10_n20357 ) );
NAND2_X1 _u10_U9002  ( .A1(_u10_n20356 ), .A2(_u10_n20357 ), .ZN(adr1[8]) );
NAND2_X1 _u10_U9001  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20352 ) );
NAND2_X1 _u10_U9000  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20353 ) );
NAND2_X1 _u10_U8999  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20354 ) );
NAND2_X1 _u10_U8998  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20355 ) );
NAND4_X1 _u10_U8997  ( .A1(_u10_n20352 ), .A2(_u10_n20353 ), .A3(_u10_n20354 ), .A4(_u10_n20355 ), .ZN(_u10_n20337 ) );
NAND2_X1 _u10_U8996  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20348 ) );
NAND2_X1 _u10_U8995  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20349 ) );
NAND2_X1 _u10_U8994  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20350 ) );
NAND2_X1 _u10_U8993  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20351 ) );
NAND4_X1 _u10_U8992  ( .A1(_u10_n20348 ), .A2(_u10_n20349 ), .A3(_u10_n20350 ), .A4(_u10_n20351 ), .ZN(_u10_n20338 ) );
NAND2_X1 _u10_U8991  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20344 ) );
NAND2_X1 _u10_U8990  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20345 ) );
NAND2_X1 _u10_U8989  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20346 ) );
NAND2_X1 _u10_U8988  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20347 ) );
NAND4_X1 _u10_U8987  ( .A1(_u10_n20344 ), .A2(_u10_n20345 ), .A3(_u10_n20346 ), .A4(_u10_n20347 ), .ZN(_u10_n20339 ) );
NAND2_X1 _u10_U8986  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20341 ) );
NAND2_X1 _u10_U8985  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20342 ) );
NAND2_X1 _u10_U8984  ( .A1(ch0_adr1[9]), .A2(_u10_n12004 ), .ZN(_u10_n20343 ) );
NAND3_X1 _u10_U8983  ( .A1(_u10_n20341 ), .A2(_u10_n20342 ), .A3(_u10_n20343 ), .ZN(_u10_n20340 ) );
NOR4_X1 _u10_U8982  ( .A1(_u10_n20337 ), .A2(_u10_n20338 ), .A3(_u10_n20339 ), .A4(_u10_n20340 ), .ZN(_u10_n20315 ) );
NAND2_X1 _u10_U8981  ( .A1(1'b0), .A2(_u10_n11994 ), .ZN(_u10_n20333 ) );
NAND2_X1 _u10_U8980  ( .A1(1'b0), .A2(_u10_n11975 ), .ZN(_u10_n20334 ) );
NAND2_X1 _u10_U8979  ( .A1(1'b0), .A2(_u10_n11951 ), .ZN(_u10_n20335 ) );
NAND2_X1 _u10_U8978  ( .A1(1'b0), .A2(_u10_n11927 ), .ZN(_u10_n20336 ) );
NAND4_X1 _u10_U8977  ( .A1(_u10_n20333 ), .A2(_u10_n20334 ), .A3(_u10_n20335 ), .A4(_u10_n20336 ), .ZN(_u10_n20317 ) );
NAND2_X1 _u10_U8976  ( .A1(1'b0), .A2(_u10_n11898 ), .ZN(_u10_n20329 ) );
NAND2_X1 _u10_U8975  ( .A1(1'b0), .A2(_u10_n11874 ), .ZN(_u10_n20330 ) );
NAND2_X1 _u10_U8974  ( .A1(1'b0), .A2(_u10_n11850 ), .ZN(_u10_n20331 ) );
NAND2_X1 _u10_U8973  ( .A1(1'b0), .A2(_u10_n11826 ), .ZN(_u10_n20332 ) );
NAND4_X1 _u10_U8972  ( .A1(_u10_n20329 ), .A2(_u10_n20330 ), .A3(_u10_n20331 ), .A4(_u10_n20332 ), .ZN(_u10_n20318 ) );
NAND2_X1 _u10_U8971  ( .A1(1'b0), .A2(_u10_n11802 ), .ZN(_u10_n20325 ) );
NAND2_X1 _u10_U8970  ( .A1(1'b0), .A2(_u10_n11778 ), .ZN(_u10_n20326 ) );
NAND2_X1 _u10_U8969  ( .A1(1'b0), .A2(_u10_n11754 ), .ZN(_u10_n20327 ) );
NAND2_X1 _u10_U8968  ( .A1(1'b0), .A2(_u10_n11730 ), .ZN(_u10_n20328 ) );
NAND4_X1 _u10_U8967  ( .A1(_u10_n20325 ), .A2(_u10_n20326 ), .A3(_u10_n20327 ), .A4(_u10_n20328 ), .ZN(_u10_n20319 ) );
NAND2_X1 _u10_U8966  ( .A1(1'b0), .A2(_u10_n11706 ), .ZN(_u10_n20321 ) );
NAND2_X1 _u10_U8965  ( .A1(1'b0), .A2(_u10_n11682 ), .ZN(_u10_n20322 ) );
NAND2_X1 _u10_U8964  ( .A1(1'b0), .A2(_u10_n11658 ), .ZN(_u10_n20323 ) );
NAND2_X1 _u10_U8963  ( .A1(1'b0), .A2(_u10_n11634 ), .ZN(_u10_n20324 ) );
NAND4_X1 _u10_U8962  ( .A1(_u10_n20321 ), .A2(_u10_n20322 ), .A3(_u10_n20323 ), .A4(_u10_n20324 ), .ZN(_u10_n20320 ) );
NOR4_X1 _u10_U8961  ( .A1(_u10_n20317 ), .A2(_u10_n20318 ), .A3(_u10_n20319 ), .A4(_u10_n20320 ), .ZN(_u10_n20316 ) );
NAND2_X1 _u10_U8960  ( .A1(_u10_n20315 ), .A2(_u10_n20316 ), .ZN(adr1[9]) );
NAND2_X1 _u10_U8959  ( .A1(1'b0), .A2(_u10_n12335 ), .ZN(_u10_n20311 ) );
NAND2_X1 _u10_U8958  ( .A1(1'b0), .A2(_u10_n12311 ), .ZN(_u10_n20312 ) );
NAND2_X1 _u10_U8957  ( .A1(1'b0), .A2(_u10_n12287 ), .ZN(_u10_n20313 ) );
NAND2_X1 _u10_U8956  ( .A1(1'b0), .A2(_u10_n12263 ), .ZN(_u10_n20314 ) );
NAND4_X1 _u10_U8955  ( .A1(_u10_n20311 ), .A2(_u10_n20312 ), .A3(_u10_n20313 ), .A4(_u10_n20314 ), .ZN(_u10_n20296 ) );
NAND2_X1 _u10_U8954  ( .A1(1'b0), .A2(_u10_n12239 ), .ZN(_u10_n20307 ) );
NAND2_X1 _u10_U8953  ( .A1(1'b0), .A2(_u10_n12215 ), .ZN(_u10_n20308 ) );
NAND2_X1 _u10_U8952  ( .A1(1'b0), .A2(_u10_n12191 ), .ZN(_u10_n20309 ) );
NAND2_X1 _u10_U8951  ( .A1(1'b0), .A2(_u10_n12167 ), .ZN(_u10_n20310 ) );
NAND4_X1 _u10_U8950  ( .A1(_u10_n20307 ), .A2(_u10_n20308 ), .A3(_u10_n20309 ), .A4(_u10_n20310 ), .ZN(_u10_n20297 ) );
NAND2_X1 _u10_U8949  ( .A1(1'b0), .A2(_u10_n12143 ), .ZN(_u10_n20303 ) );
NAND2_X1 _u10_U8948  ( .A1(1'b0), .A2(_u10_n12119 ), .ZN(_u10_n20304 ) );
NAND2_X1 _u10_U8947  ( .A1(1'b0), .A2(_u10_n12095 ), .ZN(_u10_n20305 ) );
NAND2_X1 _u10_U8946  ( .A1(1'b0), .A2(_u10_n12071 ), .ZN(_u10_n20306 ) );
NAND4_X1 _u10_U8945  ( .A1(_u10_n20303 ), .A2(_u10_n20304 ), .A3(_u10_n20305 ), .A4(_u10_n20306 ), .ZN(_u10_n20298 ) );
NAND2_X1 _u10_U8944  ( .A1(1'b0), .A2(_u10_n12047 ), .ZN(_u10_n20300 ) );
NAND2_X1 _u10_U8943  ( .A1(1'b0), .A2(_u10_n12023 ), .ZN(_u10_n20301 ) );
NAND2_X1 _u10_U8942  ( .A1(1'b0), .A2(_u10_n12004 ), .ZN(_u10_n20302 ) );
NAND3_X1 _u10_U8941  ( .A1(_u10_n20300 ), .A2(_u10_n20301 ), .A3(_u10_n20302 ), .ZN(_u10_n20299 ) );
NOR4_X1 _u10_U8940  ( .A1(_u10_n20296 ), .A2(_u10_n20297 ), .A3(_u10_n20298 ), .A4(_u10_n20299 ), .ZN(_u10_n20274 ) );
NAND2_X1 _u10_U8939  ( .A1(1'b0), .A2(_u10_n11995 ), .ZN(_u10_n20292 ) );
NAND2_X1 _u10_U8938  ( .A1(1'b0), .A2(_u10_n11973 ), .ZN(_u10_n20293 ) );
NAND2_X1 _u10_U8937  ( .A1(1'b0), .A2(_u10_n11949 ), .ZN(_u10_n20294 ) );
NAND2_X1 _u10_U8936  ( .A1(1'b0), .A2(_u10_n11925 ), .ZN(_u10_n20295 ) );
NAND4_X1 _u10_U8935  ( .A1(_u10_n20292 ), .A2(_u10_n20293 ), .A3(_u10_n20294 ), .A4(_u10_n20295 ), .ZN(_u10_n20276 ) );
NAND2_X1 _u10_U8934  ( .A1(1'b0), .A2(_u10_n11899 ), .ZN(_u10_n20288 ) );
NAND2_X1 _u10_U8933  ( .A1(1'b0), .A2(_u10_n11875 ), .ZN(_u10_n20289 ) );
NAND2_X1 _u10_U8932  ( .A1(1'b0), .A2(_u10_n11851 ), .ZN(_u10_n20290 ) );
NAND2_X1 _u10_U8931  ( .A1(1'b0), .A2(_u10_n11827 ), .ZN(_u10_n20291 ) );
NAND4_X1 _u10_U8930  ( .A1(_u10_n20288 ), .A2(_u10_n20289 ), .A3(_u10_n20290 ), .A4(_u10_n20291 ), .ZN(_u10_n20277 ) );
NAND2_X1 _u10_U8929  ( .A1(1'b0), .A2(_u10_n11803 ), .ZN(_u10_n20284 ) );
NAND2_X1 _u10_U8928  ( .A1(1'b0), .A2(_u10_n11779 ), .ZN(_u10_n20285 ) );
NAND2_X1 _u10_U8927  ( .A1(1'b0), .A2(_u10_n11755 ), .ZN(_u10_n20286 ) );
NAND2_X1 _u10_U8926  ( .A1(1'b0), .A2(_u10_n11731 ), .ZN(_u10_n20287 ) );
NAND4_X1 _u10_U8925  ( .A1(_u10_n20284 ), .A2(_u10_n20285 ), .A3(_u10_n20286 ), .A4(_u10_n20287 ), .ZN(_u10_n20278 ) );
NAND2_X1 _u10_U8924  ( .A1(1'b0), .A2(_u10_n11707 ), .ZN(_u10_n20280 ) );
NAND2_X1 _u10_U8923  ( .A1(1'b0), .A2(_u10_n11683 ), .ZN(_u10_n20281 ) );
NAND2_X1 _u10_U8922  ( .A1(1'b0), .A2(_u10_n11659 ), .ZN(_u10_n20282 ) );
NAND2_X1 _u10_U8921  ( .A1(1'b0), .A2(_u10_n11635 ), .ZN(_u10_n20283 ) );
NAND4_X1 _u10_U8920  ( .A1(_u10_n20280 ), .A2(_u10_n20281 ), .A3(_u10_n20282 ), .A4(_u10_n20283 ), .ZN(_u10_n20279 ) );
NOR4_X1 _u10_U8919  ( .A1(_u10_n20276 ), .A2(_u10_n20277 ), .A3(_u10_n20278 ), .A4(_u10_n20279 ), .ZN(_u10_n20275 ) );
NAND2_X1 _u10_U8918  ( .A1(_u10_n20274 ), .A2(_u10_n20275 ), .ZN(am0[0]) );
NAND2_X1 _u10_U8917  ( .A1(1'b1), .A2(_u10_n12335 ), .ZN(_u10_n20270 ) );
NAND2_X1 _u10_U8916  ( .A1(1'b1), .A2(_u10_n12311 ), .ZN(_u10_n20271 ) );
NAND2_X1 _u10_U8915  ( .A1(1'b1), .A2(_u10_n12287 ), .ZN(_u10_n20272 ) );
NAND2_X1 _u10_U8914  ( .A1(1'b1), .A2(_u10_n12263 ), .ZN(_u10_n20273 ) );
NAND4_X1 _u10_U8913  ( .A1(_u10_n20270 ), .A2(_u10_n20271 ), .A3(_u10_n20272 ), .A4(_u10_n20273 ), .ZN(_u10_n20255 ) );
NAND2_X1 _u10_U8912  ( .A1(1'b1), .A2(_u10_n12239 ), .ZN(_u10_n20266 ) );
NAND2_X1 _u10_U8911  ( .A1(1'b1), .A2(_u10_n12215 ), .ZN(_u10_n20267 ) );
NAND2_X1 _u10_U8910  ( .A1(1'b1), .A2(_u10_n12191 ), .ZN(_u10_n20268 ) );
NAND2_X1 _u10_U8909  ( .A1(1'b1), .A2(_u10_n12167 ), .ZN(_u10_n20269 ) );
NAND4_X1 _u10_U8908  ( .A1(_u10_n20266 ), .A2(_u10_n20267 ), .A3(_u10_n20268 ), .A4(_u10_n20269 ), .ZN(_u10_n20256 ) );
NAND2_X1 _u10_U8907  ( .A1(1'b1), .A2(_u10_n12143 ), .ZN(_u10_n20262 ) );
NAND2_X1 _u10_U8906  ( .A1(1'b1), .A2(_u10_n12119 ), .ZN(_u10_n20263 ) );
NAND2_X1 _u10_U8905  ( .A1(1'b1), .A2(_u10_n12095 ), .ZN(_u10_n20264 ) );
NAND2_X1 _u10_U8904  ( .A1(1'b1), .A2(_u10_n12071 ), .ZN(_u10_n20265 ) );
NAND4_X1 _u10_U8903  ( .A1(_u10_n20262 ), .A2(_u10_n20263 ), .A3(_u10_n20264 ), .A4(_u10_n20265 ), .ZN(_u10_n20257 ) );
NAND2_X1 _u10_U8902  ( .A1(1'b1), .A2(_u10_n12047 ), .ZN(_u10_n20259 ) );
NAND2_X1 _u10_U8901  ( .A1(1'b1), .A2(_u10_n12023 ), .ZN(_u10_n20260 ) );
NAND2_X1 _u10_U8900  ( .A1(1'b1), .A2(_u10_n12004 ), .ZN(_u10_n20261 ) );
NAND3_X1 _u10_U8899  ( .A1(_u10_n20259 ), .A2(_u10_n20260 ), .A3(_u10_n20261 ), .ZN(_u10_n20258 ) );
NOR4_X1 _u10_U8898  ( .A1(_u10_n20255 ), .A2(_u10_n20256 ), .A3(_u10_n20257 ), .A4(_u10_n20258 ), .ZN(_u10_n20233 ) );
NAND2_X1 _u10_U8897  ( .A1(1'b1), .A2(_u10_n11994 ), .ZN(_u10_n20251 ) );
NAND2_X1 _u10_U8896  ( .A1(1'b1), .A2(_u10_n11970 ), .ZN(_u10_n20252 ) );
NAND2_X1 _u10_U8895  ( .A1(1'b1), .A2(_u10_n11946 ), .ZN(_u10_n20253 ) );
NAND2_X1 _u10_U8894  ( .A1(1'b1), .A2(_u10_n11922 ), .ZN(_u10_n20254 ) );
NAND4_X1 _u10_U8893  ( .A1(_u10_n20251 ), .A2(_u10_n20252 ), .A3(_u10_n20253 ), .A4(_u10_n20254 ), .ZN(_u10_n20235 ) );
NAND2_X1 _u10_U8892  ( .A1(1'b1), .A2(_u10_n11902 ), .ZN(_u10_n20247 ) );
NAND2_X1 _u10_U8891  ( .A1(1'b1), .A2(_u10_n11874 ), .ZN(_u10_n20248 ) );
NAND2_X1 _u10_U8890  ( .A1(1'b1), .A2(_u10_n11854 ), .ZN(_u10_n20249 ) );
NAND2_X1 _u10_U8889  ( .A1(1'b1), .A2(_u10_n11830 ), .ZN(_u10_n20250 ) );
NAND4_X1 _u10_U8888  ( .A1(_u10_n20247 ), .A2(_u10_n20248 ), .A3(_u10_n20249 ), .A4(_u10_n20250 ), .ZN(_u10_n20236 ) );
NAND2_X1 _u10_U8887  ( .A1(1'b1), .A2(_u10_n11802 ), .ZN(_u10_n20243 ) );
NAND2_X1 _u10_U8886  ( .A1(1'b1), .A2(_u10_n11780 ), .ZN(_u10_n20244 ) );
NAND2_X1 _u10_U8885  ( .A1(1'b1), .A2(_u10_n11758 ), .ZN(_u10_n20245 ) );
NAND2_X1 _u10_U8884  ( .A1(1'b1), .A2(_u10_n11734 ), .ZN(_u10_n20246 ) );
NAND4_X1 _u10_U8883  ( .A1(_u10_n20243 ), .A2(_u10_n20244 ), .A3(_u10_n20245 ), .A4(_u10_n20246 ), .ZN(_u10_n20237 ) );
NAND2_X1 _u10_U8882  ( .A1(1'b1), .A2(_u10_n11710 ), .ZN(_u10_n20239 ) );
NAND2_X1 _u10_U8881  ( .A1(1'b1), .A2(_u10_n11686 ), .ZN(_u10_n20240 ) );
NAND2_X1 _u10_U8880  ( .A1(1'b1), .A2(_u10_n11662 ), .ZN(_u10_n20241 ) );
NAND2_X1 _u10_U8879  ( .A1(1'b1), .A2(_u10_n11638 ), .ZN(_u10_n20242 ) );
NAND4_X1 _u10_U8878  ( .A1(_u10_n20239 ), .A2(_u10_n20240 ), .A3(_u10_n20241 ), .A4(_u10_n20242 ), .ZN(_u10_n20238 ) );
NOR4_X1 _u10_U8877  ( .A1(_u10_n20235 ), .A2(_u10_n20236 ), .A3(_u10_n20237 ), .A4(_u10_n20238 ), .ZN(_u10_n20234 ) );
NAND2_X1 _u10_U8876  ( .A1(_u10_n20233 ), .A2(_u10_n20234 ), .ZN(am0[10]) );
NAND2_X1 _u10_U8875  ( .A1(1'b1), .A2(_u10_n12353 ), .ZN(_u10_n20229 ) );
NAND2_X1 _u10_U8874  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n20230 ) );
NAND2_X1 _u10_U8873  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n20231 ) );
NAND2_X1 _u10_U8872  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n20232 ) );
NAND4_X1 _u10_U8871  ( .A1(_u10_n20229 ), .A2(_u10_n20230 ), .A3(_u10_n20231 ), .A4(_u10_n20232 ), .ZN(_u10_n20214 ) );
NAND2_X1 _u10_U8870  ( .A1(1'b1), .A2(_u10_n12257 ), .ZN(_u10_n20225 ) );
NAND2_X1 _u10_U8869  ( .A1(1'b1), .A2(_u10_n12233 ), .ZN(_u10_n20226 ) );
NAND2_X1 _u10_U8868  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n20227 ) );
NAND2_X1 _u10_U8867  ( .A1(1'b1), .A2(_u10_n12185 ), .ZN(_u10_n20228 ) );
NAND4_X1 _u10_U8866  ( .A1(_u10_n20225 ), .A2(_u10_n20226 ), .A3(_u10_n20227 ), .A4(_u10_n20228 ), .ZN(_u10_n20215 ) );
NAND2_X1 _u10_U8865  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n20221 ) );
NAND2_X1 _u10_U8864  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n20222 ) );
NAND2_X1 _u10_U8863  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n20223 ) );
NAND2_X1 _u10_U8862  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n20224 ) );
NAND4_X1 _u10_U8861  ( .A1(_u10_n20221 ), .A2(_u10_n20222 ), .A3(_u10_n20223 ), .A4(_u10_n20224 ), .ZN(_u10_n20216 ) );
NAND2_X1 _u10_U8860  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n20218 ) );
NAND2_X1 _u10_U8859  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n20219 ) );
NAND2_X1 _u10_U8858  ( .A1(1'b1), .A2(_u10_n12004 ), .ZN(_u10_n20220 ) );
NAND3_X1 _u10_U8857  ( .A1(_u10_n20218 ), .A2(_u10_n20219 ), .A3(_u10_n20220 ), .ZN(_u10_n20217 ) );
NOR4_X1 _u10_U8856  ( .A1(_u10_n20214 ), .A2(_u10_n20215 ), .A3(_u10_n20216 ), .A4(_u10_n20217 ), .ZN(_u10_n20192 ) );
NAND2_X1 _u10_U8855  ( .A1(1'b1), .A2(_u10_n11998 ), .ZN(_u10_n20210 ) );
NAND2_X1 _u10_U8854  ( .A1(1'b1), .A2(_u10_n11973 ), .ZN(_u10_n20211 ) );
NAND2_X1 _u10_U8853  ( .A1(1'b1), .A2(_u10_n11949 ), .ZN(_u10_n20212 ) );
NAND2_X1 _u10_U8852  ( .A1(1'b1), .A2(_u10_n11925 ), .ZN(_u10_n20213 ) );
NAND4_X1 _u10_U8851  ( .A1(_u10_n20210 ), .A2(_u10_n20211 ), .A3(_u10_n20212 ), .A4(_u10_n20213 ), .ZN(_u10_n20194 ) );
NAND2_X1 _u10_U8850  ( .A1(1'b1), .A2(_u10_n11900 ), .ZN(_u10_n20206 ) );
NAND2_X1 _u10_U8849  ( .A1(1'b1), .A2(_u10_n11878 ), .ZN(_u10_n20207 ) );
NAND2_X1 _u10_U8848  ( .A1(1'b1), .A2(_u10_n11852 ), .ZN(_u10_n20208 ) );
NAND2_X1 _u10_U8847  ( .A1(1'b1), .A2(_u10_n11828 ), .ZN(_u10_n20209 ) );
NAND4_X1 _u10_U8846  ( .A1(_u10_n20206 ), .A2(_u10_n20207 ), .A3(_u10_n20208 ), .A4(_u10_n20209 ), .ZN(_u10_n20195 ) );
NAND2_X1 _u10_U8845  ( .A1(1'b1), .A2(_u10_n11806 ), .ZN(_u10_n20202 ) );
NAND2_X1 _u10_U8844  ( .A1(1'b1), .A2(_u10_n11782 ), .ZN(_u10_n20203 ) );
NAND2_X1 _u10_U8843  ( .A1(1'b1), .A2(_u10_n11759 ), .ZN(_u10_n20204 ) );
NAND2_X1 _u10_U8842  ( .A1(1'b1), .A2(_u10_n11735 ), .ZN(_u10_n20205 ) );
NAND4_X1 _u10_U8841  ( .A1(_u10_n20202 ), .A2(_u10_n20203 ), .A3(_u10_n20204 ), .A4(_u10_n20205 ), .ZN(_u10_n20196 ) );
NAND2_X1 _u10_U8840  ( .A1(1'b1), .A2(_u10_n11711 ), .ZN(_u10_n20198 ) );
NAND2_X1 _u10_U8839  ( .A1(1'b1), .A2(_u10_n11687 ), .ZN(_u10_n20199 ) );
NAND2_X1 _u10_U8838  ( .A1(1'b1), .A2(_u10_n11660 ), .ZN(_u10_n20200 ) );
NAND2_X1 _u10_U8837  ( .A1(1'b1), .A2(_u10_n11636 ), .ZN(_u10_n20201 ) );
NAND4_X1 _u10_U8836  ( .A1(_u10_n20198 ), .A2(_u10_n20199 ), .A3(_u10_n20200 ), .A4(_u10_n20201 ), .ZN(_u10_n20197 ) );
NOR4_X1 _u10_U8835  ( .A1(_u10_n20194 ), .A2(_u10_n20195 ), .A3(_u10_n20196 ), .A4(_u10_n20197 ), .ZN(_u10_n20193 ) );
NAND2_X1 _u10_U8834  ( .A1(_u10_n20192 ), .A2(_u10_n20193 ), .ZN(am0[11]) );
NAND2_X1 _u10_U8833  ( .A1(1'b1), .A2(_u10_n12430 ), .ZN(_u10_n20188 ) );
NAND2_X1 _u10_U8832  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n20189 ) );
NAND2_X1 _u10_U8831  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n20190 ) );
NAND2_X1 _u10_U8830  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n20191 ) );
NAND4_X1 _u10_U8829  ( .A1(_u10_n20188 ), .A2(_u10_n20189 ), .A3(_u10_n20190 ), .A4(_u10_n20191 ), .ZN(_u10_n20173 ) );
NAND2_X1 _u10_U8828  ( .A1(1'b1), .A2(_u10_n12422 ), .ZN(_u10_n20184 ) );
NAND2_X1 _u10_U8827  ( .A1(1'b1), .A2(_u10_n12421 ), .ZN(_u10_n20185 ) );
NAND2_X1 _u10_U8826  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n20186 ) );
NAND2_X1 _u10_U8825  ( .A1(1'b1), .A2(_u10_n12419 ), .ZN(_u10_n20187 ) );
NAND4_X1 _u10_U8824  ( .A1(_u10_n20184 ), .A2(_u10_n20185 ), .A3(_u10_n20186 ), .A4(_u10_n20187 ), .ZN(_u10_n20174 ) );
NAND2_X1 _u10_U8823  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n20180 ) );
NAND2_X1 _u10_U8822  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n20181 ) );
NAND2_X1 _u10_U8821  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n20182 ) );
NAND2_X1 _u10_U8820  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n20183 ) );
NAND4_X1 _u10_U8819  ( .A1(_u10_n20180 ), .A2(_u10_n20181 ), .A3(_u10_n20182 ), .A4(_u10_n20183 ), .ZN(_u10_n20175 ) );
NAND2_X1 _u10_U8818  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n20177 ) );
NAND2_X1 _u10_U8817  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n20178 ) );
NAND2_X1 _u10_U8816  ( .A1(1'b1), .A2(_u10_n12004 ), .ZN(_u10_n20179 ) );
NAND3_X1 _u10_U8815  ( .A1(_u10_n20177 ), .A2(_u10_n20178 ), .A3(_u10_n20179 ), .ZN(_u10_n20176 ) );
NOR4_X1 _u10_U8814  ( .A1(_u10_n20173 ), .A2(_u10_n20174 ), .A3(_u10_n20175 ), .A4(_u10_n20176 ), .ZN(_u10_n20151 ) );
NAND2_X1 _u10_U8813  ( .A1(1'b1), .A2(_u10_n11999 ), .ZN(_u10_n20169 ) );
NAND2_X1 _u10_U8812  ( .A1(1'b1), .A2(_u10_n11974 ), .ZN(_u10_n20170 ) );
NAND2_X1 _u10_U8811  ( .A1(1'b1), .A2(_u10_n11945 ), .ZN(_u10_n20171 ) );
NAND2_X1 _u10_U8810  ( .A1(1'b1), .A2(_u10_n11921 ), .ZN(_u10_n20172 ) );
NAND4_X1 _u10_U8809  ( .A1(_u10_n20169 ), .A2(_u10_n20170 ), .A3(_u10_n20171 ), .A4(_u10_n20172 ), .ZN(_u10_n20153 ) );
NAND2_X1 _u10_U8808  ( .A1(1'b1), .A2(_u10_n11903 ), .ZN(_u10_n20165 ) );
NAND2_X1 _u10_U8807  ( .A1(1'b1), .A2(_u10_n11879 ), .ZN(_u10_n20166 ) );
NAND2_X1 _u10_U8806  ( .A1(1'b1), .A2(_u10_n11852 ), .ZN(_u10_n20167 ) );
NAND2_X1 _u10_U8805  ( .A1(1'b1), .A2(_u10_n11831 ), .ZN(_u10_n20168 ) );
NAND4_X1 _u10_U8804  ( .A1(_u10_n20165 ), .A2(_u10_n20166 ), .A3(_u10_n20167 ), .A4(_u10_n20168 ), .ZN(_u10_n20154 ) );
NAND2_X1 _u10_U8803  ( .A1(1'b1), .A2(_u10_n11807 ), .ZN(_u10_n20161 ) );
NAND2_X1 _u10_U8802  ( .A1(1'b1), .A2(_u10_n11783 ), .ZN(_u10_n20162 ) );
NAND2_X1 _u10_U8801  ( .A1(1'b1), .A2(_u10_n11757 ), .ZN(_u10_n20163 ) );
NAND2_X1 _u10_U8800  ( .A1(1'b1), .A2(_u10_n11733 ), .ZN(_u10_n20164 ) );
NAND4_X1 _u10_U8799  ( .A1(_u10_n20161 ), .A2(_u10_n20162 ), .A3(_u10_n20163 ), .A4(_u10_n20164 ), .ZN(_u10_n20155 ) );
NAND2_X1 _u10_U8798  ( .A1(1'b1), .A2(_u10_n11709 ), .ZN(_u10_n20157 ) );
NAND2_X1 _u10_U8797  ( .A1(1'b1), .A2(_u10_n11685 ), .ZN(_u10_n20158 ) );
NAND2_X1 _u10_U8796  ( .A1(1'b1), .A2(_u10_n11660 ), .ZN(_u10_n20159 ) );
NAND2_X1 _u10_U8795  ( .A1(1'b1), .A2(_u10_n11636 ), .ZN(_u10_n20160 ) );
NAND4_X1 _u10_U8794  ( .A1(_u10_n20157 ), .A2(_u10_n20158 ), .A3(_u10_n20159 ), .A4(_u10_n20160 ), .ZN(_u10_n20156 ) );
NOR4_X1 _u10_U8793  ( .A1(_u10_n20153 ), .A2(_u10_n20154 ), .A3(_u10_n20155 ), .A4(_u10_n20156 ), .ZN(_u10_n20152 ) );
NAND2_X1 _u10_U8792  ( .A1(_u10_n20151 ), .A2(_u10_n20152 ), .ZN(am0[12]) );
NAND2_X1 _u10_U8791  ( .A1(1'b1), .A2(_u10_n12352 ), .ZN(_u10_n20147 ) );
NAND2_X1 _u10_U8790  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n20148 ) );
NAND2_X1 _u10_U8789  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n20149 ) );
NAND2_X1 _u10_U8788  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n20150 ) );
NAND4_X1 _u10_U8787  ( .A1(_u10_n20147 ), .A2(_u10_n20148 ), .A3(_u10_n20149 ), .A4(_u10_n20150 ), .ZN(_u10_n20132 ) );
NAND2_X1 _u10_U8786  ( .A1(1'b1), .A2(_u10_n12256 ), .ZN(_u10_n20143 ) );
NAND2_X1 _u10_U8785  ( .A1(1'b1), .A2(_u10_n12232 ), .ZN(_u10_n20144 ) );
NAND2_X1 _u10_U8784  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n20145 ) );
NAND2_X1 _u10_U8783  ( .A1(1'b1), .A2(_u10_n12184 ), .ZN(_u10_n20146 ) );
NAND4_X1 _u10_U8782  ( .A1(_u10_n20143 ), .A2(_u10_n20144 ), .A3(_u10_n20145 ), .A4(_u10_n20146 ), .ZN(_u10_n20133 ) );
NAND2_X1 _u10_U8781  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n20139 ) );
NAND2_X1 _u10_U8780  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n20140 ) );
NAND2_X1 _u10_U8779  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n20141 ) );
NAND2_X1 _u10_U8778  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n20142 ) );
NAND4_X1 _u10_U8777  ( .A1(_u10_n20139 ), .A2(_u10_n20140 ), .A3(_u10_n20141 ), .A4(_u10_n20142 ), .ZN(_u10_n20134 ) );
NAND2_X1 _u10_U8776  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n20136 ) );
NAND2_X1 _u10_U8775  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n20137 ) );
NAND2_X1 _u10_U8774  ( .A1(1'b1), .A2(_u10_n12004 ), .ZN(_u10_n20138 ) );
NAND3_X1 _u10_U8773  ( .A1(_u10_n20136 ), .A2(_u10_n20137 ), .A3(_u10_n20138 ), .ZN(_u10_n20135 ) );
NOR4_X1 _u10_U8772  ( .A1(_u10_n20132 ), .A2(_u10_n20133 ), .A3(_u10_n20134 ), .A4(_u10_n20135 ), .ZN(_u10_n20110 ) );
NAND2_X1 _u10_U8771  ( .A1(1'b1), .A2(_u10_n11997 ), .ZN(_u10_n20128 ) );
NAND2_X1 _u10_U8770  ( .A1(1'b1), .A2(_u10_n11972 ), .ZN(_u10_n20129 ) );
NAND2_X1 _u10_U8769  ( .A1(1'b1), .A2(_u10_n11950 ), .ZN(_u10_n20130 ) );
NAND2_X1 _u10_U8768  ( .A1(1'b1), .A2(_u10_n11926 ), .ZN(_u10_n20131 ) );
NAND4_X1 _u10_U8767  ( .A1(_u10_n20128 ), .A2(_u10_n20129 ), .A3(_u10_n20130 ), .A4(_u10_n20131 ), .ZN(_u10_n20112 ) );
NAND2_X1 _u10_U8766  ( .A1(1'b1), .A2(_u10_n11901 ), .ZN(_u10_n20124 ) );
NAND2_X1 _u10_U8765  ( .A1(1'b1), .A2(_u10_n11877 ), .ZN(_u10_n20125 ) );
NAND2_X1 _u10_U8764  ( .A1(1'b1), .A2(_u10_n11855 ), .ZN(_u10_n20126 ) );
NAND2_X1 _u10_U8763  ( .A1(1'b1), .A2(_u10_n11829 ), .ZN(_u10_n20127 ) );
NAND4_X1 _u10_U8762  ( .A1(_u10_n20124 ), .A2(_u10_n20125 ), .A3(_u10_n20126 ), .A4(_u10_n20127 ), .ZN(_u10_n20113 ) );
NAND2_X1 _u10_U8761  ( .A1(1'b1), .A2(_u10_n11805 ), .ZN(_u10_n20120 ) );
NAND2_X1 _u10_U8760  ( .A1(1'b1), .A2(_u10_n11781 ), .ZN(_u10_n20121 ) );
NAND2_X1 _u10_U8759  ( .A1(1'b1), .A2(_u10_n11753 ), .ZN(_u10_n20122 ) );
NAND2_X1 _u10_U8758  ( .A1(1'b1), .A2(_u10_n11729 ), .ZN(_u10_n20123 ) );
NAND4_X1 _u10_U8757  ( .A1(_u10_n20120 ), .A2(_u10_n20121 ), .A3(_u10_n20122 ), .A4(_u10_n20123 ), .ZN(_u10_n20114 ) );
NAND2_X1 _u10_U8756  ( .A1(1'b1), .A2(_u10_n11705 ), .ZN(_u10_n20116 ) );
NAND2_X1 _u10_U8755  ( .A1(1'b1), .A2(_u10_n11681 ), .ZN(_u10_n20117 ) );
NAND2_X1 _u10_U8754  ( .A1(1'b1), .A2(_u10_n11663 ), .ZN(_u10_n20118 ) );
NAND2_X1 _u10_U8753  ( .A1(1'b1), .A2(_u10_n11639 ), .ZN(_u10_n20119 ) );
NAND4_X1 _u10_U8752  ( .A1(_u10_n20116 ), .A2(_u10_n20117 ), .A3(_u10_n20118 ), .A4(_u10_n20119 ), .ZN(_u10_n20115 ) );
NOR4_X1 _u10_U8751  ( .A1(_u10_n20112 ), .A2(_u10_n20113 ), .A3(_u10_n20114 ), .A4(_u10_n20115 ), .ZN(_u10_n20111 ) );
NAND2_X1 _u10_U8750  ( .A1(_u10_n20110 ), .A2(_u10_n20111 ), .ZN(am0[13]) );
NAND2_X1 _u10_U8749  ( .A1(1'b1), .A2(_u10_n12353 ), .ZN(_u10_n20106 ) );
NAND2_X1 _u10_U8748  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n20107 ) );
NAND2_X1 _u10_U8747  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n20108 ) );
NAND2_X1 _u10_U8746  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n20109 ) );
NAND4_X1 _u10_U8745  ( .A1(_u10_n20106 ), .A2(_u10_n20107 ), .A3(_u10_n20108 ), .A4(_u10_n20109 ), .ZN(_u10_n20091 ) );
NAND2_X1 _u10_U8744  ( .A1(1'b1), .A2(_u10_n12257 ), .ZN(_u10_n20102 ) );
NAND2_X1 _u10_U8743  ( .A1(1'b1), .A2(_u10_n12233 ), .ZN(_u10_n20103 ) );
NAND2_X1 _u10_U8742  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n20104 ) );
NAND2_X1 _u10_U8741  ( .A1(1'b1), .A2(_u10_n12185 ), .ZN(_u10_n20105 ) );
NAND4_X1 _u10_U8740  ( .A1(_u10_n20102 ), .A2(_u10_n20103 ), .A3(_u10_n20104 ), .A4(_u10_n20105 ), .ZN(_u10_n20092 ) );
NAND2_X1 _u10_U8739  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n20098 ) );
NAND2_X1 _u10_U8738  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n20099 ) );
NAND2_X1 _u10_U8737  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n20100 ) );
NAND2_X1 _u10_U8736  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n20101 ) );
NAND4_X1 _u10_U8735  ( .A1(_u10_n20098 ), .A2(_u10_n20099 ), .A3(_u10_n20100 ), .A4(_u10_n20101 ), .ZN(_u10_n20093 ) );
NAND2_X1 _u10_U8734  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n20095 ) );
NAND2_X1 _u10_U8733  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n20096 ) );
NAND2_X1 _u10_U8732  ( .A1(1'b1), .A2(_u10_n12004 ), .ZN(_u10_n20097 ) );
NAND3_X1 _u10_U8731  ( .A1(_u10_n20095 ), .A2(_u10_n20096 ), .A3(_u10_n20097 ), .ZN(_u10_n20094 ) );
NOR4_X1 _u10_U8730  ( .A1(_u10_n20091 ), .A2(_u10_n20092 ), .A3(_u10_n20093 ), .A4(_u10_n20094 ), .ZN(_u10_n20069 ) );
NAND2_X1 _u10_U8729  ( .A1(1'b1), .A2(_u10_n11996 ), .ZN(_u10_n20087 ) );
NAND2_X1 _u10_U8728  ( .A1(1'b1), .A2(_u10_n11972 ), .ZN(_u10_n20088 ) );
NAND2_X1 _u10_U8727  ( .A1(1'b1), .A2(_u10_n11948 ), .ZN(_u10_n20089 ) );
NAND2_X1 _u10_U8726  ( .A1(1'b1), .A2(_u10_n11924 ), .ZN(_u10_n20090 ) );
NAND4_X1 _u10_U8725  ( .A1(_u10_n20087 ), .A2(_u10_n20088 ), .A3(_u10_n20089 ), .A4(_u10_n20090 ), .ZN(_u10_n20071 ) );
NAND2_X1 _u10_U8724  ( .A1(1'b1), .A2(_u10_n11900 ), .ZN(_u10_n20083 ) );
NAND2_X1 _u10_U8723  ( .A1(1'b1), .A2(_u10_n11876 ), .ZN(_u10_n20084 ) );
NAND2_X1 _u10_U8722  ( .A1(1'b1), .A2(_u10_n11852 ), .ZN(_u10_n20085 ) );
NAND2_X1 _u10_U8721  ( .A1(1'b1), .A2(_u10_n11828 ), .ZN(_u10_n20086 ) );
NAND4_X1 _u10_U8720  ( .A1(_u10_n20083 ), .A2(_u10_n20084 ), .A3(_u10_n20085 ), .A4(_u10_n20086 ), .ZN(_u10_n20072 ) );
NAND2_X1 _u10_U8719  ( .A1(1'b1), .A2(_u10_n11804 ), .ZN(_u10_n20079 ) );
NAND2_X1 _u10_U8718  ( .A1(1'b1), .A2(_u10_n11780 ), .ZN(_u10_n20080 ) );
NAND2_X1 _u10_U8717  ( .A1(1'b1), .A2(_u10_n11756 ), .ZN(_u10_n20081 ) );
NAND2_X1 _u10_U8716  ( .A1(1'b1), .A2(_u10_n11732 ), .ZN(_u10_n20082 ) );
NAND4_X1 _u10_U8715  ( .A1(_u10_n20079 ), .A2(_u10_n20080 ), .A3(_u10_n20081 ), .A4(_u10_n20082 ), .ZN(_u10_n20073 ) );
NAND2_X1 _u10_U8714  ( .A1(1'b1), .A2(_u10_n11708 ), .ZN(_u10_n20075 ) );
NAND2_X1 _u10_U8713  ( .A1(1'b1), .A2(_u10_n11684 ), .ZN(_u10_n20076 ) );
NAND2_X1 _u10_U8712  ( .A1(1'b1), .A2(_u10_n11660 ), .ZN(_u10_n20077 ) );
NAND2_X1 _u10_U8711  ( .A1(1'b1), .A2(_u10_n11636 ), .ZN(_u10_n20078 ) );
NAND4_X1 _u10_U8710  ( .A1(_u10_n20075 ), .A2(_u10_n20076 ), .A3(_u10_n20077 ), .A4(_u10_n20078 ), .ZN(_u10_n20074 ) );
NOR4_X1 _u10_U8709  ( .A1(_u10_n20071 ), .A2(_u10_n20072 ), .A3(_u10_n20073 ), .A4(_u10_n20074 ), .ZN(_u10_n20070 ) );
NAND2_X1 _u10_U8708  ( .A1(_u10_n20069 ), .A2(_u10_n20070 ), .ZN(am0[14]) );
NAND2_X1 _u10_U8707  ( .A1(1'b1), .A2(_u10_n12356 ), .ZN(_u10_n20065 ) );
NAND2_X1 _u10_U8706  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n20066 ) );
NAND2_X1 _u10_U8705  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n20067 ) );
NAND2_X1 _u10_U8704  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n20068 ) );
NAND4_X1 _u10_U8703  ( .A1(_u10_n20065 ), .A2(_u10_n20066 ), .A3(_u10_n20067 ), .A4(_u10_n20068 ), .ZN(_u10_n20050 ) );
NAND2_X1 _u10_U8702  ( .A1(1'b1), .A2(_u10_n12260 ), .ZN(_u10_n20061 ) );
NAND2_X1 _u10_U8701  ( .A1(1'b1), .A2(_u10_n12236 ), .ZN(_u10_n20062 ) );
NAND2_X1 _u10_U8700  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n20063 ) );
NAND2_X1 _u10_U8699  ( .A1(1'b1), .A2(_u10_n12188 ), .ZN(_u10_n20064 ) );
NAND4_X1 _u10_U8698  ( .A1(_u10_n20061 ), .A2(_u10_n20062 ), .A3(_u10_n20063 ), .A4(_u10_n20064 ), .ZN(_u10_n20051 ) );
NAND2_X1 _u10_U8697  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n20057 ) );
NAND2_X1 _u10_U8696  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n20058 ) );
NAND2_X1 _u10_U8695  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n20059 ) );
NAND2_X1 _u10_U8694  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n20060 ) );
NAND4_X1 _u10_U8693  ( .A1(_u10_n20057 ), .A2(_u10_n20058 ), .A3(_u10_n20059 ), .A4(_u10_n20060 ), .ZN(_u10_n20052 ) );
NAND2_X1 _u10_U8692  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n20054 ) );
NAND2_X1 _u10_U8691  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n20055 ) );
NAND2_X1 _u10_U8690  ( .A1(1'b1), .A2(_u10_n12004 ), .ZN(_u10_n20056 ) );
NAND3_X1 _u10_U8689  ( .A1(_u10_n20054 ), .A2(_u10_n20055 ), .A3(_u10_n20056 ), .ZN(_u10_n20053 ) );
NOR4_X1 _u10_U8688  ( .A1(_u10_n20050 ), .A2(_u10_n20051 ), .A3(_u10_n20052 ), .A4(_u10_n20053 ), .ZN(_u10_n20028 ) );
NAND2_X1 _u10_U8687  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n20046 ) );
NAND2_X1 _u10_U8686  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n20047 ) );
NAND2_X1 _u10_U8685  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n20048 ) );
NAND2_X1 _u10_U8684  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n20049 ) );
NAND4_X1 _u10_U8683  ( .A1(_u10_n20046 ), .A2(_u10_n20047 ), .A3(_u10_n20048 ), .A4(_u10_n20049 ), .ZN(_u10_n20030 ) );
NAND2_X1 _u10_U8682  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n20042 ) );
NAND2_X1 _u10_U8681  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n20043 ) );
NAND2_X1 _u10_U8680  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n20044 ) );
NAND2_X1 _u10_U8679  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n20045 ) );
NAND4_X1 _u10_U8678  ( .A1(_u10_n20042 ), .A2(_u10_n20043 ), .A3(_u10_n20044 ), .A4(_u10_n20045 ), .ZN(_u10_n20031 ) );
NAND2_X1 _u10_U8677  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n20038 ) );
NAND2_X1 _u10_U8676  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n20039 ) );
NAND2_X1 _u10_U8675  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n20040 ) );
NAND2_X1 _u10_U8674  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n20041 ) );
NAND4_X1 _u10_U8673  ( .A1(_u10_n20038 ), .A2(_u10_n20039 ), .A3(_u10_n20040 ), .A4(_u10_n20041 ), .ZN(_u10_n20032 ) );
NAND2_X1 _u10_U8672  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n20034 ) );
NAND2_X1 _u10_U8671  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n20035 ) );
NAND2_X1 _u10_U8670  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n20036 ) );
NAND2_X1 _u10_U8669  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n20037 ) );
NAND4_X1 _u10_U8668  ( .A1(_u10_n20034 ), .A2(_u10_n20035 ), .A3(_u10_n20036 ), .A4(_u10_n20037 ), .ZN(_u10_n20033 ) );
NOR4_X1 _u10_U8667  ( .A1(_u10_n20030 ), .A2(_u10_n20031 ), .A3(_u10_n20032 ), .A4(_u10_n20033 ), .ZN(_u10_n20029 ) );
NAND2_X1 _u10_U8666  ( .A1(_u10_n20028 ), .A2(_u10_n20029 ), .ZN(am0[15]) );
NAND2_X1 _u10_U8665  ( .A1(1'b1), .A2(_u10_n12354 ), .ZN(_u10_n20024 ) );
NAND2_X1 _u10_U8664  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n20025 ) );
NAND2_X1 _u10_U8663  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n20026 ) );
NAND2_X1 _u10_U8662  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n20027 ) );
NAND4_X1 _u10_U8661  ( .A1(_u10_n20024 ), .A2(_u10_n20025 ), .A3(_u10_n20026 ), .A4(_u10_n20027 ), .ZN(_u10_n20009 ) );
NAND2_X1 _u10_U8660  ( .A1(1'b1), .A2(_u10_n12258 ), .ZN(_u10_n20020 ) );
NAND2_X1 _u10_U8659  ( .A1(1'b1), .A2(_u10_n12234 ), .ZN(_u10_n20021 ) );
NAND2_X1 _u10_U8658  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n20022 ) );
NAND2_X1 _u10_U8657  ( .A1(1'b1), .A2(_u10_n12186 ), .ZN(_u10_n20023 ) );
NAND4_X1 _u10_U8656  ( .A1(_u10_n20020 ), .A2(_u10_n20021 ), .A3(_u10_n20022 ), .A4(_u10_n20023 ), .ZN(_u10_n20010 ) );
NAND2_X1 _u10_U8655  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n20016 ) );
NAND2_X1 _u10_U8654  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n20017 ) );
NAND2_X1 _u10_U8653  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n20018 ) );
NAND2_X1 _u10_U8652  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n20019 ) );
NAND4_X1 _u10_U8651  ( .A1(_u10_n20016 ), .A2(_u10_n20017 ), .A3(_u10_n20018 ), .A4(_u10_n20019 ), .ZN(_u10_n20011 ) );
NAND2_X1 _u10_U8650  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n20013 ) );
NAND2_X1 _u10_U8649  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n20014 ) );
NAND2_X1 _u10_U8648  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n20015 ) );
NAND3_X1 _u10_U8647  ( .A1(_u10_n20013 ), .A2(_u10_n20014 ), .A3(_u10_n20015 ), .ZN(_u10_n20012 ) );
NOR4_X1 _u10_U8646  ( .A1(_u10_n20009 ), .A2(_u10_n20010 ), .A3(_u10_n20011 ), .A4(_u10_n20012 ), .ZN(_u10_n19987 ) );
NAND2_X1 _u10_U8645  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n20005 ) );
NAND2_X1 _u10_U8644  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n20006 ) );
NAND2_X1 _u10_U8643  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n20007 ) );
NAND2_X1 _u10_U8642  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n20008 ) );
NAND4_X1 _u10_U8641  ( .A1(_u10_n20005 ), .A2(_u10_n20006 ), .A3(_u10_n20007 ), .A4(_u10_n20008 ), .ZN(_u10_n19989 ) );
NAND2_X1 _u10_U8640  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n20001 ) );
NAND2_X1 _u10_U8639  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n20002 ) );
NAND2_X1 _u10_U8638  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n20003 ) );
NAND2_X1 _u10_U8637  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n20004 ) );
NAND4_X1 _u10_U8636  ( .A1(_u10_n20001 ), .A2(_u10_n20002 ), .A3(_u10_n20003 ), .A4(_u10_n20004 ), .ZN(_u10_n19990 ) );
NAND2_X1 _u10_U8635  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n19997 ) );
NAND2_X1 _u10_U8634  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n19998 ) );
NAND2_X1 _u10_U8633  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n19999 ) );
NAND2_X1 _u10_U8632  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n20000 ) );
NAND4_X1 _u10_U8631  ( .A1(_u10_n19997 ), .A2(_u10_n19998 ), .A3(_u10_n19999 ), .A4(_u10_n20000 ), .ZN(_u10_n19991 ) );
NAND2_X1 _u10_U8630  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n19993 ) );
NAND2_X1 _u10_U8629  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n19994 ) );
NAND2_X1 _u10_U8628  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n19995 ) );
NAND2_X1 _u10_U8627  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n19996 ) );
NAND4_X1 _u10_U8626  ( .A1(_u10_n19993 ), .A2(_u10_n19994 ), .A3(_u10_n19995 ), .A4(_u10_n19996 ), .ZN(_u10_n19992 ) );
NOR4_X1 _u10_U8625  ( .A1(_u10_n19989 ), .A2(_u10_n19990 ), .A3(_u10_n19991 ), .A4(_u10_n19992 ), .ZN(_u10_n19988 ) );
NAND2_X1 _u10_U8624  ( .A1(_u10_n19987 ), .A2(_u10_n19988 ), .ZN(am0[16]) );
NAND2_X1 _u10_U8623  ( .A1(1'b1), .A2(_u10_n12355 ), .ZN(_u10_n19983 ) );
NAND2_X1 _u10_U8622  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n19984 ) );
NAND2_X1 _u10_U8621  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n19985 ) );
NAND2_X1 _u10_U8620  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n19986 ) );
NAND4_X1 _u10_U8619  ( .A1(_u10_n19983 ), .A2(_u10_n19984 ), .A3(_u10_n19985 ), .A4(_u10_n19986 ), .ZN(_u10_n19968 ) );
NAND2_X1 _u10_U8618  ( .A1(1'b1), .A2(_u10_n12259 ), .ZN(_u10_n19979 ) );
NAND2_X1 _u10_U8617  ( .A1(1'b1), .A2(_u10_n12235 ), .ZN(_u10_n19980 ) );
NAND2_X1 _u10_U8616  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n19981 ) );
NAND2_X1 _u10_U8615  ( .A1(1'b1), .A2(_u10_n12187 ), .ZN(_u10_n19982 ) );
NAND4_X1 _u10_U8614  ( .A1(_u10_n19979 ), .A2(_u10_n19980 ), .A3(_u10_n19981 ), .A4(_u10_n19982 ), .ZN(_u10_n19969 ) );
NAND2_X1 _u10_U8613  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n19975 ) );
NAND2_X1 _u10_U8612  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n19976 ) );
NAND2_X1 _u10_U8611  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n19977 ) );
NAND2_X1 _u10_U8610  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n19978 ) );
NAND4_X1 _u10_U8609  ( .A1(_u10_n19975 ), .A2(_u10_n19976 ), .A3(_u10_n19977 ), .A4(_u10_n19978 ), .ZN(_u10_n19970 ) );
NAND2_X1 _u10_U8608  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n19972 ) );
NAND2_X1 _u10_U8607  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n19973 ) );
NAND2_X1 _u10_U8606  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19974 ) );
NAND3_X1 _u10_U8605  ( .A1(_u10_n19972 ), .A2(_u10_n19973 ), .A3(_u10_n19974 ), .ZN(_u10_n19971 ) );
NOR4_X1 _u10_U8604  ( .A1(_u10_n19968 ), .A2(_u10_n19969 ), .A3(_u10_n19970 ), .A4(_u10_n19971 ), .ZN(_u10_n19946 ) );
NAND2_X1 _u10_U8603  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n19964 ) );
NAND2_X1 _u10_U8602  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n19965 ) );
NAND2_X1 _u10_U8601  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n19966 ) );
NAND2_X1 _u10_U8600  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n19967 ) );
NAND4_X1 _u10_U8599  ( .A1(_u10_n19964 ), .A2(_u10_n19965 ), .A3(_u10_n19966 ), .A4(_u10_n19967 ), .ZN(_u10_n19948 ) );
NAND2_X1 _u10_U8598  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n19960 ) );
NAND2_X1 _u10_U8597  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n19961 ) );
NAND2_X1 _u10_U8596  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n19962 ) );
NAND2_X1 _u10_U8595  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n19963 ) );
NAND4_X1 _u10_U8594  ( .A1(_u10_n19960 ), .A2(_u10_n19961 ), .A3(_u10_n19962 ), .A4(_u10_n19963 ), .ZN(_u10_n19949 ) );
NAND2_X1 _u10_U8593  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n19956 ) );
NAND2_X1 _u10_U8592  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n19957 ) );
NAND2_X1 _u10_U8591  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n19958 ) );
NAND2_X1 _u10_U8590  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n19959 ) );
NAND4_X1 _u10_U8589  ( .A1(_u10_n19956 ), .A2(_u10_n19957 ), .A3(_u10_n19958 ), .A4(_u10_n19959 ), .ZN(_u10_n19950 ) );
NAND2_X1 _u10_U8588  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n19952 ) );
NAND2_X1 _u10_U8587  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n19953 ) );
NAND2_X1 _u10_U8586  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n19954 ) );
NAND2_X1 _u10_U8585  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n19955 ) );
NAND4_X1 _u10_U8584  ( .A1(_u10_n19952 ), .A2(_u10_n19953 ), .A3(_u10_n19954 ), .A4(_u10_n19955 ), .ZN(_u10_n19951 ) );
NOR4_X1 _u10_U8583  ( .A1(_u10_n19948 ), .A2(_u10_n19949 ), .A3(_u10_n19950 ), .A4(_u10_n19951 ), .ZN(_u10_n19947 ) );
NAND2_X1 _u10_U8582  ( .A1(_u10_n19946 ), .A2(_u10_n19947 ), .ZN(am0[17]) );
NAND2_X1 _u10_U8581  ( .A1(1'b1), .A2(_u10_n12353 ), .ZN(_u10_n19942 ) );
NAND2_X1 _u10_U8580  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n19943 ) );
NAND2_X1 _u10_U8579  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n19944 ) );
NAND2_X1 _u10_U8578  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n19945 ) );
NAND4_X1 _u10_U8577  ( .A1(_u10_n19942 ), .A2(_u10_n19943 ), .A3(_u10_n19944 ), .A4(_u10_n19945 ), .ZN(_u10_n19927 ) );
NAND2_X1 _u10_U8576  ( .A1(1'b1), .A2(_u10_n12257 ), .ZN(_u10_n19938 ) );
NAND2_X1 _u10_U8575  ( .A1(1'b1), .A2(_u10_n12233 ), .ZN(_u10_n19939 ) );
NAND2_X1 _u10_U8574  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n19940 ) );
NAND2_X1 _u10_U8573  ( .A1(1'b1), .A2(_u10_n12185 ), .ZN(_u10_n19941 ) );
NAND4_X1 _u10_U8572  ( .A1(_u10_n19938 ), .A2(_u10_n19939 ), .A3(_u10_n19940 ), .A4(_u10_n19941 ), .ZN(_u10_n19928 ) );
NAND2_X1 _u10_U8571  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n19934 ) );
NAND2_X1 _u10_U8570  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n19935 ) );
NAND2_X1 _u10_U8569  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n19936 ) );
NAND2_X1 _u10_U8568  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n19937 ) );
NAND4_X1 _u10_U8567  ( .A1(_u10_n19934 ), .A2(_u10_n19935 ), .A3(_u10_n19936 ), .A4(_u10_n19937 ), .ZN(_u10_n19929 ) );
NAND2_X1 _u10_U8566  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n19931 ) );
NAND2_X1 _u10_U8565  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n19932 ) );
NAND2_X1 _u10_U8564  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19933 ) );
NAND3_X1 _u10_U8563  ( .A1(_u10_n19931 ), .A2(_u10_n19932 ), .A3(_u10_n19933 ), .ZN(_u10_n19930 ) );
NOR4_X1 _u10_U8562  ( .A1(_u10_n19927 ), .A2(_u10_n19928 ), .A3(_u10_n19929 ), .A4(_u10_n19930 ), .ZN(_u10_n19905 ) );
NAND2_X1 _u10_U8561  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n19923 ) );
NAND2_X1 _u10_U8560  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n19924 ) );
NAND2_X1 _u10_U8559  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n19925 ) );
NAND2_X1 _u10_U8558  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n19926 ) );
NAND4_X1 _u10_U8557  ( .A1(_u10_n19923 ), .A2(_u10_n19924 ), .A3(_u10_n19925 ), .A4(_u10_n19926 ), .ZN(_u10_n19907 ) );
NAND2_X1 _u10_U8556  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n19919 ) );
NAND2_X1 _u10_U8555  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n19920 ) );
NAND2_X1 _u10_U8554  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n19921 ) );
NAND2_X1 _u10_U8553  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n19922 ) );
NAND4_X1 _u10_U8552  ( .A1(_u10_n19919 ), .A2(_u10_n19920 ), .A3(_u10_n19921 ), .A4(_u10_n19922 ), .ZN(_u10_n19908 ) );
NAND2_X1 _u10_U8551  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n19915 ) );
NAND2_X1 _u10_U8550  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n19916 ) );
NAND2_X1 _u10_U8549  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n19917 ) );
NAND2_X1 _u10_U8548  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n19918 ) );
NAND4_X1 _u10_U8547  ( .A1(_u10_n19915 ), .A2(_u10_n19916 ), .A3(_u10_n19917 ), .A4(_u10_n19918 ), .ZN(_u10_n19909 ) );
NAND2_X1 _u10_U8546  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n19911 ) );
NAND2_X1 _u10_U8545  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n19912 ) );
NAND2_X1 _u10_U8544  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n19913 ) );
NAND2_X1 _u10_U8543  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n19914 ) );
NAND4_X1 _u10_U8542  ( .A1(_u10_n19911 ), .A2(_u10_n19912 ), .A3(_u10_n19913 ), .A4(_u10_n19914 ), .ZN(_u10_n19910 ) );
NOR4_X1 _u10_U8541  ( .A1(_u10_n19907 ), .A2(_u10_n19908 ), .A3(_u10_n19909 ), .A4(_u10_n19910 ), .ZN(_u10_n19906 ) );
NAND2_X1 _u10_U8540  ( .A1(_u10_n19905 ), .A2(_u10_n19906 ), .ZN(am0[18]) );
NAND2_X1 _u10_U8539  ( .A1(1'b1), .A2(_u10_n12430 ), .ZN(_u10_n19901 ) );
NAND2_X1 _u10_U8538  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n19902 ) );
NAND2_X1 _u10_U8537  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n19903 ) );
NAND2_X1 _u10_U8536  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n19904 ) );
NAND4_X1 _u10_U8535  ( .A1(_u10_n19901 ), .A2(_u10_n19902 ), .A3(_u10_n19903 ), .A4(_u10_n19904 ), .ZN(_u10_n19886 ) );
NAND2_X1 _u10_U8534  ( .A1(1'b1), .A2(_u10_n12422 ), .ZN(_u10_n19897 ) );
NAND2_X1 _u10_U8533  ( .A1(1'b1), .A2(_u10_n12421 ), .ZN(_u10_n19898 ) );
NAND2_X1 _u10_U8532  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n19899 ) );
NAND2_X1 _u10_U8531  ( .A1(1'b1), .A2(_u10_n12419 ), .ZN(_u10_n19900 ) );
NAND4_X1 _u10_U8530  ( .A1(_u10_n19897 ), .A2(_u10_n19898 ), .A3(_u10_n19899 ), .A4(_u10_n19900 ), .ZN(_u10_n19887 ) );
NAND2_X1 _u10_U8529  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n19893 ) );
NAND2_X1 _u10_U8528  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n19894 ) );
NAND2_X1 _u10_U8527  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n19895 ) );
NAND2_X1 _u10_U8526  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n19896 ) );
NAND4_X1 _u10_U8525  ( .A1(_u10_n19893 ), .A2(_u10_n19894 ), .A3(_u10_n19895 ), .A4(_u10_n19896 ), .ZN(_u10_n19888 ) );
NAND2_X1 _u10_U8524  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n19890 ) );
NAND2_X1 _u10_U8523  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n19891 ) );
NAND2_X1 _u10_U8522  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19892 ) );
NAND3_X1 _u10_U8521  ( .A1(_u10_n19890 ), .A2(_u10_n19891 ), .A3(_u10_n19892 ), .ZN(_u10_n19889 ) );
NOR4_X1 _u10_U8520  ( .A1(_u10_n19886 ), .A2(_u10_n19887 ), .A3(_u10_n19888 ), .A4(_u10_n19889 ), .ZN(_u10_n19864 ) );
NAND2_X1 _u10_U8519  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n19882 ) );
NAND2_X1 _u10_U8518  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n19883 ) );
NAND2_X1 _u10_U8517  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n19884 ) );
NAND2_X1 _u10_U8516  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n19885 ) );
NAND4_X1 _u10_U8515  ( .A1(_u10_n19882 ), .A2(_u10_n19883 ), .A3(_u10_n19884 ), .A4(_u10_n19885 ), .ZN(_u10_n19866 ) );
NAND2_X1 _u10_U8514  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n19878 ) );
NAND2_X1 _u10_U8513  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n19879 ) );
NAND2_X1 _u10_U8512  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n19880 ) );
NAND2_X1 _u10_U8511  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n19881 ) );
NAND4_X1 _u10_U8510  ( .A1(_u10_n19878 ), .A2(_u10_n19879 ), .A3(_u10_n19880 ), .A4(_u10_n19881 ), .ZN(_u10_n19867 ) );
NAND2_X1 _u10_U8509  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n19874 ) );
NAND2_X1 _u10_U8508  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n19875 ) );
NAND2_X1 _u10_U8507  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n19876 ) );
NAND2_X1 _u10_U8506  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n19877 ) );
NAND4_X1 _u10_U8505  ( .A1(_u10_n19874 ), .A2(_u10_n19875 ), .A3(_u10_n19876 ), .A4(_u10_n19877 ), .ZN(_u10_n19868 ) );
NAND2_X1 _u10_U8504  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n19870 ) );
NAND2_X1 _u10_U8503  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n19871 ) );
NAND2_X1 _u10_U8502  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n19872 ) );
NAND2_X1 _u10_U8501  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n19873 ) );
NAND4_X1 _u10_U8500  ( .A1(_u10_n19870 ), .A2(_u10_n19871 ), .A3(_u10_n19872 ), .A4(_u10_n19873 ), .ZN(_u10_n19869 ) );
NOR4_X1 _u10_U8499  ( .A1(_u10_n19866 ), .A2(_u10_n19867 ), .A3(_u10_n19868 ), .A4(_u10_n19869 ), .ZN(_u10_n19865 ) );
NAND2_X1 _u10_U8498  ( .A1(_u10_n19864 ), .A2(_u10_n19865 ), .ZN(am0[19]) );
NAND2_X1 _u10_U8497  ( .A1(1'b0), .A2(_u10_n12352 ), .ZN(_u10_n19860 ) );
NAND2_X1 _u10_U8496  ( .A1(1'b0), .A2(_u10_n12312 ), .ZN(_u10_n19861 ) );
NAND2_X1 _u10_U8495  ( .A1(1'b0), .A2(_u10_n12288 ), .ZN(_u10_n19862 ) );
NAND2_X1 _u10_U8494  ( .A1(1'b0), .A2(_u10_n12264 ), .ZN(_u10_n19863 ) );
NAND4_X1 _u10_U8493  ( .A1(_u10_n19860 ), .A2(_u10_n19861 ), .A3(_u10_n19862 ), .A4(_u10_n19863 ), .ZN(_u10_n19845 ) );
NAND2_X1 _u10_U8492  ( .A1(1'b0), .A2(_u10_n12256 ), .ZN(_u10_n19856 ) );
NAND2_X1 _u10_U8491  ( .A1(1'b0), .A2(_u10_n12232 ), .ZN(_u10_n19857 ) );
NAND2_X1 _u10_U8490  ( .A1(1'b0), .A2(_u10_n12192 ), .ZN(_u10_n19858 ) );
NAND2_X1 _u10_U8489  ( .A1(1'b0), .A2(_u10_n12184 ), .ZN(_u10_n19859 ) );
NAND4_X1 _u10_U8488  ( .A1(_u10_n19856 ), .A2(_u10_n19857 ), .A3(_u10_n19858 ), .A4(_u10_n19859 ), .ZN(_u10_n19846 ) );
NAND2_X1 _u10_U8487  ( .A1(1'b0), .A2(_u10_n12144 ), .ZN(_u10_n19852 ) );
NAND2_X1 _u10_U8486  ( .A1(1'b0), .A2(_u10_n12120 ), .ZN(_u10_n19853 ) );
NAND2_X1 _u10_U8485  ( .A1(1'b0), .A2(_u10_n12096 ), .ZN(_u10_n19854 ) );
NAND2_X1 _u10_U8484  ( .A1(1'b0), .A2(_u10_n12072 ), .ZN(_u10_n19855 ) );
NAND4_X1 _u10_U8483  ( .A1(_u10_n19852 ), .A2(_u10_n19853 ), .A3(_u10_n19854 ), .A4(_u10_n19855 ), .ZN(_u10_n19847 ) );
NAND2_X1 _u10_U8482  ( .A1(1'b0), .A2(_u10_n12048 ), .ZN(_u10_n19849 ) );
NAND2_X1 _u10_U8481  ( .A1(1'b0), .A2(_u10_n12024 ), .ZN(_u10_n19850 ) );
NAND2_X1 _u10_U8480  ( .A1(1'b0), .A2(_u10_n12005 ), .ZN(_u10_n19851 ) );
NAND3_X1 _u10_U8479  ( .A1(_u10_n19849 ), .A2(_u10_n19850 ), .A3(_u10_n19851 ), .ZN(_u10_n19848 ) );
NOR4_X1 _u10_U8478  ( .A1(_u10_n19845 ), .A2(_u10_n19846 ), .A3(_u10_n19847 ), .A4(_u10_n19848 ), .ZN(_u10_n19823 ) );
NAND2_X1 _u10_U8477  ( .A1(1'b0), .A2(_u10_n11988 ), .ZN(_u10_n19841 ) );
NAND2_X1 _u10_U8476  ( .A1(1'b0), .A2(_u10_n11964 ), .ZN(_u10_n19842 ) );
NAND2_X1 _u10_U8475  ( .A1(1'b0), .A2(_u10_n11940 ), .ZN(_u10_n19843 ) );
NAND2_X1 _u10_U8474  ( .A1(1'b0), .A2(_u10_n11916 ), .ZN(_u10_n19844 ) );
NAND4_X1 _u10_U8473  ( .A1(_u10_n19841 ), .A2(_u10_n19842 ), .A3(_u10_n19843 ), .A4(_u10_n19844 ), .ZN(_u10_n19825 ) );
NAND2_X1 _u10_U8472  ( .A1(1'b0), .A2(_u10_n11892 ), .ZN(_u10_n19837 ) );
NAND2_X1 _u10_U8471  ( .A1(1'b0), .A2(_u10_n11868 ), .ZN(_u10_n19838 ) );
NAND2_X1 _u10_U8470  ( .A1(1'b0), .A2(_u10_n11844 ), .ZN(_u10_n19839 ) );
NAND2_X1 _u10_U8469  ( .A1(1'b0), .A2(_u10_n11820 ), .ZN(_u10_n19840 ) );
NAND4_X1 _u10_U8468  ( .A1(_u10_n19837 ), .A2(_u10_n19838 ), .A3(_u10_n19839 ), .A4(_u10_n19840 ), .ZN(_u10_n19826 ) );
NAND2_X1 _u10_U8467  ( .A1(1'b0), .A2(_u10_n11796 ), .ZN(_u10_n19833 ) );
NAND2_X1 _u10_U8466  ( .A1(1'b0), .A2(_u10_n11772 ), .ZN(_u10_n19834 ) );
NAND2_X1 _u10_U8465  ( .A1(1'b0), .A2(_u10_n11748 ), .ZN(_u10_n19835 ) );
NAND2_X1 _u10_U8464  ( .A1(1'b0), .A2(_u10_n11724 ), .ZN(_u10_n19836 ) );
NAND4_X1 _u10_U8463  ( .A1(_u10_n19833 ), .A2(_u10_n19834 ), .A3(_u10_n19835 ), .A4(_u10_n19836 ), .ZN(_u10_n19827 ) );
NAND2_X1 _u10_U8462  ( .A1(1'b0), .A2(_u10_n11700 ), .ZN(_u10_n19829 ) );
NAND2_X1 _u10_U8461  ( .A1(1'b0), .A2(_u10_n11676 ), .ZN(_u10_n19830 ) );
NAND2_X1 _u10_U8460  ( .A1(1'b0), .A2(_u10_n11652 ), .ZN(_u10_n19831 ) );
NAND2_X1 _u10_U8459  ( .A1(1'b0), .A2(_u10_n11628 ), .ZN(_u10_n19832 ) );
NAND4_X1 _u10_U8458  ( .A1(_u10_n19829 ), .A2(_u10_n19830 ), .A3(_u10_n19831 ), .A4(_u10_n19832 ), .ZN(_u10_n19828 ) );
NOR4_X1 _u10_U8457  ( .A1(_u10_n19825 ), .A2(_u10_n19826 ), .A3(_u10_n19827 ), .A4(_u10_n19828 ), .ZN(_u10_n19824 ) );
NAND2_X1 _u10_U8456  ( .A1(_u10_n19823 ), .A2(_u10_n19824 ), .ZN(am0[1]) );
NAND2_X1 _u10_U8455  ( .A1(1'b1), .A2(_u10_n12430 ), .ZN(_u10_n19819 ) );
NAND2_X1 _u10_U8454  ( .A1(1'b1), .A2(_u10_n12312 ), .ZN(_u10_n19820 ) );
NAND2_X1 _u10_U8453  ( .A1(1'b1), .A2(_u10_n12288 ), .ZN(_u10_n19821 ) );
NAND2_X1 _u10_U8452  ( .A1(1'b1), .A2(_u10_n12264 ), .ZN(_u10_n19822 ) );
NAND4_X1 _u10_U8451  ( .A1(_u10_n19819 ), .A2(_u10_n19820 ), .A3(_u10_n19821 ), .A4(_u10_n19822 ), .ZN(_u10_n19804 ) );
NAND2_X1 _u10_U8450  ( .A1(1'b1), .A2(_u10_n12422 ), .ZN(_u10_n19815 ) );
NAND2_X1 _u10_U8449  ( .A1(1'b1), .A2(_u10_n12421 ), .ZN(_u10_n19816 ) );
NAND2_X1 _u10_U8448  ( .A1(1'b1), .A2(_u10_n12192 ), .ZN(_u10_n19817 ) );
NAND2_X1 _u10_U8447  ( .A1(1'b1), .A2(_u10_n12419 ), .ZN(_u10_n19818 ) );
NAND4_X1 _u10_U8446  ( .A1(_u10_n19815 ), .A2(_u10_n19816 ), .A3(_u10_n19817 ), .A4(_u10_n19818 ), .ZN(_u10_n19805 ) );
NAND2_X1 _u10_U8445  ( .A1(1'b1), .A2(_u10_n12144 ), .ZN(_u10_n19811 ) );
NAND2_X1 _u10_U8444  ( .A1(1'b1), .A2(_u10_n12120 ), .ZN(_u10_n19812 ) );
NAND2_X1 _u10_U8443  ( .A1(1'b1), .A2(_u10_n12096 ), .ZN(_u10_n19813 ) );
NAND2_X1 _u10_U8442  ( .A1(1'b1), .A2(_u10_n12072 ), .ZN(_u10_n19814 ) );
NAND4_X1 _u10_U8441  ( .A1(_u10_n19811 ), .A2(_u10_n19812 ), .A3(_u10_n19813 ), .A4(_u10_n19814 ), .ZN(_u10_n19806 ) );
NAND2_X1 _u10_U8440  ( .A1(1'b1), .A2(_u10_n12048 ), .ZN(_u10_n19808 ) );
NAND2_X1 _u10_U8439  ( .A1(1'b1), .A2(_u10_n12024 ), .ZN(_u10_n19809 ) );
NAND2_X1 _u10_U8438  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19810 ) );
NAND3_X1 _u10_U8437  ( .A1(_u10_n19808 ), .A2(_u10_n19809 ), .A3(_u10_n19810 ), .ZN(_u10_n19807 ) );
NOR4_X1 _u10_U8436  ( .A1(_u10_n19804 ), .A2(_u10_n19805 ), .A3(_u10_n19806 ), .A4(_u10_n19807 ), .ZN(_u10_n19782 ) );
NAND2_X1 _u10_U8435  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n19800 ) );
NAND2_X1 _u10_U8434  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n19801 ) );
NAND2_X1 _u10_U8433  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n19802 ) );
NAND2_X1 _u10_U8432  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n19803 ) );
NAND4_X1 _u10_U8431  ( .A1(_u10_n19800 ), .A2(_u10_n19801 ), .A3(_u10_n19802 ), .A4(_u10_n19803 ), .ZN(_u10_n19784 ) );
NAND2_X1 _u10_U8430  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n19796 ) );
NAND2_X1 _u10_U8429  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n19797 ) );
NAND2_X1 _u10_U8428  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n19798 ) );
NAND2_X1 _u10_U8427  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n19799 ) );
NAND4_X1 _u10_U8426  ( .A1(_u10_n19796 ), .A2(_u10_n19797 ), .A3(_u10_n19798 ), .A4(_u10_n19799 ), .ZN(_u10_n19785 ) );
NAND2_X1 _u10_U8425  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n19792 ) );
NAND2_X1 _u10_U8424  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n19793 ) );
NAND2_X1 _u10_U8423  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n19794 ) );
NAND2_X1 _u10_U8422  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n19795 ) );
NAND4_X1 _u10_U8421  ( .A1(_u10_n19792 ), .A2(_u10_n19793 ), .A3(_u10_n19794 ), .A4(_u10_n19795 ), .ZN(_u10_n19786 ) );
NAND2_X1 _u10_U8420  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n19788 ) );
NAND2_X1 _u10_U8419  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n19789 ) );
NAND2_X1 _u10_U8418  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n19790 ) );
NAND2_X1 _u10_U8417  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n19791 ) );
NAND4_X1 _u10_U8416  ( .A1(_u10_n19788 ), .A2(_u10_n19789 ), .A3(_u10_n19790 ), .A4(_u10_n19791 ), .ZN(_u10_n19787 ) );
NOR4_X1 _u10_U8415  ( .A1(_u10_n19784 ), .A2(_u10_n19785 ), .A3(_u10_n19786 ), .A4(_u10_n19787 ), .ZN(_u10_n19783 ) );
NAND2_X1 _u10_U8414  ( .A1(_u10_n19782 ), .A2(_u10_n19783 ), .ZN(am0[20]) );
NAND2_X1 _u10_U8413  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19778 ) );
NAND2_X1 _u10_U8412  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19779 ) );
NAND2_X1 _u10_U8411  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19780 ) );
NAND2_X1 _u10_U8410  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19781 ) );
NAND4_X1 _u10_U8409  ( .A1(_u10_n19778 ), .A2(_u10_n19779 ), .A3(_u10_n19780 ), .A4(_u10_n19781 ), .ZN(_u10_n19763 ) );
NAND2_X1 _u10_U8408  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19774 ) );
NAND2_X1 _u10_U8407  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19775 ) );
NAND2_X1 _u10_U8406  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19776 ) );
NAND2_X1 _u10_U8405  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19777 ) );
NAND4_X1 _u10_U8404  ( .A1(_u10_n19774 ), .A2(_u10_n19775 ), .A3(_u10_n19776 ), .A4(_u10_n19777 ), .ZN(_u10_n19764 ) );
NAND2_X1 _u10_U8403  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19770 ) );
NAND2_X1 _u10_U8402  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19771 ) );
NAND2_X1 _u10_U8401  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19772 ) );
NAND2_X1 _u10_U8400  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19773 ) );
NAND4_X1 _u10_U8399  ( .A1(_u10_n19770 ), .A2(_u10_n19771 ), .A3(_u10_n19772 ), .A4(_u10_n19773 ), .ZN(_u10_n19765 ) );
NAND2_X1 _u10_U8398  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19767 ) );
NAND2_X1 _u10_U8397  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19768 ) );
NAND2_X1 _u10_U8396  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19769 ) );
NAND3_X1 _u10_U8395  ( .A1(_u10_n19767 ), .A2(_u10_n19768 ), .A3(_u10_n19769 ), .ZN(_u10_n19766 ) );
NOR4_X1 _u10_U8394  ( .A1(_u10_n19763 ), .A2(_u10_n19764 ), .A3(_u10_n19765 ), .A4(_u10_n19766 ), .ZN(_u10_n19741 ) );
NAND2_X1 _u10_U8393  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n19759 ) );
NAND2_X1 _u10_U8392  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n19760 ) );
NAND2_X1 _u10_U8391  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n19761 ) );
NAND2_X1 _u10_U8390  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n19762 ) );
NAND4_X1 _u10_U8389  ( .A1(_u10_n19759 ), .A2(_u10_n19760 ), .A3(_u10_n19761 ), .A4(_u10_n19762 ), .ZN(_u10_n19743 ) );
NAND2_X1 _u10_U8388  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n19755 ) );
NAND2_X1 _u10_U8387  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n19756 ) );
NAND2_X1 _u10_U8386  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n19757 ) );
NAND2_X1 _u10_U8385  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n19758 ) );
NAND4_X1 _u10_U8384  ( .A1(_u10_n19755 ), .A2(_u10_n19756 ), .A3(_u10_n19757 ), .A4(_u10_n19758 ), .ZN(_u10_n19744 ) );
NAND2_X1 _u10_U8383  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n19751 ) );
NAND2_X1 _u10_U8382  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n19752 ) );
NAND2_X1 _u10_U8381  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n19753 ) );
NAND2_X1 _u10_U8380  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n19754 ) );
NAND4_X1 _u10_U8379  ( .A1(_u10_n19751 ), .A2(_u10_n19752 ), .A3(_u10_n19753 ), .A4(_u10_n19754 ), .ZN(_u10_n19745 ) );
NAND2_X1 _u10_U8378  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n19747 ) );
NAND2_X1 _u10_U8377  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n19748 ) );
NAND2_X1 _u10_U8376  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n19749 ) );
NAND2_X1 _u10_U8375  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n19750 ) );
NAND4_X1 _u10_U8374  ( .A1(_u10_n19747 ), .A2(_u10_n19748 ), .A3(_u10_n19749 ), .A4(_u10_n19750 ), .ZN(_u10_n19746 ) );
NOR4_X1 _u10_U8373  ( .A1(_u10_n19743 ), .A2(_u10_n19744 ), .A3(_u10_n19745 ), .A4(_u10_n19746 ), .ZN(_u10_n19742 ) );
NAND2_X1 _u10_U8372  ( .A1(_u10_n19741 ), .A2(_u10_n19742 ), .ZN(am0[21]) );
NAND2_X1 _u10_U8371  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19737 ) );
NAND2_X1 _u10_U8370  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19738 ) );
NAND2_X1 _u10_U8369  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19739 ) );
NAND2_X1 _u10_U8368  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19740 ) );
NAND4_X1 _u10_U8367  ( .A1(_u10_n19737 ), .A2(_u10_n19738 ), .A3(_u10_n19739 ), .A4(_u10_n19740 ), .ZN(_u10_n19722 ) );
NAND2_X1 _u10_U8366  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19733 ) );
NAND2_X1 _u10_U8365  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19734 ) );
NAND2_X1 _u10_U8364  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19735 ) );
NAND2_X1 _u10_U8363  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19736 ) );
NAND4_X1 _u10_U8362  ( .A1(_u10_n19733 ), .A2(_u10_n19734 ), .A3(_u10_n19735 ), .A4(_u10_n19736 ), .ZN(_u10_n19723 ) );
NAND2_X1 _u10_U8361  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19729 ) );
NAND2_X1 _u10_U8360  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19730 ) );
NAND2_X1 _u10_U8359  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19731 ) );
NAND2_X1 _u10_U8358  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19732 ) );
NAND4_X1 _u10_U8357  ( .A1(_u10_n19729 ), .A2(_u10_n19730 ), .A3(_u10_n19731 ), .A4(_u10_n19732 ), .ZN(_u10_n19724 ) );
NAND2_X1 _u10_U8356  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19726 ) );
NAND2_X1 _u10_U8355  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19727 ) );
NAND2_X1 _u10_U8354  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19728 ) );
NAND3_X1 _u10_U8353  ( .A1(_u10_n19726 ), .A2(_u10_n19727 ), .A3(_u10_n19728 ), .ZN(_u10_n19725 ) );
NOR4_X1 _u10_U8352  ( .A1(_u10_n19722 ), .A2(_u10_n19723 ), .A3(_u10_n19724 ), .A4(_u10_n19725 ), .ZN(_u10_n19700 ) );
NAND2_X1 _u10_U8351  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n19718 ) );
NAND2_X1 _u10_U8350  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n19719 ) );
NAND2_X1 _u10_U8349  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n19720 ) );
NAND2_X1 _u10_U8348  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n19721 ) );
NAND4_X1 _u10_U8347  ( .A1(_u10_n19718 ), .A2(_u10_n19719 ), .A3(_u10_n19720 ), .A4(_u10_n19721 ), .ZN(_u10_n19702 ) );
NAND2_X1 _u10_U8346  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n19714 ) );
NAND2_X1 _u10_U8345  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n19715 ) );
NAND2_X1 _u10_U8344  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n19716 ) );
NAND2_X1 _u10_U8343  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n19717 ) );
NAND4_X1 _u10_U8342  ( .A1(_u10_n19714 ), .A2(_u10_n19715 ), .A3(_u10_n19716 ), .A4(_u10_n19717 ), .ZN(_u10_n19703 ) );
NAND2_X1 _u10_U8341  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n19710 ) );
NAND2_X1 _u10_U8340  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n19711 ) );
NAND2_X1 _u10_U8339  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n19712 ) );
NAND2_X1 _u10_U8338  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n19713 ) );
NAND4_X1 _u10_U8337  ( .A1(_u10_n19710 ), .A2(_u10_n19711 ), .A3(_u10_n19712 ), .A4(_u10_n19713 ), .ZN(_u10_n19704 ) );
NAND2_X1 _u10_U8336  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n19706 ) );
NAND2_X1 _u10_U8335  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n19707 ) );
NAND2_X1 _u10_U8334  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n19708 ) );
NAND2_X1 _u10_U8333  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n19709 ) );
NAND4_X1 _u10_U8332  ( .A1(_u10_n19706 ), .A2(_u10_n19707 ), .A3(_u10_n19708 ), .A4(_u10_n19709 ), .ZN(_u10_n19705 ) );
NOR4_X1 _u10_U8331  ( .A1(_u10_n19702 ), .A2(_u10_n19703 ), .A3(_u10_n19704 ), .A4(_u10_n19705 ), .ZN(_u10_n19701 ) );
NAND2_X1 _u10_U8330  ( .A1(_u10_n19700 ), .A2(_u10_n19701 ), .ZN(am0[22]) );
NAND2_X1 _u10_U8329  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19696 ) );
NAND2_X1 _u10_U8328  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19697 ) );
NAND2_X1 _u10_U8327  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19698 ) );
NAND2_X1 _u10_U8326  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19699 ) );
NAND4_X1 _u10_U8325  ( .A1(_u10_n19696 ), .A2(_u10_n19697 ), .A3(_u10_n19698 ), .A4(_u10_n19699 ), .ZN(_u10_n19681 ) );
NAND2_X1 _u10_U8324  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19692 ) );
NAND2_X1 _u10_U8323  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19693 ) );
NAND2_X1 _u10_U8322  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19694 ) );
NAND2_X1 _u10_U8321  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19695 ) );
NAND4_X1 _u10_U8320  ( .A1(_u10_n19692 ), .A2(_u10_n19693 ), .A3(_u10_n19694 ), .A4(_u10_n19695 ), .ZN(_u10_n19682 ) );
NAND2_X1 _u10_U8319  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19688 ) );
NAND2_X1 _u10_U8318  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19689 ) );
NAND2_X1 _u10_U8317  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19690 ) );
NAND2_X1 _u10_U8316  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19691 ) );
NAND4_X1 _u10_U8315  ( .A1(_u10_n19688 ), .A2(_u10_n19689 ), .A3(_u10_n19690 ), .A4(_u10_n19691 ), .ZN(_u10_n19683 ) );
NAND2_X1 _u10_U8314  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19685 ) );
NAND2_X1 _u10_U8313  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19686 ) );
NAND2_X1 _u10_U8312  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19687 ) );
NAND3_X1 _u10_U8311  ( .A1(_u10_n19685 ), .A2(_u10_n19686 ), .A3(_u10_n19687 ), .ZN(_u10_n19684 ) );
NOR4_X1 _u10_U8310  ( .A1(_u10_n19681 ), .A2(_u10_n19682 ), .A3(_u10_n19683 ), .A4(_u10_n19684 ), .ZN(_u10_n19659 ) );
NAND2_X1 _u10_U8309  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n19677 ) );
NAND2_X1 _u10_U8308  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n19678 ) );
NAND2_X1 _u10_U8307  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n19679 ) );
NAND2_X1 _u10_U8306  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n19680 ) );
NAND4_X1 _u10_U8305  ( .A1(_u10_n19677 ), .A2(_u10_n19678 ), .A3(_u10_n19679 ), .A4(_u10_n19680 ), .ZN(_u10_n19661 ) );
NAND2_X1 _u10_U8304  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n19673 ) );
NAND2_X1 _u10_U8303  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n19674 ) );
NAND2_X1 _u10_U8302  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n19675 ) );
NAND2_X1 _u10_U8301  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n19676 ) );
NAND4_X1 _u10_U8300  ( .A1(_u10_n19673 ), .A2(_u10_n19674 ), .A3(_u10_n19675 ), .A4(_u10_n19676 ), .ZN(_u10_n19662 ) );
NAND2_X1 _u10_U8299  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n19669 ) );
NAND2_X1 _u10_U8298  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n19670 ) );
NAND2_X1 _u10_U8297  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n19671 ) );
NAND2_X1 _u10_U8296  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n19672 ) );
NAND4_X1 _u10_U8295  ( .A1(_u10_n19669 ), .A2(_u10_n19670 ), .A3(_u10_n19671 ), .A4(_u10_n19672 ), .ZN(_u10_n19663 ) );
NAND2_X1 _u10_U8294  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n19665 ) );
NAND2_X1 _u10_U8293  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n19666 ) );
NAND2_X1 _u10_U8292  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n19667 ) );
NAND2_X1 _u10_U8291  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n19668 ) );
NAND4_X1 _u10_U8290  ( .A1(_u10_n19665 ), .A2(_u10_n19666 ), .A3(_u10_n19667 ), .A4(_u10_n19668 ), .ZN(_u10_n19664 ) );
NOR4_X1 _u10_U8289  ( .A1(_u10_n19661 ), .A2(_u10_n19662 ), .A3(_u10_n19663 ), .A4(_u10_n19664 ), .ZN(_u10_n19660 ) );
NAND2_X1 _u10_U8288  ( .A1(_u10_n19659 ), .A2(_u10_n19660 ), .ZN(am0[23]) );
NAND2_X1 _u10_U8287  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19655 ) );
NAND2_X1 _u10_U8286  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19656 ) );
NAND2_X1 _u10_U8285  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19657 ) );
NAND2_X1 _u10_U8284  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19658 ) );
NAND4_X1 _u10_U8283  ( .A1(_u10_n19655 ), .A2(_u10_n19656 ), .A3(_u10_n19657 ), .A4(_u10_n19658 ), .ZN(_u10_n19640 ) );
NAND2_X1 _u10_U8282  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19651 ) );
NAND2_X1 _u10_U8281  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19652 ) );
NAND2_X1 _u10_U8280  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19653 ) );
NAND2_X1 _u10_U8279  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19654 ) );
NAND4_X1 _u10_U8278  ( .A1(_u10_n19651 ), .A2(_u10_n19652 ), .A3(_u10_n19653 ), .A4(_u10_n19654 ), .ZN(_u10_n19641 ) );
NAND2_X1 _u10_U8277  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19647 ) );
NAND2_X1 _u10_U8276  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19648 ) );
NAND2_X1 _u10_U8275  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19649 ) );
NAND2_X1 _u10_U8274  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19650 ) );
NAND4_X1 _u10_U8273  ( .A1(_u10_n19647 ), .A2(_u10_n19648 ), .A3(_u10_n19649 ), .A4(_u10_n19650 ), .ZN(_u10_n19642 ) );
NAND2_X1 _u10_U8272  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19644 ) );
NAND2_X1 _u10_U8271  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19645 ) );
NAND2_X1 _u10_U8270  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19646 ) );
NAND3_X1 _u10_U8269  ( .A1(_u10_n19644 ), .A2(_u10_n19645 ), .A3(_u10_n19646 ), .ZN(_u10_n19643 ) );
NOR4_X1 _u10_U8268  ( .A1(_u10_n19640 ), .A2(_u10_n19641 ), .A3(_u10_n19642 ), .A4(_u10_n19643 ), .ZN(_u10_n19618 ) );
NAND2_X1 _u10_U8267  ( .A1(1'b1), .A2(_u10_n11988 ), .ZN(_u10_n19636 ) );
NAND2_X1 _u10_U8266  ( .A1(1'b1), .A2(_u10_n11964 ), .ZN(_u10_n19637 ) );
NAND2_X1 _u10_U8265  ( .A1(1'b1), .A2(_u10_n11940 ), .ZN(_u10_n19638 ) );
NAND2_X1 _u10_U8264  ( .A1(1'b1), .A2(_u10_n11916 ), .ZN(_u10_n19639 ) );
NAND4_X1 _u10_U8263  ( .A1(_u10_n19636 ), .A2(_u10_n19637 ), .A3(_u10_n19638 ), .A4(_u10_n19639 ), .ZN(_u10_n19620 ) );
NAND2_X1 _u10_U8262  ( .A1(1'b1), .A2(_u10_n11892 ), .ZN(_u10_n19632 ) );
NAND2_X1 _u10_U8261  ( .A1(1'b1), .A2(_u10_n11868 ), .ZN(_u10_n19633 ) );
NAND2_X1 _u10_U8260  ( .A1(1'b1), .A2(_u10_n11844 ), .ZN(_u10_n19634 ) );
NAND2_X1 _u10_U8259  ( .A1(1'b1), .A2(_u10_n11820 ), .ZN(_u10_n19635 ) );
NAND4_X1 _u10_U8258  ( .A1(_u10_n19632 ), .A2(_u10_n19633 ), .A3(_u10_n19634 ), .A4(_u10_n19635 ), .ZN(_u10_n19621 ) );
NAND2_X1 _u10_U8257  ( .A1(1'b1), .A2(_u10_n11796 ), .ZN(_u10_n19628 ) );
NAND2_X1 _u10_U8256  ( .A1(1'b1), .A2(_u10_n11772 ), .ZN(_u10_n19629 ) );
NAND2_X1 _u10_U8255  ( .A1(1'b1), .A2(_u10_n11748 ), .ZN(_u10_n19630 ) );
NAND2_X1 _u10_U8254  ( .A1(1'b1), .A2(_u10_n11724 ), .ZN(_u10_n19631 ) );
NAND4_X1 _u10_U8253  ( .A1(_u10_n19628 ), .A2(_u10_n19629 ), .A3(_u10_n19630 ), .A4(_u10_n19631 ), .ZN(_u10_n19622 ) );
NAND2_X1 _u10_U8252  ( .A1(1'b1), .A2(_u10_n11700 ), .ZN(_u10_n19624 ) );
NAND2_X1 _u10_U8251  ( .A1(1'b1), .A2(_u10_n11676 ), .ZN(_u10_n19625 ) );
NAND2_X1 _u10_U8250  ( .A1(1'b1), .A2(_u10_n11652 ), .ZN(_u10_n19626 ) );
NAND2_X1 _u10_U8249  ( .A1(1'b1), .A2(_u10_n11628 ), .ZN(_u10_n19627 ) );
NAND4_X1 _u10_U8248  ( .A1(_u10_n19624 ), .A2(_u10_n19625 ), .A3(_u10_n19626 ), .A4(_u10_n19627 ), .ZN(_u10_n19623 ) );
NOR4_X1 _u10_U8247  ( .A1(_u10_n19620 ), .A2(_u10_n19621 ), .A3(_u10_n19622 ), .A4(_u10_n19623 ), .ZN(_u10_n19619 ) );
NAND2_X1 _u10_U8246  ( .A1(_u10_n19618 ), .A2(_u10_n19619 ), .ZN(am0[24]) );
NAND2_X1 _u10_U8245  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19614 ) );
NAND2_X1 _u10_U8244  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19615 ) );
NAND2_X1 _u10_U8243  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19616 ) );
NAND2_X1 _u10_U8242  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19617 ) );
NAND4_X1 _u10_U8241  ( .A1(_u10_n19614 ), .A2(_u10_n19615 ), .A3(_u10_n19616 ), .A4(_u10_n19617 ), .ZN(_u10_n19599 ) );
NAND2_X1 _u10_U8240  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19610 ) );
NAND2_X1 _u10_U8239  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19611 ) );
NAND2_X1 _u10_U8238  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19612 ) );
NAND2_X1 _u10_U8237  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19613 ) );
NAND4_X1 _u10_U8236  ( .A1(_u10_n19610 ), .A2(_u10_n19611 ), .A3(_u10_n19612 ), .A4(_u10_n19613 ), .ZN(_u10_n19600 ) );
NAND2_X1 _u10_U8235  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19606 ) );
NAND2_X1 _u10_U8234  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19607 ) );
NAND2_X1 _u10_U8233  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19608 ) );
NAND2_X1 _u10_U8232  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19609 ) );
NAND4_X1 _u10_U8231  ( .A1(_u10_n19606 ), .A2(_u10_n19607 ), .A3(_u10_n19608 ), .A4(_u10_n19609 ), .ZN(_u10_n19601 ) );
NAND2_X1 _u10_U8230  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19603 ) );
NAND2_X1 _u10_U8229  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19604 ) );
NAND2_X1 _u10_U8228  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19605 ) );
NAND3_X1 _u10_U8227  ( .A1(_u10_n19603 ), .A2(_u10_n19604 ), .A3(_u10_n19605 ), .ZN(_u10_n19602 ) );
NOR4_X1 _u10_U8226  ( .A1(_u10_n19599 ), .A2(_u10_n19600 ), .A3(_u10_n19601 ), .A4(_u10_n19602 ), .ZN(_u10_n19577 ) );
NAND2_X1 _u10_U8225  ( .A1(1'b1), .A2(_u10_n11989 ), .ZN(_u10_n19595 ) );
NAND2_X1 _u10_U8224  ( .A1(1'b1), .A2(_u10_n11965 ), .ZN(_u10_n19596 ) );
NAND2_X1 _u10_U8223  ( .A1(1'b1), .A2(_u10_n11941 ), .ZN(_u10_n19597 ) );
NAND2_X1 _u10_U8222  ( .A1(1'b1), .A2(_u10_n11917 ), .ZN(_u10_n19598 ) );
NAND4_X1 _u10_U8221  ( .A1(_u10_n19595 ), .A2(_u10_n19596 ), .A3(_u10_n19597 ), .A4(_u10_n19598 ), .ZN(_u10_n19579 ) );
NAND2_X1 _u10_U8220  ( .A1(1'b1), .A2(_u10_n11893 ), .ZN(_u10_n19591 ) );
NAND2_X1 _u10_U8219  ( .A1(1'b1), .A2(_u10_n11869 ), .ZN(_u10_n19592 ) );
NAND2_X1 _u10_U8218  ( .A1(1'b1), .A2(_u10_n11845 ), .ZN(_u10_n19593 ) );
NAND2_X1 _u10_U8217  ( .A1(1'b1), .A2(_u10_n11821 ), .ZN(_u10_n19594 ) );
NAND4_X1 _u10_U8216  ( .A1(_u10_n19591 ), .A2(_u10_n19592 ), .A3(_u10_n19593 ), .A4(_u10_n19594 ), .ZN(_u10_n19580 ) );
NAND2_X1 _u10_U8215  ( .A1(1'b1), .A2(_u10_n11797 ), .ZN(_u10_n19587 ) );
NAND2_X1 _u10_U8214  ( .A1(1'b1), .A2(_u10_n11773 ), .ZN(_u10_n19588 ) );
NAND2_X1 _u10_U8213  ( .A1(1'b1), .A2(_u10_n11749 ), .ZN(_u10_n19589 ) );
NAND2_X1 _u10_U8212  ( .A1(1'b1), .A2(_u10_n11725 ), .ZN(_u10_n19590 ) );
NAND4_X1 _u10_U8211  ( .A1(_u10_n19587 ), .A2(_u10_n19588 ), .A3(_u10_n19589 ), .A4(_u10_n19590 ), .ZN(_u10_n19581 ) );
NAND2_X1 _u10_U8210  ( .A1(1'b1), .A2(_u10_n11701 ), .ZN(_u10_n19583 ) );
NAND2_X1 _u10_U8209  ( .A1(1'b1), .A2(_u10_n11677 ), .ZN(_u10_n19584 ) );
NAND2_X1 _u10_U8208  ( .A1(1'b1), .A2(_u10_n11653 ), .ZN(_u10_n19585 ) );
NAND2_X1 _u10_U8207  ( .A1(1'b1), .A2(_u10_n11629 ), .ZN(_u10_n19586 ) );
NAND4_X1 _u10_U8206  ( .A1(_u10_n19583 ), .A2(_u10_n19584 ), .A3(_u10_n19585 ), .A4(_u10_n19586 ), .ZN(_u10_n19582 ) );
NOR4_X1 _u10_U8205  ( .A1(_u10_n19579 ), .A2(_u10_n19580 ), .A3(_u10_n19581 ), .A4(_u10_n19582 ), .ZN(_u10_n19578 ) );
NAND2_X1 _u10_U8204  ( .A1(_u10_n19577 ), .A2(_u10_n19578 ), .ZN(am0[25]) );
NAND2_X1 _u10_U8203  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19573 ) );
NAND2_X1 _u10_U8202  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19574 ) );
NAND2_X1 _u10_U8201  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19575 ) );
NAND2_X1 _u10_U8200  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19576 ) );
NAND4_X1 _u10_U8199  ( .A1(_u10_n19573 ), .A2(_u10_n19574 ), .A3(_u10_n19575 ), .A4(_u10_n19576 ), .ZN(_u10_n19558 ) );
NAND2_X1 _u10_U8198  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19569 ) );
NAND2_X1 _u10_U8197  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19570 ) );
NAND2_X1 _u10_U8196  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19571 ) );
NAND2_X1 _u10_U8195  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19572 ) );
NAND4_X1 _u10_U8194  ( .A1(_u10_n19569 ), .A2(_u10_n19570 ), .A3(_u10_n19571 ), .A4(_u10_n19572 ), .ZN(_u10_n19559 ) );
NAND2_X1 _u10_U8193  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19565 ) );
NAND2_X1 _u10_U8192  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19566 ) );
NAND2_X1 _u10_U8191  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19567 ) );
NAND2_X1 _u10_U8190  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19568 ) );
NAND4_X1 _u10_U8189  ( .A1(_u10_n19565 ), .A2(_u10_n19566 ), .A3(_u10_n19567 ), .A4(_u10_n19568 ), .ZN(_u10_n19560 ) );
NAND2_X1 _u10_U8188  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19562 ) );
NAND2_X1 _u10_U8187  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19563 ) );
NAND2_X1 _u10_U8186  ( .A1(1'b1), .A2(_u10_n12005 ), .ZN(_u10_n19564 ) );
NAND3_X1 _u10_U8185  ( .A1(_u10_n19562 ), .A2(_u10_n19563 ), .A3(_u10_n19564 ), .ZN(_u10_n19561 ) );
NOR4_X1 _u10_U8184  ( .A1(_u10_n19558 ), .A2(_u10_n19559 ), .A3(_u10_n19560 ), .A4(_u10_n19561 ), .ZN(_u10_n19536 ) );
NAND2_X1 _u10_U8183  ( .A1(1'b1), .A2(_u10_n11989 ), .ZN(_u10_n19554 ) );
NAND2_X1 _u10_U8182  ( .A1(1'b1), .A2(_u10_n11965 ), .ZN(_u10_n19555 ) );
NAND2_X1 _u10_U8181  ( .A1(1'b1), .A2(_u10_n11941 ), .ZN(_u10_n19556 ) );
NAND2_X1 _u10_U8180  ( .A1(1'b1), .A2(_u10_n11917 ), .ZN(_u10_n19557 ) );
NAND4_X1 _u10_U8179  ( .A1(_u10_n19554 ), .A2(_u10_n19555 ), .A3(_u10_n19556 ), .A4(_u10_n19557 ), .ZN(_u10_n19538 ) );
NAND2_X1 _u10_U8178  ( .A1(1'b1), .A2(_u10_n11893 ), .ZN(_u10_n19550 ) );
NAND2_X1 _u10_U8177  ( .A1(1'b1), .A2(_u10_n11869 ), .ZN(_u10_n19551 ) );
NAND2_X1 _u10_U8176  ( .A1(1'b1), .A2(_u10_n11845 ), .ZN(_u10_n19552 ) );
NAND2_X1 _u10_U8175  ( .A1(1'b1), .A2(_u10_n11821 ), .ZN(_u10_n19553 ) );
NAND4_X1 _u10_U8174  ( .A1(_u10_n19550 ), .A2(_u10_n19551 ), .A3(_u10_n19552 ), .A4(_u10_n19553 ), .ZN(_u10_n19539 ) );
NAND2_X1 _u10_U8173  ( .A1(1'b1), .A2(_u10_n11797 ), .ZN(_u10_n19546 ) );
NAND2_X1 _u10_U8172  ( .A1(1'b1), .A2(_u10_n11773 ), .ZN(_u10_n19547 ) );
NAND2_X1 _u10_U8171  ( .A1(1'b1), .A2(_u10_n11749 ), .ZN(_u10_n19548 ) );
NAND2_X1 _u10_U8170  ( .A1(1'b1), .A2(_u10_n11725 ), .ZN(_u10_n19549 ) );
NAND4_X1 _u10_U8169  ( .A1(_u10_n19546 ), .A2(_u10_n19547 ), .A3(_u10_n19548 ), .A4(_u10_n19549 ), .ZN(_u10_n19540 ) );
NAND2_X1 _u10_U8168  ( .A1(1'b1), .A2(_u10_n11701 ), .ZN(_u10_n19542 ) );
NAND2_X1 _u10_U8167  ( .A1(1'b1), .A2(_u10_n11677 ), .ZN(_u10_n19543 ) );
NAND2_X1 _u10_U8166  ( .A1(1'b1), .A2(_u10_n11653 ), .ZN(_u10_n19544 ) );
NAND2_X1 _u10_U8165  ( .A1(1'b1), .A2(_u10_n11629 ), .ZN(_u10_n19545 ) );
NAND4_X1 _u10_U8164  ( .A1(_u10_n19542 ), .A2(_u10_n19543 ), .A3(_u10_n19544 ), .A4(_u10_n19545 ), .ZN(_u10_n19541 ) );
NOR4_X1 _u10_U8163  ( .A1(_u10_n19538 ), .A2(_u10_n19539 ), .A3(_u10_n19540 ), .A4(_u10_n19541 ), .ZN(_u10_n19537 ) );
NAND2_X1 _u10_U8162  ( .A1(_u10_n19536 ), .A2(_u10_n19537 ), .ZN(am0[26]) );
NAND2_X1 _u10_U8161  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19532 ) );
NAND2_X1 _u10_U8160  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19533 ) );
NAND2_X1 _u10_U8159  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19534 ) );
NAND2_X1 _u10_U8158  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19535 ) );
NAND4_X1 _u10_U8157  ( .A1(_u10_n19532 ), .A2(_u10_n19533 ), .A3(_u10_n19534 ), .A4(_u10_n19535 ), .ZN(_u10_n19517 ) );
NAND2_X1 _u10_U8156  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19528 ) );
NAND2_X1 _u10_U8155  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19529 ) );
NAND2_X1 _u10_U8154  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19530 ) );
NAND2_X1 _u10_U8153  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19531 ) );
NAND4_X1 _u10_U8152  ( .A1(_u10_n19528 ), .A2(_u10_n19529 ), .A3(_u10_n19530 ), .A4(_u10_n19531 ), .ZN(_u10_n19518 ) );
NAND2_X1 _u10_U8151  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19524 ) );
NAND2_X1 _u10_U8150  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19525 ) );
NAND2_X1 _u10_U8149  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19526 ) );
NAND2_X1 _u10_U8148  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19527 ) );
NAND4_X1 _u10_U8147  ( .A1(_u10_n19524 ), .A2(_u10_n19525 ), .A3(_u10_n19526 ), .A4(_u10_n19527 ), .ZN(_u10_n19519 ) );
NAND2_X1 _u10_U8146  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19521 ) );
NAND2_X1 _u10_U8145  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19522 ) );
NAND2_X1 _u10_U8144  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19523 ) );
NAND3_X1 _u10_U8143  ( .A1(_u10_n19521 ), .A2(_u10_n19522 ), .A3(_u10_n19523 ), .ZN(_u10_n19520 ) );
NOR4_X1 _u10_U8142  ( .A1(_u10_n19517 ), .A2(_u10_n19518 ), .A3(_u10_n19519 ), .A4(_u10_n19520 ), .ZN(_u10_n19495 ) );
NAND2_X1 _u10_U8141  ( .A1(1'b1), .A2(_u10_n11989 ), .ZN(_u10_n19513 ) );
NAND2_X1 _u10_U8140  ( .A1(1'b1), .A2(_u10_n11965 ), .ZN(_u10_n19514 ) );
NAND2_X1 _u10_U8139  ( .A1(1'b1), .A2(_u10_n11941 ), .ZN(_u10_n19515 ) );
NAND2_X1 _u10_U8138  ( .A1(1'b1), .A2(_u10_n11917 ), .ZN(_u10_n19516 ) );
NAND4_X1 _u10_U8137  ( .A1(_u10_n19513 ), .A2(_u10_n19514 ), .A3(_u10_n19515 ), .A4(_u10_n19516 ), .ZN(_u10_n19497 ) );
NAND2_X1 _u10_U8136  ( .A1(1'b1), .A2(_u10_n11893 ), .ZN(_u10_n19509 ) );
NAND2_X1 _u10_U8135  ( .A1(1'b1), .A2(_u10_n11869 ), .ZN(_u10_n19510 ) );
NAND2_X1 _u10_U8134  ( .A1(1'b1), .A2(_u10_n11845 ), .ZN(_u10_n19511 ) );
NAND2_X1 _u10_U8133  ( .A1(1'b1), .A2(_u10_n11821 ), .ZN(_u10_n19512 ) );
NAND4_X1 _u10_U8132  ( .A1(_u10_n19509 ), .A2(_u10_n19510 ), .A3(_u10_n19511 ), .A4(_u10_n19512 ), .ZN(_u10_n19498 ) );
NAND2_X1 _u10_U8131  ( .A1(1'b1), .A2(_u10_n11797 ), .ZN(_u10_n19505 ) );
NAND2_X1 _u10_U8130  ( .A1(1'b1), .A2(_u10_n11773 ), .ZN(_u10_n19506 ) );
NAND2_X1 _u10_U8129  ( .A1(1'b1), .A2(_u10_n11749 ), .ZN(_u10_n19507 ) );
NAND2_X1 _u10_U8128  ( .A1(1'b1), .A2(_u10_n11725 ), .ZN(_u10_n19508 ) );
NAND4_X1 _u10_U8127  ( .A1(_u10_n19505 ), .A2(_u10_n19506 ), .A3(_u10_n19507 ), .A4(_u10_n19508 ), .ZN(_u10_n19499 ) );
NAND2_X1 _u10_U8126  ( .A1(1'b1), .A2(_u10_n11701 ), .ZN(_u10_n19501 ) );
NAND2_X1 _u10_U8125  ( .A1(1'b1), .A2(_u10_n11677 ), .ZN(_u10_n19502 ) );
NAND2_X1 _u10_U8124  ( .A1(1'b1), .A2(_u10_n11653 ), .ZN(_u10_n19503 ) );
NAND2_X1 _u10_U8123  ( .A1(1'b1), .A2(_u10_n11629 ), .ZN(_u10_n19504 ) );
NAND4_X1 _u10_U8122  ( .A1(_u10_n19501 ), .A2(_u10_n19502 ), .A3(_u10_n19503 ), .A4(_u10_n19504 ), .ZN(_u10_n19500 ) );
NOR4_X1 _u10_U8121  ( .A1(_u10_n19497 ), .A2(_u10_n19498 ), .A3(_u10_n19499 ), .A4(_u10_n19500 ), .ZN(_u10_n19496 ) );
NAND2_X1 _u10_U8120  ( .A1(_u10_n19495 ), .A2(_u10_n19496 ), .ZN(am0[27]) );
NAND2_X1 _u10_U8119  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19491 ) );
NAND2_X1 _u10_U8118  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19492 ) );
NAND2_X1 _u10_U8117  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19493 ) );
NAND2_X1 _u10_U8116  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19494 ) );
NAND4_X1 _u10_U8115  ( .A1(_u10_n19491 ), .A2(_u10_n19492 ), .A3(_u10_n19493 ), .A4(_u10_n19494 ), .ZN(_u10_n19476 ) );
NAND2_X1 _u10_U8114  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19487 ) );
NAND2_X1 _u10_U8113  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19488 ) );
NAND2_X1 _u10_U8112  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19489 ) );
NAND2_X1 _u10_U8111  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19490 ) );
NAND4_X1 _u10_U8110  ( .A1(_u10_n19487 ), .A2(_u10_n19488 ), .A3(_u10_n19489 ), .A4(_u10_n19490 ), .ZN(_u10_n19477 ) );
NAND2_X1 _u10_U8109  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19483 ) );
NAND2_X1 _u10_U8108  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19484 ) );
NAND2_X1 _u10_U8107  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19485 ) );
NAND2_X1 _u10_U8106  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19486 ) );
NAND4_X1 _u10_U8105  ( .A1(_u10_n19483 ), .A2(_u10_n19484 ), .A3(_u10_n19485 ), .A4(_u10_n19486 ), .ZN(_u10_n19478 ) );
NAND2_X1 _u10_U8104  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19480 ) );
NAND2_X1 _u10_U8103  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19481 ) );
NAND2_X1 _u10_U8102  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19482 ) );
NAND3_X1 _u10_U8101  ( .A1(_u10_n19480 ), .A2(_u10_n19481 ), .A3(_u10_n19482 ), .ZN(_u10_n19479 ) );
NOR4_X1 _u10_U8100  ( .A1(_u10_n19476 ), .A2(_u10_n19477 ), .A3(_u10_n19478 ), .A4(_u10_n19479 ), .ZN(_u10_n19454 ) );
NAND2_X1 _u10_U8099  ( .A1(1'b1), .A2(_u10_n11989 ), .ZN(_u10_n19472 ) );
NAND2_X1 _u10_U8098  ( .A1(1'b1), .A2(_u10_n11965 ), .ZN(_u10_n19473 ) );
NAND2_X1 _u10_U8097  ( .A1(1'b1), .A2(_u10_n11941 ), .ZN(_u10_n19474 ) );
NAND2_X1 _u10_U8096  ( .A1(1'b1), .A2(_u10_n11917 ), .ZN(_u10_n19475 ) );
NAND4_X1 _u10_U8095  ( .A1(_u10_n19472 ), .A2(_u10_n19473 ), .A3(_u10_n19474 ), .A4(_u10_n19475 ), .ZN(_u10_n19456 ) );
NAND2_X1 _u10_U8094  ( .A1(1'b1), .A2(_u10_n11893 ), .ZN(_u10_n19468 ) );
NAND2_X1 _u10_U8093  ( .A1(1'b1), .A2(_u10_n11869 ), .ZN(_u10_n19469 ) );
NAND2_X1 _u10_U8092  ( .A1(1'b1), .A2(_u10_n11845 ), .ZN(_u10_n19470 ) );
NAND2_X1 _u10_U8091  ( .A1(1'b1), .A2(_u10_n11821 ), .ZN(_u10_n19471 ) );
NAND4_X1 _u10_U8090  ( .A1(_u10_n19468 ), .A2(_u10_n19469 ), .A3(_u10_n19470 ), .A4(_u10_n19471 ), .ZN(_u10_n19457 ) );
NAND2_X1 _u10_U8089  ( .A1(1'b1), .A2(_u10_n11797 ), .ZN(_u10_n19464 ) );
NAND2_X1 _u10_U8088  ( .A1(1'b1), .A2(_u10_n11773 ), .ZN(_u10_n19465 ) );
NAND2_X1 _u10_U8087  ( .A1(1'b1), .A2(_u10_n11749 ), .ZN(_u10_n19466 ) );
NAND2_X1 _u10_U8086  ( .A1(1'b1), .A2(_u10_n11725 ), .ZN(_u10_n19467 ) );
NAND4_X1 _u10_U8085  ( .A1(_u10_n19464 ), .A2(_u10_n19465 ), .A3(_u10_n19466 ), .A4(_u10_n19467 ), .ZN(_u10_n19458 ) );
NAND2_X1 _u10_U8084  ( .A1(1'b1), .A2(_u10_n11701 ), .ZN(_u10_n19460 ) );
NAND2_X1 _u10_U8083  ( .A1(1'b1), .A2(_u10_n11677 ), .ZN(_u10_n19461 ) );
NAND2_X1 _u10_U8082  ( .A1(1'b1), .A2(_u10_n11653 ), .ZN(_u10_n19462 ) );
NAND2_X1 _u10_U8081  ( .A1(1'b1), .A2(_u10_n11629 ), .ZN(_u10_n19463 ) );
NAND4_X1 _u10_U8080  ( .A1(_u10_n19460 ), .A2(_u10_n19461 ), .A3(_u10_n19462 ), .A4(_u10_n19463 ), .ZN(_u10_n19459 ) );
NOR4_X1 _u10_U8079  ( .A1(_u10_n19456 ), .A2(_u10_n19457 ), .A3(_u10_n19458 ), .A4(_u10_n19459 ), .ZN(_u10_n19455 ) );
NAND2_X1 _u10_U8078  ( .A1(_u10_n19454 ), .A2(_u10_n19455 ), .ZN(am0[28]) );
NAND2_X1 _u10_U8077  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19450 ) );
NAND2_X1 _u10_U8076  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19451 ) );
NAND2_X1 _u10_U8075  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19452 ) );
NAND2_X1 _u10_U8074  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19453 ) );
NAND4_X1 _u10_U8073  ( .A1(_u10_n19450 ), .A2(_u10_n19451 ), .A3(_u10_n19452 ), .A4(_u10_n19453 ), .ZN(_u10_n19435 ) );
NAND2_X1 _u10_U8072  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19446 ) );
NAND2_X1 _u10_U8071  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19447 ) );
NAND2_X1 _u10_U8070  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19448 ) );
NAND2_X1 _u10_U8069  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19449 ) );
NAND4_X1 _u10_U8068  ( .A1(_u10_n19446 ), .A2(_u10_n19447 ), .A3(_u10_n19448 ), .A4(_u10_n19449 ), .ZN(_u10_n19436 ) );
NAND2_X1 _u10_U8067  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19442 ) );
NAND2_X1 _u10_U8066  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19443 ) );
NAND2_X1 _u10_U8065  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19444 ) );
NAND2_X1 _u10_U8064  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19445 ) );
NAND4_X1 _u10_U8063  ( .A1(_u10_n19442 ), .A2(_u10_n19443 ), .A3(_u10_n19444 ), .A4(_u10_n19445 ), .ZN(_u10_n19437 ) );
NAND2_X1 _u10_U8062  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19439 ) );
NAND2_X1 _u10_U8061  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19440 ) );
NAND2_X1 _u10_U8060  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19441 ) );
NAND3_X1 _u10_U8059  ( .A1(_u10_n19439 ), .A2(_u10_n19440 ), .A3(_u10_n19441 ), .ZN(_u10_n19438 ) );
NOR4_X1 _u10_U8058  ( .A1(_u10_n19435 ), .A2(_u10_n19436 ), .A3(_u10_n19437 ), .A4(_u10_n19438 ), .ZN(_u10_n19413 ) );
NAND2_X1 _u10_U8057  ( .A1(1'b1), .A2(_u10_n11989 ), .ZN(_u10_n19431 ) );
NAND2_X1 _u10_U8056  ( .A1(1'b1), .A2(_u10_n11965 ), .ZN(_u10_n19432 ) );
NAND2_X1 _u10_U8055  ( .A1(1'b1), .A2(_u10_n11941 ), .ZN(_u10_n19433 ) );
NAND2_X1 _u10_U8054  ( .A1(1'b1), .A2(_u10_n11917 ), .ZN(_u10_n19434 ) );
NAND4_X1 _u10_U8053  ( .A1(_u10_n19431 ), .A2(_u10_n19432 ), .A3(_u10_n19433 ), .A4(_u10_n19434 ), .ZN(_u10_n19415 ) );
NAND2_X1 _u10_U8052  ( .A1(1'b1), .A2(_u10_n11893 ), .ZN(_u10_n19427 ) );
NAND2_X1 _u10_U8051  ( .A1(1'b1), .A2(_u10_n11869 ), .ZN(_u10_n19428 ) );
NAND2_X1 _u10_U8050  ( .A1(1'b1), .A2(_u10_n11845 ), .ZN(_u10_n19429 ) );
NAND2_X1 _u10_U8049  ( .A1(1'b1), .A2(_u10_n11821 ), .ZN(_u10_n19430 ) );
NAND4_X1 _u10_U8048  ( .A1(_u10_n19427 ), .A2(_u10_n19428 ), .A3(_u10_n19429 ), .A4(_u10_n19430 ), .ZN(_u10_n19416 ) );
NAND2_X1 _u10_U8047  ( .A1(1'b1), .A2(_u10_n11797 ), .ZN(_u10_n19423 ) );
NAND2_X1 _u10_U8046  ( .A1(1'b1), .A2(_u10_n11773 ), .ZN(_u10_n19424 ) );
NAND2_X1 _u10_U8045  ( .A1(1'b1), .A2(_u10_n11749 ), .ZN(_u10_n19425 ) );
NAND2_X1 _u10_U8044  ( .A1(1'b1), .A2(_u10_n11725 ), .ZN(_u10_n19426 ) );
NAND4_X1 _u10_U8043  ( .A1(_u10_n19423 ), .A2(_u10_n19424 ), .A3(_u10_n19425 ), .A4(_u10_n19426 ), .ZN(_u10_n19417 ) );
NAND2_X1 _u10_U8042  ( .A1(1'b1), .A2(_u10_n11701 ), .ZN(_u10_n19419 ) );
NAND2_X1 _u10_U8041  ( .A1(1'b1), .A2(_u10_n11677 ), .ZN(_u10_n19420 ) );
NAND2_X1 _u10_U8040  ( .A1(1'b1), .A2(_u10_n11653 ), .ZN(_u10_n19421 ) );
NAND2_X1 _u10_U8039  ( .A1(1'b1), .A2(_u10_n11629 ), .ZN(_u10_n19422 ) );
NAND4_X1 _u10_U8038  ( .A1(_u10_n19419 ), .A2(_u10_n19420 ), .A3(_u10_n19421 ), .A4(_u10_n19422 ), .ZN(_u10_n19418 ) );
NOR4_X1 _u10_U8037  ( .A1(_u10_n19415 ), .A2(_u10_n19416 ), .A3(_u10_n19417 ), .A4(_u10_n19418 ), .ZN(_u10_n19414 ) );
NAND2_X1 _u10_U8036  ( .A1(_u10_n19413 ), .A2(_u10_n19414 ), .ZN(am0[29]) );
NAND2_X1 _u10_U8035  ( .A1(1'b0), .A2(_u10_n12336 ), .ZN(_u10_n19409 ) );
NAND2_X1 _u10_U8034  ( .A1(1'b0), .A2(_u10_n12313 ), .ZN(_u10_n19410 ) );
NAND2_X1 _u10_U8033  ( .A1(1'b0), .A2(_u10_n12289 ), .ZN(_u10_n19411 ) );
NAND2_X1 _u10_U8032  ( .A1(1'b0), .A2(_u10_n12265 ), .ZN(_u10_n19412 ) );
NAND4_X1 _u10_U8031  ( .A1(_u10_n19409 ), .A2(_u10_n19410 ), .A3(_u10_n19411 ), .A4(_u10_n19412 ), .ZN(_u10_n19394 ) );
NAND2_X1 _u10_U8030  ( .A1(1'b0), .A2(_u10_n12240 ), .ZN(_u10_n19405 ) );
NAND2_X1 _u10_U8029  ( .A1(1'b0), .A2(_u10_n12216 ), .ZN(_u10_n19406 ) );
NAND2_X1 _u10_U8028  ( .A1(1'b0), .A2(_u10_n12193 ), .ZN(_u10_n19407 ) );
NAND2_X1 _u10_U8027  ( .A1(1'b0), .A2(_u10_n12168 ), .ZN(_u10_n19408 ) );
NAND4_X1 _u10_U8026  ( .A1(_u10_n19405 ), .A2(_u10_n19406 ), .A3(_u10_n19407 ), .A4(_u10_n19408 ), .ZN(_u10_n19395 ) );
NAND2_X1 _u10_U8025  ( .A1(1'b0), .A2(_u10_n12145 ), .ZN(_u10_n19401 ) );
NAND2_X1 _u10_U8024  ( .A1(1'b0), .A2(_u10_n12121 ), .ZN(_u10_n19402 ) );
NAND2_X1 _u10_U8023  ( .A1(1'b0), .A2(_u10_n12097 ), .ZN(_u10_n19403 ) );
NAND2_X1 _u10_U8022  ( .A1(1'b0), .A2(_u10_n12073 ), .ZN(_u10_n19404 ) );
NAND4_X1 _u10_U8021  ( .A1(_u10_n19401 ), .A2(_u10_n19402 ), .A3(_u10_n19403 ), .A4(_u10_n19404 ), .ZN(_u10_n19396 ) );
NAND2_X1 _u10_U8020  ( .A1(1'b0), .A2(_u10_n12049 ), .ZN(_u10_n19398 ) );
NAND2_X1 _u10_U8019  ( .A1(1'b0), .A2(_u10_n12025 ), .ZN(_u10_n19399 ) );
NAND2_X1 _u10_U8018  ( .A1(1'b0), .A2(_u10_n12006 ), .ZN(_u10_n19400 ) );
NAND3_X1 _u10_U8017  ( .A1(_u10_n19398 ), .A2(_u10_n19399 ), .A3(_u10_n19400 ), .ZN(_u10_n19397 ) );
NOR4_X1 _u10_U8016  ( .A1(_u10_n19394 ), .A2(_u10_n19395 ), .A3(_u10_n19396 ), .A4(_u10_n19397 ), .ZN(_u10_n19372 ) );
NAND2_X1 _u10_U8015  ( .A1(1'b0), .A2(_u10_n11989 ), .ZN(_u10_n19390 ) );
NAND2_X1 _u10_U8014  ( .A1(1'b0), .A2(_u10_n11965 ), .ZN(_u10_n19391 ) );
NAND2_X1 _u10_U8013  ( .A1(1'b0), .A2(_u10_n11941 ), .ZN(_u10_n19392 ) );
NAND2_X1 _u10_U8012  ( .A1(1'b0), .A2(_u10_n11917 ), .ZN(_u10_n19393 ) );
NAND4_X1 _u10_U8011  ( .A1(_u10_n19390 ), .A2(_u10_n19391 ), .A3(_u10_n19392 ), .A4(_u10_n19393 ), .ZN(_u10_n19374 ) );
NAND2_X1 _u10_U8010  ( .A1(1'b0), .A2(_u10_n11893 ), .ZN(_u10_n19386 ) );
NAND2_X1 _u10_U8009  ( .A1(1'b0), .A2(_u10_n11869 ), .ZN(_u10_n19387 ) );
NAND2_X1 _u10_U8008  ( .A1(1'b0), .A2(_u10_n11845 ), .ZN(_u10_n19388 ) );
NAND2_X1 _u10_U8007  ( .A1(1'b0), .A2(_u10_n11821 ), .ZN(_u10_n19389 ) );
NAND4_X1 _u10_U8006  ( .A1(_u10_n19386 ), .A2(_u10_n19387 ), .A3(_u10_n19388 ), .A4(_u10_n19389 ), .ZN(_u10_n19375 ) );
NAND2_X1 _u10_U8005  ( .A1(1'b0), .A2(_u10_n11797 ), .ZN(_u10_n19382 ) );
NAND2_X1 _u10_U8004  ( .A1(1'b0), .A2(_u10_n11773 ), .ZN(_u10_n19383 ) );
NAND2_X1 _u10_U8003  ( .A1(1'b0), .A2(_u10_n11749 ), .ZN(_u10_n19384 ) );
NAND2_X1 _u10_U8002  ( .A1(1'b0), .A2(_u10_n11725 ), .ZN(_u10_n19385 ) );
NAND4_X1 _u10_U8001  ( .A1(_u10_n19382 ), .A2(_u10_n19383 ), .A3(_u10_n19384 ), .A4(_u10_n19385 ), .ZN(_u10_n19376 ) );
NAND2_X1 _u10_U8000  ( .A1(1'b0), .A2(_u10_n11701 ), .ZN(_u10_n19378 ) );
NAND2_X1 _u10_U7999  ( .A1(1'b0), .A2(_u10_n11677 ), .ZN(_u10_n19379 ) );
NAND2_X1 _u10_U7998  ( .A1(1'b0), .A2(_u10_n11653 ), .ZN(_u10_n19380 ) );
NAND2_X1 _u10_U7997  ( .A1(1'b0), .A2(_u10_n11629 ), .ZN(_u10_n19381 ) );
NAND4_X1 _u10_U7996  ( .A1(_u10_n19378 ), .A2(_u10_n19379 ), .A3(_u10_n19380 ), .A4(_u10_n19381 ), .ZN(_u10_n19377 ) );
NOR4_X1 _u10_U7995  ( .A1(_u10_n19374 ), .A2(_u10_n19375 ), .A3(_u10_n19376 ), .A4(_u10_n19377 ), .ZN(_u10_n19373 ) );
NAND2_X1 _u10_U7994  ( .A1(_u10_n19372 ), .A2(_u10_n19373 ), .ZN(am0[2]) );
NAND2_X1 _u10_U7993  ( .A1(1'b1), .A2(_u10_n12336 ), .ZN(_u10_n19368 ) );
NAND2_X1 _u10_U7992  ( .A1(1'b1), .A2(_u10_n12313 ), .ZN(_u10_n19369 ) );
NAND2_X1 _u10_U7991  ( .A1(1'b1), .A2(_u10_n12289 ), .ZN(_u10_n19370 ) );
NAND2_X1 _u10_U7990  ( .A1(1'b1), .A2(_u10_n12265 ), .ZN(_u10_n19371 ) );
NAND4_X1 _u10_U7989  ( .A1(_u10_n19368 ), .A2(_u10_n19369 ), .A3(_u10_n19370 ), .A4(_u10_n19371 ), .ZN(_u10_n19353 ) );
NAND2_X1 _u10_U7988  ( .A1(1'b1), .A2(_u10_n12240 ), .ZN(_u10_n19364 ) );
NAND2_X1 _u10_U7987  ( .A1(1'b1), .A2(_u10_n12216 ), .ZN(_u10_n19365 ) );
NAND2_X1 _u10_U7986  ( .A1(1'b1), .A2(_u10_n12193 ), .ZN(_u10_n19366 ) );
NAND2_X1 _u10_U7985  ( .A1(1'b1), .A2(_u10_n12168 ), .ZN(_u10_n19367 ) );
NAND4_X1 _u10_U7984  ( .A1(_u10_n19364 ), .A2(_u10_n19365 ), .A3(_u10_n19366 ), .A4(_u10_n19367 ), .ZN(_u10_n19354 ) );
NAND2_X1 _u10_U7983  ( .A1(1'b1), .A2(_u10_n12145 ), .ZN(_u10_n19360 ) );
NAND2_X1 _u10_U7982  ( .A1(1'b1), .A2(_u10_n12121 ), .ZN(_u10_n19361 ) );
NAND2_X1 _u10_U7981  ( .A1(1'b1), .A2(_u10_n12097 ), .ZN(_u10_n19362 ) );
NAND2_X1 _u10_U7980  ( .A1(1'b1), .A2(_u10_n12073 ), .ZN(_u10_n19363 ) );
NAND4_X1 _u10_U7979  ( .A1(_u10_n19360 ), .A2(_u10_n19361 ), .A3(_u10_n19362 ), .A4(_u10_n19363 ), .ZN(_u10_n19355 ) );
NAND2_X1 _u10_U7978  ( .A1(1'b1), .A2(_u10_n12049 ), .ZN(_u10_n19357 ) );
NAND2_X1 _u10_U7977  ( .A1(1'b1), .A2(_u10_n12025 ), .ZN(_u10_n19358 ) );
NAND2_X1 _u10_U7976  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19359 ) );
NAND3_X1 _u10_U7975  ( .A1(_u10_n19357 ), .A2(_u10_n19358 ), .A3(_u10_n19359 ), .ZN(_u10_n19356 ) );
NOR4_X1 _u10_U7974  ( .A1(_u10_n19353 ), .A2(_u10_n19354 ), .A3(_u10_n19355 ), .A4(_u10_n19356 ), .ZN(_u10_n19331 ) );
NAND2_X1 _u10_U7973  ( .A1(1'b1), .A2(_u10_n11989 ), .ZN(_u10_n19349 ) );
NAND2_X1 _u10_U7972  ( .A1(1'b1), .A2(_u10_n11965 ), .ZN(_u10_n19350 ) );
NAND2_X1 _u10_U7971  ( .A1(1'b1), .A2(_u10_n11941 ), .ZN(_u10_n19351 ) );
NAND2_X1 _u10_U7970  ( .A1(1'b1), .A2(_u10_n11917 ), .ZN(_u10_n19352 ) );
NAND4_X1 _u10_U7969  ( .A1(_u10_n19349 ), .A2(_u10_n19350 ), .A3(_u10_n19351 ), .A4(_u10_n19352 ), .ZN(_u10_n19333 ) );
NAND2_X1 _u10_U7968  ( .A1(1'b1), .A2(_u10_n11893 ), .ZN(_u10_n19345 ) );
NAND2_X1 _u10_U7967  ( .A1(1'b1), .A2(_u10_n11869 ), .ZN(_u10_n19346 ) );
NAND2_X1 _u10_U7966  ( .A1(1'b1), .A2(_u10_n11845 ), .ZN(_u10_n19347 ) );
NAND2_X1 _u10_U7965  ( .A1(1'b1), .A2(_u10_n11821 ), .ZN(_u10_n19348 ) );
NAND4_X1 _u10_U7964  ( .A1(_u10_n19345 ), .A2(_u10_n19346 ), .A3(_u10_n19347 ), .A4(_u10_n19348 ), .ZN(_u10_n19334 ) );
NAND2_X1 _u10_U7963  ( .A1(1'b1), .A2(_u10_n11797 ), .ZN(_u10_n19341 ) );
NAND2_X1 _u10_U7962  ( .A1(1'b1), .A2(_u10_n11773 ), .ZN(_u10_n19342 ) );
NAND2_X1 _u10_U7961  ( .A1(1'b1), .A2(_u10_n11749 ), .ZN(_u10_n19343 ) );
NAND2_X1 _u10_U7960  ( .A1(1'b1), .A2(_u10_n11725 ), .ZN(_u10_n19344 ) );
NAND4_X1 _u10_U7959  ( .A1(_u10_n19341 ), .A2(_u10_n19342 ), .A3(_u10_n19343 ), .A4(_u10_n19344 ), .ZN(_u10_n19335 ) );
NAND2_X1 _u10_U7958  ( .A1(1'b1), .A2(_u10_n11701 ), .ZN(_u10_n19337 ) );
NAND2_X1 _u10_U7957  ( .A1(1'b1), .A2(_u10_n11677 ), .ZN(_u10_n19338 ) );
NAND2_X1 _u10_U7956  ( .A1(1'b1), .A2(_u10_n11653 ), .ZN(_u10_n19339 ) );
NAND2_X1 _u10_U7955  ( .A1(1'b1), .A2(_u10_n11629 ), .ZN(_u10_n19340 ) );
NAND4_X1 _u10_U7954  ( .A1(_u10_n19337 ), .A2(_u10_n19338 ), .A3(_u10_n19339 ), .A4(_u10_n19340 ), .ZN(_u10_n19336 ) );
NOR4_X1 _u10_U7953  ( .A1(_u10_n19333 ), .A2(_u10_n19334 ), .A3(_u10_n19335 ), .A4(_u10_n19336 ), .ZN(_u10_n19332 ) );
NAND2_X1 _u10_U7952  ( .A1(_u10_n19331 ), .A2(_u10_n19332 ), .ZN(am0[30]) );
NAND2_X1 _u10_U7951  ( .A1(1'b1), .A2(_u10_n12337 ), .ZN(_u10_n19327 ) );
NAND2_X1 _u10_U7950  ( .A1(1'b1), .A2(_u10_n12314 ), .ZN(_u10_n19328 ) );
NAND2_X1 _u10_U7949  ( .A1(1'b1), .A2(_u10_n12290 ), .ZN(_u10_n19329 ) );
NAND2_X1 _u10_U7948  ( .A1(1'b1), .A2(_u10_n12266 ), .ZN(_u10_n19330 ) );
NAND4_X1 _u10_U7947  ( .A1(_u10_n19327 ), .A2(_u10_n19328 ), .A3(_u10_n19329 ), .A4(_u10_n19330 ), .ZN(_u10_n19312 ) );
NAND2_X1 _u10_U7946  ( .A1(1'b1), .A2(_u10_n12241 ), .ZN(_u10_n19323 ) );
NAND2_X1 _u10_U7945  ( .A1(1'b1), .A2(_u10_n12217 ), .ZN(_u10_n19324 ) );
NAND2_X1 _u10_U7944  ( .A1(1'b1), .A2(_u10_n12194 ), .ZN(_u10_n19325 ) );
NAND2_X1 _u10_U7943  ( .A1(1'b1), .A2(_u10_n12169 ), .ZN(_u10_n19326 ) );
NAND4_X1 _u10_U7942  ( .A1(_u10_n19323 ), .A2(_u10_n19324 ), .A3(_u10_n19325 ), .A4(_u10_n19326 ), .ZN(_u10_n19313 ) );
NAND2_X1 _u10_U7941  ( .A1(1'b1), .A2(_u10_n12146 ), .ZN(_u10_n19319 ) );
NAND2_X1 _u10_U7940  ( .A1(1'b1), .A2(_u10_n12122 ), .ZN(_u10_n19320 ) );
NAND2_X1 _u10_U7939  ( .A1(1'b1), .A2(_u10_n12098 ), .ZN(_u10_n19321 ) );
NAND2_X1 _u10_U7938  ( .A1(1'b1), .A2(_u10_n12074 ), .ZN(_u10_n19322 ) );
NAND4_X1 _u10_U7937  ( .A1(_u10_n19319 ), .A2(_u10_n19320 ), .A3(_u10_n19321 ), .A4(_u10_n19322 ), .ZN(_u10_n19314 ) );
NAND2_X1 _u10_U7936  ( .A1(1'b1), .A2(_u10_n12050 ), .ZN(_u10_n19316 ) );
NAND2_X1 _u10_U7935  ( .A1(1'b1), .A2(_u10_n12026 ), .ZN(_u10_n19317 ) );
NAND2_X1 _u10_U7934  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19318 ) );
NAND3_X1 _u10_U7933  ( .A1(_u10_n19316 ), .A2(_u10_n19317 ), .A3(_u10_n19318 ), .ZN(_u10_n19315 ) );
NOR4_X1 _u10_U7932  ( .A1(_u10_n19312 ), .A2(_u10_n19313 ), .A3(_u10_n19314 ), .A4(_u10_n19315 ), .ZN(_u10_n19290 ) );
NAND2_X1 _u10_U7931  ( .A1(1'b1), .A2(_u10_n11989 ), .ZN(_u10_n19308 ) );
NAND2_X1 _u10_U7930  ( .A1(1'b1), .A2(_u10_n11965 ), .ZN(_u10_n19309 ) );
NAND2_X1 _u10_U7929  ( .A1(1'b1), .A2(_u10_n11941 ), .ZN(_u10_n19310 ) );
NAND2_X1 _u10_U7928  ( .A1(1'b1), .A2(_u10_n11917 ), .ZN(_u10_n19311 ) );
NAND4_X1 _u10_U7927  ( .A1(_u10_n19308 ), .A2(_u10_n19309 ), .A3(_u10_n19310 ), .A4(_u10_n19311 ), .ZN(_u10_n19292 ) );
NAND2_X1 _u10_U7926  ( .A1(1'b1), .A2(_u10_n11893 ), .ZN(_u10_n19304 ) );
NAND2_X1 _u10_U7925  ( .A1(1'b1), .A2(_u10_n11869 ), .ZN(_u10_n19305 ) );
NAND2_X1 _u10_U7924  ( .A1(1'b1), .A2(_u10_n11845 ), .ZN(_u10_n19306 ) );
NAND2_X1 _u10_U7923  ( .A1(1'b1), .A2(_u10_n11821 ), .ZN(_u10_n19307 ) );
NAND4_X1 _u10_U7922  ( .A1(_u10_n19304 ), .A2(_u10_n19305 ), .A3(_u10_n19306 ), .A4(_u10_n19307 ), .ZN(_u10_n19293 ) );
NAND2_X1 _u10_U7921  ( .A1(1'b1), .A2(_u10_n11797 ), .ZN(_u10_n19300 ) );
NAND2_X1 _u10_U7920  ( .A1(1'b1), .A2(_u10_n11773 ), .ZN(_u10_n19301 ) );
NAND2_X1 _u10_U7919  ( .A1(1'b1), .A2(_u10_n11749 ), .ZN(_u10_n19302 ) );
NAND2_X1 _u10_U7918  ( .A1(1'b1), .A2(_u10_n11725 ), .ZN(_u10_n19303 ) );
NAND4_X1 _u10_U7917  ( .A1(_u10_n19300 ), .A2(_u10_n19301 ), .A3(_u10_n19302 ), .A4(_u10_n19303 ), .ZN(_u10_n19294 ) );
NAND2_X1 _u10_U7916  ( .A1(1'b1), .A2(_u10_n11701 ), .ZN(_u10_n19296 ) );
NAND2_X1 _u10_U7915  ( .A1(1'b1), .A2(_u10_n11677 ), .ZN(_u10_n19297 ) );
NAND2_X1 _u10_U7914  ( .A1(1'b1), .A2(_u10_n11653 ), .ZN(_u10_n19298 ) );
NAND2_X1 _u10_U7913  ( .A1(1'b1), .A2(_u10_n11629 ), .ZN(_u10_n19299 ) );
NAND4_X1 _u10_U7912  ( .A1(_u10_n19296 ), .A2(_u10_n19297 ), .A3(_u10_n19298 ), .A4(_u10_n19299 ), .ZN(_u10_n19295 ) );
NOR4_X1 _u10_U7911  ( .A1(_u10_n19292 ), .A2(_u10_n19293 ), .A3(_u10_n19294 ), .A4(_u10_n19295 ), .ZN(_u10_n19291 ) );
NAND2_X1 _u10_U7910  ( .A1(_u10_n19290 ), .A2(_u10_n19291 ), .ZN(am0[31]) );
NAND2_X1 _u10_U7909  ( .A1(1'b0), .A2(_u10_n12337 ), .ZN(_u10_n19286 ) );
NAND2_X1 _u10_U7908  ( .A1(1'b0), .A2(_u10_n12314 ), .ZN(_u10_n19287 ) );
NAND2_X1 _u10_U7907  ( .A1(1'b0), .A2(_u10_n12290 ), .ZN(_u10_n19288 ) );
NAND2_X1 _u10_U7906  ( .A1(1'b0), .A2(_u10_n12266 ), .ZN(_u10_n19289 ) );
NAND4_X1 _u10_U7905  ( .A1(_u10_n19286 ), .A2(_u10_n19287 ), .A3(_u10_n19288 ), .A4(_u10_n19289 ), .ZN(_u10_n19271 ) );
NAND2_X1 _u10_U7904  ( .A1(1'b0), .A2(_u10_n12241 ), .ZN(_u10_n19282 ) );
NAND2_X1 _u10_U7903  ( .A1(1'b0), .A2(_u10_n12217 ), .ZN(_u10_n19283 ) );
NAND2_X1 _u10_U7902  ( .A1(1'b0), .A2(_u10_n12194 ), .ZN(_u10_n19284 ) );
NAND2_X1 _u10_U7901  ( .A1(1'b0), .A2(_u10_n12169 ), .ZN(_u10_n19285 ) );
NAND4_X1 _u10_U7900  ( .A1(_u10_n19282 ), .A2(_u10_n19283 ), .A3(_u10_n19284 ), .A4(_u10_n19285 ), .ZN(_u10_n19272 ) );
NAND2_X1 _u10_U7899  ( .A1(1'b0), .A2(_u10_n12146 ), .ZN(_u10_n19278 ) );
NAND2_X1 _u10_U7898  ( .A1(1'b0), .A2(_u10_n12122 ), .ZN(_u10_n19279 ) );
NAND2_X1 _u10_U7897  ( .A1(1'b0), .A2(_u10_n12098 ), .ZN(_u10_n19280 ) );
NAND2_X1 _u10_U7896  ( .A1(1'b0), .A2(_u10_n12074 ), .ZN(_u10_n19281 ) );
NAND4_X1 _u10_U7895  ( .A1(_u10_n19278 ), .A2(_u10_n19279 ), .A3(_u10_n19280 ), .A4(_u10_n19281 ), .ZN(_u10_n19273 ) );
NAND2_X1 _u10_U7894  ( .A1(1'b0), .A2(_u10_n12050 ), .ZN(_u10_n19275 ) );
NAND2_X1 _u10_U7893  ( .A1(1'b0), .A2(_u10_n12026 ), .ZN(_u10_n19276 ) );
NAND2_X1 _u10_U7892  ( .A1(1'b0), .A2(_u10_n12006 ), .ZN(_u10_n19277 ) );
NAND3_X1 _u10_U7891  ( .A1(_u10_n19275 ), .A2(_u10_n19276 ), .A3(_u10_n19277 ), .ZN(_u10_n19274 ) );
NOR4_X1 _u10_U7890  ( .A1(_u10_n19271 ), .A2(_u10_n19272 ), .A3(_u10_n19273 ), .A4(_u10_n19274 ), .ZN(_u10_n19249 ) );
NAND2_X1 _u10_U7889  ( .A1(1'b0), .A2(_u10_n11989 ), .ZN(_u10_n19267 ) );
NAND2_X1 _u10_U7888  ( .A1(1'b0), .A2(_u10_n11965 ), .ZN(_u10_n19268 ) );
NAND2_X1 _u10_U7887  ( .A1(1'b0), .A2(_u10_n11941 ), .ZN(_u10_n19269 ) );
NAND2_X1 _u10_U7886  ( .A1(1'b0), .A2(_u10_n11917 ), .ZN(_u10_n19270 ) );
NAND4_X1 _u10_U7885  ( .A1(_u10_n19267 ), .A2(_u10_n19268 ), .A3(_u10_n19269 ), .A4(_u10_n19270 ), .ZN(_u10_n19251 ) );
NAND2_X1 _u10_U7884  ( .A1(1'b0), .A2(_u10_n11893 ), .ZN(_u10_n19263 ) );
NAND2_X1 _u10_U7883  ( .A1(1'b0), .A2(_u10_n11869 ), .ZN(_u10_n19264 ) );
NAND2_X1 _u10_U7882  ( .A1(1'b0), .A2(_u10_n11845 ), .ZN(_u10_n19265 ) );
NAND2_X1 _u10_U7881  ( .A1(1'b0), .A2(_u10_n11821 ), .ZN(_u10_n19266 ) );
NAND4_X1 _u10_U7880  ( .A1(_u10_n19263 ), .A2(_u10_n19264 ), .A3(_u10_n19265 ), .A4(_u10_n19266 ), .ZN(_u10_n19252 ) );
NAND2_X1 _u10_U7879  ( .A1(1'b0), .A2(_u10_n11797 ), .ZN(_u10_n19259 ) );
NAND2_X1 _u10_U7878  ( .A1(1'b0), .A2(_u10_n11773 ), .ZN(_u10_n19260 ) );
NAND2_X1 _u10_U7877  ( .A1(1'b0), .A2(_u10_n11749 ), .ZN(_u10_n19261 ) );
NAND2_X1 _u10_U7876  ( .A1(1'b0), .A2(_u10_n11725 ), .ZN(_u10_n19262 ) );
NAND4_X1 _u10_U7875  ( .A1(_u10_n19259 ), .A2(_u10_n19260 ), .A3(_u10_n19261 ), .A4(_u10_n19262 ), .ZN(_u10_n19253 ) );
NAND2_X1 _u10_U7874  ( .A1(1'b0), .A2(_u10_n11701 ), .ZN(_u10_n19255 ) );
NAND2_X1 _u10_U7873  ( .A1(1'b0), .A2(_u10_n11677 ), .ZN(_u10_n19256 ) );
NAND2_X1 _u10_U7872  ( .A1(1'b0), .A2(_u10_n11653 ), .ZN(_u10_n19257 ) );
NAND2_X1 _u10_U7871  ( .A1(1'b0), .A2(_u10_n11629 ), .ZN(_u10_n19258 ) );
NAND4_X1 _u10_U7870  ( .A1(_u10_n19255 ), .A2(_u10_n19256 ), .A3(_u10_n19257 ), .A4(_u10_n19258 ), .ZN(_u10_n19254 ) );
NOR4_X1 _u10_U7869  ( .A1(_u10_n19251 ), .A2(_u10_n19252 ), .A3(_u10_n19253 ), .A4(_u10_n19254 ), .ZN(_u10_n19250 ) );
NAND2_X1 _u10_U7868  ( .A1(_u10_n19249 ), .A2(_u10_n19250 ), .ZN(am0[3]) );
NAND2_X1 _u10_U7867  ( .A1(1'b1), .A2(_u10_n12337 ), .ZN(_u10_n19245 ) );
NAND2_X1 _u10_U7866  ( .A1(1'b1), .A2(_u10_n12314 ), .ZN(_u10_n19246 ) );
NAND2_X1 _u10_U7865  ( .A1(1'b1), .A2(_u10_n12290 ), .ZN(_u10_n19247 ) );
NAND2_X1 _u10_U7864  ( .A1(1'b1), .A2(_u10_n12266 ), .ZN(_u10_n19248 ) );
NAND4_X1 _u10_U7863  ( .A1(_u10_n19245 ), .A2(_u10_n19246 ), .A3(_u10_n19247 ), .A4(_u10_n19248 ), .ZN(_u10_n19230 ) );
NAND2_X1 _u10_U7862  ( .A1(1'b1), .A2(_u10_n12241 ), .ZN(_u10_n19241 ) );
NAND2_X1 _u10_U7861  ( .A1(1'b1), .A2(_u10_n12217 ), .ZN(_u10_n19242 ) );
NAND2_X1 _u10_U7860  ( .A1(1'b1), .A2(_u10_n12194 ), .ZN(_u10_n19243 ) );
NAND2_X1 _u10_U7859  ( .A1(1'b1), .A2(_u10_n12169 ), .ZN(_u10_n19244 ) );
NAND4_X1 _u10_U7858  ( .A1(_u10_n19241 ), .A2(_u10_n19242 ), .A3(_u10_n19243 ), .A4(_u10_n19244 ), .ZN(_u10_n19231 ) );
NAND2_X1 _u10_U7857  ( .A1(1'b1), .A2(_u10_n12146 ), .ZN(_u10_n19237 ) );
NAND2_X1 _u10_U7856  ( .A1(1'b1), .A2(_u10_n12122 ), .ZN(_u10_n19238 ) );
NAND2_X1 _u10_U7855  ( .A1(1'b1), .A2(_u10_n12098 ), .ZN(_u10_n19239 ) );
NAND2_X1 _u10_U7854  ( .A1(1'b1), .A2(_u10_n12074 ), .ZN(_u10_n19240 ) );
NAND4_X1 _u10_U7853  ( .A1(_u10_n19237 ), .A2(_u10_n19238 ), .A3(_u10_n19239 ), .A4(_u10_n19240 ), .ZN(_u10_n19232 ) );
NAND2_X1 _u10_U7852  ( .A1(1'b1), .A2(_u10_n12050 ), .ZN(_u10_n19234 ) );
NAND2_X1 _u10_U7851  ( .A1(1'b1), .A2(_u10_n12026 ), .ZN(_u10_n19235 ) );
NAND2_X1 _u10_U7850  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19236 ) );
NAND3_X1 _u10_U7849  ( .A1(_u10_n19234 ), .A2(_u10_n19235 ), .A3(_u10_n19236 ), .ZN(_u10_n19233 ) );
NOR4_X1 _u10_U7848  ( .A1(_u10_n19230 ), .A2(_u10_n19231 ), .A3(_u10_n19232 ), .A4(_u10_n19233 ), .ZN(_u10_n19208 ) );
NAND2_X1 _u10_U7847  ( .A1(1'b1), .A2(_u10_n11989 ), .ZN(_u10_n19226 ) );
NAND2_X1 _u10_U7846  ( .A1(1'b1), .A2(_u10_n11965 ), .ZN(_u10_n19227 ) );
NAND2_X1 _u10_U7845  ( .A1(1'b1), .A2(_u10_n11941 ), .ZN(_u10_n19228 ) );
NAND2_X1 _u10_U7844  ( .A1(1'b1), .A2(_u10_n11917 ), .ZN(_u10_n19229 ) );
NAND4_X1 _u10_U7843  ( .A1(_u10_n19226 ), .A2(_u10_n19227 ), .A3(_u10_n19228 ), .A4(_u10_n19229 ), .ZN(_u10_n19210 ) );
NAND2_X1 _u10_U7842  ( .A1(1'b1), .A2(_u10_n11893 ), .ZN(_u10_n19222 ) );
NAND2_X1 _u10_U7841  ( .A1(1'b1), .A2(_u10_n11869 ), .ZN(_u10_n19223 ) );
NAND2_X1 _u10_U7840  ( .A1(1'b1), .A2(_u10_n11845 ), .ZN(_u10_n19224 ) );
NAND2_X1 _u10_U7839  ( .A1(1'b1), .A2(_u10_n11821 ), .ZN(_u10_n19225 ) );
NAND4_X1 _u10_U7838  ( .A1(_u10_n19222 ), .A2(_u10_n19223 ), .A3(_u10_n19224 ), .A4(_u10_n19225 ), .ZN(_u10_n19211 ) );
NAND2_X1 _u10_U7837  ( .A1(1'b1), .A2(_u10_n11797 ), .ZN(_u10_n19218 ) );
NAND2_X1 _u10_U7836  ( .A1(1'b1), .A2(_u10_n11773 ), .ZN(_u10_n19219 ) );
NAND2_X1 _u10_U7835  ( .A1(1'b1), .A2(_u10_n11749 ), .ZN(_u10_n19220 ) );
NAND2_X1 _u10_U7834  ( .A1(1'b1), .A2(_u10_n11725 ), .ZN(_u10_n19221 ) );
NAND4_X1 _u10_U7833  ( .A1(_u10_n19218 ), .A2(_u10_n19219 ), .A3(_u10_n19220 ), .A4(_u10_n19221 ), .ZN(_u10_n19212 ) );
NAND2_X1 _u10_U7832  ( .A1(1'b1), .A2(_u10_n11701 ), .ZN(_u10_n19214 ) );
NAND2_X1 _u10_U7831  ( .A1(1'b1), .A2(_u10_n11677 ), .ZN(_u10_n19215 ) );
NAND2_X1 _u10_U7830  ( .A1(1'b1), .A2(_u10_n11653 ), .ZN(_u10_n19216 ) );
NAND2_X1 _u10_U7829  ( .A1(1'b1), .A2(_u10_n11629 ), .ZN(_u10_n19217 ) );
NAND4_X1 _u10_U7828  ( .A1(_u10_n19214 ), .A2(_u10_n19215 ), .A3(_u10_n19216 ), .A4(_u10_n19217 ), .ZN(_u10_n19213 ) );
NOR4_X1 _u10_U7827  ( .A1(_u10_n19210 ), .A2(_u10_n19211 ), .A3(_u10_n19212 ), .A4(_u10_n19213 ), .ZN(_u10_n19209 ) );
NAND2_X1 _u10_U7826  ( .A1(_u10_n19208 ), .A2(_u10_n19209 ), .ZN(am0[4]) );
NAND2_X1 _u10_U7825  ( .A1(1'b1), .A2(_u10_n12337 ), .ZN(_u10_n19204 ) );
NAND2_X1 _u10_U7824  ( .A1(1'b1), .A2(_u10_n12314 ), .ZN(_u10_n19205 ) );
NAND2_X1 _u10_U7823  ( .A1(1'b1), .A2(_u10_n12290 ), .ZN(_u10_n19206 ) );
NAND2_X1 _u10_U7822  ( .A1(1'b1), .A2(_u10_n12266 ), .ZN(_u10_n19207 ) );
NAND4_X1 _u10_U7821  ( .A1(_u10_n19204 ), .A2(_u10_n19205 ), .A3(_u10_n19206 ), .A4(_u10_n19207 ), .ZN(_u10_n19189 ) );
NAND2_X1 _u10_U7820  ( .A1(1'b1), .A2(_u10_n12241 ), .ZN(_u10_n19200 ) );
NAND2_X1 _u10_U7819  ( .A1(1'b1), .A2(_u10_n12217 ), .ZN(_u10_n19201 ) );
NAND2_X1 _u10_U7818  ( .A1(1'b1), .A2(_u10_n12194 ), .ZN(_u10_n19202 ) );
NAND2_X1 _u10_U7817  ( .A1(1'b1), .A2(_u10_n12169 ), .ZN(_u10_n19203 ) );
NAND4_X1 _u10_U7816  ( .A1(_u10_n19200 ), .A2(_u10_n19201 ), .A3(_u10_n19202 ), .A4(_u10_n19203 ), .ZN(_u10_n19190 ) );
NAND2_X1 _u10_U7815  ( .A1(1'b1), .A2(_u10_n12146 ), .ZN(_u10_n19196 ) );
NAND2_X1 _u10_U7814  ( .A1(1'b1), .A2(_u10_n12122 ), .ZN(_u10_n19197 ) );
NAND2_X1 _u10_U7813  ( .A1(1'b1), .A2(_u10_n12098 ), .ZN(_u10_n19198 ) );
NAND2_X1 _u10_U7812  ( .A1(1'b1), .A2(_u10_n12074 ), .ZN(_u10_n19199 ) );
NAND4_X1 _u10_U7811  ( .A1(_u10_n19196 ), .A2(_u10_n19197 ), .A3(_u10_n19198 ), .A4(_u10_n19199 ), .ZN(_u10_n19191 ) );
NAND2_X1 _u10_U7810  ( .A1(1'b1), .A2(_u10_n12050 ), .ZN(_u10_n19193 ) );
NAND2_X1 _u10_U7809  ( .A1(1'b1), .A2(_u10_n12026 ), .ZN(_u10_n19194 ) );
NAND2_X1 _u10_U7808  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19195 ) );
NAND3_X1 _u10_U7807  ( .A1(_u10_n19193 ), .A2(_u10_n19194 ), .A3(_u10_n19195 ), .ZN(_u10_n19192 ) );
NOR4_X1 _u10_U7806  ( .A1(_u10_n19189 ), .A2(_u10_n19190 ), .A3(_u10_n19191 ), .A4(_u10_n19192 ), .ZN(_u10_n19167 ) );
NAND2_X1 _u10_U7805  ( .A1(1'b1), .A2(_u10_n11989 ), .ZN(_u10_n19185 ) );
NAND2_X1 _u10_U7804  ( .A1(1'b1), .A2(_u10_n11965 ), .ZN(_u10_n19186 ) );
NAND2_X1 _u10_U7803  ( .A1(1'b1), .A2(_u10_n11941 ), .ZN(_u10_n19187 ) );
NAND2_X1 _u10_U7802  ( .A1(1'b1), .A2(_u10_n11917 ), .ZN(_u10_n19188 ) );
NAND4_X1 _u10_U7801  ( .A1(_u10_n19185 ), .A2(_u10_n19186 ), .A3(_u10_n19187 ), .A4(_u10_n19188 ), .ZN(_u10_n19169 ) );
NAND2_X1 _u10_U7800  ( .A1(1'b1), .A2(_u10_n11893 ), .ZN(_u10_n19181 ) );
NAND2_X1 _u10_U7799  ( .A1(1'b1), .A2(_u10_n11869 ), .ZN(_u10_n19182 ) );
NAND2_X1 _u10_U7798  ( .A1(1'b1), .A2(_u10_n11845 ), .ZN(_u10_n19183 ) );
NAND2_X1 _u10_U7797  ( .A1(1'b1), .A2(_u10_n11821 ), .ZN(_u10_n19184 ) );
NAND4_X1 _u10_U7796  ( .A1(_u10_n19181 ), .A2(_u10_n19182 ), .A3(_u10_n19183 ), .A4(_u10_n19184 ), .ZN(_u10_n19170 ) );
NAND2_X1 _u10_U7795  ( .A1(1'b1), .A2(_u10_n11797 ), .ZN(_u10_n19177 ) );
NAND2_X1 _u10_U7794  ( .A1(1'b1), .A2(_u10_n11773 ), .ZN(_u10_n19178 ) );
NAND2_X1 _u10_U7793  ( .A1(1'b1), .A2(_u10_n11749 ), .ZN(_u10_n19179 ) );
NAND2_X1 _u10_U7792  ( .A1(1'b1), .A2(_u10_n11725 ), .ZN(_u10_n19180 ) );
NAND4_X1 _u10_U7791  ( .A1(_u10_n19177 ), .A2(_u10_n19178 ), .A3(_u10_n19179 ), .A4(_u10_n19180 ), .ZN(_u10_n19171 ) );
NAND2_X1 _u10_U7790  ( .A1(1'b1), .A2(_u10_n11701 ), .ZN(_u10_n19173 ) );
NAND2_X1 _u10_U7789  ( .A1(1'b1), .A2(_u10_n11677 ), .ZN(_u10_n19174 ) );
NAND2_X1 _u10_U7788  ( .A1(1'b1), .A2(_u10_n11653 ), .ZN(_u10_n19175 ) );
NAND2_X1 _u10_U7787  ( .A1(1'b1), .A2(_u10_n11629 ), .ZN(_u10_n19176 ) );
NAND4_X1 _u10_U7786  ( .A1(_u10_n19173 ), .A2(_u10_n19174 ), .A3(_u10_n19175 ), .A4(_u10_n19176 ), .ZN(_u10_n19172 ) );
NOR4_X1 _u10_U7785  ( .A1(_u10_n19169 ), .A2(_u10_n19170 ), .A3(_u10_n19171 ), .A4(_u10_n19172 ), .ZN(_u10_n19168 ) );
NAND2_X1 _u10_U7784  ( .A1(_u10_n19167 ), .A2(_u10_n19168 ), .ZN(am0[5]) );
NAND2_X1 _u10_U7783  ( .A1(1'b1), .A2(_u10_n12337 ), .ZN(_u10_n19163 ) );
NAND2_X1 _u10_U7782  ( .A1(1'b1), .A2(_u10_n12314 ), .ZN(_u10_n19164 ) );
NAND2_X1 _u10_U7781  ( .A1(1'b1), .A2(_u10_n12290 ), .ZN(_u10_n19165 ) );
NAND2_X1 _u10_U7780  ( .A1(1'b1), .A2(_u10_n12266 ), .ZN(_u10_n19166 ) );
NAND4_X1 _u10_U7779  ( .A1(_u10_n19163 ), .A2(_u10_n19164 ), .A3(_u10_n19165 ), .A4(_u10_n19166 ), .ZN(_u10_n19148 ) );
NAND2_X1 _u10_U7778  ( .A1(1'b1), .A2(_u10_n12241 ), .ZN(_u10_n19159 ) );
NAND2_X1 _u10_U7777  ( .A1(1'b1), .A2(_u10_n12217 ), .ZN(_u10_n19160 ) );
NAND2_X1 _u10_U7776  ( .A1(1'b1), .A2(_u10_n12194 ), .ZN(_u10_n19161 ) );
NAND2_X1 _u10_U7775  ( .A1(1'b1), .A2(_u10_n12169 ), .ZN(_u10_n19162 ) );
NAND4_X1 _u10_U7774  ( .A1(_u10_n19159 ), .A2(_u10_n19160 ), .A3(_u10_n19161 ), .A4(_u10_n19162 ), .ZN(_u10_n19149 ) );
NAND2_X1 _u10_U7773  ( .A1(1'b1), .A2(_u10_n12146 ), .ZN(_u10_n19155 ) );
NAND2_X1 _u10_U7772  ( .A1(1'b1), .A2(_u10_n12122 ), .ZN(_u10_n19156 ) );
NAND2_X1 _u10_U7771  ( .A1(1'b1), .A2(_u10_n12098 ), .ZN(_u10_n19157 ) );
NAND2_X1 _u10_U7770  ( .A1(1'b1), .A2(_u10_n12074 ), .ZN(_u10_n19158 ) );
NAND4_X1 _u10_U7769  ( .A1(_u10_n19155 ), .A2(_u10_n19156 ), .A3(_u10_n19157 ), .A4(_u10_n19158 ), .ZN(_u10_n19150 ) );
NAND2_X1 _u10_U7768  ( .A1(1'b1), .A2(_u10_n12050 ), .ZN(_u10_n19152 ) );
NAND2_X1 _u10_U7767  ( .A1(1'b1), .A2(_u10_n12026 ), .ZN(_u10_n19153 ) );
NAND2_X1 _u10_U7766  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19154 ) );
NAND3_X1 _u10_U7765  ( .A1(_u10_n19152 ), .A2(_u10_n19153 ), .A3(_u10_n19154 ), .ZN(_u10_n19151 ) );
NOR4_X1 _u10_U7764  ( .A1(_u10_n19148 ), .A2(_u10_n19149 ), .A3(_u10_n19150 ), .A4(_u10_n19151 ), .ZN(_u10_n19126 ) );
NAND2_X1 _u10_U7763  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n19144 ) );
NAND2_X1 _u10_U7762  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n19145 ) );
NAND2_X1 _u10_U7761  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n19146 ) );
NAND2_X1 _u10_U7760  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n19147 ) );
NAND4_X1 _u10_U7759  ( .A1(_u10_n19144 ), .A2(_u10_n19145 ), .A3(_u10_n19146 ), .A4(_u10_n19147 ), .ZN(_u10_n19128 ) );
NAND2_X1 _u10_U7758  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n19140 ) );
NAND2_X1 _u10_U7757  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n19141 ) );
NAND2_X1 _u10_U7756  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n19142 ) );
NAND2_X1 _u10_U7755  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n19143 ) );
NAND4_X1 _u10_U7754  ( .A1(_u10_n19140 ), .A2(_u10_n19141 ), .A3(_u10_n19142 ), .A4(_u10_n19143 ), .ZN(_u10_n19129 ) );
NAND2_X1 _u10_U7753  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n19136 ) );
NAND2_X1 _u10_U7752  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n19137 ) );
NAND2_X1 _u10_U7751  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n19138 ) );
NAND2_X1 _u10_U7750  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n19139 ) );
NAND4_X1 _u10_U7749  ( .A1(_u10_n19136 ), .A2(_u10_n19137 ), .A3(_u10_n19138 ), .A4(_u10_n19139 ), .ZN(_u10_n19130 ) );
NAND2_X1 _u10_U7748  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n19132 ) );
NAND2_X1 _u10_U7747  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n19133 ) );
NAND2_X1 _u10_U7746  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n19134 ) );
NAND2_X1 _u10_U7745  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n19135 ) );
NAND4_X1 _u10_U7744  ( .A1(_u10_n19132 ), .A2(_u10_n19133 ), .A3(_u10_n19134 ), .A4(_u10_n19135 ), .ZN(_u10_n19131 ) );
NOR4_X1 _u10_U7743  ( .A1(_u10_n19128 ), .A2(_u10_n19129 ), .A3(_u10_n19130 ), .A4(_u10_n19131 ), .ZN(_u10_n19127 ) );
NAND2_X1 _u10_U7742  ( .A1(_u10_n19126 ), .A2(_u10_n19127 ), .ZN(am0[6]) );
NAND2_X1 _u10_U7741  ( .A1(1'b1), .A2(_u10_n12337 ), .ZN(_u10_n19122 ) );
NAND2_X1 _u10_U7740  ( .A1(1'b1), .A2(_u10_n12314 ), .ZN(_u10_n19123 ) );
NAND2_X1 _u10_U7739  ( .A1(1'b1), .A2(_u10_n12290 ), .ZN(_u10_n19124 ) );
NAND2_X1 _u10_U7738  ( .A1(1'b1), .A2(_u10_n12266 ), .ZN(_u10_n19125 ) );
NAND4_X1 _u10_U7737  ( .A1(_u10_n19122 ), .A2(_u10_n19123 ), .A3(_u10_n19124 ), .A4(_u10_n19125 ), .ZN(_u10_n19107 ) );
NAND2_X1 _u10_U7736  ( .A1(1'b1), .A2(_u10_n12241 ), .ZN(_u10_n19118 ) );
NAND2_X1 _u10_U7735  ( .A1(1'b1), .A2(_u10_n12217 ), .ZN(_u10_n19119 ) );
NAND2_X1 _u10_U7734  ( .A1(1'b1), .A2(_u10_n12194 ), .ZN(_u10_n19120 ) );
NAND2_X1 _u10_U7733  ( .A1(1'b1), .A2(_u10_n12169 ), .ZN(_u10_n19121 ) );
NAND4_X1 _u10_U7732  ( .A1(_u10_n19118 ), .A2(_u10_n19119 ), .A3(_u10_n19120 ), .A4(_u10_n19121 ), .ZN(_u10_n19108 ) );
NAND2_X1 _u10_U7731  ( .A1(1'b1), .A2(_u10_n12146 ), .ZN(_u10_n19114 ) );
NAND2_X1 _u10_U7730  ( .A1(1'b1), .A2(_u10_n12122 ), .ZN(_u10_n19115 ) );
NAND2_X1 _u10_U7729  ( .A1(1'b1), .A2(_u10_n12098 ), .ZN(_u10_n19116 ) );
NAND2_X1 _u10_U7728  ( .A1(1'b1), .A2(_u10_n12074 ), .ZN(_u10_n19117 ) );
NAND4_X1 _u10_U7727  ( .A1(_u10_n19114 ), .A2(_u10_n19115 ), .A3(_u10_n19116 ), .A4(_u10_n19117 ), .ZN(_u10_n19109 ) );
NAND2_X1 _u10_U7726  ( .A1(1'b1), .A2(_u10_n12050 ), .ZN(_u10_n19111 ) );
NAND2_X1 _u10_U7725  ( .A1(1'b1), .A2(_u10_n12026 ), .ZN(_u10_n19112 ) );
NAND2_X1 _u10_U7724  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19113 ) );
NAND3_X1 _u10_U7723  ( .A1(_u10_n19111 ), .A2(_u10_n19112 ), .A3(_u10_n19113 ), .ZN(_u10_n19110 ) );
NOR4_X1 _u10_U7722  ( .A1(_u10_n19107 ), .A2(_u10_n19108 ), .A3(_u10_n19109 ), .A4(_u10_n19110 ), .ZN(_u10_n19085 ) );
NAND2_X1 _u10_U7721  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n19103 ) );
NAND2_X1 _u10_U7720  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n19104 ) );
NAND2_X1 _u10_U7719  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n19105 ) );
NAND2_X1 _u10_U7718  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n19106 ) );
NAND4_X1 _u10_U7717  ( .A1(_u10_n19103 ), .A2(_u10_n19104 ), .A3(_u10_n19105 ), .A4(_u10_n19106 ), .ZN(_u10_n19087 ) );
NAND2_X1 _u10_U7716  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n19099 ) );
NAND2_X1 _u10_U7715  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n19100 ) );
NAND2_X1 _u10_U7714  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n19101 ) );
NAND2_X1 _u10_U7713  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n19102 ) );
NAND4_X1 _u10_U7712  ( .A1(_u10_n19099 ), .A2(_u10_n19100 ), .A3(_u10_n19101 ), .A4(_u10_n19102 ), .ZN(_u10_n19088 ) );
NAND2_X1 _u10_U7711  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n19095 ) );
NAND2_X1 _u10_U7710  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n19096 ) );
NAND2_X1 _u10_U7709  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n19097 ) );
NAND2_X1 _u10_U7708  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n19098 ) );
NAND4_X1 _u10_U7707  ( .A1(_u10_n19095 ), .A2(_u10_n19096 ), .A3(_u10_n19097 ), .A4(_u10_n19098 ), .ZN(_u10_n19089 ) );
NAND2_X1 _u10_U7706  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n19091 ) );
NAND2_X1 _u10_U7705  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n19092 ) );
NAND2_X1 _u10_U7704  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n19093 ) );
NAND2_X1 _u10_U7703  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n19094 ) );
NAND4_X1 _u10_U7702  ( .A1(_u10_n19091 ), .A2(_u10_n19092 ), .A3(_u10_n19093 ), .A4(_u10_n19094 ), .ZN(_u10_n19090 ) );
NOR4_X1 _u10_U7701  ( .A1(_u10_n19087 ), .A2(_u10_n19088 ), .A3(_u10_n19089 ), .A4(_u10_n19090 ), .ZN(_u10_n19086 ) );
NAND2_X1 _u10_U7700  ( .A1(_u10_n19085 ), .A2(_u10_n19086 ), .ZN(am0[7]) );
NAND2_X1 _u10_U7699  ( .A1(1'b1), .A2(_u10_n12337 ), .ZN(_u10_n19081 ) );
NAND2_X1 _u10_U7698  ( .A1(1'b1), .A2(_u10_n12314 ), .ZN(_u10_n19082 ) );
NAND2_X1 _u10_U7697  ( .A1(1'b1), .A2(_u10_n12290 ), .ZN(_u10_n19083 ) );
NAND2_X1 _u10_U7696  ( .A1(1'b1), .A2(_u10_n12266 ), .ZN(_u10_n19084 ) );
NAND4_X1 _u10_U7695  ( .A1(_u10_n19081 ), .A2(_u10_n19082 ), .A3(_u10_n19083 ), .A4(_u10_n19084 ), .ZN(_u10_n19066 ) );
NAND2_X1 _u10_U7694  ( .A1(1'b1), .A2(_u10_n12241 ), .ZN(_u10_n19077 ) );
NAND2_X1 _u10_U7693  ( .A1(1'b1), .A2(_u10_n12217 ), .ZN(_u10_n19078 ) );
NAND2_X1 _u10_U7692  ( .A1(1'b1), .A2(_u10_n12194 ), .ZN(_u10_n19079 ) );
NAND2_X1 _u10_U7691  ( .A1(1'b1), .A2(_u10_n12169 ), .ZN(_u10_n19080 ) );
NAND4_X1 _u10_U7690  ( .A1(_u10_n19077 ), .A2(_u10_n19078 ), .A3(_u10_n19079 ), .A4(_u10_n19080 ), .ZN(_u10_n19067 ) );
NAND2_X1 _u10_U7689  ( .A1(1'b1), .A2(_u10_n12146 ), .ZN(_u10_n19073 ) );
NAND2_X1 _u10_U7688  ( .A1(1'b1), .A2(_u10_n12122 ), .ZN(_u10_n19074 ) );
NAND2_X1 _u10_U7687  ( .A1(1'b1), .A2(_u10_n12098 ), .ZN(_u10_n19075 ) );
NAND2_X1 _u10_U7686  ( .A1(1'b1), .A2(_u10_n12074 ), .ZN(_u10_n19076 ) );
NAND4_X1 _u10_U7685  ( .A1(_u10_n19073 ), .A2(_u10_n19074 ), .A3(_u10_n19075 ), .A4(_u10_n19076 ), .ZN(_u10_n19068 ) );
NAND2_X1 _u10_U7684  ( .A1(1'b1), .A2(_u10_n12050 ), .ZN(_u10_n19070 ) );
NAND2_X1 _u10_U7683  ( .A1(1'b1), .A2(_u10_n12026 ), .ZN(_u10_n19071 ) );
NAND2_X1 _u10_U7682  ( .A1(1'b1), .A2(_u10_n12006 ), .ZN(_u10_n19072 ) );
NAND3_X1 _u10_U7681  ( .A1(_u10_n19070 ), .A2(_u10_n19071 ), .A3(_u10_n19072 ), .ZN(_u10_n19069 ) );
NOR4_X1 _u10_U7680  ( .A1(_u10_n19066 ), .A2(_u10_n19067 ), .A3(_u10_n19068 ), .A4(_u10_n19069 ), .ZN(_u10_n19044 ) );
NAND2_X1 _u10_U7679  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n19062 ) );
NAND2_X1 _u10_U7678  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n19063 ) );
NAND2_X1 _u10_U7677  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n19064 ) );
NAND2_X1 _u10_U7676  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n19065 ) );
NAND4_X1 _u10_U7675  ( .A1(_u10_n19062 ), .A2(_u10_n19063 ), .A3(_u10_n19064 ), .A4(_u10_n19065 ), .ZN(_u10_n19046 ) );
NAND2_X1 _u10_U7674  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n19058 ) );
NAND2_X1 _u10_U7673  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n19059 ) );
NAND2_X1 _u10_U7672  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n19060 ) );
NAND2_X1 _u10_U7671  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n19061 ) );
NAND4_X1 _u10_U7670  ( .A1(_u10_n19058 ), .A2(_u10_n19059 ), .A3(_u10_n19060 ), .A4(_u10_n19061 ), .ZN(_u10_n19047 ) );
NAND2_X1 _u10_U7669  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n19054 ) );
NAND2_X1 _u10_U7668  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n19055 ) );
NAND2_X1 _u10_U7667  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n19056 ) );
NAND2_X1 _u10_U7666  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n19057 ) );
NAND4_X1 _u10_U7665  ( .A1(_u10_n19054 ), .A2(_u10_n19055 ), .A3(_u10_n19056 ), .A4(_u10_n19057 ), .ZN(_u10_n19048 ) );
NAND2_X1 _u10_U7664  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n19050 ) );
NAND2_X1 _u10_U7663  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n19051 ) );
NAND2_X1 _u10_U7662  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n19052 ) );
NAND2_X1 _u10_U7661  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n19053 ) );
NAND4_X1 _u10_U7660  ( .A1(_u10_n19050 ), .A2(_u10_n19051 ), .A3(_u10_n19052 ), .A4(_u10_n19053 ), .ZN(_u10_n19049 ) );
NOR4_X1 _u10_U7659  ( .A1(_u10_n19046 ), .A2(_u10_n19047 ), .A3(_u10_n19048 ), .A4(_u10_n19049 ), .ZN(_u10_n19045 ) );
NAND2_X1 _u10_U7658  ( .A1(_u10_n19044 ), .A2(_u10_n19045 ), .ZN(am0[8]) );
NAND2_X1 _u10_U7657  ( .A1(1'b1), .A2(_u10_n12337 ), .ZN(_u10_n19040 ) );
NAND2_X1 _u10_U7656  ( .A1(1'b1), .A2(_u10_n12314 ), .ZN(_u10_n19041 ) );
NAND2_X1 _u10_U7655  ( .A1(1'b1), .A2(_u10_n12290 ), .ZN(_u10_n19042 ) );
NAND2_X1 _u10_U7654  ( .A1(1'b1), .A2(_u10_n12266 ), .ZN(_u10_n19043 ) );
NAND4_X1 _u10_U7653  ( .A1(_u10_n19040 ), .A2(_u10_n19041 ), .A3(_u10_n19042 ), .A4(_u10_n19043 ), .ZN(_u10_n19025 ) );
NAND2_X1 _u10_U7652  ( .A1(1'b1), .A2(_u10_n12241 ), .ZN(_u10_n19036 ) );
NAND2_X1 _u10_U7651  ( .A1(1'b1), .A2(_u10_n12217 ), .ZN(_u10_n19037 ) );
NAND2_X1 _u10_U7650  ( .A1(1'b1), .A2(_u10_n12194 ), .ZN(_u10_n19038 ) );
NAND2_X1 _u10_U7649  ( .A1(1'b1), .A2(_u10_n12169 ), .ZN(_u10_n19039 ) );
NAND4_X1 _u10_U7648  ( .A1(_u10_n19036 ), .A2(_u10_n19037 ), .A3(_u10_n19038 ), .A4(_u10_n19039 ), .ZN(_u10_n19026 ) );
NAND2_X1 _u10_U7647  ( .A1(1'b1), .A2(_u10_n12146 ), .ZN(_u10_n19032 ) );
NAND2_X1 _u10_U7646  ( .A1(1'b1), .A2(_u10_n12122 ), .ZN(_u10_n19033 ) );
NAND2_X1 _u10_U7645  ( .A1(1'b1), .A2(_u10_n12098 ), .ZN(_u10_n19034 ) );
NAND2_X1 _u10_U7644  ( .A1(1'b1), .A2(_u10_n12074 ), .ZN(_u10_n19035 ) );
NAND4_X1 _u10_U7643  ( .A1(_u10_n19032 ), .A2(_u10_n19033 ), .A3(_u10_n19034 ), .A4(_u10_n19035 ), .ZN(_u10_n19027 ) );
NAND2_X1 _u10_U7642  ( .A1(1'b1), .A2(_u10_n12050 ), .ZN(_u10_n19029 ) );
NAND2_X1 _u10_U7641  ( .A1(1'b1), .A2(_u10_n12026 ), .ZN(_u10_n19030 ) );
NAND2_X1 _u10_U7640  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n19031 ) );
NAND3_X1 _u10_U7639  ( .A1(_u10_n19029 ), .A2(_u10_n19030 ), .A3(_u10_n19031 ), .ZN(_u10_n19028 ) );
NOR4_X1 _u10_U7638  ( .A1(_u10_n19025 ), .A2(_u10_n19026 ), .A3(_u10_n19027 ), .A4(_u10_n19028 ), .ZN(_u10_n19003 ) );
NAND2_X1 _u10_U7637  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n19021 ) );
NAND2_X1 _u10_U7636  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n19022 ) );
NAND2_X1 _u10_U7635  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n19023 ) );
NAND2_X1 _u10_U7634  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n19024 ) );
NAND4_X1 _u10_U7633  ( .A1(_u10_n19021 ), .A2(_u10_n19022 ), .A3(_u10_n19023 ), .A4(_u10_n19024 ), .ZN(_u10_n19005 ) );
NAND2_X1 _u10_U7632  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n19017 ) );
NAND2_X1 _u10_U7631  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n19018 ) );
NAND2_X1 _u10_U7630  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n19019 ) );
NAND2_X1 _u10_U7629  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n19020 ) );
NAND4_X1 _u10_U7628  ( .A1(_u10_n19017 ), .A2(_u10_n19018 ), .A3(_u10_n19019 ), .A4(_u10_n19020 ), .ZN(_u10_n19006 ) );
NAND2_X1 _u10_U7627  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n19013 ) );
NAND2_X1 _u10_U7626  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n19014 ) );
NAND2_X1 _u10_U7625  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n19015 ) );
NAND2_X1 _u10_U7624  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n19016 ) );
NAND4_X1 _u10_U7623  ( .A1(_u10_n19013 ), .A2(_u10_n19014 ), .A3(_u10_n19015 ), .A4(_u10_n19016 ), .ZN(_u10_n19007 ) );
NAND2_X1 _u10_U7622  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n19009 ) );
NAND2_X1 _u10_U7621  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n19010 ) );
NAND2_X1 _u10_U7620  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n19011 ) );
NAND2_X1 _u10_U7619  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n19012 ) );
NAND4_X1 _u10_U7618  ( .A1(_u10_n19009 ), .A2(_u10_n19010 ), .A3(_u10_n19011 ), .A4(_u10_n19012 ), .ZN(_u10_n19008 ) );
NOR4_X1 _u10_U7617  ( .A1(_u10_n19005 ), .A2(_u10_n19006 ), .A3(_u10_n19007 ), .A4(_u10_n19008 ), .ZN(_u10_n19004 ) );
NAND2_X1 _u10_U7616  ( .A1(_u10_n19003 ), .A2(_u10_n19004 ), .ZN(am0[9]) );
NAND2_X1 _u10_U7615  ( .A1(1'b0), .A2(_u10_n12337 ), .ZN(_u10_n18999 ) );
NAND2_X1 _u10_U7614  ( .A1(1'b0), .A2(_u10_n12314 ), .ZN(_u10_n19000 ) );
NAND2_X1 _u10_U7613  ( .A1(1'b0), .A2(_u10_n12290 ), .ZN(_u10_n19001 ) );
NAND2_X1 _u10_U7612  ( .A1(1'b0), .A2(_u10_n12266 ), .ZN(_u10_n19002 ) );
NAND4_X1 _u10_U7611  ( .A1(_u10_n18999 ), .A2(_u10_n19000 ), .A3(_u10_n19001 ), .A4(_u10_n19002 ), .ZN(_u10_n18984 ) );
NAND2_X1 _u10_U7610  ( .A1(1'b0), .A2(_u10_n12241 ), .ZN(_u10_n18995 ) );
NAND2_X1 _u10_U7609  ( .A1(1'b0), .A2(_u10_n12217 ), .ZN(_u10_n18996 ) );
NAND2_X1 _u10_U7608  ( .A1(1'b0), .A2(_u10_n12194 ), .ZN(_u10_n18997 ) );
NAND2_X1 _u10_U7607  ( .A1(1'b0), .A2(_u10_n12169 ), .ZN(_u10_n18998 ) );
NAND4_X1 _u10_U7606  ( .A1(_u10_n18995 ), .A2(_u10_n18996 ), .A3(_u10_n18997 ), .A4(_u10_n18998 ), .ZN(_u10_n18985 ) );
NAND2_X1 _u10_U7605  ( .A1(1'b0), .A2(_u10_n12146 ), .ZN(_u10_n18991 ) );
NAND2_X1 _u10_U7604  ( .A1(1'b0), .A2(_u10_n12122 ), .ZN(_u10_n18992 ) );
NAND2_X1 _u10_U7603  ( .A1(1'b0), .A2(_u10_n12098 ), .ZN(_u10_n18993 ) );
NAND2_X1 _u10_U7602  ( .A1(1'b0), .A2(_u10_n12074 ), .ZN(_u10_n18994 ) );
NAND4_X1 _u10_U7601  ( .A1(_u10_n18991 ), .A2(_u10_n18992 ), .A3(_u10_n18993 ), .A4(_u10_n18994 ), .ZN(_u10_n18986 ) );
NAND2_X1 _u10_U7600  ( .A1(1'b0), .A2(_u10_n12050 ), .ZN(_u10_n18988 ) );
NAND2_X1 _u10_U7599  ( .A1(1'b0), .A2(_u10_n12026 ), .ZN(_u10_n18989 ) );
NAND2_X1 _u10_U7598  ( .A1(1'b0), .A2(_u10_n12007 ), .ZN(_u10_n18990 ) );
NAND3_X1 _u10_U7597  ( .A1(_u10_n18988 ), .A2(_u10_n18989 ), .A3(_u10_n18990 ), .ZN(_u10_n18987 ) );
NOR4_X1 _u10_U7596  ( .A1(_u10_n18984 ), .A2(_u10_n18985 ), .A3(_u10_n18986 ), .A4(_u10_n18987 ), .ZN(_u10_n18962 ) );
NAND2_X1 _u10_U7595  ( .A1(1'b0), .A2(_u10_n11990 ), .ZN(_u10_n18980 ) );
NAND2_X1 _u10_U7594  ( .A1(1'b0), .A2(_u10_n11966 ), .ZN(_u10_n18981 ) );
NAND2_X1 _u10_U7593  ( .A1(1'b0), .A2(_u10_n11942 ), .ZN(_u10_n18982 ) );
NAND2_X1 _u10_U7592  ( .A1(1'b0), .A2(_u10_n11918 ), .ZN(_u10_n18983 ) );
NAND4_X1 _u10_U7591  ( .A1(_u10_n18980 ), .A2(_u10_n18981 ), .A3(_u10_n18982 ), .A4(_u10_n18983 ), .ZN(_u10_n18964 ) );
NAND2_X1 _u10_U7590  ( .A1(1'b0), .A2(_u10_n11894 ), .ZN(_u10_n18976 ) );
NAND2_X1 _u10_U7589  ( .A1(1'b0), .A2(_u10_n11870 ), .ZN(_u10_n18977 ) );
NAND2_X1 _u10_U7588  ( .A1(1'b0), .A2(_u10_n11846 ), .ZN(_u10_n18978 ) );
NAND2_X1 _u10_U7587  ( .A1(1'b0), .A2(_u10_n11822 ), .ZN(_u10_n18979 ) );
NAND4_X1 _u10_U7586  ( .A1(_u10_n18976 ), .A2(_u10_n18977 ), .A3(_u10_n18978 ), .A4(_u10_n18979 ), .ZN(_u10_n18965 ) );
NAND2_X1 _u10_U7585  ( .A1(1'b0), .A2(_u10_n11798 ), .ZN(_u10_n18972 ) );
NAND2_X1 _u10_U7584  ( .A1(1'b0), .A2(_u10_n11774 ), .ZN(_u10_n18973 ) );
NAND2_X1 _u10_U7583  ( .A1(1'b0), .A2(_u10_n11750 ), .ZN(_u10_n18974 ) );
NAND2_X1 _u10_U7582  ( .A1(1'b0), .A2(_u10_n11726 ), .ZN(_u10_n18975 ) );
NAND4_X1 _u10_U7581  ( .A1(_u10_n18972 ), .A2(_u10_n18973 ), .A3(_u10_n18974 ), .A4(_u10_n18975 ), .ZN(_u10_n18966 ) );
NAND2_X1 _u10_U7580  ( .A1(1'b0), .A2(_u10_n11702 ), .ZN(_u10_n18968 ) );
NAND2_X1 _u10_U7579  ( .A1(1'b0), .A2(_u10_n11678 ), .ZN(_u10_n18969 ) );
NAND2_X1 _u10_U7578  ( .A1(1'b0), .A2(_u10_n11654 ), .ZN(_u10_n18970 ) );
NAND2_X1 _u10_U7577  ( .A1(1'b0), .A2(_u10_n11630 ), .ZN(_u10_n18971 ) );
NAND4_X1 _u10_U7576  ( .A1(_u10_n18968 ), .A2(_u10_n18969 ), .A3(_u10_n18970 ), .A4(_u10_n18971 ), .ZN(_u10_n18967 ) );
NOR4_X1 _u10_U7575  ( .A1(_u10_n18964 ), .A2(_u10_n18965 ), .A3(_u10_n18966 ), .A4(_u10_n18967 ), .ZN(_u10_n18963 ) );
NAND2_X1 _u10_U7574  ( .A1(_u10_n18962 ), .A2(_u10_n18963 ), .ZN(am1[0]) );
NAND2_X1 _u10_U7573  ( .A1(1'b1), .A2(_u10_n12337 ), .ZN(_u10_n18958 ) );
NAND2_X1 _u10_U7572  ( .A1(1'b1), .A2(_u10_n12314 ), .ZN(_u10_n18959 ) );
NAND2_X1 _u10_U7571  ( .A1(1'b1), .A2(_u10_n12290 ), .ZN(_u10_n18960 ) );
NAND2_X1 _u10_U7570  ( .A1(1'b1), .A2(_u10_n12266 ), .ZN(_u10_n18961 ) );
NAND4_X1 _u10_U7569  ( .A1(_u10_n18958 ), .A2(_u10_n18959 ), .A3(_u10_n18960 ), .A4(_u10_n18961 ), .ZN(_u10_n18943 ) );
NAND2_X1 _u10_U7568  ( .A1(1'b1), .A2(_u10_n12241 ), .ZN(_u10_n18954 ) );
NAND2_X1 _u10_U7567  ( .A1(1'b1), .A2(_u10_n12217 ), .ZN(_u10_n18955 ) );
NAND2_X1 _u10_U7566  ( .A1(1'b1), .A2(_u10_n12194 ), .ZN(_u10_n18956 ) );
NAND2_X1 _u10_U7565  ( .A1(1'b1), .A2(_u10_n12169 ), .ZN(_u10_n18957 ) );
NAND4_X1 _u10_U7564  ( .A1(_u10_n18954 ), .A2(_u10_n18955 ), .A3(_u10_n18956 ), .A4(_u10_n18957 ), .ZN(_u10_n18944 ) );
NAND2_X1 _u10_U7563  ( .A1(1'b1), .A2(_u10_n12146 ), .ZN(_u10_n18950 ) );
NAND2_X1 _u10_U7562  ( .A1(1'b1), .A2(_u10_n12122 ), .ZN(_u10_n18951 ) );
NAND2_X1 _u10_U7561  ( .A1(1'b1), .A2(_u10_n12098 ), .ZN(_u10_n18952 ) );
NAND2_X1 _u10_U7560  ( .A1(1'b1), .A2(_u10_n12074 ), .ZN(_u10_n18953 ) );
NAND4_X1 _u10_U7559  ( .A1(_u10_n18950 ), .A2(_u10_n18951 ), .A3(_u10_n18952 ), .A4(_u10_n18953 ), .ZN(_u10_n18945 ) );
NAND2_X1 _u10_U7558  ( .A1(1'b1), .A2(_u10_n12050 ), .ZN(_u10_n18947 ) );
NAND2_X1 _u10_U7557  ( .A1(1'b1), .A2(_u10_n12026 ), .ZN(_u10_n18948 ) );
NAND2_X1 _u10_U7556  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18949 ) );
NAND3_X1 _u10_U7555  ( .A1(_u10_n18947 ), .A2(_u10_n18948 ), .A3(_u10_n18949 ), .ZN(_u10_n18946 ) );
NOR4_X1 _u10_U7554  ( .A1(_u10_n18943 ), .A2(_u10_n18944 ), .A3(_u10_n18945 ), .A4(_u10_n18946 ), .ZN(_u10_n18921 ) );
NAND2_X1 _u10_U7553  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n18939 ) );
NAND2_X1 _u10_U7552  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n18940 ) );
NAND2_X1 _u10_U7551  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n18941 ) );
NAND2_X1 _u10_U7550  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n18942 ) );
NAND4_X1 _u10_U7549  ( .A1(_u10_n18939 ), .A2(_u10_n18940 ), .A3(_u10_n18941 ), .A4(_u10_n18942 ), .ZN(_u10_n18923 ) );
NAND2_X1 _u10_U7548  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n18935 ) );
NAND2_X1 _u10_U7547  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n18936 ) );
NAND2_X1 _u10_U7546  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n18937 ) );
NAND2_X1 _u10_U7545  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n18938 ) );
NAND4_X1 _u10_U7544  ( .A1(_u10_n18935 ), .A2(_u10_n18936 ), .A3(_u10_n18937 ), .A4(_u10_n18938 ), .ZN(_u10_n18924 ) );
NAND2_X1 _u10_U7543  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n18931 ) );
NAND2_X1 _u10_U7542  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n18932 ) );
NAND2_X1 _u10_U7541  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n18933 ) );
NAND2_X1 _u10_U7540  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n18934 ) );
NAND4_X1 _u10_U7539  ( .A1(_u10_n18931 ), .A2(_u10_n18932 ), .A3(_u10_n18933 ), .A4(_u10_n18934 ), .ZN(_u10_n18925 ) );
NAND2_X1 _u10_U7538  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n18927 ) );
NAND2_X1 _u10_U7537  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n18928 ) );
NAND2_X1 _u10_U7536  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n18929 ) );
NAND2_X1 _u10_U7535  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n18930 ) );
NAND4_X1 _u10_U7534  ( .A1(_u10_n18927 ), .A2(_u10_n18928 ), .A3(_u10_n18929 ), .A4(_u10_n18930 ), .ZN(_u10_n18926 ) );
NOR4_X1 _u10_U7533  ( .A1(_u10_n18923 ), .A2(_u10_n18924 ), .A3(_u10_n18925 ), .A4(_u10_n18926 ), .ZN(_u10_n18922 ) );
NAND2_X1 _u10_U7532  ( .A1(_u10_n18921 ), .A2(_u10_n18922 ), .ZN(am1[10]) );
NAND2_X1 _u10_U7531  ( .A1(1'b1), .A2(_u10_n12337 ), .ZN(_u10_n18917 ) );
NAND2_X1 _u10_U7530  ( .A1(1'b1), .A2(_u10_n12314 ), .ZN(_u10_n18918 ) );
NAND2_X1 _u10_U7529  ( .A1(1'b1), .A2(_u10_n12290 ), .ZN(_u10_n18919 ) );
NAND2_X1 _u10_U7528  ( .A1(1'b1), .A2(_u10_n12266 ), .ZN(_u10_n18920 ) );
NAND4_X1 _u10_U7527  ( .A1(_u10_n18917 ), .A2(_u10_n18918 ), .A3(_u10_n18919 ), .A4(_u10_n18920 ), .ZN(_u10_n18902 ) );
NAND2_X1 _u10_U7526  ( .A1(1'b1), .A2(_u10_n12241 ), .ZN(_u10_n18913 ) );
NAND2_X1 _u10_U7525  ( .A1(1'b1), .A2(_u10_n12217 ), .ZN(_u10_n18914 ) );
NAND2_X1 _u10_U7524  ( .A1(1'b1), .A2(_u10_n12194 ), .ZN(_u10_n18915 ) );
NAND2_X1 _u10_U7523  ( .A1(1'b1), .A2(_u10_n12169 ), .ZN(_u10_n18916 ) );
NAND4_X1 _u10_U7522  ( .A1(_u10_n18913 ), .A2(_u10_n18914 ), .A3(_u10_n18915 ), .A4(_u10_n18916 ), .ZN(_u10_n18903 ) );
NAND2_X1 _u10_U7521  ( .A1(1'b1), .A2(_u10_n12146 ), .ZN(_u10_n18909 ) );
NAND2_X1 _u10_U7520  ( .A1(1'b1), .A2(_u10_n12122 ), .ZN(_u10_n18910 ) );
NAND2_X1 _u10_U7519  ( .A1(1'b1), .A2(_u10_n12098 ), .ZN(_u10_n18911 ) );
NAND2_X1 _u10_U7518  ( .A1(1'b1), .A2(_u10_n12074 ), .ZN(_u10_n18912 ) );
NAND4_X1 _u10_U7517  ( .A1(_u10_n18909 ), .A2(_u10_n18910 ), .A3(_u10_n18911 ), .A4(_u10_n18912 ), .ZN(_u10_n18904 ) );
NAND2_X1 _u10_U7516  ( .A1(1'b1), .A2(_u10_n12050 ), .ZN(_u10_n18906 ) );
NAND2_X1 _u10_U7515  ( .A1(1'b1), .A2(_u10_n12026 ), .ZN(_u10_n18907 ) );
NAND2_X1 _u10_U7514  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18908 ) );
NAND3_X1 _u10_U7513  ( .A1(_u10_n18906 ), .A2(_u10_n18907 ), .A3(_u10_n18908 ), .ZN(_u10_n18905 ) );
NOR4_X1 _u10_U7512  ( .A1(_u10_n18902 ), .A2(_u10_n18903 ), .A3(_u10_n18904 ), .A4(_u10_n18905 ), .ZN(_u10_n18880 ) );
NAND2_X1 _u10_U7511  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n18898 ) );
NAND2_X1 _u10_U7510  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n18899 ) );
NAND2_X1 _u10_U7509  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n18900 ) );
NAND2_X1 _u10_U7508  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n18901 ) );
NAND4_X1 _u10_U7507  ( .A1(_u10_n18898 ), .A2(_u10_n18899 ), .A3(_u10_n18900 ), .A4(_u10_n18901 ), .ZN(_u10_n18882 ) );
NAND2_X1 _u10_U7506  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n18894 ) );
NAND2_X1 _u10_U7505  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n18895 ) );
NAND2_X1 _u10_U7504  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n18896 ) );
NAND2_X1 _u10_U7503  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n18897 ) );
NAND4_X1 _u10_U7502  ( .A1(_u10_n18894 ), .A2(_u10_n18895 ), .A3(_u10_n18896 ), .A4(_u10_n18897 ), .ZN(_u10_n18883 ) );
NAND2_X1 _u10_U7501  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n18890 ) );
NAND2_X1 _u10_U7500  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n18891 ) );
NAND2_X1 _u10_U7499  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n18892 ) );
NAND2_X1 _u10_U7498  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n18893 ) );
NAND4_X1 _u10_U7497  ( .A1(_u10_n18890 ), .A2(_u10_n18891 ), .A3(_u10_n18892 ), .A4(_u10_n18893 ), .ZN(_u10_n18884 ) );
NAND2_X1 _u10_U7496  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n18886 ) );
NAND2_X1 _u10_U7495  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n18887 ) );
NAND2_X1 _u10_U7494  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n18888 ) );
NAND2_X1 _u10_U7493  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n18889 ) );
NAND4_X1 _u10_U7492  ( .A1(_u10_n18886 ), .A2(_u10_n18887 ), .A3(_u10_n18888 ), .A4(_u10_n18889 ), .ZN(_u10_n18885 ) );
NOR4_X1 _u10_U7491  ( .A1(_u10_n18882 ), .A2(_u10_n18883 ), .A3(_u10_n18884 ), .A4(_u10_n18885 ), .ZN(_u10_n18881 ) );
NAND2_X1 _u10_U7490  ( .A1(_u10_n18880 ), .A2(_u10_n18881 ), .ZN(am1[11]) );
NAND2_X1 _u10_U7489  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18876 ) );
NAND2_X1 _u10_U7488  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18877 ) );
NAND2_X1 _u10_U7487  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18878 ) );
NAND2_X1 _u10_U7486  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18879 ) );
NAND4_X1 _u10_U7485  ( .A1(_u10_n18876 ), .A2(_u10_n18877 ), .A3(_u10_n18878 ), .A4(_u10_n18879 ), .ZN(_u10_n18861 ) );
NAND2_X1 _u10_U7484  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18872 ) );
NAND2_X1 _u10_U7483  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18873 ) );
NAND2_X1 _u10_U7482  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18874 ) );
NAND2_X1 _u10_U7481  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18875 ) );
NAND4_X1 _u10_U7480  ( .A1(_u10_n18872 ), .A2(_u10_n18873 ), .A3(_u10_n18874 ), .A4(_u10_n18875 ), .ZN(_u10_n18862 ) );
NAND2_X1 _u10_U7479  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18868 ) );
NAND2_X1 _u10_U7478  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18869 ) );
NAND2_X1 _u10_U7477  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18870 ) );
NAND2_X1 _u10_U7476  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18871 ) );
NAND4_X1 _u10_U7475  ( .A1(_u10_n18868 ), .A2(_u10_n18869 ), .A3(_u10_n18870 ), .A4(_u10_n18871 ), .ZN(_u10_n18863 ) );
NAND2_X1 _u10_U7474  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18865 ) );
NAND2_X1 _u10_U7473  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18866 ) );
NAND2_X1 _u10_U7472  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18867 ) );
NAND3_X1 _u10_U7471  ( .A1(_u10_n18865 ), .A2(_u10_n18866 ), .A3(_u10_n18867 ), .ZN(_u10_n18864 ) );
NOR4_X1 _u10_U7470  ( .A1(_u10_n18861 ), .A2(_u10_n18862 ), .A3(_u10_n18863 ), .A4(_u10_n18864 ), .ZN(_u10_n18839 ) );
NAND2_X1 _u10_U7469  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n18857 ) );
NAND2_X1 _u10_U7468  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n18858 ) );
NAND2_X1 _u10_U7467  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n18859 ) );
NAND2_X1 _u10_U7466  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n18860 ) );
NAND4_X1 _u10_U7465  ( .A1(_u10_n18857 ), .A2(_u10_n18858 ), .A3(_u10_n18859 ), .A4(_u10_n18860 ), .ZN(_u10_n18841 ) );
NAND2_X1 _u10_U7464  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n18853 ) );
NAND2_X1 _u10_U7463  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n18854 ) );
NAND2_X1 _u10_U7462  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n18855 ) );
NAND2_X1 _u10_U7461  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n18856 ) );
NAND4_X1 _u10_U7460  ( .A1(_u10_n18853 ), .A2(_u10_n18854 ), .A3(_u10_n18855 ), .A4(_u10_n18856 ), .ZN(_u10_n18842 ) );
NAND2_X1 _u10_U7459  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n18849 ) );
NAND2_X1 _u10_U7458  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n18850 ) );
NAND2_X1 _u10_U7457  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n18851 ) );
NAND2_X1 _u10_U7456  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n18852 ) );
NAND4_X1 _u10_U7455  ( .A1(_u10_n18849 ), .A2(_u10_n18850 ), .A3(_u10_n18851 ), .A4(_u10_n18852 ), .ZN(_u10_n18843 ) );
NAND2_X1 _u10_U7454  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n18845 ) );
NAND2_X1 _u10_U7453  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n18846 ) );
NAND2_X1 _u10_U7452  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n18847 ) );
NAND2_X1 _u10_U7451  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n18848 ) );
NAND4_X1 _u10_U7450  ( .A1(_u10_n18845 ), .A2(_u10_n18846 ), .A3(_u10_n18847 ), .A4(_u10_n18848 ), .ZN(_u10_n18844 ) );
NOR4_X1 _u10_U7449  ( .A1(_u10_n18841 ), .A2(_u10_n18842 ), .A3(_u10_n18843 ), .A4(_u10_n18844 ), .ZN(_u10_n18840 ) );
NAND2_X1 _u10_U7448  ( .A1(_u10_n18839 ), .A2(_u10_n18840 ), .ZN(am1[12]) );
NAND2_X1 _u10_U7447  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18835 ) );
NAND2_X1 _u10_U7446  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18836 ) );
NAND2_X1 _u10_U7445  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18837 ) );
NAND2_X1 _u10_U7444  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18838 ) );
NAND4_X1 _u10_U7443  ( .A1(_u10_n18835 ), .A2(_u10_n18836 ), .A3(_u10_n18837 ), .A4(_u10_n18838 ), .ZN(_u10_n18820 ) );
NAND2_X1 _u10_U7442  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18831 ) );
NAND2_X1 _u10_U7441  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18832 ) );
NAND2_X1 _u10_U7440  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18833 ) );
NAND2_X1 _u10_U7439  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18834 ) );
NAND4_X1 _u10_U7438  ( .A1(_u10_n18831 ), .A2(_u10_n18832 ), .A3(_u10_n18833 ), .A4(_u10_n18834 ), .ZN(_u10_n18821 ) );
NAND2_X1 _u10_U7437  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18827 ) );
NAND2_X1 _u10_U7436  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18828 ) );
NAND2_X1 _u10_U7435  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18829 ) );
NAND2_X1 _u10_U7434  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18830 ) );
NAND4_X1 _u10_U7433  ( .A1(_u10_n18827 ), .A2(_u10_n18828 ), .A3(_u10_n18829 ), .A4(_u10_n18830 ), .ZN(_u10_n18822 ) );
NAND2_X1 _u10_U7432  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18824 ) );
NAND2_X1 _u10_U7431  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18825 ) );
NAND2_X1 _u10_U7430  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18826 ) );
NAND3_X1 _u10_U7429  ( .A1(_u10_n18824 ), .A2(_u10_n18825 ), .A3(_u10_n18826 ), .ZN(_u10_n18823 ) );
NOR4_X1 _u10_U7428  ( .A1(_u10_n18820 ), .A2(_u10_n18821 ), .A3(_u10_n18822 ), .A4(_u10_n18823 ), .ZN(_u10_n18798 ) );
NAND2_X1 _u10_U7427  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n18816 ) );
NAND2_X1 _u10_U7426  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n18817 ) );
NAND2_X1 _u10_U7425  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n18818 ) );
NAND2_X1 _u10_U7424  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n18819 ) );
NAND4_X1 _u10_U7423  ( .A1(_u10_n18816 ), .A2(_u10_n18817 ), .A3(_u10_n18818 ), .A4(_u10_n18819 ), .ZN(_u10_n18800 ) );
NAND2_X1 _u10_U7422  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n18812 ) );
NAND2_X1 _u10_U7421  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n18813 ) );
NAND2_X1 _u10_U7420  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n18814 ) );
NAND2_X1 _u10_U7419  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n18815 ) );
NAND4_X1 _u10_U7418  ( .A1(_u10_n18812 ), .A2(_u10_n18813 ), .A3(_u10_n18814 ), .A4(_u10_n18815 ), .ZN(_u10_n18801 ) );
NAND2_X1 _u10_U7417  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n18808 ) );
NAND2_X1 _u10_U7416  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n18809 ) );
NAND2_X1 _u10_U7415  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n18810 ) );
NAND2_X1 _u10_U7414  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n18811 ) );
NAND4_X1 _u10_U7413  ( .A1(_u10_n18808 ), .A2(_u10_n18809 ), .A3(_u10_n18810 ), .A4(_u10_n18811 ), .ZN(_u10_n18802 ) );
NAND2_X1 _u10_U7412  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n18804 ) );
NAND2_X1 _u10_U7411  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n18805 ) );
NAND2_X1 _u10_U7410  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n18806 ) );
NAND2_X1 _u10_U7409  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n18807 ) );
NAND4_X1 _u10_U7408  ( .A1(_u10_n18804 ), .A2(_u10_n18805 ), .A3(_u10_n18806 ), .A4(_u10_n18807 ), .ZN(_u10_n18803 ) );
NOR4_X1 _u10_U7407  ( .A1(_u10_n18800 ), .A2(_u10_n18801 ), .A3(_u10_n18802 ), .A4(_u10_n18803 ), .ZN(_u10_n18799 ) );
NAND2_X1 _u10_U7406  ( .A1(_u10_n18798 ), .A2(_u10_n18799 ), .ZN(am1[13]) );
NAND2_X1 _u10_U7405  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18794 ) );
NAND2_X1 _u10_U7404  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18795 ) );
NAND2_X1 _u10_U7403  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18796 ) );
NAND2_X1 _u10_U7402  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18797 ) );
NAND4_X1 _u10_U7401  ( .A1(_u10_n18794 ), .A2(_u10_n18795 ), .A3(_u10_n18796 ), .A4(_u10_n18797 ), .ZN(_u10_n18779 ) );
NAND2_X1 _u10_U7400  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18790 ) );
NAND2_X1 _u10_U7399  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18791 ) );
NAND2_X1 _u10_U7398  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18792 ) );
NAND2_X1 _u10_U7397  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18793 ) );
NAND4_X1 _u10_U7396  ( .A1(_u10_n18790 ), .A2(_u10_n18791 ), .A3(_u10_n18792 ), .A4(_u10_n18793 ), .ZN(_u10_n18780 ) );
NAND2_X1 _u10_U7395  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18786 ) );
NAND2_X1 _u10_U7394  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18787 ) );
NAND2_X1 _u10_U7393  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18788 ) );
NAND2_X1 _u10_U7392  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18789 ) );
NAND4_X1 _u10_U7391  ( .A1(_u10_n18786 ), .A2(_u10_n18787 ), .A3(_u10_n18788 ), .A4(_u10_n18789 ), .ZN(_u10_n18781 ) );
NAND2_X1 _u10_U7390  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18783 ) );
NAND2_X1 _u10_U7389  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18784 ) );
NAND2_X1 _u10_U7388  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18785 ) );
NAND3_X1 _u10_U7387  ( .A1(_u10_n18783 ), .A2(_u10_n18784 ), .A3(_u10_n18785 ), .ZN(_u10_n18782 ) );
NOR4_X1 _u10_U7386  ( .A1(_u10_n18779 ), .A2(_u10_n18780 ), .A3(_u10_n18781 ), .A4(_u10_n18782 ), .ZN(_u10_n18757 ) );
NAND2_X1 _u10_U7385  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n18775 ) );
NAND2_X1 _u10_U7384  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n18776 ) );
NAND2_X1 _u10_U7383  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n18777 ) );
NAND2_X1 _u10_U7382  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n18778 ) );
NAND4_X1 _u10_U7381  ( .A1(_u10_n18775 ), .A2(_u10_n18776 ), .A3(_u10_n18777 ), .A4(_u10_n18778 ), .ZN(_u10_n18759 ) );
NAND2_X1 _u10_U7380  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n18771 ) );
NAND2_X1 _u10_U7379  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n18772 ) );
NAND2_X1 _u10_U7378  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n18773 ) );
NAND2_X1 _u10_U7377  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n18774 ) );
NAND4_X1 _u10_U7376  ( .A1(_u10_n18771 ), .A2(_u10_n18772 ), .A3(_u10_n18773 ), .A4(_u10_n18774 ), .ZN(_u10_n18760 ) );
NAND2_X1 _u10_U7375  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n18767 ) );
NAND2_X1 _u10_U7374  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n18768 ) );
NAND2_X1 _u10_U7373  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n18769 ) );
NAND2_X1 _u10_U7372  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n18770 ) );
NAND4_X1 _u10_U7371  ( .A1(_u10_n18767 ), .A2(_u10_n18768 ), .A3(_u10_n18769 ), .A4(_u10_n18770 ), .ZN(_u10_n18761 ) );
NAND2_X1 _u10_U7370  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n18763 ) );
NAND2_X1 _u10_U7369  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n18764 ) );
NAND2_X1 _u10_U7368  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n18765 ) );
NAND2_X1 _u10_U7367  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n18766 ) );
NAND4_X1 _u10_U7366  ( .A1(_u10_n18763 ), .A2(_u10_n18764 ), .A3(_u10_n18765 ), .A4(_u10_n18766 ), .ZN(_u10_n18762 ) );
NOR4_X1 _u10_U7365  ( .A1(_u10_n18759 ), .A2(_u10_n18760 ), .A3(_u10_n18761 ), .A4(_u10_n18762 ), .ZN(_u10_n18758 ) );
NAND2_X1 _u10_U7364  ( .A1(_u10_n18757 ), .A2(_u10_n18758 ), .ZN(am1[14]) );
NAND2_X1 _u10_U7363  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18753 ) );
NAND2_X1 _u10_U7362  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18754 ) );
NAND2_X1 _u10_U7361  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18755 ) );
NAND2_X1 _u10_U7360  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18756 ) );
NAND4_X1 _u10_U7359  ( .A1(_u10_n18753 ), .A2(_u10_n18754 ), .A3(_u10_n18755 ), .A4(_u10_n18756 ), .ZN(_u10_n18738 ) );
NAND2_X1 _u10_U7358  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18749 ) );
NAND2_X1 _u10_U7357  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18750 ) );
NAND2_X1 _u10_U7356  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18751 ) );
NAND2_X1 _u10_U7355  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18752 ) );
NAND4_X1 _u10_U7354  ( .A1(_u10_n18749 ), .A2(_u10_n18750 ), .A3(_u10_n18751 ), .A4(_u10_n18752 ), .ZN(_u10_n18739 ) );
NAND2_X1 _u10_U7353  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18745 ) );
NAND2_X1 _u10_U7352  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18746 ) );
NAND2_X1 _u10_U7351  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18747 ) );
NAND2_X1 _u10_U7350  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18748 ) );
NAND4_X1 _u10_U7349  ( .A1(_u10_n18745 ), .A2(_u10_n18746 ), .A3(_u10_n18747 ), .A4(_u10_n18748 ), .ZN(_u10_n18740 ) );
NAND2_X1 _u10_U7348  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18742 ) );
NAND2_X1 _u10_U7347  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18743 ) );
NAND2_X1 _u10_U7346  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18744 ) );
NAND3_X1 _u10_U7345  ( .A1(_u10_n18742 ), .A2(_u10_n18743 ), .A3(_u10_n18744 ), .ZN(_u10_n18741 ) );
NOR4_X1 _u10_U7344  ( .A1(_u10_n18738 ), .A2(_u10_n18739 ), .A3(_u10_n18740 ), .A4(_u10_n18741 ), .ZN(_u10_n18716 ) );
NAND2_X1 _u10_U7343  ( .A1(1'b1), .A2(_u10_n11990 ), .ZN(_u10_n18734 ) );
NAND2_X1 _u10_U7342  ( .A1(1'b1), .A2(_u10_n11966 ), .ZN(_u10_n18735 ) );
NAND2_X1 _u10_U7341  ( .A1(1'b1), .A2(_u10_n11942 ), .ZN(_u10_n18736 ) );
NAND2_X1 _u10_U7340  ( .A1(1'b1), .A2(_u10_n11918 ), .ZN(_u10_n18737 ) );
NAND4_X1 _u10_U7339  ( .A1(_u10_n18734 ), .A2(_u10_n18735 ), .A3(_u10_n18736 ), .A4(_u10_n18737 ), .ZN(_u10_n18718 ) );
NAND2_X1 _u10_U7338  ( .A1(1'b1), .A2(_u10_n11894 ), .ZN(_u10_n18730 ) );
NAND2_X1 _u10_U7337  ( .A1(1'b1), .A2(_u10_n11870 ), .ZN(_u10_n18731 ) );
NAND2_X1 _u10_U7336  ( .A1(1'b1), .A2(_u10_n11846 ), .ZN(_u10_n18732 ) );
NAND2_X1 _u10_U7335  ( .A1(1'b1), .A2(_u10_n11822 ), .ZN(_u10_n18733 ) );
NAND4_X1 _u10_U7334  ( .A1(_u10_n18730 ), .A2(_u10_n18731 ), .A3(_u10_n18732 ), .A4(_u10_n18733 ), .ZN(_u10_n18719 ) );
NAND2_X1 _u10_U7333  ( .A1(1'b1), .A2(_u10_n11798 ), .ZN(_u10_n18726 ) );
NAND2_X1 _u10_U7332  ( .A1(1'b1), .A2(_u10_n11774 ), .ZN(_u10_n18727 ) );
NAND2_X1 _u10_U7331  ( .A1(1'b1), .A2(_u10_n11750 ), .ZN(_u10_n18728 ) );
NAND2_X1 _u10_U7330  ( .A1(1'b1), .A2(_u10_n11726 ), .ZN(_u10_n18729 ) );
NAND4_X1 _u10_U7329  ( .A1(_u10_n18726 ), .A2(_u10_n18727 ), .A3(_u10_n18728 ), .A4(_u10_n18729 ), .ZN(_u10_n18720 ) );
NAND2_X1 _u10_U7328  ( .A1(1'b1), .A2(_u10_n11702 ), .ZN(_u10_n18722 ) );
NAND2_X1 _u10_U7327  ( .A1(1'b1), .A2(_u10_n11678 ), .ZN(_u10_n18723 ) );
NAND2_X1 _u10_U7326  ( .A1(1'b1), .A2(_u10_n11654 ), .ZN(_u10_n18724 ) );
NAND2_X1 _u10_U7325  ( .A1(1'b1), .A2(_u10_n11630 ), .ZN(_u10_n18725 ) );
NAND4_X1 _u10_U7324  ( .A1(_u10_n18722 ), .A2(_u10_n18723 ), .A3(_u10_n18724 ), .A4(_u10_n18725 ), .ZN(_u10_n18721 ) );
NOR4_X1 _u10_U7323  ( .A1(_u10_n18718 ), .A2(_u10_n18719 ), .A3(_u10_n18720 ), .A4(_u10_n18721 ), .ZN(_u10_n18717 ) );
NAND2_X1 _u10_U7322  ( .A1(_u10_n18716 ), .A2(_u10_n18717 ), .ZN(am1[15]) );
NAND2_X1 _u10_U7321  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18712 ) );
NAND2_X1 _u10_U7320  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18713 ) );
NAND2_X1 _u10_U7319  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18714 ) );
NAND2_X1 _u10_U7318  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18715 ) );
NAND4_X1 _u10_U7317  ( .A1(_u10_n18712 ), .A2(_u10_n18713 ), .A3(_u10_n18714 ), .A4(_u10_n18715 ), .ZN(_u10_n18697 ) );
NAND2_X1 _u10_U7316  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18708 ) );
NAND2_X1 _u10_U7315  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18709 ) );
NAND2_X1 _u10_U7314  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18710 ) );
NAND2_X1 _u10_U7313  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18711 ) );
NAND4_X1 _u10_U7312  ( .A1(_u10_n18708 ), .A2(_u10_n18709 ), .A3(_u10_n18710 ), .A4(_u10_n18711 ), .ZN(_u10_n18698 ) );
NAND2_X1 _u10_U7311  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18704 ) );
NAND2_X1 _u10_U7310  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18705 ) );
NAND2_X1 _u10_U7309  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18706 ) );
NAND2_X1 _u10_U7308  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18707 ) );
NAND4_X1 _u10_U7307  ( .A1(_u10_n18704 ), .A2(_u10_n18705 ), .A3(_u10_n18706 ), .A4(_u10_n18707 ), .ZN(_u10_n18699 ) );
NAND2_X1 _u10_U7306  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18701 ) );
NAND2_X1 _u10_U7305  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18702 ) );
NAND2_X1 _u10_U7304  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18703 ) );
NAND3_X1 _u10_U7303  ( .A1(_u10_n18701 ), .A2(_u10_n18702 ), .A3(_u10_n18703 ), .ZN(_u10_n18700 ) );
NOR4_X1 _u10_U7302  ( .A1(_u10_n18697 ), .A2(_u10_n18698 ), .A3(_u10_n18699 ), .A4(_u10_n18700 ), .ZN(_u10_n18675 ) );
NAND2_X1 _u10_U7301  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18693 ) );
NAND2_X1 _u10_U7300  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18694 ) );
NAND2_X1 _u10_U7299  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18695 ) );
NAND2_X1 _u10_U7298  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18696 ) );
NAND4_X1 _u10_U7297  ( .A1(_u10_n18693 ), .A2(_u10_n18694 ), .A3(_u10_n18695 ), .A4(_u10_n18696 ), .ZN(_u10_n18677 ) );
NAND2_X1 _u10_U7296  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18689 ) );
NAND2_X1 _u10_U7295  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18690 ) );
NAND2_X1 _u10_U7294  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18691 ) );
NAND2_X1 _u10_U7293  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18692 ) );
NAND4_X1 _u10_U7292  ( .A1(_u10_n18689 ), .A2(_u10_n18690 ), .A3(_u10_n18691 ), .A4(_u10_n18692 ), .ZN(_u10_n18678 ) );
NAND2_X1 _u10_U7291  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18685 ) );
NAND2_X1 _u10_U7290  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18686 ) );
NAND2_X1 _u10_U7289  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18687 ) );
NAND2_X1 _u10_U7288  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18688 ) );
NAND4_X1 _u10_U7287  ( .A1(_u10_n18685 ), .A2(_u10_n18686 ), .A3(_u10_n18687 ), .A4(_u10_n18688 ), .ZN(_u10_n18679 ) );
NAND2_X1 _u10_U7286  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18681 ) );
NAND2_X1 _u10_U7285  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18682 ) );
NAND2_X1 _u10_U7284  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18683 ) );
NAND2_X1 _u10_U7283  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18684 ) );
NAND4_X1 _u10_U7282  ( .A1(_u10_n18681 ), .A2(_u10_n18682 ), .A3(_u10_n18683 ), .A4(_u10_n18684 ), .ZN(_u10_n18680 ) );
NOR4_X1 _u10_U7281  ( .A1(_u10_n18677 ), .A2(_u10_n18678 ), .A3(_u10_n18679 ), .A4(_u10_n18680 ), .ZN(_u10_n18676 ) );
NAND2_X1 _u10_U7280  ( .A1(_u10_n18675 ), .A2(_u10_n18676 ), .ZN(am1[16]) );
NAND2_X1 _u10_U7279  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18671 ) );
NAND2_X1 _u10_U7278  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18672 ) );
NAND2_X1 _u10_U7277  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18673 ) );
NAND2_X1 _u10_U7276  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18674 ) );
NAND4_X1 _u10_U7275  ( .A1(_u10_n18671 ), .A2(_u10_n18672 ), .A3(_u10_n18673 ), .A4(_u10_n18674 ), .ZN(_u10_n18656 ) );
NAND2_X1 _u10_U7274  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18667 ) );
NAND2_X1 _u10_U7273  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18668 ) );
NAND2_X1 _u10_U7272  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18669 ) );
NAND2_X1 _u10_U7271  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18670 ) );
NAND4_X1 _u10_U7270  ( .A1(_u10_n18667 ), .A2(_u10_n18668 ), .A3(_u10_n18669 ), .A4(_u10_n18670 ), .ZN(_u10_n18657 ) );
NAND2_X1 _u10_U7269  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18663 ) );
NAND2_X1 _u10_U7268  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18664 ) );
NAND2_X1 _u10_U7267  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18665 ) );
NAND2_X1 _u10_U7266  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18666 ) );
NAND4_X1 _u10_U7265  ( .A1(_u10_n18663 ), .A2(_u10_n18664 ), .A3(_u10_n18665 ), .A4(_u10_n18666 ), .ZN(_u10_n18658 ) );
NAND2_X1 _u10_U7264  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18660 ) );
NAND2_X1 _u10_U7263  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18661 ) );
NAND2_X1 _u10_U7262  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18662 ) );
NAND3_X1 _u10_U7261  ( .A1(_u10_n18660 ), .A2(_u10_n18661 ), .A3(_u10_n18662 ), .ZN(_u10_n18659 ) );
NOR4_X1 _u10_U7260  ( .A1(_u10_n18656 ), .A2(_u10_n18657 ), .A3(_u10_n18658 ), .A4(_u10_n18659 ), .ZN(_u10_n18634 ) );
NAND2_X1 _u10_U7259  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18652 ) );
NAND2_X1 _u10_U7258  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18653 ) );
NAND2_X1 _u10_U7257  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18654 ) );
NAND2_X1 _u10_U7256  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18655 ) );
NAND4_X1 _u10_U7255  ( .A1(_u10_n18652 ), .A2(_u10_n18653 ), .A3(_u10_n18654 ), .A4(_u10_n18655 ), .ZN(_u10_n18636 ) );
NAND2_X1 _u10_U7254  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18648 ) );
NAND2_X1 _u10_U7253  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18649 ) );
NAND2_X1 _u10_U7252  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18650 ) );
NAND2_X1 _u10_U7251  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18651 ) );
NAND4_X1 _u10_U7250  ( .A1(_u10_n18648 ), .A2(_u10_n18649 ), .A3(_u10_n18650 ), .A4(_u10_n18651 ), .ZN(_u10_n18637 ) );
NAND2_X1 _u10_U7249  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18644 ) );
NAND2_X1 _u10_U7248  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18645 ) );
NAND2_X1 _u10_U7247  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18646 ) );
NAND2_X1 _u10_U7246  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18647 ) );
NAND4_X1 _u10_U7245  ( .A1(_u10_n18644 ), .A2(_u10_n18645 ), .A3(_u10_n18646 ), .A4(_u10_n18647 ), .ZN(_u10_n18638 ) );
NAND2_X1 _u10_U7244  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18640 ) );
NAND2_X1 _u10_U7243  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18641 ) );
NAND2_X1 _u10_U7242  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18642 ) );
NAND2_X1 _u10_U7241  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18643 ) );
NAND4_X1 _u10_U7240  ( .A1(_u10_n18640 ), .A2(_u10_n18641 ), .A3(_u10_n18642 ), .A4(_u10_n18643 ), .ZN(_u10_n18639 ) );
NOR4_X1 _u10_U7239  ( .A1(_u10_n18636 ), .A2(_u10_n18637 ), .A3(_u10_n18638 ), .A4(_u10_n18639 ), .ZN(_u10_n18635 ) );
NAND2_X1 _u10_U7238  ( .A1(_u10_n18634 ), .A2(_u10_n18635 ), .ZN(am1[17]) );
NAND2_X1 _u10_U7237  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18630 ) );
NAND2_X1 _u10_U7236  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18631 ) );
NAND2_X1 _u10_U7235  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18632 ) );
NAND2_X1 _u10_U7234  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18633 ) );
NAND4_X1 _u10_U7233  ( .A1(_u10_n18630 ), .A2(_u10_n18631 ), .A3(_u10_n18632 ), .A4(_u10_n18633 ), .ZN(_u10_n18615 ) );
NAND2_X1 _u10_U7232  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18626 ) );
NAND2_X1 _u10_U7231  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18627 ) );
NAND2_X1 _u10_U7230  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18628 ) );
NAND2_X1 _u10_U7229  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18629 ) );
NAND4_X1 _u10_U7228  ( .A1(_u10_n18626 ), .A2(_u10_n18627 ), .A3(_u10_n18628 ), .A4(_u10_n18629 ), .ZN(_u10_n18616 ) );
NAND2_X1 _u10_U7227  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18622 ) );
NAND2_X1 _u10_U7226  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18623 ) );
NAND2_X1 _u10_U7225  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18624 ) );
NAND2_X1 _u10_U7224  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18625 ) );
NAND4_X1 _u10_U7223  ( .A1(_u10_n18622 ), .A2(_u10_n18623 ), .A3(_u10_n18624 ), .A4(_u10_n18625 ), .ZN(_u10_n18617 ) );
NAND2_X1 _u10_U7222  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18619 ) );
NAND2_X1 _u10_U7221  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18620 ) );
NAND2_X1 _u10_U7220  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18621 ) );
NAND3_X1 _u10_U7219  ( .A1(_u10_n18619 ), .A2(_u10_n18620 ), .A3(_u10_n18621 ), .ZN(_u10_n18618 ) );
NOR4_X1 _u10_U7218  ( .A1(_u10_n18615 ), .A2(_u10_n18616 ), .A3(_u10_n18617 ), .A4(_u10_n18618 ), .ZN(_u10_n18593 ) );
NAND2_X1 _u10_U7217  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18611 ) );
NAND2_X1 _u10_U7216  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18612 ) );
NAND2_X1 _u10_U7215  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18613 ) );
NAND2_X1 _u10_U7214  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18614 ) );
NAND4_X1 _u10_U7213  ( .A1(_u10_n18611 ), .A2(_u10_n18612 ), .A3(_u10_n18613 ), .A4(_u10_n18614 ), .ZN(_u10_n18595 ) );
NAND2_X1 _u10_U7212  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18607 ) );
NAND2_X1 _u10_U7211  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18608 ) );
NAND2_X1 _u10_U7210  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18609 ) );
NAND2_X1 _u10_U7209  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18610 ) );
NAND4_X1 _u10_U7208  ( .A1(_u10_n18607 ), .A2(_u10_n18608 ), .A3(_u10_n18609 ), .A4(_u10_n18610 ), .ZN(_u10_n18596 ) );
NAND2_X1 _u10_U7207  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18603 ) );
NAND2_X1 _u10_U7206  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18604 ) );
NAND2_X1 _u10_U7205  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18605 ) );
NAND2_X1 _u10_U7204  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18606 ) );
NAND4_X1 _u10_U7203  ( .A1(_u10_n18603 ), .A2(_u10_n18604 ), .A3(_u10_n18605 ), .A4(_u10_n18606 ), .ZN(_u10_n18597 ) );
NAND2_X1 _u10_U7202  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18599 ) );
NAND2_X1 _u10_U7201  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18600 ) );
NAND2_X1 _u10_U7200  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18601 ) );
NAND2_X1 _u10_U7199  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18602 ) );
NAND4_X1 _u10_U7198  ( .A1(_u10_n18599 ), .A2(_u10_n18600 ), .A3(_u10_n18601 ), .A4(_u10_n18602 ), .ZN(_u10_n18598 ) );
NOR4_X1 _u10_U7197  ( .A1(_u10_n18595 ), .A2(_u10_n18596 ), .A3(_u10_n18597 ), .A4(_u10_n18598 ), .ZN(_u10_n18594 ) );
NAND2_X1 _u10_U7196  ( .A1(_u10_n18593 ), .A2(_u10_n18594 ), .ZN(am1[18]) );
NAND2_X1 _u10_U7195  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18589 ) );
NAND2_X1 _u10_U7194  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18590 ) );
NAND2_X1 _u10_U7193  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18591 ) );
NAND2_X1 _u10_U7192  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18592 ) );
NAND4_X1 _u10_U7191  ( .A1(_u10_n18589 ), .A2(_u10_n18590 ), .A3(_u10_n18591 ), .A4(_u10_n18592 ), .ZN(_u10_n18574 ) );
NAND2_X1 _u10_U7190  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18585 ) );
NAND2_X1 _u10_U7189  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18586 ) );
NAND2_X1 _u10_U7188  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18587 ) );
NAND2_X1 _u10_U7187  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18588 ) );
NAND4_X1 _u10_U7186  ( .A1(_u10_n18585 ), .A2(_u10_n18586 ), .A3(_u10_n18587 ), .A4(_u10_n18588 ), .ZN(_u10_n18575 ) );
NAND2_X1 _u10_U7185  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18581 ) );
NAND2_X1 _u10_U7184  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18582 ) );
NAND2_X1 _u10_U7183  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18583 ) );
NAND2_X1 _u10_U7182  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18584 ) );
NAND4_X1 _u10_U7181  ( .A1(_u10_n18581 ), .A2(_u10_n18582 ), .A3(_u10_n18583 ), .A4(_u10_n18584 ), .ZN(_u10_n18576 ) );
NAND2_X1 _u10_U7180  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18578 ) );
NAND2_X1 _u10_U7179  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18579 ) );
NAND2_X1 _u10_U7178  ( .A1(1'b1), .A2(_u10_n12007 ), .ZN(_u10_n18580 ) );
NAND3_X1 _u10_U7177  ( .A1(_u10_n18578 ), .A2(_u10_n18579 ), .A3(_u10_n18580 ), .ZN(_u10_n18577 ) );
NOR4_X1 _u10_U7176  ( .A1(_u10_n18574 ), .A2(_u10_n18575 ), .A3(_u10_n18576 ), .A4(_u10_n18577 ), .ZN(_u10_n18552 ) );
NAND2_X1 _u10_U7175  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18570 ) );
NAND2_X1 _u10_U7174  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18571 ) );
NAND2_X1 _u10_U7173  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18572 ) );
NAND2_X1 _u10_U7172  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18573 ) );
NAND4_X1 _u10_U7171  ( .A1(_u10_n18570 ), .A2(_u10_n18571 ), .A3(_u10_n18572 ), .A4(_u10_n18573 ), .ZN(_u10_n18554 ) );
NAND2_X1 _u10_U7170  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18566 ) );
NAND2_X1 _u10_U7169  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18567 ) );
NAND2_X1 _u10_U7168  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18568 ) );
NAND2_X1 _u10_U7167  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18569 ) );
NAND4_X1 _u10_U7166  ( .A1(_u10_n18566 ), .A2(_u10_n18567 ), .A3(_u10_n18568 ), .A4(_u10_n18569 ), .ZN(_u10_n18555 ) );
NAND2_X1 _u10_U7165  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18562 ) );
NAND2_X1 _u10_U7164  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18563 ) );
NAND2_X1 _u10_U7163  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18564 ) );
NAND2_X1 _u10_U7162  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18565 ) );
NAND4_X1 _u10_U7161  ( .A1(_u10_n18562 ), .A2(_u10_n18563 ), .A3(_u10_n18564 ), .A4(_u10_n18565 ), .ZN(_u10_n18556 ) );
NAND2_X1 _u10_U7160  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18558 ) );
NAND2_X1 _u10_U7159  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18559 ) );
NAND2_X1 _u10_U7158  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18560 ) );
NAND2_X1 _u10_U7157  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18561 ) );
NAND4_X1 _u10_U7156  ( .A1(_u10_n18558 ), .A2(_u10_n18559 ), .A3(_u10_n18560 ), .A4(_u10_n18561 ), .ZN(_u10_n18557 ) );
NOR4_X1 _u10_U7155  ( .A1(_u10_n18554 ), .A2(_u10_n18555 ), .A3(_u10_n18556 ), .A4(_u10_n18557 ), .ZN(_u10_n18553 ) );
NAND2_X1 _u10_U7154  ( .A1(_u10_n18552 ), .A2(_u10_n18553 ), .ZN(am1[19]) );
NAND2_X1 _u10_U7153  ( .A1(1'b0), .A2(_u10_n12338 ), .ZN(_u10_n18548 ) );
NAND2_X1 _u10_U7152  ( .A1(1'b0), .A2(_u10_n12315 ), .ZN(_u10_n18549 ) );
NAND2_X1 _u10_U7151  ( .A1(1'b0), .A2(_u10_n12291 ), .ZN(_u10_n18550 ) );
NAND2_X1 _u10_U7150  ( .A1(1'b0), .A2(_u10_n12267 ), .ZN(_u10_n18551 ) );
NAND4_X1 _u10_U7149  ( .A1(_u10_n18548 ), .A2(_u10_n18549 ), .A3(_u10_n18550 ), .A4(_u10_n18551 ), .ZN(_u10_n18533 ) );
NAND2_X1 _u10_U7148  ( .A1(1'b0), .A2(_u10_n12242 ), .ZN(_u10_n18544 ) );
NAND2_X1 _u10_U7147  ( .A1(1'b0), .A2(_u10_n12218 ), .ZN(_u10_n18545 ) );
NAND2_X1 _u10_U7146  ( .A1(1'b0), .A2(_u10_n12195 ), .ZN(_u10_n18546 ) );
NAND2_X1 _u10_U7145  ( .A1(1'b0), .A2(_u10_n12170 ), .ZN(_u10_n18547 ) );
NAND4_X1 _u10_U7144  ( .A1(_u10_n18544 ), .A2(_u10_n18545 ), .A3(_u10_n18546 ), .A4(_u10_n18547 ), .ZN(_u10_n18534 ) );
NAND2_X1 _u10_U7143  ( .A1(1'b0), .A2(_u10_n12147 ), .ZN(_u10_n18540 ) );
NAND2_X1 _u10_U7142  ( .A1(1'b0), .A2(_u10_n12123 ), .ZN(_u10_n18541 ) );
NAND2_X1 _u10_U7141  ( .A1(1'b0), .A2(_u10_n12099 ), .ZN(_u10_n18542 ) );
NAND2_X1 _u10_U7140  ( .A1(1'b0), .A2(_u10_n12075 ), .ZN(_u10_n18543 ) );
NAND4_X1 _u10_U7139  ( .A1(_u10_n18540 ), .A2(_u10_n18541 ), .A3(_u10_n18542 ), .A4(_u10_n18543 ), .ZN(_u10_n18535 ) );
NAND2_X1 _u10_U7138  ( .A1(1'b0), .A2(_u10_n12051 ), .ZN(_u10_n18537 ) );
NAND2_X1 _u10_U7137  ( .A1(1'b0), .A2(_u10_n12027 ), .ZN(_u10_n18538 ) );
NAND2_X1 _u10_U7136  ( .A1(1'b0), .A2(_u10_n12008 ), .ZN(_u10_n18539 ) );
NAND3_X1 _u10_U7135  ( .A1(_u10_n18537 ), .A2(_u10_n18538 ), .A3(_u10_n18539 ), .ZN(_u10_n18536 ) );
NOR4_X1 _u10_U7134  ( .A1(_u10_n18533 ), .A2(_u10_n18534 ), .A3(_u10_n18535 ), .A4(_u10_n18536 ), .ZN(_u10_n18511 ) );
NAND2_X1 _u10_U7133  ( .A1(1'b0), .A2(_u10_n11991 ), .ZN(_u10_n18529 ) );
NAND2_X1 _u10_U7132  ( .A1(1'b0), .A2(_u10_n11967 ), .ZN(_u10_n18530 ) );
NAND2_X1 _u10_U7131  ( .A1(1'b0), .A2(_u10_n11943 ), .ZN(_u10_n18531 ) );
NAND2_X1 _u10_U7130  ( .A1(1'b0), .A2(_u10_n11919 ), .ZN(_u10_n18532 ) );
NAND4_X1 _u10_U7129  ( .A1(_u10_n18529 ), .A2(_u10_n18530 ), .A3(_u10_n18531 ), .A4(_u10_n18532 ), .ZN(_u10_n18513 ) );
NAND2_X1 _u10_U7128  ( .A1(1'b0), .A2(_u10_n11895 ), .ZN(_u10_n18525 ) );
NAND2_X1 _u10_U7127  ( .A1(1'b0), .A2(_u10_n11871 ), .ZN(_u10_n18526 ) );
NAND2_X1 _u10_U7126  ( .A1(1'b0), .A2(_u10_n11847 ), .ZN(_u10_n18527 ) );
NAND2_X1 _u10_U7125  ( .A1(1'b0), .A2(_u10_n11823 ), .ZN(_u10_n18528 ) );
NAND4_X1 _u10_U7124  ( .A1(_u10_n18525 ), .A2(_u10_n18526 ), .A3(_u10_n18527 ), .A4(_u10_n18528 ), .ZN(_u10_n18514 ) );
NAND2_X1 _u10_U7123  ( .A1(1'b0), .A2(_u10_n11799 ), .ZN(_u10_n18521 ) );
NAND2_X1 _u10_U7122  ( .A1(1'b0), .A2(_u10_n11775 ), .ZN(_u10_n18522 ) );
NAND2_X1 _u10_U7121  ( .A1(1'b0), .A2(_u10_n11751 ), .ZN(_u10_n18523 ) );
NAND2_X1 _u10_U7120  ( .A1(1'b0), .A2(_u10_n11727 ), .ZN(_u10_n18524 ) );
NAND4_X1 _u10_U7119  ( .A1(_u10_n18521 ), .A2(_u10_n18522 ), .A3(_u10_n18523 ), .A4(_u10_n18524 ), .ZN(_u10_n18515 ) );
NAND2_X1 _u10_U7118  ( .A1(1'b0), .A2(_u10_n11703 ), .ZN(_u10_n18517 ) );
NAND2_X1 _u10_U7117  ( .A1(1'b0), .A2(_u10_n11679 ), .ZN(_u10_n18518 ) );
NAND2_X1 _u10_U7116  ( .A1(1'b0), .A2(_u10_n11655 ), .ZN(_u10_n18519 ) );
NAND2_X1 _u10_U7115  ( .A1(1'b0), .A2(_u10_n11631 ), .ZN(_u10_n18520 ) );
NAND4_X1 _u10_U7114  ( .A1(_u10_n18517 ), .A2(_u10_n18518 ), .A3(_u10_n18519 ), .A4(_u10_n18520 ), .ZN(_u10_n18516 ) );
NOR4_X1 _u10_U7113  ( .A1(_u10_n18513 ), .A2(_u10_n18514 ), .A3(_u10_n18515 ), .A4(_u10_n18516 ), .ZN(_u10_n18512 ) );
NAND2_X1 _u10_U7112  ( .A1(_u10_n18511 ), .A2(_u10_n18512 ), .ZN(am1[1]) );
NAND2_X1 _u10_U7111  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18507 ) );
NAND2_X1 _u10_U7110  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18508 ) );
NAND2_X1 _u10_U7109  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18509 ) );
NAND2_X1 _u10_U7108  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18510 ) );
NAND4_X1 _u10_U7107  ( .A1(_u10_n18507 ), .A2(_u10_n18508 ), .A3(_u10_n18509 ), .A4(_u10_n18510 ), .ZN(_u10_n18492 ) );
NAND2_X1 _u10_U7106  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18503 ) );
NAND2_X1 _u10_U7105  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18504 ) );
NAND2_X1 _u10_U7104  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18505 ) );
NAND2_X1 _u10_U7103  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18506 ) );
NAND4_X1 _u10_U7102  ( .A1(_u10_n18503 ), .A2(_u10_n18504 ), .A3(_u10_n18505 ), .A4(_u10_n18506 ), .ZN(_u10_n18493 ) );
NAND2_X1 _u10_U7101  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18499 ) );
NAND2_X1 _u10_U7100  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18500 ) );
NAND2_X1 _u10_U7099  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18501 ) );
NAND2_X1 _u10_U7098  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18502 ) );
NAND4_X1 _u10_U7097  ( .A1(_u10_n18499 ), .A2(_u10_n18500 ), .A3(_u10_n18501 ), .A4(_u10_n18502 ), .ZN(_u10_n18494 ) );
NAND2_X1 _u10_U7096  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18496 ) );
NAND2_X1 _u10_U7095  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18497 ) );
NAND2_X1 _u10_U7094  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18498 ) );
NAND3_X1 _u10_U7093  ( .A1(_u10_n18496 ), .A2(_u10_n18497 ), .A3(_u10_n18498 ), .ZN(_u10_n18495 ) );
NOR4_X1 _u10_U7092  ( .A1(_u10_n18492 ), .A2(_u10_n18493 ), .A3(_u10_n18494 ), .A4(_u10_n18495 ), .ZN(_u10_n18470 ) );
NAND2_X1 _u10_U7091  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18488 ) );
NAND2_X1 _u10_U7090  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18489 ) );
NAND2_X1 _u10_U7089  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18490 ) );
NAND2_X1 _u10_U7088  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18491 ) );
NAND4_X1 _u10_U7087  ( .A1(_u10_n18488 ), .A2(_u10_n18489 ), .A3(_u10_n18490 ), .A4(_u10_n18491 ), .ZN(_u10_n18472 ) );
NAND2_X1 _u10_U7086  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18484 ) );
NAND2_X1 _u10_U7085  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18485 ) );
NAND2_X1 _u10_U7084  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18486 ) );
NAND2_X1 _u10_U7083  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18487 ) );
NAND4_X1 _u10_U7082  ( .A1(_u10_n18484 ), .A2(_u10_n18485 ), .A3(_u10_n18486 ), .A4(_u10_n18487 ), .ZN(_u10_n18473 ) );
NAND2_X1 _u10_U7081  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18480 ) );
NAND2_X1 _u10_U7080  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18481 ) );
NAND2_X1 _u10_U7079  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18482 ) );
NAND2_X1 _u10_U7078  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18483 ) );
NAND4_X1 _u10_U7077  ( .A1(_u10_n18480 ), .A2(_u10_n18481 ), .A3(_u10_n18482 ), .A4(_u10_n18483 ), .ZN(_u10_n18474 ) );
NAND2_X1 _u10_U7076  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18476 ) );
NAND2_X1 _u10_U7075  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18477 ) );
NAND2_X1 _u10_U7074  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18478 ) );
NAND2_X1 _u10_U7073  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18479 ) );
NAND4_X1 _u10_U7072  ( .A1(_u10_n18476 ), .A2(_u10_n18477 ), .A3(_u10_n18478 ), .A4(_u10_n18479 ), .ZN(_u10_n18475 ) );
NOR4_X1 _u10_U7071  ( .A1(_u10_n18472 ), .A2(_u10_n18473 ), .A3(_u10_n18474 ), .A4(_u10_n18475 ), .ZN(_u10_n18471 ) );
NAND2_X1 _u10_U7070  ( .A1(_u10_n18470 ), .A2(_u10_n18471 ), .ZN(am1[20]) );
NAND2_X1 _u10_U7069  ( .A1(1'b1), .A2(_u10_n12338 ), .ZN(_u10_n18466 ) );
NAND2_X1 _u10_U7068  ( .A1(1'b1), .A2(_u10_n12315 ), .ZN(_u10_n18467 ) );
NAND2_X1 _u10_U7067  ( .A1(1'b1), .A2(_u10_n12291 ), .ZN(_u10_n18468 ) );
NAND2_X1 _u10_U7066  ( .A1(1'b1), .A2(_u10_n12267 ), .ZN(_u10_n18469 ) );
NAND4_X1 _u10_U7065  ( .A1(_u10_n18466 ), .A2(_u10_n18467 ), .A3(_u10_n18468 ), .A4(_u10_n18469 ), .ZN(_u10_n18451 ) );
NAND2_X1 _u10_U7064  ( .A1(1'b1), .A2(_u10_n12242 ), .ZN(_u10_n18462 ) );
NAND2_X1 _u10_U7063  ( .A1(1'b1), .A2(_u10_n12218 ), .ZN(_u10_n18463 ) );
NAND2_X1 _u10_U7062  ( .A1(1'b1), .A2(_u10_n12195 ), .ZN(_u10_n18464 ) );
NAND2_X1 _u10_U7061  ( .A1(1'b1), .A2(_u10_n12170 ), .ZN(_u10_n18465 ) );
NAND4_X1 _u10_U7060  ( .A1(_u10_n18462 ), .A2(_u10_n18463 ), .A3(_u10_n18464 ), .A4(_u10_n18465 ), .ZN(_u10_n18452 ) );
NAND2_X1 _u10_U7059  ( .A1(1'b1), .A2(_u10_n12147 ), .ZN(_u10_n18458 ) );
NAND2_X1 _u10_U7058  ( .A1(1'b1), .A2(_u10_n12123 ), .ZN(_u10_n18459 ) );
NAND2_X1 _u10_U7057  ( .A1(1'b1), .A2(_u10_n12099 ), .ZN(_u10_n18460 ) );
NAND2_X1 _u10_U7056  ( .A1(1'b1), .A2(_u10_n12075 ), .ZN(_u10_n18461 ) );
NAND4_X1 _u10_U7055  ( .A1(_u10_n18458 ), .A2(_u10_n18459 ), .A3(_u10_n18460 ), .A4(_u10_n18461 ), .ZN(_u10_n18453 ) );
NAND2_X1 _u10_U7054  ( .A1(1'b1), .A2(_u10_n12051 ), .ZN(_u10_n18455 ) );
NAND2_X1 _u10_U7053  ( .A1(1'b1), .A2(_u10_n12027 ), .ZN(_u10_n18456 ) );
NAND2_X1 _u10_U7052  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18457 ) );
NAND3_X1 _u10_U7051  ( .A1(_u10_n18455 ), .A2(_u10_n18456 ), .A3(_u10_n18457 ), .ZN(_u10_n18454 ) );
NOR4_X1 _u10_U7050  ( .A1(_u10_n18451 ), .A2(_u10_n18452 ), .A3(_u10_n18453 ), .A4(_u10_n18454 ), .ZN(_u10_n18429 ) );
NAND2_X1 _u10_U7049  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18447 ) );
NAND2_X1 _u10_U7048  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18448 ) );
NAND2_X1 _u10_U7047  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18449 ) );
NAND2_X1 _u10_U7046  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18450 ) );
NAND4_X1 _u10_U7045  ( .A1(_u10_n18447 ), .A2(_u10_n18448 ), .A3(_u10_n18449 ), .A4(_u10_n18450 ), .ZN(_u10_n18431 ) );
NAND2_X1 _u10_U7044  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18443 ) );
NAND2_X1 _u10_U7043  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18444 ) );
NAND2_X1 _u10_U7042  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18445 ) );
NAND2_X1 _u10_U7041  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18446 ) );
NAND4_X1 _u10_U7040  ( .A1(_u10_n18443 ), .A2(_u10_n18444 ), .A3(_u10_n18445 ), .A4(_u10_n18446 ), .ZN(_u10_n18432 ) );
NAND2_X1 _u10_U7039  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18439 ) );
NAND2_X1 _u10_U7038  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18440 ) );
NAND2_X1 _u10_U7037  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18441 ) );
NAND2_X1 _u10_U7036  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18442 ) );
NAND4_X1 _u10_U7035  ( .A1(_u10_n18439 ), .A2(_u10_n18440 ), .A3(_u10_n18441 ), .A4(_u10_n18442 ), .ZN(_u10_n18433 ) );
NAND2_X1 _u10_U7034  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18435 ) );
NAND2_X1 _u10_U7033  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18436 ) );
NAND2_X1 _u10_U7032  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18437 ) );
NAND2_X1 _u10_U7031  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18438 ) );
NAND4_X1 _u10_U7030  ( .A1(_u10_n18435 ), .A2(_u10_n18436 ), .A3(_u10_n18437 ), .A4(_u10_n18438 ), .ZN(_u10_n18434 ) );
NOR4_X1 _u10_U7029  ( .A1(_u10_n18431 ), .A2(_u10_n18432 ), .A3(_u10_n18433 ), .A4(_u10_n18434 ), .ZN(_u10_n18430 ) );
NAND2_X1 _u10_U7028  ( .A1(_u10_n18429 ), .A2(_u10_n18430 ), .ZN(am1[21]) );
NAND2_X1 _u10_U7027  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18425 ) );
NAND2_X1 _u10_U7026  ( .A1(1'b1), .A2(_u10_n12329 ), .ZN(_u10_n18426 ) );
NAND2_X1 _u10_U7025  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18427 ) );
NAND2_X1 _u10_U7024  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18428 ) );
NAND4_X1 _u10_U7023  ( .A1(_u10_n18425 ), .A2(_u10_n18426 ), .A3(_u10_n18427 ), .A4(_u10_n18428 ), .ZN(_u10_n18410 ) );
NAND2_X1 _u10_U7022  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18421 ) );
NAND2_X1 _u10_U7021  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18422 ) );
NAND2_X1 _u10_U7020  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18423 ) );
NAND2_X1 _u10_U7019  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18424 ) );
NAND4_X1 _u10_U7018  ( .A1(_u10_n18421 ), .A2(_u10_n18422 ), .A3(_u10_n18423 ), .A4(_u10_n18424 ), .ZN(_u10_n18411 ) );
NAND2_X1 _u10_U7017  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18417 ) );
NAND2_X1 _u10_U7016  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18418 ) );
NAND2_X1 _u10_U7015  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18419 ) );
NAND2_X1 _u10_U7014  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18420 ) );
NAND4_X1 _u10_U7013  ( .A1(_u10_n18417 ), .A2(_u10_n18418 ), .A3(_u10_n18419 ), .A4(_u10_n18420 ), .ZN(_u10_n18412 ) );
NAND2_X1 _u10_U7012  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18414 ) );
NAND2_X1 _u10_U7011  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18415 ) );
NAND2_X1 _u10_U7010  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18416 ) );
NAND3_X1 _u10_U7009  ( .A1(_u10_n18414 ), .A2(_u10_n18415 ), .A3(_u10_n18416 ), .ZN(_u10_n18413 ) );
NOR4_X1 _u10_U7008  ( .A1(_u10_n18410 ), .A2(_u10_n18411 ), .A3(_u10_n18412 ), .A4(_u10_n18413 ), .ZN(_u10_n18388 ) );
NAND2_X1 _u10_U7007  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18406 ) );
NAND2_X1 _u10_U7006  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18407 ) );
NAND2_X1 _u10_U7005  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18408 ) );
NAND2_X1 _u10_U7004  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18409 ) );
NAND4_X1 _u10_U7003  ( .A1(_u10_n18406 ), .A2(_u10_n18407 ), .A3(_u10_n18408 ), .A4(_u10_n18409 ), .ZN(_u10_n18390 ) );
NAND2_X1 _u10_U7002  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18402 ) );
NAND2_X1 _u10_U7001  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18403 ) );
NAND2_X1 _u10_U7000  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18404 ) );
NAND2_X1 _u10_U6999  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18405 ) );
NAND4_X1 _u10_U6998  ( .A1(_u10_n18402 ), .A2(_u10_n18403 ), .A3(_u10_n18404 ), .A4(_u10_n18405 ), .ZN(_u10_n18391 ) );
NAND2_X1 _u10_U6997  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18398 ) );
NAND2_X1 _u10_U6996  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18399 ) );
NAND2_X1 _u10_U6995  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18400 ) );
NAND2_X1 _u10_U6994  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18401 ) );
NAND4_X1 _u10_U6993  ( .A1(_u10_n18398 ), .A2(_u10_n18399 ), .A3(_u10_n18400 ), .A4(_u10_n18401 ), .ZN(_u10_n18392 ) );
NAND2_X1 _u10_U6992  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18394 ) );
NAND2_X1 _u10_U6991  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18395 ) );
NAND2_X1 _u10_U6990  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18396 ) );
NAND2_X1 _u10_U6989  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18397 ) );
NAND4_X1 _u10_U6988  ( .A1(_u10_n18394 ), .A2(_u10_n18395 ), .A3(_u10_n18396 ), .A4(_u10_n18397 ), .ZN(_u10_n18393 ) );
NOR4_X1 _u10_U6987  ( .A1(_u10_n18390 ), .A2(_u10_n18391 ), .A3(_u10_n18392 ), .A4(_u10_n18393 ), .ZN(_u10_n18389 ) );
NAND2_X1 _u10_U6986  ( .A1(_u10_n18388 ), .A2(_u10_n18389 ), .ZN(am1[22]) );
NAND2_X1 _u10_U6985  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18384 ) );
NAND2_X1 _u10_U6984  ( .A1(1'b1), .A2(_u10_n12328 ), .ZN(_u10_n18385 ) );
NAND2_X1 _u10_U6983  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18386 ) );
NAND2_X1 _u10_U6982  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18387 ) );
NAND4_X1 _u10_U6981  ( .A1(_u10_n18384 ), .A2(_u10_n18385 ), .A3(_u10_n18386 ), .A4(_u10_n18387 ), .ZN(_u10_n18369 ) );
NAND2_X1 _u10_U6980  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18380 ) );
NAND2_X1 _u10_U6979  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18381 ) );
NAND2_X1 _u10_U6978  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18382 ) );
NAND2_X1 _u10_U6977  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18383 ) );
NAND4_X1 _u10_U6976  ( .A1(_u10_n18380 ), .A2(_u10_n18381 ), .A3(_u10_n18382 ), .A4(_u10_n18383 ), .ZN(_u10_n18370 ) );
NAND2_X1 _u10_U6975  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18376 ) );
NAND2_X1 _u10_U6974  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18377 ) );
NAND2_X1 _u10_U6973  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18378 ) );
NAND2_X1 _u10_U6972  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18379 ) );
NAND4_X1 _u10_U6971  ( .A1(_u10_n18376 ), .A2(_u10_n18377 ), .A3(_u10_n18378 ), .A4(_u10_n18379 ), .ZN(_u10_n18371 ) );
NAND2_X1 _u10_U6970  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18373 ) );
NAND2_X1 _u10_U6969  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18374 ) );
NAND2_X1 _u10_U6968  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18375 ) );
NAND3_X1 _u10_U6967  ( .A1(_u10_n18373 ), .A2(_u10_n18374 ), .A3(_u10_n18375 ), .ZN(_u10_n18372 ) );
NOR4_X1 _u10_U6966  ( .A1(_u10_n18369 ), .A2(_u10_n18370 ), .A3(_u10_n18371 ), .A4(_u10_n18372 ), .ZN(_u10_n18347 ) );
NAND2_X1 _u10_U6965  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18365 ) );
NAND2_X1 _u10_U6964  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18366 ) );
NAND2_X1 _u10_U6963  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18367 ) );
NAND2_X1 _u10_U6962  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18368 ) );
NAND4_X1 _u10_U6961  ( .A1(_u10_n18365 ), .A2(_u10_n18366 ), .A3(_u10_n18367 ), .A4(_u10_n18368 ), .ZN(_u10_n18349 ) );
NAND2_X1 _u10_U6960  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18361 ) );
NAND2_X1 _u10_U6959  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18362 ) );
NAND2_X1 _u10_U6958  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18363 ) );
NAND2_X1 _u10_U6957  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18364 ) );
NAND4_X1 _u10_U6956  ( .A1(_u10_n18361 ), .A2(_u10_n18362 ), .A3(_u10_n18363 ), .A4(_u10_n18364 ), .ZN(_u10_n18350 ) );
NAND2_X1 _u10_U6955  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18357 ) );
NAND2_X1 _u10_U6954  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18358 ) );
NAND2_X1 _u10_U6953  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18359 ) );
NAND2_X1 _u10_U6952  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18360 ) );
NAND4_X1 _u10_U6951  ( .A1(_u10_n18357 ), .A2(_u10_n18358 ), .A3(_u10_n18359 ), .A4(_u10_n18360 ), .ZN(_u10_n18351 ) );
NAND2_X1 _u10_U6950  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18353 ) );
NAND2_X1 _u10_U6949  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18354 ) );
NAND2_X1 _u10_U6948  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18355 ) );
NAND2_X1 _u10_U6947  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18356 ) );
NAND4_X1 _u10_U6946  ( .A1(_u10_n18353 ), .A2(_u10_n18354 ), .A3(_u10_n18355 ), .A4(_u10_n18356 ), .ZN(_u10_n18352 ) );
NOR4_X1 _u10_U6945  ( .A1(_u10_n18349 ), .A2(_u10_n18350 ), .A3(_u10_n18351 ), .A4(_u10_n18352 ), .ZN(_u10_n18348 ) );
NAND2_X1 _u10_U6944  ( .A1(_u10_n18347 ), .A2(_u10_n18348 ), .ZN(am1[23]) );
NAND2_X1 _u10_U6943  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18343 ) );
NAND2_X1 _u10_U6942  ( .A1(1'b1), .A2(_u10_n12330 ), .ZN(_u10_n18344 ) );
NAND2_X1 _u10_U6941  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18345 ) );
NAND2_X1 _u10_U6940  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18346 ) );
NAND4_X1 _u10_U6939  ( .A1(_u10_n18343 ), .A2(_u10_n18344 ), .A3(_u10_n18345 ), .A4(_u10_n18346 ), .ZN(_u10_n18328 ) );
NAND2_X1 _u10_U6938  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18339 ) );
NAND2_X1 _u10_U6937  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18340 ) );
NAND2_X1 _u10_U6936  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18341 ) );
NAND2_X1 _u10_U6935  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18342 ) );
NAND4_X1 _u10_U6934  ( .A1(_u10_n18339 ), .A2(_u10_n18340 ), .A3(_u10_n18341 ), .A4(_u10_n18342 ), .ZN(_u10_n18329 ) );
NAND2_X1 _u10_U6933  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18335 ) );
NAND2_X1 _u10_U6932  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18336 ) );
NAND2_X1 _u10_U6931  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18337 ) );
NAND2_X1 _u10_U6930  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18338 ) );
NAND4_X1 _u10_U6929  ( .A1(_u10_n18335 ), .A2(_u10_n18336 ), .A3(_u10_n18337 ), .A4(_u10_n18338 ), .ZN(_u10_n18330 ) );
NAND2_X1 _u10_U6928  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18332 ) );
NAND2_X1 _u10_U6927  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18333 ) );
NAND2_X1 _u10_U6926  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18334 ) );
NAND3_X1 _u10_U6925  ( .A1(_u10_n18332 ), .A2(_u10_n18333 ), .A3(_u10_n18334 ), .ZN(_u10_n18331 ) );
NOR4_X1 _u10_U6924  ( .A1(_u10_n18328 ), .A2(_u10_n18329 ), .A3(_u10_n18330 ), .A4(_u10_n18331 ), .ZN(_u10_n18306 ) );
NAND2_X1 _u10_U6923  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18324 ) );
NAND2_X1 _u10_U6922  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18325 ) );
NAND2_X1 _u10_U6921  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18326 ) );
NAND2_X1 _u10_U6920  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18327 ) );
NAND4_X1 _u10_U6919  ( .A1(_u10_n18324 ), .A2(_u10_n18325 ), .A3(_u10_n18326 ), .A4(_u10_n18327 ), .ZN(_u10_n18308 ) );
NAND2_X1 _u10_U6918  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18320 ) );
NAND2_X1 _u10_U6917  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18321 ) );
NAND2_X1 _u10_U6916  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18322 ) );
NAND2_X1 _u10_U6915  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18323 ) );
NAND4_X1 _u10_U6914  ( .A1(_u10_n18320 ), .A2(_u10_n18321 ), .A3(_u10_n18322 ), .A4(_u10_n18323 ), .ZN(_u10_n18309 ) );
NAND2_X1 _u10_U6913  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18316 ) );
NAND2_X1 _u10_U6912  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18317 ) );
NAND2_X1 _u10_U6911  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18318 ) );
NAND2_X1 _u10_U6910  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18319 ) );
NAND4_X1 _u10_U6909  ( .A1(_u10_n18316 ), .A2(_u10_n18317 ), .A3(_u10_n18318 ), .A4(_u10_n18319 ), .ZN(_u10_n18310 ) );
NAND2_X1 _u10_U6908  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18312 ) );
NAND2_X1 _u10_U6907  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18313 ) );
NAND2_X1 _u10_U6906  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18314 ) );
NAND2_X1 _u10_U6905  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18315 ) );
NAND4_X1 _u10_U6904  ( .A1(_u10_n18312 ), .A2(_u10_n18313 ), .A3(_u10_n18314 ), .A4(_u10_n18315 ), .ZN(_u10_n18311 ) );
NOR4_X1 _u10_U6903  ( .A1(_u10_n18308 ), .A2(_u10_n18309 ), .A3(_u10_n18310 ), .A4(_u10_n18311 ), .ZN(_u10_n18307 ) );
NAND2_X1 _u10_U6902  ( .A1(_u10_n18306 ), .A2(_u10_n18307 ), .ZN(am1[24]) );
NAND2_X1 _u10_U6901  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18302 ) );
NAND2_X1 _u10_U6900  ( .A1(1'b1), .A2(_u10_n12331 ), .ZN(_u10_n18303 ) );
NAND2_X1 _u10_U6899  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18304 ) );
NAND2_X1 _u10_U6898  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18305 ) );
NAND4_X1 _u10_U6897  ( .A1(_u10_n18302 ), .A2(_u10_n18303 ), .A3(_u10_n18304 ), .A4(_u10_n18305 ), .ZN(_u10_n18287 ) );
NAND2_X1 _u10_U6896  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18298 ) );
NAND2_X1 _u10_U6895  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18299 ) );
NAND2_X1 _u10_U6894  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18300 ) );
NAND2_X1 _u10_U6893  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18301 ) );
NAND4_X1 _u10_U6892  ( .A1(_u10_n18298 ), .A2(_u10_n18299 ), .A3(_u10_n18300 ), .A4(_u10_n18301 ), .ZN(_u10_n18288 ) );
NAND2_X1 _u10_U6891  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18294 ) );
NAND2_X1 _u10_U6890  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18295 ) );
NAND2_X1 _u10_U6889  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18296 ) );
NAND2_X1 _u10_U6888  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18297 ) );
NAND4_X1 _u10_U6887  ( .A1(_u10_n18294 ), .A2(_u10_n18295 ), .A3(_u10_n18296 ), .A4(_u10_n18297 ), .ZN(_u10_n18289 ) );
NAND2_X1 _u10_U6886  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18291 ) );
NAND2_X1 _u10_U6885  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18292 ) );
NAND2_X1 _u10_U6884  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18293 ) );
NAND3_X1 _u10_U6883  ( .A1(_u10_n18291 ), .A2(_u10_n18292 ), .A3(_u10_n18293 ), .ZN(_u10_n18290 ) );
NOR4_X1 _u10_U6882  ( .A1(_u10_n18287 ), .A2(_u10_n18288 ), .A3(_u10_n18289 ), .A4(_u10_n18290 ), .ZN(_u10_n18265 ) );
NAND2_X1 _u10_U6881  ( .A1(1'b1), .A2(_u10_n11991 ), .ZN(_u10_n18283 ) );
NAND2_X1 _u10_U6880  ( .A1(1'b1), .A2(_u10_n11967 ), .ZN(_u10_n18284 ) );
NAND2_X1 _u10_U6879  ( .A1(1'b1), .A2(_u10_n11943 ), .ZN(_u10_n18285 ) );
NAND2_X1 _u10_U6878  ( .A1(1'b1), .A2(_u10_n11919 ), .ZN(_u10_n18286 ) );
NAND4_X1 _u10_U6877  ( .A1(_u10_n18283 ), .A2(_u10_n18284 ), .A3(_u10_n18285 ), .A4(_u10_n18286 ), .ZN(_u10_n18267 ) );
NAND2_X1 _u10_U6876  ( .A1(1'b1), .A2(_u10_n11895 ), .ZN(_u10_n18279 ) );
NAND2_X1 _u10_U6875  ( .A1(1'b1), .A2(_u10_n11871 ), .ZN(_u10_n18280 ) );
NAND2_X1 _u10_U6874  ( .A1(1'b1), .A2(_u10_n11847 ), .ZN(_u10_n18281 ) );
NAND2_X1 _u10_U6873  ( .A1(1'b1), .A2(_u10_n11823 ), .ZN(_u10_n18282 ) );
NAND4_X1 _u10_U6872  ( .A1(_u10_n18279 ), .A2(_u10_n18280 ), .A3(_u10_n18281 ), .A4(_u10_n18282 ), .ZN(_u10_n18268 ) );
NAND2_X1 _u10_U6871  ( .A1(1'b1), .A2(_u10_n11799 ), .ZN(_u10_n18275 ) );
NAND2_X1 _u10_U6870  ( .A1(1'b1), .A2(_u10_n11775 ), .ZN(_u10_n18276 ) );
NAND2_X1 _u10_U6869  ( .A1(1'b1), .A2(_u10_n11751 ), .ZN(_u10_n18277 ) );
NAND2_X1 _u10_U6868  ( .A1(1'b1), .A2(_u10_n11727 ), .ZN(_u10_n18278 ) );
NAND4_X1 _u10_U6867  ( .A1(_u10_n18275 ), .A2(_u10_n18276 ), .A3(_u10_n18277 ), .A4(_u10_n18278 ), .ZN(_u10_n18269 ) );
NAND2_X1 _u10_U6866  ( .A1(1'b1), .A2(_u10_n11703 ), .ZN(_u10_n18271 ) );
NAND2_X1 _u10_U6865  ( .A1(1'b1), .A2(_u10_n11679 ), .ZN(_u10_n18272 ) );
NAND2_X1 _u10_U6864  ( .A1(1'b1), .A2(_u10_n11655 ), .ZN(_u10_n18273 ) );
NAND2_X1 _u10_U6863  ( .A1(1'b1), .A2(_u10_n11631 ), .ZN(_u10_n18274 ) );
NAND4_X1 _u10_U6862  ( .A1(_u10_n18271 ), .A2(_u10_n18272 ), .A3(_u10_n18273 ), .A4(_u10_n18274 ), .ZN(_u10_n18270 ) );
NOR4_X1 _u10_U6861  ( .A1(_u10_n18267 ), .A2(_u10_n18268 ), .A3(_u10_n18269 ), .A4(_u10_n18270 ), .ZN(_u10_n18266 ) );
NAND2_X1 _u10_U6860  ( .A1(_u10_n18265 ), .A2(_u10_n18266 ), .ZN(am1[25]) );
NAND2_X1 _u10_U6859  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18261 ) );
NAND2_X1 _u10_U6858  ( .A1(1'b1), .A2(_u10_n12429 ), .ZN(_u10_n18262 ) );
NAND2_X1 _u10_U6857  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18263 ) );
NAND2_X1 _u10_U6856  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18264 ) );
NAND4_X1 _u10_U6855  ( .A1(_u10_n18261 ), .A2(_u10_n18262 ), .A3(_u10_n18263 ), .A4(_u10_n18264 ), .ZN(_u10_n18246 ) );
NAND2_X1 _u10_U6854  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18257 ) );
NAND2_X1 _u10_U6853  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18258 ) );
NAND2_X1 _u10_U6852  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18259 ) );
NAND2_X1 _u10_U6851  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18260 ) );
NAND4_X1 _u10_U6850  ( .A1(_u10_n18257 ), .A2(_u10_n18258 ), .A3(_u10_n18259 ), .A4(_u10_n18260 ), .ZN(_u10_n18247 ) );
NAND2_X1 _u10_U6849  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18253 ) );
NAND2_X1 _u10_U6848  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18254 ) );
NAND2_X1 _u10_U6847  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18255 ) );
NAND2_X1 _u10_U6846  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18256 ) );
NAND4_X1 _u10_U6845  ( .A1(_u10_n18253 ), .A2(_u10_n18254 ), .A3(_u10_n18255 ), .A4(_u10_n18256 ), .ZN(_u10_n18248 ) );
NAND2_X1 _u10_U6844  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18250 ) );
NAND2_X1 _u10_U6843  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18251 ) );
NAND2_X1 _u10_U6842  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18252 ) );
NAND3_X1 _u10_U6841  ( .A1(_u10_n18250 ), .A2(_u10_n18251 ), .A3(_u10_n18252 ), .ZN(_u10_n18249 ) );
NOR4_X1 _u10_U6840  ( .A1(_u10_n18246 ), .A2(_u10_n18247 ), .A3(_u10_n18248 ), .A4(_u10_n18249 ), .ZN(_u10_n18224 ) );
NAND2_X1 _u10_U6839  ( .A1(1'b1), .A2(_u10_n11992 ), .ZN(_u10_n18242 ) );
NAND2_X1 _u10_U6838  ( .A1(1'b1), .A2(_u10_n11968 ), .ZN(_u10_n18243 ) );
NAND2_X1 _u10_U6837  ( .A1(1'b1), .A2(_u10_n11944 ), .ZN(_u10_n18244 ) );
NAND2_X1 _u10_U6836  ( .A1(1'b1), .A2(_u10_n11920 ), .ZN(_u10_n18245 ) );
NAND4_X1 _u10_U6835  ( .A1(_u10_n18242 ), .A2(_u10_n18243 ), .A3(_u10_n18244 ), .A4(_u10_n18245 ), .ZN(_u10_n18226 ) );
NAND2_X1 _u10_U6834  ( .A1(1'b1), .A2(_u10_n11896 ), .ZN(_u10_n18238 ) );
NAND2_X1 _u10_U6833  ( .A1(1'b1), .A2(_u10_n11872 ), .ZN(_u10_n18239 ) );
NAND2_X1 _u10_U6832  ( .A1(1'b1), .A2(_u10_n11848 ), .ZN(_u10_n18240 ) );
NAND2_X1 _u10_U6831  ( .A1(1'b1), .A2(_u10_n11824 ), .ZN(_u10_n18241 ) );
NAND4_X1 _u10_U6830  ( .A1(_u10_n18238 ), .A2(_u10_n18239 ), .A3(_u10_n18240 ), .A4(_u10_n18241 ), .ZN(_u10_n18227 ) );
NAND2_X1 _u10_U6829  ( .A1(1'b1), .A2(_u10_n11800 ), .ZN(_u10_n18234 ) );
NAND2_X1 _u10_U6828  ( .A1(1'b1), .A2(_u10_n11776 ), .ZN(_u10_n18235 ) );
NAND2_X1 _u10_U6827  ( .A1(1'b1), .A2(_u10_n11752 ), .ZN(_u10_n18236 ) );
NAND2_X1 _u10_U6826  ( .A1(1'b1), .A2(_u10_n11728 ), .ZN(_u10_n18237 ) );
NAND4_X1 _u10_U6825  ( .A1(_u10_n18234 ), .A2(_u10_n18235 ), .A3(_u10_n18236 ), .A4(_u10_n18237 ), .ZN(_u10_n18228 ) );
NAND2_X1 _u10_U6824  ( .A1(1'b1), .A2(_u10_n11704 ), .ZN(_u10_n18230 ) );
NAND2_X1 _u10_U6823  ( .A1(1'b1), .A2(_u10_n11680 ), .ZN(_u10_n18231 ) );
NAND2_X1 _u10_U6822  ( .A1(1'b1), .A2(_u10_n11656 ), .ZN(_u10_n18232 ) );
NAND2_X1 _u10_U6821  ( .A1(1'b1), .A2(_u10_n11632 ), .ZN(_u10_n18233 ) );
NAND4_X1 _u10_U6820  ( .A1(_u10_n18230 ), .A2(_u10_n18231 ), .A3(_u10_n18232 ), .A4(_u10_n18233 ), .ZN(_u10_n18229 ) );
NOR4_X1 _u10_U6819  ( .A1(_u10_n18226 ), .A2(_u10_n18227 ), .A3(_u10_n18228 ), .A4(_u10_n18229 ), .ZN(_u10_n18225 ) );
NAND2_X1 _u10_U6818  ( .A1(_u10_n18224 ), .A2(_u10_n18225 ), .ZN(am1[26]) );
NAND2_X1 _u10_U6817  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18220 ) );
NAND2_X1 _u10_U6816  ( .A1(1'b1), .A2(_u10_n12332 ), .ZN(_u10_n18221 ) );
NAND2_X1 _u10_U6815  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18222 ) );
NAND2_X1 _u10_U6814  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18223 ) );
NAND4_X1 _u10_U6813  ( .A1(_u10_n18220 ), .A2(_u10_n18221 ), .A3(_u10_n18222 ), .A4(_u10_n18223 ), .ZN(_u10_n18205 ) );
NAND2_X1 _u10_U6812  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18216 ) );
NAND2_X1 _u10_U6811  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18217 ) );
NAND2_X1 _u10_U6810  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18218 ) );
NAND2_X1 _u10_U6809  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18219 ) );
NAND4_X1 _u10_U6808  ( .A1(_u10_n18216 ), .A2(_u10_n18217 ), .A3(_u10_n18218 ), .A4(_u10_n18219 ), .ZN(_u10_n18206 ) );
NAND2_X1 _u10_U6807  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18212 ) );
NAND2_X1 _u10_U6806  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18213 ) );
NAND2_X1 _u10_U6805  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18214 ) );
NAND2_X1 _u10_U6804  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18215 ) );
NAND4_X1 _u10_U6803  ( .A1(_u10_n18212 ), .A2(_u10_n18213 ), .A3(_u10_n18214 ), .A4(_u10_n18215 ), .ZN(_u10_n18207 ) );
NAND2_X1 _u10_U6802  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18209 ) );
NAND2_X1 _u10_U6801  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18210 ) );
NAND2_X1 _u10_U6800  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18211 ) );
NAND3_X1 _u10_U6799  ( .A1(_u10_n18209 ), .A2(_u10_n18210 ), .A3(_u10_n18211 ), .ZN(_u10_n18208 ) );
NOR4_X1 _u10_U6798  ( .A1(_u10_n18205 ), .A2(_u10_n18206 ), .A3(_u10_n18207 ), .A4(_u10_n18208 ), .ZN(_u10_n18183 ) );
NAND2_X1 _u10_U6797  ( .A1(1'b1), .A2(_u10_n11992 ), .ZN(_u10_n18201 ) );
NAND2_X1 _u10_U6796  ( .A1(1'b1), .A2(_u10_n11968 ), .ZN(_u10_n18202 ) );
NAND2_X1 _u10_U6795  ( .A1(1'b1), .A2(_u10_n11944 ), .ZN(_u10_n18203 ) );
NAND2_X1 _u10_U6794  ( .A1(1'b1), .A2(_u10_n11920 ), .ZN(_u10_n18204 ) );
NAND4_X1 _u10_U6793  ( .A1(_u10_n18201 ), .A2(_u10_n18202 ), .A3(_u10_n18203 ), .A4(_u10_n18204 ), .ZN(_u10_n18185 ) );
NAND2_X1 _u10_U6792  ( .A1(1'b1), .A2(_u10_n11896 ), .ZN(_u10_n18197 ) );
NAND2_X1 _u10_U6791  ( .A1(1'b1), .A2(_u10_n11872 ), .ZN(_u10_n18198 ) );
NAND2_X1 _u10_U6790  ( .A1(1'b1), .A2(_u10_n11848 ), .ZN(_u10_n18199 ) );
NAND2_X1 _u10_U6789  ( .A1(1'b1), .A2(_u10_n11824 ), .ZN(_u10_n18200 ) );
NAND4_X1 _u10_U6788  ( .A1(_u10_n18197 ), .A2(_u10_n18198 ), .A3(_u10_n18199 ), .A4(_u10_n18200 ), .ZN(_u10_n18186 ) );
NAND2_X1 _u10_U6787  ( .A1(1'b1), .A2(_u10_n11800 ), .ZN(_u10_n18193 ) );
NAND2_X1 _u10_U6786  ( .A1(1'b1), .A2(_u10_n11776 ), .ZN(_u10_n18194 ) );
NAND2_X1 _u10_U6785  ( .A1(1'b1), .A2(_u10_n11752 ), .ZN(_u10_n18195 ) );
NAND2_X1 _u10_U6784  ( .A1(1'b1), .A2(_u10_n11728 ), .ZN(_u10_n18196 ) );
NAND4_X1 _u10_U6783  ( .A1(_u10_n18193 ), .A2(_u10_n18194 ), .A3(_u10_n18195 ), .A4(_u10_n18196 ), .ZN(_u10_n18187 ) );
NAND2_X1 _u10_U6782  ( .A1(1'b1), .A2(_u10_n11704 ), .ZN(_u10_n18189 ) );
NAND2_X1 _u10_U6781  ( .A1(1'b1), .A2(_u10_n11680 ), .ZN(_u10_n18190 ) );
NAND2_X1 _u10_U6780  ( .A1(1'b1), .A2(_u10_n11656 ), .ZN(_u10_n18191 ) );
NAND2_X1 _u10_U6779  ( .A1(1'b1), .A2(_u10_n11632 ), .ZN(_u10_n18192 ) );
NAND4_X1 _u10_U6778  ( .A1(_u10_n18189 ), .A2(_u10_n18190 ), .A3(_u10_n18191 ), .A4(_u10_n18192 ), .ZN(_u10_n18188 ) );
NOR4_X1 _u10_U6777  ( .A1(_u10_n18185 ), .A2(_u10_n18186 ), .A3(_u10_n18187 ), .A4(_u10_n18188 ), .ZN(_u10_n18184 ) );
NAND2_X1 _u10_U6776  ( .A1(_u10_n18183 ), .A2(_u10_n18184 ), .ZN(am1[27]) );
NAND2_X1 _u10_U6775  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18179 ) );
NAND2_X1 _u10_U6774  ( .A1(1'b1), .A2(_u10_n12329 ), .ZN(_u10_n18180 ) );
NAND2_X1 _u10_U6773  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18181 ) );
NAND2_X1 _u10_U6772  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18182 ) );
NAND4_X1 _u10_U6771  ( .A1(_u10_n18179 ), .A2(_u10_n18180 ), .A3(_u10_n18181 ), .A4(_u10_n18182 ), .ZN(_u10_n18164 ) );
NAND2_X1 _u10_U6770  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18175 ) );
NAND2_X1 _u10_U6769  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18176 ) );
NAND2_X1 _u10_U6768  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18177 ) );
NAND2_X1 _u10_U6767  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18178 ) );
NAND4_X1 _u10_U6766  ( .A1(_u10_n18175 ), .A2(_u10_n18176 ), .A3(_u10_n18177 ), .A4(_u10_n18178 ), .ZN(_u10_n18165 ) );
NAND2_X1 _u10_U6765  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18171 ) );
NAND2_X1 _u10_U6764  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18172 ) );
NAND2_X1 _u10_U6763  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18173 ) );
NAND2_X1 _u10_U6762  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18174 ) );
NAND4_X1 _u10_U6761  ( .A1(_u10_n18171 ), .A2(_u10_n18172 ), .A3(_u10_n18173 ), .A4(_u10_n18174 ), .ZN(_u10_n18166 ) );
NAND2_X1 _u10_U6760  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18168 ) );
NAND2_X1 _u10_U6759  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18169 ) );
NAND2_X1 _u10_U6758  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18170 ) );
NAND3_X1 _u10_U6757  ( .A1(_u10_n18168 ), .A2(_u10_n18169 ), .A3(_u10_n18170 ), .ZN(_u10_n18167 ) );
NOR4_X1 _u10_U6756  ( .A1(_u10_n18164 ), .A2(_u10_n18165 ), .A3(_u10_n18166 ), .A4(_u10_n18167 ), .ZN(_u10_n18142 ) );
NAND2_X1 _u10_U6755  ( .A1(1'b1), .A2(_u10_n11992 ), .ZN(_u10_n18160 ) );
NAND2_X1 _u10_U6754  ( .A1(1'b1), .A2(_u10_n11968 ), .ZN(_u10_n18161 ) );
NAND2_X1 _u10_U6753  ( .A1(1'b1), .A2(_u10_n11944 ), .ZN(_u10_n18162 ) );
NAND2_X1 _u10_U6752  ( .A1(1'b1), .A2(_u10_n11920 ), .ZN(_u10_n18163 ) );
NAND4_X1 _u10_U6751  ( .A1(_u10_n18160 ), .A2(_u10_n18161 ), .A3(_u10_n18162 ), .A4(_u10_n18163 ), .ZN(_u10_n18144 ) );
NAND2_X1 _u10_U6750  ( .A1(1'b1), .A2(_u10_n11896 ), .ZN(_u10_n18156 ) );
NAND2_X1 _u10_U6749  ( .A1(1'b1), .A2(_u10_n11872 ), .ZN(_u10_n18157 ) );
NAND2_X1 _u10_U6748  ( .A1(1'b1), .A2(_u10_n11848 ), .ZN(_u10_n18158 ) );
NAND2_X1 _u10_U6747  ( .A1(1'b1), .A2(_u10_n11824 ), .ZN(_u10_n18159 ) );
NAND4_X1 _u10_U6746  ( .A1(_u10_n18156 ), .A2(_u10_n18157 ), .A3(_u10_n18158 ), .A4(_u10_n18159 ), .ZN(_u10_n18145 ) );
NAND2_X1 _u10_U6745  ( .A1(1'b1), .A2(_u10_n11800 ), .ZN(_u10_n18152 ) );
NAND2_X1 _u10_U6744  ( .A1(1'b1), .A2(_u10_n11776 ), .ZN(_u10_n18153 ) );
NAND2_X1 _u10_U6743  ( .A1(1'b1), .A2(_u10_n11752 ), .ZN(_u10_n18154 ) );
NAND2_X1 _u10_U6742  ( .A1(1'b1), .A2(_u10_n11728 ), .ZN(_u10_n18155 ) );
NAND4_X1 _u10_U6741  ( .A1(_u10_n18152 ), .A2(_u10_n18153 ), .A3(_u10_n18154 ), .A4(_u10_n18155 ), .ZN(_u10_n18146 ) );
NAND2_X1 _u10_U6740  ( .A1(1'b1), .A2(_u10_n11704 ), .ZN(_u10_n18148 ) );
NAND2_X1 _u10_U6739  ( .A1(1'b1), .A2(_u10_n11680 ), .ZN(_u10_n18149 ) );
NAND2_X1 _u10_U6738  ( .A1(1'b1), .A2(_u10_n11656 ), .ZN(_u10_n18150 ) );
NAND2_X1 _u10_U6737  ( .A1(1'b1), .A2(_u10_n11632 ), .ZN(_u10_n18151 ) );
NAND4_X1 _u10_U6736  ( .A1(_u10_n18148 ), .A2(_u10_n18149 ), .A3(_u10_n18150 ), .A4(_u10_n18151 ), .ZN(_u10_n18147 ) );
NOR4_X1 _u10_U6735  ( .A1(_u10_n18144 ), .A2(_u10_n18145 ), .A3(_u10_n18146 ), .A4(_u10_n18147 ), .ZN(_u10_n18143 ) );
NAND2_X1 _u10_U6734  ( .A1(_u10_n18142 ), .A2(_u10_n18143 ), .ZN(am1[28]) );
NAND2_X1 _u10_U6733  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18138 ) );
NAND2_X1 _u10_U6732  ( .A1(1'b1), .A2(_u10_n12328 ), .ZN(_u10_n18139 ) );
NAND2_X1 _u10_U6731  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18140 ) );
NAND2_X1 _u10_U6730  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18141 ) );
NAND4_X1 _u10_U6729  ( .A1(_u10_n18138 ), .A2(_u10_n18139 ), .A3(_u10_n18140 ), .A4(_u10_n18141 ), .ZN(_u10_n18123 ) );
NAND2_X1 _u10_U6728  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18134 ) );
NAND2_X1 _u10_U6727  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18135 ) );
NAND2_X1 _u10_U6726  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18136 ) );
NAND2_X1 _u10_U6725  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18137 ) );
NAND4_X1 _u10_U6724  ( .A1(_u10_n18134 ), .A2(_u10_n18135 ), .A3(_u10_n18136 ), .A4(_u10_n18137 ), .ZN(_u10_n18124 ) );
NAND2_X1 _u10_U6723  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18130 ) );
NAND2_X1 _u10_U6722  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18131 ) );
NAND2_X1 _u10_U6721  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18132 ) );
NAND2_X1 _u10_U6720  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18133 ) );
NAND4_X1 _u10_U6719  ( .A1(_u10_n18130 ), .A2(_u10_n18131 ), .A3(_u10_n18132 ), .A4(_u10_n18133 ), .ZN(_u10_n18125 ) );
NAND2_X1 _u10_U6718  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18127 ) );
NAND2_X1 _u10_U6717  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18128 ) );
NAND2_X1 _u10_U6716  ( .A1(1'b1), .A2(_u10_n12008 ), .ZN(_u10_n18129 ) );
NAND3_X1 _u10_U6715  ( .A1(_u10_n18127 ), .A2(_u10_n18128 ), .A3(_u10_n18129 ), .ZN(_u10_n18126 ) );
NOR4_X1 _u10_U6714  ( .A1(_u10_n18123 ), .A2(_u10_n18124 ), .A3(_u10_n18125 ), .A4(_u10_n18126 ), .ZN(_u10_n18101 ) );
NAND2_X1 _u10_U6713  ( .A1(1'b1), .A2(_u10_n11992 ), .ZN(_u10_n18119 ) );
NAND2_X1 _u10_U6712  ( .A1(1'b1), .A2(_u10_n11968 ), .ZN(_u10_n18120 ) );
NAND2_X1 _u10_U6711  ( .A1(1'b1), .A2(_u10_n11944 ), .ZN(_u10_n18121 ) );
NAND2_X1 _u10_U6710  ( .A1(1'b1), .A2(_u10_n11920 ), .ZN(_u10_n18122 ) );
NAND4_X1 _u10_U6709  ( .A1(_u10_n18119 ), .A2(_u10_n18120 ), .A3(_u10_n18121 ), .A4(_u10_n18122 ), .ZN(_u10_n18103 ) );
NAND2_X1 _u10_U6708  ( .A1(1'b1), .A2(_u10_n11896 ), .ZN(_u10_n18115 ) );
NAND2_X1 _u10_U6707  ( .A1(1'b1), .A2(_u10_n11872 ), .ZN(_u10_n18116 ) );
NAND2_X1 _u10_U6706  ( .A1(1'b1), .A2(_u10_n11848 ), .ZN(_u10_n18117 ) );
NAND2_X1 _u10_U6705  ( .A1(1'b1), .A2(_u10_n11824 ), .ZN(_u10_n18118 ) );
NAND4_X1 _u10_U6704  ( .A1(_u10_n18115 ), .A2(_u10_n18116 ), .A3(_u10_n18117 ), .A4(_u10_n18118 ), .ZN(_u10_n18104 ) );
NAND2_X1 _u10_U6703  ( .A1(1'b1), .A2(_u10_n11800 ), .ZN(_u10_n18111 ) );
NAND2_X1 _u10_U6702  ( .A1(1'b1), .A2(_u10_n11776 ), .ZN(_u10_n18112 ) );
NAND2_X1 _u10_U6701  ( .A1(1'b1), .A2(_u10_n11752 ), .ZN(_u10_n18113 ) );
NAND2_X1 _u10_U6700  ( .A1(1'b1), .A2(_u10_n11728 ), .ZN(_u10_n18114 ) );
NAND4_X1 _u10_U6699  ( .A1(_u10_n18111 ), .A2(_u10_n18112 ), .A3(_u10_n18113 ), .A4(_u10_n18114 ), .ZN(_u10_n18105 ) );
NAND2_X1 _u10_U6698  ( .A1(1'b1), .A2(_u10_n11704 ), .ZN(_u10_n18107 ) );
NAND2_X1 _u10_U6697  ( .A1(1'b1), .A2(_u10_n11680 ), .ZN(_u10_n18108 ) );
NAND2_X1 _u10_U6696  ( .A1(1'b1), .A2(_u10_n11656 ), .ZN(_u10_n18109 ) );
NAND2_X1 _u10_U6695  ( .A1(1'b1), .A2(_u10_n11632 ), .ZN(_u10_n18110 ) );
NAND4_X1 _u10_U6694  ( .A1(_u10_n18107 ), .A2(_u10_n18108 ), .A3(_u10_n18109 ), .A4(_u10_n18110 ), .ZN(_u10_n18106 ) );
NOR4_X1 _u10_U6693  ( .A1(_u10_n18103 ), .A2(_u10_n18104 ), .A3(_u10_n18105 ), .A4(_u10_n18106 ), .ZN(_u10_n18102 ) );
NAND2_X1 _u10_U6692  ( .A1(_u10_n18101 ), .A2(_u10_n18102 ), .ZN(am1[29]) );
NAND2_X1 _u10_U6691  ( .A1(1'b0), .A2(_u10_n12339 ), .ZN(_u10_n18097 ) );
NAND2_X1 _u10_U6690  ( .A1(1'b0), .A2(_u10_n12330 ), .ZN(_u10_n18098 ) );
NAND2_X1 _u10_U6689  ( .A1(1'b0), .A2(_u10_n12292 ), .ZN(_u10_n18099 ) );
NAND2_X1 _u10_U6688  ( .A1(1'b0), .A2(_u10_n12268 ), .ZN(_u10_n18100 ) );
NAND4_X1 _u10_U6687  ( .A1(_u10_n18097 ), .A2(_u10_n18098 ), .A3(_u10_n18099 ), .A4(_u10_n18100 ), .ZN(_u10_n18082 ) );
NAND2_X1 _u10_U6686  ( .A1(1'b0), .A2(_u10_n12243 ), .ZN(_u10_n18093 ) );
NAND2_X1 _u10_U6685  ( .A1(1'b0), .A2(_u10_n12219 ), .ZN(_u10_n18094 ) );
NAND2_X1 _u10_U6684  ( .A1(1'b0), .A2(_u10_n12196 ), .ZN(_u10_n18095 ) );
NAND2_X1 _u10_U6683  ( .A1(1'b0), .A2(_u10_n12171 ), .ZN(_u10_n18096 ) );
NAND4_X1 _u10_U6682  ( .A1(_u10_n18093 ), .A2(_u10_n18094 ), .A3(_u10_n18095 ), .A4(_u10_n18096 ), .ZN(_u10_n18083 ) );
NAND2_X1 _u10_U6681  ( .A1(1'b0), .A2(_u10_n12148 ), .ZN(_u10_n18089 ) );
NAND2_X1 _u10_U6680  ( .A1(1'b0), .A2(_u10_n12124 ), .ZN(_u10_n18090 ) );
NAND2_X1 _u10_U6679  ( .A1(1'b0), .A2(_u10_n12100 ), .ZN(_u10_n18091 ) );
NAND2_X1 _u10_U6678  ( .A1(1'b0), .A2(_u10_n12076 ), .ZN(_u10_n18092 ) );
NAND4_X1 _u10_U6677  ( .A1(_u10_n18089 ), .A2(_u10_n18090 ), .A3(_u10_n18091 ), .A4(_u10_n18092 ), .ZN(_u10_n18084 ) );
NAND2_X1 _u10_U6676  ( .A1(1'b0), .A2(_u10_n12052 ), .ZN(_u10_n18086 ) );
NAND2_X1 _u10_U6675  ( .A1(1'b0), .A2(_u10_n12028 ), .ZN(_u10_n18087 ) );
NAND2_X1 _u10_U6674  ( .A1(1'b0), .A2(_u10_n12008 ), .ZN(_u10_n18088 ) );
NAND3_X1 _u10_U6673  ( .A1(_u10_n18086 ), .A2(_u10_n18087 ), .A3(_u10_n18088 ), .ZN(_u10_n18085 ) );
NOR4_X1 _u10_U6672  ( .A1(_u10_n18082 ), .A2(_u10_n18083 ), .A3(_u10_n18084 ), .A4(_u10_n18085 ), .ZN(_u10_n18060 ) );
NAND2_X1 _u10_U6671  ( .A1(1'b0), .A2(_u10_n11992 ), .ZN(_u10_n18078 ) );
NAND2_X1 _u10_U6670  ( .A1(1'b0), .A2(_u10_n11968 ), .ZN(_u10_n18079 ) );
NAND2_X1 _u10_U6669  ( .A1(1'b0), .A2(_u10_n11944 ), .ZN(_u10_n18080 ) );
NAND2_X1 _u10_U6668  ( .A1(1'b0), .A2(_u10_n11920 ), .ZN(_u10_n18081 ) );
NAND4_X1 _u10_U6667  ( .A1(_u10_n18078 ), .A2(_u10_n18079 ), .A3(_u10_n18080 ), .A4(_u10_n18081 ), .ZN(_u10_n18062 ) );
NAND2_X1 _u10_U6666  ( .A1(1'b0), .A2(_u10_n11896 ), .ZN(_u10_n18074 ) );
NAND2_X1 _u10_U6665  ( .A1(1'b0), .A2(_u10_n11872 ), .ZN(_u10_n18075 ) );
NAND2_X1 _u10_U6664  ( .A1(1'b0), .A2(_u10_n11848 ), .ZN(_u10_n18076 ) );
NAND2_X1 _u10_U6663  ( .A1(1'b0), .A2(_u10_n11824 ), .ZN(_u10_n18077 ) );
NAND4_X1 _u10_U6662  ( .A1(_u10_n18074 ), .A2(_u10_n18075 ), .A3(_u10_n18076 ), .A4(_u10_n18077 ), .ZN(_u10_n18063 ) );
NAND2_X1 _u10_U6661  ( .A1(1'b0), .A2(_u10_n11800 ), .ZN(_u10_n18070 ) );
NAND2_X1 _u10_U6660  ( .A1(1'b0), .A2(_u10_n11776 ), .ZN(_u10_n18071 ) );
NAND2_X1 _u10_U6659  ( .A1(1'b0), .A2(_u10_n11752 ), .ZN(_u10_n18072 ) );
NAND2_X1 _u10_U6658  ( .A1(1'b0), .A2(_u10_n11728 ), .ZN(_u10_n18073 ) );
NAND4_X1 _u10_U6657  ( .A1(_u10_n18070 ), .A2(_u10_n18071 ), .A3(_u10_n18072 ), .A4(_u10_n18073 ), .ZN(_u10_n18064 ) );
NAND2_X1 _u10_U6656  ( .A1(1'b0), .A2(_u10_n11704 ), .ZN(_u10_n18066 ) );
NAND2_X1 _u10_U6655  ( .A1(1'b0), .A2(_u10_n11680 ), .ZN(_u10_n18067 ) );
NAND2_X1 _u10_U6654  ( .A1(1'b0), .A2(_u10_n11656 ), .ZN(_u10_n18068 ) );
NAND2_X1 _u10_U6653  ( .A1(1'b0), .A2(_u10_n11632 ), .ZN(_u10_n18069 ) );
NAND4_X1 _u10_U6652  ( .A1(_u10_n18066 ), .A2(_u10_n18067 ), .A3(_u10_n18068 ), .A4(_u10_n18069 ), .ZN(_u10_n18065 ) );
NOR4_X1 _u10_U6651  ( .A1(_u10_n18062 ), .A2(_u10_n18063 ), .A3(_u10_n18064 ), .A4(_u10_n18065 ), .ZN(_u10_n18061 ) );
NAND2_X1 _u10_U6650  ( .A1(_u10_n18060 ), .A2(_u10_n18061 ), .ZN(am1[2]) );
NAND2_X1 _u10_U6649  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18056 ) );
NAND2_X1 _u10_U6648  ( .A1(1'b1), .A2(_u10_n12331 ), .ZN(_u10_n18057 ) );
NAND2_X1 _u10_U6647  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18058 ) );
NAND2_X1 _u10_U6646  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18059 ) );
NAND4_X1 _u10_U6645  ( .A1(_u10_n18056 ), .A2(_u10_n18057 ), .A3(_u10_n18058 ), .A4(_u10_n18059 ), .ZN(_u10_n18041 ) );
NAND2_X1 _u10_U6644  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18052 ) );
NAND2_X1 _u10_U6643  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18053 ) );
NAND2_X1 _u10_U6642  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18054 ) );
NAND2_X1 _u10_U6641  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18055 ) );
NAND4_X1 _u10_U6640  ( .A1(_u10_n18052 ), .A2(_u10_n18053 ), .A3(_u10_n18054 ), .A4(_u10_n18055 ), .ZN(_u10_n18042 ) );
NAND2_X1 _u10_U6639  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18048 ) );
NAND2_X1 _u10_U6638  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18049 ) );
NAND2_X1 _u10_U6637  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18050 ) );
NAND2_X1 _u10_U6636  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18051 ) );
NAND4_X1 _u10_U6635  ( .A1(_u10_n18048 ), .A2(_u10_n18049 ), .A3(_u10_n18050 ), .A4(_u10_n18051 ), .ZN(_u10_n18043 ) );
NAND2_X1 _u10_U6634  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18045 ) );
NAND2_X1 _u10_U6633  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18046 ) );
NAND2_X1 _u10_U6632  ( .A1(1'b1), .A2(_u10_n12009 ), .ZN(_u10_n18047 ) );
NAND3_X1 _u10_U6631  ( .A1(_u10_n18045 ), .A2(_u10_n18046 ), .A3(_u10_n18047 ), .ZN(_u10_n18044 ) );
NOR4_X1 _u10_U6630  ( .A1(_u10_n18041 ), .A2(_u10_n18042 ), .A3(_u10_n18043 ), .A4(_u10_n18044 ), .ZN(_u10_n18019 ) );
NAND2_X1 _u10_U6629  ( .A1(1'b1), .A2(_u10_n11992 ), .ZN(_u10_n18037 ) );
NAND2_X1 _u10_U6628  ( .A1(1'b1), .A2(_u10_n11968 ), .ZN(_u10_n18038 ) );
NAND2_X1 _u10_U6627  ( .A1(1'b1), .A2(_u10_n11944 ), .ZN(_u10_n18039 ) );
NAND2_X1 _u10_U6626  ( .A1(1'b1), .A2(_u10_n11920 ), .ZN(_u10_n18040 ) );
NAND4_X1 _u10_U6625  ( .A1(_u10_n18037 ), .A2(_u10_n18038 ), .A3(_u10_n18039 ), .A4(_u10_n18040 ), .ZN(_u10_n18021 ) );
NAND2_X1 _u10_U6624  ( .A1(1'b1), .A2(_u10_n11896 ), .ZN(_u10_n18033 ) );
NAND2_X1 _u10_U6623  ( .A1(1'b1), .A2(_u10_n11872 ), .ZN(_u10_n18034 ) );
NAND2_X1 _u10_U6622  ( .A1(1'b1), .A2(_u10_n11848 ), .ZN(_u10_n18035 ) );
NAND2_X1 _u10_U6621  ( .A1(1'b1), .A2(_u10_n11824 ), .ZN(_u10_n18036 ) );
NAND4_X1 _u10_U6620  ( .A1(_u10_n18033 ), .A2(_u10_n18034 ), .A3(_u10_n18035 ), .A4(_u10_n18036 ), .ZN(_u10_n18022 ) );
NAND2_X1 _u10_U6619  ( .A1(1'b1), .A2(_u10_n11800 ), .ZN(_u10_n18029 ) );
NAND2_X1 _u10_U6618  ( .A1(1'b1), .A2(_u10_n11776 ), .ZN(_u10_n18030 ) );
NAND2_X1 _u10_U6617  ( .A1(1'b1), .A2(_u10_n11752 ), .ZN(_u10_n18031 ) );
NAND2_X1 _u10_U6616  ( .A1(1'b1), .A2(_u10_n11728 ), .ZN(_u10_n18032 ) );
NAND4_X1 _u10_U6615  ( .A1(_u10_n18029 ), .A2(_u10_n18030 ), .A3(_u10_n18031 ), .A4(_u10_n18032 ), .ZN(_u10_n18023 ) );
NAND2_X1 _u10_U6614  ( .A1(1'b1), .A2(_u10_n11704 ), .ZN(_u10_n18025 ) );
NAND2_X1 _u10_U6613  ( .A1(1'b1), .A2(_u10_n11680 ), .ZN(_u10_n18026 ) );
NAND2_X1 _u10_U6612  ( .A1(1'b1), .A2(_u10_n11656 ), .ZN(_u10_n18027 ) );
NAND2_X1 _u10_U6611  ( .A1(1'b1), .A2(_u10_n11632 ), .ZN(_u10_n18028 ) );
NAND4_X1 _u10_U6610  ( .A1(_u10_n18025 ), .A2(_u10_n18026 ), .A3(_u10_n18027 ), .A4(_u10_n18028 ), .ZN(_u10_n18024 ) );
NOR4_X1 _u10_U6609  ( .A1(_u10_n18021 ), .A2(_u10_n18022 ), .A3(_u10_n18023 ), .A4(_u10_n18024 ), .ZN(_u10_n18020 ) );
NAND2_X1 _u10_U6608  ( .A1(_u10_n18019 ), .A2(_u10_n18020 ), .ZN(am1[30]) );
NAND2_X1 _u10_U6607  ( .A1(1'b1), .A2(_u10_n12339 ), .ZN(_u10_n18015 ) );
NAND2_X1 _u10_U6606  ( .A1(1'b1), .A2(_u10_n12329 ), .ZN(_u10_n18016 ) );
NAND2_X1 _u10_U6605  ( .A1(1'b1), .A2(_u10_n12292 ), .ZN(_u10_n18017 ) );
NAND2_X1 _u10_U6604  ( .A1(1'b1), .A2(_u10_n12268 ), .ZN(_u10_n18018 ) );
NAND4_X1 _u10_U6603  ( .A1(_u10_n18015 ), .A2(_u10_n18016 ), .A3(_u10_n18017 ), .A4(_u10_n18018 ), .ZN(_u10_n18000 ) );
NAND2_X1 _u10_U6602  ( .A1(1'b1), .A2(_u10_n12243 ), .ZN(_u10_n18011 ) );
NAND2_X1 _u10_U6601  ( .A1(1'b1), .A2(_u10_n12219 ), .ZN(_u10_n18012 ) );
NAND2_X1 _u10_U6600  ( .A1(1'b1), .A2(_u10_n12196 ), .ZN(_u10_n18013 ) );
NAND2_X1 _u10_U6599  ( .A1(1'b1), .A2(_u10_n12171 ), .ZN(_u10_n18014 ) );
NAND4_X1 _u10_U6598  ( .A1(_u10_n18011 ), .A2(_u10_n18012 ), .A3(_u10_n18013 ), .A4(_u10_n18014 ), .ZN(_u10_n18001 ) );
NAND2_X1 _u10_U6597  ( .A1(1'b1), .A2(_u10_n12148 ), .ZN(_u10_n18007 ) );
NAND2_X1 _u10_U6596  ( .A1(1'b1), .A2(_u10_n12124 ), .ZN(_u10_n18008 ) );
NAND2_X1 _u10_U6595  ( .A1(1'b1), .A2(_u10_n12100 ), .ZN(_u10_n18009 ) );
NAND2_X1 _u10_U6594  ( .A1(1'b1), .A2(_u10_n12076 ), .ZN(_u10_n18010 ) );
NAND4_X1 _u10_U6593  ( .A1(_u10_n18007 ), .A2(_u10_n18008 ), .A3(_u10_n18009 ), .A4(_u10_n18010 ), .ZN(_u10_n18002 ) );
NAND2_X1 _u10_U6592  ( .A1(1'b1), .A2(_u10_n12052 ), .ZN(_u10_n18004 ) );
NAND2_X1 _u10_U6591  ( .A1(1'b1), .A2(_u10_n12028 ), .ZN(_u10_n18005 ) );
NAND2_X1 _u10_U6590  ( .A1(1'b1), .A2(_u10_n12009 ), .ZN(_u10_n18006 ) );
NAND3_X1 _u10_U6589  ( .A1(_u10_n18004 ), .A2(_u10_n18005 ), .A3(_u10_n18006 ), .ZN(_u10_n18003 ) );
NOR4_X1 _u10_U6588  ( .A1(_u10_n18000 ), .A2(_u10_n18001 ), .A3(_u10_n18002 ), .A4(_u10_n18003 ), .ZN(_u10_n17978 ) );
NAND2_X1 _u10_U6587  ( .A1(1'b1), .A2(_u10_n11992 ), .ZN(_u10_n17996 ) );
NAND2_X1 _u10_U6586  ( .A1(1'b1), .A2(_u10_n11968 ), .ZN(_u10_n17997 ) );
NAND2_X1 _u10_U6585  ( .A1(1'b1), .A2(_u10_n11944 ), .ZN(_u10_n17998 ) );
NAND2_X1 _u10_U6584  ( .A1(1'b1), .A2(_u10_n11920 ), .ZN(_u10_n17999 ) );
NAND4_X1 _u10_U6583  ( .A1(_u10_n17996 ), .A2(_u10_n17997 ), .A3(_u10_n17998 ), .A4(_u10_n17999 ), .ZN(_u10_n17980 ) );
NAND2_X1 _u10_U6582  ( .A1(1'b1), .A2(_u10_n11896 ), .ZN(_u10_n17992 ) );
NAND2_X1 _u10_U6581  ( .A1(1'b1), .A2(_u10_n11872 ), .ZN(_u10_n17993 ) );
NAND2_X1 _u10_U6580  ( .A1(1'b1), .A2(_u10_n11848 ), .ZN(_u10_n17994 ) );
NAND2_X1 _u10_U6579  ( .A1(1'b1), .A2(_u10_n11824 ), .ZN(_u10_n17995 ) );
NAND4_X1 _u10_U6578  ( .A1(_u10_n17992 ), .A2(_u10_n17993 ), .A3(_u10_n17994 ), .A4(_u10_n17995 ), .ZN(_u10_n17981 ) );
NAND2_X1 _u10_U6577  ( .A1(1'b1), .A2(_u10_n11800 ), .ZN(_u10_n17988 ) );
NAND2_X1 _u10_U6576  ( .A1(1'b1), .A2(_u10_n11776 ), .ZN(_u10_n17989 ) );
NAND2_X1 _u10_U6575  ( .A1(1'b1), .A2(_u10_n11752 ), .ZN(_u10_n17990 ) );
NAND2_X1 _u10_U6574  ( .A1(1'b1), .A2(_u10_n11728 ), .ZN(_u10_n17991 ) );
NAND4_X1 _u10_U6573  ( .A1(_u10_n17988 ), .A2(_u10_n17989 ), .A3(_u10_n17990 ), .A4(_u10_n17991 ), .ZN(_u10_n17982 ) );
NAND2_X1 _u10_U6572  ( .A1(1'b1), .A2(_u10_n11704 ), .ZN(_u10_n17984 ) );
NAND2_X1 _u10_U6571  ( .A1(1'b1), .A2(_u10_n11680 ), .ZN(_u10_n17985 ) );
NAND2_X1 _u10_U6570  ( .A1(1'b1), .A2(_u10_n11656 ), .ZN(_u10_n17986 ) );
NAND2_X1 _u10_U6569  ( .A1(1'b1), .A2(_u10_n11632 ), .ZN(_u10_n17987 ) );
NAND4_X1 _u10_U6568  ( .A1(_u10_n17984 ), .A2(_u10_n17985 ), .A3(_u10_n17986 ), .A4(_u10_n17987 ), .ZN(_u10_n17983 ) );
NOR4_X1 _u10_U6567  ( .A1(_u10_n17980 ), .A2(_u10_n17981 ), .A3(_u10_n17982 ), .A4(_u10_n17983 ), .ZN(_u10_n17979 ) );
NAND2_X1 _u10_U6566  ( .A1(_u10_n17978 ), .A2(_u10_n17979 ), .ZN(am1[31]) );
NAND2_X1 _u10_U6565  ( .A1(1'b0), .A2(_u10_n12340 ), .ZN(_u10_n17974 ) );
NAND2_X1 _u10_U6564  ( .A1(1'b0), .A2(_u10_n12316 ), .ZN(_u10_n17975 ) );
NAND2_X1 _u10_U6563  ( .A1(1'b0), .A2(_u10_n12293 ), .ZN(_u10_n17976 ) );
NAND2_X1 _u10_U6562  ( .A1(1'b0), .A2(_u10_n12269 ), .ZN(_u10_n17977 ) );
NAND4_X1 _u10_U6561  ( .A1(_u10_n17974 ), .A2(_u10_n17975 ), .A3(_u10_n17976 ), .A4(_u10_n17977 ), .ZN(_u10_n17959 ) );
NAND2_X1 _u10_U6560  ( .A1(1'b0), .A2(_u10_n12244 ), .ZN(_u10_n17970 ) );
NAND2_X1 _u10_U6559  ( .A1(1'b0), .A2(_u10_n12220 ), .ZN(_u10_n17971 ) );
NAND2_X1 _u10_U6558  ( .A1(1'b0), .A2(_u10_n12197 ), .ZN(_u10_n17972 ) );
NAND2_X1 _u10_U6557  ( .A1(1'b0), .A2(_u10_n12172 ), .ZN(_u10_n17973 ) );
NAND4_X1 _u10_U6556  ( .A1(_u10_n17970 ), .A2(_u10_n17971 ), .A3(_u10_n17972 ), .A4(_u10_n17973 ), .ZN(_u10_n17960 ) );
NAND2_X1 _u10_U6555  ( .A1(1'b0), .A2(_u10_n12149 ), .ZN(_u10_n17966 ) );
NAND2_X1 _u10_U6554  ( .A1(1'b0), .A2(_u10_n12125 ), .ZN(_u10_n17967 ) );
NAND2_X1 _u10_U6553  ( .A1(1'b0), .A2(_u10_n12101 ), .ZN(_u10_n17968 ) );
NAND2_X1 _u10_U6552  ( .A1(1'b0), .A2(_u10_n12077 ), .ZN(_u10_n17969 ) );
NAND4_X1 _u10_U6551  ( .A1(_u10_n17966 ), .A2(_u10_n17967 ), .A3(_u10_n17968 ), .A4(_u10_n17969 ), .ZN(_u10_n17961 ) );
NAND2_X1 _u10_U6550  ( .A1(1'b0), .A2(_u10_n12053 ), .ZN(_u10_n17963 ) );
NAND2_X1 _u10_U6549  ( .A1(1'b0), .A2(_u10_n12029 ), .ZN(_u10_n17964 ) );
NAND2_X1 _u10_U6548  ( .A1(1'b0), .A2(_u10_n12009 ), .ZN(_u10_n17965 ) );
NAND3_X1 _u10_U6547  ( .A1(_u10_n17963 ), .A2(_u10_n17964 ), .A3(_u10_n17965 ), .ZN(_u10_n17962 ) );
NOR4_X1 _u10_U6546  ( .A1(_u10_n17959 ), .A2(_u10_n17960 ), .A3(_u10_n17961 ), .A4(_u10_n17962 ), .ZN(_u10_n17937 ) );
NAND2_X1 _u10_U6545  ( .A1(1'b0), .A2(_u10_n11992 ), .ZN(_u10_n17955 ) );
NAND2_X1 _u10_U6544  ( .A1(1'b0), .A2(_u10_n11968 ), .ZN(_u10_n17956 ) );
NAND2_X1 _u10_U6543  ( .A1(1'b0), .A2(_u10_n11944 ), .ZN(_u10_n17957 ) );
NAND2_X1 _u10_U6542  ( .A1(1'b0), .A2(_u10_n11920 ), .ZN(_u10_n17958 ) );
NAND4_X1 _u10_U6541  ( .A1(_u10_n17955 ), .A2(_u10_n17956 ), .A3(_u10_n17957 ), .A4(_u10_n17958 ), .ZN(_u10_n17939 ) );
NAND2_X1 _u10_U6540  ( .A1(1'b0), .A2(_u10_n11896 ), .ZN(_u10_n17951 ) );
NAND2_X1 _u10_U6539  ( .A1(1'b0), .A2(_u10_n11872 ), .ZN(_u10_n17952 ) );
NAND2_X1 _u10_U6538  ( .A1(1'b0), .A2(_u10_n11848 ), .ZN(_u10_n17953 ) );
NAND2_X1 _u10_U6537  ( .A1(1'b0), .A2(_u10_n11824 ), .ZN(_u10_n17954 ) );
NAND4_X1 _u10_U6536  ( .A1(_u10_n17951 ), .A2(_u10_n17952 ), .A3(_u10_n17953 ), .A4(_u10_n17954 ), .ZN(_u10_n17940 ) );
NAND2_X1 _u10_U6535  ( .A1(1'b0), .A2(_u10_n11800 ), .ZN(_u10_n17947 ) );
NAND2_X1 _u10_U6534  ( .A1(1'b0), .A2(_u10_n11776 ), .ZN(_u10_n17948 ) );
NAND2_X1 _u10_U6533  ( .A1(1'b0), .A2(_u10_n11752 ), .ZN(_u10_n17949 ) );
NAND2_X1 _u10_U6532  ( .A1(1'b0), .A2(_u10_n11728 ), .ZN(_u10_n17950 ) );
NAND4_X1 _u10_U6531  ( .A1(_u10_n17947 ), .A2(_u10_n17948 ), .A3(_u10_n17949 ), .A4(_u10_n17950 ), .ZN(_u10_n17941 ) );
NAND2_X1 _u10_U6530  ( .A1(1'b0), .A2(_u10_n11704 ), .ZN(_u10_n17943 ) );
NAND2_X1 _u10_U6529  ( .A1(1'b0), .A2(_u10_n11680 ), .ZN(_u10_n17944 ) );
NAND2_X1 _u10_U6528  ( .A1(1'b0), .A2(_u10_n11656 ), .ZN(_u10_n17945 ) );
NAND2_X1 _u10_U6527  ( .A1(1'b0), .A2(_u10_n11632 ), .ZN(_u10_n17946 ) );
NAND4_X1 _u10_U6526  ( .A1(_u10_n17943 ), .A2(_u10_n17944 ), .A3(_u10_n17945 ), .A4(_u10_n17946 ), .ZN(_u10_n17942 ) );
NOR4_X1 _u10_U6525  ( .A1(_u10_n17939 ), .A2(_u10_n17940 ), .A3(_u10_n17941 ), .A4(_u10_n17942 ), .ZN(_u10_n17938 ) );
NAND2_X1 _u10_U6524  ( .A1(_u10_n17937 ), .A2(_u10_n17938 ), .ZN(am1[3]) );
NAND2_X1 _u10_U6523  ( .A1(1'b1), .A2(_u10_n12340 ), .ZN(_u10_n17933 ) );
NAND2_X1 _u10_U6522  ( .A1(1'b1), .A2(_u10_n12316 ), .ZN(_u10_n17934 ) );
NAND2_X1 _u10_U6521  ( .A1(1'b1), .A2(_u10_n12293 ), .ZN(_u10_n17935 ) );
NAND2_X1 _u10_U6520  ( .A1(1'b1), .A2(_u10_n12269 ), .ZN(_u10_n17936 ) );
NAND4_X1 _u10_U6519  ( .A1(_u10_n17933 ), .A2(_u10_n17934 ), .A3(_u10_n17935 ), .A4(_u10_n17936 ), .ZN(_u10_n17918 ) );
NAND2_X1 _u10_U6518  ( .A1(1'b1), .A2(_u10_n12244 ), .ZN(_u10_n17929 ) );
NAND2_X1 _u10_U6517  ( .A1(1'b1), .A2(_u10_n12220 ), .ZN(_u10_n17930 ) );
NAND2_X1 _u10_U6516  ( .A1(1'b1), .A2(_u10_n12197 ), .ZN(_u10_n17931 ) );
NAND2_X1 _u10_U6515  ( .A1(1'b1), .A2(_u10_n12172 ), .ZN(_u10_n17932 ) );
NAND4_X1 _u10_U6514  ( .A1(_u10_n17929 ), .A2(_u10_n17930 ), .A3(_u10_n17931 ), .A4(_u10_n17932 ), .ZN(_u10_n17919 ) );
NAND2_X1 _u10_U6513  ( .A1(1'b1), .A2(_u10_n12149 ), .ZN(_u10_n17925 ) );
NAND2_X1 _u10_U6512  ( .A1(1'b1), .A2(_u10_n12125 ), .ZN(_u10_n17926 ) );
NAND2_X1 _u10_U6511  ( .A1(1'b1), .A2(_u10_n12101 ), .ZN(_u10_n17927 ) );
NAND2_X1 _u10_U6510  ( .A1(1'b1), .A2(_u10_n12077 ), .ZN(_u10_n17928 ) );
NAND4_X1 _u10_U6509  ( .A1(_u10_n17925 ), .A2(_u10_n17926 ), .A3(_u10_n17927 ), .A4(_u10_n17928 ), .ZN(_u10_n17920 ) );
NAND2_X1 _u10_U6508  ( .A1(1'b1), .A2(_u10_n12053 ), .ZN(_u10_n17922 ) );
NAND2_X1 _u10_U6507  ( .A1(1'b1), .A2(_u10_n12029 ), .ZN(_u10_n17923 ) );
NAND2_X1 _u10_U6506  ( .A1(1'b1), .A2(_u10_n12009 ), .ZN(_u10_n17924 ) );
NAND3_X1 _u10_U6505  ( .A1(_u10_n17922 ), .A2(_u10_n17923 ), .A3(_u10_n17924 ), .ZN(_u10_n17921 ) );
NOR4_X1 _u10_U6504  ( .A1(_u10_n17918 ), .A2(_u10_n17919 ), .A3(_u10_n17920 ), .A4(_u10_n17921 ), .ZN(_u10_n17896 ) );
NAND2_X1 _u10_U6503  ( .A1(1'b1), .A2(_u10_n11992 ), .ZN(_u10_n17914 ) );
NAND2_X1 _u10_U6502  ( .A1(1'b1), .A2(_u10_n11968 ), .ZN(_u10_n17915 ) );
NAND2_X1 _u10_U6501  ( .A1(1'b1), .A2(_u10_n11944 ), .ZN(_u10_n17916 ) );
NAND2_X1 _u10_U6500  ( .A1(1'b1), .A2(_u10_n11920 ), .ZN(_u10_n17917 ) );
NAND4_X1 _u10_U6499  ( .A1(_u10_n17914 ), .A2(_u10_n17915 ), .A3(_u10_n17916 ), .A4(_u10_n17917 ), .ZN(_u10_n17898 ) );
NAND2_X1 _u10_U6498  ( .A1(1'b1), .A2(_u10_n11896 ), .ZN(_u10_n17910 ) );
NAND2_X1 _u10_U6497  ( .A1(1'b1), .A2(_u10_n11872 ), .ZN(_u10_n17911 ) );
NAND2_X1 _u10_U6496  ( .A1(1'b1), .A2(_u10_n11848 ), .ZN(_u10_n17912 ) );
NAND2_X1 _u10_U6495  ( .A1(1'b1), .A2(_u10_n11824 ), .ZN(_u10_n17913 ) );
NAND4_X1 _u10_U6494  ( .A1(_u10_n17910 ), .A2(_u10_n17911 ), .A3(_u10_n17912 ), .A4(_u10_n17913 ), .ZN(_u10_n17899 ) );
NAND2_X1 _u10_U6493  ( .A1(1'b1), .A2(_u10_n11800 ), .ZN(_u10_n17906 ) );
NAND2_X1 _u10_U6492  ( .A1(1'b1), .A2(_u10_n11776 ), .ZN(_u10_n17907 ) );
NAND2_X1 _u10_U6491  ( .A1(1'b1), .A2(_u10_n11752 ), .ZN(_u10_n17908 ) );
NAND2_X1 _u10_U6490  ( .A1(1'b1), .A2(_u10_n11728 ), .ZN(_u10_n17909 ) );
NAND4_X1 _u10_U6489  ( .A1(_u10_n17906 ), .A2(_u10_n17907 ), .A3(_u10_n17908 ), .A4(_u10_n17909 ), .ZN(_u10_n17900 ) );
NAND2_X1 _u10_U6488  ( .A1(1'b1), .A2(_u10_n11704 ), .ZN(_u10_n17902 ) );
NAND2_X1 _u10_U6487  ( .A1(1'b1), .A2(_u10_n11680 ), .ZN(_u10_n17903 ) );
NAND2_X1 _u10_U6486  ( .A1(1'b1), .A2(_u10_n11656 ), .ZN(_u10_n17904 ) );
NAND2_X1 _u10_U6485  ( .A1(1'b1), .A2(_u10_n11632 ), .ZN(_u10_n17905 ) );
NAND4_X1 _u10_U6484  ( .A1(_u10_n17902 ), .A2(_u10_n17903 ), .A3(_u10_n17904 ), .A4(_u10_n17905 ), .ZN(_u10_n17901 ) );
NOR4_X1 _u10_U6483  ( .A1(_u10_n17898 ), .A2(_u10_n17899 ), .A3(_u10_n17900 ), .A4(_u10_n17901 ), .ZN(_u10_n17897 ) );
NAND2_X1 _u10_U6482  ( .A1(_u10_n17896 ), .A2(_u10_n17897 ), .ZN(am1[4]) );
NAND2_X1 _u10_U6481  ( .A1(1'b1), .A2(_u10_n12340 ), .ZN(_u10_n17892 ) );
NAND2_X1 _u10_U6480  ( .A1(1'b1), .A2(_u10_n12316 ), .ZN(_u10_n17893 ) );
NAND2_X1 _u10_U6479  ( .A1(1'b1), .A2(_u10_n12293 ), .ZN(_u10_n17894 ) );
NAND2_X1 _u10_U6478  ( .A1(1'b1), .A2(_u10_n12269 ), .ZN(_u10_n17895 ) );
NAND4_X1 _u10_U6477  ( .A1(_u10_n17892 ), .A2(_u10_n17893 ), .A3(_u10_n17894 ), .A4(_u10_n17895 ), .ZN(_u10_n17877 ) );
NAND2_X1 _u10_U6476  ( .A1(1'b1), .A2(_u10_n12244 ), .ZN(_u10_n17888 ) );
NAND2_X1 _u10_U6475  ( .A1(1'b1), .A2(_u10_n12220 ), .ZN(_u10_n17889 ) );
NAND2_X1 _u10_U6474  ( .A1(1'b1), .A2(_u10_n12197 ), .ZN(_u10_n17890 ) );
NAND2_X1 _u10_U6473  ( .A1(1'b1), .A2(_u10_n12172 ), .ZN(_u10_n17891 ) );
NAND4_X1 _u10_U6472  ( .A1(_u10_n17888 ), .A2(_u10_n17889 ), .A3(_u10_n17890 ), .A4(_u10_n17891 ), .ZN(_u10_n17878 ) );
NAND2_X1 _u10_U6471  ( .A1(1'b1), .A2(_u10_n12149 ), .ZN(_u10_n17884 ) );
NAND2_X1 _u10_U6470  ( .A1(1'b1), .A2(_u10_n12125 ), .ZN(_u10_n17885 ) );
NAND2_X1 _u10_U6469  ( .A1(1'b1), .A2(_u10_n12101 ), .ZN(_u10_n17886 ) );
NAND2_X1 _u10_U6468  ( .A1(1'b1), .A2(_u10_n12077 ), .ZN(_u10_n17887 ) );
NAND4_X1 _u10_U6467  ( .A1(_u10_n17884 ), .A2(_u10_n17885 ), .A3(_u10_n17886 ), .A4(_u10_n17887 ), .ZN(_u10_n17879 ) );
NAND2_X1 _u10_U6466  ( .A1(1'b1), .A2(_u10_n12053 ), .ZN(_u10_n17881 ) );
NAND2_X1 _u10_U6465  ( .A1(1'b1), .A2(_u10_n12029 ), .ZN(_u10_n17882 ) );
NAND2_X1 _u10_U6464  ( .A1(1'b1), .A2(_u10_n12009 ), .ZN(_u10_n17883 ) );
NAND3_X1 _u10_U6463  ( .A1(_u10_n17881 ), .A2(_u10_n17882 ), .A3(_u10_n17883 ), .ZN(_u10_n17880 ) );
NOR4_X1 _u10_U6462  ( .A1(_u10_n17877 ), .A2(_u10_n17878 ), .A3(_u10_n17879 ), .A4(_u10_n17880 ), .ZN(_u10_n17855 ) );
NAND2_X1 _u10_U6461  ( .A1(1'b1), .A2(_u10_n11992 ), .ZN(_u10_n17873 ) );
NAND2_X1 _u10_U6460  ( .A1(1'b1), .A2(_u10_n11968 ), .ZN(_u10_n17874 ) );
NAND2_X1 _u10_U6459  ( .A1(1'b1), .A2(_u10_n11944 ), .ZN(_u10_n17875 ) );
NAND2_X1 _u10_U6458  ( .A1(1'b1), .A2(_u10_n11920 ), .ZN(_u10_n17876 ) );
NAND4_X1 _u10_U6457  ( .A1(_u10_n17873 ), .A2(_u10_n17874 ), .A3(_u10_n17875 ), .A4(_u10_n17876 ), .ZN(_u10_n17857 ) );
NAND2_X1 _u10_U6456  ( .A1(1'b1), .A2(_u10_n11896 ), .ZN(_u10_n17869 ) );
NAND2_X1 _u10_U6455  ( .A1(1'b1), .A2(_u10_n11872 ), .ZN(_u10_n17870 ) );
NAND2_X1 _u10_U6454  ( .A1(1'b1), .A2(_u10_n11848 ), .ZN(_u10_n17871 ) );
NAND2_X1 _u10_U6453  ( .A1(1'b1), .A2(_u10_n11824 ), .ZN(_u10_n17872 ) );
NAND4_X1 _u10_U6452  ( .A1(_u10_n17869 ), .A2(_u10_n17870 ), .A3(_u10_n17871 ), .A4(_u10_n17872 ), .ZN(_u10_n17858 ) );
NAND2_X1 _u10_U6451  ( .A1(1'b1), .A2(_u10_n11800 ), .ZN(_u10_n17865 ) );
NAND2_X1 _u10_U6450  ( .A1(1'b1), .A2(_u10_n11776 ), .ZN(_u10_n17866 ) );
NAND2_X1 _u10_U6449  ( .A1(1'b1), .A2(_u10_n11752 ), .ZN(_u10_n17867 ) );
NAND2_X1 _u10_U6448  ( .A1(1'b1), .A2(_u10_n11728 ), .ZN(_u10_n17868 ) );
NAND4_X1 _u10_U6447  ( .A1(_u10_n17865 ), .A2(_u10_n17866 ), .A3(_u10_n17867 ), .A4(_u10_n17868 ), .ZN(_u10_n17859 ) );
NAND2_X1 _u10_U6446  ( .A1(1'b1), .A2(_u10_n11704 ), .ZN(_u10_n17861 ) );
NAND2_X1 _u10_U6445  ( .A1(1'b1), .A2(_u10_n11680 ), .ZN(_u10_n17862 ) );
NAND2_X1 _u10_U6444  ( .A1(1'b1), .A2(_u10_n11656 ), .ZN(_u10_n17863 ) );
NAND2_X1 _u10_U6443  ( .A1(1'b1), .A2(_u10_n11632 ), .ZN(_u10_n17864 ) );
NAND4_X1 _u10_U6442  ( .A1(_u10_n17861 ), .A2(_u10_n17862 ), .A3(_u10_n17863 ), .A4(_u10_n17864 ), .ZN(_u10_n17860 ) );
NOR4_X1 _u10_U6441  ( .A1(_u10_n17857 ), .A2(_u10_n17858 ), .A3(_u10_n17859 ), .A4(_u10_n17860 ), .ZN(_u10_n17856 ) );
NAND2_X1 _u10_U6440  ( .A1(_u10_n17855 ), .A2(_u10_n17856 ), .ZN(am1[5]) );
NAND2_X1 _u10_U6439  ( .A1(1'b1), .A2(_u10_n12340 ), .ZN(_u10_n17851 ) );
NAND2_X1 _u10_U6438  ( .A1(1'b1), .A2(_u10_n12316 ), .ZN(_u10_n17852 ) );
NAND2_X1 _u10_U6437  ( .A1(1'b1), .A2(_u10_n12293 ), .ZN(_u10_n17853 ) );
NAND2_X1 _u10_U6436  ( .A1(1'b1), .A2(_u10_n12269 ), .ZN(_u10_n17854 ) );
NAND4_X1 _u10_U6435  ( .A1(_u10_n17851 ), .A2(_u10_n17852 ), .A3(_u10_n17853 ), .A4(_u10_n17854 ), .ZN(_u10_n17836 ) );
NAND2_X1 _u10_U6434  ( .A1(1'b1), .A2(_u10_n12244 ), .ZN(_u10_n17847 ) );
NAND2_X1 _u10_U6433  ( .A1(1'b1), .A2(_u10_n12220 ), .ZN(_u10_n17848 ) );
NAND2_X1 _u10_U6432  ( .A1(1'b1), .A2(_u10_n12197 ), .ZN(_u10_n17849 ) );
NAND2_X1 _u10_U6431  ( .A1(1'b1), .A2(_u10_n12172 ), .ZN(_u10_n17850 ) );
NAND4_X1 _u10_U6430  ( .A1(_u10_n17847 ), .A2(_u10_n17848 ), .A3(_u10_n17849 ), .A4(_u10_n17850 ), .ZN(_u10_n17837 ) );
NAND2_X1 _u10_U6429  ( .A1(1'b1), .A2(_u10_n12149 ), .ZN(_u10_n17843 ) );
NAND2_X1 _u10_U6428  ( .A1(1'b1), .A2(_u10_n12125 ), .ZN(_u10_n17844 ) );
NAND2_X1 _u10_U6427  ( .A1(1'b1), .A2(_u10_n12101 ), .ZN(_u10_n17845 ) );
NAND2_X1 _u10_U6426  ( .A1(1'b1), .A2(_u10_n12077 ), .ZN(_u10_n17846 ) );
NAND4_X1 _u10_U6425  ( .A1(_u10_n17843 ), .A2(_u10_n17844 ), .A3(_u10_n17845 ), .A4(_u10_n17846 ), .ZN(_u10_n17838 ) );
NAND2_X1 _u10_U6424  ( .A1(1'b1), .A2(_u10_n12053 ), .ZN(_u10_n17840 ) );
NAND2_X1 _u10_U6423  ( .A1(1'b1), .A2(_u10_n12029 ), .ZN(_u10_n17841 ) );
NAND2_X1 _u10_U6422  ( .A1(1'b1), .A2(_u10_n12009 ), .ZN(_u10_n17842 ) );
NAND3_X1 _u10_U6421  ( .A1(_u10_n17840 ), .A2(_u10_n17841 ), .A3(_u10_n17842 ), .ZN(_u10_n17839 ) );
NOR4_X1 _u10_U6420  ( .A1(_u10_n17836 ), .A2(_u10_n17837 ), .A3(_u10_n17838 ), .A4(_u10_n17839 ), .ZN(_u10_n17814 ) );
NAND2_X1 _u10_U6419  ( .A1(1'b1), .A2(_u10_n11992 ), .ZN(_u10_n17832 ) );
NAND2_X1 _u10_U6418  ( .A1(1'b1), .A2(_u10_n11968 ), .ZN(_u10_n17833 ) );
NAND2_X1 _u10_U6417  ( .A1(1'b1), .A2(_u10_n11944 ), .ZN(_u10_n17834 ) );
NAND2_X1 _u10_U6416  ( .A1(1'b1), .A2(_u10_n11920 ), .ZN(_u10_n17835 ) );
NAND4_X1 _u10_U6415  ( .A1(_u10_n17832 ), .A2(_u10_n17833 ), .A3(_u10_n17834 ), .A4(_u10_n17835 ), .ZN(_u10_n17816 ) );
NAND2_X1 _u10_U6414  ( .A1(1'b1), .A2(_u10_n11896 ), .ZN(_u10_n17828 ) );
NAND2_X1 _u10_U6413  ( .A1(1'b1), .A2(_u10_n11872 ), .ZN(_u10_n17829 ) );
NAND2_X1 _u10_U6412  ( .A1(1'b1), .A2(_u10_n11848 ), .ZN(_u10_n17830 ) );
NAND2_X1 _u10_U6411  ( .A1(1'b1), .A2(_u10_n11824 ), .ZN(_u10_n17831 ) );
NAND4_X1 _u10_U6410  ( .A1(_u10_n17828 ), .A2(_u10_n17829 ), .A3(_u10_n17830 ), .A4(_u10_n17831 ), .ZN(_u10_n17817 ) );
NAND2_X1 _u10_U6409  ( .A1(1'b1), .A2(_u10_n11800 ), .ZN(_u10_n17824 ) );
NAND2_X1 _u10_U6408  ( .A1(1'b1), .A2(_u10_n11776 ), .ZN(_u10_n17825 ) );
NAND2_X1 _u10_U6407  ( .A1(1'b1), .A2(_u10_n11752 ), .ZN(_u10_n17826 ) );
NAND2_X1 _u10_U6406  ( .A1(1'b1), .A2(_u10_n11728 ), .ZN(_u10_n17827 ) );
NAND4_X1 _u10_U6405  ( .A1(_u10_n17824 ), .A2(_u10_n17825 ), .A3(_u10_n17826 ), .A4(_u10_n17827 ), .ZN(_u10_n17818 ) );
NAND2_X1 _u10_U6404  ( .A1(1'b1), .A2(_u10_n11704 ), .ZN(_u10_n17820 ) );
NAND2_X1 _u10_U6403  ( .A1(1'b1), .A2(_u10_n11680 ), .ZN(_u10_n17821 ) );
NAND2_X1 _u10_U6402  ( .A1(1'b1), .A2(_u10_n11656 ), .ZN(_u10_n17822 ) );
NAND2_X1 _u10_U6401  ( .A1(1'b1), .A2(_u10_n11632 ), .ZN(_u10_n17823 ) );
NAND4_X1 _u10_U6400  ( .A1(_u10_n17820 ), .A2(_u10_n17821 ), .A3(_u10_n17822 ), .A4(_u10_n17823 ), .ZN(_u10_n17819 ) );
NOR4_X1 _u10_U6399  ( .A1(_u10_n17816 ), .A2(_u10_n17817 ), .A3(_u10_n17818 ), .A4(_u10_n17819 ), .ZN(_u10_n17815 ) );
NAND2_X1 _u10_U6398  ( .A1(_u10_n17814 ), .A2(_u10_n17815 ), .ZN(am1[6]) );
NAND2_X1 _u10_U6397  ( .A1(1'b1), .A2(_u10_n12340 ), .ZN(_u10_n17810 ) );
NAND2_X1 _u10_U6396  ( .A1(1'b1), .A2(_u10_n12316 ), .ZN(_u10_n17811 ) );
NAND2_X1 _u10_U6395  ( .A1(1'b1), .A2(_u10_n12293 ), .ZN(_u10_n17812 ) );
NAND2_X1 _u10_U6394  ( .A1(1'b1), .A2(_u10_n12269 ), .ZN(_u10_n17813 ) );
NAND4_X1 _u10_U6393  ( .A1(_u10_n17810 ), .A2(_u10_n17811 ), .A3(_u10_n17812 ), .A4(_u10_n17813 ), .ZN(_u10_n17795 ) );
NAND2_X1 _u10_U6392  ( .A1(1'b1), .A2(_u10_n12244 ), .ZN(_u10_n17806 ) );
NAND2_X1 _u10_U6391  ( .A1(1'b1), .A2(_u10_n12220 ), .ZN(_u10_n17807 ) );
NAND2_X1 _u10_U6390  ( .A1(1'b1), .A2(_u10_n12197 ), .ZN(_u10_n17808 ) );
NAND2_X1 _u10_U6389  ( .A1(1'b1), .A2(_u10_n12172 ), .ZN(_u10_n17809 ) );
NAND4_X1 _u10_U6388  ( .A1(_u10_n17806 ), .A2(_u10_n17807 ), .A3(_u10_n17808 ), .A4(_u10_n17809 ), .ZN(_u10_n17796 ) );
NAND2_X1 _u10_U6387  ( .A1(1'b1), .A2(_u10_n12149 ), .ZN(_u10_n17802 ) );
NAND2_X1 _u10_U6386  ( .A1(1'b1), .A2(_u10_n12125 ), .ZN(_u10_n17803 ) );
NAND2_X1 _u10_U6385  ( .A1(1'b1), .A2(_u10_n12101 ), .ZN(_u10_n17804 ) );
NAND2_X1 _u10_U6384  ( .A1(1'b1), .A2(_u10_n12077 ), .ZN(_u10_n17805 ) );
NAND4_X1 _u10_U6383  ( .A1(_u10_n17802 ), .A2(_u10_n17803 ), .A3(_u10_n17804 ), .A4(_u10_n17805 ), .ZN(_u10_n17797 ) );
NAND2_X1 _u10_U6382  ( .A1(1'b1), .A2(_u10_n12053 ), .ZN(_u10_n17799 ) );
NAND2_X1 _u10_U6381  ( .A1(1'b1), .A2(_u10_n12029 ), .ZN(_u10_n17800 ) );
NAND2_X1 _u10_U6380  ( .A1(1'b1), .A2(_u10_n12009 ), .ZN(_u10_n17801 ) );
NAND3_X1 _u10_U6379  ( .A1(_u10_n17799 ), .A2(_u10_n17800 ), .A3(_u10_n17801 ), .ZN(_u10_n17798 ) );
NOR4_X1 _u10_U6378  ( .A1(_u10_n17795 ), .A2(_u10_n17796 ), .A3(_u10_n17797 ), .A4(_u10_n17798 ), .ZN(_u10_n17773 ) );
NAND2_X1 _u10_U6377  ( .A1(1'b1), .A2(_u10_n11993 ), .ZN(_u10_n17791 ) );
NAND2_X1 _u10_U6376  ( .A1(1'b1), .A2(_u10_n11969 ), .ZN(_u10_n17792 ) );
NAND2_X1 _u10_U6375  ( .A1(1'b1), .A2(_u10_n11945 ), .ZN(_u10_n17793 ) );
NAND2_X1 _u10_U6374  ( .A1(1'b1), .A2(_u10_n11921 ), .ZN(_u10_n17794 ) );
NAND4_X1 _u10_U6373  ( .A1(_u10_n17791 ), .A2(_u10_n17792 ), .A3(_u10_n17793 ), .A4(_u10_n17794 ), .ZN(_u10_n17775 ) );
NAND2_X1 _u10_U6372  ( .A1(1'b1), .A2(_u10_n11897 ), .ZN(_u10_n17787 ) );
NAND2_X1 _u10_U6371  ( .A1(1'b1), .A2(_u10_n11873 ), .ZN(_u10_n17788 ) );
NAND2_X1 _u10_U6370  ( .A1(1'b1), .A2(_u10_n11849 ), .ZN(_u10_n17789 ) );
NAND2_X1 _u10_U6369  ( .A1(1'b1), .A2(_u10_n11825 ), .ZN(_u10_n17790 ) );
NAND4_X1 _u10_U6368  ( .A1(_u10_n17787 ), .A2(_u10_n17788 ), .A3(_u10_n17789 ), .A4(_u10_n17790 ), .ZN(_u10_n17776 ) );
NAND2_X1 _u10_U6367  ( .A1(1'b1), .A2(_u10_n11801 ), .ZN(_u10_n17783 ) );
NAND2_X1 _u10_U6366  ( .A1(1'b1), .A2(_u10_n11777 ), .ZN(_u10_n17784 ) );
NAND2_X1 _u10_U6365  ( .A1(1'b1), .A2(_u10_n11753 ), .ZN(_u10_n17785 ) );
NAND2_X1 _u10_U6364  ( .A1(1'b1), .A2(_u10_n11729 ), .ZN(_u10_n17786 ) );
NAND4_X1 _u10_U6363  ( .A1(_u10_n17783 ), .A2(_u10_n17784 ), .A3(_u10_n17785 ), .A4(_u10_n17786 ), .ZN(_u10_n17777 ) );
NAND2_X1 _u10_U6362  ( .A1(1'b1), .A2(_u10_n11705 ), .ZN(_u10_n17779 ) );
NAND2_X1 _u10_U6361  ( .A1(1'b1), .A2(_u10_n11681 ), .ZN(_u10_n17780 ) );
NAND2_X1 _u10_U6360  ( .A1(1'b1), .A2(_u10_n11657 ), .ZN(_u10_n17781 ) );
NAND2_X1 _u10_U6359  ( .A1(1'b1), .A2(_u10_n11633 ), .ZN(_u10_n17782 ) );
NAND4_X1 _u10_U6358  ( .A1(_u10_n17779 ), .A2(_u10_n17780 ), .A3(_u10_n17781 ), .A4(_u10_n17782 ), .ZN(_u10_n17778 ) );
NOR4_X1 _u10_U6357  ( .A1(_u10_n17775 ), .A2(_u10_n17776 ), .A3(_u10_n17777 ), .A4(_u10_n17778 ), .ZN(_u10_n17774 ) );
NAND2_X1 _u10_U6356  ( .A1(_u10_n17773 ), .A2(_u10_n17774 ), .ZN(am1[7]) );
NAND2_X1 _u10_U6355  ( .A1(1'b1), .A2(_u10_n12340 ), .ZN(_u10_n17769 ) );
NAND2_X1 _u10_U6354  ( .A1(1'b1), .A2(_u10_n12316 ), .ZN(_u10_n17770 ) );
NAND2_X1 _u10_U6353  ( .A1(1'b1), .A2(_u10_n12293 ), .ZN(_u10_n17771 ) );
NAND2_X1 _u10_U6352  ( .A1(1'b1), .A2(_u10_n12269 ), .ZN(_u10_n17772 ) );
NAND4_X1 _u10_U6351  ( .A1(_u10_n17769 ), .A2(_u10_n17770 ), .A3(_u10_n17771 ), .A4(_u10_n17772 ), .ZN(_u10_n17754 ) );
NAND2_X1 _u10_U6350  ( .A1(1'b1), .A2(_u10_n12244 ), .ZN(_u10_n17765 ) );
NAND2_X1 _u10_U6349  ( .A1(1'b1), .A2(_u10_n12220 ), .ZN(_u10_n17766 ) );
NAND2_X1 _u10_U6348  ( .A1(1'b1), .A2(_u10_n12197 ), .ZN(_u10_n17767 ) );
NAND2_X1 _u10_U6347  ( .A1(1'b1), .A2(_u10_n12172 ), .ZN(_u10_n17768 ) );
NAND4_X1 _u10_U6346  ( .A1(_u10_n17765 ), .A2(_u10_n17766 ), .A3(_u10_n17767 ), .A4(_u10_n17768 ), .ZN(_u10_n17755 ) );
NAND2_X1 _u10_U6345  ( .A1(1'b1), .A2(_u10_n12149 ), .ZN(_u10_n17761 ) );
NAND2_X1 _u10_U6344  ( .A1(1'b1), .A2(_u10_n12125 ), .ZN(_u10_n17762 ) );
NAND2_X1 _u10_U6343  ( .A1(1'b1), .A2(_u10_n12101 ), .ZN(_u10_n17763 ) );
NAND2_X1 _u10_U6342  ( .A1(1'b1), .A2(_u10_n12077 ), .ZN(_u10_n17764 ) );
NAND4_X1 _u10_U6341  ( .A1(_u10_n17761 ), .A2(_u10_n17762 ), .A3(_u10_n17763 ), .A4(_u10_n17764 ), .ZN(_u10_n17756 ) );
NAND2_X1 _u10_U6340  ( .A1(1'b1), .A2(_u10_n12053 ), .ZN(_u10_n17758 ) );
NAND2_X1 _u10_U6339  ( .A1(1'b1), .A2(_u10_n12029 ), .ZN(_u10_n17759 ) );
NAND2_X1 _u10_U6338  ( .A1(1'b1), .A2(_u10_n12009 ), .ZN(_u10_n17760 ) );
NAND3_X1 _u10_U6337  ( .A1(_u10_n17758 ), .A2(_u10_n17759 ), .A3(_u10_n17760 ), .ZN(_u10_n17757 ) );
NOR4_X1 _u10_U6336  ( .A1(_u10_n17754 ), .A2(_u10_n17755 ), .A3(_u10_n17756 ), .A4(_u10_n17757 ), .ZN(_u10_n17732 ) );
NAND2_X1 _u10_U6335  ( .A1(1'b1), .A2(_u10_n11993 ), .ZN(_u10_n17750 ) );
NAND2_X1 _u10_U6334  ( .A1(1'b1), .A2(_u10_n11969 ), .ZN(_u10_n17751 ) );
NAND2_X1 _u10_U6333  ( .A1(1'b1), .A2(_u10_n11945 ), .ZN(_u10_n17752 ) );
NAND2_X1 _u10_U6332  ( .A1(1'b1), .A2(_u10_n11921 ), .ZN(_u10_n17753 ) );
NAND4_X1 _u10_U6331  ( .A1(_u10_n17750 ), .A2(_u10_n17751 ), .A3(_u10_n17752 ), .A4(_u10_n17753 ), .ZN(_u10_n17734 ) );
NAND2_X1 _u10_U6330  ( .A1(1'b1), .A2(_u10_n11897 ), .ZN(_u10_n17746 ) );
NAND2_X1 _u10_U6329  ( .A1(1'b1), .A2(_u10_n11873 ), .ZN(_u10_n17747 ) );
NAND2_X1 _u10_U6328  ( .A1(1'b1), .A2(_u10_n11849 ), .ZN(_u10_n17748 ) );
NAND2_X1 _u10_U6327  ( .A1(1'b1), .A2(_u10_n11825 ), .ZN(_u10_n17749 ) );
NAND4_X1 _u10_U6326  ( .A1(_u10_n17746 ), .A2(_u10_n17747 ), .A3(_u10_n17748 ), .A4(_u10_n17749 ), .ZN(_u10_n17735 ) );
NAND2_X1 _u10_U6325  ( .A1(1'b1), .A2(_u10_n11801 ), .ZN(_u10_n17742 ) );
NAND2_X1 _u10_U6324  ( .A1(1'b1), .A2(_u10_n11777 ), .ZN(_u10_n17743 ) );
NAND2_X1 _u10_U6323  ( .A1(1'b1), .A2(_u10_n11753 ), .ZN(_u10_n17744 ) );
NAND2_X1 _u10_U6322  ( .A1(1'b1), .A2(_u10_n11729 ), .ZN(_u10_n17745 ) );
NAND4_X1 _u10_U6321  ( .A1(_u10_n17742 ), .A2(_u10_n17743 ), .A3(_u10_n17744 ), .A4(_u10_n17745 ), .ZN(_u10_n17736 ) );
NAND2_X1 _u10_U6320  ( .A1(1'b1), .A2(_u10_n11705 ), .ZN(_u10_n17738 ) );
NAND2_X1 _u10_U6319  ( .A1(1'b1), .A2(_u10_n11681 ), .ZN(_u10_n17739 ) );
NAND2_X1 _u10_U6318  ( .A1(1'b1), .A2(_u10_n11657 ), .ZN(_u10_n17740 ) );
NAND2_X1 _u10_U6317  ( .A1(1'b1), .A2(_u10_n11633 ), .ZN(_u10_n17741 ) );
NAND4_X1 _u10_U6316  ( .A1(_u10_n17738 ), .A2(_u10_n17739 ), .A3(_u10_n17740 ), .A4(_u10_n17741 ), .ZN(_u10_n17737 ) );
NOR4_X1 _u10_U6315  ( .A1(_u10_n17734 ), .A2(_u10_n17735 ), .A3(_u10_n17736 ), .A4(_u10_n17737 ), .ZN(_u10_n17733 ) );
NAND2_X1 _u10_U6314  ( .A1(_u10_n17732 ), .A2(_u10_n17733 ), .ZN(am1[8]) );
NAND2_X1 _u10_U6313  ( .A1(1'b1), .A2(_u10_n12340 ), .ZN(_u10_n17728 ) );
NAND2_X1 _u10_U6312  ( .A1(1'b1), .A2(_u10_n12316 ), .ZN(_u10_n17729 ) );
NAND2_X1 _u10_U6311  ( .A1(1'b1), .A2(_u10_n12293 ), .ZN(_u10_n17730 ) );
NAND2_X1 _u10_U6310  ( .A1(1'b1), .A2(_u10_n12269 ), .ZN(_u10_n17731 ) );
NAND4_X1 _u10_U6309  ( .A1(_u10_n17728 ), .A2(_u10_n17729 ), .A3(_u10_n17730 ), .A4(_u10_n17731 ), .ZN(_u10_n17713 ) );
NAND2_X1 _u10_U6308  ( .A1(1'b1), .A2(_u10_n12244 ), .ZN(_u10_n17724 ) );
NAND2_X1 _u10_U6307  ( .A1(1'b1), .A2(_u10_n12220 ), .ZN(_u10_n17725 ) );
NAND2_X1 _u10_U6306  ( .A1(1'b1), .A2(_u10_n12197 ), .ZN(_u10_n17726 ) );
NAND2_X1 _u10_U6305  ( .A1(1'b1), .A2(_u10_n12172 ), .ZN(_u10_n17727 ) );
NAND4_X1 _u10_U6304  ( .A1(_u10_n17724 ), .A2(_u10_n17725 ), .A3(_u10_n17726 ), .A4(_u10_n17727 ), .ZN(_u10_n17714 ) );
NAND2_X1 _u10_U6303  ( .A1(1'b1), .A2(_u10_n12149 ), .ZN(_u10_n17720 ) );
NAND2_X1 _u10_U6302  ( .A1(1'b1), .A2(_u10_n12125 ), .ZN(_u10_n17721 ) );
NAND2_X1 _u10_U6301  ( .A1(1'b1), .A2(_u10_n12101 ), .ZN(_u10_n17722 ) );
NAND2_X1 _u10_U6300  ( .A1(1'b1), .A2(_u10_n12077 ), .ZN(_u10_n17723 ) );
NAND4_X1 _u10_U6299  ( .A1(_u10_n17720 ), .A2(_u10_n17721 ), .A3(_u10_n17722 ), .A4(_u10_n17723 ), .ZN(_u10_n17715 ) );
NAND2_X1 _u10_U6298  ( .A1(1'b1), .A2(_u10_n12053 ), .ZN(_u10_n17717 ) );
NAND2_X1 _u10_U6297  ( .A1(1'b1), .A2(_u10_n12029 ), .ZN(_u10_n17718 ) );
NAND2_X1 _u10_U6296  ( .A1(1'b1), .A2(_u10_n12009 ), .ZN(_u10_n17719 ) );
NAND3_X1 _u10_U6295  ( .A1(_u10_n17717 ), .A2(_u10_n17718 ), .A3(_u10_n17719 ), .ZN(_u10_n17716 ) );
NOR4_X1 _u10_U6294  ( .A1(_u10_n17713 ), .A2(_u10_n17714 ), .A3(_u10_n17715 ), .A4(_u10_n17716 ), .ZN(_u10_n17691 ) );
NAND2_X1 _u10_U6293  ( .A1(1'b1), .A2(_u10_n11993 ), .ZN(_u10_n17709 ) );
NAND2_X1 _u10_U6292  ( .A1(1'b1), .A2(_u10_n11969 ), .ZN(_u10_n17710 ) );
NAND2_X1 _u10_U6291  ( .A1(1'b1), .A2(_u10_n11945 ), .ZN(_u10_n17711 ) );
NAND2_X1 _u10_U6290  ( .A1(1'b1), .A2(_u10_n11921 ), .ZN(_u10_n17712 ) );
NAND4_X1 _u10_U6289  ( .A1(_u10_n17709 ), .A2(_u10_n17710 ), .A3(_u10_n17711 ), .A4(_u10_n17712 ), .ZN(_u10_n17693 ) );
NAND2_X1 _u10_U6288  ( .A1(1'b1), .A2(_u10_n11897 ), .ZN(_u10_n17705 ) );
NAND2_X1 _u10_U6287  ( .A1(1'b1), .A2(_u10_n11873 ), .ZN(_u10_n17706 ) );
NAND2_X1 _u10_U6286  ( .A1(1'b1), .A2(_u10_n11849 ), .ZN(_u10_n17707 ) );
NAND2_X1 _u10_U6285  ( .A1(1'b1), .A2(_u10_n11825 ), .ZN(_u10_n17708 ) );
NAND4_X1 _u10_U6284  ( .A1(_u10_n17705 ), .A2(_u10_n17706 ), .A3(_u10_n17707 ), .A4(_u10_n17708 ), .ZN(_u10_n17694 ) );
NAND2_X1 _u10_U6283  ( .A1(1'b1), .A2(_u10_n11801 ), .ZN(_u10_n17701 ) );
NAND2_X1 _u10_U6282  ( .A1(1'b1), .A2(_u10_n11777 ), .ZN(_u10_n17702 ) );
NAND2_X1 _u10_U6281  ( .A1(1'b1), .A2(_u10_n11753 ), .ZN(_u10_n17703 ) );
NAND2_X1 _u10_U6280  ( .A1(1'b1), .A2(_u10_n11729 ), .ZN(_u10_n17704 ) );
NAND4_X1 _u10_U6279  ( .A1(_u10_n17701 ), .A2(_u10_n17702 ), .A3(_u10_n17703 ), .A4(_u10_n17704 ), .ZN(_u10_n17695 ) );
NAND2_X1 _u10_U6278  ( .A1(1'b1), .A2(_u10_n11705 ), .ZN(_u10_n17697 ) );
NAND2_X1 _u10_U6277  ( .A1(1'b1), .A2(_u10_n11681 ), .ZN(_u10_n17698 ) );
NAND2_X1 _u10_U6276  ( .A1(1'b1), .A2(_u10_n11657 ), .ZN(_u10_n17699 ) );
NAND2_X1 _u10_U6275  ( .A1(1'b1), .A2(_u10_n11633 ), .ZN(_u10_n17700 ) );
NAND4_X1 _u10_U6274  ( .A1(_u10_n17697 ), .A2(_u10_n17698 ), .A3(_u10_n17699 ), .A4(_u10_n17700 ), .ZN(_u10_n17696 ) );
NOR4_X1 _u10_U6273  ( .A1(_u10_n17693 ), .A2(_u10_n17694 ), .A3(_u10_n17695 ), .A4(_u10_n17696 ), .ZN(_u10_n17692 ) );
NAND2_X1 _u10_U6272  ( .A1(_u10_n17691 ), .A2(_u10_n17692 ), .ZN(am1[9]) );
NAND2_X1 _u10_U6271  ( .A1(1'b0), .A2(_u10_n12340 ), .ZN(_u10_n17687 ) );
NAND2_X1 _u10_U6270  ( .A1(1'b0), .A2(_u10_n12316 ), .ZN(_u10_n17688 ) );
NAND2_X1 _u10_U6269  ( .A1(1'b0), .A2(_u10_n12293 ), .ZN(_u10_n17689 ) );
NAND2_X1 _u10_U6268  ( .A1(1'b0), .A2(_u10_n12269 ), .ZN(_u10_n17690 ) );
NAND4_X1 _u10_U6267  ( .A1(_u10_n17687 ), .A2(_u10_n17688 ), .A3(_u10_n17689 ), .A4(_u10_n17690 ), .ZN(_u10_n17672 ) );
NAND2_X1 _u10_U6266  ( .A1(1'b0), .A2(_u10_n12244 ), .ZN(_u10_n17683 ) );
NAND2_X1 _u10_U6265  ( .A1(1'b0), .A2(_u10_n12220 ), .ZN(_u10_n17684 ) );
NAND2_X1 _u10_U6264  ( .A1(1'b0), .A2(_u10_n12197 ), .ZN(_u10_n17685 ) );
NAND2_X1 _u10_U6263  ( .A1(1'b0), .A2(_u10_n12172 ), .ZN(_u10_n17686 ) );
NAND4_X1 _u10_U6262  ( .A1(_u10_n17683 ), .A2(_u10_n17684 ), .A3(_u10_n17685 ), .A4(_u10_n17686 ), .ZN(_u10_n17673 ) );
NAND2_X1 _u10_U6261  ( .A1(1'b0), .A2(_u10_n12149 ), .ZN(_u10_n17679 ) );
NAND2_X1 _u10_U6260  ( .A1(1'b0), .A2(_u10_n12125 ), .ZN(_u10_n17680 ) );
NAND2_X1 _u10_U6259  ( .A1(1'b0), .A2(_u10_n12101 ), .ZN(_u10_n17681 ) );
NAND2_X1 _u10_U6258  ( .A1(1'b0), .A2(_u10_n12077 ), .ZN(_u10_n17682 ) );
NAND4_X1 _u10_U6257  ( .A1(_u10_n17679 ), .A2(_u10_n17680 ), .A3(_u10_n17681 ), .A4(_u10_n17682 ), .ZN(_u10_n17674 ) );
NAND2_X1 _u10_U6256  ( .A1(1'b0), .A2(_u10_n12053 ), .ZN(_u10_n17676 ) );
NAND2_X1 _u10_U6255  ( .A1(1'b0), .A2(_u10_n12029 ), .ZN(_u10_n17677 ) );
NAND2_X1 _u10_U6254  ( .A1(ch0_csr[0]), .A2(_u10_n12009 ), .ZN(_u10_n17678 ));
NAND3_X1 _u10_U6253  ( .A1(_u10_n17676 ), .A2(_u10_n17677 ), .A3(_u10_n17678 ), .ZN(_u10_n17675 ) );
NOR4_X1 _u10_U6252  ( .A1(_u10_n17672 ), .A2(_u10_n17673 ), .A3(_u10_n17674 ), .A4(_u10_n17675 ), .ZN(_u10_n17650 ) );
NAND2_X1 _u10_U6251  ( .A1(1'b0), .A2(_u10_n11993 ), .ZN(_u10_n17668 ) );
NAND2_X1 _u10_U6250  ( .A1(1'b0), .A2(_u10_n11969 ), .ZN(_u10_n17669 ) );
NAND2_X1 _u10_U6249  ( .A1(1'b0), .A2(_u10_n11945 ), .ZN(_u10_n17670 ) );
NAND2_X1 _u10_U6248  ( .A1(1'b0), .A2(_u10_n11921 ), .ZN(_u10_n17671 ) );
NAND4_X1 _u10_U6247  ( .A1(_u10_n17668 ), .A2(_u10_n17669 ), .A3(_u10_n17670 ), .A4(_u10_n17671 ), .ZN(_u10_n17652 ) );
NAND2_X1 _u10_U6246  ( .A1(1'b0), .A2(_u10_n11897 ), .ZN(_u10_n17664 ) );
NAND2_X1 _u10_U6245  ( .A1(1'b0), .A2(_u10_n11873 ), .ZN(_u10_n17665 ) );
NAND2_X1 _u10_U6244  ( .A1(1'b0), .A2(_u10_n11849 ), .ZN(_u10_n17666 ) );
NAND2_X1 _u10_U6243  ( .A1(1'b0), .A2(_u10_n11825 ), .ZN(_u10_n17667 ) );
NAND4_X1 _u10_U6242  ( .A1(_u10_n17664 ), .A2(_u10_n17665 ), .A3(_u10_n17666 ), .A4(_u10_n17667 ), .ZN(_u10_n17653 ) );
NAND2_X1 _u10_U6241  ( .A1(1'b0), .A2(_u10_n11801 ), .ZN(_u10_n17660 ) );
NAND2_X1 _u10_U6240  ( .A1(1'b0), .A2(_u10_n11777 ), .ZN(_u10_n17661 ) );
NAND2_X1 _u10_U6239  ( .A1(1'b0), .A2(_u10_n11753 ), .ZN(_u10_n17662 ) );
NAND2_X1 _u10_U6238  ( .A1(1'b0), .A2(_u10_n11729 ), .ZN(_u10_n17663 ) );
NAND4_X1 _u10_U6237  ( .A1(_u10_n17660 ), .A2(_u10_n17661 ), .A3(_u10_n17662 ), .A4(_u10_n17663 ), .ZN(_u10_n17654 ) );
NAND2_X1 _u10_U6236  ( .A1(1'b0), .A2(_u10_n11705 ), .ZN(_u10_n17656 ) );
NAND2_X1 _u10_U6235  ( .A1(1'b0), .A2(_u10_n11681 ), .ZN(_u10_n17657 ) );
NAND2_X1 _u10_U6234  ( .A1(1'b0), .A2(_u10_n11657 ), .ZN(_u10_n17658 ) );
NAND2_X1 _u10_U6233  ( .A1(1'b0), .A2(_u10_n11633 ), .ZN(_u10_n17659 ) );
NAND4_X1 _u10_U6232  ( .A1(_u10_n17656 ), .A2(_u10_n17657 ), .A3(_u10_n17658 ), .A4(_u10_n17659 ), .ZN(_u10_n17655 ) );
NOR4_X1 _u10_U6231  ( .A1(_u10_n17652 ), .A2(_u10_n17653 ), .A3(_u10_n17654 ), .A4(_u10_n17655 ), .ZN(_u10_n17651 ) );
NAND2_X1 _u10_U6230  ( .A1(_u10_n17650 ), .A2(_u10_n17651 ), .ZN(csr[0]) );
NAND2_X1 _u10_U6229  ( .A1(1'b0), .A2(_u10_n12340 ), .ZN(_u10_n17646 ) );
NAND2_X1 _u10_U6228  ( .A1(1'b0), .A2(_u10_n12316 ), .ZN(_u10_n17647 ) );
NAND2_X1 _u10_U6227  ( .A1(1'b0), .A2(_u10_n12293 ), .ZN(_u10_n17648 ) );
NAND2_X1 _u10_U6226  ( .A1(1'b0), .A2(_u10_n12269 ), .ZN(_u10_n17649 ) );
NAND4_X1 _u10_U6225  ( .A1(_u10_n17646 ), .A2(_u10_n17647 ), .A3(_u10_n17648 ), .A4(_u10_n17649 ), .ZN(_u10_n17631 ) );
NAND2_X1 _u10_U6224  ( .A1(1'b0), .A2(_u10_n12244 ), .ZN(_u10_n17642 ) );
NAND2_X1 _u10_U6223  ( .A1(1'b0), .A2(_u10_n12220 ), .ZN(_u10_n17643 ) );
NAND2_X1 _u10_U6222  ( .A1(1'b0), .A2(_u10_n12197 ), .ZN(_u10_n17644 ) );
NAND2_X1 _u10_U6221  ( .A1(1'b0), .A2(_u10_n12172 ), .ZN(_u10_n17645 ) );
NAND4_X1 _u10_U6220  ( .A1(_u10_n17642 ), .A2(_u10_n17643 ), .A3(_u10_n17644 ), .A4(_u10_n17645 ), .ZN(_u10_n17632 ) );
NAND2_X1 _u10_U6219  ( .A1(1'b0), .A2(_u10_n12149 ), .ZN(_u10_n17638 ) );
NAND2_X1 _u10_U6218  ( .A1(1'b0), .A2(_u10_n12125 ), .ZN(_u10_n17639 ) );
NAND2_X1 _u10_U6217  ( .A1(1'b0), .A2(_u10_n12101 ), .ZN(_u10_n17640 ) );
NAND2_X1 _u10_U6216  ( .A1(1'b0), .A2(_u10_n12077 ), .ZN(_u10_n17641 ) );
NAND4_X1 _u10_U6215  ( .A1(_u10_n17638 ), .A2(_u10_n17639 ), .A3(_u10_n17640 ), .A4(_u10_n17641 ), .ZN(_u10_n17633 ) );
NAND2_X1 _u10_U6214  ( .A1(1'b0), .A2(_u10_n12053 ), .ZN(_u10_n17635 ) );
NAND2_X1 _u10_U6213  ( .A1(1'b0), .A2(_u10_n12029 ), .ZN(_u10_n17636 ) );
NAND2_X1 _u10_U6212  ( .A1(ch0_csr[10]), .A2(_u10_n12009 ), .ZN(_u10_n17637 ) );
NAND3_X1 _u10_U6211  ( .A1(_u10_n17635 ), .A2(_u10_n17636 ), .A3(_u10_n17637 ), .ZN(_u10_n17634 ) );
NOR4_X1 _u10_U6210  ( .A1(_u10_n17631 ), .A2(_u10_n17632 ), .A3(_u10_n17633 ), .A4(_u10_n17634 ), .ZN(_u10_n17609 ) );
NAND2_X1 _u10_U6209  ( .A1(1'b0), .A2(_u10_n11998 ), .ZN(_u10_n17627 ) );
NAND2_X1 _u10_U6208  ( .A1(1'b0), .A2(_u10_n11970 ), .ZN(_u10_n17628 ) );
NAND2_X1 _u10_U6207  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n17629 ) );
NAND2_X1 _u10_U6206  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n17630 ) );
NAND4_X1 _u10_U6205  ( .A1(_u10_n17627 ), .A2(_u10_n17628 ), .A3(_u10_n17629 ), .A4(_u10_n17630 ), .ZN(_u10_n17611 ) );
NAND2_X1 _u10_U6204  ( .A1(1'b0), .A2(_u10_n11902 ), .ZN(_u10_n17623 ) );
NAND2_X1 _u10_U6203  ( .A1(1'b0), .A2(_u10_n11878 ), .ZN(_u10_n17624 ) );
NAND2_X1 _u10_U6202  ( .A1(1'b0), .A2(_u10_n11851 ), .ZN(_u10_n17625 ) );
NAND2_X1 _u10_U6201  ( .A1(1'b0), .A2(_u10_n11830 ), .ZN(_u10_n17626 ) );
NAND4_X1 _u10_U6200  ( .A1(_u10_n17623 ), .A2(_u10_n17624 ), .A3(_u10_n17625 ), .A4(_u10_n17626 ), .ZN(_u10_n17612 ) );
NAND2_X1 _u10_U6199  ( .A1(1'b0), .A2(_u10_n11806 ), .ZN(_u10_n17619 ) );
NAND2_X1 _u10_U6198  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n17620 ) );
NAND2_X1 _u10_U6197  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n17621 ) );
NAND2_X1 _u10_U6196  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n17622 ) );
NAND4_X1 _u10_U6195  ( .A1(_u10_n17619 ), .A2(_u10_n17620 ), .A3(_u10_n17621 ), .A4(_u10_n17622 ), .ZN(_u10_n17613 ) );
NAND2_X1 _u10_U6194  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n17615 ) );
NAND2_X1 _u10_U6193  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n17616 ) );
NAND2_X1 _u10_U6192  ( .A1(1'b0), .A2(_u10_n11659 ), .ZN(_u10_n17617 ) );
NAND2_X1 _u10_U6191  ( .A1(1'b0), .A2(_u10_n11635 ), .ZN(_u10_n17618 ) );
NAND4_X1 _u10_U6190  ( .A1(_u10_n17615 ), .A2(_u10_n17616 ), .A3(_u10_n17617 ), .A4(_u10_n17618 ), .ZN(_u10_n17614 ) );
NOR4_X1 _u10_U6189  ( .A1(_u10_n17611 ), .A2(_u10_n17612 ), .A3(_u10_n17613 ), .A4(_u10_n17614 ), .ZN(_u10_n17610 ) );
NAND2_X1 _u10_U6188  ( .A1(_u10_n17609 ), .A2(_u10_n17610 ), .ZN(csr[10]) );
NAND2_X1 _u10_U6187  ( .A1(1'b0), .A2(_u10_n12340 ), .ZN(_u10_n17605 ) );
NAND2_X1 _u10_U6186  ( .A1(1'b0), .A2(_u10_n12316 ), .ZN(_u10_n17606 ) );
NAND2_X1 _u10_U6185  ( .A1(1'b0), .A2(_u10_n12293 ), .ZN(_u10_n17607 ) );
NAND2_X1 _u10_U6184  ( .A1(1'b0), .A2(_u10_n12269 ), .ZN(_u10_n17608 ) );
NAND4_X1 _u10_U6183  ( .A1(_u10_n17605 ), .A2(_u10_n17606 ), .A3(_u10_n17607 ), .A4(_u10_n17608 ), .ZN(_u10_n17590 ) );
NAND2_X1 _u10_U6182  ( .A1(1'b0), .A2(_u10_n12244 ), .ZN(_u10_n17601 ) );
NAND2_X1 _u10_U6181  ( .A1(1'b0), .A2(_u10_n12220 ), .ZN(_u10_n17602 ) );
NAND2_X1 _u10_U6180  ( .A1(1'b0), .A2(_u10_n12197 ), .ZN(_u10_n17603 ) );
NAND2_X1 _u10_U6179  ( .A1(1'b0), .A2(_u10_n12172 ), .ZN(_u10_n17604 ) );
NAND4_X1 _u10_U6178  ( .A1(_u10_n17601 ), .A2(_u10_n17602 ), .A3(_u10_n17603 ), .A4(_u10_n17604 ), .ZN(_u10_n17591 ) );
NAND2_X1 _u10_U6177  ( .A1(1'b0), .A2(_u10_n12149 ), .ZN(_u10_n17597 ) );
NAND2_X1 _u10_U6176  ( .A1(1'b0), .A2(_u10_n12125 ), .ZN(_u10_n17598 ) );
NAND2_X1 _u10_U6175  ( .A1(1'b0), .A2(_u10_n12101 ), .ZN(_u10_n17599 ) );
NAND2_X1 _u10_U6174  ( .A1(1'b0), .A2(_u10_n12077 ), .ZN(_u10_n17600 ) );
NAND4_X1 _u10_U6173  ( .A1(_u10_n17597 ), .A2(_u10_n17598 ), .A3(_u10_n17599 ), .A4(_u10_n17600 ), .ZN(_u10_n17592 ) );
NAND2_X1 _u10_U6172  ( .A1(1'b0), .A2(_u10_n12053 ), .ZN(_u10_n17594 ) );
NAND2_X1 _u10_U6171  ( .A1(1'b0), .A2(_u10_n12029 ), .ZN(_u10_n17595 ) );
NAND2_X1 _u10_U6170  ( .A1(ch0_csr[11]), .A2(_u10_n12009 ), .ZN(_u10_n17596 ) );
NAND3_X1 _u10_U6169  ( .A1(_u10_n17594 ), .A2(_u10_n17595 ), .A3(_u10_n17596 ), .ZN(_u10_n17593 ) );
NOR4_X1 _u10_U6168  ( .A1(_u10_n17590 ), .A2(_u10_n17591 ), .A3(_u10_n17592 ), .A4(_u10_n17593 ), .ZN(_u10_n17568 ) );
NAND2_X1 _u10_U6167  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n17586 ) );
NAND2_X1 _u10_U6166  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n17587 ) );
NAND2_X1 _u10_U6165  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n17588 ) );
NAND2_X1 _u10_U6164  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n17589 ) );
NAND4_X1 _u10_U6163  ( .A1(_u10_n17586 ), .A2(_u10_n17587 ), .A3(_u10_n17588 ), .A4(_u10_n17589 ), .ZN(_u10_n17570 ) );
NAND2_X1 _u10_U6162  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n17582 ) );
NAND2_X1 _u10_U6161  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n17583 ) );
NAND2_X1 _u10_U6160  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n17584 ) );
NAND2_X1 _u10_U6159  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n17585 ) );
NAND4_X1 _u10_U6158  ( .A1(_u10_n17582 ), .A2(_u10_n17583 ), .A3(_u10_n17584 ), .A4(_u10_n17585 ), .ZN(_u10_n17571 ) );
NAND2_X1 _u10_U6157  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n17578 ) );
NAND2_X1 _u10_U6156  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n17579 ) );
NAND2_X1 _u10_U6155  ( .A1(1'b0), .A2(_u10_n11754 ), .ZN(_u10_n17580 ) );
NAND2_X1 _u10_U6154  ( .A1(1'b0), .A2(_u10_n11731 ), .ZN(_u10_n17581 ) );
NAND4_X1 _u10_U6153  ( .A1(_u10_n17578 ), .A2(_u10_n17579 ), .A3(_u10_n17580 ), .A4(_u10_n17581 ), .ZN(_u10_n17572 ) );
NAND2_X1 _u10_U6152  ( .A1(1'b0), .A2(_u10_n11706 ), .ZN(_u10_n17574 ) );
NAND2_X1 _u10_U6151  ( .A1(1'b0), .A2(_u10_n11683 ), .ZN(_u10_n17575 ) );
NAND2_X1 _u10_U6150  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n17576 ) );
NAND2_X1 _u10_U6149  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n17577 ) );
NAND4_X1 _u10_U6148  ( .A1(_u10_n17574 ), .A2(_u10_n17575 ), .A3(_u10_n17576 ), .A4(_u10_n17577 ), .ZN(_u10_n17573 ) );
NOR4_X1 _u10_U6147  ( .A1(_u10_n17570 ), .A2(_u10_n17571 ), .A3(_u10_n17572 ), .A4(_u10_n17573 ), .ZN(_u10_n17569 ) );
NAND2_X1 _u10_U6146  ( .A1(_u10_n17568 ), .A2(_u10_n17569 ), .ZN(csr[11]) );
NAND2_X1 _u10_U6145  ( .A1(1'b0), .A2(_u10_n12340 ), .ZN(_u10_n17564 ) );
NAND2_X1 _u10_U6144  ( .A1(1'b0), .A2(_u10_n12316 ), .ZN(_u10_n17565 ) );
NAND2_X1 _u10_U6143  ( .A1(1'b0), .A2(_u10_n12293 ), .ZN(_u10_n17566 ) );
NAND2_X1 _u10_U6142  ( .A1(1'b0), .A2(_u10_n12269 ), .ZN(_u10_n17567 ) );
NAND4_X1 _u10_U6141  ( .A1(_u10_n17564 ), .A2(_u10_n17565 ), .A3(_u10_n17566 ), .A4(_u10_n17567 ), .ZN(_u10_n17549 ) );
NAND2_X1 _u10_U6140  ( .A1(1'b0), .A2(_u10_n12244 ), .ZN(_u10_n17560 ) );
NAND2_X1 _u10_U6139  ( .A1(1'b0), .A2(_u10_n12220 ), .ZN(_u10_n17561 ) );
NAND2_X1 _u10_U6138  ( .A1(1'b0), .A2(_u10_n12197 ), .ZN(_u10_n17562 ) );
NAND2_X1 _u10_U6137  ( .A1(1'b0), .A2(_u10_n12172 ), .ZN(_u10_n17563 ) );
NAND4_X1 _u10_U6136  ( .A1(_u10_n17560 ), .A2(_u10_n17561 ), .A3(_u10_n17562 ), .A4(_u10_n17563 ), .ZN(_u10_n17550 ) );
NAND2_X1 _u10_U6135  ( .A1(1'b0), .A2(_u10_n12149 ), .ZN(_u10_n17556 ) );
NAND2_X1 _u10_U6134  ( .A1(1'b0), .A2(_u10_n12125 ), .ZN(_u10_n17557 ) );
NAND2_X1 _u10_U6133  ( .A1(1'b0), .A2(_u10_n12101 ), .ZN(_u10_n17558 ) );
NAND2_X1 _u10_U6132  ( .A1(1'b0), .A2(_u10_n12077 ), .ZN(_u10_n17559 ) );
NAND4_X1 _u10_U6131  ( .A1(_u10_n17556 ), .A2(_u10_n17557 ), .A3(_u10_n17558 ), .A4(_u10_n17559 ), .ZN(_u10_n17551 ) );
NAND2_X1 _u10_U6130  ( .A1(1'b0), .A2(_u10_n12053 ), .ZN(_u10_n17553 ) );
NAND2_X1 _u10_U6129  ( .A1(1'b0), .A2(_u10_n12029 ), .ZN(_u10_n17554 ) );
NAND2_X1 _u10_U6128  ( .A1(ch0_csr[12]), .A2(_u10_n12010 ), .ZN(_u10_n17555 ) );
NAND3_X1 _u10_U6127  ( .A1(_u10_n17553 ), .A2(_u10_n17554 ), .A3(_u10_n17555 ), .ZN(_u10_n17552 ) );
NOR4_X1 _u10_U6126  ( .A1(_u10_n17549 ), .A2(_u10_n17550 ), .A3(_u10_n17551 ), .A4(_u10_n17552 ), .ZN(_u10_n17527 ) );
NAND2_X1 _u10_U6125  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n17545 ) );
NAND2_X1 _u10_U6124  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n17546 ) );
NAND2_X1 _u10_U6123  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n17547 ) );
NAND2_X1 _u10_U6122  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n17548 ) );
NAND4_X1 _u10_U6121  ( .A1(_u10_n17545 ), .A2(_u10_n17546 ), .A3(_u10_n17547 ), .A4(_u10_n17548 ), .ZN(_u10_n17529 ) );
NAND2_X1 _u10_U6120  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n17541 ) );
NAND2_X1 _u10_U6119  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n17542 ) );
NAND2_X1 _u10_U6118  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n17543 ) );
NAND2_X1 _u10_U6117  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n17544 ) );
NAND4_X1 _u10_U6116  ( .A1(_u10_n17541 ), .A2(_u10_n17542 ), .A3(_u10_n17543 ), .A4(_u10_n17544 ), .ZN(_u10_n17530 ) );
NAND2_X1 _u10_U6115  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n17537 ) );
NAND2_X1 _u10_U6114  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n17538 ) );
NAND2_X1 _u10_U6113  ( .A1(1'b0), .A2(_u10_n11759 ), .ZN(_u10_n17539 ) );
NAND2_X1 _u10_U6112  ( .A1(1'b0), .A2(_u10_n11730 ), .ZN(_u10_n17540 ) );
NAND4_X1 _u10_U6111  ( .A1(_u10_n17537 ), .A2(_u10_n17538 ), .A3(_u10_n17539 ), .A4(_u10_n17540 ), .ZN(_u10_n17531 ) );
NAND2_X1 _u10_U6110  ( .A1(1'b0), .A2(_u10_n11711 ), .ZN(_u10_n17533 ) );
NAND2_X1 _u10_U6109  ( .A1(1'b0), .A2(_u10_n11682 ), .ZN(_u10_n17534 ) );
NAND2_X1 _u10_U6108  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n17535 ) );
NAND2_X1 _u10_U6107  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n17536 ) );
NAND4_X1 _u10_U6106  ( .A1(_u10_n17533 ), .A2(_u10_n17534 ), .A3(_u10_n17535 ), .A4(_u10_n17536 ), .ZN(_u10_n17532 ) );
NOR4_X1 _u10_U6105  ( .A1(_u10_n17529 ), .A2(_u10_n17530 ), .A3(_u10_n17531 ), .A4(_u10_n17532 ), .ZN(_u10_n17528 ) );
NAND2_X1 _u10_U6104  ( .A1(_u10_n17527 ), .A2(_u10_n17528 ), .ZN(csr[12]) );
NAND2_X1 _u10_U6103  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17523 ) );
NAND2_X1 _u10_U6102  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17524 ) );
NAND2_X1 _u10_U6101  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17525 ) );
NAND2_X1 _u10_U6100  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17526 ) );
NAND4_X1 _u10_U6099  ( .A1(_u10_n17523 ), .A2(_u10_n17524 ), .A3(_u10_n17525 ), .A4(_u10_n17526 ), .ZN(_u10_n17508 ) );
NAND2_X1 _u10_U6098  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17519 ) );
NAND2_X1 _u10_U6097  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17520 ) );
NAND2_X1 _u10_U6096  ( .A1(1'b0), .A2(_u10_n12420 ), .ZN(_u10_n17521 ) );
NAND2_X1 _u10_U6095  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17522 ) );
NAND4_X1 _u10_U6094  ( .A1(_u10_n17519 ), .A2(_u10_n17520 ), .A3(_u10_n17521 ), .A4(_u10_n17522 ), .ZN(_u10_n17509 ) );
NAND2_X1 _u10_U6093  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17515 ) );
NAND2_X1 _u10_U6092  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17516 ) );
NAND2_X1 _u10_U6091  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17517 ) );
NAND2_X1 _u10_U6090  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17518 ) );
NAND4_X1 _u10_U6089  ( .A1(_u10_n17515 ), .A2(_u10_n17516 ), .A3(_u10_n17517 ), .A4(_u10_n17518 ), .ZN(_u10_n17510 ) );
NAND2_X1 _u10_U6088  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17512 ) );
NAND2_X1 _u10_U6087  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17513 ) );
NAND2_X1 _u10_U6086  ( .A1(ch0_csr[13]), .A2(_u10_n12010 ), .ZN(_u10_n17514 ) );
NAND3_X1 _u10_U6085  ( .A1(_u10_n17512 ), .A2(_u10_n17513 ), .A3(_u10_n17514 ), .ZN(_u10_n17511 ) );
NOR4_X1 _u10_U6084  ( .A1(_u10_n17508 ), .A2(_u10_n17509 ), .A3(_u10_n17510 ), .A4(_u10_n17511 ), .ZN(_u10_n17486 ) );
NAND2_X1 _u10_U6083  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n17504 ) );
NAND2_X1 _u10_U6082  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n17505 ) );
NAND2_X1 _u10_U6081  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n17506 ) );
NAND2_X1 _u10_U6080  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n17507 ) );
NAND4_X1 _u10_U6079  ( .A1(_u10_n17504 ), .A2(_u10_n17505 ), .A3(_u10_n17506 ), .A4(_u10_n17507 ), .ZN(_u10_n17488 ) );
NAND2_X1 _u10_U6078  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n17500 ) );
NAND2_X1 _u10_U6077  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n17501 ) );
NAND2_X1 _u10_U6076  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n17502 ) );
NAND2_X1 _u10_U6075  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n17503 ) );
NAND4_X1 _u10_U6074  ( .A1(_u10_n17500 ), .A2(_u10_n17501 ), .A3(_u10_n17502 ), .A4(_u10_n17503 ), .ZN(_u10_n17489 ) );
NAND2_X1 _u10_U6073  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n17496 ) );
NAND2_X1 _u10_U6072  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n17497 ) );
NAND2_X1 _u10_U6071  ( .A1(1'b0), .A2(_u10_n12378 ), .ZN(_u10_n17498 ) );
NAND2_X1 _u10_U6070  ( .A1(1'b0), .A2(_u10_n12377 ), .ZN(_u10_n17499 ) );
NAND4_X1 _u10_U6069  ( .A1(_u10_n17496 ), .A2(_u10_n17497 ), .A3(_u10_n17498 ), .A4(_u10_n17499 ), .ZN(_u10_n17490 ) );
NAND2_X1 _u10_U6068  ( .A1(1'b0), .A2(_u10_n12372 ), .ZN(_u10_n17492 ) );
NAND2_X1 _u10_U6067  ( .A1(1'b0), .A2(_u10_n12371 ), .ZN(_u10_n17493 ) );
NAND2_X1 _u10_U6066  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n17494 ) );
NAND2_X1 _u10_U6065  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n17495 ) );
NAND4_X1 _u10_U6064  ( .A1(_u10_n17492 ), .A2(_u10_n17493 ), .A3(_u10_n17494 ), .A4(_u10_n17495 ), .ZN(_u10_n17491 ) );
NOR4_X1 _u10_U6063  ( .A1(_u10_n17488 ), .A2(_u10_n17489 ), .A3(_u10_n17490 ), .A4(_u10_n17491 ), .ZN(_u10_n17487 ) );
NAND2_X1 _u10_U6062  ( .A1(_u10_n17486 ), .A2(_u10_n17487 ), .ZN(csr[13]) );
NAND2_X1 _u10_U6061  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17482 ) );
NAND2_X1 _u10_U6060  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17483 ) );
NAND2_X1 _u10_U6059  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17484 ) );
NAND2_X1 _u10_U6058  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17485 ) );
NAND4_X1 _u10_U6057  ( .A1(_u10_n17482 ), .A2(_u10_n17483 ), .A3(_u10_n17484 ), .A4(_u10_n17485 ), .ZN(_u10_n17467 ) );
NAND2_X1 _u10_U6056  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17478 ) );
NAND2_X1 _u10_U6055  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17479 ) );
NAND2_X1 _u10_U6054  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n17480 ) );
NAND2_X1 _u10_U6053  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17481 ) );
NAND4_X1 _u10_U6052  ( .A1(_u10_n17478 ), .A2(_u10_n17479 ), .A3(_u10_n17480 ), .A4(_u10_n17481 ), .ZN(_u10_n17468 ) );
NAND2_X1 _u10_U6051  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17474 ) );
NAND2_X1 _u10_U6050  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17475 ) );
NAND2_X1 _u10_U6049  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17476 ) );
NAND2_X1 _u10_U6048  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17477 ) );
NAND4_X1 _u10_U6047  ( .A1(_u10_n17474 ), .A2(_u10_n17475 ), .A3(_u10_n17476 ), .A4(_u10_n17477 ), .ZN(_u10_n17469 ) );
NAND2_X1 _u10_U6046  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17471 ) );
NAND2_X1 _u10_U6045  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17472 ) );
NAND2_X1 _u10_U6044  ( .A1(ch0_csr[14]), .A2(_u10_n12010 ), .ZN(_u10_n17473 ) );
NAND3_X1 _u10_U6043  ( .A1(_u10_n17471 ), .A2(_u10_n17472 ), .A3(_u10_n17473 ), .ZN(_u10_n17470 ) );
NOR4_X1 _u10_U6042  ( .A1(_u10_n17467 ), .A2(_u10_n17468 ), .A3(_u10_n17469 ), .A4(_u10_n17470 ), .ZN(_u10_n17445 ) );
NAND2_X1 _u10_U6041  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n17463 ) );
NAND2_X1 _u10_U6040  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n17464 ) );
NAND2_X1 _u10_U6039  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n17465 ) );
NAND2_X1 _u10_U6038  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n17466 ) );
NAND4_X1 _u10_U6037  ( .A1(_u10_n17463 ), .A2(_u10_n17464 ), .A3(_u10_n17465 ), .A4(_u10_n17466 ), .ZN(_u10_n17447 ) );
NAND2_X1 _u10_U6036  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n17459 ) );
NAND2_X1 _u10_U6035  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n17460 ) );
NAND2_X1 _u10_U6034  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n17461 ) );
NAND2_X1 _u10_U6033  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n17462 ) );
NAND4_X1 _u10_U6032  ( .A1(_u10_n17459 ), .A2(_u10_n17460 ), .A3(_u10_n17461 ), .A4(_u10_n17462 ), .ZN(_u10_n17448 ) );
NAND2_X1 _u10_U6031  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n17455 ) );
NAND2_X1 _u10_U6030  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n17456 ) );
NAND2_X1 _u10_U6029  ( .A1(1'b0), .A2(_u10_n11755 ), .ZN(_u10_n17457 ) );
NAND2_X1 _u10_U6028  ( .A1(1'b0), .A2(_u10_n11735 ), .ZN(_u10_n17458 ) );
NAND4_X1 _u10_U6027  ( .A1(_u10_n17455 ), .A2(_u10_n17456 ), .A3(_u10_n17457 ), .A4(_u10_n17458 ), .ZN(_u10_n17449 ) );
NAND2_X1 _u10_U6026  ( .A1(1'b0), .A2(_u10_n11707 ), .ZN(_u10_n17451 ) );
NAND2_X1 _u10_U6025  ( .A1(1'b0), .A2(_u10_n11687 ), .ZN(_u10_n17452 ) );
NAND2_X1 _u10_U6024  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n17453 ) );
NAND2_X1 _u10_U6023  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n17454 ) );
NAND4_X1 _u10_U6022  ( .A1(_u10_n17451 ), .A2(_u10_n17452 ), .A3(_u10_n17453 ), .A4(_u10_n17454 ), .ZN(_u10_n17450 ) );
NOR4_X1 _u10_U6021  ( .A1(_u10_n17447 ), .A2(_u10_n17448 ), .A3(_u10_n17449 ), .A4(_u10_n17450 ), .ZN(_u10_n17446 ) );
NAND2_X1 _u10_U6020  ( .A1(_u10_n17445 ), .A2(_u10_n17446 ), .ZN(csr[14]) );
NAND2_X1 _u10_U6019  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17441 ) );
NAND2_X1 _u10_U6018  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17442 ) );
NAND2_X1 _u10_U6017  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17443 ) );
NAND2_X1 _u10_U6016  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17444 ) );
NAND4_X1 _u10_U6015  ( .A1(_u10_n17441 ), .A2(_u10_n17442 ), .A3(_u10_n17443 ), .A4(_u10_n17444 ), .ZN(_u10_n17426 ) );
NAND2_X1 _u10_U6014  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17437 ) );
NAND2_X1 _u10_U6013  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17438 ) );
NAND2_X1 _u10_U6012  ( .A1(1'b0), .A2(_u10_n12206 ), .ZN(_u10_n17439 ) );
NAND2_X1 _u10_U6011  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17440 ) );
NAND4_X1 _u10_U6010  ( .A1(_u10_n17437 ), .A2(_u10_n17438 ), .A3(_u10_n17439 ), .A4(_u10_n17440 ), .ZN(_u10_n17427 ) );
NAND2_X1 _u10_U6009  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17433 ) );
NAND2_X1 _u10_U6008  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17434 ) );
NAND2_X1 _u10_U6007  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17435 ) );
NAND2_X1 _u10_U6006  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17436 ) );
NAND4_X1 _u10_U6005  ( .A1(_u10_n17433 ), .A2(_u10_n17434 ), .A3(_u10_n17435 ), .A4(_u10_n17436 ), .ZN(_u10_n17428 ) );
NAND2_X1 _u10_U6004  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17430 ) );
NAND2_X1 _u10_U6003  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17431 ) );
NAND2_X1 _u10_U6002  ( .A1(ch0_csr[15]), .A2(_u10_n12010 ), .ZN(_u10_n17432 ) );
NAND3_X1 _u10_U6001  ( .A1(_u10_n17430 ), .A2(_u10_n17431 ), .A3(_u10_n17432 ), .ZN(_u10_n17429 ) );
NOR4_X1 _u10_U6000  ( .A1(_u10_n17426 ), .A2(_u10_n17427 ), .A3(_u10_n17428 ), .A4(_u10_n17429 ), .ZN(_u10_n17404 ) );
NAND2_X1 _u10_U5999  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n17422 ) );
NAND2_X1 _u10_U5998  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n17423 ) );
NAND2_X1 _u10_U5997  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n17424 ) );
NAND2_X1 _u10_U5996  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n17425 ) );
NAND4_X1 _u10_U5995  ( .A1(_u10_n17422 ), .A2(_u10_n17423 ), .A3(_u10_n17424 ), .A4(_u10_n17425 ), .ZN(_u10_n17406 ) );
NAND2_X1 _u10_U5994  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n17418 ) );
NAND2_X1 _u10_U5993  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n17419 ) );
NAND2_X1 _u10_U5992  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n17420 ) );
NAND2_X1 _u10_U5991  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n17421 ) );
NAND4_X1 _u10_U5990  ( .A1(_u10_n17418 ), .A2(_u10_n17419 ), .A3(_u10_n17420 ), .A4(_u10_n17421 ), .ZN(_u10_n17407 ) );
NAND2_X1 _u10_U5989  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n17414 ) );
NAND2_X1 _u10_U5988  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n17415 ) );
NAND2_X1 _u10_U5987  ( .A1(1'b0), .A2(_u10_n11753 ), .ZN(_u10_n17416 ) );
NAND2_X1 _u10_U5986  ( .A1(1'b0), .A2(_u10_n11729 ), .ZN(_u10_n17417 ) );
NAND4_X1 _u10_U5985  ( .A1(_u10_n17414 ), .A2(_u10_n17415 ), .A3(_u10_n17416 ), .A4(_u10_n17417 ), .ZN(_u10_n17408 ) );
NAND2_X1 _u10_U5984  ( .A1(1'b0), .A2(_u10_n11705 ), .ZN(_u10_n17410 ) );
NAND2_X1 _u10_U5983  ( .A1(1'b0), .A2(_u10_n11681 ), .ZN(_u10_n17411 ) );
NAND2_X1 _u10_U5982  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n17412 ) );
NAND2_X1 _u10_U5981  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n17413 ) );
NAND4_X1 _u10_U5980  ( .A1(_u10_n17410 ), .A2(_u10_n17411 ), .A3(_u10_n17412 ), .A4(_u10_n17413 ), .ZN(_u10_n17409 ) );
NOR4_X1 _u10_U5979  ( .A1(_u10_n17406 ), .A2(_u10_n17407 ), .A3(_u10_n17408 ), .A4(_u10_n17409 ), .ZN(_u10_n17405 ) );
NAND2_X1 _u10_U5978  ( .A1(_u10_n17404 ), .A2(_u10_n17405 ), .ZN(csr[15]) );
NAND2_X1 _u10_U5977  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17400 ) );
NAND2_X1 _u10_U5976  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17401 ) );
NAND2_X1 _u10_U5975  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17402 ) );
NAND2_X1 _u10_U5974  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17403 ) );
NAND4_X1 _u10_U5973  ( .A1(_u10_n17400 ), .A2(_u10_n17401 ), .A3(_u10_n17402 ), .A4(_u10_n17403 ), .ZN(_u10_n17385 ) );
NAND2_X1 _u10_U5972  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17396 ) );
NAND2_X1 _u10_U5971  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17397 ) );
NAND2_X1 _u10_U5970  ( .A1(1'b0), .A2(_u10_n12209 ), .ZN(_u10_n17398 ) );
NAND2_X1 _u10_U5969  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17399 ) );
NAND4_X1 _u10_U5968  ( .A1(_u10_n17396 ), .A2(_u10_n17397 ), .A3(_u10_n17398 ), .A4(_u10_n17399 ), .ZN(_u10_n17386 ) );
NAND2_X1 _u10_U5967  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17392 ) );
NAND2_X1 _u10_U5966  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17393 ) );
NAND2_X1 _u10_U5965  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17394 ) );
NAND2_X1 _u10_U5964  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17395 ) );
NAND4_X1 _u10_U5963  ( .A1(_u10_n17392 ), .A2(_u10_n17393 ), .A3(_u10_n17394 ), .A4(_u10_n17395 ), .ZN(_u10_n17387 ) );
NAND2_X1 _u10_U5962  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17389 ) );
NAND2_X1 _u10_U5961  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17390 ) );
NAND2_X1 _u10_U5960  ( .A1(ch0_csr[16]), .A2(_u10_n12010 ), .ZN(_u10_n17391 ) );
NAND3_X1 _u10_U5959  ( .A1(_u10_n17389 ), .A2(_u10_n17390 ), .A3(_u10_n17391 ), .ZN(_u10_n17388 ) );
NOR4_X1 _u10_U5958  ( .A1(_u10_n17385 ), .A2(_u10_n17386 ), .A3(_u10_n17387 ), .A4(_u10_n17388 ), .ZN(_u10_n17363 ) );
NAND2_X1 _u10_U5957  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n17381 ) );
NAND2_X1 _u10_U5956  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n17382 ) );
NAND2_X1 _u10_U5955  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n17383 ) );
NAND2_X1 _u10_U5954  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n17384 ) );
NAND4_X1 _u10_U5953  ( .A1(_u10_n17381 ), .A2(_u10_n17382 ), .A3(_u10_n17383 ), .A4(_u10_n17384 ), .ZN(_u10_n17365 ) );
NAND2_X1 _u10_U5952  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n17377 ) );
NAND2_X1 _u10_U5951  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n17378 ) );
NAND2_X1 _u10_U5950  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n17379 ) );
NAND2_X1 _u10_U5949  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n17380 ) );
NAND4_X1 _u10_U5948  ( .A1(_u10_n17377 ), .A2(_u10_n17378 ), .A3(_u10_n17379 ), .A4(_u10_n17380 ), .ZN(_u10_n17366 ) );
NAND2_X1 _u10_U5947  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n17373 ) );
NAND2_X1 _u10_U5946  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n17374 ) );
NAND2_X1 _u10_U5945  ( .A1(1'b0), .A2(_u10_n11755 ), .ZN(_u10_n17375 ) );
NAND2_X1 _u10_U5944  ( .A1(1'b0), .A2(_u10_n11731 ), .ZN(_u10_n17376 ) );
NAND4_X1 _u10_U5943  ( .A1(_u10_n17373 ), .A2(_u10_n17374 ), .A3(_u10_n17375 ), .A4(_u10_n17376 ), .ZN(_u10_n17367 ) );
NAND2_X1 _u10_U5942  ( .A1(1'b0), .A2(_u10_n11707 ), .ZN(_u10_n17369 ) );
NAND2_X1 _u10_U5941  ( .A1(1'b0), .A2(_u10_n11683 ), .ZN(_u10_n17370 ) );
NAND2_X1 _u10_U5940  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n17371 ) );
NAND2_X1 _u10_U5939  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n17372 ) );
NAND4_X1 _u10_U5938  ( .A1(_u10_n17369 ), .A2(_u10_n17370 ), .A3(_u10_n17371 ), .A4(_u10_n17372 ), .ZN(_u10_n17368 ) );
NOR4_X1 _u10_U5937  ( .A1(_u10_n17365 ), .A2(_u10_n17366 ), .A3(_u10_n17367 ), .A4(_u10_n17368 ), .ZN(_u10_n17364 ) );
NAND2_X1 _u10_U5936  ( .A1(_u10_n17363 ), .A2(_u10_n17364 ), .ZN(csr[16]) );
NAND2_X1 _u10_U5935  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17359 ) );
NAND2_X1 _u10_U5934  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17360 ) );
NAND2_X1 _u10_U5933  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17361 ) );
NAND2_X1 _u10_U5932  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17362 ) );
NAND4_X1 _u10_U5931  ( .A1(_u10_n17359 ), .A2(_u10_n17360 ), .A3(_u10_n17361 ), .A4(_u10_n17362 ), .ZN(_u10_n17344 ) );
NAND2_X1 _u10_U5930  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17355 ) );
NAND2_X1 _u10_U5929  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17356 ) );
NAND2_X1 _u10_U5928  ( .A1(1'b0), .A2(_u10_n12211 ), .ZN(_u10_n17357 ) );
NAND2_X1 _u10_U5927  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17358 ) );
NAND4_X1 _u10_U5926  ( .A1(_u10_n17355 ), .A2(_u10_n17356 ), .A3(_u10_n17357 ), .A4(_u10_n17358 ), .ZN(_u10_n17345 ) );
NAND2_X1 _u10_U5925  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17351 ) );
NAND2_X1 _u10_U5924  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17352 ) );
NAND2_X1 _u10_U5923  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17353 ) );
NAND2_X1 _u10_U5922  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17354 ) );
NAND4_X1 _u10_U5921  ( .A1(_u10_n17351 ), .A2(_u10_n17352 ), .A3(_u10_n17353 ), .A4(_u10_n17354 ), .ZN(_u10_n17346 ) );
NAND2_X1 _u10_U5920  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17348 ) );
NAND2_X1 _u10_U5919  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17349 ) );
NAND2_X1 _u10_U5918  ( .A1(ch0_csr[17]), .A2(_u10_n12010 ), .ZN(_u10_n17350 ) );
NAND3_X1 _u10_U5917  ( .A1(_u10_n17348 ), .A2(_u10_n17349 ), .A3(_u10_n17350 ), .ZN(_u10_n17347 ) );
NOR4_X1 _u10_U5916  ( .A1(_u10_n17344 ), .A2(_u10_n17345 ), .A3(_u10_n17346 ), .A4(_u10_n17347 ), .ZN(_u10_n17322 ) );
NAND2_X1 _u10_U5915  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n17340 ) );
NAND2_X1 _u10_U5914  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n17341 ) );
NAND2_X1 _u10_U5913  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n17342 ) );
NAND2_X1 _u10_U5912  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n17343 ) );
NAND4_X1 _u10_U5911  ( .A1(_u10_n17340 ), .A2(_u10_n17341 ), .A3(_u10_n17342 ), .A4(_u10_n17343 ), .ZN(_u10_n17324 ) );
NAND2_X1 _u10_U5910  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n17336 ) );
NAND2_X1 _u10_U5909  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n17337 ) );
NAND2_X1 _u10_U5908  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n17338 ) );
NAND2_X1 _u10_U5907  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n17339 ) );
NAND4_X1 _u10_U5906  ( .A1(_u10_n17336 ), .A2(_u10_n17337 ), .A3(_u10_n17338 ), .A4(_u10_n17339 ), .ZN(_u10_n17325 ) );
NAND2_X1 _u10_U5905  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n17332 ) );
NAND2_X1 _u10_U5904  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n17333 ) );
NAND2_X1 _u10_U5903  ( .A1(1'b0), .A2(_u10_n11757 ), .ZN(_u10_n17334 ) );
NAND2_X1 _u10_U5902  ( .A1(1'b0), .A2(_u10_n11732 ), .ZN(_u10_n17335 ) );
NAND4_X1 _u10_U5901  ( .A1(_u10_n17332 ), .A2(_u10_n17333 ), .A3(_u10_n17334 ), .A4(_u10_n17335 ), .ZN(_u10_n17326 ) );
NAND2_X1 _u10_U5900  ( .A1(1'b0), .A2(_u10_n11709 ), .ZN(_u10_n17328 ) );
NAND2_X1 _u10_U5899  ( .A1(1'b0), .A2(_u10_n11684 ), .ZN(_u10_n17329 ) );
NAND2_X1 _u10_U5898  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n17330 ) );
NAND2_X1 _u10_U5897  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n17331 ) );
NAND4_X1 _u10_U5896  ( .A1(_u10_n17328 ), .A2(_u10_n17329 ), .A3(_u10_n17330 ), .A4(_u10_n17331 ), .ZN(_u10_n17327 ) );
NOR4_X1 _u10_U5895  ( .A1(_u10_n17324 ), .A2(_u10_n17325 ), .A3(_u10_n17326 ), .A4(_u10_n17327 ), .ZN(_u10_n17323 ) );
NAND2_X1 _u10_U5894  ( .A1(_u10_n17322 ), .A2(_u10_n17323 ), .ZN(csr[17]) );
NAND2_X1 _u10_U5893  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17318 ) );
NAND2_X1 _u10_U5892  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17319 ) );
NAND2_X1 _u10_U5891  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17320 ) );
NAND2_X1 _u10_U5890  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17321 ) );
NAND4_X1 _u10_U5889  ( .A1(_u10_n17318 ), .A2(_u10_n17319 ), .A3(_u10_n17320 ), .A4(_u10_n17321 ), .ZN(_u10_n17303 ) );
NAND2_X1 _u10_U5888  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17314 ) );
NAND2_X1 _u10_U5887  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17315 ) );
NAND2_X1 _u10_U5886  ( .A1(1'b0), .A2(_u10_n12210 ), .ZN(_u10_n17316 ) );
NAND2_X1 _u10_U5885  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17317 ) );
NAND4_X1 _u10_U5884  ( .A1(_u10_n17314 ), .A2(_u10_n17315 ), .A3(_u10_n17316 ), .A4(_u10_n17317 ), .ZN(_u10_n17304 ) );
NAND2_X1 _u10_U5883  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17310 ) );
NAND2_X1 _u10_U5882  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17311 ) );
NAND2_X1 _u10_U5881  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17312 ) );
NAND2_X1 _u10_U5880  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17313 ) );
NAND4_X1 _u10_U5879  ( .A1(_u10_n17310 ), .A2(_u10_n17311 ), .A3(_u10_n17312 ), .A4(_u10_n17313 ), .ZN(_u10_n17305 ) );
NAND2_X1 _u10_U5878  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17307 ) );
NAND2_X1 _u10_U5877  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17308 ) );
NAND2_X1 _u10_U5876  ( .A1(ch0_csr[18]), .A2(_u10_n12010 ), .ZN(_u10_n17309 ) );
NAND3_X1 _u10_U5875  ( .A1(_u10_n17307 ), .A2(_u10_n17308 ), .A3(_u10_n17309 ), .ZN(_u10_n17306 ) );
NOR4_X1 _u10_U5874  ( .A1(_u10_n17303 ), .A2(_u10_n17304 ), .A3(_u10_n17305 ), .A4(_u10_n17306 ), .ZN(_u10_n17281 ) );
NAND2_X1 _u10_U5873  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n17299 ) );
NAND2_X1 _u10_U5872  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n17300 ) );
NAND2_X1 _u10_U5871  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n17301 ) );
NAND2_X1 _u10_U5870  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n17302 ) );
NAND4_X1 _u10_U5869  ( .A1(_u10_n17299 ), .A2(_u10_n17300 ), .A3(_u10_n17301 ), .A4(_u10_n17302 ), .ZN(_u10_n17283 ) );
NAND2_X1 _u10_U5868  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n17295 ) );
NAND2_X1 _u10_U5867  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n17296 ) );
NAND2_X1 _u10_U5866  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n17297 ) );
NAND2_X1 _u10_U5865  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n17298 ) );
NAND4_X1 _u10_U5864  ( .A1(_u10_n17295 ), .A2(_u10_n17296 ), .A3(_u10_n17297 ), .A4(_u10_n17298 ), .ZN(_u10_n17284 ) );
NAND2_X1 _u10_U5863  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n17291 ) );
NAND2_X1 _u10_U5862  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n17292 ) );
NAND2_X1 _u10_U5861  ( .A1(1'b0), .A2(_u10_n11756 ), .ZN(_u10_n17293 ) );
NAND2_X1 _u10_U5860  ( .A1(1'b0), .A2(_u10_n11734 ), .ZN(_u10_n17294 ) );
NAND4_X1 _u10_U5859  ( .A1(_u10_n17291 ), .A2(_u10_n17292 ), .A3(_u10_n17293 ), .A4(_u10_n17294 ), .ZN(_u10_n17285 ) );
NAND2_X1 _u10_U5858  ( .A1(1'b0), .A2(_u10_n11708 ), .ZN(_u10_n17287 ) );
NAND2_X1 _u10_U5857  ( .A1(1'b0), .A2(_u10_n11686 ), .ZN(_u10_n17288 ) );
NAND2_X1 _u10_U5856  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n17289 ) );
NAND2_X1 _u10_U5855  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n17290 ) );
NAND4_X1 _u10_U5854  ( .A1(_u10_n17287 ), .A2(_u10_n17288 ), .A3(_u10_n17289 ), .A4(_u10_n17290 ), .ZN(_u10_n17286 ) );
NOR4_X1 _u10_U5853  ( .A1(_u10_n17283 ), .A2(_u10_n17284 ), .A3(_u10_n17285 ), .A4(_u10_n17286 ), .ZN(_u10_n17282 ) );
NAND2_X1 _u10_U5852  ( .A1(_u10_n17281 ), .A2(_u10_n17282 ), .ZN(csr[18]) );
NAND2_X1 _u10_U5851  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17277 ) );
NAND2_X1 _u10_U5850  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17278 ) );
NAND2_X1 _u10_U5849  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17279 ) );
NAND2_X1 _u10_U5848  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17280 ) );
NAND4_X1 _u10_U5847  ( .A1(_u10_n17277 ), .A2(_u10_n17278 ), .A3(_u10_n17279 ), .A4(_u10_n17280 ), .ZN(_u10_n17262 ) );
NAND2_X1 _u10_U5846  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17273 ) );
NAND2_X1 _u10_U5845  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17274 ) );
NAND2_X1 _u10_U5844  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n17275 ) );
NAND2_X1 _u10_U5843  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17276 ) );
NAND4_X1 _u10_U5842  ( .A1(_u10_n17273 ), .A2(_u10_n17274 ), .A3(_u10_n17275 ), .A4(_u10_n17276 ), .ZN(_u10_n17263 ) );
NAND2_X1 _u10_U5841  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17269 ) );
NAND2_X1 _u10_U5840  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17270 ) );
NAND2_X1 _u10_U5839  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17271 ) );
NAND2_X1 _u10_U5838  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17272 ) );
NAND4_X1 _u10_U5837  ( .A1(_u10_n17269 ), .A2(_u10_n17270 ), .A3(_u10_n17271 ), .A4(_u10_n17272 ), .ZN(_u10_n17264 ) );
NAND2_X1 _u10_U5836  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17266 ) );
NAND2_X1 _u10_U5835  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17267 ) );
NAND2_X1 _u10_U5834  ( .A1(ch0_csr[19]), .A2(_u10_n12010 ), .ZN(_u10_n17268 ) );
NAND3_X1 _u10_U5833  ( .A1(_u10_n17266 ), .A2(_u10_n17267 ), .A3(_u10_n17268 ), .ZN(_u10_n17265 ) );
NOR4_X1 _u10_U5832  ( .A1(_u10_n17262 ), .A2(_u10_n17263 ), .A3(_u10_n17264 ), .A4(_u10_n17265 ), .ZN(_u10_n17240 ) );
NAND2_X1 _u10_U5831  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n17258 ) );
NAND2_X1 _u10_U5830  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n17259 ) );
NAND2_X1 _u10_U5829  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n17260 ) );
NAND2_X1 _u10_U5828  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n17261 ) );
NAND4_X1 _u10_U5827  ( .A1(_u10_n17258 ), .A2(_u10_n17259 ), .A3(_u10_n17260 ), .A4(_u10_n17261 ), .ZN(_u10_n17242 ) );
NAND2_X1 _u10_U5826  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n17254 ) );
NAND2_X1 _u10_U5825  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n17255 ) );
NAND2_X1 _u10_U5824  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n17256 ) );
NAND2_X1 _u10_U5823  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n17257 ) );
NAND4_X1 _u10_U5822  ( .A1(_u10_n17254 ), .A2(_u10_n17255 ), .A3(_u10_n17256 ), .A4(_u10_n17257 ), .ZN(_u10_n17243 ) );
NAND2_X1 _u10_U5821  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n17250 ) );
NAND2_X1 _u10_U5820  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n17251 ) );
NAND2_X1 _u10_U5819  ( .A1(1'b0), .A2(_u10_n11759 ), .ZN(_u10_n17252 ) );
NAND2_X1 _u10_U5818  ( .A1(1'b0), .A2(_u10_n11735 ), .ZN(_u10_n17253 ) );
NAND4_X1 _u10_U5817  ( .A1(_u10_n17250 ), .A2(_u10_n17251 ), .A3(_u10_n17252 ), .A4(_u10_n17253 ), .ZN(_u10_n17244 ) );
NAND2_X1 _u10_U5816  ( .A1(1'b0), .A2(_u10_n11711 ), .ZN(_u10_n17246 ) );
NAND2_X1 _u10_U5815  ( .A1(1'b0), .A2(_u10_n11687 ), .ZN(_u10_n17247 ) );
NAND2_X1 _u10_U5814  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n17248 ) );
NAND2_X1 _u10_U5813  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n17249 ) );
NAND4_X1 _u10_U5812  ( .A1(_u10_n17246 ), .A2(_u10_n17247 ), .A3(_u10_n17248 ), .A4(_u10_n17249 ), .ZN(_u10_n17245 ) );
NOR4_X1 _u10_U5811  ( .A1(_u10_n17242 ), .A2(_u10_n17243 ), .A3(_u10_n17244 ), .A4(_u10_n17245 ), .ZN(_u10_n17241 ) );
NAND2_X1 _u10_U5810  ( .A1(_u10_n17240 ), .A2(_u10_n17241 ), .ZN(csr[19]) );
NAND2_X1 _u10_U5809  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17236 ) );
NAND2_X1 _u10_U5808  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17237 ) );
NAND2_X1 _u10_U5807  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17238 ) );
NAND2_X1 _u10_U5806  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17239 ) );
NAND4_X1 _u10_U5805  ( .A1(_u10_n17236 ), .A2(_u10_n17237 ), .A3(_u10_n17238 ), .A4(_u10_n17239 ), .ZN(_u10_n17221 ) );
NAND2_X1 _u10_U5804  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17232 ) );
NAND2_X1 _u10_U5803  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17233 ) );
NAND2_X1 _u10_U5802  ( .A1(1'b0), .A2(_u10_n12207 ), .ZN(_u10_n17234 ) );
NAND2_X1 _u10_U5801  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17235 ) );
NAND4_X1 _u10_U5800  ( .A1(_u10_n17232 ), .A2(_u10_n17233 ), .A3(_u10_n17234 ), .A4(_u10_n17235 ), .ZN(_u10_n17222 ) );
NAND2_X1 _u10_U5799  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17228 ) );
NAND2_X1 _u10_U5798  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17229 ) );
NAND2_X1 _u10_U5797  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17230 ) );
NAND2_X1 _u10_U5796  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17231 ) );
NAND4_X1 _u10_U5795  ( .A1(_u10_n17228 ), .A2(_u10_n17229 ), .A3(_u10_n17230 ), .A4(_u10_n17231 ), .ZN(_u10_n17223 ) );
NAND2_X1 _u10_U5794  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17225 ) );
NAND2_X1 _u10_U5793  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17226 ) );
NAND2_X1 _u10_U5792  ( .A1(ch0_csr[1]), .A2(_u10_n12010 ), .ZN(_u10_n17227 ));
NAND3_X1 _u10_U5791  ( .A1(_u10_n17225 ), .A2(_u10_n17226 ), .A3(_u10_n17227 ), .ZN(_u10_n17224 ) );
NOR4_X1 _u10_U5790  ( .A1(_u10_n17221 ), .A2(_u10_n17222 ), .A3(_u10_n17223 ), .A4(_u10_n17224 ), .ZN(_u10_n17199 ) );
NAND2_X1 _u10_U5789  ( .A1(1'b0), .A2(_u10_n11976 ), .ZN(_u10_n17217 ) );
NAND2_X1 _u10_U5788  ( .A1(1'b0), .A2(_u10_n11952 ), .ZN(_u10_n17218 ) );
NAND2_X1 _u10_U5787  ( .A1(1'b0), .A2(_u10_n11928 ), .ZN(_u10_n17219 ) );
NAND2_X1 _u10_U5786  ( .A1(1'b0), .A2(_u10_n11904 ), .ZN(_u10_n17220 ) );
NAND4_X1 _u10_U5785  ( .A1(_u10_n17217 ), .A2(_u10_n17218 ), .A3(_u10_n17219 ), .A4(_u10_n17220 ), .ZN(_u10_n17201 ) );
NAND2_X1 _u10_U5784  ( .A1(1'b0), .A2(_u10_n11880 ), .ZN(_u10_n17213 ) );
NAND2_X1 _u10_U5783  ( .A1(1'b0), .A2(_u10_n11856 ), .ZN(_u10_n17214 ) );
NAND2_X1 _u10_U5782  ( .A1(1'b0), .A2(_u10_n11832 ), .ZN(_u10_n17215 ) );
NAND2_X1 _u10_U5781  ( .A1(1'b0), .A2(_u10_n11808 ), .ZN(_u10_n17216 ) );
NAND4_X1 _u10_U5780  ( .A1(_u10_n17213 ), .A2(_u10_n17214 ), .A3(_u10_n17215 ), .A4(_u10_n17216 ), .ZN(_u10_n17202 ) );
NAND2_X1 _u10_U5779  ( .A1(1'b0), .A2(_u10_n11784 ), .ZN(_u10_n17209 ) );
NAND2_X1 _u10_U5778  ( .A1(1'b0), .A2(_u10_n11760 ), .ZN(_u10_n17210 ) );
NAND2_X1 _u10_U5777  ( .A1(1'b0), .A2(_u10_n11758 ), .ZN(_u10_n17211 ) );
NAND2_X1 _u10_U5776  ( .A1(1'b0), .A2(_u10_n11733 ), .ZN(_u10_n17212 ) );
NAND4_X1 _u10_U5775  ( .A1(_u10_n17209 ), .A2(_u10_n17210 ), .A3(_u10_n17211 ), .A4(_u10_n17212 ), .ZN(_u10_n17203 ) );
NAND2_X1 _u10_U5774  ( .A1(1'b0), .A2(_u10_n11710 ), .ZN(_u10_n17205 ) );
NAND2_X1 _u10_U5773  ( .A1(1'b0), .A2(_u10_n11685 ), .ZN(_u10_n17206 ) );
NAND2_X1 _u10_U5772  ( .A1(1'b0), .A2(_u10_n11640 ), .ZN(_u10_n17207 ) );
NAND2_X1 _u10_U5771  ( .A1(1'b0), .A2(_u10_n11616 ), .ZN(_u10_n17208 ) );
NAND4_X1 _u10_U5770  ( .A1(_u10_n17205 ), .A2(_u10_n17206 ), .A3(_u10_n17207 ), .A4(_u10_n17208 ), .ZN(_u10_n17204 ) );
NOR4_X1 _u10_U5769  ( .A1(_u10_n17201 ), .A2(_u10_n17202 ), .A3(_u10_n17203 ), .A4(_u10_n17204 ), .ZN(_u10_n17200 ) );
NAND2_X1 _u10_U5768  ( .A1(_u10_n17199 ), .A2(_u10_n17200 ), .ZN(csr[1]) );
NAND2_X1 _u10_U5767  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17195 ) );
NAND2_X1 _u10_U5766  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17196 ) );
NAND2_X1 _u10_U5765  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17197 ) );
NAND2_X1 _u10_U5764  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17198 ) );
NAND4_X1 _u10_U5763  ( .A1(_u10_n17195 ), .A2(_u10_n17196 ), .A3(_u10_n17197 ), .A4(_u10_n17198 ), .ZN(_u10_n17180 ) );
NAND2_X1 _u10_U5762  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17191 ) );
NAND2_X1 _u10_U5761  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17192 ) );
NAND2_X1 _u10_U5760  ( .A1(1'b0), .A2(_u10_n12420 ), .ZN(_u10_n17193 ) );
NAND2_X1 _u10_U5759  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17194 ) );
NAND4_X1 _u10_U5758  ( .A1(_u10_n17191 ), .A2(_u10_n17192 ), .A3(_u10_n17193 ), .A4(_u10_n17194 ), .ZN(_u10_n17181 ) );
NAND2_X1 _u10_U5757  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17187 ) );
NAND2_X1 _u10_U5756  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17188 ) );
NAND2_X1 _u10_U5755  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17189 ) );
NAND2_X1 _u10_U5754  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17190 ) );
NAND4_X1 _u10_U5753  ( .A1(_u10_n17187 ), .A2(_u10_n17188 ), .A3(_u10_n17189 ), .A4(_u10_n17190 ), .ZN(_u10_n17182 ) );
NAND2_X1 _u10_U5752  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17184 ) );
NAND2_X1 _u10_U5751  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17185 ) );
NAND2_X1 _u10_U5750  ( .A1(ch0_csr[20]), .A2(_u10_n12010 ), .ZN(_u10_n17186 ) );
NAND3_X1 _u10_U5749  ( .A1(_u10_n17184 ), .A2(_u10_n17185 ), .A3(_u10_n17186 ), .ZN(_u10_n17183 ) );
NOR4_X1 _u10_U5748  ( .A1(_u10_n17180 ), .A2(_u10_n17181 ), .A3(_u10_n17182 ), .A4(_u10_n17183 ), .ZN(_u10_n17158 ) );
NAND2_X1 _u10_U5747  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n17176 ) );
NAND2_X1 _u10_U5746  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n17177 ) );
NAND2_X1 _u10_U5745  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n17178 ) );
NAND2_X1 _u10_U5744  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n17179 ) );
NAND4_X1 _u10_U5743  ( .A1(_u10_n17176 ), .A2(_u10_n17177 ), .A3(_u10_n17178 ), .A4(_u10_n17179 ), .ZN(_u10_n17160 ) );
NAND2_X1 _u10_U5742  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n17172 ) );
NAND2_X1 _u10_U5741  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n17173 ) );
NAND2_X1 _u10_U5740  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n17174 ) );
NAND2_X1 _u10_U5739  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n17175 ) );
NAND4_X1 _u10_U5738  ( .A1(_u10_n17172 ), .A2(_u10_n17173 ), .A3(_u10_n17174 ), .A4(_u10_n17175 ), .ZN(_u10_n17161 ) );
NAND2_X1 _u10_U5737  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n17168 ) );
NAND2_X1 _u10_U5736  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n17169 ) );
NAND2_X1 _u10_U5735  ( .A1(1'b0), .A2(_u10_n12378 ), .ZN(_u10_n17170 ) );
NAND2_X1 _u10_U5734  ( .A1(1'b0), .A2(_u10_n12377 ), .ZN(_u10_n17171 ) );
NAND4_X1 _u10_U5733  ( .A1(_u10_n17168 ), .A2(_u10_n17169 ), .A3(_u10_n17170 ), .A4(_u10_n17171 ), .ZN(_u10_n17162 ) );
NAND2_X1 _u10_U5732  ( .A1(1'b0), .A2(_u10_n12372 ), .ZN(_u10_n17164 ) );
NAND2_X1 _u10_U5731  ( .A1(1'b0), .A2(_u10_n12371 ), .ZN(_u10_n17165 ) );
NAND2_X1 _u10_U5730  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n17166 ) );
NAND2_X1 _u10_U5729  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n17167 ) );
NAND4_X1 _u10_U5728  ( .A1(_u10_n17164 ), .A2(_u10_n17165 ), .A3(_u10_n17166 ), .A4(_u10_n17167 ), .ZN(_u10_n17163 ) );
NOR4_X1 _u10_U5727  ( .A1(_u10_n17160 ), .A2(_u10_n17161 ), .A3(_u10_n17162 ), .A4(_u10_n17163 ), .ZN(_u10_n17159 ) );
NAND2_X1 _u10_U5726  ( .A1(_u10_n17158 ), .A2(_u10_n17159 ), .ZN(csr[20]) );
NAND2_X1 _u10_U5725  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17154 ) );
NAND2_X1 _u10_U5724  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17155 ) );
NAND2_X1 _u10_U5723  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17156 ) );
NAND2_X1 _u10_U5722  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17157 ) );
NAND4_X1 _u10_U5721  ( .A1(_u10_n17154 ), .A2(_u10_n17155 ), .A3(_u10_n17156 ), .A4(_u10_n17157 ), .ZN(_u10_n17139 ) );
NAND2_X1 _u10_U5720  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17150 ) );
NAND2_X1 _u10_U5719  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17151 ) );
NAND2_X1 _u10_U5718  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n17152 ) );
NAND2_X1 _u10_U5717  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17153 ) );
NAND4_X1 _u10_U5716  ( .A1(_u10_n17150 ), .A2(_u10_n17151 ), .A3(_u10_n17152 ), .A4(_u10_n17153 ), .ZN(_u10_n17140 ) );
NAND2_X1 _u10_U5715  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17146 ) );
NAND2_X1 _u10_U5714  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17147 ) );
NAND2_X1 _u10_U5713  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17148 ) );
NAND2_X1 _u10_U5712  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17149 ) );
NAND4_X1 _u10_U5711  ( .A1(_u10_n17146 ), .A2(_u10_n17147 ), .A3(_u10_n17148 ), .A4(_u10_n17149 ), .ZN(_u10_n17141 ) );
NAND2_X1 _u10_U5710  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17143 ) );
NAND2_X1 _u10_U5709  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17144 ) );
NAND2_X1 _u10_U5708  ( .A1(ch0_csr[21]), .A2(_u10_n12010 ), .ZN(_u10_n17145 ) );
NAND3_X1 _u10_U5707  ( .A1(_u10_n17143 ), .A2(_u10_n17144 ), .A3(_u10_n17145 ), .ZN(_u10_n17142 ) );
NOR4_X1 _u10_U5706  ( .A1(_u10_n17139 ), .A2(_u10_n17140 ), .A3(_u10_n17141 ), .A4(_u10_n17142 ), .ZN(_u10_n17117 ) );
NAND2_X1 _u10_U5705  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n17135 ) );
NAND2_X1 _u10_U5704  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n17136 ) );
NAND2_X1 _u10_U5703  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n17137 ) );
NAND2_X1 _u10_U5702  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n17138 ) );
NAND4_X1 _u10_U5701  ( .A1(_u10_n17135 ), .A2(_u10_n17136 ), .A3(_u10_n17137 ), .A4(_u10_n17138 ), .ZN(_u10_n17119 ) );
NAND2_X1 _u10_U5700  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n17131 ) );
NAND2_X1 _u10_U5699  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n17132 ) );
NAND2_X1 _u10_U5698  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n17133 ) );
NAND2_X1 _u10_U5697  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n17134 ) );
NAND4_X1 _u10_U5696  ( .A1(_u10_n17131 ), .A2(_u10_n17132 ), .A3(_u10_n17133 ), .A4(_u10_n17134 ), .ZN(_u10_n17120 ) );
NAND2_X1 _u10_U5695  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n17127 ) );
NAND2_X1 _u10_U5694  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n17128 ) );
NAND2_X1 _u10_U5693  ( .A1(1'b0), .A2(_u10_n11757 ), .ZN(_u10_n17129 ) );
NAND2_X1 _u10_U5692  ( .A1(1'b0), .A2(_u10_n11733 ), .ZN(_u10_n17130 ) );
NAND4_X1 _u10_U5691  ( .A1(_u10_n17127 ), .A2(_u10_n17128 ), .A3(_u10_n17129 ), .A4(_u10_n17130 ), .ZN(_u10_n17121 ) );
NAND2_X1 _u10_U5690  ( .A1(1'b0), .A2(_u10_n11709 ), .ZN(_u10_n17123 ) );
NAND2_X1 _u10_U5689  ( .A1(1'b0), .A2(_u10_n11685 ), .ZN(_u10_n17124 ) );
NAND2_X1 _u10_U5688  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n17125 ) );
NAND2_X1 _u10_U5687  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n17126 ) );
NAND4_X1 _u10_U5686  ( .A1(_u10_n17123 ), .A2(_u10_n17124 ), .A3(_u10_n17125 ), .A4(_u10_n17126 ), .ZN(_u10_n17122 ) );
NOR4_X1 _u10_U5685  ( .A1(_u10_n17119 ), .A2(_u10_n17120 ), .A3(_u10_n17121 ), .A4(_u10_n17122 ), .ZN(_u10_n17118 ) );
NAND2_X1 _u10_U5684  ( .A1(_u10_n17117 ), .A2(_u10_n17118 ), .ZN(csr[21]) );
NAND2_X1 _u10_U5683  ( .A1(1'b0), .A2(_u10_n12341 ), .ZN(_u10_n17113 ) );
NAND2_X1 _u10_U5682  ( .A1(1'b0), .A2(_u10_n12317 ), .ZN(_u10_n17114 ) );
NAND2_X1 _u10_U5681  ( .A1(1'b0), .A2(_u10_n12294 ), .ZN(_u10_n17115 ) );
NAND2_X1 _u10_U5680  ( .A1(1'b0), .A2(_u10_n12270 ), .ZN(_u10_n17116 ) );
NAND4_X1 _u10_U5679  ( .A1(_u10_n17113 ), .A2(_u10_n17114 ), .A3(_u10_n17115 ), .A4(_u10_n17116 ), .ZN(_u10_n17098 ) );
NAND2_X1 _u10_U5678  ( .A1(1'b0), .A2(_u10_n12245 ), .ZN(_u10_n17109 ) );
NAND2_X1 _u10_U5677  ( .A1(1'b0), .A2(_u10_n12221 ), .ZN(_u10_n17110 ) );
NAND2_X1 _u10_U5676  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n17111 ) );
NAND2_X1 _u10_U5675  ( .A1(1'b0), .A2(_u10_n12173 ), .ZN(_u10_n17112 ) );
NAND4_X1 _u10_U5674  ( .A1(_u10_n17109 ), .A2(_u10_n17110 ), .A3(_u10_n17111 ), .A4(_u10_n17112 ), .ZN(_u10_n17099 ) );
NAND2_X1 _u10_U5673  ( .A1(1'b0), .A2(_u10_n12150 ), .ZN(_u10_n17105 ) );
NAND2_X1 _u10_U5672  ( .A1(1'b0), .A2(_u10_n12126 ), .ZN(_u10_n17106 ) );
NAND2_X1 _u10_U5671  ( .A1(1'b0), .A2(_u10_n12102 ), .ZN(_u10_n17107 ) );
NAND2_X1 _u10_U5670  ( .A1(1'b0), .A2(_u10_n12078 ), .ZN(_u10_n17108 ) );
NAND4_X1 _u10_U5669  ( .A1(_u10_n17105 ), .A2(_u10_n17106 ), .A3(_u10_n17107 ), .A4(_u10_n17108 ), .ZN(_u10_n17100 ) );
NAND2_X1 _u10_U5668  ( .A1(1'b0), .A2(_u10_n12054 ), .ZN(_u10_n17102 ) );
NAND2_X1 _u10_U5667  ( .A1(1'b0), .A2(_u10_n12030 ), .ZN(_u10_n17103 ) );
NAND2_X1 _u10_U5666  ( .A1(ch0_csr[22]), .A2(_u10_n12010 ), .ZN(_u10_n17104 ) );
NAND3_X1 _u10_U5665  ( .A1(_u10_n17102 ), .A2(_u10_n17103 ), .A3(_u10_n17104 ), .ZN(_u10_n17101 ) );
NOR4_X1 _u10_U5664  ( .A1(_u10_n17098 ), .A2(_u10_n17099 ), .A3(_u10_n17100 ), .A4(_u10_n17101 ), .ZN(_u10_n17076 ) );
NAND2_X1 _u10_U5663  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n17094 ) );
NAND2_X1 _u10_U5662  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n17095 ) );
NAND2_X1 _u10_U5661  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n17096 ) );
NAND2_X1 _u10_U5660  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n17097 ) );
NAND4_X1 _u10_U5659  ( .A1(_u10_n17094 ), .A2(_u10_n17095 ), .A3(_u10_n17096 ), .A4(_u10_n17097 ), .ZN(_u10_n17078 ) );
NAND2_X1 _u10_U5658  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n17090 ) );
NAND2_X1 _u10_U5657  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n17091 ) );
NAND2_X1 _u10_U5656  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n17092 ) );
NAND2_X1 _u10_U5655  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n17093 ) );
NAND4_X1 _u10_U5654  ( .A1(_u10_n17090 ), .A2(_u10_n17091 ), .A3(_u10_n17092 ), .A4(_u10_n17093 ), .ZN(_u10_n17079 ) );
NAND2_X1 _u10_U5653  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n17086 ) );
NAND2_X1 _u10_U5652  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n17087 ) );
NAND2_X1 _u10_U5651  ( .A1(1'b0), .A2(_u10_n11756 ), .ZN(_u10_n17088 ) );
NAND2_X1 _u10_U5650  ( .A1(1'b0), .A2(_u10_n11732 ), .ZN(_u10_n17089 ) );
NAND4_X1 _u10_U5649  ( .A1(_u10_n17086 ), .A2(_u10_n17087 ), .A3(_u10_n17088 ), .A4(_u10_n17089 ), .ZN(_u10_n17080 ) );
NAND2_X1 _u10_U5648  ( .A1(1'b0), .A2(_u10_n11708 ), .ZN(_u10_n17082 ) );
NAND2_X1 _u10_U5647  ( .A1(1'b0), .A2(_u10_n11684 ), .ZN(_u10_n17083 ) );
NAND2_X1 _u10_U5646  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n17084 ) );
NAND2_X1 _u10_U5645  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n17085 ) );
NAND4_X1 _u10_U5644  ( .A1(_u10_n17082 ), .A2(_u10_n17083 ), .A3(_u10_n17084 ), .A4(_u10_n17085 ), .ZN(_u10_n17081 ) );
NOR4_X1 _u10_U5643  ( .A1(_u10_n17078 ), .A2(_u10_n17079 ), .A3(_u10_n17080 ), .A4(_u10_n17081 ), .ZN(_u10_n17077 ) );
NAND2_X1 _u10_U5642  ( .A1(_u10_n17076 ), .A2(_u10_n17077 ), .ZN(csr[22]) );
NAND2_X1 _u10_U5641  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n17072 ) );
NAND2_X1 _u10_U5640  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n17073 ) );
NAND2_X1 _u10_U5639  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n17074 ) );
NAND2_X1 _u10_U5638  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n17075 ) );
NAND4_X1 _u10_U5637  ( .A1(_u10_n17072 ), .A2(_u10_n17073 ), .A3(_u10_n17074 ), .A4(_u10_n17075 ), .ZN(_u10_n17057 ) );
NAND2_X1 _u10_U5636  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n17068 ) );
NAND2_X1 _u10_U5635  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n17069 ) );
NAND2_X1 _u10_U5634  ( .A1(1'b0), .A2(_u10_n12209 ), .ZN(_u10_n17070 ) );
NAND2_X1 _u10_U5633  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n17071 ) );
NAND4_X1 _u10_U5632  ( .A1(_u10_n17068 ), .A2(_u10_n17069 ), .A3(_u10_n17070 ), .A4(_u10_n17071 ), .ZN(_u10_n17058 ) );
NAND2_X1 _u10_U5631  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n17064 ) );
NAND2_X1 _u10_U5630  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n17065 ) );
NAND2_X1 _u10_U5629  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n17066 ) );
NAND2_X1 _u10_U5628  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n17067 ) );
NAND4_X1 _u10_U5627  ( .A1(_u10_n17064 ), .A2(_u10_n17065 ), .A3(_u10_n17066 ), .A4(_u10_n17067 ), .ZN(_u10_n17059 ) );
NAND2_X1 _u10_U5626  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n17061 ) );
NAND2_X1 _u10_U5625  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n17062 ) );
NAND2_X1 _u10_U5624  ( .A1(1'b0), .A2(_u10_n12011 ), .ZN(_u10_n17063 ) );
NAND3_X1 _u10_U5623  ( .A1(_u10_n17061 ), .A2(_u10_n17062 ), .A3(_u10_n17063 ), .ZN(_u10_n17060 ) );
NOR4_X1 _u10_U5622  ( .A1(_u10_n17057 ), .A2(_u10_n17058 ), .A3(_u10_n17059 ), .A4(_u10_n17060 ), .ZN(_u10_n17035 ) );
NAND2_X1 _u10_U5621  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n17053 ) );
NAND2_X1 _u10_U5620  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n17054 ) );
NAND2_X1 _u10_U5619  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n17055 ) );
NAND2_X1 _u10_U5618  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n17056 ) );
NAND4_X1 _u10_U5617  ( .A1(_u10_n17053 ), .A2(_u10_n17054 ), .A3(_u10_n17055 ), .A4(_u10_n17056 ), .ZN(_u10_n17037 ) );
NAND2_X1 _u10_U5616  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n17049 ) );
NAND2_X1 _u10_U5615  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n17050 ) );
NAND2_X1 _u10_U5614  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n17051 ) );
NAND2_X1 _u10_U5613  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n17052 ) );
NAND4_X1 _u10_U5612  ( .A1(_u10_n17049 ), .A2(_u10_n17050 ), .A3(_u10_n17051 ), .A4(_u10_n17052 ), .ZN(_u10_n17038 ) );
NAND2_X1 _u10_U5611  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n17045 ) );
NAND2_X1 _u10_U5610  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n17046 ) );
NAND2_X1 _u10_U5609  ( .A1(1'b0), .A2(_u10_n11753 ), .ZN(_u10_n17047 ) );
NAND2_X1 _u10_U5608  ( .A1(1'b0), .A2(_u10_n11729 ), .ZN(_u10_n17048 ) );
NAND4_X1 _u10_U5607  ( .A1(_u10_n17045 ), .A2(_u10_n17046 ), .A3(_u10_n17047 ), .A4(_u10_n17048 ), .ZN(_u10_n17039 ) );
NAND2_X1 _u10_U5606  ( .A1(1'b0), .A2(_u10_n11705 ), .ZN(_u10_n17041 ) );
NAND2_X1 _u10_U5605  ( .A1(1'b0), .A2(_u10_n11681 ), .ZN(_u10_n17042 ) );
NAND2_X1 _u10_U5604  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n17043 ) );
NAND2_X1 _u10_U5603  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n17044 ) );
NAND4_X1 _u10_U5602  ( .A1(_u10_n17041 ), .A2(_u10_n17042 ), .A3(_u10_n17043 ), .A4(_u10_n17044 ), .ZN(_u10_n17040 ) );
NOR4_X1 _u10_U5601  ( .A1(_u10_n17037 ), .A2(_u10_n17038 ), .A3(_u10_n17039 ), .A4(_u10_n17040 ), .ZN(_u10_n17036 ) );
NAND2_X1 _u10_U5600  ( .A1(_u10_n17035 ), .A2(_u10_n17036 ), .ZN(csr[23]) );
NAND2_X1 _u10_U5599  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n17031 ) );
NAND2_X1 _u10_U5598  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n17032 ) );
NAND2_X1 _u10_U5597  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n17033 ) );
NAND2_X1 _u10_U5596  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n17034 ) );
NAND4_X1 _u10_U5595  ( .A1(_u10_n17031 ), .A2(_u10_n17032 ), .A3(_u10_n17033 ), .A4(_u10_n17034 ), .ZN(_u10_n17016 ) );
NAND2_X1 _u10_U5594  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n17027 ) );
NAND2_X1 _u10_U5593  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n17028 ) );
NAND2_X1 _u10_U5592  ( .A1(1'b0), .A2(_u10_n12211 ), .ZN(_u10_n17029 ) );
NAND2_X1 _u10_U5591  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n17030 ) );
NAND4_X1 _u10_U5590  ( .A1(_u10_n17027 ), .A2(_u10_n17028 ), .A3(_u10_n17029 ), .A4(_u10_n17030 ), .ZN(_u10_n17017 ) );
NAND2_X1 _u10_U5589  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n17023 ) );
NAND2_X1 _u10_U5588  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n17024 ) );
NAND2_X1 _u10_U5587  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n17025 ) );
NAND2_X1 _u10_U5586  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n17026 ) );
NAND4_X1 _u10_U5585  ( .A1(_u10_n17023 ), .A2(_u10_n17024 ), .A3(_u10_n17025 ), .A4(_u10_n17026 ), .ZN(_u10_n17018 ) );
NAND2_X1 _u10_U5584  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n17020 ) );
NAND2_X1 _u10_U5583  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n17021 ) );
NAND2_X1 _u10_U5582  ( .A1(1'b0), .A2(_u10_n12011 ), .ZN(_u10_n17022 ) );
NAND3_X1 _u10_U5581  ( .A1(_u10_n17020 ), .A2(_u10_n17021 ), .A3(_u10_n17022 ), .ZN(_u10_n17019 ) );
NOR4_X1 _u10_U5580  ( .A1(_u10_n17016 ), .A2(_u10_n17017 ), .A3(_u10_n17018 ), .A4(_u10_n17019 ), .ZN(_u10_n16994 ) );
NAND2_X1 _u10_U5579  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n17012 ) );
NAND2_X1 _u10_U5578  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n17013 ) );
NAND2_X1 _u10_U5577  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n17014 ) );
NAND2_X1 _u10_U5576  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n17015 ) );
NAND4_X1 _u10_U5575  ( .A1(_u10_n17012 ), .A2(_u10_n17013 ), .A3(_u10_n17014 ), .A4(_u10_n17015 ), .ZN(_u10_n16996 ) );
NAND2_X1 _u10_U5574  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n17008 ) );
NAND2_X1 _u10_U5573  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n17009 ) );
NAND2_X1 _u10_U5572  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n17010 ) );
NAND2_X1 _u10_U5571  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n17011 ) );
NAND4_X1 _u10_U5570  ( .A1(_u10_n17008 ), .A2(_u10_n17009 ), .A3(_u10_n17010 ), .A4(_u10_n17011 ), .ZN(_u10_n16997 ) );
NAND2_X1 _u10_U5569  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n17004 ) );
NAND2_X1 _u10_U5568  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n17005 ) );
NAND2_X1 _u10_U5567  ( .A1(1'b0), .A2(_u10_n11758 ), .ZN(_u10_n17006 ) );
NAND2_X1 _u10_U5566  ( .A1(1'b0), .A2(_u10_n11734 ), .ZN(_u10_n17007 ) );
NAND4_X1 _u10_U5565  ( .A1(_u10_n17004 ), .A2(_u10_n17005 ), .A3(_u10_n17006 ), .A4(_u10_n17007 ), .ZN(_u10_n16998 ) );
NAND2_X1 _u10_U5564  ( .A1(1'b0), .A2(_u10_n11710 ), .ZN(_u10_n17000 ) );
NAND2_X1 _u10_U5563  ( .A1(1'b0), .A2(_u10_n11686 ), .ZN(_u10_n17001 ) );
NAND2_X1 _u10_U5562  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n17002 ) );
NAND2_X1 _u10_U5561  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n17003 ) );
NAND4_X1 _u10_U5560  ( .A1(_u10_n17000 ), .A2(_u10_n17001 ), .A3(_u10_n17002 ), .A4(_u10_n17003 ), .ZN(_u10_n16999 ) );
NOR4_X1 _u10_U5559  ( .A1(_u10_n16996 ), .A2(_u10_n16997 ), .A3(_u10_n16998 ), .A4(_u10_n16999 ), .ZN(_u10_n16995 ) );
NAND2_X1 _u10_U5558  ( .A1(_u10_n16994 ), .A2(_u10_n16995 ), .ZN(csr[24]) );
NAND2_X1 _u10_U5557  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n16990 ) );
NAND2_X1 _u10_U5556  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n16991 ) );
NAND2_X1 _u10_U5555  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n16992 ) );
NAND2_X1 _u10_U5554  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n16993 ) );
NAND4_X1 _u10_U5553  ( .A1(_u10_n16990 ), .A2(_u10_n16991 ), .A3(_u10_n16992 ), .A4(_u10_n16993 ), .ZN(_u10_n16975 ) );
NAND2_X1 _u10_U5552  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n16986 ) );
NAND2_X1 _u10_U5551  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n16987 ) );
NAND2_X1 _u10_U5550  ( .A1(1'b0), .A2(_u10_n12210 ), .ZN(_u10_n16988 ) );
NAND2_X1 _u10_U5549  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n16989 ) );
NAND4_X1 _u10_U5548  ( .A1(_u10_n16986 ), .A2(_u10_n16987 ), .A3(_u10_n16988 ), .A4(_u10_n16989 ), .ZN(_u10_n16976 ) );
NAND2_X1 _u10_U5547  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n16982 ) );
NAND2_X1 _u10_U5546  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n16983 ) );
NAND2_X1 _u10_U5545  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n16984 ) );
NAND2_X1 _u10_U5544  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n16985 ) );
NAND4_X1 _u10_U5543  ( .A1(_u10_n16982 ), .A2(_u10_n16983 ), .A3(_u10_n16984 ), .A4(_u10_n16985 ), .ZN(_u10_n16977 ) );
NAND2_X1 _u10_U5542  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n16979 ) );
NAND2_X1 _u10_U5541  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n16980 ) );
NAND2_X1 _u10_U5540  ( .A1(1'b0), .A2(_u10_n12011 ), .ZN(_u10_n16981 ) );
NAND3_X1 _u10_U5539  ( .A1(_u10_n16979 ), .A2(_u10_n16980 ), .A3(_u10_n16981 ), .ZN(_u10_n16978 ) );
NOR4_X1 _u10_U5538  ( .A1(_u10_n16975 ), .A2(_u10_n16976 ), .A3(_u10_n16977 ), .A4(_u10_n16978 ), .ZN(_u10_n16953 ) );
NAND2_X1 _u10_U5537  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n16971 ) );
NAND2_X1 _u10_U5536  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n16972 ) );
NAND2_X1 _u10_U5535  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n16973 ) );
NAND2_X1 _u10_U5534  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n16974 ) );
NAND4_X1 _u10_U5533  ( .A1(_u10_n16971 ), .A2(_u10_n16972 ), .A3(_u10_n16973 ), .A4(_u10_n16974 ), .ZN(_u10_n16955 ) );
NAND2_X1 _u10_U5532  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n16967 ) );
NAND2_X1 _u10_U5531  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n16968 ) );
NAND2_X1 _u10_U5530  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n16969 ) );
NAND2_X1 _u10_U5529  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n16970 ) );
NAND4_X1 _u10_U5528  ( .A1(_u10_n16967 ), .A2(_u10_n16968 ), .A3(_u10_n16969 ), .A4(_u10_n16970 ), .ZN(_u10_n16956 ) );
NAND2_X1 _u10_U5527  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n16963 ) );
NAND2_X1 _u10_U5526  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n16964 ) );
NAND2_X1 _u10_U5525  ( .A1(1'b0), .A2(_u10_n11757 ), .ZN(_u10_n16965 ) );
NAND2_X1 _u10_U5524  ( .A1(1'b0), .A2(_u10_n11733 ), .ZN(_u10_n16966 ) );
NAND4_X1 _u10_U5523  ( .A1(_u10_n16963 ), .A2(_u10_n16964 ), .A3(_u10_n16965 ), .A4(_u10_n16966 ), .ZN(_u10_n16957 ) );
NAND2_X1 _u10_U5522  ( .A1(1'b0), .A2(_u10_n11709 ), .ZN(_u10_n16959 ) );
NAND2_X1 _u10_U5521  ( .A1(1'b0), .A2(_u10_n11685 ), .ZN(_u10_n16960 ) );
NAND2_X1 _u10_U5520  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n16961 ) );
NAND2_X1 _u10_U5519  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n16962 ) );
NAND4_X1 _u10_U5518  ( .A1(_u10_n16959 ), .A2(_u10_n16960 ), .A3(_u10_n16961 ), .A4(_u10_n16962 ), .ZN(_u10_n16958 ) );
NOR4_X1 _u10_U5517  ( .A1(_u10_n16955 ), .A2(_u10_n16956 ), .A3(_u10_n16957 ), .A4(_u10_n16958 ), .ZN(_u10_n16954 ) );
NAND2_X1 _u10_U5516  ( .A1(_u10_n16953 ), .A2(_u10_n16954 ), .ZN(csr[25]) );
NAND2_X1 _u10_U5515  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n16949 ) );
NAND2_X1 _u10_U5514  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n16950 ) );
NAND2_X1 _u10_U5513  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n16951 ) );
NAND2_X1 _u10_U5512  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n16952 ) );
NAND4_X1 _u10_U5511  ( .A1(_u10_n16949 ), .A2(_u10_n16950 ), .A3(_u10_n16951 ), .A4(_u10_n16952 ), .ZN(_u10_n16934 ) );
NAND2_X1 _u10_U5510  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n16945 ) );
NAND2_X1 _u10_U5509  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n16946 ) );
NAND2_X1 _u10_U5508  ( .A1(1'b0), .A2(_u10_n12207 ), .ZN(_u10_n16947 ) );
NAND2_X1 _u10_U5507  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n16948 ) );
NAND4_X1 _u10_U5506  ( .A1(_u10_n16945 ), .A2(_u10_n16946 ), .A3(_u10_n16947 ), .A4(_u10_n16948 ), .ZN(_u10_n16935 ) );
NAND2_X1 _u10_U5505  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n16941 ) );
NAND2_X1 _u10_U5504  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n16942 ) );
NAND2_X1 _u10_U5503  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n16943 ) );
NAND2_X1 _u10_U5502  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n16944 ) );
NAND4_X1 _u10_U5501  ( .A1(_u10_n16941 ), .A2(_u10_n16942 ), .A3(_u10_n16943 ), .A4(_u10_n16944 ), .ZN(_u10_n16936 ) );
NAND2_X1 _u10_U5500  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n16938 ) );
NAND2_X1 _u10_U5499  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n16939 ) );
NAND2_X1 _u10_U5498  ( .A1(1'b0), .A2(_u10_n12011 ), .ZN(_u10_n16940 ) );
NAND3_X1 _u10_U5497  ( .A1(_u10_n16938 ), .A2(_u10_n16939 ), .A3(_u10_n16940 ), .ZN(_u10_n16937 ) );
NOR4_X1 _u10_U5496  ( .A1(_u10_n16934 ), .A2(_u10_n16935 ), .A3(_u10_n16936 ), .A4(_u10_n16937 ), .ZN(_u10_n16912 ) );
NAND2_X1 _u10_U5495  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n16930 ) );
NAND2_X1 _u10_U5494  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n16931 ) );
NAND2_X1 _u10_U5493  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n16932 ) );
NAND2_X1 _u10_U5492  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n16933 ) );
NAND4_X1 _u10_U5491  ( .A1(_u10_n16930 ), .A2(_u10_n16931 ), .A3(_u10_n16932 ), .A4(_u10_n16933 ), .ZN(_u10_n16914 ) );
NAND2_X1 _u10_U5490  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n16926 ) );
NAND2_X1 _u10_U5489  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n16927 ) );
NAND2_X1 _u10_U5488  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n16928 ) );
NAND2_X1 _u10_U5487  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n16929 ) );
NAND4_X1 _u10_U5486  ( .A1(_u10_n16926 ), .A2(_u10_n16927 ), .A3(_u10_n16928 ), .A4(_u10_n16929 ), .ZN(_u10_n16915 ) );
NAND2_X1 _u10_U5485  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n16922 ) );
NAND2_X1 _u10_U5484  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n16923 ) );
NAND2_X1 _u10_U5483  ( .A1(1'b0), .A2(_u10_n11755 ), .ZN(_u10_n16924 ) );
NAND2_X1 _u10_U5482  ( .A1(1'b0), .A2(_u10_n11731 ), .ZN(_u10_n16925 ) );
NAND4_X1 _u10_U5481  ( .A1(_u10_n16922 ), .A2(_u10_n16923 ), .A3(_u10_n16924 ), .A4(_u10_n16925 ), .ZN(_u10_n16916 ) );
NAND2_X1 _u10_U5480  ( .A1(1'b0), .A2(_u10_n11707 ), .ZN(_u10_n16918 ) );
NAND2_X1 _u10_U5479  ( .A1(1'b0), .A2(_u10_n11683 ), .ZN(_u10_n16919 ) );
NAND2_X1 _u10_U5478  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n16920 ) );
NAND2_X1 _u10_U5477  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n16921 ) );
NAND4_X1 _u10_U5476  ( .A1(_u10_n16918 ), .A2(_u10_n16919 ), .A3(_u10_n16920 ), .A4(_u10_n16921 ), .ZN(_u10_n16917 ) );
NOR4_X1 _u10_U5475  ( .A1(_u10_n16914 ), .A2(_u10_n16915 ), .A3(_u10_n16916 ), .A4(_u10_n16917 ), .ZN(_u10_n16913 ) );
NAND2_X1 _u10_U5474  ( .A1(_u10_n16912 ), .A2(_u10_n16913 ), .ZN(csr[26]) );
NAND2_X1 _u10_U5473  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n16908 ) );
NAND2_X1 _u10_U5472  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n16909 ) );
NAND2_X1 _u10_U5471  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n16910 ) );
NAND2_X1 _u10_U5470  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n16911 ) );
NAND4_X1 _u10_U5469  ( .A1(_u10_n16908 ), .A2(_u10_n16909 ), .A3(_u10_n16910 ), .A4(_u10_n16911 ), .ZN(_u10_n16893 ) );
NAND2_X1 _u10_U5468  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n16904 ) );
NAND2_X1 _u10_U5467  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n16905 ) );
NAND2_X1 _u10_U5466  ( .A1(1'b0), .A2(_u10_n12420 ), .ZN(_u10_n16906 ) );
NAND2_X1 _u10_U5465  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n16907 ) );
NAND4_X1 _u10_U5464  ( .A1(_u10_n16904 ), .A2(_u10_n16905 ), .A3(_u10_n16906 ), .A4(_u10_n16907 ), .ZN(_u10_n16894 ) );
NAND2_X1 _u10_U5463  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n16900 ) );
NAND2_X1 _u10_U5462  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n16901 ) );
NAND2_X1 _u10_U5461  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n16902 ) );
NAND2_X1 _u10_U5460  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n16903 ) );
NAND4_X1 _u10_U5459  ( .A1(_u10_n16900 ), .A2(_u10_n16901 ), .A3(_u10_n16902 ), .A4(_u10_n16903 ), .ZN(_u10_n16895 ) );
NAND2_X1 _u10_U5458  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n16897 ) );
NAND2_X1 _u10_U5457  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n16898 ) );
NAND2_X1 _u10_U5456  ( .A1(1'b0), .A2(_u10_n12011 ), .ZN(_u10_n16899 ) );
NAND3_X1 _u10_U5455  ( .A1(_u10_n16897 ), .A2(_u10_n16898 ), .A3(_u10_n16899 ), .ZN(_u10_n16896 ) );
NOR4_X1 _u10_U5454  ( .A1(_u10_n16893 ), .A2(_u10_n16894 ), .A3(_u10_n16895 ), .A4(_u10_n16896 ), .ZN(_u10_n16871 ) );
NAND2_X1 _u10_U5453  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n16889 ) );
NAND2_X1 _u10_U5452  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n16890 ) );
NAND2_X1 _u10_U5451  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n16891 ) );
NAND2_X1 _u10_U5450  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n16892 ) );
NAND4_X1 _u10_U5449  ( .A1(_u10_n16889 ), .A2(_u10_n16890 ), .A3(_u10_n16891 ), .A4(_u10_n16892 ), .ZN(_u10_n16873 ) );
NAND2_X1 _u10_U5448  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n16885 ) );
NAND2_X1 _u10_U5447  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n16886 ) );
NAND2_X1 _u10_U5446  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n16887 ) );
NAND2_X1 _u10_U5445  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n16888 ) );
NAND4_X1 _u10_U5444  ( .A1(_u10_n16885 ), .A2(_u10_n16886 ), .A3(_u10_n16887 ), .A4(_u10_n16888 ), .ZN(_u10_n16874 ) );
NAND2_X1 _u10_U5443  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n16881 ) );
NAND2_X1 _u10_U5442  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n16882 ) );
NAND2_X1 _u10_U5441  ( .A1(1'b0), .A2(_u10_n11754 ), .ZN(_u10_n16883 ) );
NAND2_X1 _u10_U5440  ( .A1(1'b0), .A2(_u10_n11730 ), .ZN(_u10_n16884 ) );
NAND4_X1 _u10_U5439  ( .A1(_u10_n16881 ), .A2(_u10_n16882 ), .A3(_u10_n16883 ), .A4(_u10_n16884 ), .ZN(_u10_n16875 ) );
NAND2_X1 _u10_U5438  ( .A1(1'b0), .A2(_u10_n11706 ), .ZN(_u10_n16877 ) );
NAND2_X1 _u10_U5437  ( .A1(1'b0), .A2(_u10_n11682 ), .ZN(_u10_n16878 ) );
NAND2_X1 _u10_U5436  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n16879 ) );
NAND2_X1 _u10_U5435  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n16880 ) );
NAND4_X1 _u10_U5434  ( .A1(_u10_n16877 ), .A2(_u10_n16878 ), .A3(_u10_n16879 ), .A4(_u10_n16880 ), .ZN(_u10_n16876 ) );
NOR4_X1 _u10_U5433  ( .A1(_u10_n16873 ), .A2(_u10_n16874 ), .A3(_u10_n16875 ), .A4(_u10_n16876 ), .ZN(_u10_n16872 ) );
NAND2_X1 _u10_U5432  ( .A1(_u10_n16871 ), .A2(_u10_n16872 ), .ZN(csr[27]) );
NAND2_X1 _u10_U5431  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n16867 ) );
NAND2_X1 _u10_U5430  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n16868 ) );
NAND2_X1 _u10_U5429  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n16869 ) );
NAND2_X1 _u10_U5428  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n16870 ) );
NAND4_X1 _u10_U5427  ( .A1(_u10_n16867 ), .A2(_u10_n16868 ), .A3(_u10_n16869 ), .A4(_u10_n16870 ), .ZN(_u10_n16852 ) );
NAND2_X1 _u10_U5426  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n16863 ) );
NAND2_X1 _u10_U5425  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n16864 ) );
NAND2_X1 _u10_U5424  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n16865 ) );
NAND2_X1 _u10_U5423  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n16866 ) );
NAND4_X1 _u10_U5422  ( .A1(_u10_n16863 ), .A2(_u10_n16864 ), .A3(_u10_n16865 ), .A4(_u10_n16866 ), .ZN(_u10_n16853 ) );
NAND2_X1 _u10_U5421  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n16859 ) );
NAND2_X1 _u10_U5420  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n16860 ) );
NAND2_X1 _u10_U5419  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n16861 ) );
NAND2_X1 _u10_U5418  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n16862 ) );
NAND4_X1 _u10_U5417  ( .A1(_u10_n16859 ), .A2(_u10_n16860 ), .A3(_u10_n16861 ), .A4(_u10_n16862 ), .ZN(_u10_n16854 ) );
NAND2_X1 _u10_U5416  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n16856 ) );
NAND2_X1 _u10_U5415  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n16857 ) );
NAND2_X1 _u10_U5414  ( .A1(1'b0), .A2(_u10_n12011 ), .ZN(_u10_n16858 ) );
NAND3_X1 _u10_U5413  ( .A1(_u10_n16856 ), .A2(_u10_n16857 ), .A3(_u10_n16858 ), .ZN(_u10_n16855 ) );
NOR4_X1 _u10_U5412  ( .A1(_u10_n16852 ), .A2(_u10_n16853 ), .A3(_u10_n16854 ), .A4(_u10_n16855 ), .ZN(_u10_n16830 ) );
NAND2_X1 _u10_U5411  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n16848 ) );
NAND2_X1 _u10_U5410  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n16849 ) );
NAND2_X1 _u10_U5409  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n16850 ) );
NAND2_X1 _u10_U5408  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n16851 ) );
NAND4_X1 _u10_U5407  ( .A1(_u10_n16848 ), .A2(_u10_n16849 ), .A3(_u10_n16850 ), .A4(_u10_n16851 ), .ZN(_u10_n16832 ) );
NAND2_X1 _u10_U5406  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n16844 ) );
NAND2_X1 _u10_U5405  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n16845 ) );
NAND2_X1 _u10_U5404  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n16846 ) );
NAND2_X1 _u10_U5403  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n16847 ) );
NAND4_X1 _u10_U5402  ( .A1(_u10_n16844 ), .A2(_u10_n16845 ), .A3(_u10_n16846 ), .A4(_u10_n16847 ), .ZN(_u10_n16833 ) );
NAND2_X1 _u10_U5401  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n16840 ) );
NAND2_X1 _u10_U5400  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n16841 ) );
NAND2_X1 _u10_U5399  ( .A1(1'b0), .A2(_u10_n11758 ), .ZN(_u10_n16842 ) );
NAND2_X1 _u10_U5398  ( .A1(1'b0), .A2(_u10_n11734 ), .ZN(_u10_n16843 ) );
NAND4_X1 _u10_U5397  ( .A1(_u10_n16840 ), .A2(_u10_n16841 ), .A3(_u10_n16842 ), .A4(_u10_n16843 ), .ZN(_u10_n16834 ) );
NAND2_X1 _u10_U5396  ( .A1(1'b0), .A2(_u10_n11710 ), .ZN(_u10_n16836 ) );
NAND2_X1 _u10_U5395  ( .A1(1'b0), .A2(_u10_n11686 ), .ZN(_u10_n16837 ) );
NAND2_X1 _u10_U5394  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n16838 ) );
NAND2_X1 _u10_U5393  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n16839 ) );
NAND4_X1 _u10_U5392  ( .A1(_u10_n16836 ), .A2(_u10_n16837 ), .A3(_u10_n16838 ), .A4(_u10_n16839 ), .ZN(_u10_n16835 ) );
NOR4_X1 _u10_U5391  ( .A1(_u10_n16832 ), .A2(_u10_n16833 ), .A3(_u10_n16834 ), .A4(_u10_n16835 ), .ZN(_u10_n16831 ) );
NAND2_X1 _u10_U5390  ( .A1(_u10_n16830 ), .A2(_u10_n16831 ), .ZN(csr[28]) );
NAND2_X1 _u10_U5389  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n16826 ) );
NAND2_X1 _u10_U5388  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n16827 ) );
NAND2_X1 _u10_U5387  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n16828 ) );
NAND2_X1 _u10_U5386  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n16829 ) );
NAND4_X1 _u10_U5385  ( .A1(_u10_n16826 ), .A2(_u10_n16827 ), .A3(_u10_n16828 ), .A4(_u10_n16829 ), .ZN(_u10_n16811 ) );
NAND2_X1 _u10_U5384  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n16822 ) );
NAND2_X1 _u10_U5383  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n16823 ) );
NAND2_X1 _u10_U5382  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n16824 ) );
NAND2_X1 _u10_U5381  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n16825 ) );
NAND4_X1 _u10_U5380  ( .A1(_u10_n16822 ), .A2(_u10_n16823 ), .A3(_u10_n16824 ), .A4(_u10_n16825 ), .ZN(_u10_n16812 ) );
NAND2_X1 _u10_U5379  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n16818 ) );
NAND2_X1 _u10_U5378  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n16819 ) );
NAND2_X1 _u10_U5377  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n16820 ) );
NAND2_X1 _u10_U5376  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n16821 ) );
NAND4_X1 _u10_U5375  ( .A1(_u10_n16818 ), .A2(_u10_n16819 ), .A3(_u10_n16820 ), .A4(_u10_n16821 ), .ZN(_u10_n16813 ) );
NAND2_X1 _u10_U5374  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n16815 ) );
NAND2_X1 _u10_U5373  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n16816 ) );
NAND2_X1 _u10_U5372  ( .A1(1'b0), .A2(_u10_n12011 ), .ZN(_u10_n16817 ) );
NAND3_X1 _u10_U5371  ( .A1(_u10_n16815 ), .A2(_u10_n16816 ), .A3(_u10_n16817 ), .ZN(_u10_n16814 ) );
NOR4_X1 _u10_U5370  ( .A1(_u10_n16811 ), .A2(_u10_n16812 ), .A3(_u10_n16813 ), .A4(_u10_n16814 ), .ZN(_u10_n16789 ) );
NAND2_X1 _u10_U5369  ( .A1(1'b0), .A2(_u10_n11977 ), .ZN(_u10_n16807 ) );
NAND2_X1 _u10_U5368  ( .A1(1'b0), .A2(_u10_n11953 ), .ZN(_u10_n16808 ) );
NAND2_X1 _u10_U5367  ( .A1(1'b0), .A2(_u10_n11929 ), .ZN(_u10_n16809 ) );
NAND2_X1 _u10_U5366  ( .A1(1'b0), .A2(_u10_n11905 ), .ZN(_u10_n16810 ) );
NAND4_X1 _u10_U5365  ( .A1(_u10_n16807 ), .A2(_u10_n16808 ), .A3(_u10_n16809 ), .A4(_u10_n16810 ), .ZN(_u10_n16791 ) );
NAND2_X1 _u10_U5364  ( .A1(1'b0), .A2(_u10_n11881 ), .ZN(_u10_n16803 ) );
NAND2_X1 _u10_U5363  ( .A1(1'b0), .A2(_u10_n11857 ), .ZN(_u10_n16804 ) );
NAND2_X1 _u10_U5362  ( .A1(1'b0), .A2(_u10_n11833 ), .ZN(_u10_n16805 ) );
NAND2_X1 _u10_U5361  ( .A1(1'b0), .A2(_u10_n11809 ), .ZN(_u10_n16806 ) );
NAND4_X1 _u10_U5360  ( .A1(_u10_n16803 ), .A2(_u10_n16804 ), .A3(_u10_n16805 ), .A4(_u10_n16806 ), .ZN(_u10_n16792 ) );
NAND2_X1 _u10_U5359  ( .A1(1'b0), .A2(_u10_n11785 ), .ZN(_u10_n16799 ) );
NAND2_X1 _u10_U5358  ( .A1(1'b0), .A2(_u10_n11761 ), .ZN(_u10_n16800 ) );
NAND2_X1 _u10_U5357  ( .A1(1'b0), .A2(_u10_n11759 ), .ZN(_u10_n16801 ) );
NAND2_X1 _u10_U5356  ( .A1(1'b0), .A2(_u10_n11735 ), .ZN(_u10_n16802 ) );
NAND4_X1 _u10_U5355  ( .A1(_u10_n16799 ), .A2(_u10_n16800 ), .A3(_u10_n16801 ), .A4(_u10_n16802 ), .ZN(_u10_n16793 ) );
NAND2_X1 _u10_U5354  ( .A1(1'b0), .A2(_u10_n11711 ), .ZN(_u10_n16795 ) );
NAND2_X1 _u10_U5353  ( .A1(1'b0), .A2(_u10_n11687 ), .ZN(_u10_n16796 ) );
NAND2_X1 _u10_U5352  ( .A1(1'b0), .A2(_u10_n11641 ), .ZN(_u10_n16797 ) );
NAND2_X1 _u10_U5351  ( .A1(1'b0), .A2(_u10_n11617 ), .ZN(_u10_n16798 ) );
NAND4_X1 _u10_U5350  ( .A1(_u10_n16795 ), .A2(_u10_n16796 ), .A3(_u10_n16797 ), .A4(_u10_n16798 ), .ZN(_u10_n16794 ) );
NOR4_X1 _u10_U5349  ( .A1(_u10_n16791 ), .A2(_u10_n16792 ), .A3(_u10_n16793 ), .A4(_u10_n16794 ), .ZN(_u10_n16790 ) );
NAND2_X1 _u10_U5348  ( .A1(_u10_n16789 ), .A2(_u10_n16790 ), .ZN(csr[29]) );
NAND2_X1 _u10_U5347  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n16785 ) );
NAND2_X1 _u10_U5346  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n16786 ) );
NAND2_X1 _u10_U5345  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n16787 ) );
NAND2_X1 _u10_U5344  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n16788 ) );
NAND4_X1 _u10_U5343  ( .A1(_u10_n16785 ), .A2(_u10_n16786 ), .A3(_u10_n16787 ), .A4(_u10_n16788 ), .ZN(_u10_n16770 ) );
NAND2_X1 _u10_U5342  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n16781 ) );
NAND2_X1 _u10_U5341  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n16782 ) );
NAND2_X1 _u10_U5340  ( .A1(1'b0), .A2(_u10_n12206 ), .ZN(_u10_n16783 ) );
NAND2_X1 _u10_U5339  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n16784 ) );
NAND4_X1 _u10_U5338  ( .A1(_u10_n16781 ), .A2(_u10_n16782 ), .A3(_u10_n16783 ), .A4(_u10_n16784 ), .ZN(_u10_n16771 ) );
NAND2_X1 _u10_U5337  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n16777 ) );
NAND2_X1 _u10_U5336  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n16778 ) );
NAND2_X1 _u10_U5335  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n16779 ) );
NAND2_X1 _u10_U5334  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n16780 ) );
NAND4_X1 _u10_U5333  ( .A1(_u10_n16777 ), .A2(_u10_n16778 ), .A3(_u10_n16779 ), .A4(_u10_n16780 ), .ZN(_u10_n16772 ) );
NAND2_X1 _u10_U5332  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n16774 ) );
NAND2_X1 _u10_U5331  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n16775 ) );
NAND2_X1 _u10_U5330  ( .A1(ch0_csr[2]), .A2(_u10_n12011 ), .ZN(_u10_n16776 ));
NAND3_X1 _u10_U5329  ( .A1(_u10_n16774 ), .A2(_u10_n16775 ), .A3(_u10_n16776 ), .ZN(_u10_n16773 ) );
NOR4_X1 _u10_U5328  ( .A1(_u10_n16770 ), .A2(_u10_n16771 ), .A3(_u10_n16772 ), .A4(_u10_n16773 ), .ZN(_u10_n16748 ) );
NAND2_X1 _u10_U5327  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16766 ) );
NAND2_X1 _u10_U5326  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16767 ) );
NAND2_X1 _u10_U5325  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16768 ) );
NAND2_X1 _u10_U5324  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16769 ) );
NAND4_X1 _u10_U5323  ( .A1(_u10_n16766 ), .A2(_u10_n16767 ), .A3(_u10_n16768 ), .A4(_u10_n16769 ), .ZN(_u10_n16750 ) );
NAND2_X1 _u10_U5322  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16762 ) );
NAND2_X1 _u10_U5321  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16763 ) );
NAND2_X1 _u10_U5320  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16764 ) );
NAND2_X1 _u10_U5319  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16765 ) );
NAND4_X1 _u10_U5318  ( .A1(_u10_n16762 ), .A2(_u10_n16763 ), .A3(_u10_n16764 ), .A4(_u10_n16765 ), .ZN(_u10_n16751 ) );
NAND2_X1 _u10_U5317  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16758 ) );
NAND2_X1 _u10_U5316  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16759 ) );
NAND2_X1 _u10_U5315  ( .A1(1'b0), .A2(_u10_n11755 ), .ZN(_u10_n16760 ) );
NAND2_X1 _u10_U5314  ( .A1(1'b0), .A2(_u10_n11731 ), .ZN(_u10_n16761 ) );
NAND4_X1 _u10_U5313  ( .A1(_u10_n16758 ), .A2(_u10_n16759 ), .A3(_u10_n16760 ), .A4(_u10_n16761 ), .ZN(_u10_n16752 ) );
NAND2_X1 _u10_U5312  ( .A1(1'b0), .A2(_u10_n11707 ), .ZN(_u10_n16754 ) );
NAND2_X1 _u10_U5311  ( .A1(1'b0), .A2(_u10_n11683 ), .ZN(_u10_n16755 ) );
NAND2_X1 _u10_U5310  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16756 ) );
NAND2_X1 _u10_U5309  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16757 ) );
NAND4_X1 _u10_U5308  ( .A1(_u10_n16754 ), .A2(_u10_n16755 ), .A3(_u10_n16756 ), .A4(_u10_n16757 ), .ZN(_u10_n16753 ) );
NOR4_X1 _u10_U5307  ( .A1(_u10_n16750 ), .A2(_u10_n16751 ), .A3(_u10_n16752 ), .A4(_u10_n16753 ), .ZN(_u10_n16749 ) );
NAND2_X1 _u10_U5306  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n16744 ) );
NAND2_X1 _u10_U5305  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n16745 ) );
NAND2_X1 _u10_U5304  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n16746 ) );
NAND2_X1 _u10_U5303  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n16747 ) );
NAND4_X1 _u10_U5302  ( .A1(_u10_n16744 ), .A2(_u10_n16745 ), .A3(_u10_n16746 ), .A4(_u10_n16747 ), .ZN(_u10_n16729 ) );
NAND2_X1 _u10_U5301  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n16740 ) );
NAND2_X1 _u10_U5300  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n16741 ) );
NAND2_X1 _u10_U5299  ( .A1(1'b0), .A2(_u10_n12209 ), .ZN(_u10_n16742 ) );
NAND2_X1 _u10_U5298  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n16743 ) );
NAND4_X1 _u10_U5297  ( .A1(_u10_n16740 ), .A2(_u10_n16741 ), .A3(_u10_n16742 ), .A4(_u10_n16743 ), .ZN(_u10_n16730 ) );
NAND2_X1 _u10_U5296  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n16736 ) );
NAND2_X1 _u10_U5295  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n16737 ) );
NAND2_X1 _u10_U5294  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n16738 ) );
NAND2_X1 _u10_U5293  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n16739 ) );
NAND4_X1 _u10_U5292  ( .A1(_u10_n16736 ), .A2(_u10_n16737 ), .A3(_u10_n16738 ), .A4(_u10_n16739 ), .ZN(_u10_n16731 ) );
NAND2_X1 _u10_U5291  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n16733 ) );
NAND2_X1 _u10_U5290  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n16734 ) );
NAND2_X1 _u10_U5289  ( .A1(1'b0), .A2(_u10_n12011 ), .ZN(_u10_n16735 ) );
NAND3_X1 _u10_U5288  ( .A1(_u10_n16733 ), .A2(_u10_n16734 ), .A3(_u10_n16735 ), .ZN(_u10_n16732 ) );
NOR4_X1 _u10_U5287  ( .A1(_u10_n16729 ), .A2(_u10_n16730 ), .A3(_u10_n16731 ), .A4(_u10_n16732 ), .ZN(_u10_n16707 ) );
NAND2_X1 _u10_U5286  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16725 ) );
NAND2_X1 _u10_U5285  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16726 ) );
NAND2_X1 _u10_U5284  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16727 ) );
NAND2_X1 _u10_U5283  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16728 ) );
NAND4_X1 _u10_U5282  ( .A1(_u10_n16725 ), .A2(_u10_n16726 ), .A3(_u10_n16727 ), .A4(_u10_n16728 ), .ZN(_u10_n16709 ) );
NAND2_X1 _u10_U5281  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16721 ) );
NAND2_X1 _u10_U5280  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16722 ) );
NAND2_X1 _u10_U5279  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16723 ) );
NAND2_X1 _u10_U5278  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16724 ) );
NAND4_X1 _u10_U5277  ( .A1(_u10_n16721 ), .A2(_u10_n16722 ), .A3(_u10_n16723 ), .A4(_u10_n16724 ), .ZN(_u10_n16710 ) );
NAND2_X1 _u10_U5276  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16717 ) );
NAND2_X1 _u10_U5275  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16718 ) );
NAND2_X1 _u10_U5274  ( .A1(1'b0), .A2(_u10_n11754 ), .ZN(_u10_n16719 ) );
NAND2_X1 _u10_U5273  ( .A1(1'b0), .A2(_u10_n11730 ), .ZN(_u10_n16720 ) );
NAND4_X1 _u10_U5272  ( .A1(_u10_n16717 ), .A2(_u10_n16718 ), .A3(_u10_n16719 ), .A4(_u10_n16720 ), .ZN(_u10_n16711 ) );
NAND2_X1 _u10_U5271  ( .A1(1'b0), .A2(_u10_n11706 ), .ZN(_u10_n16713 ) );
NAND2_X1 _u10_U5270  ( .A1(1'b0), .A2(_u10_n11682 ), .ZN(_u10_n16714 ) );
NAND2_X1 _u10_U5269  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16715 ) );
NAND2_X1 _u10_U5268  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16716 ) );
NAND4_X1 _u10_U5267  ( .A1(_u10_n16713 ), .A2(_u10_n16714 ), .A3(_u10_n16715 ), .A4(_u10_n16716 ), .ZN(_u10_n16712 ) );
NOR4_X1 _u10_U5266  ( .A1(_u10_n16709 ), .A2(_u10_n16710 ), .A3(_u10_n16711 ), .A4(_u10_n16712 ), .ZN(_u10_n16708 ) );
NAND2_X1 _u10_U5265  ( .A1(_u10_n16707 ), .A2(_u10_n16708 ), .ZN(csr[30]) );
NAND2_X1 _u10_U5264  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n16703 ) );
NAND2_X1 _u10_U5263  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n16704 ) );
NAND2_X1 _u10_U5262  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n16705 ) );
NAND2_X1 _u10_U5261  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n16706 ) );
NAND4_X1 _u10_U5260  ( .A1(_u10_n16703 ), .A2(_u10_n16704 ), .A3(_u10_n16705 ), .A4(_u10_n16706 ), .ZN(_u10_n16688 ) );
NAND2_X1 _u10_U5259  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n16699 ) );
NAND2_X1 _u10_U5258  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n16700 ) );
NAND2_X1 _u10_U5257  ( .A1(1'b0), .A2(_u10_n12211 ), .ZN(_u10_n16701 ) );
NAND2_X1 _u10_U5256  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n16702 ) );
NAND4_X1 _u10_U5255  ( .A1(_u10_n16699 ), .A2(_u10_n16700 ), .A3(_u10_n16701 ), .A4(_u10_n16702 ), .ZN(_u10_n16689 ) );
NAND2_X1 _u10_U5254  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n16695 ) );
NAND2_X1 _u10_U5253  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n16696 ) );
NAND2_X1 _u10_U5252  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n16697 ) );
NAND2_X1 _u10_U5251  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n16698 ) );
NAND4_X1 _u10_U5250  ( .A1(_u10_n16695 ), .A2(_u10_n16696 ), .A3(_u10_n16697 ), .A4(_u10_n16698 ), .ZN(_u10_n16690 ) );
NAND2_X1 _u10_U5249  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n16692 ) );
NAND2_X1 _u10_U5248  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n16693 ) );
NAND2_X1 _u10_U5247  ( .A1(1'b0), .A2(_u10_n12011 ), .ZN(_u10_n16694 ) );
NAND3_X1 _u10_U5246  ( .A1(_u10_n16692 ), .A2(_u10_n16693 ), .A3(_u10_n16694 ), .ZN(_u10_n16691 ) );
NOR4_X1 _u10_U5245  ( .A1(_u10_n16688 ), .A2(_u10_n16689 ), .A3(_u10_n16690 ), .A4(_u10_n16691 ), .ZN(_u10_n16666 ) );
NAND2_X1 _u10_U5244  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16684 ) );
NAND2_X1 _u10_U5243  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16685 ) );
NAND2_X1 _u10_U5242  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16686 ) );
NAND2_X1 _u10_U5241  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16687 ) );
NAND4_X1 _u10_U5240  ( .A1(_u10_n16684 ), .A2(_u10_n16685 ), .A3(_u10_n16686 ), .A4(_u10_n16687 ), .ZN(_u10_n16668 ) );
NAND2_X1 _u10_U5239  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16680 ) );
NAND2_X1 _u10_U5238  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16681 ) );
NAND2_X1 _u10_U5237  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16682 ) );
NAND2_X1 _u10_U5236  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16683 ) );
NAND4_X1 _u10_U5235  ( .A1(_u10_n16680 ), .A2(_u10_n16681 ), .A3(_u10_n16682 ), .A4(_u10_n16683 ), .ZN(_u10_n16669 ) );
NAND2_X1 _u10_U5234  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16676 ) );
NAND2_X1 _u10_U5233  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16677 ) );
NAND2_X1 _u10_U5232  ( .A1(1'b0), .A2(_u10_n12378 ), .ZN(_u10_n16678 ) );
NAND2_X1 _u10_U5231  ( .A1(1'b0), .A2(_u10_n12377 ), .ZN(_u10_n16679 ) );
NAND4_X1 _u10_U5230  ( .A1(_u10_n16676 ), .A2(_u10_n16677 ), .A3(_u10_n16678 ), .A4(_u10_n16679 ), .ZN(_u10_n16670 ) );
NAND2_X1 _u10_U5229  ( .A1(1'b0), .A2(_u10_n12372 ), .ZN(_u10_n16672 ) );
NAND2_X1 _u10_U5228  ( .A1(1'b0), .A2(_u10_n12371 ), .ZN(_u10_n16673 ) );
NAND2_X1 _u10_U5227  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16674 ) );
NAND2_X1 _u10_U5226  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16675 ) );
NAND4_X1 _u10_U5225  ( .A1(_u10_n16672 ), .A2(_u10_n16673 ), .A3(_u10_n16674 ), .A4(_u10_n16675 ), .ZN(_u10_n16671 ) );
NOR4_X1 _u10_U5224  ( .A1(_u10_n16668 ), .A2(_u10_n16669 ), .A3(_u10_n16670 ), .A4(_u10_n16671 ), .ZN(_u10_n16667 ) );
NAND2_X1 _u10_U5223  ( .A1(_u10_n16666 ), .A2(_u10_n16667 ), .ZN(csr[31]) );
NAND2_X1 _u10_U5222  ( .A1(1'b0), .A2(_u10_n12342 ), .ZN(_u10_n16662 ) );
NAND2_X1 _u10_U5221  ( .A1(1'b0), .A2(_u10_n12318 ), .ZN(_u10_n16663 ) );
NAND2_X1 _u10_U5220  ( .A1(1'b0), .A2(_u10_n12295 ), .ZN(_u10_n16664 ) );
NAND2_X1 _u10_U5219  ( .A1(1'b0), .A2(_u10_n12271 ), .ZN(_u10_n16665 ) );
NAND4_X1 _u10_U5218  ( .A1(_u10_n16662 ), .A2(_u10_n16663 ), .A3(_u10_n16664 ), .A4(_u10_n16665 ), .ZN(_u10_n16647 ) );
NAND2_X1 _u10_U5217  ( .A1(1'b0), .A2(_u10_n12246 ), .ZN(_u10_n16658 ) );
NAND2_X1 _u10_U5216  ( .A1(1'b0), .A2(_u10_n12222 ), .ZN(_u10_n16659 ) );
NAND2_X1 _u10_U5215  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n16660 ) );
NAND2_X1 _u10_U5214  ( .A1(1'b0), .A2(_u10_n12174 ), .ZN(_u10_n16661 ) );
NAND4_X1 _u10_U5213  ( .A1(_u10_n16658 ), .A2(_u10_n16659 ), .A3(_u10_n16660 ), .A4(_u10_n16661 ), .ZN(_u10_n16648 ) );
NAND2_X1 _u10_U5212  ( .A1(1'b0), .A2(_u10_n12151 ), .ZN(_u10_n16654 ) );
NAND2_X1 _u10_U5211  ( .A1(1'b0), .A2(_u10_n12127 ), .ZN(_u10_n16655 ) );
NAND2_X1 _u10_U5210  ( .A1(1'b0), .A2(_u10_n12103 ), .ZN(_u10_n16656 ) );
NAND2_X1 _u10_U5209  ( .A1(1'b0), .A2(_u10_n12079 ), .ZN(_u10_n16657 ) );
NAND4_X1 _u10_U5208  ( .A1(_u10_n16654 ), .A2(_u10_n16655 ), .A3(_u10_n16656 ), .A4(_u10_n16657 ), .ZN(_u10_n16649 ) );
NAND2_X1 _u10_U5207  ( .A1(1'b0), .A2(_u10_n12055 ), .ZN(_u10_n16651 ) );
NAND2_X1 _u10_U5206  ( .A1(1'b0), .A2(_u10_n12031 ), .ZN(_u10_n16652 ) );
NAND2_X1 _u10_U5205  ( .A1(ch0_csr[3]), .A2(_u10_n12011 ), .ZN(_u10_n16653 ));
NAND3_X1 _u10_U5204  ( .A1(_u10_n16651 ), .A2(_u10_n16652 ), .A3(_u10_n16653 ), .ZN(_u10_n16650 ) );
NOR4_X1 _u10_U5203  ( .A1(_u10_n16647 ), .A2(_u10_n16648 ), .A3(_u10_n16649 ), .A4(_u10_n16650 ), .ZN(_u10_n16625 ) );
NAND2_X1 _u10_U5202  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16643 ) );
NAND2_X1 _u10_U5201  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16644 ) );
NAND2_X1 _u10_U5200  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16645 ) );
NAND2_X1 _u10_U5199  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16646 ) );
NAND4_X1 _u10_U5198  ( .A1(_u10_n16643 ), .A2(_u10_n16644 ), .A3(_u10_n16645 ), .A4(_u10_n16646 ), .ZN(_u10_n16627 ) );
NAND2_X1 _u10_U5197  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16639 ) );
NAND2_X1 _u10_U5196  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16640 ) );
NAND2_X1 _u10_U5195  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16641 ) );
NAND2_X1 _u10_U5194  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16642 ) );
NAND4_X1 _u10_U5193  ( .A1(_u10_n16639 ), .A2(_u10_n16640 ), .A3(_u10_n16641 ), .A4(_u10_n16642 ), .ZN(_u10_n16628 ) );
NAND2_X1 _u10_U5192  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16635 ) );
NAND2_X1 _u10_U5191  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16636 ) );
NAND2_X1 _u10_U5190  ( .A1(1'b0), .A2(_u10_n11759 ), .ZN(_u10_n16637 ) );
NAND2_X1 _u10_U5189  ( .A1(1'b0), .A2(_u10_n11735 ), .ZN(_u10_n16638 ) );
NAND4_X1 _u10_U5188  ( .A1(_u10_n16635 ), .A2(_u10_n16636 ), .A3(_u10_n16637 ), .A4(_u10_n16638 ), .ZN(_u10_n16629 ) );
NAND2_X1 _u10_U5187  ( .A1(1'b0), .A2(_u10_n11711 ), .ZN(_u10_n16631 ) );
NAND2_X1 _u10_U5186  ( .A1(1'b0), .A2(_u10_n11687 ), .ZN(_u10_n16632 ) );
NAND2_X1 _u10_U5185  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16633 ) );
NAND2_X1 _u10_U5184  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16634 ) );
NAND4_X1 _u10_U5183  ( .A1(_u10_n16631 ), .A2(_u10_n16632 ), .A3(_u10_n16633 ), .A4(_u10_n16634 ), .ZN(_u10_n16630 ) );
NOR4_X1 _u10_U5182  ( .A1(_u10_n16627 ), .A2(_u10_n16628 ), .A3(_u10_n16629 ), .A4(_u10_n16630 ), .ZN(_u10_n16626 ) );
NAND2_X1 _u10_U5181  ( .A1(_u10_n16625 ), .A2(_u10_n16626 ), .ZN(csr[3]) );
NAND2_X1 _u10_U5180  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16621 ) );
NAND2_X1 _u10_U5179  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16622 ) );
NAND2_X1 _u10_U5178  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16623 ) );
NAND2_X1 _u10_U5177  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16624 ) );
NAND4_X1 _u10_U5176  ( .A1(_u10_n16621 ), .A2(_u10_n16622 ), .A3(_u10_n16623 ), .A4(_u10_n16624 ), .ZN(_u10_n16606 ) );
NAND2_X1 _u10_U5175  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16617 ) );
NAND2_X1 _u10_U5174  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16618 ) );
NAND2_X1 _u10_U5173  ( .A1(1'b0), .A2(_u10_n12210 ), .ZN(_u10_n16619 ) );
NAND2_X1 _u10_U5172  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16620 ) );
NAND4_X1 _u10_U5171  ( .A1(_u10_n16617 ), .A2(_u10_n16618 ), .A3(_u10_n16619 ), .A4(_u10_n16620 ), .ZN(_u10_n16607 ) );
NAND2_X1 _u10_U5170  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16613 ) );
NAND2_X1 _u10_U5169  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16614 ) );
NAND2_X1 _u10_U5168  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16615 ) );
NAND2_X1 _u10_U5167  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16616 ) );
NAND4_X1 _u10_U5166  ( .A1(_u10_n16613 ), .A2(_u10_n16614 ), .A3(_u10_n16615 ), .A4(_u10_n16616 ), .ZN(_u10_n16608 ) );
NAND2_X1 _u10_U5165  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16610 ) );
NAND2_X1 _u10_U5164  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16611 ) );
NAND2_X1 _u10_U5163  ( .A1(ch0_csr[4]), .A2(_u10_n12011 ), .ZN(_u10_n16612 ));
NAND3_X1 _u10_U5162  ( .A1(_u10_n16610 ), .A2(_u10_n16611 ), .A3(_u10_n16612 ), .ZN(_u10_n16609 ) );
NOR4_X1 _u10_U5161  ( .A1(_u10_n16606 ), .A2(_u10_n16607 ), .A3(_u10_n16608 ), .A4(_u10_n16609 ), .ZN(_u10_n16584 ) );
NAND2_X1 _u10_U5160  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16602 ) );
NAND2_X1 _u10_U5159  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16603 ) );
NAND2_X1 _u10_U5158  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16604 ) );
NAND2_X1 _u10_U5157  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16605 ) );
NAND4_X1 _u10_U5156  ( .A1(_u10_n16602 ), .A2(_u10_n16603 ), .A3(_u10_n16604 ), .A4(_u10_n16605 ), .ZN(_u10_n16586 ) );
NAND2_X1 _u10_U5155  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16598 ) );
NAND2_X1 _u10_U5154  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16599 ) );
NAND2_X1 _u10_U5153  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16600 ) );
NAND2_X1 _u10_U5152  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16601 ) );
NAND4_X1 _u10_U5151  ( .A1(_u10_n16598 ), .A2(_u10_n16599 ), .A3(_u10_n16600 ), .A4(_u10_n16601 ), .ZN(_u10_n16587 ) );
NAND2_X1 _u10_U5150  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16594 ) );
NAND2_X1 _u10_U5149  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16595 ) );
NAND2_X1 _u10_U5148  ( .A1(1'b0), .A2(_u10_n11756 ), .ZN(_u10_n16596 ) );
NAND2_X1 _u10_U5147  ( .A1(1'b0), .A2(_u10_n11732 ), .ZN(_u10_n16597 ) );
NAND4_X1 _u10_U5146  ( .A1(_u10_n16594 ), .A2(_u10_n16595 ), .A3(_u10_n16596 ), .A4(_u10_n16597 ), .ZN(_u10_n16588 ) );
NAND2_X1 _u10_U5145  ( .A1(1'b0), .A2(_u10_n11708 ), .ZN(_u10_n16590 ) );
NAND2_X1 _u10_U5144  ( .A1(1'b0), .A2(_u10_n11684 ), .ZN(_u10_n16591 ) );
NAND2_X1 _u10_U5143  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16592 ) );
NAND2_X1 _u10_U5142  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16593 ) );
NAND4_X1 _u10_U5141  ( .A1(_u10_n16590 ), .A2(_u10_n16591 ), .A3(_u10_n16592 ), .A4(_u10_n16593 ), .ZN(_u10_n16589 ) );
NOR4_X1 _u10_U5140  ( .A1(_u10_n16586 ), .A2(_u10_n16587 ), .A3(_u10_n16588 ), .A4(_u10_n16589 ), .ZN(_u10_n16585 ) );
NAND2_X1 _u10_U5139  ( .A1(_u10_n16584 ), .A2(_u10_n16585 ), .ZN(csr[4]) );
NAND2_X1 _u10_U5138  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16580 ) );
NAND2_X1 _u10_U5137  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16581 ) );
NAND2_X1 _u10_U5136  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16582 ) );
NAND2_X1 _u10_U5135  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16583 ) );
NAND4_X1 _u10_U5134  ( .A1(_u10_n16580 ), .A2(_u10_n16581 ), .A3(_u10_n16582 ), .A4(_u10_n16583 ), .ZN(_u10_n16565 ) );
NAND2_X1 _u10_U5133  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16576 ) );
NAND2_X1 _u10_U5132  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16577 ) );
NAND2_X1 _u10_U5131  ( .A1(1'b0), .A2(_u10_n12207 ), .ZN(_u10_n16578 ) );
NAND2_X1 _u10_U5130  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16579 ) );
NAND4_X1 _u10_U5129  ( .A1(_u10_n16576 ), .A2(_u10_n16577 ), .A3(_u10_n16578 ), .A4(_u10_n16579 ), .ZN(_u10_n16566 ) );
NAND2_X1 _u10_U5128  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16572 ) );
NAND2_X1 _u10_U5127  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16573 ) );
NAND2_X1 _u10_U5126  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16574 ) );
NAND2_X1 _u10_U5125  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16575 ) );
NAND4_X1 _u10_U5124  ( .A1(_u10_n16572 ), .A2(_u10_n16573 ), .A3(_u10_n16574 ), .A4(_u10_n16575 ), .ZN(_u10_n16567 ) );
NAND2_X1 _u10_U5123  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16569 ) );
NAND2_X1 _u10_U5122  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16570 ) );
NAND2_X1 _u10_U5121  ( .A1(ch0_csr[5]), .A2(_u10_n12012 ), .ZN(_u10_n16571 ));
NAND3_X1 _u10_U5120  ( .A1(_u10_n16569 ), .A2(_u10_n16570 ), .A3(_u10_n16571 ), .ZN(_u10_n16568 ) );
NOR4_X1 _u10_U5119  ( .A1(_u10_n16565 ), .A2(_u10_n16566 ), .A3(_u10_n16567 ), .A4(_u10_n16568 ), .ZN(_u10_n16543 ) );
NAND2_X1 _u10_U5118  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16561 ) );
NAND2_X1 _u10_U5117  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16562 ) );
NAND2_X1 _u10_U5116  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16563 ) );
NAND2_X1 _u10_U5115  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16564 ) );
NAND4_X1 _u10_U5114  ( .A1(_u10_n16561 ), .A2(_u10_n16562 ), .A3(_u10_n16563 ), .A4(_u10_n16564 ), .ZN(_u10_n16545 ) );
NAND2_X1 _u10_U5113  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16557 ) );
NAND2_X1 _u10_U5112  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16558 ) );
NAND2_X1 _u10_U5111  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16559 ) );
NAND2_X1 _u10_U5110  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16560 ) );
NAND4_X1 _u10_U5109  ( .A1(_u10_n16557 ), .A2(_u10_n16558 ), .A3(_u10_n16559 ), .A4(_u10_n16560 ), .ZN(_u10_n16546 ) );
NAND2_X1 _u10_U5108  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16553 ) );
NAND2_X1 _u10_U5107  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16554 ) );
NAND2_X1 _u10_U5106  ( .A1(1'b0), .A2(_u10_n11753 ), .ZN(_u10_n16555 ) );
NAND2_X1 _u10_U5105  ( .A1(1'b0), .A2(_u10_n11729 ), .ZN(_u10_n16556 ) );
NAND4_X1 _u10_U5104  ( .A1(_u10_n16553 ), .A2(_u10_n16554 ), .A3(_u10_n16555 ), .A4(_u10_n16556 ), .ZN(_u10_n16547 ) );
NAND2_X1 _u10_U5103  ( .A1(1'b0), .A2(_u10_n11705 ), .ZN(_u10_n16549 ) );
NAND2_X1 _u10_U5102  ( .A1(1'b0), .A2(_u10_n11681 ), .ZN(_u10_n16550 ) );
NAND2_X1 _u10_U5101  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16551 ) );
NAND2_X1 _u10_U5100  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16552 ) );
NAND4_X1 _u10_U5099  ( .A1(_u10_n16549 ), .A2(_u10_n16550 ), .A3(_u10_n16551 ), .A4(_u10_n16552 ), .ZN(_u10_n16548 ) );
NOR4_X1 _u10_U5098  ( .A1(_u10_n16545 ), .A2(_u10_n16546 ), .A3(_u10_n16547 ), .A4(_u10_n16548 ), .ZN(_u10_n16544 ) );
NAND2_X1 _u10_U5097  ( .A1(_u10_n16543 ), .A2(_u10_n16544 ), .ZN(csr[5]) );
NAND2_X1 _u10_U5096  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16539 ) );
NAND2_X1 _u10_U5095  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16540 ) );
NAND2_X1 _u10_U5094  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16541 ) );
NAND2_X1 _u10_U5093  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16542 ) );
NAND4_X1 _u10_U5092  ( .A1(_u10_n16539 ), .A2(_u10_n16540 ), .A3(_u10_n16541 ), .A4(_u10_n16542 ), .ZN(_u10_n16524 ) );
NAND2_X1 _u10_U5091  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16535 ) );
NAND2_X1 _u10_U5090  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16536 ) );
NAND2_X1 _u10_U5089  ( .A1(1'b0), .A2(_u10_n12420 ), .ZN(_u10_n16537 ) );
NAND2_X1 _u10_U5088  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16538 ) );
NAND4_X1 _u10_U5087  ( .A1(_u10_n16535 ), .A2(_u10_n16536 ), .A3(_u10_n16537 ), .A4(_u10_n16538 ), .ZN(_u10_n16525 ) );
NAND2_X1 _u10_U5086  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16531 ) );
NAND2_X1 _u10_U5085  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16532 ) );
NAND2_X1 _u10_U5084  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16533 ) );
NAND2_X1 _u10_U5083  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16534 ) );
NAND4_X1 _u10_U5082  ( .A1(_u10_n16531 ), .A2(_u10_n16532 ), .A3(_u10_n16533 ), .A4(_u10_n16534 ), .ZN(_u10_n16526 ) );
NAND2_X1 _u10_U5081  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16528 ) );
NAND2_X1 _u10_U5080  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16529 ) );
NAND2_X1 _u10_U5079  ( .A1(ch0_csr[6]), .A2(_u10_n12012 ), .ZN(_u10_n16530 ));
NAND3_X1 _u10_U5078  ( .A1(_u10_n16528 ), .A2(_u10_n16529 ), .A3(_u10_n16530 ), .ZN(_u10_n16527 ) );
NOR4_X1 _u10_U5077  ( .A1(_u10_n16524 ), .A2(_u10_n16525 ), .A3(_u10_n16526 ), .A4(_u10_n16527 ), .ZN(_u10_n16502 ) );
NAND2_X1 _u10_U5076  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16520 ) );
NAND2_X1 _u10_U5075  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16521 ) );
NAND2_X1 _u10_U5074  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16522 ) );
NAND2_X1 _u10_U5073  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16523 ) );
NAND4_X1 _u10_U5072  ( .A1(_u10_n16520 ), .A2(_u10_n16521 ), .A3(_u10_n16522 ), .A4(_u10_n16523 ), .ZN(_u10_n16504 ) );
NAND2_X1 _u10_U5071  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16516 ) );
NAND2_X1 _u10_U5070  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16517 ) );
NAND2_X1 _u10_U5069  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16518 ) );
NAND2_X1 _u10_U5068  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16519 ) );
NAND4_X1 _u10_U5067  ( .A1(_u10_n16516 ), .A2(_u10_n16517 ), .A3(_u10_n16518 ), .A4(_u10_n16519 ), .ZN(_u10_n16505 ) );
NAND2_X1 _u10_U5066  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16512 ) );
NAND2_X1 _u10_U5065  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16513 ) );
NAND2_X1 _u10_U5064  ( .A1(1'b0), .A2(_u10_n11758 ), .ZN(_u10_n16514 ) );
NAND2_X1 _u10_U5063  ( .A1(1'b0), .A2(_u10_n11734 ), .ZN(_u10_n16515 ) );
NAND4_X1 _u10_U5062  ( .A1(_u10_n16512 ), .A2(_u10_n16513 ), .A3(_u10_n16514 ), .A4(_u10_n16515 ), .ZN(_u10_n16506 ) );
NAND2_X1 _u10_U5061  ( .A1(1'b0), .A2(_u10_n11710 ), .ZN(_u10_n16508 ) );
NAND2_X1 _u10_U5060  ( .A1(1'b0), .A2(_u10_n11686 ), .ZN(_u10_n16509 ) );
NAND2_X1 _u10_U5059  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16510 ) );
NAND2_X1 _u10_U5058  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16511 ) );
NAND4_X1 _u10_U5057  ( .A1(_u10_n16508 ), .A2(_u10_n16509 ), .A3(_u10_n16510 ), .A4(_u10_n16511 ), .ZN(_u10_n16507 ) );
NOR4_X1 _u10_U5056  ( .A1(_u10_n16504 ), .A2(_u10_n16505 ), .A3(_u10_n16506 ), .A4(_u10_n16507 ), .ZN(_u10_n16503 ) );
NAND2_X1 _u10_U5055  ( .A1(_u10_n16502 ), .A2(_u10_n16503 ), .ZN(csr[6]) );
NAND2_X1 _u10_U5054  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16498 ) );
NAND2_X1 _u10_U5053  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16499 ) );
NAND2_X1 _u10_U5052  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16500 ) );
NAND2_X1 _u10_U5051  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16501 ) );
NAND4_X1 _u10_U5050  ( .A1(_u10_n16498 ), .A2(_u10_n16499 ), .A3(_u10_n16500 ), .A4(_u10_n16501 ), .ZN(_u10_n16483 ) );
NAND2_X1 _u10_U5049  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16494 ) );
NAND2_X1 _u10_U5048  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16495 ) );
NAND2_X1 _u10_U5047  ( .A1(1'b0), .A2(_u10_n12212 ), .ZN(_u10_n16496 ) );
NAND2_X1 _u10_U5046  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16497 ) );
NAND4_X1 _u10_U5045  ( .A1(_u10_n16494 ), .A2(_u10_n16495 ), .A3(_u10_n16496 ), .A4(_u10_n16497 ), .ZN(_u10_n16484 ) );
NAND2_X1 _u10_U5044  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16490 ) );
NAND2_X1 _u10_U5043  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16491 ) );
NAND2_X1 _u10_U5042  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16492 ) );
NAND2_X1 _u10_U5041  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16493 ) );
NAND4_X1 _u10_U5040  ( .A1(_u10_n16490 ), .A2(_u10_n16491 ), .A3(_u10_n16492 ), .A4(_u10_n16493 ), .ZN(_u10_n16485 ) );
NAND2_X1 _u10_U5039  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16487 ) );
NAND2_X1 _u10_U5038  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16488 ) );
NAND2_X1 _u10_U5037  ( .A1(ch0_csr[7]), .A2(_u10_n12012 ), .ZN(_u10_n16489 ));
NAND3_X1 _u10_U5036  ( .A1(_u10_n16487 ), .A2(_u10_n16488 ), .A3(_u10_n16489 ), .ZN(_u10_n16486 ) );
NOR4_X1 _u10_U5035  ( .A1(_u10_n16483 ), .A2(_u10_n16484 ), .A3(_u10_n16485 ), .A4(_u10_n16486 ), .ZN(_u10_n16461 ) );
NAND2_X1 _u10_U5034  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16479 ) );
NAND2_X1 _u10_U5033  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16480 ) );
NAND2_X1 _u10_U5032  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16481 ) );
NAND2_X1 _u10_U5031  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16482 ) );
NAND4_X1 _u10_U5030  ( .A1(_u10_n16479 ), .A2(_u10_n16480 ), .A3(_u10_n16481 ), .A4(_u10_n16482 ), .ZN(_u10_n16463 ) );
NAND2_X1 _u10_U5029  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16475 ) );
NAND2_X1 _u10_U5028  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16476 ) );
NAND2_X1 _u10_U5027  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16477 ) );
NAND2_X1 _u10_U5026  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16478 ) );
NAND4_X1 _u10_U5025  ( .A1(_u10_n16475 ), .A2(_u10_n16476 ), .A3(_u10_n16477 ), .A4(_u10_n16478 ), .ZN(_u10_n16464 ) );
NAND2_X1 _u10_U5024  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16471 ) );
NAND2_X1 _u10_U5023  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16472 ) );
NAND2_X1 _u10_U5022  ( .A1(1'b0), .A2(_u10_n11757 ), .ZN(_u10_n16473 ) );
NAND2_X1 _u10_U5021  ( .A1(1'b0), .A2(_u10_n11733 ), .ZN(_u10_n16474 ) );
NAND4_X1 _u10_U5020  ( .A1(_u10_n16471 ), .A2(_u10_n16472 ), .A3(_u10_n16473 ), .A4(_u10_n16474 ), .ZN(_u10_n16465 ) );
NAND2_X1 _u10_U5019  ( .A1(1'b0), .A2(_u10_n11709 ), .ZN(_u10_n16467 ) );
NAND2_X1 _u10_U5018  ( .A1(1'b0), .A2(_u10_n11685 ), .ZN(_u10_n16468 ) );
NAND2_X1 _u10_U5017  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16469 ) );
NAND2_X1 _u10_U5016  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16470 ) );
NAND4_X1 _u10_U5015  ( .A1(_u10_n16467 ), .A2(_u10_n16468 ), .A3(_u10_n16469 ), .A4(_u10_n16470 ), .ZN(_u10_n16466 ) );
NOR4_X1 _u10_U5014  ( .A1(_u10_n16463 ), .A2(_u10_n16464 ), .A3(_u10_n16465 ), .A4(_u10_n16466 ), .ZN(_u10_n16462 ) );
NAND2_X1 _u10_U5013  ( .A1(_u10_n16461 ), .A2(_u10_n16462 ), .ZN(csr[7]) );
NAND2_X1 _u10_U5012  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16457 ) );
NAND2_X1 _u10_U5011  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16458 ) );
NAND2_X1 _u10_U5010  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16459 ) );
NAND2_X1 _u10_U5009  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16460 ) );
NAND4_X1 _u10_U5008  ( .A1(_u10_n16457 ), .A2(_u10_n16458 ), .A3(_u10_n16459 ), .A4(_u10_n16460 ), .ZN(_u10_n16442 ) );
NAND2_X1 _u10_U5007  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16453 ) );
NAND2_X1 _u10_U5006  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16454 ) );
NAND2_X1 _u10_U5005  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n16455 ) );
NAND2_X1 _u10_U5004  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16456 ) );
NAND4_X1 _u10_U5003  ( .A1(_u10_n16453 ), .A2(_u10_n16454 ), .A3(_u10_n16455 ), .A4(_u10_n16456 ), .ZN(_u10_n16443 ) );
NAND2_X1 _u10_U5002  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16449 ) );
NAND2_X1 _u10_U5001  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16450 ) );
NAND2_X1 _u10_U5000  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16451 ) );
NAND2_X1 _u10_U4999  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16452 ) );
NAND4_X1 _u10_U4998  ( .A1(_u10_n16449 ), .A2(_u10_n16450 ), .A3(_u10_n16451 ), .A4(_u10_n16452 ), .ZN(_u10_n16444 ) );
NAND2_X1 _u10_U4997  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16446 ) );
NAND2_X1 _u10_U4996  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16447 ) );
NAND2_X1 _u10_U4995  ( .A1(ch0_csr[8]), .A2(_u10_n12012 ), .ZN(_u10_n16448 ));
NAND3_X1 _u10_U4994  ( .A1(_u10_n16446 ), .A2(_u10_n16447 ), .A3(_u10_n16448 ), .ZN(_u10_n16445 ) );
NOR4_X1 _u10_U4993  ( .A1(_u10_n16442 ), .A2(_u10_n16443 ), .A3(_u10_n16444 ), .A4(_u10_n16445 ), .ZN(_u10_n16420 ) );
NAND2_X1 _u10_U4992  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16438 ) );
NAND2_X1 _u10_U4991  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16439 ) );
NAND2_X1 _u10_U4990  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16440 ) );
NAND2_X1 _u10_U4989  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16441 ) );
NAND4_X1 _u10_U4988  ( .A1(_u10_n16438 ), .A2(_u10_n16439 ), .A3(_u10_n16440 ), .A4(_u10_n16441 ), .ZN(_u10_n16422 ) );
NAND2_X1 _u10_U4987  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16434 ) );
NAND2_X1 _u10_U4986  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16435 ) );
NAND2_X1 _u10_U4985  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16436 ) );
NAND2_X1 _u10_U4984  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16437 ) );
NAND4_X1 _u10_U4983  ( .A1(_u10_n16434 ), .A2(_u10_n16435 ), .A3(_u10_n16436 ), .A4(_u10_n16437 ), .ZN(_u10_n16423 ) );
NAND2_X1 _u10_U4982  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16430 ) );
NAND2_X1 _u10_U4981  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16431 ) );
NAND2_X1 _u10_U4980  ( .A1(1'b0), .A2(_u10_n11754 ), .ZN(_u10_n16432 ) );
NAND2_X1 _u10_U4979  ( .A1(1'b0), .A2(_u10_n11730 ), .ZN(_u10_n16433 ) );
NAND4_X1 _u10_U4978  ( .A1(_u10_n16430 ), .A2(_u10_n16431 ), .A3(_u10_n16432 ), .A4(_u10_n16433 ), .ZN(_u10_n16424 ) );
NAND2_X1 _u10_U4977  ( .A1(1'b0), .A2(_u10_n11706 ), .ZN(_u10_n16426 ) );
NAND2_X1 _u10_U4976  ( .A1(1'b0), .A2(_u10_n11682 ), .ZN(_u10_n16427 ) );
NAND2_X1 _u10_U4975  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16428 ) );
NAND2_X1 _u10_U4974  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16429 ) );
NAND4_X1 _u10_U4973  ( .A1(_u10_n16426 ), .A2(_u10_n16427 ), .A3(_u10_n16428 ), .A4(_u10_n16429 ), .ZN(_u10_n16425 ) );
NOR4_X1 _u10_U4972  ( .A1(_u10_n16422 ), .A2(_u10_n16423 ), .A3(_u10_n16424 ), .A4(_u10_n16425 ), .ZN(_u10_n16421 ) );
NAND2_X1 _u10_U4971  ( .A1(_u10_n16420 ), .A2(_u10_n16421 ), .ZN(csr[8]) );
NAND2_X1 _u10_U4970  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16416 ) );
NAND2_X1 _u10_U4969  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16417 ) );
NAND2_X1 _u10_U4968  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16418 ) );
NAND2_X1 _u10_U4967  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16419 ) );
NAND4_X1 _u10_U4966  ( .A1(_u10_n16416 ), .A2(_u10_n16417 ), .A3(_u10_n16418 ), .A4(_u10_n16419 ), .ZN(_u10_n16401 ) );
NAND2_X1 _u10_U4965  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16412 ) );
NAND2_X1 _u10_U4964  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16413 ) );
NAND2_X1 _u10_U4963  ( .A1(1'b0), .A2(_u10_n12206 ), .ZN(_u10_n16414 ) );
NAND2_X1 _u10_U4962  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16415 ) );
NAND4_X1 _u10_U4961  ( .A1(_u10_n16412 ), .A2(_u10_n16413 ), .A3(_u10_n16414 ), .A4(_u10_n16415 ), .ZN(_u10_n16402 ) );
NAND2_X1 _u10_U4960  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16408 ) );
NAND2_X1 _u10_U4959  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16409 ) );
NAND2_X1 _u10_U4958  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16410 ) );
NAND2_X1 _u10_U4957  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16411 ) );
NAND4_X1 _u10_U4956  ( .A1(_u10_n16408 ), .A2(_u10_n16409 ), .A3(_u10_n16410 ), .A4(_u10_n16411 ), .ZN(_u10_n16403 ) );
NAND2_X1 _u10_U4955  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16405 ) );
NAND2_X1 _u10_U4954  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16406 ) );
NAND2_X1 _u10_U4953  ( .A1(1'b0), .A2(_u10_n12012 ), .ZN(_u10_n16407 ) );
NAND3_X1 _u10_U4952  ( .A1(_u10_n16405 ), .A2(_u10_n16406 ), .A3(_u10_n16407 ), .ZN(_u10_n16404 ) );
NOR4_X1 _u10_U4951  ( .A1(_u10_n16401 ), .A2(_u10_n16402 ), .A3(_u10_n16403 ), .A4(_u10_n16404 ), .ZN(_u10_n16379 ) );
NAND2_X1 _u10_U4950  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16397 ) );
NAND2_X1 _u10_U4949  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16398 ) );
NAND2_X1 _u10_U4948  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16399 ) );
NAND2_X1 _u10_U4947  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16400 ) );
NAND4_X1 _u10_U4946  ( .A1(_u10_n16397 ), .A2(_u10_n16398 ), .A3(_u10_n16399 ), .A4(_u10_n16400 ), .ZN(_u10_n16381 ) );
NAND2_X1 _u10_U4945  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16393 ) );
NAND2_X1 _u10_U4944  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16394 ) );
NAND2_X1 _u10_U4943  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16395 ) );
NAND2_X1 _u10_U4942  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16396 ) );
NAND4_X1 _u10_U4941  ( .A1(_u10_n16393 ), .A2(_u10_n16394 ), .A3(_u10_n16395 ), .A4(_u10_n16396 ), .ZN(_u10_n16382 ) );
NAND2_X1 _u10_U4940  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16389 ) );
NAND2_X1 _u10_U4939  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16390 ) );
NAND2_X1 _u10_U4938  ( .A1(1'b0), .A2(_u10_n11754 ), .ZN(_u10_n16391 ) );
NAND2_X1 _u10_U4937  ( .A1(1'b0), .A2(_u10_n11730 ), .ZN(_u10_n16392 ) );
NAND4_X1 _u10_U4936  ( .A1(_u10_n16389 ), .A2(_u10_n16390 ), .A3(_u10_n16391 ), .A4(_u10_n16392 ), .ZN(_u10_n16383 ) );
NAND2_X1 _u10_U4935  ( .A1(1'b0), .A2(_u10_n11706 ), .ZN(_u10_n16385 ) );
NAND2_X1 _u10_U4934  ( .A1(1'b0), .A2(_u10_n11682 ), .ZN(_u10_n16386 ) );
NAND2_X1 _u10_U4933  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16387 ) );
NAND2_X1 _u10_U4932  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16388 ) );
NAND4_X1 _u10_U4931  ( .A1(_u10_n16385 ), .A2(_u10_n16386 ), .A3(_u10_n16387 ), .A4(_u10_n16388 ), .ZN(_u10_n16384 ) );
NOR4_X1 _u10_U4930  ( .A1(_u10_n16381 ), .A2(_u10_n16382 ), .A3(_u10_n16383 ), .A4(_u10_n16384 ), .ZN(_u10_n16380 ) );
NAND2_X1 _u10_U4929  ( .A1(_u10_n16379 ), .A2(_u10_n16380 ), .ZN(csr[9]) );
NAND2_X1 _u10_U4928  ( .A1(_u10_n11552 ), .A2(_u10_n11551 ), .ZN(_u10_n16378 ) );
NAND2_X1 _u10_U4927  ( .A1(_u10_n11550 ), .A2(_u10_n16378 ), .ZN(de_start));
MUX2_X1 _u10_U4926  ( .A(_u10_n22999 ), .B(_u10_gnt_p0_d[4] ), .S(de_start),.Z(_u10_n10672 ) );
MUX2_X1 _u10_U4925  ( .A(_u10_n22998 ), .B(_u10_gnt_p0_d[3] ), .S(de_start),.Z(_u10_n10673 ) );
MUX2_X1 _u10_U4924  ( .A(_u10_n22997 ), .B(_u10_gnt_p0_d[2] ), .S(de_start),.Z(_u10_n10674 ) );
MUX2_X1 _u10_U4923  ( .A(_u10_n22996 ), .B(_u10_gnt_p0_d[1] ), .S(de_start),.Z(_u10_n10675 ) );
MUX2_X1 _u10_U4922  ( .A(_u10_n23000 ), .B(_u10_gnt_p0_d[0] ), .S(de_start),.Z(_u10_n10676 ) );
INV_X1 _u10_U4921  ( .A(_u10_n13702 ), .ZN(_u10_n24 ) );
NOR2_X1 _u10_U4920  ( .A1(_u10_n22990 ), .A2(_u10_n16377 ), .ZN(_u10_n16370 ) );
NOR2_X1 _u10_U4919  ( .A1(_u10_n22991 ), .A2(_u10_n16376 ), .ZN(_u10_n16371 ) );
NOR2_X1 _u10_U4918  ( .A1(_u10_n16375 ), .A2(_u10_n10664 ), .ZN(_u10_n16372 ) );
NOR2_X1 _u10_U4917  ( .A1(_u10_n16374 ), .A2(_u10_n10665 ), .ZN(_u10_n16373 ) );
NOR4_X1 _u10_U4916  ( .A1(_u10_n16370 ), .A2(_u10_n16371 ), .A3(_u10_n16372 ), .A4(_u10_n16373 ), .ZN(_u10_n16327 ) );
NOR2_X1 _u10_U4915  ( .A1(_u10_n16369 ), .A2(_u10_n11542 ), .ZN(_u10_n16362 ) );
NOR2_X1 _u10_U4914  ( .A1(_u10_n16368 ), .A2(_u10_n11543 ), .ZN(_u10_n16363 ) );
NOR2_X1 _u10_U4913  ( .A1(_u10_n22988 ), .A2(_u10_n16367 ), .ZN(_u10_n16364 ) );
NOR2_X1 _u10_U4912  ( .A1(_u10_n22989 ), .A2(_u10_n16366 ), .ZN(_u10_n16365 ) );
NOR4_X1 _u10_U4911  ( .A1(_u10_n16362 ), .A2(_u10_n16363 ), .A3(_u10_n16364 ), .A4(_u10_n16365 ), .ZN(_u10_n16328 ) );
NAND2_X1 _u10_U4910  ( .A1(_u10_n22992 ), .A2(_u10_n12152 ), .ZN(_u10_n16358 ) );
NAND2_X1 _u10_U4909  ( .A1(_u10_n22993 ), .A2(_u10_n12128 ), .ZN(_u10_n16359 ) );
NAND2_X1 _u10_U4908  ( .A1(_u10_n22994 ), .A2(_u10_n12104 ), .ZN(_u10_n16360 ) );
NAND2_X1 _u10_U4907  ( .A1(_u10_n22995 ), .A2(_u10_n12080 ), .ZN(_u10_n16361 ) );
NAND4_X1 _u10_U4906  ( .A1(_u10_n16358 ), .A2(_u10_n16359 ), .A3(_u10_n16360 ), .A4(_u10_n16361 ), .ZN(_u10_n16351 ) );
NOR2_X1 _u10_U4905  ( .A1(_u10_n16357 ), .A2(_u10_n11539 ), .ZN(_u10_n16352 ) );
NOR2_X1 _u10_U4904  ( .A1(_u10_n16356 ), .A2(_u10_n10662 ), .ZN(_u10_n16353 ) );
NOR2_X1 _u10_U4903  ( .A1(_u10_n16355 ), .A2(_u10_n10663 ), .ZN(_u10_n16354 ) );
NOR4_X1 _u10_U4902  ( .A1(_u10_n16351 ), .A2(_u10_n16352 ), .A3(_u10_n16353 ), .A4(_u10_n16354 ), .ZN(_u10_n16329 ) );
NAND2_X1 _u10_U4901  ( .A1(_u10_n11976 ), .A2(_u10_ndr_r[15]), .ZN(_u10_n16347 ) );
NAND2_X1 _u10_U4900  ( .A1(_u10_n11952 ), .A2(_u10_ndr_r[16]), .ZN(_u10_n16348 ) );
NAND2_X1 _u10_U4899  ( .A1(_u10_n11928 ), .A2(_u10_ndr_r[17]), .ZN(_u10_n16349 ) );
NAND2_X1 _u10_U4898  ( .A1(_u10_n11904 ), .A2(_u10_ndr_r[18]), .ZN(_u10_n16350 ) );
NAND4_X1 _u10_U4897  ( .A1(_u10_n16347 ), .A2(_u10_n16348 ), .A3(_u10_n16349 ), .A4(_u10_n16350 ), .ZN(_u10_n16331 ) );
NAND2_X1 _u10_U4896  ( .A1(_u10_n11880 ), .A2(_u10_ndr_r[19]), .ZN(_u10_n16343 ) );
NAND2_X1 _u10_U4895  ( .A1(_u10_n11856 ), .A2(_u10_ndr_r[20]), .ZN(_u10_n16344 ) );
NAND2_X1 _u10_U4894  ( .A1(_u10_n11832 ), .A2(_u10_ndr_r[21]), .ZN(_u10_n16345 ) );
NAND2_X1 _u10_U4893  ( .A1(_u10_n11808 ), .A2(_u10_ndr_r[22]), .ZN(_u10_n16346 ) );
NAND4_X1 _u10_U4892  ( .A1(_u10_n16343 ), .A2(_u10_n16344 ), .A3(_u10_n16345 ), .A4(_u10_n16346 ), .ZN(_u10_n16332 ) );
NAND2_X1 _u10_U4891  ( .A1(_u10_n11784 ), .A2(_u10_ndr_r[23]), .ZN(_u10_n16339 ) );
NAND2_X1 _u10_U4890  ( .A1(_u10_n11760 ), .A2(_u10_ndr_r[24]), .ZN(_u10_n16340 ) );
NAND2_X1 _u10_U4889  ( .A1(_u10_n12378 ), .A2(_u10_ndr_r[25]), .ZN(_u10_n16341 ) );
NAND2_X1 _u10_U4888  ( .A1(_u10_n12377 ), .A2(_u10_ndr_r[26]), .ZN(_u10_n16342 ) );
NAND4_X1 _u10_U4887  ( .A1(_u10_n16339 ), .A2(_u10_n16340 ), .A3(_u10_n16341 ), .A4(_u10_n16342 ), .ZN(_u10_n16333 ) );
NAND2_X1 _u10_U4886  ( .A1(_u10_n12372 ), .A2(_u10_ndr_r[27]), .ZN(_u10_n16335 ) );
NAND2_X1 _u10_U4885  ( .A1(_u10_n12371 ), .A2(_u10_ndr_r[28]), .ZN(_u10_n16336 ) );
NAND2_X1 _u10_U4884  ( .A1(_u10_n11640 ), .A2(_u10_ndr_r[29]), .ZN(_u10_n16337 ) );
NAND2_X1 _u10_U4883  ( .A1(_u10_n11616 ), .A2(_u10_ndr_r[30]), .ZN(_u10_n16338 ) );
NAND4_X1 _u10_U4882  ( .A1(_u10_n16335 ), .A2(_u10_n16336 ), .A3(_u10_n16337 ), .A4(_u10_n16338 ), .ZN(_u10_n16334 ) );
NOR4_X1 _u10_U4881  ( .A1(_u10_n16331 ), .A2(_u10_n16332 ), .A3(_u10_n16333 ), .A4(_u10_n16334 ), .ZN(_u10_n16330 ) );
NAND4_X1 _u10_U4880  ( .A1(_u10_n16327 ), .A2(_u10_n16328 ), .A3(_u10_n16329 ), .A4(_u10_n16330 ), .ZN(ndr) );
NAND2_X1 _u10_U4879  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16323 ) );
NAND2_X1 _u10_U4878  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16324 ) );
NAND2_X1 _u10_U4877  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16325 ) );
NAND2_X1 _u10_U4876  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16326 ) );
NAND4_X1 _u10_U4875  ( .A1(_u10_n16323 ), .A2(_u10_n16324 ), .A3(_u10_n16325 ), .A4(_u10_n16326 ), .ZN(_u10_n16308 ) );
NAND2_X1 _u10_U4874  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16319 ) );
NAND2_X1 _u10_U4873  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16320 ) );
NAND2_X1 _u10_U4872  ( .A1(1'b0), .A2(_u10_n12209 ), .ZN(_u10_n16321 ) );
NAND2_X1 _u10_U4871  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16322 ) );
NAND4_X1 _u10_U4870  ( .A1(_u10_n16319 ), .A2(_u10_n16320 ), .A3(_u10_n16321 ), .A4(_u10_n16322 ), .ZN(_u10_n16309 ) );
NAND2_X1 _u10_U4869  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16315 ) );
NAND2_X1 _u10_U4868  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16316 ) );
NAND2_X1 _u10_U4867  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16317 ) );
NAND2_X1 _u10_U4866  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16318 ) );
NAND4_X1 _u10_U4865  ( .A1(_u10_n16315 ), .A2(_u10_n16316 ), .A3(_u10_n16317 ), .A4(_u10_n16318 ), .ZN(_u10_n16310 ) );
NAND2_X1 _u10_U4864  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16312 ) );
NAND2_X1 _u10_U4863  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16313 ) );
NAND2_X1 _u10_U4862  ( .A1(1'b0), .A2(_u10_n12012 ), .ZN(_u10_n16314 ) );
NAND3_X1 _u10_U4861  ( .A1(_u10_n16312 ), .A2(_u10_n16313 ), .A3(_u10_n16314 ), .ZN(_u10_n16311 ) );
NOR4_X1 _u10_U4860  ( .A1(_u10_n16308 ), .A2(_u10_n16309 ), .A3(_u10_n16310 ), .A4(_u10_n16311 ), .ZN(_u10_n16286 ) );
NAND2_X1 _u10_U4859  ( .A1(1'b0), .A2(_u10_n11978 ), .ZN(_u10_n16304 ) );
NAND2_X1 _u10_U4858  ( .A1(1'b0), .A2(_u10_n11954 ), .ZN(_u10_n16305 ) );
NAND2_X1 _u10_U4857  ( .A1(1'b0), .A2(_u10_n11930 ), .ZN(_u10_n16306 ) );
NAND2_X1 _u10_U4856  ( .A1(1'b0), .A2(_u10_n11906 ), .ZN(_u10_n16307 ) );
NAND4_X1 _u10_U4855  ( .A1(_u10_n16304 ), .A2(_u10_n16305 ), .A3(_u10_n16306 ), .A4(_u10_n16307 ), .ZN(_u10_n16288 ) );
NAND2_X1 _u10_U4854  ( .A1(1'b0), .A2(_u10_n11882 ), .ZN(_u10_n16300 ) );
NAND2_X1 _u10_U4853  ( .A1(1'b0), .A2(_u10_n11858 ), .ZN(_u10_n16301 ) );
NAND2_X1 _u10_U4852  ( .A1(1'b0), .A2(_u10_n11834 ), .ZN(_u10_n16302 ) );
NAND2_X1 _u10_U4851  ( .A1(1'b0), .A2(_u10_n11810 ), .ZN(_u10_n16303 ) );
NAND4_X1 _u10_U4850  ( .A1(_u10_n16300 ), .A2(_u10_n16301 ), .A3(_u10_n16302 ), .A4(_u10_n16303 ), .ZN(_u10_n16289 ) );
NAND2_X1 _u10_U4849  ( .A1(1'b0), .A2(_u10_n11786 ), .ZN(_u10_n16296 ) );
NAND2_X1 _u10_U4848  ( .A1(1'b0), .A2(_u10_n11762 ), .ZN(_u10_n16297 ) );
NAND2_X1 _u10_U4847  ( .A1(1'b0), .A2(_u10_n11755 ), .ZN(_u10_n16298 ) );
NAND2_X1 _u10_U4846  ( .A1(1'b0), .A2(_u10_n11731 ), .ZN(_u10_n16299 ) );
NAND4_X1 _u10_U4845  ( .A1(_u10_n16296 ), .A2(_u10_n16297 ), .A3(_u10_n16298 ), .A4(_u10_n16299 ), .ZN(_u10_n16290 ) );
NAND2_X1 _u10_U4844  ( .A1(1'b0), .A2(_u10_n11707 ), .ZN(_u10_n16292 ) );
NAND2_X1 _u10_U4843  ( .A1(1'b0), .A2(_u10_n11683 ), .ZN(_u10_n16293 ) );
NAND2_X1 _u10_U4842  ( .A1(1'b0), .A2(_u10_n11642 ), .ZN(_u10_n16294 ) );
NAND2_X1 _u10_U4841  ( .A1(1'b0), .A2(_u10_n11618 ), .ZN(_u10_n16295 ) );
NAND4_X1 _u10_U4840  ( .A1(_u10_n16292 ), .A2(_u10_n16293 ), .A3(_u10_n16294 ), .A4(_u10_n16295 ), .ZN(_u10_n16291 ) );
NOR4_X1 _u10_U4839  ( .A1(_u10_n16288 ), .A2(_u10_n16289 ), .A3(_u10_n16290 ), .A4(_u10_n16291 ), .ZN(_u10_n16287 ) );
NAND2_X1 _u10_U4838  ( .A1(_u10_n16286 ), .A2(_u10_n16287 ), .ZN(pointer[0]));
NAND2_X1 _u10_U4837  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16282 ) );
NAND2_X1 _u10_U4836  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16283 ) );
NAND2_X1 _u10_U4835  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16284 ) );
NAND2_X1 _u10_U4834  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16285 ) );
NAND4_X1 _u10_U4833  ( .A1(_u10_n16282 ), .A2(_u10_n16283 ), .A3(_u10_n16284 ), .A4(_u10_n16285 ), .ZN(_u10_n16267 ) );
NAND2_X1 _u10_U4832  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16278 ) );
NAND2_X1 _u10_U4831  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16279 ) );
NAND2_X1 _u10_U4830  ( .A1(1'b0), .A2(_u10_n12211 ), .ZN(_u10_n16280 ) );
NAND2_X1 _u10_U4829  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16281 ) );
NAND4_X1 _u10_U4828  ( .A1(_u10_n16278 ), .A2(_u10_n16279 ), .A3(_u10_n16280 ), .A4(_u10_n16281 ), .ZN(_u10_n16268 ) );
NAND2_X1 _u10_U4827  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16274 ) );
NAND2_X1 _u10_U4826  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16275 ) );
NAND2_X1 _u10_U4825  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16276 ) );
NAND2_X1 _u10_U4824  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16277 ) );
NAND4_X1 _u10_U4823  ( .A1(_u10_n16274 ), .A2(_u10_n16275 ), .A3(_u10_n16276 ), .A4(_u10_n16277 ), .ZN(_u10_n16269 ) );
NAND2_X1 _u10_U4822  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16271 ) );
NAND2_X1 _u10_U4821  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16272 ) );
NAND2_X1 _u10_U4820  ( .A1(1'b0), .A2(_u10_n12012 ), .ZN(_u10_n16273 ) );
NAND3_X1 _u10_U4819  ( .A1(_u10_n16271 ), .A2(_u10_n16272 ), .A3(_u10_n16273 ), .ZN(_u10_n16270 ) );
NOR4_X1 _u10_U4818  ( .A1(_u10_n16267 ), .A2(_u10_n16268 ), .A3(_u10_n16269 ), .A4(_u10_n16270 ), .ZN(_u10_n16245 ) );
NAND2_X1 _u10_U4817  ( .A1(1'b0), .A2(_u10_n11997 ), .ZN(_u10_n16263 ) );
NAND2_X1 _u10_U4816  ( .A1(1'b0), .A2(_u10_n11971 ), .ZN(_u10_n16264 ) );
NAND2_X1 _u10_U4815  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n16265 ) );
NAND2_X1 _u10_U4814  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n16266 ) );
NAND4_X1 _u10_U4813  ( .A1(_u10_n16263 ), .A2(_u10_n16264 ), .A3(_u10_n16265 ), .A4(_u10_n16266 ), .ZN(_u10_n16247 ) );
NAND2_X1 _u10_U4812  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n16259 ) );
NAND2_X1 _u10_U4811  ( .A1(1'b0), .A2(_u10_n11877 ), .ZN(_u10_n16260 ) );
NAND2_X1 _u10_U4810  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n16261 ) );
NAND2_X1 _u10_U4809  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n16262 ) );
NAND4_X1 _u10_U4808  ( .A1(_u10_n16259 ), .A2(_u10_n16260 ), .A3(_u10_n16261 ), .A4(_u10_n16262 ), .ZN(_u10_n16248 ) );
NAND2_X1 _u10_U4807  ( .A1(1'b0), .A2(_u10_n11805 ), .ZN(_u10_n16255 ) );
NAND2_X1 _u10_U4806  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n16256 ) );
NAND2_X1 _u10_U4805  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n16257 ) );
NAND2_X1 _u10_U4804  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n16258 ) );
NAND4_X1 _u10_U4803  ( .A1(_u10_n16255 ), .A2(_u10_n16256 ), .A3(_u10_n16257 ), .A4(_u10_n16258 ), .ZN(_u10_n16249 ) );
NAND2_X1 _u10_U4802  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n16251 ) );
NAND2_X1 _u10_U4801  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n16252 ) );
NAND2_X1 _u10_U4800  ( .A1(1'b0), .A2(_u10_n11662 ), .ZN(_u10_n16253 ) );
NAND2_X1 _u10_U4799  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n16254 ) );
NAND4_X1 _u10_U4798  ( .A1(_u10_n16251 ), .A2(_u10_n16252 ), .A3(_u10_n16253 ), .A4(_u10_n16254 ), .ZN(_u10_n16250 ) );
NOR4_X1 _u10_U4797  ( .A1(_u10_n16247 ), .A2(_u10_n16248 ), .A3(_u10_n16249 ), .A4(_u10_n16250 ), .ZN(_u10_n16246 ) );
NAND2_X1 _u10_U4796  ( .A1(_u10_n16245 ), .A2(_u10_n16246 ), .ZN(pointer[10]) );
NAND2_X1 _u10_U4795  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16241 ) );
NAND2_X1 _u10_U4794  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16242 ) );
NAND2_X1 _u10_U4793  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16243 ) );
NAND2_X1 _u10_U4792  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16244 ) );
NAND4_X1 _u10_U4791  ( .A1(_u10_n16241 ), .A2(_u10_n16242 ), .A3(_u10_n16243 ), .A4(_u10_n16244 ), .ZN(_u10_n16226 ) );
NAND2_X1 _u10_U4790  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16237 ) );
NAND2_X1 _u10_U4789  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16238 ) );
NAND2_X1 _u10_U4788  ( .A1(1'b0), .A2(_u10_n12210 ), .ZN(_u10_n16239 ) );
NAND2_X1 _u10_U4787  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16240 ) );
NAND4_X1 _u10_U4786  ( .A1(_u10_n16237 ), .A2(_u10_n16238 ), .A3(_u10_n16239 ), .A4(_u10_n16240 ), .ZN(_u10_n16227 ) );
NAND2_X1 _u10_U4785  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16233 ) );
NAND2_X1 _u10_U4784  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16234 ) );
NAND2_X1 _u10_U4783  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16235 ) );
NAND2_X1 _u10_U4782  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16236 ) );
NAND4_X1 _u10_U4781  ( .A1(_u10_n16233 ), .A2(_u10_n16234 ), .A3(_u10_n16235 ), .A4(_u10_n16236 ), .ZN(_u10_n16228 ) );
NAND2_X1 _u10_U4780  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16230 ) );
NAND2_X1 _u10_U4779  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16231 ) );
NAND2_X1 _u10_U4778  ( .A1(1'b0), .A2(_u10_n12012 ), .ZN(_u10_n16232 ) );
NAND3_X1 _u10_U4777  ( .A1(_u10_n16230 ), .A2(_u10_n16231 ), .A3(_u10_n16232 ), .ZN(_u10_n16229 ) );
NOR4_X1 _u10_U4776  ( .A1(_u10_n16226 ), .A2(_u10_n16227 ), .A3(_u10_n16228 ), .A4(_u10_n16229 ), .ZN(_u10_n16204 ) );
NAND2_X1 _u10_U4775  ( .A1(1'b0), .A2(_u10_n11998 ), .ZN(_u10_n16222 ) );
NAND2_X1 _u10_U4774  ( .A1(1'b0), .A2(_u10_n11970 ), .ZN(_u10_n16223 ) );
NAND2_X1 _u10_U4773  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n16224 ) );
NAND2_X1 _u10_U4772  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n16225 ) );
NAND4_X1 _u10_U4771  ( .A1(_u10_n16222 ), .A2(_u10_n16223 ), .A3(_u10_n16224 ), .A4(_u10_n16225 ), .ZN(_u10_n16206 ) );
NAND2_X1 _u10_U4770  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n16218 ) );
NAND2_X1 _u10_U4769  ( .A1(1'b0), .A2(_u10_n11878 ), .ZN(_u10_n16219 ) );
NAND2_X1 _u10_U4768  ( .A1(1'b0), .A2(_u10_n11850 ), .ZN(_u10_n16220 ) );
NAND2_X1 _u10_U4767  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n16221 ) );
NAND4_X1 _u10_U4766  ( .A1(_u10_n16218 ), .A2(_u10_n16219 ), .A3(_u10_n16220 ), .A4(_u10_n16221 ), .ZN(_u10_n16207 ) );
NAND2_X1 _u10_U4765  ( .A1(1'b0), .A2(_u10_n11806 ), .ZN(_u10_n16214 ) );
NAND2_X1 _u10_U4764  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n16215 ) );
NAND2_X1 _u10_U4763  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n16216 ) );
NAND2_X1 _u10_U4762  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n16217 ) );
NAND4_X1 _u10_U4761  ( .A1(_u10_n16214 ), .A2(_u10_n16215 ), .A3(_u10_n16216 ), .A4(_u10_n16217 ), .ZN(_u10_n16208 ) );
NAND2_X1 _u10_U4760  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n16210 ) );
NAND2_X1 _u10_U4759  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n16211 ) );
NAND2_X1 _u10_U4758  ( .A1(1'b0), .A2(_u10_n11658 ), .ZN(_u10_n16212 ) );
NAND2_X1 _u10_U4757  ( .A1(1'b0), .A2(_u10_n11634 ), .ZN(_u10_n16213 ) );
NAND4_X1 _u10_U4756  ( .A1(_u10_n16210 ), .A2(_u10_n16211 ), .A3(_u10_n16212 ), .A4(_u10_n16213 ), .ZN(_u10_n16209 ) );
NOR4_X1 _u10_U4755  ( .A1(_u10_n16206 ), .A2(_u10_n16207 ), .A3(_u10_n16208 ), .A4(_u10_n16209 ), .ZN(_u10_n16205 ) );
NAND2_X1 _u10_U4754  ( .A1(_u10_n16204 ), .A2(_u10_n16205 ), .ZN(pointer[11]) );
NAND2_X1 _u10_U4753  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16200 ) );
NAND2_X1 _u10_U4752  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16201 ) );
NAND2_X1 _u10_U4751  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16202 ) );
NAND2_X1 _u10_U4750  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16203 ) );
NAND4_X1 _u10_U4749  ( .A1(_u10_n16200 ), .A2(_u10_n16201 ), .A3(_u10_n16202 ), .A4(_u10_n16203 ), .ZN(_u10_n16185 ) );
NAND2_X1 _u10_U4748  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16196 ) );
NAND2_X1 _u10_U4747  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16197 ) );
NAND2_X1 _u10_U4746  ( .A1(1'b0), .A2(_u10_n12207 ), .ZN(_u10_n16198 ) );
NAND2_X1 _u10_U4745  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16199 ) );
NAND4_X1 _u10_U4744  ( .A1(_u10_n16196 ), .A2(_u10_n16197 ), .A3(_u10_n16198 ), .A4(_u10_n16199 ), .ZN(_u10_n16186 ) );
NAND2_X1 _u10_U4743  ( .A1(1'b0), .A2(_u10_n12152 ), .ZN(_u10_n16192 ) );
NAND2_X1 _u10_U4742  ( .A1(1'b0), .A2(_u10_n12128 ), .ZN(_u10_n16193 ) );
NAND2_X1 _u10_U4741  ( .A1(1'b0), .A2(_u10_n12104 ), .ZN(_u10_n16194 ) );
NAND2_X1 _u10_U4740  ( .A1(1'b0), .A2(_u10_n12080 ), .ZN(_u10_n16195 ) );
NAND4_X1 _u10_U4739  ( .A1(_u10_n16192 ), .A2(_u10_n16193 ), .A3(_u10_n16194 ), .A4(_u10_n16195 ), .ZN(_u10_n16187 ) );
NAND2_X1 _u10_U4738  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16189 ) );
NAND2_X1 _u10_U4737  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16190 ) );
NAND2_X1 _u10_U4736  ( .A1(1'b0), .A2(_u10_n12012 ), .ZN(_u10_n16191 ) );
NAND3_X1 _u10_U4735  ( .A1(_u10_n16189 ), .A2(_u10_n16190 ), .A3(_u10_n16191 ), .ZN(_u10_n16188 ) );
NOR4_X1 _u10_U4734  ( .A1(_u10_n16185 ), .A2(_u10_n16186 ), .A3(_u10_n16187 ), .A4(_u10_n16188 ), .ZN(_u10_n16163 ) );
NAND2_X1 _u10_U4733  ( .A1(1'b0), .A2(_u10_n11994 ), .ZN(_u10_n16181 ) );
NAND2_X1 _u10_U4732  ( .A1(1'b0), .A2(_u10_n11974 ), .ZN(_u10_n16182 ) );
NAND2_X1 _u10_U4731  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n16183 ) );
NAND2_X1 _u10_U4730  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n16184 ) );
NAND4_X1 _u10_U4729  ( .A1(_u10_n16181 ), .A2(_u10_n16182 ), .A3(_u10_n16183 ), .A4(_u10_n16184 ), .ZN(_u10_n16165 ) );
NAND2_X1 _u10_U4728  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n16177 ) );
NAND2_X1 _u10_U4727  ( .A1(1'b0), .A2(_u10_n11874 ), .ZN(_u10_n16178 ) );
NAND2_X1 _u10_U4726  ( .A1(1'b0), .A2(_u10_n11851 ), .ZN(_u10_n16179 ) );
NAND2_X1 _u10_U4725  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n16180 ) );
NAND4_X1 _u10_U4724  ( .A1(_u10_n16177 ), .A2(_u10_n16178 ), .A3(_u10_n16179 ), .A4(_u10_n16180 ), .ZN(_u10_n16166 ) );
NAND2_X1 _u10_U4723  ( .A1(1'b0), .A2(_u10_n11802 ), .ZN(_u10_n16173 ) );
NAND2_X1 _u10_U4722  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n16174 ) );
NAND2_X1 _u10_U4721  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n16175 ) );
NAND2_X1 _u10_U4720  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n16176 ) );
NAND4_X1 _u10_U4719  ( .A1(_u10_n16173 ), .A2(_u10_n16174 ), .A3(_u10_n16175 ), .A4(_u10_n16176 ), .ZN(_u10_n16167 ) );
NAND2_X1 _u10_U4718  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n16169 ) );
NAND2_X1 _u10_U4717  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n16170 ) );
NAND2_X1 _u10_U4716  ( .A1(1'b0), .A2(_u10_n11659 ), .ZN(_u10_n16171 ) );
NAND2_X1 _u10_U4715  ( .A1(1'b0), .A2(_u10_n11635 ), .ZN(_u10_n16172 ) );
NAND4_X1 _u10_U4714  ( .A1(_u10_n16169 ), .A2(_u10_n16170 ), .A3(_u10_n16171 ), .A4(_u10_n16172 ), .ZN(_u10_n16168 ) );
NOR4_X1 _u10_U4713  ( .A1(_u10_n16165 ), .A2(_u10_n16166 ), .A3(_u10_n16167 ), .A4(_u10_n16168 ), .ZN(_u10_n16164 ) );
NAND2_X1 _u10_U4712  ( .A1(_u10_n16163 ), .A2(_u10_n16164 ), .ZN(pointer[12]) );
NAND2_X1 _u10_U4711  ( .A1(1'b0), .A2(_u10_n12343 ), .ZN(_u10_n16159 ) );
NAND2_X1 _u10_U4710  ( .A1(1'b0), .A2(_u10_n12319 ), .ZN(_u10_n16160 ) );
NAND2_X1 _u10_U4709  ( .A1(1'b0), .A2(_u10_n12296 ), .ZN(_u10_n16161 ) );
NAND2_X1 _u10_U4708  ( .A1(1'b0), .A2(_u10_n12272 ), .ZN(_u10_n16162 ) );
NAND4_X1 _u10_U4707  ( .A1(_u10_n16159 ), .A2(_u10_n16160 ), .A3(_u10_n16161 ), .A4(_u10_n16162 ), .ZN(_u10_n16144 ) );
NAND2_X1 _u10_U4706  ( .A1(1'b0), .A2(_u10_n12247 ), .ZN(_u10_n16155 ) );
NAND2_X1 _u10_U4705  ( .A1(1'b0), .A2(_u10_n12223 ), .ZN(_u10_n16156 ) );
NAND2_X1 _u10_U4704  ( .A1(1'b0), .A2(_u10_n12208 ), .ZN(_u10_n16157 ) );
NAND2_X1 _u10_U4703  ( .A1(1'b0), .A2(_u10_n12175 ), .ZN(_u10_n16158 ) );
NAND4_X1 _u10_U4702  ( .A1(_u10_n16155 ), .A2(_u10_n16156 ), .A3(_u10_n16157 ), .A4(_u10_n16158 ), .ZN(_u10_n16145 ) );
NAND2_X1 _u10_U4701  ( .A1(1'b0), .A2(_u10_n12162 ), .ZN(_u10_n16151 ) );
NAND2_X1 _u10_U4700  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n16152 ) );
NAND2_X1 _u10_U4699  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n16153 ) );
NAND2_X1 _u10_U4698  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n16154 ) );
NAND4_X1 _u10_U4697  ( .A1(_u10_n16151 ), .A2(_u10_n16152 ), .A3(_u10_n16153 ), .A4(_u10_n16154 ), .ZN(_u10_n16146 ) );
NAND2_X1 _u10_U4696  ( .A1(1'b0), .A2(_u10_n12056 ), .ZN(_u10_n16148 ) );
NAND2_X1 _u10_U4695  ( .A1(1'b0), .A2(_u10_n12032 ), .ZN(_u10_n16149 ) );
NAND2_X1 _u10_U4694  ( .A1(1'b0), .A2(_u10_n12012 ), .ZN(_u10_n16150 ) );
NAND3_X1 _u10_U4693  ( .A1(_u10_n16148 ), .A2(_u10_n16149 ), .A3(_u10_n16150 ), .ZN(_u10_n16147 ) );
NOR4_X1 _u10_U4692  ( .A1(_u10_n16144 ), .A2(_u10_n16145 ), .A3(_u10_n16146 ), .A4(_u10_n16147 ), .ZN(_u10_n16122 ) );
NAND2_X1 _u10_U4691  ( .A1(1'b0), .A2(_u10_n11995 ), .ZN(_u10_n16140 ) );
NAND2_X1 _u10_U4690  ( .A1(1'b0), .A2(_u10_n12395 ), .ZN(_u10_n16141 ) );
NAND2_X1 _u10_U4689  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n16142 ) );
NAND2_X1 _u10_U4688  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n16143 ) );
NAND4_X1 _u10_U4687  ( .A1(_u10_n16140 ), .A2(_u10_n16141 ), .A3(_u10_n16142 ), .A4(_u10_n16143 ), .ZN(_u10_n16124 ) );
NAND2_X1 _u10_U4686  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n16136 ) );
NAND2_X1 _u10_U4685  ( .A1(1'b0), .A2(_u10_n11875 ), .ZN(_u10_n16137 ) );
NAND2_X1 _u10_U4684  ( .A1(1'b0), .A2(_u10_n11855 ), .ZN(_u10_n16138 ) );
NAND2_X1 _u10_U4683  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n16139 ) );
NAND4_X1 _u10_U4682  ( .A1(_u10_n16136 ), .A2(_u10_n16137 ), .A3(_u10_n16138 ), .A4(_u10_n16139 ), .ZN(_u10_n16125 ) );
NAND2_X1 _u10_U4681  ( .A1(1'b0), .A2(_u10_n11803 ), .ZN(_u10_n16132 ) );
NAND2_X1 _u10_U4680  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n16133 ) );
NAND2_X1 _u10_U4679  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n16134 ) );
NAND2_X1 _u10_U4678  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n16135 ) );
NAND4_X1 _u10_U4677  ( .A1(_u10_n16132 ), .A2(_u10_n16133 ), .A3(_u10_n16134 ), .A4(_u10_n16135 ), .ZN(_u10_n16126 ) );
NAND2_X1 _u10_U4676  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n16128 ) );
NAND2_X1 _u10_U4675  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n16129 ) );
NAND2_X1 _u10_U4674  ( .A1(1'b0), .A2(_u10_n11663 ), .ZN(_u10_n16130 ) );
NAND2_X1 _u10_U4673  ( .A1(1'b0), .A2(_u10_n11639 ), .ZN(_u10_n16131 ) );
NAND4_X1 _u10_U4672  ( .A1(_u10_n16128 ), .A2(_u10_n16129 ), .A3(_u10_n16130 ), .A4(_u10_n16131 ), .ZN(_u10_n16127 ) );
NOR4_X1 _u10_U4671  ( .A1(_u10_n16124 ), .A2(_u10_n16125 ), .A3(_u10_n16126 ), .A4(_u10_n16127 ), .ZN(_u10_n16123 ) );
NAND2_X1 _u10_U4670  ( .A1(_u10_n16122 ), .A2(_u10_n16123 ), .ZN(pointer[13]) );
NAND2_X1 _u10_U4669  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n16118 ) );
NAND2_X1 _u10_U4668  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n16119 ) );
NAND2_X1 _u10_U4667  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n16120 ) );
NAND2_X1 _u10_U4666  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n16121 ) );
NAND4_X1 _u10_U4665  ( .A1(_u10_n16118 ), .A2(_u10_n16119 ), .A3(_u10_n16120 ), .A4(_u10_n16121 ), .ZN(_u10_n16103 ) );
NAND2_X1 _u10_U4664  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n16114 ) );
NAND2_X1 _u10_U4663  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n16115 ) );
NAND2_X1 _u10_U4662  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n16116 ) );
NAND2_X1 _u10_U4661  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n16117 ) );
NAND4_X1 _u10_U4660  ( .A1(_u10_n16114 ), .A2(_u10_n16115 ), .A3(_u10_n16116 ), .A4(_u10_n16117 ), .ZN(_u10_n16104 ) );
NAND2_X1 _u10_U4659  ( .A1(1'b0), .A2(_u10_n12159 ), .ZN(_u10_n16110 ) );
NAND2_X1 _u10_U4658  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n16111 ) );
NAND2_X1 _u10_U4657  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n16112 ) );
NAND2_X1 _u10_U4656  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n16113 ) );
NAND4_X1 _u10_U4655  ( .A1(_u10_n16110 ), .A2(_u10_n16111 ), .A3(_u10_n16112 ), .A4(_u10_n16113 ), .ZN(_u10_n16105 ) );
NAND2_X1 _u10_U4654  ( .A1(1'b0), .A2(_u10_n12067 ), .ZN(_u10_n16107 ) );
NAND2_X1 _u10_U4653  ( .A1(1'b0), .A2(_u10_n12043 ), .ZN(_u10_n16108 ) );
NAND2_X1 _u10_U4652  ( .A1(1'b0), .A2(_u10_n12012 ), .ZN(_u10_n16109 ) );
NAND3_X1 _u10_U4651  ( .A1(_u10_n16107 ), .A2(_u10_n16108 ), .A3(_u10_n16109 ), .ZN(_u10_n16106 ) );
NOR4_X1 _u10_U4650  ( .A1(_u10_n16103 ), .A2(_u10_n16104 ), .A3(_u10_n16105 ), .A4(_u10_n16106 ), .ZN(_u10_n16081 ) );
NAND2_X1 _u10_U4649  ( .A1(1'b0), .A2(_u10_n12396 ), .ZN(_u10_n16099 ) );
NAND2_X1 _u10_U4648  ( .A1(1'b0), .A2(_u10_n11969 ), .ZN(_u10_n16100 ) );
NAND2_X1 _u10_U4647  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n16101 ) );
NAND2_X1 _u10_U4646  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n16102 ) );
NAND4_X1 _u10_U4645  ( .A1(_u10_n16099 ), .A2(_u10_n16100 ), .A3(_u10_n16101 ), .A4(_u10_n16102 ), .ZN(_u10_n16083 ) );
NAND2_X1 _u10_U4644  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n16095 ) );
NAND2_X1 _u10_U4643  ( .A1(1'b0), .A2(_u10_n12387 ), .ZN(_u10_n16096 ) );
NAND2_X1 _u10_U4642  ( .A1(1'b0), .A2(_u10_n12386 ), .ZN(_u10_n16097 ) );
NAND2_X1 _u10_U4641  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n16098 ) );
NAND4_X1 _u10_U4640  ( .A1(_u10_n16095 ), .A2(_u10_n16096 ), .A3(_u10_n16097 ), .A4(_u10_n16098 ), .ZN(_u10_n16084 ) );
NAND2_X1 _u10_U4639  ( .A1(1'b0), .A2(_u10_n12380 ), .ZN(_u10_n16091 ) );
NAND2_X1 _u10_U4638  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n16092 ) );
NAND2_X1 _u10_U4637  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n16093 ) );
NAND2_X1 _u10_U4636  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n16094 ) );
NAND4_X1 _u10_U4635  ( .A1(_u10_n16091 ), .A2(_u10_n16092 ), .A3(_u10_n16093 ), .A4(_u10_n16094 ), .ZN(_u10_n16085 ) );
NAND2_X1 _u10_U4634  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n16087 ) );
NAND2_X1 _u10_U4633  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n16088 ) );
NAND2_X1 _u10_U4632  ( .A1(1'b0), .A2(_u10_n12370 ), .ZN(_u10_n16089 ) );
NAND2_X1 _u10_U4631  ( .A1(1'b0), .A2(_u10_n12369 ), .ZN(_u10_n16090 ) );
NAND4_X1 _u10_U4630  ( .A1(_u10_n16087 ), .A2(_u10_n16088 ), .A3(_u10_n16089 ), .A4(_u10_n16090 ), .ZN(_u10_n16086 ) );
NOR4_X1 _u10_U4629  ( .A1(_u10_n16083 ), .A2(_u10_n16084 ), .A3(_u10_n16085 ), .A4(_u10_n16086 ), .ZN(_u10_n16082 ) );
NAND2_X1 _u10_U4628  ( .A1(_u10_n16081 ), .A2(_u10_n16082 ), .ZN(pointer[14]) );
NAND2_X1 _u10_U4627  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n16077 ) );
NAND2_X1 _u10_U4626  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n16078 ) );
NAND2_X1 _u10_U4625  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n16079 ) );
NAND2_X1 _u10_U4624  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n16080 ) );
NAND4_X1 _u10_U4623  ( .A1(_u10_n16077 ), .A2(_u10_n16078 ), .A3(_u10_n16079 ), .A4(_u10_n16080 ), .ZN(_u10_n16062 ) );
NAND2_X1 _u10_U4622  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n16073 ) );
NAND2_X1 _u10_U4621  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n16074 ) );
NAND2_X1 _u10_U4620  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n16075 ) );
NAND2_X1 _u10_U4619  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n16076 ) );
NAND4_X1 _u10_U4618  ( .A1(_u10_n16073 ), .A2(_u10_n16074 ), .A3(_u10_n16075 ), .A4(_u10_n16076 ), .ZN(_u10_n16063 ) );
NAND2_X1 _u10_U4617  ( .A1(1'b0), .A2(_u10_n12160 ), .ZN(_u10_n16069 ) );
NAND2_X1 _u10_U4616  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n16070 ) );
NAND2_X1 _u10_U4615  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n16071 ) );
NAND2_X1 _u10_U4614  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n16072 ) );
NAND4_X1 _u10_U4613  ( .A1(_u10_n16069 ), .A2(_u10_n16070 ), .A3(_u10_n16071 ), .A4(_u10_n16072 ), .ZN(_u10_n16064 ) );
NAND2_X1 _u10_U4612  ( .A1(1'b0), .A2(_u10_n12066 ), .ZN(_u10_n16066 ) );
NAND2_X1 _u10_U4611  ( .A1(1'b0), .A2(_u10_n12042 ), .ZN(_u10_n16067 ) );
NAND2_X1 _u10_U4610  ( .A1(1'b0), .A2(_u10_n12012 ), .ZN(_u10_n16068 ) );
NAND3_X1 _u10_U4609  ( .A1(_u10_n16066 ), .A2(_u10_n16067 ), .A3(_u10_n16068 ), .ZN(_u10_n16065 ) );
NOR4_X1 _u10_U4608  ( .A1(_u10_n16062 ), .A2(_u10_n16063 ), .A3(_u10_n16064 ), .A4(_u10_n16065 ), .ZN(_u10_n16040 ) );
NAND2_X1 _u10_U4607  ( .A1(1'b0), .A2(_u10_n11993 ), .ZN(_u10_n16058 ) );
NAND2_X1 _u10_U4606  ( .A1(1'b0), .A2(_u10_n11973 ), .ZN(_u10_n16059 ) );
NAND2_X1 _u10_U4605  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n16060 ) );
NAND2_X1 _u10_U4604  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n16061 ) );
NAND4_X1 _u10_U4603  ( .A1(_u10_n16058 ), .A2(_u10_n16059 ), .A3(_u10_n16060 ), .A4(_u10_n16061 ), .ZN(_u10_n16042 ) );
NAND2_X1 _u10_U4602  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n16054 ) );
NAND2_X1 _u10_U4601  ( .A1(1'b0), .A2(_u10_n11873 ), .ZN(_u10_n16055 ) );
NAND2_X1 _u10_U4600  ( .A1(1'b0), .A2(_u10_n11855 ), .ZN(_u10_n16056 ) );
NAND2_X1 _u10_U4599  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n16057 ) );
NAND4_X1 _u10_U4598  ( .A1(_u10_n16054 ), .A2(_u10_n16055 ), .A3(_u10_n16056 ), .A4(_u10_n16057 ), .ZN(_u10_n16043 ) );
NAND2_X1 _u10_U4597  ( .A1(1'b0), .A2(_u10_n11801 ), .ZN(_u10_n16050 ) );
NAND2_X1 _u10_U4596  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n16051 ) );
NAND2_X1 _u10_U4595  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n16052 ) );
NAND2_X1 _u10_U4594  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n16053 ) );
NAND4_X1 _u10_U4593  ( .A1(_u10_n16050 ), .A2(_u10_n16051 ), .A3(_u10_n16052 ), .A4(_u10_n16053 ), .ZN(_u10_n16044 ) );
NAND2_X1 _u10_U4592  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n16046 ) );
NAND2_X1 _u10_U4591  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n16047 ) );
NAND2_X1 _u10_U4590  ( .A1(1'b0), .A2(_u10_n11663 ), .ZN(_u10_n16048 ) );
NAND2_X1 _u10_U4589  ( .A1(1'b0), .A2(_u10_n11639 ), .ZN(_u10_n16049 ) );
NAND4_X1 _u10_U4588  ( .A1(_u10_n16046 ), .A2(_u10_n16047 ), .A3(_u10_n16048 ), .A4(_u10_n16049 ), .ZN(_u10_n16045 ) );
NOR4_X1 _u10_U4587  ( .A1(_u10_n16042 ), .A2(_u10_n16043 ), .A3(_u10_n16044 ), .A4(_u10_n16045 ), .ZN(_u10_n16041 ) );
NAND2_X1 _u10_U4586  ( .A1(_u10_n16040 ), .A2(_u10_n16041 ), .ZN(pointer[15]) );
NAND2_X1 _u10_U4585  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n16036 ) );
NAND2_X1 _u10_U4584  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n16037 ) );
NAND2_X1 _u10_U4583  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n16038 ) );
NAND2_X1 _u10_U4582  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n16039 ) );
NAND4_X1 _u10_U4581  ( .A1(_u10_n16036 ), .A2(_u10_n16037 ), .A3(_u10_n16038 ), .A4(_u10_n16039 ), .ZN(_u10_n16021 ) );
NAND2_X1 _u10_U4580  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n16032 ) );
NAND2_X1 _u10_U4579  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n16033 ) );
NAND2_X1 _u10_U4578  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n16034 ) );
NAND2_X1 _u10_U4577  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n16035 ) );
NAND4_X1 _u10_U4576  ( .A1(_u10_n16032 ), .A2(_u10_n16033 ), .A3(_u10_n16034 ), .A4(_u10_n16035 ), .ZN(_u10_n16022 ) );
NAND2_X1 _u10_U4575  ( .A1(1'b0), .A2(_u10_n12414 ), .ZN(_u10_n16028 ) );
NAND2_X1 _u10_U4574  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n16029 ) );
NAND2_X1 _u10_U4573  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n16030 ) );
NAND2_X1 _u10_U4572  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n16031 ) );
NAND4_X1 _u10_U4571  ( .A1(_u10_n16028 ), .A2(_u10_n16029 ), .A3(_u10_n16030 ), .A4(_u10_n16031 ), .ZN(_u10_n16023 ) );
NAND2_X1 _u10_U4570  ( .A1(1'b0), .A2(_u10_n12063 ), .ZN(_u10_n16025 ) );
NAND2_X1 _u10_U4569  ( .A1(1'b0), .A2(_u10_n12039 ), .ZN(_u10_n16026 ) );
NAND2_X1 _u10_U4568  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n16027 ) );
NAND3_X1 _u10_U4567  ( .A1(_u10_n16025 ), .A2(_u10_n16026 ), .A3(_u10_n16027 ), .ZN(_u10_n16024 ) );
NOR4_X1 _u10_U4566  ( .A1(_u10_n16021 ), .A2(_u10_n16022 ), .A3(_u10_n16023 ), .A4(_u10_n16024 ), .ZN(_u10_n15999 ) );
NAND2_X1 _u10_U4565  ( .A1(1'b0), .A2(_u10_n11999 ), .ZN(_u10_n16017 ) );
NAND2_X1 _u10_U4564  ( .A1(1'b0), .A2(_u10_n11971 ), .ZN(_u10_n16018 ) );
NAND2_X1 _u10_U4563  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n16019 ) );
NAND2_X1 _u10_U4562  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n16020 ) );
NAND4_X1 _u10_U4561  ( .A1(_u10_n16017 ), .A2(_u10_n16018 ), .A3(_u10_n16019 ), .A4(_u10_n16020 ), .ZN(_u10_n16001 ) );
NAND2_X1 _u10_U4560  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n16013 ) );
NAND2_X1 _u10_U4559  ( .A1(1'b0), .A2(_u10_n11879 ), .ZN(_u10_n16014 ) );
NAND2_X1 _u10_U4558  ( .A1(1'b0), .A2(_u10_n11849 ), .ZN(_u10_n16015 ) );
NAND2_X1 _u10_U4557  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n16016 ) );
NAND4_X1 _u10_U4556  ( .A1(_u10_n16013 ), .A2(_u10_n16014 ), .A3(_u10_n16015 ), .A4(_u10_n16016 ), .ZN(_u10_n16002 ) );
NAND2_X1 _u10_U4555  ( .A1(1'b0), .A2(_u10_n11807 ), .ZN(_u10_n16009 ) );
NAND2_X1 _u10_U4554  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n16010 ) );
NAND2_X1 _u10_U4553  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n16011 ) );
NAND2_X1 _u10_U4552  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n16012 ) );
NAND4_X1 _u10_U4551  ( .A1(_u10_n16009 ), .A2(_u10_n16010 ), .A3(_u10_n16011 ), .A4(_u10_n16012 ), .ZN(_u10_n16003 ) );
NAND2_X1 _u10_U4550  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n16005 ) );
NAND2_X1 _u10_U4549  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n16006 ) );
NAND2_X1 _u10_U4548  ( .A1(1'b0), .A2(_u10_n11657 ), .ZN(_u10_n16007 ) );
NAND2_X1 _u10_U4547  ( .A1(1'b0), .A2(_u10_n11633 ), .ZN(_u10_n16008 ) );
NAND4_X1 _u10_U4546  ( .A1(_u10_n16005 ), .A2(_u10_n16006 ), .A3(_u10_n16007 ), .A4(_u10_n16008 ), .ZN(_u10_n16004 ) );
NOR4_X1 _u10_U4545  ( .A1(_u10_n16001 ), .A2(_u10_n16002 ), .A3(_u10_n16003 ), .A4(_u10_n16004 ), .ZN(_u10_n16000 ) );
NAND2_X1 _u10_U4544  ( .A1(_u10_n15999 ), .A2(_u10_n16000 ), .ZN(pointer[16]) );
NAND2_X1 _u10_U4543  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n15995 ) );
NAND2_X1 _u10_U4542  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n15996 ) );
NAND2_X1 _u10_U4541  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n15997 ) );
NAND2_X1 _u10_U4540  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n15998 ) );
NAND4_X1 _u10_U4539  ( .A1(_u10_n15995 ), .A2(_u10_n15996 ), .A3(_u10_n15997 ), .A4(_u10_n15998 ), .ZN(_u10_n15980 ) );
NAND2_X1 _u10_U4538  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n15991 ) );
NAND2_X1 _u10_U4537  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n15992 ) );
NAND2_X1 _u10_U4536  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n15993 ) );
NAND2_X1 _u10_U4535  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n15994 ) );
NAND4_X1 _u10_U4534  ( .A1(_u10_n15991 ), .A2(_u10_n15992 ), .A3(_u10_n15993 ), .A4(_u10_n15994 ), .ZN(_u10_n15981 ) );
NAND2_X1 _u10_U4533  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n15987 ) );
NAND2_X1 _u10_U4532  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n15988 ) );
NAND2_X1 _u10_U4531  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n15989 ) );
NAND2_X1 _u10_U4530  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n15990 ) );
NAND4_X1 _u10_U4529  ( .A1(_u10_n15987 ), .A2(_u10_n15988 ), .A3(_u10_n15989 ), .A4(_u10_n15990 ), .ZN(_u10_n15982 ) );
NAND2_X1 _u10_U4528  ( .A1(1'b0), .A2(_u10_n12065 ), .ZN(_u10_n15984 ) );
NAND2_X1 _u10_U4527  ( .A1(1'b0), .A2(_u10_n12041 ), .ZN(_u10_n15985 ) );
NAND2_X1 _u10_U4526  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15986 ) );
NAND3_X1 _u10_U4525  ( .A1(_u10_n15984 ), .A2(_u10_n15985 ), .A3(_u10_n15986 ), .ZN(_u10_n15983 ) );
NOR4_X1 _u10_U4524  ( .A1(_u10_n15980 ), .A2(_u10_n15981 ), .A3(_u10_n15982 ), .A4(_u10_n15983 ), .ZN(_u10_n15958 ) );
NAND2_X1 _u10_U4523  ( .A1(1'b0), .A2(_u10_n11996 ), .ZN(_u10_n15976 ) );
NAND2_X1 _u10_U4522  ( .A1(1'b0), .A2(_u10_n11972 ), .ZN(_u10_n15977 ) );
NAND2_X1 _u10_U4521  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n15978 ) );
NAND2_X1 _u10_U4520  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n15979 ) );
NAND4_X1 _u10_U4519  ( .A1(_u10_n15976 ), .A2(_u10_n15977 ), .A3(_u10_n15978 ), .A4(_u10_n15979 ), .ZN(_u10_n15960 ) );
NAND2_X1 _u10_U4518  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n15972 ) );
NAND2_X1 _u10_U4517  ( .A1(1'b0), .A2(_u10_n11876 ), .ZN(_u10_n15973 ) );
NAND2_X1 _u10_U4516  ( .A1(1'b0), .A2(_u10_n11854 ), .ZN(_u10_n15974 ) );
NAND2_X1 _u10_U4515  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n15975 ) );
NAND4_X1 _u10_U4514  ( .A1(_u10_n15972 ), .A2(_u10_n15973 ), .A3(_u10_n15974 ), .A4(_u10_n15975 ), .ZN(_u10_n15961 ) );
NAND2_X1 _u10_U4513  ( .A1(1'b0), .A2(_u10_n11804 ), .ZN(_u10_n15968 ) );
NAND2_X1 _u10_U4512  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n15969 ) );
NAND2_X1 _u10_U4511  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n15970 ) );
NAND2_X1 _u10_U4510  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n15971 ) );
NAND4_X1 _u10_U4509  ( .A1(_u10_n15968 ), .A2(_u10_n15969 ), .A3(_u10_n15970 ), .A4(_u10_n15971 ), .ZN(_u10_n15962 ) );
NAND2_X1 _u10_U4508  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n15964 ) );
NAND2_X1 _u10_U4507  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n15965 ) );
NAND2_X1 _u10_U4506  ( .A1(1'b0), .A2(_u10_n11660 ), .ZN(_u10_n15966 ) );
NAND2_X1 _u10_U4505  ( .A1(1'b0), .A2(_u10_n11638 ), .ZN(_u10_n15967 ) );
NAND4_X1 _u10_U4504  ( .A1(_u10_n15964 ), .A2(_u10_n15965 ), .A3(_u10_n15966 ), .A4(_u10_n15967 ), .ZN(_u10_n15963 ) );
NOR4_X1 _u10_U4503  ( .A1(_u10_n15960 ), .A2(_u10_n15961 ), .A3(_u10_n15962 ), .A4(_u10_n15963 ), .ZN(_u10_n15959 ) );
NAND2_X1 _u10_U4502  ( .A1(_u10_n15958 ), .A2(_u10_n15959 ), .ZN(pointer[17]) );
NAND2_X1 _u10_U4501  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n15954 ) );
NAND2_X1 _u10_U4500  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n15955 ) );
NAND2_X1 _u10_U4499  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n15956 ) );
NAND2_X1 _u10_U4498  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n15957 ) );
NAND4_X1 _u10_U4497  ( .A1(_u10_n15954 ), .A2(_u10_n15955 ), .A3(_u10_n15956 ), .A4(_u10_n15957 ), .ZN(_u10_n15939 ) );
NAND2_X1 _u10_U4496  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n15950 ) );
NAND2_X1 _u10_U4495  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n15951 ) );
NAND2_X1 _u10_U4494  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n15952 ) );
NAND2_X1 _u10_U4493  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n15953 ) );
NAND4_X1 _u10_U4492  ( .A1(_u10_n15950 ), .A2(_u10_n15951 ), .A3(_u10_n15952 ), .A4(_u10_n15953 ), .ZN(_u10_n15940 ) );
NAND2_X1 _u10_U4491  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n15946 ) );
NAND2_X1 _u10_U4490  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n15947 ) );
NAND2_X1 _u10_U4489  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n15948 ) );
NAND2_X1 _u10_U4488  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n15949 ) );
NAND4_X1 _u10_U4487  ( .A1(_u10_n15946 ), .A2(_u10_n15947 ), .A3(_u10_n15948 ), .A4(_u10_n15949 ), .ZN(_u10_n15941 ) );
NAND2_X1 _u10_U4486  ( .A1(1'b0), .A2(_u10_n12406 ), .ZN(_u10_n15943 ) );
NAND2_X1 _u10_U4485  ( .A1(1'b0), .A2(_u10_n12405 ), .ZN(_u10_n15944 ) );
NAND2_X1 _u10_U4484  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15945 ) );
NAND3_X1 _u10_U4483  ( .A1(_u10_n15943 ), .A2(_u10_n15944 ), .A3(_u10_n15945 ), .ZN(_u10_n15942 ) );
NOR4_X1 _u10_U4482  ( .A1(_u10_n15939 ), .A2(_u10_n15940 ), .A3(_u10_n15941 ), .A4(_u10_n15942 ), .ZN(_u10_n15917 ) );
NAND2_X1 _u10_U4481  ( .A1(1'b0), .A2(_u10_n11997 ), .ZN(_u10_n15935 ) );
NAND2_X1 _u10_U4480  ( .A1(1'b0), .A2(_u10_n11975 ), .ZN(_u10_n15936 ) );
NAND2_X1 _u10_U4479  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n15937 ) );
NAND2_X1 _u10_U4478  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n15938 ) );
NAND4_X1 _u10_U4477  ( .A1(_u10_n15935 ), .A2(_u10_n15936 ), .A3(_u10_n15937 ), .A4(_u10_n15938 ), .ZN(_u10_n15919 ) );
NAND2_X1 _u10_U4476  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n15931 ) );
NAND2_X1 _u10_U4475  ( .A1(1'b0), .A2(_u10_n11877 ), .ZN(_u10_n15932 ) );
NAND2_X1 _u10_U4474  ( .A1(1'b0), .A2(_u10_n11852 ), .ZN(_u10_n15933 ) );
NAND2_X1 _u10_U4473  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n15934 ) );
NAND4_X1 _u10_U4472  ( .A1(_u10_n15931 ), .A2(_u10_n15932 ), .A3(_u10_n15933 ), .A4(_u10_n15934 ), .ZN(_u10_n15920 ) );
NAND2_X1 _u10_U4471  ( .A1(1'b0), .A2(_u10_n11805 ), .ZN(_u10_n15927 ) );
NAND2_X1 _u10_U4470  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n15928 ) );
NAND2_X1 _u10_U4469  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n15929 ) );
NAND2_X1 _u10_U4468  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n15930 ) );
NAND4_X1 _u10_U4467  ( .A1(_u10_n15927 ), .A2(_u10_n15928 ), .A3(_u10_n15929 ), .A4(_u10_n15930 ), .ZN(_u10_n15921 ) );
NAND2_X1 _u10_U4466  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n15923 ) );
NAND2_X1 _u10_U4465  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n15924 ) );
NAND2_X1 _u10_U4464  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n15925 ) );
NAND2_X1 _u10_U4463  ( .A1(1'b0), .A2(_u10_n11636 ), .ZN(_u10_n15926 ) );
NAND4_X1 _u10_U4462  ( .A1(_u10_n15923 ), .A2(_u10_n15924 ), .A3(_u10_n15925 ), .A4(_u10_n15926 ), .ZN(_u10_n15922 ) );
NOR4_X1 _u10_U4461  ( .A1(_u10_n15919 ), .A2(_u10_n15920 ), .A3(_u10_n15921 ), .A4(_u10_n15922 ), .ZN(_u10_n15918 ) );
NAND2_X1 _u10_U4460  ( .A1(_u10_n15917 ), .A2(_u10_n15918 ), .ZN(pointer[18]) );
NAND2_X1 _u10_U4459  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n15913 ) );
NAND2_X1 _u10_U4458  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n15914 ) );
NAND2_X1 _u10_U4457  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n15915 ) );
NAND2_X1 _u10_U4456  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n15916 ) );
NAND4_X1 _u10_U4455  ( .A1(_u10_n15913 ), .A2(_u10_n15914 ), .A3(_u10_n15915 ), .A4(_u10_n15916 ), .ZN(_u10_n15898 ) );
NAND2_X1 _u10_U4454  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n15909 ) );
NAND2_X1 _u10_U4453  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n15910 ) );
NAND2_X1 _u10_U4452  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n15911 ) );
NAND2_X1 _u10_U4451  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n15912 ) );
NAND4_X1 _u10_U4450  ( .A1(_u10_n15909 ), .A2(_u10_n15910 ), .A3(_u10_n15911 ), .A4(_u10_n15912 ), .ZN(_u10_n15899 ) );
NAND2_X1 _u10_U4449  ( .A1(1'b0), .A2(_u10_n12162 ), .ZN(_u10_n15905 ) );
NAND2_X1 _u10_U4448  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n15906 ) );
NAND2_X1 _u10_U4447  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n15907 ) );
NAND2_X1 _u10_U4446  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n15908 ) );
NAND4_X1 _u10_U4445  ( .A1(_u10_n15905 ), .A2(_u10_n15906 ), .A3(_u10_n15907 ), .A4(_u10_n15908 ), .ZN(_u10_n15900 ) );
NAND2_X1 _u10_U4444  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n15902 ) );
NAND2_X1 _u10_U4443  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n15903 ) );
NAND2_X1 _u10_U4442  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15904 ) );
NAND3_X1 _u10_U4441  ( .A1(_u10_n15902 ), .A2(_u10_n15903 ), .A3(_u10_n15904 ), .ZN(_u10_n15901 ) );
NOR4_X1 _u10_U4440  ( .A1(_u10_n15898 ), .A2(_u10_n15899 ), .A3(_u10_n15900 ), .A4(_u10_n15901 ), .ZN(_u10_n15876 ) );
NAND2_X1 _u10_U4439  ( .A1(1'b0), .A2(_u10_n12396 ), .ZN(_u10_n15894 ) );
NAND2_X1 _u10_U4438  ( .A1(1'b0), .A2(_u10_n11971 ), .ZN(_u10_n15895 ) );
NAND2_X1 _u10_U4437  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n15896 ) );
NAND2_X1 _u10_U4436  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n15897 ) );
NAND4_X1 _u10_U4435  ( .A1(_u10_n15894 ), .A2(_u10_n15895 ), .A3(_u10_n15896 ), .A4(_u10_n15897 ), .ZN(_u10_n15878 ) );
NAND2_X1 _u10_U4434  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n15890 ) );
NAND2_X1 _u10_U4433  ( .A1(1'b0), .A2(_u10_n12387 ), .ZN(_u10_n15891 ) );
NAND2_X1 _u10_U4432  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n15892 ) );
NAND2_X1 _u10_U4431  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n15893 ) );
NAND4_X1 _u10_U4430  ( .A1(_u10_n15890 ), .A2(_u10_n15891 ), .A3(_u10_n15892 ), .A4(_u10_n15893 ), .ZN(_u10_n15879 ) );
NAND2_X1 _u10_U4429  ( .A1(1'b0), .A2(_u10_n12380 ), .ZN(_u10_n15886 ) );
NAND2_X1 _u10_U4428  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n15887 ) );
NAND2_X1 _u10_U4427  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n15888 ) );
NAND2_X1 _u10_U4426  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n15889 ) );
NAND4_X1 _u10_U4425  ( .A1(_u10_n15886 ), .A2(_u10_n15887 ), .A3(_u10_n15888 ), .A4(_u10_n15889 ), .ZN(_u10_n15880 ) );
NAND2_X1 _u10_U4424  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n15882 ) );
NAND2_X1 _u10_U4423  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n15883 ) );
NAND2_X1 _u10_U4422  ( .A1(1'b0), .A2(_u10_n11662 ), .ZN(_u10_n15884 ) );
NAND2_X1 _u10_U4421  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n15885 ) );
NAND4_X1 _u10_U4420  ( .A1(_u10_n15882 ), .A2(_u10_n15883 ), .A3(_u10_n15884 ), .A4(_u10_n15885 ), .ZN(_u10_n15881 ) );
NOR4_X1 _u10_U4419  ( .A1(_u10_n15878 ), .A2(_u10_n15879 ), .A3(_u10_n15880 ), .A4(_u10_n15881 ), .ZN(_u10_n15877 ) );
NAND2_X1 _u10_U4418  ( .A1(_u10_n15876 ), .A2(_u10_n15877 ), .ZN(pointer[19]) );
NAND2_X1 _u10_U4417  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n15872 ) );
NAND2_X1 _u10_U4416  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n15873 ) );
NAND2_X1 _u10_U4415  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n15874 ) );
NAND2_X1 _u10_U4414  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n15875 ) );
NAND4_X1 _u10_U4413  ( .A1(_u10_n15872 ), .A2(_u10_n15873 ), .A3(_u10_n15874 ), .A4(_u10_n15875 ), .ZN(_u10_n15857 ) );
NAND2_X1 _u10_U4412  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n15868 ) );
NAND2_X1 _u10_U4411  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n15869 ) );
NAND2_X1 _u10_U4410  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n15870 ) );
NAND2_X1 _u10_U4409  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n15871 ) );
NAND4_X1 _u10_U4408  ( .A1(_u10_n15868 ), .A2(_u10_n15869 ), .A3(_u10_n15870 ), .A4(_u10_n15871 ), .ZN(_u10_n15858 ) );
NAND2_X1 _u10_U4407  ( .A1(1'b0), .A2(_u10_n12161 ), .ZN(_u10_n15864 ) );
NAND2_X1 _u10_U4406  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n15865 ) );
NAND2_X1 _u10_U4405  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n15866 ) );
NAND2_X1 _u10_U4404  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n15867 ) );
NAND4_X1 _u10_U4403  ( .A1(_u10_n15864 ), .A2(_u10_n15865 ), .A3(_u10_n15866 ), .A4(_u10_n15867 ), .ZN(_u10_n15859 ) );
NAND2_X1 _u10_U4402  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n15861 ) );
NAND2_X1 _u10_U4401  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n15862 ) );
NAND2_X1 _u10_U4400  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15863 ) );
NAND3_X1 _u10_U4399  ( .A1(_u10_n15861 ), .A2(_u10_n15862 ), .A3(_u10_n15863 ), .ZN(_u10_n15860 ) );
NOR4_X1 _u10_U4398  ( .A1(_u10_n15857 ), .A2(_u10_n15858 ), .A3(_u10_n15859 ), .A4(_u10_n15860 ), .ZN(_u10_n15835 ) );
NAND2_X1 _u10_U4397  ( .A1(1'b0), .A2(_u10_n11999 ), .ZN(_u10_n15853 ) );
NAND2_X1 _u10_U4396  ( .A1(1'b0), .A2(_u10_n11970 ), .ZN(_u10_n15854 ) );
NAND2_X1 _u10_U4395  ( .A1(1'b0), .A2(_u10_n11931 ), .ZN(_u10_n15855 ) );
NAND2_X1 _u10_U4394  ( .A1(1'b0), .A2(_u10_n11907 ), .ZN(_u10_n15856 ) );
NAND4_X1 _u10_U4393  ( .A1(_u10_n15853 ), .A2(_u10_n15854 ), .A3(_u10_n15855 ), .A4(_u10_n15856 ), .ZN(_u10_n15837 ) );
NAND2_X1 _u10_U4392  ( .A1(1'b0), .A2(_u10_n11883 ), .ZN(_u10_n15849 ) );
NAND2_X1 _u10_U4391  ( .A1(1'b0), .A2(_u10_n11879 ), .ZN(_u10_n15850 ) );
NAND2_X1 _u10_U4390  ( .A1(1'b0), .A2(_u10_n12386 ), .ZN(_u10_n15851 ) );
NAND2_X1 _u10_U4389  ( .A1(1'b0), .A2(_u10_n11811 ), .ZN(_u10_n15852 ) );
NAND4_X1 _u10_U4388  ( .A1(_u10_n15849 ), .A2(_u10_n15850 ), .A3(_u10_n15851 ), .A4(_u10_n15852 ), .ZN(_u10_n15838 ) );
NAND2_X1 _u10_U4387  ( .A1(1'b0), .A2(_u10_n11807 ), .ZN(_u10_n15845 ) );
NAND2_X1 _u10_U4386  ( .A1(1'b0), .A2(_u10_n11763 ), .ZN(_u10_n15846 ) );
NAND2_X1 _u10_U4385  ( .A1(1'b0), .A2(_u10_n11736 ), .ZN(_u10_n15847 ) );
NAND2_X1 _u10_U4384  ( .A1(1'b0), .A2(_u10_n11712 ), .ZN(_u10_n15848 ) );
NAND4_X1 _u10_U4383  ( .A1(_u10_n15845 ), .A2(_u10_n15846 ), .A3(_u10_n15847 ), .A4(_u10_n15848 ), .ZN(_u10_n15839 ) );
NAND2_X1 _u10_U4382  ( .A1(1'b0), .A2(_u10_n11688 ), .ZN(_u10_n15841 ) );
NAND2_X1 _u10_U4381  ( .A1(1'b0), .A2(_u10_n11664 ), .ZN(_u10_n15842 ) );
NAND2_X1 _u10_U4380  ( .A1(1'b0), .A2(_u10_n12370 ), .ZN(_u10_n15843 ) );
NAND2_X1 _u10_U4379  ( .A1(1'b0), .A2(_u10_n12369 ), .ZN(_u10_n15844 ) );
NAND4_X1 _u10_U4378  ( .A1(_u10_n15841 ), .A2(_u10_n15842 ), .A3(_u10_n15843 ), .A4(_u10_n15844 ), .ZN(_u10_n15840 ) );
NOR4_X1 _u10_U4377  ( .A1(_u10_n15837 ), .A2(_u10_n15838 ), .A3(_u10_n15839 ), .A4(_u10_n15840 ), .ZN(_u10_n15836 ) );
NAND2_X1 _u10_U4376  ( .A1(_u10_n15835 ), .A2(_u10_n15836 ), .ZN(pointer[1]));
NAND2_X1 _u10_U4375  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n15831 ) );
NAND2_X1 _u10_U4374  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n15832 ) );
NAND2_X1 _u10_U4373  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n15833 ) );
NAND2_X1 _u10_U4372  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n15834 ) );
NAND4_X1 _u10_U4371  ( .A1(_u10_n15831 ), .A2(_u10_n15832 ), .A3(_u10_n15833 ), .A4(_u10_n15834 ), .ZN(_u10_n15816 ) );
NAND2_X1 _u10_U4370  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n15827 ) );
NAND2_X1 _u10_U4369  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n15828 ) );
NAND2_X1 _u10_U4368  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n15829 ) );
NAND2_X1 _u10_U4367  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n15830 ) );
NAND4_X1 _u10_U4366  ( .A1(_u10_n15827 ), .A2(_u10_n15828 ), .A3(_u10_n15829 ), .A4(_u10_n15830 ), .ZN(_u10_n15817 ) );
NAND2_X1 _u10_U4365  ( .A1(1'b0), .A2(_u10_n12163 ), .ZN(_u10_n15823 ) );
NAND2_X1 _u10_U4364  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n15824 ) );
NAND2_X1 _u10_U4363  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n15825 ) );
NAND2_X1 _u10_U4362  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n15826 ) );
NAND4_X1 _u10_U4361  ( .A1(_u10_n15823 ), .A2(_u10_n15824 ), .A3(_u10_n15825 ), .A4(_u10_n15826 ), .ZN(_u10_n15818 ) );
NAND2_X1 _u10_U4360  ( .A1(1'b0), .A2(_u10_n12068 ), .ZN(_u10_n15820 ) );
NAND2_X1 _u10_U4359  ( .A1(1'b0), .A2(_u10_n12044 ), .ZN(_u10_n15821 ) );
NAND2_X1 _u10_U4358  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15822 ) );
NAND3_X1 _u10_U4357  ( .A1(_u10_n15820 ), .A2(_u10_n15821 ), .A3(_u10_n15822 ), .ZN(_u10_n15819 ) );
NOR4_X1 _u10_U4356  ( .A1(_u10_n15816 ), .A2(_u10_n15817 ), .A3(_u10_n15818 ), .A4(_u10_n15819 ), .ZN(_u10_n15794 ) );
NAND2_X1 _u10_U4355  ( .A1(1'b0), .A2(_u10_n11994 ), .ZN(_u10_n15812 ) );
NAND2_X1 _u10_U4354  ( .A1(1'b0), .A2(_u10_n11970 ), .ZN(_u10_n15813 ) );
NAND2_X1 _u10_U4353  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15814 ) );
NAND2_X1 _u10_U4352  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15815 ) );
NAND4_X1 _u10_U4351  ( .A1(_u10_n15812 ), .A2(_u10_n15813 ), .A3(_u10_n15814 ), .A4(_u10_n15815 ), .ZN(_u10_n15796 ) );
NAND2_X1 _u10_U4350  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15808 ) );
NAND2_X1 _u10_U4349  ( .A1(1'b0), .A2(_u10_n11874 ), .ZN(_u10_n15809 ) );
NAND2_X1 _u10_U4348  ( .A1(1'b0), .A2(_u10_n11850 ), .ZN(_u10_n15810 ) );
NAND2_X1 _u10_U4347  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15811 ) );
NAND4_X1 _u10_U4346  ( .A1(_u10_n15808 ), .A2(_u10_n15809 ), .A3(_u10_n15810 ), .A4(_u10_n15811 ), .ZN(_u10_n15797 ) );
NAND2_X1 _u10_U4345  ( .A1(1'b0), .A2(_u10_n11802 ), .ZN(_u10_n15804 ) );
NAND2_X1 _u10_U4344  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15805 ) );
NAND2_X1 _u10_U4343  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15806 ) );
NAND2_X1 _u10_U4342  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15807 ) );
NAND4_X1 _u10_U4341  ( .A1(_u10_n15804 ), .A2(_u10_n15805 ), .A3(_u10_n15806 ), .A4(_u10_n15807 ), .ZN(_u10_n15798 ) );
NAND2_X1 _u10_U4340  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15800 ) );
NAND2_X1 _u10_U4339  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15801 ) );
NAND2_X1 _u10_U4338  ( .A1(1'b0), .A2(_u10_n11658 ), .ZN(_u10_n15802 ) );
NAND2_X1 _u10_U4337  ( .A1(1'b0), .A2(_u10_n11634 ), .ZN(_u10_n15803 ) );
NAND4_X1 _u10_U4336  ( .A1(_u10_n15800 ), .A2(_u10_n15801 ), .A3(_u10_n15802 ), .A4(_u10_n15803 ), .ZN(_u10_n15799 ) );
NOR4_X1 _u10_U4335  ( .A1(_u10_n15796 ), .A2(_u10_n15797 ), .A3(_u10_n15798 ), .A4(_u10_n15799 ), .ZN(_u10_n15795 ) );
NAND2_X1 _u10_U4334  ( .A1(_u10_n15794 ), .A2(_u10_n15795 ), .ZN(pointer[20]) );
NAND2_X1 _u10_U4333  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n15790 ) );
NAND2_X1 _u10_U4332  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n15791 ) );
NAND2_X1 _u10_U4331  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n15792 ) );
NAND2_X1 _u10_U4330  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n15793 ) );
NAND4_X1 _u10_U4329  ( .A1(_u10_n15790 ), .A2(_u10_n15791 ), .A3(_u10_n15792 ), .A4(_u10_n15793 ), .ZN(_u10_n15775 ) );
NAND2_X1 _u10_U4328  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n15786 ) );
NAND2_X1 _u10_U4327  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n15787 ) );
NAND2_X1 _u10_U4326  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n15788 ) );
NAND2_X1 _u10_U4325  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n15789 ) );
NAND4_X1 _u10_U4324  ( .A1(_u10_n15786 ), .A2(_u10_n15787 ), .A3(_u10_n15788 ), .A4(_u10_n15789 ), .ZN(_u10_n15776 ) );
NAND2_X1 _u10_U4323  ( .A1(1'b0), .A2(_u10_n12162 ), .ZN(_u10_n15782 ) );
NAND2_X1 _u10_U4322  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n15783 ) );
NAND2_X1 _u10_U4321  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n15784 ) );
NAND2_X1 _u10_U4320  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n15785 ) );
NAND4_X1 _u10_U4319  ( .A1(_u10_n15782 ), .A2(_u10_n15783 ), .A3(_u10_n15784 ), .A4(_u10_n15785 ), .ZN(_u10_n15777 ) );
NAND2_X1 _u10_U4318  ( .A1(1'b0), .A2(_u10_n12067 ), .ZN(_u10_n15779 ) );
NAND2_X1 _u10_U4317  ( .A1(1'b0), .A2(_u10_n12043 ), .ZN(_u10_n15780 ) );
NAND2_X1 _u10_U4316  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15781 ) );
NAND3_X1 _u10_U4315  ( .A1(_u10_n15779 ), .A2(_u10_n15780 ), .A3(_u10_n15781 ), .ZN(_u10_n15778 ) );
NOR4_X1 _u10_U4314  ( .A1(_u10_n15775 ), .A2(_u10_n15776 ), .A3(_u10_n15777 ), .A4(_u10_n15778 ), .ZN(_u10_n15753 ) );
NAND2_X1 _u10_U4313  ( .A1(1'b0), .A2(_u10_n11995 ), .ZN(_u10_n15771 ) );
NAND2_X1 _u10_U4312  ( .A1(1'b0), .A2(_u10_n11975 ), .ZN(_u10_n15772 ) );
NAND2_X1 _u10_U4311  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15773 ) );
NAND2_X1 _u10_U4310  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15774 ) );
NAND4_X1 _u10_U4309  ( .A1(_u10_n15771 ), .A2(_u10_n15772 ), .A3(_u10_n15773 ), .A4(_u10_n15774 ), .ZN(_u10_n15755 ) );
NAND2_X1 _u10_U4308  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15767 ) );
NAND2_X1 _u10_U4307  ( .A1(1'b0), .A2(_u10_n11875 ), .ZN(_u10_n15768 ) );
NAND2_X1 _u10_U4306  ( .A1(1'b0), .A2(_u10_n11851 ), .ZN(_u10_n15769 ) );
NAND2_X1 _u10_U4305  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15770 ) );
NAND4_X1 _u10_U4304  ( .A1(_u10_n15767 ), .A2(_u10_n15768 ), .A3(_u10_n15769 ), .A4(_u10_n15770 ), .ZN(_u10_n15756 ) );
NAND2_X1 _u10_U4303  ( .A1(1'b0), .A2(_u10_n11803 ), .ZN(_u10_n15763 ) );
NAND2_X1 _u10_U4302  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15764 ) );
NAND2_X1 _u10_U4301  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15765 ) );
NAND2_X1 _u10_U4300  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15766 ) );
NAND4_X1 _u10_U4299  ( .A1(_u10_n15763 ), .A2(_u10_n15764 ), .A3(_u10_n15765 ), .A4(_u10_n15766 ), .ZN(_u10_n15757 ) );
NAND2_X1 _u10_U4298  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15759 ) );
NAND2_X1 _u10_U4297  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15760 ) );
NAND2_X1 _u10_U4296  ( .A1(1'b0), .A2(_u10_n11659 ), .ZN(_u10_n15761 ) );
NAND2_X1 _u10_U4295  ( .A1(1'b0), .A2(_u10_n11635 ), .ZN(_u10_n15762 ) );
NAND4_X1 _u10_U4294  ( .A1(_u10_n15759 ), .A2(_u10_n15760 ), .A3(_u10_n15761 ), .A4(_u10_n15762 ), .ZN(_u10_n15758 ) );
NOR4_X1 _u10_U4293  ( .A1(_u10_n15755 ), .A2(_u10_n15756 ), .A3(_u10_n15757 ), .A4(_u10_n15758 ), .ZN(_u10_n15754 ) );
NAND2_X1 _u10_U4292  ( .A1(_u10_n15753 ), .A2(_u10_n15754 ), .ZN(pointer[21]) );
NAND2_X1 _u10_U4291  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n15749 ) );
NAND2_X1 _u10_U4290  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n15750 ) );
NAND2_X1 _u10_U4289  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n15751 ) );
NAND2_X1 _u10_U4288  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n15752 ) );
NAND4_X1 _u10_U4287  ( .A1(_u10_n15749 ), .A2(_u10_n15750 ), .A3(_u10_n15751 ), .A4(_u10_n15752 ), .ZN(_u10_n15734 ) );
NAND2_X1 _u10_U4286  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n15745 ) );
NAND2_X1 _u10_U4285  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n15746 ) );
NAND2_X1 _u10_U4284  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n15747 ) );
NAND2_X1 _u10_U4283  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n15748 ) );
NAND4_X1 _u10_U4282  ( .A1(_u10_n15745 ), .A2(_u10_n15746 ), .A3(_u10_n15747 ), .A4(_u10_n15748 ), .ZN(_u10_n15735 ) );
NAND2_X1 _u10_U4281  ( .A1(1'b0), .A2(_u10_n12159 ), .ZN(_u10_n15741 ) );
NAND2_X1 _u10_U4280  ( .A1(1'b0), .A2(_u10_n12129 ), .ZN(_u10_n15742 ) );
NAND2_X1 _u10_U4279  ( .A1(1'b0), .A2(_u10_n12105 ), .ZN(_u10_n15743 ) );
NAND2_X1 _u10_U4278  ( .A1(1'b0), .A2(_u10_n12081 ), .ZN(_u10_n15744 ) );
NAND4_X1 _u10_U4277  ( .A1(_u10_n15741 ), .A2(_u10_n15742 ), .A3(_u10_n15743 ), .A4(_u10_n15744 ), .ZN(_u10_n15736 ) );
NAND2_X1 _u10_U4276  ( .A1(1'b0), .A2(_u10_n12066 ), .ZN(_u10_n15738 ) );
NAND2_X1 _u10_U4275  ( .A1(1'b0), .A2(_u10_n12042 ), .ZN(_u10_n15739 ) );
NAND2_X1 _u10_U4274  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15740 ) );
NAND3_X1 _u10_U4273  ( .A1(_u10_n15738 ), .A2(_u10_n15739 ), .A3(_u10_n15740 ), .ZN(_u10_n15737 ) );
NOR4_X1 _u10_U4272  ( .A1(_u10_n15734 ), .A2(_u10_n15735 ), .A3(_u10_n15736 ), .A4(_u10_n15737 ), .ZN(_u10_n15712 ) );
NAND2_X1 _u10_U4271  ( .A1(1'b0), .A2(_u10_n11998 ), .ZN(_u10_n15730 ) );
NAND2_X1 _u10_U4270  ( .A1(1'b0), .A2(_u10_n11971 ), .ZN(_u10_n15731 ) );
NAND2_X1 _u10_U4269  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15732 ) );
NAND2_X1 _u10_U4268  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15733 ) );
NAND4_X1 _u10_U4267  ( .A1(_u10_n15730 ), .A2(_u10_n15731 ), .A3(_u10_n15732 ), .A4(_u10_n15733 ), .ZN(_u10_n15714 ) );
NAND2_X1 _u10_U4266  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15726 ) );
NAND2_X1 _u10_U4265  ( .A1(1'b0), .A2(_u10_n11878 ), .ZN(_u10_n15727 ) );
NAND2_X1 _u10_U4264  ( .A1(1'b0), .A2(_u10_n11855 ), .ZN(_u10_n15728 ) );
NAND2_X1 _u10_U4263  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15729 ) );
NAND4_X1 _u10_U4262  ( .A1(_u10_n15726 ), .A2(_u10_n15727 ), .A3(_u10_n15728 ), .A4(_u10_n15729 ), .ZN(_u10_n15715 ) );
NAND2_X1 _u10_U4261  ( .A1(1'b0), .A2(_u10_n11806 ), .ZN(_u10_n15722 ) );
NAND2_X1 _u10_U4260  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15723 ) );
NAND2_X1 _u10_U4259  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15724 ) );
NAND2_X1 _u10_U4258  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15725 ) );
NAND4_X1 _u10_U4257  ( .A1(_u10_n15722 ), .A2(_u10_n15723 ), .A3(_u10_n15724 ), .A4(_u10_n15725 ), .ZN(_u10_n15716 ) );
NAND2_X1 _u10_U4256  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15718 ) );
NAND2_X1 _u10_U4255  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15719 ) );
NAND2_X1 _u10_U4254  ( .A1(1'b0), .A2(_u10_n11663 ), .ZN(_u10_n15720 ) );
NAND2_X1 _u10_U4253  ( .A1(1'b0), .A2(_u10_n11639 ), .ZN(_u10_n15721 ) );
NAND4_X1 _u10_U4252  ( .A1(_u10_n15718 ), .A2(_u10_n15719 ), .A3(_u10_n15720 ), .A4(_u10_n15721 ), .ZN(_u10_n15717 ) );
NOR4_X1 _u10_U4251  ( .A1(_u10_n15714 ), .A2(_u10_n15715 ), .A3(_u10_n15716 ), .A4(_u10_n15717 ), .ZN(_u10_n15713 ) );
NAND2_X1 _u10_U4250  ( .A1(_u10_n15712 ), .A2(_u10_n15713 ), .ZN(pointer[22]) );
NAND2_X1 _u10_U4249  ( .A1(1'b0), .A2(_u10_n12344 ), .ZN(_u10_n15708 ) );
NAND2_X1 _u10_U4248  ( .A1(1'b0), .A2(_u10_n12320 ), .ZN(_u10_n15709 ) );
NAND2_X1 _u10_U4247  ( .A1(1'b0), .A2(_u10_n12297 ), .ZN(_u10_n15710 ) );
NAND2_X1 _u10_U4246  ( .A1(1'b0), .A2(_u10_n12273 ), .ZN(_u10_n15711 ) );
NAND4_X1 _u10_U4245  ( .A1(_u10_n15708 ), .A2(_u10_n15709 ), .A3(_u10_n15710 ), .A4(_u10_n15711 ), .ZN(_u10_n15693 ) );
NAND2_X1 _u10_U4244  ( .A1(1'b0), .A2(_u10_n12248 ), .ZN(_u10_n15704 ) );
NAND2_X1 _u10_U4243  ( .A1(1'b0), .A2(_u10_n12224 ), .ZN(_u10_n15705 ) );
NAND2_X1 _u10_U4242  ( .A1(1'b0), .A2(_u10_n12198 ), .ZN(_u10_n15706 ) );
NAND2_X1 _u10_U4241  ( .A1(1'b0), .A2(_u10_n12176 ), .ZN(_u10_n15707 ) );
NAND4_X1 _u10_U4240  ( .A1(_u10_n15704 ), .A2(_u10_n15705 ), .A3(_u10_n15706 ), .A4(_u10_n15707 ), .ZN(_u10_n15694 ) );
NAND2_X1 _u10_U4239  ( .A1(1'b0), .A2(_u10_n12159 ), .ZN(_u10_n15700 ) );
NAND2_X1 _u10_U4238  ( .A1(1'b0), .A2(_u10_n12137 ), .ZN(_u10_n15701 ) );
NAND2_X1 _u10_U4237  ( .A1(1'b0), .A2(_u10_n12113 ), .ZN(_u10_n15702 ) );
NAND2_X1 _u10_U4236  ( .A1(1'b0), .A2(_u10_n12089 ), .ZN(_u10_n15703 ) );
NAND4_X1 _u10_U4235  ( .A1(_u10_n15700 ), .A2(_u10_n15701 ), .A3(_u10_n15702 ), .A4(_u10_n15703 ), .ZN(_u10_n15695 ) );
NAND2_X1 _u10_U4234  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n15697 ) );
NAND2_X1 _u10_U4233  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n15698 ) );
NAND2_X1 _u10_U4232  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15699 ) );
NAND3_X1 _u10_U4231  ( .A1(_u10_n15697 ), .A2(_u10_n15698 ), .A3(_u10_n15699 ), .ZN(_u10_n15696 ) );
NOR4_X1 _u10_U4230  ( .A1(_u10_n15693 ), .A2(_u10_n15694 ), .A3(_u10_n15695 ), .A4(_u10_n15696 ), .ZN(_u10_n15671 ) );
NAND2_X1 _u10_U4229  ( .A1(1'b0), .A2(_u10_n12396 ), .ZN(_u10_n15689 ) );
NAND2_X1 _u10_U4228  ( .A1(1'b0), .A2(_u10_n11974 ), .ZN(_u10_n15690 ) );
NAND2_X1 _u10_U4227  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15691 ) );
NAND2_X1 _u10_U4226  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15692 ) );
NAND4_X1 _u10_U4225  ( .A1(_u10_n15689 ), .A2(_u10_n15690 ), .A3(_u10_n15691 ), .A4(_u10_n15692 ), .ZN(_u10_n15673 ) );
NAND2_X1 _u10_U4224  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15685 ) );
NAND2_X1 _u10_U4223  ( .A1(1'b0), .A2(_u10_n12387 ), .ZN(_u10_n15686 ) );
NAND2_X1 _u10_U4222  ( .A1(1'b0), .A2(_u10_n12386 ), .ZN(_u10_n15687 ) );
NAND2_X1 _u10_U4221  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15688 ) );
NAND4_X1 _u10_U4220  ( .A1(_u10_n15685 ), .A2(_u10_n15686 ), .A3(_u10_n15687 ), .A4(_u10_n15688 ), .ZN(_u10_n15674 ) );
NAND2_X1 _u10_U4219  ( .A1(1'b0), .A2(_u10_n12380 ), .ZN(_u10_n15681 ) );
NAND2_X1 _u10_U4218  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15682 ) );
NAND2_X1 _u10_U4217  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15683 ) );
NAND2_X1 _u10_U4216  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15684 ) );
NAND4_X1 _u10_U4215  ( .A1(_u10_n15681 ), .A2(_u10_n15682 ), .A3(_u10_n15683 ), .A4(_u10_n15684 ), .ZN(_u10_n15675 ) );
NAND2_X1 _u10_U4214  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15677 ) );
NAND2_X1 _u10_U4213  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15678 ) );
NAND2_X1 _u10_U4212  ( .A1(1'b0), .A2(_u10_n12370 ), .ZN(_u10_n15679 ) );
NAND2_X1 _u10_U4211  ( .A1(1'b0), .A2(_u10_n12369 ), .ZN(_u10_n15680 ) );
NAND4_X1 _u10_U4210  ( .A1(_u10_n15677 ), .A2(_u10_n15678 ), .A3(_u10_n15679 ), .A4(_u10_n15680 ), .ZN(_u10_n15676 ) );
NOR4_X1 _u10_U4209  ( .A1(_u10_n15673 ), .A2(_u10_n15674 ), .A3(_u10_n15675 ), .A4(_u10_n15676 ), .ZN(_u10_n15672 ) );
NAND2_X1 _u10_U4208  ( .A1(_u10_n15671 ), .A2(_u10_n15672 ), .ZN(pointer[23]) );
NAND2_X1 _u10_U4207  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15667 ) );
NAND2_X1 _u10_U4206  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15668 ) );
NAND2_X1 _u10_U4205  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15669 ) );
NAND2_X1 _u10_U4204  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15670 ) );
NAND4_X1 _u10_U4203  ( .A1(_u10_n15667 ), .A2(_u10_n15668 ), .A3(_u10_n15669 ), .A4(_u10_n15670 ), .ZN(_u10_n15652 ) );
NAND2_X1 _u10_U4202  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15663 ) );
NAND2_X1 _u10_U4201  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15664 ) );
NAND2_X1 _u10_U4200  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15665 ) );
NAND2_X1 _u10_U4199  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15666 ) );
NAND4_X1 _u10_U4198  ( .A1(_u10_n15663 ), .A2(_u10_n15664 ), .A3(_u10_n15665 ), .A4(_u10_n15666 ), .ZN(_u10_n15653 ) );
NAND2_X1 _u10_U4197  ( .A1(1'b0), .A2(_u10_n12160 ), .ZN(_u10_n15659 ) );
NAND2_X1 _u10_U4196  ( .A1(1'b0), .A2(_u10_n12139 ), .ZN(_u10_n15660 ) );
NAND2_X1 _u10_U4195  ( .A1(1'b0), .A2(_u10_n12115 ), .ZN(_u10_n15661 ) );
NAND2_X1 _u10_U4194  ( .A1(1'b0), .A2(_u10_n12091 ), .ZN(_u10_n15662 ) );
NAND4_X1 _u10_U4193  ( .A1(_u10_n15659 ), .A2(_u10_n15660 ), .A3(_u10_n15661 ), .A4(_u10_n15662 ), .ZN(_u10_n15654 ) );
NAND2_X1 _u10_U4192  ( .A1(1'b0), .A2(_u10_n12063 ), .ZN(_u10_n15656 ) );
NAND2_X1 _u10_U4191  ( .A1(1'b0), .A2(_u10_n12039 ), .ZN(_u10_n15657 ) );
NAND2_X1 _u10_U4190  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15658 ) );
NAND3_X1 _u10_U4189  ( .A1(_u10_n15656 ), .A2(_u10_n15657 ), .A3(_u10_n15658 ), .ZN(_u10_n15655 ) );
NOR4_X1 _u10_U4188  ( .A1(_u10_n15652 ), .A2(_u10_n15653 ), .A3(_u10_n15654 ), .A4(_u10_n15655 ), .ZN(_u10_n15630 ) );
NAND2_X1 _u10_U4187  ( .A1(1'b0), .A2(_u10_n11993 ), .ZN(_u10_n15648 ) );
NAND2_X1 _u10_U4186  ( .A1(1'b0), .A2(_u10_n12395 ), .ZN(_u10_n15649 ) );
NAND2_X1 _u10_U4185  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15650 ) );
NAND2_X1 _u10_U4184  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15651 ) );
NAND4_X1 _u10_U4183  ( .A1(_u10_n15648 ), .A2(_u10_n15649 ), .A3(_u10_n15650 ), .A4(_u10_n15651 ), .ZN(_u10_n15632 ) );
NAND2_X1 _u10_U4182  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15644 ) );
NAND2_X1 _u10_U4181  ( .A1(1'b0), .A2(_u10_n11873 ), .ZN(_u10_n15645 ) );
NAND2_X1 _u10_U4180  ( .A1(1'b0), .A2(_u10_n11849 ), .ZN(_u10_n15646 ) );
NAND2_X1 _u10_U4179  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15647 ) );
NAND4_X1 _u10_U4178  ( .A1(_u10_n15644 ), .A2(_u10_n15645 ), .A3(_u10_n15646 ), .A4(_u10_n15647 ), .ZN(_u10_n15633 ) );
NAND2_X1 _u10_U4177  ( .A1(1'b0), .A2(_u10_n11801 ), .ZN(_u10_n15640 ) );
NAND2_X1 _u10_U4176  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15641 ) );
NAND2_X1 _u10_U4175  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15642 ) );
NAND2_X1 _u10_U4174  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15643 ) );
NAND4_X1 _u10_U4173  ( .A1(_u10_n15640 ), .A2(_u10_n15641 ), .A3(_u10_n15642 ), .A4(_u10_n15643 ), .ZN(_u10_n15634 ) );
NAND2_X1 _u10_U4172  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15636 ) );
NAND2_X1 _u10_U4171  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15637 ) );
NAND2_X1 _u10_U4170  ( .A1(1'b0), .A2(_u10_n11657 ), .ZN(_u10_n15638 ) );
NAND2_X1 _u10_U4169  ( .A1(1'b0), .A2(_u10_n11633 ), .ZN(_u10_n15639 ) );
NAND4_X1 _u10_U4168  ( .A1(_u10_n15636 ), .A2(_u10_n15637 ), .A3(_u10_n15638 ), .A4(_u10_n15639 ), .ZN(_u10_n15635 ) );
NOR4_X1 _u10_U4167  ( .A1(_u10_n15632 ), .A2(_u10_n15633 ), .A3(_u10_n15634 ), .A4(_u10_n15635 ), .ZN(_u10_n15631 ) );
NAND2_X1 _u10_U4166  ( .A1(_u10_n15630 ), .A2(_u10_n15631 ), .ZN(pointer[24]) );
NAND2_X1 _u10_U4165  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15626 ) );
NAND2_X1 _u10_U4164  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15627 ) );
NAND2_X1 _u10_U4163  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15628 ) );
NAND2_X1 _u10_U4162  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15629 ) );
NAND4_X1 _u10_U4161  ( .A1(_u10_n15626 ), .A2(_u10_n15627 ), .A3(_u10_n15628 ), .A4(_u10_n15629 ), .ZN(_u10_n15611 ) );
NAND2_X1 _u10_U4160  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15622 ) );
NAND2_X1 _u10_U4159  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15623 ) );
NAND2_X1 _u10_U4158  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15624 ) );
NAND2_X1 _u10_U4157  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15625 ) );
NAND4_X1 _u10_U4156  ( .A1(_u10_n15622 ), .A2(_u10_n15623 ), .A3(_u10_n15624 ), .A4(_u10_n15625 ), .ZN(_u10_n15612 ) );
NAND2_X1 _u10_U4155  ( .A1(1'b0), .A2(_u10_n12414 ), .ZN(_u10_n15618 ) );
NAND2_X1 _u10_U4154  ( .A1(1'b0), .A2(_u10_n12135 ), .ZN(_u10_n15619 ) );
NAND2_X1 _u10_U4153  ( .A1(1'b0), .A2(_u10_n12111 ), .ZN(_u10_n15620 ) );
NAND2_X1 _u10_U4152  ( .A1(1'b0), .A2(_u10_n12087 ), .ZN(_u10_n15621 ) );
NAND4_X1 _u10_U4151  ( .A1(_u10_n15618 ), .A2(_u10_n15619 ), .A3(_u10_n15620 ), .A4(_u10_n15621 ), .ZN(_u10_n15613 ) );
NAND2_X1 _u10_U4150  ( .A1(1'b0), .A2(_u10_n12065 ), .ZN(_u10_n15615 ) );
NAND2_X1 _u10_U4149  ( .A1(1'b0), .A2(_u10_n12041 ), .ZN(_u10_n15616 ) );
NAND2_X1 _u10_U4148  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15617 ) );
NAND3_X1 _u10_U4147  ( .A1(_u10_n15615 ), .A2(_u10_n15616 ), .A3(_u10_n15617 ), .ZN(_u10_n15614 ) );
NOR4_X1 _u10_U4146  ( .A1(_u10_n15611 ), .A2(_u10_n15612 ), .A3(_u10_n15613 ), .A4(_u10_n15614 ), .ZN(_u10_n15589 ) );
NAND2_X1 _u10_U4145  ( .A1(1'b0), .A2(_u10_n11996 ), .ZN(_u10_n15607 ) );
NAND2_X1 _u10_U4144  ( .A1(1'b0), .A2(_u10_n11974 ), .ZN(_u10_n15608 ) );
NAND2_X1 _u10_U4143  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15609 ) );
NAND2_X1 _u10_U4142  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15610 ) );
NAND4_X1 _u10_U4141  ( .A1(_u10_n15607 ), .A2(_u10_n15608 ), .A3(_u10_n15609 ), .A4(_u10_n15610 ), .ZN(_u10_n15591 ) );
NAND2_X1 _u10_U4140  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15603 ) );
NAND2_X1 _u10_U4139  ( .A1(1'b0), .A2(_u10_n11876 ), .ZN(_u10_n15604 ) );
NAND2_X1 _u10_U4138  ( .A1(1'b0), .A2(_u10_n11850 ), .ZN(_u10_n15605 ) );
NAND2_X1 _u10_U4137  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15606 ) );
NAND4_X1 _u10_U4136  ( .A1(_u10_n15603 ), .A2(_u10_n15604 ), .A3(_u10_n15605 ), .A4(_u10_n15606 ), .ZN(_u10_n15592 ) );
NAND2_X1 _u10_U4135  ( .A1(1'b0), .A2(_u10_n11804 ), .ZN(_u10_n15599 ) );
NAND2_X1 _u10_U4134  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15600 ) );
NAND2_X1 _u10_U4133  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15601 ) );
NAND2_X1 _u10_U4132  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15602 ) );
NAND4_X1 _u10_U4131  ( .A1(_u10_n15599 ), .A2(_u10_n15600 ), .A3(_u10_n15601 ), .A4(_u10_n15602 ), .ZN(_u10_n15593 ) );
NAND2_X1 _u10_U4130  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15595 ) );
NAND2_X1 _u10_U4129  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15596 ) );
NAND2_X1 _u10_U4128  ( .A1(1'b0), .A2(_u10_n11658 ), .ZN(_u10_n15597 ) );
NAND2_X1 _u10_U4127  ( .A1(1'b0), .A2(_u10_n11634 ), .ZN(_u10_n15598 ) );
NAND4_X1 _u10_U4126  ( .A1(_u10_n15595 ), .A2(_u10_n15596 ), .A3(_u10_n15597 ), .A4(_u10_n15598 ), .ZN(_u10_n15594 ) );
NOR4_X1 _u10_U4125  ( .A1(_u10_n15591 ), .A2(_u10_n15592 ), .A3(_u10_n15593 ), .A4(_u10_n15594 ), .ZN(_u10_n15590 ) );
NAND2_X1 _u10_U4124  ( .A1(_u10_n15589 ), .A2(_u10_n15590 ), .ZN(pointer[25]) );
NAND2_X1 _u10_U4123  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15585 ) );
NAND2_X1 _u10_U4122  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15586 ) );
NAND2_X1 _u10_U4121  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15587 ) );
NAND2_X1 _u10_U4120  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15588 ) );
NAND4_X1 _u10_U4119  ( .A1(_u10_n15585 ), .A2(_u10_n15586 ), .A3(_u10_n15587 ), .A4(_u10_n15588 ), .ZN(_u10_n15570 ) );
NAND2_X1 _u10_U4118  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15581 ) );
NAND2_X1 _u10_U4117  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15582 ) );
NAND2_X1 _u10_U4116  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15583 ) );
NAND2_X1 _u10_U4115  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15584 ) );
NAND4_X1 _u10_U4114  ( .A1(_u10_n15581 ), .A2(_u10_n15582 ), .A3(_u10_n15583 ), .A4(_u10_n15584 ), .ZN(_u10_n15571 ) );
NAND2_X1 _u10_U4113  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n15577 ) );
NAND2_X1 _u10_U4112  ( .A1(1'b0), .A2(_u10_n12136 ), .ZN(_u10_n15578 ) );
NAND2_X1 _u10_U4111  ( .A1(1'b0), .A2(_u10_n12112 ), .ZN(_u10_n15579 ) );
NAND2_X1 _u10_U4110  ( .A1(1'b0), .A2(_u10_n12088 ), .ZN(_u10_n15580 ) );
NAND4_X1 _u10_U4109  ( .A1(_u10_n15577 ), .A2(_u10_n15578 ), .A3(_u10_n15579 ), .A4(_u10_n15580 ), .ZN(_u10_n15572 ) );
NAND2_X1 _u10_U4108  ( .A1(1'b0), .A2(_u10_n12406 ), .ZN(_u10_n15574 ) );
NAND2_X1 _u10_U4107  ( .A1(1'b0), .A2(_u10_n12405 ), .ZN(_u10_n15575 ) );
NAND2_X1 _u10_U4106  ( .A1(1'b0), .A2(_u10_n12013 ), .ZN(_u10_n15576 ) );
NAND3_X1 _u10_U4105  ( .A1(_u10_n15574 ), .A2(_u10_n15575 ), .A3(_u10_n15576 ), .ZN(_u10_n15573 ) );
NOR4_X1 _u10_U4104  ( .A1(_u10_n15570 ), .A2(_u10_n15571 ), .A3(_u10_n15572 ), .A4(_u10_n15573 ), .ZN(_u10_n15548 ) );
NAND2_X1 _u10_U4103  ( .A1(1'b0), .A2(_u10_n11997 ), .ZN(_u10_n15566 ) );
NAND2_X1 _u10_U4102  ( .A1(1'b0), .A2(_u10_n11969 ), .ZN(_u10_n15567 ) );
NAND2_X1 _u10_U4101  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15568 ) );
NAND2_X1 _u10_U4100  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15569 ) );
NAND4_X1 _u10_U4099  ( .A1(_u10_n15566 ), .A2(_u10_n15567 ), .A3(_u10_n15568 ), .A4(_u10_n15569 ), .ZN(_u10_n15550 ) );
NAND2_X1 _u10_U4098  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15562 ) );
NAND2_X1 _u10_U4097  ( .A1(1'b0), .A2(_u10_n11877 ), .ZN(_u10_n15563 ) );
NAND2_X1 _u10_U4096  ( .A1(1'b0), .A2(_u10_n11852 ), .ZN(_u10_n15564 ) );
NAND2_X1 _u10_U4095  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15565 ) );
NAND4_X1 _u10_U4094  ( .A1(_u10_n15562 ), .A2(_u10_n15563 ), .A3(_u10_n15564 ), .A4(_u10_n15565 ), .ZN(_u10_n15551 ) );
NAND2_X1 _u10_U4093  ( .A1(1'b0), .A2(_u10_n11805 ), .ZN(_u10_n15558 ) );
NAND2_X1 _u10_U4092  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15559 ) );
NAND2_X1 _u10_U4091  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15560 ) );
NAND2_X1 _u10_U4090  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15561 ) );
NAND4_X1 _u10_U4089  ( .A1(_u10_n15558 ), .A2(_u10_n15559 ), .A3(_u10_n15560 ), .A4(_u10_n15561 ), .ZN(_u10_n15552 ) );
NAND2_X1 _u10_U4088  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15554 ) );
NAND2_X1 _u10_U4087  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15555 ) );
NAND2_X1 _u10_U4086  ( .A1(1'b0), .A2(_u10_n11660 ), .ZN(_u10_n15556 ) );
NAND2_X1 _u10_U4085  ( .A1(1'b0), .A2(_u10_n11636 ), .ZN(_u10_n15557 ) );
NAND4_X1 _u10_U4084  ( .A1(_u10_n15554 ), .A2(_u10_n15555 ), .A3(_u10_n15556 ), .A4(_u10_n15557 ), .ZN(_u10_n15553 ) );
NOR4_X1 _u10_U4083  ( .A1(_u10_n15550 ), .A2(_u10_n15551 ), .A3(_u10_n15552 ), .A4(_u10_n15553 ), .ZN(_u10_n15549 ) );
NAND2_X1 _u10_U4082  ( .A1(_u10_n15548 ), .A2(_u10_n15549 ), .ZN(pointer[26]) );
NAND2_X1 _u10_U4081  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15544 ) );
NAND2_X1 _u10_U4080  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15545 ) );
NAND2_X1 _u10_U4079  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15546 ) );
NAND2_X1 _u10_U4078  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15547 ) );
NAND4_X1 _u10_U4077  ( .A1(_u10_n15544 ), .A2(_u10_n15545 ), .A3(_u10_n15546 ), .A4(_u10_n15547 ), .ZN(_u10_n15529 ) );
NAND2_X1 _u10_U4076  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15540 ) );
NAND2_X1 _u10_U4075  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15541 ) );
NAND2_X1 _u10_U4074  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15542 ) );
NAND2_X1 _u10_U4073  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15543 ) );
NAND4_X1 _u10_U4072  ( .A1(_u10_n15540 ), .A2(_u10_n15541 ), .A3(_u10_n15542 ), .A4(_u10_n15543 ), .ZN(_u10_n15530 ) );
NAND2_X1 _u10_U4071  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n15536 ) );
NAND2_X1 _u10_U4070  ( .A1(1'b0), .A2(_u10_n12138 ), .ZN(_u10_n15537 ) );
NAND2_X1 _u10_U4069  ( .A1(1'b0), .A2(_u10_n12114 ), .ZN(_u10_n15538 ) );
NAND2_X1 _u10_U4068  ( .A1(1'b0), .A2(_u10_n12090 ), .ZN(_u10_n15539 ) );
NAND4_X1 _u10_U4067  ( .A1(_u10_n15536 ), .A2(_u10_n15537 ), .A3(_u10_n15538 ), .A4(_u10_n15539 ), .ZN(_u10_n15531 ) );
NAND2_X1 _u10_U4066  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n15533 ) );
NAND2_X1 _u10_U4065  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n15534 ) );
NAND2_X1 _u10_U4064  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15535 ) );
NAND3_X1 _u10_U4063  ( .A1(_u10_n15533 ), .A2(_u10_n15534 ), .A3(_u10_n15535 ), .ZN(_u10_n15532 ) );
NOR4_X1 _u10_U4062  ( .A1(_u10_n15529 ), .A2(_u10_n15530 ), .A3(_u10_n15531 ), .A4(_u10_n15532 ), .ZN(_u10_n15507 ) );
NAND2_X1 _u10_U4061  ( .A1(1'b0), .A2(_u10_n11996 ), .ZN(_u10_n15525 ) );
NAND2_X1 _u10_U4060  ( .A1(1'b0), .A2(_u10_n11973 ), .ZN(_u10_n15526 ) );
NAND2_X1 _u10_U4059  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15527 ) );
NAND2_X1 _u10_U4058  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15528 ) );
NAND4_X1 _u10_U4057  ( .A1(_u10_n15525 ), .A2(_u10_n15526 ), .A3(_u10_n15527 ), .A4(_u10_n15528 ), .ZN(_u10_n15509 ) );
NAND2_X1 _u10_U4056  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15521 ) );
NAND2_X1 _u10_U4055  ( .A1(1'b0), .A2(_u10_n11876 ), .ZN(_u10_n15522 ) );
NAND2_X1 _u10_U4054  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n15523 ) );
NAND2_X1 _u10_U4053  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15524 ) );
NAND4_X1 _u10_U4052  ( .A1(_u10_n15521 ), .A2(_u10_n15522 ), .A3(_u10_n15523 ), .A4(_u10_n15524 ), .ZN(_u10_n15510 ) );
NAND2_X1 _u10_U4051  ( .A1(1'b0), .A2(_u10_n11804 ), .ZN(_u10_n15517 ) );
NAND2_X1 _u10_U4050  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15518 ) );
NAND2_X1 _u10_U4049  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15519 ) );
NAND2_X1 _u10_U4048  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15520 ) );
NAND4_X1 _u10_U4047  ( .A1(_u10_n15517 ), .A2(_u10_n15518 ), .A3(_u10_n15519 ), .A4(_u10_n15520 ), .ZN(_u10_n15511 ) );
NAND2_X1 _u10_U4046  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15513 ) );
NAND2_X1 _u10_U4045  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15514 ) );
NAND2_X1 _u10_U4044  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n15515 ) );
NAND2_X1 _u10_U4043  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n15516 ) );
NAND4_X1 _u10_U4042  ( .A1(_u10_n15513 ), .A2(_u10_n15514 ), .A3(_u10_n15515 ), .A4(_u10_n15516 ), .ZN(_u10_n15512 ) );
NOR4_X1 _u10_U4041  ( .A1(_u10_n15509 ), .A2(_u10_n15510 ), .A3(_u10_n15511 ), .A4(_u10_n15512 ), .ZN(_u10_n15508 ) );
NAND2_X1 _u10_U4040  ( .A1(_u10_n15507 ), .A2(_u10_n15508 ), .ZN(pointer[27]) );
NAND2_X1 _u10_U4039  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15503 ) );
NAND2_X1 _u10_U4038  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15504 ) );
NAND2_X1 _u10_U4037  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15505 ) );
NAND2_X1 _u10_U4036  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15506 ) );
NAND4_X1 _u10_U4035  ( .A1(_u10_n15503 ), .A2(_u10_n15504 ), .A3(_u10_n15505 ), .A4(_u10_n15506 ), .ZN(_u10_n15488 ) );
NAND2_X1 _u10_U4034  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15499 ) );
NAND2_X1 _u10_U4033  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15500 ) );
NAND2_X1 _u10_U4032  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15501 ) );
NAND2_X1 _u10_U4031  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15502 ) );
NAND4_X1 _u10_U4030  ( .A1(_u10_n15499 ), .A2(_u10_n15500 ), .A3(_u10_n15501 ), .A4(_u10_n15502 ), .ZN(_u10_n15489 ) );
NAND2_X1 _u10_U4029  ( .A1(1'b0), .A2(_u10_n12161 ), .ZN(_u10_n15495 ) );
NAND2_X1 _u10_U4028  ( .A1(1'b0), .A2(_u10_n12413 ), .ZN(_u10_n15496 ) );
NAND2_X1 _u10_U4027  ( .A1(1'b0), .A2(_u10_n12412 ), .ZN(_u10_n15497 ) );
NAND2_X1 _u10_U4026  ( .A1(1'b0), .A2(_u10_n12411 ), .ZN(_u10_n15498 ) );
NAND4_X1 _u10_U4025  ( .A1(_u10_n15495 ), .A2(_u10_n15496 ), .A3(_u10_n15497 ), .A4(_u10_n15498 ), .ZN(_u10_n15490 ) );
NAND2_X1 _u10_U4024  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n15492 ) );
NAND2_X1 _u10_U4023  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n15493 ) );
NAND2_X1 _u10_U4022  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15494 ) );
NAND3_X1 _u10_U4021  ( .A1(_u10_n15492 ), .A2(_u10_n15493 ), .A3(_u10_n15494 ), .ZN(_u10_n15491 ) );
NOR4_X1 _u10_U4020  ( .A1(_u10_n15488 ), .A2(_u10_n15489 ), .A3(_u10_n15490 ), .A4(_u10_n15491 ), .ZN(_u10_n15466 ) );
NAND2_X1 _u10_U4019  ( .A1(1'b0), .A2(_u10_n11999 ), .ZN(_u10_n15484 ) );
NAND2_X1 _u10_U4018  ( .A1(1'b0), .A2(_u10_n11972 ), .ZN(_u10_n15485 ) );
NAND2_X1 _u10_U4017  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15486 ) );
NAND2_X1 _u10_U4016  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15487 ) );
NAND4_X1 _u10_U4015  ( .A1(_u10_n15484 ), .A2(_u10_n15485 ), .A3(_u10_n15486 ), .A4(_u10_n15487 ), .ZN(_u10_n15468 ) );
NAND2_X1 _u10_U4014  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15480 ) );
NAND2_X1 _u10_U4013  ( .A1(1'b0), .A2(_u10_n11879 ), .ZN(_u10_n15481 ) );
NAND2_X1 _u10_U4012  ( .A1(1'b0), .A2(_u10_n11854 ), .ZN(_u10_n15482 ) );
NAND2_X1 _u10_U4011  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15483 ) );
NAND4_X1 _u10_U4010  ( .A1(_u10_n15480 ), .A2(_u10_n15481 ), .A3(_u10_n15482 ), .A4(_u10_n15483 ), .ZN(_u10_n15469 ) );
NAND2_X1 _u10_U4009  ( .A1(1'b0), .A2(_u10_n11807 ), .ZN(_u10_n15476 ) );
NAND2_X1 _u10_U4008  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15477 ) );
NAND2_X1 _u10_U4007  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15478 ) );
NAND2_X1 _u10_U4006  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15479 ) );
NAND4_X1 _u10_U4005  ( .A1(_u10_n15476 ), .A2(_u10_n15477 ), .A3(_u10_n15478 ), .A4(_u10_n15479 ), .ZN(_u10_n15470 ) );
NAND2_X1 _u10_U4004  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15472 ) );
NAND2_X1 _u10_U4003  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15473 ) );
NAND2_X1 _u10_U4002  ( .A1(1'b0), .A2(_u10_n11662 ), .ZN(_u10_n15474 ) );
NAND2_X1 _u10_U4001  ( .A1(1'b0), .A2(_u10_n11638 ), .ZN(_u10_n15475 ) );
NAND4_X1 _u10_U4000  ( .A1(_u10_n15472 ), .A2(_u10_n15473 ), .A3(_u10_n15474 ), .A4(_u10_n15475 ), .ZN(_u10_n15471 ) );
NOR4_X1 _u10_U3999  ( .A1(_u10_n15468 ), .A2(_u10_n15469 ), .A3(_u10_n15470 ), .A4(_u10_n15471 ), .ZN(_u10_n15467 ) );
NAND2_X1 _u10_U3998  ( .A1(_u10_n15466 ), .A2(_u10_n15467 ), .ZN(pointer[28]) );
NAND2_X1 _u10_U3997  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15462 ) );
NAND2_X1 _u10_U3996  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15463 ) );
NAND2_X1 _u10_U3995  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15464 ) );
NAND2_X1 _u10_U3994  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15465 ) );
NAND4_X1 _u10_U3993  ( .A1(_u10_n15462 ), .A2(_u10_n15463 ), .A3(_u10_n15464 ), .A4(_u10_n15465 ), .ZN(_u10_n15447 ) );
NAND2_X1 _u10_U3992  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15458 ) );
NAND2_X1 _u10_U3991  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15459 ) );
NAND2_X1 _u10_U3990  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15460 ) );
NAND2_X1 _u10_U3989  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15461 ) );
NAND4_X1 _u10_U3988  ( .A1(_u10_n15458 ), .A2(_u10_n15459 ), .A3(_u10_n15460 ), .A4(_u10_n15461 ), .ZN(_u10_n15448 ) );
NAND2_X1 _u10_U3987  ( .A1(1'b0), .A2(_u10_n12161 ), .ZN(_u10_n15454 ) );
NAND2_X1 _u10_U3986  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n15455 ) );
NAND2_X1 _u10_U3985  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n15456 ) );
NAND2_X1 _u10_U3984  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n15457 ) );
NAND4_X1 _u10_U3983  ( .A1(_u10_n15454 ), .A2(_u10_n15455 ), .A3(_u10_n15456 ), .A4(_u10_n15457 ), .ZN(_u10_n15449 ) );
NAND2_X1 _u10_U3982  ( .A1(1'b0), .A2(_u10_n12068 ), .ZN(_u10_n15451 ) );
NAND2_X1 _u10_U3981  ( .A1(1'b0), .A2(_u10_n12044 ), .ZN(_u10_n15452 ) );
NAND2_X1 _u10_U3980  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15453 ) );
NAND3_X1 _u10_U3979  ( .A1(_u10_n15451 ), .A2(_u10_n15452 ), .A3(_u10_n15453 ), .ZN(_u10_n15450 ) );
NOR4_X1 _u10_U3978  ( .A1(_u10_n15447 ), .A2(_u10_n15448 ), .A3(_u10_n15449 ), .A4(_u10_n15450 ), .ZN(_u10_n15425 ) );
NAND2_X1 _u10_U3977  ( .A1(1'b0), .A2(_u10_n11994 ), .ZN(_u10_n15443 ) );
NAND2_X1 _u10_U3976  ( .A1(1'b0), .A2(_u10_n11975 ), .ZN(_u10_n15444 ) );
NAND2_X1 _u10_U3975  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15445 ) );
NAND2_X1 _u10_U3974  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15446 ) );
NAND4_X1 _u10_U3973  ( .A1(_u10_n15443 ), .A2(_u10_n15444 ), .A3(_u10_n15445 ), .A4(_u10_n15446 ), .ZN(_u10_n15427 ) );
NAND2_X1 _u10_U3972  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15439 ) );
NAND2_X1 _u10_U3971  ( .A1(1'b0), .A2(_u10_n11874 ), .ZN(_u10_n15440 ) );
NAND2_X1 _u10_U3970  ( .A1(1'b0), .A2(_u10_n11850 ), .ZN(_u10_n15441 ) );
NAND2_X1 _u10_U3969  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15442 ) );
NAND4_X1 _u10_U3968  ( .A1(_u10_n15439 ), .A2(_u10_n15440 ), .A3(_u10_n15441 ), .A4(_u10_n15442 ), .ZN(_u10_n15428 ) );
NAND2_X1 _u10_U3967  ( .A1(1'b0), .A2(_u10_n11802 ), .ZN(_u10_n15435 ) );
NAND2_X1 _u10_U3966  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15436 ) );
NAND2_X1 _u10_U3965  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15437 ) );
NAND2_X1 _u10_U3964  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15438 ) );
NAND4_X1 _u10_U3963  ( .A1(_u10_n15435 ), .A2(_u10_n15436 ), .A3(_u10_n15437 ), .A4(_u10_n15438 ), .ZN(_u10_n15429 ) );
NAND2_X1 _u10_U3962  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15431 ) );
NAND2_X1 _u10_U3961  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15432 ) );
NAND2_X1 _u10_U3960  ( .A1(1'b0), .A2(_u10_n11658 ), .ZN(_u10_n15433 ) );
NAND2_X1 _u10_U3959  ( .A1(1'b0), .A2(_u10_n11634 ), .ZN(_u10_n15434 ) );
NAND4_X1 _u10_U3958  ( .A1(_u10_n15431 ), .A2(_u10_n15432 ), .A3(_u10_n15433 ), .A4(_u10_n15434 ), .ZN(_u10_n15430 ) );
NOR4_X1 _u10_U3957  ( .A1(_u10_n15427 ), .A2(_u10_n15428 ), .A3(_u10_n15429 ), .A4(_u10_n15430 ), .ZN(_u10_n15426 ) );
NAND2_X1 _u10_U3956  ( .A1(_u10_n15425 ), .A2(_u10_n15426 ), .ZN(pointer[29]) );
NAND2_X1 _u10_U3955  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15421 ) );
NAND2_X1 _u10_U3954  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15422 ) );
NAND2_X1 _u10_U3953  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15423 ) );
NAND2_X1 _u10_U3952  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15424 ) );
NAND4_X1 _u10_U3951  ( .A1(_u10_n15421 ), .A2(_u10_n15422 ), .A3(_u10_n15423 ), .A4(_u10_n15424 ), .ZN(_u10_n15406 ) );
NAND2_X1 _u10_U3950  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15417 ) );
NAND2_X1 _u10_U3949  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15418 ) );
NAND2_X1 _u10_U3948  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15419 ) );
NAND2_X1 _u10_U3947  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15420 ) );
NAND4_X1 _u10_U3946  ( .A1(_u10_n15417 ), .A2(_u10_n15418 ), .A3(_u10_n15419 ), .A4(_u10_n15420 ), .ZN(_u10_n15407 ) );
NAND2_X1 _u10_U3945  ( .A1(1'b0), .A2(_u10_n12163 ), .ZN(_u10_n15413 ) );
NAND2_X1 _u10_U3944  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n15414 ) );
NAND2_X1 _u10_U3943  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n15415 ) );
NAND2_X1 _u10_U3942  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n15416 ) );
NAND4_X1 _u10_U3941  ( .A1(_u10_n15413 ), .A2(_u10_n15414 ), .A3(_u10_n15415 ), .A4(_u10_n15416 ), .ZN(_u10_n15408 ) );
NAND2_X1 _u10_U3940  ( .A1(1'b0), .A2(_u10_n12067 ), .ZN(_u10_n15410 ) );
NAND2_X1 _u10_U3939  ( .A1(1'b0), .A2(_u10_n12043 ), .ZN(_u10_n15411 ) );
NAND2_X1 _u10_U3938  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15412 ) );
NAND3_X1 _u10_U3937  ( .A1(_u10_n15410 ), .A2(_u10_n15411 ), .A3(_u10_n15412 ), .ZN(_u10_n15409 ) );
NOR4_X1 _u10_U3936  ( .A1(_u10_n15406 ), .A2(_u10_n15407 ), .A3(_u10_n15408 ), .A4(_u10_n15409 ), .ZN(_u10_n15384 ) );
NAND2_X1 _u10_U3935  ( .A1(1'b0), .A2(_u10_n11995 ), .ZN(_u10_n15402 ) );
NAND2_X1 _u10_U3934  ( .A1(1'b0), .A2(_u10_n12395 ), .ZN(_u10_n15403 ) );
NAND2_X1 _u10_U3933  ( .A1(1'b0), .A2(_u10_n11932 ), .ZN(_u10_n15404 ) );
NAND2_X1 _u10_U3932  ( .A1(1'b0), .A2(_u10_n11908 ), .ZN(_u10_n15405 ) );
NAND4_X1 _u10_U3931  ( .A1(_u10_n15402 ), .A2(_u10_n15403 ), .A3(_u10_n15404 ), .A4(_u10_n15405 ), .ZN(_u10_n15386 ) );
NAND2_X1 _u10_U3930  ( .A1(1'b0), .A2(_u10_n11884 ), .ZN(_u10_n15398 ) );
NAND2_X1 _u10_U3929  ( .A1(1'b0), .A2(_u10_n11875 ), .ZN(_u10_n15399 ) );
NAND2_X1 _u10_U3928  ( .A1(1'b0), .A2(_u10_n11851 ), .ZN(_u10_n15400 ) );
NAND2_X1 _u10_U3927  ( .A1(1'b0), .A2(_u10_n11812 ), .ZN(_u10_n15401 ) );
NAND4_X1 _u10_U3926  ( .A1(_u10_n15398 ), .A2(_u10_n15399 ), .A3(_u10_n15400 ), .A4(_u10_n15401 ), .ZN(_u10_n15387 ) );
NAND2_X1 _u10_U3925  ( .A1(1'b0), .A2(_u10_n11803 ), .ZN(_u10_n15394 ) );
NAND2_X1 _u10_U3924  ( .A1(1'b0), .A2(_u10_n11764 ), .ZN(_u10_n15395 ) );
NAND2_X1 _u10_U3923  ( .A1(1'b0), .A2(_u10_n11737 ), .ZN(_u10_n15396 ) );
NAND2_X1 _u10_U3922  ( .A1(1'b0), .A2(_u10_n11713 ), .ZN(_u10_n15397 ) );
NAND4_X1 _u10_U3921  ( .A1(_u10_n15394 ), .A2(_u10_n15395 ), .A3(_u10_n15396 ), .A4(_u10_n15397 ), .ZN(_u10_n15388 ) );
NAND2_X1 _u10_U3920  ( .A1(1'b0), .A2(_u10_n11689 ), .ZN(_u10_n15390 ) );
NAND2_X1 _u10_U3919  ( .A1(1'b0), .A2(_u10_n11665 ), .ZN(_u10_n15391 ) );
NAND2_X1 _u10_U3918  ( .A1(1'b0), .A2(_u10_n11659 ), .ZN(_u10_n15392 ) );
NAND2_X1 _u10_U3917  ( .A1(1'b0), .A2(_u10_n11635 ), .ZN(_u10_n15393 ) );
NAND4_X1 _u10_U3916  ( .A1(_u10_n15390 ), .A2(_u10_n15391 ), .A3(_u10_n15392 ), .A4(_u10_n15393 ), .ZN(_u10_n15389 ) );
NOR4_X1 _u10_U3915  ( .A1(_u10_n15386 ), .A2(_u10_n15387 ), .A3(_u10_n15388 ), .A4(_u10_n15389 ), .ZN(_u10_n15385 ) );
NAND2_X1 _u10_U3914  ( .A1(_u10_n15384 ), .A2(_u10_n15385 ), .ZN(pointer[2]));
NAND2_X1 _u10_U3913  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15380 ) );
NAND2_X1 _u10_U3912  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15381 ) );
NAND2_X1 _u10_U3911  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15382 ) );
NAND2_X1 _u10_U3910  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15383 ) );
NAND4_X1 _u10_U3909  ( .A1(_u10_n15380 ), .A2(_u10_n15381 ), .A3(_u10_n15382 ), .A4(_u10_n15383 ), .ZN(_u10_n15365 ) );
NAND2_X1 _u10_U3908  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15376 ) );
NAND2_X1 _u10_U3907  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15377 ) );
NAND2_X1 _u10_U3906  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15378 ) );
NAND2_X1 _u10_U3905  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15379 ) );
NAND4_X1 _u10_U3904  ( .A1(_u10_n15376 ), .A2(_u10_n15377 ), .A3(_u10_n15378 ), .A4(_u10_n15379 ), .ZN(_u10_n15366 ) );
NAND2_X1 _u10_U3903  ( .A1(1'b0), .A2(_u10_n12162 ), .ZN(_u10_n15372 ) );
NAND2_X1 _u10_U3902  ( .A1(1'b0), .A2(_u10_n12137 ), .ZN(_u10_n15373 ) );
NAND2_X1 _u10_U3901  ( .A1(1'b0), .A2(_u10_n12113 ), .ZN(_u10_n15374 ) );
NAND2_X1 _u10_U3900  ( .A1(1'b0), .A2(_u10_n12089 ), .ZN(_u10_n15375 ) );
NAND4_X1 _u10_U3899  ( .A1(_u10_n15372 ), .A2(_u10_n15373 ), .A3(_u10_n15374 ), .A4(_u10_n15375 ), .ZN(_u10_n15367 ) );
NAND2_X1 _u10_U3898  ( .A1(1'b0), .A2(_u10_n12066 ), .ZN(_u10_n15369 ) );
NAND2_X1 _u10_U3897  ( .A1(1'b0), .A2(_u10_n12042 ), .ZN(_u10_n15370 ) );
NAND2_X1 _u10_U3896  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15371 ) );
NAND3_X1 _u10_U3895  ( .A1(_u10_n15369 ), .A2(_u10_n15370 ), .A3(_u10_n15371 ), .ZN(_u10_n15368 ) );
NOR4_X1 _u10_U3894  ( .A1(_u10_n15365 ), .A2(_u10_n15366 ), .A3(_u10_n15367 ), .A4(_u10_n15368 ), .ZN(_u10_n15343 ) );
NAND2_X1 _u10_U3893  ( .A1(1'b0), .A2(_u10_n11998 ), .ZN(_u10_n15361 ) );
NAND2_X1 _u10_U3892  ( .A1(1'b0), .A2(_u10_n11970 ), .ZN(_u10_n15362 ) );
NAND2_X1 _u10_U3891  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n15363 ) );
NAND2_X1 _u10_U3890  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n15364 ) );
NAND4_X1 _u10_U3889  ( .A1(_u10_n15361 ), .A2(_u10_n15362 ), .A3(_u10_n15363 ), .A4(_u10_n15364 ), .ZN(_u10_n15345 ) );
NAND2_X1 _u10_U3888  ( .A1(1'b0), .A2(_u10_n11901 ), .ZN(_u10_n15357 ) );
NAND2_X1 _u10_U3887  ( .A1(1'b0), .A2(_u10_n11878 ), .ZN(_u10_n15358 ) );
NAND2_X1 _u10_U3886  ( .A1(1'b0), .A2(_u10_n11851 ), .ZN(_u10_n15359 ) );
NAND2_X1 _u10_U3885  ( .A1(1'b0), .A2(_u10_n11829 ), .ZN(_u10_n15360 ) );
NAND4_X1 _u10_U3884  ( .A1(_u10_n15357 ), .A2(_u10_n15358 ), .A3(_u10_n15359 ), .A4(_u10_n15360 ), .ZN(_u10_n15346 ) );
NAND2_X1 _u10_U3883  ( .A1(1'b0), .A2(_u10_n11806 ), .ZN(_u10_n15353 ) );
NAND2_X1 _u10_U3882  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n15354 ) );
NAND2_X1 _u10_U3881  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n15355 ) );
NAND2_X1 _u10_U3880  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n15356 ) );
NAND4_X1 _u10_U3879  ( .A1(_u10_n15353 ), .A2(_u10_n15354 ), .A3(_u10_n15355 ), .A4(_u10_n15356 ), .ZN(_u10_n15347 ) );
NAND2_X1 _u10_U3878  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n15349 ) );
NAND2_X1 _u10_U3877  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n15350 ) );
NAND2_X1 _u10_U3876  ( .A1(1'b0), .A2(_u10_n11659 ), .ZN(_u10_n15351 ) );
NAND2_X1 _u10_U3875  ( .A1(1'b0), .A2(_u10_n11635 ), .ZN(_u10_n15352 ) );
NAND4_X1 _u10_U3874  ( .A1(_u10_n15349 ), .A2(_u10_n15350 ), .A3(_u10_n15351 ), .A4(_u10_n15352 ), .ZN(_u10_n15348 ) );
NOR4_X1 _u10_U3873  ( .A1(_u10_n15345 ), .A2(_u10_n15346 ), .A3(_u10_n15347 ), .A4(_u10_n15348 ), .ZN(_u10_n15344 ) );
NAND2_X1 _u10_U3872  ( .A1(_u10_n15343 ), .A2(_u10_n15344 ), .ZN(pointer[30]) );
NAND2_X1 _u10_U3871  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15339 ) );
NAND2_X1 _u10_U3870  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15340 ) );
NAND2_X1 _u10_U3869  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15341 ) );
NAND2_X1 _u10_U3868  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15342 ) );
NAND4_X1 _u10_U3867  ( .A1(_u10_n15339 ), .A2(_u10_n15340 ), .A3(_u10_n15341 ), .A4(_u10_n15342 ), .ZN(_u10_n15324 ) );
NAND2_X1 _u10_U3866  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15335 ) );
NAND2_X1 _u10_U3865  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15336 ) );
NAND2_X1 _u10_U3864  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15337 ) );
NAND2_X1 _u10_U3863  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15338 ) );
NAND4_X1 _u10_U3862  ( .A1(_u10_n15335 ), .A2(_u10_n15336 ), .A3(_u10_n15337 ), .A4(_u10_n15338 ), .ZN(_u10_n15325 ) );
NAND2_X1 _u10_U3861  ( .A1(1'b0), .A2(_u10_n12159 ), .ZN(_u10_n15331 ) );
NAND2_X1 _u10_U3860  ( .A1(1'b0), .A2(_u10_n12139 ), .ZN(_u10_n15332 ) );
NAND2_X1 _u10_U3859  ( .A1(1'b0), .A2(_u10_n12115 ), .ZN(_u10_n15333 ) );
NAND2_X1 _u10_U3858  ( .A1(1'b0), .A2(_u10_n12091 ), .ZN(_u10_n15334 ) );
NAND4_X1 _u10_U3857  ( .A1(_u10_n15331 ), .A2(_u10_n15332 ), .A3(_u10_n15333 ), .A4(_u10_n15334 ), .ZN(_u10_n15326 ) );
NAND2_X1 _u10_U3856  ( .A1(1'b0), .A2(_u10_n12063 ), .ZN(_u10_n15328 ) );
NAND2_X1 _u10_U3855  ( .A1(1'b0), .A2(_u10_n12039 ), .ZN(_u10_n15329 ) );
NAND2_X1 _u10_U3854  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15330 ) );
NAND3_X1 _u10_U3853  ( .A1(_u10_n15328 ), .A2(_u10_n15329 ), .A3(_u10_n15330 ), .ZN(_u10_n15327 ) );
NOR4_X1 _u10_U3852  ( .A1(_u10_n15324 ), .A2(_u10_n15325 ), .A3(_u10_n15326 ), .A4(_u10_n15327 ), .ZN(_u10_n15302 ) );
NAND2_X1 _u10_U3851  ( .A1(1'b0), .A2(_u10_n11999 ), .ZN(_u10_n15320 ) );
NAND2_X1 _u10_U3850  ( .A1(1'b0), .A2(_u10_n11974 ), .ZN(_u10_n15321 ) );
NAND2_X1 _u10_U3849  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n15322 ) );
NAND2_X1 _u10_U3848  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n15323 ) );
NAND4_X1 _u10_U3847  ( .A1(_u10_n15320 ), .A2(_u10_n15321 ), .A3(_u10_n15322 ), .A4(_u10_n15323 ), .ZN(_u10_n15304 ) );
NAND2_X1 _u10_U3846  ( .A1(1'b0), .A2(_u10_n11902 ), .ZN(_u10_n15316 ) );
NAND2_X1 _u10_U3845  ( .A1(1'b0), .A2(_u10_n11879 ), .ZN(_u10_n15317 ) );
NAND2_X1 _u10_U3844  ( .A1(1'b0), .A2(_u10_n11855 ), .ZN(_u10_n15318 ) );
NAND2_X1 _u10_U3843  ( .A1(1'b0), .A2(_u10_n11830 ), .ZN(_u10_n15319 ) );
NAND4_X1 _u10_U3842  ( .A1(_u10_n15316 ), .A2(_u10_n15317 ), .A3(_u10_n15318 ), .A4(_u10_n15319 ), .ZN(_u10_n15305 ) );
NAND2_X1 _u10_U3841  ( .A1(1'b0), .A2(_u10_n11807 ), .ZN(_u10_n15312 ) );
NAND2_X1 _u10_U3840  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n15313 ) );
NAND2_X1 _u10_U3839  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n15314 ) );
NAND2_X1 _u10_U3838  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n15315 ) );
NAND4_X1 _u10_U3837  ( .A1(_u10_n15312 ), .A2(_u10_n15313 ), .A3(_u10_n15314 ), .A4(_u10_n15315 ), .ZN(_u10_n15306 ) );
NAND2_X1 _u10_U3836  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n15308 ) );
NAND2_X1 _u10_U3835  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n15309 ) );
NAND2_X1 _u10_U3834  ( .A1(1'b0), .A2(_u10_n11663 ), .ZN(_u10_n15310 ) );
NAND2_X1 _u10_U3833  ( .A1(1'b0), .A2(_u10_n11639 ), .ZN(_u10_n15311 ) );
NAND4_X1 _u10_U3832  ( .A1(_u10_n15308 ), .A2(_u10_n15309 ), .A3(_u10_n15310 ), .A4(_u10_n15311 ), .ZN(_u10_n15307 ) );
NOR4_X1 _u10_U3831  ( .A1(_u10_n15304 ), .A2(_u10_n15305 ), .A3(_u10_n15306 ), .A4(_u10_n15307 ), .ZN(_u10_n15303 ) );
NAND2_X1 _u10_U3830  ( .A1(_u10_n15302 ), .A2(_u10_n15303 ), .ZN(pointer[31]) );
NAND2_X1 _u10_U3829  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15298 ) );
NAND2_X1 _u10_U3828  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15299 ) );
NAND2_X1 _u10_U3827  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15300 ) );
NAND2_X1 _u10_U3826  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15301 ) );
NAND4_X1 _u10_U3825  ( .A1(_u10_n15298 ), .A2(_u10_n15299 ), .A3(_u10_n15300 ), .A4(_u10_n15301 ), .ZN(_u10_n15283 ) );
NAND2_X1 _u10_U3824  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15294 ) );
NAND2_X1 _u10_U3823  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15295 ) );
NAND2_X1 _u10_U3822  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15296 ) );
NAND2_X1 _u10_U3821  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15297 ) );
NAND4_X1 _u10_U3820  ( .A1(_u10_n15294 ), .A2(_u10_n15295 ), .A3(_u10_n15296 ), .A4(_u10_n15297 ), .ZN(_u10_n15284 ) );
NAND2_X1 _u10_U3819  ( .A1(1'b0), .A2(_u10_n12163 ), .ZN(_u10_n15290 ) );
NAND2_X1 _u10_U3818  ( .A1(1'b0), .A2(_u10_n12136 ), .ZN(_u10_n15291 ) );
NAND2_X1 _u10_U3817  ( .A1(1'b0), .A2(_u10_n12112 ), .ZN(_u10_n15292 ) );
NAND2_X1 _u10_U3816  ( .A1(1'b0), .A2(_u10_n12088 ), .ZN(_u10_n15293 ) );
NAND4_X1 _u10_U3815  ( .A1(_u10_n15290 ), .A2(_u10_n15291 ), .A3(_u10_n15292 ), .A4(_u10_n15293 ), .ZN(_u10_n15285 ) );
NAND2_X1 _u10_U3814  ( .A1(1'b0), .A2(_u10_n12065 ), .ZN(_u10_n15287 ) );
NAND2_X1 _u10_U3813  ( .A1(1'b0), .A2(_u10_n12041 ), .ZN(_u10_n15288 ) );
NAND2_X1 _u10_U3812  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15289 ) );
NAND3_X1 _u10_U3811  ( .A1(_u10_n15287 ), .A2(_u10_n15288 ), .A3(_u10_n15289 ), .ZN(_u10_n15286 ) );
NOR4_X1 _u10_U3810  ( .A1(_u10_n15283 ), .A2(_u10_n15284 ), .A3(_u10_n15285 ), .A4(_u10_n15286 ), .ZN(_u10_n15261 ) );
NAND2_X1 _u10_U3809  ( .A1(1'b0), .A2(_u10_n12396 ), .ZN(_u10_n15279 ) );
NAND2_X1 _u10_U3808  ( .A1(1'b0), .A2(_u10_n12395 ), .ZN(_u10_n15280 ) );
NAND2_X1 _u10_U3807  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n15281 ) );
NAND2_X1 _u10_U3806  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n15282 ) );
NAND4_X1 _u10_U3805  ( .A1(_u10_n15279 ), .A2(_u10_n15280 ), .A3(_u10_n15281 ), .A4(_u10_n15282 ), .ZN(_u10_n15263 ) );
NAND2_X1 _u10_U3804  ( .A1(1'b0), .A2(_u10_n11898 ), .ZN(_u10_n15275 ) );
NAND2_X1 _u10_U3803  ( .A1(1'b0), .A2(_u10_n12387 ), .ZN(_u10_n15276 ) );
NAND2_X1 _u10_U3802  ( .A1(1'b0), .A2(_u10_n12386 ), .ZN(_u10_n15277 ) );
NAND2_X1 _u10_U3801  ( .A1(1'b0), .A2(_u10_n11826 ), .ZN(_u10_n15278 ) );
NAND4_X1 _u10_U3800  ( .A1(_u10_n15275 ), .A2(_u10_n15276 ), .A3(_u10_n15277 ), .A4(_u10_n15278 ), .ZN(_u10_n15264 ) );
NAND2_X1 _u10_U3799  ( .A1(1'b0), .A2(_u10_n12380 ), .ZN(_u10_n15271 ) );
NAND2_X1 _u10_U3798  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n15272 ) );
NAND2_X1 _u10_U3797  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n15273 ) );
NAND2_X1 _u10_U3796  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n15274 ) );
NAND4_X1 _u10_U3795  ( .A1(_u10_n15271 ), .A2(_u10_n15272 ), .A3(_u10_n15273 ), .A4(_u10_n15274 ), .ZN(_u10_n15265 ) );
NAND2_X1 _u10_U3794  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n15267 ) );
NAND2_X1 _u10_U3793  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n15268 ) );
NAND2_X1 _u10_U3792  ( .A1(1'b0), .A2(_u10_n12370 ), .ZN(_u10_n15269 ) );
NAND2_X1 _u10_U3791  ( .A1(1'b0), .A2(_u10_n12369 ), .ZN(_u10_n15270 ) );
NAND4_X1 _u10_U3790  ( .A1(_u10_n15267 ), .A2(_u10_n15268 ), .A3(_u10_n15269 ), .A4(_u10_n15270 ), .ZN(_u10_n15266 ) );
NOR4_X1 _u10_U3789  ( .A1(_u10_n15263 ), .A2(_u10_n15264 ), .A3(_u10_n15265 ), .A4(_u10_n15266 ), .ZN(_u10_n15262 ) );
NAND2_X1 _u10_U3788  ( .A1(_u10_n15261 ), .A2(_u10_n15262 ), .ZN(pointer[3]));
NAND2_X1 _u10_U3787  ( .A1(1'b0), .A2(_u10_n12345 ), .ZN(_u10_n15257 ) );
NAND2_X1 _u10_U3786  ( .A1(1'b0), .A2(_u10_n12321 ), .ZN(_u10_n15258 ) );
NAND2_X1 _u10_U3785  ( .A1(1'b0), .A2(_u10_n12298 ), .ZN(_u10_n15259 ) );
NAND2_X1 _u10_U3784  ( .A1(1'b0), .A2(_u10_n12274 ), .ZN(_u10_n15260 ) );
NAND4_X1 _u10_U3783  ( .A1(_u10_n15257 ), .A2(_u10_n15258 ), .A3(_u10_n15259 ), .A4(_u10_n15260 ), .ZN(_u10_n15242 ) );
NAND2_X1 _u10_U3782  ( .A1(1'b0), .A2(_u10_n12249 ), .ZN(_u10_n15253 ) );
NAND2_X1 _u10_U3781  ( .A1(1'b0), .A2(_u10_n12225 ), .ZN(_u10_n15254 ) );
NAND2_X1 _u10_U3780  ( .A1(1'b0), .A2(_u10_n12199 ), .ZN(_u10_n15255 ) );
NAND2_X1 _u10_U3779  ( .A1(1'b0), .A2(_u10_n12177 ), .ZN(_u10_n15256 ) );
NAND4_X1 _u10_U3778  ( .A1(_u10_n15253 ), .A2(_u10_n15254 ), .A3(_u10_n15255 ), .A4(_u10_n15256 ), .ZN(_u10_n15243 ) );
NAND2_X1 _u10_U3777  ( .A1(1'b0), .A2(_u10_n12163 ), .ZN(_u10_n15249 ) );
NAND2_X1 _u10_U3776  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n15250 ) );
NAND2_X1 _u10_U3775  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n15251 ) );
NAND2_X1 _u10_U3774  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n15252 ) );
NAND4_X1 _u10_U3773  ( .A1(_u10_n15249 ), .A2(_u10_n15250 ), .A3(_u10_n15251 ), .A4(_u10_n15252 ), .ZN(_u10_n15244 ) );
NAND2_X1 _u10_U3772  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n15246 ) );
NAND2_X1 _u10_U3771  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n15247 ) );
NAND2_X1 _u10_U3770  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15248 ) );
NAND3_X1 _u10_U3769  ( .A1(_u10_n15246 ), .A2(_u10_n15247 ), .A3(_u10_n15248 ), .ZN(_u10_n15245 ) );
NOR4_X1 _u10_U3768  ( .A1(_u10_n15242 ), .A2(_u10_n15243 ), .A3(_u10_n15244 ), .A4(_u10_n15245 ), .ZN(_u10_n15220 ) );
NAND2_X1 _u10_U3767  ( .A1(1'b0), .A2(_u10_n11993 ), .ZN(_u10_n15238 ) );
NAND2_X1 _u10_U3766  ( .A1(1'b0), .A2(_u10_n11973 ), .ZN(_u10_n15239 ) );
NAND2_X1 _u10_U3765  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n15240 ) );
NAND2_X1 _u10_U3764  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n15241 ) );
NAND4_X1 _u10_U3763  ( .A1(_u10_n15238 ), .A2(_u10_n15239 ), .A3(_u10_n15240 ), .A4(_u10_n15241 ), .ZN(_u10_n15222 ) );
NAND2_X1 _u10_U3762  ( .A1(1'b0), .A2(_u10_n11903 ), .ZN(_u10_n15234 ) );
NAND2_X1 _u10_U3761  ( .A1(1'b0), .A2(_u10_n11873 ), .ZN(_u10_n15235 ) );
NAND2_X1 _u10_U3760  ( .A1(1'b0), .A2(_u10_n11849 ), .ZN(_u10_n15236 ) );
NAND2_X1 _u10_U3759  ( .A1(1'b0), .A2(_u10_n11831 ), .ZN(_u10_n15237 ) );
NAND4_X1 _u10_U3758  ( .A1(_u10_n15234 ), .A2(_u10_n15235 ), .A3(_u10_n15236 ), .A4(_u10_n15237 ), .ZN(_u10_n15223 ) );
NAND2_X1 _u10_U3757  ( .A1(1'b0), .A2(_u10_n11801 ), .ZN(_u10_n15230 ) );
NAND2_X1 _u10_U3756  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n15231 ) );
NAND2_X1 _u10_U3755  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n15232 ) );
NAND2_X1 _u10_U3754  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n15233 ) );
NAND4_X1 _u10_U3753  ( .A1(_u10_n15230 ), .A2(_u10_n15231 ), .A3(_u10_n15232 ), .A4(_u10_n15233 ), .ZN(_u10_n15224 ) );
NAND2_X1 _u10_U3752  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n15226 ) );
NAND2_X1 _u10_U3751  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n15227 ) );
NAND2_X1 _u10_U3750  ( .A1(1'b0), .A2(_u10_n11657 ), .ZN(_u10_n15228 ) );
NAND2_X1 _u10_U3749  ( .A1(1'b0), .A2(_u10_n11633 ), .ZN(_u10_n15229 ) );
NAND4_X1 _u10_U3748  ( .A1(_u10_n15226 ), .A2(_u10_n15227 ), .A3(_u10_n15228 ), .A4(_u10_n15229 ), .ZN(_u10_n15225 ) );
NOR4_X1 _u10_U3747  ( .A1(_u10_n15222 ), .A2(_u10_n15223 ), .A3(_u10_n15224 ), .A4(_u10_n15225 ), .ZN(_u10_n15221 ) );
NAND2_X1 _u10_U3746  ( .A1(_u10_n15220 ), .A2(_u10_n15221 ), .ZN(pointer[4]));
NAND2_X1 _u10_U3745  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n15216 ) );
NAND2_X1 _u10_U3744  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n15217 ) );
NAND2_X1 _u10_U3743  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n15218 ) );
NAND2_X1 _u10_U3742  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n15219 ) );
NAND4_X1 _u10_U3741  ( .A1(_u10_n15216 ), .A2(_u10_n15217 ), .A3(_u10_n15218 ), .A4(_u10_n15219 ), .ZN(_u10_n15201 ) );
NAND2_X1 _u10_U3740  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n15212 ) );
NAND2_X1 _u10_U3739  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n15213 ) );
NAND2_X1 _u10_U3738  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n15214 ) );
NAND2_X1 _u10_U3737  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n15215 ) );
NAND4_X1 _u10_U3736  ( .A1(_u10_n15212 ), .A2(_u10_n15213 ), .A3(_u10_n15214 ), .A4(_u10_n15215 ), .ZN(_u10_n15202 ) );
NAND2_X1 _u10_U3735  ( .A1(1'b0), .A2(_u10_n12162 ), .ZN(_u10_n15208 ) );
NAND2_X1 _u10_U3734  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n15209 ) );
NAND2_X1 _u10_U3733  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n15210 ) );
NAND2_X1 _u10_U3732  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n15211 ) );
NAND4_X1 _u10_U3731  ( .A1(_u10_n15208 ), .A2(_u10_n15209 ), .A3(_u10_n15210 ), .A4(_u10_n15211 ), .ZN(_u10_n15203 ) );
NAND2_X1 _u10_U3730  ( .A1(1'b0), .A2(_u10_n12406 ), .ZN(_u10_n15205 ) );
NAND2_X1 _u10_U3729  ( .A1(1'b0), .A2(_u10_n12405 ), .ZN(_u10_n15206 ) );
NAND2_X1 _u10_U3728  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15207 ) );
NAND3_X1 _u10_U3727  ( .A1(_u10_n15205 ), .A2(_u10_n15206 ), .A3(_u10_n15207 ), .ZN(_u10_n15204 ) );
NOR4_X1 _u10_U3726  ( .A1(_u10_n15201 ), .A2(_u10_n15202 ), .A3(_u10_n15203 ), .A4(_u10_n15204 ), .ZN(_u10_n15179 ) );
NAND2_X1 _u10_U3725  ( .A1(1'b0), .A2(_u10_n11996 ), .ZN(_u10_n15197 ) );
NAND2_X1 _u10_U3724  ( .A1(1'b0), .A2(_u10_n11969 ), .ZN(_u10_n15198 ) );
NAND2_X1 _u10_U3723  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n15199 ) );
NAND2_X1 _u10_U3722  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n15200 ) );
NAND4_X1 _u10_U3721  ( .A1(_u10_n15197 ), .A2(_u10_n15198 ), .A3(_u10_n15199 ), .A4(_u10_n15200 ), .ZN(_u10_n15181 ) );
NAND2_X1 _u10_U3720  ( .A1(1'b0), .A2(_u10_n11899 ), .ZN(_u10_n15193 ) );
NAND2_X1 _u10_U3719  ( .A1(1'b0), .A2(_u10_n11876 ), .ZN(_u10_n15194 ) );
NAND2_X1 _u10_U3718  ( .A1(1'b0), .A2(_u10_n11852 ), .ZN(_u10_n15195 ) );
NAND2_X1 _u10_U3717  ( .A1(1'b0), .A2(_u10_n11827 ), .ZN(_u10_n15196 ) );
NAND4_X1 _u10_U3716  ( .A1(_u10_n15193 ), .A2(_u10_n15194 ), .A3(_u10_n15195 ), .A4(_u10_n15196 ), .ZN(_u10_n15182 ) );
NAND2_X1 _u10_U3715  ( .A1(1'b0), .A2(_u10_n11804 ), .ZN(_u10_n15189 ) );
NAND2_X1 _u10_U3714  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n15190 ) );
NAND2_X1 _u10_U3713  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n15191 ) );
NAND2_X1 _u10_U3712  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n15192 ) );
NAND4_X1 _u10_U3711  ( .A1(_u10_n15189 ), .A2(_u10_n15190 ), .A3(_u10_n15191 ), .A4(_u10_n15192 ), .ZN(_u10_n15183 ) );
NAND2_X1 _u10_U3710  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n15185 ) );
NAND2_X1 _u10_U3709  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n15186 ) );
NAND2_X1 _u10_U3708  ( .A1(1'b0), .A2(_u10_n11660 ), .ZN(_u10_n15187 ) );
NAND2_X1 _u10_U3707  ( .A1(1'b0), .A2(_u10_n11636 ), .ZN(_u10_n15188 ) );
NAND4_X1 _u10_U3706  ( .A1(_u10_n15185 ), .A2(_u10_n15186 ), .A3(_u10_n15187 ), .A4(_u10_n15188 ), .ZN(_u10_n15184 ) );
NOR4_X1 _u10_U3705  ( .A1(_u10_n15181 ), .A2(_u10_n15182 ), .A3(_u10_n15183 ), .A4(_u10_n15184 ), .ZN(_u10_n15180 ) );
NAND2_X1 _u10_U3704  ( .A1(_u10_n15179 ), .A2(_u10_n15180 ), .ZN(pointer[5]));
NAND2_X1 _u10_U3703  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n15175 ) );
NAND2_X1 _u10_U3702  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n15176 ) );
NAND2_X1 _u10_U3701  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n15177 ) );
NAND2_X1 _u10_U3700  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n15178 ) );
NAND4_X1 _u10_U3699  ( .A1(_u10_n15175 ), .A2(_u10_n15176 ), .A3(_u10_n15177 ), .A4(_u10_n15178 ), .ZN(_u10_n15160 ) );
NAND2_X1 _u10_U3698  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n15171 ) );
NAND2_X1 _u10_U3697  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n15172 ) );
NAND2_X1 _u10_U3696  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n15173 ) );
NAND2_X1 _u10_U3695  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n15174 ) );
NAND4_X1 _u10_U3694  ( .A1(_u10_n15171 ), .A2(_u10_n15172 ), .A3(_u10_n15173 ), .A4(_u10_n15174 ), .ZN(_u10_n15161 ) );
NAND2_X1 _u10_U3693  ( .A1(1'b0), .A2(_u10_n12159 ), .ZN(_u10_n15167 ) );
NAND2_X1 _u10_U3692  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n15168 ) );
NAND2_X1 _u10_U3691  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n15169 ) );
NAND2_X1 _u10_U3690  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n15170 ) );
NAND4_X1 _u10_U3689  ( .A1(_u10_n15167 ), .A2(_u10_n15168 ), .A3(_u10_n15169 ), .A4(_u10_n15170 ), .ZN(_u10_n15162 ) );
NAND2_X1 _u10_U3688  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n15164 ) );
NAND2_X1 _u10_U3687  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n15165 ) );
NAND2_X1 _u10_U3686  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15166 ) );
NAND3_X1 _u10_U3685  ( .A1(_u10_n15164 ), .A2(_u10_n15165 ), .A3(_u10_n15166 ), .ZN(_u10_n15163 ) );
NOR4_X1 _u10_U3684  ( .A1(_u10_n15160 ), .A2(_u10_n15161 ), .A3(_u10_n15162 ), .A4(_u10_n15163 ), .ZN(_u10_n15138 ) );
NAND2_X1 _u10_U3683  ( .A1(1'b0), .A2(_u10_n11997 ), .ZN(_u10_n15156 ) );
NAND2_X1 _u10_U3682  ( .A1(1'b0), .A2(_u10_n11972 ), .ZN(_u10_n15157 ) );
NAND2_X1 _u10_U3681  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n15158 ) );
NAND2_X1 _u10_U3680  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n15159 ) );
NAND4_X1 _u10_U3679  ( .A1(_u10_n15156 ), .A2(_u10_n15157 ), .A3(_u10_n15158 ), .A4(_u10_n15159 ), .ZN(_u10_n15140 ) );
NAND2_X1 _u10_U3678  ( .A1(1'b0), .A2(_u10_n12388 ), .ZN(_u10_n15152 ) );
NAND2_X1 _u10_U3677  ( .A1(1'b0), .A2(_u10_n11877 ), .ZN(_u10_n15153 ) );
NAND2_X1 _u10_U3676  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n15154 ) );
NAND2_X1 _u10_U3675  ( .A1(1'b0), .A2(_u10_n12385 ), .ZN(_u10_n15155 ) );
NAND4_X1 _u10_U3674  ( .A1(_u10_n15152 ), .A2(_u10_n15153 ), .A3(_u10_n15154 ), .A4(_u10_n15155 ), .ZN(_u10_n15141 ) );
NAND2_X1 _u10_U3673  ( .A1(1'b0), .A2(_u10_n11805 ), .ZN(_u10_n15148 ) );
NAND2_X1 _u10_U3672  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n15149 ) );
NAND2_X1 _u10_U3671  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n15150 ) );
NAND2_X1 _u10_U3670  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n15151 ) );
NAND4_X1 _u10_U3669  ( .A1(_u10_n15148 ), .A2(_u10_n15149 ), .A3(_u10_n15150 ), .A4(_u10_n15151 ), .ZN(_u10_n15142 ) );
NAND2_X1 _u10_U3668  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n15144 ) );
NAND2_X1 _u10_U3667  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n15145 ) );
NAND2_X1 _u10_U3666  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n15146 ) );
NAND2_X1 _u10_U3665  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n15147 ) );
NAND4_X1 _u10_U3664  ( .A1(_u10_n15144 ), .A2(_u10_n15145 ), .A3(_u10_n15146 ), .A4(_u10_n15147 ), .ZN(_u10_n15143 ) );
NOR4_X1 _u10_U3663  ( .A1(_u10_n15140 ), .A2(_u10_n15141 ), .A3(_u10_n15142 ), .A4(_u10_n15143 ), .ZN(_u10_n15139 ) );
NAND2_X1 _u10_U3662  ( .A1(_u10_n15138 ), .A2(_u10_n15139 ), .ZN(pointer[6]));
NAND2_X1 _u10_U3661  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n15134 ) );
NAND2_X1 _u10_U3660  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n15135 ) );
NAND2_X1 _u10_U3659  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n15136 ) );
NAND2_X1 _u10_U3658  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n15137 ) );
NAND4_X1 _u10_U3657  ( .A1(_u10_n15134 ), .A2(_u10_n15135 ), .A3(_u10_n15136 ), .A4(_u10_n15137 ), .ZN(_u10_n15119 ) );
NAND2_X1 _u10_U3656  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n15130 ) );
NAND2_X1 _u10_U3655  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n15131 ) );
NAND2_X1 _u10_U3654  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n15132 ) );
NAND2_X1 _u10_U3653  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n15133 ) );
NAND4_X1 _u10_U3652  ( .A1(_u10_n15130 ), .A2(_u10_n15131 ), .A3(_u10_n15132 ), .A4(_u10_n15133 ), .ZN(_u10_n15120 ) );
NAND2_X1 _u10_U3651  ( .A1(1'b0), .A2(_u10_n12160 ), .ZN(_u10_n15126 ) );
NAND2_X1 _u10_U3650  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n15127 ) );
NAND2_X1 _u10_U3649  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n15128 ) );
NAND2_X1 _u10_U3648  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n15129 ) );
NAND4_X1 _u10_U3647  ( .A1(_u10_n15126 ), .A2(_u10_n15127 ), .A3(_u10_n15128 ), .A4(_u10_n15129 ), .ZN(_u10_n15121 ) );
NAND2_X1 _u10_U3646  ( .A1(1'b0), .A2(_u10_n12068 ), .ZN(_u10_n15123 ) );
NAND2_X1 _u10_U3645  ( .A1(1'b0), .A2(_u10_n12044 ), .ZN(_u10_n15124 ) );
NAND2_X1 _u10_U3644  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15125 ) );
NAND3_X1 _u10_U3643  ( .A1(_u10_n15123 ), .A2(_u10_n15124 ), .A3(_u10_n15125 ), .ZN(_u10_n15122 ) );
NOR4_X1 _u10_U3642  ( .A1(_u10_n15119 ), .A2(_u10_n15120 ), .A3(_u10_n15121 ), .A4(_u10_n15122 ), .ZN(_u10_n15097 ) );
NAND2_X1 _u10_U3641  ( .A1(1'b0), .A2(_u10_n11999 ), .ZN(_u10_n15115 ) );
NAND2_X1 _u10_U3640  ( .A1(1'b0), .A2(_u10_n11972 ), .ZN(_u10_n15116 ) );
NAND2_X1 _u10_U3639  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n15117 ) );
NAND2_X1 _u10_U3638  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n15118 ) );
NAND4_X1 _u10_U3637  ( .A1(_u10_n15115 ), .A2(_u10_n15116 ), .A3(_u10_n15117 ), .A4(_u10_n15118 ), .ZN(_u10_n15099 ) );
NAND2_X1 _u10_U3636  ( .A1(1'b0), .A2(_u10_n11897 ), .ZN(_u10_n15111 ) );
NAND2_X1 _u10_U3635  ( .A1(1'b0), .A2(_u10_n11879 ), .ZN(_u10_n15112 ) );
NAND2_X1 _u10_U3634  ( .A1(1'b0), .A2(_u10_n11854 ), .ZN(_u10_n15113 ) );
NAND2_X1 _u10_U3633  ( .A1(1'b0), .A2(_u10_n11825 ), .ZN(_u10_n15114 ) );
NAND4_X1 _u10_U3632  ( .A1(_u10_n15111 ), .A2(_u10_n15112 ), .A3(_u10_n15113 ), .A4(_u10_n15114 ), .ZN(_u10_n15100 ) );
NAND2_X1 _u10_U3631  ( .A1(1'b0), .A2(_u10_n11807 ), .ZN(_u10_n15107 ) );
NAND2_X1 _u10_U3630  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n15108 ) );
NAND2_X1 _u10_U3629  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n15109 ) );
NAND2_X1 _u10_U3628  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n15110 ) );
NAND4_X1 _u10_U3627  ( .A1(_u10_n15107 ), .A2(_u10_n15108 ), .A3(_u10_n15109 ), .A4(_u10_n15110 ), .ZN(_u10_n15101 ) );
NAND2_X1 _u10_U3626  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n15103 ) );
NAND2_X1 _u10_U3625  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n15104 ) );
NAND2_X1 _u10_U3624  ( .A1(1'b0), .A2(_u10_n11662 ), .ZN(_u10_n15105 ) );
NAND2_X1 _u10_U3623  ( .A1(1'b0), .A2(_u10_n11638 ), .ZN(_u10_n15106 ) );
NAND4_X1 _u10_U3622  ( .A1(_u10_n15103 ), .A2(_u10_n15104 ), .A3(_u10_n15105 ), .A4(_u10_n15106 ), .ZN(_u10_n15102 ) );
NOR4_X1 _u10_U3621  ( .A1(_u10_n15099 ), .A2(_u10_n15100 ), .A3(_u10_n15101 ), .A4(_u10_n15102 ), .ZN(_u10_n15098 ) );
NAND2_X1 _u10_U3620  ( .A1(_u10_n15097 ), .A2(_u10_n15098 ), .ZN(pointer[7]));
NAND2_X1 _u10_U3619  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n15093 ) );
NAND2_X1 _u10_U3618  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n15094 ) );
NAND2_X1 _u10_U3617  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n15095 ) );
NAND2_X1 _u10_U3616  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n15096 ) );
NAND4_X1 _u10_U3615  ( .A1(_u10_n15093 ), .A2(_u10_n15094 ), .A3(_u10_n15095 ), .A4(_u10_n15096 ), .ZN(_u10_n15078 ) );
NAND2_X1 _u10_U3614  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n15089 ) );
NAND2_X1 _u10_U3613  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n15090 ) );
NAND2_X1 _u10_U3612  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n15091 ) );
NAND2_X1 _u10_U3611  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n15092 ) );
NAND4_X1 _u10_U3610  ( .A1(_u10_n15089 ), .A2(_u10_n15090 ), .A3(_u10_n15091 ), .A4(_u10_n15092 ), .ZN(_u10_n15079 ) );
NAND2_X1 _u10_U3609  ( .A1(1'b0), .A2(_u10_n12414 ), .ZN(_u10_n15085 ) );
NAND2_X1 _u10_U3608  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n15086 ) );
NAND2_X1 _u10_U3607  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n15087 ) );
NAND2_X1 _u10_U3606  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n15088 ) );
NAND4_X1 _u10_U3605  ( .A1(_u10_n15085 ), .A2(_u10_n15086 ), .A3(_u10_n15087 ), .A4(_u10_n15088 ), .ZN(_u10_n15080 ) );
NAND2_X1 _u10_U3604  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n15082 ) );
NAND2_X1 _u10_U3603  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n15083 ) );
NAND2_X1 _u10_U3602  ( .A1(1'b0), .A2(_u10_n12014 ), .ZN(_u10_n15084 ) );
NAND3_X1 _u10_U3601  ( .A1(_u10_n15082 ), .A2(_u10_n15083 ), .A3(_u10_n15084 ), .ZN(_u10_n15081 ) );
NOR4_X1 _u10_U3600  ( .A1(_u10_n15078 ), .A2(_u10_n15079 ), .A3(_u10_n15080 ), .A4(_u10_n15081 ), .ZN(_u10_n15056 ) );
NAND2_X1 _u10_U3599  ( .A1(1'b0), .A2(_u10_n11994 ), .ZN(_u10_n15074 ) );
NAND2_X1 _u10_U3598  ( .A1(1'b0), .A2(_u10_n11975 ), .ZN(_u10_n15075 ) );
NAND2_X1 _u10_U3597  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n15076 ) );
NAND2_X1 _u10_U3596  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n15077 ) );
NAND4_X1 _u10_U3595  ( .A1(_u10_n15074 ), .A2(_u10_n15075 ), .A3(_u10_n15076 ), .A4(_u10_n15077 ), .ZN(_u10_n15058 ) );
NAND2_X1 _u10_U3594  ( .A1(1'b0), .A2(_u10_n11900 ), .ZN(_u10_n15070 ) );
NAND2_X1 _u10_U3593  ( .A1(1'b0), .A2(_u10_n11874 ), .ZN(_u10_n15071 ) );
NAND2_X1 _u10_U3592  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n15072 ) );
NAND2_X1 _u10_U3591  ( .A1(1'b0), .A2(_u10_n11828 ), .ZN(_u10_n15073 ) );
NAND4_X1 _u10_U3590  ( .A1(_u10_n15070 ), .A2(_u10_n15071 ), .A3(_u10_n15072 ), .A4(_u10_n15073 ), .ZN(_u10_n15059 ) );
NAND2_X1 _u10_U3589  ( .A1(1'b0), .A2(_u10_n11802 ), .ZN(_u10_n15066 ) );
NAND2_X1 _u10_U3588  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n15067 ) );
NAND2_X1 _u10_U3587  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n15068 ) );
NAND2_X1 _u10_U3586  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n15069 ) );
NAND4_X1 _u10_U3585  ( .A1(_u10_n15066 ), .A2(_u10_n15067 ), .A3(_u10_n15068 ), .A4(_u10_n15069 ), .ZN(_u10_n15060 ) );
NAND2_X1 _u10_U3584  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n15062 ) );
NAND2_X1 _u10_U3583  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n15063 ) );
NAND2_X1 _u10_U3582  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n15064 ) );
NAND2_X1 _u10_U3581  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n15065 ) );
NAND4_X1 _u10_U3580  ( .A1(_u10_n15062 ), .A2(_u10_n15063 ), .A3(_u10_n15064 ), .A4(_u10_n15065 ), .ZN(_u10_n15061 ) );
NOR4_X1 _u10_U3579  ( .A1(_u10_n15058 ), .A2(_u10_n15059 ), .A3(_u10_n15060 ), .A4(_u10_n15061 ), .ZN(_u10_n15057 ) );
NAND2_X1 _u10_U3578  ( .A1(_u10_n15056 ), .A2(_u10_n15057 ), .ZN(pointer[8]));
NAND2_X1 _u10_U3577  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n15052 ) );
NAND2_X1 _u10_U3576  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n15053 ) );
NAND2_X1 _u10_U3575  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n15054 ) );
NAND2_X1 _u10_U3574  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n15055 ) );
NAND4_X1 _u10_U3573  ( .A1(_u10_n15052 ), .A2(_u10_n15053 ), .A3(_u10_n15054 ), .A4(_u10_n15055 ), .ZN(_u10_n15037 ) );
NAND2_X1 _u10_U3572  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n15048 ) );
NAND2_X1 _u10_U3571  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n15049 ) );
NAND2_X1 _u10_U3570  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n15050 ) );
NAND2_X1 _u10_U3569  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n15051 ) );
NAND4_X1 _u10_U3568  ( .A1(_u10_n15048 ), .A2(_u10_n15049 ), .A3(_u10_n15050 ), .A4(_u10_n15051 ), .ZN(_u10_n15038 ) );
NAND2_X1 _u10_U3567  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n15044 ) );
NAND2_X1 _u10_U3566  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n15045 ) );
NAND2_X1 _u10_U3565  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n15046 ) );
NAND2_X1 _u10_U3564  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n15047 ) );
NAND4_X1 _u10_U3563  ( .A1(_u10_n15044 ), .A2(_u10_n15045 ), .A3(_u10_n15046 ), .A4(_u10_n15047 ), .ZN(_u10_n15039 ) );
NAND2_X1 _u10_U3562  ( .A1(1'b0), .A2(_u10_n12067 ), .ZN(_u10_n15041 ) );
NAND2_X1 _u10_U3561  ( .A1(1'b0), .A2(_u10_n12043 ), .ZN(_u10_n15042 ) );
NAND2_X1 _u10_U3560  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n15043 ) );
NAND3_X1 _u10_U3559  ( .A1(_u10_n15041 ), .A2(_u10_n15042 ), .A3(_u10_n15043 ), .ZN(_u10_n15040 ) );
NOR4_X1 _u10_U3558  ( .A1(_u10_n15037 ), .A2(_u10_n15038 ), .A3(_u10_n15039 ), .A4(_u10_n15040 ), .ZN(_u10_n15015 ) );
NAND2_X1 _u10_U3557  ( .A1(1'b0), .A2(_u10_n11995 ), .ZN(_u10_n15033 ) );
NAND2_X1 _u10_U3556  ( .A1(1'b0), .A2(_u10_n11971 ), .ZN(_u10_n15034 ) );
NAND2_X1 _u10_U3555  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n15035 ) );
NAND2_X1 _u10_U3554  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n15036 ) );
NAND4_X1 _u10_U3553  ( .A1(_u10_n15033 ), .A2(_u10_n15034 ), .A3(_u10_n15035 ), .A4(_u10_n15036 ), .ZN(_u10_n15017 ) );
NAND2_X1 _u10_U3552  ( .A1(1'b0), .A2(_u10_n11901 ), .ZN(_u10_n15029 ) );
NAND2_X1 _u10_U3551  ( .A1(1'b0), .A2(_u10_n11875 ), .ZN(_u10_n15030 ) );
NAND2_X1 _u10_U3550  ( .A1(1'b0), .A2(_u10_n11850 ), .ZN(_u10_n15031 ) );
NAND2_X1 _u10_U3549  ( .A1(1'b0), .A2(_u10_n11829 ), .ZN(_u10_n15032 ) );
NAND4_X1 _u10_U3548  ( .A1(_u10_n15029 ), .A2(_u10_n15030 ), .A3(_u10_n15031 ), .A4(_u10_n15032 ), .ZN(_u10_n15018 ) );
NAND2_X1 _u10_U3547  ( .A1(1'b0), .A2(_u10_n11803 ), .ZN(_u10_n15025 ) );
NAND2_X1 _u10_U3546  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n15026 ) );
NAND2_X1 _u10_U3545  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n15027 ) );
NAND2_X1 _u10_U3544  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n15028 ) );
NAND4_X1 _u10_U3543  ( .A1(_u10_n15025 ), .A2(_u10_n15026 ), .A3(_u10_n15027 ), .A4(_u10_n15028 ), .ZN(_u10_n15019 ) );
NAND2_X1 _u10_U3542  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n15021 ) );
NAND2_X1 _u10_U3541  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n15022 ) );
NAND2_X1 _u10_U3540  ( .A1(1'b0), .A2(_u10_n11658 ), .ZN(_u10_n15023 ) );
NAND2_X1 _u10_U3539  ( .A1(1'b0), .A2(_u10_n11634 ), .ZN(_u10_n15024 ) );
NAND4_X1 _u10_U3538  ( .A1(_u10_n15021 ), .A2(_u10_n15022 ), .A3(_u10_n15023 ), .A4(_u10_n15024 ), .ZN(_u10_n15020 ) );
NOR4_X1 _u10_U3537  ( .A1(_u10_n15017 ), .A2(_u10_n15018 ), .A3(_u10_n15019 ), .A4(_u10_n15020 ), .ZN(_u10_n15016 ) );
NAND2_X1 _u10_U3536  ( .A1(_u10_n15015 ), .A2(_u10_n15016 ), .ZN(pointer[9]));
NAND2_X1 _u10_U3535  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n15011 ) );
NAND2_X1 _u10_U3534  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n15012 ) );
NAND2_X1 _u10_U3533  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n15013 ) );
NAND2_X1 _u10_U3532  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n15014 ) );
NAND4_X1 _u10_U3531  ( .A1(_u10_n15011 ), .A2(_u10_n15012 ), .A3(_u10_n15013 ), .A4(_u10_n15014 ), .ZN(_u10_n14996 ) );
NAND2_X1 _u10_U3530  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n15007 ) );
NAND2_X1 _u10_U3529  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n15008 ) );
NAND2_X1 _u10_U3528  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n15009 ) );
NAND2_X1 _u10_U3527  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n15010 ) );
NAND4_X1 _u10_U3526  ( .A1(_u10_n15007 ), .A2(_u10_n15008 ), .A3(_u10_n15009 ), .A4(_u10_n15010 ), .ZN(_u10_n14997 ) );
NAND2_X1 _u10_U3525  ( .A1(1'b0), .A2(_u10_n12160 ), .ZN(_u10_n15003 ) );
NAND2_X1 _u10_U3524  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n15004 ) );
NAND2_X1 _u10_U3523  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n15005 ) );
NAND2_X1 _u10_U3522  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n15006 ) );
NAND4_X1 _u10_U3521  ( .A1(_u10_n15003 ), .A2(_u10_n15004 ), .A3(_u10_n15005 ), .A4(_u10_n15006 ), .ZN(_u10_n14998 ) );
NAND2_X1 _u10_U3520  ( .A1(1'b0), .A2(_u10_n12066 ), .ZN(_u10_n15000 ) );
NAND2_X1 _u10_U3519  ( .A1(1'b0), .A2(_u10_n12042 ), .ZN(_u10_n15001 ) );
NAND2_X1 _u10_U3518  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n15002 ) );
NAND3_X1 _u10_U3517  ( .A1(_u10_n15000 ), .A2(_u10_n15001 ), .A3(_u10_n15002 ), .ZN(_u10_n14999 ) );
NOR4_X1 _u10_U3516  ( .A1(_u10_n14996 ), .A2(_u10_n14997 ), .A3(_u10_n14998 ), .A4(_u10_n14999 ), .ZN(_u10_n14974 ) );
NAND2_X1 _u10_U3515  ( .A1(1'b0), .A2(_u10_n11999 ), .ZN(_u10_n14992 ) );
NAND2_X1 _u10_U3514  ( .A1(1'b0), .A2(_u10_n11975 ), .ZN(_u10_n14993 ) );
NAND2_X1 _u10_U3513  ( .A1(1'b0), .A2(_u10_n11933 ), .ZN(_u10_n14994 ) );
NAND2_X1 _u10_U3512  ( .A1(1'b0), .A2(_u10_n11909 ), .ZN(_u10_n14995 ) );
NAND4_X1 _u10_U3511  ( .A1(_u10_n14992 ), .A2(_u10_n14993 ), .A3(_u10_n14994 ), .A4(_u10_n14995 ), .ZN(_u10_n14976 ) );
NAND2_X1 _u10_U3510  ( .A1(1'b0), .A2(_u10_n11903 ), .ZN(_u10_n14988 ) );
NAND2_X1 _u10_U3509  ( .A1(1'b0), .A2(_u10_n11879 ), .ZN(_u10_n14989 ) );
NAND2_X1 _u10_U3508  ( .A1(1'b0), .A2(_u10_n11854 ), .ZN(_u10_n14990 ) );
NAND2_X1 _u10_U3507  ( .A1(1'b0), .A2(_u10_n11831 ), .ZN(_u10_n14991 ) );
NAND4_X1 _u10_U3506  ( .A1(_u10_n14988 ), .A2(_u10_n14989 ), .A3(_u10_n14990 ), .A4(_u10_n14991 ), .ZN(_u10_n14977 ) );
NAND2_X1 _u10_U3505  ( .A1(1'b0), .A2(_u10_n11807 ), .ZN(_u10_n14984 ) );
NAND2_X1 _u10_U3504  ( .A1(1'b0), .A2(_u10_n11765 ), .ZN(_u10_n14985 ) );
NAND2_X1 _u10_U3503  ( .A1(1'b0), .A2(_u10_n11738 ), .ZN(_u10_n14986 ) );
NAND2_X1 _u10_U3502  ( .A1(1'b0), .A2(_u10_n11714 ), .ZN(_u10_n14987 ) );
NAND4_X1 _u10_U3501  ( .A1(_u10_n14984 ), .A2(_u10_n14985 ), .A3(_u10_n14986 ), .A4(_u10_n14987 ), .ZN(_u10_n14978 ) );
NAND2_X1 _u10_U3500  ( .A1(1'b0), .A2(_u10_n11690 ), .ZN(_u10_n14980 ) );
NAND2_X1 _u10_U3499  ( .A1(1'b0), .A2(_u10_n11666 ), .ZN(_u10_n14981 ) );
NAND2_X1 _u10_U3498  ( .A1(1'b0), .A2(_u10_n11662 ), .ZN(_u10_n14982 ) );
NAND2_X1 _u10_U3497  ( .A1(1'b0), .A2(_u10_n11638 ), .ZN(_u10_n14983 ) );
NAND4_X1 _u10_U3496  ( .A1(_u10_n14980 ), .A2(_u10_n14981 ), .A3(_u10_n14982 ), .A4(_u10_n14983 ), .ZN(_u10_n14979 ) );
NOR4_X1 _u10_U3495  ( .A1(_u10_n14976 ), .A2(_u10_n14977 ), .A3(_u10_n14978 ), .A4(_u10_n14979 ), .ZN(_u10_n14975 ) );
NAND2_X1 _u10_U3494  ( .A1(_u10_n14974 ), .A2(_u10_n14975 ), .ZN(pointer_s[0]) );
NAND2_X1 _u10_U3493  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n14970 ) );
NAND2_X1 _u10_U3492  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n14971 ) );
NAND2_X1 _u10_U3491  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n14972 ) );
NAND2_X1 _u10_U3490  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n14973 ) );
NAND4_X1 _u10_U3489  ( .A1(_u10_n14970 ), .A2(_u10_n14971 ), .A3(_u10_n14972 ), .A4(_u10_n14973 ), .ZN(_u10_n14955 ) );
NAND2_X1 _u10_U3488  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n14966 ) );
NAND2_X1 _u10_U3487  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n14967 ) );
NAND2_X1 _u10_U3486  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n14968 ) );
NAND2_X1 _u10_U3485  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n14969 ) );
NAND4_X1 _u10_U3484  ( .A1(_u10_n14966 ), .A2(_u10_n14967 ), .A3(_u10_n14968 ), .A4(_u10_n14969 ), .ZN(_u10_n14956 ) );
NAND2_X1 _u10_U3483  ( .A1(1'b0), .A2(_u10_n12164 ), .ZN(_u10_n14962 ) );
NAND2_X1 _u10_U3482  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n14963 ) );
NAND2_X1 _u10_U3481  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n14964 ) );
NAND2_X1 _u10_U3480  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n14965 ) );
NAND4_X1 _u10_U3479  ( .A1(_u10_n14962 ), .A2(_u10_n14963 ), .A3(_u10_n14964 ), .A4(_u10_n14965 ), .ZN(_u10_n14957 ) );
NAND2_X1 _u10_U3478  ( .A1(1'b0), .A2(_u10_n12063 ), .ZN(_u10_n14959 ) );
NAND2_X1 _u10_U3477  ( .A1(1'b0), .A2(_u10_n12039 ), .ZN(_u10_n14960 ) );
NAND2_X1 _u10_U3476  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14961 ) );
NAND3_X1 _u10_U3475  ( .A1(_u10_n14959 ), .A2(_u10_n14960 ), .A3(_u10_n14961 ), .ZN(_u10_n14958 ) );
NOR4_X1 _u10_U3474  ( .A1(_u10_n14955 ), .A2(_u10_n14956 ), .A3(_u10_n14957 ), .A4(_u10_n14958 ), .ZN(_u10_n14933 ) );
NAND2_X1 _u10_U3473  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14951 ) );
NAND2_X1 _u10_U3472  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14952 ) );
NAND2_X1 _u10_U3471  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14953 ) );
NAND2_X1 _u10_U3470  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14954 ) );
NAND4_X1 _u10_U3469  ( .A1(_u10_n14951 ), .A2(_u10_n14952 ), .A3(_u10_n14953 ), .A4(_u10_n14954 ), .ZN(_u10_n14935 ) );
NAND2_X1 _u10_U3468  ( .A1(1'b0), .A2(_u10_n11899 ), .ZN(_u10_n14947 ) );
NAND2_X1 _u10_U3467  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14948 ) );
NAND2_X1 _u10_U3466  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14949 ) );
NAND2_X1 _u10_U3465  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14950 ) );
NAND4_X1 _u10_U3464  ( .A1(_u10_n14947 ), .A2(_u10_n14948 ), .A3(_u10_n14949 ), .A4(_u10_n14950 ), .ZN(_u10_n14936 ) );
NAND2_X1 _u10_U3463  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14943 ) );
NAND2_X1 _u10_U3462  ( .A1(1'b0), .A2(_u10_n11778 ), .ZN(_u10_n14944 ) );
NAND2_X1 _u10_U3461  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14945 ) );
NAND2_X1 _u10_U3460  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14946 ) );
NAND4_X1 _u10_U3459  ( .A1(_u10_n14943 ), .A2(_u10_n14944 ), .A3(_u10_n14945 ), .A4(_u10_n14946 ), .ZN(_u10_n14937 ) );
NAND2_X1 _u10_U3458  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14939 ) );
NAND2_X1 _u10_U3457  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14940 ) );
NAND2_X1 _u10_U3456  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14941 ) );
NAND2_X1 _u10_U3455  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14942 ) );
NAND4_X1 _u10_U3454  ( .A1(_u10_n14939 ), .A2(_u10_n14940 ), .A3(_u10_n14941 ), .A4(_u10_n14942 ), .ZN(_u10_n14938 ) );
NOR4_X1 _u10_U3453  ( .A1(_u10_n14935 ), .A2(_u10_n14936 ), .A3(_u10_n14937 ), .A4(_u10_n14938 ), .ZN(_u10_n14934 ) );
NAND2_X1 _u10_U3452  ( .A1(_u10_n14933 ), .A2(_u10_n14934 ), .ZN(pointer_s[10]) );
NAND2_X1 _u10_U3451  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n14929 ) );
NAND2_X1 _u10_U3450  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n14930 ) );
NAND2_X1 _u10_U3449  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n14931 ) );
NAND2_X1 _u10_U3448  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n14932 ) );
NAND4_X1 _u10_U3447  ( .A1(_u10_n14929 ), .A2(_u10_n14930 ), .A3(_u10_n14931 ), .A4(_u10_n14932 ), .ZN(_u10_n14914 ) );
NAND2_X1 _u10_U3446  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n14925 ) );
NAND2_X1 _u10_U3445  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n14926 ) );
NAND2_X1 _u10_U3444  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n14927 ) );
NAND2_X1 _u10_U3443  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n14928 ) );
NAND4_X1 _u10_U3442  ( .A1(_u10_n14925 ), .A2(_u10_n14926 ), .A3(_u10_n14927 ), .A4(_u10_n14928 ), .ZN(_u10_n14915 ) );
NAND2_X1 _u10_U3441  ( .A1(1'b0), .A2(_u10_n12161 ), .ZN(_u10_n14921 ) );
NAND2_X1 _u10_U3440  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n14922 ) );
NAND2_X1 _u10_U3439  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n14923 ) );
NAND2_X1 _u10_U3438  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n14924 ) );
NAND4_X1 _u10_U3437  ( .A1(_u10_n14921 ), .A2(_u10_n14922 ), .A3(_u10_n14923 ), .A4(_u10_n14924 ), .ZN(_u10_n14916 ) );
NAND2_X1 _u10_U3436  ( .A1(1'b0), .A2(_u10_n12065 ), .ZN(_u10_n14918 ) );
NAND2_X1 _u10_U3435  ( .A1(1'b0), .A2(_u10_n12041 ), .ZN(_u10_n14919 ) );
NAND2_X1 _u10_U3434  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14920 ) );
NAND3_X1 _u10_U3433  ( .A1(_u10_n14918 ), .A2(_u10_n14919 ), .A3(_u10_n14920 ), .ZN(_u10_n14917 ) );
NOR4_X1 _u10_U3432  ( .A1(_u10_n14914 ), .A2(_u10_n14915 ), .A3(_u10_n14916 ), .A4(_u10_n14917 ), .ZN(_u10_n14892 ) );
NAND2_X1 _u10_U3431  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14910 ) );
NAND2_X1 _u10_U3430  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14911 ) );
NAND2_X1 _u10_U3429  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14912 ) );
NAND2_X1 _u10_U3428  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14913 ) );
NAND4_X1 _u10_U3427  ( .A1(_u10_n14910 ), .A2(_u10_n14911 ), .A3(_u10_n14912 ), .A4(_u10_n14913 ), .ZN(_u10_n14894 ) );
NAND2_X1 _u10_U3426  ( .A1(1'b0), .A2(_u10_n11898 ), .ZN(_u10_n14906 ) );
NAND2_X1 _u10_U3425  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14907 ) );
NAND2_X1 _u10_U3424  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14908 ) );
NAND2_X1 _u10_U3423  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14909 ) );
NAND4_X1 _u10_U3422  ( .A1(_u10_n14906 ), .A2(_u10_n14907 ), .A3(_u10_n14908 ), .A4(_u10_n14909 ), .ZN(_u10_n14895 ) );
NAND2_X1 _u10_U3421  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14902 ) );
NAND2_X1 _u10_U3420  ( .A1(1'b0), .A2(_u10_n11779 ), .ZN(_u10_n14903 ) );
NAND2_X1 _u10_U3419  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14904 ) );
NAND2_X1 _u10_U3418  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14905 ) );
NAND4_X1 _u10_U3417  ( .A1(_u10_n14902 ), .A2(_u10_n14903 ), .A3(_u10_n14904 ), .A4(_u10_n14905 ), .ZN(_u10_n14896 ) );
NAND2_X1 _u10_U3416  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14898 ) );
NAND2_X1 _u10_U3415  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14899 ) );
NAND2_X1 _u10_U3414  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14900 ) );
NAND2_X1 _u10_U3413  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14901 ) );
NAND4_X1 _u10_U3412  ( .A1(_u10_n14898 ), .A2(_u10_n14899 ), .A3(_u10_n14900 ), .A4(_u10_n14901 ), .ZN(_u10_n14897 ) );
NOR4_X1 _u10_U3411  ( .A1(_u10_n14894 ), .A2(_u10_n14895 ), .A3(_u10_n14896 ), .A4(_u10_n14897 ), .ZN(_u10_n14893 ) );
NAND2_X1 _u10_U3410  ( .A1(_u10_n14892 ), .A2(_u10_n14893 ), .ZN(pointer_s[11]) );
NAND2_X1 _u10_U3409  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n14888 ) );
NAND2_X1 _u10_U3408  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n14889 ) );
NAND2_X1 _u10_U3407  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n14890 ) );
NAND2_X1 _u10_U3406  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n14891 ) );
NAND4_X1 _u10_U3405  ( .A1(_u10_n14888 ), .A2(_u10_n14889 ), .A3(_u10_n14890 ), .A4(_u10_n14891 ), .ZN(_u10_n14873 ) );
NAND2_X1 _u10_U3404  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n14884 ) );
NAND2_X1 _u10_U3403  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n14885 ) );
NAND2_X1 _u10_U3402  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n14886 ) );
NAND2_X1 _u10_U3401  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n14887 ) );
NAND4_X1 _u10_U3400  ( .A1(_u10_n14884 ), .A2(_u10_n14885 ), .A3(_u10_n14886 ), .A4(_u10_n14887 ), .ZN(_u10_n14874 ) );
NAND2_X1 _u10_U3399  ( .A1(1'b0), .A2(_u10_n12163 ), .ZN(_u10_n14880 ) );
NAND2_X1 _u10_U3398  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n14881 ) );
NAND2_X1 _u10_U3397  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n14882 ) );
NAND2_X1 _u10_U3396  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n14883 ) );
NAND4_X1 _u10_U3395  ( .A1(_u10_n14880 ), .A2(_u10_n14881 ), .A3(_u10_n14882 ), .A4(_u10_n14883 ), .ZN(_u10_n14875 ) );
NAND2_X1 _u10_U3394  ( .A1(1'b0), .A2(_u10_n12406 ), .ZN(_u10_n14877 ) );
NAND2_X1 _u10_U3393  ( .A1(1'b0), .A2(_u10_n12405 ), .ZN(_u10_n14878 ) );
NAND2_X1 _u10_U3392  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14879 ) );
NAND3_X1 _u10_U3391  ( .A1(_u10_n14877 ), .A2(_u10_n14878 ), .A3(_u10_n14879 ), .ZN(_u10_n14876 ) );
NOR4_X1 _u10_U3390  ( .A1(_u10_n14873 ), .A2(_u10_n14874 ), .A3(_u10_n14875 ), .A4(_u10_n14876 ), .ZN(_u10_n14851 ) );
NAND2_X1 _u10_U3389  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14869 ) );
NAND2_X1 _u10_U3388  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14870 ) );
NAND2_X1 _u10_U3387  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14871 ) );
NAND2_X1 _u10_U3386  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14872 ) );
NAND4_X1 _u10_U3385  ( .A1(_u10_n14869 ), .A2(_u10_n14870 ), .A3(_u10_n14871 ), .A4(_u10_n14872 ), .ZN(_u10_n14853 ) );
NAND2_X1 _u10_U3384  ( .A1(1'b0), .A2(_u10_n11903 ), .ZN(_u10_n14865 ) );
NAND2_X1 _u10_U3383  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14866 ) );
NAND2_X1 _u10_U3382  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14867 ) );
NAND2_X1 _u10_U3381  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14868 ) );
NAND4_X1 _u10_U3380  ( .A1(_u10_n14865 ), .A2(_u10_n14866 ), .A3(_u10_n14867 ), .A4(_u10_n14868 ), .ZN(_u10_n14854 ) );
NAND2_X1 _u10_U3379  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14861 ) );
NAND2_X1 _u10_U3378  ( .A1(1'b0), .A2(_u10_n11783 ), .ZN(_u10_n14862 ) );
NAND2_X1 _u10_U3377  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14863 ) );
NAND2_X1 _u10_U3376  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14864 ) );
NAND4_X1 _u10_U3375  ( .A1(_u10_n14861 ), .A2(_u10_n14862 ), .A3(_u10_n14863 ), .A4(_u10_n14864 ), .ZN(_u10_n14855 ) );
NAND2_X1 _u10_U3374  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14857 ) );
NAND2_X1 _u10_U3373  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14858 ) );
NAND2_X1 _u10_U3372  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14859 ) );
NAND2_X1 _u10_U3371  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14860 ) );
NAND4_X1 _u10_U3370  ( .A1(_u10_n14857 ), .A2(_u10_n14858 ), .A3(_u10_n14859 ), .A4(_u10_n14860 ), .ZN(_u10_n14856 ) );
NOR4_X1 _u10_U3369  ( .A1(_u10_n14853 ), .A2(_u10_n14854 ), .A3(_u10_n14855 ), .A4(_u10_n14856 ), .ZN(_u10_n14852 ) );
NAND2_X1 _u10_U3368  ( .A1(_u10_n14851 ), .A2(_u10_n14852 ), .ZN(pointer_s[12]) );
NAND2_X1 _u10_U3367  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n14847 ) );
NAND2_X1 _u10_U3366  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n14848 ) );
NAND2_X1 _u10_U3365  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n14849 ) );
NAND2_X1 _u10_U3364  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n14850 ) );
NAND4_X1 _u10_U3363  ( .A1(_u10_n14847 ), .A2(_u10_n14848 ), .A3(_u10_n14849 ), .A4(_u10_n14850 ), .ZN(_u10_n14832 ) );
NAND2_X1 _u10_U3362  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n14843 ) );
NAND2_X1 _u10_U3361  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n14844 ) );
NAND2_X1 _u10_U3360  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n14845 ) );
NAND2_X1 _u10_U3359  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n14846 ) );
NAND4_X1 _u10_U3358  ( .A1(_u10_n14843 ), .A2(_u10_n14844 ), .A3(_u10_n14845 ), .A4(_u10_n14846 ), .ZN(_u10_n14833 ) );
NAND2_X1 _u10_U3357  ( .A1(1'b0), .A2(_u10_n12414 ), .ZN(_u10_n14839 ) );
NAND2_X1 _u10_U3356  ( .A1(1'b0), .A2(_u10_n12130 ), .ZN(_u10_n14840 ) );
NAND2_X1 _u10_U3355  ( .A1(1'b0), .A2(_u10_n12106 ), .ZN(_u10_n14841 ) );
NAND2_X1 _u10_U3354  ( .A1(1'b0), .A2(_u10_n12082 ), .ZN(_u10_n14842 ) );
NAND4_X1 _u10_U3353  ( .A1(_u10_n14839 ), .A2(_u10_n14840 ), .A3(_u10_n14841 ), .A4(_u10_n14842 ), .ZN(_u10_n14834 ) );
NAND2_X1 _u10_U3352  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n14836 ) );
NAND2_X1 _u10_U3351  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n14837 ) );
NAND2_X1 _u10_U3350  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14838 ) );
NAND3_X1 _u10_U3349  ( .A1(_u10_n14836 ), .A2(_u10_n14837 ), .A3(_u10_n14838 ), .ZN(_u10_n14835 ) );
NOR4_X1 _u10_U3348  ( .A1(_u10_n14832 ), .A2(_u10_n14833 ), .A3(_u10_n14834 ), .A4(_u10_n14835 ), .ZN(_u10_n14810 ) );
NAND2_X1 _u10_U3347  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14828 ) );
NAND2_X1 _u10_U3346  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14829 ) );
NAND2_X1 _u10_U3345  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14830 ) );
NAND2_X1 _u10_U3344  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14831 ) );
NAND4_X1 _u10_U3343  ( .A1(_u10_n14828 ), .A2(_u10_n14829 ), .A3(_u10_n14830 ), .A4(_u10_n14831 ), .ZN(_u10_n14812 ) );
NAND2_X1 _u10_U3342  ( .A1(1'b0), .A2(_u10_n12388 ), .ZN(_u10_n14824 ) );
NAND2_X1 _u10_U3341  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14825 ) );
NAND2_X1 _u10_U3340  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14826 ) );
NAND2_X1 _u10_U3339  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14827 ) );
NAND4_X1 _u10_U3338  ( .A1(_u10_n14824 ), .A2(_u10_n14825 ), .A3(_u10_n14826 ), .A4(_u10_n14827 ), .ZN(_u10_n14813 ) );
NAND2_X1 _u10_U3337  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14820 ) );
NAND2_X1 _u10_U3336  ( .A1(1'b0), .A2(_u10_n12379 ), .ZN(_u10_n14821 ) );
NAND2_X1 _u10_U3335  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14822 ) );
NAND2_X1 _u10_U3334  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14823 ) );
NAND4_X1 _u10_U3333  ( .A1(_u10_n14820 ), .A2(_u10_n14821 ), .A3(_u10_n14822 ), .A4(_u10_n14823 ), .ZN(_u10_n14814 ) );
NAND2_X1 _u10_U3332  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14816 ) );
NAND2_X1 _u10_U3331  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14817 ) );
NAND2_X1 _u10_U3330  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14818 ) );
NAND2_X1 _u10_U3329  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14819 ) );
NAND4_X1 _u10_U3328  ( .A1(_u10_n14816 ), .A2(_u10_n14817 ), .A3(_u10_n14818 ), .A4(_u10_n14819 ), .ZN(_u10_n14815 ) );
NOR4_X1 _u10_U3327  ( .A1(_u10_n14812 ), .A2(_u10_n14813 ), .A3(_u10_n14814 ), .A4(_u10_n14815 ), .ZN(_u10_n14811 ) );
NAND2_X1 _u10_U3326  ( .A1(_u10_n14810 ), .A2(_u10_n14811 ), .ZN(pointer_s[13]) );
NAND2_X1 _u10_U3325  ( .A1(1'b0), .A2(_u10_n12346 ), .ZN(_u10_n14806 ) );
NAND2_X1 _u10_U3324  ( .A1(1'b0), .A2(_u10_n12322 ), .ZN(_u10_n14807 ) );
NAND2_X1 _u10_U3323  ( .A1(1'b0), .A2(_u10_n12299 ), .ZN(_u10_n14808 ) );
NAND2_X1 _u10_U3322  ( .A1(1'b0), .A2(_u10_n12275 ), .ZN(_u10_n14809 ) );
NAND4_X1 _u10_U3321  ( .A1(_u10_n14806 ), .A2(_u10_n14807 ), .A3(_u10_n14808 ), .A4(_u10_n14809 ), .ZN(_u10_n14791 ) );
NAND2_X1 _u10_U3320  ( .A1(1'b0), .A2(_u10_n12250 ), .ZN(_u10_n14802 ) );
NAND2_X1 _u10_U3319  ( .A1(1'b0), .A2(_u10_n12226 ), .ZN(_u10_n14803 ) );
NAND2_X1 _u10_U3318  ( .A1(1'b0), .A2(_u10_n12200 ), .ZN(_u10_n14804 ) );
NAND2_X1 _u10_U3317  ( .A1(1'b0), .A2(_u10_n12178 ), .ZN(_u10_n14805 ) );
NAND4_X1 _u10_U3316  ( .A1(_u10_n14802 ), .A2(_u10_n14803 ), .A3(_u10_n14804 ), .A4(_u10_n14805 ), .ZN(_u10_n14792 ) );
NAND2_X1 _u10_U3315  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14798 ) );
NAND2_X1 _u10_U3314  ( .A1(1'b0), .A2(_u10_n12135 ), .ZN(_u10_n14799 ) );
NAND2_X1 _u10_U3313  ( .A1(1'b0), .A2(_u10_n12111 ), .ZN(_u10_n14800 ) );
NAND2_X1 _u10_U3312  ( .A1(1'b0), .A2(_u10_n12087 ), .ZN(_u10_n14801 ) );
NAND4_X1 _u10_U3311  ( .A1(_u10_n14798 ), .A2(_u10_n14799 ), .A3(_u10_n14800 ), .A4(_u10_n14801 ), .ZN(_u10_n14793 ) );
NAND2_X1 _u10_U3310  ( .A1(1'b0), .A2(_u10_n12064 ), .ZN(_u10_n14795 ) );
NAND2_X1 _u10_U3309  ( .A1(1'b0), .A2(_u10_n12040 ), .ZN(_u10_n14796 ) );
NAND2_X1 _u10_U3308  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14797 ) );
NAND3_X1 _u10_U3307  ( .A1(_u10_n14795 ), .A2(_u10_n14796 ), .A3(_u10_n14797 ), .ZN(_u10_n14794 ) );
NOR4_X1 _u10_U3306  ( .A1(_u10_n14791 ), .A2(_u10_n14792 ), .A3(_u10_n14793 ), .A4(_u10_n14794 ), .ZN(_u10_n14769 ) );
NAND2_X1 _u10_U3305  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14787 ) );
NAND2_X1 _u10_U3304  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14788 ) );
NAND2_X1 _u10_U3303  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14789 ) );
NAND2_X1 _u10_U3302  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14790 ) );
NAND4_X1 _u10_U3301  ( .A1(_u10_n14787 ), .A2(_u10_n14788 ), .A3(_u10_n14789 ), .A4(_u10_n14790 ), .ZN(_u10_n14771 ) );
NAND2_X1 _u10_U3300  ( .A1(1'b0), .A2(_u10_n11897 ), .ZN(_u10_n14783 ) );
NAND2_X1 _u10_U3299  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14784 ) );
NAND2_X1 _u10_U3298  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14785 ) );
NAND2_X1 _u10_U3297  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14786 ) );
NAND4_X1 _u10_U3296  ( .A1(_u10_n14783 ), .A2(_u10_n14784 ), .A3(_u10_n14785 ), .A4(_u10_n14786 ), .ZN(_u10_n14772 ) );
NAND2_X1 _u10_U3295  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14779 ) );
NAND2_X1 _u10_U3294  ( .A1(1'b0), .A2(_u10_n11777 ), .ZN(_u10_n14780 ) );
NAND2_X1 _u10_U3293  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14781 ) );
NAND2_X1 _u10_U3292  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14782 ) );
NAND4_X1 _u10_U3291  ( .A1(_u10_n14779 ), .A2(_u10_n14780 ), .A3(_u10_n14781 ), .A4(_u10_n14782 ), .ZN(_u10_n14773 ) );
NAND2_X1 _u10_U3290  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14775 ) );
NAND2_X1 _u10_U3289  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14776 ) );
NAND2_X1 _u10_U3288  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14777 ) );
NAND2_X1 _u10_U3287  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14778 ) );
NAND4_X1 _u10_U3286  ( .A1(_u10_n14775 ), .A2(_u10_n14776 ), .A3(_u10_n14777 ), .A4(_u10_n14778 ), .ZN(_u10_n14774 ) );
NOR4_X1 _u10_U3285  ( .A1(_u10_n14771 ), .A2(_u10_n14772 ), .A3(_u10_n14773 ), .A4(_u10_n14774 ), .ZN(_u10_n14770 ) );
NAND2_X1 _u10_U3284  ( .A1(_u10_n14769 ), .A2(_u10_n14770 ), .ZN(pointer_s[14]) );
NAND2_X1 _u10_U3283  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14765 ) );
NAND2_X1 _u10_U3282  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14766 ) );
NAND2_X1 _u10_U3281  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14767 ) );
NAND2_X1 _u10_U3280  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14768 ) );
NAND4_X1 _u10_U3279  ( .A1(_u10_n14765 ), .A2(_u10_n14766 ), .A3(_u10_n14767 ), .A4(_u10_n14768 ), .ZN(_u10_n14750 ) );
NAND2_X1 _u10_U3278  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14761 ) );
NAND2_X1 _u10_U3277  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14762 ) );
NAND2_X1 _u10_U3276  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14763 ) );
NAND2_X1 _u10_U3275  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14764 ) );
NAND4_X1 _u10_U3274  ( .A1(_u10_n14761 ), .A2(_u10_n14762 ), .A3(_u10_n14763 ), .A4(_u10_n14764 ), .ZN(_u10_n14751 ) );
NAND2_X1 _u10_U3273  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14757 ) );
NAND2_X1 _u10_U3272  ( .A1(1'b0), .A2(_u10_n12136 ), .ZN(_u10_n14758 ) );
NAND2_X1 _u10_U3271  ( .A1(1'b0), .A2(_u10_n12112 ), .ZN(_u10_n14759 ) );
NAND2_X1 _u10_U3270  ( .A1(1'b0), .A2(_u10_n12088 ), .ZN(_u10_n14760 ) );
NAND4_X1 _u10_U3269  ( .A1(_u10_n14757 ), .A2(_u10_n14758 ), .A3(_u10_n14759 ), .A4(_u10_n14760 ), .ZN(_u10_n14752 ) );
NAND2_X1 _u10_U3268  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14754 ) );
NAND2_X1 _u10_U3267  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14755 ) );
NAND2_X1 _u10_U3266  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14756 ) );
NAND3_X1 _u10_U3265  ( .A1(_u10_n14754 ), .A2(_u10_n14755 ), .A3(_u10_n14756 ), .ZN(_u10_n14753 ) );
NOR4_X1 _u10_U3264  ( .A1(_u10_n14750 ), .A2(_u10_n14751 ), .A3(_u10_n14752 ), .A4(_u10_n14753 ), .ZN(_u10_n14728 ) );
NAND2_X1 _u10_U3263  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14746 ) );
NAND2_X1 _u10_U3262  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14747 ) );
NAND2_X1 _u10_U3261  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14748 ) );
NAND2_X1 _u10_U3260  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14749 ) );
NAND4_X1 _u10_U3259  ( .A1(_u10_n14746 ), .A2(_u10_n14747 ), .A3(_u10_n14748 ), .A4(_u10_n14749 ), .ZN(_u10_n14730 ) );
NAND2_X1 _u10_U3258  ( .A1(1'b0), .A2(_u10_n12388 ), .ZN(_u10_n14742 ) );
NAND2_X1 _u10_U3257  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14743 ) );
NAND2_X1 _u10_U3256  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14744 ) );
NAND2_X1 _u10_U3255  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14745 ) );
NAND4_X1 _u10_U3254  ( .A1(_u10_n14742 ), .A2(_u10_n14743 ), .A3(_u10_n14744 ), .A4(_u10_n14745 ), .ZN(_u10_n14731 ) );
NAND2_X1 _u10_U3253  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14738 ) );
NAND2_X1 _u10_U3252  ( .A1(1'b0), .A2(_u10_n11782 ), .ZN(_u10_n14739 ) );
NAND2_X1 _u10_U3251  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14740 ) );
NAND2_X1 _u10_U3250  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14741 ) );
NAND4_X1 _u10_U3249  ( .A1(_u10_n14738 ), .A2(_u10_n14739 ), .A3(_u10_n14740 ), .A4(_u10_n14741 ), .ZN(_u10_n14732 ) );
NAND2_X1 _u10_U3248  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14734 ) );
NAND2_X1 _u10_U3247  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14735 ) );
NAND2_X1 _u10_U3246  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14736 ) );
NAND2_X1 _u10_U3245  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14737 ) );
NAND4_X1 _u10_U3244  ( .A1(_u10_n14734 ), .A2(_u10_n14735 ), .A3(_u10_n14736 ), .A4(_u10_n14737 ), .ZN(_u10_n14733 ) );
NOR4_X1 _u10_U3243  ( .A1(_u10_n14730 ), .A2(_u10_n14731 ), .A3(_u10_n14732 ), .A4(_u10_n14733 ), .ZN(_u10_n14729 ) );
NAND2_X1 _u10_U3242  ( .A1(_u10_n14728 ), .A2(_u10_n14729 ), .ZN(pointer_s[15]) );
NAND2_X1 _u10_U3241  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14724 ) );
NAND2_X1 _u10_U3240  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14725 ) );
NAND2_X1 _u10_U3239  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14726 ) );
NAND2_X1 _u10_U3238  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14727 ) );
NAND4_X1 _u10_U3237  ( .A1(_u10_n14724 ), .A2(_u10_n14725 ), .A3(_u10_n14726 ), .A4(_u10_n14727 ), .ZN(_u10_n14709 ) );
NAND2_X1 _u10_U3236  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14720 ) );
NAND2_X1 _u10_U3235  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14721 ) );
NAND2_X1 _u10_U3234  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14722 ) );
NAND2_X1 _u10_U3233  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14723 ) );
NAND4_X1 _u10_U3232  ( .A1(_u10_n14720 ), .A2(_u10_n14721 ), .A3(_u10_n14722 ), .A4(_u10_n14723 ), .ZN(_u10_n14710 ) );
NAND2_X1 _u10_U3231  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14716 ) );
NAND2_X1 _u10_U3230  ( .A1(1'b0), .A2(_u10_n12413 ), .ZN(_u10_n14717 ) );
NAND2_X1 _u10_U3229  ( .A1(1'b0), .A2(_u10_n12412 ), .ZN(_u10_n14718 ) );
NAND2_X1 _u10_U3228  ( .A1(1'b0), .A2(_u10_n12411 ), .ZN(_u10_n14719 ) );
NAND4_X1 _u10_U3227  ( .A1(_u10_n14716 ), .A2(_u10_n14717 ), .A3(_u10_n14718 ), .A4(_u10_n14719 ), .ZN(_u10_n14711 ) );
NAND2_X1 _u10_U3226  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14713 ) );
NAND2_X1 _u10_U3225  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14714 ) );
NAND2_X1 _u10_U3224  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14715 ) );
NAND3_X1 _u10_U3223  ( .A1(_u10_n14713 ), .A2(_u10_n14714 ), .A3(_u10_n14715 ), .ZN(_u10_n14712 ) );
NOR4_X1 _u10_U3222  ( .A1(_u10_n14709 ), .A2(_u10_n14710 ), .A3(_u10_n14711 ), .A4(_u10_n14712 ), .ZN(_u10_n14687 ) );
NAND2_X1 _u10_U3221  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14705 ) );
NAND2_X1 _u10_U3220  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14706 ) );
NAND2_X1 _u10_U3219  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14707 ) );
NAND2_X1 _u10_U3218  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14708 ) );
NAND4_X1 _u10_U3217  ( .A1(_u10_n14705 ), .A2(_u10_n14706 ), .A3(_u10_n14707 ), .A4(_u10_n14708 ), .ZN(_u10_n14689 ) );
NAND2_X1 _u10_U3216  ( .A1(1'b0), .A2(_u10_n11900 ), .ZN(_u10_n14701 ) );
NAND2_X1 _u10_U3215  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14702 ) );
NAND2_X1 _u10_U3214  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14703 ) );
NAND2_X1 _u10_U3213  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14704 ) );
NAND4_X1 _u10_U3212  ( .A1(_u10_n14701 ), .A2(_u10_n14702 ), .A3(_u10_n14703 ), .A4(_u10_n14704 ), .ZN(_u10_n14690 ) );
NAND2_X1 _u10_U3211  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14697 ) );
NAND2_X1 _u10_U3210  ( .A1(1'b0), .A2(_u10_n11780 ), .ZN(_u10_n14698 ) );
NAND2_X1 _u10_U3209  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14699 ) );
NAND2_X1 _u10_U3208  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14700 ) );
NAND4_X1 _u10_U3207  ( .A1(_u10_n14697 ), .A2(_u10_n14698 ), .A3(_u10_n14699 ), .A4(_u10_n14700 ), .ZN(_u10_n14691 ) );
NAND2_X1 _u10_U3206  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14693 ) );
NAND2_X1 _u10_U3205  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14694 ) );
NAND2_X1 _u10_U3204  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14695 ) );
NAND2_X1 _u10_U3203  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14696 ) );
NAND4_X1 _u10_U3202  ( .A1(_u10_n14693 ), .A2(_u10_n14694 ), .A3(_u10_n14695 ), .A4(_u10_n14696 ), .ZN(_u10_n14692 ) );
NOR4_X1 _u10_U3201  ( .A1(_u10_n14689 ), .A2(_u10_n14690 ), .A3(_u10_n14691 ), .A4(_u10_n14692 ), .ZN(_u10_n14688 ) );
NAND2_X1 _u10_U3200  ( .A1(_u10_n14687 ), .A2(_u10_n14688 ), .ZN(pointer_s[16]) );
NAND2_X1 _u10_U3199  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14683 ) );
NAND2_X1 _u10_U3198  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14684 ) );
NAND2_X1 _u10_U3197  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14685 ) );
NAND2_X1 _u10_U3196  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14686 ) );
NAND4_X1 _u10_U3195  ( .A1(_u10_n14683 ), .A2(_u10_n14684 ), .A3(_u10_n14685 ), .A4(_u10_n14686 ), .ZN(_u10_n14668 ) );
NAND2_X1 _u10_U3194  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14679 ) );
NAND2_X1 _u10_U3193  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14680 ) );
NAND2_X1 _u10_U3192  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14681 ) );
NAND2_X1 _u10_U3191  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14682 ) );
NAND4_X1 _u10_U3190  ( .A1(_u10_n14679 ), .A2(_u10_n14680 ), .A3(_u10_n14681 ), .A4(_u10_n14682 ), .ZN(_u10_n14669 ) );
NAND2_X1 _u10_U3189  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14675 ) );
NAND2_X1 _u10_U3188  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n14676 ) );
NAND2_X1 _u10_U3187  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n14677 ) );
NAND2_X1 _u10_U3186  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n14678 ) );
NAND4_X1 _u10_U3185  ( .A1(_u10_n14675 ), .A2(_u10_n14676 ), .A3(_u10_n14677 ), .A4(_u10_n14678 ), .ZN(_u10_n14670 ) );
NAND2_X1 _u10_U3184  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14672 ) );
NAND2_X1 _u10_U3183  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14673 ) );
NAND2_X1 _u10_U3182  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14674 ) );
NAND3_X1 _u10_U3181  ( .A1(_u10_n14672 ), .A2(_u10_n14673 ), .A3(_u10_n14674 ), .ZN(_u10_n14671 ) );
NOR4_X1 _u10_U3180  ( .A1(_u10_n14668 ), .A2(_u10_n14669 ), .A3(_u10_n14670 ), .A4(_u10_n14671 ), .ZN(_u10_n14646 ) );
NAND2_X1 _u10_U3179  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14664 ) );
NAND2_X1 _u10_U3178  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14665 ) );
NAND2_X1 _u10_U3177  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14666 ) );
NAND2_X1 _u10_U3176  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14667 ) );
NAND4_X1 _u10_U3175  ( .A1(_u10_n14664 ), .A2(_u10_n14665 ), .A3(_u10_n14666 ), .A4(_u10_n14667 ), .ZN(_u10_n14648 ) );
NAND2_X1 _u10_U3174  ( .A1(1'b0), .A2(_u10_n11901 ), .ZN(_u10_n14660 ) );
NAND2_X1 _u10_U3173  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14661 ) );
NAND2_X1 _u10_U3172  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14662 ) );
NAND2_X1 _u10_U3171  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14663 ) );
NAND4_X1 _u10_U3170  ( .A1(_u10_n14660 ), .A2(_u10_n14661 ), .A3(_u10_n14662 ), .A4(_u10_n14663 ), .ZN(_u10_n14649 ) );
NAND2_X1 _u10_U3169  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14656 ) );
NAND2_X1 _u10_U3168  ( .A1(1'b0), .A2(_u10_n11781 ), .ZN(_u10_n14657 ) );
NAND2_X1 _u10_U3167  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14658 ) );
NAND2_X1 _u10_U3166  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14659 ) );
NAND4_X1 _u10_U3165  ( .A1(_u10_n14656 ), .A2(_u10_n14657 ), .A3(_u10_n14658 ), .A4(_u10_n14659 ), .ZN(_u10_n14650 ) );
NAND2_X1 _u10_U3164  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14652 ) );
NAND2_X1 _u10_U3163  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14653 ) );
NAND2_X1 _u10_U3162  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14654 ) );
NAND2_X1 _u10_U3161  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14655 ) );
NAND4_X1 _u10_U3160  ( .A1(_u10_n14652 ), .A2(_u10_n14653 ), .A3(_u10_n14654 ), .A4(_u10_n14655 ), .ZN(_u10_n14651 ) );
NOR4_X1 _u10_U3159  ( .A1(_u10_n14648 ), .A2(_u10_n14649 ), .A3(_u10_n14650 ), .A4(_u10_n14651 ), .ZN(_u10_n14647 ) );
NAND2_X1 _u10_U3158  ( .A1(_u10_n14646 ), .A2(_u10_n14647 ), .ZN(pointer_s[17]) );
NAND2_X1 _u10_U3157  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14642 ) );
NAND2_X1 _u10_U3156  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14643 ) );
NAND2_X1 _u10_U3155  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14644 ) );
NAND2_X1 _u10_U3154  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14645 ) );
NAND4_X1 _u10_U3153  ( .A1(_u10_n14642 ), .A2(_u10_n14643 ), .A3(_u10_n14644 ), .A4(_u10_n14645 ), .ZN(_u10_n14627 ) );
NAND2_X1 _u10_U3152  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14638 ) );
NAND2_X1 _u10_U3151  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14639 ) );
NAND2_X1 _u10_U3150  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14640 ) );
NAND2_X1 _u10_U3149  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14641 ) );
NAND4_X1 _u10_U3148  ( .A1(_u10_n14638 ), .A2(_u10_n14639 ), .A3(_u10_n14640 ), .A4(_u10_n14641 ), .ZN(_u10_n14628 ) );
NAND2_X1 _u10_U3147  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14634 ) );
NAND2_X1 _u10_U3146  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n14635 ) );
NAND2_X1 _u10_U3145  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n14636 ) );
NAND2_X1 _u10_U3144  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n14637 ) );
NAND4_X1 _u10_U3143  ( .A1(_u10_n14634 ), .A2(_u10_n14635 ), .A3(_u10_n14636 ), .A4(_u10_n14637 ), .ZN(_u10_n14629 ) );
NAND2_X1 _u10_U3142  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14631 ) );
NAND2_X1 _u10_U3141  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14632 ) );
NAND2_X1 _u10_U3140  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14633 ) );
NAND3_X1 _u10_U3139  ( .A1(_u10_n14631 ), .A2(_u10_n14632 ), .A3(_u10_n14633 ), .ZN(_u10_n14630 ) );
NOR4_X1 _u10_U3138  ( .A1(_u10_n14627 ), .A2(_u10_n14628 ), .A3(_u10_n14629 ), .A4(_u10_n14630 ), .ZN(_u10_n14605 ) );
NAND2_X1 _u10_U3137  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14623 ) );
NAND2_X1 _u10_U3136  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14624 ) );
NAND2_X1 _u10_U3135  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14625 ) );
NAND2_X1 _u10_U3134  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14626 ) );
NAND4_X1 _u10_U3133  ( .A1(_u10_n14623 ), .A2(_u10_n14624 ), .A3(_u10_n14625 ), .A4(_u10_n14626 ), .ZN(_u10_n14607 ) );
NAND2_X1 _u10_U3132  ( .A1(1'b0), .A2(_u10_n11902 ), .ZN(_u10_n14619 ) );
NAND2_X1 _u10_U3131  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14620 ) );
NAND2_X1 _u10_U3130  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14621 ) );
NAND2_X1 _u10_U3129  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14622 ) );
NAND4_X1 _u10_U3128  ( .A1(_u10_n14619 ), .A2(_u10_n14620 ), .A3(_u10_n14621 ), .A4(_u10_n14622 ), .ZN(_u10_n14608 ) );
NAND2_X1 _u10_U3127  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14615 ) );
NAND2_X1 _u10_U3126  ( .A1(1'b0), .A2(_u10_n11778 ), .ZN(_u10_n14616 ) );
NAND2_X1 _u10_U3125  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14617 ) );
NAND2_X1 _u10_U3124  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14618 ) );
NAND4_X1 _u10_U3123  ( .A1(_u10_n14615 ), .A2(_u10_n14616 ), .A3(_u10_n14617 ), .A4(_u10_n14618 ), .ZN(_u10_n14609 ) );
NAND2_X1 _u10_U3122  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14611 ) );
NAND2_X1 _u10_U3121  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14612 ) );
NAND2_X1 _u10_U3120  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14613 ) );
NAND2_X1 _u10_U3119  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14614 ) );
NAND4_X1 _u10_U3118  ( .A1(_u10_n14611 ), .A2(_u10_n14612 ), .A3(_u10_n14613 ), .A4(_u10_n14614 ), .ZN(_u10_n14610 ) );
NOR4_X1 _u10_U3117  ( .A1(_u10_n14607 ), .A2(_u10_n14608 ), .A3(_u10_n14609 ), .A4(_u10_n14610 ), .ZN(_u10_n14606 ) );
NAND2_X1 _u10_U3116  ( .A1(_u10_n14605 ), .A2(_u10_n14606 ), .ZN(pointer_s[18]) );
NAND2_X1 _u10_U3115  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14601 ) );
NAND2_X1 _u10_U3114  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14602 ) );
NAND2_X1 _u10_U3113  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14603 ) );
NAND2_X1 _u10_U3112  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14604 ) );
NAND4_X1 _u10_U3111  ( .A1(_u10_n14601 ), .A2(_u10_n14602 ), .A3(_u10_n14603 ), .A4(_u10_n14604 ), .ZN(_u10_n14586 ) );
NAND2_X1 _u10_U3110  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14597 ) );
NAND2_X1 _u10_U3109  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14598 ) );
NAND2_X1 _u10_U3108  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14599 ) );
NAND2_X1 _u10_U3107  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14600 ) );
NAND4_X1 _u10_U3106  ( .A1(_u10_n14597 ), .A2(_u10_n14598 ), .A3(_u10_n14599 ), .A4(_u10_n14600 ), .ZN(_u10_n14587 ) );
NAND2_X1 _u10_U3105  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14593 ) );
NAND2_X1 _u10_U3104  ( .A1(1'b0), .A2(_u10_n12135 ), .ZN(_u10_n14594 ) );
NAND2_X1 _u10_U3103  ( .A1(1'b0), .A2(_u10_n12111 ), .ZN(_u10_n14595 ) );
NAND2_X1 _u10_U3102  ( .A1(1'b0), .A2(_u10_n12087 ), .ZN(_u10_n14596 ) );
NAND4_X1 _u10_U3101  ( .A1(_u10_n14593 ), .A2(_u10_n14594 ), .A3(_u10_n14595 ), .A4(_u10_n14596 ), .ZN(_u10_n14588 ) );
NAND2_X1 _u10_U3100  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14590 ) );
NAND2_X1 _u10_U3099  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14591 ) );
NAND2_X1 _u10_U3098  ( .A1(1'b0), .A2(_u10_n12015 ), .ZN(_u10_n14592 ) );
NAND3_X1 _u10_U3097  ( .A1(_u10_n14590 ), .A2(_u10_n14591 ), .A3(_u10_n14592 ), .ZN(_u10_n14589 ) );
NOR4_X1 _u10_U3096  ( .A1(_u10_n14586 ), .A2(_u10_n14587 ), .A3(_u10_n14588 ), .A4(_u10_n14589 ), .ZN(_u10_n14564 ) );
NAND2_X1 _u10_U3095  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14582 ) );
NAND2_X1 _u10_U3094  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14583 ) );
NAND2_X1 _u10_U3093  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14584 ) );
NAND2_X1 _u10_U3092  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14585 ) );
NAND4_X1 _u10_U3091  ( .A1(_u10_n14582 ), .A2(_u10_n14583 ), .A3(_u10_n14584 ), .A4(_u10_n14585 ), .ZN(_u10_n14566 ) );
NAND2_X1 _u10_U3090  ( .A1(1'b0), .A2(_u10_n11899 ), .ZN(_u10_n14578 ) );
NAND2_X1 _u10_U3089  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14579 ) );
NAND2_X1 _u10_U3088  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14580 ) );
NAND2_X1 _u10_U3087  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14581 ) );
NAND4_X1 _u10_U3086  ( .A1(_u10_n14578 ), .A2(_u10_n14579 ), .A3(_u10_n14580 ), .A4(_u10_n14581 ), .ZN(_u10_n14567 ) );
NAND2_X1 _u10_U3085  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14574 ) );
NAND2_X1 _u10_U3084  ( .A1(1'b0), .A2(_u10_n11779 ), .ZN(_u10_n14575 ) );
NAND2_X1 _u10_U3083  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14576 ) );
NAND2_X1 _u10_U3082  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14577 ) );
NAND4_X1 _u10_U3081  ( .A1(_u10_n14574 ), .A2(_u10_n14575 ), .A3(_u10_n14576 ), .A4(_u10_n14577 ), .ZN(_u10_n14568 ) );
NAND2_X1 _u10_U3080  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14570 ) );
NAND2_X1 _u10_U3079  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14571 ) );
NAND2_X1 _u10_U3078  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14572 ) );
NAND2_X1 _u10_U3077  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14573 ) );
NAND4_X1 _u10_U3076  ( .A1(_u10_n14570 ), .A2(_u10_n14571 ), .A3(_u10_n14572 ), .A4(_u10_n14573 ), .ZN(_u10_n14569 ) );
NOR4_X1 _u10_U3075  ( .A1(_u10_n14566 ), .A2(_u10_n14567 ), .A3(_u10_n14568 ), .A4(_u10_n14569 ), .ZN(_u10_n14565 ) );
NAND2_X1 _u10_U3074  ( .A1(_u10_n14564 ), .A2(_u10_n14565 ), .ZN(pointer_s[19]) );
NAND2_X1 _u10_U3073  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14560 ) );
NAND2_X1 _u10_U3072  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14561 ) );
NAND2_X1 _u10_U3071  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14562 ) );
NAND2_X1 _u10_U3070  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14563 ) );
NAND4_X1 _u10_U3069  ( .A1(_u10_n14560 ), .A2(_u10_n14561 ), .A3(_u10_n14562 ), .A4(_u10_n14563 ), .ZN(_u10_n14545 ) );
NAND2_X1 _u10_U3068  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14556 ) );
NAND2_X1 _u10_U3067  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14557 ) );
NAND2_X1 _u10_U3066  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14558 ) );
NAND2_X1 _u10_U3065  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14559 ) );
NAND4_X1 _u10_U3064  ( .A1(_u10_n14556 ), .A2(_u10_n14557 ), .A3(_u10_n14558 ), .A4(_u10_n14559 ), .ZN(_u10_n14546 ) );
NAND2_X1 _u10_U3063  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14552 ) );
NAND2_X1 _u10_U3062  ( .A1(1'b0), .A2(_u10_n12137 ), .ZN(_u10_n14553 ) );
NAND2_X1 _u10_U3061  ( .A1(1'b0), .A2(_u10_n12113 ), .ZN(_u10_n14554 ) );
NAND2_X1 _u10_U3060  ( .A1(1'b0), .A2(_u10_n12089 ), .ZN(_u10_n14555 ) );
NAND4_X1 _u10_U3059  ( .A1(_u10_n14552 ), .A2(_u10_n14553 ), .A3(_u10_n14554 ), .A4(_u10_n14555 ), .ZN(_u10_n14547 ) );
NAND2_X1 _u10_U3058  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14549 ) );
NAND2_X1 _u10_U3057  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14550 ) );
NAND2_X1 _u10_U3056  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14551 ) );
NAND3_X1 _u10_U3055  ( .A1(_u10_n14549 ), .A2(_u10_n14550 ), .A3(_u10_n14551 ), .ZN(_u10_n14548 ) );
NOR4_X1 _u10_U3054  ( .A1(_u10_n14545 ), .A2(_u10_n14546 ), .A3(_u10_n14547 ), .A4(_u10_n14548 ), .ZN(_u10_n14523 ) );
NAND2_X1 _u10_U3053  ( .A1(1'b0), .A2(_u10_n11979 ), .ZN(_u10_n14541 ) );
NAND2_X1 _u10_U3052  ( .A1(1'b0), .A2(_u10_n11955 ), .ZN(_u10_n14542 ) );
NAND2_X1 _u10_U3051  ( .A1(1'b0), .A2(_u10_n11934 ), .ZN(_u10_n14543 ) );
NAND2_X1 _u10_U3050  ( .A1(1'b0), .A2(_u10_n11910 ), .ZN(_u10_n14544 ) );
NAND4_X1 _u10_U3049  ( .A1(_u10_n14541 ), .A2(_u10_n14542 ), .A3(_u10_n14543 ), .A4(_u10_n14544 ), .ZN(_u10_n14525 ) );
NAND2_X1 _u10_U3048  ( .A1(1'b0), .A2(_u10_n11897 ), .ZN(_u10_n14537 ) );
NAND2_X1 _u10_U3047  ( .A1(1'b0), .A2(_u10_n11859 ), .ZN(_u10_n14538 ) );
NAND2_X1 _u10_U3046  ( .A1(1'b0), .A2(_u10_n11835 ), .ZN(_u10_n14539 ) );
NAND2_X1 _u10_U3045  ( .A1(1'b0), .A2(_u10_n11813 ), .ZN(_u10_n14540 ) );
NAND4_X1 _u10_U3044  ( .A1(_u10_n14537 ), .A2(_u10_n14538 ), .A3(_u10_n14539 ), .A4(_u10_n14540 ), .ZN(_u10_n14526 ) );
NAND2_X1 _u10_U3043  ( .A1(1'b0), .A2(_u10_n11787 ), .ZN(_u10_n14533 ) );
NAND2_X1 _u10_U3042  ( .A1(1'b0), .A2(_u10_n11782 ), .ZN(_u10_n14534 ) );
NAND2_X1 _u10_U3041  ( .A1(1'b0), .A2(_u10_n11739 ), .ZN(_u10_n14535 ) );
NAND2_X1 _u10_U3040  ( .A1(1'b0), .A2(_u10_n11715 ), .ZN(_u10_n14536 ) );
NAND4_X1 _u10_U3039  ( .A1(_u10_n14533 ), .A2(_u10_n14534 ), .A3(_u10_n14535 ), .A4(_u10_n14536 ), .ZN(_u10_n14527 ) );
NAND2_X1 _u10_U3038  ( .A1(1'b0), .A2(_u10_n11691 ), .ZN(_u10_n14529 ) );
NAND2_X1 _u10_U3037  ( .A1(1'b0), .A2(_u10_n11667 ), .ZN(_u10_n14530 ) );
NAND2_X1 _u10_U3036  ( .A1(1'b0), .A2(_u10_n11643 ), .ZN(_u10_n14531 ) );
NAND2_X1 _u10_U3035  ( .A1(1'b0), .A2(_u10_n11619 ), .ZN(_u10_n14532 ) );
NAND4_X1 _u10_U3034  ( .A1(_u10_n14529 ), .A2(_u10_n14530 ), .A3(_u10_n14531 ), .A4(_u10_n14532 ), .ZN(_u10_n14528 ) );
NOR4_X1 _u10_U3033  ( .A1(_u10_n14525 ), .A2(_u10_n14526 ), .A3(_u10_n14527 ), .A4(_u10_n14528 ), .ZN(_u10_n14524 ) );
NAND2_X1 _u10_U3032  ( .A1(_u10_n14523 ), .A2(_u10_n14524 ), .ZN(pointer_s[1]) );
NAND2_X1 _u10_U3031  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14519 ) );
NAND2_X1 _u10_U3030  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14520 ) );
NAND2_X1 _u10_U3029  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14521 ) );
NAND2_X1 _u10_U3028  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14522 ) );
NAND4_X1 _u10_U3027  ( .A1(_u10_n14519 ), .A2(_u10_n14520 ), .A3(_u10_n14521 ), .A4(_u10_n14522 ), .ZN(_u10_n14504 ) );
NAND2_X1 _u10_U3026  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14515 ) );
NAND2_X1 _u10_U3025  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14516 ) );
NAND2_X1 _u10_U3024  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14517 ) );
NAND2_X1 _u10_U3023  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14518 ) );
NAND4_X1 _u10_U3022  ( .A1(_u10_n14515 ), .A2(_u10_n14516 ), .A3(_u10_n14517 ), .A4(_u10_n14518 ), .ZN(_u10_n14505 ) );
NAND2_X1 _u10_U3021  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14511 ) );
NAND2_X1 _u10_U3020  ( .A1(1'b0), .A2(_u10_n12139 ), .ZN(_u10_n14512 ) );
NAND2_X1 _u10_U3019  ( .A1(1'b0), .A2(_u10_n12115 ), .ZN(_u10_n14513 ) );
NAND2_X1 _u10_U3018  ( .A1(1'b0), .A2(_u10_n12091 ), .ZN(_u10_n14514 ) );
NAND4_X1 _u10_U3017  ( .A1(_u10_n14511 ), .A2(_u10_n14512 ), .A3(_u10_n14513 ), .A4(_u10_n14514 ), .ZN(_u10_n14506 ) );
NAND2_X1 _u10_U3016  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14508 ) );
NAND2_X1 _u10_U3015  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14509 ) );
NAND2_X1 _u10_U3014  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14510 ) );
NAND3_X1 _u10_U3013  ( .A1(_u10_n14508 ), .A2(_u10_n14509 ), .A3(_u10_n14510 ), .ZN(_u10_n14507 ) );
NOR4_X1 _u10_U3012  ( .A1(_u10_n14504 ), .A2(_u10_n14505 ), .A3(_u10_n14506 ), .A4(_u10_n14507 ), .ZN(_u10_n14482 ) );
NAND2_X1 _u10_U3011  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14500 ) );
NAND2_X1 _u10_U3010  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14501 ) );
NAND2_X1 _u10_U3009  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14502 ) );
NAND2_X1 _u10_U3008  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14503 ) );
NAND4_X1 _u10_U3007  ( .A1(_u10_n14500 ), .A2(_u10_n14501 ), .A3(_u10_n14502 ), .A4(_u10_n14503 ), .ZN(_u10_n14484 ) );
NAND2_X1 _u10_U3006  ( .A1(1'b0), .A2(_u10_n11898 ), .ZN(_u10_n14496 ) );
NAND2_X1 _u10_U3005  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14497 ) );
NAND2_X1 _u10_U3004  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14498 ) );
NAND2_X1 _u10_U3003  ( .A1(1'b0), .A2(_u10_n11827 ), .ZN(_u10_n14499 ) );
NAND4_X1 _u10_U3002  ( .A1(_u10_n14496 ), .A2(_u10_n14497 ), .A3(_u10_n14498 ), .A4(_u10_n14499 ), .ZN(_u10_n14485 ) );
NAND2_X1 _u10_U3001  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14492 ) );
NAND2_X1 _u10_U3000  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14493 ) );
NAND2_X1 _u10_U2999  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14494 ) );
NAND2_X1 _u10_U2998  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14495 ) );
NAND4_X1 _u10_U2997  ( .A1(_u10_n14492 ), .A2(_u10_n14493 ), .A3(_u10_n14494 ), .A4(_u10_n14495 ), .ZN(_u10_n14486 ) );
NAND2_X1 _u10_U2996  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14488 ) );
NAND2_X1 _u10_U2995  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14489 ) );
NAND2_X1 _u10_U2994  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14490 ) );
NAND2_X1 _u10_U2993  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14491 ) );
NAND4_X1 _u10_U2992  ( .A1(_u10_n14488 ), .A2(_u10_n14489 ), .A3(_u10_n14490 ), .A4(_u10_n14491 ), .ZN(_u10_n14487 ) );
NOR4_X1 _u10_U2991  ( .A1(_u10_n14484 ), .A2(_u10_n14485 ), .A3(_u10_n14486 ), .A4(_u10_n14487 ), .ZN(_u10_n14483 ) );
NAND2_X1 _u10_U2990  ( .A1(_u10_n14482 ), .A2(_u10_n14483 ), .ZN(pointer_s[20]) );
NAND2_X1 _u10_U2989  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14478 ) );
NAND2_X1 _u10_U2988  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14479 ) );
NAND2_X1 _u10_U2987  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14480 ) );
NAND2_X1 _u10_U2986  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14481 ) );
NAND4_X1 _u10_U2985  ( .A1(_u10_n14478 ), .A2(_u10_n14479 ), .A3(_u10_n14480 ), .A4(_u10_n14481 ), .ZN(_u10_n14463 ) );
NAND2_X1 _u10_U2984  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14474 ) );
NAND2_X1 _u10_U2983  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14475 ) );
NAND2_X1 _u10_U2982  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14476 ) );
NAND2_X1 _u10_U2981  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14477 ) );
NAND4_X1 _u10_U2980  ( .A1(_u10_n14474 ), .A2(_u10_n14475 ), .A3(_u10_n14476 ), .A4(_u10_n14477 ), .ZN(_u10_n14464 ) );
NAND2_X1 _u10_U2979  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14470 ) );
NAND2_X1 _u10_U2978  ( .A1(1'b0), .A2(_u10_n12138 ), .ZN(_u10_n14471 ) );
NAND2_X1 _u10_U2977  ( .A1(1'b0), .A2(_u10_n12114 ), .ZN(_u10_n14472 ) );
NAND2_X1 _u10_U2976  ( .A1(1'b0), .A2(_u10_n12090 ), .ZN(_u10_n14473 ) );
NAND4_X1 _u10_U2975  ( .A1(_u10_n14470 ), .A2(_u10_n14471 ), .A3(_u10_n14472 ), .A4(_u10_n14473 ), .ZN(_u10_n14465 ) );
NAND2_X1 _u10_U2974  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14467 ) );
NAND2_X1 _u10_U2973  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14468 ) );
NAND2_X1 _u10_U2972  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14469 ) );
NAND3_X1 _u10_U2971  ( .A1(_u10_n14467 ), .A2(_u10_n14468 ), .A3(_u10_n14469 ), .ZN(_u10_n14466 ) );
NOR4_X1 _u10_U2970  ( .A1(_u10_n14463 ), .A2(_u10_n14464 ), .A3(_u10_n14465 ), .A4(_u10_n14466 ), .ZN(_u10_n14441 ) );
NAND2_X1 _u10_U2969  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14459 ) );
NAND2_X1 _u10_U2968  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14460 ) );
NAND2_X1 _u10_U2967  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14461 ) );
NAND2_X1 _u10_U2966  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14462 ) );
NAND4_X1 _u10_U2965  ( .A1(_u10_n14459 ), .A2(_u10_n14460 ), .A3(_u10_n14461 ), .A4(_u10_n14462 ), .ZN(_u10_n14443 ) );
NAND2_X1 _u10_U2964  ( .A1(1'b0), .A2(_u10_n11903 ), .ZN(_u10_n14455 ) );
NAND2_X1 _u10_U2963  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14456 ) );
NAND2_X1 _u10_U2962  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14457 ) );
NAND2_X1 _u10_U2961  ( .A1(1'b0), .A2(_u10_n11826 ), .ZN(_u10_n14458 ) );
NAND4_X1 _u10_U2960  ( .A1(_u10_n14455 ), .A2(_u10_n14456 ), .A3(_u10_n14457 ), .A4(_u10_n14458 ), .ZN(_u10_n14444 ) );
NAND2_X1 _u10_U2959  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14451 ) );
NAND2_X1 _u10_U2958  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14452 ) );
NAND2_X1 _u10_U2957  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14453 ) );
NAND2_X1 _u10_U2956  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14454 ) );
NAND4_X1 _u10_U2955  ( .A1(_u10_n14451 ), .A2(_u10_n14452 ), .A3(_u10_n14453 ), .A4(_u10_n14454 ), .ZN(_u10_n14445 ) );
NAND2_X1 _u10_U2954  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14447 ) );
NAND2_X1 _u10_U2953  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14448 ) );
NAND2_X1 _u10_U2952  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14449 ) );
NAND2_X1 _u10_U2951  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14450 ) );
NAND4_X1 _u10_U2950  ( .A1(_u10_n14447 ), .A2(_u10_n14448 ), .A3(_u10_n14449 ), .A4(_u10_n14450 ), .ZN(_u10_n14446 ) );
NOR4_X1 _u10_U2949  ( .A1(_u10_n14443 ), .A2(_u10_n14444 ), .A3(_u10_n14445 ), .A4(_u10_n14446 ), .ZN(_u10_n14442 ) );
NAND2_X1 _u10_U2948  ( .A1(_u10_n14441 ), .A2(_u10_n14442 ), .ZN(pointer_s[21]) );
NAND2_X1 _u10_U2947  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14437 ) );
NAND2_X1 _u10_U2946  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14438 ) );
NAND2_X1 _u10_U2945  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14439 ) );
NAND2_X1 _u10_U2944  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14440 ) );
NAND4_X1 _u10_U2943  ( .A1(_u10_n14437 ), .A2(_u10_n14438 ), .A3(_u10_n14439 ), .A4(_u10_n14440 ), .ZN(_u10_n14422 ) );
NAND2_X1 _u10_U2942  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14433 ) );
NAND2_X1 _u10_U2941  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14434 ) );
NAND2_X1 _u10_U2940  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14435 ) );
NAND2_X1 _u10_U2939  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14436 ) );
NAND4_X1 _u10_U2938  ( .A1(_u10_n14433 ), .A2(_u10_n14434 ), .A3(_u10_n14435 ), .A4(_u10_n14436 ), .ZN(_u10_n14423 ) );
NAND2_X1 _u10_U2937  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14429 ) );
NAND2_X1 _u10_U2936  ( .A1(1'b0), .A2(_u10_n12135 ), .ZN(_u10_n14430 ) );
NAND2_X1 _u10_U2935  ( .A1(1'b0), .A2(_u10_n12111 ), .ZN(_u10_n14431 ) );
NAND2_X1 _u10_U2934  ( .A1(1'b0), .A2(_u10_n12087 ), .ZN(_u10_n14432 ) );
NAND4_X1 _u10_U2933  ( .A1(_u10_n14429 ), .A2(_u10_n14430 ), .A3(_u10_n14431 ), .A4(_u10_n14432 ), .ZN(_u10_n14424 ) );
NAND2_X1 _u10_U2932  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14426 ) );
NAND2_X1 _u10_U2931  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14427 ) );
NAND2_X1 _u10_U2930  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14428 ) );
NAND3_X1 _u10_U2929  ( .A1(_u10_n14426 ), .A2(_u10_n14427 ), .A3(_u10_n14428 ), .ZN(_u10_n14425 ) );
NOR4_X1 _u10_U2928  ( .A1(_u10_n14422 ), .A2(_u10_n14423 ), .A3(_u10_n14424 ), .A4(_u10_n14425 ), .ZN(_u10_n14400 ) );
NAND2_X1 _u10_U2927  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14418 ) );
NAND2_X1 _u10_U2926  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14419 ) );
NAND2_X1 _u10_U2925  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14420 ) );
NAND2_X1 _u10_U2924  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14421 ) );
NAND4_X1 _u10_U2923  ( .A1(_u10_n14418 ), .A2(_u10_n14419 ), .A3(_u10_n14420 ), .A4(_u10_n14421 ), .ZN(_u10_n14402 ) );
NAND2_X1 _u10_U2922  ( .A1(1'b0), .A2(_u10_n12388 ), .ZN(_u10_n14414 ) );
NAND2_X1 _u10_U2921  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14415 ) );
NAND2_X1 _u10_U2920  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14416 ) );
NAND2_X1 _u10_U2919  ( .A1(1'b0), .A2(_u10_n11831 ), .ZN(_u10_n14417 ) );
NAND4_X1 _u10_U2918  ( .A1(_u10_n14414 ), .A2(_u10_n14415 ), .A3(_u10_n14416 ), .A4(_u10_n14417 ), .ZN(_u10_n14403 ) );
NAND2_X1 _u10_U2917  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14410 ) );
NAND2_X1 _u10_U2916  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14411 ) );
NAND2_X1 _u10_U2915  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14412 ) );
NAND2_X1 _u10_U2914  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14413 ) );
NAND4_X1 _u10_U2913  ( .A1(_u10_n14410 ), .A2(_u10_n14411 ), .A3(_u10_n14412 ), .A4(_u10_n14413 ), .ZN(_u10_n14404 ) );
NAND2_X1 _u10_U2912  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14406 ) );
NAND2_X1 _u10_U2911  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14407 ) );
NAND2_X1 _u10_U2910  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14408 ) );
NAND2_X1 _u10_U2909  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14409 ) );
NAND4_X1 _u10_U2908  ( .A1(_u10_n14406 ), .A2(_u10_n14407 ), .A3(_u10_n14408 ), .A4(_u10_n14409 ), .ZN(_u10_n14405 ) );
NOR4_X1 _u10_U2907  ( .A1(_u10_n14402 ), .A2(_u10_n14403 ), .A3(_u10_n14404 ), .A4(_u10_n14405 ), .ZN(_u10_n14401 ) );
NAND2_X1 _u10_U2906  ( .A1(_u10_n14400 ), .A2(_u10_n14401 ), .ZN(pointer_s[22]) );
NAND2_X1 _u10_U2905  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14396 ) );
NAND2_X1 _u10_U2904  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14397 ) );
NAND2_X1 _u10_U2903  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14398 ) );
NAND2_X1 _u10_U2902  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14399 ) );
NAND4_X1 _u10_U2901  ( .A1(_u10_n14396 ), .A2(_u10_n14397 ), .A3(_u10_n14398 ), .A4(_u10_n14399 ), .ZN(_u10_n14381 ) );
NAND2_X1 _u10_U2900  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14392 ) );
NAND2_X1 _u10_U2899  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14393 ) );
NAND2_X1 _u10_U2898  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14394 ) );
NAND2_X1 _u10_U2897  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14395 ) );
NAND4_X1 _u10_U2896  ( .A1(_u10_n14392 ), .A2(_u10_n14393 ), .A3(_u10_n14394 ), .A4(_u10_n14395 ), .ZN(_u10_n14382 ) );
NAND2_X1 _u10_U2895  ( .A1(1'b0), .A2(_u10_n12153 ), .ZN(_u10_n14388 ) );
NAND2_X1 _u10_U2894  ( .A1(1'b0), .A2(_u10_n12136 ), .ZN(_u10_n14389 ) );
NAND2_X1 _u10_U2893  ( .A1(1'b0), .A2(_u10_n12112 ), .ZN(_u10_n14390 ) );
NAND2_X1 _u10_U2892  ( .A1(1'b0), .A2(_u10_n12088 ), .ZN(_u10_n14391 ) );
NAND4_X1 _u10_U2891  ( .A1(_u10_n14388 ), .A2(_u10_n14389 ), .A3(_u10_n14390 ), .A4(_u10_n14391 ), .ZN(_u10_n14383 ) );
NAND2_X1 _u10_U2890  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14385 ) );
NAND2_X1 _u10_U2889  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14386 ) );
NAND2_X1 _u10_U2888  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14387 ) );
NAND3_X1 _u10_U2887  ( .A1(_u10_n14385 ), .A2(_u10_n14386 ), .A3(_u10_n14387 ), .ZN(_u10_n14384 ) );
NOR4_X1 _u10_U2886  ( .A1(_u10_n14381 ), .A2(_u10_n14382 ), .A3(_u10_n14383 ), .A4(_u10_n14384 ), .ZN(_u10_n14359 ) );
NAND2_X1 _u10_U2885  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14377 ) );
NAND2_X1 _u10_U2884  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14378 ) );
NAND2_X1 _u10_U2883  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14379 ) );
NAND2_X1 _u10_U2882  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14380 ) );
NAND4_X1 _u10_U2881  ( .A1(_u10_n14377 ), .A2(_u10_n14378 ), .A3(_u10_n14379 ), .A4(_u10_n14380 ), .ZN(_u10_n14361 ) );
NAND2_X1 _u10_U2880  ( .A1(1'b0), .A2(_u10_n11897 ), .ZN(_u10_n14373 ) );
NAND2_X1 _u10_U2879  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14374 ) );
NAND2_X1 _u10_U2878  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14375 ) );
NAND2_X1 _u10_U2877  ( .A1(1'b0), .A2(_u10_n12385 ), .ZN(_u10_n14376 ) );
NAND4_X1 _u10_U2876  ( .A1(_u10_n14373 ), .A2(_u10_n14374 ), .A3(_u10_n14375 ), .A4(_u10_n14376 ), .ZN(_u10_n14362 ) );
NAND2_X1 _u10_U2875  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14369 ) );
NAND2_X1 _u10_U2874  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14370 ) );
NAND2_X1 _u10_U2873  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14371 ) );
NAND2_X1 _u10_U2872  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14372 ) );
NAND4_X1 _u10_U2871  ( .A1(_u10_n14369 ), .A2(_u10_n14370 ), .A3(_u10_n14371 ), .A4(_u10_n14372 ), .ZN(_u10_n14363 ) );
NAND2_X1 _u10_U2870  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14365 ) );
NAND2_X1 _u10_U2869  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14366 ) );
NAND2_X1 _u10_U2868  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14367 ) );
NAND2_X1 _u10_U2867  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14368 ) );
NAND4_X1 _u10_U2866  ( .A1(_u10_n14365 ), .A2(_u10_n14366 ), .A3(_u10_n14367 ), .A4(_u10_n14368 ), .ZN(_u10_n14364 ) );
NOR4_X1 _u10_U2865  ( .A1(_u10_n14361 ), .A2(_u10_n14362 ), .A3(_u10_n14363 ), .A4(_u10_n14364 ), .ZN(_u10_n14360 ) );
NAND2_X1 _u10_U2864  ( .A1(_u10_n14359 ), .A2(_u10_n14360 ), .ZN(pointer_s[23]) );
NAND2_X1 _u10_U2863  ( .A1(1'b0), .A2(_u10_n12347 ), .ZN(_u10_n14355 ) );
NAND2_X1 _u10_U2862  ( .A1(1'b0), .A2(_u10_n12323 ), .ZN(_u10_n14356 ) );
NAND2_X1 _u10_U2861  ( .A1(1'b0), .A2(_u10_n12300 ), .ZN(_u10_n14357 ) );
NAND2_X1 _u10_U2860  ( .A1(1'b0), .A2(_u10_n12276 ), .ZN(_u10_n14358 ) );
NAND4_X1 _u10_U2859  ( .A1(_u10_n14355 ), .A2(_u10_n14356 ), .A3(_u10_n14357 ), .A4(_u10_n14358 ), .ZN(_u10_n14340 ) );
NAND2_X1 _u10_U2858  ( .A1(1'b0), .A2(_u10_n12251 ), .ZN(_u10_n14351 ) );
NAND2_X1 _u10_U2857  ( .A1(1'b0), .A2(_u10_n12227 ), .ZN(_u10_n14352 ) );
NAND2_X1 _u10_U2856  ( .A1(1'b0), .A2(_u10_n12201 ), .ZN(_u10_n14353 ) );
NAND2_X1 _u10_U2855  ( .A1(1'b0), .A2(_u10_n12179 ), .ZN(_u10_n14354 ) );
NAND4_X1 _u10_U2854  ( .A1(_u10_n14351 ), .A2(_u10_n14352 ), .A3(_u10_n14353 ), .A4(_u10_n14354 ), .ZN(_u10_n14341 ) );
NAND2_X1 _u10_U2853  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n14347 ) );
NAND2_X1 _u10_U2852  ( .A1(1'b0), .A2(_u10_n12138 ), .ZN(_u10_n14348 ) );
NAND2_X1 _u10_U2851  ( .A1(1'b0), .A2(_u10_n12114 ), .ZN(_u10_n14349 ) );
NAND2_X1 _u10_U2850  ( .A1(1'b0), .A2(_u10_n12090 ), .ZN(_u10_n14350 ) );
NAND4_X1 _u10_U2849  ( .A1(_u10_n14347 ), .A2(_u10_n14348 ), .A3(_u10_n14349 ), .A4(_u10_n14350 ), .ZN(_u10_n14342 ) );
NAND2_X1 _u10_U2848  ( .A1(1'b0), .A2(_u10_n12057 ), .ZN(_u10_n14344 ) );
NAND2_X1 _u10_U2847  ( .A1(1'b0), .A2(_u10_n12033 ), .ZN(_u10_n14345 ) );
NAND2_X1 _u10_U2846  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14346 ) );
NAND3_X1 _u10_U2845  ( .A1(_u10_n14344 ), .A2(_u10_n14345 ), .A3(_u10_n14346 ), .ZN(_u10_n14343 ) );
NOR4_X1 _u10_U2844  ( .A1(_u10_n14340 ), .A2(_u10_n14341 ), .A3(_u10_n14342 ), .A4(_u10_n14343 ), .ZN(_u10_n14318 ) );
NAND2_X1 _u10_U2843  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14336 ) );
NAND2_X1 _u10_U2842  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14337 ) );
NAND2_X1 _u10_U2841  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14338 ) );
NAND2_X1 _u10_U2840  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14339 ) );
NAND4_X1 _u10_U2839  ( .A1(_u10_n14336 ), .A2(_u10_n14337 ), .A3(_u10_n14338 ), .A4(_u10_n14339 ), .ZN(_u10_n14320 ) );
NAND2_X1 _u10_U2838  ( .A1(1'b0), .A2(_u10_n11900 ), .ZN(_u10_n14332 ) );
NAND2_X1 _u10_U2837  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14333 ) );
NAND2_X1 _u10_U2836  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14334 ) );
NAND2_X1 _u10_U2835  ( .A1(1'b0), .A2(_u10_n11825 ), .ZN(_u10_n14335 ) );
NAND4_X1 _u10_U2834  ( .A1(_u10_n14332 ), .A2(_u10_n14333 ), .A3(_u10_n14334 ), .A4(_u10_n14335 ), .ZN(_u10_n14321 ) );
NAND2_X1 _u10_U2833  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14328 ) );
NAND2_X1 _u10_U2832  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14329 ) );
NAND2_X1 _u10_U2831  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14330 ) );
NAND2_X1 _u10_U2830  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14331 ) );
NAND4_X1 _u10_U2829  ( .A1(_u10_n14328 ), .A2(_u10_n14329 ), .A3(_u10_n14330 ), .A4(_u10_n14331 ), .ZN(_u10_n14322 ) );
NAND2_X1 _u10_U2828  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14324 ) );
NAND2_X1 _u10_U2827  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14325 ) );
NAND2_X1 _u10_U2826  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14326 ) );
NAND2_X1 _u10_U2825  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14327 ) );
NAND4_X1 _u10_U2824  ( .A1(_u10_n14324 ), .A2(_u10_n14325 ), .A3(_u10_n14326 ), .A4(_u10_n14327 ), .ZN(_u10_n14323 ) );
NOR4_X1 _u10_U2823  ( .A1(_u10_n14320 ), .A2(_u10_n14321 ), .A3(_u10_n14322 ), .A4(_u10_n14323 ), .ZN(_u10_n14319 ) );
NAND2_X1 _u10_U2822  ( .A1(_u10_n14318 ), .A2(_u10_n14319 ), .ZN(pointer_s[24]) );
NAND2_X1 _u10_U2821  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n14314 ) );
NAND2_X1 _u10_U2820  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n14315 ) );
NAND2_X1 _u10_U2819  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n14316 ) );
NAND2_X1 _u10_U2818  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n14317 ) );
NAND4_X1 _u10_U2817  ( .A1(_u10_n14314 ), .A2(_u10_n14315 ), .A3(_u10_n14316 ), .A4(_u10_n14317 ), .ZN(_u10_n14299 ) );
NAND2_X1 _u10_U2816  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n14310 ) );
NAND2_X1 _u10_U2815  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n14311 ) );
NAND2_X1 _u10_U2814  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n14312 ) );
NAND2_X1 _u10_U2813  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n14313 ) );
NAND4_X1 _u10_U2812  ( .A1(_u10_n14310 ), .A2(_u10_n14311 ), .A3(_u10_n14312 ), .A4(_u10_n14313 ), .ZN(_u10_n14300 ) );
NAND2_X1 _u10_U2811  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n14306 ) );
NAND2_X1 _u10_U2810  ( .A1(1'b0), .A2(_u10_n12135 ), .ZN(_u10_n14307 ) );
NAND2_X1 _u10_U2809  ( .A1(1'b0), .A2(_u10_n12111 ), .ZN(_u10_n14308 ) );
NAND2_X1 _u10_U2808  ( .A1(1'b0), .A2(_u10_n12087 ), .ZN(_u10_n14309 ) );
NAND4_X1 _u10_U2807  ( .A1(_u10_n14306 ), .A2(_u10_n14307 ), .A3(_u10_n14308 ), .A4(_u10_n14309 ), .ZN(_u10_n14301 ) );
NAND2_X1 _u10_U2806  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n14303 ) );
NAND2_X1 _u10_U2805  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n14304 ) );
NAND2_X1 _u10_U2804  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14305 ) );
NAND3_X1 _u10_U2803  ( .A1(_u10_n14303 ), .A2(_u10_n14304 ), .A3(_u10_n14305 ), .ZN(_u10_n14302 ) );
NOR4_X1 _u10_U2802  ( .A1(_u10_n14299 ), .A2(_u10_n14300 ), .A3(_u10_n14301 ), .A4(_u10_n14302 ), .ZN(_u10_n14277 ) );
NAND2_X1 _u10_U2801  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14295 ) );
NAND2_X1 _u10_U2800  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14296 ) );
NAND2_X1 _u10_U2799  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14297 ) );
NAND2_X1 _u10_U2798  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14298 ) );
NAND4_X1 _u10_U2797  ( .A1(_u10_n14295 ), .A2(_u10_n14296 ), .A3(_u10_n14297 ), .A4(_u10_n14298 ), .ZN(_u10_n14279 ) );
NAND2_X1 _u10_U2796  ( .A1(1'b0), .A2(_u10_n11901 ), .ZN(_u10_n14291 ) );
NAND2_X1 _u10_U2795  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14292 ) );
NAND2_X1 _u10_U2794  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14293 ) );
NAND2_X1 _u10_U2793  ( .A1(1'b0), .A2(_u10_n12385 ), .ZN(_u10_n14294 ) );
NAND4_X1 _u10_U2792  ( .A1(_u10_n14291 ), .A2(_u10_n14292 ), .A3(_u10_n14293 ), .A4(_u10_n14294 ), .ZN(_u10_n14280 ) );
NAND2_X1 _u10_U2791  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14287 ) );
NAND2_X1 _u10_U2790  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14288 ) );
NAND2_X1 _u10_U2789  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14289 ) );
NAND2_X1 _u10_U2788  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14290 ) );
NAND4_X1 _u10_U2787  ( .A1(_u10_n14287 ), .A2(_u10_n14288 ), .A3(_u10_n14289 ), .A4(_u10_n14290 ), .ZN(_u10_n14281 ) );
NAND2_X1 _u10_U2786  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14283 ) );
NAND2_X1 _u10_U2785  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14284 ) );
NAND2_X1 _u10_U2784  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14285 ) );
NAND2_X1 _u10_U2783  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14286 ) );
NAND4_X1 _u10_U2782  ( .A1(_u10_n14283 ), .A2(_u10_n14284 ), .A3(_u10_n14285 ), .A4(_u10_n14286 ), .ZN(_u10_n14282 ) );
NOR4_X1 _u10_U2781  ( .A1(_u10_n14279 ), .A2(_u10_n14280 ), .A3(_u10_n14281 ), .A4(_u10_n14282 ), .ZN(_u10_n14278 ) );
NAND2_X1 _u10_U2780  ( .A1(_u10_n14277 ), .A2(_u10_n14278 ), .ZN(pointer_s[25]) );
NAND2_X1 _u10_U2779  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n14273 ) );
NAND2_X1 _u10_U2778  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n14274 ) );
NAND2_X1 _u10_U2777  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n14275 ) );
NAND2_X1 _u10_U2776  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n14276 ) );
NAND4_X1 _u10_U2775  ( .A1(_u10_n14273 ), .A2(_u10_n14274 ), .A3(_u10_n14275 ), .A4(_u10_n14276 ), .ZN(_u10_n14258 ) );
NAND2_X1 _u10_U2774  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n14269 ) );
NAND2_X1 _u10_U2773  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n14270 ) );
NAND2_X1 _u10_U2772  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n14271 ) );
NAND2_X1 _u10_U2771  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n14272 ) );
NAND4_X1 _u10_U2770  ( .A1(_u10_n14269 ), .A2(_u10_n14270 ), .A3(_u10_n14271 ), .A4(_u10_n14272 ), .ZN(_u10_n14259 ) );
NAND2_X1 _u10_U2769  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n14265 ) );
NAND2_X1 _u10_U2768  ( .A1(1'b0), .A2(_u10_n12136 ), .ZN(_u10_n14266 ) );
NAND2_X1 _u10_U2767  ( .A1(1'b0), .A2(_u10_n12112 ), .ZN(_u10_n14267 ) );
NAND2_X1 _u10_U2766  ( .A1(1'b0), .A2(_u10_n12088 ), .ZN(_u10_n14268 ) );
NAND4_X1 _u10_U2765  ( .A1(_u10_n14265 ), .A2(_u10_n14266 ), .A3(_u10_n14267 ), .A4(_u10_n14268 ), .ZN(_u10_n14260 ) );
NAND2_X1 _u10_U2764  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n14262 ) );
NAND2_X1 _u10_U2763  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n14263 ) );
NAND2_X1 _u10_U2762  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14264 ) );
NAND3_X1 _u10_U2761  ( .A1(_u10_n14262 ), .A2(_u10_n14263 ), .A3(_u10_n14264 ), .ZN(_u10_n14261 ) );
NOR4_X1 _u10_U2760  ( .A1(_u10_n14258 ), .A2(_u10_n14259 ), .A3(_u10_n14260 ), .A4(_u10_n14261 ), .ZN(_u10_n14236 ) );
NAND2_X1 _u10_U2759  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14254 ) );
NAND2_X1 _u10_U2758  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14255 ) );
NAND2_X1 _u10_U2757  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14256 ) );
NAND2_X1 _u10_U2756  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14257 ) );
NAND4_X1 _u10_U2755  ( .A1(_u10_n14254 ), .A2(_u10_n14255 ), .A3(_u10_n14256 ), .A4(_u10_n14257 ), .ZN(_u10_n14238 ) );
NAND2_X1 _u10_U2754  ( .A1(1'b0), .A2(_u10_n11902 ), .ZN(_u10_n14250 ) );
NAND2_X1 _u10_U2753  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14251 ) );
NAND2_X1 _u10_U2752  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14252 ) );
NAND2_X1 _u10_U2751  ( .A1(1'b0), .A2(_u10_n11828 ), .ZN(_u10_n14253 ) );
NAND4_X1 _u10_U2750  ( .A1(_u10_n14250 ), .A2(_u10_n14251 ), .A3(_u10_n14252 ), .A4(_u10_n14253 ), .ZN(_u10_n14239 ) );
NAND2_X1 _u10_U2749  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14246 ) );
NAND2_X1 _u10_U2748  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14247 ) );
NAND2_X1 _u10_U2747  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14248 ) );
NAND2_X1 _u10_U2746  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14249 ) );
NAND4_X1 _u10_U2745  ( .A1(_u10_n14246 ), .A2(_u10_n14247 ), .A3(_u10_n14248 ), .A4(_u10_n14249 ), .ZN(_u10_n14240 ) );
NAND2_X1 _u10_U2744  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14242 ) );
NAND2_X1 _u10_U2743  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14243 ) );
NAND2_X1 _u10_U2742  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14244 ) );
NAND2_X1 _u10_U2741  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14245 ) );
NAND4_X1 _u10_U2740  ( .A1(_u10_n14242 ), .A2(_u10_n14243 ), .A3(_u10_n14244 ), .A4(_u10_n14245 ), .ZN(_u10_n14241 ) );
NOR4_X1 _u10_U2739  ( .A1(_u10_n14238 ), .A2(_u10_n14239 ), .A3(_u10_n14240 ), .A4(_u10_n14241 ), .ZN(_u10_n14237 ) );
NAND2_X1 _u10_U2738  ( .A1(_u10_n14236 ), .A2(_u10_n14237 ), .ZN(pointer_s[26]) );
NAND2_X1 _u10_U2737  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n14232 ) );
NAND2_X1 _u10_U2736  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n14233 ) );
NAND2_X1 _u10_U2735  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n14234 ) );
NAND2_X1 _u10_U2734  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n14235 ) );
NAND4_X1 _u10_U2733  ( .A1(_u10_n14232 ), .A2(_u10_n14233 ), .A3(_u10_n14234 ), .A4(_u10_n14235 ), .ZN(_u10_n14217 ) );
NAND2_X1 _u10_U2732  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n14228 ) );
NAND2_X1 _u10_U2731  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n14229 ) );
NAND2_X1 _u10_U2730  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n14230 ) );
NAND2_X1 _u10_U2729  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n14231 ) );
NAND4_X1 _u10_U2728  ( .A1(_u10_n14228 ), .A2(_u10_n14229 ), .A3(_u10_n14230 ), .A4(_u10_n14231 ), .ZN(_u10_n14218 ) );
NAND2_X1 _u10_U2727  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n14224 ) );
NAND2_X1 _u10_U2726  ( .A1(1'b0), .A2(_u10_n12413 ), .ZN(_u10_n14225 ) );
NAND2_X1 _u10_U2725  ( .A1(1'b0), .A2(_u10_n12412 ), .ZN(_u10_n14226 ) );
NAND2_X1 _u10_U2724  ( .A1(1'b0), .A2(_u10_n12411 ), .ZN(_u10_n14227 ) );
NAND4_X1 _u10_U2723  ( .A1(_u10_n14224 ), .A2(_u10_n14225 ), .A3(_u10_n14226 ), .A4(_u10_n14227 ), .ZN(_u10_n14219 ) );
NAND2_X1 _u10_U2722  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n14221 ) );
NAND2_X1 _u10_U2721  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n14222 ) );
NAND2_X1 _u10_U2720  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14223 ) );
NAND3_X1 _u10_U2719  ( .A1(_u10_n14221 ), .A2(_u10_n14222 ), .A3(_u10_n14223 ), .ZN(_u10_n14220 ) );
NOR4_X1 _u10_U2718  ( .A1(_u10_n14217 ), .A2(_u10_n14218 ), .A3(_u10_n14219 ), .A4(_u10_n14220 ), .ZN(_u10_n14195 ) );
NAND2_X1 _u10_U2717  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14213 ) );
NAND2_X1 _u10_U2716  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14214 ) );
NAND2_X1 _u10_U2715  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14215 ) );
NAND2_X1 _u10_U2714  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14216 ) );
NAND4_X1 _u10_U2713  ( .A1(_u10_n14213 ), .A2(_u10_n14214 ), .A3(_u10_n14215 ), .A4(_u10_n14216 ), .ZN(_u10_n14197 ) );
NAND2_X1 _u10_U2712  ( .A1(1'b0), .A2(_u10_n11898 ), .ZN(_u10_n14209 ) );
NAND2_X1 _u10_U2711  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14210 ) );
NAND2_X1 _u10_U2710  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14211 ) );
NAND2_X1 _u10_U2709  ( .A1(1'b0), .A2(_u10_n11829 ), .ZN(_u10_n14212 ) );
NAND4_X1 _u10_U2708  ( .A1(_u10_n14209 ), .A2(_u10_n14210 ), .A3(_u10_n14211 ), .A4(_u10_n14212 ), .ZN(_u10_n14198 ) );
NAND2_X1 _u10_U2707  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14205 ) );
NAND2_X1 _u10_U2706  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14206 ) );
NAND2_X1 _u10_U2705  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14207 ) );
NAND2_X1 _u10_U2704  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14208 ) );
NAND4_X1 _u10_U2703  ( .A1(_u10_n14205 ), .A2(_u10_n14206 ), .A3(_u10_n14207 ), .A4(_u10_n14208 ), .ZN(_u10_n14199 ) );
NAND2_X1 _u10_U2702  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14201 ) );
NAND2_X1 _u10_U2701  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14202 ) );
NAND2_X1 _u10_U2700  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14203 ) );
NAND2_X1 _u10_U2699  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14204 ) );
NAND4_X1 _u10_U2698  ( .A1(_u10_n14201 ), .A2(_u10_n14202 ), .A3(_u10_n14203 ), .A4(_u10_n14204 ), .ZN(_u10_n14200 ) );
NOR4_X1 _u10_U2697  ( .A1(_u10_n14197 ), .A2(_u10_n14198 ), .A3(_u10_n14199 ), .A4(_u10_n14200 ), .ZN(_u10_n14196 ) );
NAND2_X1 _u10_U2696  ( .A1(_u10_n14195 ), .A2(_u10_n14196 ), .ZN(pointer_s[27]) );
NAND2_X1 _u10_U2695  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n14191 ) );
NAND2_X1 _u10_U2694  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n14192 ) );
NAND2_X1 _u10_U2693  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n14193 ) );
NAND2_X1 _u10_U2692  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n14194 ) );
NAND4_X1 _u10_U2691  ( .A1(_u10_n14191 ), .A2(_u10_n14192 ), .A3(_u10_n14193 ), .A4(_u10_n14194 ), .ZN(_u10_n14176 ) );
NAND2_X1 _u10_U2690  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n14187 ) );
NAND2_X1 _u10_U2689  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n14188 ) );
NAND2_X1 _u10_U2688  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n14189 ) );
NAND2_X1 _u10_U2687  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n14190 ) );
NAND4_X1 _u10_U2686  ( .A1(_u10_n14187 ), .A2(_u10_n14188 ), .A3(_u10_n14189 ), .A4(_u10_n14190 ), .ZN(_u10_n14177 ) );
NAND2_X1 _u10_U2685  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n14183 ) );
NAND2_X1 _u10_U2684  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n14184 ) );
NAND2_X1 _u10_U2683  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n14185 ) );
NAND2_X1 _u10_U2682  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n14186 ) );
NAND4_X1 _u10_U2681  ( .A1(_u10_n14183 ), .A2(_u10_n14184 ), .A3(_u10_n14185 ), .A4(_u10_n14186 ), .ZN(_u10_n14178 ) );
NAND2_X1 _u10_U2680  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n14180 ) );
NAND2_X1 _u10_U2679  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n14181 ) );
NAND2_X1 _u10_U2678  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14182 ) );
NAND3_X1 _u10_U2677  ( .A1(_u10_n14180 ), .A2(_u10_n14181 ), .A3(_u10_n14182 ), .ZN(_u10_n14179 ) );
NOR4_X1 _u10_U2676  ( .A1(_u10_n14176 ), .A2(_u10_n14177 ), .A3(_u10_n14178 ), .A4(_u10_n14179 ), .ZN(_u10_n14154 ) );
NAND2_X1 _u10_U2675  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14172 ) );
NAND2_X1 _u10_U2674  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14173 ) );
NAND2_X1 _u10_U2673  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14174 ) );
NAND2_X1 _u10_U2672  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14175 ) );
NAND4_X1 _u10_U2671  ( .A1(_u10_n14172 ), .A2(_u10_n14173 ), .A3(_u10_n14174 ), .A4(_u10_n14175 ), .ZN(_u10_n14156 ) );
NAND2_X1 _u10_U2670  ( .A1(1'b0), .A2(_u10_n11899 ), .ZN(_u10_n14168 ) );
NAND2_X1 _u10_U2669  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14169 ) );
NAND2_X1 _u10_U2668  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14170 ) );
NAND2_X1 _u10_U2667  ( .A1(1'b0), .A2(_u10_n11830 ), .ZN(_u10_n14171 ) );
NAND4_X1 _u10_U2666  ( .A1(_u10_n14168 ), .A2(_u10_n14169 ), .A3(_u10_n14170 ), .A4(_u10_n14171 ), .ZN(_u10_n14157 ) );
NAND2_X1 _u10_U2665  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14164 ) );
NAND2_X1 _u10_U2664  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14165 ) );
NAND2_X1 _u10_U2663  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14166 ) );
NAND2_X1 _u10_U2662  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14167 ) );
NAND4_X1 _u10_U2661  ( .A1(_u10_n14164 ), .A2(_u10_n14165 ), .A3(_u10_n14166 ), .A4(_u10_n14167 ), .ZN(_u10_n14158 ) );
NAND2_X1 _u10_U2660  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14160 ) );
NAND2_X1 _u10_U2659  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14161 ) );
NAND2_X1 _u10_U2658  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14162 ) );
NAND2_X1 _u10_U2657  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14163 ) );
NAND4_X1 _u10_U2656  ( .A1(_u10_n14160 ), .A2(_u10_n14161 ), .A3(_u10_n14162 ), .A4(_u10_n14163 ), .ZN(_u10_n14159 ) );
NOR4_X1 _u10_U2655  ( .A1(_u10_n14156 ), .A2(_u10_n14157 ), .A3(_u10_n14158 ), .A4(_u10_n14159 ), .ZN(_u10_n14155 ) );
NAND2_X1 _u10_U2654  ( .A1(_u10_n14154 ), .A2(_u10_n14155 ), .ZN(pointer_s[28]) );
NAND2_X1 _u10_U2653  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n14150 ) );
NAND2_X1 _u10_U2652  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n14151 ) );
NAND2_X1 _u10_U2651  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n14152 ) );
NAND2_X1 _u10_U2650  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n14153 ) );
NAND4_X1 _u10_U2649  ( .A1(_u10_n14150 ), .A2(_u10_n14151 ), .A3(_u10_n14152 ), .A4(_u10_n14153 ), .ZN(_u10_n14135 ) );
NAND2_X1 _u10_U2648  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n14146 ) );
NAND2_X1 _u10_U2647  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n14147 ) );
NAND2_X1 _u10_U2646  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n14148 ) );
NAND2_X1 _u10_U2645  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n14149 ) );
NAND4_X1 _u10_U2644  ( .A1(_u10_n14146 ), .A2(_u10_n14147 ), .A3(_u10_n14148 ), .A4(_u10_n14149 ), .ZN(_u10_n14136 ) );
NAND2_X1 _u10_U2643  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n14142 ) );
NAND2_X1 _u10_U2642  ( .A1(1'b0), .A2(_u10_n12140 ), .ZN(_u10_n14143 ) );
NAND2_X1 _u10_U2641  ( .A1(1'b0), .A2(_u10_n12116 ), .ZN(_u10_n14144 ) );
NAND2_X1 _u10_U2640  ( .A1(1'b0), .A2(_u10_n12092 ), .ZN(_u10_n14145 ) );
NAND4_X1 _u10_U2639  ( .A1(_u10_n14142 ), .A2(_u10_n14143 ), .A3(_u10_n14144 ), .A4(_u10_n14145 ), .ZN(_u10_n14137 ) );
NAND2_X1 _u10_U2638  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n14139 ) );
NAND2_X1 _u10_U2637  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n14140 ) );
NAND2_X1 _u10_U2636  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14141 ) );
NAND3_X1 _u10_U2635  ( .A1(_u10_n14139 ), .A2(_u10_n14140 ), .A3(_u10_n14141 ), .ZN(_u10_n14138 ) );
NOR4_X1 _u10_U2634  ( .A1(_u10_n14135 ), .A2(_u10_n14136 ), .A3(_u10_n14137 ), .A4(_u10_n14138 ), .ZN(_u10_n14113 ) );
NAND2_X1 _u10_U2633  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14131 ) );
NAND2_X1 _u10_U2632  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14132 ) );
NAND2_X1 _u10_U2631  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14133 ) );
NAND2_X1 _u10_U2630  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14134 ) );
NAND4_X1 _u10_U2629  ( .A1(_u10_n14131 ), .A2(_u10_n14132 ), .A3(_u10_n14133 ), .A4(_u10_n14134 ), .ZN(_u10_n14115 ) );
NAND2_X1 _u10_U2628  ( .A1(1'b0), .A2(_u10_n11898 ), .ZN(_u10_n14127 ) );
NAND2_X1 _u10_U2627  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14128 ) );
NAND2_X1 _u10_U2626  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14129 ) );
NAND2_X1 _u10_U2625  ( .A1(1'b0), .A2(_u10_n11827 ), .ZN(_u10_n14130 ) );
NAND4_X1 _u10_U2624  ( .A1(_u10_n14127 ), .A2(_u10_n14128 ), .A3(_u10_n14129 ), .A4(_u10_n14130 ), .ZN(_u10_n14116 ) );
NAND2_X1 _u10_U2623  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14123 ) );
NAND2_X1 _u10_U2622  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14124 ) );
NAND2_X1 _u10_U2621  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14125 ) );
NAND2_X1 _u10_U2620  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14126 ) );
NAND4_X1 _u10_U2619  ( .A1(_u10_n14123 ), .A2(_u10_n14124 ), .A3(_u10_n14125 ), .A4(_u10_n14126 ), .ZN(_u10_n14117 ) );
NAND2_X1 _u10_U2618  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14119 ) );
NAND2_X1 _u10_U2617  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14120 ) );
NAND2_X1 _u10_U2616  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14121 ) );
NAND2_X1 _u10_U2615  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14122 ) );
NAND4_X1 _u10_U2614  ( .A1(_u10_n14119 ), .A2(_u10_n14120 ), .A3(_u10_n14121 ), .A4(_u10_n14122 ), .ZN(_u10_n14118 ) );
NOR4_X1 _u10_U2613  ( .A1(_u10_n14115 ), .A2(_u10_n14116 ), .A3(_u10_n14117 ), .A4(_u10_n14118 ), .ZN(_u10_n14114 ) );
NAND2_X1 _u10_U2612  ( .A1(_u10_n14113 ), .A2(_u10_n14114 ), .ZN(pointer_s[29]) );
NAND2_X1 _u10_U2611  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n14109 ) );
NAND2_X1 _u10_U2610  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n14110 ) );
NAND2_X1 _u10_U2609  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n14111 ) );
NAND2_X1 _u10_U2608  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n14112 ) );
NAND4_X1 _u10_U2607  ( .A1(_u10_n14109 ), .A2(_u10_n14110 ), .A3(_u10_n14111 ), .A4(_u10_n14112 ), .ZN(_u10_n14094 ) );
NAND2_X1 _u10_U2606  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n14105 ) );
NAND2_X1 _u10_U2605  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n14106 ) );
NAND2_X1 _u10_U2604  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n14107 ) );
NAND2_X1 _u10_U2603  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n14108 ) );
NAND4_X1 _u10_U2602  ( .A1(_u10_n14105 ), .A2(_u10_n14106 ), .A3(_u10_n14107 ), .A4(_u10_n14108 ), .ZN(_u10_n14095 ) );
NAND2_X1 _u10_U2601  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n14101 ) );
NAND2_X1 _u10_U2600  ( .A1(1'b0), .A2(_u10_n12413 ), .ZN(_u10_n14102 ) );
NAND2_X1 _u10_U2599  ( .A1(1'b0), .A2(_u10_n12412 ), .ZN(_u10_n14103 ) );
NAND2_X1 _u10_U2598  ( .A1(1'b0), .A2(_u10_n12411 ), .ZN(_u10_n14104 ) );
NAND4_X1 _u10_U2597  ( .A1(_u10_n14101 ), .A2(_u10_n14102 ), .A3(_u10_n14103 ), .A4(_u10_n14104 ), .ZN(_u10_n14096 ) );
NAND2_X1 _u10_U2596  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n14098 ) );
NAND2_X1 _u10_U2595  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n14099 ) );
NAND2_X1 _u10_U2594  ( .A1(1'b0), .A2(_u10_n12016 ), .ZN(_u10_n14100 ) );
NAND3_X1 _u10_U2593  ( .A1(_u10_n14098 ), .A2(_u10_n14099 ), .A3(_u10_n14100 ), .ZN(_u10_n14097 ) );
NOR4_X1 _u10_U2592  ( .A1(_u10_n14094 ), .A2(_u10_n14095 ), .A3(_u10_n14096 ), .A4(_u10_n14097 ), .ZN(_u10_n14072 ) );
NAND2_X1 _u10_U2591  ( .A1(1'b0), .A2(_u10_n11980 ), .ZN(_u10_n14090 ) );
NAND2_X1 _u10_U2590  ( .A1(1'b0), .A2(_u10_n11956 ), .ZN(_u10_n14091 ) );
NAND2_X1 _u10_U2589  ( .A1(1'b0), .A2(_u10_n11935 ), .ZN(_u10_n14092 ) );
NAND2_X1 _u10_U2588  ( .A1(1'b0), .A2(_u10_n11911 ), .ZN(_u10_n14093 ) );
NAND4_X1 _u10_U2587  ( .A1(_u10_n14090 ), .A2(_u10_n14091 ), .A3(_u10_n14092 ), .A4(_u10_n14093 ), .ZN(_u10_n14074 ) );
NAND2_X1 _u10_U2586  ( .A1(1'b0), .A2(_u10_n11903 ), .ZN(_u10_n14086 ) );
NAND2_X1 _u10_U2585  ( .A1(1'b0), .A2(_u10_n11860 ), .ZN(_u10_n14087 ) );
NAND2_X1 _u10_U2584  ( .A1(1'b0), .A2(_u10_n11836 ), .ZN(_u10_n14088 ) );
NAND2_X1 _u10_U2583  ( .A1(1'b0), .A2(_u10_n11825 ), .ZN(_u10_n14089 ) );
NAND4_X1 _u10_U2582  ( .A1(_u10_n14086 ), .A2(_u10_n14087 ), .A3(_u10_n14088 ), .A4(_u10_n14089 ), .ZN(_u10_n14075 ) );
NAND2_X1 _u10_U2581  ( .A1(1'b0), .A2(_u10_n11788 ), .ZN(_u10_n14082 ) );
NAND2_X1 _u10_U2580  ( .A1(1'b0), .A2(_u10_n11766 ), .ZN(_u10_n14083 ) );
NAND2_X1 _u10_U2579  ( .A1(1'b0), .A2(_u10_n11740 ), .ZN(_u10_n14084 ) );
NAND2_X1 _u10_U2578  ( .A1(1'b0), .A2(_u10_n11716 ), .ZN(_u10_n14085 ) );
NAND4_X1 _u10_U2577  ( .A1(_u10_n14082 ), .A2(_u10_n14083 ), .A3(_u10_n14084 ), .A4(_u10_n14085 ), .ZN(_u10_n14076 ) );
NAND2_X1 _u10_U2576  ( .A1(1'b0), .A2(_u10_n11692 ), .ZN(_u10_n14078 ) );
NAND2_X1 _u10_U2575  ( .A1(1'b0), .A2(_u10_n11668 ), .ZN(_u10_n14079 ) );
NAND2_X1 _u10_U2574  ( .A1(1'b0), .A2(_u10_n11644 ), .ZN(_u10_n14080 ) );
NAND2_X1 _u10_U2573  ( .A1(1'b0), .A2(_u10_n11620 ), .ZN(_u10_n14081 ) );
NAND4_X1 _u10_U2572  ( .A1(_u10_n14078 ), .A2(_u10_n14079 ), .A3(_u10_n14080 ), .A4(_u10_n14081 ), .ZN(_u10_n14077 ) );
NOR4_X1 _u10_U2571  ( .A1(_u10_n14074 ), .A2(_u10_n14075 ), .A3(_u10_n14076 ), .A4(_u10_n14077 ), .ZN(_u10_n14073 ) );
NAND2_X1 _u10_U2570  ( .A1(_u10_n14072 ), .A2(_u10_n14073 ), .ZN(pointer_s[2]) );
NAND2_X1 _u10_U2569  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n14068 ) );
NAND2_X1 _u10_U2568  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n14069 ) );
NAND2_X1 _u10_U2567  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n14070 ) );
NAND2_X1 _u10_U2566  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n14071 ) );
NAND4_X1 _u10_U2565  ( .A1(_u10_n14068 ), .A2(_u10_n14069 ), .A3(_u10_n14070 ), .A4(_u10_n14071 ), .ZN(_u10_n14053 ) );
NAND2_X1 _u10_U2564  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n14064 ) );
NAND2_X1 _u10_U2563  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n14065 ) );
NAND2_X1 _u10_U2562  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n14066 ) );
NAND2_X1 _u10_U2561  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n14067 ) );
NAND4_X1 _u10_U2560  ( .A1(_u10_n14064 ), .A2(_u10_n14065 ), .A3(_u10_n14066 ), .A4(_u10_n14067 ), .ZN(_u10_n14054 ) );
NAND2_X1 _u10_U2559  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n14060 ) );
NAND2_X1 _u10_U2558  ( .A1(1'b0), .A2(_u10_n12137 ), .ZN(_u10_n14061 ) );
NAND2_X1 _u10_U2557  ( .A1(1'b0), .A2(_u10_n12113 ), .ZN(_u10_n14062 ) );
NAND2_X1 _u10_U2556  ( .A1(1'b0), .A2(_u10_n12089 ), .ZN(_u10_n14063 ) );
NAND4_X1 _u10_U2555  ( .A1(_u10_n14060 ), .A2(_u10_n14061 ), .A3(_u10_n14062 ), .A4(_u10_n14063 ), .ZN(_u10_n14055 ) );
NAND2_X1 _u10_U2554  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n14057 ) );
NAND2_X1 _u10_U2553  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n14058 ) );
NAND2_X1 _u10_U2552  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n14059 ) );
NAND3_X1 _u10_U2551  ( .A1(_u10_n14057 ), .A2(_u10_n14058 ), .A3(_u10_n14059 ), .ZN(_u10_n14056 ) );
NOR4_X1 _u10_U2550  ( .A1(_u10_n14053 ), .A2(_u10_n14054 ), .A3(_u10_n14055 ), .A4(_u10_n14056 ), .ZN(_u10_n14031 ) );
NAND2_X1 _u10_U2549  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n14049 ) );
NAND2_X1 _u10_U2548  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n14050 ) );
NAND2_X1 _u10_U2547  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n14051 ) );
NAND2_X1 _u10_U2546  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n14052 ) );
NAND4_X1 _u10_U2545  ( .A1(_u10_n14049 ), .A2(_u10_n14050 ), .A3(_u10_n14051 ), .A4(_u10_n14052 ), .ZN(_u10_n14033 ) );
NAND2_X1 _u10_U2544  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n14045 ) );
NAND2_X1 _u10_U2543  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n14046 ) );
NAND2_X1 _u10_U2542  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n14047 ) );
NAND2_X1 _u10_U2541  ( .A1(1'b0), .A2(_u10_n11826 ), .ZN(_u10_n14048 ) );
NAND4_X1 _u10_U2540  ( .A1(_u10_n14045 ), .A2(_u10_n14046 ), .A3(_u10_n14047 ), .A4(_u10_n14048 ), .ZN(_u10_n14034 ) );
NAND2_X1 _u10_U2539  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n14041 ) );
NAND2_X1 _u10_U2538  ( .A1(1'b0), .A2(_u10_n11780 ), .ZN(_u10_n14042 ) );
NAND2_X1 _u10_U2537  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n14043 ) );
NAND2_X1 _u10_U2536  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n14044 ) );
NAND4_X1 _u10_U2535  ( .A1(_u10_n14041 ), .A2(_u10_n14042 ), .A3(_u10_n14043 ), .A4(_u10_n14044 ), .ZN(_u10_n14035 ) );
NAND2_X1 _u10_U2534  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n14037 ) );
NAND2_X1 _u10_U2533  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n14038 ) );
NAND2_X1 _u10_U2532  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n14039 ) );
NAND2_X1 _u10_U2531  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n14040 ) );
NAND4_X1 _u10_U2530  ( .A1(_u10_n14037 ), .A2(_u10_n14038 ), .A3(_u10_n14039 ), .A4(_u10_n14040 ), .ZN(_u10_n14036 ) );
NOR4_X1 _u10_U2529  ( .A1(_u10_n14033 ), .A2(_u10_n14034 ), .A3(_u10_n14035 ), .A4(_u10_n14036 ), .ZN(_u10_n14032 ) );
NAND2_X1 _u10_U2528  ( .A1(_u10_n14031 ), .A2(_u10_n14032 ), .ZN(pointer_s[30]) );
NAND2_X1 _u10_U2527  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n14027 ) );
NAND2_X1 _u10_U2526  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n14028 ) );
NAND2_X1 _u10_U2525  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n14029 ) );
NAND2_X1 _u10_U2524  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n14030 ) );
NAND4_X1 _u10_U2523  ( .A1(_u10_n14027 ), .A2(_u10_n14028 ), .A3(_u10_n14029 ), .A4(_u10_n14030 ), .ZN(_u10_n14012 ) );
NAND2_X1 _u10_U2522  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n14023 ) );
NAND2_X1 _u10_U2521  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n14024 ) );
NAND2_X1 _u10_U2520  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n14025 ) );
NAND2_X1 _u10_U2519  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n14026 ) );
NAND4_X1 _u10_U2518  ( .A1(_u10_n14023 ), .A2(_u10_n14024 ), .A3(_u10_n14025 ), .A4(_u10_n14026 ), .ZN(_u10_n14013 ) );
NAND2_X1 _u10_U2517  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n14019 ) );
NAND2_X1 _u10_U2516  ( .A1(1'b0), .A2(_u10_n12139 ), .ZN(_u10_n14020 ) );
NAND2_X1 _u10_U2515  ( .A1(1'b0), .A2(_u10_n12115 ), .ZN(_u10_n14021 ) );
NAND2_X1 _u10_U2514  ( .A1(1'b0), .A2(_u10_n12091 ), .ZN(_u10_n14022 ) );
NAND4_X1 _u10_U2513  ( .A1(_u10_n14019 ), .A2(_u10_n14020 ), .A3(_u10_n14021 ), .A4(_u10_n14022 ), .ZN(_u10_n14014 ) );
NAND2_X1 _u10_U2512  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n14016 ) );
NAND2_X1 _u10_U2511  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n14017 ) );
NAND2_X1 _u10_U2510  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n14018 ) );
NAND3_X1 _u10_U2509  ( .A1(_u10_n14016 ), .A2(_u10_n14017 ), .A3(_u10_n14018 ), .ZN(_u10_n14015 ) );
NOR4_X1 _u10_U2508  ( .A1(_u10_n14012 ), .A2(_u10_n14013 ), .A3(_u10_n14014 ), .A4(_u10_n14015 ), .ZN(_u10_n13990 ) );
NAND2_X1 _u10_U2507  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n14008 ) );
NAND2_X1 _u10_U2506  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n14009 ) );
NAND2_X1 _u10_U2505  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n14010 ) );
NAND2_X1 _u10_U2504  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n14011 ) );
NAND4_X1 _u10_U2503  ( .A1(_u10_n14008 ), .A2(_u10_n14009 ), .A3(_u10_n14010 ), .A4(_u10_n14011 ), .ZN(_u10_n13992 ) );
NAND2_X1 _u10_U2502  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n14004 ) );
NAND2_X1 _u10_U2501  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n14005 ) );
NAND2_X1 _u10_U2500  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n14006 ) );
NAND2_X1 _u10_U2499  ( .A1(1'b0), .A2(_u10_n11831 ), .ZN(_u10_n14007 ) );
NAND4_X1 _u10_U2498  ( .A1(_u10_n14004 ), .A2(_u10_n14005 ), .A3(_u10_n14006 ), .A4(_u10_n14007 ), .ZN(_u10_n13993 ) );
NAND2_X1 _u10_U2497  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n14000 ) );
NAND2_X1 _u10_U2496  ( .A1(1'b0), .A2(_u10_n11781 ), .ZN(_u10_n14001 ) );
NAND2_X1 _u10_U2495  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n14002 ) );
NAND2_X1 _u10_U2494  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n14003 ) );
NAND4_X1 _u10_U2493  ( .A1(_u10_n14000 ), .A2(_u10_n14001 ), .A3(_u10_n14002 ), .A4(_u10_n14003 ), .ZN(_u10_n13994 ) );
NAND2_X1 _u10_U2492  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13996 ) );
NAND2_X1 _u10_U2491  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13997 ) );
NAND2_X1 _u10_U2490  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13998 ) );
NAND2_X1 _u10_U2489  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13999 ) );
NAND4_X1 _u10_U2488  ( .A1(_u10_n13996 ), .A2(_u10_n13997 ), .A3(_u10_n13998 ), .A4(_u10_n13999 ), .ZN(_u10_n13995 ) );
NOR4_X1 _u10_U2487  ( .A1(_u10_n13992 ), .A2(_u10_n13993 ), .A3(_u10_n13994 ), .A4(_u10_n13995 ), .ZN(_u10_n13991 ) );
NAND2_X1 _u10_U2486  ( .A1(_u10_n13990 ), .A2(_u10_n13991 ), .ZN(pointer_s[31]) );
NAND2_X1 _u10_U2485  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n13986 ) );
NAND2_X1 _u10_U2484  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n13987 ) );
NAND2_X1 _u10_U2483  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n13988 ) );
NAND2_X1 _u10_U2482  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n13989 ) );
NAND4_X1 _u10_U2481  ( .A1(_u10_n13986 ), .A2(_u10_n13987 ), .A3(_u10_n13988 ), .A4(_u10_n13989 ), .ZN(_u10_n13971 ) );
NAND2_X1 _u10_U2480  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n13982 ) );
NAND2_X1 _u10_U2479  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n13983 ) );
NAND2_X1 _u10_U2478  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n13984 ) );
NAND2_X1 _u10_U2477  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n13985 ) );
NAND4_X1 _u10_U2476  ( .A1(_u10_n13982 ), .A2(_u10_n13983 ), .A3(_u10_n13984 ), .A4(_u10_n13985 ), .ZN(_u10_n13972 ) );
NAND2_X1 _u10_U2475  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n13978 ) );
NAND2_X1 _u10_U2474  ( .A1(1'b0), .A2(_u10_n12138 ), .ZN(_u10_n13979 ) );
NAND2_X1 _u10_U2473  ( .A1(1'b0), .A2(_u10_n12114 ), .ZN(_u10_n13980 ) );
NAND2_X1 _u10_U2472  ( .A1(1'b0), .A2(_u10_n12090 ), .ZN(_u10_n13981 ) );
NAND4_X1 _u10_U2471  ( .A1(_u10_n13978 ), .A2(_u10_n13979 ), .A3(_u10_n13980 ), .A4(_u10_n13981 ), .ZN(_u10_n13973 ) );
NAND2_X1 _u10_U2470  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n13975 ) );
NAND2_X1 _u10_U2469  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n13976 ) );
NAND2_X1 _u10_U2468  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n13977 ) );
NAND3_X1 _u10_U2467  ( .A1(_u10_n13975 ), .A2(_u10_n13976 ), .A3(_u10_n13977 ), .ZN(_u10_n13974 ) );
NOR4_X1 _u10_U2466  ( .A1(_u10_n13971 ), .A2(_u10_n13972 ), .A3(_u10_n13973 ), .A4(_u10_n13974 ), .ZN(_u10_n13949 ) );
NAND2_X1 _u10_U2465  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n13967 ) );
NAND2_X1 _u10_U2464  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n13968 ) );
NAND2_X1 _u10_U2463  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n13969 ) );
NAND2_X1 _u10_U2462  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n13970 ) );
NAND4_X1 _u10_U2461  ( .A1(_u10_n13967 ), .A2(_u10_n13968 ), .A3(_u10_n13969 ), .A4(_u10_n13970 ), .ZN(_u10_n13951 ) );
NAND2_X1 _u10_U2460  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n13963 ) );
NAND2_X1 _u10_U2459  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n13964 ) );
NAND2_X1 _u10_U2458  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n13965 ) );
NAND2_X1 _u10_U2457  ( .A1(1'b0), .A2(_u10_n12385 ), .ZN(_u10_n13966 ) );
NAND4_X1 _u10_U2456  ( .A1(_u10_n13963 ), .A2(_u10_n13964 ), .A3(_u10_n13965 ), .A4(_u10_n13966 ), .ZN(_u10_n13952 ) );
NAND2_X1 _u10_U2455  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n13959 ) );
NAND2_X1 _u10_U2454  ( .A1(1'b0), .A2(_u10_n11778 ), .ZN(_u10_n13960 ) );
NAND2_X1 _u10_U2453  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n13961 ) );
NAND2_X1 _u10_U2452  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n13962 ) );
NAND4_X1 _u10_U2451  ( .A1(_u10_n13959 ), .A2(_u10_n13960 ), .A3(_u10_n13961 ), .A4(_u10_n13962 ), .ZN(_u10_n13953 ) );
NAND2_X1 _u10_U2450  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13955 ) );
NAND2_X1 _u10_U2449  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13956 ) );
NAND2_X1 _u10_U2448  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13957 ) );
NAND2_X1 _u10_U2447  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13958 ) );
NAND4_X1 _u10_U2446  ( .A1(_u10_n13955 ), .A2(_u10_n13956 ), .A3(_u10_n13957 ), .A4(_u10_n13958 ), .ZN(_u10_n13954 ) );
NOR4_X1 _u10_U2445  ( .A1(_u10_n13951 ), .A2(_u10_n13952 ), .A3(_u10_n13953 ), .A4(_u10_n13954 ), .ZN(_u10_n13950 ) );
NAND2_X1 _u10_U2444  ( .A1(_u10_n13949 ), .A2(_u10_n13950 ), .ZN(pointer_s[3]) );
NAND2_X1 _u10_U2443  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n13945 ) );
NAND2_X1 _u10_U2442  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n13946 ) );
NAND2_X1 _u10_U2441  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n13947 ) );
NAND2_X1 _u10_U2440  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n13948 ) );
NAND4_X1 _u10_U2439  ( .A1(_u10_n13945 ), .A2(_u10_n13946 ), .A3(_u10_n13947 ), .A4(_u10_n13948 ), .ZN(_u10_n13930 ) );
NAND2_X1 _u10_U2438  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n13941 ) );
NAND2_X1 _u10_U2437  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n13942 ) );
NAND2_X1 _u10_U2436  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n13943 ) );
NAND2_X1 _u10_U2435  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n13944 ) );
NAND4_X1 _u10_U2434  ( .A1(_u10_n13941 ), .A2(_u10_n13942 ), .A3(_u10_n13943 ), .A4(_u10_n13944 ), .ZN(_u10_n13931 ) );
NAND2_X1 _u10_U2433  ( .A1(1'b0), .A2(_u10_n12154 ), .ZN(_u10_n13937 ) );
NAND2_X1 _u10_U2432  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n13938 ) );
NAND2_X1 _u10_U2431  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n13939 ) );
NAND2_X1 _u10_U2430  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n13940 ) );
NAND4_X1 _u10_U2429  ( .A1(_u10_n13937 ), .A2(_u10_n13938 ), .A3(_u10_n13939 ), .A4(_u10_n13940 ), .ZN(_u10_n13932 ) );
NAND2_X1 _u10_U2428  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n13934 ) );
NAND2_X1 _u10_U2427  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n13935 ) );
NAND2_X1 _u10_U2426  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n13936 ) );
NAND3_X1 _u10_U2425  ( .A1(_u10_n13934 ), .A2(_u10_n13935 ), .A3(_u10_n13936 ), .ZN(_u10_n13933 ) );
NOR4_X1 _u10_U2424  ( .A1(_u10_n13930 ), .A2(_u10_n13931 ), .A3(_u10_n13932 ), .A4(_u10_n13933 ), .ZN(_u10_n13908 ) );
NAND2_X1 _u10_U2423  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n13926 ) );
NAND2_X1 _u10_U2422  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n13927 ) );
NAND2_X1 _u10_U2421  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n13928 ) );
NAND2_X1 _u10_U2420  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n13929 ) );
NAND4_X1 _u10_U2419  ( .A1(_u10_n13926 ), .A2(_u10_n13927 ), .A3(_u10_n13928 ), .A4(_u10_n13929 ), .ZN(_u10_n13910 ) );
NAND2_X1 _u10_U2418  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n13922 ) );
NAND2_X1 _u10_U2417  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n13923 ) );
NAND2_X1 _u10_U2416  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n13924 ) );
NAND2_X1 _u10_U2415  ( .A1(1'b0), .A2(_u10_n11825 ), .ZN(_u10_n13925 ) );
NAND4_X1 _u10_U2414  ( .A1(_u10_n13922 ), .A2(_u10_n13923 ), .A3(_u10_n13924 ), .A4(_u10_n13925 ), .ZN(_u10_n13911 ) );
NAND2_X1 _u10_U2413  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n13918 ) );
NAND2_X1 _u10_U2412  ( .A1(1'b0), .A2(_u10_n11779 ), .ZN(_u10_n13919 ) );
NAND2_X1 _u10_U2411  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n13920 ) );
NAND2_X1 _u10_U2410  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n13921 ) );
NAND4_X1 _u10_U2409  ( .A1(_u10_n13918 ), .A2(_u10_n13919 ), .A3(_u10_n13920 ), .A4(_u10_n13921 ), .ZN(_u10_n13912 ) );
NAND2_X1 _u10_U2408  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13914 ) );
NAND2_X1 _u10_U2407  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13915 ) );
NAND2_X1 _u10_U2406  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13916 ) );
NAND2_X1 _u10_U2405  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13917 ) );
NAND4_X1 _u10_U2404  ( .A1(_u10_n13914 ), .A2(_u10_n13915 ), .A3(_u10_n13916 ), .A4(_u10_n13917 ), .ZN(_u10_n13913 ) );
NOR4_X1 _u10_U2403  ( .A1(_u10_n13910 ), .A2(_u10_n13911 ), .A3(_u10_n13912 ), .A4(_u10_n13913 ), .ZN(_u10_n13909 ) );
NAND2_X1 _u10_U2402  ( .A1(_u10_n13908 ), .A2(_u10_n13909 ), .ZN(pointer_s[4]) );
NAND2_X1 _u10_U2401  ( .A1(1'b0), .A2(_u10_n12348 ), .ZN(_u10_n13904 ) );
NAND2_X1 _u10_U2400  ( .A1(1'b0), .A2(_u10_n12324 ), .ZN(_u10_n13905 ) );
NAND2_X1 _u10_U2399  ( .A1(1'b0), .A2(_u10_n12301 ), .ZN(_u10_n13906 ) );
NAND2_X1 _u10_U2398  ( .A1(1'b0), .A2(_u10_n12277 ), .ZN(_u10_n13907 ) );
NAND4_X1 _u10_U2397  ( .A1(_u10_n13904 ), .A2(_u10_n13905 ), .A3(_u10_n13906 ), .A4(_u10_n13907 ), .ZN(_u10_n13889 ) );
NAND2_X1 _u10_U2396  ( .A1(1'b0), .A2(_u10_n12252 ), .ZN(_u10_n13900 ) );
NAND2_X1 _u10_U2395  ( .A1(1'b0), .A2(_u10_n12228 ), .ZN(_u10_n13901 ) );
NAND2_X1 _u10_U2394  ( .A1(1'b0), .A2(_u10_n12202 ), .ZN(_u10_n13902 ) );
NAND2_X1 _u10_U2393  ( .A1(1'b0), .A2(_u10_n12180 ), .ZN(_u10_n13903 ) );
NAND4_X1 _u10_U2392  ( .A1(_u10_n13900 ), .A2(_u10_n13901 ), .A3(_u10_n13902 ), .A4(_u10_n13903 ), .ZN(_u10_n13890 ) );
NAND2_X1 _u10_U2391  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13896 ) );
NAND2_X1 _u10_U2390  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13897 ) );
NAND2_X1 _u10_U2389  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13898 ) );
NAND2_X1 _u10_U2388  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13899 ) );
NAND4_X1 _u10_U2387  ( .A1(_u10_n13896 ), .A2(_u10_n13897 ), .A3(_u10_n13898 ), .A4(_u10_n13899 ), .ZN(_u10_n13891 ) );
NAND2_X1 _u10_U2386  ( .A1(1'b0), .A2(_u10_n12058 ), .ZN(_u10_n13893 ) );
NAND2_X1 _u10_U2385  ( .A1(1'b0), .A2(_u10_n12034 ), .ZN(_u10_n13894 ) );
NAND2_X1 _u10_U2384  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n13895 ) );
NAND3_X1 _u10_U2383  ( .A1(_u10_n13893 ), .A2(_u10_n13894 ), .A3(_u10_n13895 ), .ZN(_u10_n13892 ) );
NOR4_X1 _u10_U2382  ( .A1(_u10_n13889 ), .A2(_u10_n13890 ), .A3(_u10_n13891 ), .A4(_u10_n13892 ), .ZN(_u10_n13867 ) );
NAND2_X1 _u10_U2381  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n13885 ) );
NAND2_X1 _u10_U2380  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n13886 ) );
NAND2_X1 _u10_U2379  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n13887 ) );
NAND2_X1 _u10_U2378  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n13888 ) );
NAND4_X1 _u10_U2377  ( .A1(_u10_n13885 ), .A2(_u10_n13886 ), .A3(_u10_n13887 ), .A4(_u10_n13888 ), .ZN(_u10_n13869 ) );
NAND2_X1 _u10_U2376  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n13881 ) );
NAND2_X1 _u10_U2375  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n13882 ) );
NAND2_X1 _u10_U2374  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n13883 ) );
NAND2_X1 _u10_U2373  ( .A1(1'b0), .A2(_u10_n11828 ), .ZN(_u10_n13884 ) );
NAND4_X1 _u10_U2372  ( .A1(_u10_n13881 ), .A2(_u10_n13882 ), .A3(_u10_n13883 ), .A4(_u10_n13884 ), .ZN(_u10_n13870 ) );
NAND2_X1 _u10_U2371  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n13877 ) );
NAND2_X1 _u10_U2370  ( .A1(1'b0), .A2(_u10_n11783 ), .ZN(_u10_n13878 ) );
NAND2_X1 _u10_U2369  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n13879 ) );
NAND2_X1 _u10_U2368  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n13880 ) );
NAND4_X1 _u10_U2367  ( .A1(_u10_n13877 ), .A2(_u10_n13878 ), .A3(_u10_n13879 ), .A4(_u10_n13880 ), .ZN(_u10_n13871 ) );
NAND2_X1 _u10_U2366  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13873 ) );
NAND2_X1 _u10_U2365  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13874 ) );
NAND2_X1 _u10_U2364  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13875 ) );
NAND2_X1 _u10_U2363  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13876 ) );
NAND4_X1 _u10_U2362  ( .A1(_u10_n13873 ), .A2(_u10_n13874 ), .A3(_u10_n13875 ), .A4(_u10_n13876 ), .ZN(_u10_n13872 ) );
NOR4_X1 _u10_U2361  ( .A1(_u10_n13869 ), .A2(_u10_n13870 ), .A3(_u10_n13871 ), .A4(_u10_n13872 ), .ZN(_u10_n13868 ) );
NAND2_X1 _u10_U2360  ( .A1(_u10_n13867 ), .A2(_u10_n13868 ), .ZN(pointer_s[5]) );
NAND2_X1 _u10_U2359  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13863 ) );
NAND2_X1 _u10_U2358  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13864 ) );
NAND2_X1 _u10_U2357  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13865 ) );
NAND2_X1 _u10_U2356  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13866 ) );
NAND4_X1 _u10_U2355  ( .A1(_u10_n13863 ), .A2(_u10_n13864 ), .A3(_u10_n13865 ), .A4(_u10_n13866 ), .ZN(_u10_n13848 ) );
NAND2_X1 _u10_U2354  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13859 ) );
NAND2_X1 _u10_U2353  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13860 ) );
NAND2_X1 _u10_U2352  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13861 ) );
NAND2_X1 _u10_U2351  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13862 ) );
NAND4_X1 _u10_U2350  ( .A1(_u10_n13859 ), .A2(_u10_n13860 ), .A3(_u10_n13861 ), .A4(_u10_n13862 ), .ZN(_u10_n13849 ) );
NAND2_X1 _u10_U2349  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13855 ) );
NAND2_X1 _u10_U2348  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13856 ) );
NAND2_X1 _u10_U2347  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13857 ) );
NAND2_X1 _u10_U2346  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13858 ) );
NAND4_X1 _u10_U2345  ( .A1(_u10_n13855 ), .A2(_u10_n13856 ), .A3(_u10_n13857 ), .A4(_u10_n13858 ), .ZN(_u10_n13850 ) );
NAND2_X1 _u10_U2344  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13852 ) );
NAND2_X1 _u10_U2343  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13853 ) );
NAND2_X1 _u10_U2342  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n13854 ) );
NAND3_X1 _u10_U2341  ( .A1(_u10_n13852 ), .A2(_u10_n13853 ), .A3(_u10_n13854 ), .ZN(_u10_n13851 ) );
NOR4_X1 _u10_U2340  ( .A1(_u10_n13848 ), .A2(_u10_n13849 ), .A3(_u10_n13850 ), .A4(_u10_n13851 ), .ZN(_u10_n13826 ) );
NAND2_X1 _u10_U2339  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n13844 ) );
NAND2_X1 _u10_U2338  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n13845 ) );
NAND2_X1 _u10_U2337  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n13846 ) );
NAND2_X1 _u10_U2336  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n13847 ) );
NAND4_X1 _u10_U2335  ( .A1(_u10_n13844 ), .A2(_u10_n13845 ), .A3(_u10_n13846 ), .A4(_u10_n13847 ), .ZN(_u10_n13828 ) );
NAND2_X1 _u10_U2334  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n13840 ) );
NAND2_X1 _u10_U2333  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n13841 ) );
NAND2_X1 _u10_U2332  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n13842 ) );
NAND2_X1 _u10_U2331  ( .A1(1'b0), .A2(_u10_n11829 ), .ZN(_u10_n13843 ) );
NAND4_X1 _u10_U2330  ( .A1(_u10_n13840 ), .A2(_u10_n13841 ), .A3(_u10_n13842 ), .A4(_u10_n13843 ), .ZN(_u10_n13829 ) );
NAND2_X1 _u10_U2329  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n13836 ) );
NAND2_X1 _u10_U2328  ( .A1(1'b0), .A2(_u10_n12379 ), .ZN(_u10_n13837 ) );
NAND2_X1 _u10_U2327  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n13838 ) );
NAND2_X1 _u10_U2326  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n13839 ) );
NAND4_X1 _u10_U2325  ( .A1(_u10_n13836 ), .A2(_u10_n13837 ), .A3(_u10_n13838 ), .A4(_u10_n13839 ), .ZN(_u10_n13830 ) );
NAND2_X1 _u10_U2324  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13832 ) );
NAND2_X1 _u10_U2323  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13833 ) );
NAND2_X1 _u10_U2322  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13834 ) );
NAND2_X1 _u10_U2321  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13835 ) );
NAND4_X1 _u10_U2320  ( .A1(_u10_n13832 ), .A2(_u10_n13833 ), .A3(_u10_n13834 ), .A4(_u10_n13835 ), .ZN(_u10_n13831 ) );
NOR4_X1 _u10_U2319  ( .A1(_u10_n13828 ), .A2(_u10_n13829 ), .A3(_u10_n13830 ), .A4(_u10_n13831 ), .ZN(_u10_n13827 ) );
NAND2_X1 _u10_U2318  ( .A1(_u10_n13826 ), .A2(_u10_n13827 ), .ZN(pointer_s[6]) );
NAND2_X1 _u10_U2317  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13822 ) );
NAND2_X1 _u10_U2316  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13823 ) );
NAND2_X1 _u10_U2315  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13824 ) );
NAND2_X1 _u10_U2314  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13825 ) );
NAND4_X1 _u10_U2313  ( .A1(_u10_n13822 ), .A2(_u10_n13823 ), .A3(_u10_n13824 ), .A4(_u10_n13825 ), .ZN(_u10_n13807 ) );
NAND2_X1 _u10_U2312  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13818 ) );
NAND2_X1 _u10_U2311  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13819 ) );
NAND2_X1 _u10_U2310  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13820 ) );
NAND2_X1 _u10_U2309  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13821 ) );
NAND4_X1 _u10_U2308  ( .A1(_u10_n13818 ), .A2(_u10_n13819 ), .A3(_u10_n13820 ), .A4(_u10_n13821 ), .ZN(_u10_n13808 ) );
NAND2_X1 _u10_U2307  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13814 ) );
NAND2_X1 _u10_U2306  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13815 ) );
NAND2_X1 _u10_U2305  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13816 ) );
NAND2_X1 _u10_U2304  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13817 ) );
NAND4_X1 _u10_U2303  ( .A1(_u10_n13814 ), .A2(_u10_n13815 ), .A3(_u10_n13816 ), .A4(_u10_n13817 ), .ZN(_u10_n13809 ) );
NAND2_X1 _u10_U2302  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13811 ) );
NAND2_X1 _u10_U2301  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13812 ) );
NAND2_X1 _u10_U2300  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n13813 ) );
NAND3_X1 _u10_U2299  ( .A1(_u10_n13811 ), .A2(_u10_n13812 ), .A3(_u10_n13813 ), .ZN(_u10_n13810 ) );
NOR4_X1 _u10_U2298  ( .A1(_u10_n13807 ), .A2(_u10_n13808 ), .A3(_u10_n13809 ), .A4(_u10_n13810 ), .ZN(_u10_n13785 ) );
NAND2_X1 _u10_U2297  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n13803 ) );
NAND2_X1 _u10_U2296  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n13804 ) );
NAND2_X1 _u10_U2295  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n13805 ) );
NAND2_X1 _u10_U2294  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n13806 ) );
NAND4_X1 _u10_U2293  ( .A1(_u10_n13803 ), .A2(_u10_n13804 ), .A3(_u10_n13805 ), .A4(_u10_n13806 ), .ZN(_u10_n13787 ) );
NAND2_X1 _u10_U2292  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n13799 ) );
NAND2_X1 _u10_U2291  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n13800 ) );
NAND2_X1 _u10_U2290  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n13801 ) );
NAND2_X1 _u10_U2289  ( .A1(1'b0), .A2(_u10_n11830 ), .ZN(_u10_n13802 ) );
NAND4_X1 _u10_U2288  ( .A1(_u10_n13799 ), .A2(_u10_n13800 ), .A3(_u10_n13801 ), .A4(_u10_n13802 ), .ZN(_u10_n13788 ) );
NAND2_X1 _u10_U2287  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n13795 ) );
NAND2_X1 _u10_U2286  ( .A1(1'b0), .A2(_u10_n11777 ), .ZN(_u10_n13796 ) );
NAND2_X1 _u10_U2285  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n13797 ) );
NAND2_X1 _u10_U2284  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n13798 ) );
NAND4_X1 _u10_U2283  ( .A1(_u10_n13795 ), .A2(_u10_n13796 ), .A3(_u10_n13797 ), .A4(_u10_n13798 ), .ZN(_u10_n13789 ) );
NAND2_X1 _u10_U2282  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13791 ) );
NAND2_X1 _u10_U2281  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13792 ) );
NAND2_X1 _u10_U2280  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13793 ) );
NAND2_X1 _u10_U2279  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13794 ) );
NAND4_X1 _u10_U2278  ( .A1(_u10_n13791 ), .A2(_u10_n13792 ), .A3(_u10_n13793 ), .A4(_u10_n13794 ), .ZN(_u10_n13790 ) );
NOR4_X1 _u10_U2277  ( .A1(_u10_n13787 ), .A2(_u10_n13788 ), .A3(_u10_n13789 ), .A4(_u10_n13790 ), .ZN(_u10_n13786 ) );
NAND2_X1 _u10_U2276  ( .A1(_u10_n13785 ), .A2(_u10_n13786 ), .ZN(pointer_s[7]) );
NAND2_X1 _u10_U2275  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13781 ) );
NAND2_X1 _u10_U2274  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13782 ) );
NAND2_X1 _u10_U2273  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13783 ) );
NAND2_X1 _u10_U2272  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13784 ) );
NAND4_X1 _u10_U2271  ( .A1(_u10_n13781 ), .A2(_u10_n13782 ), .A3(_u10_n13783 ), .A4(_u10_n13784 ), .ZN(_u10_n13766 ) );
NAND2_X1 _u10_U2270  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13777 ) );
NAND2_X1 _u10_U2269  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13778 ) );
NAND2_X1 _u10_U2268  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13779 ) );
NAND2_X1 _u10_U2267  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13780 ) );
NAND4_X1 _u10_U2266  ( .A1(_u10_n13777 ), .A2(_u10_n13778 ), .A3(_u10_n13779 ), .A4(_u10_n13780 ), .ZN(_u10_n13767 ) );
NAND2_X1 _u10_U2265  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13773 ) );
NAND2_X1 _u10_U2264  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13774 ) );
NAND2_X1 _u10_U2263  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13775 ) );
NAND2_X1 _u10_U2262  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13776 ) );
NAND4_X1 _u10_U2261  ( .A1(_u10_n13773 ), .A2(_u10_n13774 ), .A3(_u10_n13775 ), .A4(_u10_n13776 ), .ZN(_u10_n13768 ) );
NAND2_X1 _u10_U2260  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13770 ) );
NAND2_X1 _u10_U2259  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13771 ) );
NAND2_X1 _u10_U2258  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n13772 ) );
NAND3_X1 _u10_U2257  ( .A1(_u10_n13770 ), .A2(_u10_n13771 ), .A3(_u10_n13772 ), .ZN(_u10_n13769 ) );
NOR4_X1 _u10_U2256  ( .A1(_u10_n13766 ), .A2(_u10_n13767 ), .A3(_u10_n13768 ), .A4(_u10_n13769 ), .ZN(_u10_n13744 ) );
NAND2_X1 _u10_U2255  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n13762 ) );
NAND2_X1 _u10_U2254  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n13763 ) );
NAND2_X1 _u10_U2253  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n13764 ) );
NAND2_X1 _u10_U2252  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n13765 ) );
NAND4_X1 _u10_U2251  ( .A1(_u10_n13762 ), .A2(_u10_n13763 ), .A3(_u10_n13764 ), .A4(_u10_n13765 ), .ZN(_u10_n13746 ) );
NAND2_X1 _u10_U2250  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n13758 ) );
NAND2_X1 _u10_U2249  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n13759 ) );
NAND2_X1 _u10_U2248  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n13760 ) );
NAND2_X1 _u10_U2247  ( .A1(1'b0), .A2(_u10_n11826 ), .ZN(_u10_n13761 ) );
NAND4_X1 _u10_U2246  ( .A1(_u10_n13758 ), .A2(_u10_n13759 ), .A3(_u10_n13760 ), .A4(_u10_n13761 ), .ZN(_u10_n13747 ) );
NAND2_X1 _u10_U2245  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n13754 ) );
NAND2_X1 _u10_U2244  ( .A1(1'b0), .A2(_u10_n11782 ), .ZN(_u10_n13755 ) );
NAND2_X1 _u10_U2243  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n13756 ) );
NAND2_X1 _u10_U2242  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n13757 ) );
NAND4_X1 _u10_U2241  ( .A1(_u10_n13754 ), .A2(_u10_n13755 ), .A3(_u10_n13756 ), .A4(_u10_n13757 ), .ZN(_u10_n13748 ) );
NAND2_X1 _u10_U2240  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13750 ) );
NAND2_X1 _u10_U2239  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13751 ) );
NAND2_X1 _u10_U2238  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13752 ) );
NAND2_X1 _u10_U2237  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13753 ) );
NAND4_X1 _u10_U2236  ( .A1(_u10_n13750 ), .A2(_u10_n13751 ), .A3(_u10_n13752 ), .A4(_u10_n13753 ), .ZN(_u10_n13749 ) );
NOR4_X1 _u10_U2235  ( .A1(_u10_n13746 ), .A2(_u10_n13747 ), .A3(_u10_n13748 ), .A4(_u10_n13749 ), .ZN(_u10_n13745 ) );
NAND2_X1 _u10_U2234  ( .A1(_u10_n13744 ), .A2(_u10_n13745 ), .ZN(pointer_s[8]) );
NAND2_X1 _u10_U2233  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13740 ) );
NAND2_X1 _u10_U2232  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13741 ) );
NAND2_X1 _u10_U2231  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13742 ) );
NAND2_X1 _u10_U2230  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13743 ) );
NAND4_X1 _u10_U2229  ( .A1(_u10_n13740 ), .A2(_u10_n13741 ), .A3(_u10_n13742 ), .A4(_u10_n13743 ), .ZN(_u10_n13725 ) );
NAND2_X1 _u10_U2228  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13736 ) );
NAND2_X1 _u10_U2227  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13737 ) );
NAND2_X1 _u10_U2226  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13738 ) );
NAND2_X1 _u10_U2225  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13739 ) );
NAND4_X1 _u10_U2224  ( .A1(_u10_n13736 ), .A2(_u10_n13737 ), .A3(_u10_n13738 ), .A4(_u10_n13739 ), .ZN(_u10_n13726 ) );
NAND2_X1 _u10_U2223  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13732 ) );
NAND2_X1 _u10_U2222  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13733 ) );
NAND2_X1 _u10_U2221  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13734 ) );
NAND2_X1 _u10_U2220  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13735 ) );
NAND4_X1 _u10_U2219  ( .A1(_u10_n13732 ), .A2(_u10_n13733 ), .A3(_u10_n13734 ), .A4(_u10_n13735 ), .ZN(_u10_n13727 ) );
NAND2_X1 _u10_U2218  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13729 ) );
NAND2_X1 _u10_U2217  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13730 ) );
NAND2_X1 _u10_U2216  ( .A1(1'b0), .A2(_u10_n12017 ), .ZN(_u10_n13731 ) );
NAND3_X1 _u10_U2215  ( .A1(_u10_n13729 ), .A2(_u10_n13730 ), .A3(_u10_n13731 ), .ZN(_u10_n13728 ) );
NOR4_X1 _u10_U2214  ( .A1(_u10_n13725 ), .A2(_u10_n13726 ), .A3(_u10_n13727 ), .A4(_u10_n13728 ), .ZN(_u10_n13703 ) );
NAND2_X1 _u10_U2213  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n13721 ) );
NAND2_X1 _u10_U2212  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n13722 ) );
NAND2_X1 _u10_U2211  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n13723 ) );
NAND2_X1 _u10_U2210  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n13724 ) );
NAND4_X1 _u10_U2209  ( .A1(_u10_n13721 ), .A2(_u10_n13722 ), .A3(_u10_n13723 ), .A4(_u10_n13724 ), .ZN(_u10_n13705 ) );
NAND2_X1 _u10_U2208  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n13717 ) );
NAND2_X1 _u10_U2207  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n13718 ) );
NAND2_X1 _u10_U2206  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n13719 ) );
NAND2_X1 _u10_U2205  ( .A1(1'b0), .A2(_u10_n11827 ), .ZN(_u10_n13720 ) );
NAND4_X1 _u10_U2204  ( .A1(_u10_n13717 ), .A2(_u10_n13718 ), .A3(_u10_n13719 ), .A4(_u10_n13720 ), .ZN(_u10_n13706 ) );
NAND2_X1 _u10_U2203  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n13713 ) );
NAND2_X1 _u10_U2202  ( .A1(1'b0), .A2(_u10_n11780 ), .ZN(_u10_n13714 ) );
NAND2_X1 _u10_U2201  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n13715 ) );
NAND2_X1 _u10_U2200  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n13716 ) );
NAND4_X1 _u10_U2199  ( .A1(_u10_n13713 ), .A2(_u10_n13714 ), .A3(_u10_n13715 ), .A4(_u10_n13716 ), .ZN(_u10_n13707 ) );
NAND2_X1 _u10_U2198  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13709 ) );
NAND2_X1 _u10_U2197  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13710 ) );
NAND2_X1 _u10_U2196  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13711 ) );
NAND2_X1 _u10_U2195  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13712 ) );
NAND4_X1 _u10_U2194  ( .A1(_u10_n13709 ), .A2(_u10_n13710 ), .A3(_u10_n13711 ), .A4(_u10_n13712 ), .ZN(_u10_n13708 ) );
NOR4_X1 _u10_U2193  ( .A1(_u10_n13705 ), .A2(_u10_n13706 ), .A3(_u10_n13707 ), .A4(_u10_n13708 ), .ZN(_u10_n13704 ) );
NAND2_X1 _u10_U2192  ( .A1(_u10_n13703 ), .A2(_u10_n13704 ), .ZN(pointer_s[9]) );
NOR2_X1 _u10_U2191  ( .A1(ch0_csr[13]), .A2(_u10_n13702 ), .ZN(_u10_req_p0_0_ ) );
AND2_X1 _u10_U2190  ( .A1(_u10_n24 ), .A2(ch0_csr[13]), .ZN(_u10_req_p1_0_ ));
NAND2_X1 _u10_U2189  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13698 ) );
NAND2_X1 _u10_U2188  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13699 ) );
NAND2_X1 _u10_U2187  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13700 ) );
NAND2_X1 _u10_U2186  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13701 ) );
NAND4_X1 _u10_U2185  ( .A1(_u10_n13698 ), .A2(_u10_n13699 ), .A3(_u10_n13700 ), .A4(_u10_n13701 ), .ZN(_u10_n13683 ) );
NAND2_X1 _u10_U2184  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13694 ) );
NAND2_X1 _u10_U2183  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13695 ) );
NAND2_X1 _u10_U2182  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13696 ) );
NAND2_X1 _u10_U2181  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13697 ) );
NAND4_X1 _u10_U2180  ( .A1(_u10_n13694 ), .A2(_u10_n13695 ), .A3(_u10_n13696 ), .A4(_u10_n13697 ), .ZN(_u10_n13684 ) );
NAND2_X1 _u10_U2179  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13690 ) );
NAND2_X1 _u10_U2178  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13691 ) );
NAND2_X1 _u10_U2177  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13692 ) );
NAND2_X1 _u10_U2176  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13693 ) );
NAND4_X1 _u10_U2175  ( .A1(_u10_n13690 ), .A2(_u10_n13691 ), .A3(_u10_n13692 ), .A4(_u10_n13693 ), .ZN(_u10_n13685 ) );
NAND2_X1 _u10_U2174  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13687 ) );
NAND2_X1 _u10_U2173  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13688 ) );
NAND2_X1 _u10_U2172  ( .A1(ch0_txsz[0]), .A2(_u10_n12017 ), .ZN(_u10_n13689 ) );
NAND3_X1 _u10_U2171  ( .A1(_u10_n13687 ), .A2(_u10_n13688 ), .A3(_u10_n13689 ), .ZN(_u10_n13686 ) );
NOR4_X1 _u10_U2170  ( .A1(_u10_n13683 ), .A2(_u10_n13684 ), .A3(_u10_n13685 ), .A4(_u10_n13686 ), .ZN(_u10_n13661 ) );
NAND2_X1 _u10_U2169  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n13679 ) );
NAND2_X1 _u10_U2168  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n13680 ) );
NAND2_X1 _u10_U2167  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n13681 ) );
NAND2_X1 _u10_U2166  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n13682 ) );
NAND4_X1 _u10_U2165  ( .A1(_u10_n13679 ), .A2(_u10_n13680 ), .A3(_u10_n13681 ), .A4(_u10_n13682 ), .ZN(_u10_n13663 ) );
NAND2_X1 _u10_U2164  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n13675 ) );
NAND2_X1 _u10_U2163  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n13676 ) );
NAND2_X1 _u10_U2162  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n13677 ) );
NAND2_X1 _u10_U2161  ( .A1(1'b0), .A2(_u10_n11826 ), .ZN(_u10_n13678 ) );
NAND4_X1 _u10_U2160  ( .A1(_u10_n13675 ), .A2(_u10_n13676 ), .A3(_u10_n13677 ), .A4(_u10_n13678 ), .ZN(_u10_n13664 ) );
NAND2_X1 _u10_U2159  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n13671 ) );
NAND2_X1 _u10_U2158  ( .A1(1'b0), .A2(_u10_n11781 ), .ZN(_u10_n13672 ) );
NAND2_X1 _u10_U2157  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n13673 ) );
NAND2_X1 _u10_U2156  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n13674 ) );
NAND4_X1 _u10_U2155  ( .A1(_u10_n13671 ), .A2(_u10_n13672 ), .A3(_u10_n13673 ), .A4(_u10_n13674 ), .ZN(_u10_n13665 ) );
NAND2_X1 _u10_U2154  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13667 ) );
NAND2_X1 _u10_U2153  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13668 ) );
NAND2_X1 _u10_U2152  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13669 ) );
NAND2_X1 _u10_U2151  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13670 ) );
NAND4_X1 _u10_U2150  ( .A1(_u10_n13667 ), .A2(_u10_n13668 ), .A3(_u10_n13669 ), .A4(_u10_n13670 ), .ZN(_u10_n13666 ) );
NOR4_X1 _u10_U2149  ( .A1(_u10_n13663 ), .A2(_u10_n13664 ), .A3(_u10_n13665 ), .A4(_u10_n13666 ), .ZN(_u10_n13662 ) );
NAND2_X1 _u10_U2148  ( .A1(_u10_n13661 ), .A2(_u10_n13662 ), .ZN(txsz[0]) );
NAND2_X1 _u10_U2147  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13657 ) );
NAND2_X1 _u10_U2146  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13658 ) );
NAND2_X1 _u10_U2145  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13659 ) );
NAND2_X1 _u10_U2144  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13660 ) );
NAND4_X1 _u10_U2143  ( .A1(_u10_n13657 ), .A2(_u10_n13658 ), .A3(_u10_n13659 ), .A4(_u10_n13660 ), .ZN(_u10_n13642 ) );
NAND2_X1 _u10_U2142  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13653 ) );
NAND2_X1 _u10_U2141  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13654 ) );
NAND2_X1 _u10_U2140  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13655 ) );
NAND2_X1 _u10_U2139  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13656 ) );
NAND4_X1 _u10_U2138  ( .A1(_u10_n13653 ), .A2(_u10_n13654 ), .A3(_u10_n13655 ), .A4(_u10_n13656 ), .ZN(_u10_n13643 ) );
NAND2_X1 _u10_U2137  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13649 ) );
NAND2_X1 _u10_U2136  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13650 ) );
NAND2_X1 _u10_U2135  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13651 ) );
NAND2_X1 _u10_U2134  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13652 ) );
NAND4_X1 _u10_U2133  ( .A1(_u10_n13649 ), .A2(_u10_n13650 ), .A3(_u10_n13651 ), .A4(_u10_n13652 ), .ZN(_u10_n13644 ) );
NAND2_X1 _u10_U2132  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13646 ) );
NAND2_X1 _u10_U2131  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13647 ) );
NAND2_X1 _u10_U2130  ( .A1(ch0_txsz[10]), .A2(_u10_n12017 ), .ZN(_u10_n13648 ) );
NAND3_X1 _u10_U2129  ( .A1(_u10_n13646 ), .A2(_u10_n13647 ), .A3(_u10_n13648 ), .ZN(_u10_n13645 ) );
NOR4_X1 _u10_U2128  ( .A1(_u10_n13642 ), .A2(_u10_n13643 ), .A3(_u10_n13644 ), .A4(_u10_n13645 ), .ZN(_u10_n13620 ) );
NAND2_X1 _u10_U2127  ( .A1(1'b0), .A2(_u10_n11981 ), .ZN(_u10_n13638 ) );
NAND2_X1 _u10_U2126  ( .A1(1'b0), .A2(_u10_n11957 ), .ZN(_u10_n13639 ) );
NAND2_X1 _u10_U2125  ( .A1(1'b0), .A2(_u10_n11936 ), .ZN(_u10_n13640 ) );
NAND2_X1 _u10_U2124  ( .A1(1'b0), .A2(_u10_n11912 ), .ZN(_u10_n13641 ) );
NAND4_X1 _u10_U2123  ( .A1(_u10_n13638 ), .A2(_u10_n13639 ), .A3(_u10_n13640 ), .A4(_u10_n13641 ), .ZN(_u10_n13622 ) );
NAND2_X1 _u10_U2122  ( .A1(1'b0), .A2(_u10_n11885 ), .ZN(_u10_n13634 ) );
NAND2_X1 _u10_U2121  ( .A1(1'b0), .A2(_u10_n11861 ), .ZN(_u10_n13635 ) );
NAND2_X1 _u10_U2120  ( .A1(1'b0), .A2(_u10_n11837 ), .ZN(_u10_n13636 ) );
NAND2_X1 _u10_U2119  ( .A1(1'b0), .A2(_u10_n11831 ), .ZN(_u10_n13637 ) );
NAND4_X1 _u10_U2118  ( .A1(_u10_n13634 ), .A2(_u10_n13635 ), .A3(_u10_n13636 ), .A4(_u10_n13637 ), .ZN(_u10_n13623 ) );
NAND2_X1 _u10_U2117  ( .A1(1'b0), .A2(_u10_n11789 ), .ZN(_u10_n13630 ) );
NAND2_X1 _u10_U2116  ( .A1(1'b0), .A2(_u10_n11782 ), .ZN(_u10_n13631 ) );
NAND2_X1 _u10_U2115  ( .A1(1'b0), .A2(_u10_n11741 ), .ZN(_u10_n13632 ) );
NAND2_X1 _u10_U2114  ( .A1(1'b0), .A2(_u10_n11717 ), .ZN(_u10_n13633 ) );
NAND4_X1 _u10_U2113  ( .A1(_u10_n13630 ), .A2(_u10_n13631 ), .A3(_u10_n13632 ), .A4(_u10_n13633 ), .ZN(_u10_n13624 ) );
NAND2_X1 _u10_U2112  ( .A1(1'b0), .A2(_u10_n11693 ), .ZN(_u10_n13626 ) );
NAND2_X1 _u10_U2111  ( .A1(1'b0), .A2(_u10_n11669 ), .ZN(_u10_n13627 ) );
NAND2_X1 _u10_U2110  ( .A1(1'b0), .A2(_u10_n11645 ), .ZN(_u10_n13628 ) );
NAND2_X1 _u10_U2109  ( .A1(1'b0), .A2(_u10_n11621 ), .ZN(_u10_n13629 ) );
NAND4_X1 _u10_U2108  ( .A1(_u10_n13626 ), .A2(_u10_n13627 ), .A3(_u10_n13628 ), .A4(_u10_n13629 ), .ZN(_u10_n13625 ) );
NOR4_X1 _u10_U2107  ( .A1(_u10_n13622 ), .A2(_u10_n13623 ), .A3(_u10_n13624 ), .A4(_u10_n13625 ), .ZN(_u10_n13621 ) );
NAND2_X1 _u10_U2106  ( .A1(_u10_n13620 ), .A2(_u10_n13621 ), .ZN(txsz[10]));
NAND2_X1 _u10_U2105  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13616 ) );
NAND2_X1 _u10_U2104  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13617 ) );
NAND2_X1 _u10_U2103  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13618 ) );
NAND2_X1 _u10_U2102  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13619 ) );
NAND4_X1 _u10_U2101  ( .A1(_u10_n13616 ), .A2(_u10_n13617 ), .A3(_u10_n13618 ), .A4(_u10_n13619 ), .ZN(_u10_n13601 ) );
NAND2_X1 _u10_U2100  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13612 ) );
NAND2_X1 _u10_U2099  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13613 ) );
NAND2_X1 _u10_U2098  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13614 ) );
NAND2_X1 _u10_U2097  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13615 ) );
NAND4_X1 _u10_U2096  ( .A1(_u10_n13612 ), .A2(_u10_n13613 ), .A3(_u10_n13614 ), .A4(_u10_n13615 ), .ZN(_u10_n13602 ) );
NAND2_X1 _u10_U2095  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13608 ) );
NAND2_X1 _u10_U2094  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13609 ) );
NAND2_X1 _u10_U2093  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13610 ) );
NAND2_X1 _u10_U2092  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13611 ) );
NAND4_X1 _u10_U2091  ( .A1(_u10_n13608 ), .A2(_u10_n13609 ), .A3(_u10_n13610 ), .A4(_u10_n13611 ), .ZN(_u10_n13603 ) );
NAND2_X1 _u10_U2090  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13605 ) );
NAND2_X1 _u10_U2089  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13606 ) );
NAND2_X1 _u10_U2088  ( .A1(ch0_txsz[11]), .A2(_u10_n12017 ), .ZN(_u10_n13607 ) );
NAND3_X1 _u10_U2087  ( .A1(_u10_n13605 ), .A2(_u10_n13606 ), .A3(_u10_n13607 ), .ZN(_u10_n13604 ) );
NOR4_X1 _u10_U2086  ( .A1(_u10_n13601 ), .A2(_u10_n13602 ), .A3(_u10_n13603 ), .A4(_u10_n13604 ), .ZN(_u10_n13579 ) );
NAND2_X1 _u10_U2085  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13597 ) );
NAND2_X1 _u10_U2084  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13598 ) );
NAND2_X1 _u10_U2083  ( .A1(1'b0), .A2(_u10_n11946 ), .ZN(_u10_n13599 ) );
NAND2_X1 _u10_U2082  ( .A1(1'b0), .A2(_u10_n11922 ), .ZN(_u10_n13600 ) );
NAND4_X1 _u10_U2081  ( .A1(_u10_n13597 ), .A2(_u10_n13598 ), .A3(_u10_n13599 ), .A4(_u10_n13600 ), .ZN(_u10_n13581 ) );
NAND2_X1 _u10_U2080  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13593 ) );
NAND2_X1 _u10_U2079  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13594 ) );
NAND2_X1 _u10_U2078  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13595 ) );
NAND2_X1 _u10_U2077  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13596 ) );
NAND4_X1 _u10_U2076  ( .A1(_u10_n13593 ), .A2(_u10_n13594 ), .A3(_u10_n13595 ), .A4(_u10_n13596 ), .ZN(_u10_n13582 ) );
NAND2_X1 _u10_U2075  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13589 ) );
NAND2_X1 _u10_U2074  ( .A1(1'b0), .A2(_u10_n11782 ), .ZN(_u10_n13590 ) );
NAND2_X1 _u10_U2073  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13591 ) );
NAND2_X1 _u10_U2072  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13592 ) );
NAND4_X1 _u10_U2071  ( .A1(_u10_n13589 ), .A2(_u10_n13590 ), .A3(_u10_n13591 ), .A4(_u10_n13592 ), .ZN(_u10_n13583 ) );
NAND2_X1 _u10_U2070  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13585 ) );
NAND2_X1 _u10_U2069  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13586 ) );
NAND2_X1 _u10_U2068  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13587 ) );
NAND2_X1 _u10_U2067  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13588 ) );
NAND4_X1 _u10_U2066  ( .A1(_u10_n13585 ), .A2(_u10_n13586 ), .A3(_u10_n13587 ), .A4(_u10_n13588 ), .ZN(_u10_n13584 ) );
NOR4_X1 _u10_U2065  ( .A1(_u10_n13581 ), .A2(_u10_n13582 ), .A3(_u10_n13583 ), .A4(_u10_n13584 ), .ZN(_u10_n13580 ) );
NAND2_X1 _u10_U2064  ( .A1(_u10_n13579 ), .A2(_u10_n13580 ), .ZN(txsz[11]));
NAND2_X1 _u10_U2063  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13575 ) );
NAND2_X1 _u10_U2062  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13576 ) );
NAND2_X1 _u10_U2061  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13577 ) );
NAND2_X1 _u10_U2060  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13578 ) );
NAND4_X1 _u10_U2059  ( .A1(_u10_n13575 ), .A2(_u10_n13576 ), .A3(_u10_n13577 ), .A4(_u10_n13578 ), .ZN(_u10_n13560 ) );
NAND2_X1 _u10_U2058  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13571 ) );
NAND2_X1 _u10_U2057  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13572 ) );
NAND2_X1 _u10_U2056  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13573 ) );
NAND2_X1 _u10_U2055  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13574 ) );
NAND4_X1 _u10_U2054  ( .A1(_u10_n13571 ), .A2(_u10_n13572 ), .A3(_u10_n13573 ), .A4(_u10_n13574 ), .ZN(_u10_n13561 ) );
NAND2_X1 _u10_U2053  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13567 ) );
NAND2_X1 _u10_U2052  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13568 ) );
NAND2_X1 _u10_U2051  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13569 ) );
NAND2_X1 _u10_U2050  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13570 ) );
NAND4_X1 _u10_U2049  ( .A1(_u10_n13567 ), .A2(_u10_n13568 ), .A3(_u10_n13569 ), .A4(_u10_n13570 ), .ZN(_u10_n13562 ) );
NAND2_X1 _u10_U2048  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13564 ) );
NAND2_X1 _u10_U2047  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13565 ) );
NAND2_X1 _u10_U2046  ( .A1(1'b0), .A2(_u10_n12018 ), .ZN(_u10_n13566 ) );
NAND3_X1 _u10_U2045  ( .A1(_u10_n13564 ), .A2(_u10_n13565 ), .A3(_u10_n13566 ), .ZN(_u10_n13563 ) );
NOR4_X1 _u10_U2044  ( .A1(_u10_n13560 ), .A2(_u10_n13561 ), .A3(_u10_n13562 ), .A4(_u10_n13563 ), .ZN(_u10_n13538 ) );
NAND2_X1 _u10_U2043  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13556 ) );
NAND2_X1 _u10_U2042  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13557 ) );
NAND2_X1 _u10_U2041  ( .A1(1'b0), .A2(_u10_n11950 ), .ZN(_u10_n13558 ) );
NAND2_X1 _u10_U2040  ( .A1(1'b0), .A2(_u10_n11926 ), .ZN(_u10_n13559 ) );
NAND4_X1 _u10_U2039  ( .A1(_u10_n13556 ), .A2(_u10_n13557 ), .A3(_u10_n13558 ), .A4(_u10_n13559 ), .ZN(_u10_n13540 ) );
NAND2_X1 _u10_U2038  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13552 ) );
NAND2_X1 _u10_U2037  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13553 ) );
NAND2_X1 _u10_U2036  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13554 ) );
NAND2_X1 _u10_U2035  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13555 ) );
NAND4_X1 _u10_U2034  ( .A1(_u10_n13552 ), .A2(_u10_n13553 ), .A3(_u10_n13554 ), .A4(_u10_n13555 ), .ZN(_u10_n13541 ) );
NAND2_X1 _u10_U2033  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13548 ) );
NAND2_X1 _u10_U2032  ( .A1(1'b0), .A2(_u10_n11783 ), .ZN(_u10_n13549 ) );
NAND2_X1 _u10_U2031  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13550 ) );
NAND2_X1 _u10_U2030  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13551 ) );
NAND4_X1 _u10_U2029  ( .A1(_u10_n13548 ), .A2(_u10_n13549 ), .A3(_u10_n13550 ), .A4(_u10_n13551 ), .ZN(_u10_n13542 ) );
NAND2_X1 _u10_U2028  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13544 ) );
NAND2_X1 _u10_U2027  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13545 ) );
NAND2_X1 _u10_U2026  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13546 ) );
NAND2_X1 _u10_U2025  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13547 ) );
NAND4_X1 _u10_U2024  ( .A1(_u10_n13544 ), .A2(_u10_n13545 ), .A3(_u10_n13546 ), .A4(_u10_n13547 ), .ZN(_u10_n13543 ) );
NOR4_X1 _u10_U2023  ( .A1(_u10_n13540 ), .A2(_u10_n13541 ), .A3(_u10_n13542 ), .A4(_u10_n13543 ), .ZN(_u10_n13539 ) );
NAND2_X1 _u10_U2022  ( .A1(_u10_n13538 ), .A2(_u10_n13539 ), .ZN(txsz[12]));
NAND2_X1 _u10_U2021  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13534 ) );
NAND2_X1 _u10_U2020  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13535 ) );
NAND2_X1 _u10_U2019  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13536 ) );
NAND2_X1 _u10_U2018  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13537 ) );
NAND4_X1 _u10_U2017  ( .A1(_u10_n13534 ), .A2(_u10_n13535 ), .A3(_u10_n13536 ), .A4(_u10_n13537 ), .ZN(_u10_n13519 ) );
NAND2_X1 _u10_U2016  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13530 ) );
NAND2_X1 _u10_U2015  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13531 ) );
NAND2_X1 _u10_U2014  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13532 ) );
NAND2_X1 _u10_U2013  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13533 ) );
NAND4_X1 _u10_U2012  ( .A1(_u10_n13530 ), .A2(_u10_n13531 ), .A3(_u10_n13532 ), .A4(_u10_n13533 ), .ZN(_u10_n13520 ) );
NAND2_X1 _u10_U2011  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13526 ) );
NAND2_X1 _u10_U2010  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13527 ) );
NAND2_X1 _u10_U2009  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13528 ) );
NAND2_X1 _u10_U2008  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13529 ) );
NAND4_X1 _u10_U2007  ( .A1(_u10_n13526 ), .A2(_u10_n13527 ), .A3(_u10_n13528 ), .A4(_u10_n13529 ), .ZN(_u10_n13521 ) );
NAND2_X1 _u10_U2006  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13523 ) );
NAND2_X1 _u10_U2005  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13524 ) );
NAND2_X1 _u10_U2004  ( .A1(1'b0), .A2(_u10_n12018 ), .ZN(_u10_n13525 ) );
NAND3_X1 _u10_U2003  ( .A1(_u10_n13523 ), .A2(_u10_n13524 ), .A3(_u10_n13525 ), .ZN(_u10_n13522 ) );
NOR4_X1 _u10_U2002  ( .A1(_u10_n13519 ), .A2(_u10_n13520 ), .A3(_u10_n13521 ), .A4(_u10_n13522 ), .ZN(_u10_n13497 ) );
NAND2_X1 _u10_U2001  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13515 ) );
NAND2_X1 _u10_U2000  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13516 ) );
NAND2_X1 _u10_U1999  ( .A1(1'b0), .A2(_u10_n12394 ), .ZN(_u10_n13517 ) );
NAND2_X1 _u10_U1998  ( .A1(1'b0), .A2(_u10_n12393 ), .ZN(_u10_n13518 ) );
NAND4_X1 _u10_U1997  ( .A1(_u10_n13515 ), .A2(_u10_n13516 ), .A3(_u10_n13517 ), .A4(_u10_n13518 ), .ZN(_u10_n13499 ) );
NAND2_X1 _u10_U1996  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13511 ) );
NAND2_X1 _u10_U1995  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13512 ) );
NAND2_X1 _u10_U1994  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13513 ) );
NAND2_X1 _u10_U1993  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13514 ) );
NAND4_X1 _u10_U1992  ( .A1(_u10_n13511 ), .A2(_u10_n13512 ), .A3(_u10_n13513 ), .A4(_u10_n13514 ), .ZN(_u10_n13500 ) );
NAND2_X1 _u10_U1991  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13507 ) );
NAND2_X1 _u10_U1990  ( .A1(1'b0), .A2(_u10_n12379 ), .ZN(_u10_n13508 ) );
NAND2_X1 _u10_U1989  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13509 ) );
NAND2_X1 _u10_U1988  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13510 ) );
NAND4_X1 _u10_U1987  ( .A1(_u10_n13507 ), .A2(_u10_n13508 ), .A3(_u10_n13509 ), .A4(_u10_n13510 ), .ZN(_u10_n13501 ) );
NAND2_X1 _u10_U1986  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13503 ) );
NAND2_X1 _u10_U1985  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13504 ) );
NAND2_X1 _u10_U1984  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13505 ) );
NAND2_X1 _u10_U1983  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13506 ) );
NAND4_X1 _u10_U1982  ( .A1(_u10_n13503 ), .A2(_u10_n13504 ), .A3(_u10_n13505 ), .A4(_u10_n13506 ), .ZN(_u10_n13502 ) );
NOR4_X1 _u10_U1981  ( .A1(_u10_n13499 ), .A2(_u10_n13500 ), .A3(_u10_n13501 ), .A4(_u10_n13502 ), .ZN(_u10_n13498 ) );
NAND2_X1 _u10_U1980  ( .A1(_u10_n13497 ), .A2(_u10_n13498 ), .ZN(txsz[13]));
NAND2_X1 _u10_U1979  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13493 ) );
NAND2_X1 _u10_U1978  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13494 ) );
NAND2_X1 _u10_U1977  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13495 ) );
NAND2_X1 _u10_U1976  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13496 ) );
NAND4_X1 _u10_U1975  ( .A1(_u10_n13493 ), .A2(_u10_n13494 ), .A3(_u10_n13495 ), .A4(_u10_n13496 ), .ZN(_u10_n13478 ) );
NAND2_X1 _u10_U1974  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13489 ) );
NAND2_X1 _u10_U1973  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13490 ) );
NAND2_X1 _u10_U1972  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13491 ) );
NAND2_X1 _u10_U1971  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13492 ) );
NAND4_X1 _u10_U1970  ( .A1(_u10_n13489 ), .A2(_u10_n13490 ), .A3(_u10_n13491 ), .A4(_u10_n13492 ), .ZN(_u10_n13479 ) );
NAND2_X1 _u10_U1969  ( .A1(1'b0), .A2(_u10_n12155 ), .ZN(_u10_n13485 ) );
NAND2_X1 _u10_U1968  ( .A1(1'b0), .A2(_u10_n12131 ), .ZN(_u10_n13486 ) );
NAND2_X1 _u10_U1967  ( .A1(1'b0), .A2(_u10_n12107 ), .ZN(_u10_n13487 ) );
NAND2_X1 _u10_U1966  ( .A1(1'b0), .A2(_u10_n12083 ), .ZN(_u10_n13488 ) );
NAND4_X1 _u10_U1965  ( .A1(_u10_n13485 ), .A2(_u10_n13486 ), .A3(_u10_n13487 ), .A4(_u10_n13488 ), .ZN(_u10_n13480 ) );
NAND2_X1 _u10_U1964  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13482 ) );
NAND2_X1 _u10_U1963  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13483 ) );
NAND2_X1 _u10_U1962  ( .A1(1'b0), .A2(_u10_n12018 ), .ZN(_u10_n13484 ) );
NAND3_X1 _u10_U1961  ( .A1(_u10_n13482 ), .A2(_u10_n13483 ), .A3(_u10_n13484 ), .ZN(_u10_n13481 ) );
NOR4_X1 _u10_U1960  ( .A1(_u10_n13478 ), .A2(_u10_n13479 ), .A3(_u10_n13480 ), .A4(_u10_n13481 ), .ZN(_u10_n13456 ) );
NAND2_X1 _u10_U1959  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13474 ) );
NAND2_X1 _u10_U1958  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13475 ) );
NAND2_X1 _u10_U1957  ( .A1(1'b0), .A2(_u10_n11949 ), .ZN(_u10_n13476 ) );
NAND2_X1 _u10_U1956  ( .A1(1'b0), .A2(_u10_n11925 ), .ZN(_u10_n13477 ) );
NAND4_X1 _u10_U1955  ( .A1(_u10_n13474 ), .A2(_u10_n13475 ), .A3(_u10_n13476 ), .A4(_u10_n13477 ), .ZN(_u10_n13458 ) );
NAND2_X1 _u10_U1954  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13470 ) );
NAND2_X1 _u10_U1953  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13471 ) );
NAND2_X1 _u10_U1952  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13472 ) );
NAND2_X1 _u10_U1951  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13473 ) );
NAND4_X1 _u10_U1950  ( .A1(_u10_n13470 ), .A2(_u10_n13471 ), .A3(_u10_n13472 ), .A4(_u10_n13473 ), .ZN(_u10_n13459 ) );
NAND2_X1 _u10_U1949  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13466 ) );
NAND2_X1 _u10_U1948  ( .A1(1'b0), .A2(_u10_n11777 ), .ZN(_u10_n13467 ) );
NAND2_X1 _u10_U1947  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13468 ) );
NAND2_X1 _u10_U1946  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13469 ) );
NAND4_X1 _u10_U1945  ( .A1(_u10_n13466 ), .A2(_u10_n13467 ), .A3(_u10_n13468 ), .A4(_u10_n13469 ), .ZN(_u10_n13460 ) );
NAND2_X1 _u10_U1944  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13462 ) );
NAND2_X1 _u10_U1943  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13463 ) );
NAND2_X1 _u10_U1942  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13464 ) );
NAND2_X1 _u10_U1941  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13465 ) );
NAND4_X1 _u10_U1940  ( .A1(_u10_n13462 ), .A2(_u10_n13463 ), .A3(_u10_n13464 ), .A4(_u10_n13465 ), .ZN(_u10_n13461 ) );
NOR4_X1 _u10_U1939  ( .A1(_u10_n13458 ), .A2(_u10_n13459 ), .A3(_u10_n13460 ), .A4(_u10_n13461 ), .ZN(_u10_n13457 ) );
NAND2_X1 _u10_U1938  ( .A1(_u10_n13456 ), .A2(_u10_n13457 ), .ZN(txsz[14]));
NAND2_X1 _u10_U1937  ( .A1(1'b0), .A2(_u10_n12349 ), .ZN(_u10_n13452 ) );
NAND2_X1 _u10_U1936  ( .A1(1'b0), .A2(_u10_n12325 ), .ZN(_u10_n13453 ) );
NAND2_X1 _u10_U1935  ( .A1(1'b0), .A2(_u10_n12302 ), .ZN(_u10_n13454 ) );
NAND2_X1 _u10_U1934  ( .A1(1'b0), .A2(_u10_n12278 ), .ZN(_u10_n13455 ) );
NAND4_X1 _u10_U1933  ( .A1(_u10_n13452 ), .A2(_u10_n13453 ), .A3(_u10_n13454 ), .A4(_u10_n13455 ), .ZN(_u10_n13437 ) );
NAND2_X1 _u10_U1932  ( .A1(1'b0), .A2(_u10_n12253 ), .ZN(_u10_n13448 ) );
NAND2_X1 _u10_U1931  ( .A1(1'b0), .A2(_u10_n12229 ), .ZN(_u10_n13449 ) );
NAND2_X1 _u10_U1930  ( .A1(1'b0), .A2(_u10_n12203 ), .ZN(_u10_n13450 ) );
NAND2_X1 _u10_U1929  ( .A1(1'b0), .A2(_u10_n12181 ), .ZN(_u10_n13451 ) );
NAND4_X1 _u10_U1928  ( .A1(_u10_n13448 ), .A2(_u10_n13449 ), .A3(_u10_n13450 ), .A4(_u10_n13451 ), .ZN(_u10_n13438 ) );
NAND2_X1 _u10_U1927  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13444 ) );
NAND2_X1 _u10_U1926  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13445 ) );
NAND2_X1 _u10_U1925  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13446 ) );
NAND2_X1 _u10_U1924  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13447 ) );
NAND4_X1 _u10_U1923  ( .A1(_u10_n13444 ), .A2(_u10_n13445 ), .A3(_u10_n13446 ), .A4(_u10_n13447 ), .ZN(_u10_n13439 ) );
NAND2_X1 _u10_U1922  ( .A1(1'b0), .A2(_u10_n12059 ), .ZN(_u10_n13441 ) );
NAND2_X1 _u10_U1921  ( .A1(1'b0), .A2(_u10_n12035 ), .ZN(_u10_n13442 ) );
NAND2_X1 _u10_U1920  ( .A1(ch0_txsz[15]), .A2(_u10_n12018 ), .ZN(_u10_n13443 ) );
NAND3_X1 _u10_U1919  ( .A1(_u10_n13441 ), .A2(_u10_n13442 ), .A3(_u10_n13443 ), .ZN(_u10_n13440 ) );
NOR4_X1 _u10_U1918  ( .A1(_u10_n13437 ), .A2(_u10_n13438 ), .A3(_u10_n13439 ), .A4(_u10_n13440 ), .ZN(_u10_n13415 ) );
NAND2_X1 _u10_U1917  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13433 ) );
NAND2_X1 _u10_U1916  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13434 ) );
NAND2_X1 _u10_U1915  ( .A1(1'b0), .A2(_u10_n11945 ), .ZN(_u10_n13435 ) );
NAND2_X1 _u10_U1914  ( .A1(1'b0), .A2(_u10_n11921 ), .ZN(_u10_n13436 ) );
NAND4_X1 _u10_U1913  ( .A1(_u10_n13433 ), .A2(_u10_n13434 ), .A3(_u10_n13435 ), .A4(_u10_n13436 ), .ZN(_u10_n13417 ) );
NAND2_X1 _u10_U1912  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13429 ) );
NAND2_X1 _u10_U1911  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13430 ) );
NAND2_X1 _u10_U1910  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13431 ) );
NAND2_X1 _u10_U1909  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13432 ) );
NAND4_X1 _u10_U1908  ( .A1(_u10_n13429 ), .A2(_u10_n13430 ), .A3(_u10_n13431 ), .A4(_u10_n13432 ), .ZN(_u10_n13418 ) );
NAND2_X1 _u10_U1907  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13425 ) );
NAND2_X1 _u10_U1906  ( .A1(1'b0), .A2(_u10_n12379 ), .ZN(_u10_n13426 ) );
NAND2_X1 _u10_U1905  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13427 ) );
NAND2_X1 _u10_U1904  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13428 ) );
NAND4_X1 _u10_U1903  ( .A1(_u10_n13425 ), .A2(_u10_n13426 ), .A3(_u10_n13427 ), .A4(_u10_n13428 ), .ZN(_u10_n13419 ) );
NAND2_X1 _u10_U1902  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13421 ) );
NAND2_X1 _u10_U1901  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13422 ) );
NAND2_X1 _u10_U1900  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13423 ) );
NAND2_X1 _u10_U1899  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13424 ) );
NAND4_X1 _u10_U1898  ( .A1(_u10_n13421 ), .A2(_u10_n13422 ), .A3(_u10_n13423 ), .A4(_u10_n13424 ), .ZN(_u10_n13420 ) );
NOR4_X1 _u10_U1897  ( .A1(_u10_n13417 ), .A2(_u10_n13418 ), .A3(_u10_n13419 ), .A4(_u10_n13420 ), .ZN(_u10_n13416 ) );
NAND2_X1 _u10_U1896  ( .A1(_u10_n13415 ), .A2(_u10_n13416 ), .ZN(txsz[15]));
NAND2_X1 _u10_U1895  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13411 ) );
NAND2_X1 _u10_U1894  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13412 ) );
NAND2_X1 _u10_U1893  ( .A1(1'b0), .A2(_u10_n12428 ), .ZN(_u10_n13413 ) );
NAND2_X1 _u10_U1892  ( .A1(1'b0), .A2(_u10_n12427 ), .ZN(_u10_n13414 ) );
NAND4_X1 _u10_U1891  ( .A1(_u10_n13411 ), .A2(_u10_n13412 ), .A3(_u10_n13413 ), .A4(_u10_n13414 ), .ZN(_u10_n13396 ) );
NAND2_X1 _u10_U1890  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13407 ) );
NAND2_X1 _u10_U1889  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13408 ) );
NAND2_X1 _u10_U1888  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13409 ) );
NAND2_X1 _u10_U1887  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13410 ) );
NAND4_X1 _u10_U1886  ( .A1(_u10_n13407 ), .A2(_u10_n13408 ), .A3(_u10_n13409 ), .A4(_u10_n13410 ), .ZN(_u10_n13397 ) );
NAND2_X1 _u10_U1885  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13403 ) );
NAND2_X1 _u10_U1884  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13404 ) );
NAND2_X1 _u10_U1883  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13405 ) );
NAND2_X1 _u10_U1882  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13406 ) );
NAND4_X1 _u10_U1881  ( .A1(_u10_n13403 ), .A2(_u10_n13404 ), .A3(_u10_n13405 ), .A4(_u10_n13406 ), .ZN(_u10_n13398 ) );
NAND2_X1 _u10_U1880  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13400 ) );
NAND2_X1 _u10_U1879  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13401 ) );
NAND2_X1 _u10_U1878  ( .A1(ch0_txsz[16]), .A2(_u10_n12018 ), .ZN(_u10_n13402 ) );
NAND3_X1 _u10_U1877  ( .A1(_u10_n13400 ), .A2(_u10_n13401 ), .A3(_u10_n13402 ), .ZN(_u10_n13399 ) );
NOR4_X1 _u10_U1876  ( .A1(_u10_n13396 ), .A2(_u10_n13397 ), .A3(_u10_n13398 ), .A4(_u10_n13399 ), .ZN(_u10_n13374 ) );
NAND2_X1 _u10_U1875  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13392 ) );
NAND2_X1 _u10_U1874  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13393 ) );
NAND2_X1 _u10_U1873  ( .A1(1'b0), .A2(_u10_n11948 ), .ZN(_u10_n13394 ) );
NAND2_X1 _u10_U1872  ( .A1(1'b0), .A2(_u10_n11924 ), .ZN(_u10_n13395 ) );
NAND4_X1 _u10_U1871  ( .A1(_u10_n13392 ), .A2(_u10_n13393 ), .A3(_u10_n13394 ), .A4(_u10_n13395 ), .ZN(_u10_n13376 ) );
NAND2_X1 _u10_U1870  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13388 ) );
NAND2_X1 _u10_U1869  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13389 ) );
NAND2_X1 _u10_U1868  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13390 ) );
NAND2_X1 _u10_U1867  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13391 ) );
NAND4_X1 _u10_U1866  ( .A1(_u10_n13388 ), .A2(_u10_n13389 ), .A3(_u10_n13390 ), .A4(_u10_n13391 ), .ZN(_u10_n13377 ) );
NAND2_X1 _u10_U1865  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13384 ) );
NAND2_X1 _u10_U1864  ( .A1(1'b0), .A2(_u10_n11780 ), .ZN(_u10_n13385 ) );
NAND2_X1 _u10_U1863  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13386 ) );
NAND2_X1 _u10_U1862  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13387 ) );
NAND4_X1 _u10_U1861  ( .A1(_u10_n13384 ), .A2(_u10_n13385 ), .A3(_u10_n13386 ), .A4(_u10_n13387 ), .ZN(_u10_n13378 ) );
NAND2_X1 _u10_U1860  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13380 ) );
NAND2_X1 _u10_U1859  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13381 ) );
NAND2_X1 _u10_U1858  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13382 ) );
NAND2_X1 _u10_U1857  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13383 ) );
NAND4_X1 _u10_U1856  ( .A1(_u10_n13380 ), .A2(_u10_n13381 ), .A3(_u10_n13382 ), .A4(_u10_n13383 ), .ZN(_u10_n13379 ) );
NOR4_X1 _u10_U1855  ( .A1(_u10_n13376 ), .A2(_u10_n13377 ), .A3(_u10_n13378 ), .A4(_u10_n13379 ), .ZN(_u10_n13375 ) );
NAND2_X1 _u10_U1854  ( .A1(_u10_n13374 ), .A2(_u10_n13375 ), .ZN(txsz[16]));
NAND2_X1 _u10_U1853  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13370 ) );
NAND2_X1 _u10_U1852  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13371 ) );
NAND2_X1 _u10_U1851  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n13372 ) );
NAND2_X1 _u10_U1850  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n13373 ) );
NAND4_X1 _u10_U1849  ( .A1(_u10_n13370 ), .A2(_u10_n13371 ), .A3(_u10_n13372 ), .A4(_u10_n13373 ), .ZN(_u10_n13355 ) );
NAND2_X1 _u10_U1848  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13366 ) );
NAND2_X1 _u10_U1847  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13367 ) );
NAND2_X1 _u10_U1846  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13368 ) );
NAND2_X1 _u10_U1845  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13369 ) );
NAND4_X1 _u10_U1844  ( .A1(_u10_n13366 ), .A2(_u10_n13367 ), .A3(_u10_n13368 ), .A4(_u10_n13369 ), .ZN(_u10_n13356 ) );
NAND2_X1 _u10_U1843  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13362 ) );
NAND2_X1 _u10_U1842  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13363 ) );
NAND2_X1 _u10_U1841  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13364 ) );
NAND2_X1 _u10_U1840  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13365 ) );
NAND4_X1 _u10_U1839  ( .A1(_u10_n13362 ), .A2(_u10_n13363 ), .A3(_u10_n13364 ), .A4(_u10_n13365 ), .ZN(_u10_n13357 ) );
NAND2_X1 _u10_U1838  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13359 ) );
NAND2_X1 _u10_U1837  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13360 ) );
NAND2_X1 _u10_U1836  ( .A1(ch0_txsz[17]), .A2(_u10_n12018 ), .ZN(_u10_n13361 ) );
NAND3_X1 _u10_U1835  ( .A1(_u10_n13359 ), .A2(_u10_n13360 ), .A3(_u10_n13361 ), .ZN(_u10_n13358 ) );
NOR4_X1 _u10_U1834  ( .A1(_u10_n13355 ), .A2(_u10_n13356 ), .A3(_u10_n13357 ), .A4(_u10_n13358 ), .ZN(_u10_n13333 ) );
NAND2_X1 _u10_U1833  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13351 ) );
NAND2_X1 _u10_U1832  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13352 ) );
NAND2_X1 _u10_U1831  ( .A1(1'b0), .A2(_u10_n11948 ), .ZN(_u10_n13353 ) );
NAND2_X1 _u10_U1830  ( .A1(1'b0), .A2(_u10_n11924 ), .ZN(_u10_n13354 ) );
NAND4_X1 _u10_U1829  ( .A1(_u10_n13351 ), .A2(_u10_n13352 ), .A3(_u10_n13353 ), .A4(_u10_n13354 ), .ZN(_u10_n13335 ) );
NAND2_X1 _u10_U1828  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13347 ) );
NAND2_X1 _u10_U1827  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13348 ) );
NAND2_X1 _u10_U1826  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13349 ) );
NAND2_X1 _u10_U1825  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13350 ) );
NAND4_X1 _u10_U1824  ( .A1(_u10_n13347 ), .A2(_u10_n13348 ), .A3(_u10_n13349 ), .A4(_u10_n13350 ), .ZN(_u10_n13336 ) );
NAND2_X1 _u10_U1823  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13343 ) );
NAND2_X1 _u10_U1822  ( .A1(1'b0), .A2(_u10_n11781 ), .ZN(_u10_n13344 ) );
NAND2_X1 _u10_U1821  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13345 ) );
NAND2_X1 _u10_U1820  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13346 ) );
NAND4_X1 _u10_U1819  ( .A1(_u10_n13343 ), .A2(_u10_n13344 ), .A3(_u10_n13345 ), .A4(_u10_n13346 ), .ZN(_u10_n13337 ) );
NAND2_X1 _u10_U1818  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13339 ) );
NAND2_X1 _u10_U1817  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13340 ) );
NAND2_X1 _u10_U1816  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13341 ) );
NAND2_X1 _u10_U1815  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13342 ) );
NAND4_X1 _u10_U1814  ( .A1(_u10_n13339 ), .A2(_u10_n13340 ), .A3(_u10_n13341 ), .A4(_u10_n13342 ), .ZN(_u10_n13338 ) );
NOR4_X1 _u10_U1813  ( .A1(_u10_n13335 ), .A2(_u10_n13336 ), .A3(_u10_n13337 ), .A4(_u10_n13338 ), .ZN(_u10_n13334 ) );
NAND2_X1 _u10_U1812  ( .A1(_u10_n13333 ), .A2(_u10_n13334 ), .ZN(txsz[17]));
NAND2_X1 _u10_U1811  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13329 ) );
NAND2_X1 _u10_U1810  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13330 ) );
NAND2_X1 _u10_U1809  ( .A1(1'b0), .A2(_u10_n12305 ), .ZN(_u10_n13331 ) );
NAND2_X1 _u10_U1808  ( .A1(1'b0), .A2(_u10_n12281 ), .ZN(_u10_n13332 ) );
NAND4_X1 _u10_U1807  ( .A1(_u10_n13329 ), .A2(_u10_n13330 ), .A3(_u10_n13331 ), .A4(_u10_n13332 ), .ZN(_u10_n13314 ) );
NAND2_X1 _u10_U1806  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13325 ) );
NAND2_X1 _u10_U1805  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13326 ) );
NAND2_X1 _u10_U1804  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13327 ) );
NAND2_X1 _u10_U1803  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13328 ) );
NAND4_X1 _u10_U1802  ( .A1(_u10_n13325 ), .A2(_u10_n13326 ), .A3(_u10_n13327 ), .A4(_u10_n13328 ), .ZN(_u10_n13315 ) );
NAND2_X1 _u10_U1801  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13321 ) );
NAND2_X1 _u10_U1800  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13322 ) );
NAND2_X1 _u10_U1799  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13323 ) );
NAND2_X1 _u10_U1798  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13324 ) );
NAND4_X1 _u10_U1797  ( .A1(_u10_n13321 ), .A2(_u10_n13322 ), .A3(_u10_n13323 ), .A4(_u10_n13324 ), .ZN(_u10_n13316 ) );
NAND2_X1 _u10_U1796  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13318 ) );
NAND2_X1 _u10_U1795  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13319 ) );
NAND2_X1 _u10_U1794  ( .A1(ch0_txsz[18]), .A2(_u10_n12018 ), .ZN(_u10_n13320 ) );
NAND3_X1 _u10_U1793  ( .A1(_u10_n13318 ), .A2(_u10_n13319 ), .A3(_u10_n13320 ), .ZN(_u10_n13317 ) );
NOR4_X1 _u10_U1792  ( .A1(_u10_n13314 ), .A2(_u10_n13315 ), .A3(_u10_n13316 ), .A4(_u10_n13317 ), .ZN(_u10_n13292 ) );
NAND2_X1 _u10_U1791  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13310 ) );
NAND2_X1 _u10_U1790  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13311 ) );
NAND2_X1 _u10_U1789  ( .A1(1'b0), .A2(_u10_n11951 ), .ZN(_u10_n13312 ) );
NAND2_X1 _u10_U1788  ( .A1(1'b0), .A2(_u10_n11927 ), .ZN(_u10_n13313 ) );
NAND4_X1 _u10_U1787  ( .A1(_u10_n13310 ), .A2(_u10_n13311 ), .A3(_u10_n13312 ), .A4(_u10_n13313 ), .ZN(_u10_n13294 ) );
NAND2_X1 _u10_U1786  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13306 ) );
NAND2_X1 _u10_U1785  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13307 ) );
NAND2_X1 _u10_U1784  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13308 ) );
NAND2_X1 _u10_U1783  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13309 ) );
NAND4_X1 _u10_U1782  ( .A1(_u10_n13306 ), .A2(_u10_n13307 ), .A3(_u10_n13308 ), .A4(_u10_n13309 ), .ZN(_u10_n13295 ) );
NAND2_X1 _u10_U1781  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13302 ) );
NAND2_X1 _u10_U1780  ( .A1(1'b0), .A2(_u10_n11778 ), .ZN(_u10_n13303 ) );
NAND2_X1 _u10_U1779  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13304 ) );
NAND2_X1 _u10_U1778  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13305 ) );
NAND4_X1 _u10_U1777  ( .A1(_u10_n13302 ), .A2(_u10_n13303 ), .A3(_u10_n13304 ), .A4(_u10_n13305 ), .ZN(_u10_n13296 ) );
NAND2_X1 _u10_U1776  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13298 ) );
NAND2_X1 _u10_U1775  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13299 ) );
NAND2_X1 _u10_U1774  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13300 ) );
NAND2_X1 _u10_U1773  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13301 ) );
NAND4_X1 _u10_U1772  ( .A1(_u10_n13298 ), .A2(_u10_n13299 ), .A3(_u10_n13300 ), .A4(_u10_n13301 ), .ZN(_u10_n13297 ) );
NOR4_X1 _u10_U1771  ( .A1(_u10_n13294 ), .A2(_u10_n13295 ), .A3(_u10_n13296 ), .A4(_u10_n13297 ), .ZN(_u10_n13293 ) );
NAND2_X1 _u10_U1770  ( .A1(_u10_n13292 ), .A2(_u10_n13293 ), .ZN(txsz[18]));
NAND2_X1 _u10_U1769  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13288 ) );
NAND2_X1 _u10_U1768  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13289 ) );
NAND2_X1 _u10_U1767  ( .A1(1'b0), .A2(_u10_n12307 ), .ZN(_u10_n13290 ) );
NAND2_X1 _u10_U1766  ( .A1(1'b0), .A2(_u10_n12283 ), .ZN(_u10_n13291 ) );
NAND4_X1 _u10_U1765  ( .A1(_u10_n13288 ), .A2(_u10_n13289 ), .A3(_u10_n13290 ), .A4(_u10_n13291 ), .ZN(_u10_n13273 ) );
NAND2_X1 _u10_U1764  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13284 ) );
NAND2_X1 _u10_U1763  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13285 ) );
NAND2_X1 _u10_U1762  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13286 ) );
NAND2_X1 _u10_U1761  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13287 ) );
NAND4_X1 _u10_U1760  ( .A1(_u10_n13284 ), .A2(_u10_n13285 ), .A3(_u10_n13286 ), .A4(_u10_n13287 ), .ZN(_u10_n13274 ) );
NAND2_X1 _u10_U1759  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13280 ) );
NAND2_X1 _u10_U1758  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13281 ) );
NAND2_X1 _u10_U1757  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13282 ) );
NAND2_X1 _u10_U1756  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13283 ) );
NAND4_X1 _u10_U1755  ( .A1(_u10_n13280 ), .A2(_u10_n13281 ), .A3(_u10_n13282 ), .A4(_u10_n13283 ), .ZN(_u10_n13275 ) );
NAND2_X1 _u10_U1754  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13277 ) );
NAND2_X1 _u10_U1753  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13278 ) );
NAND2_X1 _u10_U1752  ( .A1(ch0_txsz[19]), .A2(_u10_n12018 ), .ZN(_u10_n13279 ) );
NAND3_X1 _u10_U1751  ( .A1(_u10_n13277 ), .A2(_u10_n13278 ), .A3(_u10_n13279 ), .ZN(_u10_n13276 ) );
NOR4_X1 _u10_U1750  ( .A1(_u10_n13273 ), .A2(_u10_n13274 ), .A3(_u10_n13275 ), .A4(_u10_n13276 ), .ZN(_u10_n13251 ) );
NAND2_X1 _u10_U1749  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13269 ) );
NAND2_X1 _u10_U1748  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13270 ) );
NAND2_X1 _u10_U1747  ( .A1(1'b0), .A2(_u10_n11947 ), .ZN(_u10_n13271 ) );
NAND2_X1 _u10_U1746  ( .A1(1'b0), .A2(_u10_n11923 ), .ZN(_u10_n13272 ) );
NAND4_X1 _u10_U1745  ( .A1(_u10_n13269 ), .A2(_u10_n13270 ), .A3(_u10_n13271 ), .A4(_u10_n13272 ), .ZN(_u10_n13253 ) );
NAND2_X1 _u10_U1744  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13265 ) );
NAND2_X1 _u10_U1743  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13266 ) );
NAND2_X1 _u10_U1742  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13267 ) );
NAND2_X1 _u10_U1741  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13268 ) );
NAND4_X1 _u10_U1740  ( .A1(_u10_n13265 ), .A2(_u10_n13266 ), .A3(_u10_n13267 ), .A4(_u10_n13268 ), .ZN(_u10_n13254 ) );
NAND2_X1 _u10_U1739  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13261 ) );
NAND2_X1 _u10_U1738  ( .A1(1'b0), .A2(_u10_n11779 ), .ZN(_u10_n13262 ) );
NAND2_X1 _u10_U1737  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13263 ) );
NAND2_X1 _u10_U1736  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13264 ) );
NAND4_X1 _u10_U1735  ( .A1(_u10_n13261 ), .A2(_u10_n13262 ), .A3(_u10_n13263 ), .A4(_u10_n13264 ), .ZN(_u10_n13255 ) );
NAND2_X1 _u10_U1734  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13257 ) );
NAND2_X1 _u10_U1733  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13258 ) );
NAND2_X1 _u10_U1732  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13259 ) );
NAND2_X1 _u10_U1731  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13260 ) );
NAND4_X1 _u10_U1730  ( .A1(_u10_n13257 ), .A2(_u10_n13258 ), .A3(_u10_n13259 ), .A4(_u10_n13260 ), .ZN(_u10_n13256 ) );
NOR4_X1 _u10_U1729  ( .A1(_u10_n13253 ), .A2(_u10_n13254 ), .A3(_u10_n13255 ), .A4(_u10_n13256 ), .ZN(_u10_n13252 ) );
NAND2_X1 _u10_U1728  ( .A1(_u10_n13251 ), .A2(_u10_n13252 ), .ZN(txsz[19]));
NAND2_X1 _u10_U1727  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13247 ) );
NAND2_X1 _u10_U1726  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13248 ) );
NAND2_X1 _u10_U1725  ( .A1(1'b0), .A2(_u10_n12306 ), .ZN(_u10_n13249 ) );
NAND2_X1 _u10_U1724  ( .A1(1'b0), .A2(_u10_n12282 ), .ZN(_u10_n13250 ) );
NAND4_X1 _u10_U1723  ( .A1(_u10_n13247 ), .A2(_u10_n13248 ), .A3(_u10_n13249 ), .A4(_u10_n13250 ), .ZN(_u10_n13232 ) );
NAND2_X1 _u10_U1722  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13243 ) );
NAND2_X1 _u10_U1721  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13244 ) );
NAND2_X1 _u10_U1720  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13245 ) );
NAND2_X1 _u10_U1719  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13246 ) );
NAND4_X1 _u10_U1718  ( .A1(_u10_n13243 ), .A2(_u10_n13244 ), .A3(_u10_n13245 ), .A4(_u10_n13246 ), .ZN(_u10_n13233 ) );
NAND2_X1 _u10_U1717  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13239 ) );
NAND2_X1 _u10_U1716  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13240 ) );
NAND2_X1 _u10_U1715  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13241 ) );
NAND2_X1 _u10_U1714  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13242 ) );
NAND4_X1 _u10_U1713  ( .A1(_u10_n13239 ), .A2(_u10_n13240 ), .A3(_u10_n13241 ), .A4(_u10_n13242 ), .ZN(_u10_n13234 ) );
NAND2_X1 _u10_U1712  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13236 ) );
NAND2_X1 _u10_U1711  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13237 ) );
NAND2_X1 _u10_U1710  ( .A1(ch0_txsz[1]), .A2(_u10_n12018 ), .ZN(_u10_n13238 ) );
NAND3_X1 _u10_U1709  ( .A1(_u10_n13236 ), .A2(_u10_n13237 ), .A3(_u10_n13238 ), .ZN(_u10_n13235 ) );
NOR4_X1 _u10_U1708  ( .A1(_u10_n13232 ), .A2(_u10_n13233 ), .A3(_u10_n13234 ), .A4(_u10_n13235 ), .ZN(_u10_n13210 ) );
NAND2_X1 _u10_U1707  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13228 ) );
NAND2_X1 _u10_U1706  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13229 ) );
NAND2_X1 _u10_U1705  ( .A1(1'b0), .A2(_u10_n11946 ), .ZN(_u10_n13230 ) );
NAND2_X1 _u10_U1704  ( .A1(1'b0), .A2(_u10_n11922 ), .ZN(_u10_n13231 ) );
NAND4_X1 _u10_U1703  ( .A1(_u10_n13228 ), .A2(_u10_n13229 ), .A3(_u10_n13230 ), .A4(_u10_n13231 ), .ZN(_u10_n13212 ) );
NAND2_X1 _u10_U1702  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13224 ) );
NAND2_X1 _u10_U1701  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13225 ) );
NAND2_X1 _u10_U1700  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13226 ) );
NAND2_X1 _u10_U1699  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13227 ) );
NAND4_X1 _u10_U1698  ( .A1(_u10_n13224 ), .A2(_u10_n13225 ), .A3(_u10_n13226 ), .A4(_u10_n13227 ), .ZN(_u10_n13213 ) );
NAND2_X1 _u10_U1697  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13220 ) );
NAND2_X1 _u10_U1696  ( .A1(1'b0), .A2(_u10_n11782 ), .ZN(_u10_n13221 ) );
NAND2_X1 _u10_U1695  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13222 ) );
NAND2_X1 _u10_U1694  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13223 ) );
NAND4_X1 _u10_U1693  ( .A1(_u10_n13220 ), .A2(_u10_n13221 ), .A3(_u10_n13222 ), .A4(_u10_n13223 ), .ZN(_u10_n13214 ) );
NAND2_X1 _u10_U1692  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13216 ) );
NAND2_X1 _u10_U1691  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13217 ) );
NAND2_X1 _u10_U1690  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13218 ) );
NAND2_X1 _u10_U1689  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13219 ) );
NAND4_X1 _u10_U1688  ( .A1(_u10_n13216 ), .A2(_u10_n13217 ), .A3(_u10_n13218 ), .A4(_u10_n13219 ), .ZN(_u10_n13215 ) );
NOR4_X1 _u10_U1687  ( .A1(_u10_n13212 ), .A2(_u10_n13213 ), .A3(_u10_n13214 ), .A4(_u10_n13215 ), .ZN(_u10_n13211 ) );
NAND2_X1 _u10_U1686  ( .A1(_u10_n13210 ), .A2(_u10_n13211 ), .ZN(txsz[1]) );
NAND2_X1 _u10_U1685  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13206 ) );
NAND2_X1 _u10_U1684  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13207 ) );
NAND2_X1 _u10_U1683  ( .A1(1'b0), .A2(_u10_n12305 ), .ZN(_u10_n13208 ) );
NAND2_X1 _u10_U1682  ( .A1(1'b0), .A2(_u10_n12281 ), .ZN(_u10_n13209 ) );
NAND4_X1 _u10_U1681  ( .A1(_u10_n13206 ), .A2(_u10_n13207 ), .A3(_u10_n13208 ), .A4(_u10_n13209 ), .ZN(_u10_n13191 ) );
NAND2_X1 _u10_U1680  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13202 ) );
NAND2_X1 _u10_U1679  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13203 ) );
NAND2_X1 _u10_U1678  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13204 ) );
NAND2_X1 _u10_U1677  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13205 ) );
NAND4_X1 _u10_U1676  ( .A1(_u10_n13202 ), .A2(_u10_n13203 ), .A3(_u10_n13204 ), .A4(_u10_n13205 ), .ZN(_u10_n13192 ) );
NAND2_X1 _u10_U1675  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13198 ) );
NAND2_X1 _u10_U1674  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13199 ) );
NAND2_X1 _u10_U1673  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13200 ) );
NAND2_X1 _u10_U1672  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13201 ) );
NAND4_X1 _u10_U1671  ( .A1(_u10_n13198 ), .A2(_u10_n13199 ), .A3(_u10_n13200 ), .A4(_u10_n13201 ), .ZN(_u10_n13193 ) );
NAND2_X1 _u10_U1670  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13195 ) );
NAND2_X1 _u10_U1669  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13196 ) );
NAND2_X1 _u10_U1668  ( .A1(ch0_txsz[20]), .A2(_u10_n12018 ), .ZN(_u10_n13197 ) );
NAND3_X1 _u10_U1667  ( .A1(_u10_n13195 ), .A2(_u10_n13196 ), .A3(_u10_n13197 ), .ZN(_u10_n13194 ) );
NOR4_X1 _u10_U1666  ( .A1(_u10_n13191 ), .A2(_u10_n13192 ), .A3(_u10_n13193 ), .A4(_u10_n13194 ), .ZN(_u10_n13169 ) );
NAND2_X1 _u10_U1665  ( .A1(1'b0), .A2(_u10_n11982 ), .ZN(_u10_n13187 ) );
NAND2_X1 _u10_U1664  ( .A1(1'b0), .A2(_u10_n11958 ), .ZN(_u10_n13188 ) );
NAND2_X1 _u10_U1663  ( .A1(1'b0), .A2(_u10_n11951 ), .ZN(_u10_n13189 ) );
NAND2_X1 _u10_U1662  ( .A1(1'b0), .A2(_u10_n11927 ), .ZN(_u10_n13190 ) );
NAND4_X1 _u10_U1661  ( .A1(_u10_n13187 ), .A2(_u10_n13188 ), .A3(_u10_n13189 ), .A4(_u10_n13190 ), .ZN(_u10_n13171 ) );
NAND2_X1 _u10_U1660  ( .A1(1'b0), .A2(_u10_n11886 ), .ZN(_u10_n13183 ) );
NAND2_X1 _u10_U1659  ( .A1(1'b0), .A2(_u10_n11862 ), .ZN(_u10_n13184 ) );
NAND2_X1 _u10_U1658  ( .A1(1'b0), .A2(_u10_n11838 ), .ZN(_u10_n13185 ) );
NAND2_X1 _u10_U1657  ( .A1(1'b0), .A2(_u10_n11814 ), .ZN(_u10_n13186 ) );
NAND4_X1 _u10_U1656  ( .A1(_u10_n13183 ), .A2(_u10_n13184 ), .A3(_u10_n13185 ), .A4(_u10_n13186 ), .ZN(_u10_n13172 ) );
NAND2_X1 _u10_U1655  ( .A1(1'b0), .A2(_u10_n11790 ), .ZN(_u10_n13179 ) );
NAND2_X1 _u10_U1654  ( .A1(1'b0), .A2(_u10_n11777 ), .ZN(_u10_n13180 ) );
NAND2_X1 _u10_U1653  ( .A1(1'b0), .A2(_u10_n11742 ), .ZN(_u10_n13181 ) );
NAND2_X1 _u10_U1652  ( .A1(1'b0), .A2(_u10_n11718 ), .ZN(_u10_n13182 ) );
NAND4_X1 _u10_U1651  ( .A1(_u10_n13179 ), .A2(_u10_n13180 ), .A3(_u10_n13181 ), .A4(_u10_n13182 ), .ZN(_u10_n13173 ) );
NAND2_X1 _u10_U1650  ( .A1(1'b0), .A2(_u10_n11694 ), .ZN(_u10_n13175 ) );
NAND2_X1 _u10_U1649  ( .A1(1'b0), .A2(_u10_n11670 ), .ZN(_u10_n13176 ) );
NAND2_X1 _u10_U1648  ( .A1(1'b0), .A2(_u10_n11646 ), .ZN(_u10_n13177 ) );
NAND2_X1 _u10_U1647  ( .A1(1'b0), .A2(_u10_n11622 ), .ZN(_u10_n13178 ) );
NAND4_X1 _u10_U1646  ( .A1(_u10_n13175 ), .A2(_u10_n13176 ), .A3(_u10_n13177 ), .A4(_u10_n13178 ), .ZN(_u10_n13174 ) );
NOR4_X1 _u10_U1645  ( .A1(_u10_n13171 ), .A2(_u10_n13172 ), .A3(_u10_n13173 ), .A4(_u10_n13174 ), .ZN(_u10_n13170 ) );
NAND2_X1 _u10_U1644  ( .A1(_u10_n13169 ), .A2(_u10_n13170 ), .ZN(txsz[20]));
NAND2_X1 _u10_U1643  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13165 ) );
NAND2_X1 _u10_U1642  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13166 ) );
NAND2_X1 _u10_U1641  ( .A1(1'b0), .A2(_u10_n12304 ), .ZN(_u10_n13167 ) );
NAND2_X1 _u10_U1640  ( .A1(1'b0), .A2(_u10_n12280 ), .ZN(_u10_n13168 ) );
NAND4_X1 _u10_U1639  ( .A1(_u10_n13165 ), .A2(_u10_n13166 ), .A3(_u10_n13167 ), .A4(_u10_n13168 ), .ZN(_u10_n13150 ) );
NAND2_X1 _u10_U1638  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13161 ) );
NAND2_X1 _u10_U1637  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13162 ) );
NAND2_X1 _u10_U1636  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13163 ) );
NAND2_X1 _u10_U1635  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13164 ) );
NAND4_X1 _u10_U1634  ( .A1(_u10_n13161 ), .A2(_u10_n13162 ), .A3(_u10_n13163 ), .A4(_u10_n13164 ), .ZN(_u10_n13151 ) );
NAND2_X1 _u10_U1633  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13157 ) );
NAND2_X1 _u10_U1632  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13158 ) );
NAND2_X1 _u10_U1631  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13159 ) );
NAND2_X1 _u10_U1630  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13160 ) );
NAND4_X1 _u10_U1629  ( .A1(_u10_n13157 ), .A2(_u10_n13158 ), .A3(_u10_n13159 ), .A4(_u10_n13160 ), .ZN(_u10_n13152 ) );
NAND2_X1 _u10_U1628  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13154 ) );
NAND2_X1 _u10_U1627  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13155 ) );
NAND2_X1 _u10_U1626  ( .A1(ch0_txsz[21]), .A2(_u10_n12018 ), .ZN(_u10_n13156 ) );
NAND3_X1 _u10_U1625  ( .A1(_u10_n13154 ), .A2(_u10_n13155 ), .A3(_u10_n13156 ), .ZN(_u10_n13153 ) );
NOR4_X1 _u10_U1624  ( .A1(_u10_n13150 ), .A2(_u10_n13151 ), .A3(_u10_n13152 ), .A4(_u10_n13153 ), .ZN(_u10_n13128 ) );
NAND2_X1 _u10_U1623  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n13146 ) );
NAND2_X1 _u10_U1622  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n13147 ) );
NAND2_X1 _u10_U1621  ( .A1(1'b0), .A2(_u10_n11947 ), .ZN(_u10_n13148 ) );
NAND2_X1 _u10_U1620  ( .A1(1'b0), .A2(_u10_n11923 ), .ZN(_u10_n13149 ) );
NAND4_X1 _u10_U1619  ( .A1(_u10_n13146 ), .A2(_u10_n13147 ), .A3(_u10_n13148 ), .A4(_u10_n13149 ), .ZN(_u10_n13130 ) );
NAND2_X1 _u10_U1618  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n13142 ) );
NAND2_X1 _u10_U1617  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n13143 ) );
NAND2_X1 _u10_U1616  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n13144 ) );
NAND2_X1 _u10_U1615  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n13145 ) );
NAND4_X1 _u10_U1614  ( .A1(_u10_n13142 ), .A2(_u10_n13143 ), .A3(_u10_n13144 ), .A4(_u10_n13145 ), .ZN(_u10_n13131 ) );
NAND2_X1 _u10_U1613  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n13138 ) );
NAND2_X1 _u10_U1612  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n13139 ) );
NAND2_X1 _u10_U1611  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n13140 ) );
NAND2_X1 _u10_U1610  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n13141 ) );
NAND4_X1 _u10_U1609  ( .A1(_u10_n13138 ), .A2(_u10_n13139 ), .A3(_u10_n13140 ), .A4(_u10_n13141 ), .ZN(_u10_n13132 ) );
NAND2_X1 _u10_U1608  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n13134 ) );
NAND2_X1 _u10_U1607  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n13135 ) );
NAND2_X1 _u10_U1606  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n13136 ) );
NAND2_X1 _u10_U1605  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n13137 ) );
NAND4_X1 _u10_U1604  ( .A1(_u10_n13134 ), .A2(_u10_n13135 ), .A3(_u10_n13136 ), .A4(_u10_n13137 ), .ZN(_u10_n13133 ) );
NOR4_X1 _u10_U1603  ( .A1(_u10_n13130 ), .A2(_u10_n13131 ), .A3(_u10_n13132 ), .A4(_u10_n13133 ), .ZN(_u10_n13129 ) );
NAND2_X1 _u10_U1602  ( .A1(_u10_n13128 ), .A2(_u10_n13129 ), .ZN(txsz[21]));
NAND2_X1 _u10_U1601  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13124 ) );
NAND2_X1 _u10_U1600  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13125 ) );
NAND2_X1 _u10_U1599  ( .A1(1'b0), .A2(_u10_n12303 ), .ZN(_u10_n13126 ) );
NAND2_X1 _u10_U1598  ( .A1(1'b0), .A2(_u10_n12279 ), .ZN(_u10_n13127 ) );
NAND4_X1 _u10_U1597  ( .A1(_u10_n13124 ), .A2(_u10_n13125 ), .A3(_u10_n13126 ), .A4(_u10_n13127 ), .ZN(_u10_n13109 ) );
NAND2_X1 _u10_U1596  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13120 ) );
NAND2_X1 _u10_U1595  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13121 ) );
NAND2_X1 _u10_U1594  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13122 ) );
NAND2_X1 _u10_U1593  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13123 ) );
NAND4_X1 _u10_U1592  ( .A1(_u10_n13120 ), .A2(_u10_n13121 ), .A3(_u10_n13122 ), .A4(_u10_n13123 ), .ZN(_u10_n13110 ) );
NAND2_X1 _u10_U1591  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13116 ) );
NAND2_X1 _u10_U1590  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13117 ) );
NAND2_X1 _u10_U1589  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13118 ) );
NAND2_X1 _u10_U1588  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13119 ) );
NAND4_X1 _u10_U1587  ( .A1(_u10_n13116 ), .A2(_u10_n13117 ), .A3(_u10_n13118 ), .A4(_u10_n13119 ), .ZN(_u10_n13111 ) );
NAND2_X1 _u10_U1586  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13113 ) );
NAND2_X1 _u10_U1585  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13114 ) );
NAND2_X1 _u10_U1584  ( .A1(ch0_txsz[22]), .A2(_u10_n12018 ), .ZN(_u10_n13115 ) );
NAND3_X1 _u10_U1583  ( .A1(_u10_n13113 ), .A2(_u10_n13114 ), .A3(_u10_n13115 ), .ZN(_u10_n13112 ) );
NOR4_X1 _u10_U1582  ( .A1(_u10_n13109 ), .A2(_u10_n13110 ), .A3(_u10_n13111 ), .A4(_u10_n13112 ), .ZN(_u10_n13087 ) );
NAND2_X1 _u10_U1581  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n13105 ) );
NAND2_X1 _u10_U1580  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n13106 ) );
NAND2_X1 _u10_U1579  ( .A1(1'b0), .A2(_u10_n11946 ), .ZN(_u10_n13107 ) );
NAND2_X1 _u10_U1578  ( .A1(1'b0), .A2(_u10_n11922 ), .ZN(_u10_n13108 ) );
NAND4_X1 _u10_U1577  ( .A1(_u10_n13105 ), .A2(_u10_n13106 ), .A3(_u10_n13107 ), .A4(_u10_n13108 ), .ZN(_u10_n13089 ) );
NAND2_X1 _u10_U1576  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n13101 ) );
NAND2_X1 _u10_U1575  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n13102 ) );
NAND2_X1 _u10_U1574  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n13103 ) );
NAND2_X1 _u10_U1573  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n13104 ) );
NAND4_X1 _u10_U1572  ( .A1(_u10_n13101 ), .A2(_u10_n13102 ), .A3(_u10_n13103 ), .A4(_u10_n13104 ), .ZN(_u10_n13090 ) );
NAND2_X1 _u10_U1571  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n13097 ) );
NAND2_X1 _u10_U1570  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n13098 ) );
NAND2_X1 _u10_U1569  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n13099 ) );
NAND2_X1 _u10_U1568  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n13100 ) );
NAND4_X1 _u10_U1567  ( .A1(_u10_n13097 ), .A2(_u10_n13098 ), .A3(_u10_n13099 ), .A4(_u10_n13100 ), .ZN(_u10_n13091 ) );
NAND2_X1 _u10_U1566  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n13093 ) );
NAND2_X1 _u10_U1565  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n13094 ) );
NAND2_X1 _u10_U1564  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n13095 ) );
NAND2_X1 _u10_U1563  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n13096 ) );
NAND4_X1 _u10_U1562  ( .A1(_u10_n13093 ), .A2(_u10_n13094 ), .A3(_u10_n13095 ), .A4(_u10_n13096 ), .ZN(_u10_n13092 ) );
NOR4_X1 _u10_U1561  ( .A1(_u10_n13089 ), .A2(_u10_n13090 ), .A3(_u10_n13091 ), .A4(_u10_n13092 ), .ZN(_u10_n13088 ) );
NAND2_X1 _u10_U1560  ( .A1(_u10_n13087 ), .A2(_u10_n13088 ), .ZN(txsz[22]));
NAND2_X1 _u10_U1559  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13083 ) );
NAND2_X1 _u10_U1558  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13084 ) );
NAND2_X1 _u10_U1557  ( .A1(1'b0), .A2(_u10_n12428 ), .ZN(_u10_n13085 ) );
NAND2_X1 _u10_U1556  ( .A1(1'b0), .A2(_u10_n12427 ), .ZN(_u10_n13086 ) );
NAND4_X1 _u10_U1555  ( .A1(_u10_n13083 ), .A2(_u10_n13084 ), .A3(_u10_n13085 ), .A4(_u10_n13086 ), .ZN(_u10_n13068 ) );
NAND2_X1 _u10_U1554  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13079 ) );
NAND2_X1 _u10_U1553  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13080 ) );
NAND2_X1 _u10_U1552  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13081 ) );
NAND2_X1 _u10_U1551  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13082 ) );
NAND4_X1 _u10_U1550  ( .A1(_u10_n13079 ), .A2(_u10_n13080 ), .A3(_u10_n13081 ), .A4(_u10_n13082 ), .ZN(_u10_n13069 ) );
NAND2_X1 _u10_U1549  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13075 ) );
NAND2_X1 _u10_U1548  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13076 ) );
NAND2_X1 _u10_U1547  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13077 ) );
NAND2_X1 _u10_U1546  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13078 ) );
NAND4_X1 _u10_U1545  ( .A1(_u10_n13075 ), .A2(_u10_n13076 ), .A3(_u10_n13077 ), .A4(_u10_n13078 ), .ZN(_u10_n13070 ) );
NAND2_X1 _u10_U1544  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13072 ) );
NAND2_X1 _u10_U1543  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13073 ) );
NAND2_X1 _u10_U1542  ( .A1(ch0_txsz[23]), .A2(_u10_n12019 ), .ZN(_u10_n13074 ) );
NAND3_X1 _u10_U1541  ( .A1(_u10_n13072 ), .A2(_u10_n13073 ), .A3(_u10_n13074 ), .ZN(_u10_n13071 ) );
NOR4_X1 _u10_U1540  ( .A1(_u10_n13068 ), .A2(_u10_n13069 ), .A3(_u10_n13070 ), .A4(_u10_n13071 ), .ZN(_u10_n13046 ) );
NAND2_X1 _u10_U1539  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n13064 ) );
NAND2_X1 _u10_U1538  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n13065 ) );
NAND2_X1 _u10_U1537  ( .A1(1'b0), .A2(_u10_n11950 ), .ZN(_u10_n13066 ) );
NAND2_X1 _u10_U1536  ( .A1(1'b0), .A2(_u10_n11926 ), .ZN(_u10_n13067 ) );
NAND4_X1 _u10_U1535  ( .A1(_u10_n13064 ), .A2(_u10_n13065 ), .A3(_u10_n13066 ), .A4(_u10_n13067 ), .ZN(_u10_n13048 ) );
NAND2_X1 _u10_U1534  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n13060 ) );
NAND2_X1 _u10_U1533  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n13061 ) );
NAND2_X1 _u10_U1532  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n13062 ) );
NAND2_X1 _u10_U1531  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n13063 ) );
NAND4_X1 _u10_U1530  ( .A1(_u10_n13060 ), .A2(_u10_n13061 ), .A3(_u10_n13062 ), .A4(_u10_n13063 ), .ZN(_u10_n13049 ) );
NAND2_X1 _u10_U1529  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n13056 ) );
NAND2_X1 _u10_U1528  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n13057 ) );
NAND2_X1 _u10_U1527  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n13058 ) );
NAND2_X1 _u10_U1526  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n13059 ) );
NAND4_X1 _u10_U1525  ( .A1(_u10_n13056 ), .A2(_u10_n13057 ), .A3(_u10_n13058 ), .A4(_u10_n13059 ), .ZN(_u10_n13050 ) );
NAND2_X1 _u10_U1524  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n13052 ) );
NAND2_X1 _u10_U1523  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n13053 ) );
NAND2_X1 _u10_U1522  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n13054 ) );
NAND2_X1 _u10_U1521  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n13055 ) );
NAND4_X1 _u10_U1520  ( .A1(_u10_n13052 ), .A2(_u10_n13053 ), .A3(_u10_n13054 ), .A4(_u10_n13055 ), .ZN(_u10_n13051 ) );
NOR4_X1 _u10_U1519  ( .A1(_u10_n13048 ), .A2(_u10_n13049 ), .A3(_u10_n13050 ), .A4(_u10_n13051 ), .ZN(_u10_n13047 ) );
NAND2_X1 _u10_U1518  ( .A1(_u10_n13046 ), .A2(_u10_n13047 ), .ZN(txsz[23]));
NAND2_X1 _u10_U1517  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13042 ) );
NAND2_X1 _u10_U1516  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13043 ) );
NAND2_X1 _u10_U1515  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n13044 ) );
NAND2_X1 _u10_U1514  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n13045 ) );
NAND4_X1 _u10_U1513  ( .A1(_u10_n13042 ), .A2(_u10_n13043 ), .A3(_u10_n13044 ), .A4(_u10_n13045 ), .ZN(_u10_n13027 ) );
NAND2_X1 _u10_U1512  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n13038 ) );
NAND2_X1 _u10_U1511  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n13039 ) );
NAND2_X1 _u10_U1510  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n13040 ) );
NAND2_X1 _u10_U1509  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13041 ) );
NAND4_X1 _u10_U1508  ( .A1(_u10_n13038 ), .A2(_u10_n13039 ), .A3(_u10_n13040 ), .A4(_u10_n13041 ), .ZN(_u10_n13028 ) );
NAND2_X1 _u10_U1507  ( .A1(1'b0), .A2(_u10_n12156 ), .ZN(_u10_n13034 ) );
NAND2_X1 _u10_U1506  ( .A1(1'b0), .A2(_u10_n12132 ), .ZN(_u10_n13035 ) );
NAND2_X1 _u10_U1505  ( .A1(1'b0), .A2(_u10_n12108 ), .ZN(_u10_n13036 ) );
NAND2_X1 _u10_U1504  ( .A1(1'b0), .A2(_u10_n12084 ), .ZN(_u10_n13037 ) );
NAND4_X1 _u10_U1503  ( .A1(_u10_n13034 ), .A2(_u10_n13035 ), .A3(_u10_n13036 ), .A4(_u10_n13037 ), .ZN(_u10_n13029 ) );
NAND2_X1 _u10_U1502  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n13031 ) );
NAND2_X1 _u10_U1501  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n13032 ) );
NAND2_X1 _u10_U1500  ( .A1(ch0_txsz[24]), .A2(_u10_n12019 ), .ZN(_u10_n13033 ) );
NAND3_X1 _u10_U1499  ( .A1(_u10_n13031 ), .A2(_u10_n13032 ), .A3(_u10_n13033 ), .ZN(_u10_n13030 ) );
NOR4_X1 _u10_U1498  ( .A1(_u10_n13027 ), .A2(_u10_n13028 ), .A3(_u10_n13029 ), .A4(_u10_n13030 ), .ZN(_u10_n13005 ) );
NAND2_X1 _u10_U1497  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n13023 ) );
NAND2_X1 _u10_U1496  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n13024 ) );
NAND2_X1 _u10_U1495  ( .A1(1'b0), .A2(_u10_n12394 ), .ZN(_u10_n13025 ) );
NAND2_X1 _u10_U1494  ( .A1(1'b0), .A2(_u10_n12393 ), .ZN(_u10_n13026 ) );
NAND4_X1 _u10_U1493  ( .A1(_u10_n13023 ), .A2(_u10_n13024 ), .A3(_u10_n13025 ), .A4(_u10_n13026 ), .ZN(_u10_n13007 ) );
NAND2_X1 _u10_U1492  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n13019 ) );
NAND2_X1 _u10_U1491  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n13020 ) );
NAND2_X1 _u10_U1490  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n13021 ) );
NAND2_X1 _u10_U1489  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n13022 ) );
NAND4_X1 _u10_U1488  ( .A1(_u10_n13019 ), .A2(_u10_n13020 ), .A3(_u10_n13021 ), .A4(_u10_n13022 ), .ZN(_u10_n13008 ) );
NAND2_X1 _u10_U1487  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n13015 ) );
NAND2_X1 _u10_U1486  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n13016 ) );
NAND2_X1 _u10_U1485  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n13017 ) );
NAND2_X1 _u10_U1484  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n13018 ) );
NAND4_X1 _u10_U1483  ( .A1(_u10_n13015 ), .A2(_u10_n13016 ), .A3(_u10_n13017 ), .A4(_u10_n13018 ), .ZN(_u10_n13009 ) );
NAND2_X1 _u10_U1482  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n13011 ) );
NAND2_X1 _u10_U1481  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n13012 ) );
NAND2_X1 _u10_U1480  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n13013 ) );
NAND2_X1 _u10_U1479  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n13014 ) );
NAND4_X1 _u10_U1478  ( .A1(_u10_n13011 ), .A2(_u10_n13012 ), .A3(_u10_n13013 ), .A4(_u10_n13014 ), .ZN(_u10_n13010 ) );
NOR4_X1 _u10_U1477  ( .A1(_u10_n13007 ), .A2(_u10_n13008 ), .A3(_u10_n13009 ), .A4(_u10_n13010 ), .ZN(_u10_n13006 ) );
NAND2_X1 _u10_U1476  ( .A1(_u10_n13005 ), .A2(_u10_n13006 ), .ZN(txsz[24]));
NAND2_X1 _u10_U1475  ( .A1(1'b0), .A2(_u10_n12350 ), .ZN(_u10_n13001 ) );
NAND2_X1 _u10_U1474  ( .A1(1'b0), .A2(_u10_n12326 ), .ZN(_u10_n13002 ) );
NAND2_X1 _u10_U1473  ( .A1(1'b0), .A2(_u10_n12303 ), .ZN(_u10_n13003 ) );
NAND2_X1 _u10_U1472  ( .A1(1'b0), .A2(_u10_n12279 ), .ZN(_u10_n13004 ) );
NAND4_X1 _u10_U1471  ( .A1(_u10_n13001 ), .A2(_u10_n13002 ), .A3(_u10_n13003 ), .A4(_u10_n13004 ), .ZN(_u10_n12986 ) );
NAND2_X1 _u10_U1470  ( .A1(1'b0), .A2(_u10_n12254 ), .ZN(_u10_n12997 ) );
NAND2_X1 _u10_U1469  ( .A1(1'b0), .A2(_u10_n12230 ), .ZN(_u10_n12998 ) );
NAND2_X1 _u10_U1468  ( .A1(1'b0), .A2(_u10_n12204 ), .ZN(_u10_n12999 ) );
NAND2_X1 _u10_U1467  ( .A1(1'b0), .A2(_u10_n12182 ), .ZN(_u10_n13000 ) );
NAND4_X1 _u10_U1466  ( .A1(_u10_n12997 ), .A2(_u10_n12998 ), .A3(_u10_n12999 ), .A4(_u10_n13000 ), .ZN(_u10_n12987 ) );
NAND2_X1 _u10_U1465  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12993 ) );
NAND2_X1 _u10_U1464  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12994 ) );
NAND2_X1 _u10_U1463  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12995 ) );
NAND2_X1 _u10_U1462  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12996 ) );
NAND4_X1 _u10_U1461  ( .A1(_u10_n12993 ), .A2(_u10_n12994 ), .A3(_u10_n12995 ), .A4(_u10_n12996 ), .ZN(_u10_n12988 ) );
NAND2_X1 _u10_U1460  ( .A1(1'b0), .A2(_u10_n12060 ), .ZN(_u10_n12990 ) );
NAND2_X1 _u10_U1459  ( .A1(1'b0), .A2(_u10_n12036 ), .ZN(_u10_n12991 ) );
NAND2_X1 _u10_U1458  ( .A1(ch0_txsz[25]), .A2(_u10_n12019 ), .ZN(_u10_n12992 ) );
NAND3_X1 _u10_U1457  ( .A1(_u10_n12990 ), .A2(_u10_n12991 ), .A3(_u10_n12992 ), .ZN(_u10_n12989 ) );
NOR4_X1 _u10_U1456  ( .A1(_u10_n12986 ), .A2(_u10_n12987 ), .A3(_u10_n12988 ), .A4(_u10_n12989 ), .ZN(_u10_n12964 ) );
NAND2_X1 _u10_U1455  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n12982 ) );
NAND2_X1 _u10_U1454  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n12983 ) );
NAND2_X1 _u10_U1453  ( .A1(1'b0), .A2(_u10_n11949 ), .ZN(_u10_n12984 ) );
NAND2_X1 _u10_U1452  ( .A1(1'b0), .A2(_u10_n11925 ), .ZN(_u10_n12985 ) );
NAND4_X1 _u10_U1451  ( .A1(_u10_n12982 ), .A2(_u10_n12983 ), .A3(_u10_n12984 ), .A4(_u10_n12985 ), .ZN(_u10_n12966 ) );
NAND2_X1 _u10_U1450  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n12978 ) );
NAND2_X1 _u10_U1449  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n12979 ) );
NAND2_X1 _u10_U1448  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n12980 ) );
NAND2_X1 _u10_U1447  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n12981 ) );
NAND4_X1 _u10_U1446  ( .A1(_u10_n12978 ), .A2(_u10_n12979 ), .A3(_u10_n12980 ), .A4(_u10_n12981 ), .ZN(_u10_n12967 ) );
NAND2_X1 _u10_U1445  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n12974 ) );
NAND2_X1 _u10_U1444  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n12975 ) );
NAND2_X1 _u10_U1443  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n12976 ) );
NAND2_X1 _u10_U1442  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n12977 ) );
NAND4_X1 _u10_U1441  ( .A1(_u10_n12974 ), .A2(_u10_n12975 ), .A3(_u10_n12976 ), .A4(_u10_n12977 ), .ZN(_u10_n12968 ) );
NAND2_X1 _u10_U1440  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n12970 ) );
NAND2_X1 _u10_U1439  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n12971 ) );
NAND2_X1 _u10_U1438  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n12972 ) );
NAND2_X1 _u10_U1437  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n12973 ) );
NAND4_X1 _u10_U1436  ( .A1(_u10_n12970 ), .A2(_u10_n12971 ), .A3(_u10_n12972 ), .A4(_u10_n12973 ), .ZN(_u10_n12969 ) );
NOR4_X1 _u10_U1435  ( .A1(_u10_n12966 ), .A2(_u10_n12967 ), .A3(_u10_n12968 ), .A4(_u10_n12969 ), .ZN(_u10_n12965 ) );
NAND2_X1 _u10_U1434  ( .A1(_u10_n12964 ), .A2(_u10_n12965 ), .ZN(txsz[25]));
NAND2_X1 _u10_U1433  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12960 ) );
NAND2_X1 _u10_U1432  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12961 ) );
NAND2_X1 _u10_U1431  ( .A1(1'b0), .A2(_u10_n12305 ), .ZN(_u10_n12962 ) );
NAND2_X1 _u10_U1430  ( .A1(1'b0), .A2(_u10_n12281 ), .ZN(_u10_n12963 ) );
NAND4_X1 _u10_U1429  ( .A1(_u10_n12960 ), .A2(_u10_n12961 ), .A3(_u10_n12962 ), .A4(_u10_n12963 ), .ZN(_u10_n12945 ) );
NAND2_X1 _u10_U1428  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12956 ) );
NAND2_X1 _u10_U1427  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12957 ) );
NAND2_X1 _u10_U1426  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12958 ) );
NAND2_X1 _u10_U1425  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12959 ) );
NAND4_X1 _u10_U1424  ( .A1(_u10_n12956 ), .A2(_u10_n12957 ), .A3(_u10_n12958 ), .A4(_u10_n12959 ), .ZN(_u10_n12946 ) );
NAND2_X1 _u10_U1423  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12952 ) );
NAND2_X1 _u10_U1422  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12953 ) );
NAND2_X1 _u10_U1421  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12954 ) );
NAND2_X1 _u10_U1420  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12955 ) );
NAND4_X1 _u10_U1419  ( .A1(_u10_n12952 ), .A2(_u10_n12953 ), .A3(_u10_n12954 ), .A4(_u10_n12955 ), .ZN(_u10_n12947 ) );
NAND2_X1 _u10_U1418  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12949 ) );
NAND2_X1 _u10_U1417  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12950 ) );
NAND2_X1 _u10_U1416  ( .A1(ch0_txsz[26]), .A2(_u10_n12019 ), .ZN(_u10_n12951 ) );
NAND3_X1 _u10_U1415  ( .A1(_u10_n12949 ), .A2(_u10_n12950 ), .A3(_u10_n12951 ), .ZN(_u10_n12948 ) );
NOR4_X1 _u10_U1414  ( .A1(_u10_n12945 ), .A2(_u10_n12946 ), .A3(_u10_n12947 ), .A4(_u10_n12948 ), .ZN(_u10_n12923 ) );
NAND2_X1 _u10_U1413  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n12941 ) );
NAND2_X1 _u10_U1412  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n12942 ) );
NAND2_X1 _u10_U1411  ( .A1(1'b0), .A2(_u10_n11945 ), .ZN(_u10_n12943 ) );
NAND2_X1 _u10_U1410  ( .A1(1'b0), .A2(_u10_n11921 ), .ZN(_u10_n12944 ) );
NAND4_X1 _u10_U1409  ( .A1(_u10_n12941 ), .A2(_u10_n12942 ), .A3(_u10_n12943 ), .A4(_u10_n12944 ), .ZN(_u10_n12925 ) );
NAND2_X1 _u10_U1408  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n12937 ) );
NAND2_X1 _u10_U1407  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n12938 ) );
NAND2_X1 _u10_U1406  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n12939 ) );
NAND2_X1 _u10_U1405  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n12940 ) );
NAND4_X1 _u10_U1404  ( .A1(_u10_n12937 ), .A2(_u10_n12938 ), .A3(_u10_n12939 ), .A4(_u10_n12940 ), .ZN(_u10_n12926 ) );
NAND2_X1 _u10_U1403  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n12933 ) );
NAND2_X1 _u10_U1402  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n12934 ) );
NAND2_X1 _u10_U1401  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n12935 ) );
NAND2_X1 _u10_U1400  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n12936 ) );
NAND4_X1 _u10_U1399  ( .A1(_u10_n12933 ), .A2(_u10_n12934 ), .A3(_u10_n12935 ), .A4(_u10_n12936 ), .ZN(_u10_n12927 ) );
NAND2_X1 _u10_U1398  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n12929 ) );
NAND2_X1 _u10_U1397  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n12930 ) );
NAND2_X1 _u10_U1396  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n12931 ) );
NAND2_X1 _u10_U1395  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n12932 ) );
NAND4_X1 _u10_U1394  ( .A1(_u10_n12929 ), .A2(_u10_n12930 ), .A3(_u10_n12931 ), .A4(_u10_n12932 ), .ZN(_u10_n12928 ) );
NOR4_X1 _u10_U1393  ( .A1(_u10_n12925 ), .A2(_u10_n12926 ), .A3(_u10_n12927 ), .A4(_u10_n12928 ), .ZN(_u10_n12924 ) );
NAND2_X1 _u10_U1392  ( .A1(_u10_n12923 ), .A2(_u10_n12924 ), .ZN(txsz[26]));
NAND2_X1 _u10_U1391  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12919 ) );
NAND2_X1 _u10_U1390  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12920 ) );
NAND2_X1 _u10_U1389  ( .A1(1'b0), .A2(_u10_n12303 ), .ZN(_u10_n12921 ) );
NAND2_X1 _u10_U1388  ( .A1(1'b0), .A2(_u10_n12279 ), .ZN(_u10_n12922 ) );
NAND4_X1 _u10_U1387  ( .A1(_u10_n12919 ), .A2(_u10_n12920 ), .A3(_u10_n12921 ), .A4(_u10_n12922 ), .ZN(_u10_n12904 ) );
NAND2_X1 _u10_U1386  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12915 ) );
NAND2_X1 _u10_U1385  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12916 ) );
NAND2_X1 _u10_U1384  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12917 ) );
NAND2_X1 _u10_U1383  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12918 ) );
NAND4_X1 _u10_U1382  ( .A1(_u10_n12915 ), .A2(_u10_n12916 ), .A3(_u10_n12917 ), .A4(_u10_n12918 ), .ZN(_u10_n12905 ) );
NAND2_X1 _u10_U1381  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12911 ) );
NAND2_X1 _u10_U1380  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12912 ) );
NAND2_X1 _u10_U1379  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12913 ) );
NAND2_X1 _u10_U1378  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12914 ) );
NAND4_X1 _u10_U1377  ( .A1(_u10_n12911 ), .A2(_u10_n12912 ), .A3(_u10_n12913 ), .A4(_u10_n12914 ), .ZN(_u10_n12906 ) );
NAND2_X1 _u10_U1376  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12908 ) );
NAND2_X1 _u10_U1375  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12909 ) );
NAND2_X1 _u10_U1374  ( .A1(1'b0), .A2(_u10_n12019 ), .ZN(_u10_n12910 ) );
NAND3_X1 _u10_U1373  ( .A1(_u10_n12908 ), .A2(_u10_n12909 ), .A3(_u10_n12910 ), .ZN(_u10_n12907 ) );
NOR4_X1 _u10_U1372  ( .A1(_u10_n12904 ), .A2(_u10_n12905 ), .A3(_u10_n12906 ), .A4(_u10_n12907 ), .ZN(_u10_n12882 ) );
NAND2_X1 _u10_U1371  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n12900 ) );
NAND2_X1 _u10_U1370  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n12901 ) );
NAND2_X1 _u10_U1369  ( .A1(1'b0), .A2(_u10_n11947 ), .ZN(_u10_n12902 ) );
NAND2_X1 _u10_U1368  ( .A1(1'b0), .A2(_u10_n11923 ), .ZN(_u10_n12903 ) );
NAND4_X1 _u10_U1367  ( .A1(_u10_n12900 ), .A2(_u10_n12901 ), .A3(_u10_n12902 ), .A4(_u10_n12903 ), .ZN(_u10_n12884 ) );
NAND2_X1 _u10_U1366  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n12896 ) );
NAND2_X1 _u10_U1365  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n12897 ) );
NAND2_X1 _u10_U1364  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n12898 ) );
NAND2_X1 _u10_U1363  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n12899 ) );
NAND4_X1 _u10_U1362  ( .A1(_u10_n12896 ), .A2(_u10_n12897 ), .A3(_u10_n12898 ), .A4(_u10_n12899 ), .ZN(_u10_n12885 ) );
NAND2_X1 _u10_U1361  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n12892 ) );
NAND2_X1 _u10_U1360  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n12893 ) );
NAND2_X1 _u10_U1359  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n12894 ) );
NAND2_X1 _u10_U1358  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n12895 ) );
NAND4_X1 _u10_U1357  ( .A1(_u10_n12892 ), .A2(_u10_n12893 ), .A3(_u10_n12894 ), .A4(_u10_n12895 ), .ZN(_u10_n12886 ) );
NAND2_X1 _u10_U1356  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n12888 ) );
NAND2_X1 _u10_U1355  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n12889 ) );
NAND2_X1 _u10_U1354  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n12890 ) );
NAND2_X1 _u10_U1353  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n12891 ) );
NAND4_X1 _u10_U1352  ( .A1(_u10_n12888 ), .A2(_u10_n12889 ), .A3(_u10_n12890 ), .A4(_u10_n12891 ), .ZN(_u10_n12887 ) );
NOR4_X1 _u10_U1351  ( .A1(_u10_n12884 ), .A2(_u10_n12885 ), .A3(_u10_n12886 ), .A4(_u10_n12887 ), .ZN(_u10_n12883 ) );
NAND2_X1 _u10_U1350  ( .A1(_u10_n12882 ), .A2(_u10_n12883 ), .ZN(txsz[27]));
NAND2_X1 _u10_U1349  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12878 ) );
NAND2_X1 _u10_U1348  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12879 ) );
NAND2_X1 _u10_U1347  ( .A1(1'b0), .A2(_u10_n12428 ), .ZN(_u10_n12880 ) );
NAND2_X1 _u10_U1346  ( .A1(1'b0), .A2(_u10_n12427 ), .ZN(_u10_n12881 ) );
NAND4_X1 _u10_U1345  ( .A1(_u10_n12878 ), .A2(_u10_n12879 ), .A3(_u10_n12880 ), .A4(_u10_n12881 ), .ZN(_u10_n12863 ) );
NAND2_X1 _u10_U1344  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12874 ) );
NAND2_X1 _u10_U1343  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12875 ) );
NAND2_X1 _u10_U1342  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12876 ) );
NAND2_X1 _u10_U1341  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12877 ) );
NAND4_X1 _u10_U1340  ( .A1(_u10_n12874 ), .A2(_u10_n12875 ), .A3(_u10_n12876 ), .A4(_u10_n12877 ), .ZN(_u10_n12864 ) );
NAND2_X1 _u10_U1339  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12870 ) );
NAND2_X1 _u10_U1338  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12871 ) );
NAND2_X1 _u10_U1337  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12872 ) );
NAND2_X1 _u10_U1336  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12873 ) );
NAND4_X1 _u10_U1335  ( .A1(_u10_n12870 ), .A2(_u10_n12871 ), .A3(_u10_n12872 ), .A4(_u10_n12873 ), .ZN(_u10_n12865 ) );
NAND2_X1 _u10_U1334  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12867 ) );
NAND2_X1 _u10_U1333  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12868 ) );
NAND2_X1 _u10_U1332  ( .A1(1'b0), .A2(_u10_n12019 ), .ZN(_u10_n12869 ) );
NAND3_X1 _u10_U1331  ( .A1(_u10_n12867 ), .A2(_u10_n12868 ), .A3(_u10_n12869 ), .ZN(_u10_n12866 ) );
NOR4_X1 _u10_U1330  ( .A1(_u10_n12863 ), .A2(_u10_n12864 ), .A3(_u10_n12865 ), .A4(_u10_n12866 ), .ZN(_u10_n12841 ) );
NAND2_X1 _u10_U1329  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n12859 ) );
NAND2_X1 _u10_U1328  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n12860 ) );
NAND2_X1 _u10_U1327  ( .A1(1'b0), .A2(_u10_n11948 ), .ZN(_u10_n12861 ) );
NAND2_X1 _u10_U1326  ( .A1(1'b0), .A2(_u10_n11924 ), .ZN(_u10_n12862 ) );
NAND4_X1 _u10_U1325  ( .A1(_u10_n12859 ), .A2(_u10_n12860 ), .A3(_u10_n12861 ), .A4(_u10_n12862 ), .ZN(_u10_n12843 ) );
NAND2_X1 _u10_U1324  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n12855 ) );
NAND2_X1 _u10_U1323  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n12856 ) );
NAND2_X1 _u10_U1322  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n12857 ) );
NAND2_X1 _u10_U1321  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n12858 ) );
NAND4_X1 _u10_U1320  ( .A1(_u10_n12855 ), .A2(_u10_n12856 ), .A3(_u10_n12857 ), .A4(_u10_n12858 ), .ZN(_u10_n12844 ) );
NAND2_X1 _u10_U1319  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n12851 ) );
NAND2_X1 _u10_U1318  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n12852 ) );
NAND2_X1 _u10_U1317  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n12853 ) );
NAND2_X1 _u10_U1316  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n12854 ) );
NAND4_X1 _u10_U1315  ( .A1(_u10_n12851 ), .A2(_u10_n12852 ), .A3(_u10_n12853 ), .A4(_u10_n12854 ), .ZN(_u10_n12845 ) );
NAND2_X1 _u10_U1314  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n12847 ) );
NAND2_X1 _u10_U1313  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n12848 ) );
NAND2_X1 _u10_U1312  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n12849 ) );
NAND2_X1 _u10_U1311  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n12850 ) );
NAND4_X1 _u10_U1310  ( .A1(_u10_n12847 ), .A2(_u10_n12848 ), .A3(_u10_n12849 ), .A4(_u10_n12850 ), .ZN(_u10_n12846 ) );
NOR4_X1 _u10_U1309  ( .A1(_u10_n12843 ), .A2(_u10_n12844 ), .A3(_u10_n12845 ), .A4(_u10_n12846 ), .ZN(_u10_n12842 ) );
NAND2_X1 _u10_U1308  ( .A1(_u10_n12841 ), .A2(_u10_n12842 ), .ZN(txsz[28]));
NAND2_X1 _u10_U1307  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12837 ) );
NAND2_X1 _u10_U1306  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12838 ) );
NAND2_X1 _u10_U1305  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n12839 ) );
NAND2_X1 _u10_U1304  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n12840 ) );
NAND4_X1 _u10_U1303  ( .A1(_u10_n12837 ), .A2(_u10_n12838 ), .A3(_u10_n12839 ), .A4(_u10_n12840 ), .ZN(_u10_n12822 ) );
NAND2_X1 _u10_U1302  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12833 ) );
NAND2_X1 _u10_U1301  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12834 ) );
NAND2_X1 _u10_U1300  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12835 ) );
NAND2_X1 _u10_U1299  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12836 ) );
NAND4_X1 _u10_U1298  ( .A1(_u10_n12833 ), .A2(_u10_n12834 ), .A3(_u10_n12835 ), .A4(_u10_n12836 ), .ZN(_u10_n12823 ) );
NAND2_X1 _u10_U1297  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12829 ) );
NAND2_X1 _u10_U1296  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12830 ) );
NAND2_X1 _u10_U1295  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12831 ) );
NAND2_X1 _u10_U1294  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12832 ) );
NAND4_X1 _u10_U1293  ( .A1(_u10_n12829 ), .A2(_u10_n12830 ), .A3(_u10_n12831 ), .A4(_u10_n12832 ), .ZN(_u10_n12824 ) );
NAND2_X1 _u10_U1292  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12826 ) );
NAND2_X1 _u10_U1291  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12827 ) );
NAND2_X1 _u10_U1290  ( .A1(1'b0), .A2(_u10_n12019 ), .ZN(_u10_n12828 ) );
NAND3_X1 _u10_U1289  ( .A1(_u10_n12826 ), .A2(_u10_n12827 ), .A3(_u10_n12828 ), .ZN(_u10_n12825 ) );
NOR4_X1 _u10_U1288  ( .A1(_u10_n12822 ), .A2(_u10_n12823 ), .A3(_u10_n12824 ), .A4(_u10_n12825 ), .ZN(_u10_n12800 ) );
NAND2_X1 _u10_U1287  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n12818 ) );
NAND2_X1 _u10_U1286  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n12819 ) );
NAND2_X1 _u10_U1285  ( .A1(1'b0), .A2(_u10_n11951 ), .ZN(_u10_n12820 ) );
NAND2_X1 _u10_U1284  ( .A1(1'b0), .A2(_u10_n11927 ), .ZN(_u10_n12821 ) );
NAND4_X1 _u10_U1283  ( .A1(_u10_n12818 ), .A2(_u10_n12819 ), .A3(_u10_n12820 ), .A4(_u10_n12821 ), .ZN(_u10_n12802 ) );
NAND2_X1 _u10_U1282  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n12814 ) );
NAND2_X1 _u10_U1281  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n12815 ) );
NAND2_X1 _u10_U1280  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n12816 ) );
NAND2_X1 _u10_U1279  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n12817 ) );
NAND4_X1 _u10_U1278  ( .A1(_u10_n12814 ), .A2(_u10_n12815 ), .A3(_u10_n12816 ), .A4(_u10_n12817 ), .ZN(_u10_n12803 ) );
NAND2_X1 _u10_U1277  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n12810 ) );
NAND2_X1 _u10_U1276  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n12811 ) );
NAND2_X1 _u10_U1275  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n12812 ) );
NAND2_X1 _u10_U1274  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n12813 ) );
NAND4_X1 _u10_U1273  ( .A1(_u10_n12810 ), .A2(_u10_n12811 ), .A3(_u10_n12812 ), .A4(_u10_n12813 ), .ZN(_u10_n12804 ) );
NAND2_X1 _u10_U1272  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n12806 ) );
NAND2_X1 _u10_U1271  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n12807 ) );
NAND2_X1 _u10_U1270  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n12808 ) );
NAND2_X1 _u10_U1269  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n12809 ) );
NAND4_X1 _u10_U1268  ( .A1(_u10_n12806 ), .A2(_u10_n12807 ), .A3(_u10_n12808 ), .A4(_u10_n12809 ), .ZN(_u10_n12805 ) );
NOR4_X1 _u10_U1267  ( .A1(_u10_n12802 ), .A2(_u10_n12803 ), .A3(_u10_n12804 ), .A4(_u10_n12805 ), .ZN(_u10_n12801 ) );
NAND2_X1 _u10_U1266  ( .A1(_u10_n12800 ), .A2(_u10_n12801 ), .ZN(txsz[29]));
NAND2_X1 _u10_U1265  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12796 ) );
NAND2_X1 _u10_U1264  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12797 ) );
NAND2_X1 _u10_U1263  ( .A1(1'b0), .A2(_u10_n12428 ), .ZN(_u10_n12798 ) );
NAND2_X1 _u10_U1262  ( .A1(1'b0), .A2(_u10_n12427 ), .ZN(_u10_n12799 ) );
NAND4_X1 _u10_U1261  ( .A1(_u10_n12796 ), .A2(_u10_n12797 ), .A3(_u10_n12798 ), .A4(_u10_n12799 ), .ZN(_u10_n12781 ) );
NAND2_X1 _u10_U1260  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12792 ) );
NAND2_X1 _u10_U1259  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12793 ) );
NAND2_X1 _u10_U1258  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12794 ) );
NAND2_X1 _u10_U1257  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12795 ) );
NAND4_X1 _u10_U1256  ( .A1(_u10_n12792 ), .A2(_u10_n12793 ), .A3(_u10_n12794 ), .A4(_u10_n12795 ), .ZN(_u10_n12782 ) );
NAND2_X1 _u10_U1255  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12788 ) );
NAND2_X1 _u10_U1254  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12789 ) );
NAND2_X1 _u10_U1253  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12790 ) );
NAND2_X1 _u10_U1252  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12791 ) );
NAND4_X1 _u10_U1251  ( .A1(_u10_n12788 ), .A2(_u10_n12789 ), .A3(_u10_n12790 ), .A4(_u10_n12791 ), .ZN(_u10_n12783 ) );
NAND2_X1 _u10_U1250  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12785 ) );
NAND2_X1 _u10_U1249  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12786 ) );
NAND2_X1 _u10_U1248  ( .A1(ch0_txsz[2]), .A2(_u10_n12019 ), .ZN(_u10_n12787 ) );
NAND3_X1 _u10_U1247  ( .A1(_u10_n12785 ), .A2(_u10_n12786 ), .A3(_u10_n12787 ), .ZN(_u10_n12784 ) );
NOR4_X1 _u10_U1246  ( .A1(_u10_n12781 ), .A2(_u10_n12782 ), .A3(_u10_n12783 ), .A4(_u10_n12784 ), .ZN(_u10_n12759 ) );
NAND2_X1 _u10_U1245  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n12777 ) );
NAND2_X1 _u10_U1244  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n12778 ) );
NAND2_X1 _u10_U1243  ( .A1(1'b0), .A2(_u10_n11947 ), .ZN(_u10_n12779 ) );
NAND2_X1 _u10_U1242  ( .A1(1'b0), .A2(_u10_n11923 ), .ZN(_u10_n12780 ) );
NAND4_X1 _u10_U1241  ( .A1(_u10_n12777 ), .A2(_u10_n12778 ), .A3(_u10_n12779 ), .A4(_u10_n12780 ), .ZN(_u10_n12761 ) );
NAND2_X1 _u10_U1240  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n12773 ) );
NAND2_X1 _u10_U1239  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n12774 ) );
NAND2_X1 _u10_U1238  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n12775 ) );
NAND2_X1 _u10_U1237  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n12776 ) );
NAND4_X1 _u10_U1236  ( .A1(_u10_n12773 ), .A2(_u10_n12774 ), .A3(_u10_n12775 ), .A4(_u10_n12776 ), .ZN(_u10_n12762 ) );
NAND2_X1 _u10_U1235  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n12769 ) );
NAND2_X1 _u10_U1234  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n12770 ) );
NAND2_X1 _u10_U1233  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n12771 ) );
NAND2_X1 _u10_U1232  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n12772 ) );
NAND4_X1 _u10_U1231  ( .A1(_u10_n12769 ), .A2(_u10_n12770 ), .A3(_u10_n12771 ), .A4(_u10_n12772 ), .ZN(_u10_n12763 ) );
NAND2_X1 _u10_U1230  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n12765 ) );
NAND2_X1 _u10_U1229  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n12766 ) );
NAND2_X1 _u10_U1228  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n12767 ) );
NAND2_X1 _u10_U1227  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n12768 ) );
NAND4_X1 _u10_U1226  ( .A1(_u10_n12765 ), .A2(_u10_n12766 ), .A3(_u10_n12767 ), .A4(_u10_n12768 ), .ZN(_u10_n12764 ) );
NOR4_X1 _u10_U1225  ( .A1(_u10_n12761 ), .A2(_u10_n12762 ), .A3(_u10_n12763 ), .A4(_u10_n12764 ), .ZN(_u10_n12760 ) );
NAND2_X1 _u10_U1224  ( .A1(_u10_n12759 ), .A2(_u10_n12760 ), .ZN(txsz[2]) );
NAND2_X1 _u10_U1223  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12755 ) );
NAND2_X1 _u10_U1222  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12756 ) );
NAND2_X1 _u10_U1221  ( .A1(1'b0), .A2(_u10_n12304 ), .ZN(_u10_n12757 ) );
NAND2_X1 _u10_U1220  ( .A1(1'b0), .A2(_u10_n12280 ), .ZN(_u10_n12758 ) );
NAND4_X1 _u10_U1219  ( .A1(_u10_n12755 ), .A2(_u10_n12756 ), .A3(_u10_n12757 ), .A4(_u10_n12758 ), .ZN(_u10_n12740 ) );
NAND2_X1 _u10_U1218  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12751 ) );
NAND2_X1 _u10_U1217  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12752 ) );
NAND2_X1 _u10_U1216  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12753 ) );
NAND2_X1 _u10_U1215  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12754 ) );
NAND4_X1 _u10_U1214  ( .A1(_u10_n12751 ), .A2(_u10_n12752 ), .A3(_u10_n12753 ), .A4(_u10_n12754 ), .ZN(_u10_n12741 ) );
NAND2_X1 _u10_U1213  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12747 ) );
NAND2_X1 _u10_U1212  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12748 ) );
NAND2_X1 _u10_U1211  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12749 ) );
NAND2_X1 _u10_U1210  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12750 ) );
NAND4_X1 _u10_U1209  ( .A1(_u10_n12747 ), .A2(_u10_n12748 ), .A3(_u10_n12749 ), .A4(_u10_n12750 ), .ZN(_u10_n12742 ) );
NAND2_X1 _u10_U1208  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12744 ) );
NAND2_X1 _u10_U1207  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12745 ) );
NAND2_X1 _u10_U1206  ( .A1(1'b0), .A2(_u10_n12019 ), .ZN(_u10_n12746 ) );
NAND3_X1 _u10_U1205  ( .A1(_u10_n12744 ), .A2(_u10_n12745 ), .A3(_u10_n12746 ), .ZN(_u10_n12743 ) );
NOR4_X1 _u10_U1204  ( .A1(_u10_n12740 ), .A2(_u10_n12741 ), .A3(_u10_n12742 ), .A4(_u10_n12743 ), .ZN(_u10_n12718 ) );
NAND2_X1 _u10_U1203  ( .A1(1'b0), .A2(_u10_n11983 ), .ZN(_u10_n12736 ) );
NAND2_X1 _u10_U1202  ( .A1(1'b0), .A2(_u10_n11959 ), .ZN(_u10_n12737 ) );
NAND2_X1 _u10_U1201  ( .A1(1'b0), .A2(_u10_n11946 ), .ZN(_u10_n12738 ) );
NAND2_X1 _u10_U1200  ( .A1(1'b0), .A2(_u10_n11922 ), .ZN(_u10_n12739 ) );
NAND4_X1 _u10_U1199  ( .A1(_u10_n12736 ), .A2(_u10_n12737 ), .A3(_u10_n12738 ), .A4(_u10_n12739 ), .ZN(_u10_n12720 ) );
NAND2_X1 _u10_U1198  ( .A1(1'b0), .A2(_u10_n11887 ), .ZN(_u10_n12732 ) );
NAND2_X1 _u10_U1197  ( .A1(1'b0), .A2(_u10_n11863 ), .ZN(_u10_n12733 ) );
NAND2_X1 _u10_U1196  ( .A1(1'b0), .A2(_u10_n11839 ), .ZN(_u10_n12734 ) );
NAND2_X1 _u10_U1195  ( .A1(1'b0), .A2(_u10_n11815 ), .ZN(_u10_n12735 ) );
NAND4_X1 _u10_U1194  ( .A1(_u10_n12732 ), .A2(_u10_n12733 ), .A3(_u10_n12734 ), .A4(_u10_n12735 ), .ZN(_u10_n12721 ) );
NAND2_X1 _u10_U1193  ( .A1(1'b0), .A2(_u10_n11791 ), .ZN(_u10_n12728 ) );
NAND2_X1 _u10_U1192  ( .A1(1'b0), .A2(_u10_n11767 ), .ZN(_u10_n12729 ) );
NAND2_X1 _u10_U1191  ( .A1(1'b0), .A2(_u10_n11743 ), .ZN(_u10_n12730 ) );
NAND2_X1 _u10_U1190  ( .A1(1'b0), .A2(_u10_n11719 ), .ZN(_u10_n12731 ) );
NAND4_X1 _u10_U1189  ( .A1(_u10_n12728 ), .A2(_u10_n12729 ), .A3(_u10_n12730 ), .A4(_u10_n12731 ), .ZN(_u10_n12722 ) );
NAND2_X1 _u10_U1188  ( .A1(1'b0), .A2(_u10_n11695 ), .ZN(_u10_n12724 ) );
NAND2_X1 _u10_U1187  ( .A1(1'b0), .A2(_u10_n11671 ), .ZN(_u10_n12725 ) );
NAND2_X1 _u10_U1186  ( .A1(1'b0), .A2(_u10_n11647 ), .ZN(_u10_n12726 ) );
NAND2_X1 _u10_U1185  ( .A1(1'b0), .A2(_u10_n11623 ), .ZN(_u10_n12727 ) );
NAND4_X1 _u10_U1184  ( .A1(_u10_n12724 ), .A2(_u10_n12725 ), .A3(_u10_n12726 ), .A4(_u10_n12727 ), .ZN(_u10_n12723 ) );
NOR4_X1 _u10_U1183  ( .A1(_u10_n12720 ), .A2(_u10_n12721 ), .A3(_u10_n12722 ), .A4(_u10_n12723 ), .ZN(_u10_n12719 ) );
NAND2_X1 _u10_U1182  ( .A1(_u10_n12718 ), .A2(_u10_n12719 ), .ZN(txsz[30]));
NAND2_X1 _u10_U1181  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12714 ) );
NAND2_X1 _u10_U1180  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12715 ) );
NAND2_X1 _u10_U1179  ( .A1(1'b0), .A2(_u10_n12307 ), .ZN(_u10_n12716 ) );
NAND2_X1 _u10_U1178  ( .A1(1'b0), .A2(_u10_n12283 ), .ZN(_u10_n12717 ) );
NAND4_X1 _u10_U1177  ( .A1(_u10_n12714 ), .A2(_u10_n12715 ), .A3(_u10_n12716 ), .A4(_u10_n12717 ), .ZN(_u10_n12699 ) );
NAND2_X1 _u10_U1176  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12710 ) );
NAND2_X1 _u10_U1175  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12711 ) );
NAND2_X1 _u10_U1174  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12712 ) );
NAND2_X1 _u10_U1173  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12713 ) );
NAND4_X1 _u10_U1172  ( .A1(_u10_n12710 ), .A2(_u10_n12711 ), .A3(_u10_n12712 ), .A4(_u10_n12713 ), .ZN(_u10_n12700 ) );
NAND2_X1 _u10_U1171  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12706 ) );
NAND2_X1 _u10_U1170  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12707 ) );
NAND2_X1 _u10_U1169  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12708 ) );
NAND2_X1 _u10_U1168  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12709 ) );
NAND4_X1 _u10_U1167  ( .A1(_u10_n12706 ), .A2(_u10_n12707 ), .A3(_u10_n12708 ), .A4(_u10_n12709 ), .ZN(_u10_n12701 ) );
NAND2_X1 _u10_U1166  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12703 ) );
NAND2_X1 _u10_U1165  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12704 ) );
NAND2_X1 _u10_U1164  ( .A1(1'b0), .A2(_u10_n12019 ), .ZN(_u10_n12705 ) );
NAND3_X1 _u10_U1163  ( .A1(_u10_n12703 ), .A2(_u10_n12704 ), .A3(_u10_n12705 ), .ZN(_u10_n12702 ) );
NOR4_X1 _u10_U1162  ( .A1(_u10_n12699 ), .A2(_u10_n12700 ), .A3(_u10_n12701 ), .A4(_u10_n12702 ), .ZN(_u10_n12677 ) );
NAND2_X1 _u10_U1161  ( .A1(1'b0), .A2(_u10_n11998 ), .ZN(_u10_n12695 ) );
NAND2_X1 _u10_U1160  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n12696 ) );
NAND2_X1 _u10_U1159  ( .A1(1'b0), .A2(_u10_n11951 ), .ZN(_u10_n12697 ) );
NAND2_X1 _u10_U1158  ( .A1(1'b0), .A2(_u10_n11927 ), .ZN(_u10_n12698 ) );
NAND4_X1 _u10_U1157  ( .A1(_u10_n12695 ), .A2(_u10_n12696 ), .A3(_u10_n12697 ), .A4(_u10_n12698 ), .ZN(_u10_n12679 ) );
NAND2_X1 _u10_U1156  ( .A1(1'b0), .A2(_u10_n11901 ), .ZN(_u10_n12691 ) );
NAND2_X1 _u10_U1155  ( .A1(1'b0), .A2(_u10_n11878 ), .ZN(_u10_n12692 ) );
NAND2_X1 _u10_U1154  ( .A1(1'b0), .A2(_u10_n11853 ), .ZN(_u10_n12693 ) );
NAND2_X1 _u10_U1153  ( .A1(1'b0), .A2(_u10_n11829 ), .ZN(_u10_n12694 ) );
NAND4_X1 _u10_U1152  ( .A1(_u10_n12691 ), .A2(_u10_n12692 ), .A3(_u10_n12693 ), .A4(_u10_n12694 ), .ZN(_u10_n12680 ) );
NAND2_X1 _u10_U1151  ( .A1(1'b0), .A2(_u10_n11806 ), .ZN(_u10_n12687 ) );
NAND2_X1 _u10_U1150  ( .A1(1'b0), .A2(_u10_n11782 ), .ZN(_u10_n12688 ) );
NAND2_X1 _u10_U1149  ( .A1(1'b0), .A2(_u10_n11759 ), .ZN(_u10_n12689 ) );
NAND2_X1 _u10_U1148  ( .A1(1'b0), .A2(_u10_n11735 ), .ZN(_u10_n12690 ) );
NAND4_X1 _u10_U1147  ( .A1(_u10_n12687 ), .A2(_u10_n12688 ), .A3(_u10_n12689 ), .A4(_u10_n12690 ), .ZN(_u10_n12681 ) );
NAND2_X1 _u10_U1146  ( .A1(1'b0), .A2(_u10_n11711 ), .ZN(_u10_n12683 ) );
NAND2_X1 _u10_U1145  ( .A1(1'b0), .A2(_u10_n11687 ), .ZN(_u10_n12684 ) );
NAND2_X1 _u10_U1144  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n12685 ) );
NAND2_X1 _u10_U1143  ( .A1(1'b0), .A2(_u10_n11637 ), .ZN(_u10_n12686 ) );
NAND4_X1 _u10_U1142  ( .A1(_u10_n12683 ), .A2(_u10_n12684 ), .A3(_u10_n12685 ), .A4(_u10_n12686 ), .ZN(_u10_n12682 ) );
NOR4_X1 _u10_U1141  ( .A1(_u10_n12679 ), .A2(_u10_n12680 ), .A3(_u10_n12681 ), .A4(_u10_n12682 ), .ZN(_u10_n12678 ) );
NAND2_X1 _u10_U1140  ( .A1(_u10_n12677 ), .A2(_u10_n12678 ), .ZN(txsz[31]));
NAND2_X1 _u10_U1139  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12673 ) );
NAND2_X1 _u10_U1138  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12674 ) );
NAND2_X1 _u10_U1137  ( .A1(1'b0), .A2(_u10_n12306 ), .ZN(_u10_n12675 ) );
NAND2_X1 _u10_U1136  ( .A1(1'b0), .A2(_u10_n12282 ), .ZN(_u10_n12676 ) );
NAND4_X1 _u10_U1135  ( .A1(_u10_n12673 ), .A2(_u10_n12674 ), .A3(_u10_n12675 ), .A4(_u10_n12676 ), .ZN(_u10_n12658 ) );
NAND2_X1 _u10_U1134  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12669 ) );
NAND2_X1 _u10_U1133  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12670 ) );
NAND2_X1 _u10_U1132  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12671 ) );
NAND2_X1 _u10_U1131  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12672 ) );
NAND4_X1 _u10_U1130  ( .A1(_u10_n12669 ), .A2(_u10_n12670 ), .A3(_u10_n12671 ), .A4(_u10_n12672 ), .ZN(_u10_n12659 ) );
NAND2_X1 _u10_U1129  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12665 ) );
NAND2_X1 _u10_U1128  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12666 ) );
NAND2_X1 _u10_U1127  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12667 ) );
NAND2_X1 _u10_U1126  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12668 ) );
NAND4_X1 _u10_U1125  ( .A1(_u10_n12665 ), .A2(_u10_n12666 ), .A3(_u10_n12667 ), .A4(_u10_n12668 ), .ZN(_u10_n12660 ) );
NAND2_X1 _u10_U1124  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12662 ) );
NAND2_X1 _u10_U1123  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12663 ) );
NAND2_X1 _u10_U1122  ( .A1(ch0_txsz[3]), .A2(_u10_n12019 ), .ZN(_u10_n12664 ) );
NAND3_X1 _u10_U1121  ( .A1(_u10_n12662 ), .A2(_u10_n12663 ), .A3(_u10_n12664 ), .ZN(_u10_n12661 ) );
NOR4_X1 _u10_U1120  ( .A1(_u10_n12658 ), .A2(_u10_n12659 ), .A3(_u10_n12660 ), .A4(_u10_n12661 ), .ZN(_u10_n12636 ) );
NAND2_X1 _u10_U1119  ( .A1(1'b0), .A2(_u10_n11999 ), .ZN(_u10_n12654 ) );
NAND2_X1 _u10_U1118  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n12655 ) );
NAND2_X1 _u10_U1117  ( .A1(1'b0), .A2(_u10_n11947 ), .ZN(_u10_n12656 ) );
NAND2_X1 _u10_U1116  ( .A1(1'b0), .A2(_u10_n11923 ), .ZN(_u10_n12657 ) );
NAND4_X1 _u10_U1115  ( .A1(_u10_n12654 ), .A2(_u10_n12655 ), .A3(_u10_n12656 ), .A4(_u10_n12657 ), .ZN(_u10_n12638 ) );
NAND2_X1 _u10_U1114  ( .A1(1'b0), .A2(_u10_n11903 ), .ZN(_u10_n12650 ) );
NAND2_X1 _u10_U1113  ( .A1(1'b0), .A2(_u10_n11879 ), .ZN(_u10_n12651 ) );
NAND2_X1 _u10_U1112  ( .A1(1'b0), .A2(_u10_n11854 ), .ZN(_u10_n12652 ) );
NAND2_X1 _u10_U1111  ( .A1(1'b0), .A2(_u10_n11831 ), .ZN(_u10_n12653 ) );
NAND4_X1 _u10_U1110  ( .A1(_u10_n12650 ), .A2(_u10_n12651 ), .A3(_u10_n12652 ), .A4(_u10_n12653 ), .ZN(_u10_n12639 ) );
NAND2_X1 _u10_U1109  ( .A1(1'b0), .A2(_u10_n11807 ), .ZN(_u10_n12646 ) );
NAND2_X1 _u10_U1108  ( .A1(1'b0), .A2(_u10_n11783 ), .ZN(_u10_n12647 ) );
NAND2_X1 _u10_U1107  ( .A1(1'b0), .A2(_u10_n11758 ), .ZN(_u10_n12648 ) );
NAND2_X1 _u10_U1106  ( .A1(1'b0), .A2(_u10_n11734 ), .ZN(_u10_n12649 ) );
NAND4_X1 _u10_U1105  ( .A1(_u10_n12646 ), .A2(_u10_n12647 ), .A3(_u10_n12648 ), .A4(_u10_n12649 ), .ZN(_u10_n12640 ) );
NAND2_X1 _u10_U1104  ( .A1(1'b0), .A2(_u10_n11710 ), .ZN(_u10_n12642 ) );
NAND2_X1 _u10_U1103  ( .A1(1'b0), .A2(_u10_n11686 ), .ZN(_u10_n12643 ) );
NAND2_X1 _u10_U1102  ( .A1(1'b0), .A2(_u10_n11661 ), .ZN(_u10_n12644 ) );
NAND2_X1 _u10_U1101  ( .A1(1'b0), .A2(_u10_n11638 ), .ZN(_u10_n12645 ) );
NAND4_X1 _u10_U1100  ( .A1(_u10_n12642 ), .A2(_u10_n12643 ), .A3(_u10_n12644 ), .A4(_u10_n12645 ), .ZN(_u10_n12641 ) );
NOR4_X1 _u10_U1099  ( .A1(_u10_n12638 ), .A2(_u10_n12639 ), .A3(_u10_n12640 ), .A4(_u10_n12641 ), .ZN(_u10_n12637 ) );
NAND2_X1 _u10_U1098  ( .A1(_u10_n12636 ), .A2(_u10_n12637 ), .ZN(txsz[3]) );
NAND2_X1 _u10_U1097  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12632 ) );
NAND2_X1 _u10_U1096  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12633 ) );
NAND2_X1 _u10_U1095  ( .A1(1'b0), .A2(_u10_n12305 ), .ZN(_u10_n12634 ) );
NAND2_X1 _u10_U1094  ( .A1(1'b0), .A2(_u10_n12281 ), .ZN(_u10_n12635 ) );
NAND4_X1 _u10_U1093  ( .A1(_u10_n12632 ), .A2(_u10_n12633 ), .A3(_u10_n12634 ), .A4(_u10_n12635 ), .ZN(_u10_n12617 ) );
NAND2_X1 _u10_U1092  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12628 ) );
NAND2_X1 _u10_U1091  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12629 ) );
NAND2_X1 _u10_U1090  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12630 ) );
NAND2_X1 _u10_U1089  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12631 ) );
NAND4_X1 _u10_U1088  ( .A1(_u10_n12628 ), .A2(_u10_n12629 ), .A3(_u10_n12630 ), .A4(_u10_n12631 ), .ZN(_u10_n12618 ) );
NAND2_X1 _u10_U1087  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12624 ) );
NAND2_X1 _u10_U1086  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12625 ) );
NAND2_X1 _u10_U1085  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12626 ) );
NAND2_X1 _u10_U1084  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12627 ) );
NAND4_X1 _u10_U1083  ( .A1(_u10_n12624 ), .A2(_u10_n12625 ), .A3(_u10_n12626 ), .A4(_u10_n12627 ), .ZN(_u10_n12619 ) );
NAND2_X1 _u10_U1082  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12621 ) );
NAND2_X1 _u10_U1081  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12622 ) );
NAND2_X1 _u10_U1080  ( .A1(ch0_txsz[4]), .A2(_u10_n12019 ), .ZN(_u10_n12623 ) );
NAND3_X1 _u10_U1079  ( .A1(_u10_n12621 ), .A2(_u10_n12622 ), .A3(_u10_n12623 ), .ZN(_u10_n12620 ) );
NOR4_X1 _u10_U1078  ( .A1(_u10_n12617 ), .A2(_u10_n12618 ), .A3(_u10_n12619 ), .A4(_u10_n12620 ), .ZN(_u10_n12595 ) );
NAND2_X1 _u10_U1077  ( .A1(1'b0), .A2(_u10_n11993 ), .ZN(_u10_n12613 ) );
NAND2_X1 _u10_U1076  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n12614 ) );
NAND2_X1 _u10_U1075  ( .A1(1'b0), .A2(_u10_n11946 ), .ZN(_u10_n12615 ) );
NAND2_X1 _u10_U1074  ( .A1(1'b0), .A2(_u10_n11922 ), .ZN(_u10_n12616 ) );
NAND4_X1 _u10_U1073  ( .A1(_u10_n12613 ), .A2(_u10_n12614 ), .A3(_u10_n12615 ), .A4(_u10_n12616 ), .ZN(_u10_n12597 ) );
NAND2_X1 _u10_U1072  ( .A1(1'b0), .A2(_u10_n11902 ), .ZN(_u10_n12609 ) );
NAND2_X1 _u10_U1071  ( .A1(1'b0), .A2(_u10_n11873 ), .ZN(_u10_n12610 ) );
NAND2_X1 _u10_U1070  ( .A1(1'b0), .A2(_u10_n11855 ), .ZN(_u10_n12611 ) );
NAND2_X1 _u10_U1069  ( .A1(1'b0), .A2(_u10_n11830 ), .ZN(_u10_n12612 ) );
NAND4_X1 _u10_U1068  ( .A1(_u10_n12609 ), .A2(_u10_n12610 ), .A3(_u10_n12611 ), .A4(_u10_n12612 ), .ZN(_u10_n12598 ) );
NAND2_X1 _u10_U1067  ( .A1(1'b0), .A2(_u10_n11801 ), .ZN(_u10_n12605 ) );
NAND2_X1 _u10_U1066  ( .A1(1'b0), .A2(_u10_n12379 ), .ZN(_u10_n12606 ) );
NAND2_X1 _u10_U1065  ( .A1(1'b0), .A2(_u10_n11756 ), .ZN(_u10_n12607 ) );
NAND2_X1 _u10_U1064  ( .A1(1'b0), .A2(_u10_n11732 ), .ZN(_u10_n12608 ) );
NAND4_X1 _u10_U1063  ( .A1(_u10_n12605 ), .A2(_u10_n12606 ), .A3(_u10_n12607 ), .A4(_u10_n12608 ), .ZN(_u10_n12599 ) );
NAND2_X1 _u10_U1062  ( .A1(1'b0), .A2(_u10_n11708 ), .ZN(_u10_n12601 ) );
NAND2_X1 _u10_U1061  ( .A1(1'b0), .A2(_u10_n11684 ), .ZN(_u10_n12602 ) );
NAND2_X1 _u10_U1060  ( .A1(1'b0), .A2(_u10_n11663 ), .ZN(_u10_n12603 ) );
NAND2_X1 _u10_U1059  ( .A1(1'b0), .A2(_u10_n11639 ), .ZN(_u10_n12604 ) );
NAND4_X1 _u10_U1058  ( .A1(_u10_n12601 ), .A2(_u10_n12602 ), .A3(_u10_n12603 ), .A4(_u10_n12604 ), .ZN(_u10_n12600 ) );
NOR4_X1 _u10_U1057  ( .A1(_u10_n12597 ), .A2(_u10_n12598 ), .A3(_u10_n12599 ), .A4(_u10_n12600 ), .ZN(_u10_n12596 ) );
NAND2_X1 _u10_U1056  ( .A1(_u10_n12595 ), .A2(_u10_n12596 ), .ZN(txsz[4]) );
NAND2_X1 _u10_U1055  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12591 ) );
NAND2_X1 _u10_U1054  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12592 ) );
NAND2_X1 _u10_U1053  ( .A1(1'b0), .A2(_u10_n12303 ), .ZN(_u10_n12593 ) );
NAND2_X1 _u10_U1052  ( .A1(1'b0), .A2(_u10_n12279 ), .ZN(_u10_n12594 ) );
NAND4_X1 _u10_U1051  ( .A1(_u10_n12591 ), .A2(_u10_n12592 ), .A3(_u10_n12593 ), .A4(_u10_n12594 ), .ZN(_u10_n12576 ) );
NAND2_X1 _u10_U1050  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12587 ) );
NAND2_X1 _u10_U1049  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12588 ) );
NAND2_X1 _u10_U1048  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12589 ) );
NAND2_X1 _u10_U1047  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12590 ) );
NAND4_X1 _u10_U1046  ( .A1(_u10_n12587 ), .A2(_u10_n12588 ), .A3(_u10_n12589 ), .A4(_u10_n12590 ), .ZN(_u10_n12577 ) );
NAND2_X1 _u10_U1045  ( .A1(1'b0), .A2(_u10_n12157 ), .ZN(_u10_n12583 ) );
NAND2_X1 _u10_U1044  ( .A1(1'b0), .A2(_u10_n12133 ), .ZN(_u10_n12584 ) );
NAND2_X1 _u10_U1043  ( .A1(1'b0), .A2(_u10_n12109 ), .ZN(_u10_n12585 ) );
NAND2_X1 _u10_U1042  ( .A1(1'b0), .A2(_u10_n12085 ), .ZN(_u10_n12586 ) );
NAND4_X1 _u10_U1041  ( .A1(_u10_n12583 ), .A2(_u10_n12584 ), .A3(_u10_n12585 ), .A4(_u10_n12586 ), .ZN(_u10_n12578 ) );
NAND2_X1 _u10_U1040  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12580 ) );
NAND2_X1 _u10_U1039  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12581 ) );
NAND2_X1 _u10_U1038  ( .A1(ch0_txsz[5]), .A2(_u10_n12020 ), .ZN(_u10_n12582 ) );
NAND3_X1 _u10_U1037  ( .A1(_u10_n12580 ), .A2(_u10_n12581 ), .A3(_u10_n12582 ), .ZN(_u10_n12579 ) );
NOR4_X1 _u10_U1036  ( .A1(_u10_n12576 ), .A2(_u10_n12577 ), .A3(_u10_n12578 ), .A4(_u10_n12579 ), .ZN(_u10_n12554 ) );
NAND2_X1 _u10_U1035  ( .A1(1'b0), .A2(_u10_n11993 ), .ZN(_u10_n12572 ) );
NAND2_X1 _u10_U1034  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n12573 ) );
NAND2_X1 _u10_U1033  ( .A1(1'b0), .A2(_u10_n11950 ), .ZN(_u10_n12574 ) );
NAND2_X1 _u10_U1032  ( .A1(1'b0), .A2(_u10_n11926 ), .ZN(_u10_n12575 ) );
NAND4_X1 _u10_U1031  ( .A1(_u10_n12572 ), .A2(_u10_n12573 ), .A3(_u10_n12574 ), .A4(_u10_n12575 ), .ZN(_u10_n12556 ) );
NAND2_X1 _u10_U1030  ( .A1(1'b0), .A2(_u10_n11897 ), .ZN(_u10_n12568 ) );
NAND2_X1 _u10_U1029  ( .A1(1'b0), .A2(_u10_n11873 ), .ZN(_u10_n12569 ) );
NAND2_X1 _u10_U1028  ( .A1(1'b0), .A2(_u10_n11849 ), .ZN(_u10_n12570 ) );
NAND2_X1 _u10_U1027  ( .A1(1'b0), .A2(_u10_n11825 ), .ZN(_u10_n12571 ) );
NAND4_X1 _u10_U1026  ( .A1(_u10_n12568 ), .A2(_u10_n12569 ), .A3(_u10_n12570 ), .A4(_u10_n12571 ), .ZN(_u10_n12557 ) );
NAND2_X1 _u10_U1025  ( .A1(1'b0), .A2(_u10_n11801 ), .ZN(_u10_n12564 ) );
NAND2_X1 _u10_U1024  ( .A1(1'b0), .A2(_u10_n11777 ), .ZN(_u10_n12565 ) );
NAND2_X1 _u10_U1023  ( .A1(1'b0), .A2(_u10_n11753 ), .ZN(_u10_n12566 ) );
NAND2_X1 _u10_U1022  ( .A1(1'b0), .A2(_u10_n11729 ), .ZN(_u10_n12567 ) );
NAND4_X1 _u10_U1021  ( .A1(_u10_n12564 ), .A2(_u10_n12565 ), .A3(_u10_n12566 ), .A4(_u10_n12567 ), .ZN(_u10_n12558 ) );
NAND2_X1 _u10_U1020  ( .A1(1'b0), .A2(_u10_n11705 ), .ZN(_u10_n12560 ) );
NAND2_X1 _u10_U1019  ( .A1(1'b0), .A2(_u10_n11681 ), .ZN(_u10_n12561 ) );
NAND2_X1 _u10_U1018  ( .A1(1'b0), .A2(_u10_n11657 ), .ZN(_u10_n12562 ) );
NAND2_X1 _u10_U1017  ( .A1(1'b0), .A2(_u10_n11633 ), .ZN(_u10_n12563 ) );
NAND4_X1 _u10_U1016  ( .A1(_u10_n12560 ), .A2(_u10_n12561 ), .A3(_u10_n12562 ), .A4(_u10_n12563 ), .ZN(_u10_n12559 ) );
NOR4_X1 _u10_U1015  ( .A1(_u10_n12556 ), .A2(_u10_n12557 ), .A3(_u10_n12558 ), .A4(_u10_n12559 ), .ZN(_u10_n12555 ) );
NAND2_X1 _u10_U1014  ( .A1(_u10_n12554 ), .A2(_u10_n12555 ), .ZN(txsz[5]) );
NAND2_X1 _u10_U1013  ( .A1(1'b0), .A2(_u10_n12351 ), .ZN(_u10_n12550 ) );
NAND2_X1 _u10_U1012  ( .A1(1'b0), .A2(_u10_n12327 ), .ZN(_u10_n12551 ) );
NAND2_X1 _u10_U1011  ( .A1(1'b0), .A2(_u10_n12308 ), .ZN(_u10_n12552 ) );
NAND2_X1 _u10_U1010  ( .A1(1'b0), .A2(_u10_n12284 ), .ZN(_u10_n12553 ) );
NAND4_X1 _u10_U1009  ( .A1(_u10_n12550 ), .A2(_u10_n12551 ), .A3(_u10_n12552 ), .A4(_u10_n12553 ), .ZN(_u10_n12535 ) );
NAND2_X1 _u10_U1008  ( .A1(1'b0), .A2(_u10_n12255 ), .ZN(_u10_n12546 ) );
NAND2_X1 _u10_U1007  ( .A1(1'b0), .A2(_u10_n12231 ), .ZN(_u10_n12547 ) );
NAND2_X1 _u10_U1006  ( .A1(1'b0), .A2(_u10_n12205 ), .ZN(_u10_n12548 ) );
NAND2_X1 _u10_U1005  ( .A1(1'b0), .A2(_u10_n12183 ), .ZN(_u10_n12549 ) );
NAND4_X1 _u10_U1004  ( .A1(_u10_n12546 ), .A2(_u10_n12547 ), .A3(_u10_n12548 ), .A4(_u10_n12549 ), .ZN(_u10_n12536 ) );
NAND2_X1 _u10_U1003  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n12542 ) );
NAND2_X1 _u10_U1002  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n12543 ) );
NAND2_X1 _u10_U1001  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n12544 ) );
NAND2_X1 _u10_U1000  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n12545 ) );
NAND4_X1 _u10_U999  ( .A1(_u10_n12542 ), .A2(_u10_n12543 ), .A3(_u10_n12544 ), .A4(_u10_n12545 ), .ZN(_u10_n12537 ) );
NAND2_X1 _u10_U998  ( .A1(1'b0), .A2(_u10_n12061 ), .ZN(_u10_n12539 ) );
NAND2_X1 _u10_U997  ( .A1(1'b0), .A2(_u10_n12037 ), .ZN(_u10_n12540 ) );
NAND2_X1 _u10_U996  ( .A1(ch0_txsz[6]), .A2(_u10_n12020 ), .ZN(_u10_n12541 ));
NAND3_X1 _u10_U995  ( .A1(_u10_n12539 ), .A2(_u10_n12540 ), .A3(_u10_n12541 ), .ZN(_u10_n12538 ) );
NOR4_X1 _u10_U994  ( .A1(_u10_n12535 ), .A2(_u10_n12536 ), .A3(_u10_n12537 ),.A4(_u10_n12538 ), .ZN(_u10_n12513 ) );
NAND2_X1 _u10_U993  ( .A1(1'b0), .A2(_u10_n11995 ), .ZN(_u10_n12531 ) );
NAND2_X1 _u10_U992  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n12532 ) );
NAND2_X1 _u10_U991  ( .A1(1'b0), .A2(_u10_n12394 ), .ZN(_u10_n12533 ) );
NAND2_X1 _u10_U990  ( .A1(1'b0), .A2(_u10_n12393 ), .ZN(_u10_n12534 ) );
NAND4_X1 _u10_U989  ( .A1(_u10_n12531 ), .A2(_u10_n12532 ), .A3(_u10_n12533 ), .A4(_u10_n12534 ), .ZN(_u10_n12515 ) );
NAND2_X1 _u10_U988  ( .A1(1'b0), .A2(_u10_n11902 ), .ZN(_u10_n12527 ) );
NAND2_X1 _u10_U987  ( .A1(1'b0), .A2(_u10_n11875 ), .ZN(_u10_n12528 ) );
NAND2_X1 _u10_U986  ( .A1(1'b0), .A2(_u10_n11854 ), .ZN(_u10_n12529 ) );
NAND2_X1 _u10_U985  ( .A1(1'b0), .A2(_u10_n11830 ), .ZN(_u10_n12530 ) );
NAND4_X1 _u10_U984  ( .A1(_u10_n12527 ), .A2(_u10_n12528 ), .A3(_u10_n12529 ), .A4(_u10_n12530 ), .ZN(_u10_n12516 ) );
NAND2_X1 _u10_U983  ( .A1(1'b0), .A2(_u10_n11803 ), .ZN(_u10_n12523 ) );
NAND2_X1 _u10_U982  ( .A1(1'b0), .A2(_u10_n11781 ), .ZN(_u10_n12524 ) );
NAND2_X1 _u10_U981  ( .A1(1'b0), .A2(_u10_n11758 ), .ZN(_u10_n12525 ) );
NAND2_X1 _u10_U980  ( .A1(1'b0), .A2(_u10_n11734 ), .ZN(_u10_n12526 ) );
NAND4_X1 _u10_U979  ( .A1(_u10_n12523 ), .A2(_u10_n12524 ), .A3(_u10_n12525 ), .A4(_u10_n12526 ), .ZN(_u10_n12517 ) );
NAND2_X1 _u10_U978  ( .A1(1'b0), .A2(_u10_n11710 ), .ZN(_u10_n12519 ) );
NAND2_X1 _u10_U977  ( .A1(1'b0), .A2(_u10_n11686 ), .ZN(_u10_n12520 ) );
NAND2_X1 _u10_U976  ( .A1(1'b0), .A2(_u10_n11662 ), .ZN(_u10_n12521 ) );
NAND2_X1 _u10_U975  ( .A1(1'b0), .A2(_u10_n11638 ), .ZN(_u10_n12522 ) );
NAND4_X1 _u10_U974  ( .A1(_u10_n12519 ), .A2(_u10_n12520 ), .A3(_u10_n12521 ), .A4(_u10_n12522 ), .ZN(_u10_n12518 ) );
NOR4_X1 _u10_U973  ( .A1(_u10_n12515 ), .A2(_u10_n12516 ), .A3(_u10_n12517 ),.A4(_u10_n12518 ), .ZN(_u10_n12514 ) );
NAND2_X1 _u10_U972  ( .A1(_u10_n12513 ), .A2(_u10_n12514 ), .ZN(txsz[6]) );
NAND2_X1 _u10_U971  ( .A1(1'b0), .A2(_u10_n12352 ), .ZN(_u10_n12509 ) );
NAND2_X1 _u10_U970  ( .A1(1'b0), .A2(_u10_n12332 ), .ZN(_u10_n12510 ) );
NAND2_X1 _u10_U969  ( .A1(1'b0), .A2(_u10_n12307 ), .ZN(_u10_n12511 ) );
NAND2_X1 _u10_U968  ( .A1(1'b0), .A2(_u10_n12283 ), .ZN(_u10_n12512 ) );
NAND4_X1 _u10_U967  ( .A1(_u10_n12509 ), .A2(_u10_n12510 ), .A3(_u10_n12511 ), .A4(_u10_n12512 ), .ZN(_u10_n12494 ) );
NAND2_X1 _u10_U966  ( .A1(1'b0), .A2(_u10_n12256 ), .ZN(_u10_n12505 ) );
NAND2_X1 _u10_U965  ( .A1(1'b0), .A2(_u10_n12232 ), .ZN(_u10_n12506 ) );
NAND2_X1 _u10_U964  ( .A1(1'b0), .A2(_u10_n12206 ), .ZN(_u10_n12507 ) );
NAND2_X1 _u10_U963  ( .A1(1'b0), .A2(_u10_n12184 ), .ZN(_u10_n12508 ) );
NAND4_X1 _u10_U962  ( .A1(_u10_n12505 ), .A2(_u10_n12506 ), .A3(_u10_n12507 ), .A4(_u10_n12508 ), .ZN(_u10_n12495 ) );
NAND2_X1 _u10_U961  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n12501 ) );
NAND2_X1 _u10_U960  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n12502 ) );
NAND2_X1 _u10_U959  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n12503 ) );
NAND2_X1 _u10_U958  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n12504 ) );
NAND4_X1 _u10_U957  ( .A1(_u10_n12501 ), .A2(_u10_n12502 ), .A3(_u10_n12503 ), .A4(_u10_n12504 ), .ZN(_u10_n12496 ) );
NAND2_X1 _u10_U956  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n12498 ) );
NAND2_X1 _u10_U955  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n12499 ) );
NAND2_X1 _u10_U954  ( .A1(ch0_txsz[7]), .A2(_u10_n12020 ), .ZN(_u10_n12500 ));
NAND3_X1 _u10_U953  ( .A1(_u10_n12498 ), .A2(_u10_n12499 ), .A3(_u10_n12500 ), .ZN(_u10_n12497 ) );
NOR4_X1 _u10_U952  ( .A1(_u10_n12494 ), .A2(_u10_n12495 ), .A3(_u10_n12496 ),.A4(_u10_n12497 ), .ZN(_u10_n12472 ) );
NAND2_X1 _u10_U951  ( .A1(1'b0), .A2(_u10_n11996 ), .ZN(_u10_n12490 ) );
NAND2_X1 _u10_U950  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n12491 ) );
NAND2_X1 _u10_U949  ( .A1(1'b0), .A2(_u10_n11950 ), .ZN(_u10_n12492 ) );
NAND2_X1 _u10_U948  ( .A1(1'b0), .A2(_u10_n11926 ), .ZN(_u10_n12493 ) );
NAND4_X1 _u10_U947  ( .A1(_u10_n12490 ), .A2(_u10_n12491 ), .A3(_u10_n12492 ), .A4(_u10_n12493 ), .ZN(_u10_n12474 ) );
NAND2_X1 _u10_U946  ( .A1(1'b0), .A2(_u10_n11900 ), .ZN(_u10_n12486 ) );
NAND2_X1 _u10_U945  ( .A1(1'b0), .A2(_u10_n11876 ), .ZN(_u10_n12487 ) );
NAND2_X1 _u10_U944  ( .A1(1'b0), .A2(_u10_n11852 ), .ZN(_u10_n12488 ) );
NAND2_X1 _u10_U943  ( .A1(1'b0), .A2(_u10_n11828 ), .ZN(_u10_n12489 ) );
NAND4_X1 _u10_U942  ( .A1(_u10_n12486 ), .A2(_u10_n12487 ), .A3(_u10_n12488 ), .A4(_u10_n12489 ), .ZN(_u10_n12475 ) );
NAND2_X1 _u10_U941  ( .A1(1'b0), .A2(_u10_n11804 ), .ZN(_u10_n12482 ) );
NAND2_X1 _u10_U940  ( .A1(1'b0), .A2(_u10_n11780 ), .ZN(_u10_n12483 ) );
NAND2_X1 _u10_U939  ( .A1(1'b0), .A2(_u10_n11756 ), .ZN(_u10_n12484 ) );
NAND2_X1 _u10_U938  ( .A1(1'b0), .A2(_u10_n11732 ), .ZN(_u10_n12485 ) );
NAND4_X1 _u10_U937  ( .A1(_u10_n12482 ), .A2(_u10_n12483 ), .A3(_u10_n12484 ), .A4(_u10_n12485 ), .ZN(_u10_n12476 ) );
NAND2_X1 _u10_U936  ( .A1(1'b0), .A2(_u10_n11708 ), .ZN(_u10_n12478 ) );
NAND2_X1 _u10_U935  ( .A1(1'b0), .A2(_u10_n11684 ), .ZN(_u10_n12479 ) );
NAND2_X1 _u10_U934  ( .A1(1'b0), .A2(_u10_n11660 ), .ZN(_u10_n12480 ) );
NAND2_X1 _u10_U933  ( .A1(1'b0), .A2(_u10_n11636 ), .ZN(_u10_n12481 ) );
NAND4_X1 _u10_U932  ( .A1(_u10_n12478 ), .A2(_u10_n12479 ), .A3(_u10_n12480 ), .A4(_u10_n12481 ), .ZN(_u10_n12477 ) );
NOR4_X1 _u10_U931  ( .A1(_u10_n12474 ), .A2(_u10_n12475 ), .A3(_u10_n12476 ),.A4(_u10_n12477 ), .ZN(_u10_n12473 ) );
NAND2_X1 _u10_U930  ( .A1(_u10_n12472 ), .A2(_u10_n12473 ), .ZN(txsz[7]) );
NAND2_X1 _u10_U929  ( .A1(1'b0), .A2(_u10_n12352 ), .ZN(_u10_n12468 ) );
NAND2_X1 _u10_U928  ( .A1(1'b0), .A2(_u10_n12331 ), .ZN(_u10_n12469 ) );
NAND2_X1 _u10_U927  ( .A1(1'b0), .A2(_u10_n12306 ), .ZN(_u10_n12470 ) );
NAND2_X1 _u10_U926  ( .A1(1'b0), .A2(_u10_n12282 ), .ZN(_u10_n12471 ) );
NAND4_X1 _u10_U925  ( .A1(_u10_n12468 ), .A2(_u10_n12469 ), .A3(_u10_n12470 ), .A4(_u10_n12471 ), .ZN(_u10_n12453 ) );
NAND2_X1 _u10_U924  ( .A1(1'b0), .A2(_u10_n12256 ), .ZN(_u10_n12464 ) );
NAND2_X1 _u10_U923  ( .A1(1'b0), .A2(_u10_n12232 ), .ZN(_u10_n12465 ) );
NAND2_X1 _u10_U922  ( .A1(1'b0), .A2(_u10_n12206 ), .ZN(_u10_n12466 ) );
NAND2_X1 _u10_U921  ( .A1(1'b0), .A2(_u10_n12184 ), .ZN(_u10_n12467 ) );
NAND4_X1 _u10_U920  ( .A1(_u10_n12464 ), .A2(_u10_n12465 ), .A3(_u10_n12466 ), .A4(_u10_n12467 ), .ZN(_u10_n12454 ) );
NAND2_X1 _u10_U919  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n12460 ) );
NAND2_X1 _u10_U918  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n12461 ) );
NAND2_X1 _u10_U917  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n12462 ) );
NAND2_X1 _u10_U916  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n12463 ) );
NAND4_X1 _u10_U915  ( .A1(_u10_n12460 ), .A2(_u10_n12461 ), .A3(_u10_n12462 ), .A4(_u10_n12463 ), .ZN(_u10_n12455 ) );
NAND2_X1 _u10_U914  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n12457 ) );
NAND2_X1 _u10_U913  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n12458 ) );
NAND2_X1 _u10_U912  ( .A1(ch0_txsz[8]), .A2(_u10_n12020 ), .ZN(_u10_n12459 ));
NAND3_X1 _u10_U911  ( .A1(_u10_n12457 ), .A2(_u10_n12458 ), .A3(_u10_n12459 ), .ZN(_u10_n12456 ) );
NOR4_X1 _u10_U910  ( .A1(_u10_n12453 ), .A2(_u10_n12454 ), .A3(_u10_n12455 ),.A4(_u10_n12456 ), .ZN(_u10_n12431 ) );
NAND2_X1 _u10_U909  ( .A1(1'b0), .A2(_u10_n11994 ), .ZN(_u10_n12449 ) );
NAND2_X1 _u10_U908  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n12450 ) );
NAND2_X1 _u10_U907  ( .A1(1'b0), .A2(_u10_n11949 ), .ZN(_u10_n12451 ) );
NAND2_X1 _u10_U906  ( .A1(1'b0), .A2(_u10_n11925 ), .ZN(_u10_n12452 ) );
NAND4_X1 _u10_U905  ( .A1(_u10_n12449 ), .A2(_u10_n12450 ), .A3(_u10_n12451 ), .A4(_u10_n12452 ), .ZN(_u10_n12433 ) );
NAND2_X1 _u10_U904  ( .A1(1'b0), .A2(_u10_n11898 ), .ZN(_u10_n12445 ) );
NAND2_X1 _u10_U903  ( .A1(1'b0), .A2(_u10_n11874 ), .ZN(_u10_n12446 ) );
NAND2_X1 _u10_U902  ( .A1(1'b0), .A2(_u10_n11850 ), .ZN(_u10_n12447 ) );
NAND2_X1 _u10_U901  ( .A1(1'b0), .A2(_u10_n11826 ), .ZN(_u10_n12448 ) );
NAND4_X1 _u10_U900  ( .A1(_u10_n12445 ), .A2(_u10_n12446 ), .A3(_u10_n12447 ), .A4(_u10_n12448 ), .ZN(_u10_n12434 ) );
NAND2_X1 _u10_U899  ( .A1(1'b0), .A2(_u10_n11802 ), .ZN(_u10_n12441 ) );
NAND2_X1 _u10_U898  ( .A1(1'b0), .A2(_u10_n11778 ), .ZN(_u10_n12442 ) );
NAND2_X1 _u10_U897  ( .A1(1'b0), .A2(_u10_n11754 ), .ZN(_u10_n12443 ) );
NAND2_X1 _u10_U896  ( .A1(1'b0), .A2(_u10_n11730 ), .ZN(_u10_n12444 ) );
NAND4_X1 _u10_U895  ( .A1(_u10_n12441 ), .A2(_u10_n12442 ), .A3(_u10_n12443 ), .A4(_u10_n12444 ), .ZN(_u10_n12435 ) );
NAND2_X1 _u10_U894  ( .A1(1'b0), .A2(_u10_n11706 ), .ZN(_u10_n12437 ) );
NAND2_X1 _u10_U893  ( .A1(1'b0), .A2(_u10_n11682 ), .ZN(_u10_n12438 ) );
NAND2_X1 _u10_U892  ( .A1(1'b0), .A2(_u10_n11658 ), .ZN(_u10_n12439 ) );
NAND2_X1 _u10_U891  ( .A1(1'b0), .A2(_u10_n11634 ), .ZN(_u10_n12440 ) );
NAND4_X1 _u10_U890  ( .A1(_u10_n12437 ), .A2(_u10_n12438 ), .A3(_u10_n12439 ), .A4(_u10_n12440 ), .ZN(_u10_n12436 ) );
NOR4_X1 _u10_U889  ( .A1(_u10_n12433 ), .A2(_u10_n12434 ), .A3(_u10_n12435 ),.A4(_u10_n12436 ), .ZN(_u10_n12432 ) );
NAND2_X1 _u10_U888  ( .A1(_u10_n12431 ), .A2(_u10_n12432 ), .ZN(txsz[8]) );
NAND2_X1 _u10_U887  ( .A1(1'b0), .A2(_u10_n12352 ), .ZN(_u10_n12423 ) );
NAND2_X1 _u10_U886  ( .A1(1'b0), .A2(_u10_n12331 ), .ZN(_u10_n12424 ) );
NAND2_X1 _u10_U885  ( .A1(1'b0), .A2(_u10_n12305 ), .ZN(_u10_n12425 ) );
NAND2_X1 _u10_U884  ( .A1(1'b0), .A2(_u10_n12281 ), .ZN(_u10_n12426 ) );
NAND4_X1 _u10_U883  ( .A1(_u10_n12423 ), .A2(_u10_n12424 ), .A3(_u10_n12425 ), .A4(_u10_n12426 ), .ZN(_u10_n12397 ) );
NAND2_X1 _u10_U882  ( .A1(1'b0), .A2(_u10_n12256 ), .ZN(_u10_n12415 ) );
NAND2_X1 _u10_U881  ( .A1(1'b0), .A2(_u10_n12232 ), .ZN(_u10_n12416 ) );
NAND2_X1 _u10_U880  ( .A1(1'b0), .A2(_u10_n12206 ), .ZN(_u10_n12417 ) );
NAND2_X1 _u10_U879  ( .A1(1'b0), .A2(_u10_n12184 ), .ZN(_u10_n12418 ) );
NAND4_X1 _u10_U878  ( .A1(_u10_n12415 ), .A2(_u10_n12416 ), .A3(_u10_n12417 ), .A4(_u10_n12418 ), .ZN(_u10_n12398 ) );
NAND2_X1 _u10_U877  ( .A1(1'b0), .A2(_u10_n12158 ), .ZN(_u10_n12407 ) );
NAND2_X1 _u10_U876  ( .A1(1'b0), .A2(_u10_n12134 ), .ZN(_u10_n12408 ) );
NAND2_X1 _u10_U875  ( .A1(1'b0), .A2(_u10_n12110 ), .ZN(_u10_n12409 ) );
NAND2_X1 _u10_U874  ( .A1(1'b0), .A2(_u10_n12086 ), .ZN(_u10_n12410 ) );
NAND4_X1 _u10_U873  ( .A1(_u10_n12407 ), .A2(_u10_n12408 ), .A3(_u10_n12409 ), .A4(_u10_n12410 ), .ZN(_u10_n12399 ) );
NAND2_X1 _u10_U872  ( .A1(1'b0), .A2(_u10_n12062 ), .ZN(_u10_n12401 ) );
NAND2_X1 _u10_U871  ( .A1(1'b0), .A2(_u10_n12038 ), .ZN(_u10_n12402 ) );
NAND2_X1 _u10_U870  ( .A1(ch0_txsz[9]), .A2(_u10_n12020 ), .ZN(_u10_n12403 ));
NAND3_X1 _u10_U869  ( .A1(_u10_n12401 ), .A2(_u10_n12402 ), .A3(_u10_n12403 ), .ZN(_u10_n12400 ) );
NOR4_X1 _u10_U868  ( .A1(_u10_n12397 ), .A2(_u10_n12398 ), .A3(_u10_n12399 ),.A4(_u10_n12400 ), .ZN(_u10_n12359 ) );
NAND2_X1 _u10_U867  ( .A1(1'b0), .A2(_u10_n11995 ), .ZN(_u10_n12389 ) );
NAND2_X1 _u10_U866  ( .A1(1'b0), .A2(_u10_n11960 ), .ZN(_u10_n12390 ) );
NAND2_X1 _u10_U865  ( .A1(1'b0), .A2(_u10_n11945 ), .ZN(_u10_n12391 ) );
NAND2_X1 _u10_U864  ( .A1(1'b0), .A2(_u10_n11921 ), .ZN(_u10_n12392 ) );
NAND4_X1 _u10_U863  ( .A1(_u10_n12389 ), .A2(_u10_n12390 ), .A3(_u10_n12391 ), .A4(_u10_n12392 ), .ZN(_u10_n12361 ) );
NAND2_X1 _u10_U862  ( .A1(1'b0), .A2(_u10_n11899 ), .ZN(_u10_n12381 ) );
NAND2_X1 _u10_U861  ( .A1(1'b0), .A2(_u10_n11875 ), .ZN(_u10_n12382 ) );
NAND2_X1 _u10_U860  ( .A1(1'b0), .A2(_u10_n11851 ), .ZN(_u10_n12383 ) );
NAND2_X1 _u10_U859  ( .A1(1'b0), .A2(_u10_n11827 ), .ZN(_u10_n12384 ) );
NAND4_X1 _u10_U858  ( .A1(_u10_n12381 ), .A2(_u10_n12382 ), .A3(_u10_n12383 ), .A4(_u10_n12384 ), .ZN(_u10_n12362 ) );
NAND2_X1 _u10_U857  ( .A1(1'b0), .A2(_u10_n11803 ), .ZN(_u10_n12373 ) );
NAND2_X1 _u10_U856  ( .A1(1'b0), .A2(_u10_n11779 ), .ZN(_u10_n12374 ) );
NAND2_X1 _u10_U855  ( .A1(1'b0), .A2(_u10_n11755 ), .ZN(_u10_n12375 ) );
NAND2_X1 _u10_U854  ( .A1(1'b0), .A2(_u10_n11731 ), .ZN(_u10_n12376 ) );
NAND4_X1 _u10_U853  ( .A1(_u10_n12373 ), .A2(_u10_n12374 ), .A3(_u10_n12375 ), .A4(_u10_n12376 ), .ZN(_u10_n12363 ) );
NAND2_X1 _u10_U852  ( .A1(1'b0), .A2(_u10_n11707 ), .ZN(_u10_n12365 ) );
NAND2_X1 _u10_U851  ( .A1(1'b0), .A2(_u10_n11683 ), .ZN(_u10_n12366 ) );
NAND2_X1 _u10_U850  ( .A1(1'b0), .A2(_u10_n11659 ), .ZN(_u10_n12367 ) );
NAND2_X1 _u10_U849  ( .A1(1'b0), .A2(_u10_n11635 ), .ZN(_u10_n12368 ) );
NAND4_X1 _u10_U848  ( .A1(_u10_n12365 ), .A2(_u10_n12366 ), .A3(_u10_n12367 ), .A4(_u10_n12368 ), .ZN(_u10_n12364 ) );
NOR4_X1 _u10_U847  ( .A1(_u10_n12361 ), .A2(_u10_n12362 ), .A3(_u10_n12363 ),.A4(_u10_n12364 ), .ZN(_u10_n12360 ) );
NAND2_X1 _u10_U846  ( .A1(_u10_n12359 ), .A2(_u10_n12360 ), .ZN(txsz[9]) );
INV_X4 _u10_U845  ( .A(n5), .ZN(_u10_n12358 ) );
INV_X8 _u10_U844  ( .A(_u10_n12358 ), .ZN(_u10_n12357 ) );
BUF_X4 _u10_U843  ( .A(_u10_n12369 ), .Z(_u10_n11634 ) );
BUF_X4 _u10_U842  ( .A(_u10_n12370 ), .Z(_u10_n11658 ) );
BUF_X4 _u10_U841  ( .A(_u10_n12380 ), .Z(_u10_n11802 ) );
BUF_X4 _u10_U840  ( .A(_u10_n12396 ), .Z(_u10_n11994 ) );
BUF_X4 _u10_U839  ( .A(_u10_n12369 ), .Z(_u10_n11636 ) );
BUF_X4 _u10_U838  ( .A(_u10_n12370 ), .Z(_u10_n11660 ) );
BUF_X4 _u10_U837  ( .A(_u10_n12380 ), .Z(_u10_n11804 ) );
BUF_X4 _u10_U836  ( .A(_u10_n12396 ), .Z(_u10_n11996 ) );
BUF_X4 _u10_U835  ( .A(_u10_n12369 ), .Z(_u10_n11635 ) );
BUF_X4 _u10_U834  ( .A(_u10_n12370 ), .Z(_u10_n11659 ) );
BUF_X4 _u10_U833  ( .A(_u10_n12380 ), .Z(_u10_n11803 ) );
BUF_X4 _u10_U832  ( .A(_u10_n12396 ), .Z(_u10_n11995 ) );
BUF_X4 _u10_U831  ( .A(_u10_n12369 ), .Z(_u10_n11637 ) );
BUF_X4 _u10_U830  ( .A(_u10_n12370 ), .Z(_u10_n11661 ) );
BUF_X4 _u10_U829  ( .A(_u10_n12380 ), .Z(_u10_n11805 ) );
BUF_X4 _u10_U828  ( .A(_u10_n12396 ), .Z(_u10_n11997 ) );
BUF_X4 _u10_U827  ( .A(_u10_n12369 ), .Z(_u10_n11638 ) );
BUF_X4 _u10_U826  ( .A(_u10_n12370 ), .Z(_u10_n11662 ) );
BUF_X4 _u10_U825  ( .A(_u10_n12380 ), .Z(_u10_n11806 ) );
BUF_X4 _u10_U824  ( .A(_u10_n12396 ), .Z(_u10_n11998 ) );
BUF_X4 _u10_U823  ( .A(_u10_n12380 ), .Z(_u10_n11807 ) );
BUF_X4 _u10_U822  ( .A(_u10_n12396 ), .Z(_u10_n11999 ) );
BUF_X4 _u10_U821  ( .A(_u10_n12369 ), .Z(_u10_n11639 ) );
BUF_X4 _u10_U820  ( .A(_u10_n12370 ), .Z(_u10_n11663 ) );
BUF_X4 _u10_U819  ( .A(_u10_n12393 ), .Z(_u10_n11927 ) );
BUF_X4 _u10_U818  ( .A(_u10_n12395 ), .Z(_u10_n11975 ) );
BUF_X4 _u10_U817  ( .A(_u10_n12394 ), .Z(_u10_n11951 ) );
BUF_X4 _u10_U816  ( .A(_u10_n12393 ), .Z(_u10_n11925 ) );
BUF_X4 _u10_U815  ( .A(_u10_n12395 ), .Z(_u10_n11973 ) );
BUF_X4 _u10_U814  ( .A(_u10_n12394 ), .Z(_u10_n11949 ) );
BUF_X4 _u10_U813  ( .A(_u10_n12393 ), .Z(_u10_n11924 ) );
BUF_X4 _u10_U812  ( .A(_u10_n12395 ), .Z(_u10_n11972 ) );
BUF_X4 _u10_U811  ( .A(_u10_n12394 ), .Z(_u10_n11948 ) );
BUF_X4 _u10_U810  ( .A(_u10_n12393 ), .Z(_u10_n11923 ) );
BUF_X4 _u10_U809  ( .A(_u10_n12395 ), .Z(_u10_n11971 ) );
BUF_X4 _u10_U808  ( .A(_u10_n12394 ), .Z(_u10_n11947 ) );
BUF_X4 _u10_U807  ( .A(_u10_n12393 ), .Z(_u10_n11922 ) );
BUF_X4 _u10_U806  ( .A(_u10_n12395 ), .Z(_u10_n11970 ) );
BUF_X4 _u10_U805  ( .A(_u10_n12394 ), .Z(_u10_n11946 ) );
BUF_X4 _u10_U804  ( .A(_u10_n12395 ), .Z(_u10_n11974 ) );
BUF_X4 _u10_U803  ( .A(_u10_n12371 ), .Z(_u10_n11682 ) );
BUF_X4 _u10_U802  ( .A(_u10_n12372 ), .Z(_u10_n11706 ) );
BUF_X4 _u10_U801  ( .A(_u10_n12377 ), .Z(_u10_n11730 ) );
BUF_X4 _u10_U800  ( .A(_u10_n12379 ), .Z(_u10_n11778 ) );
BUF_X4 _u10_U799  ( .A(_u10_n12378 ), .Z(_u10_n11754 ) );
BUF_X4 _u10_U798  ( .A(_u10_n12385 ), .Z(_u10_n11826 ) );
BUF_X4 _u10_U797  ( .A(_u10_n12387 ), .Z(_u10_n11874 ) );
BUF_X4 _u10_U796  ( .A(_u10_n12386 ), .Z(_u10_n11850 ) );
BUF_X4 _u10_U795  ( .A(_u10_n12388 ), .Z(_u10_n11898 ) );
BUF_X4 _u10_U794  ( .A(_u10_n12411 ), .Z(_u10_n12089 ) );
BUF_X4 _u10_U793  ( .A(_u10_n12413 ), .Z(_u10_n12137 ) );
BUF_X4 _u10_U792  ( .A(_u10_n12412 ), .Z(_u10_n12113 ) );
BUF_X4 _u10_U791  ( .A(_u10_n12414 ), .Z(_u10_n12161 ) );
BUF_X4 _u10_U790  ( .A(_u10_n12371 ), .Z(_u10_n11684 ) );
BUF_X4 _u10_U789  ( .A(_u10_n12372 ), .Z(_u10_n11708 ) );
BUF_X4 _u10_U788  ( .A(_u10_n12377 ), .Z(_u10_n11732 ) );
BUF_X4 _u10_U787  ( .A(_u10_n12379 ), .Z(_u10_n11780 ) );
BUF_X4 _u10_U786  ( .A(_u10_n12378 ), .Z(_u10_n11756 ) );
BUF_X4 _u10_U785  ( .A(_u10_n12385 ), .Z(_u10_n11828 ) );
BUF_X4 _u10_U784  ( .A(_u10_n12387 ), .Z(_u10_n11876 ) );
BUF_X4 _u10_U783  ( .A(_u10_n12386 ), .Z(_u10_n11852 ) );
BUF_X4 _u10_U782  ( .A(_u10_n12388 ), .Z(_u10_n11900 ) );
BUF_X4 _u10_U781  ( .A(_u10_n12411 ), .Z(_u10_n12091 ) );
BUF_X4 _u10_U780  ( .A(_u10_n12413 ), .Z(_u10_n12139 ) );
BUF_X4 _u10_U779  ( .A(_u10_n12412 ), .Z(_u10_n12115 ) );
BUF_X4 _u10_U778  ( .A(_u10_n12414 ), .Z(_u10_n12163 ) );
BUF_X4 _u10_U777  ( .A(_u10_n12371 ), .Z(_u10_n11683 ) );
BUF_X4 _u10_U776  ( .A(_u10_n12372 ), .Z(_u10_n11707 ) );
BUF_X4 _u10_U775  ( .A(_u10_n12377 ), .Z(_u10_n11731 ) );
BUF_X4 _u10_U774  ( .A(_u10_n12379 ), .Z(_u10_n11779 ) );
BUF_X4 _u10_U773  ( .A(_u10_n12378 ), .Z(_u10_n11755 ) );
BUF_X4 _u10_U772  ( .A(_u10_n12385 ), .Z(_u10_n11827 ) );
BUF_X4 _u10_U771  ( .A(_u10_n12387 ), .Z(_u10_n11875 ) );
BUF_X4 _u10_U770  ( .A(_u10_n12386 ), .Z(_u10_n11851 ) );
BUF_X4 _u10_U769  ( .A(_u10_n12388 ), .Z(_u10_n11899 ) );
BUF_X4 _u10_U768  ( .A(_u10_n12411 ), .Z(_u10_n12090 ) );
BUF_X4 _u10_U767  ( .A(_u10_n12413 ), .Z(_u10_n12138 ) );
BUF_X4 _u10_U766  ( .A(_u10_n12412 ), .Z(_u10_n12114 ) );
BUF_X4 _u10_U765  ( .A(_u10_n12414 ), .Z(_u10_n12162 ) );
BUF_X4 _u10_U764  ( .A(_u10_n12371 ), .Z(_u10_n11685 ) );
BUF_X4 _u10_U763  ( .A(_u10_n12372 ), .Z(_u10_n11709 ) );
BUF_X4 _u10_U762  ( .A(_u10_n12377 ), .Z(_u10_n11733 ) );
BUF_X4 _u10_U761  ( .A(_u10_n12379 ), .Z(_u10_n11781 ) );
BUF_X4 _u10_U760  ( .A(_u10_n12378 ), .Z(_u10_n11757 ) );
BUF_X4 _u10_U759  ( .A(_u10_n12385 ), .Z(_u10_n11829 ) );
BUF_X4 _u10_U758  ( .A(_u10_n12387 ), .Z(_u10_n11877 ) );
BUF_X4 _u10_U757  ( .A(_u10_n12386 ), .Z(_u10_n11853 ) );
BUF_X4 _u10_U756  ( .A(_u10_n12388 ), .Z(_u10_n11901 ) );
BUF_X4 _u10_U755  ( .A(_u10_n12411 ), .Z(_u10_n12092 ) );
BUF_X4 _u10_U754  ( .A(_u10_n12413 ), .Z(_u10_n12140 ) );
BUF_X4 _u10_U753  ( .A(_u10_n12412 ), .Z(_u10_n12116 ) );
BUF_X4 _u10_U752  ( .A(_u10_n12414 ), .Z(_u10_n12164 ) );
BUF_X4 _u10_U751  ( .A(_u10_n12411 ), .Z(_u10_n12087 ) );
BUF_X4 _u10_U750  ( .A(_u10_n12413 ), .Z(_u10_n12135 ) );
BUF_X4 _u10_U749  ( .A(_u10_n12412 ), .Z(_u10_n12111 ) );
BUF_X4 _u10_U748  ( .A(_u10_n12414 ), .Z(_u10_n12159 ) );
BUF_X4 _u10_U747  ( .A(_u10_n12371 ), .Z(_u10_n11686 ) );
BUF_X4 _u10_U746  ( .A(_u10_n12372 ), .Z(_u10_n11710 ) );
BUF_X4 _u10_U745  ( .A(_u10_n12377 ), .Z(_u10_n11734 ) );
BUF_X4 _u10_U744  ( .A(_u10_n12378 ), .Z(_u10_n11758 ) );
BUF_X4 _u10_U743  ( .A(_u10_n12385 ), .Z(_u10_n11830 ) );
BUF_X4 _u10_U742  ( .A(_u10_n12386 ), .Z(_u10_n11854 ) );
BUF_X4 _u10_U741  ( .A(_u10_n12388 ), .Z(_u10_n11902 ) );
BUF_X4 _u10_U740  ( .A(_u10_n12371 ), .Z(_u10_n11687 ) );
BUF_X4 _u10_U739  ( .A(_u10_n12372 ), .Z(_u10_n11711 ) );
BUF_X4 _u10_U738  ( .A(_u10_n12377 ), .Z(_u10_n11735 ) );
BUF_X4 _u10_U737  ( .A(_u10_n12379 ), .Z(_u10_n11782 ) );
BUF_X4 _u10_U736  ( .A(_u10_n12378 ), .Z(_u10_n11759 ) );
BUF_X4 _u10_U735  ( .A(_u10_n12387 ), .Z(_u10_n11878 ) );
BUF_X4 _u10_U734  ( .A(_u10_n12393 ), .Z(_u10_n11926 ) );
BUF_X4 _u10_U733  ( .A(_u10_n12394 ), .Z(_u10_n11950 ) );
BUF_X4 _u10_U732  ( .A(_u10_n12379 ), .Z(_u10_n11783 ) );
BUF_X4 _u10_U731  ( .A(_u10_n12385 ), .Z(_u10_n11831 ) );
BUF_X4 _u10_U730  ( .A(_u10_n12387 ), .Z(_u10_n11879 ) );
BUF_X4 _u10_U729  ( .A(_u10_n12388 ), .Z(_u10_n11903 ) );
BUF_X4 _u10_U728  ( .A(_u10_n12411 ), .Z(_u10_n12088 ) );
BUF_X4 _u10_U727  ( .A(_u10_n12413 ), .Z(_u10_n12136 ) );
BUF_X4 _u10_U726  ( .A(_u10_n12412 ), .Z(_u10_n12112 ) );
BUF_X4 _u10_U725  ( .A(_u10_n12414 ), .Z(_u10_n12160 ) );
BUF_X4 _u10_U724  ( .A(_u10_n12386 ), .Z(_u10_n11855 ) );
BUF_X4 _u10_U723  ( .A(_u10_n11634 ), .Z(_u10_n11633 ) );
BUF_X4 _u10_U722  ( .A(_u10_n11658 ), .Z(_u10_n11657 ) );
BUF_X4 _u10_U721  ( .A(_u10_n11802 ), .Z(_u10_n11801 ) );
BUF_X4 _u10_U720  ( .A(_u10_n11994 ), .Z(_u10_n11993 ) );
BUF_X4 _u10_U719  ( .A(_u10_n11639 ), .Z(_u10_n11617 ) );
BUF_X4 _u10_U718  ( .A(_u10_n11663 ), .Z(_u10_n11641 ) );
BUF_X4 _u10_U717  ( .A(_u10_n11807 ), .Z(_u10_n11785 ) );
BUF_X4 _u10_U716  ( .A(_u10_n11999 ), .Z(_u10_n11977 ) );
BUF_X4 _u10_U715  ( .A(_u10_n11638 ), .Z(_u10_n11623 ) );
BUF_X4 _u10_U714  ( .A(_u10_n11662 ), .Z(_u10_n11647 ) );
BUF_X4 _u10_U713  ( .A(_u10_n11804 ), .Z(_u10_n11791 ) );
BUF_X4 _u10_U712  ( .A(_u10_n11996 ), .Z(_u10_n11983 ) );
BUF_X4 _u10_U711  ( .A(_u10_n11639 ), .Z(_u10_n11619 ) );
BUF_X4 _u10_U710  ( .A(_u10_n11663 ), .Z(_u10_n11643 ) );
BUF_X4 _u10_U709  ( .A(_u10_n11634 ), .Z(_u10_n11632 ) );
BUF_X4 _u10_U708  ( .A(_u10_n11658 ), .Z(_u10_n11656 ) );
BUF_X4 _u10_U707  ( .A(_u10_n11802 ), .Z(_u10_n11800 ) );
BUF_X4 _u10_U706  ( .A(_u10_n11994 ), .Z(_u10_n11992 ) );
BUF_X4 _u10_U705  ( .A(_u10_n11636 ), .Z(_u10_n11627 ) );
BUF_X4 _u10_U704  ( .A(_u10_n11660 ), .Z(_u10_n11651 ) );
BUF_X4 _u10_U703  ( .A(_u10_n11804 ), .Z(_u10_n11795 ) );
BUF_X4 _u10_U702  ( .A(_u10_n11996 ), .Z(_u10_n11987 ) );
BUF_X4 _u10_U701  ( .A(_u10_n11635 ), .Z(_u10_n11629 ) );
BUF_X4 _u10_U700  ( .A(_u10_n11659 ), .Z(_u10_n11653 ) );
BUF_X4 _u10_U699  ( .A(_u10_n11803 ), .Z(_u10_n11797 ) );
BUF_X4 _u10_U698  ( .A(_u10_n11995 ), .Z(_u10_n11989 ) );
BUF_X4 _u10_U697  ( .A(_u10_n11637 ), .Z(_u10_n11624 ) );
BUF_X4 _u10_U696  ( .A(_u10_n11661 ), .Z(_u10_n11648 ) );
BUF_X4 _u10_U695  ( .A(_u10_n11805 ), .Z(_u10_n11792 ) );
BUF_X4 _u10_U694  ( .A(_u10_n11997 ), .Z(_u10_n11984 ) );
BUF_X4 _u10_U693  ( .A(_u10_n11638 ), .Z(_u10_n11622 ) );
BUF_X4 _u10_U692  ( .A(_u10_n11662 ), .Z(_u10_n11646 ) );
BUF_X4 _u10_U691  ( .A(_u10_n11805 ), .Z(_u10_n11790 ) );
BUF_X4 _u10_U690  ( .A(_u10_n11997 ), .Z(_u10_n11982 ) );
BUF_X4 _u10_U689  ( .A(_u10_n11635 ), .Z(_u10_n11628 ) );
BUF_X4 _u10_U688  ( .A(_u10_n11659 ), .Z(_u10_n11652 ) );
BUF_X4 _u10_U687  ( .A(_u10_n11803 ), .Z(_u10_n11796 ) );
BUF_X4 _u10_U686  ( .A(_u10_n11995 ), .Z(_u10_n11988 ) );
BUF_X4 _u10_U685  ( .A(_u10_n11635 ), .Z(_u10_n11630 ) );
BUF_X4 _u10_U684  ( .A(_u10_n11659 ), .Z(_u10_n11654 ) );
BUF_X4 _u10_U683  ( .A(_u10_n11803 ), .Z(_u10_n11798 ) );
BUF_X4 _u10_U682  ( .A(_u10_n11995 ), .Z(_u10_n11990 ) );
BUF_X4 _u10_U681  ( .A(_u10_n11637 ), .Z(_u10_n11625 ) );
BUF_X4 _u10_U680  ( .A(_u10_n11661 ), .Z(_u10_n11649 ) );
BUF_X4 _u10_U679  ( .A(_u10_n11805 ), .Z(_u10_n11793 ) );
BUF_X4 _u10_U678  ( .A(_u10_n11997 ), .Z(_u10_n11985 ) );
BUF_X4 _u10_U677  ( .A(_u10_n11634 ), .Z(_u10_n11631 ) );
BUF_X4 _u10_U676  ( .A(_u10_n11658 ), .Z(_u10_n11655 ) );
BUF_X4 _u10_U675  ( .A(_u10_n11802 ), .Z(_u10_n11799 ) );
BUF_X4 _u10_U674  ( .A(_u10_n11994 ), .Z(_u10_n11991 ) );
BUF_X4 _u10_U673  ( .A(_u10_n11636 ), .Z(_u10_n11626 ) );
BUF_X4 _u10_U672  ( .A(_u10_n11660 ), .Z(_u10_n11650 ) );
BUF_X4 _u10_U671  ( .A(_u10_n11804 ), .Z(_u10_n11794 ) );
BUF_X4 _u10_U670  ( .A(_u10_n11996 ), .Z(_u10_n11986 ) );
BUF_X4 _u10_U669  ( .A(_u10_n12369 ), .Z(_u10_n11621 ) );
BUF_X4 _u10_U668  ( .A(_u10_n12370 ), .Z(_u10_n11645 ) );
BUF_X4 _u10_U667  ( .A(_u10_n11806 ), .Z(_u10_n11789 ) );
BUF_X4 _u10_U666  ( .A(_u10_n11998 ), .Z(_u10_n11981 ) );
BUF_X4 _u10_U665  ( .A(_u10_n11633 ), .Z(_u10_n11620 ) );
BUF_X4 _u10_U664  ( .A(_u10_n11657 ), .Z(_u10_n11644 ) );
BUF_X4 _u10_U663  ( .A(_u10_n11806 ), .Z(_u10_n11788 ) );
BUF_X4 _u10_U662  ( .A(_u10_n11998 ), .Z(_u10_n11980 ) );
BUF_X4 _u10_U661  ( .A(_u10_n11806 ), .Z(_u10_n11787 ) );
BUF_X4 _u10_U660  ( .A(_u10_n11998 ), .Z(_u10_n11979 ) );
BUF_X4 _u10_U659  ( .A(_u10_n11639 ), .Z(_u10_n11618 ) );
BUF_X4 _u10_U658  ( .A(_u10_n11663 ), .Z(_u10_n11642 ) );
BUF_X4 _u10_U657  ( .A(_u10_n12380 ), .Z(_u10_n11786 ) );
BUF_X4 _u10_U656  ( .A(_u10_n12396 ), .Z(_u10_n11978 ) );
BUF_X4 _u10_U655  ( .A(_u10_n11639 ), .Z(_u10_n11616 ) );
BUF_X4 _u10_U654  ( .A(_u10_n11663 ), .Z(_u10_n11640 ) );
BUF_X4 _u10_U653  ( .A(_u10_n11801 ), .Z(_u10_n11784 ) );
BUF_X4 _u10_U652  ( .A(_u10_n11993 ), .Z(_u10_n11976 ) );
BUF_X4 _u10_U651  ( .A(_u10_n12427 ), .Z(_u10_n12284 ) );
BUF_X4 _u10_U650  ( .A(_u10_n12429 ), .Z(_u10_n12332 ) );
BUF_X4 _u10_U649  ( .A(_u10_n12428 ), .Z(_u10_n12308 ) );
BUF_X4 _u10_U648  ( .A(_u10_n12427 ), .Z(_u10_n12283 ) );
BUF_X4 _u10_U647  ( .A(_u10_n12429 ), .Z(_u10_n12331 ) );
BUF_X4 _u10_U646  ( .A(_u10_n12428 ), .Z(_u10_n12307 ) );
BUF_X4 _u10_U645  ( .A(_u10_n12427 ), .Z(_u10_n12282 ) );
BUF_X4 _u10_U644  ( .A(_u10_n12429 ), .Z(_u10_n12330 ) );
BUF_X4 _u10_U643  ( .A(_u10_n12428 ), .Z(_u10_n12306 ) );
BUF_X4 _u10_U642  ( .A(_u10_n12427 ), .Z(_u10_n12281 ) );
BUF_X4 _u10_U641  ( .A(_u10_n12429 ), .Z(_u10_n12329 ) );
BUF_X4 _u10_U640  ( .A(_u10_n12428 ), .Z(_u10_n12305 ) );
BUF_X4 _u10_U639  ( .A(_u10_n12427 ), .Z(_u10_n12280 ) );
BUF_X4 _u10_U638  ( .A(_u10_n12429 ), .Z(_u10_n12328 ) );
BUF_X4 _u10_U637  ( .A(_u10_n12428 ), .Z(_u10_n12304 ) );
BUF_X4 _u10_U636  ( .A(_u10_n12405 ), .Z(_u10_n12041 ) );
BUF_X4 _u10_U635  ( .A(_u10_n12406 ), .Z(_u10_n12065 ) );
BUF_X4 _u10_U634  ( .A(_u10_n12419 ), .Z(_u10_n12186 ) );
BUF_X4 _u10_U633  ( .A(_u10_n12421 ), .Z(_u10_n12234 ) );
BUF_X4 _u10_U632  ( .A(_u10_n12420 ), .Z(_u10_n12209 ) );
BUF_X4 _u10_U631  ( .A(_u10_n12422 ), .Z(_u10_n12258 ) );
BUF_X4 _u10_U630  ( .A(_u10_n12430 ), .Z(_u10_n12354 ) );
BUF_X4 _u10_U629  ( .A(_u10_n12405 ), .Z(_u10_n12043 ) );
BUF_X4 _u10_U628  ( .A(_u10_n12406 ), .Z(_u10_n12067 ) );
BUF_X4 _u10_U627  ( .A(_u10_n12419 ), .Z(_u10_n12187 ) );
BUF_X4 _u10_U626  ( .A(_u10_n12421 ), .Z(_u10_n12235 ) );
BUF_X4 _u10_U625  ( .A(_u10_n12420 ), .Z(_u10_n12211 ) );
BUF_X4 _u10_U624  ( .A(_u10_n12422 ), .Z(_u10_n12259 ) );
BUF_X4 _u10_U623  ( .A(_u10_n12430 ), .Z(_u10_n12355 ) );
BUF_X4 _u10_U622  ( .A(_u10_n12405 ), .Z(_u10_n12042 ) );
BUF_X4 _u10_U621  ( .A(_u10_n12406 ), .Z(_u10_n12066 ) );
BUF_X4 _u10_U620  ( .A(_u10_n12420 ), .Z(_u10_n12210 ) );
BUF_X4 _u10_U619  ( .A(_u10_n12405 ), .Z(_u10_n12044 ) );
BUF_X4 _u10_U618  ( .A(_u10_n12406 ), .Z(_u10_n12068 ) );
BUF_X4 _u10_U617  ( .A(_u10_n12419 ), .Z(_u10_n12188 ) );
BUF_X4 _u10_U616  ( .A(_u10_n12421 ), .Z(_u10_n12236 ) );
BUF_X4 _u10_U615  ( .A(_u10_n12420 ), .Z(_u10_n12212 ) );
BUF_X4 _u10_U614  ( .A(_u10_n12422 ), .Z(_u10_n12260 ) );
BUF_X4 _u10_U613  ( .A(_u10_n12430 ), .Z(_u10_n12356 ) );
BUF_X4 _u10_U612  ( .A(_u10_n12405 ), .Z(_u10_n12039 ) );
BUF_X4 _u10_U611  ( .A(_u10_n12406 ), .Z(_u10_n12063 ) );
BUF_X4 _u10_U610  ( .A(_u10_n12419 ), .Z(_u10_n12185 ) );
BUF_X4 _u10_U609  ( .A(_u10_n12421 ), .Z(_u10_n12233 ) );
BUF_X4 _u10_U608  ( .A(_u10_n12420 ), .Z(_u10_n12207 ) );
BUF_X4 _u10_U607  ( .A(_u10_n12422 ), .Z(_u10_n12257 ) );
BUF_X4 _u10_U606  ( .A(_u10_n12430 ), .Z(_u10_n12353 ) );
BUF_X4 _u10_U605  ( .A(_u10_n12427 ), .Z(_u10_n12279 ) );
BUF_X4 _u10_U604  ( .A(_u10_n12428 ), .Z(_u10_n12303 ) );
BUF_X4 _u10_U603  ( .A(_u10_n12405 ), .Z(_u10_n12040 ) );
BUF_X4 _u10_U602  ( .A(_u10_n12406 ), .Z(_u10_n12064 ) );
BUF_X4 _u10_U601  ( .A(_u10_n12420 ), .Z(_u10_n12208 ) );
BUF_X4 _u10_U600  ( .A(_u10_n11922 ), .Z(_u10_n11921 ) );
BUF_X4 _u10_U599  ( .A(_u10_n11970 ), .Z(_u10_n11969 ) );
BUF_X4 _u10_U598  ( .A(_u10_n11946 ), .Z(_u10_n11945 ) );
BUF_X4 _u10_U597  ( .A(_u10_n11682 ), .Z(_u10_n11681 ) );
BUF_X4 _u10_U596  ( .A(_u10_n11706 ), .Z(_u10_n11705 ) );
BUF_X4 _u10_U595  ( .A(_u10_n11730 ), .Z(_u10_n11729 ) );
BUF_X4 _u10_U594  ( .A(_u10_n11778 ), .Z(_u10_n11777 ) );
BUF_X4 _u10_U593  ( .A(_u10_n11754 ), .Z(_u10_n11753 ) );
BUF_X4 _u10_U592  ( .A(_u10_n11826 ), .Z(_u10_n11825 ) );
BUF_X4 _u10_U591  ( .A(_u10_n11874 ), .Z(_u10_n11873 ) );
BUF_X4 _u10_U590  ( .A(_u10_n11850 ), .Z(_u10_n11849 ) );
BUF_X4 _u10_U589  ( .A(_u10_n11898 ), .Z(_u10_n11897 ) );
BUF_X4 _u10_U588  ( .A(_u10_n12087 ), .Z(_u10_n12086 ) );
BUF_X4 _u10_U587  ( .A(_u10_n12135 ), .Z(_u10_n12134 ) );
BUF_X4 _u10_U586  ( .A(_u10_n12111 ), .Z(_u10_n12110 ) );
BUF_X4 _u10_U585  ( .A(_u10_n12159 ), .Z(_u10_n12158 ) );
BUF_X4 _u10_U584  ( .A(_u10_n12404 ), .Z(_u10_n12020 ) );
BUF_X4 _u10_U583  ( .A(_u10_n11925 ), .Z(_u10_n11913 ) );
BUF_X4 _u10_U582  ( .A(_u10_n11973 ), .Z(_u10_n11961 ) );
BUF_X4 _u10_U581  ( .A(_u10_n11949 ), .Z(_u10_n11937 ) );
BUF_X4 _u10_U580  ( .A(_u10_n11924 ), .Z(_u10_n11914 ) );
BUF_X4 _u10_U579  ( .A(_u10_n11972 ), .Z(_u10_n11962 ) );
BUF_X4 _u10_U578  ( .A(_u10_n11948 ), .Z(_u10_n11938 ) );
BUF_X4 _u10_U577  ( .A(_u10_n11923 ), .Z(_u10_n11916 ) );
BUF_X4 _u10_U576  ( .A(_u10_n11971 ), .Z(_u10_n11964 ) );
BUF_X4 _u10_U575  ( .A(_u10_n11947 ), .Z(_u10_n11940 ) );
BUF_X4 _u10_U574  ( .A(_u10_n11923 ), .Z(_u10_n11917 ) );
BUF_X4 _u10_U573  ( .A(_u10_n11971 ), .Z(_u10_n11965 ) );
BUF_X4 _u10_U572  ( .A(_u10_n11947 ), .Z(_u10_n11941 ) );
BUF_X4 _u10_U571  ( .A(_u10_n11923 ), .Z(_u10_n11918 ) );
BUF_X4 _u10_U570  ( .A(_u10_n11971 ), .Z(_u10_n11966 ) );
BUF_X4 _u10_U569  ( .A(_u10_n11947 ), .Z(_u10_n11942 ) );
BUF_X4 _u10_U568  ( .A(_u10_n11922 ), .Z(_u10_n11919 ) );
BUF_X4 _u10_U567  ( .A(_u10_n11970 ), .Z(_u10_n11967 ) );
BUF_X4 _u10_U566  ( .A(_u10_n11946 ), .Z(_u10_n11943 ) );
BUF_X4 _u10_U565  ( .A(_u10_n11922 ), .Z(_u10_n11920 ) );
BUF_X4 _u10_U564  ( .A(_u10_n11970 ), .Z(_u10_n11968 ) );
BUF_X4 _u10_U563  ( .A(_u10_n11946 ), .Z(_u10_n11944 ) );
BUF_X4 _u10_U562  ( .A(_u10_n11926 ), .Z(_u10_n11909 ) );
BUF_X4 _u10_U561  ( .A(_u10_n11950 ), .Z(_u10_n11933 ) );
BUF_X4 _u10_U560  ( .A(_u10_n12088 ), .Z(_u10_n12078 ) );
BUF_X4 _u10_U559  ( .A(_u10_n12136 ), .Z(_u10_n12126 ) );
BUF_X4 _u10_U558  ( .A(_u10_n12112 ), .Z(_u10_n12102 ) );
BUF_X4 _u10_U557  ( .A(_u10_n12160 ), .Z(_u10_n12150 ) );
BUF_X4 _u10_U556  ( .A(_u10_n11783 ), .Z(_u10_n11761 ) );
BUF_X4 _u10_U555  ( .A(_u10_n11831 ), .Z(_u10_n11809 ) );
BUF_X4 _u10_U554  ( .A(_u10_n11879 ), .Z(_u10_n11857 ) );
BUF_X4 _u10_U553  ( .A(_u10_n11855 ), .Z(_u10_n11833 ) );
BUF_X4 _u10_U552  ( .A(_u10_n11903 ), .Z(_u10_n11881 ) );
BUF_X4 _u10_U551  ( .A(_u10_n11927 ), .Z(_u10_n11905 ) );
BUF_X4 _u10_U550  ( .A(_u10_n11975 ), .Z(_u10_n11953 ) );
BUF_X4 _u10_U549  ( .A(_u10_n11951 ), .Z(_u10_n11929 ) );
BUF_X4 _u10_U548  ( .A(_u10_n11927 ), .Z(_u10_n11906 ) );
BUF_X4 _u10_U547  ( .A(_u10_n11975 ), .Z(_u10_n11954 ) );
BUF_X4 _u10_U546  ( .A(_u10_n11951 ), .Z(_u10_n11930 ) );
BUF_X4 _u10_U545  ( .A(_u10_n12393 ), .Z(_u10_n11907 ) );
BUF_X4 _u10_U544  ( .A(_u10_n12394 ), .Z(_u10_n11931 ) );
BUF_X4 _u10_U543  ( .A(_u10_n11921 ), .Z(_u10_n11908 ) );
BUF_X4 _u10_U542  ( .A(_u10_n11945 ), .Z(_u10_n11932 ) );
BUF_X4 _u10_U541  ( .A(_u10_n12090 ), .Z(_u10_n12083 ) );
BUF_X4 _u10_U540  ( .A(_u10_n12138 ), .Z(_u10_n12131 ) );
BUF_X4 _u10_U539  ( .A(_u10_n12114 ), .Z(_u10_n12107 ) );
BUF_X4 _u10_U538  ( .A(_u10_n12160 ), .Z(_u10_n12155 ) );
BUF_X4 _u10_U537  ( .A(_u10_n11974 ), .Z(_u10_n11958 ) );
BUF_X4 _u10_U536  ( .A(_u10_n11686 ), .Z(_u10_n11671 ) );
BUF_X4 _u10_U535  ( .A(_u10_n11710 ), .Z(_u10_n11695 ) );
BUF_X4 _u10_U534  ( .A(_u10_n11734 ), .Z(_u10_n11719 ) );
BUF_X4 _u10_U533  ( .A(_u10_n11783 ), .Z(_u10_n11767 ) );
BUF_X4 _u10_U532  ( .A(_u10_n11758 ), .Z(_u10_n11743 ) );
BUF_X4 _u10_U531  ( .A(_u10_n11830 ), .Z(_u10_n11815 ) );
BUF_X4 _u10_U530  ( .A(_u10_n11876 ), .Z(_u10_n11863 ) );
BUF_X4 _u10_U529  ( .A(_u10_n11854 ), .Z(_u10_n11839 ) );
BUF_X4 _u10_U528  ( .A(_u10_n11902 ), .Z(_u10_n11887 ) );
BUF_X4 _u10_U527  ( .A(_u10_n11974 ), .Z(_u10_n11959 ) );
BUF_X4 _u10_U526  ( .A(_u10_n11974 ), .Z(_u10_n11960 ) );
BUF_X4 _u10_U525  ( .A(_u10_n11687 ), .Z(_u10_n11667 ) );
BUF_X4 _u10_U524  ( .A(_u10_n11735 ), .Z(_u10_n11715 ) );
BUF_X4 _u10_U523  ( .A(_u10_n11759 ), .Z(_u10_n11739 ) );
BUF_X4 _u10_U522  ( .A(_u10_n11827 ), .Z(_u10_n11813 ) );
BUF_X4 _u10_U521  ( .A(_u10_n11878 ), .Z(_u10_n11859 ) );
BUF_X4 _u10_U520  ( .A(_u10_n11855 ), .Z(_u10_n11835 ) );
BUF_X4 _u10_U519  ( .A(_u10_n11926 ), .Z(_u10_n11910 ) );
BUF_X4 _u10_U518  ( .A(_u10_n11974 ), .Z(_u10_n11955 ) );
BUF_X4 _u10_U517  ( .A(_u10_n11950 ), .Z(_u10_n11934 ) );
BUF_X4 _u10_U516  ( .A(_u10_n11684 ), .Z(_u10_n11666 ) );
BUF_X4 _u10_U515  ( .A(_u10_n11708 ), .Z(_u10_n11690 ) );
BUF_X4 _u10_U514  ( .A(_u10_n11732 ), .Z(_u10_n11714 ) );
BUF_X4 _u10_U513  ( .A(_u10_n11783 ), .Z(_u10_n11765 ) );
BUF_X4 _u10_U512  ( .A(_u10_n11756 ), .Z(_u10_n11738 ) );
BUF_X4 _u10_U511  ( .A(_u10_n12088 ), .Z(_u10_n12082 ) );
BUF_X4 _u10_U510  ( .A(_u10_n12136 ), .Z(_u10_n12130 ) );
BUF_X4 _u10_U509  ( .A(_u10_n12112 ), .Z(_u10_n12106 ) );
BUF_X4 _u10_U508  ( .A(_u10_n11682 ), .Z(_u10_n11680 ) );
BUF_X4 _u10_U507  ( .A(_u10_n11706 ), .Z(_u10_n11704 ) );
BUF_X4 _u10_U506  ( .A(_u10_n11730 ), .Z(_u10_n11728 ) );
BUF_X4 _u10_U505  ( .A(_u10_n11778 ), .Z(_u10_n11776 ) );
BUF_X4 _u10_U504  ( .A(_u10_n11754 ), .Z(_u10_n11752 ) );
BUF_X4 _u10_U503  ( .A(_u10_n11826 ), .Z(_u10_n11824 ) );
BUF_X4 _u10_U502  ( .A(_u10_n11874 ), .Z(_u10_n11872 ) );
BUF_X4 _u10_U501  ( .A(_u10_n11850 ), .Z(_u10_n11848 ) );
BUF_X4 _u10_U500  ( .A(_u10_n11898 ), .Z(_u10_n11896 ) );
BUF_X4 _u10_U499  ( .A(_u10_n12089 ), .Z(_u10_n12076 ) );
BUF_X4 _u10_U498  ( .A(_u10_n12137 ), .Z(_u10_n12124 ) );
BUF_X4 _u10_U497  ( .A(_u10_n12113 ), .Z(_u10_n12100 ) );
BUF_X4 _u10_U496  ( .A(_u10_n12161 ), .Z(_u10_n12148 ) );
BUF_X4 _u10_U495  ( .A(_u10_n11684 ), .Z(_u10_n11675 ) );
BUF_X4 _u10_U494  ( .A(_u10_n11708 ), .Z(_u10_n11699 ) );
BUF_X4 _u10_U493  ( .A(_u10_n11732 ), .Z(_u10_n11723 ) );
BUF_X4 _u10_U492  ( .A(_u10_n11780 ), .Z(_u10_n11771 ) );
BUF_X4 _u10_U491  ( .A(_u10_n11756 ), .Z(_u10_n11747 ) );
BUF_X4 _u10_U490  ( .A(_u10_n11828 ), .Z(_u10_n11819 ) );
BUF_X4 _u10_U489  ( .A(_u10_n11876 ), .Z(_u10_n11867 ) );
BUF_X4 _u10_U488  ( .A(_u10_n11852 ), .Z(_u10_n11843 ) );
BUF_X4 _u10_U487  ( .A(_u10_n11900 ), .Z(_u10_n11891 ) );
BUF_X4 _u10_U486  ( .A(_u10_n11924 ), .Z(_u10_n11915 ) );
BUF_X4 _u10_U485  ( .A(_u10_n11972 ), .Z(_u10_n11963 ) );
BUF_X4 _u10_U484  ( .A(_u10_n11948 ), .Z(_u10_n11939 ) );
BUF_X4 _u10_U483  ( .A(_u10_n12091 ), .Z(_u10_n12071 ) );
BUF_X4 _u10_U482  ( .A(_u10_n12139 ), .Z(_u10_n12119 ) );
BUF_X4 _u10_U481  ( .A(_u10_n12115 ), .Z(_u10_n12095 ) );
BUF_X4 _u10_U480  ( .A(_u10_n12163 ), .Z(_u10_n12143 ) );
BUF_X4 _u10_U479  ( .A(_u10_n11683 ), .Z(_u10_n11677 ) );
BUF_X4 _u10_U478  ( .A(_u10_n11707 ), .Z(_u10_n11701 ) );
BUF_X4 _u10_U477  ( .A(_u10_n11731 ), .Z(_u10_n11725 ) );
BUF_X4 _u10_U476  ( .A(_u10_n11779 ), .Z(_u10_n11773 ) );
BUF_X4 _u10_U475  ( .A(_u10_n11755 ), .Z(_u10_n11749 ) );
BUF_X4 _u10_U474  ( .A(_u10_n11827 ), .Z(_u10_n11821 ) );
BUF_X4 _u10_U473  ( .A(_u10_n11875 ), .Z(_u10_n11869 ) );
BUF_X4 _u10_U472  ( .A(_u10_n11851 ), .Z(_u10_n11845 ) );
BUF_X4 _u10_U471  ( .A(_u10_n11899 ), .Z(_u10_n11893 ) );
BUF_X4 _u10_U470  ( .A(_u10_n12090 ), .Z(_u10_n12074 ) );
BUF_X4 _u10_U469  ( .A(_u10_n12138 ), .Z(_u10_n12122 ) );
BUF_X4 _u10_U468  ( .A(_u10_n12114 ), .Z(_u10_n12098 ) );
BUF_X4 _u10_U467  ( .A(_u10_n12162 ), .Z(_u10_n12146 ) );
BUF_X4 _u10_U466  ( .A(_u10_n11685 ), .Z(_u10_n11672 ) );
BUF_X4 _u10_U465  ( .A(_u10_n11709 ), .Z(_u10_n11696 ) );
BUF_X4 _u10_U464  ( .A(_u10_n11733 ), .Z(_u10_n11720 ) );
BUF_X4 _u10_U463  ( .A(_u10_n11781 ), .Z(_u10_n11768 ) );
BUF_X4 _u10_U462  ( .A(_u10_n11757 ), .Z(_u10_n11744 ) );
BUF_X4 _u10_U461  ( .A(_u10_n11829 ), .Z(_u10_n11816 ) );
BUF_X4 _u10_U460  ( .A(_u10_n11877 ), .Z(_u10_n11864 ) );
BUF_X4 _u10_U459  ( .A(_u10_n11853 ), .Z(_u10_n11840 ) );
BUF_X4 _u10_U458  ( .A(_u10_n11901 ), .Z(_u10_n11888 ) );
BUF_X4 _u10_U457  ( .A(_u10_n12087 ), .Z(_u10_n12084 ) );
BUF_X4 _u10_U456  ( .A(_u10_n12135 ), .Z(_u10_n12132 ) );
BUF_X4 _u10_U455  ( .A(_u10_n12111 ), .Z(_u10_n12108 ) );
BUF_X4 _u10_U454  ( .A(_u10_n12159 ), .Z(_u10_n12156 ) );
BUF_X4 _u10_U453  ( .A(_u10_n11686 ), .Z(_u10_n11670 ) );
BUF_X4 _u10_U452  ( .A(_u10_n11710 ), .Z(_u10_n11694 ) );
BUF_X4 _u10_U451  ( .A(_u10_n11734 ), .Z(_u10_n11718 ) );
BUF_X4 _u10_U450  ( .A(_u10_n11758 ), .Z(_u10_n11742 ) );
BUF_X4 _u10_U449  ( .A(_u10_n11830 ), .Z(_u10_n11814 ) );
BUF_X4 _u10_U448  ( .A(_u10_n11877 ), .Z(_u10_n11862 ) );
BUF_X4 _u10_U447  ( .A(_u10_n11854 ), .Z(_u10_n11838 ) );
BUF_X4 _u10_U446  ( .A(_u10_n11902 ), .Z(_u10_n11886 ) );
BUF_X4 _u10_U445  ( .A(_u10_n12090 ), .Z(_u10_n12073 ) );
BUF_X4 _u10_U444  ( .A(_u10_n12138 ), .Z(_u10_n12121 ) );
BUF_X4 _u10_U443  ( .A(_u10_n12114 ), .Z(_u10_n12097 ) );
BUF_X4 _u10_U442  ( .A(_u10_n12162 ), .Z(_u10_n12145 ) );
BUF_X4 _u10_U441  ( .A(_u10_n11683 ), .Z(_u10_n11676 ) );
BUF_X4 _u10_U440  ( .A(_u10_n11707 ), .Z(_u10_n11700 ) );
BUF_X4 _u10_U439  ( .A(_u10_n11731 ), .Z(_u10_n11724 ) );
BUF_X4 _u10_U438  ( .A(_u10_n11779 ), .Z(_u10_n11772 ) );
BUF_X4 _u10_U437  ( .A(_u10_n11755 ), .Z(_u10_n11748 ) );
BUF_X4 _u10_U436  ( .A(_u10_n11827 ), .Z(_u10_n11820 ) );
BUF_X4 _u10_U435  ( .A(_u10_n11875 ), .Z(_u10_n11868 ) );
BUF_X4 _u10_U434  ( .A(_u10_n11851 ), .Z(_u10_n11844 ) );
BUF_X4 _u10_U433  ( .A(_u10_n11899 ), .Z(_u10_n11892 ) );
BUF_X4 _u10_U432  ( .A(_u10_n12090 ), .Z(_u10_n12072 ) );
BUF_X4 _u10_U431  ( .A(_u10_n12138 ), .Z(_u10_n12120 ) );
BUF_X4 _u10_U430  ( .A(_u10_n12114 ), .Z(_u10_n12096 ) );
BUF_X4 _u10_U429  ( .A(_u10_n12162 ), .Z(_u10_n12144 ) );
BUF_X4 _u10_U428  ( .A(_u10_n11683 ), .Z(_u10_n11678 ) );
BUF_X4 _u10_U427  ( .A(_u10_n11707 ), .Z(_u10_n11702 ) );
BUF_X4 _u10_U426  ( .A(_u10_n11731 ), .Z(_u10_n11726 ) );
BUF_X4 _u10_U425  ( .A(_u10_n11779 ), .Z(_u10_n11774 ) );
BUF_X4 _u10_U424  ( .A(_u10_n11755 ), .Z(_u10_n11750 ) );
BUF_X4 _u10_U423  ( .A(_u10_n11827 ), .Z(_u10_n11822 ) );
BUF_X4 _u10_U422  ( .A(_u10_n11875 ), .Z(_u10_n11870 ) );
BUF_X4 _u10_U421  ( .A(_u10_n11851 ), .Z(_u10_n11846 ) );
BUF_X4 _u10_U420  ( .A(_u10_n11899 ), .Z(_u10_n11894 ) );
BUF_X4 _u10_U419  ( .A(_u10_n11685 ), .Z(_u10_n11673 ) );
BUF_X4 _u10_U418  ( .A(_u10_n11709 ), .Z(_u10_n11697 ) );
BUF_X4 _u10_U417  ( .A(_u10_n11733 ), .Z(_u10_n11721 ) );
BUF_X4 _u10_U416  ( .A(_u10_n11781 ), .Z(_u10_n11769 ) );
BUF_X4 _u10_U415  ( .A(_u10_n11757 ), .Z(_u10_n11745 ) );
BUF_X4 _u10_U414  ( .A(_u10_n11829 ), .Z(_u10_n11817 ) );
BUF_X4 _u10_U413  ( .A(_u10_n11877 ), .Z(_u10_n11865 ) );
BUF_X4 _u10_U412  ( .A(_u10_n11853 ), .Z(_u10_n11841 ) );
BUF_X4 _u10_U411  ( .A(_u10_n11901 ), .Z(_u10_n11889 ) );
BUF_X4 _u10_U410  ( .A(_u10_n12091 ), .Z(_u10_n12070 ) );
BUF_X4 _u10_U409  ( .A(_u10_n12139 ), .Z(_u10_n12118 ) );
BUF_X4 _u10_U408  ( .A(_u10_n12115 ), .Z(_u10_n12094 ) );
BUF_X4 _u10_U407  ( .A(_u10_n12163 ), .Z(_u10_n12142 ) );
BUF_X4 _u10_U406  ( .A(_u10_n11682 ), .Z(_u10_n11679 ) );
BUF_X4 _u10_U405  ( .A(_u10_n11706 ), .Z(_u10_n11703 ) );
BUF_X4 _u10_U404  ( .A(_u10_n11730 ), .Z(_u10_n11727 ) );
BUF_X4 _u10_U403  ( .A(_u10_n11778 ), .Z(_u10_n11775 ) );
BUF_X4 _u10_U402  ( .A(_u10_n11754 ), .Z(_u10_n11751 ) );
BUF_X4 _u10_U401  ( .A(_u10_n11826 ), .Z(_u10_n11823 ) );
BUF_X4 _u10_U400  ( .A(_u10_n11874 ), .Z(_u10_n11871 ) );
BUF_X4 _u10_U399  ( .A(_u10_n11850 ), .Z(_u10_n11847 ) );
BUF_X4 _u10_U398  ( .A(_u10_n11898 ), .Z(_u10_n11895 ) );
BUF_X4 _u10_U397  ( .A(_u10_n11684 ), .Z(_u10_n11674 ) );
BUF_X4 _u10_U396  ( .A(_u10_n11708 ), .Z(_u10_n11698 ) );
BUF_X4 _u10_U395  ( .A(_u10_n11732 ), .Z(_u10_n11722 ) );
BUF_X4 _u10_U394  ( .A(_u10_n11780 ), .Z(_u10_n11770 ) );
BUF_X4 _u10_U393  ( .A(_u10_n11756 ), .Z(_u10_n11746 ) );
BUF_X4 _u10_U392  ( .A(_u10_n11828 ), .Z(_u10_n11818 ) );
BUF_X4 _u10_U391  ( .A(_u10_n11876 ), .Z(_u10_n11866 ) );
BUF_X4 _u10_U390  ( .A(_u10_n11852 ), .Z(_u10_n11842 ) );
BUF_X4 _u10_U389  ( .A(_u10_n11900 ), .Z(_u10_n11890 ) );
BUF_X4 _u10_U388  ( .A(_u10_n12089 ), .Z(_u10_n12075 ) );
BUF_X4 _u10_U387  ( .A(_u10_n12137 ), .Z(_u10_n12123 ) );
BUF_X4 _u10_U386  ( .A(_u10_n12113 ), .Z(_u10_n12099 ) );
BUF_X4 _u10_U385  ( .A(_u10_n12161 ), .Z(_u10_n12147 ) );
BUF_X4 _u10_U384  ( .A(_u10_n12091 ), .Z(_u10_n12069 ) );
BUF_X4 _u10_U383  ( .A(_u10_n12139 ), .Z(_u10_n12117 ) );
BUF_X4 _u10_U382  ( .A(_u10_n12115 ), .Z(_u10_n12093 ) );
BUF_X4 _u10_U381  ( .A(_u10_n12163 ), .Z(_u10_n12141 ) );
BUF_X4 _u10_U380  ( .A(_u10_n12089 ), .Z(_u10_n12077 ) );
BUF_X4 _u10_U379  ( .A(_u10_n12137 ), .Z(_u10_n12125 ) );
BUF_X4 _u10_U378  ( .A(_u10_n12113 ), .Z(_u10_n12101 ) );
BUF_X4 _u10_U377  ( .A(_u10_n11687 ), .Z(_u10_n11669 ) );
BUF_X4 _u10_U376  ( .A(_u10_n11711 ), .Z(_u10_n11693 ) );
BUF_X4 _u10_U375  ( .A(_u10_n11735 ), .Z(_u10_n11717 ) );
BUF_X4 _u10_U374  ( .A(_u10_n11759 ), .Z(_u10_n11741 ) );
BUF_X4 _u10_U373  ( .A(_u10_n11878 ), .Z(_u10_n11861 ) );
BUF_X4 _u10_U372  ( .A(_u10_n12386 ), .Z(_u10_n11837 ) );
BUF_X4 _u10_U371  ( .A(_u10_n11899 ), .Z(_u10_n11885 ) );
BUF_X4 _u10_U370  ( .A(_u10_n11926 ), .Z(_u10_n11912 ) );
BUF_X4 _u10_U369  ( .A(_u10_n12395 ), .Z(_u10_n11957 ) );
BUF_X4 _u10_U368  ( .A(_u10_n11950 ), .Z(_u10_n11936 ) );
BUF_X4 _u10_U367  ( .A(_u10_n12087 ), .Z(_u10_n12085 ) );
BUF_X4 _u10_U366  ( .A(_u10_n12135 ), .Z(_u10_n12133 ) );
BUF_X4 _u10_U365  ( .A(_u10_n12111 ), .Z(_u10_n12109 ) );
BUF_X4 _u10_U364  ( .A(_u10_n12159 ), .Z(_u10_n12157 ) );
BUF_X4 _u10_U363  ( .A(_u10_n12414 ), .Z(_u10_n12154 ) );
BUF_X4 _u10_U362  ( .A(_u10_n11687 ), .Z(_u10_n11668 ) );
BUF_X4 _u10_U361  ( .A(_u10_n11711 ), .Z(_u10_n11692 ) );
BUF_X4 _u10_U360  ( .A(_u10_n11735 ), .Z(_u10_n11716 ) );
BUF_X4 _u10_U359  ( .A(_u10_n11782 ), .Z(_u10_n11766 ) );
BUF_X4 _u10_U358  ( .A(_u10_n11759 ), .Z(_u10_n11740 ) );
BUF_X4 _u10_U357  ( .A(_u10_n11878 ), .Z(_u10_n11860 ) );
BUF_X4 _u10_U356  ( .A(_u10_n11849 ), .Z(_u10_n11836 ) );
BUF_X4 _u10_U355  ( .A(_u10_n11926 ), .Z(_u10_n11911 ) );
BUF_X4 _u10_U354  ( .A(_u10_n11969 ), .Z(_u10_n11956 ) );
BUF_X4 _u10_U353  ( .A(_u10_n11950 ), .Z(_u10_n11935 ) );
BUF_X4 _u10_U352  ( .A(_u10_n12371 ), .Z(_u10_n11665 ) );
BUF_X4 _u10_U351  ( .A(_u10_n12372 ), .Z(_u10_n11689 ) );
BUF_X4 _u10_U350  ( .A(_u10_n12377 ), .Z(_u10_n11713 ) );
BUF_X4 _u10_U349  ( .A(_u10_n11783 ), .Z(_u10_n11764 ) );
BUF_X4 _u10_U348  ( .A(_u10_n12378 ), .Z(_u10_n11737 ) );
BUF_X4 _u10_U347  ( .A(_u10_n11831 ), .Z(_u10_n11812 ) );
BUF_X4 _u10_U346  ( .A(_u10_n11903 ), .Z(_u10_n11884 ) );
BUF_X4 _u10_U345  ( .A(_u10_n12164 ), .Z(_u10_n12153 ) );
BUF_X4 _u10_U344  ( .A(_u10_n12088 ), .Z(_u10_n12081 ) );
BUF_X4 _u10_U343  ( .A(_u10_n12136 ), .Z(_u10_n12129 ) );
BUF_X4 _u10_U342  ( .A(_u10_n12112 ), .Z(_u10_n12105 ) );
BUF_X4 _u10_U341  ( .A(_u10_n11711 ), .Z(_u10_n11691 ) );
BUF_X4 _u10_U340  ( .A(_u10_n11681 ), .Z(_u10_n11664 ) );
BUF_X4 _u10_U339  ( .A(_u10_n11705 ), .Z(_u10_n11688 ) );
BUF_X4 _u10_U338  ( .A(_u10_n11729 ), .Z(_u10_n11712 ) );
BUF_X4 _u10_U337  ( .A(_u10_n11783 ), .Z(_u10_n11763 ) );
BUF_X4 _u10_U336  ( .A(_u10_n11753 ), .Z(_u10_n11736 ) );
BUF_X4 _u10_U335  ( .A(_u10_n11831 ), .Z(_u10_n11811 ) );
BUF_X4 _u10_U334  ( .A(_u10_n11903 ), .Z(_u10_n11883 ) );
BUF_X4 _u10_U333  ( .A(_u10_n12411 ), .Z(_u10_n12080 ) );
BUF_X4 _u10_U332  ( .A(_u10_n12413 ), .Z(_u10_n12128 ) );
BUF_X4 _u10_U331  ( .A(_u10_n12412 ), .Z(_u10_n12104 ) );
BUF_X4 _u10_U330  ( .A(_u10_n12160 ), .Z(_u10_n12152 ) );
BUF_X4 _u10_U329  ( .A(_u10_n12379 ), .Z(_u10_n11762 ) );
BUF_X4 _u10_U328  ( .A(_u10_n12385 ), .Z(_u10_n11810 ) );
BUF_X4 _u10_U327  ( .A(_u10_n12387 ), .Z(_u10_n11858 ) );
BUF_X4 _u10_U326  ( .A(_u10_n11855 ), .Z(_u10_n11834 ) );
BUF_X4 _u10_U325  ( .A(_u10_n12092 ), .Z(_u10_n12079 ) );
BUF_X4 _u10_U324  ( .A(_u10_n12140 ), .Z(_u10_n12127 ) );
BUF_X4 _u10_U323  ( .A(_u10_n12116 ), .Z(_u10_n12103 ) );
BUF_X4 _u10_U322  ( .A(_u10_n12160 ), .Z(_u10_n12151 ) );
BUF_X4 _u10_U321  ( .A(_u10_n12388 ), .Z(_u10_n11882 ) );
BUF_X4 _u10_U320  ( .A(_u10_n12161 ), .Z(_u10_n12149 ) );
BUF_X4 _u10_U319  ( .A(_u10_n11927 ), .Z(_u10_n11904 ) );
BUF_X4 _u10_U318  ( .A(_u10_n11975 ), .Z(_u10_n11952 ) );
BUF_X4 _u10_U317  ( .A(_u10_n11951 ), .Z(_u10_n11928 ) );
BUF_X4 _u10_U316  ( .A(_u10_n11777 ), .Z(_u10_n11760 ) );
BUF_X4 _u10_U315  ( .A(_u10_n11825 ), .Z(_u10_n11808 ) );
BUF_X4 _u10_U314  ( .A(_u10_n11873 ), .Z(_u10_n11856 ) );
BUF_X4 _u10_U313  ( .A(_u10_n11855 ), .Z(_u10_n11832 ) );
BUF_X4 _u10_U312  ( .A(_u10_n11897 ), .Z(_u10_n11880 ) );
BUF_X4 _u10_U311  ( .A(_u10_n12404 ), .Z(_u10_n12008 ) );
BUF_X4 _u10_U310  ( .A(_u10_n12404 ), .Z(_u10_n12009 ) );
BUF_X4 _u10_U309  ( .A(_u10_n12404 ), .Z(_u10_n12010 ) );
BUF_X4 _u10_U308  ( .A(_u10_n12404 ), .Z(_u10_n12016 ) );
BUF_X4 _u10_U307  ( .A(_u10_n12404 ), .Z(_u10_n12015 ) );
BUF_X4 _u10_U306  ( .A(_u10_n12404 ), .Z(_u10_n12003 ) );
BUF_X4 _u10_U305  ( .A(_u10_n12404 ), .Z(_u10_n12006 ) );
BUF_X4 _u10_U304  ( .A(_u10_n12404 ), .Z(_u10_n12001 ) );
BUF_X4 _u10_U303  ( .A(_u10_n12404 ), .Z(_u10_n12018 ) );
BUF_X4 _u10_U302  ( .A(_u10_n12404 ), .Z(_u10_n12019 ) );
BUF_X4 _u10_U301  ( .A(_u10_n12404 ), .Z(_u10_n12005 ) );
BUF_X4 _u10_U300  ( .A(_u10_n12404 ), .Z(_u10_n12004 ) );
BUF_X4 _u10_U299  ( .A(_u10_n12404 ), .Z(_u10_n12007 ) );
BUF_X4 _u10_U298  ( .A(_u10_n12404 ), .Z(_u10_n12002 ) );
BUF_X4 _u10_U297  ( .A(_u10_n12404 ), .Z(_u10_n12017 ) );
BUF_X4 _u10_U296  ( .A(_u10_n12404 ), .Z(_u10_n12014 ) );
BUF_X4 _u10_U295  ( .A(_u10_n12404 ), .Z(_u10_n12013 ) );
BUF_X4 _u10_U294  ( .A(_u10_n12404 ), .Z(_u10_n12012 ) );
BUF_X4 _u10_U293  ( .A(_u10_n12404 ), .Z(_u10_n12011 ) );
BUF_X4 _u10_U292  ( .A(_u10_n12404 ), .Z(_u10_n12000 ) );
BUF_X4 _u10_U291  ( .A(_u10_n12039 ), .Z(_u10_n12038 ) );
BUF_X4 _u10_U290  ( .A(_u10_n12063 ), .Z(_u10_n12062 ) );
BUF_X4 _u10_U289  ( .A(_u10_n12185 ), .Z(_u10_n12184 ) );
BUF_X4 _u10_U288  ( .A(_u10_n12233 ), .Z(_u10_n12232 ) );
BUF_X4 _u10_U287  ( .A(_u10_n12207 ), .Z(_u10_n12206 ) );
BUF_X4 _u10_U286  ( .A(_u10_n12257 ), .Z(_u10_n12256 ) );
BUF_X4 _u10_U285  ( .A(_u10_n12353 ), .Z(_u10_n12352 ) );
BUF_X4 _u10_U284  ( .A(_u10_n12283 ), .Z(_u10_n12261 ) );
BUF_X4 _u10_U283  ( .A(_u10_n12331 ), .Z(_u10_n12309 ) );
BUF_X4 _u10_U282  ( .A(_u10_n12307 ), .Z(_u10_n12285 ) );
BUF_X4 _u10_U281  ( .A(_u10_n12283 ), .Z(_u10_n12263 ) );
BUF_X4 _u10_U280  ( .A(_u10_n12331 ), .Z(_u10_n12311 ) );
BUF_X4 _u10_U279  ( .A(_u10_n12307 ), .Z(_u10_n12287 ) );
BUF_X4 _u10_U278  ( .A(_u10_n12282 ), .Z(_u10_n12264 ) );
BUF_X4 _u10_U277  ( .A(_u10_n12330 ), .Z(_u10_n12312 ) );
BUF_X4 _u10_U276  ( .A(_u10_n12306 ), .Z(_u10_n12288 ) );
BUF_X4 _u10_U275  ( .A(_u10_n12282 ), .Z(_u10_n12265 ) );
BUF_X4 _u10_U274  ( .A(_u10_n12330 ), .Z(_u10_n12313 ) );
BUF_X4 _u10_U273  ( .A(_u10_n12306 ), .Z(_u10_n12289 ) );
BUF_X4 _u10_U272  ( .A(_u10_n12282 ), .Z(_u10_n12266 ) );
BUF_X4 _u10_U271  ( .A(_u10_n12330 ), .Z(_u10_n12314 ) );
BUF_X4 _u10_U270  ( .A(_u10_n12306 ), .Z(_u10_n12290 ) );
BUF_X4 _u10_U269  ( .A(_u10_n12281 ), .Z(_u10_n12267 ) );
BUF_X4 _u10_U268  ( .A(_u10_n12329 ), .Z(_u10_n12315 ) );
BUF_X4 _u10_U267  ( .A(_u10_n12305 ), .Z(_u10_n12291 ) );
BUF_X4 _u10_U266  ( .A(_u10_n12281 ), .Z(_u10_n12268 ) );
BUF_X4 _u10_U265  ( .A(_u10_n12305 ), .Z(_u10_n12292 ) );
BUF_X4 _u10_U264  ( .A(_u10_n12281 ), .Z(_u10_n12269 ) );
BUF_X4 _u10_U263  ( .A(_u10_n12329 ), .Z(_u10_n12316 ) );
BUF_X4 _u10_U262  ( .A(_u10_n12305 ), .Z(_u10_n12293 ) );
BUF_X4 _u10_U261  ( .A(_u10_n12405 ), .Z(_u10_n12030 ) );
BUF_X4 _u10_U260  ( .A(_u10_n12406 ), .Z(_u10_n12054 ) );
BUF_X4 _u10_U259  ( .A(_u10_n12188 ), .Z(_u10_n12173 ) );
BUF_X4 _u10_U258  ( .A(_u10_n12236 ), .Z(_u10_n12221 ) );
BUF_X4 _u10_U257  ( .A(_u10_n12260 ), .Z(_u10_n12245 ) );
BUF_X4 _u10_U256  ( .A(_u10_n12280 ), .Z(_u10_n12270 ) );
BUF_X4 _u10_U255  ( .A(_u10_n12328 ), .Z(_u10_n12317 ) );
BUF_X4 _u10_U254  ( .A(_u10_n12304 ), .Z(_u10_n12294 ) );
BUF_X4 _u10_U253  ( .A(_u10_n12356 ), .Z(_u10_n12341 ) );
BUF_X4 _u10_U252  ( .A(_u10_n12280 ), .Z(_u10_n12271 ) );
BUF_X4 _u10_U251  ( .A(_u10_n12328 ), .Z(_u10_n12318 ) );
BUF_X4 _u10_U250  ( .A(_u10_n12304 ), .Z(_u10_n12295 ) );
BUF_X4 _u10_U249  ( .A(_u10_n12280 ), .Z(_u10_n12272 ) );
BUF_X4 _u10_U248  ( .A(_u10_n12328 ), .Z(_u10_n12319 ) );
BUF_X4 _u10_U247  ( .A(_u10_n12304 ), .Z(_u10_n12296 ) );
BUF_X4 _u10_U246  ( .A(_u10_n12427 ), .Z(_u10_n12273 ) );
BUF_X4 _u10_U245  ( .A(_u10_n12328 ), .Z(_u10_n12320 ) );
BUF_X4 _u10_U244  ( .A(_u10_n12428 ), .Z(_u10_n12297 ) );
BUF_X4 _u10_U243  ( .A(_u10_n12284 ), .Z(_u10_n12274 ) );
BUF_X4 _u10_U242  ( .A(_u10_n12429 ), .Z(_u10_n12321 ) );
BUF_X4 _u10_U241  ( .A(_u10_n12308 ), .Z(_u10_n12298 ) );
BUF_X4 _u10_U240  ( .A(_u10_n12279 ), .Z(_u10_n12278 ) );
BUF_X4 _u10_U239  ( .A(_u10_n12332 ), .Z(_u10_n12325 ) );
BUF_X4 _u10_U238  ( .A(_u10_n12303 ), .Z(_u10_n12302 ) );
BUF_X4 _u10_U237  ( .A(_u10_n12330 ), .Z(_u10_n12326 ) );
BUF_X4 _u10_U236  ( .A(_u10_n12329 ), .Z(_u10_n12327 ) );
BUF_X4 _u10_U235  ( .A(_u10_n12044 ), .Z(_u10_n12033 ) );
BUF_X4 _u10_U234  ( .A(_u10_n12068 ), .Z(_u10_n12057 ) );
BUF_X4 _u10_U233  ( .A(_u10_n12419 ), .Z(_u10_n12179 ) );
BUF_X4 _u10_U232  ( .A(_u10_n12421 ), .Z(_u10_n12227 ) );
BUF_X4 _u10_U231  ( .A(_u10_n12420 ), .Z(_u10_n12201 ) );
BUF_X4 _u10_U230  ( .A(_u10_n12279 ), .Z(_u10_n12276 ) );
BUF_X4 _u10_U229  ( .A(_u10_n12331 ), .Z(_u10_n12323 ) );
BUF_X4 _u10_U228  ( .A(_u10_n12303 ), .Z(_u10_n12300 ) );
BUF_X4 _u10_U227  ( .A(_u10_n12188 ), .Z(_u10_n12178 ) );
BUF_X4 _u10_U226  ( .A(_u10_n12236 ), .Z(_u10_n12226 ) );
BUF_X4 _u10_U225  ( .A(_u10_n12206 ), .Z(_u10_n12200 ) );
BUF_X4 _u10_U224  ( .A(_u10_n12280 ), .Z(_u10_n12275 ) );
BUF_X4 _u10_U223  ( .A(_u10_n12331 ), .Z(_u10_n12322 ) );
BUF_X4 _u10_U222  ( .A(_u10_n12304 ), .Z(_u10_n12299 ) );
BUF_X4 _u10_U221  ( .A(_u10_n12041 ), .Z(_u10_n12028 ) );
BUF_X4 _u10_U220  ( .A(_u10_n12065 ), .Z(_u10_n12052 ) );
BUF_X4 _u10_U219  ( .A(_u10_n12186 ), .Z(_u10_n12171 ) );
BUF_X4 _u10_U218  ( .A(_u10_n12234 ), .Z(_u10_n12219 ) );
BUF_X4 _u10_U217  ( .A(_u10_n12209 ), .Z(_u10_n12196 ) );
BUF_X4 _u10_U216  ( .A(_u10_n12258 ), .Z(_u10_n12243 ) );
BUF_X4 _u10_U215  ( .A(_u10_n12354 ), .Z(_u10_n12339 ) );
BUF_X4 _u10_U214  ( .A(_u10_n12043 ), .Z(_u10_n12023 ) );
BUF_X4 _u10_U213  ( .A(_u10_n12067 ), .Z(_u10_n12047 ) );
BUF_X4 _u10_U212  ( .A(_u10_n12187 ), .Z(_u10_n12167 ) );
BUF_X4 _u10_U211  ( .A(_u10_n12235 ), .Z(_u10_n12215 ) );
BUF_X4 _u10_U210  ( .A(_u10_n12211 ), .Z(_u10_n12191 ) );
BUF_X4 _u10_U209  ( .A(_u10_n12259 ), .Z(_u10_n12239 ) );
BUF_X4 _u10_U208  ( .A(_u10_n12355 ), .Z(_u10_n12335 ) );
BUF_X4 _u10_U207  ( .A(_u10_n12042 ), .Z(_u10_n12026 ) );
BUF_X4 _u10_U206  ( .A(_u10_n12066 ), .Z(_u10_n12050 ) );
BUF_X4 _u10_U205  ( .A(_u10_n12188 ), .Z(_u10_n12169 ) );
BUF_X4 _u10_U204  ( .A(_u10_n12236 ), .Z(_u10_n12217 ) );
BUF_X4 _u10_U203  ( .A(_u10_n12210 ), .Z(_u10_n12194 ) );
BUF_X4 _u10_U202  ( .A(_u10_n12260 ), .Z(_u10_n12241 ) );
BUF_X4 _u10_U201  ( .A(_u10_n12356 ), .Z(_u10_n12337 ) );
BUF_X4 _u10_U200  ( .A(_u10_n12039 ), .Z(_u10_n12036 ) );
BUF_X4 _u10_U199  ( .A(_u10_n12063 ), .Z(_u10_n12060 ) );
BUF_X4 _u10_U198  ( .A(_u10_n12185 ), .Z(_u10_n12182 ) );
BUF_X4 _u10_U197  ( .A(_u10_n12233 ), .Z(_u10_n12230 ) );
BUF_X4 _u10_U196  ( .A(_u10_n12207 ), .Z(_u10_n12204 ) );
BUF_X4 _u10_U195  ( .A(_u10_n12257 ), .Z(_u10_n12254 ) );
BUF_X4 _u10_U194  ( .A(_u10_n12353 ), .Z(_u10_n12350 ) );
BUF_X4 _u10_U193  ( .A(_u10_n12042 ), .Z(_u10_n12025 ) );
BUF_X4 _u10_U192  ( .A(_u10_n12066 ), .Z(_u10_n12049 ) );
BUF_X4 _u10_U191  ( .A(_u10_n12186 ), .Z(_u10_n12168 ) );
BUF_X4 _u10_U190  ( .A(_u10_n12234 ), .Z(_u10_n12216 ) );
BUF_X4 _u10_U189  ( .A(_u10_n12210 ), .Z(_u10_n12193 ) );
BUF_X4 _u10_U188  ( .A(_u10_n12258 ), .Z(_u10_n12240 ) );
BUF_X4 _u10_U187  ( .A(_u10_n12354 ), .Z(_u10_n12336 ) );
BUF_X4 _u10_U186  ( .A(_u10_n12042 ), .Z(_u10_n12024 ) );
BUF_X4 _u10_U185  ( .A(_u10_n12066 ), .Z(_u10_n12048 ) );
BUF_X4 _u10_U184  ( .A(_u10_n12210 ), .Z(_u10_n12192 ) );
BUF_X4 _u10_U183  ( .A(_u10_n12043 ), .Z(_u10_n12022 ) );
BUF_X4 _u10_U182  ( .A(_u10_n12067 ), .Z(_u10_n12046 ) );
BUF_X4 _u10_U181  ( .A(_u10_n12187 ), .Z(_u10_n12166 ) );
BUF_X4 _u10_U180  ( .A(_u10_n12235 ), .Z(_u10_n12214 ) );
BUF_X4 _u10_U179  ( .A(_u10_n12211 ), .Z(_u10_n12190 ) );
BUF_X4 _u10_U178  ( .A(_u10_n12259 ), .Z(_u10_n12238 ) );
BUF_X4 _u10_U177  ( .A(_u10_n12283 ), .Z(_u10_n12262 ) );
BUF_X4 _u10_U176  ( .A(_u10_n12331 ), .Z(_u10_n12310 ) );
BUF_X4 _u10_U175  ( .A(_u10_n12307 ), .Z(_u10_n12286 ) );
BUF_X4 _u10_U174  ( .A(_u10_n12355 ), .Z(_u10_n12334 ) );
BUF_X4 _u10_U173  ( .A(_u10_n12041 ), .Z(_u10_n12027 ) );
BUF_X4 _u10_U172  ( .A(_u10_n12065 ), .Z(_u10_n12051 ) );
BUF_X4 _u10_U171  ( .A(_u10_n12186 ), .Z(_u10_n12170 ) );
BUF_X4 _u10_U170  ( .A(_u10_n12234 ), .Z(_u10_n12218 ) );
BUF_X4 _u10_U169  ( .A(_u10_n12209 ), .Z(_u10_n12195 ) );
BUF_X4 _u10_U168  ( .A(_u10_n12258 ), .Z(_u10_n12242 ) );
BUF_X4 _u10_U167  ( .A(_u10_n12354 ), .Z(_u10_n12338 ) );
BUF_X4 _u10_U166  ( .A(_u10_n12043 ), .Z(_u10_n12021 ) );
BUF_X4 _u10_U165  ( .A(_u10_n12067 ), .Z(_u10_n12045 ) );
BUF_X4 _u10_U164  ( .A(_u10_n12187 ), .Z(_u10_n12165 ) );
BUF_X4 _u10_U163  ( .A(_u10_n12235 ), .Z(_u10_n12213 ) );
BUF_X4 _u10_U162  ( .A(_u10_n12211 ), .Z(_u10_n12189 ) );
BUF_X4 _u10_U161  ( .A(_u10_n12259 ), .Z(_u10_n12237 ) );
BUF_X4 _u10_U160  ( .A(_u10_n12355 ), .Z(_u10_n12333 ) );
BUF_X4 _u10_U159  ( .A(_u10_n12041 ), .Z(_u10_n12029 ) );
BUF_X4 _u10_U158  ( .A(_u10_n12065 ), .Z(_u10_n12053 ) );
BUF_X4 _u10_U157  ( .A(_u10_n12186 ), .Z(_u10_n12172 ) );
BUF_X4 _u10_U156  ( .A(_u10_n12234 ), .Z(_u10_n12220 ) );
BUF_X4 _u10_U155  ( .A(_u10_n12209 ), .Z(_u10_n12197 ) );
BUF_X4 _u10_U154  ( .A(_u10_n12040 ), .Z(_u10_n12035 ) );
BUF_X4 _u10_U153  ( .A(_u10_n12064 ), .Z(_u10_n12059 ) );
BUF_X4 _u10_U152  ( .A(_u10_n12184 ), .Z(_u10_n12181 ) );
BUF_X4 _u10_U151  ( .A(_u10_n12232 ), .Z(_u10_n12229 ) );
BUF_X4 _u10_U150  ( .A(_u10_n12212 ), .Z(_u10_n12203 ) );
BUF_X4 _u10_U149  ( .A(_u10_n12039 ), .Z(_u10_n12037 ) );
BUF_X4 _u10_U148  ( .A(_u10_n12063 ), .Z(_u10_n12061 ) );
BUF_X4 _u10_U147  ( .A(_u10_n12185 ), .Z(_u10_n12183 ) );
BUF_X4 _u10_U146  ( .A(_u10_n12233 ), .Z(_u10_n12231 ) );
BUF_X4 _u10_U145  ( .A(_u10_n12207 ), .Z(_u10_n12205 ) );
BUF_X4 _u10_U144  ( .A(_u10_n12257 ), .Z(_u10_n12255 ) );
BUF_X4 _u10_U143  ( .A(_u10_n12353 ), .Z(_u10_n12351 ) );
BUF_X4 _u10_U142  ( .A(_u10_n12041 ), .Z(_u10_n12034 ) );
BUF_X4 _u10_U141  ( .A(_u10_n12065 ), .Z(_u10_n12058 ) );
BUF_X4 _u10_U140  ( .A(_u10_n12188 ), .Z(_u10_n12180 ) );
BUF_X4 _u10_U139  ( .A(_u10_n12236 ), .Z(_u10_n12228 ) );
BUF_X4 _u10_U138  ( .A(_u10_n12206 ), .Z(_u10_n12202 ) );
BUF_X4 _u10_U137  ( .A(_u10_n12422 ), .Z(_u10_n12252 ) );
BUF_X4 _u10_U136  ( .A(_u10_n12279 ), .Z(_u10_n12277 ) );
BUF_X4 _u10_U135  ( .A(_u10_n12330 ), .Z(_u10_n12324 ) );
BUF_X4 _u10_U134  ( .A(_u10_n12303 ), .Z(_u10_n12301 ) );
BUF_X4 _u10_U133  ( .A(_u10_n12430 ), .Z(_u10_n12348 ) );
BUF_X4 _u10_U132  ( .A(_u10_n12186 ), .Z(_u10_n12177 ) );
BUF_X4 _u10_U131  ( .A(_u10_n12234 ), .Z(_u10_n12225 ) );
BUF_X4 _u10_U130  ( .A(_u10_n12207 ), .Z(_u10_n12199 ) );
BUF_X4 _u10_U129  ( .A(_u10_n12260 ), .Z(_u10_n12249 ) );
BUF_X4 _u10_U128  ( .A(_u10_n12356 ), .Z(_u10_n12345 ) );
BUF_X4 _u10_U127  ( .A(_u10_n12256 ), .Z(_u10_n12251 ) );
BUF_X4 _u10_U126  ( .A(_u10_n12352 ), .Z(_u10_n12347 ) );
BUF_X4 _u10_U125  ( .A(_u10_n12185 ), .Z(_u10_n12176 ) );
BUF_X4 _u10_U124  ( .A(_u10_n12233 ), .Z(_u10_n12224 ) );
BUF_X4 _u10_U123  ( .A(_u10_n12208 ), .Z(_u10_n12198 ) );
BUF_X4 _u10_U122  ( .A(_u10_n12258 ), .Z(_u10_n12248 ) );
BUF_X4 _u10_U121  ( .A(_u10_n12354 ), .Z(_u10_n12344 ) );
BUF_X4 _u10_U120  ( .A(_u10_n12257 ), .Z(_u10_n12250 ) );
BUF_X4 _u10_U119  ( .A(_u10_n12353 ), .Z(_u10_n12346 ) );
BUF_X4 _u10_U118  ( .A(_u10_n12038 ), .Z(_u10_n12032 ) );
BUF_X4 _u10_U117  ( .A(_u10_n12062 ), .Z(_u10_n12056 ) );
BUF_X4 _u10_U116  ( .A(_u10_n12187 ), .Z(_u10_n12175 ) );
BUF_X4 _u10_U115  ( .A(_u10_n12235 ), .Z(_u10_n12223 ) );
BUF_X4 _u10_U114  ( .A(_u10_n12259 ), .Z(_u10_n12247 ) );
BUF_X4 _u10_U113  ( .A(_u10_n12355 ), .Z(_u10_n12343 ) );
BUF_X4 _u10_U112  ( .A(_u10_n12044 ), .Z(_u10_n12031 ) );
BUF_X4 _u10_U111  ( .A(_u10_n12068 ), .Z(_u10_n12055 ) );
BUF_X4 _u10_U110  ( .A(_u10_n12187 ), .Z(_u10_n12174 ) );
BUF_X4 _u10_U109  ( .A(_u10_n12235 ), .Z(_u10_n12222 ) );
BUF_X4 _u10_U108  ( .A(_u10_n12259 ), .Z(_u10_n12246 ) );
BUF_X4 _u10_U107  ( .A(_u10_n12355 ), .Z(_u10_n12342 ) );
BUF_X4 _u10_U106  ( .A(_u10_n12258 ), .Z(_u10_n12244 ) );
BUF_X4 _u10_U105  ( .A(_u10_n12354 ), .Z(_u10_n12340 ) );
BUF_X4 _u10_U104  ( .A(_u10_n12260 ), .Z(_u10_n12253 ) );
BUF_X4 _u10_U103  ( .A(_u10_n12356 ), .Z(_u10_n12349 ) );
NAND2_X4 _u10_U102  ( .A1(_u10_n16748 ), .A2(_u10_n16749 ), .ZN(csr[2]) );
MUX2_X2 _u10_U101  ( .A(_u10_gnt_p0_d[4] ), .B(_u10_n22999 ), .S(dma_busy),.Z(ch_sel[4]) );
AND3_X4 _u10_U100  ( .A1(_u10_n22925 ), .A2(ch_sel[4]), .A3(ch_sel[2]), .ZN(_u10_n22924 ) );
AND3_X4 _u10_U99  ( .A1(ch_sel[2]), .A2(ch_sel[4]), .A3(_u10_n22911 ), .ZN(_u10_n12380 ) );
MUX2_X2 _u10_U98  ( .A(_u10_gnt_p0_d[2] ), .B(_u10_n22997 ), .S(dma_busy),.Z(ch_sel[2]) );
AND3_X4 _u10_U97  ( .A1(ch_sel[2]), .A2(ch_sel[3]), .A3(_u10_n22911 ), .ZN(_u10_n12396 ) );
MUX2_X2 _u10_U96  ( .A(_u10_gnt_p0_d[0] ), .B(_u10_n23000 ), .S(dma_busy),.Z(ch_sel[0]) );
MUX2_X2 _u10_U95  ( .A(_u10_gnt_p0_d[1] ), .B(_u10_n22996 ), .S(dma_busy),.Z(ch_sel[1]) );
MUX2_X2 _u10_U94  ( .A(_u10_gnt_p0_d[3] ), .B(_u10_n22998 ), .S(dma_busy),.Z(ch_sel[3]) );
INV_X4 _u10_U92  ( .A(1'b1), .ZN(_u10_ack_o[30] ) );
INV_X4 _u10_U90  ( .A(1'b1), .ZN(_u10_ack_o[29] ) );
INV_X4 _u10_U88  ( .A(1'b1), .ZN(_u10_ack_o[28] ) );
INV_X4 _u10_U86  ( .A(1'b1), .ZN(_u10_ack_o[27] ) );
INV_X4 _u10_U84  ( .A(1'b1), .ZN(_u10_ack_o[26] ) );
INV_X4 _u10_U82  ( .A(1'b1), .ZN(_u10_ack_o[25] ) );
INV_X4 _u10_U80  ( .A(1'b1), .ZN(_u10_ack_o[24] ) );
INV_X4 _u10_U78  ( .A(1'b1), .ZN(_u10_ack_o[23] ) );
INV_X4 _u10_U76  ( .A(1'b1), .ZN(_u10_ack_o[22] ) );
INV_X4 _u10_U74  ( .A(1'b1), .ZN(_u10_ack_o[21] ) );
INV_X4 _u10_U72  ( .A(1'b1), .ZN(_u10_ack_o[20] ) );
INV_X4 _u10_U70  ( .A(1'b1), .ZN(_u10_ack_o[19] ) );
INV_X4 _u10_U68  ( .A(1'b1), .ZN(_u10_ack_o[18] ) );
INV_X4 _u10_U66  ( .A(1'b1), .ZN(_u10_ack_o[17] ) );
INV_X4 _u10_U64  ( .A(1'b1), .ZN(_u10_ack_o[16] ) );
INV_X4 _u10_U62  ( .A(1'b1), .ZN(_u10_ack_o[15] ) );
INV_X4 _u10_U60  ( .A(1'b1), .ZN(_u10_ack_o[14] ) );
INV_X4 _u10_U58  ( .A(1'b1), .ZN(_u10_ack_o[13] ) );
INV_X4 _u10_U56  ( .A(1'b1), .ZN(_u10_ack_o[12] ) );
INV_X4 _u10_U54  ( .A(1'b1), .ZN(_u10_ack_o[11] ) );
INV_X4 _u10_U52  ( .A(1'b1), .ZN(_u10_ack_o[10] ) );
INV_X4 _u10_U50  ( .A(1'b1), .ZN(_u10_ack_o[9] ) );
INV_X4 _u10_U48  ( .A(1'b1), .ZN(_u10_ack_o[8] ) );
INV_X4 _u10_U46  ( .A(1'b1), .ZN(_u10_ack_o[7] ) );
INV_X4 _u10_U44  ( .A(1'b1), .ZN(_u10_ack_o[6] ) );
INV_X4 _u10_U42  ( .A(1'b1), .ZN(_u10_ack_o[5] ) );
INV_X4 _u10_U40  ( .A(1'b1), .ZN(_u10_ack_o[4] ) );
INV_X4 _u10_U38  ( .A(1'b1), .ZN(_u10_ack_o[3] ) );
INV_X4 _u10_U36  ( .A(1'b1), .ZN(_u10_ack_o[2] ) );
INV_X4 _u10_U34  ( .A(1'b1), .ZN(_u10_ack_o[1] ) );
DFF_X2 _u10_next_start_reg  ( .D(_u10_N1033 ), .CK(clk_i), .Q(), .QN(_u10_n11550 ) );
DFF_X2 _u10_de_start_r_reg  ( .D(_u10_n11552 ), .CK(clk_i), .Q(), .QN(_u10_n11551 ) );
DFF_X2 _u10_req_r_reg_0_  ( .D(_u10_N967 ), .CK(clk_i), .Q(_u10_req_r_0_ ),.QN() );
DFF_X2 _u10_ack_o_reg_0_  ( .D(_u10_N1034 ), .CK(clk_i), .Q(dma_ack_o[0]),.QN(_u10_n5 ) );
DFF_X2 _u10_ndnr_reg_0_  ( .D(_u10_N1032 ), .CK(clk_i), .Q(ndnr[0]), .QN());
DFF_X2 _u10_ndnr_reg_1_  ( .D(_u10_N1031 ), .CK(clk_i), .Q(ndnr[1]), .QN());
DFF_X2 _u10_ndnr_reg_2_  ( .D(_u10_N1030 ), .CK(clk_i), .Q(ndnr[2]), .QN());
DFF_X2 _u10_ndnr_reg_3_  ( .D(_u10_N1029 ), .CK(clk_i), .Q(ndnr[3]), .QN());
DFF_X2 _u10_ndnr_reg_4_  ( .D(_u10_N1028 ), .CK(clk_i), .Q(ndnr[4]), .QN());
DFF_X2 _u10_ndnr_reg_5_  ( .D(_u10_N1027 ), .CK(clk_i), .Q(ndnr[5]), .QN());
DFF_X2 _u10_ndnr_reg_6_  ( .D(_u10_N1026 ), .CK(clk_i), .Q(ndnr[6]), .QN());
DFF_X2 _u10_ndnr_reg_7_  ( .D(_u10_N1025 ), .CK(clk_i), .Q(ndnr[7]), .QN());
DFF_X2 _u10_ndnr_reg_8_  ( .D(_u10_N1024 ), .CK(clk_i), .Q(ndnr[8]), .QN());
DFF_X2 _u10_ndnr_reg_9_  ( .D(_u10_N1023 ), .CK(clk_i), .Q(ndnr[9]), .QN());
DFF_X2 _u10_ndnr_reg_10_  ( .D(_u10_N1022 ), .CK(clk_i), .Q(ndnr[10]), .QN());
DFF_X2 _u10_ndnr_reg_11_  ( .D(_u10_N1021 ), .CK(clk_i), .Q(ndnr[11]), .QN());
DFF_X2 _u10_ndnr_reg_12_  ( .D(_u10_N1020 ), .CK(clk_i), .Q(ndnr[12]), .QN());
DFF_X2 _u10_ndnr_reg_13_  ( .D(_u10_N1019 ), .CK(clk_i), .Q(ndnr[13]), .QN());
DFF_X2 _u10_ndnr_reg_14_  ( .D(_u10_N1018 ), .CK(clk_i), .Q(ndnr[14]), .QN());
DFF_X2 _u10_ndnr_reg_15_  ( .D(_u10_N1017 ), .CK(clk_i), .Q(ndnr[15]), .QN());
DFF_X2 _u10_ndnr_reg_16_  ( .D(_u10_N1016 ), .CK(clk_i), .Q(ndnr[16]), .QN());
DFF_X2 _u10_ndnr_reg_17_  ( .D(_u10_N1015 ), .CK(clk_i), .Q(ndnr[17]), .QN());
DFF_X2 _u10_ndnr_reg_18_  ( .D(_u10_N1014 ), .CK(clk_i), .Q(ndnr[18]), .QN());
DFF_X2 _u10_ndnr_reg_19_  ( .D(_u10_N1013 ), .CK(clk_i), .Q(ndnr[19]), .QN());
DFF_X2 _u10_ndnr_reg_20_  ( .D(_u10_N1012 ), .CK(clk_i), .Q(ndnr[20]), .QN());
DFF_X2 _u10_ndnr_reg_21_  ( .D(_u10_N1011 ), .CK(clk_i), .Q(ndnr[21]), .QN());
DFF_X2 _u10_ndnr_reg_22_  ( .D(_u10_N1010 ), .CK(clk_i), .Q(ndnr[22]), .QN());
DFF_X2 _u10_ndnr_reg_23_  ( .D(_u10_N1009 ), .CK(clk_i), .Q(ndnr[23]), .QN());
DFF_X2 _u10_ndnr_reg_24_  ( .D(_u10_N1008 ), .CK(clk_i), .Q(ndnr[24]), .QN());
DFF_X2 _u10_ndnr_reg_25_  ( .D(_u10_N1007 ), .CK(clk_i), .Q(ndnr[25]), .QN());
DFF_X2 _u10_ndnr_reg_26_  ( .D(_u10_N1006 ), .CK(clk_i), .Q(ndnr[26]), .QN());
DFF_X2 _u10_ndnr_reg_27_  ( .D(_u10_N1005 ), .CK(clk_i), .Q(ndnr[27]), .QN());
DFF_X2 _u10_ndnr_reg_28_  ( .D(_u10_N1004 ), .CK(clk_i), .Q(ndnr[28]), .QN());
DFF_X2 _u10_ndnr_reg_29_  ( .D(_u10_N1003 ), .CK(clk_i), .Q(ndnr[29]), .QN());
DFF_X2 _u10_ndnr_reg_30_  ( .D(_u10_N1002 ), .CK(clk_i), .Q(ndnr[30]), .QN());
DFF_X2 _u10_ndr_r_reg_1_  ( .D(_u10_N1000 ), .CK(clk_i), .Q(), .QN(_u10_n22991 ) );
DFF_X2 _u10_ndr_r_reg_2_  ( .D(_u10_N999 ), .CK(clk_i), .Q(), .QN(_u10_n22990 ) );
DFF_X2 _u10_ndr_r_reg_3_  ( .D(_u10_N998 ), .CK(clk_i), .Q(_u10_n22994 ),.QN() );
DFF_X2 _u10_ndr_r_reg_4_  ( .D(_u10_N997 ), .CK(clk_i), .Q(_u10_n22995 ),.QN() );
DFF_X2 _u10_ndr_r_reg_5_  ( .D(_u10_N996 ), .CK(clk_i), .Q(), .QN(_u10_n11543 ) );
DFF_X2 _u10_ndr_r_reg_6_  ( .D(_u10_N995 ), .CK(clk_i), .Q(), .QN(_u10_n11542 ) );
DFF_X2 _u10_ndr_r_reg_7_  ( .D(_u10_N994 ), .CK(clk_i), .Q(), .QN(_u10_n10663 ) );
DFF_X2 _u10_ndr_r_reg_8_  ( .D(_u10_N993 ), .CK(clk_i), .Q(), .QN(_u10_n10662 ) );
DFF_X2 _u10_ndr_r_reg_9_  ( .D(_u10_N992 ), .CK(clk_i), .Q(), .QN(_u10_n22989 ) );
DFF_X2 _u10_ndr_r_reg_10_  ( .D(_u10_N991 ), .CK(clk_i), .Q(), .QN(_u10_n22988 ) );
DFF_X2 _u10_ndr_r_reg_11_  ( .D(_u10_N990 ), .CK(clk_i), .Q(_u10_n22992 ),.QN() );
DFF_X2 _u10_ndr_r_reg_12_  ( .D(_u10_N989 ), .CK(clk_i), .Q(_u10_n22993 ),.QN() );
DFF_X2 _u10_ndr_r_reg_13_  ( .D(_u10_N988 ), .CK(clk_i), .Q(), .QN(_u10_n10665 ) );
DFF_X2 _u10_ndr_r_reg_14_  ( .D(_u10_N987 ), .CK(clk_i), .Q(), .QN(_u10_n10664 ) );
DFF_X2 _u10_ndr_r_reg_15_  ( .D(_u10_N986 ), .CK(clk_i), .Q(_u10_ndr_r[15]),.QN() );
DFF_X2 _u10_ndr_r_reg_16_  ( .D(_u10_N985 ), .CK(clk_i), .Q(_u10_ndr_r[16]),.QN() );
DFF_X2 _u10_ndr_r_reg_17_  ( .D(_u10_N984 ), .CK(clk_i), .Q(_u10_ndr_r[17]),.QN() );
DFF_X2 _u10_ndr_r_reg_18_  ( .D(_u10_N983 ), .CK(clk_i), .Q(_u10_ndr_r[18]),.QN() );
DFF_X2 _u10_ndr_r_reg_19_  ( .D(_u10_N982 ), .CK(clk_i), .Q(_u10_ndr_r[19]),.QN() );
DFF_X2 _u10_ndr_r_reg_20_  ( .D(_u10_N981 ), .CK(clk_i), .Q(_u10_ndr_r[20]),.QN() );
DFF_X2 _u10_ndr_r_reg_21_  ( .D(_u10_N980 ), .CK(clk_i), .Q(_u10_ndr_r[21]),.QN() );
DFF_X2 _u10_ndr_r_reg_22_  ( .D(_u10_N979 ), .CK(clk_i), .Q(_u10_ndr_r[22]),.QN() );
DFF_X2 _u10_ndr_r_reg_23_  ( .D(_u10_N978 ), .CK(clk_i), .Q(_u10_ndr_r[23]),.QN() );
DFF_X2 _u10_ndr_r_reg_24_  ( .D(_u10_N977 ), .CK(clk_i), .Q(_u10_ndr_r[24]),.QN() );
DFF_X2 _u10_ndr_r_reg_25_  ( .D(_u10_N976 ), .CK(clk_i), .Q(_u10_ndr_r[25]),.QN() );
DFF_X2 _u10_ndr_r_reg_26_  ( .D(_u10_N975 ), .CK(clk_i), .Q(_u10_ndr_r[26]),.QN() );
DFF_X2 _u10_ndr_r_reg_27_  ( .D(_u10_N974 ), .CK(clk_i), .Q(_u10_ndr_r[27]),.QN() );
DFF_X2 _u10_ndr_r_reg_28_  ( .D(_u10_N973 ), .CK(clk_i), .Q(_u10_ndr_r[28]),.QN() );
DFF_X2 _u10_ndr_r_reg_29_  ( .D(_u10_N972 ), .CK(clk_i), .Q(_u10_ndr_r[29]),.QN() );
DFF_X2 _u10_ndr_r_reg_30_  ( .D(_u10_N971 ), .CK(clk_i), .Q(_u10_ndr_r[30]),.QN() );
DFFR_X1 _u10_ch_sel_r_reg_1_  ( .D(_u10_n10675 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_n22996 ), .QN() );
DFFR_X1 _u10_ch_sel_r_reg_2_  ( .D(_u10_n10674 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_n22997 ), .QN() );
DFFR_X1 _u10_ch_sel_r_reg_3_  ( .D(_u10_n10673 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_n22998 ), .QN() );
DFFR_X1 _u10_ch_sel_r_reg_4_  ( .D(_u10_n10672 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_n22999 ), .QN() );
DFFR_X1 _u10_ch_sel_r_reg_0_  ( .D(_u10_n10676 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_n23000 ), .QN() );
SDFF_X2 _u10_ndr_r_reg_0_  ( .D(dma_nd_i[0]), .SI(1'b0), .SE(_u10_n23001 ),.CK(clk_i), .Q(), .QN(_u10_n11539 ) );
INV_X4 _u10_u0_U100  ( .A(1'b1), .ZN(_u10_u0_pri_out[2] ) );
INV_X4 _u10_u0_U80  ( .A(1'b1), .ZN(_u10_u0_pri_out[1] ) );
INV_X4 _u10_u0_U60  ( .A(1'b1), .ZN(_u10_u0_pri_out[0] ) );
INV_X4 _u10_u0_u0_U16  ( .A(1'b1), .ZN(_u10_u0_u0_pri_out[7] ) );
INV_X4 _u10_u0_u0_U14  ( .A(1'b1), .ZN(_u10_u0_u0_pri_out[6] ) );
INV_X4 _u10_u0_u0_U12  ( .A(1'b1), .ZN(_u10_u0_u0_pri_out[5] ) );
INV_X4 _u10_u0_u0_U10  ( .A(1'b1), .ZN(_u10_u0_u0_pri_out[4] ) );
INV_X4 _u10_u0_u0_U8  ( .A(1'b1), .ZN(_u10_u0_u0_pri_out[3] ) );
INV_X4 _u10_u0_u0_U6  ( .A(1'b1), .ZN(_u10_u0_u0_pri_out[2] ) );
INV_X4 _u10_u0_u0_U4  ( .A(1'b1), .ZN(_u10_u0_u0_pri_out[1] ) );
INV_X4 _u10_u0_u0_U2  ( .A(1'b1), .ZN(_u10_u0_u0_pri_out[0] ) );
INV_X4 _u10_u0_u1_U16  ( .A(1'b1), .ZN(_u10_u0_u1_pri_out[7] ) );
INV_X4 _u10_u0_u1_U14  ( .A(1'b1), .ZN(_u10_u0_u1_pri_out[6] ) );
INV_X4 _u10_u0_u1_U12  ( .A(1'b1), .ZN(_u10_u0_u1_pri_out[5] ) );
INV_X4 _u10_u0_u1_U10  ( .A(1'b1), .ZN(_u10_u0_u1_pri_out[4] ) );
INV_X4 _u10_u0_u1_U8  ( .A(1'b1), .ZN(_u10_u0_u1_pri_out[3] ) );
INV_X4 _u10_u0_u1_U6  ( .A(1'b1), .ZN(_u10_u0_u1_pri_out[2] ) );
INV_X4 _u10_u0_u1_U4  ( .A(1'b1), .ZN(_u10_u0_u1_pri_out[1] ) );
INV_X4 _u10_u0_u1_U2  ( .A(1'b1), .ZN(_u10_u0_u1_pri_out[0] ) );
INV_X4 _u10_u0_u2_U16  ( .A(1'b1), .ZN(_u10_u0_u2_pri_out[7] ) );
INV_X4 _u10_u0_u2_U14  ( .A(1'b1), .ZN(_u10_u0_u2_pri_out[6] ) );
INV_X4 _u10_u0_u2_U12  ( .A(1'b1), .ZN(_u10_u0_u2_pri_out[5] ) );
INV_X4 _u10_u0_u2_U10  ( .A(1'b1), .ZN(_u10_u0_u2_pri_out[4] ) );
INV_X4 _u10_u0_u2_U8  ( .A(1'b1), .ZN(_u10_u0_u2_pri_out[3] ) );
INV_X4 _u10_u0_u2_U6  ( .A(1'b1), .ZN(_u10_u0_u2_pri_out[2] ) );
INV_X4 _u10_u0_u2_U4  ( .A(1'b1), .ZN(_u10_u0_u2_pri_out[1] ) );
INV_X4 _u10_u0_u2_U2  ( .A(1'b1), .ZN(_u10_u0_u2_pri_out[0] ) );
INV_X4 _u10_u0_u3_U16  ( .A(1'b1), .ZN(_u10_u0_u3_pri_out[7] ) );
INV_X4 _u10_u0_u3_U14  ( .A(1'b1), .ZN(_u10_u0_u3_pri_out[6] ) );
INV_X4 _u10_u0_u3_U12  ( .A(1'b1), .ZN(_u10_u0_u3_pri_out[5] ) );
INV_X4 _u10_u0_u3_U10  ( .A(1'b1), .ZN(_u10_u0_u3_pri_out[4] ) );
INV_X4 _u10_u0_u3_U8  ( .A(1'b1), .ZN(_u10_u0_u3_pri_out[3] ) );
INV_X4 _u10_u0_u3_U6  ( .A(1'b1), .ZN(_u10_u0_u3_pri_out[2] ) );
INV_X4 _u10_u0_u3_U4  ( .A(1'b1), .ZN(_u10_u0_u3_pri_out[1] ) );
INV_X4 _u10_u0_u3_U2  ( .A(1'b1), .ZN(_u10_u0_u3_pri_out[0] ) );
INV_X4 _u10_u0_u4_U16  ( .A(1'b1), .ZN(_u10_u0_u4_pri_out[7] ) );
INV_X4 _u10_u0_u4_U14  ( .A(1'b1), .ZN(_u10_u0_u4_pri_out[6] ) );
INV_X4 _u10_u0_u4_U12  ( .A(1'b1), .ZN(_u10_u0_u4_pri_out[5] ) );
INV_X4 _u10_u0_u4_U10  ( .A(1'b1), .ZN(_u10_u0_u4_pri_out[4] ) );
INV_X4 _u10_u0_u4_U8  ( .A(1'b1), .ZN(_u10_u0_u4_pri_out[3] ) );
INV_X4 _u10_u0_u4_U6  ( .A(1'b1), .ZN(_u10_u0_u4_pri_out[2] ) );
INV_X4 _u10_u0_u4_U4  ( .A(1'b1), .ZN(_u10_u0_u4_pri_out[1] ) );
INV_X4 _u10_u0_u4_U2  ( .A(1'b1), .ZN(_u10_u0_u4_pri_out[0] ) );
INV_X4 _u10_u0_u5_U16  ( .A(1'b1), .ZN(_u10_u0_u5_pri_out[7] ) );
INV_X4 _u10_u0_u5_U14  ( .A(1'b1), .ZN(_u10_u0_u5_pri_out[6] ) );
INV_X4 _u10_u0_u5_U12  ( .A(1'b1), .ZN(_u10_u0_u5_pri_out[5] ) );
INV_X4 _u10_u0_u5_U10  ( .A(1'b1), .ZN(_u10_u0_u5_pri_out[4] ) );
INV_X4 _u10_u0_u5_U8  ( .A(1'b1), .ZN(_u10_u0_u5_pri_out[3] ) );
INV_X4 _u10_u0_u5_U6  ( .A(1'b1), .ZN(_u10_u0_u5_pri_out[2] ) );
INV_X4 _u10_u0_u5_U4  ( .A(1'b1), .ZN(_u10_u0_u5_pri_out[1] ) );
INV_X4 _u10_u0_u5_U2  ( .A(1'b1), .ZN(_u10_u0_u5_pri_out[0] ) );
INV_X4 _u10_u0_u6_U16  ( .A(1'b1), .ZN(_u10_u0_u6_pri_out[7] ) );
INV_X4 _u10_u0_u6_U14  ( .A(1'b1), .ZN(_u10_u0_u6_pri_out[6] ) );
INV_X4 _u10_u0_u6_U12  ( .A(1'b1), .ZN(_u10_u0_u6_pri_out[5] ) );
INV_X4 _u10_u0_u6_U10  ( .A(1'b1), .ZN(_u10_u0_u6_pri_out[4] ) );
INV_X4 _u10_u0_u6_U8  ( .A(1'b1), .ZN(_u10_u0_u6_pri_out[3] ) );
INV_X4 _u10_u0_u6_U6  ( .A(1'b1), .ZN(_u10_u0_u6_pri_out[2] ) );
INV_X4 _u10_u0_u6_U4  ( .A(1'b1), .ZN(_u10_u0_u6_pri_out[1] ) );
INV_X4 _u10_u0_u6_U2  ( .A(1'b1), .ZN(_u10_u0_u6_pri_out[0] ) );
INV_X4 _u10_u0_u7_U16  ( .A(1'b1), .ZN(_u10_u0_u7_pri_out[7] ) );
INV_X4 _u10_u0_u7_U14  ( .A(1'b1), .ZN(_u10_u0_u7_pri_out[6] ) );
INV_X4 _u10_u0_u7_U12  ( .A(1'b1), .ZN(_u10_u0_u7_pri_out[5] ) );
INV_X4 _u10_u0_u7_U10  ( .A(1'b1), .ZN(_u10_u0_u7_pri_out[4] ) );
INV_X4 _u10_u0_u7_U8  ( .A(1'b1), .ZN(_u10_u0_u7_pri_out[3] ) );
INV_X4 _u10_u0_u7_U6  ( .A(1'b1), .ZN(_u10_u0_u7_pri_out[2] ) );
INV_X4 _u10_u0_u7_U4  ( .A(1'b1), .ZN(_u10_u0_u7_pri_out[1] ) );
INV_X4 _u10_u0_u7_U2  ( .A(1'b1), .ZN(_u10_u0_u7_pri_out[0] ) );
INV_X4 _u10_u0_u8_U16  ( .A(1'b1), .ZN(_u10_u0_u8_pri_out[7] ) );
INV_X4 _u10_u0_u8_U14  ( .A(1'b1), .ZN(_u10_u0_u8_pri_out[6] ) );
INV_X4 _u10_u0_u8_U12  ( .A(1'b1), .ZN(_u10_u0_u8_pri_out[5] ) );
INV_X4 _u10_u0_u8_U10  ( .A(1'b1), .ZN(_u10_u0_u8_pri_out[4] ) );
INV_X4 _u10_u0_u8_U8  ( .A(1'b1), .ZN(_u10_u0_u8_pri_out[3] ) );
INV_X4 _u10_u0_u8_U6  ( .A(1'b1), .ZN(_u10_u0_u8_pri_out[2] ) );
INV_X4 _u10_u0_u8_U4  ( .A(1'b1), .ZN(_u10_u0_u8_pri_out[1] ) );
INV_X4 _u10_u0_u8_U2  ( .A(1'b1), .ZN(_u10_u0_u8_pri_out[0] ) );
INV_X4 _u10_u0_u9_U16  ( .A(1'b1), .ZN(_u10_u0_u9_pri_out[7] ) );
INV_X4 _u10_u0_u9_U14  ( .A(1'b1), .ZN(_u10_u0_u9_pri_out[6] ) );
INV_X4 _u10_u0_u9_U12  ( .A(1'b1), .ZN(_u10_u0_u9_pri_out[5] ) );
INV_X4 _u10_u0_u9_U10  ( .A(1'b1), .ZN(_u10_u0_u9_pri_out[4] ) );
INV_X4 _u10_u0_u9_U8  ( .A(1'b1), .ZN(_u10_u0_u9_pri_out[3] ) );
INV_X4 _u10_u0_u9_U6  ( .A(1'b1), .ZN(_u10_u0_u9_pri_out[2] ) );
INV_X4 _u10_u0_u9_U4  ( .A(1'b1), .ZN(_u10_u0_u9_pri_out[1] ) );
INV_X4 _u10_u0_u9_U2  ( .A(1'b1), .ZN(_u10_u0_u9_pri_out[0] ) );
INV_X4 _u10_u0_u10_U16  ( .A(1'b1), .ZN(_u10_u0_u10_pri_out[7] ) );
INV_X4 _u10_u0_u10_U14  ( .A(1'b1), .ZN(_u10_u0_u10_pri_out[6] ) );
INV_X4 _u10_u0_u10_U12  ( .A(1'b1), .ZN(_u10_u0_u10_pri_out[5] ) );
INV_X4 _u10_u0_u10_U10  ( .A(1'b1), .ZN(_u10_u0_u10_pri_out[4] ) );
INV_X4 _u10_u0_u10_U8  ( .A(1'b1), .ZN(_u10_u0_u10_pri_out[3] ) );
INV_X4 _u10_u0_u10_U6  ( .A(1'b1), .ZN(_u10_u0_u10_pri_out[2] ) );
INV_X4 _u10_u0_u10_U4  ( .A(1'b1), .ZN(_u10_u0_u10_pri_out[1] ) );
INV_X4 _u10_u0_u10_U2  ( .A(1'b1), .ZN(_u10_u0_u10_pri_out[0] ) );
INV_X4 _u10_u0_u11_U16  ( .A(1'b1), .ZN(_u10_u0_u11_pri_out[7] ) );
INV_X4 _u10_u0_u11_U14  ( .A(1'b1), .ZN(_u10_u0_u11_pri_out[6] ) );
INV_X4 _u10_u0_u11_U12  ( .A(1'b1), .ZN(_u10_u0_u11_pri_out[5] ) );
INV_X4 _u10_u0_u11_U10  ( .A(1'b1), .ZN(_u10_u0_u11_pri_out[4] ) );
INV_X4 _u10_u0_u11_U8  ( .A(1'b1), .ZN(_u10_u0_u11_pri_out[3] ) );
INV_X4 _u10_u0_u11_U6  ( .A(1'b1), .ZN(_u10_u0_u11_pri_out[2] ) );
INV_X4 _u10_u0_u11_U4  ( .A(1'b1), .ZN(_u10_u0_u11_pri_out[1] ) );
INV_X4 _u10_u0_u11_U2  ( .A(1'b1), .ZN(_u10_u0_u11_pri_out[0] ) );
INV_X4 _u10_u0_u12_U16  ( .A(1'b1), .ZN(_u10_u0_u12_pri_out[7] ) );
INV_X4 _u10_u0_u12_U14  ( .A(1'b1), .ZN(_u10_u0_u12_pri_out[6] ) );
INV_X4 _u10_u0_u12_U12  ( .A(1'b1), .ZN(_u10_u0_u12_pri_out[5] ) );
INV_X4 _u10_u0_u12_U10  ( .A(1'b1), .ZN(_u10_u0_u12_pri_out[4] ) );
INV_X4 _u10_u0_u12_U8  ( .A(1'b1), .ZN(_u10_u0_u12_pri_out[3] ) );
INV_X4 _u10_u0_u12_U6  ( .A(1'b1), .ZN(_u10_u0_u12_pri_out[2] ) );
INV_X4 _u10_u0_u12_U4  ( .A(1'b1), .ZN(_u10_u0_u12_pri_out[1] ) );
INV_X4 _u10_u0_u12_U2  ( .A(1'b1), .ZN(_u10_u0_u12_pri_out[0] ) );
INV_X4 _u10_u0_u13_U16  ( .A(1'b1), .ZN(_u10_u0_u13_pri_out[7] ) );
INV_X4 _u10_u0_u13_U14  ( .A(1'b1), .ZN(_u10_u0_u13_pri_out[6] ) );
INV_X4 _u10_u0_u13_U12  ( .A(1'b1), .ZN(_u10_u0_u13_pri_out[5] ) );
INV_X4 _u10_u0_u13_U10  ( .A(1'b1), .ZN(_u10_u0_u13_pri_out[4] ) );
INV_X4 _u10_u0_u13_U8  ( .A(1'b1), .ZN(_u10_u0_u13_pri_out[3] ) );
INV_X4 _u10_u0_u13_U6  ( .A(1'b1), .ZN(_u10_u0_u13_pri_out[2] ) );
INV_X4 _u10_u0_u13_U4  ( .A(1'b1), .ZN(_u10_u0_u13_pri_out[1] ) );
INV_X4 _u10_u0_u13_U2  ( .A(1'b1), .ZN(_u10_u0_u13_pri_out[0] ) );
INV_X4 _u10_u0_u14_U16  ( .A(1'b1), .ZN(_u10_u0_u14_pri_out[7] ) );
INV_X4 _u10_u0_u14_U14  ( .A(1'b1), .ZN(_u10_u0_u14_pri_out[6] ) );
INV_X4 _u10_u0_u14_U12  ( .A(1'b1), .ZN(_u10_u0_u14_pri_out[5] ) );
INV_X4 _u10_u0_u14_U10  ( .A(1'b1), .ZN(_u10_u0_u14_pri_out[4] ) );
INV_X4 _u10_u0_u14_U8  ( .A(1'b1), .ZN(_u10_u0_u14_pri_out[3] ) );
INV_X4 _u10_u0_u14_U6  ( .A(1'b1), .ZN(_u10_u0_u14_pri_out[2] ) );
INV_X4 _u10_u0_u14_U4  ( .A(1'b1), .ZN(_u10_u0_u14_pri_out[1] ) );
INV_X4 _u10_u0_u14_U2  ( .A(1'b1), .ZN(_u10_u0_u14_pri_out[0] ) );
INV_X4 _u10_u0_u15_U16  ( .A(1'b1), .ZN(_u10_u0_u15_pri_out[7] ) );
INV_X4 _u10_u0_u15_U14  ( .A(1'b1), .ZN(_u10_u0_u15_pri_out[6] ) );
INV_X4 _u10_u0_u15_U12  ( .A(1'b1), .ZN(_u10_u0_u15_pri_out[5] ) );
INV_X4 _u10_u0_u15_U10  ( .A(1'b1), .ZN(_u10_u0_u15_pri_out[4] ) );
INV_X4 _u10_u0_u15_U8  ( .A(1'b1), .ZN(_u10_u0_u15_pri_out[3] ) );
INV_X4 _u10_u0_u15_U6  ( .A(1'b1), .ZN(_u10_u0_u15_pri_out[2] ) );
INV_X4 _u10_u0_u15_U4  ( .A(1'b1), .ZN(_u10_u0_u15_pri_out[1] ) );
INV_X4 _u10_u0_u15_U2  ( .A(1'b1), .ZN(_u10_u0_u15_pri_out[0] ) );
INV_X4 _u10_u0_u16_U16  ( .A(1'b1), .ZN(_u10_u0_u16_pri_out[7] ) );
INV_X4 _u10_u0_u16_U14  ( .A(1'b1), .ZN(_u10_u0_u16_pri_out[6] ) );
INV_X4 _u10_u0_u16_U12  ( .A(1'b1), .ZN(_u10_u0_u16_pri_out[5] ) );
INV_X4 _u10_u0_u16_U10  ( .A(1'b1), .ZN(_u10_u0_u16_pri_out[4] ) );
INV_X4 _u10_u0_u16_U8  ( .A(1'b1), .ZN(_u10_u0_u16_pri_out[3] ) );
INV_X4 _u10_u0_u16_U6  ( .A(1'b1), .ZN(_u10_u0_u16_pri_out[2] ) );
INV_X4 _u10_u0_u16_U4  ( .A(1'b1), .ZN(_u10_u0_u16_pri_out[1] ) );
INV_X4 _u10_u0_u16_U2  ( .A(1'b1), .ZN(_u10_u0_u16_pri_out[0] ) );
INV_X4 _u10_u0_u17_U16  ( .A(1'b1), .ZN(_u10_u0_u17_pri_out[7] ) );
INV_X4 _u10_u0_u17_U14  ( .A(1'b1), .ZN(_u10_u0_u17_pri_out[6] ) );
INV_X4 _u10_u0_u17_U12  ( .A(1'b1), .ZN(_u10_u0_u17_pri_out[5] ) );
INV_X4 _u10_u0_u17_U10  ( .A(1'b1), .ZN(_u10_u0_u17_pri_out[4] ) );
INV_X4 _u10_u0_u17_U8  ( .A(1'b1), .ZN(_u10_u0_u17_pri_out[3] ) );
INV_X4 _u10_u0_u17_U6  ( .A(1'b1), .ZN(_u10_u0_u17_pri_out[2] ) );
INV_X4 _u10_u0_u17_U4  ( .A(1'b1), .ZN(_u10_u0_u17_pri_out[1] ) );
INV_X4 _u10_u0_u17_U2  ( .A(1'b1), .ZN(_u10_u0_u17_pri_out[0] ) );
INV_X4 _u10_u0_u18_U16  ( .A(1'b1), .ZN(_u10_u0_u18_pri_out[7] ) );
INV_X4 _u10_u0_u18_U14  ( .A(1'b1), .ZN(_u10_u0_u18_pri_out[6] ) );
INV_X4 _u10_u0_u18_U12  ( .A(1'b1), .ZN(_u10_u0_u18_pri_out[5] ) );
INV_X4 _u10_u0_u18_U10  ( .A(1'b1), .ZN(_u10_u0_u18_pri_out[4] ) );
INV_X4 _u10_u0_u18_U8  ( .A(1'b1), .ZN(_u10_u0_u18_pri_out[3] ) );
INV_X4 _u10_u0_u18_U6  ( .A(1'b1), .ZN(_u10_u0_u18_pri_out[2] ) );
INV_X4 _u10_u0_u18_U4  ( .A(1'b1), .ZN(_u10_u0_u18_pri_out[1] ) );
INV_X4 _u10_u0_u18_U2  ( .A(1'b1), .ZN(_u10_u0_u18_pri_out[0] ) );
INV_X4 _u10_u0_u19_U16  ( .A(1'b1), .ZN(_u10_u0_u19_pri_out[7] ) );
INV_X4 _u10_u0_u19_U14  ( .A(1'b1), .ZN(_u10_u0_u19_pri_out[6] ) );
INV_X4 _u10_u0_u19_U12  ( .A(1'b1), .ZN(_u10_u0_u19_pri_out[5] ) );
INV_X4 _u10_u0_u19_U10  ( .A(1'b1), .ZN(_u10_u0_u19_pri_out[4] ) );
INV_X4 _u10_u0_u19_U8  ( .A(1'b1), .ZN(_u10_u0_u19_pri_out[3] ) );
INV_X4 _u10_u0_u19_U6  ( .A(1'b1), .ZN(_u10_u0_u19_pri_out[2] ) );
INV_X4 _u10_u0_u19_U4  ( .A(1'b1), .ZN(_u10_u0_u19_pri_out[1] ) );
INV_X4 _u10_u0_u19_U2  ( .A(1'b1), .ZN(_u10_u0_u19_pri_out[0] ) );
INV_X4 _u10_u0_u20_U16  ( .A(1'b1), .ZN(_u10_u0_u20_pri_out[7] ) );
INV_X4 _u10_u0_u20_U14  ( .A(1'b1), .ZN(_u10_u0_u20_pri_out[6] ) );
INV_X4 _u10_u0_u20_U12  ( .A(1'b1), .ZN(_u10_u0_u20_pri_out[5] ) );
INV_X4 _u10_u0_u20_U10  ( .A(1'b1), .ZN(_u10_u0_u20_pri_out[4] ) );
INV_X4 _u10_u0_u20_U8  ( .A(1'b1), .ZN(_u10_u0_u20_pri_out[3] ) );
INV_X4 _u10_u0_u20_U6  ( .A(1'b1), .ZN(_u10_u0_u20_pri_out[2] ) );
INV_X4 _u10_u0_u20_U4  ( .A(1'b1), .ZN(_u10_u0_u20_pri_out[1] ) );
INV_X4 _u10_u0_u20_U2  ( .A(1'b1), .ZN(_u10_u0_u20_pri_out[0] ) );
INV_X4 _u10_u0_u21_U16  ( .A(1'b1), .ZN(_u10_u0_u21_pri_out[7] ) );
INV_X4 _u10_u0_u21_U14  ( .A(1'b1), .ZN(_u10_u0_u21_pri_out[6] ) );
INV_X4 _u10_u0_u21_U12  ( .A(1'b1), .ZN(_u10_u0_u21_pri_out[5] ) );
INV_X4 _u10_u0_u21_U10  ( .A(1'b1), .ZN(_u10_u0_u21_pri_out[4] ) );
INV_X4 _u10_u0_u21_U8  ( .A(1'b1), .ZN(_u10_u0_u21_pri_out[3] ) );
INV_X4 _u10_u0_u21_U6  ( .A(1'b1), .ZN(_u10_u0_u21_pri_out[2] ) );
INV_X4 _u10_u0_u21_U4  ( .A(1'b1), .ZN(_u10_u0_u21_pri_out[1] ) );
INV_X4 _u10_u0_u21_U2  ( .A(1'b1), .ZN(_u10_u0_u21_pri_out[0] ) );
INV_X4 _u10_u0_u22_U16  ( .A(1'b1), .ZN(_u10_u0_u22_pri_out[7] ) );
INV_X4 _u10_u0_u22_U14  ( .A(1'b1), .ZN(_u10_u0_u22_pri_out[6] ) );
INV_X4 _u10_u0_u22_U12  ( .A(1'b1), .ZN(_u10_u0_u22_pri_out[5] ) );
INV_X4 _u10_u0_u22_U10  ( .A(1'b1), .ZN(_u10_u0_u22_pri_out[4] ) );
INV_X4 _u10_u0_u22_U8  ( .A(1'b1), .ZN(_u10_u0_u22_pri_out[3] ) );
INV_X4 _u10_u0_u22_U6  ( .A(1'b1), .ZN(_u10_u0_u22_pri_out[2] ) );
INV_X4 _u10_u0_u22_U4  ( .A(1'b1), .ZN(_u10_u0_u22_pri_out[1] ) );
INV_X4 _u10_u0_u22_U2  ( .A(1'b1), .ZN(_u10_u0_u22_pri_out[0] ) );
INV_X4 _u10_u0_u23_U16  ( .A(1'b1), .ZN(_u10_u0_u23_pri_out[7] ) );
INV_X4 _u10_u0_u23_U14  ( .A(1'b1), .ZN(_u10_u0_u23_pri_out[6] ) );
INV_X4 _u10_u0_u23_U12  ( .A(1'b1), .ZN(_u10_u0_u23_pri_out[5] ) );
INV_X4 _u10_u0_u23_U10  ( .A(1'b1), .ZN(_u10_u0_u23_pri_out[4] ) );
INV_X4 _u10_u0_u23_U8  ( .A(1'b1), .ZN(_u10_u0_u23_pri_out[3] ) );
INV_X4 _u10_u0_u23_U6  ( .A(1'b1), .ZN(_u10_u0_u23_pri_out[2] ) );
INV_X4 _u10_u0_u23_U4  ( .A(1'b1), .ZN(_u10_u0_u23_pri_out[1] ) );
INV_X4 _u10_u0_u23_U2  ( .A(1'b1), .ZN(_u10_u0_u23_pri_out[0] ) );
INV_X4 _u10_u0_u24_U16  ( .A(1'b1), .ZN(_u10_u0_u24_pri_out[7] ) );
INV_X4 _u10_u0_u24_U14  ( .A(1'b1), .ZN(_u10_u0_u24_pri_out[6] ) );
INV_X4 _u10_u0_u24_U12  ( .A(1'b1), .ZN(_u10_u0_u24_pri_out[5] ) );
INV_X4 _u10_u0_u24_U10  ( .A(1'b1), .ZN(_u10_u0_u24_pri_out[4] ) );
INV_X4 _u10_u0_u24_U8  ( .A(1'b1), .ZN(_u10_u0_u24_pri_out[3] ) );
INV_X4 _u10_u0_u24_U6  ( .A(1'b1), .ZN(_u10_u0_u24_pri_out[2] ) );
INV_X4 _u10_u0_u24_U4  ( .A(1'b1), .ZN(_u10_u0_u24_pri_out[1] ) );
INV_X4 _u10_u0_u24_U2  ( .A(1'b1), .ZN(_u10_u0_u24_pri_out[0] ) );
INV_X4 _u10_u0_u25_U16  ( .A(1'b1), .ZN(_u10_u0_u25_pri_out[7] ) );
INV_X4 _u10_u0_u25_U14  ( .A(1'b1), .ZN(_u10_u0_u25_pri_out[6] ) );
INV_X4 _u10_u0_u25_U12  ( .A(1'b1), .ZN(_u10_u0_u25_pri_out[5] ) );
INV_X4 _u10_u0_u25_U10  ( .A(1'b1), .ZN(_u10_u0_u25_pri_out[4] ) );
INV_X4 _u10_u0_u25_U8  ( .A(1'b1), .ZN(_u10_u0_u25_pri_out[3] ) );
INV_X4 _u10_u0_u25_U6  ( .A(1'b1), .ZN(_u10_u0_u25_pri_out[2] ) );
INV_X4 _u10_u0_u25_U4  ( .A(1'b1), .ZN(_u10_u0_u25_pri_out[1] ) );
INV_X4 _u10_u0_u25_U2  ( .A(1'b1), .ZN(_u10_u0_u25_pri_out[0] ) );
INV_X4 _u10_u0_u26_U16  ( .A(1'b1), .ZN(_u10_u0_u26_pri_out[7] ) );
INV_X4 _u10_u0_u26_U14  ( .A(1'b1), .ZN(_u10_u0_u26_pri_out[6] ) );
INV_X4 _u10_u0_u26_U12  ( .A(1'b1), .ZN(_u10_u0_u26_pri_out[5] ) );
INV_X4 _u10_u0_u26_U10  ( .A(1'b1), .ZN(_u10_u0_u26_pri_out[4] ) );
INV_X4 _u10_u0_u26_U8  ( .A(1'b1), .ZN(_u10_u0_u26_pri_out[3] ) );
INV_X4 _u10_u0_u26_U6  ( .A(1'b1), .ZN(_u10_u0_u26_pri_out[2] ) );
INV_X4 _u10_u0_u26_U4  ( .A(1'b1), .ZN(_u10_u0_u26_pri_out[1] ) );
INV_X4 _u10_u0_u26_U2  ( .A(1'b1), .ZN(_u10_u0_u26_pri_out[0] ) );
INV_X4 _u10_u0_u27_U16  ( .A(1'b1), .ZN(_u10_u0_u27_pri_out[7] ) );
INV_X4 _u10_u0_u27_U14  ( .A(1'b1), .ZN(_u10_u0_u27_pri_out[6] ) );
INV_X4 _u10_u0_u27_U12  ( .A(1'b1), .ZN(_u10_u0_u27_pri_out[5] ) );
INV_X4 _u10_u0_u27_U10  ( .A(1'b1), .ZN(_u10_u0_u27_pri_out[4] ) );
INV_X4 _u10_u0_u27_U8  ( .A(1'b1), .ZN(_u10_u0_u27_pri_out[3] ) );
INV_X4 _u10_u0_u27_U6  ( .A(1'b1), .ZN(_u10_u0_u27_pri_out[2] ) );
INV_X4 _u10_u0_u27_U4  ( .A(1'b1), .ZN(_u10_u0_u27_pri_out[1] ) );
INV_X4 _u10_u0_u27_U2  ( .A(1'b1), .ZN(_u10_u0_u27_pri_out[0] ) );
INV_X4 _u10_u0_u28_U16  ( .A(1'b1), .ZN(_u10_u0_u28_pri_out[7] ) );
INV_X4 _u10_u0_u28_U14  ( .A(1'b1), .ZN(_u10_u0_u28_pri_out[6] ) );
INV_X4 _u10_u0_u28_U12  ( .A(1'b1), .ZN(_u10_u0_u28_pri_out[5] ) );
INV_X4 _u10_u0_u28_U10  ( .A(1'b1), .ZN(_u10_u0_u28_pri_out[4] ) );
INV_X4 _u10_u0_u28_U8  ( .A(1'b1), .ZN(_u10_u0_u28_pri_out[3] ) );
INV_X4 _u10_u0_u28_U6  ( .A(1'b1), .ZN(_u10_u0_u28_pri_out[2] ) );
INV_X4 _u10_u0_u28_U4  ( .A(1'b1), .ZN(_u10_u0_u28_pri_out[1] ) );
INV_X4 _u10_u0_u28_U2  ( .A(1'b1), .ZN(_u10_u0_u28_pri_out[0] ) );
INV_X4 _u10_u0_u29_U16  ( .A(1'b1), .ZN(_u10_u0_u29_pri_out[7] ) );
INV_X4 _u10_u0_u29_U14  ( .A(1'b1), .ZN(_u10_u0_u29_pri_out[6] ) );
INV_X4 _u10_u0_u29_U12  ( .A(1'b1), .ZN(_u10_u0_u29_pri_out[5] ) );
INV_X4 _u10_u0_u29_U10  ( .A(1'b1), .ZN(_u10_u0_u29_pri_out[4] ) );
INV_X4 _u10_u0_u29_U8  ( .A(1'b1), .ZN(_u10_u0_u29_pri_out[3] ) );
INV_X4 _u10_u0_u29_U6  ( .A(1'b1), .ZN(_u10_u0_u29_pri_out[2] ) );
INV_X4 _u10_u0_u29_U4  ( .A(1'b1), .ZN(_u10_u0_u29_pri_out[1] ) );
INV_X4 _u10_u0_u29_U2  ( .A(1'b1), .ZN(_u10_u0_u29_pri_out[0] ) );
INV_X4 _u10_u0_u30_U16  ( .A(1'b1), .ZN(_u10_u0_u30_pri_out[7] ) );
INV_X4 _u10_u0_u30_U14  ( .A(1'b1), .ZN(_u10_u0_u30_pri_out[6] ) );
INV_X4 _u10_u0_u30_U12  ( .A(1'b1), .ZN(_u10_u0_u30_pri_out[5] ) );
INV_X4 _u10_u0_u30_U10  ( .A(1'b1), .ZN(_u10_u0_u30_pri_out[4] ) );
INV_X4 _u10_u0_u30_U8  ( .A(1'b1), .ZN(_u10_u0_u30_pri_out[3] ) );
INV_X4 _u10_u0_u30_U6  ( .A(1'b1), .ZN(_u10_u0_u30_pri_out[2] ) );
INV_X4 _u10_u0_u30_U4  ( .A(1'b1), .ZN(_u10_u0_u30_pri_out[1] ) );
INV_X4 _u10_u0_u30_U2  ( .A(1'b1), .ZN(_u10_u0_u30_pri_out[0] ) );
INV_X1 _u10_u1_U1603  ( .A(1'b0), .ZN(_u10_u1_n2136 ) );
INV_X1 _u10_u1_U1602  ( .A(1'b0), .ZN(_u10_u1_n2139 ) );
NAND2_X1 _u10_u1_U1601  ( .A1(_u10_u1_n2136 ), .A2(_u10_u1_n2139 ), .ZN(_u10_u1_n2435 ) );
INV_X1 _u10_u1_U1600  ( .A(_u10_u1_n2435 ), .ZN(_u10_u1_n2483 ) );
INV_X1 _u10_u1_U1599  ( .A(1'b0), .ZN(_u10_u1_n2014 ) );
INV_X1 _u10_u1_U1598  ( .A(1'b0), .ZN(_u10_u1_n1844 ) );
NAND2_X1 _u10_u1_U1597  ( .A1(_u10_u1_n2014 ), .A2(_u10_u1_n1844 ), .ZN(_u10_u1_n2650 ) );
INV_X1 _u10_u1_U1596  ( .A(_u10_u1_n2650 ), .ZN(_u10_u1_n2023 ) );
INV_X1 _u10_u1_U1595  ( .A(1'b0), .ZN(_u10_u1_n2022 ) );
NAND2_X1 _u10_u1_U1594  ( .A1(_u10_u1_n2023 ), .A2(_u10_u1_n2022 ), .ZN(_u10_u1_n3278 ) );
INV_X1 _u10_u1_U1593  ( .A(_u10_u1_n3278 ), .ZN(_u10_u1_n3356 ) );
INV_X1 _u10_u1_U1592  ( .A(1'b0), .ZN(_u10_u1_n2068 ) );
INV_X1 _u10_u1_U1591  ( .A(1'b0), .ZN(_u10_u1_n2065 ) );
NAND2_X1 _u10_u1_U1590  ( .A1(_u10_u1_n2068 ), .A2(_u10_u1_n2065 ), .ZN(_u10_u1_n2287 ) );
INV_X1 _u10_u1_U1589  ( .A(_u10_u1_n2287 ), .ZN(_u10_u1_n2074 ) );
INV_X1 _u10_u1_U1588  ( .A(1'b0), .ZN(_u10_u1_n3024 ) );
INV_X1 _u10_u1_U1587  ( .A(1'b0), .ZN(_u10_u1_n1875 ) );
INV_X1 _u10_u1_U1586  ( .A(1'b0), .ZN(_u10_u1_n1857 ) );
NAND2_X1 _u10_u1_U1585  ( .A1(_u10_u1_n1875 ), .A2(_u10_u1_n1857 ), .ZN(_u10_u1_n2225 ) );
INV_X1 _u10_u1_U1584  ( .A(_u10_u1_n2225 ), .ZN(_u10_u1_n2990 ) );
INV_X1 _u10_u1_U1583  ( .A(1'b0), .ZN(_u10_u1_n1849 ) );
NAND2_X1 _u10_u1_U1582  ( .A1(_u10_u1_n2990 ), .A2(_u10_u1_n1849 ), .ZN(_u10_u1_n2216 ) );
INV_X1 _u10_u1_U1581  ( .A(_u10_u1_n2216 ), .ZN(_u10_u1_n2439 ) );
NAND3_X1 _u10_u1_U1580  ( .A1(_u10_u1_n2074 ), .A2(_u10_u1_n3024 ), .A3(_u10_u1_n2439 ), .ZN(_u10_u1_n2888 ) );
INV_X1 _u10_u1_U1579  ( .A(_u10_u1_n2888 ), .ZN(_u10_u1_n2380 ) );
INV_X1 _u10_u1_U1578  ( .A(1'b0), .ZN(_u10_u1_n2418 ) );
NAND2_X1 _u10_u1_U1577  ( .A1(_u10_u1_n2380 ), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n2960 ) );
INV_X1 _u10_u1_U1576  ( .A(_u10_u1_n2960 ), .ZN(_u10_u1_n2398 ) );
INV_X1 _u10_u1_U1575  ( .A(1'b0), .ZN(_u10_u1_n2878 ) );
INV_X1 _u10_u1_U1574  ( .A(1'b0), .ZN(_u10_u1_n2495 ) );
NAND2_X1 _u10_u1_U1573  ( .A1(_u10_u1_n2878 ), .A2(_u10_u1_n2495 ), .ZN(_u10_u1_n3060 ) );
INV_X1 _u10_u1_U1572  ( .A(_u10_u1_n3060 ), .ZN(_u10_u1_n3316 ) );
INV_X1 _u10_u1_U1571  ( .A(1'b0), .ZN(_u10_u1_n1907 ) );
NAND2_X1 _u10_u1_U1570  ( .A1(_u10_u1_n3316 ), .A2(_u10_u1_n1907 ), .ZN(_u10_u1_n2482 ) );
INV_X1 _u10_u1_U1569  ( .A(_u10_u1_n2482 ), .ZN(_u10_u1_n1894 ) );
INV_X1 _u10_u1_U1568  ( .A(1'b0), .ZN(_u10_u1_n1892 ) );
INV_X1 _u10_u1_U1567  ( .A(1'b0), .ZN(_u10_u1_n2619 ) );
NAND2_X1 _u10_u1_U1566  ( .A1(_u10_u1_n1892 ), .A2(_u10_u1_n2619 ), .ZN(_u10_u1_n2780 ) );
INV_X1 _u10_u1_U1565  ( .A(_u10_u1_n2780 ), .ZN(_u10_u1_n2294 ) );
NAND2_X1 _u10_u1_U1564  ( .A1(_u10_u1_n1894 ), .A2(_u10_u1_n2294 ), .ZN(_u10_u1_n2157 ) );
INV_X1 _u10_u1_U1563  ( .A(_u10_u1_n2157 ), .ZN(_u10_u1_n2815 ) );
INV_X1 _u10_u1_U1562  ( .A(1'b0), .ZN(_u10_u1_n1955 ) );
INV_X1 _u10_u1_U1561  ( .A(1'b0), .ZN(_u10_u1_n2063 ) );
NAND2_X1 _u10_u1_U1560  ( .A1(_u10_u1_n1955 ), .A2(_u10_u1_n2063 ), .ZN(_u10_u1_n2694 ) );
INV_X1 _u10_u1_U1559  ( .A(_u10_u1_n2694 ), .ZN(_u10_u1_n2105 ) );
INV_X1 _u10_u1_U1558  ( .A(1'b0), .ZN(_u10_u1_n2106 ) );
NAND2_X1 _u10_u1_U1557  ( .A1(_u10_u1_n2105 ), .A2(_u10_u1_n2106 ), .ZN(_u10_u1_n2574 ) );
INV_X1 _u10_u1_U1556  ( .A(1'b0), .ZN(_u10_u1_n2740 ) );
INV_X1 _u10_u1_U1555  ( .A(1'b0), .ZN(_u10_u1_n2155 ) );
NAND2_X1 _u10_u1_U1554  ( .A1(_u10_u1_n2740 ), .A2(_u10_u1_n2155 ), .ZN(_u10_u1_n2268 ) );
NOR2_X1 _u10_u1_U1553  ( .A1(_u10_u1_n2574 ), .A2(_u10_u1_n2268 ), .ZN(_u10_u1_n1885 ) );
INV_X1 _u10_u1_U1552  ( .A(_u10_req_p0_0_ ), .ZN(_u10_u1_n1845 ) );
INV_X1 _u10_u1_U1551  ( .A(1'b0), .ZN(_u10_u1_n2043 ) );
NAND2_X1 _u10_u1_U1550  ( .A1(_u10_u1_n1845 ), .A2(_u10_u1_n2043 ), .ZN(_u10_u1_n3086 ) );
INV_X1 _u10_u1_U1549  ( .A(_u10_u1_n3086 ), .ZN(_u10_u1_n3065 ) );
NAND2_X1 _u10_u1_U1548  ( .A1(1'b0), .A2(_u10_u1_n3065 ), .ZN(_u10_u1_n3358 ) );
INV_X1 _u10_u1_U1547  ( .A(_u10_u1_n3358 ), .ZN(_u10_u1_n3073 ) );
NAND3_X1 _u10_u1_U1546  ( .A1(_u10_u1_n2815 ), .A2(_u10_u1_n1885 ), .A3(_u10_u1_n3073 ), .ZN(_u10_u1_n3087 ) );
INV_X1 _u10_u1_U1545  ( .A(_u10_u1_n3087 ), .ZN(_u10_u1_n3134 ) );
NAND3_X1 _u10_u1_U1544  ( .A1(_u10_u1_n3356 ), .A2(_u10_u1_n2398 ), .A3(_u10_u1_n3134 ), .ZN(_u10_u1_n3408 ) );
INV_X1 _u10_u1_U1543  ( .A(1'b0), .ZN(_u10_u1_n2017 ) );
NAND2_X1 _u10_u1_U1542  ( .A1(_u10_u1_n3408 ), .A2(_u10_u1_n2017 ), .ZN(_u10_u1_n3407 ) );
AND2_X1 _u10_u1_U1541  ( .A1(_u10_u1_n2483 ), .A2(_u10_u1_n3407 ), .ZN(_u10_u1_n3390 ) );
NOR3_X1 _u10_u1_U1540  ( .A1(_u10_gnt_p0_d[3] ), .A2(_u10_gnt_p0_d[4] ),.A3(_u10_gnt_p0_d[0] ), .ZN(_u10_u1_n3391 ) );
NOR2_X1 _u10_u1_U1539  ( .A1(_u10_u1_n13 ), .A2(_u10_u1_n14 ), .ZN(_u10_u1_n3257 ) );
NAND2_X1 _u10_u1_U1538  ( .A1(_u10_u1_n3391 ), .A2(_u10_u1_n3257 ), .ZN(_u10_u1_n3248 ) );
NOR3_X1 _u10_u1_U1537  ( .A1(_u10_gnt_p0_d[4] ), .A2(_u10_u1_n15 ), .A3(_u10_gnt_p0_d[3] ), .ZN(_u10_u1_n3371 ) );
NAND2_X1 _u10_u1_U1536  ( .A1(_u10_u1_n3371 ), .A2(_u10_u1_n3257 ), .ZN(_u10_u1_n2932 ) );
NAND2_X1 _u10_u1_U1535  ( .A1(_u10_u1_n3248 ), .A2(_u10_u1_n2932 ), .ZN(_u10_u1_n2796 ) );
NAND2_X1 _u10_u1_U1534  ( .A1(_u10_u1_n3390 ), .A2(_u10_u1_n2796 ), .ZN(_u10_u1_n3375 ) );
NOR2_X1 _u10_u1_U1533  ( .A1(_u10_u1_n12 ), .A2(_u10_u1_n10 ), .ZN(_u10_u1_n3369 ) );
AND2_X1 _u10_u1_U1532  ( .A1(_u10_u1_n3369 ), .A2(_u10_u1_n15 ), .ZN(_u10_u1_n3355 ) );
NOR2_X1 _u10_u1_U1531  ( .A1(_u10_gnt_p0_d[2] ), .A2(_u10_u1_n14 ), .ZN(_u10_u1_n3298 ) );
NAND2_X1 _u10_u1_U1530  ( .A1(_u10_u1_n3355 ), .A2(_u10_u1_n3298 ), .ZN(_u10_u1_n2966 ) );
INV_X1 _u10_u1_U1529  ( .A(_u10_u1_n2966 ), .ZN(_u10_u1_n2146 ) );
NAND2_X1 _u10_u1_U1528  ( .A1(_u10_u1_n2483 ), .A2(_u10_u1_n2017 ), .ZN(_u10_u1_n2506 ) );
INV_X1 _u10_u1_U1527  ( .A(1'b0), .ZN(_u10_u1_n3007 ) );
INV_X1 _u10_u1_U1526  ( .A(1'b0), .ZN(_u10_u1_n1846 ) );
NAND2_X1 _u10_u1_U1525  ( .A1(_u10_u1_n3007 ), .A2(_u10_u1_n1846 ), .ZN(_u10_u1_n1933 ) );
INV_X1 _u10_u1_U1524  ( .A(_u10_u1_n1933 ), .ZN(_u10_u1_n2024 ) );
NAND2_X1 _u10_u1_U1523  ( .A1(_u10_u1_n3065 ), .A2(_u10_u1_n2024 ), .ZN(_u10_u1_n2663 ) );
INV_X1 _u10_u1_U1522  ( .A(_u10_u1_n2663 ), .ZN(_u10_u1_n2008 ) );
INV_X1 _u10_u1_U1521  ( .A(1'b0), .ZN(_u10_u1_n3033 ) );
INV_X1 _u10_u1_U1520  ( .A(1'b0), .ZN(_u10_u1_n1903 ) );
NAND2_X1 _u10_u1_U1519  ( .A1(_u10_u1_n3033 ), .A2(_u10_u1_n1903 ), .ZN(_u10_u1_n2861 ) );
NOR2_X1 _u10_u1_U1518  ( .A1(_u10_u1_n2861 ), .A2(1'b0), .ZN(_u10_u1_n2662 ));
INV_X1 _u10_u1_U1517  ( .A(1'b0), .ZN(_u10_u1_n2505 ) );
NAND2_X1 _u10_u1_U1516  ( .A1(_u10_u1_n2662 ), .A2(_u10_u1_n2505 ), .ZN(_u10_u1_n2621 ) );
INV_X1 _u10_u1_U1515  ( .A(_u10_u1_n2621 ), .ZN(_u10_u1_n2430 ) );
NAND2_X1 _u10_u1_U1514  ( .A1(_u10_u1_n2008 ), .A2(_u10_u1_n2430 ), .ZN(_u10_u1_n2007 ) );
NOR3_X1 _u10_u1_U1513  ( .A1(_u10_u1_n2506 ), .A2(1'b0), .A3(_u10_u1_n2007 ),.ZN(_u10_u1_n1843 ) );
NAND2_X1 _u10_u1_U1512  ( .A1(_u10_u1_n1843 ), .A2(_u10_u1_n2023 ), .ZN(_u10_u1_n1919 ) );
INV_X1 _u10_u1_U1511  ( .A(_u10_u1_n1919 ), .ZN(_u10_u1_n2354 ) );
NAND3_X1 _u10_u1_U1510  ( .A1(_u10_u1_n2878 ), .A2(_u10_u1_n1907 ), .A3(_u10_u1_n2354 ), .ZN(_u10_u1_n2010 ) );
INV_X1 _u10_u1_U1509  ( .A(_u10_u1_n2010 ), .ZN(_u10_u1_n2227 ) );
NAND2_X1 _u10_u1_U1508  ( .A1(_u10_u1_n2227 ), .A2(_u10_u1_n2495 ), .ZN(_u10_u1_n2478 ) );
INV_X1 _u10_u1_U1507  ( .A(_u10_u1_n2478 ), .ZN(_u10_u1_n2486 ) );
NAND2_X1 _u10_u1_U1506  ( .A1(_u10_u1_n2486 ), .A2(_u10_u1_n1892 ), .ZN(_u10_u1_n1895 ) );
INV_X1 _u10_u1_U1505  ( .A(_u10_u1_n1895 ), .ZN(_u10_u1_n2295 ) );
NAND2_X1 _u10_u1_U1504  ( .A1(1'b0), .A2(_u10_u1_n2990 ), .ZN(_u10_u1_n3406 ) );
NAND2_X1 _u10_u1_U1503  ( .A1(_u10_u1_n2418 ), .A2(_u10_u1_n3406 ), .ZN(_u10_u1_n3101 ) );
NAND2_X1 _u10_u1_U1502  ( .A1(1'b0), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n2045 ) );
INV_X1 _u10_u1_U1501  ( .A(_u10_u1_n2045 ), .ZN(_u10_u1_n2133 ) );
NOR2_X1 _u10_u1_U1500  ( .A1(_u10_u1_n3101 ), .A2(_u10_u1_n2133 ), .ZN(_u10_u1_n3373 ) );
NOR2_X1 _u10_u1_U1499  ( .A1(_u10_u1_n2065 ), .A2(_u10_u1_n2216 ), .ZN(_u10_u1_n3340 ) );
NAND2_X1 _u10_u1_U1498  ( .A1(_u10_u1_n3024 ), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n2314 ) );
INV_X1 _u10_u1_U1497  ( .A(_u10_u1_n2314 ), .ZN(_u10_u1_n2209 ) );
NAND2_X1 _u10_u1_U1496  ( .A1(_u10_u1_n3340 ), .A2(_u10_u1_n2209 ), .ZN(_u10_u1_n2356 ) );
NAND2_X1 _u10_u1_U1495  ( .A1(_u10_u1_n3373 ), .A2(_u10_u1_n2356 ), .ZN(_u10_u1_n3405 ) );
NAND2_X1 _u10_u1_U1494  ( .A1(_u10_u1_n2295 ), .A2(_u10_u1_n3405 ), .ZN(_u10_u1_n3404 ) );
NAND2_X1 _u10_u1_U1493  ( .A1(1'b0), .A2(_u10_u1_n2662 ), .ZN(_u10_u1_n1929 ) );
NOR2_X1 _u10_u1_U1492  ( .A1(_u10_u1_n1929 ), .A2(_u10_u1_n2663 ), .ZN(_u10_u1_n1916 ) );
NAND2_X1 _u10_u1_U1491  ( .A1(_u10_u1_n1916 ), .A2(_u10_u1_n1894 ), .ZN(_u10_u1_n2974 ) );
INV_X1 _u10_u1_U1490  ( .A(_u10_u1_n2506 ), .ZN(_u10_u1_n2370 ) );
NAND2_X1 _u10_u1_U1489  ( .A1(1'b0), .A2(_u10_u1_n2370 ), .ZN(_u10_u1_n1979 ) );
NOR3_X1 _u10_u1_U1488  ( .A1(_u10_u1_n2007 ), .A2(1'b0), .A3(_u10_u1_n1979 ),.ZN(_u10_u1_n2608 ) );
NAND2_X1 _u10_u1_U1487  ( .A1(_u10_u1_n3316 ), .A2(_u10_u1_n2608 ), .ZN(_u10_u1_n1891 ) );
INV_X1 _u10_u1_U1486  ( .A(_u10_u1_n1891 ), .ZN(_u10_u1_n3343 ) );
NOR3_X1 _u10_u1_U1485  ( .A1(_u10_u1_n2007 ), .A2(_u10_u1_n2435 ), .A3(_u10_u1_n2017 ), .ZN(_u10_u1_n3157 ) );
AND2_X1 _u10_u1_U1484  ( .A1(_u10_u1_n3157 ), .A2(_u10_u1_n1894 ), .ZN(_u10_u1_n3056 ) );
NOR2_X1 _u10_u1_U1483  ( .A1(_u10_u1_n3343 ), .A2(_u10_u1_n3056 ), .ZN(_u10_u1_n2471 ) );
NAND3_X1 _u10_u1_U1482  ( .A1(_u10_u1_n3404 ), .A2(_u10_u1_n2974 ), .A3(_u10_u1_n2471 ), .ZN(_u10_u1_n3403 ) );
NAND2_X1 _u10_u1_U1481  ( .A1(_u10_u1_n2146 ), .A2(_u10_u1_n3403 ), .ZN(_u10_u1_n3376 ) );
NOR3_X1 _u10_u1_U1480  ( .A1(_u10_gnt_p0_d[4] ), .A2(_u10_u1_n12 ), .A3(_u10_gnt_p0_d[0] ), .ZN(_u10_u1_n3297 ) );
NAND2_X1 _u10_u1_U1479  ( .A1(_u10_u1_n3297 ), .A2(_u10_u1_n3298 ), .ZN(_u10_u1_n3195 ) );
INV_X1 _u10_u1_U1478  ( .A(_u10_u1_n3195 ), .ZN(_u10_u1_n2012 ) );
NAND3_X1 _u10_u1_U1477  ( .A1(_u10_u1_n2398 ), .A2(_u10_u1_n2023 ), .A3(_u10_u1_n3134 ), .ZN(_u10_u1_n3402 ) );
NAND2_X1 _u10_u1_U1476  ( .A1(_u10_u1_n2022 ), .A2(_u10_u1_n3402 ), .ZN(_u10_u1_n3131 ) );
NAND2_X1 _u10_u1_U1475  ( .A1(_u10_u1_n2012 ), .A2(_u10_u1_n3131 ), .ZN(_u10_u1_n3377 ) );
NAND2_X1 _u10_u1_U1474  ( .A1(_u10_u1_n3391 ), .A2(_u10_u1_n3298 ), .ZN(_u10_u1_n3143 ) );
NAND2_X1 _u10_u1_U1473  ( .A1(_u10_u1_n3356 ), .A2(_u10_u1_n2017 ), .ZN(_u10_u1_n2632 ) );
INV_X1 _u10_u1_U1472  ( .A(_u10_u1_n2632 ), .ZN(_u10_u1_n2140 ) );
NAND2_X1 _u10_u1_U1471  ( .A1(_u10_u1_n2140 ), .A2(_u10_u1_n2483 ), .ZN(_u10_u1_n2811 ) );
INV_X1 _u10_u1_U1470  ( .A(_u10_u1_n2811 ), .ZN(_u10_u1_n3227 ) );
NAND2_X1 _u10_u1_U1469  ( .A1(_u10_u1_n3227 ), .A2(_u10_u1_n2505 ), .ZN(_u10_u1_n2979 ) );
NOR2_X1 _u10_u1_U1468  ( .A1(_u10_u1_n2979 ), .A2(1'b0), .ZN(_u10_u1_n1904 ));
INV_X1 _u10_u1_U1467  ( .A(_u10_u1_n2861 ), .ZN(_u10_u1_n2837 ) );
NAND2_X1 _u10_u1_U1466  ( .A1(_u10_u1_n1904 ), .A2(_u10_u1_n2837 ), .ZN(_u10_u1_n2131 ) );
NOR3_X1 _u10_u1_U1465  ( .A1(_u10_u1_n3143 ), .A2(1'b0), .A3(_u10_u1_n2131 ),.ZN(_u10_u1_n3155 ) );
NOR2_X1 _u10_u1_U1464  ( .A1(_u10_gnt_p0_d[1] ), .A2(_u10_gnt_p0_d[2] ),.ZN(_u10_u1_n3149 ) );
NAND2_X1 _u10_u1_U1463  ( .A1(_u10_u1_n3391 ), .A2(_u10_u1_n3149 ), .ZN(_u10_u1_n2042 ) );
NOR4_X1 _u10_u1_U1462  ( .A1(_u10_u1_n2131 ), .A2(_u10_u1_n1933 ), .A3(_u10_u1_n2042 ), .A4(1'b0), .ZN(_u10_u1_n3401 ) );
NOR2_X1 _u10_u1_U1461  ( .A1(_u10_u1_n3155 ), .A2(_u10_u1_n3401 ), .ZN(_u10_u1_n2274 ) );
NAND2_X1 _u10_u1_U1460  ( .A1(_u10_u1_n3371 ), .A2(_u10_u1_n3149 ), .ZN(_u10_u1_n3027 ) );
NOR3_X1 _u10_u1_U1459  ( .A1(_u10_u1_n1933 ), .A2(_u10_u1_n3027 ), .A3(_u10_u1_n2131 ), .ZN(_u10_u1_n2299 ) );
INV_X1 _u10_u1_U1458  ( .A(_u10_u1_n2299 ), .ZN(_u10_u1_n1935 ) );
NAND2_X1 _u10_u1_U1457  ( .A1(_u10_u1_n2274 ), .A2(_u10_u1_n1935 ), .ZN(_u10_u1_n2826 ) );
NAND2_X1 _u10_u1_U1456  ( .A1(_u10_u1_n3369 ), .A2(_u10_u1_n3257 ), .ZN(_u10_u1_n2353 ) );
INV_X1 _u10_u1_U1455  ( .A(_u10_u1_n2353 ), .ZN(_u10_u1_n1837 ) );
NAND2_X1 _u10_u1_U1454  ( .A1(_u10_u1_n2354 ), .A2(_u10_u1_n1837 ), .ZN(_u10_u1_n2877 ) );
INV_X1 _u10_u1_U1453  ( .A(_u10_u1_n2877 ), .ZN(_u10_u1_n2631 ) );
NOR2_X1 _u10_u1_U1452  ( .A1(_u10_u1_n2826 ), .A2(_u10_u1_n2631 ), .ZN(_u10_u1_n2219 ) );
NOR2_X1 _u10_u1_U1451  ( .A1(_u10_u1_n2219 ), .A2(_u10_u1_n2356 ), .ZN(_u10_u1_n3379 ) );
NAND3_X1 _u10_u1_U1450  ( .A1(_u10_u1_n2008 ), .A2(_u10_u1_n2837 ), .A3(1'b0), .ZN(_u10_u1_n2725 ) );
INV_X1 _u10_u1_U1449  ( .A(_u10_u1_n2725 ), .ZN(_u10_u1_n2836 ) );
INV_X1 _u10_u1_U1448  ( .A(_u10_u1_n2268 ), .ZN(_u10_u1_n1963 ) );
NAND2_X1 _u10_u1_U1447  ( .A1(_u10_u1_n2815 ), .A2(_u10_u1_n1963 ), .ZN(_u10_u1_n3365 ) );
INV_X1 _u10_u1_U1446  ( .A(_u10_u1_n3365 ), .ZN(_u10_u1_n2804 ) );
NAND2_X1 _u10_u1_U1445  ( .A1(_u10_u1_n2836 ), .A2(_u10_u1_n2804 ), .ZN(_u10_u1_n2769 ) );
INV_X1 _u10_u1_U1444  ( .A(_u10_u1_n2769 ), .ZN(_u10_u1_n2778 ) );
NAND2_X1 _u10_u1_U1443  ( .A1(_u10_u1_n1894 ), .A2(_u10_u1_n1892 ), .ZN(_u10_u1_n2620 ) );
NOR2_X1 _u10_u1_U1442  ( .A1(_u10_u1_n2620 ), .A2(_u10_u1_n3358 ), .ZN(_u10_u1_n3400 ) );
NOR2_X1 _u10_u1_U1441  ( .A1(_u10_u1_n3400 ), .A2(1'b0), .ZN(_u10_u1_n3399 ));
NOR2_X1 _u10_u1_U1440  ( .A1(_u10_u1_n3399 ), .A2(_u10_u1_n2268 ), .ZN(_u10_u1_n3393 ) );
INV_X1 _u10_u1_U1439  ( .A(_u10_u1_n2356 ), .ZN(_u10_u1_n2046 ) );
NAND3_X1 _u10_u1_U1438  ( .A1(_u10_u1_n2990 ), .A2(_u10_u1_n2209 ), .A3(1'b0), .ZN(_u10_u1_n3243 ) );
INV_X1 _u10_u1_U1437  ( .A(_u10_u1_n3243 ), .ZN(_u10_u1_n2170 ) );
NOR2_X1 _u10_u1_U1436  ( .A1(_u10_u1_n2046 ), .A2(_u10_u1_n2170 ), .ZN(_u10_u1_n3091 ) );
NOR2_X1 _u10_u1_U1435  ( .A1(_u10_u1_n1895 ), .A2(1'b0), .ZN(_u10_u1_n2397 ));
NAND2_X1 _u10_u1_U1434  ( .A1(_u10_u1_n2397 ), .A2(_u10_u1_n2740 ), .ZN(_u10_u1_n2989 ) );
INV_X1 _u10_u1_U1433  ( .A(_u10_u1_n2989 ), .ZN(_u10_u1_n2522 ) );
NAND2_X1 _u10_u1_U1432  ( .A1(_u10_u1_n2522 ), .A2(_u10_u1_n2155 ), .ZN(_u10_u1_n2315 ) );
NOR2_X1 _u10_u1_U1431  ( .A1(_u10_u1_n3091 ), .A2(_u10_u1_n2315 ), .ZN(_u10_u1_n3394 ) );
INV_X1 _u10_u1_U1430  ( .A(_u10_u1_n2315 ), .ZN(_u10_u1_n2152 ) );
NAND2_X1 _u10_u1_U1429  ( .A1(1'b0), .A2(_u10_u1_n2152 ), .ZN(_u10_u1_n3396 ) );
NOR3_X1 _u10_u1_U1428  ( .A1(_u10_u1_n3060 ), .A2(1'b0), .A3(_u10_u1_n1907 ),.ZN(_u10_u1_n2497 ) );
NAND2_X1 _u10_u1_U1427  ( .A1(_u10_u1_n2497 ), .A2(_u10_u1_n2619 ), .ZN(_u10_u1_n2293 ) );
NOR2_X1 _u10_u1_U1426  ( .A1(_u10_u1_n2293 ), .A2(1'b0), .ZN(_u10_u1_n2312 ));
INV_X1 _u10_u1_U1425  ( .A(_u10_u1_n2312 ), .ZN(_u10_u1_n2737 ) );
NAND2_X1 _u10_u1_U1424  ( .A1(_u10_u1_n2133 ), .A2(_u10_u1_n2522 ), .ZN(_u10_u1_n3398 ) );
NAND2_X1 _u10_u1_U1423  ( .A1(_u10_u1_n2737 ), .A2(_u10_u1_n3398 ), .ZN(_u10_u1_n3386 ) );
NAND2_X1 _u10_u1_U1422  ( .A1(_u10_u1_n3386 ), .A2(_u10_u1_n2155 ), .ZN(_u10_u1_n3397 ) );
AND2_X1 _u10_u1_U1421  ( .A1(_u10_u1_n3396 ), .A2(_u10_u1_n3397 ), .ZN(_u10_u1_n2774 ) );
NAND2_X1 _u10_u1_U1420  ( .A1(_u10_u1_n3056 ), .A2(_u10_u1_n2740 ), .ZN(_u10_u1_n2526 ) );
INV_X1 _u10_u1_U1419  ( .A(_u10_u1_n2526 ), .ZN(_u10_u1_n3307 ) );
NAND2_X1 _u10_u1_U1418  ( .A1(_u10_u1_n3307 ), .A2(_u10_u1_n2155 ), .ZN(_u10_u1_n3395 ) );
NAND2_X1 _u10_u1_U1417  ( .A1(_u10_u1_n2774 ), .A2(_u10_u1_n3395 ), .ZN(_u10_u1_n2531 ) );
NOR4_X1 _u10_u1_U1416  ( .A1(_u10_u1_n2778 ), .A2(_u10_u1_n3393 ), .A3(_u10_u1_n3394 ), .A4(_u10_u1_n2531 ), .ZN(_u10_u1_n3392 ) );
NAND3_X1 _u10_u1_U1415  ( .A1(_u10_gnt_p0_d[4] ), .A2(_u10_gnt_p0_d[0] ),.A3(_u10_u1_n3257 ), .ZN(_u10_u1_n2529 ) );
NOR2_X1 _u10_u1_U1414  ( .A1(_u10_u1_n3392 ), .A2(_u10_u1_n2529 ), .ZN(_u10_u1_n3380 ) );
NOR2_X1 _u10_u1_U1413  ( .A1(_u10_gnt_p0_d[1] ), .A2(_u10_u1_n13 ), .ZN(_u10_u1_n3324 ) );
NAND2_X1 _u10_u1_U1412  ( .A1(_u10_u1_n3324 ), .A2(_u10_u1_n3371 ), .ZN(_u10_u1_n2868 ) );
INV_X1 _u10_u1_U1411  ( .A(_u10_u1_n2868 ), .ZN(_u10_u1_n2703 ) );
AND2_X1 _u10_u1_U1410  ( .A1(_u10_u1_n3391 ), .A2(_u10_u1_n3324 ), .ZN(_u10_u1_n2702 ) );
NAND2_X1 _u10_u1_U1409  ( .A1(_u10_u1_n2702 ), .A2(_u10_u1_n3033 ), .ZN(_u10_u1_n2869 ) );
INV_X1 _u10_u1_U1408  ( .A(_u10_u1_n2869 ), .ZN(_u10_u1_n3372 ) );
NOR2_X1 _u10_u1_U1407  ( .A1(_u10_u1_n2703 ), .A2(_u10_u1_n3372 ), .ZN(_u10_u1_n2400 ) );
INV_X1 _u10_u1_U1406  ( .A(_u10_u1_n1979 ), .ZN(_u10_u1_n2507 ) );
NAND3_X1 _u10_u1_U1405  ( .A1(_u10_u1_n3065 ), .A2(_u10_u1_n1846 ), .A3(1'b0), .ZN(_u10_u1_n1912 ) );
INV_X1 _u10_u1_U1404  ( .A(_u10_u1_n1912 ), .ZN(_u10_u1_n1897 ) );
NAND3_X1 _u10_u1_U1403  ( .A1(_u10_u1_n1897 ), .A2(_u10_u1_n2105 ), .A3(_u10_u1_n2804 ), .ZN(_u10_u1_n2119 ) );
NOR3_X1 _u10_u1_U1402  ( .A1(_u10_u1_n2960 ), .A2(_u10_u1_n2650 ), .A3(_u10_u1_n2119 ), .ZN(_u10_u1_n3127 ) );
AND2_X1 _u10_u1_U1401  ( .A1(_u10_u1_n3127 ), .A2(_u10_u1_n2370 ), .ZN(_u10_u1_n1984 ) );
INV_X1 _u10_u1_U1400  ( .A(1'b0), .ZN(_u10_u1_n2867 ) );
NAND2_X1 _u10_u1_U1399  ( .A1(_u10_u1_n2505 ), .A2(_u10_u1_n2867 ), .ZN(_u10_u1_n1980 ) );
NOR4_X1 _u10_u1_U1398  ( .A1(_u10_u1_n2507 ), .A2(_u10_u1_n3390 ), .A3(_u10_u1_n1984 ), .A4(_u10_u1_n1980 ), .ZN(_u10_u1_n3389 ) );
NOR2_X1 _u10_u1_U1397  ( .A1(_u10_u1_n2400 ), .A2(_u10_u1_n3389 ), .ZN(_u10_u1_n3381 ) );
NOR2_X1 _u10_u1_U1396  ( .A1(_u10_u1_n2157 ), .A2(_u10_u1_n1912 ), .ZN(_u10_u1_n1833 ) );
NOR2_X1 _u10_u1_U1395  ( .A1(_u10_u1_n2482 ), .A2(_u10_u1_n3358 ), .ZN(_u10_u1_n3388 ) );
NOR3_X1 _u10_u1_U1394  ( .A1(_u10_u1_n1833 ), .A2(_u10_u1_n3343 ), .A3(_u10_u1_n3388 ), .ZN(_u10_u1_n3387 ) );
NOR2_X1 _u10_u1_U1393  ( .A1(1'b0), .A2(_u10_u1_n3387 ), .ZN(_u10_u1_n3384 ));
NAND2_X1 _u10_u1_U1392  ( .A1(_u10_u1_n2074 ), .A2(_u10_u1_n1849 ), .ZN(_u10_u1_n2198 ) );
INV_X1 _u10_u1_U1391  ( .A(_u10_u1_n2198 ), .ZN(_u10_u1_n1886 ) );
NAND3_X1 _u10_u1_U1390  ( .A1(_u10_u1_n1886 ), .A2(_u10_u1_n2063 ), .A3(1'b0), .ZN(_u10_u1_n2193 ) );
INV_X1 _u10_u1_U1389  ( .A(_u10_u1_n2193 ), .ZN(_u10_u1_n2666 ) );
NAND2_X1 _u10_u1_U1388  ( .A1(_u10_u1_n2666 ), .A2(_u10_u1_n1875 ), .ZN(_u10_u1_n2191 ) );
NAND2_X1 _u10_u1_U1387  ( .A1(_u10_u1_n2209 ), .A2(_u10_u1_n1857 ), .ZN(_u10_u1_n1883 ) );
NOR2_X1 _u10_u1_U1386  ( .A1(_u10_u1_n2191 ), .A2(_u10_u1_n1883 ), .ZN(_u10_u1_n2171 ) );
NOR2_X1 _u10_u1_U1385  ( .A1(_u10_u1_n2694 ), .A2(1'b0), .ZN(_u10_u1_n2265 ));
NAND2_X1 _u10_u1_U1384  ( .A1(1'b0), .A2(_u10_u1_n2265 ), .ZN(_u10_u1_n2072 ) );
NAND2_X1 _u10_u1_U1383  ( .A1(_u10_u1_n2065 ), .A2(_u10_u1_n1849 ), .ZN(_u10_u1_n2423 ) );
NOR2_X1 _u10_u1_U1382  ( .A1(_u10_u1_n2072 ), .A2(_u10_u1_n2423 ), .ZN(_u10_u1_n2202 ) );
NAND2_X1 _u10_u1_U1381  ( .A1(_u10_u1_n2202 ), .A2(_u10_u1_n1875 ), .ZN(_u10_u1_n2189 ) );
NOR2_X1 _u10_u1_U1380  ( .A1(_u10_u1_n2189 ), .A2(_u10_u1_n1883 ), .ZN(_u10_u1_n2912 ) );
NOR2_X1 _u10_u1_U1379  ( .A1(_u10_u1_n2171 ), .A2(_u10_u1_n2912 ), .ZN(_u10_u1_n3245 ) );
NOR2_X1 _u10_u1_U1378  ( .A1(_u10_u1_n3245 ), .A2(_u10_u1_n2989 ), .ZN(_u10_u1_n3385 ) );
NOR4_X1 _u10_u1_U1377  ( .A1(_u10_u1_n3307 ), .A2(_u10_u1_n3384 ), .A3(_u10_u1_n3385 ), .A4(_u10_u1_n3386 ), .ZN(_u10_u1_n3383 ) );
NAND2_X1 _u10_u1_U1376  ( .A1(_u10_u1_n3355 ), .A2(_u10_u1_n3149 ), .ZN(_u10_u1_n1830 ) );
NOR2_X1 _u10_u1_U1375  ( .A1(_u10_u1_n3383 ), .A2(_u10_u1_n1830 ), .ZN(_u10_u1_n3382 ) );
NOR4_X1 _u10_u1_U1374  ( .A1(_u10_u1_n3379 ), .A2(_u10_u1_n3380 ), .A3(_u10_u1_n3381 ), .A4(_u10_u1_n3382 ), .ZN(_u10_u1_n3378 ) );
NAND4_X1 _u10_u1_U1373  ( .A1(_u10_u1_n3375 ), .A2(_u10_u1_n3376 ), .A3(_u10_u1_n3377 ), .A4(_u10_u1_n3378 ), .ZN(_u10_u1_n3158 ) );
NAND3_X1 _u10_u1_U1372  ( .A1(_u10_u1_n1963 ), .A2(_u10_u1_n2106 ), .A3(1'b0), .ZN(_u10_u1_n2239 ) );
INV_X1 _u10_u1_U1371  ( .A(_u10_u1_n2239 ), .ZN(_u10_u1_n2269 ) );
NAND2_X1 _u10_u1_U1370  ( .A1(_u10_u1_n2269 ), .A2(_u10_u1_n2265 ), .ZN(_u10_u1_n2596 ) );
NOR2_X1 _u10_u1_U1369  ( .A1(_u10_u1_n2596 ), .A2(_u10_u1_n2423 ), .ZN(_u10_u1_n2203 ) );
INV_X1 _u10_u1_U1368  ( .A(_u10_u1_n2203 ), .ZN(_u10_u1_n3374 ) );
NOR3_X1 _u10_u1_U1367  ( .A1(_u10_u1_n1883 ), .A2(1'b0), .A3(_u10_u1_n3374 ),.ZN(_u10_u1_n2480 ) );
NOR2_X1 _u10_u1_U1366  ( .A1(_u10_u1_n2171 ), .A2(_u10_u1_n2480 ), .ZN(_u10_u1_n3070 ) );
NAND3_X1 _u10_u1_U1365  ( .A1(_u10_u1_n1963 ), .A2(_u10_u1_n2619 ), .A3(1'b0), .ZN(_u10_u1_n3183 ) );
NOR2_X1 _u10_u1_U1364  ( .A1(_u10_u1_n3183 ), .A2(1'b0), .ZN(_u10_u1_n2407 ));
NAND2_X1 _u10_u1_U1363  ( .A1(_u10_u1_n2407 ), .A2(_u10_u1_n1955 ), .ZN(_u10_u1_n2240 ) );
INV_X1 _u10_u1_U1362  ( .A(_u10_u1_n2240 ), .ZN(_u10_u1_n3361 ) );
NAND3_X1 _u10_u1_U1361  ( .A1(_u10_u1_n2068 ), .A2(_u10_u1_n2063 ), .A3(_u10_u1_n3361 ), .ZN(_u10_u1_n2597 ) );
INV_X1 _u10_u1_U1360  ( .A(_u10_u1_n2597 ), .ZN(_u10_u1_n3093 ) );
INV_X1 _u10_u1_U1359  ( .A(_u10_u1_n2423 ), .ZN(_u10_u1_n2201 ) );
NAND3_X1 _u10_u1_U1358  ( .A1(_u10_u1_n3093 ), .A2(_u10_u1_n1875 ), .A3(_u10_u1_n2201 ), .ZN(_u10_u1_n1949 ) );
NOR2_X1 _u10_u1_U1357  ( .A1(_u10_u1_n1883 ), .A2(_u10_u1_n1949 ), .ZN(_u10_u1_n3125 ) );
NOR3_X1 _u10_u1_U1356  ( .A1(_u10_u1_n3125 ), .A2(_u10_u1_n2912 ), .A3(_u10_u1_n2046 ), .ZN(_u10_u1_n2345 ) );
NOR2_X1 _u10_u1_U1355  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u1_n2618 ) );
NAND2_X1 _u10_u1_U1354  ( .A1(_u10_u1_n2312 ), .A2(_u10_u1_n2618 ), .ZN(_u10_u1_n2403 ) );
NOR2_X1 _u10_u1_U1353  ( .A1(_u10_u1_n2403 ), .A2(1'b0), .ZN(_u10_u1_n2553 ));
NAND3_X1 _u10_u1_U1352  ( .A1(_u10_u1_n1886 ), .A2(_u10_u1_n2063 ), .A3(_u10_u1_n2553 ), .ZN(_u10_u1_n2588 ) );
NOR3_X1 _u10_u1_U1351  ( .A1(_u10_u1_n1883 ), .A2(1'b0), .A3(_u10_u1_n2588 ),.ZN(_u10_u1_n2887 ) );
INV_X1 _u10_u1_U1350  ( .A(_u10_u1_n2887 ), .ZN(_u10_u1_n2277 ) );
NAND4_X1 _u10_u1_U1349  ( .A1(_u10_u1_n3070 ), .A2(_u10_u1_n3373 ), .A3(_u10_u1_n2345 ), .A4(_u10_u1_n2277 ), .ZN(_u10_u1_n3370 ) );
NAND2_X1 _u10_u1_U1348  ( .A1(_u10_u1_n3372 ), .A2(_u10_u1_n1904 ), .ZN(_u10_u1_n2346 ) );
NAND2_X1 _u10_u1_U1347  ( .A1(_u10_u1_n1904 ), .A2(_u10_u1_n2703 ), .ZN(_u10_u1_n2343 ) );
AND2_X1 _u10_u1_U1346  ( .A1(_u10_u1_n2346 ), .A2(_u10_u1_n2343 ), .ZN(_u10_u1_n1868 ) );
NAND2_X1 _u10_u1_U1345  ( .A1(_u10_u1_n3298 ), .A2(_u10_u1_n3371 ), .ZN(_u10_u1_n2127 ) );
OR2_X1 _u10_u1_U1344  ( .A1(_u10_u1_n2131 ), .A2(_u10_u1_n2127 ), .ZN(_u10_u1_n2250 ) );
NAND2_X1 _u10_u1_U1343  ( .A1(_u10_u1_n1868 ), .A2(_u10_u1_n2250 ), .ZN(_u10_u1_n2276 ) );
NAND2_X1 _u10_u1_U1342  ( .A1(_u10_u1_n3370 ), .A2(_u10_u1_n2276 ), .ZN(_u10_u1_n3348 ) );
AND2_X1 _u10_u1_U1341  ( .A1(_u10_u1_n3369 ), .A2(_u10_gnt_p0_d[0] ), .ZN(_u10_u1_n3330 ) );
NAND2_X1 _u10_u1_U1340  ( .A1(_u10_u1_n3330 ), .A2(_u10_u1_n3149 ), .ZN(_u10_u1_n2351 ) );
INV_X1 _u10_u1_U1339  ( .A(_u10_u1_n1830 ), .ZN(_u10_u1_n2327 ) );
NAND2_X1 _u10_u1_U1338  ( .A1(_u10_u1_n2327 ), .A2(_u10_u1_n2740 ), .ZN(_u10_u1_n3368 ) );
NAND2_X1 _u10_u1_U1337  ( .A1(_u10_u1_n2351 ), .A2(_u10_u1_n3368 ), .ZN(_u10_u1_n2934 ) );
NAND2_X1 _u10_u1_U1336  ( .A1(_u10_u1_n2934 ), .A2(_u10_u1_n2780 ), .ZN(_u10_u1_n3349 ) );
NOR3_X1 _u10_u1_U1335  ( .A1(_u10_u1_n10 ), .A2(_u10_u1_n15 ), .A3(_u10_gnt_p0_d[3] ), .ZN(_u10_u1_n3148 ) );
NAND2_X1 _u10_u1_U1334  ( .A1(_u10_u1_n3324 ), .A2(_u10_u1_n3148 ), .ZN(_u10_u1_n2223 ) );
INV_X1 _u10_u1_U1333  ( .A(_u10_u1_n2223 ), .ZN(_u10_u1_n1950 ) );
NAND2_X1 _u10_u1_U1332  ( .A1(_u10_u1_n3307 ), .A2(_u10_u1_n2618 ), .ZN(_u10_u1_n3367 ) );
AND2_X1 _u10_u1_U1331  ( .A1(_u10_u1_n2239 ), .A2(_u10_u1_n3367 ), .ZN(_u10_u1_n2549 ) );
NAND3_X1 _u10_u1_U1330  ( .A1(_u10_u1_n2815 ), .A2(_u10_u1_n1963 ), .A3(_u10_u1_n1916 ), .ZN(_u10_u1_n2795 ) );
NAND2_X1 _u10_u1_U1329  ( .A1(_u10_u1_n2804 ), .A2(_u10_u1_n1897 ), .ZN(_u10_u1_n3366 ) );
NAND2_X1 _u10_u1_U1328  ( .A1(_u10_u1_n2795 ), .A2(_u10_u1_n3366 ), .ZN(_u10_u1_n3219 ) );
INV_X1 _u10_u1_U1327  ( .A(_u10_u1_n3219 ), .ZN(_u10_u1_n1956 ) );
NAND2_X1 _u10_u1_U1326  ( .A1(_u10_u1_n2152 ), .A2(_u10_u1_n2106 ), .ZN(_u10_u1_n1946 ) );
NOR2_X1 _u10_u1_U1325  ( .A1(_u10_u1_n2356 ), .A2(_u10_u1_n1946 ), .ZN(_u10_u1_n1961 ) );
INV_X1 _u10_u1_U1324  ( .A(_u10_u1_n1946 ), .ZN(_u10_u1_n2108 ) );
NAND2_X1 _u10_u1_U1323  ( .A1(_u10_u1_n2108 ), .A2(_u10_u1_n2133 ), .ZN(_u10_u1_n2794 ) );
INV_X1 _u10_u1_U1322  ( .A(_u10_u1_n2794 ), .ZN(_u10_u1_n2406 ) );
NOR2_X1 _u10_u1_U1321  ( .A1(_u10_u1_n1946 ), .A2(_u10_u1_n3243 ), .ZN(_u10_u1_n3363 ) );
NOR2_X1 _u10_u1_U1320  ( .A1(_u10_u1_n3365 ), .A2(_u10_u1_n3358 ), .ZN(_u10_u1_n3364 ) );
OR2_X1 _u10_u1_U1319  ( .A1(_u10_u1_n3363 ), .A2(_u10_u1_n3364 ), .ZN(_u10_u1_n3362 ) );
NOR4_X1 _u10_u1_U1318  ( .A1(_u10_u1_n1961 ), .A2(_u10_u1_n3361 ), .A3(_u10_u1_n2406 ), .A4(_u10_u1_n3362 ), .ZN(_u10_u1_n3069 ) );
NAND2_X1 _u10_u1_U1317  ( .A1(1'b0), .A2(_u10_u1_n2108 ), .ZN(_u10_u1_n2550 ) );
INV_X1 _u10_u1_U1316  ( .A(_u10_u1_n2550 ), .ZN(_u10_u1_n3309 ) );
NAND2_X1 _u10_u1_U1315  ( .A1(_u10_u1_n2106 ), .A2(_u10_u1_n1955 ), .ZN(_u10_u1_n2766 ) );
NOR4_X1 _u10_u1_U1314  ( .A1(_u10_u1_n2553 ), .A2(_u10_u1_n3309 ), .A3(_u10_u1_n2778 ), .A4(_u10_u1_n2766 ), .ZN(_u10_u1_n3360 ) );
NAND4_X1 _u10_u1_U1313  ( .A1(_u10_u1_n2549 ), .A2(_u10_u1_n1956 ), .A3(_u10_u1_n3069 ), .A4(_u10_u1_n3360 ), .ZN(_u10_u1_n3359 ) );
NAND2_X1 _u10_u1_U1312  ( .A1(_u10_u1_n1950 ), .A2(_u10_u1_n3359 ), .ZN(_u10_u1_n3350 ) );
NAND2_X1 _u10_u1_U1311  ( .A1(_u10_u1_n2351 ), .A2(_u10_u1_n2966 ), .ZN(_u10_u1_n2271 ) );
NAND3_X1 _u10_u1_U1310  ( .A1(_u10_u1_n2725 ), .A2(_u10_u1_n1912 ), .A3(_u10_u1_n3358 ), .ZN(_u10_u1_n3357 ) );
AND2_X1 _u10_u1_U1309  ( .A1(_u10_u1_n1894 ), .A2(_u10_u1_n3357 ), .ZN(_u10_u1_n3057 ) );
AND2_X1 _u10_u1_U1308  ( .A1(_u10_u1_n2271 ), .A2(_u10_u1_n3057 ), .ZN(_u10_u1_n3352 ) );
INV_X1 _u10_u1_U1307  ( .A(_u10_u1_n2480 ), .ZN(_u10_u1_n2321 ) );
NAND2_X1 _u10_u1_U1306  ( .A1(_u10_u1_n3091 ), .A2(_u10_u1_n2321 ), .ZN(_u10_u1_n3099 ) );
NAND2_X1 _u10_u1_U1305  ( .A1(_u10_u1_n3356 ), .A2(_u10_u1_n2012 ), .ZN(_u10_u1_n2169 ) );
INV_X1 _u10_u1_U1304  ( .A(_u10_u1_n2169 ), .ZN(_u10_u1_n2229 ) );
AND2_X1 _u10_u1_U1303  ( .A1(_u10_u1_n3099 ), .A2(_u10_u1_n2229 ), .ZN(_u10_u1_n3353 ) );
INV_X1 _u10_u1_U1302  ( .A(_u10_u1_n2979 ), .ZN(_u10_u1_n2508 ) );
INV_X1 _u10_u1_U1301  ( .A(_u10_u1_n3248 ), .ZN(_u10_u1_n2322 ) );
NAND2_X1 _u10_u1_U1300  ( .A1(_u10_u1_n2508 ), .A2(_u10_u1_n2322 ), .ZN(_u10_u1_n2275 ) );
NAND2_X1 _u10_u1_U1299  ( .A1(_u10_u1_n3355 ), .A2(_u10_u1_n3324 ), .ZN(_u10_u1_n2834 ) );
INV_X1 _u10_u1_U1298  ( .A(_u10_u1_n2834 ), .ZN(_u10_u1_n1920 ) );
NAND2_X1 _u10_u1_U1297  ( .A1(_u10_u1_n2227 ), .A2(_u10_u1_n1920 ), .ZN(_u10_u1_n2674 ) );
NAND2_X1 _u10_u1_U1296  ( .A1(_u10_u1_n2275 ), .A2(_u10_u1_n2674 ), .ZN(_u10_u1_n2088 ) );
AND2_X1 _u10_u1_U1295  ( .A1(_u10_u1_n2088 ), .A2(_u10_u1_n3125 ), .ZN(_u10_u1_n3354 ) );
NOR3_X1 _u10_u1_U1294  ( .A1(_u10_u1_n3352 ), .A2(_u10_u1_n3353 ), .A3(_u10_u1_n3354 ), .ZN(_u10_u1_n3351 ) );
NAND4_X1 _u10_u1_U1293  ( .A1(_u10_u1_n3348 ), .A2(_u10_u1_n3349 ), .A3(_u10_u1_n3350 ), .A4(_u10_u1_n3351 ), .ZN(_u10_u1_n3159 ) );
NOR3_X1 _u10_u1_U1292  ( .A1(_u10_gnt_p0_d[3] ), .A2(_u10_u1_n10 ), .A3(_u10_gnt_p0_d[0] ), .ZN(_u10_u1_n3256 ) );
NAND2_X1 _u10_u1_U1291  ( .A1(_u10_u1_n3298 ), .A2(_u10_u1_n3256 ), .ZN(_u10_u1_n2059 ) );
INV_X1 _u10_u1_U1290  ( .A(_u10_u1_n2059 ), .ZN(_u10_u1_n2234 ) );
NAND2_X1 _u10_u1_U1289  ( .A1(1'b0), .A2(_u10_u1_n2234 ), .ZN(_u10_u1_n3331 ) );
INV_X1 _u10_u1_U1288  ( .A(_u10_u1_n2529 ), .ZN(_u10_u1_n2147 ) );
NAND2_X1 _u10_u1_U1287  ( .A1(_u10_u1_n2152 ), .A2(_u10_u1_n2147 ), .ZN(_u10_u1_n3344 ) );
NAND2_X1 _u10_u1_U1286  ( .A1(_u10_u1_n3330 ), .A2(_u10_gnt_p0_d[1] ), .ZN(_u10_u1_n1994 ) );
INV_X1 _u10_u1_U1285  ( .A(_u10_u1_n1994 ), .ZN(_u10_u1_n2228 ) );
NAND2_X1 _u10_u1_U1284  ( .A1(_u10_u1_n2486 ), .A2(_u10_u1_n2228 ), .ZN(_u10_u1_n2942 ) );
NOR3_X1 _u10_u1_U1283  ( .A1(_u10_u1_n12 ), .A2(_u10_u1_n15 ), .A3(_u10_gnt_p0_d[4] ), .ZN(_u10_u1_n3299 ) );
NAND2_X1 _u10_u1_U1282  ( .A1(_u10_u1_n3324 ), .A2(_u10_u1_n3299 ), .ZN(_u10_u1_n2044 ) );
NAND2_X1 _u10_u1_U1281  ( .A1(_u10_u1_n3297 ), .A2(_u10_u1_n3324 ), .ZN(_u10_u1_n2813 ) );
INV_X1 _u10_u1_U1280  ( .A(_u10_u1_n2813 ), .ZN(_u10_u1_n2453 ) );
NAND2_X1 _u10_u1_U1279  ( .A1(_u10_u1_n2453 ), .A2(_u10_u1_n2014 ), .ZN(_u10_u1_n1826 ) );
NAND2_X1 _u10_u1_U1278  ( .A1(_u10_u1_n2044 ), .A2(_u10_u1_n1826 ), .ZN(_u10_u1_n2247 ) );
NAND2_X1 _u10_u1_U1277  ( .A1(_u10_u1_n3299 ), .A2(_u10_u1_n3149 ), .ZN(_u10_u1_n2019 ) );
INV_X1 _u10_u1_U1276  ( .A(_u10_u1_n2019 ), .ZN(_u10_u1_n3032 ) );
NAND2_X1 _u10_u1_U1275  ( .A1(_u10_u1_n2140 ), .A2(_u10_u1_n3032 ), .ZN(_u10_u1_n3346 ) );
INV_X1 _u10_u1_U1274  ( .A(_u10_u1_n2932 ), .ZN(_u10_u1_n2450 ) );
NAND2_X1 _u10_u1_U1273  ( .A1(_u10_u1_n3227 ), .A2(_u10_u1_n2450 ), .ZN(_u10_u1_n3347 ) );
NAND2_X1 _u10_u1_U1272  ( .A1(_u10_u1_n3346 ), .A2(_u10_u1_n3347 ), .ZN(_u10_u1_n3103 ) );
NOR2_X1 _u10_u1_U1271  ( .A1(_u10_u1_n2247 ), .A2(_u10_u1_n3103 ), .ZN(_u10_u1_n3211 ) );
INV_X1 _u10_u1_U1270  ( .A(_u10_u1_n3211 ), .ZN(_u10_u1_n1836 ) );
NAND2_X1 _u10_u1_U1269  ( .A1(_u10_u1_n3297 ), .A2(_u10_u1_n3149 ), .ZN(_u10_u1_n2020 ) );
INV_X1 _u10_u1_U1268  ( .A(_u10_u1_n2020 ), .ZN(_u10_u1_n2634 ) );
NAND2_X1 _u10_u1_U1267  ( .A1(_u10_u1_n2634 ), .A2(_u10_u1_n2139 ), .ZN(_u10_u1_n2733 ) );
INV_X1 _u10_u1_U1266  ( .A(_u10_u1_n2733 ), .ZN(_u10_u1_n3345 ) );
NAND2_X1 _u10_u1_U1265  ( .A1(_u10_u1_n3345 ), .A2(_u10_u1_n2140 ), .ZN(_u10_u1_n2627 ) );
INV_X1 _u10_u1_U1264  ( .A(_u10_u1_n2627 ), .ZN(_u10_u1_n2249 ) );
NOR2_X1 _u10_u1_U1263  ( .A1(_u10_u1_n1836 ), .A2(_u10_u1_n2249 ), .ZN(_u10_u1_n2298 ) );
NAND3_X1 _u10_u1_U1262  ( .A1(_u10_u1_n3344 ), .A2(_u10_u1_n2942 ), .A3(_u10_u1_n2298 ), .ZN(_u10_u1_n2049 ) );
NAND2_X1 _u10_u1_U1261  ( .A1(_u10_u1_n2171 ), .A2(_u10_u1_n2049 ), .ZN(_u10_u1_n3332 ) );
NAND2_X1 _u10_u1_U1260  ( .A1(1'b0), .A2(_u10_u1_n2322 ), .ZN(_u10_u1_n3333 ) );
INV_X1 _u10_u1_U1259  ( .A(_u10_u1_n2795 ), .ZN(_u10_u1_n2776 ) );
NAND2_X1 _u10_u1_U1258  ( .A1(_u10_u1_n2776 ), .A2(_u10_u1_n2105 ), .ZN(_u10_u1_n2122 ) );
NOR3_X1 _u10_u1_U1257  ( .A1(_u10_u1_n2198 ), .A2(_u10_u1_n2225 ), .A3(_u10_u1_n2122 ), .ZN(_u10_u1_n2707 ) );
NAND3_X1 _u10_u1_U1256  ( .A1(_u10_u1_n1963 ), .A2(_u10_u1_n2619 ), .A3(_u10_u1_n3343 ), .ZN(_u10_u1_n3182 ) );
INV_X1 _u10_u1_U1255  ( .A(_u10_u1_n3182 ), .ZN(_u10_u1_n2535 ) );
INV_X1 _u10_u1_U1254  ( .A(_u10_u1_n2766 ), .ZN(_u10_u1_n2104 ) );
NAND3_X1 _u10_u1_U1253  ( .A1(_u10_u1_n2535 ), .A2(_u10_u1_n2063 ), .A3(_u10_u1_n2104 ), .ZN(_u10_u1_n2121 ) );
NOR2_X1 _u10_u1_U1252  ( .A1(_u10_u1_n2121 ), .A2(_u10_u1_n2287 ), .ZN(_u10_u1_n3153 ) );
NAND2_X1 _u10_u1_U1251  ( .A1(_u10_u1_n3153 ), .A2(_u10_u1_n2439 ), .ZN(_u10_u1_n2383 ) );
INV_X1 _u10_u1_U1250  ( .A(_u10_u1_n2383 ), .ZN(_u10_u1_n3178 ) );
NOR2_X1 _u10_u1_U1249  ( .A1(_u10_u1_n2189 ), .A2(1'b0), .ZN(_u10_u1_n2918 ));
NOR2_X1 _u10_u1_U1248  ( .A1(1'b0), .A2(_u10_u1_n1949 ), .ZN(_u10_u1_n3342 ));
OR2_X1 _u10_u1_U1247  ( .A1(_u10_u1_n2918 ), .A2(_u10_u1_n3342 ), .ZN(_u10_u1_n3341 ) );
NOR4_X1 _u10_u1_U1246  ( .A1(_u10_u1_n2707 ), .A2(_u10_u1_n3340 ), .A3(_u10_u1_n3178 ), .A4(_u10_u1_n3341 ), .ZN(_u10_u1_n2080 ) );
NAND3_X1 _u10_u1_U1245  ( .A1(_u10_gnt_p0_d[3] ), .A2(_u10_gnt_p0_d[0] ),.A3(_u10_u1_n3257 ), .ZN(_u10_u1_n2705 ) );
NOR2_X1 _u10_u1_U1244  ( .A1(_u10_u1_n2080 ), .A2(_u10_u1_n2705 ), .ZN(_u10_u1_n3335 ) );
INV_X1 _u10_u1_U1243  ( .A(_u10_u1_n2042 ), .ZN(_u10_u1_n1988 ) );
NAND2_X1 _u10_u1_U1242  ( .A1(_u10_u1_n1988 ), .A2(_u10_u1_n2043 ), .ZN(_u10_u1_n3339 ) );
NAND2_X1 _u10_u1_U1241  ( .A1(_u10_u1_n3027 ), .A2(_u10_u1_n3339 ), .ZN(_u10_u1_n2025 ) );
AND2_X1 _u10_u1_U1240  ( .A1(_u10_u1_n1933 ), .A2(_u10_u1_n2025 ), .ZN(_u10_u1_n3336 ) );
NAND2_X1 _u10_u1_U1239  ( .A1(_u10_u1_n3256 ), .A2(_u10_u1_n3149 ), .ZN(_u10_u1_n2465 ) );
NOR2_X1 _u10_u1_U1238  ( .A1(_u10_u1_n2465 ), .A2(_u10_u1_n2189 ), .ZN(_u10_u1_n3337 ) );
NOR2_X1 _u10_u1_U1237  ( .A1(_u10_u1_n2298 ), .A2(_u10_u1_n2321 ), .ZN(_u10_u1_n3338 ) );
NOR4_X1 _u10_u1_U1236  ( .A1(_u10_u1_n3335 ), .A2(_u10_u1_n3336 ), .A3(_u10_u1_n3337 ), .A4(_u10_u1_n3338 ), .ZN(_u10_u1_n3334 ) );
NAND4_X1 _u10_u1_U1235  ( .A1(_u10_u1_n3331 ), .A2(_u10_u1_n3332 ), .A3(_u10_u1_n3333 ), .A4(_u10_u1_n3334 ), .ZN(_u10_u1_n3160 ) );
NAND2_X1 _u10_u1_U1234  ( .A1(_u10_u1_n3330 ), .A2(_u10_gnt_p0_d[2] ), .ZN(_u10_u1_n2576 ) );
NAND2_X1 _u10_u1_U1233  ( .A1(_u10_u1_n2133 ), .A2(_u10_u1_n2354 ), .ZN(_u10_u1_n1914 ) );
NOR2_X1 _u10_u1_U1232  ( .A1(_u10_u1_n2576 ), .A2(_u10_u1_n1914 ), .ZN(_u10_u1_n3318 ) );
INV_X1 _u10_u1_U1231  ( .A(_u10_u1_n3153 ), .ZN(_u10_u1_n2064 ) );
NOR2_X1 _u10_u1_U1230  ( .A1(1'b0), .A2(_u10_u1_n2064 ), .ZN(_u10_u1_n3329 ));
NAND3_X1 _u10_u1_U1229  ( .A1(_u10_u1_n2265 ), .A2(_u10_u1_n2201 ), .A3(_u10_u1_n3309 ), .ZN(_u10_u1_n3283 ) );
NAND2_X1 _u10_u1_U1228  ( .A1(_u10_u1_n2588 ), .A2(_u10_u1_n3283 ), .ZN(_u10_u1_n2742 ) );
NOR2_X1 _u10_u1_U1227  ( .A1(_u10_u1_n3329 ), .A2(_u10_u1_n2742 ), .ZN(_u10_u1_n3328 ) );
NOR2_X1 _u10_u1_U1226  ( .A1(1'b0), .A2(_u10_u1_n3328 ), .ZN(_u10_u1_n3326 ));
NAND2_X1 _u10_u1_U1225  ( .A1(_u10_u1_n2203 ), .A2(_u10_u1_n1875 ), .ZN(_u10_u1_n3327 ) );
NAND2_X1 _u10_u1_U1224  ( .A1(_u10_u1_n1949 ), .A2(_u10_u1_n3327 ), .ZN(_u10_u1_n2589 ) );
NOR2_X1 _u10_u1_U1223  ( .A1(_u10_u1_n3326 ), .A2(_u10_u1_n2589 ), .ZN(_u10_u1_n3325 ) );
NOR2_X1 _u10_u1_U1222  ( .A1(_u10_u1_n3325 ), .A2(_u10_u1_n2465 ), .ZN(_u10_u1_n3319 ) );
NAND2_X1 _u10_u1_U1221  ( .A1(_u10_u1_n3256 ), .A2(_u10_u1_n3324 ), .ZN(_u10_u1_n2096 ) );
NAND2_X1 _u10_u1_U1220  ( .A1(_u10_u1_n3298 ), .A2(_u10_u1_n3148 ), .ZN(_u10_u1_n2110 ) );
INV_X1 _u10_u1_U1219  ( .A(_u10_u1_n2110 ), .ZN(_u10_u1_n2263 ) );
NAND2_X1 _u10_u1_U1218  ( .A1(_u10_u1_n2263 ), .A2(_u10_u1_n2068 ), .ZN(_u10_u1_n3323 ) );
NAND2_X1 _u10_u1_U1217  ( .A1(_u10_u1_n2096 ), .A2(_u10_u1_n3323 ), .ZN(_u10_u1_n2428 ) );
INV_X1 _u10_u1_U1216  ( .A(_u10_u1_n2428 ), .ZN(_u10_u1_n3120 ) );
NOR2_X1 _u10_u1_U1215  ( .A1(_u10_u1_n3120 ), .A2(_u10_u1_n2121 ), .ZN(_u10_u1_n3320 ) );
NAND3_X1 _u10_u1_U1214  ( .A1(_u10_u1_n2535 ), .A2(_u10_u1_n1950 ), .A3(_u10_u1_n2104 ), .ZN(_u10_u1_n3321 ) );
INV_X1 _u10_u1_U1213  ( .A(_u10_u1_n2576 ), .ZN(_u10_u1_n1910 ) );
NAND2_X1 _u10_u1_U1212  ( .A1(_u10_u1_n2354 ), .A2(_u10_u1_n1910 ), .ZN(_u10_u1_n3210 ) );
INV_X1 _u10_u1_U1211  ( .A(_u10_u1_n3210 ), .ZN(_u10_u1_n2254 ) );
NAND3_X1 _u10_u1_U1210  ( .A1(_u10_u1_n2254 ), .A2(_u10_u1_n1907 ), .A3(_u10_u1_n3125 ), .ZN(_u10_u1_n3322 ) );
NAND2_X1 _u10_u1_U1209  ( .A1(_u10_u1_n3321 ), .A2(_u10_u1_n3322 ), .ZN(_u10_u1_n2031 ) );
NOR4_X1 _u10_u1_U1208  ( .A1(_u10_u1_n3318 ), .A2(_u10_u1_n3319 ), .A3(_u10_u1_n3320 ), .A4(_u10_u1_n2031 ), .ZN(_u10_u1_n3284 ) );
NOR2_X1 _u10_u1_U1207  ( .A1(_u10_u1_n2826 ), .A2(_u10_u1_n2229 ), .ZN(_u10_u1_n2527 ) );
INV_X1 _u10_u1_U1206  ( .A(_u10_u1_n3125 ), .ZN(_u10_u1_n2628 ) );
NOR2_X1 _u10_u1_U1205  ( .A1(_u10_u1_n2527 ), .A2(_u10_u1_n2628 ), .ZN(_u10_u1_n3312 ) );
NAND2_X1 _u10_u1_U1204  ( .A1(_u10_u1_n3309 ), .A2(_u10_u1_n2265 ), .ZN(_u10_u1_n3317 ) );
NAND3_X1 _u10_u1_U1203  ( .A1(_u10_u1_n2265 ), .A2(_u10_u1_n2418 ), .A3(_u10_u1_n2108 ), .ZN(_u10_u1_n3109 ) );
INV_X1 _u10_u1_U1202  ( .A(_u10_u1_n3109 ), .ZN(_u10_u1_n2087 ) );
NAND2_X1 _u10_u1_U1201  ( .A1(_u10_u1_n2087 ), .A2(1'b0), .ZN(_u10_u1_n2124 ) );
NAND2_X1 _u10_u1_U1200  ( .A1(_u10_u1_n3317 ), .A2(_u10_u1_n2124 ), .ZN(_u10_u1_n2755 ) );
INV_X1 _u10_u1_U1199  ( .A(_u10_u1_n2755 ), .ZN(_u10_u1_n2690 ) );
NOR2_X1 _u10_u1_U1198  ( .A1(_u10_u1_n2690 ), .A2(_u10_u1_n2110 ), .ZN(_u10_u1_n3313 ) );
AND2_X1 _u10_u1_U1197  ( .A1(_u10_u1_n1885 ), .A2(_u10_u1_n2398 ), .ZN(_u10_u1_n2141 ) );
NAND4_X1 _u10_u1_U1196  ( .A1(_u10_u1_n2141 ), .A2(_u10_u1_n2294 ), .A3(_u10_u1_n3316 ), .A4(_u10_u1_n2354 ), .ZN(_u10_u1_n1847 ) );
NOR2_X1 _u10_u1_U1195  ( .A1(_u10_u1_n2353 ), .A2(_u10_u1_n1847 ), .ZN(_u10_u1_n3314 ) );
NAND2_X1 _u10_u1_U1194  ( .A1(_u10_u1_n2887 ), .A2(_u10_u1_n2014 ), .ZN(_u10_u1_n2592 ) );
NOR2_X1 _u10_u1_U1193  ( .A1(_u10_u1_n2813 ), .A2(_u10_u1_n2592 ), .ZN(_u10_u1_n3315 ) );
NOR4_X1 _u10_u1_U1192  ( .A1(_u10_u1_n3312 ), .A2(_u10_u1_n3313 ), .A3(_u10_u1_n3314 ), .A4(_u10_u1_n3315 ), .ZN(_u10_u1_n3285 ) );
NOR2_X1 _u10_u1_U1191  ( .A1(1'b0), .A2(_u10_u1_n2690 ), .ZN(_u10_u1_n3311 ));
NOR2_X1 _u10_u1_U1190  ( .A1(_u10_u1_n3311 ), .A2(_u10_u1_n3153 ), .ZN(_u10_u1_n3310 ) );
NOR2_X1 _u10_u1_U1189  ( .A1(_u10_u1_n3310 ), .A2(_u10_u1_n2059 ), .ZN(_u10_u1_n3300 ) );
NOR2_X1 _u10_u1_U1188  ( .A1(_u10_u1_n3210 ), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n3301 ) );
NOR2_X1 _u10_u1_U1187  ( .A1(_u10_u1_n3309 ), .A2(_u10_u1_n2269 ), .ZN(_u10_u1_n3308 ) );
NOR2_X1 _u10_u1_U1186  ( .A1(_u10_u1_n3308 ), .A2(_u10_u1_n2694 ), .ZN(_u10_u1_n3305 ) );
INV_X1 _u10_u1_U1185  ( .A(_u10_u1_n2574 ), .ZN(_u10_u1_n2399 ) );
NAND3_X1 _u10_u1_U1184  ( .A1(_u10_u1_n2399 ), .A2(_u10_u1_n2155 ), .A3(_u10_u1_n3307 ), .ZN(_u10_u1_n2544 ) );
INV_X1 _u10_u1_U1183  ( .A(_u10_u1_n2544 ), .ZN(_u10_u1_n3306 ) );
NOR2_X1 _u10_u1_U1182  ( .A1(_u10_u1_n3305 ), .A2(_u10_u1_n3306 ), .ZN(_u10_u1_n3304 ) );
NOR2_X1 _u10_u1_U1181  ( .A1(_u10_u1_n3304 ), .A2(_u10_u1_n2096 ), .ZN(_u10_u1_n3302 ) );
INV_X1 _u10_u1_U1180  ( .A(_u10_u1_n2044 ), .ZN(_u10_u1_n2454 ) );
NOR2_X1 _u10_u1_U1179  ( .A1(_u10_u1_n3103 ), .A2(_u10_u1_n2454 ), .ZN(_u10_u1_n2916 ) );
NOR2_X1 _u10_u1_U1178  ( .A1(_u10_u1_n2916 ), .A2(_u10_u1_n2277 ), .ZN(_u10_u1_n3303 ) );
NOR4_X1 _u10_u1_U1177  ( .A1(_u10_u1_n3300 ), .A2(_u10_u1_n3301 ), .A3(_u10_u1_n3302 ), .A4(_u10_u1_n3303 ), .ZN(_u10_u1_n3286 ) );
NAND2_X1 _u10_u1_U1176  ( .A1(_u10_u1_n2141 ), .A2(_u10_u1_n2815 ), .ZN(_u10_u1_n1938 ) );
NOR2_X1 _u10_u1_U1175  ( .A1(_u10_u1_n1938 ), .A2(_u10_u1_n2007 ), .ZN(_u10_u1_n2415 ) );
INV_X1 _u10_u1_U1174  ( .A(_u10_u1_n2415 ), .ZN(_u10_u1_n2633 ) );
NOR3_X1 _u10_u1_U1173  ( .A1(_u10_u1_n2169 ), .A2(_u10_u1_n2435 ), .A3(_u10_u1_n2633 ), .ZN(_u10_u1_n3288 ) );
NAND2_X1 _u10_u1_U1172  ( .A1(_u10_u1_n3298 ), .A2(_u10_u1_n3299 ), .ZN(_u10_u1_n2814 ) );
NOR2_X1 _u10_u1_U1171  ( .A1(_u10_u1_n2650 ), .A2(_u10_u1_n2814 ), .ZN(_u10_u1_n2047 ) );
NAND2_X1 _u10_u1_U1170  ( .A1(_u10_u1_n3297 ), .A2(_u10_u1_n3257 ), .ZN(_u10_u1_n1877 ) );
INV_X1 _u10_u1_U1169  ( .A(_u10_u1_n1877 ), .ZN(_u10_u1_n2672 ) );
NOR3_X1 _u10_u1_U1168  ( .A1(_u10_u1_n2047 ), .A2(_u10_u1_n2672 ), .A3(_u10_u1_n2247 ), .ZN(_u10_u1_n3277 ) );
NOR3_X1 _u10_u1_U1167  ( .A1(_u10_u1_n2544 ), .A2(_u10_u1_n3277 ), .A3(_u10_u1_n2888 ), .ZN(_u10_u1_n3289 ) );
NOR3_X1 _u10_u1_U1166  ( .A1(_u10_u1_n2017 ), .A2(_u10_u1_n2621 ), .A3(_u10_u1_n2435 ), .ZN(_u10_u1_n3296 ) );
NOR3_X1 _u10_u1_U1165  ( .A1(_u10_u1_n1979 ), .A2(_u10_u1_n2861 ), .A3(_u10_u1_n1980 ), .ZN(_u10_u1_n1828 ) );
NOR2_X1 _u10_u1_U1164  ( .A1(_u10_u1_n3296 ), .A2(_u10_u1_n1828 ), .ZN(_u10_u1_n3293 ) );
INV_X1 _u10_u1_U1163  ( .A(_u10_u1_n2127 ), .ZN(_u10_u1_n2434 ) );
INV_X1 _u10_u1_U1162  ( .A(_u10_u1_n3143 ), .ZN(_u10_u1_n1898 ) );
NAND2_X1 _u10_u1_U1161  ( .A1(_u10_u1_n1898 ), .A2(_u10_u1_n3007 ), .ZN(_u10_u1_n3294 ) );
NAND2_X1 _u10_u1_U1160  ( .A1(_u10_u1_n2024 ), .A2(_u10_u1_n2025 ), .ZN(_u10_u1_n3295 ) );
NAND2_X1 _u10_u1_U1159  ( .A1(_u10_u1_n3294 ), .A2(_u10_u1_n3295 ), .ZN(_u10_u1_n1827 ) );
NOR2_X1 _u10_u1_U1158  ( .A1(_u10_u1_n2434 ), .A2(_u10_u1_n1827 ), .ZN(_u10_u1_n2821 ) );
NOR2_X1 _u10_u1_U1157  ( .A1(_u10_u1_n3293 ), .A2(_u10_u1_n2821 ), .ZN(_u10_u1_n3290 ) );
NAND2_X1 _u10_u1_U1156  ( .A1(_u10_u1_n2877 ), .A2(_u10_u1_n2674 ), .ZN(_u10_u1_n2378 ) );
NOR2_X1 _u10_u1_U1155  ( .A1(_u10_u1_n2826 ), .A2(_u10_u1_n2378 ), .ZN(_u10_u1_n3292 ) );
NOR2_X1 _u10_u1_U1154  ( .A1(_u10_u1_n3292 ), .A2(_u10_u1_n2321 ), .ZN(_u10_u1_n3291 ) );
NOR4_X1 _u10_u1_U1153  ( .A1(_u10_u1_n3288 ), .A2(_u10_u1_n3289 ), .A3(_u10_u1_n3290 ), .A4(_u10_u1_n3291 ), .ZN(_u10_u1_n3287 ) );
NAND4_X1 _u10_u1_U1152  ( .A1(_u10_u1_n3284 ), .A2(_u10_u1_n3285 ), .A3(_u10_u1_n3286 ), .A4(_u10_u1_n3287 ), .ZN(_u10_u1_n2558 ) );
NAND2_X1 _u10_u1_U1151  ( .A1(_u10_u1_n2380 ), .A2(_u10_u1_n2672 ), .ZN(_u10_u1_n2955 ) );
OR3_X1 _u10_u1_U1150  ( .A1(_u10_u1_n1946 ), .A2(_u10_u1_n2694 ), .A3(_u10_u1_n2955 ), .ZN(_u10_u1_n3281 ) );
INV_X1 _u10_u1_U1149  ( .A(_u10_u1_n2705 ), .ZN(_u10_u1_n2078 ) );
NAND2_X1 _u10_u1_U1148  ( .A1(_u10_u1_n2439 ), .A2(_u10_u1_n2065 ), .ZN(_u10_u1_n2709 ) );
INV_X1 _u10_u1_U1147  ( .A(_u10_u1_n2709 ), .ZN(_u10_u1_n2086 ) );
NAND3_X1 _u10_u1_U1146  ( .A1(_u10_u1_n2087 ), .A2(_u10_u1_n2078 ), .A3(_u10_u1_n2086 ), .ZN(_u10_u1_n2258 ) );
OR2_X1 _u10_u1_U1145  ( .A1(_u10_u1_n3283 ), .A2(_u10_u1_n2225 ), .ZN(_u10_u1_n3282 ) );
NAND3_X1 _u10_u1_U1144  ( .A1(_u10_u1_n3281 ), .A2(_u10_u1_n2258 ), .A3(_u10_u1_n3282 ), .ZN(_u10_u1_n2891 ) );
NAND2_X1 _u10_u1_U1143  ( .A1(_u10_u1_n2133 ), .A2(_u10_u1_n2397 ), .ZN(_u10_u1_n1966 ) );
AND2_X1 _u10_u1_U1142  ( .A1(_u10_u1_n1966 ), .A2(_u10_u1_n2293 ), .ZN(_u10_u1_n3280 ) );
NOR2_X1 _u10_u1_U1141  ( .A1(_u10_u1_n3280 ), .A2(_u10_u1_n2351 ), .ZN(_u10_u1_n3268 ) );
NAND3_X1 _u10_u1_U1140  ( .A1(_u10_u1_n2014 ), .A2(_u10_u1_n2418 ), .A3(_u10_u1_n2707 ), .ZN(_u10_u1_n2013 ) );
INV_X1 _u10_u1_U1139  ( .A(_u10_u1_n2013 ), .ZN(_u10_u1_n3228 ) );
INV_X1 _u10_u1_U1138  ( .A(_u10_u1_n2592 ), .ZN(_u10_u1_n2882 ) );
NOR2_X1 _u10_u1_U1137  ( .A1(_u10_u1_n3228 ), .A2(_u10_u1_n2882 ), .ZN(_u10_u1_n3279 ) );
NAND3_X1 _u10_u1_U1136  ( .A1(_u10_u1_n2022 ), .A2(_u10_u1_n1844 ), .A3(_u10_u1_n2012 ), .ZN(_u10_u1_n2593 ) );
NOR2_X1 _u10_u1_U1135  ( .A1(_u10_u1_n3279 ), .A2(_u10_u1_n2593 ), .ZN(_u10_u1_n3269 ) );
NOR2_X1 _u10_u1_U1134  ( .A1(_u10_u1_n2506 ), .A2(_u10_u1_n3278 ), .ZN(_u10_u1_n3274 ) );
NAND2_X1 _u10_u1_U1133  ( .A1(_u10_u1_n2019 ), .A2(_u10_u1_n2733 ), .ZN(_u10_u1_n2714 ) );
INV_X1 _u10_u1_U1132  ( .A(_u10_u1_n2714 ), .ZN(_u10_u1_n2963 ) );
NOR2_X1 _u10_u1_U1131  ( .A1(_u10_u1_n2963 ), .A2(_u10_u1_n2632 ), .ZN(_u10_u1_n3275 ) );
INV_X1 _u10_u1_U1130  ( .A(_u10_u1_n3277 ), .ZN(_u10_u1_n3276 ) );
NOR4_X1 _u10_u1_U1129  ( .A1(_u10_u1_n2229 ), .A2(_u10_u1_n3274 ), .A3(_u10_u1_n3275 ), .A4(_u10_u1_n3276 ), .ZN(_u10_u1_n3273 ) );
NOR2_X1 _u10_u1_U1128  ( .A1(_u10_u1_n3273 ), .A2(_u10_u1_n2888 ), .ZN(_u10_u1_n3272 ) );
INV_X1 _u10_u1_U1127  ( .A(_u10_u1_n2096 ), .ZN(_u10_u1_n2236 ) );
NOR2_X1 _u10_u1_U1126  ( .A1(_u10_u1_n3272 ), .A2(_u10_u1_n2236 ), .ZN(_u10_u1_n3271 ) );
NAND2_X1 _u10_u1_U1125  ( .A1(_u10_u1_n2778 ), .A2(_u10_u1_n2063 ), .ZN(_u10_u1_n2756 ) );
NOR2_X1 _u10_u1_U1124  ( .A1(_u10_u1_n3271 ), .A2(_u10_u1_n2756 ), .ZN(_u10_u1_n3270 ) );
NOR3_X1 _u10_u1_U1123  ( .A1(_u10_u1_n3268 ), .A2(_u10_u1_n3269 ), .A3(_u10_u1_n3270 ), .ZN(_u10_u1_n3249 ) );
NOR2_X1 _u10_u1_U1122  ( .A1(1'b0), .A2(_u10_u1_n2588 ), .ZN(_u10_u1_n3267 ));
INV_X1 _u10_u1_U1121  ( .A(_u10_u1_n2191 ), .ZN(_u10_u1_n2286 ) );
NOR2_X1 _u10_u1_U1120  ( .A1(_u10_u1_n3267 ), .A2(_u10_u1_n2286 ), .ZN(_u10_u1_n3266 ) );
NAND2_X1 _u10_u1_U1119  ( .A1(_u10_u1_n1877 ), .A2(_u10_u1_n2705 ), .ZN(_u10_u1_n3111 ) );
INV_X1 _u10_u1_U1118  ( .A(_u10_u1_n3111 ), .ZN(_u10_u1_n3110 ) );
NOR3_X1 _u10_u1_U1117  ( .A1(_u10_u1_n3266 ), .A2(1'b0), .A3(_u10_u1_n3110 ),.ZN(_u10_u1_n3261 ) );
NOR4_X1 _u10_u1_U1116  ( .A1(1'b0), .A2(_u10_u1_n1830 ), .A3(_u10_u1_n2157 ),.A4(_u10_u1_n2725 ), .ZN(_u10_u1_n3262 ) );
INV_X1 _u10_u1_U1115  ( .A(_u10_u1_n1938 ), .ZN(_u10_u1_n2948 ) );
NAND2_X1 _u10_u1_U1114  ( .A1(_u10_u1_n2948 ), .A2(_u10_u1_n2008 ), .ZN(_u10_u1_n2735 ) );
NOR2_X1 _u10_u1_U1113  ( .A1(_u10_u1_n2861 ), .A2(_u10_u1_n2735 ), .ZN(_u10_u1_n3265 ) );
NOR2_X1 _u10_u1_U1112  ( .A1(_u10_u1_n3265 ), .A2(_u10_u1_n2887 ), .ZN(_u10_u1_n3264 ) );
NOR3_X1 _u10_u1_U1111  ( .A1(_u10_u1_n2979 ), .A2(_u10_u1_n3264 ), .A3(_u10_u1_n3248 ), .ZN(_u10_u1_n3263 ) );
NOR3_X1 _u10_u1_U1110  ( .A1(_u10_u1_n3261 ), .A2(_u10_u1_n3262 ), .A3(_u10_u1_n3263 ), .ZN(_u10_u1_n3250 ) );
OR2_X1 _u10_u1_U1109  ( .A1(_u10_u1_n1929 ), .A2(_u10_u1_n2821 ), .ZN(_u10_u1_n3258 ) );
OR2_X1 _u10_u1_U1108  ( .A1(_u10_u1_n2527 ), .A2(_u10_u1_n3245 ), .ZN(_u10_u1_n3259 ) );
NAND2_X1 _u10_u1_U1107  ( .A1(_u10_u1_n2418 ), .A2(_u10_u1_n2045 ), .ZN(_u10_u1_n2671 ) );
NAND2_X1 _u10_u1_U1106  ( .A1(_u10_u1_n2229 ), .A2(_u10_u1_n2671 ), .ZN(_u10_u1_n3260 ) );
NAND3_X1 _u10_u1_U1105  ( .A1(_u10_u1_n3258 ), .A2(_u10_u1_n3259 ), .A3(_u10_u1_n3260 ), .ZN(_u10_u1_n3252 ) );
NOR2_X1 _u10_u1_U1104  ( .A1(_u10_u1_n2465 ), .A2(_u10_u1_n2191 ), .ZN(_u10_u1_n3253 ) );
NAND2_X1 _u10_u1_U1103  ( .A1(_u10_u1_n3256 ), .A2(_u10_u1_n3257 ), .ZN(_u10_u1_n1940 ) );
NOR2_X1 _u10_u1_U1102  ( .A1(_u10_u1_n1940 ), .A2(_u10_u1_n2769 ), .ZN(_u10_u1_n3254 ) );
NOR2_X1 _u10_u1_U1101  ( .A1(_u10_u1_n2209 ), .A2(_u10_u1_n2044 ), .ZN(_u10_u1_n3255 ) );
NOR4_X1 _u10_u1_U1100  ( .A1(_u10_u1_n3252 ), .A2(_u10_u1_n3253 ), .A3(_u10_u1_n3254 ), .A4(_u10_u1_n3255 ), .ZN(_u10_u1_n3251 ) );
NAND3_X1 _u10_u1_U1099  ( .A1(_u10_u1_n3249 ), .A2(_u10_u1_n3250 ), .A3(_u10_u1_n3251 ), .ZN(_u10_u1_n2841 ) );
NAND2_X1 _u10_u1_U1098  ( .A1(_u10_u1_n2912 ), .A2(_u10_u1_n2508 ), .ZN(_u10_u1_n2976 ) );
OR2_X1 _u10_u1_U1097  ( .A1(_u10_u1_n2976 ), .A2(_u10_u1_n3248 ), .ZN(_u10_u1_n3231 ) );
INV_X1 _u10_u1_U1096  ( .A(_u10_u1_n2072 ), .ZN(_u10_u1_n2692 ) );
NAND2_X1 _u10_u1_U1095  ( .A1(_u10_u1_n2692 ), .A2(_u10_u1_n2065 ), .ZN(_u10_u1_n3246 ) );
NOR2_X1 _u10_u1_U1094  ( .A1(1'b0), .A2(_u10_u1_n2553 ), .ZN(_u10_u1_n3123 ));
OR3_X1 _u10_u1_U1093  ( .A1(_u10_u1_n3123 ), .A2(1'b0), .A3(_u10_u1_n2287 ),.ZN(_u10_u1_n3247 ) );
NAND2_X1 _u10_u1_U1092  ( .A1(_u10_u1_n3246 ), .A2(_u10_u1_n3247 ), .ZN(_u10_u1_n2751 ) );
NAND2_X1 _u10_u1_U1091  ( .A1(_u10_u1_n2234 ), .A2(_u10_u1_n2751 ), .ZN(_u10_u1_n3232 ) );
INV_X1 _u10_u1_U1090  ( .A(_u10_u1_n3245 ), .ZN(_u10_u1_n3129 ) );
NOR3_X1 _u10_u1_U1089  ( .A1(_u10_u1_n3129 ), .A2(_u10_u1_n3125 ), .A3(_u10_u1_n3099 ), .ZN(_u10_u1_n3244 ) );
INV_X1 _u10_u1_U1088  ( .A(_u10_u1_n2047 ), .ZN(_u10_u1_n2173 ) );
NOR2_X1 _u10_u1_U1087  ( .A1(_u10_u1_n3244 ), .A2(_u10_u1_n2173 ), .ZN(_u10_u1_n3240 ) );
NOR2_X1 _u10_u1_U1086  ( .A1(_u10_u1_n2942 ), .A2(_u10_u1_n3243 ), .ZN(_u10_u1_n3241 ) );
NOR2_X1 _u10_u1_U1085  ( .A1(_u10_u1_n2814 ), .A2(1'b0), .ZN(_u10_u1_n2958 ));
AND2_X1 _u10_u1_U1084  ( .A1(_u10_u1_n2958 ), .A2(_u10_u1_n2882 ), .ZN(_u10_u1_n3242 ) );
NOR3_X1 _u10_u1_U1083  ( .A1(_u10_u1_n3240 ), .A2(_u10_u1_n3241 ), .A3(_u10_u1_n3242 ), .ZN(_u10_u1_n3233 ) );
NAND2_X1 _u10_u1_U1082  ( .A1(_u10_u1_n2171 ), .A2(_u10_u1_n2354 ), .ZN(_u10_u1_n2829 ) );
NOR2_X1 _u10_u1_U1081  ( .A1(_u10_u1_n2576 ), .A2(_u10_u1_n2829 ), .ZN(_u10_u1_n3235 ) );
NAND2_X1 _u10_u1_U1080  ( .A1(_u10_u1_n2295 ), .A2(_u10_u1_n2141 ), .ZN(_u10_u1_n3239 ) );
NAND2_X1 _u10_u1_U1079  ( .A1(_u10_u1_n1892 ), .A2(_u10_u1_n3239 ), .ZN(_u10_u1_n2493 ) );
AND2_X1 _u10_u1_U1078  ( .A1(_u10_u1_n2493 ), .A2(_u10_u1_n2146 ), .ZN(_u10_u1_n3236 ) );
NOR2_X1 _u10_u1_U1077  ( .A1(_u10_u1_n2110 ), .A2(_u10_u1_n2072 ), .ZN(_u10_u1_n3237 ) );
NOR2_X1 _u10_u1_U1076  ( .A1(_u10_u1_n2478 ), .A2(_u10_u1_n2321 ), .ZN(_u10_u1_n3238 ) );
NOR4_X1 _u10_u1_U1075  ( .A1(_u10_u1_n3235 ), .A2(_u10_u1_n3236 ), .A3(_u10_u1_n3237 ), .A4(_u10_u1_n3238 ), .ZN(_u10_u1_n3234 ) );
AND4_X1 _u10_u1_U1074  ( .A1(_u10_u1_n3231 ), .A2(_u10_u1_n3232 ), .A3(_u10_u1_n3233 ), .A4(_u10_u1_n3234 ), .ZN(_u10_u1_n2334 ) );
NAND2_X1 _u10_u1_U1073  ( .A1(_u10_u1_n2958 ), .A2(_u10_u1_n3228 ), .ZN(_u10_u1_n3229 ) );
NAND3_X1 _u10_u1_U1072  ( .A1(_u10_u1_n2815 ), .A2(_u10_u1_n2934 ), .A3(_u10_u1_n1916 ), .ZN(_u10_u1_n3230 ) );
AND2_X1 _u10_u1_U1071  ( .A1(_u10_u1_n3229 ), .A2(_u10_u1_n3230 ), .ZN(_u10_u1_n2943 ) );
NAND2_X1 _u10_u1_U1070  ( .A1(_u10_u1_n3228 ), .A2(_u10_u1_n2453 ), .ZN(_u10_u1_n3224 ) );
INV_X1 _u10_u1_U1069  ( .A(_u10_u1_n2735 ), .ZN(_u10_u1_n3226 ) );
NAND4_X1 _u10_u1_U1068  ( .A1(_u10_u1_n3226 ), .A2(_u10_u1_n3227 ), .A3(_u10_u1_n2662 ), .A4(_u10_u1_n2450 ), .ZN(_u10_u1_n3225 ) );
AND2_X1 _u10_u1_U1067  ( .A1(_u10_u1_n3224 ), .A2(_u10_u1_n3225 ), .ZN(_u10_u1_n2839 ) );
NAND2_X1 _u10_u1_U1066  ( .A1(_u10_u1_n2672 ), .A2(1'b0), .ZN(_u10_u1_n3222 ) );
INV_X1 _u10_u1_U1065  ( .A(_u10_u1_n1914 ), .ZN(_u10_u1_n2831 ) );
NAND2_X1 _u10_u1_U1064  ( .A1(_u10_u1_n2831 ), .A2(_u10_u1_n1837 ), .ZN(_u10_u1_n3223 ) );
NAND2_X1 _u10_u1_U1063  ( .A1(_u10_u1_n3222 ), .A2(_u10_u1_n3223 ), .ZN(_u10_u1_n2890 ) );
INV_X1 _u10_u1_U1062  ( .A(_u10_u1_n2890 ), .ZN(_u10_u1_n3221 ) );
NAND2_X1 _u10_u1_U1061  ( .A1(_u10_u1_n2839 ), .A2(_u10_u1_n3221 ), .ZN(_u10_u1_n3213 ) );
NOR2_X1 _u10_u1_U1060  ( .A1(_u10_u1_n3143 ), .A2(_u10_u1_n3007 ), .ZN(_u10_u1_n3214 ) );
NAND2_X1 _u10_u1_U1059  ( .A1(_u10_u1_n2046 ), .A2(_u10_u1_n2227 ), .ZN(_u10_u1_n2257 ) );
NOR2_X1 _u10_u1_U1058  ( .A1(_u10_u1_n2834 ), .A2(_u10_u1_n2257 ), .ZN(_u10_u1_n3215 ) );
NAND3_X1 _u10_u1_U1057  ( .A1(_u10_u1_n3182 ), .A2(_u10_u1_n2106 ), .A3(_u10_u1_n2794 ), .ZN(_u10_u1_n3218 ) );
NOR2_X1 _u10_u1_U1056  ( .A1(_u10_u1_n2407 ), .A2(_u10_u1_n1961 ), .ZN(_u10_u1_n2233 ) );
INV_X1 _u10_u1_U1055  ( .A(_u10_u1_n2233 ), .ZN(_u10_u1_n3220 ) );
NOR3_X1 _u10_u1_U1054  ( .A1(_u10_u1_n3218 ), .A2(_u10_u1_n3219 ), .A3(_u10_u1_n3220 ), .ZN(_u10_u1_n3217 ) );
NOR2_X1 _u10_u1_U1053  ( .A1(_u10_u1_n3217 ), .A2(_u10_u1_n1940 ), .ZN(_u10_u1_n3216 ) );
NOR4_X1 _u10_u1_U1052  ( .A1(_u10_u1_n3213 ), .A2(_u10_u1_n3214 ), .A3(_u10_u1_n3215 ), .A4(_u10_u1_n3216 ), .ZN(_u10_u1_n3163 ) );
OR2_X1 _u10_u1_U1051  ( .A1(_u10_u1_n1877 ), .A2(_u10_u1_n2080 ), .ZN(_u10_u1_n3212 ) );
NAND2_X1 _u10_u1_U1050  ( .A1(_u10_u1_n2631 ), .A2(_u10_u1_n3125 ), .ZN(_u10_u1_n2303 ) );
NAND2_X1 _u10_u1_U1049  ( .A1(_u10_u1_n3212 ), .A2(_u10_u1_n2303 ), .ZN(_u10_u1_n3199 ) );
NOR2_X1 _u10_u1_U1048  ( .A1(_u10_u1_n2345 ), .A2(_u10_u1_n3211 ), .ZN(_u10_u1_n3200 ) );
NOR2_X1 _u10_u1_U1047  ( .A1(1'b0), .A2(_u10_u1_n3210 ), .ZN(_u10_u1_n3209 ));
NOR3_X1 _u10_u1_U1046  ( .A1(_u10_u1_n3209 ), .A2(_u10_u1_n2631 ), .A3(_u10_u1_n2249 ), .ZN(_u10_u1_n3208 ) );
INV_X1 _u10_u1_U1045  ( .A(_u10_u1_n2912 ), .ZN(_u10_u1_n3207 ) );
NOR2_X1 _u10_u1_U1044  ( .A1(_u10_u1_n3208 ), .A2(_u10_u1_n3207 ), .ZN(_u10_u1_n3201 ) );
NAND3_X1 _u10_u1_U1043  ( .A1(_u10_u1_n2141 ), .A2(_u10_u1_n2619 ), .A3(_u10_u1_n2486 ), .ZN(_u10_u1_n2484 ) );
INV_X1 _u10_u1_U1042  ( .A(_u10_u1_n2484 ), .ZN(_u10_u1_n2719 ) );
NAND2_X1 _u10_u1_U1041  ( .A1(_u10_u1_n1891 ), .A2(_u10_u1_n2974 ), .ZN(_u10_u1_n3204 ) );
NOR2_X1 _u10_u1_U1040  ( .A1(1'b0), .A2(_u10_u1_n2257 ), .ZN(_u10_u1_n3205 ));
NOR2_X1 _u10_u1_U1039  ( .A1(_u10_u1_n2478 ), .A2(_u10_u1_n3207 ), .ZN(_u10_u1_n3206 ) );
NOR4_X1 _u10_u1_U1038  ( .A1(_u10_u1_n2719 ), .A2(_u10_u1_n3204 ), .A3(_u10_u1_n3205 ), .A4(_u10_u1_n3206 ), .ZN(_u10_u1_n3203 ) );
NOR2_X1 _u10_u1_U1037  ( .A1(_u10_u1_n3203 ), .A2(_u10_u1_n1994 ), .ZN(_u10_u1_n3202 ) );
NOR4_X1 _u10_u1_U1036  ( .A1(_u10_u1_n3199 ), .A2(_u10_u1_n3200 ), .A3(_u10_u1_n3201 ), .A4(_u10_u1_n3202 ), .ZN(_u10_u1_n3164 ) );
INV_X1 _u10_u1_U1035  ( .A(_u10_u1_n2119 ), .ZN(_u10_u1_n3196 ) );
NAND2_X1 _u10_u1_U1034  ( .A1(_u10_u1_n2398 ), .A2(_u10_u1_n2247 ), .ZN(_u10_u1_n3198 ) );
NAND2_X1 _u10_u1_U1033  ( .A1(_u10_u1_n2955 ), .A2(_u10_u1_n3198 ), .ZN(_u10_u1_n3197 ) );
NAND2_X1 _u10_u1_U1032  ( .A1(_u10_u1_n3196 ), .A2(_u10_u1_n3197 ), .ZN(_u10_u1_n3184 ) );
NAND2_X1 _u10_u1_U1031  ( .A1(_u10_u1_n3195 ), .A2(_u10_u1_n2814 ), .ZN(_u10_u1_n3194 ) );
NAND2_X1 _u10_u1_U1030  ( .A1(_u10_u1_n3127 ), .A2(_u10_u1_n3194 ), .ZN(_u10_u1_n3185 ) );
INV_X1 _u10_u1_U1029  ( .A(_u10_u1_n2275 ), .ZN(_u10_u1_n2248 ) );
NAND2_X1 _u10_u1_U1028  ( .A1(_u10_u1_n2522 ), .A2(_u10_u1_n2327 ), .ZN(_u10_u1_n2181 ) );
INV_X1 _u10_u1_U1027  ( .A(_u10_u1_n2181 ), .ZN(_u10_u1_n2949 ) );
NOR2_X1 _u10_u1_U1026  ( .A1(_u10_u1_n2248 ), .A2(_u10_u1_n2949 ), .ZN(_u10_u1_n2296 ) );
NAND2_X1 _u10_u1_U1025  ( .A1(_u10_u1_n2296 ), .A2(_u10_u1_n2627 ), .ZN(_u10_u1_n3193 ) );
NAND2_X1 _u10_u1_U1024  ( .A1(_u10_u1_n2046 ), .A2(_u10_u1_n3193 ), .ZN(_u10_u1_n3186 ) );
NOR2_X1 _u10_u1_U1023  ( .A1(_u10_u1_n1984 ), .A2(_u10_u1_n2507 ), .ZN(_u10_u1_n3191 ) );
NOR2_X1 _u10_u1_U1022  ( .A1(_u10_u1_n2450 ), .A2(_u10_u1_n2322 ), .ZN(_u10_u1_n3192 ) );
NOR2_X1 _u10_u1_U1021  ( .A1(_u10_u1_n3191 ), .A2(_u10_u1_n3192 ), .ZN(_u10_u1_n3188 ) );
NAND3_X1 _u10_u1_U1020  ( .A1(_u10_u1_n2047 ), .A2(_u10_u1_n2370 ), .A3(_u10_u1_n2415 ), .ZN(_u10_u1_n2382 ) );
INV_X1 _u10_u1_U1019  ( .A(_u10_u1_n2382 ), .ZN(_u10_u1_n3189 ) );
NOR3_X1 _u10_u1_U1018  ( .A1(_u10_u1_n1979 ), .A2(_u10_u1_n2353 ), .A3(_u10_u1_n2007 ), .ZN(_u10_u1_n3190 ) );
NOR3_X1 _u10_u1_U1017  ( .A1(_u10_u1_n3188 ), .A2(_u10_u1_n3189 ), .A3(_u10_u1_n3190 ), .ZN(_u10_u1_n3187 ) );
NAND4_X1 _u10_u1_U1016  ( .A1(_u10_u1_n3184 ), .A2(_u10_u1_n3185 ), .A3(_u10_u1_n3186 ), .A4(_u10_u1_n3187 ), .ZN(_u10_u1_n3166 ) );
NAND3_X1 _u10_u1_U1015  ( .A1(_u10_u1_n2398 ), .A2(_u10_u1_n2105 ), .A3(_u10_u1_n2152 ), .ZN(_u10_u1_n2537 ) );
NAND4_X1 _u10_u1_U1014  ( .A1(_u10_u1_n1956 ), .A2(_u10_u1_n3182 ), .A3(_u10_u1_n3183 ), .A4(_u10_u1_n2537 ), .ZN(_u10_u1_n3181 ) );
NAND2_X1 _u10_u1_U1013  ( .A1(_u10_u1_n2147 ), .A2(_u10_u1_n3181 ), .ZN(_u10_u1_n3172 ) );
INV_X1 _u10_u1_U1012  ( .A(_u10_u1_n2122 ), .ZN(_u10_u1_n2693 ) );
NAND2_X1 _u10_u1_U1011  ( .A1(_u10_u1_n2693 ), .A2(_u10_u1_n2068 ), .ZN(_u10_u1_n3180 ) );
NAND2_X1 _u10_u1_U1010  ( .A1(_u10_u1_n2597 ), .A2(_u10_u1_n3180 ), .ZN(_u10_u1_n3179 ) );
NAND2_X1 _u10_u1_U1009  ( .A1(_u10_u1_n2234 ), .A2(_u10_u1_n3179 ), .ZN(_u10_u1_n3173 ) );
NAND2_X1 _u10_u1_U1008  ( .A1(_u10_u1_n2707 ), .A2(_u10_u1_n2454 ), .ZN(_u10_u1_n3176 ) );
NAND2_X1 _u10_u1_U1007  ( .A1(_u10_u1_n3178 ), .A2(_u10_u1_n2247 ), .ZN(_u10_u1_n3177 ) );
NAND2_X1 _u10_u1_U1006  ( .A1(_u10_u1_n3176 ), .A2(_u10_u1_n3177 ), .ZN(_u10_u1_n3175 ) );
NAND2_X1 _u10_u1_U1005  ( .A1(_u10_u1_n3175 ), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n3174 ) );
NAND3_X1 _u10_u1_U1004  ( .A1(_u10_u1_n3172 ), .A2(_u10_u1_n3173 ), .A3(_u10_u1_n3174 ), .ZN(_u10_u1_n3167 ) );
INV_X1 _u10_u1_U1003  ( .A(_u10_u1_n1826 ), .ZN(_u10_u1_n3102 ) );
INV_X1 _u10_u1_U1002  ( .A(_u10_u1_n2826 ), .ZN(_u10_u1_n2320 ) );
NAND2_X1 _u10_u1_U1001  ( .A1(_u10_u1_n2320 ), .A2(_u10_u1_n2173 ), .ZN(_u10_u1_n2595 ) );
NOR4_X1 _u10_u1_U1000  ( .A1(_u10_u1_n3102 ), .A2(_u10_u1_n2595 ), .A3(_u10_u1_n2088 ), .A4(_u10_u1_n3103 ), .ZN(_u10_u1_n3171 ) );
NOR2_X1 _u10_u1_U999  ( .A1(_u10_u1_n3171 ), .A2(_u10_u1_n2045 ), .ZN(_u10_u1_n3168 ) );
NAND3_X1 _u10_u1_U998  ( .A1(_u10_u1_n2022 ), .A2(_u10_u1_n1844 ), .A3(_u10_u1_n2017 ), .ZN(_u10_u1_n2417 ) );
NOR2_X1 _u10_u1_U997  ( .A1(_u10_u1_n2417 ), .A2(_u10_u1_n2013 ), .ZN(_u10_u1_n2713 ) );
AND2_X1 _u10_u1_U996  ( .A1(_u10_u1_n3127 ), .A2(_u10_u1_n2017 ), .ZN(_u10_u1_n3170 ) );
NOR2_X1 _u10_u1_U995  ( .A1(_u10_u1_n2713 ), .A2(_u10_u1_n3170 ), .ZN(_u10_u1_n2050 ) );
NOR2_X1 _u10_u1_U994  ( .A1(_u10_u1_n2050 ), .A2(_u10_u1_n2733 ), .ZN(_u10_u1_n3169 ) );
NOR4_X1 _u10_u1_U993  ( .A1(_u10_u1_n3166 ), .A2(_u10_u1_n3167 ), .A3(_u10_u1_n3168 ), .A4(_u10_u1_n3169 ), .ZN(_u10_u1_n3165 ) );
AND3_X1 _u10_u1_U992  ( .A1(_u10_u1_n3163 ), .A2(_u10_u1_n3164 ), .A3(_u10_u1_n3165 ), .ZN(_u10_u1_n2034 ) );
NAND3_X1 _u10_u1_U991  ( .A1(_u10_u1_n2334 ), .A2(_u10_u1_n2943 ), .A3(_u10_u1_n2034 ), .ZN(_u10_u1_n3162 ) );
OR4_X1 _u10_u1_U990  ( .A1(_u10_u1_n2558 ), .A2(_u10_u1_n2891 ), .A3(_u10_u1_n2841 ), .A4(_u10_u1_n3162 ), .ZN(_u10_u1_n3161 ) );
NOR4_X1 _u10_u1_U989  ( .A1(_u10_u1_n3158 ), .A2(_u10_u1_n3159 ), .A3(_u10_u1_n3160 ), .A4(_u10_u1_n3161 ), .ZN(_u10_u1_n3042 ) );
NOR3_X1 _u10_u1_U988  ( .A1(_u10_u1_n3157 ), .A2(_u10_u1_n1916 ), .A3(_u10_u1_n3073 ), .ZN(_u10_u1_n3064 ) );
NOR2_X1 _u10_u1_U987  ( .A1(1'b0), .A2(_u10_u1_n2608 ), .ZN(_u10_u1_n3156 ));
NAND4_X1 _u10_u1_U986  ( .A1(_u10_u1_n3064 ), .A2(_u10_u1_n2725 ), .A3(_u10_u1_n3156 ), .A4(_u10_u1_n1912 ), .ZN(_u10_u1_n3098 ) );
NAND3_X1 _u10_u1_U985  ( .A1(_u10_u1_n3098 ), .A2(_u10_u1_n2878 ), .A3(_u10_u1_n1920 ), .ZN(_u10_u1_n3135 ) );
NAND3_X1 _u10_u1_U984  ( .A1(_u10_u1_n2948 ), .A2(_u10_u1_n3065 ), .A3(_u10_u1_n3155 ), .ZN(_u10_u1_n3136 ) );
NAND4_X1 _u10_u1_U983  ( .A1(_u10_u1_n3087 ), .A2(_u10_u1_n2756 ), .A3(_u10_u1_n2119 ), .A4(_u10_u1_n2544 ), .ZN(_u10_u1_n3146 ) );
NAND2_X1 _u10_u1_U982  ( .A1(_u10_u1_n2068 ), .A2(_u10_u1_n3146 ), .ZN(_u10_u1_n3151 ) );
NAND2_X1 _u10_u1_U981  ( .A1(_u10_u1_n3151 ), .A2(_u10_u1_n2596 ), .ZN(_u10_u1_n3154 ) );
NAND2_X1 _u10_u1_U980  ( .A1(_u10_u1_n2110 ), .A2(_u10_u1_n2059 ), .ZN(_u10_u1_n2306 ) );
NAND2_X1 _u10_u1_U979  ( .A1(_u10_u1_n3154 ), .A2(_u10_u1_n2306 ), .ZN(_u10_u1_n3137 ) );
AND2_X1 _u10_u1_U978  ( .A1(_u10_u1_n2497 ), .A2(_u10_u1_n2146 ), .ZN(_u10_u1_n2913 ) );
OR4_X1 _u10_u1_U977  ( .A1(_u10_u1_n3153 ), .A2(_u10_u1_n2202 ), .A3(_u10_u1_n3093 ), .A4(_u10_u1_n2203 ), .ZN(_u10_u1_n3150 ) );
NAND2_X1 _u10_u1_U976  ( .A1(_u10_u1_n2693 ), .A2(_u10_u1_n1886 ), .ZN(_u10_u1_n3152 ) );
INV_X1 _u10_u1_U975  ( .A(_u10_u1_n2124 ), .ZN(_u10_u1_n2061 ) );
NAND2_X1 _u10_u1_U974  ( .A1(_u10_u1_n2061 ), .A2(_u10_u1_n2201 ), .ZN(_u10_u1_n2540 ) );
AND2_X1 _u10_u1_U973  ( .A1(_u10_u1_n3152 ), .A2(_u10_u1_n2540 ), .ZN(_u10_u1_n2986 ) );
NAND3_X1 _u10_u1_U972  ( .A1(_u10_u1_n2201 ), .A2(_u10_u1_n3151 ), .A3(_u10_u1_n2986 ), .ZN(_u10_u1_n3083 ) );
NOR4_X1 _u10_u1_U971  ( .A1(_u10_u1_n3150 ), .A2(_u10_u1_n3083 ), .A3(_u10_u1_n2666 ), .A4(_u10_u1_n2742 ), .ZN(_u10_u1_n3147 ) );
NAND2_X1 _u10_u1_U970  ( .A1(_u10_u1_n3148 ), .A2(_u10_u1_n3149 ), .ZN(_u10_u1_n2420 ) );
NOR2_X1 _u10_u1_U969  ( .A1(_u10_u1_n3147 ), .A2(_u10_u1_n2420 ), .ZN(_u10_u1_n3139 ) );
INV_X1 _u10_u1_U968  ( .A(_u10_u1_n3146 ), .ZN(_u10_u1_n3144 ) );
NOR2_X1 _u10_u1_U967  ( .A1(_u10_u1_n2247 ), .A2(_u10_u1_n3111 ), .ZN(_u10_u1_n3145 ) );
NOR4_X1 _u10_u1_U966  ( .A1(_u10_u1_n3144 ), .A2(_u10_u1_n3145 ), .A3(_u10_u1_n2225 ), .A4(_u10_u1_n2287 ), .ZN(_u10_u1_n3140 ) );
NAND2_X1 _u10_u1_U965  ( .A1(_u10_u1_n2127 ), .A2(_u10_u1_n3143 ), .ZN(_u10_u1_n1931 ) );
NOR2_X1 _u10_u1_U964  ( .A1(_u10_u1_n1931 ), .A2(_u10_u1_n2025 ), .ZN(_u10_u1_n3142 ) );
NOR3_X1 _u10_u1_U963  ( .A1(_u10_u1_n2867 ), .A2(_u10_u1_n3142 ), .A3(_u10_u1_n2861 ), .ZN(_u10_u1_n3141 ) );
NOR4_X1 _u10_u1_U962  ( .A1(_u10_u1_n2913 ), .A2(_u10_u1_n3139 ), .A3(_u10_u1_n3140 ), .A4(_u10_u1_n3141 ), .ZN(_u10_u1_n3138 ) );
NAND4_X1 _u10_u1_U961  ( .A1(_u10_u1_n3135 ), .A2(_u10_u1_n3136 ), .A3(_u10_u1_n3137 ), .A4(_u10_u1_n3138 ), .ZN(_u10_u1_n3044 ) );
NAND2_X1 _u10_u1_U960  ( .A1(_u10_u1_n3134 ), .A2(_u10_u1_n2380 ), .ZN(_u10_u1_n3133 ) );
NAND2_X1 _u10_u1_U959  ( .A1(_u10_u1_n2418 ), .A2(_u10_u1_n3133 ), .ZN(_u10_u1_n3132 ) );
NAND2_X1 _u10_u1_U958  ( .A1(_u10_u1_n2047 ), .A2(_u10_u1_n3132 ), .ZN(_u10_u1_n3113 ) );
OR2_X1 _u10_u1_U957  ( .A1(_u10_u1_n3131 ), .A2(1'b0), .ZN(_u10_u1_n3130 ));
NAND2_X1 _u10_u1_U956  ( .A1(_u10_u1_n3130 ), .A2(_u10_u1_n2714 ), .ZN(_u10_u1_n3114 ) );
NAND2_X1 _u10_u1_U955  ( .A1(_u10_u1_n2295 ), .A2(_u10_u1_n2271 ), .ZN(_u10_u1_n2182 ) );
NAND2_X1 _u10_u1_U954  ( .A1(_u10_u1_n2674 ), .A2(_u10_u1_n2182 ), .ZN(_u10_u1_n3128 ) );
NAND2_X1 _u10_u1_U953  ( .A1(_u10_u1_n3128 ), .A2(_u10_u1_n3129 ), .ZN(_u10_u1_n3115 ) );
NOR2_X1 _u10_u1_U952  ( .A1(_u10_u1_n2713 ), .A2(_u10_u1_n3127 ), .ZN(_u10_u1_n3126 ) );
NOR2_X1 _u10_u1_U951  ( .A1(_u10_u1_n3126 ), .A2(_u10_u1_n2019 ), .ZN(_u10_u1_n3117 ) );
NOR2_X1 _u10_u1_U950  ( .A1(_u10_u1_n3125 ), .A2(_u10_u1_n2133 ), .ZN(_u10_u1_n3124 ) );
NOR2_X1 _u10_u1_U949  ( .A1(_u10_u1_n3124 ), .A2(_u10_u1_n2627 ), .ZN(_u10_u1_n3118 ) );
NOR2_X1 _u10_u1_U948  ( .A1(1'b0), .A2(_u10_u1_n3123 ), .ZN(_u10_u1_n3122 ));
NOR2_X1 _u10_u1_U947  ( .A1(_u10_u1_n3122 ), .A2(_u10_u1_n2693 ), .ZN(_u10_u1_n3121 ) );
NOR2_X1 _u10_u1_U946  ( .A1(_u10_u1_n3120 ), .A2(_u10_u1_n3121 ), .ZN(_u10_u1_n3119 ) );
NOR3_X1 _u10_u1_U945  ( .A1(_u10_u1_n3117 ), .A2(_u10_u1_n3118 ), .A3(_u10_u1_n3119 ), .ZN(_u10_u1_n3116 ) );
NAND4_X1 _u10_u1_U944  ( .A1(_u10_u1_n3113 ), .A2(_u10_u1_n3114 ), .A3(_u10_u1_n3115 ), .A4(_u10_u1_n3116 ), .ZN(_u10_u1_n3045 ) );
NAND2_X1 _u10_u1_U943  ( .A1(1'b0), .A2(_u10_u1_n2705 ), .ZN(_u10_u1_n3112 ));
NAND2_X1 _u10_u1_U942  ( .A1(_u10_u1_n3111 ), .A2(_u10_u1_n3112 ), .ZN(_u10_u1_n2284 ) );
INV_X1 _u10_u1_U941  ( .A(_u10_u1_n2284 ), .ZN(_u10_u1_n2917 ) );
NAND2_X1 _u10_u1_U940  ( .A1(_u10_u1_n2203 ), .A2(_u10_u1_n2917 ), .ZN(_u10_u1_n3105 ) );
NAND3_X1 _u10_u1_U939  ( .A1(_u10_u1_n2044 ), .A2(_u10_u1_n3109 ), .A3(_u10_u1_n3110 ), .ZN(_u10_u1_n3108 ) );
NAND2_X1 _u10_u1_U938  ( .A1(1'b0), .A2(_u10_u1_n3108 ), .ZN(_u10_u1_n3106 ));
NAND2_X1 _u10_u1_U937  ( .A1(_u10_u1_n2087 ), .A2(_u10_u1_n3024 ), .ZN(_u10_u1_n2190 ) );
INV_X1 _u10_u1_U936  ( .A(_u10_u1_n2190 ), .ZN(_u10_u1_n1856 ) );
NAND2_X1 _u10_u1_U935  ( .A1(_u10_u1_n1856 ), .A2(_u10_u1_n2234 ), .ZN(_u10_u1_n3107 ) );
NAND3_X1 _u10_u1_U934  ( .A1(_u10_u1_n3105 ), .A2(_u10_u1_n3106 ), .A3(_u10_u1_n3107 ), .ZN(_u10_u1_n3104 ) );
NAND2_X1 _u10_u1_U933  ( .A1(_u10_u1_n2990 ), .A2(_u10_u1_n3104 ), .ZN(_u10_u1_n3075 ) );
NOR2_X1 _u10_u1_U932  ( .A1(_u10_u1_n2826 ), .A2(_u10_u1_n2249 ), .ZN(_u10_u1_n3061 ) );
INV_X1 _u10_u1_U931  ( .A(_u10_u1_n3103 ), .ZN(_u10_u1_n2594 ) );
INV_X1 _u10_u1_U930  ( .A(_u10_u1_n1940 ), .ZN(_u10_u1_n2230 ) );
NAND2_X1 _u10_u1_U929  ( .A1(_u10_u1_n2108 ), .A2(_u10_u1_n2230 ), .ZN(_u10_u1_n2220 ) );
NAND4_X1 _u10_u1_U928  ( .A1(_u10_u1_n3061 ), .A2(_u10_u1_n2594 ), .A3(_u10_u1_n2296 ), .A4(_u10_u1_n2220 ), .ZN(_u10_u1_n2090 ) );
OR3_X1 _u10_u1_U927  ( .A1(_u10_u1_n2378 ), .A2(_u10_u1_n3102 ), .A3(_u10_u1_n2090 ), .ZN(_u10_u1_n3100 ) );
NAND2_X1 _u10_u1_U926  ( .A1(_u10_u1_n3100 ), .A2(_u10_u1_n3101 ), .ZN(_u10_u1_n3076 ) );
NOR2_X1 _u10_u1_U925  ( .A1(_u10_u1_n2780 ), .A2(1'b0), .ZN(_u10_u1_n2310 ));
NAND4_X1 _u10_u1_U924  ( .A1(_u10_u1_n2310 ), .A2(_u10_u1_n2141 ), .A3(_u10_u1_n2354 ), .A4(_u10_u1_n1907 ), .ZN(_u10_u1_n2649 ) );
INV_X1 _u10_u1_U923  ( .A(_u10_u1_n2649 ), .ZN(_u10_u1_n2832 ) );
NAND2_X1 _u10_u1_U922  ( .A1(_u10_u1_n2832 ), .A2(_u10_gnt_p0_d[1] ), .ZN(_u10_u1_n3095 ) );
NAND2_X1 _u10_u1_U921  ( .A1(_u10_u1_n2354 ), .A2(_u10_u1_n3099 ), .ZN(_u10_u1_n3096 ) );
INV_X1 _u10_u1_U920  ( .A(_u10_u1_n3098 ), .ZN(_u10_u1_n3097 ) );
NAND3_X1 _u10_u1_U919  ( .A1(_u10_u1_n3095 ), .A2(_u10_u1_n3096 ), .A3(_u10_u1_n3097 ), .ZN(_u10_u1_n3094 ) );
NAND2_X1 _u10_u1_U918  ( .A1(_u10_u1_n1910 ), .A2(_u10_u1_n3094 ), .ZN(_u10_u1_n3077 ) );
NOR2_X1 _u10_u1_U917  ( .A1(_u10_u1_n2216 ), .A2(_u10_u1_n2190 ), .ZN(_u10_u1_n2114 ) );
NOR2_X1 _u10_u1_U916  ( .A1(_u10_u1_n2114 ), .A2(_u10_u1_n3093 ), .ZN(_u10_u1_n3092 ) );
NOR2_X1 _u10_u1_U915  ( .A1(_u10_u1_n3092 ), .A2(_u10_u1_n2110 ), .ZN(_u10_u1_n3079 ) );
NOR2_X1 _u10_u1_U914  ( .A1(_u10_u1_n3091 ), .A2(_u10_u1_n1895 ), .ZN(_u10_u1_n3089 ) );
NAND2_X1 _u10_u1_U913  ( .A1(1'b0), .A2(_u10_u1_n2295 ), .ZN(_u10_u1_n3090 ));
NAND2_X1 _u10_u1_U912  ( .A1(_u10_u1_n2471 ), .A2(_u10_u1_n3090 ), .ZN(_u10_u1_n2396 ) );
NOR2_X1 _u10_u1_U911  ( .A1(_u10_u1_n3089 ), .A2(_u10_u1_n2396 ), .ZN(_u10_u1_n3088 ) );
NOR2_X1 _u10_u1_U910  ( .A1(_u10_u1_n3088 ), .A2(_u10_u1_n2351 ), .ZN(_u10_u1_n3080 ) );
NOR4_X1 _u10_u1_U909  ( .A1(_u10_u1_n2861 ), .A2(_u10_u1_n2960 ), .A3(_u10_u1_n2979 ), .A4(_u10_u1_n3087 ), .ZN(_u10_u1_n3085 ) );
NOR4_X1 _u10_u1_U908  ( .A1(_u10_u1_n2131 ), .A2(_u10_u1_n1938 ), .A3(_u10_u1_n3086 ), .A4(1'b0), .ZN(_u10_u1_n2134 ) );
NOR2_X1 _u10_u1_U907  ( .A1(_u10_u1_n3085 ), .A2(_u10_u1_n2134 ), .ZN(_u10_u1_n3084 ) );
NOR2_X1 _u10_u1_U906  ( .A1(_u10_u1_n3084 ), .A2(_u10_u1_n2127 ), .ZN(_u10_u1_n3081 ) );
NOR2_X1 _u10_u1_U905  ( .A1(_u10_u1_n2465 ), .A2(1'b0), .ZN(_u10_u1_n2696 ));
AND2_X1 _u10_u1_U904  ( .A1(_u10_u1_n3083 ), .A2(_u10_u1_n2696 ), .ZN(_u10_u1_n3082 ) );
NOR4_X1 _u10_u1_U903  ( .A1(_u10_u1_n3079 ), .A2(_u10_u1_n3080 ), .A3(_u10_u1_n3081 ), .A4(_u10_u1_n3082 ), .ZN(_u10_u1_n3078 ) );
NAND4_X1 _u10_u1_U902  ( .A1(_u10_u1_n3075 ), .A2(_u10_u1_n3076 ), .A3(_u10_u1_n3077 ), .A4(_u10_u1_n3078 ), .ZN(_u10_u1_n3046 ) );
NOR2_X1 _u10_u1_U901  ( .A1(_u10_u1_n1946 ), .A2(_u10_u1_n2960 ), .ZN(_u10_u1_n1960 ) );
NAND2_X1 _u10_u1_U900  ( .A1(_u10_u1_n1960 ), .A2(_u10_u1_n2063 ), .ZN(_u10_u1_n3074 ) );
AND2_X1 _u10_u1_U899  ( .A1(_u10_u1_n2403 ), .A2(_u10_u1_n3074 ), .ZN(_u10_u1_n2920 ) );
NAND2_X1 _u10_u1_U898  ( .A1(_u10_u1_n3073 ), .A2(_u10_u1_n2804 ), .ZN(_u10_u1_n3072 ) );
NAND3_X1 _u10_u1_U897  ( .A1(_u10_u1_n2920 ), .A2(_u10_u1_n3072 ), .A3(_u10_u1_n2549 ), .ZN(_u10_u1_n3071 ) );
NAND2_X1 _u10_u1_U896  ( .A1(_u10_u1_n2230 ), .A2(_u10_u1_n3071 ), .ZN(_u10_u1_n3048 ) );
OR2_X1 _u10_u1_U895  ( .A1(_u10_u1_n2275 ), .A2(_u10_u1_n3070 ), .ZN(_u10_u1_n3049 ) );
OR2_X1 _u10_u1_U894  ( .A1(_u10_u1_n3069 ), .A2(1'b0), .ZN(_u10_u1_n3067 ));
NAND2_X1 _u10_u1_U893  ( .A1(1'b0), .A2(_u10_u1_n2105 ), .ZN(_u10_u1_n3068 ));
NAND3_X1 _u10_u1_U892  ( .A1(_u10_u1_n3067 ), .A2(_u10_u1_n2119 ), .A3(_u10_u1_n3068 ), .ZN(_u10_u1_n3066 ) );
NAND2_X1 _u10_u1_U891  ( .A1(_u10_u1_n2236 ), .A2(_u10_u1_n3066 ), .ZN(_u10_u1_n3050 ) );
NAND2_X1 _u10_u1_U890  ( .A1(_u10_u1_n3065 ), .A2(1'b0), .ZN(_u10_u1_n3063 ));
AND4_X1 _u10_u1_U889  ( .A1(_u10_u1_n2829 ), .A2(_u10_u1_n2725 ), .A3(_u10_u1_n3063 ), .A4(_u10_u1_n3064 ), .ZN(_u10_u1_n3062 ) );
NOR2_X1 _u10_u1_U888  ( .A1(_u10_u1_n3062 ), .A2(_u10_u1_n2353 ), .ZN(_u10_u1_n3052 ) );
NOR2_X1 _u10_u1_U887  ( .A1(_u10_u1_n3061 ), .A2(_u10_u1_n2277 ), .ZN(_u10_u1_n3053 ) );
INV_X1 _u10_u1_U886  ( .A(_u10_u1_n2671 ), .ZN(_u10_u1_n2852 ) );
NOR2_X1 _u10_u1_U885  ( .A1(_u10_u1_n2852 ), .A2(_u10_u1_n2478 ), .ZN(_u10_u1_n3058 ) );
NOR2_X1 _u10_u1_U884  ( .A1(_u10_u1_n3060 ), .A2(_u10_u1_n1907 ), .ZN(_u10_u1_n3059 ) );
NOR4_X1 _u10_u1_U883  ( .A1(_u10_u1_n3056 ), .A2(_u10_u1_n3057 ), .A3(_u10_u1_n3058 ), .A4(_u10_u1_n3059 ), .ZN(_u10_u1_n3055 ) );
NOR2_X1 _u10_u1_U882  ( .A1(_u10_u1_n3055 ), .A2(_u10_u1_n1994 ), .ZN(_u10_u1_n3054 ) );
NOR3_X1 _u10_u1_U881  ( .A1(_u10_u1_n3052 ), .A2(_u10_u1_n3053 ), .A3(_u10_u1_n3054 ), .ZN(_u10_u1_n3051 ) );
NAND4_X1 _u10_u1_U880  ( .A1(_u10_u1_n3048 ), .A2(_u10_u1_n3049 ), .A3(_u10_u1_n3050 ), .A4(_u10_u1_n3051 ), .ZN(_u10_u1_n3047 ) );
NOR4_X1 _u10_u1_U879  ( .A1(_u10_u1_n3044 ), .A2(_u10_u1_n3045 ), .A3(_u10_u1_n3046 ), .A4(_u10_u1_n3047 ), .ZN(_u10_u1_n3043 ) );
NAND2_X1 _u10_u1_U878  ( .A1(_u10_u1_n3042 ), .A2(_u10_u1_n3043 ), .ZN(_u10_u1_n2994 ) );
NOR2_X1 _u10_u1_U877  ( .A1(1'b0), .A2(_u10_u1_n1830 ), .ZN(_u10_u1_n3038 ));
NOR2_X1 _u10_u1_U876  ( .A1(1'b0), .A2(_u10_u1_n2223 ), .ZN(_u10_u1_n3039 ));
NOR2_X1 _u10_u1_U875  ( .A1(1'b0), .A2(_u10_u1_n2576 ), .ZN(_u10_u1_n3040 ));
NOR2_X1 _u10_u1_U874  ( .A1(1'b0), .A2(_u10_u1_n2966 ), .ZN(_u10_u1_n3041 ));
NOR4_X1 _u10_u1_U873  ( .A1(_u10_u1_n3038 ), .A2(_u10_u1_n3039 ), .A3(_u10_u1_n3040 ), .A4(_u10_u1_n3041 ), .ZN(_u10_u1_n2995 ) );
NOR2_X1 _u10_u1_U872  ( .A1(1'b0), .A2(_u10_u1_n2096 ), .ZN(_u10_u1_n3034 ));
NOR2_X1 _u10_u1_U871  ( .A1(1'b0), .A2(_u10_u1_n2110 ), .ZN(_u10_u1_n3035 ));
NOR2_X1 _u10_u1_U870  ( .A1(1'b0), .A2(_u10_u1_n2834 ), .ZN(_u10_u1_n3036 ));
NOR2_X1 _u10_u1_U869  ( .A1(1'b0), .A2(_u10_u1_n2529 ), .ZN(_u10_u1_n3037 ));
NOR4_X1 _u10_u1_U868  ( .A1(_u10_u1_n3034 ), .A2(_u10_u1_n3035 ), .A3(_u10_u1_n3036 ), .A4(_u10_u1_n3037 ), .ZN(_u10_u1_n2996 ) );
NAND2_X1 _u10_u1_U867  ( .A1(_u10_u1_n2234 ), .A2(_u10_u1_n1849 ), .ZN(_u10_u1_n3028 ) );
NAND2_X1 _u10_u1_U866  ( .A1(_u10_u1_n2230 ), .A2(_u10_u1_n1955 ), .ZN(_u10_u1_n3029 ) );
NAND2_X1 _u10_u1_U865  ( .A1(_u10_u1_n2703 ), .A2(_u10_u1_n3033 ), .ZN(_u10_u1_n3030 ) );
NAND2_X1 _u10_u1_U864  ( .A1(_u10_u1_n3032 ), .A2(_u10_u1_n2139 ), .ZN(_u10_u1_n3031 ) );
NAND4_X1 _u10_u1_U863  ( .A1(_u10_u1_n3028 ), .A2(_u10_u1_n3029 ), .A3(_u10_u1_n3030 ), .A4(_u10_u1_n3031 ), .ZN(_u10_u1_n3020 ) );
INV_X1 _u10_u1_U862  ( .A(_u10_u1_n2420 ), .ZN(_u10_u1_n1852 ) );
NAND2_X1 _u10_u1_U861  ( .A1(_u10_u1_n1852 ), .A2(_u10_u1_n1875 ), .ZN(_u10_u1_n3025 ) );
INV_X1 _u10_u1_U860  ( .A(_u10_u1_n3027 ), .ZN(_u10_u1_n1987 ) );
NAND2_X1 _u10_u1_U859  ( .A1(_u10_u1_n1987 ), .A2(_u10_u1_n2043 ), .ZN(_u10_u1_n3026 ) );
NAND2_X1 _u10_u1_U858  ( .A1(_u10_u1_n3025 ), .A2(_u10_u1_n3026 ), .ZN(_u10_u1_n3021 ) );
NOR2_X1 _u10_u1_U857  ( .A1(_u10_gnt_p0_d[4] ), .A2(_u10_u1_n3024 ), .ZN(_u10_u1_n3023 ) );
NOR2_X1 _u10_u1_U856  ( .A1(_u10_u1_n3023 ), .A2(_u10_u1_n2705 ), .ZN(_u10_u1_n3022 ) );
NOR4_X1 _u10_u1_U855  ( .A1(_u10_u1_n3020 ), .A2(_u10_u1_n3021 ), .A3(next_ch), .A4(_u10_u1_n3022 ), .ZN(_u10_u1_n2997 ) );
INV_X1 _u10_u1_U854  ( .A(_u10_u1_n2465 ), .ZN(_u10_u1_n1858 ) );
NAND2_X1 _u10_u1_U853  ( .A1(_u10_u1_n1858 ), .A2(_u10_u1_n1857 ), .ZN(_u10_u1_n3016 ) );
NAND2_X1 _u10_u1_U852  ( .A1(_u10_u1_n2634 ), .A2(_u10_u1_n2136 ), .ZN(_u10_u1_n3017 ) );
NAND2_X1 _u10_u1_U851  ( .A1(_u10_u1_n2228 ), .A2(_u10_u1_n1892 ), .ZN(_u10_u1_n3018 ) );
INV_X1 _u10_u1_U850  ( .A(_u10_u1_n2351 ), .ZN(_u10_u1_n1964 ) );
NAND2_X1 _u10_u1_U849  ( .A1(_u10_u1_n1964 ), .A2(_u10_u1_n2740 ), .ZN(_u10_u1_n3019 ) );
NAND4_X1 _u10_u1_U848  ( .A1(_u10_u1_n3016 ), .A2(_u10_u1_n3017 ), .A3(_u10_u1_n3018 ), .A4(_u10_u1_n3019 ), .ZN(_u10_u1_n2999 ) );
NAND2_X1 _u10_u1_U847  ( .A1(_u10_u1_n2012 ), .A2(_u10_u1_n2017 ), .ZN(_u10_u1_n3012 ) );
OR2_X1 _u10_u1_U846  ( .A1(_u10_u1_n2814 ), .A2(1'b0), .ZN(_u10_u1_n3013 ));
NAND2_X1 _u10_u1_U845  ( .A1(_u10_u1_n2702 ), .A2(_u10_u1_n1903 ), .ZN(_u10_u1_n3014 ) );
NAND2_X1 _u10_u1_U844  ( .A1(_u10_u1_n2672 ), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n3015 ) );
NAND4_X1 _u10_u1_U843  ( .A1(_u10_u1_n3012 ), .A2(_u10_u1_n3013 ), .A3(_u10_u1_n3014 ), .A4(_u10_u1_n3015 ), .ZN(_u10_u1_n3000 ) );
NAND2_X1 _u10_u1_U842  ( .A1(_u10_u1_n2322 ), .A2(_u10_u1_n2867 ), .ZN(_u10_u1_n3008 ) );
NAND2_X1 _u10_u1_U841  ( .A1(_u10_u1_n2450 ), .A2(_u10_u1_n2505 ), .ZN(_u10_u1_n3009 ) );
NAND2_X1 _u10_u1_U840  ( .A1(_u10_u1_n1898 ), .A2(_u10_u1_n1846 ), .ZN(_u10_u1_n3010 ) );
NAND2_X1 _u10_u1_U839  ( .A1(_u10_u1_n1988 ), .A2(_u10_u1_n1845 ), .ZN(_u10_u1_n3011 ) );
NAND4_X1 _u10_u1_U838  ( .A1(_u10_u1_n3008 ), .A2(_u10_u1_n3009 ), .A3(_u10_u1_n3010 ), .A4(_u10_u1_n3011 ), .ZN(_u10_u1_n3001 ) );
NAND2_X1 _u10_u1_U837  ( .A1(_u10_u1_n2434 ), .A2(_u10_u1_n3007 ), .ZN(_u10_u1_n3003 ) );
NAND2_X1 _u10_u1_U836  ( .A1(_u10_u1_n1837 ), .A2(_u10_u1_n1907 ), .ZN(_u10_u1_n3004 ) );
NAND2_X1 _u10_u1_U835  ( .A1(_u10_u1_n2453 ), .A2(_u10_u1_n1844 ), .ZN(_u10_u1_n3005 ) );
NAND2_X1 _u10_u1_U834  ( .A1(_u10_u1_n2454 ), .A2(_u10_u1_n2014 ), .ZN(_u10_u1_n3006 ) );
NAND4_X1 _u10_u1_U833  ( .A1(_u10_u1_n3003 ), .A2(_u10_u1_n3004 ), .A3(_u10_u1_n3005 ), .A4(_u10_u1_n3006 ), .ZN(_u10_u1_n3002 ) );
NOR4_X1 _u10_u1_U832  ( .A1(_u10_u1_n2999 ), .A2(_u10_u1_n3000 ), .A3(_u10_u1_n3001 ), .A4(_u10_u1_n3002 ), .ZN(_u10_u1_n2998 ) );
AND4_X1 _u10_u1_U831  ( .A1(_u10_u1_n2995 ), .A2(_u10_u1_n2996 ), .A3(_u10_u1_n2997 ), .A4(_u10_u1_n2998 ), .ZN(_u10_u1_n1809 ) );
MUX2_X1 _u10_u1_U830  ( .A(_u10_u1_n2994 ), .B(_u10_gnt_p0_d[1] ), .S(_u10_u1_n1809 ), .Z(_u10_u1_n1998 ) );
INV_X1 _u10_u1_U829  ( .A(_u10_u1_n1843 ), .ZN(_u10_u1_n2851 ) );
NOR4_X1 _u10_u1_U828  ( .A1(_u10_u1_n2014 ), .A2(_u10_u1_n2851 ), .A3(1'b0),.A4(1'b0), .ZN(_u10_u1_n2474 ) );
NAND2_X1 _u10_u1_U827  ( .A1(_u10_u1_n2474 ), .A2(_u10_u1_n2495 ), .ZN(_u10_u1_n2973 ) );
INV_X1 _u10_u1_U826  ( .A(_u10_u1_n2973 ), .ZN(_u10_u1_n2498 ) );
NAND2_X1 _u10_u1_U825  ( .A1(_u10_u1_n2498 ), .A2(_u10_u1_n2228 ), .ZN(_u10_u1_n2991 ) );
NAND3_X1 _u10_u1_U824  ( .A1(_u10_u1_n1892 ), .A2(_u10_u1_n2495 ), .A3(1'b0),.ZN(_u10_u1_n2494 ) );
NOR3_X1 _u10_u1_U823  ( .A1(1'b0), .A2(1'b0), .A3(_u10_u1_n2494 ), .ZN(_u10_u1_n2521 ) );
NAND2_X1 _u10_u1_U822  ( .A1(_u10_u1_n2521 ), .A2(_u10_u1_n2618 ), .ZN(_u10_u1_n2643 ) );
INV_X1 _u10_u1_U821  ( .A(_u10_u1_n2643 ), .ZN(_u10_u1_n1941 ) );
NAND2_X1 _u10_u1_U820  ( .A1(_u10_u1_n1941 ), .A2(_u10_u1_n2105 ), .ZN(_u10_u1_n2752 ) );
INV_X1 _u10_u1_U819  ( .A(_u10_u1_n2752 ), .ZN(_u10_u1_n2073 ) );
NOR2_X1 _u10_u1_U818  ( .A1(_u10_u1_n2198 ), .A2(1'b0), .ZN(_u10_u1_n2184 ));
NAND2_X1 _u10_u1_U817  ( .A1(_u10_u1_n2073 ), .A2(_u10_u1_n2184 ), .ZN(_u10_u1_n2466 ) );
NAND2_X1 _u10_u1_U816  ( .A1(_u10_u1_n2184 ), .A2(1'b0), .ZN(_u10_u1_n2188 ));
NAND3_X1 _u10_u1_U815  ( .A1(_u10_u1_n2466 ), .A2(_u10_u1_n2188 ), .A3(_u10_u1_n2189 ), .ZN(_u10_u1_n2993 ) );
NAND2_X1 _u10_u1_U814  ( .A1(_u10_u1_n1858 ), .A2(_u10_u1_n2993 ), .ZN(_u10_u1_n2992 ) );
NAND2_X1 _u10_u1_U813  ( .A1(_u10_u1_n2991 ), .A2(_u10_u1_n2992 ), .ZN(_u10_u1_n2980 ) );
NAND3_X1 _u10_u1_U812  ( .A1(_u10_u1_n1886 ), .A2(_u10_u1_n2990 ), .A3(1'b0),.ZN(_u10_u1_n2938 ) );
INV_X1 _u10_u1_U811  ( .A(_u10_u1_n2938 ), .ZN(_u10_u1_n2285 ) );
NAND2_X1 _u10_u1_U810  ( .A1(_u10_u1_n2285 ), .A2(_u10_u1_n2209 ), .ZN(_u10_u1_n1945 ) );
INV_X1 _u10_u1_U809  ( .A(_u10_u1_n1945 ), .ZN(_u10_u1_n2048 ) );
NOR2_X1 _u10_u1_U808  ( .A1(_u10_u1_n2048 ), .A2(_u10_u1_n2912 ), .ZN(_u10_u1_n2056 ) );
NOR2_X1 _u10_u1_U807  ( .A1(_u10_u1_n2056 ), .A2(_u10_u1_n2989 ), .ZN(_u10_u1_n2988 ) );
NAND2_X1 _u10_u1_U806  ( .A1(1'b0), .A2(_u10_u1_n1903 ), .ZN(_u10_u1_n2009 ));
NOR3_X1 _u10_u1_U805  ( .A1(_u10_u1_n2620 ), .A2(_u10_u1_n2663 ), .A3(_u10_u1_n2009 ), .ZN(_u10_u1_n2967 ) );
AND3_X1 _u10_u1_U804  ( .A1(_u10_u1_n2740 ), .A2(_u10_u1_n2619 ), .A3(_u10_u1_n2967 ), .ZN(_u10_u1_n2941 ) );
NOR3_X1 _u10_u1_U803  ( .A1(_u10_u1_n2988 ), .A2(_u10_u1_n2521 ), .A3(_u10_u1_n2941 ), .ZN(_u10_u1_n2987 ) );
NOR2_X1 _u10_u1_U802  ( .A1(_u10_u1_n2987 ), .A2(_u10_u1_n1830 ), .ZN(_u10_u1_n2981 ) );
NAND2_X1 _u10_u1_U801  ( .A1(_u10_u1_n2498 ), .A2(_u10_u1_n2294 ), .ZN(_u10_u1_n2524 ) );
NOR2_X1 _u10_u1_U800  ( .A1(_u10_u1_n2524 ), .A2(_u10_u1_n2268 ), .ZN(_u10_u1_n2534 ) );
NAND2_X1 _u10_u1_U799  ( .A1(_u10_u1_n2534 ), .A2(_u10_u1_n2104 ), .ZN(_u10_u1_n2392 ) );
INV_X1 _u10_u1_U798  ( .A(_u10_u1_n2392 ), .ZN(_u10_u1_n2116 ) );
NAND3_X1 _u10_u1_U797  ( .A1(_u10_u1_n2074 ), .A2(_u10_u1_n2063 ), .A3(_u10_u1_n2116 ), .ZN(_u10_u1_n2607 ) );
INV_X1 _u10_u1_U796  ( .A(_u10_u1_n2607 ), .ZN(_u10_u1_n2748 ) );
NAND2_X1 _u10_u1_U795  ( .A1(_u10_u1_n2748 ), .A2(_u10_u1_n1849 ), .ZN(_u10_u1_n2541 ) );
NAND2_X1 _u10_u1_U794  ( .A1(_u10_u1_n2986 ), .A2(_u10_u1_n2541 ), .ZN(_u10_u1_n2984 ) );
NOR2_X1 _u10_u1_U793  ( .A1(_u10_u1_n2202 ), .A2(_u10_u1_n2984 ), .ZN(_u10_u1_n2985 ) );
NOR2_X1 _u10_u1_U792  ( .A1(_u10_u1_n2985 ), .A2(_u10_u1_n2420 ), .ZN(_u10_u1_n2982 ) );
AND2_X1 _u10_u1_U791  ( .A1(_u10_u1_n2984 ), .A2(_u10_u1_n2696 ), .ZN(_u10_u1_n2983 ) );
NOR4_X1 _u10_u1_U790  ( .A1(_u10_u1_n2980 ), .A2(_u10_u1_n2981 ), .A3(_u10_u1_n2982 ), .A4(_u10_u1_n2983 ), .ZN(_u10_u1_n2925 ) );
OR3_X1 _u10_u1_U789  ( .A1(_u10_u1_n2343 ), .A2(1'b0), .A3(_u10_u1_n2735 ),.ZN(_u10_u1_n2969 ) );
NAND3_X1 _u10_u1_U788  ( .A1(_u10_u1_n1955 ), .A2(_u10_u1_n2155 ), .A3(_u10_u1_n2941 ), .ZN(_u10_u1_n1952 ) );
INV_X1 _u10_u1_U787  ( .A(_u10_u1_n1952 ), .ZN(_u10_u1_n2758 ) );
INV_X1 _u10_u1_U786  ( .A(_u10_u1_n2417 ), .ZN(_u10_u1_n2464 ) );
NAND4_X1 _u10_u1_U785  ( .A1(_u10_u1_n2758 ), .A2(_u10_u1_n2464 ), .A3(_u10_u1_n2398 ), .A4(_u10_u1_n2483 ), .ZN(_u10_u1_n2933 ) );
NOR2_X1 _u10_u1_U784  ( .A1(_u10_u1_n2466 ), .A2(_u10_u1_n1883 ), .ZN(_u10_u1_n2881 ) );
NAND2_X1 _u10_u1_U783  ( .A1(_u10_u1_n2881 ), .A2(_u10_u1_n2508 ), .ZN(_u10_u1_n2977 ) );
NAND2_X1 _u10_u1_U782  ( .A1(1'b0), .A2(_u10_u1_n2464 ), .ZN(_u10_u1_n2636 ));
INV_X1 _u10_u1_U781  ( .A(_u10_u1_n2636 ), .ZN(_u10_u1_n2894 ) );
NAND3_X1 _u10_u1_U780  ( .A1(_u10_u1_n2483 ), .A2(_u10_u1_n2505 ), .A3(_u10_u1_n2894 ), .ZN(_u10_u1_n2503 ) );
INV_X1 _u10_u1_U779  ( .A(_u10_u1_n2503 ), .ZN(_u10_u1_n1983 ) );
NOR2_X1 _u10_u1_U778  ( .A1(_u10_u1_n2979 ), .A2(_u10_u1_n1945 ), .ZN(_u10_u1_n2323 ) );
NOR3_X1 _u10_u1_U777  ( .A1(_u10_u1_n1983 ), .A2(1'b0), .A3(_u10_u1_n2323 ),.ZN(_u10_u1_n2978 ) );
NAND4_X1 _u10_u1_U776  ( .A1(_u10_u1_n2976 ), .A2(_u10_u1_n2933 ), .A3(_u10_u1_n2977 ), .A4(_u10_u1_n2978 ), .ZN(_u10_u1_n2975 ) );
NAND2_X1 _u10_u1_U775  ( .A1(_u10_u1_n2322 ), .A2(_u10_u1_n2975 ), .ZN(_u10_u1_n2970 ) );
NAND2_X1 _u10_u1_U774  ( .A1(_u10_u1_n2973 ), .A2(_u10_u1_n2974 ), .ZN(_u10_u1_n2972 ) );
NAND3_X1 _u10_u1_U773  ( .A1(_u10_u1_n2972 ), .A2(_u10_u1_n1892 ), .A3(_u10_u1_n2146 ), .ZN(_u10_u1_n2971 ) );
NAND3_X1 _u10_u1_U772  ( .A1(_u10_u1_n2969 ), .A2(_u10_u1_n2970 ), .A3(_u10_u1_n2971 ), .ZN(_u10_u1_n2950 ) );
INV_X1 _u10_u1_U771  ( .A(_u10_u1_n2494 ), .ZN(_u10_u1_n2968 ) );
NOR2_X1 _u10_u1_U770  ( .A1(_u10_u1_n2967 ), .A2(_u10_u1_n2968 ), .ZN(_u10_u1_n2964 ) );
NAND2_X1 _u10_u1_U769  ( .A1(1'b0), .A2(_u10_u1_n2966 ), .ZN(_u10_u1_n2965 ));
NAND2_X1 _u10_u1_U768  ( .A1(_u10_u1_n2271 ), .A2(_u10_u1_n2965 ), .ZN(_u10_u1_n2683 ) );
NOR2_X1 _u10_u1_U767  ( .A1(_u10_u1_n2964 ), .A2(_u10_u1_n2683 ), .ZN(_u10_u1_n2951 ) );
NOR2_X1 _u10_u1_U766  ( .A1(_u10_u1_n2963 ), .A2(_u10_u1_n2417 ), .ZN(_u10_u1_n2961 ) );
INV_X1 _u10_u1_U765  ( .A(_u10_u1_n2593 ), .ZN(_u10_u1_n2962 ) );
NOR2_X1 _u10_u1_U764  ( .A1(_u10_u1_n2961 ), .A2(_u10_u1_n2962 ), .ZN(_u10_u1_n2959 ) );
NOR2_X1 _u10_u1_U763  ( .A1(_u10_u1_n2959 ), .A2(_u10_u1_n2960 ), .ZN(_u10_u1_n2954 ) );
NOR2_X1 _u10_u1_U762  ( .A1(_u10_u1_n2453 ), .A2(_u10_u1_n2958 ), .ZN(_u10_u1_n1879 ) );
NAND2_X1 _u10_u1_U761  ( .A1(_u10_u1_n1879 ), .A2(_u10_u1_n2044 ), .ZN(_u10_u1_n2957 ) );
NAND2_X1 _u10_u1_U760  ( .A1(_u10_u1_n2398 ), .A2(_u10_u1_n2957 ), .ZN(_u10_u1_n2956 ) );
NAND2_X1 _u10_u1_U759  ( .A1(_u10_u1_n2955 ), .A2(_u10_u1_n2956 ), .ZN(_u10_u1_n2617 ) );
NOR2_X1 _u10_u1_U758  ( .A1(_u10_u1_n2954 ), .A2(_u10_u1_n2617 ), .ZN(_u10_u1_n2953 ) );
NOR2_X1 _u10_u1_U757  ( .A1(_u10_u1_n2953 ), .A2(_u10_u1_n1952 ), .ZN(_u10_u1_n2952 ) );
NOR3_X1 _u10_u1_U756  ( .A1(_u10_u1_n2950 ), .A2(_u10_u1_n2951 ), .A3(_u10_u1_n2952 ), .ZN(_u10_u1_n2926 ) );
NAND2_X1 _u10_u1_U755  ( .A1(_u10_u1_n2949 ), .A2(_u10_u1_n2133 ), .ZN(_u10_u1_n2946 ) );
NAND4_X1 _u10_u1_U754  ( .A1(_u10_u1_n2948 ), .A2(_u10_u1_n1843 ), .A3(_u10_u1_n2454 ), .A4(_u10_u1_n1844 ), .ZN(_u10_u1_n2947 ) );
AND2_X1 _u10_u1_U753  ( .A1(_u10_u1_n2946 ), .A2(_u10_u1_n2947 ), .ZN(_u10_u1_n2559 ) );
NAND2_X1 _u10_u1_U752  ( .A1(1'b0), .A2(_u10_u1_n2702 ), .ZN(_u10_u1_n2944 ));
OR2_X1 _u10_u1_U751  ( .A1(_u10_u1_n2173 ), .A2(_u10_u1_n2056 ), .ZN(_u10_u1_n2945 ) );
NAND4_X1 _u10_u1_U750  ( .A1(_u10_u1_n2559 ), .A2(_u10_u1_n2943 ), .A3(_u10_u1_n2944 ), .A4(_u10_u1_n2945 ), .ZN(_u10_u1_n2928 ) );
NAND2_X1 _u10_u1_U749  ( .A1(_u10_u1_n2295 ), .A2(_u10_u1_n2146 ), .ZN(_u10_u1_n2297 ) );
NAND2_X1 _u10_u1_U748  ( .A1(_u10_u1_n2942 ), .A2(_u10_u1_n2297 ), .ZN(_u10_u1_n2342 ) );
NAND2_X1 _u10_u1_U747  ( .A1(_u10_u1_n2133 ), .A2(_u10_u1_n2342 ), .ZN(_u10_u1_n2935 ) );
AND2_X1 _u10_u1_U746  ( .A1(_u10_u1_n2941 ), .A2(_u10_u1_n2155 ), .ZN(_u10_u1_n2940 ) );
NOR2_X1 _u10_u1_U745  ( .A1(_u10_u1_n2534 ), .A2(_u10_u1_n2940 ), .ZN(_u10_u1_n2151 ) );
OR2_X1 _u10_u1_U744  ( .A1(_u10_u1_n1940 ), .A2(_u10_u1_n2151 ), .ZN(_u10_u1_n2936 ) );
OR2_X1 _u10_u1_U743  ( .A1(_u10_u1_n2466 ), .A2(1'b0), .ZN(_u10_u1_n2939 ));
NAND2_X1 _u10_u1_U742  ( .A1(_u10_u1_n2938 ), .A2(_u10_u1_n2939 ), .ZN(_u10_u1_n2706 ) );
NOR2_X1 _u10_u1_U741  ( .A1(_u10_u1_n2216 ), .A2(_u10_u1_n2607 ), .ZN(_u10_u1_n2884 ) );
NOR2_X1 _u10_u1_U740  ( .A1(_u10_u1_n2706 ), .A2(_u10_u1_n2884 ), .ZN(_u10_u1_n2081 ) );
OR2_X1 _u10_u1_U739  ( .A1(_u10_u1_n1877 ), .A2(_u10_u1_n2081 ), .ZN(_u10_u1_n2937 ) );
NAND3_X1 _u10_u1_U738  ( .A1(_u10_u1_n2935 ), .A2(_u10_u1_n2936 ), .A3(_u10_u1_n2937 ), .ZN(_u10_u1_n2929 ) );
INV_X1 _u10_u1_U737  ( .A(_u10_u1_n2934 ), .ZN(_u10_u1_n2684 ) );
NOR2_X1 _u10_u1_U736  ( .A1(_u10_u1_n2684 ), .A2(_u10_u1_n2524 ), .ZN(_u10_u1_n2930 ) );
NOR2_X1 _u10_u1_U735  ( .A1(_u10_u1_n2932 ), .A2(_u10_u1_n2933 ), .ZN(_u10_u1_n2931 ) );
NOR4_X1 _u10_u1_U734  ( .A1(_u10_u1_n2928 ), .A2(_u10_u1_n2929 ), .A3(_u10_u1_n2930 ), .A4(_u10_u1_n2931 ), .ZN(_u10_u1_n2927 ) );
NAND3_X1 _u10_u1_U733  ( .A1(_u10_u1_n2925 ), .A2(_u10_u1_n2926 ), .A3(_u10_u1_n2927 ), .ZN(_u10_u1_n2030 ) );
INV_X1 _u10_u1_U732  ( .A(_u10_u1_n2030 ), .ZN(_u10_u1_n2838 ) );
NAND2_X1 _u10_u1_U731  ( .A1(_u10_u1_n2829 ), .A2(_u10_u1_n1847 ), .ZN(_u10_u1_n2924 ) );
NAND2_X1 _u10_u1_U730  ( .A1(_u10_u1_n1837 ), .A2(_u10_u1_n2924 ), .ZN(_u10_u1_n2897 ) );
NAND3_X1 _u10_u1_U729  ( .A1(_u10_u1_n2086 ), .A2(_u10_u1_n2209 ), .A3(1'b0),.ZN(_u10_u1_n2768 ) );
NAND2_X1 _u10_u1_U728  ( .A1(_u10_u1_n2768 ), .A2(_u10_u1_n1945 ), .ZN(_u10_u1_n2923 ) );
NAND2_X1 _u10_u1_U727  ( .A1(_u10_u1_n2108 ), .A2(_u10_u1_n2923 ), .ZN(_u10_u1_n2921 ) );
NAND4_X1 _u10_u1_U726  ( .A1(1'b0), .A2(_u10_u1_n2294 ), .A3(_u10_u1_n1963 ),.A4(_u10_u1_n2106 ), .ZN(_u10_u1_n2552 ) );
INV_X1 _u10_u1_U725  ( .A(_u10_u1_n2552 ), .ZN(_u10_u1_n2764 ) );
NOR3_X1 _u10_u1_U724  ( .A1(_u10_u1_n1941 ), .A2(1'b0), .A3(_u10_u1_n2764 ),.ZN(_u10_u1_n2922 ) );
NAND3_X1 _u10_u1_U723  ( .A1(_u10_u1_n2920 ), .A2(_u10_u1_n2921 ), .A3(_u10_u1_n2922 ), .ZN(_u10_u1_n2919 ) );
NAND2_X1 _u10_u1_U722  ( .A1(_u10_u1_n2230 ), .A2(_u10_u1_n2919 ), .ZN(_u10_u1_n2898 ) );
AND2_X1 _u10_u1_U721  ( .A1(_u10_u1_n2917 ), .A2(_u10_u1_n2918 ), .ZN(_u10_u1_n2914 ) );
INV_X1 _u10_u1_U720  ( .A(_u10_u1_n2881 ), .ZN(_u10_u1_n1825 ) );
NAND2_X1 _u10_u1_U719  ( .A1(_u10_u1_n2764 ), .A2(_u10_u1_n2105 ), .ZN(_u10_u1_n2759 ) );
INV_X1 _u10_u1_U718  ( .A(_u10_u1_n2759 ), .ZN(_u10_u1_n2196 ) );
NAND2_X1 _u10_u1_U717  ( .A1(_u10_u1_n2196 ), .A2(_u10_u1_n2184 ), .ZN(_u10_u1_n2587 ) );
NOR2_X1 _u10_u1_U716  ( .A1(_u10_u1_n2587 ), .A2(_u10_u1_n1883 ), .ZN(_u10_u1_n2580 ) );
INV_X1 _u10_u1_U715  ( .A(_u10_u1_n2580 ), .ZN(_u10_u1_n2174 ) );
NAND2_X1 _u10_u1_U714  ( .A1(_u10_u1_n1825 ), .A2(_u10_u1_n2174 ), .ZN(_u10_u1_n2459 ) );
INV_X1 _u10_u1_U713  ( .A(_u10_u1_n2768 ), .ZN(_u10_u1_n2825 ) );
NOR2_X1 _u10_u1_U712  ( .A1(_u10_u1_n2171 ), .A2(_u10_u1_n2825 ), .ZN(_u10_u1_n2278 ) );
NAND2_X1 _u10_u1_U711  ( .A1(_u10_u1_n2056 ), .A2(_u10_u1_n2278 ), .ZN(_u10_u1_n2180 ) );
NOR3_X1 _u10_u1_U710  ( .A1(_u10_u1_n2459 ), .A2(_u10_u1_n2887 ), .A3(_u10_u1_n2180 ), .ZN(_u10_u1_n2741 ) );
INV_X1 _u10_u1_U709  ( .A(_u10_u1_n2741 ), .ZN(_u10_u1_n2301 ) );
NAND2_X1 _u10_u1_U708  ( .A1(_u10_u1_n2916 ), .A2(_u10_u1_n2627 ), .ZN(_u10_u1_n2373 ) );
AND2_X1 _u10_u1_U707  ( .A1(_u10_u1_n2301 ), .A2(_u10_u1_n2373 ), .ZN(_u10_u1_n2915 ) );
NOR3_X1 _u10_u1_U706  ( .A1(_u10_u1_n2913 ), .A2(_u10_u1_n2914 ), .A3(_u10_u1_n2915 ), .ZN(_u10_u1_n2899 ) );
NOR3_X1 _u10_u1_U705  ( .A1(_u10_u1_n2459 ), .A2(_u10_u1_n2912 ), .A3(_u10_u1_n2825 ), .ZN(_u10_u1_n2911 ) );
NOR2_X1 _u10_u1_U704  ( .A1(_u10_u1_n2911 ), .A2(_u10_u1_n2877 ), .ZN(_u10_u1_n2901 ) );
NOR2_X1 _u10_u1_U703  ( .A1(_u10_u1_n2459 ), .A2(_u10_u1_n2180 ), .ZN(_u10_u1_n2910 ) );
NOR2_X1 _u10_u1_U702  ( .A1(_u10_u1_n2910 ), .A2(1'b0), .ZN(_u10_u1_n2909 ));
NOR2_X1 _u10_u1_U701  ( .A1(_u10_u1_n2882 ), .A2(_u10_u1_n2909 ), .ZN(_u10_u1_n2908 ) );
NOR2_X1 _u10_u1_U700  ( .A1(_u10_u1_n2908 ), .A2(_u10_u1_n2813 ), .ZN(_u10_u1_n2902 ) );
NOR2_X1 _u10_u1_U699  ( .A1(_u10_u1_n2047 ), .A2(_u10_u1_n2229 ), .ZN(_u10_u1_n2907 ) );
NOR2_X1 _u10_u1_U698  ( .A1(_u10_u1_n2907 ), .A2(_u10_u1_n2768 ), .ZN(_u10_u1_n2903 ) );
AND2_X1 _u10_u1_U697  ( .A1(_u10_u1_n2180 ), .A2(_u10_u1_n2227 ), .ZN(_u10_u1_n2906 ) );
NOR2_X1 _u10_u1_U696  ( .A1(_u10_u1_n2906 ), .A2(_u10_u1_n2482 ), .ZN(_u10_u1_n2905 ) );
NOR2_X1 _u10_u1_U695  ( .A1(_u10_u1_n2905 ), .A2(_u10_u1_n1994 ), .ZN(_u10_u1_n2904 ) );
NOR4_X1 _u10_u1_U694  ( .A1(_u10_u1_n2901 ), .A2(_u10_u1_n2902 ), .A3(_u10_u1_n2903 ), .A4(_u10_u1_n2904 ), .ZN(_u10_u1_n2900 ) );
AND4_X1 _u10_u1_U693  ( .A1(_u10_u1_n2897 ), .A2(_u10_u1_n2898 ), .A3(_u10_u1_n2899 ), .A4(_u10_u1_n2900 ), .ZN(_u10_u1_n2333 ) );
NOR2_X1 _u10_u1_U692  ( .A1(_u10_u1_n1825 ), .A2(_u10_u1_n2169 ), .ZN(_u10_u1_n2889 ) );
NAND2_X1 _u10_u1_U691  ( .A1(_u10_u1_n2474 ), .A2(_u10_u1_n1920 ), .ZN(_u10_u1_n2892 ) );
NAND2_X1 _u10_u1_U690  ( .A1(_u10_u1_n2483 ), .A2(_u10_u1_n2450 ), .ZN(_u10_u1_n2896 ) );
NAND2_X1 _u10_u1_U689  ( .A1(_u10_u1_n2019 ), .A2(_u10_u1_n2896 ), .ZN(_u10_u1_n2895 ) );
NAND2_X1 _u10_u1_U688  ( .A1(_u10_u1_n2894 ), .A2(_u10_u1_n2895 ), .ZN(_u10_u1_n2893 ) );
NAND2_X1 _u10_u1_U687  ( .A1(_u10_u1_n2892 ), .A2(_u10_u1_n2893 ), .ZN(_u10_u1_n2039 ) );
NOR4_X1 _u10_u1_U686  ( .A1(_u10_u1_n2889 ), .A2(_u10_u1_n2890 ), .A3(_u10_u1_n2039 ), .A4(_u10_u1_n2891 ), .ZN(_u10_u1_n2842 ) );
NAND2_X1 _u10_u1_U685  ( .A1(_u10_u1_n1843 ), .A2(1'b0), .ZN(_u10_u1_n2489 ));
INV_X1 _u10_u1_U684  ( .A(_u10_u1_n2489 ), .ZN(_u10_u1_n2475 ) );
NAND2_X1 _u10_u1_U683  ( .A1(_u10_u1_n2475 ), .A2(_u10_u1_n2804 ), .ZN(_u10_u1_n2532 ) );
INV_X1 _u10_u1_U682  ( .A(_u10_u1_n2532 ), .ZN(_u10_u1_n2777 ) );
NAND2_X1 _u10_u1_U681  ( .A1(_u10_u1_n2777 ), .A2(_u10_u1_n2399 ), .ZN(_u10_u1_n2458 ) );
NOR2_X1 _u10_u1_U680  ( .A1(_u10_u1_n2888 ), .A2(_u10_u1_n2458 ), .ZN(_u10_u1_n2883 ) );
NAND2_X1 _u10_u1_U679  ( .A1(_u10_u1_n2852 ), .A2(_u10_u1_n2174 ), .ZN(_u10_u1_n2816 ) );
NOR3_X1 _u10_u1_U678  ( .A1(_u10_u1_n2881 ), .A2(_u10_u1_n2887 ), .A3(_u10_u1_n2816 ), .ZN(_u10_u1_n2451 ) );
NOR2_X1 _u10_u1_U677  ( .A1(_u10_u1_n2451 ), .A2(_u10_u1_n2320 ), .ZN(_u10_u1_n2885 ) );
NOR2_X1 _u10_u1_U676  ( .A1(_u10_u1_n2465 ), .A2(_u10_u1_n2587 ), .ZN(_u10_u1_n2886 ) );
NOR4_X1 _u10_u1_U675  ( .A1(_u10_u1_n2883 ), .A2(_u10_u1_n2884 ), .A3(_u10_u1_n2885 ), .A4(_u10_u1_n2886 ), .ZN(_u10_u1_n2843 ) );
NOR4_X1 _u10_u1_U674  ( .A1(_u10_u1_n2881 ), .A2(_u10_u1_n2882 ), .A3(_u10_u1_n2650 ), .A4(_u10_u1_n2816 ), .ZN(_u10_u1_n2880 ) );
NOR2_X1 _u10_u1_U673  ( .A1(_u10_u1_n2880 ), .A2(_u10_u1_n2814 ), .ZN(_u10_u1_n2870 ) );
NAND3_X1 _u10_u1_U672  ( .A1(_u10_u1_n2141 ), .A2(_u10_u1_n2294 ), .A3(_u10_u1_n2227 ), .ZN(_u10_u1_n2879 ) );
AND3_X1 _u10_u1_U671  ( .A1(_u10_u1_n2878 ), .A2(_u10_u1_n1907 ), .A3(_u10_u1_n2879 ), .ZN(_u10_u1_n2330 ) );
NOR2_X1 _u10_u1_U670  ( .A1(_u10_u1_n2330 ), .A2(_u10_u1_n2834 ), .ZN(_u10_u1_n2871 ) );
NOR2_X1 _u10_u1_U669  ( .A1(_u10_u1_n2877 ), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n2872 ) );
NOR2_X1 _u10_u1_U668  ( .A1(_u10_u1_n2196 ), .A2(_u10_u1_n2073 ), .ZN(_u10_u1_n2876 ) );
NOR2_X1 _u10_u1_U667  ( .A1(_u10_u1_n2876 ), .A2(_u10_u1_n2198 ), .ZN(_u10_u1_n2875 ) );
NOR2_X1 _u10_u1_U666  ( .A1(_u10_u1_n2875 ), .A2(_u10_u1_n2742 ), .ZN(_u10_u1_n2874 ) );
NOR2_X1 _u10_u1_U665  ( .A1(_u10_u1_n2874 ), .A2(_u10_u1_n2420 ), .ZN(_u10_u1_n2873 ) );
NOR4_X1 _u10_u1_U664  ( .A1(_u10_u1_n2870 ), .A2(_u10_u1_n2871 ), .A3(_u10_u1_n2872 ), .A4(_u10_u1_n2873 ), .ZN(_u10_u1_n2844 ) );
NAND2_X1 _u10_u1_U663  ( .A1(_u10_u1_n2868 ), .A2(_u10_u1_n2869 ), .ZN(_u10_u1_n2862 ) );
NAND2_X1 _u10_u1_U662  ( .A1(_u10_u1_n1983 ), .A2(_u10_u1_n2867 ), .ZN(_u10_u1_n2864 ) );
INV_X1 _u10_u1_U661  ( .A(_u10_u1_n1980 ), .ZN(_u10_u1_n2701 ) );
NAND4_X1 _u10_u1_U660  ( .A1(_u10_u1_n2701 ), .A2(_u10_u1_n2370 ), .A3(1'b0),.A4(_u10_u1_n2022 ), .ZN(_u10_u1_n2860 ) );
INV_X1 _u10_u1_U659  ( .A(_u10_u1_n2451 ), .ZN(_u10_u1_n2866 ) );
NAND2_X1 _u10_u1_U658  ( .A1(_u10_u1_n1904 ), .A2(_u10_u1_n2866 ), .ZN(_u10_u1_n2865 ) );
NAND3_X1 _u10_u1_U657  ( .A1(_u10_u1_n2864 ), .A2(_u10_u1_n2860 ), .A3(_u10_u1_n2865 ), .ZN(_u10_u1_n2863 ) );
NAND2_X1 _u10_u1_U656  ( .A1(_u10_u1_n2862 ), .A2(_u10_u1_n2863 ), .ZN(_u10_u1_n2854 ) );
NAND3_X1 _u10_u1_U655  ( .A1(_u10_u1_n1837 ), .A2(_u10_u1_n2650 ), .A3(_u10_u1_n1843 ), .ZN(_u10_u1_n2855 ) );
NAND2_X1 _u10_u1_U654  ( .A1(_u10_u1_n1983 ), .A2(_u10_u1_n2662 ), .ZN(_u10_u1_n2027 ) );
OR2_X1 _u10_u1_U653  ( .A1(_u10_u1_n2860 ), .A2(_u10_u1_n2861 ), .ZN(_u10_u1_n2859 ) );
NAND2_X1 _u10_u1_U652  ( .A1(_u10_u1_n2027 ), .A2(_u10_u1_n2859 ), .ZN(_u10_u1_n2857 ) );
INV_X1 _u10_u1_U651  ( .A(_u10_u1_n2821 ), .ZN(_u10_u1_n2858 ) );
NAND2_X1 _u10_u1_U650  ( .A1(_u10_u1_n2857 ), .A2(_u10_u1_n2858 ), .ZN(_u10_u1_n2856 ) );
NAND3_X1 _u10_u1_U649  ( .A1(_u10_u1_n2854 ), .A2(_u10_u1_n2855 ), .A3(_u10_u1_n2856 ), .ZN(_u10_u1_n2846 ) );
AND2_X1 _u10_u1_U648  ( .A1(_u10_u1_n2674 ), .A2(_u10_u1_n2594 ), .ZN(_u10_u1_n2853 ) );
NOR2_X1 _u10_u1_U647  ( .A1(_u10_u1_n2852 ), .A2(_u10_u1_n2853 ), .ZN(_u10_u1_n2847 ) );
NOR2_X1 _u10_u1_U646  ( .A1(_u10_u1_n2851 ), .A2(_u10_u1_n1938 ), .ZN(_u10_u1_n2850 ) );
NOR3_X1 _u10_u1_U645  ( .A1(_u10_u1_n2671 ), .A2(1'b0), .A3(_u10_u1_n2850 ),.ZN(_u10_u1_n2849 ) );
NOR2_X1 _u10_u1_U644  ( .A1(_u10_u1_n2849 ), .A2(_u10_u1_n2813 ), .ZN(_u10_u1_n2848 ) );
NOR3_X1 _u10_u1_U643  ( .A1(_u10_u1_n2846 ), .A2(_u10_u1_n2847 ), .A3(_u10_u1_n2848 ), .ZN(_u10_u1_n2845 ) );
NAND4_X1 _u10_u1_U642  ( .A1(_u10_u1_n2842 ), .A2(_u10_u1_n2843 ), .A3(_u10_u1_n2844 ), .A4(_u10_u1_n2845 ), .ZN(_u10_u1_n2557 ) );
NOR2_X1 _u10_u1_U641  ( .A1(_u10_u1_n2557 ), .A2(_u10_u1_n2841 ), .ZN(_u10_u1_n2840 ) );
NAND4_X1 _u10_u1_U640  ( .A1(_u10_u1_n2838 ), .A2(_u10_u1_n2839 ), .A3(_u10_u1_n2333 ), .A4(_u10_u1_n2840 ), .ZN(_u10_u1_n2817 ) );
NOR2_X1 _u10_u1_U639  ( .A1(_u10_u1_n2663 ), .A2(_u10_u1_n2837 ), .ZN(_u10_u1_n2835 ) );
NOR4_X1 _u10_u1_U638  ( .A1(_u10_u1_n2835 ), .A2(_u10_u1_n2836 ), .A3(_u10_u1_n2475 ), .A4(_u10_u1_n1916 ), .ZN(_u10_u1_n2718 ) );
OR2_X1 _u10_u1_U637  ( .A1(_u10_u1_n2834 ), .A2(_u10_u1_n2718 ), .ZN(_u10_u1_n2822 ) );
NAND4_X1 _u10_u1_U636  ( .A1(_u10_u1_n2056 ), .A2(_u10_u1_n2768 ), .A3(_u10_u1_n2174 ), .A4(_u10_u1_n2418 ), .ZN(_u10_u1_n2833 ) );
NAND2_X1 _u10_u1_U635  ( .A1(_u10_u1_n2354 ), .A2(_u10_u1_n2833 ), .ZN(_u10_u1_n2828 ) );
NOR4_X1 _u10_u1_U634  ( .A1(1'b0), .A2(_u10_u1_n2831 ), .A3(_u10_u1_n2474 ),.A4(_u10_u1_n2832 ), .ZN(_u10_u1_n2830 ) );
NAND4_X1 _u10_u1_U633  ( .A1(_u10_u1_n2828 ), .A2(_u10_u1_n2829 ), .A3(_u10_u1_n2718 ), .A4(_u10_u1_n2830 ), .ZN(_u10_u1_n2827 ) );
NAND2_X1 _u10_u1_U632  ( .A1(_u10_u1_n1910 ), .A2(_u10_u1_n2827 ), .ZN(_u10_u1_n2823 ) );
NAND2_X1 _u10_u1_U631  ( .A1(_u10_u1_n2825 ), .A2(_u10_u1_n2826 ), .ZN(_u10_u1_n2824 ) );
NAND3_X1 _u10_u1_U630  ( .A1(_u10_u1_n2822 ), .A2(_u10_u1_n2823 ), .A3(_u10_u1_n2824 ), .ZN(_u10_u1_n2818 ) );
NOR2_X1 _u10_u1_U629  ( .A1(_u10_u1_n2821 ), .A2(_u10_u1_n2662 ), .ZN(_u10_u1_n2819 ) );
AND2_X1 _u10_u1_U628  ( .A1(_u10_u1_n2047 ), .A2(_u10_u1_n2171 ), .ZN(_u10_u1_n2820 ) );
NOR4_X1 _u10_u1_U627  ( .A1(_u10_u1_n2817 ), .A2(_u10_u1_n2818 ), .A3(_u10_u1_n2819 ), .A4(_u10_u1_n2820 ), .ZN(_u10_u1_n2652 ) );
NAND2_X1 _u10_u1_U626  ( .A1(_u10_u1_n2248 ), .A2(_u10_u1_n2816 ), .ZN(_u10_u1_n2786 ) );
OR2_X1 _u10_u1_U625  ( .A1(_u10_u1_n1945 ), .A2(_u10_u1_n2219 ), .ZN(_u10_u1_n2787 ) );
AND4_X1 _u10_u1_U624  ( .A1(1'b0), .A2(_u10_u1_n2815 ), .A3(_u10_u1_n1885 ),.A4(_u10_u1_n2008 ), .ZN(_u10_u1_n2687 ) );
NAND2_X1 _u10_u1_U623  ( .A1(_u10_u1_n2086 ), .A2(_u10_u1_n2672 ), .ZN(_u10_u1_n2806 ) );
NAND2_X1 _u10_u1_U622  ( .A1(_u10_u1_n2813 ), .A2(_u10_u1_n2814 ), .ZN(_u10_u1_n2812 ) );
NAND2_X1 _u10_u1_U621  ( .A1(_u10_u1_n2380 ), .A2(_u10_u1_n2812 ), .ZN(_u10_u1_n2807 ) );
NAND3_X1 _u10_u1_U620  ( .A1(_u10_u1_n2017 ), .A2(_u10_u1_n2022 ), .A3(_u10_u1_n2714 ), .ZN(_u10_u1_n2734 ) );
NAND2_X1 _u10_u1_U619  ( .A1(_u10_u1_n2734 ), .A2(_u10_u1_n2811 ), .ZN(_u10_u1_n2810 ) );
NAND2_X1 _u10_u1_U618  ( .A1(_u10_u1_n2398 ), .A2(_u10_u1_n2810 ), .ZN(_u10_u1_n2808 ) );
NAND3_X1 _u10_u1_U617  ( .A1(_u10_u1_n2074 ), .A2(_u10_u1_n2454 ), .A3(_u10_u1_n2439 ), .ZN(_u10_u1_n2809 ) );
NAND4_X1 _u10_u1_U616  ( .A1(_u10_u1_n2806 ), .A2(_u10_u1_n2807 ), .A3(_u10_u1_n2808 ), .A4(_u10_u1_n2809 ), .ZN(_u10_u1_n2805 ) );
NAND2_X1 _u10_u1_U615  ( .A1(_u10_u1_n2687 ), .A2(_u10_u1_n2805 ), .ZN(_u10_u1_n2788 ) );
NAND3_X1 _u10_u1_U614  ( .A1(_u10_u1_n2804 ), .A2(_u10_u1_n2008 ), .A3(1'b0),.ZN(_u10_u1_n2803 ) );
AND2_X1 _u10_u1_U613  ( .A1(_u10_u1_n2803 ), .A2(_u10_u1_n2550 ), .ZN(_u10_u1_n2793 ) );
NAND2_X1 _u10_u1_U612  ( .A1(_u10_u1_n2553 ), .A2(_u10_u1_n2063 ), .ZN(_u10_u1_n2802 ) );
AND2_X1 _u10_u1_U611  ( .A1(_u10_u1_n2752 ), .A2(_u10_u1_n2802 ), .ZN(_u10_u1_n2442 ) );
AND2_X1 _u10_u1_U610  ( .A1(_u10_u1_n2442 ), .A2(_u10_u1_n2759 ), .ZN(_u10_u1_n2238 ) );
NAND2_X1 _u10_u1_U609  ( .A1(_u10_u1_n2086 ), .A2(_u10_u1_n2108 ), .ZN(_u10_u1_n2801 ) );
NAND4_X1 _u10_u1_U608  ( .A1(_u10_u1_n2793 ), .A2(_u10_u1_n2238 ), .A3(_u10_u1_n2399 ), .A4(_u10_u1_n2801 ), .ZN(_u10_u1_n2798 ) );
NAND3_X1 _u10_u1_U607  ( .A1(_u10_u1_n1952 ), .A2(_u10_u1_n2392 ), .A3(_u10_u1_n2122 ), .ZN(_u10_u1_n2799 ) );
INV_X1 _u10_u1_U606  ( .A(_u10_u1_n2458 ), .ZN(_u10_u1_n2800 ) );
NOR4_X1 _u10_u1_U605  ( .A1(_u10_u1_n2798 ), .A2(_u10_u1_n2799 ), .A3(_u10_u1_n2406 ), .A4(_u10_u1_n2800 ), .ZN(_u10_u1_n2797 ) );
NOR2_X1 _u10_u1_U604  ( .A1(_u10_u1_n2797 ), .A2(_u10_u1_n2096 ), .ZN(_u10_u1_n2790 ) );
INV_X1 _u10_u1_U603  ( .A(_u10_u1_n2796 ), .ZN(_u10_u1_n2055 ) );
NOR4_X1 _u10_u1_U602  ( .A1(1'b0), .A2(_u10_u1_n2055 ), .A3(_u10_u1_n1844 ),.A4(_u10_u1_n2506 ), .ZN(_u10_u1_n2791 ) );
NAND4_X1 _u10_u1_U601  ( .A1(_u10_u1_n2793 ), .A2(_u10_u1_n2532 ), .A3(_u10_u1_n2794 ), .A4(_u10_u1_n2795 ), .ZN(_u10_u1_n2763 ) );
AND2_X1 _u10_u1_U600  ( .A1(_u10_u1_n2763 ), .A2(_u10_u1_n2230 ), .ZN(_u10_u1_n2792 ) );
NOR3_X1 _u10_u1_U599  ( .A1(_u10_u1_n2790 ), .A2(_u10_u1_n2791 ), .A3(_u10_u1_n2792 ), .ZN(_u10_u1_n2789 ) );
NAND4_X1 _u10_u1_U598  ( .A1(_u10_u1_n2786 ), .A2(_u10_u1_n2787 ), .A3(_u10_u1_n2788 ), .A4(_u10_u1_n2789 ), .ZN(_u10_u1_n2743 ) );
OR2_X1 _u10_u1_U597  ( .A1(_u10_u1_n2278 ), .A2(_u10_u1_n2296 ), .ZN(_u10_u1_n2770 ) );
NAND2_X1 _u10_u1_U596  ( .A1(_u10_u1_n2454 ), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n2785 ) );
NAND2_X1 _u10_u1_U595  ( .A1(_u10_u1_n1877 ), .A2(_u10_u1_n2785 ), .ZN(_u10_u1_n1876 ) );
NAND2_X1 _u10_u1_U594  ( .A1(_u10_u1_n2707 ), .A2(_u10_u1_n1876 ), .ZN(_u10_u1_n2771 ) );
NAND2_X1 _u10_u1_U593  ( .A1(_u10_u1_n2278 ), .A2(_u10_u1_n1945 ), .ZN(_u10_u1_n2784 ) );
NAND2_X1 _u10_u1_U592  ( .A1(_u10_u1_n2152 ), .A2(_u10_u1_n2784 ), .ZN(_u10_u1_n2782 ) );
NAND2_X1 _u10_u1_U591  ( .A1(_u10_u1_n2521 ), .A2(_u10_u1_n2155 ), .ZN(_u10_u1_n2783 ) );
AND3_X1 _u10_u1_U590  ( .A1(_u10_u1_n2782 ), .A2(_u10_u1_n2537 ), .A3(_u10_u1_n2783 ), .ZN(_u10_u1_n2309 ) );
NAND2_X1 _u10_u1_U589  ( .A1(1'b0), .A2(_u10_u1_n2008 ), .ZN(_u10_u1_n2781 ));
NAND2_X1 _u10_u1_U588  ( .A1(_u10_u1_n2495 ), .A2(_u10_u1_n2781 ), .ZN(_u10_u1_n2739 ) );
INV_X1 _u10_u1_U587  ( .A(_u10_u1_n2739 ), .ZN(_u10_u1_n2724 ) );
NOR3_X1 _u10_u1_U586  ( .A1(_u10_u1_n2780 ), .A2(_u10_u1_n2724 ), .A3(_u10_u1_n2268 ), .ZN(_u10_u1_n2779 ) );
NOR4_X1 _u10_u1_U585  ( .A1(_u10_u1_n2776 ), .A2(_u10_u1_n2777 ), .A3(_u10_u1_n2778 ), .A4(_u10_u1_n2779 ), .ZN(_u10_u1_n2775 ) );
NAND4_X1 _u10_u1_U584  ( .A1(_u10_u1_n2309 ), .A2(_u10_u1_n2151 ), .A3(_u10_u1_n2774 ), .A4(_u10_u1_n2775 ), .ZN(_u10_u1_n2773 ) );
NAND2_X1 _u10_u1_U583  ( .A1(_u10_u1_n2147 ), .A2(_u10_u1_n2773 ), .ZN(_u10_u1_n2772 ) );
NAND3_X1 _u10_u1_U582  ( .A1(_u10_u1_n2770 ), .A2(_u10_u1_n2771 ), .A3(_u10_u1_n2772 ), .ZN(_u10_u1_n2744 ) );
NAND3_X1 _u10_u1_U581  ( .A1(_u10_u1_n1952 ), .A2(_u10_u1_n2392 ), .A3(_u10_u1_n2769 ), .ZN(_u10_u1_n2761 ) );
NOR2_X1 _u10_u1_U580  ( .A1(_u10_u1_n1946 ), .A2(_u10_u1_n2768 ), .ZN(_u10_u1_n2767 ) );
OR3_X1 _u10_u1_U579  ( .A1(_u10_u1_n2766 ), .A2(_u10_u1_n1941 ), .A3(_u10_u1_n2767 ), .ZN(_u10_u1_n2765 ) );
NOR4_X1 _u10_u1_U578  ( .A1(_u10_u1_n2764 ), .A2(_u10_u1_n2553 ), .A3(_u10_u1_n1960 ), .A4(_u10_u1_n2765 ), .ZN(_u10_u1_n2267 ) );
INV_X1 _u10_u1_U577  ( .A(_u10_u1_n2267 ), .ZN(_u10_u1_n2762 ) );
NOR3_X1 _u10_u1_U576  ( .A1(_u10_u1_n2761 ), .A2(_u10_u1_n2762 ), .A3(_u10_u1_n2763 ), .ZN(_u10_u1_n2760 ) );
NOR2_X1 _u10_u1_U575  ( .A1(_u10_u1_n2760 ), .A2(_u10_u1_n2223 ), .ZN(_u10_u1_n2745 ) );
NAND3_X1 _u10_u1_U574  ( .A1(_u10_u1_n2122 ), .A2(_u10_u1_n2063 ), .A3(_u10_u1_n2759 ), .ZN(_u10_u1_n2754 ) );
NOR3_X1 _u10_u1_U573  ( .A1(_u10_u1_n2687 ), .A2(1'b0), .A3(_u10_u1_n2758 ),.ZN(_u10_u1_n2757 ) );
NAND3_X1 _u10_u1_U572  ( .A1(_u10_u1_n2756 ), .A2(_u10_u1_n2458 ), .A3(_u10_u1_n2757 ), .ZN(_u10_u1_n2695 ) );
NOR3_X1 _u10_u1_U571  ( .A1(_u10_u1_n2754 ), .A2(_u10_u1_n2695 ), .A3(_u10_u1_n2755 ), .ZN(_u10_u1_n2753 ) );
NOR2_X1 _u10_u1_U570  ( .A1(1'b0), .A2(_u10_u1_n2753 ), .ZN(_u10_u1_n2749 ));
NOR2_X1 _u10_u1_U569  ( .A1(_u10_u1_n2287 ), .A2(_u10_u1_n2752 ), .ZN(_u10_u1_n2750 ) );
NOR4_X1 _u10_u1_U568  ( .A1(_u10_u1_n2748 ), .A2(_u10_u1_n2749 ), .A3(_u10_u1_n2750 ), .A4(_u10_u1_n2751 ), .ZN(_u10_u1_n2747 ) );
NOR2_X1 _u10_u1_U567  ( .A1(_u10_u1_n2747 ), .A2(_u10_u1_n2059 ), .ZN(_u10_u1_n2746 ) );
NOR4_X1 _u10_u1_U566  ( .A1(_u10_u1_n2743 ), .A2(_u10_u1_n2744 ), .A3(_u10_u1_n2745 ), .A4(_u10_u1_n2746 ), .ZN(_u10_u1_n2653 ) );
NAND2_X1 _u10_u1_U565  ( .A1(_u10_u1_n2696 ), .A2(_u10_u1_n2742 ), .ZN(_u10_u1_n2726 ) );
OR2_X1 _u10_u1_U564  ( .A1(_u10_u1_n2250 ), .A2(_u10_u1_n2741 ), .ZN(_u10_u1_n2727 ) );
NAND2_X1 _u10_u1_U563  ( .A1(1'b0), .A2(_u10_u1_n2522 ), .ZN(_u10_u1_n2525 ));
NAND3_X1 _u10_u1_U562  ( .A1(_u10_u1_n2739 ), .A2(_u10_u1_n2740 ), .A3(_u10_u1_n2294 ), .ZN(_u10_u1_n2738 ) );
NAND3_X1 _u10_u1_U561  ( .A1(_u10_u1_n2737 ), .A2(_u10_u1_n2525 ), .A3(_u10_u1_n2738 ), .ZN(_u10_u1_n2736 ) );
NAND2_X1 _u10_u1_U560  ( .A1(_u10_u1_n2327 ), .A2(_u10_u1_n2736 ), .ZN(_u10_u1_n2728 ) );
NOR2_X1 _u10_u1_U559  ( .A1(_u10_u1_n2735 ), .A2(_u10_u1_n2346 ), .ZN(_u10_u1_n2730 ) );
NOR2_X1 _u10_u1_U558  ( .A1(_u10_u1_n1844 ), .A2(_u10_u1_n2734 ), .ZN(_u10_u1_n2731 ) );
NOR2_X1 _u10_u1_U557  ( .A1(_u10_u1_n2636 ), .A2(_u10_u1_n2733 ), .ZN(_u10_u1_n2732 ) );
NOR3_X1 _u10_u1_U556  ( .A1(_u10_u1_n2730 ), .A2(_u10_u1_n2731 ), .A3(_u10_u1_n2732 ), .ZN(_u10_u1_n2729 ) );
NAND4_X1 _u10_u1_U555  ( .A1(_u10_u1_n2726 ), .A2(_u10_u1_n2727 ), .A3(_u10_u1_n2728 ), .A4(_u10_u1_n2729 ), .ZN(_u10_u1_n2697 ) );
NAND2_X1 _u10_u1_U554  ( .A1(_u10_u1_n2475 ), .A2(_u10_u1_n2146 ), .ZN(_u10_u1_n2721 ) );
INV_X1 _u10_u1_U553  ( .A(_u10_u1_n2683 ), .ZN(_u10_u1_n1887 ) );
NAND2_X1 _u10_u1_U552  ( .A1(_u10_u1_n2724 ), .A2(_u10_u1_n2725 ), .ZN(_u10_u1_n2723 ) );
NAND2_X1 _u10_u1_U551  ( .A1(_u10_u1_n1887 ), .A2(_u10_u1_n2723 ), .ZN(_u10_u1_n2722 ) );
NAND2_X1 _u10_u1_U550  ( .A1(_u10_u1_n2721 ), .A2(_u10_u1_n2722 ), .ZN(_u10_u1_n2720 ) );
NAND2_X1 _u10_u1_U549  ( .A1(_u10_u1_n2720 ), .A2(_u10_u1_n1892 ), .ZN(_u10_u1_n2710 ) );
NAND2_X1 _u10_u1_U548  ( .A1(1'b0), .A2(_u10_u1_n2227 ), .ZN(_u10_u1_n2716 ));
NAND2_X1 _u10_u1_U547  ( .A1(_u10_u1_n2719 ), .A2(_u10_gnt_p0_d[2] ), .ZN(_u10_u1_n2717 ) );
NAND3_X1 _u10_u1_U546  ( .A1(_u10_u1_n2716 ), .A2(_u10_u1_n2717 ), .A3(_u10_u1_n2718 ), .ZN(_u10_u1_n2715 ) );
NAND2_X1 _u10_u1_U545  ( .A1(_u10_u1_n2228 ), .A2(_u10_u1_n2715 ), .ZN(_u10_u1_n2711 ) );
NAND2_X1 _u10_u1_U544  ( .A1(_u10_u1_n2713 ), .A2(_u10_u1_n2714 ), .ZN(_u10_u1_n2712 ) );
NAND3_X1 _u10_u1_U543  ( .A1(_u10_u1_n2710 ), .A2(_u10_u1_n2711 ), .A3(_u10_u1_n2712 ), .ZN(_u10_u1_n2698 ) );
INV_X1 _u10_u1_U542  ( .A(_u10_u1_n2695 ), .ZN(_u10_u1_n2689 ) );
NOR2_X1 _u10_u1_U541  ( .A1(_u10_u1_n2689 ), .A2(_u10_u1_n2709 ), .ZN(_u10_u1_n2708 ) );
NOR3_X1 _u10_u1_U540  ( .A1(_u10_u1_n2706 ), .A2(_u10_u1_n2707 ), .A3(_u10_u1_n2708 ), .ZN(_u10_u1_n2704 ) );
NOR2_X1 _u10_u1_U539  ( .A1(_u10_u1_n2704 ), .A2(_u10_u1_n2705 ), .ZN(_u10_u1_n2699 ) );
NOR2_X1 _u10_u1_U538  ( .A1(_u10_u1_n2702 ), .A2(_u10_u1_n2703 ), .ZN(_u10_u1_n1975 ) );
NOR2_X1 _u10_u1_U537  ( .A1(_u10_u1_n2701 ), .A2(_u10_u1_n1975 ), .ZN(_u10_u1_n2700 ) );
NOR4_X1 _u10_u1_U536  ( .A1(_u10_u1_n2697 ), .A2(_u10_u1_n2698 ), .A3(_u10_u1_n2699 ), .A4(_u10_u1_n2700 ), .ZN(_u10_u1_n2654 ) );
OR2_X1 _u10_u1_U535  ( .A1(_u10_u1_n1852 ), .A2(_u10_u1_n2696 ), .ZN(_u10_u1_n2538 ) );
NAND3_X1 _u10_u1_U534  ( .A1(_u10_u1_n2695 ), .A2(_u10_u1_n2538 ), .A3(_u10_u1_n2201 ), .ZN(_u10_u1_n2676 ) );
NOR4_X1 _u10_u1_U533  ( .A1(_u10_u1_n2692 ), .A2(_u10_u1_n2116 ), .A3(_u10_u1_n2693 ), .A4(_u10_u1_n2694 ), .ZN(_u10_u1_n2691 ) );
NAND4_X1 _u10_u1_U532  ( .A1(_u10_u1_n2689 ), .A2(_u10_u1_n2238 ), .A3(_u10_u1_n2690 ), .A4(_u10_u1_n2691 ), .ZN(_u10_u1_n2688 ) );
NAND2_X1 _u10_u1_U531  ( .A1(_u10_u1_n2263 ), .A2(_u10_u1_n2688 ), .ZN(_u10_u1_n2677 ) );
NAND2_X1 _u10_u1_U530  ( .A1(_u10_u1_n2687 ), .A2(_u10_u1_n2398 ), .ZN(_u10_u1_n2686 ) );
NAND4_X1 _u10_u1_U529  ( .A1(_u10_u1_n2023 ), .A2(_u10_u1_n2686 ), .A3(_u10_u1_n1945 ), .A4(_u10_u1_n2174 ), .ZN(_u10_u1_n2685 ) );
NAND3_X1 _u10_u1_U528  ( .A1(_u10_u1_n2685 ), .A2(_u10_u1_n2022 ), .A3(_u10_u1_n2012 ), .ZN(_u10_u1_n2678 ) );
NOR3_X1 _u10_u1_U527  ( .A1(_u10_u1_n2587 ), .A2(1'b0), .A3(_u10_u1_n2284 ),.ZN(_u10_u1_n2680 ) );
NOR3_X1 _u10_u1_U526  ( .A1(_u10_u1_n2489 ), .A2(_u10_u1_n2684 ), .A3(_u10_u1_n2157 ), .ZN(_u10_u1_n2681 ) );
NOR3_X1 _u10_u1_U525  ( .A1(_u10_u1_n2418 ), .A2(_u10_u1_n1895 ), .A3(_u10_u1_n2683 ), .ZN(_u10_u1_n2682 ) );
NOR3_X1 _u10_u1_U524  ( .A1(_u10_u1_n2680 ), .A2(_u10_u1_n2681 ), .A3(_u10_u1_n2682 ), .ZN(_u10_u1_n2679 ) );
NAND4_X1 _u10_u1_U523  ( .A1(_u10_u1_n2676 ), .A2(_u10_u1_n2677 ), .A3(_u10_u1_n2678 ), .A4(_u10_u1_n2679 ), .ZN(_u10_u1_n2656 ) );
NAND2_X1 _u10_u1_U522  ( .A1(_u10_u1_n1887 ), .A2(_u10_u1_n2295 ), .ZN(_u10_u1_n2675 ) );
AND2_X1 _u10_u1_U521  ( .A1(_u10_u1_n2674 ), .A2(_u10_u1_n2675 ), .ZN(_u10_u1_n2057 ) );
NAND2_X1 _u10_u1_U520  ( .A1(_u10_u1_n2057 ), .A2(_u10_u1_n1868 ), .ZN(_u10_u1_n2673 ) );
NAND2_X1 _u10_u1_U519  ( .A1(_u10_u1_n2673 ), .A2(_u10_u1_n2180 ), .ZN(_u10_u1_n2667 ) );
NAND3_X1 _u10_u1_U518  ( .A1(_u10_u1_n2086 ), .A2(_u10_u1_n2672 ), .A3(1'b0),.ZN(_u10_u1_n2668 ) );
NAND2_X1 _u10_u1_U517  ( .A1(_u10_u1_n2627 ), .A2(_u10_u1_n2250 ), .ZN(_u10_u1_n2670 ) );
NAND2_X1 _u10_u1_U516  ( .A1(_u10_u1_n2670 ), .A2(_u10_u1_n2671 ), .ZN(_u10_u1_n2669 ) );
NAND3_X1 _u10_u1_U515  ( .A1(_u10_u1_n2667 ), .A2(_u10_u1_n2668 ), .A3(_u10_u1_n2669 ), .ZN(_u10_u1_n2657 ) );
NOR2_X1 _u10_u1_U514  ( .A1(_u10_u1_n2198 ), .A2(_u10_u1_n2063 ), .ZN(_u10_u1_n2665 ) );
NOR2_X1 _u10_u1_U513  ( .A1(_u10_u1_n2665 ), .A2(_u10_u1_n2666 ), .ZN(_u10_u1_n2664 ) );
NOR2_X1 _u10_u1_U512  ( .A1(_u10_u1_n2664 ), .A2(_u10_u1_n2420 ), .ZN(_u10_u1_n2658 ) );
NOR2_X1 _u10_u1_U511  ( .A1(_u10_u1_n2662 ), .A2(_u10_u1_n2663 ), .ZN(_u10_u1_n2661 ) );
NOR2_X1 _u10_u1_U510  ( .A1(_u10_u1_n2661 ), .A2(_u10_u1_n1916 ), .ZN(_u10_u1_n2660 ) );
NOR2_X1 _u10_u1_U509  ( .A1(_u10_u1_n2660 ), .A2(_u10_u1_n2353 ), .ZN(_u10_u1_n2659 ) );
NOR4_X1 _u10_u1_U508  ( .A1(_u10_u1_n2656 ), .A2(_u10_u1_n2657 ), .A3(_u10_u1_n2658 ), .A4(_u10_u1_n2659 ), .ZN(_u10_u1_n2655 ) );
NAND4_X1 _u10_u1_U507  ( .A1(_u10_u1_n2652 ), .A2(_u10_u1_n2653 ), .A3(_u10_u1_n2654 ), .A4(_u10_u1_n2655 ), .ZN(_u10_u1_n2651 ) );
MUX2_X1 _u10_u1_U506  ( .A(_u10_u1_n2651 ), .B(_u10_gnt_p0_d[2] ), .S(_u10_u1_n1809 ), .Z(_u10_u1_n1999 ) );
NAND2_X1 _u10_u1_U505  ( .A1(_u10_u1_n2454 ), .A2(_u10_u1_n2314 ), .ZN(_u10_u1_n2644 ) );
NAND2_X1 _u10_u1_U504  ( .A1(_u10_u1_n2012 ), .A2(_u10_u1_n2650 ), .ZN(_u10_u1_n2645 ) );
NOR2_X1 _u10_u1_U503  ( .A1(_u10_u1_n2576 ), .A2(_u10_u1_n2649 ), .ZN(_u10_u1_n2350 ) );
NOR2_X1 _u10_u1_U502  ( .A1(_u10_u1_n2173 ), .A2(_u10_u1_n2321 ), .ZN(_u10_u1_n2647 ) );
NOR2_X1 _u10_u1_U501  ( .A1(_u10_u1_n2169 ), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n2648 ) );
NOR3_X1 _u10_u1_U500  ( .A1(_u10_u1_n2350 ), .A2(_u10_u1_n2647 ), .A3(_u10_u1_n2648 ), .ZN(_u10_u1_n2646 ) );
NAND3_X1 _u10_u1_U499  ( .A1(_u10_u1_n2644 ), .A2(_u10_u1_n2645 ), .A3(_u10_u1_n2646 ), .ZN(_u10_u1_n2555 ) );
NOR2_X1 _u10_u1_U498  ( .A1(1'b0), .A2(_u10_u1_n2643 ), .ZN(_u10_u1_n2641 ));
NAND2_X1 _u10_u1_U497  ( .A1(_u10_u1_n2406 ), .A2(_u10_u1_n1955 ), .ZN(_u10_u1_n2642 ) );
NAND3_X1 _u10_u1_U496  ( .A1(_u10_u1_n2104 ), .A2(_u10_u1_n2155 ), .A3(1'b0),.ZN(_u10_u1_n2629 ) );
NAND4_X1 _u10_u1_U495  ( .A1(_u10_u1_n2642 ), .A2(_u10_u1_n2240 ), .A3(_u10_u1_n2629 ), .A4(_u10_u1_n2392 ), .ZN(_u10_u1_n2099 ) );
NOR2_X1 _u10_u1_U494  ( .A1(_u10_u1_n2641 ), .A2(_u10_u1_n2099 ), .ZN(_u10_u1_n2640 ) );
NOR2_X1 _u10_u1_U493  ( .A1(_u10_u1_n2640 ), .A2(_u10_u1_n2223 ), .ZN(_u10_u1_n2637 ) );
NOR2_X1 _u10_u1_U492  ( .A1(_u10_u1_n2474 ), .A2(_u10_u1_n2608 ), .ZN(_u10_u1_n2639 ) );
NOR2_X1 _u10_u1_U491  ( .A1(_u10_u1_n2639 ), .A2(_u10_u1_n2576 ), .ZN(_u10_u1_n2638 ) );
NOR2_X1 _u10_u1_U490  ( .A1(_u10_u1_n2637 ), .A2(_u10_u1_n2638 ), .ZN(_u10_u1_n2599 ) );
NAND2_X1 _u10_u1_U489  ( .A1(_u10_u1_n2139 ), .A2(_u10_u1_n2636 ), .ZN(_u10_u1_n2635 ) );
NAND2_X1 _u10_u1_U488  ( .A1(_u10_u1_n2634 ), .A2(_u10_u1_n2635 ), .ZN(_u10_u1_n2600 ) );
NOR4_X1 _u10_u1_U487  ( .A1(1'b0), .A2(_u10_u1_n2019 ), .A3(_u10_u1_n2632 ),.A4(_u10_u1_n2633 ), .ZN(_u10_u1_n2622 ) );
NOR3_X1 _u10_u1_U486  ( .A1(_u10_u1_n2064 ), .A2(1'b0), .A3(_u10_u1_n2420 ),.ZN(_u10_u1_n2623 ) );
NOR2_X1 _u10_u1_U485  ( .A1(_u10_u1_n2631 ), .A2(_u10_u1_n2373 ), .ZN(_u10_u1_n2630 ) );
NOR2_X1 _u10_u1_U484  ( .A1(_u10_u1_n2630 ), .A2(_u10_u1_n1825 ), .ZN(_u10_u1_n2624 ) );
NOR3_X1 _u10_u1_U483  ( .A1(1'b0), .A2(1'b0), .A3(_u10_u1_n2629 ), .ZN(_u10_u1_n2598 ) );
NAND3_X1 _u10_u1_U482  ( .A1(_u10_u1_n2201 ), .A2(_u10_u1_n1875 ), .A3(_u10_u1_n2598 ), .ZN(_u10_u1_n1878 ) );
NOR2_X1 _u10_u1_U481  ( .A1(_u10_u1_n1878 ), .A2(_u10_u1_n1883 ), .ZN(_u10_u1_n1835 ) );
INV_X1 _u10_u1_U480  ( .A(_u10_u1_n1835 ), .ZN(_u10_u1_n2500 ) );
NAND2_X1 _u10_u1_U479  ( .A1(_u10_u1_n2500 ), .A2(_u10_u1_n2628 ), .ZN(_u10_u1_n2089 ) );
NOR2_X1 _u10_u1_U478  ( .A1(_u10_u1_n2133 ), .A2(_u10_u1_n2089 ), .ZN(_u10_u1_n2626 ) );
NOR2_X1 _u10_u1_U477  ( .A1(_u10_u1_n2626 ), .A2(_u10_u1_n2627 ), .ZN(_u10_u1_n2625 ) );
NOR4_X1 _u10_u1_U476  ( .A1(_u10_u1_n2622 ), .A2(_u10_u1_n2623 ), .A3(_u10_u1_n2624 ), .A4(_u10_u1_n2625 ), .ZN(_u10_u1_n2601 ) );
NAND2_X1 _u10_u1_U475  ( .A1(1'b0), .A2(_u10_u1_n2136 ), .ZN(_u10_u1_n2006 ));
NOR3_X1 _u10_u1_U474  ( .A1(_u10_u1_n2621 ), .A2(1'b0), .A3(_u10_u1_n2006 ),.ZN(_u10_u1_n1989 ) );
NAND2_X1 _u10_u1_U473  ( .A1(_u10_u1_n1989 ), .A2(_u10_u1_n1898 ), .ZN(_u10_u1_n2609 ) );
NAND2_X1 _u10_u1_U472  ( .A1(_u10_u1_n2047 ), .A2(_u10_u1_n2089 ), .ZN(_u10_u1_n2610 ) );
NOR3_X1 _u10_u1_U471  ( .A1(_u10_u1_n2620 ), .A2(_u10_u1_n2007 ), .A3(_u10_u1_n2006 ), .ZN(_u10_u1_n2145 ) );
NAND2_X1 _u10_u1_U470  ( .A1(_u10_u1_n2145 ), .A2(_u10_u1_n2619 ), .ZN(_u10_u1_n1967 ) );
INV_X1 _u10_u1_U469  ( .A(_u10_u1_n1967 ), .ZN(_u10_u1_n1831 ) );
NAND2_X1 _u10_u1_U468  ( .A1(_u10_u1_n1831 ), .A2(_u10_u1_n2618 ), .ZN(_u10_u1_n2551 ) );
INV_X1 _u10_u1_U467  ( .A(_u10_u1_n2551 ), .ZN(_u10_u1_n1942 ) );
NAND2_X1 _u10_u1_U466  ( .A1(_u10_u1_n1942 ), .A2(_u10_u1_n2105 ), .ZN(_u10_u1_n2120 ) );
INV_X1 _u10_u1_U465  ( .A(_u10_u1_n2120 ), .ZN(_u10_u1_n2616 ) );
NAND2_X1 _u10_u1_U464  ( .A1(_u10_u1_n2616 ), .A2(_u10_u1_n2617 ), .ZN(_u10_u1_n2611 ) );
NAND3_X1 _u10_u1_U463  ( .A1(_u10_u1_n2398 ), .A2(_u10_u1_n1844 ), .A3(_u10_u1_n2616 ), .ZN(_u10_u1_n2614 ) );
NAND2_X1 _u10_u1_U462  ( .A1(_u10_u1_n2133 ), .A2(_u10_u1_n2023 ), .ZN(_u10_u1_n2615 ) );
NAND3_X1 _u10_u1_U461  ( .A1(_u10_u1_n2614 ), .A2(_u10_u1_n2022 ), .A3(_u10_u1_n2615 ), .ZN(_u10_u1_n2613 ) );
NAND2_X1 _u10_u1_U460  ( .A1(_u10_u1_n2012 ), .A2(_u10_u1_n2613 ), .ZN(_u10_u1_n2612 ) );
NAND4_X1 _u10_u1_U459  ( .A1(_u10_u1_n2609 ), .A2(_u10_u1_n2610 ), .A3(_u10_u1_n2611 ), .A4(_u10_u1_n2612 ), .ZN(_u10_u1_n2603 ) );
AND2_X1 _u10_u1_U458  ( .A1(_u10_u1_n1920 ), .A2(_u10_u1_n2608 ), .ZN(_u10_u1_n2604 ) );
NOR2_X1 _u10_u1_U457  ( .A1(_u10_u1_n2465 ), .A2(_u10_u1_n1878 ), .ZN(_u10_u1_n2605 ) );
NOR2_X1 _u10_u1_U456  ( .A1(_u10_u1_n2059 ), .A2(_u10_u1_n2607 ), .ZN(_u10_u1_n2606 ) );
NOR4_X1 _u10_u1_U455  ( .A1(_u10_u1_n2603 ), .A2(_u10_u1_n2604 ), .A3(_u10_u1_n2605 ), .A4(_u10_u1_n2606 ), .ZN(_u10_u1_n2602 ) );
AND4_X1 _u10_u1_U454  ( .A1(_u10_u1_n2599 ), .A2(_u10_u1_n2600 ), .A3(_u10_u1_n2601 ), .A4(_u10_u1_n2602 ), .ZN(_u10_u1_n2033 ) );
INV_X1 _u10_u1_U453  ( .A(_u10_u1_n2598 ), .ZN(_u10_u1_n2071 ) );
NAND2_X1 _u10_u1_U452  ( .A1(_u10_u1_n2597 ), .A2(_u10_u1_n2071 ), .ZN(_u10_u1_n2112 ) );
INV_X1 _u10_u1_U451  ( .A(_u10_u1_n2112 ), .ZN(_u10_u1_n2422 ) );
NAND2_X1 _u10_u1_U450  ( .A1(_u10_u1_n2422 ), .A2(_u10_u1_n2596 ), .ZN(_u10_u1_n2571 ) );
NAND2_X1 _u10_u1_U449  ( .A1(_u10_u1_n2263 ), .A2(_u10_u1_n2571 ), .ZN(_u10_u1_n2560 ) );
NAND3_X1 _u10_u1_U448  ( .A1(_u10_u1_n1886 ), .A2(_u10_u1_n2399 ), .A3(1'b0),.ZN(_u10_u1_n2185 ) );
NOR3_X1 _u10_u1_U447  ( .A1(_u10_u1_n2225 ), .A2(_u10_u1_n2314 ), .A3(_u10_u1_n2185 ), .ZN(_u10_u1_n2379 ) );
NAND2_X1 _u10_u1_U446  ( .A1(_u10_u1_n2379 ), .A2(_u10_u1_n2595 ), .ZN(_u10_u1_n2561 ) );
NOR2_X1 _u10_u1_U445  ( .A1(_u10_u1_n2480 ), .A2(_u10_u1_n2379 ), .ZN(_u10_u1_n2578 ) );
INV_X1 _u10_u1_U444  ( .A(_u10_u1_n2578 ), .ZN(_u10_u1_n2307 ) );
NOR2_X1 _u10_u1_U443  ( .A1(_u10_u1_n2307 ), .A2(_u10_u1_n2089 ), .ZN(_u10_u1_n2245 ) );
NOR2_X1 _u10_u1_U442  ( .A1(_u10_u1_n2594 ), .A2(_u10_u1_n2245 ), .ZN(_u10_u1_n2590 ) );
NOR2_X1 _u10_u1_U441  ( .A1(_u10_u1_n2592 ), .A2(_u10_u1_n2593 ), .ZN(_u10_u1_n2591 ) );
NOR2_X1 _u10_u1_U440  ( .A1(_u10_u1_n2590 ), .A2(_u10_u1_n2591 ), .ZN(_u10_u1_n2562 ) );
INV_X1 _u10_u1_U439  ( .A(_u10_u1_n2589 ), .ZN(_u10_u1_n2584 ) );
INV_X1 _u10_u1_U438  ( .A(_u10_u1_n2588 ), .ZN(_u10_u1_n2204 ) );
NAND2_X1 _u10_u1_U437  ( .A1(_u10_u1_n2204 ), .A2(_u10_u1_n1875 ), .ZN(_u10_u1_n2585 ) );
AND3_X1 _u10_u1_U436  ( .A1(_u10_u1_n2587 ), .A2(_u10_u1_n2466 ), .A3(_u10_u1_n1878 ), .ZN(_u10_u1_n2586 ) );
AND3_X1 _u10_u1_U435  ( .A1(_u10_u1_n2584 ), .A2(_u10_u1_n2585 ), .A3(_u10_u1_n2586 ), .ZN(_u10_u1_n2186 ) );
NOR2_X1 _u10_u1_U434  ( .A1(1'b0), .A2(_u10_u1_n2186 ), .ZN(_u10_u1_n2582 ));
NOR2_X1 _u10_u1_U433  ( .A1(_u10_u1_n2225 ), .A2(_u10_u1_n2185 ), .ZN(_u10_u1_n2583 ) );
NOR2_X1 _u10_u1_U432  ( .A1(_u10_u1_n2582 ), .A2(_u10_u1_n2583 ), .ZN(_u10_u1_n2581 ) );
NOR2_X1 _u10_u1_U431  ( .A1(_u10_u1_n2581 ), .A2(_u10_u1_n2284 ), .ZN(_u10_u1_n2564 ) );
NOR2_X1 _u10_u1_U430  ( .A1(_u10_u1_n2580 ), .A2(_u10_u1_n2307 ), .ZN(_u10_u1_n2579 ) );
NOR2_X1 _u10_u1_U429  ( .A1(_u10_u1_n2579 ), .A2(_u10_u1_n2169 ), .ZN(_u10_u1_n2565 ) );
NOR2_X1 _u10_u1_U428  ( .A1(_u10_u1_n2500 ), .A2(_u10_u1_n1919 ), .ZN(_u10_u1_n2577 ) );
NOR2_X1 _u10_u1_U427  ( .A1(_u10_u1_n1919 ), .A2(_u10_u1_n2578 ), .ZN(_u10_u1_n2332 ) );
NOR3_X1 _u10_u1_U426  ( .A1(_u10_u1_n2577 ), .A2(1'b0), .A3(_u10_u1_n2332 ),.ZN(_u10_u1_n2575 ) );
NOR2_X1 _u10_u1_U425  ( .A1(_u10_u1_n2575 ), .A2(_u10_u1_n2576 ), .ZN(_u10_u1_n2566 ) );
NOR2_X1 _u10_u1_U424  ( .A1(_u10_u1_n2574 ), .A2(_u10_u1_n2155 ), .ZN(_u10_u1_n2573 ) );
NOR2_X1 _u10_u1_U423  ( .A1(_u10_u1_n2573 ), .A2(_u10_u1_n2196 ), .ZN(_u10_u1_n2572 ) );
NOR2_X1 _u10_u1_U422  ( .A1(_u10_u1_n2572 ), .A2(_u10_u1_n2287 ), .ZN(_u10_u1_n2569 ) );
AND2_X1 _u10_u1_U421  ( .A1(_u10_u1_n2065 ), .A2(_u10_u1_n2571 ), .ZN(_u10_u1_n2570 ) );
NOR2_X1 _u10_u1_U420  ( .A1(_u10_u1_n2569 ), .A2(_u10_u1_n2570 ), .ZN(_u10_u1_n2568 ) );
NOR2_X1 _u10_u1_U419  ( .A1(_u10_u1_n2568 ), .A2(_u10_u1_n2059 ), .ZN(_u10_u1_n2567 ) );
NOR4_X1 _u10_u1_U418  ( .A1(_u10_u1_n2564 ), .A2(_u10_u1_n2565 ), .A3(_u10_u1_n2566 ), .A4(_u10_u1_n2567 ), .ZN(_u10_u1_n2563 ) );
AND4_X1 _u10_u1_U417  ( .A1(_u10_u1_n2560 ), .A2(_u10_u1_n2561 ), .A3(_u10_u1_n2562 ), .A4(_u10_u1_n2563 ), .ZN(_u10_u1_n2335 ) );
NAND3_X1 _u10_u1_U416  ( .A1(_u10_u1_n2033 ), .A2(_u10_u1_n2559 ), .A3(_u10_u1_n2335 ), .ZN(_u10_u1_n2556 ) );
NOR4_X1 _u10_u1_U415  ( .A1(_u10_u1_n2555 ), .A2(_u10_u1_n2556 ), .A3(_u10_u1_n2557 ), .A4(_u10_u1_n2558 ), .ZN(_u10_u1_n2358 ) );
NOR2_X1 _u10_u1_U414  ( .A1(_u10_u1_n1910 ), .A2(_u10_u1_n1920 ), .ZN(_u10_u1_n2371 ) );
OR2_X1 _u10_u1_U413  ( .A1(_u10_u1_n2489 ), .A2(_u10_u1_n2371 ), .ZN(_u10_u1_n2510 ) );
NOR3_X1 _u10_u1_U412  ( .A1(_u10_u1_n2157 ), .A2(_u10_u1_n2007 ), .A3(_u10_u1_n2136 ), .ZN(_u10_u1_n2381 ) );
INV_X1 _u10_u1_U411  ( .A(_u10_u1_n2381 ), .ZN(_u10_u1_n2523 ) );
NAND3_X1 _u10_u1_U410  ( .A1(_u10_u1_n2523 ), .A2(_u10_u1_n2155 ), .A3(_u10_u1_n2532 ), .ZN(_u10_u1_n2554 ) );
NAND2_X1 _u10_u1_U409  ( .A1(_u10_u1_n2104 ), .A2(_u10_u1_n2554 ), .ZN(_u10_u1_n2546 ) );
INV_X1 _u10_u1_U408  ( .A(_u10_u1_n2553 ), .ZN(_u10_u1_n2547 ) );
NAND4_X1 _u10_u1_U407  ( .A1(_u10_u1_n2549 ), .A2(_u10_u1_n2550 ), .A3(_u10_u1_n2551 ), .A4(_u10_u1_n2552 ), .ZN(_u10_u1_n2408 ) );
NAND2_X1 _u10_u1_U406  ( .A1(_u10_u1_n2408 ), .A2(_u10_u1_n1955 ), .ZN(_u10_u1_n2548 ) );
NAND3_X1 _u10_u1_U405  ( .A1(_u10_u1_n2546 ), .A2(_u10_u1_n2547 ), .A3(_u10_u1_n2548 ), .ZN(_u10_u1_n2545 ) );
NAND2_X1 _u10_u1_U404  ( .A1(_u10_u1_n1950 ), .A2(_u10_u1_n2545 ), .ZN(_u10_u1_n2511 ) );
NAND2_X1 _u10_u1_U403  ( .A1(_u10_u1_n2381 ), .A2(_u10_u1_n1885 ), .ZN(_u10_u1_n2543 ) );
NAND4_X1 _u10_u1_U402  ( .A1(_u10_u1_n2543 ), .A2(_u10_u1_n2458 ), .A3(_u10_u1_n2120 ), .A4(_u10_u1_n2544 ), .ZN(_u10_u1_n2391 ) );
NAND2_X1 _u10_u1_U401  ( .A1(_u10_u1_n1886 ), .A2(_u10_u1_n2391 ), .ZN(_u10_u1_n2542 ) );
NAND4_X1 _u10_u1_U400  ( .A1(_u10_u1_n2540 ), .A2(_u10_u1_n2541 ), .A3(_u10_u1_n2542 ), .A4(_u10_u1_n2185 ), .ZN(_u10_u1_n2539 ) );
NAND2_X1 _u10_u1_U399  ( .A1(_u10_u1_n2538 ), .A2(_u10_u1_n2539 ), .ZN(_u10_u1_n2512 ) );
OR2_X1 _u10_u1_U398  ( .A1(_u10_u1_n2537 ), .A2(_u10_u1_n12 ), .ZN(_u10_u1_n2536 ) );
NOR2_X1 _u10_u1_U397  ( .A1(_u10_u1_n2521 ), .A2(_u10_u1_n1831 ), .ZN(_u10_u1_n2156 ) );
NAND3_X1 _u10_u1_U396  ( .A1(_u10_u1_n2536 ), .A2(_u10_u1_n2156 ), .A3(_u10_u1_n2310 ), .ZN(_u10_u1_n2530 ) );
NOR3_X1 _u10_u1_U395  ( .A1(_u10_u1_n2534 ), .A2(_u10_u1_n2381 ), .A3(_u10_u1_n2535 ), .ZN(_u10_u1_n2533 ) );
NAND3_X1 _u10_u1_U394  ( .A1(_u10_u1_n1963 ), .A2(_u10_u1_n2532 ), .A3(_u10_u1_n2533 ), .ZN(_u10_u1_n2409 ) );
NOR3_X1 _u10_u1_U393  ( .A1(_u10_u1_n2530 ), .A2(_u10_u1_n2409 ), .A3(_u10_u1_n2531 ), .ZN(_u10_u1_n2528 ) );
NOR2_X1 _u10_u1_U392  ( .A1(_u10_u1_n2528 ), .A2(_u10_u1_n2529 ), .ZN(_u10_u1_n2514 ) );
NOR2_X1 _u10_u1_U391  ( .A1(_u10_u1_n2500 ), .A2(_u10_u1_n2527 ), .ZN(_u10_u1_n2515 ) );
NAND3_X1 _u10_u1_U390  ( .A1(_u10_u1_n1891 ), .A2(_u10_u1_n2525 ), .A3(_u10_u1_n2526 ), .ZN(_u10_u1_n2518 ) );
NAND4_X1 _u10_u1_U389  ( .A1(_u10_u1_n2489 ), .A2(_u10_u1_n1967 ), .A3(_u10_u1_n2523 ), .A4(_u10_u1_n2524 ), .ZN(_u10_u1_n2395 ) );
NAND3_X1 _u10_u1_U388  ( .A1(_u10_u1_n2398 ), .A2(_u10_u1_n2399 ), .A3(_u10_u1_n2522 ), .ZN(_u10_u1_n2519 ) );
NOR3_X1 _u10_u1_U387  ( .A1(_u10_u1_n2312 ), .A2(1'b0), .A3(_u10_u1_n2521 ),.ZN(_u10_u1_n2520 ) );
NAND3_X1 _u10_u1_U386  ( .A1(_u10_u1_n2310 ), .A2(_u10_u1_n2519 ), .A3(_u10_u1_n2520 ), .ZN(_u10_u1_n2328 ) );
NOR3_X1 _u10_u1_U385  ( .A1(_u10_u1_n2518 ), .A2(_u10_u1_n2395 ), .A3(_u10_u1_n2328 ), .ZN(_u10_u1_n2517 ) );
NOR2_X1 _u10_u1_U384  ( .A1(_u10_u1_n2517 ), .A2(_u10_u1_n1830 ), .ZN(_u10_u1_n2516 ) );
NOR3_X1 _u10_u1_U383  ( .A1(_u10_u1_n2514 ), .A2(_u10_u1_n2515 ), .A3(_u10_u1_n2516 ), .ZN(_u10_u1_n2513 ) );
NAND4_X1 _u10_u1_U382  ( .A1(_u10_u1_n2510 ), .A2(_u10_u1_n2511 ), .A3(_u10_u1_n2512 ), .A4(_u10_u1_n2513 ), .ZN(_u10_u1_n2460 ) );
NAND2_X1 _u10_u1_U381  ( .A1(_u10_u1_n2451 ), .A2(_u10_u1_n2245 ), .ZN(_u10_u1_n2509 ) );
NAND2_X1 _u10_u1_U380  ( .A1(_u10_u1_n2508 ), .A2(_u10_u1_n2509 ), .ZN(_u10_u1_n2502 ) );
NOR2_X1 _u10_u1_U379  ( .A1(_u10_u1_n2506 ), .A2(_u10_u1_n2507 ), .ZN(_u10_u1_n2369 ) );
NAND2_X1 _u10_u1_U378  ( .A1(_u10_u1_n2369 ), .A2(_u10_u1_n1844 ), .ZN(_u10_u1_n2449 ) );
NAND2_X1 _u10_u1_U377  ( .A1(_u10_u1_n2449 ), .A2(_u10_u1_n2505 ), .ZN(_u10_u1_n2504 ) );
NAND3_X1 _u10_u1_U376  ( .A1(_u10_u1_n2502 ), .A2(_u10_u1_n2503 ), .A3(_u10_u1_n2504 ), .ZN(_u10_u1_n2501 ) );
NAND2_X1 _u10_u1_U375  ( .A1(_u10_u1_n2322 ), .A2(_u10_u1_n2501 ), .ZN(_u10_u1_n2467 ) );
NAND2_X1 _u10_u1_U374  ( .A1(_u10_u1_n2045 ), .A2(_u10_u1_n2500 ), .ZN(_u10_u1_n2499 ) );
NAND2_X1 _u10_u1_U373  ( .A1(_u10_u1_n2295 ), .A2(_u10_u1_n2499 ), .ZN(_u10_u1_n2488 ) );
NOR3_X1 _u10_u1_U372  ( .A1(_u10_u1_n2497 ), .A2(_u10_u1_n2145 ), .A3(_u10_u1_n2498 ), .ZN(_u10_u1_n2490 ) );
NOR2_X1 _u10_u1_U371  ( .A1(_u10_u1_n2007 ), .A2(_u10_u1_n2136 ), .ZN(_u10_u1_n2492 ) );
NAND2_X1 _u10_u1_U370  ( .A1(_u10_u1_n2379 ), .A2(_u10_u1_n2295 ), .ZN(_u10_u1_n2496 ) );
NAND3_X1 _u10_u1_U369  ( .A1(_u10_u1_n2494 ), .A2(_u10_u1_n2495 ), .A3(_u10_u1_n2496 ), .ZN(_u10_u1_n2270 ) );
NOR4_X1 _u10_u1_U368  ( .A1(_u10_u1_n2492 ), .A2(_u10_u1_n2396 ), .A3(_u10_u1_n2270 ), .A4(_u10_u1_n2493 ), .ZN(_u10_u1_n2491 ) );
NAND4_X1 _u10_u1_U367  ( .A1(_u10_u1_n2488 ), .A2(_u10_u1_n2489 ), .A3(_u10_u1_n2490 ), .A4(_u10_u1_n2491 ), .ZN(_u10_u1_n2487 ) );
NAND2_X1 _u10_u1_U366  ( .A1(_u10_u1_n2146 ), .A2(_u10_u1_n2487 ), .ZN(_u10_u1_n2468 ) );
NAND2_X1 _u10_u1_U365  ( .A1(_u10_u1_n2379 ), .A2(_u10_u1_n2486 ), .ZN(_u10_u1_n2485 ) );
AND2_X1 _u10_u1_U364  ( .A1(_u10_u1_n2484 ), .A2(_u10_u1_n2485 ), .ZN(_u10_u1_n2256 ) );
NOR2_X1 _u10_u1_U363  ( .A1(_u10_u1_n2483 ), .A2(_u10_u1_n2007 ), .ZN(_u10_u1_n2481 ) );
NOR2_X1 _u10_u1_U362  ( .A1(_u10_u1_n2481 ), .A2(_u10_u1_n2482 ), .ZN(_u10_u1_n2472 ) );
NOR3_X1 _u10_u1_U361  ( .A1(_u10_u1_n1835 ), .A2(1'b0), .A3(_u10_u1_n2480 ),.ZN(_u10_u1_n2479 ) );
NOR2_X1 _u10_u1_U360  ( .A1(_u10_u1_n2479 ), .A2(_u10_u1_n2010 ), .ZN(_u10_u1_n2476 ) );
NOR2_X1 _u10_u1_U359  ( .A1(_u10_u1_n2478 ), .A2(_u10_u1_n2045 ), .ZN(_u10_u1_n2477 ) );
NOR4_X1 _u10_u1_U358  ( .A1(_u10_u1_n2474 ), .A2(_u10_u1_n2475 ), .A3(_u10_u1_n2476 ), .A4(_u10_u1_n2477 ), .ZN(_u10_u1_n2473 ) );
NAND4_X1 _u10_u1_U357  ( .A1(_u10_u1_n2471 ), .A2(_u10_u1_n2256 ), .A3(_u10_u1_n2472 ), .A4(_u10_u1_n2473 ), .ZN(_u10_u1_n2470 ) );
NAND2_X1 _u10_u1_U356  ( .A1(_u10_u1_n2228 ), .A2(_u10_u1_n2470 ), .ZN(_u10_u1_n2469 ) );
NAND3_X1 _u10_u1_U355  ( .A1(_u10_u1_n2467 ), .A2(_u10_u1_n2468 ), .A3(_u10_u1_n2469 ), .ZN(_u10_u1_n2461 ) );
NOR2_X1 _u10_u1_U354  ( .A1(_u10_u1_n2465 ), .A2(_u10_u1_n2466 ), .ZN(_u10_u1_n2462 ) );
NOR2_X1 _u10_u1_U353  ( .A1(_u10_u1_n2464 ), .A2(_u10_u1_n2019 ), .ZN(_u10_u1_n2463 ) );
NOR4_X1 _u10_u1_U352  ( .A1(_u10_u1_n2460 ), .A2(_u10_u1_n2461 ), .A3(_u10_u1_n2462 ), .A4(_u10_u1_n2463 ), .ZN(_u10_u1_n2359 ) );
NAND2_X1 _u10_u1_U351  ( .A1(_u10_u1_n2453 ), .A2(_u10_u1_n2459 ), .ZN(_u10_u1_n2443 ) );
NAND2_X1 _u10_u1_U350  ( .A1(_u10_u1_n2099 ), .A2(_u10_u1_n2063 ), .ZN(_u10_u1_n2456 ) );
NAND2_X1 _u10_u1_U349  ( .A1(_u10_u1_n2381 ), .A2(_u10_u1_n2399 ), .ZN(_u10_u1_n2457 ) );
NAND4_X1 _u10_u1_U348  ( .A1(_u10_u1_n2456 ), .A2(_u10_u1_n2457 ), .A3(_u10_u1_n2458 ), .A4(_u10_u1_n2120 ), .ZN(_u10_u1_n2455 ) );
NAND2_X1 _u10_u1_U347  ( .A1(_u10_u1_n2236 ), .A2(_u10_u1_n2455 ), .ZN(_u10_u1_n2444 ) );
NOR3_X1 _u10_u1_U346  ( .A1(_u10_u1_n2276 ), .A2(_u10_u1_n2453 ), .A3(_u10_u1_n2454 ), .ZN(_u10_u1_n2452 ) );
NOR2_X1 _u10_u1_U345  ( .A1(_u10_u1_n2245 ), .A2(_u10_u1_n2452 ), .ZN(_u10_u1_n2446 ) );
NOR2_X1 _u10_u1_U344  ( .A1(_u10_u1_n2451 ), .A2(_u10_u1_n2250 ), .ZN(_u10_u1_n2447 ) );
AND2_X1 _u10_u1_U343  ( .A1(_u10_u1_n2449 ), .A2(_u10_u1_n2450 ), .ZN(_u10_u1_n2448 ) );
NOR3_X1 _u10_u1_U342  ( .A1(_u10_u1_n2446 ), .A2(_u10_u1_n2447 ), .A3(_u10_u1_n2448 ), .ZN(_u10_u1_n2445 ) );
NAND3_X1 _u10_u1_U341  ( .A1(_u10_u1_n2443 ), .A2(_u10_u1_n2444 ), .A3(_u10_u1_n2445 ), .ZN(_u10_u1_n2410 ) );
INV_X1 _u10_u1_U340  ( .A(_u10_u1_n2391 ), .ZN(_u10_u1_n2441 ) );
NAND2_X1 _u10_u1_U339  ( .A1(_u10_u1_n2441 ), .A2(_u10_u1_n2442 ), .ZN(_u10_u1_n2440 ) );
NAND2_X1 _u10_u1_U338  ( .A1(_u10_u1_n2234 ), .A2(_u10_u1_n2440 ), .ZN(_u10_u1_n2437 ) );
NAND3_X1 _u10_u1_U337  ( .A1(_u10_u1_n2078 ), .A2(_u10_u1_n2391 ), .A3(_u10_u1_n2439 ), .ZN(_u10_u1_n2438 ) );
NAND2_X1 _u10_u1_U336  ( .A1(_u10_u1_n2437 ), .A2(_u10_u1_n2438 ), .ZN(_u10_u1_n2436 ) );
NAND2_X1 _u10_u1_U335  ( .A1(_u10_u1_n2074 ), .A2(_u10_u1_n2436 ), .ZN(_u10_u1_n2424 ) );
NAND2_X1 _u10_u1_U334  ( .A1(_u10_u1_n2434 ), .A2(_u10_u1_n2435 ), .ZN(_u10_u1_n2432 ) );
NAND2_X1 _u10_u1_U333  ( .A1(1'b0), .A2(_u10_u1_n1827 ), .ZN(_u10_u1_n2433 ));
NAND2_X1 _u10_u1_U332  ( .A1(_u10_u1_n2432 ), .A2(_u10_u1_n2433 ), .ZN(_u10_u1_n2431 ) );
NAND2_X1 _u10_u1_U331  ( .A1(_u10_u1_n2430 ), .A2(_u10_u1_n2431 ), .ZN(_u10_u1_n2425 ) );
NAND2_X1 _u10_u1_U330  ( .A1(1'b0), .A2(_u10_u1_n2399 ), .ZN(_u10_u1_n2429 ));
NAND2_X1 _u10_u1_U329  ( .A1(_u10_u1_n2238 ), .A2(_u10_u1_n2429 ), .ZN(_u10_u1_n2427 ) );
NAND2_X1 _u10_u1_U328  ( .A1(_u10_u1_n2427 ), .A2(_u10_u1_n2428 ), .ZN(_u10_u1_n2426 ) );
NAND3_X1 _u10_u1_U327  ( .A1(_u10_u1_n2424 ), .A2(_u10_u1_n2425 ), .A3(_u10_u1_n2426 ), .ZN(_u10_u1_n2411 ) );
NOR2_X1 _u10_u1_U326  ( .A1(_u10_u1_n2422 ), .A2(_u10_u1_n2423 ), .ZN(_u10_u1_n2421 ) );
NOR2_X1 _u10_u1_U325  ( .A1(_u10_u1_n2421 ), .A2(_u10_u1_n2203 ), .ZN(_u10_u1_n2419 ) );
NOR2_X1 _u10_u1_U324  ( .A1(_u10_u1_n2419 ), .A2(_u10_u1_n2420 ), .ZN(_u10_u1_n2412 ) );
NAND2_X1 _u10_u1_U323  ( .A1(_u10_u1_n2277 ), .A2(_u10_u1_n2418 ), .ZN(_u10_u1_n2416 ) );
NOR4_X1 _u10_u1_U322  ( .A1(_u10_u1_n2415 ), .A2(_u10_u1_n2416 ), .A3(_u10_u1_n2417 ), .A4(_u10_u1_n2307 ), .ZN(_u10_u1_n2414 ) );
NOR2_X1 _u10_u1_U321  ( .A1(_u10_u1_n2414 ), .A2(_u10_u1_n2020 ), .ZN(_u10_u1_n2413 ) );
NOR4_X1 _u10_u1_U320  ( .A1(_u10_u1_n2410 ), .A2(_u10_u1_n2411 ), .A3(_u10_u1_n2412 ), .A4(_u10_u1_n2413 ), .ZN(_u10_u1_n2360 ) );
NAND2_X1 _u10_u1_U319  ( .A1(_u10_u1_n2106 ), .A2(_u10_u1_n2409 ), .ZN(_u10_u1_n2402 ) );
INV_X1 _u10_u1_U318  ( .A(_u10_u1_n2408 ), .ZN(_u10_u1_n2404 ) );
NOR3_X1 _u10_u1_U317  ( .A1(_u10_u1_n2406 ), .A2(_u10_u1_n2407 ), .A3(_u10_u1_n1941 ), .ZN(_u10_u1_n2405 ) );
NAND4_X1 _u10_u1_U316  ( .A1(_u10_u1_n2402 ), .A2(_u10_u1_n2403 ), .A3(_u10_u1_n2404 ), .A4(_u10_u1_n2405 ), .ZN(_u10_u1_n2401 ) );
NAND2_X1 _u10_u1_U315  ( .A1(_u10_u1_n2230 ), .A2(_u10_u1_n2401 ), .ZN(_u10_u1_n2384 ) );
NOR3_X1 _u10_u1_U314  ( .A1(_u10_u1_n1980 ), .A2(_u10_u1_n2369 ), .A3(_u10_u1_n2400 ), .ZN(_u10_u1_n2386 ) );
NAND4_X1 _u10_u1_U313  ( .A1(_u10_u1_n2397 ), .A2(_u10_u1_n2398 ), .A3(_u10_u1_n2399 ), .A4(_u10_u1_n2155 ), .ZN(_u10_u1_n2352 ) );
NAND4_X1 _u10_u1_U312  ( .A1(_u10_u1_n2294 ), .A2(_u10_u1_n2293 ), .A3(_u10_u1_n2352 ), .A4(_u10_u1_n1966 ), .ZN(_u10_u1_n2394 ) );
NOR4_X1 _u10_u1_U311  ( .A1(_u10_u1_n2394 ), .A2(_u10_u1_n2270 ), .A3(_u10_u1_n2395 ), .A4(_u10_u1_n2396 ), .ZN(_u10_u1_n2393 ) );
NOR2_X1 _u10_u1_U310  ( .A1(_u10_u1_n2393 ), .A2(_u10_u1_n2351 ), .ZN(_u10_u1_n2387 ) );
NOR2_X1 _u10_u1_U309  ( .A1(1'b0), .A2(_u10_u1_n2392 ), .ZN(_u10_u1_n2390 ));
NOR2_X1 _u10_u1_U308  ( .A1(_u10_u1_n2390 ), .A2(_u10_u1_n2391 ), .ZN(_u10_u1_n2389 ) );
NOR3_X1 _u10_u1_U307  ( .A1(_u10_u1_n2110 ), .A2(1'b0), .A3(_u10_u1_n2389 ),.ZN(_u10_u1_n2388 ) );
NOR3_X1 _u10_u1_U306  ( .A1(_u10_u1_n2386 ), .A2(_u10_u1_n2387 ), .A3(_u10_u1_n2388 ), .ZN(_u10_u1_n2385 ) );
NAND4_X1 _u10_u1_U305  ( .A1(_u10_u1_n2382 ), .A2(_u10_u1_n2383 ), .A3(_u10_u1_n2384 ), .A4(_u10_u1_n2385 ), .ZN(_u10_u1_n2362 ) );
NAND3_X1 _u10_u1_U304  ( .A1(_u10_u1_n2025 ), .A2(_u10_u1_n1846 ), .A3(_u10_u1_n1989 ), .ZN(_u10_u1_n2374 ) );
NAND3_X1 _u10_u1_U303  ( .A1(_u10_u1_n1885 ), .A2(_u10_u1_n2380 ), .A3(_u10_u1_n2381 ), .ZN(_u10_u1_n2375 ) );
OR2_X1 _u10_u1_U302  ( .A1(_u10_u1_n2089 ), .A2(_u10_u1_n2379 ), .ZN(_u10_u1_n2377 ) );
NAND2_X1 _u10_u1_U301  ( .A1(_u10_u1_n2377 ), .A2(_u10_u1_n2378 ), .ZN(_u10_u1_n2376 ) );
NAND3_X1 _u10_u1_U300  ( .A1(_u10_u1_n2374 ), .A2(_u10_u1_n2375 ), .A3(_u10_u1_n2376 ), .ZN(_u10_u1_n2363 ) );
NOR2_X1 _u10_u1_U299  ( .A1(_u10_u1_n2354 ), .A2(_u10_u1_n2373 ), .ZN(_u10_u1_n2372 ) );
NOR2_X1 _u10_u1_U298  ( .A1(_u10_u1_n2372 ), .A2(_u10_u1_n2174 ), .ZN(_u10_u1_n2364 ) );
NOR2_X1 _u10_u1_U297  ( .A1(_u10_u1_n2370 ), .A2(_u10_u1_n2371 ), .ZN(_u10_u1_n2367 ) );
NOR2_X1 _u10_u1_U296  ( .A1(_u10_u1_n2369 ), .A2(_u10_u1_n2353 ), .ZN(_u10_u1_n2368 ) );
NOR2_X1 _u10_u1_U295  ( .A1(_u10_u1_n2367 ), .A2(_u10_u1_n2368 ), .ZN(_u10_u1_n2366 ) );
NOR2_X1 _u10_u1_U294  ( .A1(_u10_u1_n2366 ), .A2(_u10_u1_n2007 ), .ZN(_u10_u1_n2365 ) );
NOR4_X1 _u10_u1_U293  ( .A1(_u10_u1_n2362 ), .A2(_u10_u1_n2363 ), .A3(_u10_u1_n2364 ), .A4(_u10_u1_n2365 ), .ZN(_u10_u1_n2361 ) );
NAND4_X1 _u10_u1_U292  ( .A1(_u10_u1_n2358 ), .A2(_u10_u1_n2359 ), .A3(_u10_u1_n2360 ), .A4(_u10_u1_n2361 ), .ZN(_u10_u1_n2357 ) );
MUX2_X1 _u10_u1_U291  ( .A(_u10_u1_n2357 ), .B(_u10_gnt_p0_d[3] ), .S(_u10_u1_n1809 ), .Z(_u10_u1_n2000 ) );
NOR2_X1 _u10_u1_U290  ( .A1(_u10_u1_n2048 ), .A2(_u10_u1_n1835 ), .ZN(_u10_u1_n2175 ) );
NAND2_X1 _u10_u1_U289  ( .A1(_u10_u1_n2175 ), .A2(_u10_u1_n2356 ), .ZN(_u10_u1_n2355 ) );
NAND2_X1 _u10_u1_U288  ( .A1(_u10_u1_n2354 ), .A2(_u10_u1_n2355 ), .ZN(_u10_u1_n1913 ) );
NOR2_X1 _u10_u1_U287  ( .A1(_u10_u1_n2353 ), .A2(_u10_u1_n1913 ), .ZN(_u10_u1_n2347 ) );
NOR2_X1 _u10_u1_U286  ( .A1(_u10_u1_n2351 ), .A2(_u10_u1_n2352 ), .ZN(_u10_u1_n2348 ) );
NOR2_X1 _u10_u1_U285  ( .A1(_u10_u1_n1825 ), .A2(_u10_u1_n2173 ), .ZN(_u10_u1_n2349 ) );
NOR4_X1 _u10_u1_U284  ( .A1(_u10_u1_n2347 ), .A2(_u10_u1_n2348 ), .A3(_u10_u1_n2349 ), .A4(_u10_u1_n2350 ), .ZN(_u10_u1_n2336 ) );
AND3_X1 _u10_u1_U283  ( .A1(_u10_u1_n2274 ), .A2(_u10_u1_n2346 ), .A3(_u10_u1_n2169 ), .ZN(_u10_u1_n2344 ) );
NAND3_X1 _u10_u1_U282  ( .A1(_u10_u1_n2175 ), .A2(_u10_u1_n1825 ), .A3(_u10_u1_n2345 ), .ZN(_u10_u1_n1937 ) );
INV_X1 _u10_u1_U281  ( .A(_u10_u1_n1937 ), .ZN(_u10_u1_n2132 ) );
NOR2_X1 _u10_u1_U280  ( .A1(_u10_u1_n2344 ), .A2(_u10_u1_n2132 ), .ZN(_u10_u1_n2338 ) );
NOR2_X1 _u10_u1_U279  ( .A1(_u10_u1_n2132 ), .A2(_u10_u1_n2343 ), .ZN(_u10_u1_n2339 ) );
AND2_X1 _u10_u1_U278  ( .A1(_u10_u1_n2342 ), .A2(_u10_u1_n1835 ), .ZN(_u10_u1_n2340 ) );
NOR2_X1 _u10_u1_U277  ( .A1(_u10_u1_n1875 ), .A2(_u10_u1_n1883 ), .ZN(_u10_u1_n1882 ) );
INV_X1 _u10_u1_U276  ( .A(_u10_u1_n1882 ), .ZN(_u10_u1_n1918 ) );
NOR2_X1 _u10_u1_U275  ( .A1(_u10_u1_n2169 ), .A2(_u10_u1_n1918 ), .ZN(_u10_u1_n2341 ) );
NOR4_X1 _u10_u1_U274  ( .A1(_u10_u1_n2338 ), .A2(_u10_u1_n2339 ), .A3(_u10_u1_n2340 ), .A4(_u10_u1_n2341 ), .ZN(_u10_u1_n2337 ) );
AND2_X1 _u10_u1_U273  ( .A1(_u10_u1_n2336 ), .A2(_u10_u1_n2337 ), .ZN(_u10_u1_n2032 ) );
NAND4_X1 _u10_u1_U272  ( .A1(_u10_u1_n2333 ), .A2(_u10_u1_n2334 ), .A3(_u10_u1_n2335 ), .A4(_u10_u1_n2032 ), .ZN(_u10_u1_n2316 ) );
NAND2_X1 _u10_u1_U271  ( .A1(_u10_u1_n2332 ), .A2(_u10_u1_n1837 ), .ZN(_u10_u1_n2324 ) );
NAND2_X1 _u10_u1_U270  ( .A1(_u10_u1_n2227 ), .A2(_u10_u1_n2209 ), .ZN(_u10_u1_n2331 ) );
NAND2_X1 _u10_u1_U269  ( .A1(_u10_u1_n2330 ), .A2(_u10_u1_n2331 ), .ZN(_u10_u1_n2329 ) );
NAND2_X1 _u10_u1_U268  ( .A1(_u10_u1_n1920 ), .A2(_u10_u1_n2329 ), .ZN(_u10_u1_n2325 ) );
NAND2_X1 _u10_u1_U267  ( .A1(_u10_u1_n2327 ), .A2(_u10_u1_n2328 ), .ZN(_u10_u1_n2326 ) );
NAND3_X1 _u10_u1_U266  ( .A1(_u10_u1_n2324 ), .A2(_u10_u1_n2325 ), .A3(_u10_u1_n2326 ), .ZN(_u10_u1_n2317 ) );
AND2_X1 _u10_u1_U265  ( .A1(_u10_u1_n2322 ), .A2(_u10_u1_n2323 ), .ZN(_u10_u1_n2318 ) );
NOR2_X1 _u10_u1_U264  ( .A1(_u10_u1_n2320 ), .A2(_u10_u1_n2321 ), .ZN(_u10_u1_n2319 ) );
NOR4_X1 _u10_u1_U263  ( .A1(_u10_u1_n2316 ), .A2(_u10_u1_n2317 ), .A3(_u10_u1_n2318 ), .A4(_u10_u1_n2319 ), .ZN(_u10_u1_n2160 ) );
NOR2_X1 _u10_u1_U262  ( .A1(_u10_u1_n2314 ), .A2(_u10_u1_n2315 ), .ZN(_u10_u1_n2313 ) );
NOR3_X1 _u10_u1_U261  ( .A1(_u10_u1_n2268 ), .A2(_u10_u1_n2312 ), .A3(_u10_u1_n2313 ), .ZN(_u10_u1_n2311 ) );
NAND3_X1 _u10_u1_U260  ( .A1(_u10_u1_n2309 ), .A2(_u10_u1_n2310 ), .A3(_u10_u1_n2311 ), .ZN(_u10_u1_n2308 ) );
NAND2_X1 _u10_u1_U259  ( .A1(_u10_u1_n2147 ), .A2(_u10_u1_n2308 ), .ZN(_u10_u1_n2302 ) );
NAND2_X1 _u10_u1_U258  ( .A1(_u10_u1_n2276 ), .A2(_u10_u1_n2307 ), .ZN(_u10_u1_n2304 ) );
NAND2_X1 _u10_u1_U257  ( .A1(_u10_u1_n1856 ), .A2(_u10_u1_n2306 ), .ZN(_u10_u1_n2305 ) );
NAND4_X1 _u10_u1_U256  ( .A1(_u10_u1_n2302 ), .A2(_u10_u1_n2303 ), .A3(_u10_u1_n2304 ), .A4(_u10_u1_n2305 ), .ZN(_u10_u1_n2279 ) );
OR3_X1 _u10_u1_U255  ( .A1(_u10_u1_n2089 ), .A2(_u10_u1_n2046 ), .A3(_u10_u1_n2301 ), .ZN(_u10_u1_n2300 ) );
NAND2_X1 _u10_u1_U254  ( .A1(_u10_u1_n2299 ), .A2(_u10_u1_n2300 ), .ZN(_u10_u1_n2288 ) );
NAND3_X1 _u10_u1_U253  ( .A1(_u10_u1_n2296 ), .A2(_u10_u1_n2297 ), .A3(_u10_u1_n2298 ), .ZN(_u10_u1_n2221 ) );
NAND2_X1 _u10_u1_U252  ( .A1(_u10_u1_n2046 ), .A2(_u10_u1_n2221 ), .ZN(_u10_u1_n2289 ) );
NAND2_X1 _u10_u1_U251  ( .A1(_u10_u1_n2295 ), .A2(_u10_u1_n2209 ), .ZN(_u10_u1_n2292 ) );
NAND3_X1 _u10_u1_U250  ( .A1(_u10_u1_n2292 ), .A2(_u10_u1_n2293 ), .A3(_u10_u1_n2294 ), .ZN(_u10_u1_n2291 ) );
NAND2_X1 _u10_u1_U249  ( .A1(_u10_u1_n1964 ), .A2(_u10_u1_n2291 ), .ZN(_u10_u1_n2290 ) );
NAND3_X1 _u10_u1_U248  ( .A1(_u10_u1_n2288 ), .A2(_u10_u1_n2289 ), .A3(_u10_u1_n2290 ), .ZN(_u10_u1_n2280 ) );
NOR4_X1 _u10_u1_U247  ( .A1(_u10_u1_n2285 ), .A2(_u10_u1_n2286 ), .A3(_u10_u1_n2287 ), .A4(_u10_u1_n2216 ), .ZN(_u10_u1_n2283 ) );
NOR2_X1 _u10_u1_U246  ( .A1(_u10_u1_n2283 ), .A2(_u10_u1_n2284 ), .ZN(_u10_u1_n2281 ) );
NOR2_X1 _u10_u1_U245  ( .A1(_u10_u1_n1825 ), .A2(_u10_u1_n2275 ), .ZN(_u10_u1_n2282 ) );
NOR4_X1 _u10_u1_U244  ( .A1(_u10_u1_n2279 ), .A2(_u10_u1_n2280 ), .A3(_u10_u1_n2281 ), .A4(_u10_u1_n2282 ), .ZN(_u10_u1_n2161 ) );
NAND3_X1 _u10_u1_U243  ( .A1(_u10_u1_n2174 ), .A2(_u10_u1_n2277 ), .A3(_u10_u1_n2278 ), .ZN(_u10_u1_n2272 ) );
INV_X1 _u10_u1_U242  ( .A(_u10_u1_n2276 ), .ZN(_u10_u1_n2217 ) );
NAND3_X1 _u10_u1_U241  ( .A1(_u10_u1_n2274 ), .A2(_u10_u1_n2275 ), .A3(_u10_u1_n2217 ), .ZN(_u10_u1_n2273 ) );
NAND2_X1 _u10_u1_U240  ( .A1(_u10_u1_n2272 ), .A2(_u10_u1_n2273 ), .ZN(_u10_u1_n2259 ) );
NAND2_X1 _u10_u1_U239  ( .A1(_u10_u1_n2270 ), .A2(_u10_u1_n2271 ), .ZN(_u10_u1_n2260 ) );
NOR2_X1 _u10_u1_U238  ( .A1(_u10_u1_n2268 ), .A2(_u10_u1_n2269 ), .ZN(_u10_u1_n2232 ) );
NAND3_X1 _u10_u1_U237  ( .A1(_u10_u1_n2232 ), .A2(_u10_u1_n2240 ), .A3(_u10_u1_n2267 ), .ZN(_u10_u1_n2266 ) );
NAND2_X1 _u10_u1_U236  ( .A1(_u10_u1_n1950 ), .A2(_u10_u1_n2266 ), .ZN(_u10_u1_n2261 ) );
NAND3_X1 _u10_u1_U235  ( .A1(_u10_u1_n2265 ), .A2(_u10_u1_n2155 ), .A3(_u10_u1_n2238 ), .ZN(_u10_u1_n2264 ) );
NAND2_X1 _u10_u1_U234  ( .A1(_u10_u1_n2263 ), .A2(_u10_u1_n2264 ), .ZN(_u10_u1_n2262 ) );
NAND4_X1 _u10_u1_U233  ( .A1(_u10_u1_n2259 ), .A2(_u10_u1_n2260 ), .A3(_u10_u1_n2261 ), .A4(_u10_u1_n2262 ), .ZN(_u10_u1_n2241 ) );
OR2_X1 _u10_u1_U232  ( .A1(_u10_u1_n2258 ), .A2(_u10_u1_n10 ), .ZN(_u10_u1_n2251 ) );
NAND2_X1 _u10_u1_U231  ( .A1(_u10_u1_n2256 ), .A2(_u10_u1_n2257 ), .ZN(_u10_u1_n2255 ) );
NAND2_X1 _u10_u1_U230  ( .A1(_u10_u1_n2228 ), .A2(_u10_u1_n2255 ), .ZN(_u10_u1_n2252 ) );
NAND2_X1 _u10_u1_U229  ( .A1(_u10_u1_n2254 ), .A2(_u10_u1_n2209 ), .ZN(_u10_u1_n2253 ) );
NAND3_X1 _u10_u1_U228  ( .A1(_u10_u1_n2251 ), .A2(_u10_u1_n2252 ), .A3(_u10_u1_n2253 ), .ZN(_u10_u1_n2242 ) );
NOR2_X1 _u10_u1_U227  ( .A1(_u10_u1_n2132 ), .A2(_u10_u1_n2250 ), .ZN(_u10_u1_n2243 ) );
NOR3_X1 _u10_u1_U226  ( .A1(_u10_u1_n2247 ), .A2(_u10_u1_n2248 ), .A3(_u10_u1_n2249 ), .ZN(_u10_u1_n2246 ) );
NOR2_X1 _u10_u1_U225  ( .A1(_u10_u1_n2245 ), .A2(_u10_u1_n2246 ), .ZN(_u10_u1_n2244 ) );
NOR4_X1 _u10_u1_U224  ( .A1(_u10_u1_n2241 ), .A2(_u10_u1_n2242 ), .A3(_u10_u1_n2243 ), .A4(_u10_u1_n2244 ), .ZN(_u10_u1_n2162 ) );
NAND4_X1 _u10_u1_U223  ( .A1(_u10_u1_n2238 ), .A2(_u10_u1_n1885 ), .A3(_u10_u1_n2239 ), .A4(_u10_u1_n2240 ), .ZN(_u10_u1_n2237 ) );
NAND2_X1 _u10_u1_U222  ( .A1(_u10_u1_n2236 ), .A2(_u10_u1_n2237 ), .ZN(_u10_u1_n2205 ) );
NOR2_X1 _u10_u1_U221  ( .A1(1'b0), .A2(_u10_u1_n2073 ), .ZN(_u10_u1_n2123 ));
NAND2_X1 _u10_u1_U220  ( .A1(_u10_u1_n2123 ), .A2(_u10_u1_n2074 ), .ZN(_u10_u1_n2235 ) );
NAND2_X1 _u10_u1_U219  ( .A1(_u10_u1_n2234 ), .A2(_u10_u1_n2235 ), .ZN(_u10_u1_n2206 ) );
NAND2_X1 _u10_u1_U218  ( .A1(_u10_u1_n2232 ), .A2(_u10_u1_n2233 ), .ZN(_u10_u1_n2231 ) );
NAND2_X1 _u10_u1_U217  ( .A1(_u10_u1_n2230 ), .A2(_u10_u1_n2231 ), .ZN(_u10_u1_n2207 ) );
NAND2_X1 _u10_u1_U216  ( .A1(1'b0), .A2(_u10_u1_n2229 ), .ZN(_u10_u1_n2211 ));
NAND2_X1 _u10_u1_U215  ( .A1(_u10_u1_n2227 ), .A2(_u10_u1_n2228 ), .ZN(_u10_u1_n2226 ) );
NAND2_X1 _u10_u1_U214  ( .A1(_u10_u1_n2173 ), .A2(_u10_u1_n2226 ), .ZN(_u10_u1_n2224 ) );
NAND2_X1 _u10_u1_U213  ( .A1(_u10_u1_n2224 ), .A2(_u10_u1_n2225 ), .ZN(_u10_u1_n2212 ) );
NAND2_X1 _u10_u1_U212  ( .A1(_u10_u1_n2223 ), .A2(_u10_u1_n2096 ), .ZN(_u10_u1_n2222 ) );
NAND2_X1 _u10_u1_U211  ( .A1(_u10_u1_n2108 ), .A2(_u10_u1_n2222 ), .ZN(_u10_u1_n2213 ) );
INV_X1 _u10_u1_U210  ( .A(_u10_u1_n2221 ), .ZN(_u10_u1_n2218 ) );
NAND4_X1 _u10_u1_U209  ( .A1(_u10_u1_n2217 ), .A2(_u10_u1_n2218 ), .A3(_u10_u1_n2219 ), .A4(_u10_u1_n2220 ), .ZN(_u10_u1_n2215 ) );
NAND2_X1 _u10_u1_U208  ( .A1(_u10_u1_n2215 ), .A2(_u10_u1_n2216 ), .ZN(_u10_u1_n2214 ) );
NAND4_X1 _u10_u1_U207  ( .A1(_u10_u1_n2211 ), .A2(_u10_u1_n2212 ), .A3(_u10_u1_n2213 ), .A4(_u10_u1_n2214 ), .ZN(_u10_u1_n2210 ) );
NAND2_X1 _u10_u1_U206  ( .A1(_u10_u1_n2209 ), .A2(_u10_u1_n2210 ), .ZN(_u10_u1_n2208 ) );
NAND4_X1 _u10_u1_U205  ( .A1(_u10_u1_n2205 ), .A2(_u10_u1_n2206 ), .A3(_u10_u1_n2207 ), .A4(_u10_u1_n2208 ), .ZN(_u10_u1_n2164 ) );
NOR3_X1 _u10_u1_U204  ( .A1(_u10_u1_n2202 ), .A2(_u10_u1_n2203 ), .A3(_u10_u1_n2204 ), .ZN(_u10_u1_n2194 ) );
INV_X1 _u10_u1_U203  ( .A(_u10_u1_n2185 ), .ZN(_u10_u1_n2197 ) );
NAND2_X1 _u10_u1_U202  ( .A1(_u10_u1_n2201 ), .A2(_u10_u1_n2112 ), .ZN(_u10_u1_n2199 ) );
OR2_X1 _u10_u1_U201  ( .A1(_u10_u1_n2198 ), .A2(_u10_u1_n2123 ), .ZN(_u10_u1_n2200 ) );
NAND2_X1 _u10_u1_U200  ( .A1(_u10_u1_n2199 ), .A2(_u10_u1_n2200 ), .ZN(_u10_u1_n2158 ) );
NOR4_X1 _u10_u1_U199  ( .A1(_u10_u1_n2196 ), .A2(_u10_u1_n2197 ), .A3(_u10_u1_n2198 ), .A4(_u10_u1_n2158 ), .ZN(_u10_u1_n2195 ) );
NAND4_X1 _u10_u1_U198  ( .A1(_u10_u1_n2193 ), .A2(_u10_u1_n2190 ), .A3(_u10_u1_n2194 ), .A4(_u10_u1_n2195 ), .ZN(_u10_u1_n2192 ) );
NAND2_X1 _u10_u1_U197  ( .A1(_u10_u1_n1852 ), .A2(_u10_u1_n2192 ), .ZN(_u10_u1_n2176 ) );
AND4_X1 _u10_u1_U196  ( .A1(_u10_u1_n2188 ), .A2(_u10_u1_n2189 ), .A3(_u10_u1_n2190 ), .A4(_u10_u1_n2191 ), .ZN(_u10_u1_n2187 ) );
NAND4_X1 _u10_u1_U195  ( .A1(_u10_u1_n2184 ), .A2(_u10_u1_n2185 ), .A3(_u10_u1_n2186 ), .A4(_u10_u1_n2187 ), .ZN(_u10_u1_n2183 ) );
NAND2_X1 _u10_u1_U194  ( .A1(_u10_u1_n1858 ), .A2(_u10_u1_n2183 ), .ZN(_u10_u1_n2177 ) );
NAND2_X1 _u10_u1_U193  ( .A1(_u10_u1_n2181 ), .A2(_u10_u1_n2182 ), .ZN(_u10_u1_n2179 ) );
NAND2_X1 _u10_u1_U192  ( .A1(_u10_u1_n2179 ), .A2(_u10_u1_n2180 ), .ZN(_u10_u1_n2178 ) );
NAND3_X1 _u10_u1_U191  ( .A1(_u10_u1_n2176 ), .A2(_u10_u1_n2177 ), .A3(_u10_u1_n2178 ), .ZN(_u10_u1_n2165 ) );
AND2_X1 _u10_u1_U190  ( .A1(_u10_u1_n2174 ), .A2(_u10_u1_n2175 ), .ZN(_u10_u1_n2172 ) );
NOR2_X1 _u10_u1_U189  ( .A1(_u10_u1_n2172 ), .A2(_u10_u1_n2173 ), .ZN(_u10_u1_n2166 ) );
NOR2_X1 _u10_u1_U188  ( .A1(_u10_u1_n2170 ), .A2(_u10_u1_n2171 ), .ZN(_u10_u1_n2168 ) );
NOR2_X1 _u10_u1_U187  ( .A1(_u10_u1_n2168 ), .A2(_u10_u1_n2169 ), .ZN(_u10_u1_n2167 ) );
NOR4_X1 _u10_u1_U186  ( .A1(_u10_u1_n2164 ), .A2(_u10_u1_n2165 ), .A3(_u10_u1_n2166 ), .A4(_u10_u1_n2167 ), .ZN(_u10_u1_n2163 ) );
NAND4_X1 _u10_u1_U185  ( .A1(_u10_u1_n2160 ), .A2(_u10_u1_n2161 ), .A3(_u10_u1_n2162 ), .A4(_u10_u1_n2163 ), .ZN(_u10_u1_n2159 ) );
MUX2_X1 _u10_u1_U184  ( .A(_u10_u1_n2159 ), .B(_u10_gnt_p0_d[4] ), .S(_u10_u1_n1809 ), .Z(_u10_u1_n2001 ) );
NAND2_X1 _u10_u1_U183  ( .A1(_u10_u1_n1852 ), .A2(_u10_u1_n2158 ), .ZN(_u10_u1_n2142 ) );
NOR3_X1 _u10_u1_U182  ( .A1(_u10_u1_n2157 ), .A2(_u10_req_p0_0_ ), .A3(_u10_u1_n2043 ), .ZN(_u10_u1_n1884 ) );
NOR2_X1 _u10_u1_U181  ( .A1(1'b0), .A2(_u10_u1_n1884 ), .ZN(_u10_u1_n1947 ));
NAND2_X1 _u10_u1_U180  ( .A1(_u10_u1_n1947 ), .A2(_u10_u1_n2156 ), .ZN(_u10_u1_n2154 ) );
NAND2_X1 _u10_u1_U179  ( .A1(_u10_u1_n2154 ), .A2(_u10_u1_n2155 ), .ZN(_u10_u1_n2149 ) );
NOR2_X1 _u10_u1_U178  ( .A1(_u10_u1_n2046 ), .A2(_u10_u1_n1882 ), .ZN(_u10_u1_n1896 ) );
NAND2_X1 _u10_u1_U177  ( .A1(_u10_u1_n1896 ), .A2(_u10_u1_n2045 ), .ZN(_u10_u1_n2153 ) );
NAND2_X1 _u10_u1_U176  ( .A1(_u10_u1_n2152 ), .A2(_u10_u1_n2153 ), .ZN(_u10_u1_n2150 ) );
NAND3_X1 _u10_u1_U175  ( .A1(_u10_u1_n2149 ), .A2(_u10_u1_n2150 ), .A3(_u10_u1_n2151 ), .ZN(_u10_u1_n2148 ) );
NAND2_X1 _u10_u1_U174  ( .A1(_u10_u1_n2147 ), .A2(_u10_u1_n2148 ), .ZN(_u10_u1_n2143 ) );
NAND2_X1 _u10_u1_U173  ( .A1(_u10_u1_n2145 ), .A2(_u10_u1_n2146 ), .ZN(_u10_u1_n2144 ) );
NAND3_X1 _u10_u1_U172  ( .A1(_u10_u1_n2142 ), .A2(_u10_u1_n2143 ), .A3(_u10_u1_n2144 ), .ZN(_u10_u1_n2091 ) );
NAND2_X1 _u10_u1_U171  ( .A1(_u10_u1_n2141 ), .A2(_u10_u1_n1884 ), .ZN(_u10_u1_n2015 ) );
INV_X1 _u10_u1_U170  ( .A(_u10_u1_n2015 ), .ZN(_u10_u1_n1902 ) );
NAND2_X1 _u10_u1_U169  ( .A1(_u10_u1_n2140 ), .A2(_u10_u1_n1902 ), .ZN(_u10_u1_n2138 ) );
NAND2_X1 _u10_u1_U168  ( .A1(_u10_u1_n2138 ), .A2(_u10_u1_n2139 ), .ZN(_u10_u1_n2137 ) );
NAND2_X1 _u10_u1_U167  ( .A1(_u10_u1_n2136 ), .A2(_u10_u1_n2137 ), .ZN(_u10_u1_n1985 ) );
NOR3_X1 _u10_u1_U166  ( .A1(_u10_u1_n1980 ), .A2(1'b0), .A3(_u10_u1_n1985 ),.ZN(_u10_u1_n2135 ) );
OR3_X1 _u10_u1_U165  ( .A1(_u10_u1_n1828 ), .A2(_u10_u1_n2134 ), .A3(_u10_u1_n2135 ), .ZN(_u10_u1_n2128 ) );
NOR2_X1 _u10_u1_U164  ( .A1(_u10_u1_n2133 ), .A2(_u10_u1_n1882 ), .ZN(_u10_u1_n1867 ) );
AND2_X1 _u10_u1_U163  ( .A1(_u10_u1_n2132 ), .A2(_u10_u1_n1867 ), .ZN(_u10_u1_n2130 ) );
NOR2_X1 _u10_u1_U162  ( .A1(_u10_u1_n2130 ), .A2(_u10_u1_n2131 ), .ZN(_u10_u1_n2129 ) );
NAND2_X1 _u10_u1_U161  ( .A1(_u10_u1_n2009 ), .A2(_u10_u1_n2027 ), .ZN(_u10_u1_n1905 ) );
NOR3_X1 _u10_u1_U160  ( .A1(_u10_u1_n2128 ), .A2(_u10_u1_n2129 ), .A3(_u10_u1_n1905 ), .ZN(_u10_u1_n2126 ) );
NOR2_X1 _u10_u1_U159  ( .A1(_u10_u1_n2126 ), .A2(_u10_u1_n2127 ), .ZN(_u10_u1_n2092 ) );
NAND3_X1 _u10_u1_U158  ( .A1(_u10_u1_n2087 ), .A2(_u10_u1_n1857 ), .A3(1'b0),.ZN(_u10_u1_n2125 ) );
NAND3_X1 _u10_u1_U157  ( .A1(_u10_u1_n2124 ), .A2(_u10_u1_n2072 ), .A3(_u10_u1_n2125 ), .ZN(_u10_u1_n2111 ) );
NAND3_X1 _u10_u1_U156  ( .A1(_u10_u1_n2121 ), .A2(_u10_u1_n2122 ), .A3(_u10_u1_n2123 ), .ZN(_u10_u1_n2098 ) );
NAND3_X1 _u10_u1_U155  ( .A1(_u10_u1_n2119 ), .A2(_u10_u1_n1952 ), .A3(_u10_u1_n2120 ), .ZN(_u10_u1_n2100 ) );
INV_X1 _u10_u1_U154  ( .A(_u10_u1_n2100 ), .ZN(_u10_u1_n2117 ) );
NAND2_X1 _u10_u1_U153  ( .A1(_u10_u1_n1884 ), .A2(_u10_u1_n1885 ), .ZN(_u10_u1_n2118 ) );
NAND2_X1 _u10_u1_U152  ( .A1(_u10_u1_n2117 ), .A2(_u10_u1_n2118 ), .ZN(_u10_u1_n2067 ) );
NOR3_X1 _u10_u1_U151  ( .A1(_u10_u1_n2098 ), .A2(_u10_u1_n2116 ), .A3(_u10_u1_n2067 ), .ZN(_u10_u1_n2115 ) );
NOR2_X1 _u10_u1_U150  ( .A1(1'b0), .A2(_u10_u1_n2115 ), .ZN(_u10_u1_n2113 ));
NOR4_X1 _u10_u1_U149  ( .A1(_u10_u1_n2111 ), .A2(_u10_u1_n2112 ), .A3(_u10_u1_n2113 ), .A4(_u10_u1_n2114 ), .ZN(_u10_u1_n2109 ) );
NOR2_X1 _u10_u1_U148  ( .A1(_u10_u1_n2109 ), .A2(_u10_u1_n2110 ), .ZN(_u10_u1_n2093 ) );
NAND2_X1 _u10_u1_U147  ( .A1(_u10_u1_n1882 ), .A2(_u10_u1_n2108 ), .ZN(_u10_u1_n2107 ) );
NAND2_X1 _u10_u1_U146  ( .A1(_u10_u1_n2106 ), .A2(_u10_u1_n2107 ), .ZN(_u10_u1_n1962 ) );
NAND2_X1 _u10_u1_U145  ( .A1(_u10_u1_n2105 ), .A2(_u10_u1_n1962 ), .ZN(_u10_u1_n2101 ) );
NAND3_X1 _u10_u1_U144  ( .A1(_u10_u1_n2104 ), .A2(_u10_u1_n1963 ), .A3(_u10_u1_n1884 ), .ZN(_u10_u1_n2102 ) );
NAND2_X1 _u10_u1_U143  ( .A1(_u10_u1_n1961 ), .A2(_u10_u1_n1955 ), .ZN(_u10_u1_n2103 ) );
NAND3_X1 _u10_u1_U142  ( .A1(_u10_u1_n2101 ), .A2(_u10_u1_n2102 ), .A3(_u10_u1_n2103 ), .ZN(_u10_u1_n2097 ) );
NOR4_X1 _u10_u1_U141  ( .A1(_u10_u1_n2097 ), .A2(_u10_u1_n2098 ), .A3(_u10_u1_n2099 ), .A4(_u10_u1_n2100 ), .ZN(_u10_u1_n2095 ) );
NOR2_X1 _u10_u1_U140  ( .A1(_u10_u1_n2095 ), .A2(_u10_u1_n2096 ), .ZN(_u10_u1_n2094 ) );
NOR4_X1 _u10_u1_U139  ( .A1(_u10_u1_n2091 ), .A2(_u10_u1_n2092 ), .A3(_u10_u1_n2093 ), .A4(_u10_u1_n2094 ), .ZN(_u10_u1_n1810 ) );
NAND2_X1 _u10_u1_U138  ( .A1(_u10_u1_n1882 ), .A2(_u10_u1_n2090 ), .ZN(_u10_u1_n2075 ) );
NAND2_X1 _u10_u1_U137  ( .A1(_u10_u1_n2088 ), .A2(_u10_u1_n2089 ), .ZN(_u10_u1_n2076 ) );
NAND2_X1 _u10_u1_U136  ( .A1(_u10_u1_n2086 ), .A2(_u10_u1_n2087 ), .ZN(_u10_u1_n2082 ) );
NAND2_X1 _u10_u1_U135  ( .A1(_u10_u1_n1886 ), .A2(_u10_u1_n2067 ), .ZN(_u10_u1_n2085 ) );
NAND3_X1 _u10_u1_U134  ( .A1(_u10_u1_n1878 ), .A2(_u10_u1_n1875 ), .A3(_u10_u1_n2085 ), .ZN(_u10_u1_n2084 ) );
NAND2_X1 _u10_u1_U133  ( .A1(_u10_u1_n2084 ), .A2(_u10_u1_n1857 ), .ZN(_u10_u1_n2083 ) );
NAND4_X1 _u10_u1_U132  ( .A1(_u10_u1_n2080 ), .A2(_u10_u1_n2081 ), .A3(_u10_u1_n2082 ), .A4(_u10_u1_n2083 ), .ZN(_u10_u1_n2079 ) );
NAND2_X1 _u10_u1_U131  ( .A1(_u10_u1_n2078 ), .A2(_u10_u1_n2079 ), .ZN(_u10_u1_n2077 ) );
NAND3_X1 _u10_u1_U130  ( .A1(_u10_u1_n2075 ), .A2(_u10_u1_n2076 ), .A3(_u10_u1_n2077 ), .ZN(_u10_u1_n2051 ) );
NAND2_X1 _u10_u1_U129  ( .A1(_u10_u1_n2073 ), .A2(_u10_u1_n2074 ), .ZN(_u10_u1_n2069 ) );
NAND3_X1 _u10_u1_U128  ( .A1(1'b0), .A2(_u10_u1_n1857 ), .A3(_u10_u1_n1856 ),.ZN(_u10_u1_n2070 ) );
NAND4_X1 _u10_u1_U127  ( .A1(_u10_u1_n2069 ), .A2(_u10_u1_n2070 ), .A3(_u10_u1_n2071 ), .A4(_u10_u1_n2072 ), .ZN(_u10_u1_n2060 ) );
NAND2_X1 _u10_u1_U126  ( .A1(_u10_u1_n2067 ), .A2(_u10_u1_n2068 ), .ZN(_u10_u1_n2066 ) );
AND2_X1 _u10_u1_U125  ( .A1(_u10_u1_n2065 ), .A2(_u10_u1_n2066 ), .ZN(_u10_u1_n1854 ) );
NAND2_X1 _u10_u1_U124  ( .A1(_u10_u1_n1854 ), .A2(_u10_u1_n2064 ), .ZN(_u10_u1_n1859 ) );
NOR2_X1 _u10_u1_U123  ( .A1(1'b0), .A2(_u10_u1_n2063 ), .ZN(_u10_u1_n2062 ));
NOR4_X1 _u10_u1_U122  ( .A1(_u10_u1_n2060 ), .A2(_u10_u1_n1859 ), .A3(_u10_u1_n2061 ), .A4(_u10_u1_n2062 ), .ZN(_u10_u1_n2058 ) );
NOR2_X1 _u10_u1_U121  ( .A1(_u10_u1_n2058 ), .A2(_u10_u1_n2059 ), .ZN(_u10_u1_n2052 ) );
NOR2_X1 _u10_u1_U120  ( .A1(_u10_u1_n2056 ), .A2(_u10_u1_n2057 ), .ZN(_u10_u1_n2053 ) );
NOR2_X1 _u10_u1_U119  ( .A1(_u10_u1_n2055 ), .A2(_u10_u1_n1985 ), .ZN(_u10_u1_n2054 ) );
NOR4_X1 _u10_u1_U118  ( .A1(_u10_u1_n2051 ), .A2(_u10_u1_n2052 ), .A3(_u10_u1_n2053 ), .A4(_u10_u1_n2054 ), .ZN(_u10_u1_n1811 ) );
OR2_X1 _u10_u1_U117  ( .A1(_u10_u1_n2019 ), .A2(_u10_u1_n2050 ), .ZN(_u10_u1_n2035 ) );
NAND2_X1 _u10_u1_U116  ( .A1(_u10_u1_n2048 ), .A2(_u10_u1_n2049 ), .ZN(_u10_u1_n2036 ) );
NAND2_X1 _u10_u1_U115  ( .A1(_u10_u1_n2046 ), .A2(_u10_u1_n2047 ), .ZN(_u10_u1_n2037 ) );
NOR2_X1 _u10_u1_U114  ( .A1(_u10_u1_n2044 ), .A2(_u10_u1_n2045 ), .ZN(_u10_u1_n2040 ) );
NOR2_X1 _u10_u1_U113  ( .A1(_u10_u1_n2042 ), .A2(_u10_u1_n2043 ), .ZN(_u10_u1_n2041 ) );
NOR3_X1 _u10_u1_U112  ( .A1(_u10_u1_n2039 ), .A2(_u10_u1_n2040 ), .A3(_u10_u1_n2041 ), .ZN(_u10_u1_n2038 ) );
NAND4_X1 _u10_u1_U111  ( .A1(_u10_u1_n2035 ), .A2(_u10_u1_n2036 ), .A3(_u10_u1_n2037 ), .A4(_u10_u1_n2038 ), .ZN(_u10_u1_n2028 ) );
NAND3_X1 _u10_u1_U110  ( .A1(_u10_u1_n2032 ), .A2(_u10_u1_n2033 ), .A3(_u10_u1_n2034 ), .ZN(_u10_u1_n2029 ) );
NOR4_X1 _u10_u1_U109  ( .A1(_u10_u1_n2028 ), .A2(_u10_u1_n2029 ), .A3(_u10_u1_n2030 ), .A4(_u10_u1_n2031 ), .ZN(_u10_u1_n1812 ) );
INV_X1 _u10_u1_U108  ( .A(_u10_u1_n2027 ), .ZN(_u10_u1_n2026 ) );
NAND3_X1 _u10_u1_U107  ( .A1(_u10_u1_n2024 ), .A2(_u10_u1_n2025 ), .A3(_u10_u1_n2026 ), .ZN(_u10_u1_n1968 ) );
NAND2_X1 _u10_u1_U106  ( .A1(_u10_u1_n1902 ), .A2(_u10_u1_n2023 ), .ZN(_u10_u1_n2021 ) );
NAND2_X1 _u10_u1_U105  ( .A1(_u10_u1_n2021 ), .A2(_u10_u1_n2022 ), .ZN(_u10_u1_n2016 ) );
NAND2_X1 _u10_u1_U104  ( .A1(_u10_u1_n2019 ), .A2(_u10_u1_n2020 ), .ZN(_u10_u1_n2018 ) );
NAND3_X1 _u10_u1_U103  ( .A1(_u10_u1_n2016 ), .A2(_u10_u1_n2017 ), .A3(_u10_u1_n2018 ), .ZN(_u10_u1_n1969 ) );
NAND3_X1 _u10_u1_U102  ( .A1(_u10_u1_n2013 ), .A2(_u10_u1_n2014 ), .A3(_u10_u1_n2015 ), .ZN(_u10_u1_n2011 ) );
NAND3_X1 _u10_u1_U101  ( .A1(_u10_u1_n2011 ), .A2(_u10_u1_n1844 ), .A3(_u10_u1_n2012 ), .ZN(_u10_u1_n1970 ) );
NOR2_X1 _u10_u1_U100  ( .A1(_u10_u1_n2010 ), .A2(_u10_u1_n1918 ), .ZN(_u10_u1_n1995 ) );
INV_X1 _u10_u1_U99  ( .A(_u10_u1_n2009 ), .ZN(_u10_u1_n1990 ) );
NAND2_X1 _u10_u1_U98  ( .A1(_u10_u1_n1990 ), .A2(_u10_u1_n2008 ), .ZN(_u10_u1_n2003 ) );
OR2_X1 _u10_u1_U97  ( .A1(_u10_u1_n2006 ), .A2(_u10_u1_n2007 ), .ZN(_u10_u1_n2004 ) );
NAND2_X1 _u10_u1_U96  ( .A1(1'b0), .A2(_u10_u1_n1845 ), .ZN(_u10_u1_n2005 ));
NAND3_X1 _u10_u1_U95  ( .A1(_u10_u1_n2003 ), .A2(_u10_u1_n2004 ), .A3(_u10_u1_n2005 ), .ZN(_u10_u1_n1917 ) );
NOR2_X1 _u10_u1_U94  ( .A1(_u10_u1_n1897 ), .A2(_u10_u1_n1917 ), .ZN(_u10_u1_n1997 ) );
NOR2_X1 _u10_u1_U93  ( .A1(1'b0), .A2(_u10_u1_n1997 ), .ZN(_u10_u1_n1996 ));
NOR3_X1 _u10_u1_U92  ( .A1(_u10_u1_n1995 ), .A2(1'b0), .A3(_u10_u1_n1996 ),.ZN(_u10_u1_n1991 ) );
NOR2_X1 _u10_u1_U91  ( .A1(1'b0), .A2(_u10_u1_n1994 ), .ZN(_u10_u1_n1993 ));
NOR2_X1 _u10_u1_U90  ( .A1(_u10_u1_n1993 ), .A2(_u10_u1_n1920 ), .ZN(_u10_u1_n1992 ) );
NOR2_X1 _u10_u1_U89  ( .A1(_u10_u1_n1991 ), .A2(_u10_u1_n1992 ), .ZN(_u10_u1_n1972 ) );
NOR3_X1 _u10_u1_U88  ( .A1(_u10_u1_n1989 ), .A2(1'b0), .A3(_u10_u1_n1990 ),.ZN(_u10_u1_n1986 ) );
NOR2_X1 _u10_u1_U87  ( .A1(_u10_u1_n1987 ), .A2(_u10_u1_n1988 ), .ZN(_u10_u1_n1932 ) );
NOR3_X1 _u10_u1_U86  ( .A1(_u10_u1_n1986 ), .A2(1'b0), .A3(_u10_u1_n1932 ),.ZN(_u10_u1_n1973 ) );
INV_X1 _u10_u1_U85  ( .A(_u10_u1_n1985 ), .ZN(_u10_u1_n1982 ) );
NOR4_X1 _u10_u1_U84  ( .A1(1'b0), .A2(_u10_u1_n1982 ), .A3(_u10_u1_n1983 ),.A4(_u10_u1_n1984 ), .ZN(_u10_u1_n1981 ) );
NOR2_X1 _u10_u1_U83  ( .A1(1'b0), .A2(_u10_u1_n1981 ), .ZN(_u10_u1_n1977 ));
NOR2_X1 _u10_u1_U82  ( .A1(_u10_u1_n1979 ), .A2(_u10_u1_n1980 ), .ZN(_u10_u1_n1978 ) );
NOR2_X1 _u10_u1_U81  ( .A1(_u10_u1_n1977 ), .A2(_u10_u1_n1978 ), .ZN(_u10_u1_n1976 ) );
NOR2_X1 _u10_u1_U80  ( .A1(_u10_u1_n1975 ), .A2(_u10_u1_n1976 ), .ZN(_u10_u1_n1974 ) );
NOR3_X1 _u10_u1_U79  ( .A1(_u10_u1_n1972 ), .A2(_u10_u1_n1973 ), .A3(_u10_u1_n1974 ), .ZN(_u10_u1_n1971 ) );
NAND4_X1 _u10_u1_U78  ( .A1(_u10_u1_n1968 ), .A2(_u10_u1_n1969 ), .A3(_u10_u1_n1970 ), .A4(_u10_u1_n1971 ), .ZN(_u10_u1_n1814 ) );
NAND2_X1 _u10_u1_U77  ( .A1(_u10_u1_n1966 ), .A2(_u10_u1_n1967 ), .ZN(_u10_u1_n1965 ) );
NAND2_X1 _u10_u1_U76  ( .A1(_u10_u1_n1964 ), .A2(_u10_u1_n1965 ), .ZN(_u10_u1_n1921 ) );
NAND2_X1 _u10_u1_U75  ( .A1(_u10_u1_n1884 ), .A2(_u10_u1_n1963 ), .ZN(_u10_u1_n1957 ) );
INV_X1 _u10_u1_U74  ( .A(_u10_u1_n1962 ), .ZN(_u10_u1_n1958 ) );
NOR3_X1 _u10_u1_U73  ( .A1(_u10_u1_n1942 ), .A2(_u10_u1_n1960 ), .A3(_u10_u1_n1961 ), .ZN(_u10_u1_n1959 ) );
NAND4_X1 _u10_u1_U72  ( .A1(_u10_u1_n1956 ), .A2(_u10_u1_n1957 ), .A3(_u10_u1_n1958 ), .A4(_u10_u1_n1959 ), .ZN(_u10_u1_n1954 ) );
NAND2_X1 _u10_u1_U71  ( .A1(_u10_u1_n1954 ), .A2(_u10_u1_n1955 ), .ZN(_u10_u1_n1953 ) );
NAND2_X1 _u10_u1_U70  ( .A1(_u10_u1_n1952 ), .A2(_u10_u1_n1953 ), .ZN(_u10_u1_n1951 ) );
NAND2_X1 _u10_u1_U69  ( .A1(_u10_u1_n1950 ), .A2(_u10_u1_n1951 ), .ZN(_u10_u1_n1922 ) );
NAND2_X1 _u10_u1_U68  ( .A1(_u10_u1_n1875 ), .A2(_u10_u1_n1949 ), .ZN(_u10_u1_n1948 ) );
NAND2_X1 _u10_u1_U67  ( .A1(_u10_u1_n1858 ), .A2(_u10_u1_n1948 ), .ZN(_u10_u1_n1923 ) );
NOR2_X1 _u10_u1_U66  ( .A1(1'b0), .A2(_u10_u1_n1947 ), .ZN(_u10_u1_n1943 ));
NOR2_X1 _u10_u1_U65  ( .A1(_u10_u1_n1945 ), .A2(_u10_u1_n1946 ), .ZN(_u10_u1_n1944 ) );
NOR4_X1 _u10_u1_U64  ( .A1(_u10_u1_n1941 ), .A2(_u10_u1_n1942 ), .A3(_u10_u1_n1943 ), .A4(_u10_u1_n1944 ), .ZN(_u10_u1_n1939 ) );
NOR2_X1 _u10_u1_U63  ( .A1(_u10_u1_n1939 ), .A2(_u10_u1_n1940 ), .ZN(_u10_u1_n1925 ) );
NOR2_X1 _u10_u1_U62  ( .A1(_u10_req_p0_0_ ), .A2(_u10_u1_n1938 ), .ZN(_u10_u1_n1936 ) );
NOR2_X1 _u10_u1_U61  ( .A1(_u10_u1_n1936 ), .A2(_u10_u1_n1937 ), .ZN(_u10_u1_n1934 ) );
NOR2_X1 _u10_u1_U60  ( .A1(_u10_u1_n1934 ), .A2(_u10_u1_n1935 ), .ZN(_u10_u1_n1926 ) );
NOR2_X1 _u10_u1_U59  ( .A1(_u10_u1_n1932 ), .A2(_u10_u1_n1933 ), .ZN(_u10_u1_n1930 ) );
NOR2_X1 _u10_u1_U58  ( .A1(_u10_u1_n1930 ), .A2(_u10_u1_n1931 ), .ZN(_u10_u1_n1928 ) );
NOR2_X1 _u10_u1_U57  ( .A1(_u10_u1_n1928 ), .A2(_u10_u1_n1929 ), .ZN(_u10_u1_n1927 ) );
NOR3_X1 _u10_u1_U56  ( .A1(_u10_u1_n1925 ), .A2(_u10_u1_n1926 ), .A3(_u10_u1_n1927 ), .ZN(_u10_u1_n1924 ) );
NAND4_X1 _u10_u1_U55  ( .A1(_u10_u1_n1921 ), .A2(_u10_u1_n1922 ), .A3(_u10_u1_n1923 ), .A4(_u10_u1_n1924 ), .ZN(_u10_u1_n1815 ) );
NAND2_X1 _u10_u1_U54  ( .A1(_u10_u1_n1916 ), .A2(_u10_u1_n1920 ), .ZN(_u10_u1_n1908 ) );
NOR2_X1 _u10_u1_U53  ( .A1(_u10_u1_n1918 ), .A2(_u10_u1_n1919 ), .ZN(_u10_u1_n1915 ) );
NOR3_X1 _u10_u1_U52  ( .A1(_u10_u1_n1915 ), .A2(_u10_u1_n1916 ), .A3(_u10_u1_n1917 ), .ZN(_u10_u1_n1839 ) );
NAND4_X1 _u10_u1_U51  ( .A1(_u10_u1_n1839 ), .A2(_u10_u1_n1912 ), .A3(_u10_u1_n1913 ), .A4(_u10_u1_n1914 ), .ZN(_u10_u1_n1911 ) );
NAND2_X1 _u10_u1_U50  ( .A1(_u10_u1_n1910 ), .A2(_u10_u1_n1911 ), .ZN(_u10_u1_n1909 ) );
NAND2_X1 _u10_u1_U49  ( .A1(_u10_u1_n1908 ), .A2(_u10_u1_n1909 ), .ZN(_u10_u1_n1906 ) );
NAND2_X1 _u10_u1_U48  ( .A1(_u10_u1_n1906 ), .A2(_u10_u1_n1907 ), .ZN(_u10_u1_n1860 ) );
INV_X1 _u10_u1_U47  ( .A(_u10_u1_n1905 ), .ZN(_u10_u1_n1900 ) );
NAND3_X1 _u10_u1_U46  ( .A1(_u10_u1_n1902 ), .A2(_u10_u1_n1903 ), .A3(_u10_u1_n1904 ), .ZN(_u10_u1_n1901 ) );
NAND2_X1 _u10_u1_U45  ( .A1(_u10_u1_n1900 ), .A2(_u10_u1_n1901 ), .ZN(_u10_u1_n1899 ) );
NAND2_X1 _u10_u1_U44  ( .A1(_u10_u1_n1898 ), .A2(_u10_u1_n1899 ), .ZN(_u10_u1_n1861 ) );
NAND2_X1 _u10_u1_U43  ( .A1(_u10_u1_n1897 ), .A2(_u10_u1_n1894 ), .ZN(_u10_u1_n1889 ) );
OR2_X1 _u10_u1_U42  ( .A1(_u10_u1_n1895 ), .A2(_u10_u1_n1896 ), .ZN(_u10_u1_n1890 ) );
NAND3_X1 _u10_u1_U41  ( .A1(_u10_u1_n1894 ), .A2(_u10_u1_n1845 ), .A3(1'b0),.ZN(_u10_u1_n1893 ) );
AND3_X1 _u10_u1_U40  ( .A1(_u10_u1_n1891 ), .A2(_u10_u1_n1892 ), .A3(_u10_u1_n1893 ), .ZN(_u10_u1_n1834 ) );
NAND3_X1 _u10_u1_U39  ( .A1(_u10_u1_n1889 ), .A2(_u10_u1_n1890 ), .A3(_u10_u1_n1834 ), .ZN(_u10_u1_n1888 ) );
NAND2_X1 _u10_u1_U38  ( .A1(_u10_u1_n1887 ), .A2(_u10_u1_n1888 ), .ZN(_u10_u1_n1862 ) );
NAND3_X1 _u10_u1_U37  ( .A1(_u10_u1_n1884 ), .A2(_u10_u1_n1885 ), .A3(_u10_u1_n1886 ), .ZN(_u10_u1_n1874 ) );
NOR2_X1 _u10_u1_U36  ( .A1(_u10_u1_n1883 ), .A2(_u10_u1_n1874 ), .ZN(_u10_u1_n1881 ) );
NOR3_X1 _u10_u1_U35  ( .A1(_u10_u1_n1881 ), .A2(1'b0), .A3(_u10_u1_n1882 ),.ZN(_u10_u1_n1880 ) );
NOR2_X1 _u10_u1_U34  ( .A1(_u10_u1_n1879 ), .A2(_u10_u1_n1880 ), .ZN(_u10_u1_n1864 ) );
NOR2_X1 _u10_u1_U33  ( .A1(_u10_u1_n1877 ), .A2(_u10_u1_n1878 ), .ZN(_u10_u1_n1870 ) );
INV_X1 _u10_u1_U32  ( .A(_u10_u1_n1876 ), .ZN(_u10_u1_n1872 ) );
AND2_X1 _u10_u1_U31  ( .A1(_u10_u1_n1874 ), .A2(_u10_u1_n1875 ), .ZN(_u10_u1_n1873 ) );
NOR2_X1 _u10_u1_U30  ( .A1(_u10_u1_n1872 ), .A2(_u10_u1_n1873 ), .ZN(_u10_u1_n1871 ) );
NOR2_X1 _u10_u1_U29  ( .A1(_u10_u1_n1870 ), .A2(_u10_u1_n1871 ), .ZN(_u10_u1_n1869 ) );
NOR2_X1 _u10_u1_U28  ( .A1(1'b0), .A2(_u10_u1_n1869 ), .ZN(_u10_u1_n1865 ));
NOR2_X1 _u10_u1_U27  ( .A1(_u10_u1_n1867 ), .A2(_u10_u1_n1868 ), .ZN(_u10_u1_n1866 ) );
NOR3_X1 _u10_u1_U26  ( .A1(_u10_u1_n1864 ), .A2(_u10_u1_n1865 ), .A3(_u10_u1_n1866 ), .ZN(_u10_u1_n1863 ) );
NAND4_X1 _u10_u1_U25  ( .A1(_u10_u1_n1860 ), .A2(_u10_u1_n1861 ), .A3(_u10_u1_n1862 ), .A4(_u10_u1_n1863 ), .ZN(_u10_u1_n1816 ) );
NAND2_X1 _u10_u1_U24  ( .A1(_u10_u1_n1858 ), .A2(_u10_u1_n1859 ), .ZN(_u10_u1_n1850 ) );
NAND2_X1 _u10_u1_U23  ( .A1(_u10_u1_n1856 ), .A2(_u10_u1_n1857 ), .ZN(_u10_u1_n1855 ) );
NAND2_X1 _u10_u1_U22  ( .A1(_u10_u1_n1854 ), .A2(_u10_u1_n1855 ), .ZN(_u10_u1_n1853 ) );
NAND2_X1 _u10_u1_U21  ( .A1(_u10_u1_n1852 ), .A2(_u10_u1_n1853 ), .ZN(_u10_u1_n1851 ) );
NAND2_X1 _u10_u1_U20  ( .A1(_u10_u1_n1850 ), .A2(_u10_u1_n1851 ), .ZN(_u10_u1_n1848 ) );
NAND2_X1 _u10_u1_U19  ( .A1(_u10_u1_n1848 ), .A2(_u10_u1_n1849 ), .ZN(_u10_u1_n1818 ) );
OR2_X1 _u10_u1_U18  ( .A1(_u10_u1_n1847 ), .A2(_u10_u1_n15 ), .ZN(_u10_u1_n1840 ) );
NAND3_X1 _u10_u1_U17  ( .A1(_u10_u1_n1845 ), .A2(_u10_u1_n1846 ), .A3(1'b0),.ZN(_u10_u1_n1841 ) );
NAND3_X1 _u10_u1_U16  ( .A1(_u10_u1_n1843 ), .A2(_u10_u1_n1844 ), .A3(1'b0),.ZN(_u10_u1_n1842 ) );
NAND4_X1 _u10_u1_U15  ( .A1(_u10_u1_n1839 ), .A2(_u10_u1_n1840 ), .A3(_u10_u1_n1841 ), .A4(_u10_u1_n1842 ), .ZN(_u10_u1_n1838 ) );
NAND2_X1 _u10_u1_U14  ( .A1(_u10_u1_n1837 ), .A2(_u10_u1_n1838 ), .ZN(_u10_u1_n1819 ) );
NAND2_X1 _u10_u1_U13  ( .A1(_u10_u1_n1835 ), .A2(_u10_u1_n1836 ), .ZN(_u10_u1_n1820 ) );
NOR2_X1 _u10_u1_U12  ( .A1(1'b0), .A2(_u10_u1_n1834 ), .ZN(_u10_u1_n1832 ));
NOR4_X1 _u10_u1_U11  ( .A1(1'b0), .A2(_u10_u1_n1831 ), .A3(_u10_u1_n1832 ),.A4(_u10_u1_n1833 ), .ZN(_u10_u1_n1829 ) );
NOR2_X1 _u10_u1_U10  ( .A1(_u10_u1_n1829 ), .A2(_u10_u1_n1830 ), .ZN(_u10_u1_n1822 ) );
AND2_X1 _u10_u1_U9  ( .A1(_u10_u1_n1827 ), .A2(_u10_u1_n1828 ), .ZN(_u10_u1_n1823 ) );
NOR2_X1 _u10_u1_U8  ( .A1(_u10_u1_n1825 ), .A2(_u10_u1_n1826 ), .ZN(_u10_u1_n1824 ) );
NOR3_X1 _u10_u1_U7  ( .A1(_u10_u1_n1822 ), .A2(_u10_u1_n1823 ), .A3(_u10_u1_n1824 ), .ZN(_u10_u1_n1821 ) );
NAND4_X1 _u10_u1_U6  ( .A1(_u10_u1_n1818 ), .A2(_u10_u1_n1819 ), .A3(_u10_u1_n1820 ), .A4(_u10_u1_n1821 ), .ZN(_u10_u1_n1817 ) );
NOR4_X1 _u10_u1_U5  ( .A1(_u10_u1_n1814 ), .A2(_u10_u1_n1815 ), .A3(_u10_u1_n1816 ), .A4(_u10_u1_n1817 ), .ZN(_u10_u1_n1813 ) );
NAND4_X1 _u10_u1_U4  ( .A1(_u10_u1_n1810 ), .A2(_u10_u1_n1811 ), .A3(_u10_u1_n1812 ), .A4(_u10_u1_n1813 ), .ZN(_u10_u1_n1808 ) );
MUX2_X1 _u10_u1_U3  ( .A(_u10_u1_n1808 ), .B(_u10_gnt_p0_d[0] ), .S(_u10_u1_n1809 ), .Z(_u10_u1_n2002 ) );
DFFR_X1 _u10_u1_state_reg_1_  ( .D(_u10_u1_n1998 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_gnt_p0_d[1] ), .QN(_u10_u1_n14 ) );
DFFR_X1 _u10_u1_state_reg_2_  ( .D(_u10_u1_n1999 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_gnt_p0_d[2] ), .QN(_u10_u1_n13 ) );
DFFR_X1 _u10_u1_state_reg_3_  ( .D(_u10_u1_n2000 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_gnt_p0_d[3] ), .QN(_u10_u1_n12 ) );
DFFR_X1 _u10_u1_state_reg_4_  ( .D(_u10_u1_n2001 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_gnt_p0_d[4] ), .QN(_u10_u1_n10 ) );
DFFR_X1 _u10_u1_state_reg_0_  ( .D(_u10_u1_n2002 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_gnt_p0_d[0] ), .QN(_u10_u1_n15 ) );
NOR2_X1 _u10_u20_U1606  ( .A1(_u10_SYNOPSYS_UNCONNECTED_6 ), .A2(_u10_u20_n1814 ), .ZN(_u10_u20_n3174 ) );
NOR3_X1 _u10_u20_U1605  ( .A1(_u10_SYNOPSYS_UNCONNECTED_5 ), .A2(_u10_u20_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_8 ), .ZN(_u10_u20_n3328 ) );
NAND2_X1 _u10_u20_U1604  ( .A1(_u10_u20_n3174 ), .A2(_u10_u20_n3328 ), .ZN(_u10_u20_n1843 ) );
INV_X1 _u10_u20_U1603  ( .A(_u10_u20_n1843 ), .ZN(_u10_u20_n2461 ) );
INV_X1 _u10_u20_U1602  ( .A(1'b0), .ZN(_u10_u20_n2466 ) );
INV_X1 _u10_u20_U1601  ( .A(1'b0), .ZN(_u10_u20_n2305 ) );
NAND2_X1 _u10_u20_U1600  ( .A1(_u10_u20_n2466 ), .A2(_u10_u20_n2305 ), .ZN(_u10_u20_n1954 ) );
INV_X1 _u10_u20_U1599  ( .A(_u10_u20_n1954 ), .ZN(_u10_u20_n2467 ) );
INV_X1 _u10_u20_U1598  ( .A(1'b0), .ZN(_u10_u20_n1936 ) );
NOR2_X1 _u10_u20_U1597  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u20_n2223 ) );
INV_X1 _u10_u20_U1596  ( .A(1'b0), .ZN(_u10_u20_n1922 ) );
NAND2_X1 _u10_u20_U1595  ( .A1(_u10_u20_n2223 ), .A2(_u10_u20_n1922 ), .ZN(_u10_u20_n2200 ) );
NOR2_X1 _u10_u20_U1594  ( .A1(_u10_u20_n2200 ), .A2(1'b0), .ZN(_u10_u20_n2502 ) );
INV_X1 _u10_u20_U1593  ( .A(_u10_req_p1_0_ ), .ZN(_u10_u20_n2978 ) );
INV_X1 _u10_u20_U1592  ( .A(1'b0), .ZN(_u10_u20_n3000 ) );
NAND2_X1 _u10_u20_U1591  ( .A1(_u10_u20_n2978 ), .A2(_u10_u20_n3000 ), .ZN(_u10_u20_n3356 ) );
INV_X1 _u10_u20_U1590  ( .A(1'b0), .ZN(_u10_u20_n2405 ) );
INV_X1 _u10_u20_U1589  ( .A(1'b0), .ZN(_u10_u20_n2972 ) );
NAND2_X1 _u10_u20_U1588  ( .A1(_u10_u20_n2405 ), .A2(_u10_u20_n2972 ), .ZN(_u10_u20_n2008 ) );
NOR2_X1 _u10_u20_U1587  ( .A1(_u10_u20_n3356 ), .A2(_u10_u20_n2008 ), .ZN(_u10_u20_n2195 ) );
NAND2_X1 _u10_u20_U1586  ( .A1(_u10_u20_n2502 ), .A2(_u10_u20_n2195 ), .ZN(_u10_u20_n2490 ) );
INV_X1 _u10_u20_U1585  ( .A(1'b0), .ZN(_u10_u20_n3040 ) );
INV_X1 _u10_u20_U1584  ( .A(1'b0), .ZN(_u10_u20_n3006 ) );
NAND2_X1 _u10_u20_U1583  ( .A1(_u10_u20_n3040 ), .A2(_u10_u20_n3006 ), .ZN(_u10_u20_n2508 ) );
NOR2_X1 _u10_u20_U1582  ( .A1(_u10_u20_n2508 ), .A2(1'b0), .ZN(_u10_u20_n2493 ) );
INV_X1 _u10_u20_U1581  ( .A(1'b0), .ZN(_u10_u20_n2038 ) );
NAND2_X1 _u10_u20_U1580  ( .A1(_u10_u20_n2493 ), .A2(_u10_u20_n2038 ), .ZN(_u10_u20_n2174 ) );
NOR2_X1 _u10_u20_U1579  ( .A1(_u10_u20_n2490 ), .A2(_u10_u20_n2174 ), .ZN(_u10_u20_n2659 ) );
INV_X1 _u10_u20_U1578  ( .A(1'b0), .ZN(_u10_u20_n2175 ) );
NAND3_X1 _u10_u20_U1577  ( .A1(_u10_u20_n2659 ), .A2(_u10_u20_n2175 ), .A3(1'b0), .ZN(_u10_u20_n3189 ) );
NOR2_X1 _u10_u20_U1576  ( .A1(_u10_u20_n3189 ), .A2(1'b0), .ZN(_u10_u20_n2528 ) );
INV_X1 _u10_u20_U1575  ( .A(1'b0), .ZN(_u10_u20_n2837 ) );
NAND2_X1 _u10_u20_U1574  ( .A1(_u10_u20_n2528 ), .A2(_u10_u20_n2837 ), .ZN(_u10_u20_n2567 ) );
INV_X1 _u10_u20_U1573  ( .A(1'b0), .ZN(_u10_u20_n2080 ) );
INV_X1 _u10_u20_U1572  ( .A(1'b0), .ZN(_u10_u20_n2166 ) );
NAND2_X1 _u10_u20_U1571  ( .A1(_u10_u20_n2080 ), .A2(_u10_u20_n2166 ), .ZN(_u10_u20_n2840 ) );
NOR2_X1 _u10_u20_U1570  ( .A1(_u10_u20_n2567 ), .A2(_u10_u20_n2840 ), .ZN(_u10_u20_n2443 ) );
INV_X1 _u10_u20_U1569  ( .A(1'b0), .ZN(_u10_u20_n2600 ) );
INV_X1 _u10_u20_U1568  ( .A(1'b0), .ZN(_u10_u20_n2836 ) );
NAND2_X1 _u10_u20_U1567  ( .A1(_u10_u20_n2600 ), .A2(_u10_u20_n2836 ), .ZN(_u10_u20_n2428 ) );
INV_X1 _u10_u20_U1566  ( .A(_u10_u20_n2428 ), .ZN(_u10_u20_n2078 ) );
NAND2_X1 _u10_u20_U1565  ( .A1(_u10_u20_n2443 ), .A2(_u10_u20_n2078 ), .ZN(_u10_u20_n2282 ) );
INV_X1 _u10_u20_U1564  ( .A(1'b0), .ZN(_u10_u20_n2874 ) );
INV_X1 _u10_u20_U1563  ( .A(1'b0), .ZN(_u10_u20_n2031 ) );
NAND2_X1 _u10_u20_U1562  ( .A1(_u10_u20_n2874 ), .A2(_u10_u20_n2031 ), .ZN(_u10_u20_n1976 ) );
NOR2_X1 _u10_u20_U1561  ( .A1(_u10_u20_n2282 ), .A2(_u10_u20_n1976 ), .ZN(_u10_u20_n2411 ) );
NAND3_X1 _u10_u20_U1560  ( .A1(_u10_u20_n2467 ), .A2(_u10_u20_n1936 ), .A3(_u10_u20_n2411 ), .ZN(_u10_u20_n2464 ) );
NAND3_X1 _u10_u20_U1559  ( .A1(_u10_u20_n2166 ), .A2(_u10_u20_n2837 ), .A3(1'b0), .ZN(_u10_u20_n3276 ) );
INV_X1 _u10_u20_U1558  ( .A(_u10_u20_n3276 ), .ZN(_u10_u20_n2442 ) );
NAND3_X1 _u10_u20_U1557  ( .A1(_u10_u20_n2836 ), .A2(_u10_u20_n2080 ), .A3(_u10_u20_n2442 ), .ZN(_u10_u20_n2838 ) );
INV_X1 _u10_u20_U1556  ( .A(_u10_u20_n2838 ), .ZN(_u10_u20_n2850 ) );
NOR2_X1 _u10_u20_U1555  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u20_n2953 ) );
NAND2_X1 _u10_u20_U1554  ( .A1(_u10_u20_n2850 ), .A2(_u10_u20_n2953 ), .ZN(_u10_u20_n2947 ) );
INV_X1 _u10_u20_U1553  ( .A(_u10_u20_n2947 ), .ZN(_u10_u20_n2420 ) );
NAND2_X1 _u10_u20_U1552  ( .A1(_u10_u20_n1936 ), .A2(_u10_u20_n2874 ), .ZN(_u10_u20_n2030 ) );
INV_X1 _u10_u20_U1551  ( .A(_u10_u20_n2030 ), .ZN(_u10_u20_n2162 ) );
NAND2_X1 _u10_u20_U1550  ( .A1(_u10_u20_n2420 ), .A2(_u10_u20_n2162 ), .ZN(_u10_u20_n2828 ) );
INV_X1 _u10_u20_U1549  ( .A(_u10_u20_n2828 ), .ZN(_u10_u20_n2551 ) );
NAND2_X1 _u10_u20_U1548  ( .A1(_u10_u20_n2551 ), .A2(_u10_u20_n2467 ), .ZN(_u10_u20_n3416 ) );
NAND2_X1 _u10_u20_U1547  ( .A1(_u10_u20_n2464 ), .A2(_u10_u20_n3416 ), .ZN(_u10_u20_n2266 ) );
INV_X1 _u10_u20_U1546  ( .A(_u10_u20_n2266 ), .ZN(_u10_u20_n3410 ) );
NAND2_X1 _u10_u20_U1545  ( .A1(1'b0), .A2(_u10_u20_n2305 ), .ZN(_u10_u20_n3411 ) );
INV_X1 _u10_u20_U1544  ( .A(_u10_u20_n3356 ), .ZN(_u10_u20_n1983 ) );
NAND3_X1 _u10_u20_U1543  ( .A1(_u10_u20_n1983 ), .A2(_u10_u20_n2405 ), .A3(1'b0), .ZN(_u10_u20_n2022 ) );
INV_X1 _u10_u20_U1542  ( .A(_u10_u20_n2022 ), .ZN(_u10_u20_n2056 ) );
INV_X1 _u10_u20_U1541  ( .A(_u10_u20_n2840 ), .ZN(_u10_u20_n2059 ) );
INV_X1 _u10_u20_U1540  ( .A(1'b0), .ZN(_u10_u20_n1965 ) );
NAND2_X1 _u10_u20_U1539  ( .A1(_u10_u20_n2837 ), .A2(_u10_u20_n1965 ), .ZN(_u10_u20_n1852 ) );
INV_X1 _u10_u20_U1538  ( .A(_u10_u20_n1852 ), .ZN(_u10_u20_n3190 ) );
INV_X1 _u10_u20_U1537  ( .A(1'b0), .ZN(_u10_u20_n1853 ) );
NAND2_X1 _u10_u20_U1536  ( .A1(_u10_u20_n3190 ), .A2(_u10_u20_n1853 ), .ZN(_u10_u20_n2687 ) );
INV_X1 _u10_u20_U1535  ( .A(_u10_u20_n2687 ), .ZN(_u10_u20_n2019 ) );
NAND2_X1 _u10_u20_U1534  ( .A1(_u10_u20_n2059 ), .A2(_u10_u20_n2019 ), .ZN(_u10_u20_n2330 ) );
NOR2_X1 _u10_u20_U1533  ( .A1(_u10_u20_n2428 ), .A2(_u10_u20_n2330 ), .ZN(_u10_u20_n2036 ) );
NAND2_X1 _u10_u20_U1532  ( .A1(_u10_u20_n2056 ), .A2(_u10_u20_n2036 ), .ZN(_u10_u20_n3379 ) );
NOR2_X1 _u10_u20_U1531  ( .A1(_u10_u20_n3379 ), .A2(_u10_u20_n2030 ), .ZN(_u10_u20_n2026 ) );
INV_X1 _u10_u20_U1530  ( .A(1'b0), .ZN(_u10_u20_n2431 ) );
NOR2_X1 _u10_u20_U1529  ( .A1(_u10_u20_n2431 ), .A2(1'b0), .ZN(_u10_u20_n3062 ) );
NAND2_X1 _u10_u20_U1528  ( .A1(_u10_u20_n3062 ), .A2(_u10_u20_n2195 ), .ZN(_u10_u20_n3407 ) );
NOR3_X1 _u10_u20_U1527  ( .A1(_u10_u20_n2687 ), .A2(1'b0), .A3(_u10_u20_n3407 ), .ZN(_u10_u20_n3275 ) );
NAND3_X1 _u10_u20_U1526  ( .A1(_u10_u20_n2836 ), .A2(_u10_u20_n2080 ), .A3(_u10_u20_n3275 ), .ZN(_u10_u20_n3297 ) );
INV_X1 _u10_u20_U1525  ( .A(_u10_u20_n3297 ), .ZN(_u10_u20_n3172 ) );
NAND2_X1 _u10_u20_U1524  ( .A1(_u10_u20_n3172 ), .A2(_u10_u20_n2600 ), .ZN(_u10_u20_n2226 ) );
NOR2_X1 _u10_u20_U1523  ( .A1(_u10_u20_n2226 ), .A2(1'b0), .ZN(_u10_u20_n2307 ) );
INV_X1 _u10_u20_U1522  ( .A(_u10_u20_n2490 ), .ZN(_u10_u20_n2536 ) );
NAND3_X1 _u10_u20_U1521  ( .A1(_u10_u20_n2536 ), .A2(_u10_u20_n3040 ), .A3(1'b0), .ZN(_u10_u20_n3226 ) );
NOR2_X1 _u10_u20_U1520  ( .A1(_u10_u20_n3226 ), .A2(_u10_u20_n2330 ), .ZN(_u10_u20_n2441 ) );
NAND2_X1 _u10_u20_U1519  ( .A1(_u10_u20_n2441 ), .A2(_u10_u20_n2953 ), .ZN(_u10_u20_n2579 ) );
NOR2_X1 _u10_u20_U1518  ( .A1(_u10_u20_n2579 ), .A2(_u10_u20_n2030 ), .ZN(_u10_u20_n2550 ) );
NOR3_X1 _u10_u20_U1517  ( .A1(_u10_u20_n2026 ), .A2(_u10_u20_n2307 ), .A3(_u10_u20_n2550 ), .ZN(_u10_u20_n3394 ) );
NAND2_X1 _u10_u20_U1516  ( .A1(1'b0), .A2(_u10_u20_n2978 ), .ZN(_u10_u20_n3115 ) );
NOR2_X1 _u10_u20_U1515  ( .A1(_u10_u20_n3115 ), .A2(_u10_u20_n2330 ), .ZN(_u10_u20_n3126 ) );
NAND2_X1 _u10_u20_U1514  ( .A1(_u10_u20_n2162 ), .A2(_u10_u20_n2031 ), .ZN(_u10_u20_n2686 ) );
NOR2_X1 _u10_u20_U1513  ( .A1(_u10_u20_n2686 ), .A2(_u10_u20_n2428 ), .ZN(_u10_u20_n2108 ) );
NAND2_X1 _u10_u20_U1512  ( .A1(_u10_u20_n3126 ), .A2(_u10_u20_n2108 ), .ZN(_u10_u20_n3415 ) );
NAND2_X1 _u10_u20_U1511  ( .A1(_u10_u20_n3394 ), .A2(_u10_u20_n3415 ), .ZN(_u10_u20_n3089 ) );
NAND2_X1 _u10_u20_U1510  ( .A1(_u10_u20_n3089 ), .A2(_u10_u20_n2305 ), .ZN(_u10_u20_n3414 ) );
NAND2_X1 _u10_u20_U1509  ( .A1(_u10_u20_n2466 ), .A2(_u10_u20_n3414 ), .ZN(_u10_u20_n3118 ) );
NAND2_X1 _u10_u20_U1508  ( .A1(_u10_u20_n2078 ), .A2(_u10_u20_n2080 ), .ZN(_u10_u20_n2596 ) );
NAND2_X1 _u10_u20_U1507  ( .A1(1'b0), .A2(_u10_u20_n2493 ), .ZN(_u10_u20_n1961 ) );
NOR3_X1 _u10_u20_U1506  ( .A1(_u10_u20_n2490 ), .A2(1'b0), .A3(_u10_u20_n1961 ), .ZN(_u10_u20_n2054 ) );
NAND2_X1 _u10_u20_U1505  ( .A1(_u10_u20_n2054 ), .A2(_u10_u20_n3190 ), .ZN(_u10_u20_n2061 ) );
OR2_X1 _u10_u20_U1504  ( .A1(_u10_u20_n2596 ), .A2(_u10_u20_n2061 ), .ZN(_u10_u20_n1969 ) );
NOR3_X1 _u10_u20_U1503  ( .A1(_u10_u20_n1976 ), .A2(1'b0), .A3(_u10_u20_n1969 ), .ZN(_u10_u20_n2710 ) );
NAND2_X1 _u10_u20_U1502  ( .A1(_u10_u20_n2710 ), .A2(_u10_u20_n2467 ), .ZN(_u10_u20_n2545 ) );
INV_X1 _u10_u20_U1501  ( .A(_u10_u20_n2545 ), .ZN(_u10_u20_n2087 ) );
NOR2_X1 _u10_u20_U1500  ( .A1(_u10_u20_n3118 ), .A2(_u10_u20_n2087 ), .ZN(_u10_u20_n3145 ) );
NOR2_X1 _u10_u20_U1499  ( .A1(_u10_u20_n2030 ), .A2(1'b0), .ZN(_u10_u20_n2668 ) );
NAND2_X1 _u10_u20_U1498  ( .A1(1'b0), .A2(_u10_u20_n2668 ), .ZN(_u10_u20_n2163 ) );
INV_X1 _u10_u20_U1497  ( .A(_u10_u20_n2163 ), .ZN(_u10_u20_n2875 ) );
INV_X1 _u10_u20_U1496  ( .A(_u10_u20_n1976 ), .ZN(_u10_u20_n2747 ) );
NAND3_X1 _u10_u20_U1495  ( .A1(_u10_u20_n2747 ), .A2(_u10_u20_n2600 ), .A3(1'b0), .ZN(_u10_u20_n3393 ) );
NOR3_X1 _u10_u20_U1494  ( .A1(1'b0), .A2(1'b0), .A3(_u10_u20_n3393 ), .ZN(_u10_u20_n3180 ) );
INV_X1 _u10_u20_U1493  ( .A(1'b0), .ZN(_u10_u20_n2113 ) );
INV_X1 _u10_u20_U1492  ( .A(1'b0), .ZN(_u10_u20_n3066 ) );
NAND2_X1 _u10_u20_U1491  ( .A1(_u10_u20_n2175 ), .A2(_u10_u20_n3066 ), .ZN(_u10_u20_n2216 ) );
INV_X1 _u10_u20_U1490  ( .A(_u10_u20_n2659 ), .ZN(_u10_u20_n2643 ) );
NOR2_X1 _u10_u20_U1489  ( .A1(_u10_u20_n2216 ), .A2(_u10_u20_n2643 ), .ZN(_u10_u20_n2049 ) );
AND2_X1 _u10_u20_U1488  ( .A1(_u10_u20_n2049 ), .A2(_u10_u20_n1853 ), .ZN(_u10_u20_n3223 ) );
NAND2_X1 _u10_u20_U1487  ( .A1(_u10_u20_n3223 ), .A2(_u10_u20_n1965 ), .ZN(_u10_u20_n2531 ) );
NOR2_X1 _u10_u20_U1486  ( .A1(_u10_u20_n2531 ), .A2(1'b0), .ZN(_u10_u20_n2884 ) );
NAND2_X1 _u10_u20_U1485  ( .A1(_u10_u20_n2884 ), .A2(_u10_u20_n2166 ), .ZN(_u10_u20_n1841 ) );
NOR2_X1 _u10_u20_U1484  ( .A1(_u10_u20_n1841 ), .A2(1'b0), .ZN(_u10_u20_n3129 ) );
NAND2_X1 _u10_u20_U1483  ( .A1(_u10_u20_n3129 ), .A2(_u10_u20_n2836 ), .ZN(_u10_u20_n2842 ) );
INV_X1 _u10_u20_U1482  ( .A(_u10_u20_n2842 ), .ZN(_u10_u20_n2833 ) );
NAND2_X1 _u10_u20_U1481  ( .A1(_u10_u20_n2833 ), .A2(_u10_u20_n2600 ), .ZN(_u10_u20_n2853 ) );
INV_X1 _u10_u20_U1480  ( .A(_u10_u20_n2853 ), .ZN(_u10_u20_n2082 ) );
NAND2_X1 _u10_u20_U1479  ( .A1(_u10_u20_n2082 ), .A2(_u10_u20_n2031 ), .ZN(_u10_u20_n2274 ) );
INV_X1 _u10_u20_U1478  ( .A(_u10_u20_n2274 ), .ZN(_u10_u20_n2669 ) );
NAND3_X1 _u10_u20_U1477  ( .A1(_u10_u20_n2668 ), .A2(_u10_u20_n2113 ), .A3(_u10_u20_n2669 ), .ZN(_u10_u20_n1858 ) );
INV_X1 _u10_u20_U1476  ( .A(_u10_u20_n1858 ), .ZN(_u10_u20_n3067 ) );
NAND2_X1 _u10_u20_U1475  ( .A1(_u10_u20_n3067 ), .A2(1'b0), .ZN(_u10_u20_n2092 ) );
INV_X1 _u10_u20_U1474  ( .A(_u10_u20_n2092 ), .ZN(_u10_u20_n3294 ) );
INV_X1 _u10_u20_U1473  ( .A(1'b0), .ZN(_u10_u20_n2446 ) );
INV_X1 _u10_u20_U1472  ( .A(1'b0), .ZN(_u10_u20_n2996 ) );
NAND2_X1 _u10_u20_U1471  ( .A1(_u10_u20_n3067 ), .A2(_u10_u20_n2996 ), .ZN(_u10_u20_n1847 ) );
NOR3_X1 _u10_u20_U1470  ( .A1(_u10_u20_n2446 ), .A2(1'b0), .A3(_u10_u20_n1847 ), .ZN(_u10_u20_n3413 ) );
NOR4_X1 _u10_u20_U1469  ( .A1(_u10_u20_n2875 ), .A2(_u10_u20_n3180 ), .A3(_u10_u20_n3294 ), .A4(_u10_u20_n3413 ), .ZN(_u10_u20_n3412 ) );
NAND4_X1 _u10_u20_U1468  ( .A1(_u10_u20_n3410 ), .A2(_u10_u20_n3411 ), .A3(_u10_u20_n3145 ), .A4(_u10_u20_n3412 ), .ZN(_u10_u20_n3409 ) );
NAND2_X1 _u10_u20_U1467  ( .A1(_u10_u20_n2461 ), .A2(_u10_u20_n3409 ), .ZN(_u10_u20_n3380 ) );
NOR2_X1 _u10_u20_U1466  ( .A1(_u10_u20_n1817 ), .A2(_u10_u20_n1816 ), .ZN(_u10_u20_n3368 ) );
AND2_X1 _u10_u20_U1465  ( .A1(_u10_u20_n3368 ), .A2(_u10_u20_n1813 ), .ZN(_u10_u20_n3320 ) );
NOR2_X1 _u10_u20_U1464  ( .A1(_u10_SYNOPSYS_UNCONNECTED_7 ), .A2(_u10_u20_n1815 ), .ZN(_u10_u20_n3236 ) );
NAND2_X1 _u10_u20_U1463  ( .A1(_u10_u20_n3320 ), .A2(_u10_u20_n3236 ), .ZN(_u10_u20_n2607 ) );
INV_X1 _u10_u20_U1462  ( .A(_u10_u20_n2607 ), .ZN(_u10_u20_n1966 ) );
INV_X1 _u10_u20_U1461  ( .A(_u10_u20_n2200 ), .ZN(_u10_u20_n3216 ) );
NAND2_X1 _u10_u20_U1460  ( .A1(1'b0), .A2(_u10_u20_n3216 ), .ZN(_u10_u20_n2367 ) );
INV_X1 _u10_u20_U1459  ( .A(_u10_u20_n2367 ), .ZN(_u10_u20_n3183 ) );
NAND2_X1 _u10_u20_U1458  ( .A1(_u10_u20_n3183 ), .A2(_u10_u20_n2195 ), .ZN(_u10_u20_n2194 ) );
INV_X1 _u10_u20_U1457  ( .A(_u10_u20_n2194 ), .ZN(_u10_u20_n2055 ) );
NAND2_X1 _u10_u20_U1456  ( .A1(_u10_u20_n2055 ), .A2(_u10_u20_n1853 ), .ZN(_u10_u20_n3401 ) );
INV_X1 _u10_u20_U1455  ( .A(_u10_u20_n2531 ), .ZN(_u10_u20_n2190 ) );
INV_X1 _u10_u20_U1454  ( .A(1'b0), .ZN(_u10_u20_n3001 ) );
NAND2_X1 _u10_u20_U1453  ( .A1(_u10_u20_n3001 ), .A2(_u10_u20_n2466 ), .ZN(_u10_u20_n2156 ) );
NOR2_X1 _u10_u20_U1452  ( .A1(_u10_u20_n2166 ), .A2(_u10_u20_n2596 ), .ZN(_u10_u20_n2594 ) );
NAND2_X1 _u10_u20_U1451  ( .A1(_u10_u20_n2594 ), .A2(_u10_u20_n2031 ), .ZN(_u10_u20_n2752 ) );
INV_X1 _u10_u20_U1450  ( .A(_u10_u20_n2752 ), .ZN(_u10_u20_n2421 ) );
NAND2_X1 _u10_u20_U1449  ( .A1(_u10_u20_n2421 ), .A2(_u10_u20_n2874 ), .ZN(_u10_u20_n2033 ) );
INV_X1 _u10_u20_U1448  ( .A(_u10_u20_n2033 ), .ZN(_u10_u20_n2742 ) );
NAND3_X1 _u10_u20_U1447  ( .A1(_u10_u20_n2305 ), .A2(_u10_u20_n1936 ), .A3(_u10_u20_n2742 ), .ZN(_u10_u20_n1896 ) );
OR3_X1 _u10_u20_U1446  ( .A1(_u10_u20_n2156 ), .A2(1'b0), .A3(_u10_u20_n1896 ), .ZN(_u10_u20_n2905 ) );
NAND2_X1 _u10_u20_U1445  ( .A1(_u10_u20_n2113 ), .A2(_u10_u20_n2996 ), .ZN(_u10_u20_n2719 ) );
NOR2_X1 _u10_u20_U1444  ( .A1(_u10_u20_n2719 ), .A2(1'b0), .ZN(_u10_u20_n2941 ) );
INV_X1 _u10_u20_U1443  ( .A(_u10_u20_n2941 ), .ZN(_u10_u20_n2911 ) );
NOR2_X1 _u10_u20_U1442  ( .A1(_u10_u20_n2905 ), .A2(_u10_u20_n2911 ), .ZN(_u10_u20_n3222 ) );
INV_X1 _u10_u20_U1441  ( .A(_u10_u20_n3222 ), .ZN(_u10_u20_n2695 ) );
INV_X1 _u10_u20_U1440  ( .A(_u10_u20_n2156 ), .ZN(_u10_u20_n2089 ) );
NAND3_X1 _u10_u20_U1439  ( .A1(_u10_u20_n2089 ), .A2(_u10_u20_n2446 ), .A3(_u10_u20_n3180 ), .ZN(_u10_u20_n2902 ) );
NOR2_X1 _u10_u20_U1438  ( .A1(_u10_u20_n2902 ), .A2(_u10_u20_n2911 ), .ZN(_u10_u20_n2533 ) );
INV_X1 _u10_u20_U1437  ( .A(_u10_u20_n2533 ), .ZN(_u10_u20_n2485 ) );
NAND2_X1 _u10_u20_U1436  ( .A1(_u10_u20_n2695 ), .A2(_u10_u20_n2485 ), .ZN(_u10_u20_n2721 ) );
NAND2_X1 _u10_u20_U1435  ( .A1(1'b0), .A2(_u10_u20_n2113 ), .ZN(_u10_u20_n1868 ) );
INV_X1 _u10_u20_U1434  ( .A(_u10_u20_n1868 ), .ZN(_u10_u20_n2534 ) );
NOR2_X1 _u10_u20_U1433  ( .A1(_u10_u20_n2721 ), .A2(_u10_u20_n2534 ), .ZN(_u10_u20_n3231 ) );
NAND2_X1 _u10_u20_U1432  ( .A1(_u10_u20_n2467 ), .A2(_u10_u20_n3001 ), .ZN(_u10_u20_n2303 ) );
INV_X1 _u10_u20_U1431  ( .A(_u10_u20_n2303 ), .ZN(_u10_u20_n2549 ) );
INV_X1 _u10_u20_U1430  ( .A(1'b0), .ZN(_u10_u20_n2803 ) );
NAND2_X1 _u10_u20_U1429  ( .A1(_u10_u20_n2803 ), .A2(_u10_u20_n2446 ), .ZN(_u10_u20_n1846 ) );
INV_X1 _u10_u20_U1428  ( .A(_u10_u20_n1846 ), .ZN(_u10_u20_n2667 ) );
NAND3_X1 _u10_u20_U1427  ( .A1(_u10_u20_n2549 ), .A2(_u10_u20_n2667 ), .A3(1'b0), .ZN(_u10_u20_n2739 ) );
INV_X1 _u10_u20_U1426  ( .A(_u10_u20_n2739 ), .ZN(_u10_u20_n3272 ) );
INV_X1 _u10_u20_U1425  ( .A(_u10_u20_n2719 ), .ZN(_u10_u20_n2364 ) );
NAND2_X1 _u10_u20_U1424  ( .A1(_u10_u20_n3272 ), .A2(_u10_u20_n2364 ), .ZN(_u10_u20_n2852 ) );
INV_X1 _u10_u20_U1423  ( .A(_u10_u20_n2852 ), .ZN(_u10_u20_n2214 ) );
NAND2_X1 _u10_u20_U1422  ( .A1(_u10_u20_n2875 ), .A2(_u10_u20_n2089 ), .ZN(_u10_u20_n2097 ) );
INV_X1 _u10_u20_U1421  ( .A(_u10_u20_n2097 ), .ZN(_u10_u20_n2300 ) );
NAND2_X1 _u10_u20_U1420  ( .A1(_u10_u20_n2300 ), .A2(_u10_u20_n2446 ), .ZN(_u10_u20_n2001 ) );
NOR2_X1 _u10_u20_U1419  ( .A1(_u10_u20_n2001 ), .A2(_u10_u20_n2911 ), .ZN(_u10_u20_n2877 ) );
NOR2_X1 _u10_u20_U1418  ( .A1(_u10_u20_n2214 ), .A2(_u10_u20_n2877 ), .ZN(_u10_u20_n2940 ) );
NAND2_X1 _u10_u20_U1417  ( .A1(_u10_u20_n3231 ), .A2(_u10_u20_n2940 ), .ZN(_u10_u20_n3408 ) );
NAND2_X1 _u10_u20_U1416  ( .A1(_u10_u20_n2190 ), .A2(_u10_u20_n3408 ), .ZN(_u10_u20_n3402 ) );
NOR2_X1 _u10_u20_U1415  ( .A1(_u10_u20_n2446 ), .A2(_u10_u20_n2911 ), .ZN(_u10_u20_n3059 ) );
NAND2_X1 _u10_u20_U1414  ( .A1(_u10_u20_n3059 ), .A2(_u10_u20_n2190 ), .ZN(_u10_u20_n3404 ) );
AND3_X1 _u10_u20_U1413  ( .A1(_u10_u20_n3407 ), .A2(_u10_u20_n3226 ), .A3(_u10_u20_n3115 ), .ZN(_u10_u20_n3058 ) );
NAND2_X1 _u10_u20_U1412  ( .A1(_u10_u20_n3058 ), .A2(_u10_u20_n2022 ), .ZN(_u10_u20_n3406 ) );
NAND2_X1 _u10_u20_U1411  ( .A1(_u10_u20_n1853 ), .A2(_u10_u20_n3406 ), .ZN(_u10_u20_n3405 ) );
AND3_X1 _u10_u20_U1410  ( .A1(_u10_u20_n3404 ), .A2(_u10_u20_n1965 ), .A3(_u10_u20_n3405 ), .ZN(_u10_u20_n3063 ) );
NAND2_X1 _u10_u20_U1409  ( .A1(_u10_u20_n2667 ), .A2(_u10_u20_n3001 ), .ZN(_u10_u20_n1898 ) );
INV_X1 _u10_u20_U1408  ( .A(_u10_u20_n1898 ), .ZN(_u10_u20_n2835 ) );
NAND3_X1 _u10_u20_U1407  ( .A1(_u10_u20_n2364 ), .A2(_u10_u20_n2835 ), .A3(1'b0), .ZN(_u10_u20_n1869 ) );
NOR2_X1 _u10_u20_U1406  ( .A1(_u10_u20_n1869 ), .A2(_u10_u20_n2531 ), .ZN(_u10_u20_n2761 ) );
NOR3_X1 _u10_u20_U1405  ( .A1(_u10_u20_n2761 ), .A2(_u10_u20_n2528 ), .A3(_u10_u20_n2054 ), .ZN(_u10_u20_n3403 ) );
NAND4_X1 _u10_u20_U1404  ( .A1(_u10_u20_n3401 ), .A2(_u10_u20_n3402 ), .A3(_u10_u20_n3063 ), .A4(_u10_u20_n3403 ), .ZN(_u10_u20_n3400 ) );
NAND2_X1 _u10_u20_U1403  ( .A1(_u10_u20_n1966 ), .A2(_u10_u20_n3400 ), .ZN(_u10_u20_n3381 ) );
AND2_X1 _u10_u20_U1402  ( .A1(_u10_u20_n3368 ), .A2(_u10_SYNOPSYS_UNCONNECTED_8 ), .ZN(_u10_u20_n3319 ) );
NAND2_X1 _u10_u20_U1401  ( .A1(_u10_u20_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_7 ), .ZN(_u10_u20_n1849 ) );
INV_X1 _u10_u20_U1400  ( .A(_u10_u20_n1849 ), .ZN(_u10_u20_n2183 ) );
NAND2_X1 _u10_u20_U1399  ( .A1(_u10_u20_n2884 ), .A2(_u10_u20_n2183 ), .ZN(_u10_u20_n2883 ) );
INV_X1 _u10_u20_U1398  ( .A(_u10_u20_n2883 ), .ZN(_u10_u20_n1890 ) );
INV_X1 _u10_u20_U1397  ( .A(_u10_u20_n2940 ), .ZN(_u10_u20_n3278 ) );
NAND2_X1 _u10_u20_U1396  ( .A1(_u10_u20_n1890 ), .A2(_u10_u20_n3278 ), .ZN(_u10_u20_n3382 ) );
NAND2_X1 _u10_u20_U1395  ( .A1(_u10_u20_n3059 ), .A2(_u10_u20_n2669 ), .ZN(_u10_u20_n3399 ) );
NAND2_X1 _u10_u20_U1394  ( .A1(_u10_u20_n2031 ), .A2(_u10_u20_n3399 ), .ZN(_u10_u20_n3398 ) );
NAND2_X1 _u10_u20_U1393  ( .A1(_u10_u20_n2162 ), .A2(_u10_u20_n3398 ), .ZN(_u10_u20_n3395 ) );
NAND3_X1 _u10_u20_U1392  ( .A1(_u10_u20_n2747 ), .A2(_u10_u20_n2078 ), .A3(_u10_u20_n3126 ), .ZN(_u10_u20_n3396 ) );
NAND2_X1 _u10_u20_U1391  ( .A1(_u10_u20_n2055 ), .A2(_u10_u20_n2036 ), .ZN(_u10_u20_n2285 ) );
NOR2_X1 _u10_u20_U1390  ( .A1(_u10_u20_n2285 ), .A2(_u10_u20_n2030 ), .ZN(_u10_u20_n3349 ) );
INV_X1 _u10_u20_U1389  ( .A(_u10_u20_n3349 ), .ZN(_u10_u20_n1933 ) );
INV_X1 _u10_u20_U1388  ( .A(_u10_u20_n2710 ), .ZN(_u10_u20_n3397 ) );
NAND4_X1 _u10_u20_U1387  ( .A1(_u10_u20_n3395 ), .A2(_u10_u20_n3396 ), .A3(_u10_u20_n1933 ), .A4(_u10_u20_n3397 ), .ZN(_u10_u20_n3389 ) );
NAND2_X1 _u10_u20_U1386  ( .A1(_u10_u20_n1936 ), .A2(_u10_u20_n2828 ), .ZN(_u10_u20_n3141 ) );
INV_X1 _u10_u20_U1385  ( .A(_u10_u20_n3141 ), .ZN(_u10_u20_n2302 ) );
NAND2_X1 _u10_u20_U1384  ( .A1(_u10_u20_n3394 ), .A2(_u10_u20_n2302 ), .ZN(_u10_u20_n3390 ) );
NOR2_X1 _u10_u20_U1383  ( .A1(_u10_u20_n1869 ), .A2(_u10_u20_n2274 ), .ZN(_u10_u20_n3378 ) );
INV_X1 _u10_u20_U1382  ( .A(_u10_u20_n3378 ), .ZN(_u10_u20_n2748 ) );
NOR2_X1 _u10_u20_U1381  ( .A1(1'b0), .A2(_u10_u20_n2748 ), .ZN(_u10_u20_n3391 ) );
NAND2_X1 _u10_u20_U1380  ( .A1(_u10_u20_n2534 ), .A2(_u10_u20_n2669 ), .ZN(_u10_u20_n2383 ) );
INV_X1 _u10_u20_U1379  ( .A(_u10_u20_n2383 ), .ZN(_u10_u20_n1978 ) );
NAND2_X1 _u10_u20_U1378  ( .A1(_u10_u20_n1978 ), .A2(_u10_u20_n2874 ), .ZN(_u10_u20_n3392 ) );
INV_X1 _u10_u20_U1377  ( .A(_u10_u20_n2411 ), .ZN(_u10_u20_n2164 ) );
NAND4_X1 _u10_u20_U1376  ( .A1(_u10_u20_n3392 ), .A2(_u10_u20_n3393 ), .A3(_u10_u20_n2033 ), .A4(_u10_u20_n2164 ), .ZN(_u10_u20_n2476 ) );
NOR4_X1 _u10_u20_U1375  ( .A1(_u10_u20_n3389 ), .A2(_u10_u20_n3390 ), .A3(_u10_u20_n3391 ), .A4(_u10_u20_n2476 ), .ZN(_u10_u20_n3388 ) );
NAND2_X1 _u10_u20_U1374  ( .A1(_u10_u20_n3236 ), .A2(_u10_u20_n3328 ), .ZN(_u10_u20_n2025 ) );
NOR2_X1 _u10_u20_U1373  ( .A1(_u10_u20_n3388 ), .A2(_u10_u20_n2025 ), .ZN(_u10_u20_n3384 ) );
NOR2_X1 _u10_u20_U1372  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u20_n2152 ) );
NAND2_X1 _u10_u20_U1371  ( .A1(_u10_u20_n2152 ), .A2(_u10_u20_n2175 ), .ZN(_u10_u20_n2722 ) );
INV_X1 _u10_u20_U1370  ( .A(_u10_u20_n2722 ), .ZN(_u10_u20_n2588 ) );
NAND2_X1 _u10_u20_U1369  ( .A1(_u10_u20_n2549 ), .A2(_u10_u20_n3349 ), .ZN(_u10_u20_n2091 ) );
NOR2_X1 _u10_u20_U1368  ( .A1(_u10_u20_n2091 ), .A2(_u10_u20_n1846 ), .ZN(_u10_u20_n2128 ) );
NAND3_X1 _u10_u20_U1367  ( .A1(_u10_u20_n3066 ), .A2(_u10_u20_n2113 ), .A3(_u10_u20_n2128 ), .ZN(_u10_u20_n2342 ) );
INV_X1 _u10_u20_U1366  ( .A(_u10_u20_n2342 ), .ZN(_u10_u20_n3316 ) );
NAND2_X1 _u10_u20_U1365  ( .A1(_u10_u20_n2588 ), .A2(_u10_u20_n3316 ), .ZN(_u10_u20_n2142 ) );
NOR2_X1 _u10_u20_U1364  ( .A1(_u10_u20_n1954 ), .A2(_u10_u20_n1898 ), .ZN(_u10_u20_n2255 ) );
NAND2_X1 _u10_u20_U1363  ( .A1(_u10_u20_n2255 ), .A2(_u10_u20_n2996 ), .ZN(_u10_u20_n1915 ) );
INV_X1 _u10_u20_U1362  ( .A(_u10_u20_n1915 ), .ZN(_u10_u20_n2251 ) );
NAND2_X1 _u10_u20_U1361  ( .A1(_u10_u20_n2251 ), .A2(_u10_u20_n2113 ), .ZN(_u10_u20_n1925 ) );
INV_X1 _u10_u20_U1360  ( .A(_u10_u20_n2026 ), .ZN(_u10_u20_n3340 ) );
NOR3_X1 _u10_u20_U1359  ( .A1(_u10_u20_n1925 ), .A2(_u10_u20_n2216 ), .A3(_u10_u20_n3340 ), .ZN(_u10_u20_n2003 ) );
INV_X1 _u10_u20_U1358  ( .A(1'b0), .ZN(_u10_u20_n1930 ) );
NAND2_X1 _u10_u20_U1357  ( .A1(_u10_u20_n2003 ), .A2(_u10_u20_n1930 ), .ZN(_u10_u20_n3387 ) );
AND2_X1 _u10_u20_U1356  ( .A1(_u10_u20_n2142 ), .A2(_u10_u20_n3387 ), .ZN(_u10_u20_n3366 ) );
NOR3_X1 _u10_u20_U1355  ( .A1(_u10_u20_n1813 ), .A2(_u10_u20_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_4 ), .ZN(_u10_u20_n3360 ) );
NOR2_X1 _u10_u20_U1354  ( .A1(_u10_SYNOPSYS_UNCONNECTED_6 ), .A2(_u10_SYNOPSYS_UNCONNECTED_7 ), .ZN(_u10_u20_n3136 ) );
NAND2_X1 _u10_u20_U1353  ( .A1(_u10_u20_n3360 ), .A2(_u10_u20_n3136 ), .ZN(_u10_u20_n2344 ) );
NOR2_X1 _u10_u20_U1352  ( .A1(_u10_u20_n3366 ), .A2(_u10_u20_n2344 ), .ZN(_u10_u20_n3385 ) );
NOR3_X1 _u10_u20_U1351  ( .A1(_u10_SYNOPSYS_UNCONNECTED_4 ), .A2(_u10_u20_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_8 ), .ZN(_u10_u20_n3342 ) );
NAND2_X1 _u10_u20_U1350  ( .A1(_u10_u20_n3342 ), .A2(_u10_u20_n3136 ), .ZN(_u10_u20_n2584 ) );
NOR2_X1 _u10_u20_U1349  ( .A1(_u10_u20_n2584 ), .A2(1'b0), .ZN(_u10_u20_n2139 ) );
INV_X1 _u10_u20_U1348  ( .A(_u10_u20_n2216 ), .ZN(_u10_u20_n2106 ) );
AND2_X1 _u10_u20_U1347  ( .A1(_u10_u20_n2152 ), .A2(_u10_u20_n2106 ), .ZN(_u10_u20_n2336 ) );
NAND2_X1 _u10_u20_U1346  ( .A1(_u10_u20_n2139 ), .A2(_u10_u20_n2336 ), .ZN(_u10_u20_n2365 ) );
INV_X1 _u10_u20_U1345  ( .A(_u10_u20_n2365 ), .ZN(_u10_u20_n2004 ) );
AND2_X1 _u10_u20_U1344  ( .A1(_u10_u20_n2877 ), .A2(_u10_u20_n2004 ), .ZN(_u10_u20_n3386 ) );
NOR3_X1 _u10_u20_U1343  ( .A1(_u10_u20_n3384 ), .A2(_u10_u20_n3385 ), .A3(_u10_u20_n3386 ), .ZN(_u10_u20_n3383 ) );
NAND4_X1 _u10_u20_U1342  ( .A1(_u10_u20_n3380 ), .A2(_u10_u20_n3381 ), .A3(_u10_u20_n3382 ), .A4(_u10_u20_n3383 ), .ZN(_u10_u20_n3191 ) );
NAND2_X1 _u10_u20_U1341  ( .A1(_u10_u20_n2285 ), .A2(_u10_u20_n3379 ), .ZN(_u10_u20_n1975 ) );
NOR3_X1 _u10_u20_U1340  ( .A1(_u10_u20_n3378 ), .A2(1'b0), .A3(_u10_u20_n1975 ), .ZN(_u10_u20_n3122 ) );
AND4_X1 _u10_u20_U1339  ( .A1(_u10_u20_n2752 ), .A2(_u10_u20_n2383 ), .A3(_u10_u20_n1969 ), .A4(_u10_u20_n3122 ), .ZN(_u10_u20_n3377 ) );
NOR2_X1 _u10_u20_U1338  ( .A1(_u10_u20_n1814 ), .A2(_u10_u20_n1815 ), .ZN(_u10_u20_n3147 ) );
NAND2_X1 _u10_u20_U1337  ( .A1(_u10_u20_n3328 ), .A2(_u10_u20_n3147 ), .ZN(_u10_u20_n2359 ) );
NOR2_X1 _u10_u20_U1336  ( .A1(_u10_u20_n3377 ), .A2(_u10_u20_n2359 ), .ZN(_u10_u20_n3362 ) );
INV_X1 _u10_u20_U1335  ( .A(_u10_u20_n2008 ), .ZN(_u10_u20_n3097 ) );
NOR3_X1 _u10_u20_U1334  ( .A1(_u10_SYNOPSYS_UNCONNECTED_4 ), .A2(_u10_u20_n1813 ), .A3(_u10_SYNOPSYS_UNCONNECTED_5 ), .ZN(_u10_u20_n3269 ) );
NAND2_X1 _u10_u20_U1333  ( .A1(_u10_u20_n3269 ), .A2(_u10_u20_n3136 ), .ZN(_u10_u20_n3109 ) );
INV_X1 _u10_u20_U1332  ( .A(_u10_u20_n3109 ), .ZN(_u10_u20_n2999 ) );
INV_X1 _u10_u20_U1331  ( .A(_u10_u20_n2508 ), .ZN(_u10_u20_n2103 ) );
NAND2_X1 _u10_u20_U1330  ( .A1(_u10_u20_n2336 ), .A2(_u10_u20_n2103 ), .ZN(_u10_u20_n2249 ) );
NOR2_X1 _u10_u20_U1329  ( .A1(_u10_u20_n2249 ), .A2(1'b0), .ZN(_u10_u20_n1866 ) );
NAND2_X1 _u10_u20_U1328  ( .A1(_u10_u20_n1866 ), .A2(_u10_u20_n1922 ), .ZN(_u10_u20_n2632 ) );
INV_X1 _u10_u20_U1327  ( .A(_u10_u20_n2223 ), .ZN(_u10_u20_n1918 ) );
NOR2_X1 _u10_u20_U1326  ( .A1(_u10_u20_n2632 ), .A2(_u10_u20_n1918 ), .ZN(_u10_u20_n1981 ) );
NAND3_X1 _u10_u20_U1325  ( .A1(_u10_u20_n3097 ), .A2(_u10_u20_n2999 ), .A3(_u10_u20_n1981 ), .ZN(_u10_u20_n3034 ) );
NOR3_X1 _u10_u20_U1324  ( .A1(_u10_SYNOPSYS_UNCONNECTED_5 ), .A2(_u10_SYNOPSYS_UNCONNECTED_4 ), .A3(_u10_SYNOPSYS_UNCONNECTED_8 ), .ZN(_u10_u20_n3302 ) );
NAND2_X1 _u10_u20_U1323  ( .A1(_u10_u20_n3302 ), .A2(_u10_u20_n3174 ), .ZN(_u10_u20_n3162 ) );
INV_X1 _u10_u20_U1322  ( .A(_u10_u20_n3162 ), .ZN(_u10_u20_n2979 ) );
NAND2_X1 _u10_u20_U1321  ( .A1(_u10_u20_n2979 ), .A2(_u10_u20_n2972 ), .ZN(_u10_u20_n1984 ) );
AND2_X1 _u10_u20_U1320  ( .A1(_u10_u20_n3302 ), .A2(_u10_u20_n3136 ), .ZN(_u10_u20_n2977 ) );
NAND3_X1 _u10_u20_U1319  ( .A1(_u10_u20_n2977 ), .A2(_u10_u20_n3000 ), .A3(_u10_u20_n3097 ), .ZN(_u10_u20_n3376 ) );
NAND2_X1 _u10_u20_U1318  ( .A1(_u10_u20_n1984 ), .A2(_u10_u20_n3376 ), .ZN(_u10_u20_n3375 ) );
NAND2_X1 _u10_u20_U1317  ( .A1(_u10_u20_n1981 ), .A2(_u10_u20_n3375 ), .ZN(_u10_u20_n2798 ) );
NAND2_X1 _u10_u20_U1316  ( .A1(_u10_u20_n3034 ), .A2(_u10_u20_n2798 ), .ZN(_u10_u20_n2007 ) );
NAND2_X1 _u10_u20_U1315  ( .A1(_u10_u20_n3269 ), .A2(_u10_u20_n3147 ), .ZN(_u10_u20_n2102 ) );
NOR2_X1 _u10_u20_U1314  ( .A1(_u10_u20_n2249 ), .A2(_u10_u20_n2102 ), .ZN(_u10_u20_n3323 ) );
INV_X1 _u10_u20_U1313  ( .A(_u10_u20_n3323 ), .ZN(_u10_u20_n3374 ) );
INV_X1 _u10_u20_U1312  ( .A(_u10_u20_n2344 ), .ZN(_u10_u20_n2002 ) );
NAND2_X1 _u10_u20_U1311  ( .A1(_u10_u20_n2336 ), .A2(_u10_u20_n2002 ), .ZN(_u10_u20_n3225 ) );
NAND2_X1 _u10_u20_U1310  ( .A1(_u10_u20_n3374 ), .A2(_u10_u20_n3225 ), .ZN(_u10_u20_n2488 ) );
NAND2_X1 _u10_u20_U1309  ( .A1(_u10_u20_n3342 ), .A2(_u10_u20_n3236 ), .ZN(_u10_u20_n2253 ) );
NOR2_X1 _u10_u20_U1308  ( .A1(_u10_u20_n2253 ), .A2(1'b0), .ZN(_u10_u20_n1885 ) );
NAND2_X1 _u10_u20_U1307  ( .A1(_u10_u20_n3360 ), .A2(_u10_u20_n3174 ), .ZN(_u10_u20_n2254 ) );
INV_X1 _u10_u20_U1306  ( .A(_u10_u20_n2254 ), .ZN(_u10_u20_n2986 ) );
NAND2_X1 _u10_u20_U1305  ( .A1(_u10_u20_n2106 ), .A2(_u10_u20_n2986 ), .ZN(_u10_u20_n1913 ) );
INV_X1 _u10_u20_U1304  ( .A(_u10_u20_n1913 ), .ZN(_u10_u20_n2377 ) );
OR4_X1 _u10_u20_U1303  ( .A1(_u10_u20_n2007 ), .A2(_u10_u20_n2488 ), .A3(_u10_u20_n1885 ), .A4(_u10_u20_n2377 ), .ZN(_u10_u20_n3373 ) );
NAND2_X1 _u10_u20_U1302  ( .A1(_u10_u20_n2534 ), .A2(_u10_u20_n3373 ), .ZN(_u10_u20_n3370 ) );
NAND2_X1 _u10_u20_U1301  ( .A1(_u10_u20_n3342 ), .A2(_u10_u20_n3174 ), .ZN(_u10_u20_n2037 ) );
NAND2_X1 _u10_u20_U1300  ( .A1(_u10_u20_n2037 ), .A2(_u10_u20_n2254 ), .ZN(_u10_u20_n3372 ) );
NAND2_X1 _u10_u20_U1299  ( .A1(_u10_u20_n2003 ), .A2(_u10_u20_n3372 ), .ZN(_u10_u20_n3371 ) );
NAND2_X1 _u10_u20_U1298  ( .A1(_u10_u20_n3370 ), .A2(_u10_u20_n3371 ), .ZN(_u10_u20_n3363 ) );
NOR2_X1 _u10_u20_U1297  ( .A1(_u10_u20_n2490 ), .A2(_u10_u20_n1961 ), .ZN(_u10_u20_n3369 ) );
NAND2_X1 _u10_u20_U1296  ( .A1(_u10_u20_n2534 ), .A2(_u10_u20_n2049 ), .ZN(_u10_u20_n2646 ) );
INV_X1 _u10_u20_U1295  ( .A(_u10_u20_n2646 ), .ZN(_u10_u20_n3055 ) );
NOR2_X1 _u10_u20_U1294  ( .A1(_u10_u20_n3369 ), .A2(_u10_u20_n3055 ), .ZN(_u10_u20_n3367 ) );
NAND2_X1 _u10_u20_U1293  ( .A1(_u10_u20_n3368 ), .A2(_u10_u20_n3147 ), .ZN(_u10_u20_n2495 ) );
NOR2_X1 _u10_u20_U1292  ( .A1(_u10_u20_n3367 ), .A2(_u10_u20_n2495 ), .ZN(_u10_u20_n3364 ) );
INV_X1 _u10_u20_U1291  ( .A(_u10_u20_n2139 ), .ZN(_u10_u20_n3254 ) );
NOR2_X1 _u10_u20_U1290  ( .A1(_u10_u20_n3366 ), .A2(_u10_u20_n3254 ), .ZN(_u10_u20_n3365 ) );
NOR4_X1 _u10_u20_U1289  ( .A1(_u10_u20_n3362 ), .A2(_u10_u20_n3363 ), .A3(_u10_u20_n3364 ), .A4(_u10_u20_n3365 ), .ZN(_u10_u20_n3305 ) );
NAND2_X1 _u10_u20_U1288  ( .A1(_u10_u20_n3302 ), .A2(_u10_u20_n3147 ), .ZN(_u10_u20_n2980 ) );
NAND2_X1 _u10_u20_U1287  ( .A1(_u10_u20_n2102 ), .A2(_u10_u20_n2980 ), .ZN(_u10_u20_n2177 ) );
NAND2_X1 _u10_u20_U1286  ( .A1(_u10_u20_n2003 ), .A2(_u10_u20_n2493 ), .ZN(_u10_u20_n1962 ) );
NAND2_X1 _u10_u20_U1285  ( .A1(_u10_u20_n1961 ), .A2(_u10_u20_n1962 ), .ZN(_u10_u20_n3361 ) );
NAND2_X1 _u10_u20_U1284  ( .A1(_u10_u20_n2177 ), .A2(_u10_u20_n3361 ), .ZN(_u10_u20_n3357 ) );
NAND2_X1 _u10_u20_U1283  ( .A1(_u10_u20_n3236 ), .A2(_u10_u20_n3360 ), .ZN(_u10_u20_n1859 ) );
INV_X1 _u10_u20_U1282  ( .A(_u10_u20_n1859 ), .ZN(_u10_u20_n2256 ) );
NAND3_X1 _u10_u20_U1281  ( .A1(_u10_u20_n2256 ), .A2(_u10_u20_n2113 ), .A3(_u10_u20_n2128 ), .ZN(_u10_u20_n3358 ) );
NOR2_X1 _u10_u20_U1280  ( .A1(_u10_u20_n2877 ), .A2(_u10_u20_n3222 ), .ZN(_u10_u20_n3347 ) );
NAND2_X1 _u10_u20_U1279  ( .A1(_u10_u20_n3347 ), .A2(_u10_u20_n1869 ), .ZN(_u10_u20_n2005 ) );
NAND2_X1 _u10_u20_U1278  ( .A1(_u10_u20_n2488 ), .A2(_u10_u20_n2005 ), .ZN(_u10_u20_n3359 ) );
NAND3_X1 _u10_u20_U1277  ( .A1(_u10_u20_n3357 ), .A2(_u10_u20_n3358 ), .A3(_u10_u20_n3359 ), .ZN(_u10_u20_n3352 ) );
NAND2_X1 _u10_u20_U1276  ( .A1(_u10_u20_n3320 ), .A2(_u10_u20_n3136 ), .ZN(_u10_u20_n2356 ) );
INV_X1 _u10_u20_U1275  ( .A(_u10_u20_n2356 ), .ZN(_u10_u20_n2830 ) );
NAND2_X1 _u10_u20_U1274  ( .A1(_u10_u20_n2830 ), .A2(_u10_u20_n2836 ), .ZN(_u10_u20_n2291 ) );
NOR3_X1 _u10_u20_U1273  ( .A1(_u10_u20_n2291 ), .A2(_u10_u20_n2330 ), .A3(_u10_u20_n2022 ), .ZN(_u10_u20_n3353 ) );
INV_X1 _u10_u20_U1272  ( .A(_u10_u20_n1925 ), .ZN(_u10_u20_n2105 ) );
AND2_X1 _u10_u20_U1271  ( .A1(_u10_u20_n2108 ), .A2(_u10_u20_n2105 ), .ZN(_u10_u20_n2915 ) );
INV_X1 _u10_u20_U1270  ( .A(_u10_u20_n2330 ), .ZN(_u10_u20_n2107 ) );
NAND2_X1 _u10_u20_U1269  ( .A1(_u10_u20_n2915 ), .A2(_u10_u20_n2107 ), .ZN(_u10_u20_n2203 ) );
INV_X1 _u10_u20_U1268  ( .A(_u10_u20_n2203 ), .ZN(_u10_u20_n1982 ) );
NAND2_X1 _u10_u20_U1267  ( .A1(_u10_u20_n1982 ), .A2(_u10_u20_n2536 ), .ZN(_u10_u20_n2587 ) );
INV_X1 _u10_u20_U1266  ( .A(_u10_u20_n2587 ), .ZN(_u10_u20_n2697 ) );
NAND3_X1 _u10_u20_U1265  ( .A1(_u10_u20_n2697 ), .A2(_u10_u20_n2493 ), .A3(_u10_u20_n2377 ), .ZN(_u10_u20_n2412 ) );
INV_X1 _u10_u20_U1264  ( .A(_u10_u20_n2412 ), .ZN(_u10_u20_n3354 ) );
NAND2_X1 _u10_u20_U1263  ( .A1(_u10_u20_n3174 ), .A2(_u10_u20_n3269 ), .ZN(_u10_u20_n2375 ) );
INV_X1 _u10_u20_U1262  ( .A(_u10_u20_n2375 ), .ZN(_u10_u20_n2507 ) );
NAND2_X1 _u10_u20_U1261  ( .A1(_u10_u20_n1981 ), .A2(_u10_u20_n2507 ), .ZN(_u10_u20_n2621 ) );
NOR4_X1 _u10_u20_U1260  ( .A1(1'b0), .A2(_u10_u20_n3356 ), .A3(_u10_u20_n2203 ), .A4(_u10_u20_n2621 ), .ZN(_u10_u20_n3355 ) );
NOR4_X1 _u10_u20_U1259  ( .A1(_u10_u20_n3352 ), .A2(_u10_u20_n3353 ), .A3(_u10_u20_n3354 ), .A4(_u10_u20_n3355 ), .ZN(_u10_u20_n3306 ) );
NOR2_X1 _u10_u20_U1258  ( .A1(_u10_u20_n2842 ), .A2(_u10_u20_n2356 ), .ZN(_u10_u20_n1891 ) );
INV_X1 _u10_u20_U1257  ( .A(_u10_u20_n1869 ), .ZN(_u10_u20_n2885 ) );
NAND2_X1 _u10_u20_U1256  ( .A1(_u10_u20_n1891 ), .A2(_u10_u20_n2885 ), .ZN(_u10_u20_n3330 ) );
NAND2_X1 _u10_u20_U1255  ( .A1(_u10_u20_n2761 ), .A2(_u10_u20_n2837 ), .ZN(_u10_u20_n3351 ) );
NAND3_X1 _u10_u20_U1254  ( .A1(_u10_u20_n2884 ), .A2(_u10_u20_n2080 ), .A3(_u10_u20_n2915 ), .ZN(_u10_u20_n2762 ) );
NAND2_X1 _u10_u20_U1253  ( .A1(_u10_u20_n2055 ), .A2(_u10_u20_n2019 ), .ZN(_u10_u20_n3259 ) );
NAND4_X1 _u10_u20_U1252  ( .A1(_u10_u20_n3351 ), .A2(_u10_u20_n2762 ), .A3(_u10_u20_n2061 ), .A4(_u10_u20_n3259 ), .ZN(_u10_u20_n3350 ) );
NAND2_X1 _u10_u20_U1251  ( .A1(_u10_u20_n2183 ), .A2(_u10_u20_n3350 ), .ZN(_u10_u20_n3331 ) );
NAND2_X1 _u10_u20_U1250  ( .A1(_u10_u20_n3349 ), .A2(_u10_u20_n2305 ), .ZN(_u10_u20_n3348 ) );
NAND2_X1 _u10_u20_U1249  ( .A1(_u10_u20_n1896 ), .A2(_u10_u20_n3348 ), .ZN(_u10_u20_n3176 ) );
NAND2_X1 _u10_u20_U1248  ( .A1(_u10_u20_n2461 ), .A2(_u10_u20_n3176 ), .ZN(_u10_u20_n3332 ) );
INV_X1 _u10_u20_U1247  ( .A(_u10_u20_n2495 ), .ZN(_u10_u20_n2063 ) );
NAND2_X1 _u10_u20_U1246  ( .A1(_u10_u20_n2049 ), .A2(_u10_u20_n2063 ), .ZN(_u10_u20_n2886 ) );
NOR2_X1 _u10_u20_U1245  ( .A1(_u10_u20_n3347 ), .A2(_u10_u20_n2886 ), .ZN(_u10_u20_n3334 ) );
NAND2_X1 _u10_u20_U1244  ( .A1(1'b0), .A2(_u10_u20_n2835 ), .ZN(_u10_u20_n3344 ) );
NAND2_X1 _u10_u20_U1243  ( .A1(_u10_u20_n2001 ), .A2(_u10_u20_n2905 ), .ZN(_u10_u20_n3346 ) );
NAND2_X1 _u10_u20_U1242  ( .A1(_u10_u20_n3346 ), .A2(_u10_u20_n2803 ), .ZN(_u10_u20_n3345 ) );
NAND2_X1 _u10_u20_U1241  ( .A1(_u10_u20_n2087 ), .A2(_u10_u20_n2835 ), .ZN(_u10_u20_n2413 ) );
INV_X1 _u10_u20_U1240  ( .A(_u10_u20_n2128 ), .ZN(_u10_u20_n2235 ) );
NAND4_X1 _u10_u20_U1239  ( .A1(_u10_u20_n3344 ), .A2(_u10_u20_n3345 ), .A3(_u10_u20_n2413 ), .A4(_u10_u20_n2235 ), .ZN(_u10_u20_n3329 ) );
NOR2_X1 _u10_u20_U1238  ( .A1(_u10_u20_n1915 ), .A2(_u10_u20_n3340 ), .ZN(_u10_u20_n3343 ) );
NOR3_X1 _u10_u20_U1237  ( .A1(_u10_u20_n3329 ), .A2(1'b0), .A3(_u10_u20_n3343 ), .ZN(_u10_u20_n3341 ) );
NAND2_X1 _u10_u20_U1236  ( .A1(_u10_u20_n3342 ), .A2(_u10_u20_n3147 ), .ZN(_u10_u20_n2688 ) );
NOR2_X1 _u10_u20_U1235  ( .A1(_u10_u20_n3341 ), .A2(_u10_u20_n2688 ), .ZN(_u10_u20_n3335 ) );
NOR2_X1 _u10_u20_U1234  ( .A1(_u10_u20_n2256 ), .A2(_u10_u20_n1885 ), .ZN(_u10_u20_n2689 ) );
NOR2_X1 _u10_u20_U1233  ( .A1(1'b0), .A2(_u10_u20_n2413 ), .ZN(_u10_u20_n3338 ) );
NOR2_X1 _u10_u20_U1232  ( .A1(_u10_u20_n1925 ), .A2(_u10_u20_n3340 ), .ZN(_u10_u20_n3339 ) );
NOR3_X1 _u10_u20_U1231  ( .A1(_u10_u20_n2005 ), .A2(_u10_u20_n3338 ), .A3(_u10_u20_n3339 ), .ZN(_u10_u20_n3337 ) );
NOR2_X1 _u10_u20_U1230  ( .A1(_u10_u20_n2689 ), .A2(_u10_u20_n3337 ), .ZN(_u10_u20_n3336 ) );
NOR3_X1 _u10_u20_U1229  ( .A1(_u10_u20_n3334 ), .A2(_u10_u20_n3335 ), .A3(_u10_u20_n3336 ), .ZN(_u10_u20_n3333 ) );
NAND4_X1 _u10_u20_U1228  ( .A1(_u10_u20_n3330 ), .A2(_u10_u20_n3331 ), .A3(_u10_u20_n3332 ), .A4(_u10_u20_n3333 ), .ZN(_u10_u20_n3308 ) );
NAND3_X1 _u10_u20_U1227  ( .A1(_u10_SYNOPSYS_UNCONNECTED_8 ), .A2(_u10_SYNOPSYS_UNCONNECTED_5 ), .A3(_u10_u20_n3147 ), .ZN(_u10_u20_n2126 ) );
INV_X1 _u10_u20_U1226  ( .A(_u10_u20_n2126 ), .ZN(_u10_u20_n2329 ) );
NAND2_X1 _u10_u20_U1225  ( .A1(_u10_u20_n2329 ), .A2(_u10_u20_n3329 ), .ZN(_u10_u20_n3324 ) );
NAND2_X1 _u10_u20_U1224  ( .A1(_u10_u20_n3328 ), .A2(_u10_u20_n3136 ), .ZN(_u10_u20_n2000 ) );
INV_X1 _u10_u20_U1223  ( .A(_u10_u20_n2000 ), .ZN(_u10_u20_n2445 ) );
NAND3_X1 _u10_u20_U1222  ( .A1(_u10_u20_n2446 ), .A2(_u10_u20_n3001 ), .A3(_u10_u20_n2087 ), .ZN(_u10_u20_n3327 ) );
NAND2_X1 _u10_u20_U1221  ( .A1(_u10_u20_n3327 ), .A2(_u10_u20_n2905 ), .ZN(_u10_u20_n2500 ) );
NAND2_X1 _u10_u20_U1220  ( .A1(_u10_u20_n2445 ), .A2(_u10_u20_n2500 ), .ZN(_u10_u20_n3325 ) );
NAND2_X1 _u10_u20_U1219  ( .A1(1'b0), .A2(_u10_u20_n2979 ), .ZN(_u10_u20_n3326 ) );
NAND3_X1 _u10_u20_U1218  ( .A1(_u10_u20_n3324 ), .A2(_u10_u20_n3325 ), .A3(_u10_u20_n3326 ), .ZN(_u10_u20_n3309 ) );
AND2_X1 _u10_u20_U1217  ( .A1(_u10_u20_n2877 ), .A2(_u10_u20_n3223 ), .ZN(_u10_u20_n2858 ) );
NAND2_X1 _u10_u20_U1216  ( .A1(_u10_u20_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_6 ), .ZN(_u10_u20_n2346 ) );
INV_X1 _u10_u20_U1215  ( .A(_u10_u20_n2346 ), .ZN(_u10_u20_n2043 ) );
NAND2_X1 _u10_u20_U1214  ( .A1(_u10_u20_n2858 ), .A2(_u10_u20_n2043 ), .ZN(_u10_u20_n3321 ) );
NAND2_X1 _u10_u20_U1213  ( .A1(_u10_u20_n1982 ), .A2(_u10_u20_n2195 ), .ZN(_u10_u20_n3268 ) );
INV_X1 _u10_u20_U1212  ( .A(_u10_u20_n3268 ), .ZN(_u10_u20_n2222 ) );
NAND3_X1 _u10_u20_U1211  ( .A1(_u10_u20_n3323 ), .A2(_u10_u20_n3216 ), .A3(_u10_u20_n2222 ), .ZN(_u10_u20_n3322 ) );
NAND2_X1 _u10_u20_U1210  ( .A1(_u10_u20_n3321 ), .A2(_u10_u20_n3322 ), .ZN(_u10_u20_n2374 ) );
NAND2_X1 _u10_u20_U1209  ( .A1(_u10_u20_n3320 ), .A2(_u10_u20_n3174 ), .ZN(_u10_u20_n2014 ) );
NOR2_X1 _u10_u20_U1208  ( .A1(_u10_u20_n1841 ), .A2(_u10_u20_n2014 ), .ZN(_u10_u20_n2813 ) );
NAND2_X1 _u10_u20_U1207  ( .A1(_u10_u20_n2813 ), .A2(_u10_u20_n2534 ), .ZN(_u10_u20_n3310 ) );
NAND2_X1 _u10_u20_U1206  ( .A1(_u10_u20_n3319 ), .A2(_u10_u20_n3136 ), .ZN(_u10_u20_n1836 ) );
INV_X1 _u10_u20_U1205  ( .A(_u10_u20_n1836 ), .ZN(_u10_u20_n2815 ) );
NAND2_X1 _u10_u20_U1204  ( .A1(_u10_u20_n2534 ), .A2(_u10_u20_n3129 ), .ZN(_u10_u20_n2439 ) );
NAND2_X1 _u10_u20_U1203  ( .A1(_u10_u20_n2055 ), .A2(_u10_u20_n2107 ), .ZN(_u10_u20_n2062 ) );
NAND2_X1 _u10_u20_U1202  ( .A1(_u10_u20_n2439 ), .A2(_u10_u20_n2062 ), .ZN(_u10_u20_n3318 ) );
NAND2_X1 _u10_u20_U1201  ( .A1(_u10_u20_n2815 ), .A2(_u10_u20_n3318 ), .ZN(_u10_u20_n3311 ) );
NAND2_X1 _u10_u20_U1200  ( .A1(_u10_u20_n2986 ), .A2(_u10_u20_n2175 ), .ZN(_u10_u20_n3317 ) );
NAND2_X1 _u10_u20_U1199  ( .A1(_u10_u20_n2253 ), .A2(_u10_u20_n3317 ), .ZN(_u10_u20_n3157 ) );
NAND2_X1 _u10_u20_U1198  ( .A1(_u10_u20_n3316 ), .A2(_u10_u20_n3157 ), .ZN(_u10_u20_n3312 ) );
NOR2_X1 _u10_u20_U1197  ( .A1(_u10_u20_n2495 ), .A2(_u10_u20_n2194 ), .ZN(_u10_u20_n3314 ) );
NOR2_X1 _u10_u20_U1196  ( .A1(_u10_u20_n2375 ), .A2(_u10_u20_n2367 ), .ZN(_u10_u20_n3315 ) );
NOR2_X1 _u10_u20_U1195  ( .A1(_u10_u20_n3314 ), .A2(_u10_u20_n3315 ), .ZN(_u10_u20_n3313 ) );
NAND4_X1 _u10_u20_U1194  ( .A1(_u10_u20_n3310 ), .A2(_u10_u20_n3311 ), .A3(_u10_u20_n3312 ), .A4(_u10_u20_n3313 ), .ZN(_u10_u20_n2315 ) );
NOR4_X1 _u10_u20_U1193  ( .A1(_u10_u20_n3308 ), .A2(_u10_u20_n3309 ), .A3(_u10_u20_n2374 ), .A4(_u10_u20_n2315 ), .ZN(_u10_u20_n3307 ) );
NAND3_X1 _u10_u20_U1192  ( .A1(_u10_u20_n3305 ), .A2(_u10_u20_n3306 ), .A3(_u10_u20_n3307 ), .ZN(_u10_u20_n1987 ) );
AND2_X1 _u10_u20_U1191  ( .A1(1'b0), .A2(_u10_u20_n2977 ), .ZN(_u10_u20_n3240 ) );
NAND2_X1 _u10_u20_U1190  ( .A1(_u10_u20_n1891 ), .A2(_u10_u20_n2534 ), .ZN(_u10_u20_n3303 ) );
NAND4_X1 _u10_u20_U1189  ( .A1(_u10_u20_n1982 ), .A2(_u10_u20_n2659 ), .A3(_u10_u20_n2256 ), .A4(_u10_u20_n2175 ), .ZN(_u10_u20_n3304 ) );
AND2_X1 _u10_u20_U1188  ( .A1(_u10_u20_n3303 ), .A2(_u10_u20_n3304 ), .ZN(_u10_u20_n2612 ) );
NAND2_X1 _u10_u20_U1187  ( .A1(_u10_u20_n3302 ), .A2(_u10_u20_n3236 ), .ZN(_u10_u20_n2985 ) );
OR2_X1 _u10_u20_U1186  ( .A1(_u10_u20_n2431 ), .A2(_u10_u20_n2985 ), .ZN(_u10_u20_n3299 ) );
OR2_X1 _u10_u20_U1185  ( .A1(_u10_u20_n2282 ), .A2(_u10_u20_n2359 ), .ZN(_u10_u20_n3300 ) );
NAND2_X1 _u10_u20_U1184  ( .A1(_u10_u20_n1890 ), .A2(_u10_u20_n2534 ), .ZN(_u10_u20_n3301 ) );
NAND4_X1 _u10_u20_U1183  ( .A1(_u10_u20_n2612 ), .A2(_u10_u20_n3299 ), .A3(_u10_u20_n3300 ), .A4(_u10_u20_n3301 ), .ZN(_u10_u20_n3279 ) );
INV_X1 _u10_u20_U1182  ( .A(_u10_u20_n2464 ), .ZN(_u10_u20_n3295 ) );
NAND2_X1 _u10_u20_U1181  ( .A1(_u10_u20_n3295 ), .A2(_u10_u20_n2835 ), .ZN(_u10_u20_n2623 ) );
INV_X1 _u10_u20_U1180  ( .A(_u10_u20_n2623 ), .ZN(_u10_u20_n3185 ) );
INV_X1 _u10_u20_U1179  ( .A(_u10_u20_n2688 ), .ZN(_u10_u20_n2169 ) );
NAND2_X1 _u10_u20_U1178  ( .A1(_u10_u20_n3185 ), .A2(_u10_u20_n2169 ), .ZN(_u10_u20_n3286 ) );
NAND2_X1 _u10_u20_U1177  ( .A1(_u10_u20_n2833 ), .A2(_u10_u20_n3278 ), .ZN(_u10_u20_n3298 ) );
NAND3_X1 _u10_u20_U1176  ( .A1(_u10_u20_n3297 ), .A2(_u10_u20_n2838 ), .A3(_u10_u20_n3298 ), .ZN(_u10_u20_n3296 ) );
NAND2_X1 _u10_u20_U1175  ( .A1(_u10_u20_n2830 ), .A2(_u10_u20_n3296 ), .ZN(_u10_u20_n3287 ) );
NAND2_X1 _u10_u20_U1174  ( .A1(_u10_u20_n3295 ), .A2(_u10_u20_n3001 ), .ZN(_u10_u20_n3292 ) );
NAND2_X1 _u10_u20_U1173  ( .A1(_u10_u20_n3294 ), .A2(_u10_u20_n2089 ), .ZN(_u10_u20_n3293 ) );
AND2_X1 _u10_u20_U1172  ( .A1(_u10_u20_n3292 ), .A2(_u10_u20_n3293 ), .ZN(_u10_u20_n2548 ) );
NAND2_X1 _u10_u20_U1171  ( .A1(_u10_u20_n2548 ), .A2(_u10_u20_n2091 ), .ZN(_u10_u20_n2304 ) );
NAND2_X1 _u10_u20_U1170  ( .A1(_u10_u20_n2304 ), .A2(_u10_u20_n2446 ), .ZN(_u10_u20_n3290 ) );
NAND2_X1 _u10_u20_U1169  ( .A1(_u10_u20_n2549 ), .A2(_u10_u20_n2446 ), .ZN(_u10_u20_n2790 ) );
NOR2_X1 _u10_u20_U1168  ( .A1(_u10_u20_n1936 ), .A2(_u10_u20_n2790 ), .ZN(_u10_u20_n2789 ) );
INV_X1 _u10_u20_U1167  ( .A(_u10_u20_n2789 ), .ZN(_u10_u20_n3291 ) );
OR2_X1 _u10_u20_U1166  ( .A1(_u10_u20_n2828 ), .A2(_u10_u20_n2790 ), .ZN(_u10_u20_n2498 ) );
NAND4_X1 _u10_u20_U1165  ( .A1(_u10_u20_n3290 ), .A2(_u10_u20_n3291 ), .A3(_u10_u20_n2498 ), .A4(_u10_u20_n2001 ), .ZN(_u10_u20_n3289 ) );
NAND2_X1 _u10_u20_U1164  ( .A1(_u10_u20_n2445 ), .A2(_u10_u20_n3289 ), .ZN(_u10_u20_n3288 ) );
NAND3_X1 _u10_u20_U1163  ( .A1(_u10_u20_n3286 ), .A2(_u10_u20_n3287 ), .A3(_u10_u20_n3288 ), .ZN(_u10_u20_n3280 ) );
NOR2_X1 _u10_u20_U1162  ( .A1(_u10_u20_n2940 ), .A2(_u10_u20_n1913 ), .ZN(_u10_u20_n3281 ) );
INV_X1 _u10_u20_U1161  ( .A(1'b0), .ZN(_u10_u20_n1864 ) );
NAND2_X1 _u10_u20_U1160  ( .A1(1'b0), .A2(_u10_u20_n2588 ), .ZN(_u10_u20_n2141 ) );
INV_X1 _u10_u20_U1159  ( .A(_u10_u20_n2141 ), .ZN(_u10_u20_n3159 ) );
NAND3_X1 _u10_u20_U1158  ( .A1(_u10_u20_n2103 ), .A2(_u10_u20_n1864 ), .A3(_u10_u20_n3159 ), .ZN(_u10_u20_n2520 ) );
INV_X1 _u10_u20_U1157  ( .A(_u10_u20_n2520 ), .ZN(_u10_u20_n2630 ) );
INV_X1 _u10_u20_U1156  ( .A(_u10_u20_n2307 ), .ZN(_u10_u20_n2382 ) );
NOR4_X1 _u10_u20_U1155  ( .A1(_u10_u20_n2382 ), .A2(_u10_u20_n2722 ), .A3(_u10_u20_n1925 ), .A4(_u10_u20_n2508 ), .ZN(_u10_u20_n3260 ) );
NOR2_X1 _u10_u20_U1154  ( .A1(_u10_u20_n2498 ), .A2(_u10_u20_n2911 ), .ZN(_u10_u20_n2633 ) );
NOR2_X1 _u10_u20_U1153  ( .A1(_u10_u20_n2633 ), .A2(_u10_u20_n3278 ), .ZN(_u10_u20_n3285 ) );
INV_X1 _u10_u20_U1152  ( .A(_u10_u20_n1866 ), .ZN(_u10_u20_n1926 ) );
NOR2_X1 _u10_u20_U1151  ( .A1(_u10_u20_n3285 ), .A2(_u10_u20_n1926 ), .ZN(_u10_u20_n3284 ) );
NOR4_X1 _u10_u20_U1150  ( .A1(1'b0), .A2(_u10_u20_n2630 ), .A3(_u10_u20_n3260 ), .A4(_u10_u20_n3284 ), .ZN(_u10_u20_n3283 ) );
NOR2_X1 _u10_u20_U1149  ( .A1(_u10_u20_n3283 ), .A2(_u10_u20_n2980 ), .ZN(_u10_u20_n3282 ) );
NOR4_X1 _u10_u20_U1148  ( .A1(_u10_u20_n3279 ), .A2(_u10_u20_n3280 ), .A3(_u10_u20_n3281 ), .A4(_u10_u20_n3282 ), .ZN(_u10_u20_n3241 ) );
NAND2_X1 _u10_u20_U1147  ( .A1(_u10_u20_n1836 ), .A2(_u10_u20_n2291 ), .ZN(_u10_u20_n2147 ) );
NAND2_X1 _u10_u20_U1146  ( .A1(_u10_u20_n2443 ), .A2(_u10_u20_n2147 ), .ZN(_u10_u20_n3261 ) );
INV_X1 _u10_u20_U1145  ( .A(_u10_u20_n1841 ), .ZN(_u10_u20_n2571 ) );
NAND2_X1 _u10_u20_U1144  ( .A1(_u10_u20_n2571 ), .A2(_u10_u20_n3278 ), .ZN(_u10_u20_n3277 ) );
NAND2_X1 _u10_u20_U1143  ( .A1(_u10_u20_n3276 ), .A2(_u10_u20_n3277 ), .ZN(_u10_u20_n2819 ) );
OR2_X1 _u10_u20_U1142  ( .A1(_u10_u20_n2819 ), .A2(_u10_u20_n3275 ), .ZN(_u10_u20_n3273 ) );
NAND2_X1 _u10_u20_U1141  ( .A1(_u10_u20_n2815 ), .A2(_u10_u20_n2080 ), .ZN(_u10_u20_n3274 ) );
NAND2_X1 _u10_u20_U1140  ( .A1(_u10_u20_n2014 ), .A2(_u10_u20_n3274 ), .ZN(_u10_u20_n2165 ) );
NAND2_X1 _u10_u20_U1139  ( .A1(_u10_u20_n3273 ), .A2(_u10_u20_n2165 ), .ZN(_u10_u20_n3262 ) );
NAND2_X1 _u10_u20_U1138  ( .A1(_u10_u20_n2688 ), .A2(_u10_u20_n2126 ), .ZN(_u10_u20_n1956 ) );
INV_X1 _u10_u20_U1137  ( .A(_u10_u20_n1956 ), .ZN(_u10_u20_n1860 ) );
NOR2_X1 _u10_u20_U1136  ( .A1(1'b0), .A2(_u10_u20_n2498 ), .ZN(_u10_u20_n3271 ) );
NOR2_X1 _u10_u20_U1135  ( .A1(_u10_u20_n3271 ), .A2(_u10_u20_n3272 ), .ZN(_u10_u20_n3270 ) );
NOR2_X1 _u10_u20_U1134  ( .A1(_u10_u20_n1860 ), .A2(_u10_u20_n3270 ), .ZN(_u10_u20_n3264 ) );
INV_X1 _u10_u20_U1133  ( .A(_u10_u20_n2632 ), .ZN(_u10_u20_n3202 ) );
NAND2_X1 _u10_u20_U1132  ( .A1(_u10_u20_n3236 ), .A2(_u10_u20_n3269 ), .ZN(_u10_u20_n3036 ) );
INV_X1 _u10_u20_U1131  ( .A(_u10_u20_n3036 ), .ZN(_u10_u20_n1960 ) );
NAND2_X1 _u10_u20_U1130  ( .A1(_u10_u20_n3202 ), .A2(_u10_u20_n1960 ), .ZN(_u10_u20_n3079 ) );
NOR3_X1 _u10_u20_U1129  ( .A1(_u10_u20_n3079 ), .A2(1'b0), .A3(_u10_u20_n3268 ), .ZN(_u10_u20_n3265 ) );
INV_X1 _u10_u20_U1128  ( .A(_u10_u20_n2014 ), .ZN(_u10_u20_n2709 ) );
NAND2_X1 _u10_u20_U1127  ( .A1(_u10_u20_n2709 ), .A2(_u10_u20_n2166 ), .ZN(_u10_u20_n2145 ) );
INV_X1 _u10_u20_U1126  ( .A(_u10_u20_n2145 ), .ZN(_u10_u20_n3258 ) );
NOR2_X1 _u10_u20_U1125  ( .A1(_u10_u20_n3258 ), .A2(_u10_u20_n2183 ), .ZN(_u10_u20_n3267 ) );
NOR2_X1 _u10_u20_U1124  ( .A1(_u10_u20_n3267 ), .A2(_u10_u20_n2567 ), .ZN(_u10_u20_n3266 ) );
NOR3_X1 _u10_u20_U1123  ( .A1(_u10_u20_n3264 ), .A2(_u10_u20_n3265 ), .A3(_u10_u20_n3266 ), .ZN(_u10_u20_n3263 ) );
NAND3_X1 _u10_u20_U1122  ( .A1(_u10_u20_n3261 ), .A2(_u10_u20_n3262 ), .A3(_u10_u20_n3263 ), .ZN(_u10_u20_n3243 ) );
INV_X1 _u10_u20_U1121  ( .A(_u10_u20_n2102 ), .ZN(_u10_u20_n2509 ) );
NAND2_X1 _u10_u20_U1120  ( .A1(_u10_u20_n3260 ), .A2(_u10_u20_n2509 ), .ZN(_u10_u20_n3247 ) );
INV_X1 _u10_u20_U1119  ( .A(_u10_u20_n3259 ), .ZN(_u10_u20_n2015 ) );
NAND2_X1 _u10_u20_U1118  ( .A1(_u10_u20_n2015 ), .A2(_u10_u20_n3258 ), .ZN(_u10_u20_n3248 ) );
NAND2_X1 _u10_u20_U1117  ( .A1(_u10_u20_n2251 ), .A2(_u10_u20_n2169 ), .ZN(_u10_u20_n3255 ) );
OR2_X1 _u10_u20_U1116  ( .A1(_u10_u20_n3157 ), .A2(_u10_u20_n2256 ), .ZN(_u10_u20_n3257 ) );
NAND2_X1 _u10_u20_U1115  ( .A1(_u10_u20_n2105 ), .A2(_u10_u20_n3257 ), .ZN(_u10_u20_n3256 ) );
AND2_X1 _u10_u20_U1114  ( .A1(_u10_u20_n3255 ), .A2(_u10_u20_n3256 ), .ZN(_u10_u20_n3212 ) );
INV_X1 _u10_u20_U1113  ( .A(_u10_u20_n2037 ), .ZN(_u10_u20_n2987 ) );
NAND2_X1 _u10_u20_U1112  ( .A1(_u10_u20_n2987 ), .A2(_u10_u20_n2038 ), .ZN(_u10_u20_n2212 ) );
NOR2_X1 _u10_u20_U1111  ( .A1(_u10_u20_n2212 ), .A2(1'b0), .ZN(_u10_u20_n2658 ) );
INV_X1 _u10_u20_U1110  ( .A(_u10_u20_n2658 ), .ZN(_u10_u20_n2343 ) );
NAND2_X1 _u10_u20_U1109  ( .A1(_u10_u20_n2344 ), .A2(_u10_u20_n3254 ), .ZN(_u10_u20_n1928 ) );
NAND2_X1 _u10_u20_U1108  ( .A1(_u10_u20_n2588 ), .A2(_u10_u20_n1928 ), .ZN(_u10_u20_n3253 ) );
NAND2_X1 _u10_u20_U1107  ( .A1(_u10_u20_n2343 ), .A2(_u10_u20_n3253 ), .ZN(_u10_u20_n3252 ) );
NAND2_X1 _u10_u20_U1106  ( .A1(_u10_u20_n2105 ), .A2(_u10_u20_n3252 ), .ZN(_u10_u20_n3251 ) );
NAND2_X1 _u10_u20_U1105  ( .A1(_u10_u20_n3212 ), .A2(_u10_u20_n3251 ), .ZN(_u10_u20_n3250 ) );
NAND2_X1 _u10_u20_U1104  ( .A1(_u10_u20_n2307 ), .A2(_u10_u20_n3250 ), .ZN(_u10_u20_n3249 ) );
NAND3_X1 _u10_u20_U1103  ( .A1(_u10_u20_n3247 ), .A2(_u10_u20_n3248 ), .A3(_u10_u20_n3249 ), .ZN(_u10_u20_n3244 ) );
AND2_X1 _u10_u20_U1102  ( .A1(_u10_u20_n2915 ), .A2(_u10_u20_n2059 ), .ZN(_u10_u20_n2957 ) );
AND3_X1 _u10_u20_U1101  ( .A1(_u10_u20_n3223 ), .A2(_u10_u20_n2837 ), .A3(_u10_u20_n2957 ), .ZN(_u10_u20_n2051 ) );
NOR2_X1 _u10_u20_U1100  ( .A1(_u10_u20_n2528 ), .A2(_u10_u20_n2051 ), .ZN(_u10_u20_n2605 ) );
NOR2_X1 _u10_u20_U1099  ( .A1(_u10_u20_n2605 ), .A2(_u10_u20_n2346 ), .ZN(_u10_u20_n3245 ) );
NOR2_X1 _u10_u20_U1098  ( .A1(_u10_u20_n2291 ), .A2(_u10_u20_n2062 ), .ZN(_u10_u20_n3246 ) );
NOR4_X1 _u10_u20_U1097  ( .A1(_u10_u20_n3243 ), .A2(_u10_u20_n3244 ), .A3(_u10_u20_n3245 ), .A4(_u10_u20_n3246 ), .ZN(_u10_u20_n3242 ) );
NAND2_X1 _u10_u20_U1096  ( .A1(_u10_u20_n3241 ), .A2(_u10_u20_n3242 ), .ZN(_u10_u20_n2311 ) );
OR3_X1 _u10_u20_U1095  ( .A1(_u10_u20_n1987 ), .A2(_u10_u20_n3240 ), .A3(_u10_u20_n2311 ), .ZN(_u10_u20_n3192 ) );
INV_X1 _u10_u20_U1094  ( .A(_u10_u20_n2886 ), .ZN(_u10_u20_n2720 ) );
NOR2_X1 _u10_u20_U1093  ( .A1(_u10_u20_n2004 ), .A2(_u10_u20_n2720 ), .ZN(_u10_u20_n2455 ) );
INV_X1 _u10_u20_U1092  ( .A(_u10_u20_n2488 ), .ZN(_u10_u20_n2938 ) );
AND3_X1 _u10_u20_U1091  ( .A1(_u10_u20_n2455 ), .A2(_u10_u20_n1859 ), .A3(_u10_u20_n2938 ), .ZN(_u10_u20_n3239 ) );
INV_X1 _u10_u20_U1090  ( .A(_u10_u20_n2633 ), .ZN(_u10_u20_n2937 ) );
NOR2_X1 _u10_u20_U1089  ( .A1(_u10_u20_n3239 ), .A2(_u10_u20_n2937 ), .ZN(_u10_u20_n3227 ) );
NOR2_X1 _u10_u20_U1088  ( .A1(_u10_u20_n1976 ), .A2(_u10_u20_n1969 ), .ZN(_u10_u20_n3237 ) );
NOR2_X1 _u10_u20_U1087  ( .A1(1'b0), .A2(_u10_u20_n2947 ), .ZN(_u10_u20_n3238 ) );
NOR3_X1 _u10_u20_U1086  ( .A1(_u10_u20_n2476 ), .A2(_u10_u20_n3237 ), .A3(_u10_u20_n3238 ), .ZN(_u10_u20_n3235 ) );
NOR3_X1 _u10_u20_U1085  ( .A1(_u10_u20_n1813 ), .A2(_u10_u20_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_5 ), .ZN(_u10_u20_n3135 ) );
NAND2_X1 _u10_u20_U1084  ( .A1(_u10_u20_n3135 ), .A2(_u10_u20_n3236 ), .ZN(_u10_u20_n2573 ) );
NOR2_X1 _u10_u20_U1083  ( .A1(_u10_u20_n3235 ), .A2(_u10_u20_n2573 ), .ZN(_u10_u20_n3228 ) );
NOR2_X1 _u10_u20_U1082  ( .A1(_u10_u20_n2216 ), .A2(_u10_u20_n1868 ), .ZN(_u10_u20_n3233 ) );
INV_X1 _u10_u20_U1081  ( .A(_u10_u20_n2550 ), .ZN(_u10_u20_n2475 ) );
NOR3_X1 _u10_u20_U1080  ( .A1(_u10_u20_n2475 ), .A2(1'b0), .A3(_u10_u20_n1925 ), .ZN(_u10_u20_n3234 ) );
NOR3_X1 _u10_u20_U1079  ( .A1(_u10_u20_n3233 ), .A2(1'b0), .A3(_u10_u20_n3234 ), .ZN(_u10_u20_n3232 ) );
NOR2_X1 _u10_u20_U1078  ( .A1(_u10_u20_n3232 ), .A2(_u10_u20_n2037 ), .ZN(_u10_u20_n3229 ) );
NOR2_X1 _u10_u20_U1077  ( .A1(_u10_u20_n3231 ), .A2(_u10_u20_n2365 ), .ZN(_u10_u20_n3230 ) );
NOR4_X1 _u10_u20_U1076  ( .A1(_u10_u20_n3227 ), .A2(_u10_u20_n3228 ), .A3(_u10_u20_n3229 ), .A4(_u10_u20_n3230 ), .ZN(_u10_u20_n3205 ) );
NOR3_X1 _u10_u20_U1075  ( .A1(_u10_u20_n3226 ), .A2(_u10_u20_n2687 ), .A3(_u10_u20_n2145 ), .ZN(_u10_u20_n3217 ) );
NOR3_X1 _u10_u20_U1074  ( .A1(_u10_u20_n3225 ), .A2(1'b0), .A3(_u10_u20_n2587 ), .ZN(_u10_u20_n3218 ) );
NOR2_X1 _u10_u20_U1073  ( .A1(_u10_u20_n3159 ), .A2(1'b0), .ZN(_u10_u20_n3224 ) );
NOR2_X1 _u10_u20_U1072  ( .A1(_u10_u20_n3224 ), .A2(_u10_u20_n2584 ), .ZN(_u10_u20_n3219 ) );
NAND2_X1 _u10_u20_U1071  ( .A1(_u10_u20_n3222 ), .A2(_u10_u20_n3223 ), .ZN(_u10_u20_n2048 ) );
INV_X1 _u10_u20_U1070  ( .A(_u10_u20_n2048 ), .ZN(_u10_u20_n2859 ) );
NOR2_X1 _u10_u20_U1069  ( .A1(_u10_u20_n2859 ), .A2(_u10_u20_n2054 ), .ZN(_u10_u20_n3221 ) );
NOR2_X1 _u10_u20_U1068  ( .A1(_u10_u20_n3221 ), .A2(_u10_u20_n2346 ), .ZN(_u10_u20_n3220 ) );
NOR4_X1 _u10_u20_U1067  ( .A1(_u10_u20_n3217 ), .A2(_u10_u20_n3218 ), .A3(_u10_u20_n3219 ), .A4(_u10_u20_n3220 ), .ZN(_u10_u20_n3206 ) );
NAND2_X1 _u10_u20_U1066  ( .A1(_u10_u20_n2377 ), .A2(_u10_u20_n2721 ), .ZN(_u10_u20_n3213 ) );
AND4_X1 _u10_u20_U1065  ( .A1(1'b0), .A2(_u10_u20_n2502 ), .A3(_u10_u20_n2972 ), .A4(_u10_u20_n3040 ), .ZN(_u10_u20_n2406 ) );
NAND2_X1 _u10_u20_U1064  ( .A1(_u10_u20_n2406 ), .A2(_u10_u20_n2979 ), .ZN(_u10_u20_n3214 ) );
NAND2_X1 _u10_u20_U1063  ( .A1(_u10_u20_n2630 ), .A2(_u10_u20_n3216 ), .ZN(_u10_u20_n2376 ) );
INV_X1 _u10_u20_U1062  ( .A(_u10_u20_n2376 ), .ZN(_u10_u20_n3108 ) );
NAND2_X1 _u10_u20_U1061  ( .A1(_u10_u20_n3108 ), .A2(_u10_u20_n2507 ), .ZN(_u10_u20_n3215 ) );
NOR2_X1 _u10_u20_U1060  ( .A1(_u10_u20_n2937 ), .A2(1'b0), .ZN(_u10_u20_n2649 ) );
INV_X1 _u10_u20_U1059  ( .A(_u10_u20_n2253 ), .ZN(_u10_u20_n2971 ) );
NAND2_X1 _u10_u20_U1058  ( .A1(_u10_u20_n2649 ), .A2(_u10_u20_n2971 ), .ZN(_u10_u20_n2918 ) );
NAND4_X1 _u10_u20_U1057  ( .A1(_u10_u20_n3213 ), .A2(_u10_u20_n3214 ), .A3(_u10_u20_n3215 ), .A4(_u10_u20_n2918 ), .ZN(_u10_u20_n3208 ) );
NOR2_X1 _u10_u20_U1056  ( .A1(_u10_u20_n2000 ), .A2(_u10_u20_n2902 ), .ZN(_u10_u20_n3209 ) );
NOR2_X1 _u10_u20_U1055  ( .A1(_u10_u20_n3212 ), .A2(_u10_u20_n2475 ), .ZN(_u10_u20_n3210 ) );
INV_X1 _u10_u20_U1054  ( .A(_u10_u20_n2441 ), .ZN(_u10_u20_n3128 ) );
NOR2_X1 _u10_u20_U1053  ( .A1(_u10_u20_n2356 ), .A2(_u10_u20_n3128 ), .ZN(_u10_u20_n3211 ) );
NOR4_X1 _u10_u20_U1052  ( .A1(_u10_u20_n3208 ), .A2(_u10_u20_n3209 ), .A3(_u10_u20_n3210 ), .A4(_u10_u20_n3211 ), .ZN(_u10_u20_n3207 ) );
NAND3_X1 _u10_u20_U1051  ( .A1(_u10_u20_n3205 ), .A2(_u10_u20_n3206 ), .A3(_u10_u20_n3207 ), .ZN(_u10_u20_n2611 ) );
NOR2_X1 _u10_u20_U1050  ( .A1(_u10_u20_n2212 ), .A2(_u10_u20_n2216 ), .ZN(_u10_u20_n1937 ) );
NOR2_X1 _u10_u20_U1049  ( .A1(_u10_u20_n2533 ), .A2(_u10_u20_n2214 ), .ZN(_u10_u20_n2765 ) );
INV_X1 _u10_u20_U1048  ( .A(_u10_u20_n2005 ), .ZN(_u10_u20_n2111 ) );
AND2_X1 _u10_u20_U1047  ( .A1(_u10_u20_n2765 ), .A2(_u10_u20_n2111 ), .ZN(_u10_u20_n3201 ) );
INV_X1 _u10_u20_U1046  ( .A(_u10_u20_n3059 ), .ZN(_u10_u20_n3076 ) );
NAND2_X1 _u10_u20_U1045  ( .A1(_u10_u20_n3201 ), .A2(_u10_u20_n3076 ), .ZN(_u10_u20_n3204 ) );
NAND2_X1 _u10_u20_U1044  ( .A1(_u10_u20_n1937 ), .A2(_u10_u20_n3204 ), .ZN(_u10_u20_n3193 ) );
NAND2_X1 _u10_u20_U1043  ( .A1(_u10_u20_n2254 ), .A2(_u10_u20_n2212 ), .ZN(_u10_u20_n3203 ) );
NAND3_X1 _u10_u20_U1042  ( .A1(_u10_u20_n3203 ), .A2(_u10_u20_n2175 ), .A3(_u10_u20_n2649 ), .ZN(_u10_u20_n3194 ) );
NOR2_X1 _u10_u20_U1041  ( .A1(_u10_u20_n2985 ), .A2(1'b0), .ZN(_u10_u20_n1959 ) );
NAND2_X1 _u10_u20_U1040  ( .A1(_u10_u20_n1959 ), .A2(_u10_u20_n3202 ), .ZN(_u10_u20_n2202 ) );
NAND4_X1 _u10_u20_U1039  ( .A1(_u10_u20_n3079 ), .A2(_u10_u20_n2621 ), .A3(_u10_u20_n2202 ), .A4(_u10_u20_n2798 ), .ZN(_u10_u20_n3200 ) );
NAND2_X1 _u10_u20_U1038  ( .A1(_u10_u20_n3201 ), .A2(_u10_u20_n2937 ), .ZN(_u10_u20_n2772 ) );
NAND2_X1 _u10_u20_U1037  ( .A1(_u10_u20_n3200 ), .A2(_u10_u20_n2772 ), .ZN(_u10_u20_n3195 ) );
NAND2_X1 _u10_u20_U1036  ( .A1(_u10_u20_n2765 ), .A2(_u10_u20_n1869 ), .ZN(_u10_u20_n3199 ) );
NAND2_X1 _u10_u20_U1035  ( .A1(_u10_u20_n2049 ), .A2(_u10_u20_n3199 ), .ZN(_u10_u20_n3057 ) );
NOR2_X1 _u10_u20_U1034  ( .A1(_u10_u20_n2495 ), .A2(_u10_u20_n3057 ), .ZN(_u10_u20_n3197 ) );
NOR2_X1 _u10_u20_U1033  ( .A1(_u10_u20_n2883 ), .A2(_u10_u20_n2485 ), .ZN(_u10_u20_n3198 ) );
NOR2_X1 _u10_u20_U1032  ( .A1(_u10_u20_n3197 ), .A2(_u10_u20_n3198 ), .ZN(_u10_u20_n3196 ) );
NAND4_X1 _u10_u20_U1031  ( .A1(_u10_u20_n3193 ), .A2(_u10_u20_n3194 ), .A3(_u10_u20_n3195 ), .A4(_u10_u20_n3196 ), .ZN(_u10_u20_n2887 ) );
NOR4_X1 _u10_u20_U1030  ( .A1(_u10_u20_n3191 ), .A2(_u10_u20_n3192 ), .A3(_u10_u20_n2611 ), .A4(_u10_u20_n2887 ), .ZN(_u10_u20_n3015 ) );
NAND3_X1 _u10_u20_U1029  ( .A1(_u10_u20_n3190 ), .A2(_u10_u20_n2049 ), .A3(_u10_u20_n2957 ), .ZN(_u10_u20_n2699 ) );
OR2_X1 _u10_u20_U1028  ( .A1(_u10_u20_n2699 ), .A2(_u10_u20_n1813 ), .ZN(_u10_u20_n3187 ) );
NAND3_X1 _u10_u20_U1027  ( .A1(_u10_u20_n2978 ), .A2(_u10_u20_n2405 ), .A3(1'b0), .ZN(_u10_u20_n3188 ) );
NAND4_X1 _u10_u20_U1026  ( .A1(_u10_u20_n3058 ), .A2(_u10_u20_n3187 ), .A3(_u10_u20_n3188 ), .A4(_u10_u20_n3189 ), .ZN(_u10_u20_n3186 ) );
NAND2_X1 _u10_u20_U1025  ( .A1(_u10_u20_n2063 ), .A2(_u10_u20_n3186 ), .ZN(_u10_u20_n3163 ) );
NAND2_X1 _u10_u20_U1024  ( .A1(_u10_u20_n3185 ), .A2(_u10_u20_n2329 ), .ZN(_u10_u20_n3164 ) );
NAND2_X1 _u10_u20_U1023  ( .A1(_u10_u20_n2689 ), .A2(_u10_u20_n2365 ), .ZN(_u10_u20_n2736 ) );
NOR2_X1 _u10_u20_U1022  ( .A1(_u10_u20_n2736 ), .A2(_u10_u20_n2488 ), .ZN(_u10_u20_n1855 ) );
INV_X1 _u10_u20_U1021  ( .A(_u10_u20_n1855 ), .ZN(_u10_u20_n3184 ) );
NOR2_X1 _u10_u20_U1020  ( .A1(_u10_u20_n2274 ), .A2(_u10_u20_n2359 ), .ZN(_u10_u20_n2952 ) );
NOR2_X1 _u10_u20_U1019  ( .A1(_u10_u20_n3184 ), .A2(_u10_u20_n2952 ), .ZN(_u10_u20_n2776 ) );
OR2_X1 _u10_u20_U1018  ( .A1(_u10_u20_n2852 ), .A2(_u10_u20_n2776 ), .ZN(_u10_u20_n3165 ) );
NAND2_X1 _u10_u20_U1017  ( .A1(_u10_u20_n3126 ), .A2(_u10_u20_n2915 ), .ZN(_u10_u20_n3065 ) );
NOR3_X1 _u10_u20_U1016  ( .A1(_u10_u20_n3065 ), .A2(1'b0), .A3(_u10_u20_n2632 ), .ZN(_u10_u20_n3182 ) );
NOR3_X1 _u10_u20_U1015  ( .A1(_u10_u20_n3182 ), .A2(_u10_u20_n3183 ), .A3(_u10_u20_n3108 ), .ZN(_u10_u20_n3181 ) );
NOR2_X1 _u10_u20_U1014  ( .A1(_u10_u20_n3181 ), .A2(_u10_u20_n3162 ), .ZN(_u10_u20_n3167 ) );
INV_X1 _u10_u20_U1013  ( .A(_u10_u20_n3180 ), .ZN(_u10_u20_n3140 ) );
NAND3_X1 _u10_u20_U1012  ( .A1(_u10_u20_n3140 ), .A2(_u10_u20_n2163 ), .A3(_u10_u20_n2092 ), .ZN(_u10_u20_n3175 ) );
NOR4_X1 _u10_u20_U1011  ( .A1(_u10_u20_n2411 ), .A2(_u10_u20_n2710 ), .A3(_u10_u20_n3141 ), .A4(_u10_u20_n3089 ), .ZN(_u10_u20_n3179 ) );
NOR2_X1 _u10_u20_U1010  ( .A1(1'b0), .A2(_u10_u20_n3179 ), .ZN(_u10_u20_n3177 ) );
NOR2_X1 _u10_u20_U1009  ( .A1(_u10_u20_n1898 ), .A2(_u10_u20_n1847 ), .ZN(_u10_u20_n3178 ) );
NOR4_X1 _u10_u20_U1008  ( .A1(_u10_u20_n3175 ), .A2(_u10_u20_n3176 ), .A3(_u10_u20_n3177 ), .A4(_u10_u20_n3178 ), .ZN(_u10_u20_n3173 ) );
NAND2_X1 _u10_u20_U1007  ( .A1(_u10_u20_n3135 ), .A2(_u10_u20_n3174 ), .ZN(_u10_u20_n2159 ) );
NOR2_X1 _u10_u20_U1006  ( .A1(_u10_u20_n3173 ), .A2(_u10_u20_n2159 ), .ZN(_u10_u20_n3168 ) );
OR3_X1 _u10_u20_U1005  ( .A1(_u10_u20_n3172 ), .A2(1'b0), .A3(_u10_u20_n3126 ), .ZN(_u10_u20_n3171 ) );
NAND2_X1 _u10_u20_U1004  ( .A1(_u10_u20_n2600 ), .A2(_u10_u20_n3171 ), .ZN(_u10_u20_n3153 ) );
AND3_X1 _u10_u20_U1003  ( .A1(_u10_u20_n3153 ), .A2(_u10_u20_n2947 ), .A3(_u10_u20_n2579 ), .ZN(_u10_u20_n3170 ) );
NOR2_X1 _u10_u20_U1002  ( .A1(_u10_u20_n3170 ), .A2(_u10_u20_n2359 ), .ZN(_u10_u20_n3169 ) );
NOR3_X1 _u10_u20_U1001  ( .A1(_u10_u20_n3167 ), .A2(_u10_u20_n3168 ), .A3(_u10_u20_n3169 ), .ZN(_u10_u20_n3166 ) );
NAND4_X1 _u10_u20_U1000  ( .A1(_u10_u20_n3163 ), .A2(_u10_u20_n3164 ), .A3(_u10_u20_n3165 ), .A4(_u10_u20_n3166 ), .ZN(_u10_u20_n3130 ) );
NAND2_X1 _u10_u20_U999  ( .A1(_u10_u20_n2375 ), .A2(_u10_u20_n3162 ), .ZN(_u10_u20_n1923 ) );
NAND2_X1 _u10_u20_U998  ( .A1(_u10_u20_n3062 ), .A2(_u10_u20_n1923 ), .ZN(_u10_u20_n3154 ) );
NAND2_X1 _u10_u20_U997  ( .A1(_u10_u20_n2103 ), .A2(_u10_u20_n2509 ), .ZN(_u10_u20_n3161 ) );
NAND2_X1 _u10_u20_U996  ( .A1(_u10_u20_n2344 ), .A2(_u10_u20_n3161 ), .ZN(_u10_u20_n3160 ) );
NAND2_X1 _u10_u20_U995  ( .A1(_u10_u20_n3159 ), .A2(_u10_u20_n3160 ), .ZN(_u10_u20_n2635 ) );
AND3_X1 _u10_u20_U994  ( .A1(_u10_u20_n2549 ), .A2(_u10_u20_n2108 ), .A3(_u10_u20_n3126 ), .ZN(_u10_u20_n3093 ) );
NAND2_X1 _u10_u20_U993  ( .A1(_u10_u20_n3093 ), .A2(_u10_u20_n2941 ), .ZN(_u10_u20_n3158 ) );
NAND3_X1 _u10_u20_U992  ( .A1(_u10_u20_n3076 ), .A2(_u10_u20_n3066 ), .A3(_u10_u20_n3158 ), .ZN(_u10_u20_n3156 ) );
NAND2_X1 _u10_u20_U991  ( .A1(_u10_u20_n3156 ), .A2(_u10_u20_n3157 ), .ZN(_u10_u20_n3155 ) );
NAND3_X1 _u10_u20_U990  ( .A1(_u10_u20_n3154 ), .A2(_u10_u20_n2635 ), .A3(_u10_u20_n3155 ), .ZN(_u10_u20_n3131 ) );
INV_X1 _u10_u20_U989  ( .A(_u10_u20_n2594 ), .ZN(_u10_u20_n2846 ) );
NAND3_X1 _u10_u20_U988  ( .A1(_u10_u20_n2162 ), .A2(_u10_u20_n2082 ), .A3(_u10_u20_n2105 ), .ZN(_u10_u20_n2077 ) );
NAND4_X1 _u10_u20_U987  ( .A1(_u10_u20_n3153 ), .A2(_u10_u20_n1969 ), .A3(_u10_u20_n2846 ), .A4(_u10_u20_n2077 ), .ZN(_u10_u20_n3148 ) );
NAND2_X1 _u10_u20_U986  ( .A1(_u10_u20_n2838 ), .A2(_u10_u20_n3128 ), .ZN(_u10_u20_n3152 ) );
NAND2_X1 _u10_u20_U985  ( .A1(_u10_u20_n3152 ), .A2(_u10_u20_n2600 ), .ZN(_u10_u20_n3151 ) );
NAND2_X1 _u10_u20_U984  ( .A1(_u10_u20_n2282 ), .A2(_u10_u20_n3151 ), .ZN(_u10_u20_n2601 ) );
NOR4_X1 _u10_u20_U983  ( .A1(_u10_u20_n2885 ), .A2(_u10_u20_n2534 ), .A3(_u10_u20_n2214 ), .A4(_u10_u20_n3059 ), .ZN(_u10_u20_n3150 ) );
NOR2_X1 _u10_u20_U982  ( .A1(_u10_u20_n3150 ), .A2(_u10_u20_n2853 ), .ZN(_u10_u20_n3149 ) );
NOR4_X1 _u10_u20_U981  ( .A1(_u10_u20_n3148 ), .A2(_u10_u20_n2601 ), .A3(_u10_u20_n3149 ), .A4(_u10_u20_n1975 ), .ZN(_u10_u20_n3146 ) );
NAND3_X1 _u10_u20_U980  ( .A1(_u10_SYNOPSYS_UNCONNECTED_8 ), .A2(_u10_SYNOPSYS_UNCONNECTED_4 ), .A3(_u10_u20_n3147 ), .ZN(_u10_u20_n2071 ) );
NOR2_X1 _u10_u20_U979  ( .A1(_u10_u20_n3146 ), .A2(_u10_u20_n2071 ), .ZN(_u10_u20_n3132 ) );
NOR2_X1 _u10_u20_U978  ( .A1(1'b0), .A2(_u10_u20_n1847 ), .ZN(_u10_u20_n3143 ) );
INV_X1 _u10_u20_U977  ( .A(_u10_u20_n3145 ), .ZN(_u10_u20_n3144 ) );
NOR2_X1 _u10_u20_U976  ( .A1(_u10_u20_n3143 ), .A2(_u10_u20_n3144 ), .ZN(_u10_u20_n3142 ) );
NOR2_X1 _u10_u20_U975  ( .A1(1'b0), .A2(_u10_u20_n3142 ), .ZN(_u10_u20_n3137 ) );
NAND2_X1 _u10_u20_U974  ( .A1(_u10_u20_n2549 ), .A2(_u10_u20_n3141 ), .ZN(_u10_u20_n3138 ) );
NAND2_X1 _u10_u20_U973  ( .A1(_u10_u20_n1896 ), .A2(_u10_u20_n3140 ), .ZN(_u10_u20_n2544 ) );
NAND2_X1 _u10_u20_U972  ( .A1(_u10_u20_n2089 ), .A2(_u10_u20_n2544 ), .ZN(_u10_u20_n3139 ) );
NAND2_X1 _u10_u20_U971  ( .A1(_u10_u20_n3138 ), .A2(_u10_u20_n3139 ), .ZN(_u10_u20_n2795 ) );
NOR4_X1 _u10_u20_U970  ( .A1(_u10_u20_n2300 ), .A2(_u10_u20_n3137 ), .A3(_u10_u20_n2304 ), .A4(_u10_u20_n2795 ), .ZN(_u10_u20_n3134 ) );
NAND2_X1 _u10_u20_U969  ( .A1(_u10_u20_n3135 ), .A2(_u10_u20_n3136 ), .ZN(_u10_u20_n2085 ) );
NOR2_X1 _u10_u20_U968  ( .A1(_u10_u20_n3134 ), .A2(_u10_u20_n2085 ), .ZN(_u10_u20_n3133 ) );
NOR4_X1 _u10_u20_U967  ( .A1(_u10_u20_n3130 ), .A2(_u10_u20_n3131 ), .A3(_u10_u20_n3132 ), .A4(_u10_u20_n3133 ), .ZN(_u10_u20_n3016 ) );
INV_X1 _u10_u20_U966  ( .A(_u10_u20_n2686 ), .ZN(_u10_u20_n2278 ) );
NAND4_X1 _u10_u20_U965  ( .A1(_u10_u20_n2105 ), .A2(_u10_u20_n2278 ), .A3(_u10_u20_n3129 ), .A4(_u10_u20_n2600 ), .ZN(_u10_u20_n2437 ) );
NAND2_X1 _u10_u20_U964  ( .A1(_u10_u20_n3128 ), .A2(_u10_u20_n2437 ), .ZN(_u10_u20_n3127 ) );
NAND2_X1 _u10_u20_U963  ( .A1(_u10_u20_n2815 ), .A2(_u10_u20_n3127 ), .ZN(_u10_u20_n3098 ) );
INV_X1 _u10_u20_U962  ( .A(_u10_u20_n2573 ), .ZN(_u10_u20_n1967 ) );
NAND2_X1 _u10_u20_U961  ( .A1(_u10_u20_n3126 ), .A2(_u10_u20_n2078 ), .ZN(_u10_u20_n3123 ) );
NAND2_X1 _u10_u20_U960  ( .A1(_u10_u20_n3076 ), .A2(_u10_u20_n1925 ), .ZN(_u10_u20_n3125 ) );
NAND2_X1 _u10_u20_U959  ( .A1(_u10_u20_n2669 ), .A2(_u10_u20_n3125 ), .ZN(_u10_u20_n3124 ) );
NAND4_X1 _u10_u20_U958  ( .A1(_u10_u20_n3122 ), .A2(_u10_u20_n3123 ), .A3(_u10_u20_n3124 ), .A4(_u10_u20_n2579 ), .ZN(_u10_u20_n3121 ) );
NAND2_X1 _u10_u20_U957  ( .A1(_u10_u20_n3121 ), .A2(_u10_u20_n2874 ), .ZN(_u10_u20_n3120 ) );
NAND2_X1 _u10_u20_U956  ( .A1(_u10_u20_n2382 ), .A2(_u10_u20_n3120 ), .ZN(_u10_u20_n3119 ) );
NAND2_X1 _u10_u20_U955  ( .A1(_u10_u20_n1967 ), .A2(_u10_u20_n3119 ), .ZN(_u10_u20_n3099 ) );
NAND2_X1 _u10_u20_U954  ( .A1(_u10_u20_n3118 ), .A2(_u10_u20_n3001 ), .ZN(_u10_u20_n3117 ) );
NAND2_X1 _u10_u20_U953  ( .A1(_u10_u20_n2446 ), .A2(_u10_u20_n3117 ), .ZN(_u10_u20_n3116 ) );
NAND2_X1 _u10_u20_U952  ( .A1(_u10_u20_n2445 ), .A2(_u10_u20_n3116 ), .ZN(_u10_u20_n3100 ) );
OR2_X1 _u10_u20_U951  ( .A1(_u10_u20_n3115 ), .A2(_u10_u20_n2687 ), .ZN(_u10_u20_n3114 ) );
AND3_X1 _u10_u20_U950  ( .A1(_u10_u20_n2061 ), .A2(_u10_u20_n2166 ), .A3(_u10_u20_n3114 ), .ZN(_u10_u20_n3045 ) );
NOR2_X1 _u10_u20_U949  ( .A1(1'b0), .A2(_u10_u20_n3045 ), .ZN(_u10_u20_n3113 ) );
NOR2_X1 _u10_u20_U948  ( .A1(_u10_u20_n3113 ), .A2(1'b0), .ZN(_u10_u20_n3112 ) );
NOR2_X1 _u10_u20_U947  ( .A1(_u10_u20_n3112 ), .A2(_u10_u20_n2356 ), .ZN(_u10_u20_n3102 ) );
NAND2_X1 _u10_u20_U946  ( .A1(_u10_u20_n2571 ), .A2(_u10_u20_n2165 ), .ZN(_u10_u20_n3078 ) );
NAND2_X1 _u10_u20_U945  ( .A1(_u10_u20_n2365 ), .A2(_u10_u20_n3078 ), .ZN(_u10_u20_n2241 ) );
NOR2_X1 _u10_u20_U944  ( .A1(_u10_u20_n2377 ), .A2(_u10_u20_n2241 ), .ZN(_u10_u20_n3111 ) );
NOR2_X1 _u10_u20_U943  ( .A1(_u10_u20_n3111 ), .A2(_u10_u20_n1869 ), .ZN(_u10_u20_n3103 ) );
NOR2_X1 _u10_u20_U942  ( .A1(_u10_u20_n2999 ), .A2(_u10_u20_n2977 ), .ZN(_u10_u20_n3061 ) );
NOR2_X1 _u10_u20_U941  ( .A1(_u10_u20_n3061 ), .A2(_u10_u20_n2367 ), .ZN(_u10_u20_n3106 ) );
NAND2_X1 _u10_u20_U940  ( .A1(_u10_u20_n2977 ), .A2(_u10_u20_n3000 ), .ZN(_u10_u20_n3110 ) );
NAND2_X1 _u10_u20_U939  ( .A1(_u10_u20_n3109 ), .A2(_u10_u20_n3110 ), .ZN(_u10_u20_n1924 ) );
AND2_X1 _u10_u20_U938  ( .A1(_u10_u20_n1924 ), .A2(_u10_u20_n3108 ), .ZN(_u10_u20_n3107 ) );
NOR2_X1 _u10_u20_U937  ( .A1(_u10_u20_n3106 ), .A2(_u10_u20_n3107 ), .ZN(_u10_u20_n3105 ) );
NOR2_X1 _u10_u20_U936  ( .A1(_u10_u20_n3105 ), .A2(_u10_u20_n2008 ), .ZN(_u10_u20_n3104 ) );
NOR3_X1 _u10_u20_U935  ( .A1(_u10_u20_n3102 ), .A2(_u10_u20_n3103 ), .A3(_u10_u20_n3104 ), .ZN(_u10_u20_n3101 ) );
NAND4_X1 _u10_u20_U934  ( .A1(_u10_u20_n3098 ), .A2(_u10_u20_n3099 ), .A3(_u10_u20_n3100 ), .A4(_u10_u20_n3101 ), .ZN(_u10_u20_n3071 ) );
NOR2_X1 _u10_u20_U933  ( .A1(_u10_u20_n1926 ), .A2(_u10_u20_n2980 ), .ZN(_u10_u20_n2218 ) );
INV_X1 _u10_u20_U932  ( .A(_u10_u20_n2721 ), .ZN(_u10_u20_n2910 ) );
NAND2_X1 _u10_u20_U931  ( .A1(_u10_u20_n2910 ), .A2(_u10_u20_n1869 ), .ZN(_u10_u20_n2779 ) );
NAND2_X1 _u10_u20_U930  ( .A1(_u10_u20_n2218 ), .A2(_u10_u20_n2779 ), .ZN(_u10_u20_n3081 ) );
NAND2_X1 _u10_u20_U929  ( .A1(_u10_u20_n1922 ), .A2(_u10_u20_n1864 ), .ZN(_u10_u20_n2179 ) );
NOR3_X1 _u10_u20_U928  ( .A1(_u10_u20_n1961 ), .A2(_u10_u20_n1918 ), .A3(_u10_u20_n2179 ), .ZN(_u10_u20_n2693 ) );
NAND2_X1 _u10_u20_U927  ( .A1(_u10_u20_n3097 ), .A2(_u10_u20_n1924 ), .ZN(_u10_u20_n3096 ) );
NAND2_X1 _u10_u20_U926  ( .A1(_u10_u20_n1984 ), .A2(_u10_u20_n3096 ), .ZN(_u10_u20_n2506 ) );
INV_X1 _u10_u20_U925  ( .A(_u10_u20_n2506 ), .ZN(_u10_u20_n2366 ) );
NAND2_X1 _u10_u20_U924  ( .A1(_u10_u20_n2366 ), .A2(_u10_u20_n2375 ), .ZN(_u10_u20_n2236 ) );
NAND2_X1 _u10_u20_U923  ( .A1(_u10_u20_n2693 ), .A2(_u10_u20_n2236 ), .ZN(_u10_u20_n3082 ) );
NAND2_X1 _u10_u20_U922  ( .A1(1'b0), .A2(_u10_u20_n2126 ), .ZN(_u10_u20_n3095 ) );
NAND2_X1 _u10_u20_U921  ( .A1(_u10_u20_n1956 ), .A2(_u10_u20_n3095 ), .ZN(_u10_u20_n2907 ) );
OR2_X1 _u10_u20_U920  ( .A1(_u10_u20_n2902 ), .A2(_u10_u20_n2907 ), .ZN(_u10_u20_n3085 ) );
NAND2_X1 _u10_u20_U919  ( .A1(_u10_u20_n2256 ), .A2(_u10_u20_n2113 ), .ZN(_u10_u20_n3094 ) );
NAND2_X1 _u10_u20_U918  ( .A1(_u10_u20_n2688 ), .A2(_u10_u20_n3094 ), .ZN(_u10_u20_n3092 ) );
NAND2_X1 _u10_u20_U917  ( .A1(_u10_u20_n3093 ), .A2(_u10_u20_n3092 ), .ZN(_u10_u20_n3086 ) );
INV_X1 _u10_u20_U916  ( .A(_u10_u20_n2159 ), .ZN(_u10_u20_n1894 ) );
NAND2_X1 _u10_u20_U915  ( .A1(_u10_u20_n3067 ), .A2(_u10_u20_n1894 ), .ZN(_u10_u20_n3091 ) );
INV_X1 _u10_u20_U914  ( .A(_u10_u20_n3092 ), .ZN(_u10_u20_n2234 ) );
NAND3_X1 _u10_u20_U913  ( .A1(_u10_u20_n3091 ), .A2(_u10_u20_n2126 ), .A3(_u10_u20_n2234 ), .ZN(_u10_u20_n3090 ) );
NAND2_X1 _u10_u20_U912  ( .A1(1'b0), .A2(_u10_u20_n3090 ), .ZN(_u10_u20_n3087 ) );
NAND3_X1 _u10_u20_U911  ( .A1(_u10_u20_n2329 ), .A2(_u10_u20_n3089 ), .A3(_u10_u20_n2549 ), .ZN(_u10_u20_n3088 ) );
NAND4_X1 _u10_u20_U910  ( .A1(_u10_u20_n3085 ), .A2(_u10_u20_n3086 ), .A3(_u10_u20_n3087 ), .A4(_u10_u20_n3088 ), .ZN(_u10_u20_n3084 ) );
NAND2_X1 _u10_u20_U909  ( .A1(_u10_u20_n3084 ), .A2(_u10_u20_n2803 ), .ZN(_u10_u20_n3083 ) );
NAND3_X1 _u10_u20_U908  ( .A1(_u10_u20_n3081 ), .A2(_u10_u20_n3082 ), .A3(_u10_u20_n3083 ), .ZN(_u10_u20_n3072 ) );
INV_X1 _u10_u20_U907  ( .A(_u10_u20_n2689 ), .ZN(_u10_u20_n1955 ) );
NOR3_X1 _u10_u20_U906  ( .A1(_u10_u20_n1955 ), .A2(_u10_u20_n2813 ), .A3(_u10_u20_n2488 ), .ZN(_u10_u20_n3080 ) );
NOR2_X1 _u10_u20_U905  ( .A1(_u10_u20_n3080 ), .A2(_u10_u20_n2485 ), .ZN(_u10_u20_n3073 ) );
NAND3_X1 _u10_u20_U904  ( .A1(_u10_u20_n2621 ), .A2(_u10_u20_n2202 ), .A3(_u10_u20_n3079 ), .ZN(_u10_u20_n2110 ) );
NOR2_X1 _u10_u20_U903  ( .A1(_u10_u20_n2110 ), .A2(_u10_u20_n2218 ), .ZN(_u10_u20_n2775 ) );
INV_X1 _u10_u20_U902  ( .A(_u10_u20_n2775 ), .ZN(_u10_u20_n3024 ) );
INV_X1 _u10_u20_U901  ( .A(_u10_u20_n3078 ), .ZN(_u10_u20_n2133 ) );
INV_X1 _u10_u20_U900  ( .A(_u10_u20_n2007 ), .ZN(_u10_u20_n2358 ) );
NAND2_X1 _u10_u20_U899  ( .A1(_u10_u20_n2358 ), .A2(_u10_u20_n2886 ), .ZN(_u10_u20_n2240 ) );
INV_X1 _u10_u20_U898  ( .A(_u10_u20_n2240 ), .ZN(_u10_u20_n2083 ) );
NOR3_X1 _u10_u20_U897  ( .A1(_u10_u20_n2952 ), .A2(_u10_u20_n2004 ), .A3(_u10_u20_n1891 ), .ZN(_u10_u20_n3077 ) );
NAND3_X1 _u10_u20_U896  ( .A1(_u10_u20_n2083 ), .A2(_u10_u20_n2938 ), .A3(_u10_u20_n3077 ), .ZN(_u10_u20_n1886 ) );
NOR3_X1 _u10_u20_U895  ( .A1(_u10_u20_n3024 ), .A2(_u10_u20_n2133 ), .A3(_u10_u20_n1886 ), .ZN(_u10_u20_n3075 ) );
NOR2_X1 _u10_u20_U894  ( .A1(_u10_u20_n3075 ), .A2(_u10_u20_n3076 ), .ZN(_u10_u20_n3074 ) );
NOR4_X1 _u10_u20_U893  ( .A1(_u10_u20_n3071 ), .A2(_u10_u20_n3072 ), .A3(_u10_u20_n3073 ), .A4(_u10_u20_n3074 ), .ZN(_u10_u20_n3017 ) );
INV_X1 _u10_u20_U892  ( .A(_u10_u20_n3065 ), .ZN(_u10_u20_n3043 ) );
NAND2_X1 _u10_u20_U891  ( .A1(_u10_u20_n3043 ), .A2(_u10_u20_n2106 ), .ZN(_u10_u20_n3070 ) );
NAND2_X1 _u10_u20_U890  ( .A1(_u10_u20_n3070 ), .A2(_u10_u20_n2038 ), .ZN(_u10_u20_n3068 ) );
NAND2_X1 _u10_u20_U889  ( .A1(_u10_u20_n2344 ), .A2(_u10_u20_n2584 ), .ZN(_u10_u20_n3069 ) );
NAND3_X1 _u10_u20_U888  ( .A1(_u10_u20_n3068 ), .A2(_u10_u20_n1930 ), .A3(_u10_u20_n3069 ), .ZN(_u10_u20_n3047 ) );
NAND2_X1 _u10_u20_U887  ( .A1(_u10_u20_n2835 ), .A2(_u10_u20_n2466 ), .ZN(_u10_u20_n2130 ) );
INV_X1 _u10_u20_U886  ( .A(_u10_u20_n2130 ), .ZN(_u10_u20_n2168 ) );
NAND3_X1 _u10_u20_U885  ( .A1(_u10_u20_n3067 ), .A2(_u10_u20_n2329 ), .A3(_u10_u20_n2168 ), .ZN(_u10_u20_n2665 ) );
NAND3_X1 _u10_u20_U884  ( .A1(_u10_u20_n3065 ), .A2(_u10_u20_n3066 ), .A3(_u10_u20_n2342 ), .ZN(_u10_u20_n3064 ) );
NAND3_X1 _u10_u20_U883  ( .A1(_u10_u20_n3064 ), .A2(_u10_u20_n2175 ), .A3(_u10_u20_n2987 ), .ZN(_u10_u20_n3048 ) );
NOR3_X1 _u10_u20_U882  ( .A1(_u10_u20_n1849 ), .A2(1'b0), .A3(_u10_u20_n3063 ), .ZN(_u10_u20_n3050 ) );
NOR3_X1 _u10_u20_U881  ( .A1(_u10_u20_n2406 ), .A2(1'b0), .A3(_u10_u20_n3062 ), .ZN(_u10_u20_n3060 ) );
NOR3_X1 _u10_u20_U880  ( .A1(_u10_u20_n3060 ), .A2(1'b0), .A3(_u10_u20_n3061 ), .ZN(_u10_u20_n3051 ) );
NAND2_X1 _u10_u20_U879  ( .A1(_u10_u20_n3059 ), .A2(_u10_u20_n2049 ), .ZN(_u10_u20_n3056 ) );
NAND3_X1 _u10_u20_U878  ( .A1(_u10_u20_n3056 ), .A2(_u10_u20_n3057 ), .A3(_u10_u20_n3058 ), .ZN(_u10_u20_n3054 ) );
NOR4_X1 _u10_u20_U877  ( .A1(_u10_u20_n3054 ), .A2(_u10_u20_n3055 ), .A3(_u10_u20_n2055 ), .A4(_u10_u20_n2056 ), .ZN(_u10_u20_n3053 ) );
NOR3_X1 _u10_u20_U876  ( .A1(_u10_u20_n2346 ), .A2(1'b0), .A3(_u10_u20_n3053 ), .ZN(_u10_u20_n3052 ) );
NOR3_X1 _u10_u20_U875  ( .A1(_u10_u20_n3050 ), .A2(_u10_u20_n3051 ), .A3(_u10_u20_n3052 ), .ZN(_u10_u20_n3049 ) );
NAND4_X1 _u10_u20_U874  ( .A1(_u10_u20_n3047 ), .A2(_u10_u20_n2665 ), .A3(_u10_u20_n3048 ), .A4(_u10_u20_n3049 ), .ZN(_u10_u20_n3019 ) );
NAND2_X1 _u10_u20_U873  ( .A1(_u10_u20_n2056 ), .A2(_u10_u20_n2019 ), .ZN(_u10_u20_n3046 ) );
NAND2_X1 _u10_u20_U872  ( .A1(_u10_u20_n3045 ), .A2(_u10_u20_n3046 ), .ZN(_u10_u20_n3044 ) );
NAND2_X1 _u10_u20_U871  ( .A1(_u10_u20_n3044 ), .A2(_u10_u20_n2165 ), .ZN(_u10_u20_n3028 ) );
OR2_X1 _u10_u20_U870  ( .A1(_u10_u20_n2179 ), .A2(_u10_u20_n1961 ), .ZN(_u10_u20_n3037 ) );
NAND2_X1 _u10_u20_U869  ( .A1(_u10_u20_n3043 ), .A2(_u10_u20_n2336 ), .ZN(_u10_u20_n3042 ) );
NAND2_X1 _u10_u20_U868  ( .A1(_u10_u20_n3042 ), .A2(_u10_u20_n3006 ), .ZN(_u10_u20_n3041 ) );
NAND2_X1 _u10_u20_U867  ( .A1(_u10_u20_n3040 ), .A2(_u10_u20_n3041 ), .ZN(_u10_u20_n3026 ) );
NAND4_X1 _u10_u20_U866  ( .A1(_u10_u20_n3026 ), .A2(_u10_u20_n2520 ), .A3(_u10_u20_n1962 ), .A4(_u10_u20_n1864 ), .ZN(_u10_u20_n3039 ) );
NAND2_X1 _u10_u20_U865  ( .A1(_u10_u20_n3039 ), .A2(_u10_u20_n1922 ), .ZN(_u10_u20_n3038 ) );
NAND2_X1 _u10_u20_U864  ( .A1(_u10_u20_n3037 ), .A2(_u10_u20_n3038 ), .ZN(_u10_u20_n3035 ) );
NAND2_X1 _u10_u20_U863  ( .A1(_u10_u20_n2985 ), .A2(_u10_u20_n3036 ), .ZN(_u10_u20_n2432 ) );
NAND2_X1 _u10_u20_U862  ( .A1(_u10_u20_n3035 ), .A2(_u10_u20_n2432 ), .ZN(_u10_u20_n3029 ) );
INV_X1 _u10_u20_U861  ( .A(_u10_u20_n3034 ), .ZN(_u10_u20_n2777 ) );
INV_X1 _u10_u20_U860  ( .A(_u10_u20_n2772 ), .ZN(_u10_u20_n3032 ) );
NAND2_X1 _u10_u20_U859  ( .A1(_u10_u20_n1982 ), .A2(_u10_u20_n2978 ), .ZN(_u10_u20_n3033 ) );
NAND2_X1 _u10_u20_U858  ( .A1(_u10_u20_n3032 ), .A2(_u10_u20_n3033 ), .ZN(_u10_u20_n3031 ) );
NAND2_X1 _u10_u20_U857  ( .A1(_u10_u20_n2777 ), .A2(_u10_u20_n3031 ), .ZN(_u10_u20_n3030 ) );
NAND3_X1 _u10_u20_U856  ( .A1(_u10_u20_n3028 ), .A2(_u10_u20_n3029 ), .A3(_u10_u20_n3030 ), .ZN(_u10_u20_n3020 ) );
NOR3_X1 _u10_u20_U855  ( .A1(_u10_u20_n2179 ), .A2(1'b0), .A3(_u10_u20_n2375 ), .ZN(_u10_u20_n3027 ) );
NOR2_X1 _u10_u20_U854  ( .A1(_u10_u20_n3027 ), .A2(_u10_u20_n2177 ), .ZN(_u10_u20_n3025 ) );
NOR2_X1 _u10_u20_U853  ( .A1(_u10_u20_n3025 ), .A2(_u10_u20_n3026 ), .ZN(_u10_u20_n3021 ) );
NOR2_X1 _u10_u20_U852  ( .A1(_u10_u20_n2256 ), .A2(_u10_u20_n3024 ), .ZN(_u10_u20_n3023 ) );
NOR2_X1 _u10_u20_U851  ( .A1(_u10_u20_n3023 ), .A2(_u10_u20_n1868 ), .ZN(_u10_u20_n3022 ) );
NOR4_X1 _u10_u20_U850  ( .A1(_u10_u20_n3019 ), .A2(_u10_u20_n3020 ), .A3(_u10_u20_n3021 ), .A4(_u10_u20_n3022 ), .ZN(_u10_u20_n3018 ) );
NAND4_X1 _u10_u20_U849  ( .A1(_u10_u20_n3015 ), .A2(_u10_u20_n3016 ), .A3(_u10_u20_n3017 ), .A4(_u10_u20_n3018 ), .ZN(_u10_u20_n2958 ) );
NOR2_X1 _u10_u20_U848  ( .A1(1'b0), .A2(_u10_u20_n2573 ), .ZN(_u10_u20_n3011 ) );
NOR2_X1 _u10_u20_U847  ( .A1(1'b0), .A2(_u10_u20_n2359 ), .ZN(_u10_u20_n3012 ) );
NOR2_X1 _u10_u20_U846  ( .A1(1'b0), .A2(_u10_u20_n1859 ), .ZN(_u10_u20_n3013 ) );
NOR2_X1 _u10_u20_U845  ( .A1(1'b0), .A2(_u10_u20_n1836 ), .ZN(_u10_u20_n3014 ) );
NOR4_X1 _u10_u20_U844  ( .A1(_u10_u20_n3011 ), .A2(_u10_u20_n3012 ), .A3(_u10_u20_n3013 ), .A4(_u10_u20_n3014 ), .ZN(_u10_u20_n2959 ) );
NOR2_X1 _u10_u20_U843  ( .A1(1'b0), .A2(_u10_u20_n2025 ), .ZN(_u10_u20_n3007 ) );
NOR2_X1 _u10_u20_U842  ( .A1(1'b0), .A2(_u10_u20_n2085 ), .ZN(_u10_u20_n3008 ) );
NOR2_X1 _u10_u20_U841  ( .A1(1'b0), .A2(_u10_u20_n2607 ), .ZN(_u10_u20_n3009 ) );
NOR2_X1 _u10_u20_U840  ( .A1(1'b0), .A2(_u10_u20_n2071 ), .ZN(_u10_u20_n3010 ) );
NOR4_X1 _u10_u20_U839  ( .A1(_u10_u20_n3007 ), .A2(_u10_u20_n3008 ), .A3(_u10_u20_n3009 ), .A4(_u10_u20_n3010 ), .ZN(_u10_u20_n2960 ) );
NAND2_X1 _u10_u20_U838  ( .A1(_u10_u20_n1894 ), .A2(_u10_u20_n2466 ), .ZN(_u10_u20_n3002 ) );
NAND2_X1 _u10_u20_U837  ( .A1(_u10_u20_n2830 ), .A2(_u10_u20_n2600 ), .ZN(_u10_u20_n3003 ) );
NAND2_X1 _u10_u20_U836  ( .A1(_u10_u20_n1960 ), .A2(_u10_u20_n2431 ), .ZN(_u10_u20_n3004 ) );
NAND2_X1 _u10_u20_U835  ( .A1(_u10_u20_n2002 ), .A2(_u10_u20_n3006 ), .ZN(_u10_u20_n3005 ) );
NAND4_X1 _u10_u20_U834  ( .A1(_u10_u20_n3002 ), .A2(_u10_u20_n3003 ), .A3(_u10_u20_n3004 ), .A4(_u10_u20_n3005 ), .ZN(_u10_u20_n2992 ) );
NAND2_X1 _u10_u20_U833  ( .A1(_u10_u20_n2461 ), .A2(_u10_u20_n3001 ), .ZN(_u10_u20_n2997 ) );
NAND2_X1 _u10_u20_U832  ( .A1(_u10_u20_n2999 ), .A2(_u10_u20_n3000 ), .ZN(_u10_u20_n2998 ) );
NAND2_X1 _u10_u20_U831  ( .A1(_u10_u20_n2997 ), .A2(_u10_u20_n2998 ), .ZN(_u10_u20_n2993 ) );
NOR2_X1 _u10_u20_U830  ( .A1(_u10_SYNOPSYS_UNCONNECTED_4 ), .A2(_u10_u20_n2996 ), .ZN(_u10_u20_n2995 ) );
NOR2_X1 _u10_u20_U829  ( .A1(_u10_u20_n2995 ), .A2(_u10_u20_n2126 ), .ZN(_u10_u20_n2994 ) );
NOR4_X1 _u10_u20_U828  ( .A1(_u10_u20_n2992 ), .A2(_u10_u20_n2993 ), .A3(next_ch), .A4(_u10_u20_n2994 ), .ZN(_u10_u20_n2961 ) );
NAND2_X1 _u10_u20_U827  ( .A1(_u10_u20_n2445 ), .A2(_u10_u20_n2803 ), .ZN(_u10_u20_n2988 ) );
OR2_X1 _u10_u20_U826  ( .A1(_u10_u20_n2584 ), .A2(1'b0), .ZN(_u10_u20_n2989 ) );
NAND2_X1 _u10_u20_U825  ( .A1(_u10_u20_n2709 ), .A2(_u10_u20_n2080 ), .ZN(_u10_u20_n2990 ) );
NAND2_X1 _u10_u20_U824  ( .A1(_u10_u20_n2183 ), .A2(_u10_u20_n2166 ), .ZN(_u10_u20_n2991 ) );
NAND4_X1 _u10_u20_U823  ( .A1(_u10_u20_n2988 ), .A2(_u10_u20_n2989 ), .A3(_u10_u20_n2990 ), .A4(_u10_u20_n2991 ), .ZN(_u10_u20_n2963 ) );
NAND2_X1 _u10_u20_U822  ( .A1(_u10_u20_n2987 ), .A2(_u10_u20_n1930 ), .ZN(_u10_u20_n2981 ) );
NAND2_X1 _u10_u20_U821  ( .A1(_u10_u20_n2986 ), .A2(_u10_u20_n2038 ), .ZN(_u10_u20_n2982 ) );
OR2_X1 _u10_u20_U820  ( .A1(_u10_u20_n2985 ), .A2(1'b0), .ZN(_u10_u20_n2983 ) );
NAND2_X1 _u10_u20_U819  ( .A1(_u10_u20_n2169 ), .A2(_u10_u20_n2113 ), .ZN(_u10_u20_n2984 ) );
NAND4_X1 _u10_u20_U818  ( .A1(_u10_u20_n2981 ), .A2(_u10_u20_n2982 ), .A3(_u10_u20_n2983 ), .A4(_u10_u20_n2984 ), .ZN(_u10_u20_n2964 ) );
NAND2_X1 _u10_u20_U817  ( .A1(_u10_u20_n2509 ), .A2(_u10_u20_n1864 ), .ZN(_u10_u20_n2973 ) );
INV_X1 _u10_u20_U816  ( .A(_u10_u20_n2980 ), .ZN(_u10_u20_n1861 ) );
NAND2_X1 _u10_u20_U815  ( .A1(_u10_u20_n1861 ), .A2(_u10_u20_n1922 ), .ZN(_u10_u20_n2974 ) );
NAND2_X1 _u10_u20_U814  ( .A1(_u10_u20_n2979 ), .A2(_u10_u20_n2405 ), .ZN(_u10_u20_n2975 ) );
NAND2_X1 _u10_u20_U813  ( .A1(_u10_u20_n2977 ), .A2(_u10_u20_n2978 ), .ZN(_u10_u20_n2976 ) );
NAND4_X1 _u10_u20_U812  ( .A1(_u10_u20_n2973 ), .A2(_u10_u20_n2974 ), .A3(_u10_u20_n2975 ), .A4(_u10_u20_n2976 ), .ZN(_u10_u20_n2965 ) );
NAND2_X1 _u10_u20_U811  ( .A1(_u10_u20_n2507 ), .A2(_u10_u20_n2972 ), .ZN(_u10_u20_n2967 ) );
NAND2_X1 _u10_u20_U810  ( .A1(_u10_u20_n2043 ), .A2(_u10_u20_n1965 ), .ZN(_u10_u20_n2968 ) );
NAND2_X1 _u10_u20_U809  ( .A1(_u10_u20_n2063 ), .A2(_u10_u20_n1853 ), .ZN(_u10_u20_n2969 ) );
NAND2_X1 _u10_u20_U808  ( .A1(_u10_u20_n2971 ), .A2(_u10_u20_n2175 ), .ZN(_u10_u20_n2970 ) );
NAND4_X1 _u10_u20_U807  ( .A1(_u10_u20_n2967 ), .A2(_u10_u20_n2968 ), .A3(_u10_u20_n2969 ), .A4(_u10_u20_n2970 ), .ZN(_u10_u20_n2966 ) );
NOR4_X1 _u10_u20_U806  ( .A1(_u10_u20_n2963 ), .A2(_u10_u20_n2964 ), .A3(_u10_u20_n2965 ), .A4(_u10_u20_n2966 ), .ZN(_u10_u20_n2962 ) );
AND4_X1 _u10_u20_U805  ( .A1(_u10_u20_n2959 ), .A2(_u10_u20_n2960 ), .A3(_u10_u20_n2961 ), .A4(_u10_u20_n2962 ), .ZN(_u10_u20_n1819 ) );
MUX2_X1 _u10_u20_U804  ( .A(_u10_u20_n2958 ), .B(_u10_SYNOPSYS_UNCONNECTED_8 ), .S(_u10_u20_n1819 ), .Z(_u10_u20_n1808 ) );
NOR2_X1 _u10_u20_U803  ( .A1(_u10_u20_n2531 ), .A2(_u10_u20_n2607 ), .ZN(_u10_u20_n1911 ) );
NAND2_X1 _u10_u20_U802  ( .A1(_u10_u20_n1911 ), .A2(_u10_u20_n2957 ), .ZN(_u10_u20_n2954 ) );
NAND2_X1 _u10_u20_U801  ( .A1(_u10_u20_n1853 ), .A2(_u10_u20_n1965 ), .ZN(_u10_u20_n2956 ) );
NAND2_X1 _u10_u20_U800  ( .A1(_u10_u20_n1966 ), .A2(_u10_u20_n2956 ), .ZN(_u10_u20_n2955 ) );
NAND2_X1 _u10_u20_U799  ( .A1(_u10_u20_n2954 ), .A2(_u10_u20_n2955 ), .ZN(_u10_u20_n2670 ) );
NOR3_X1 _u10_u20_U798  ( .A1(_u10_u20_n1852 ), .A2(1'b0), .A3(_u10_u20_n1853 ), .ZN(_u10_u20_n2708 ) );
NAND2_X1 _u10_u20_U797  ( .A1(_u10_u20_n2708 ), .A2(_u10_u20_n2080 ), .ZN(_u10_u20_n2355 ) );
NOR2_X1 _u10_u20_U796  ( .A1(_u10_u20_n2355 ), .A2(1'b0), .ZN(_u10_u20_n2599 ) );
NAND2_X1 _u10_u20_U795  ( .A1(_u10_u20_n2953 ), .A2(_u10_u20_n2599 ), .ZN(_u10_u20_n2423 ) );
OR2_X1 _u10_u20_U794  ( .A1(_u10_u20_n2423 ), .A2(_u10_u20_n2359 ), .ZN(_u10_u20_n2949 ) );
NAND3_X1 _u10_u20_U793  ( .A1(_u10_u20_n2105 ), .A2(_u10_u20_n1936 ), .A3(_u10_u20_n2952 ), .ZN(_u10_u20_n2950 ) );
NAND3_X1 _u10_u20_U792  ( .A1(_u10_u20_n2549 ), .A2(_u10_u20_n1936 ), .A3(1'b0), .ZN(_u10_u20_n2096 ) );
INV_X1 _u10_u20_U791  ( .A(_u10_u20_n2096 ), .ZN(_u10_u20_n2301 ) );
NAND2_X1 _u10_u20_U790  ( .A1(_u10_u20_n2301 ), .A2(_u10_u20_n2446 ), .ZN(_u10_u20_n2368 ) );
INV_X1 _u10_u20_U789  ( .A(_u10_u20_n2368 ), .ZN(_u10_u20_n2326 ) );
NAND2_X1 _u10_u20_U788  ( .A1(_u10_u20_n2326 ), .A2(_u10_u20_n2941 ), .ZN(_u10_u20_n2800 ) );
INV_X1 _u10_u20_U787  ( .A(_u10_u20_n2800 ), .ZN(_u10_u20_n2081 ) );
NAND2_X1 _u10_u20_U786  ( .A1(_u10_u20_n2081 ), .A2(_u10_u20_n2049 ), .ZN(_u10_u20_n2855 ) );
INV_X1 _u10_u20_U785  ( .A(_u10_u20_n2855 ), .ZN(_u10_u20_n2347 ) );
NAND2_X1 _u10_u20_U784  ( .A1(_u10_u20_n2347 ), .A2(_u10_u20_n2063 ), .ZN(_u10_u20_n2951 ) );
NAND3_X1 _u10_u20_U783  ( .A1(_u10_u20_n2949 ), .A2(_u10_u20_n2950 ), .A3(_u10_u20_n2951 ), .ZN(_u10_u20_n1997 ) );
INV_X1 _u10_u20_U782  ( .A(_u10_u20_n1997 ), .ZN(_u10_u20_n2917 ) );
AND2_X1 _u10_u20_U781  ( .A1(_u10_u20_n2709 ), .A2(_u10_u20_n2708 ), .ZN(_u10_u20_n2942 ) );
INV_X1 _u10_u20_U780  ( .A(_u10_u20_n2907 ), .ZN(_u10_u20_n2737 ) );
NAND2_X1 _u10_u20_U779  ( .A1(_u10_u20_n2737 ), .A2(_u10_u20_n2803 ), .ZN(_u10_u20_n1888 ) );
NOR2_X1 _u10_u20_U778  ( .A1(_u10_u20_n2001 ), .A2(_u10_u20_n1888 ), .ZN(_u10_u20_n2943 ) );
NAND4_X1 _u10_u20_U777  ( .A1(1'b0), .A2(_u10_u20_n2078 ), .A3(_u10_u20_n2059 ), .A4(_u10_u20_n2031 ), .ZN(_u10_u20_n2578 ) );
NOR3_X1 _u10_u20_U776  ( .A1(_u10_u20_n2719 ), .A2(_u10_u20_n2130 ), .A3(_u10_u20_n2305 ), .ZN(_u10_u20_n2386 ) );
NAND2_X1 _u10_u20_U775  ( .A1(_u10_u20_n2386 ), .A2(_u10_u20_n2669 ), .ZN(_u10_u20_n2948 ) );
NAND3_X1 _u10_u20_U774  ( .A1(_u10_u20_n2578 ), .A2(_u10_u20_n2947 ), .A3(_u10_u20_n2948 ), .ZN(_u10_u20_n2750 ) );
NOR2_X1 _u10_u20_U773  ( .A1(_u10_u20_n2274 ), .A2(_u10_u20_n2852 ), .ZN(_u10_u20_n2946 ) );
NOR3_X1 _u10_u20_U772  ( .A1(_u10_u20_n2750 ), .A2(1'b0), .A3(_u10_u20_n2946 ), .ZN(_u10_u20_n2945 ) );
NOR2_X1 _u10_u20_U771  ( .A1(_u10_u20_n2945 ), .A2(_u10_u20_n2359 ), .ZN(_u10_u20_n2944 ) );
NOR3_X1 _u10_u20_U770  ( .A1(_u10_u20_n2942 ), .A2(_u10_u20_n2943 ), .A3(_u10_u20_n2944 ), .ZN(_u10_u20_n2919 ) );
NOR2_X1 _u10_u20_U769  ( .A1(_u10_u20_n2423 ), .A2(1'b0), .ZN(_u10_u20_n1979 ) );
NAND3_X1 _u10_u20_U768  ( .A1(_u10_u20_n2549 ), .A2(_u10_u20_n1936 ), .A3(_u10_u20_n1979 ), .ZN(_u10_u20_n2328 ) );
INV_X1 _u10_u20_U767  ( .A(_u10_u20_n2328 ), .ZN(_u10_u20_n2554 ) );
NAND3_X1 _u10_u20_U766  ( .A1(_u10_u20_n2941 ), .A2(_u10_u20_n2446 ), .A3(_u10_u20_n2554 ), .ZN(_u10_u20_n2115 ) );
NOR2_X1 _u10_u20_U765  ( .A1(_u10_u20_n2578 ), .A2(_u10_u20_n2030 ), .ZN(_u10_u20_n2553 ) );
INV_X1 _u10_u20_U764  ( .A(_u10_u20_n2553 ), .ZN(_u10_u20_n2269 ) );
NOR2_X1 _u10_u20_U763  ( .A1(_u10_u20_n2269 ), .A2(_u10_u20_n2790 ), .ZN(_u10_u20_n2657 ) );
INV_X1 _u10_u20_U762  ( .A(_u10_u20_n2657 ), .ZN(_u10_u20_n2210 ) );
NOR2_X1 _u10_u20_U761  ( .A1(_u10_u20_n2210 ), .A2(_u10_u20_n2911 ), .ZN(_u10_u20_n2213 ) );
INV_X1 _u10_u20_U760  ( .A(_u10_u20_n2213 ), .ZN(_u10_u20_n2456 ) );
NAND2_X1 _u10_u20_U759  ( .A1(_u10_u20_n2115 ), .A2(_u10_u20_n2456 ), .ZN(_u10_u20_n2634 ) );
INV_X1 _u10_u20_U758  ( .A(_u10_u20_n2634 ), .ZN(_u10_u20_n2220 ) );
NOR2_X1 _u10_u20_U757  ( .A1(_u10_u20_n2081 ), .A2(_u10_u20_n2386 ), .ZN(_u10_u20_n2131 ) );
NAND2_X1 _u10_u20_U756  ( .A1(_u10_u20_n2940 ), .A2(_u10_u20_n2131 ), .ZN(_u10_u20_n2138 ) );
INV_X1 _u10_u20_U755  ( .A(_u10_u20_n2138 ), .ZN(_u10_u20_n2927 ) );
NAND2_X1 _u10_u20_U754  ( .A1(_u10_u20_n2220 ), .A2(_u10_u20_n2927 ), .ZN(_u10_u20_n2939 ) );
NAND2_X1 _u10_u20_U753  ( .A1(_u10_u20_n1885 ), .A2(_u10_u20_n2939 ), .ZN(_u10_u20_n2931 ) );
NAND3_X1 _u10_u20_U752  ( .A1(_u10_u20_n1859 ), .A2(_u10_u20_n2365 ), .A3(_u10_u20_n2938 ), .ZN(_u10_u20_n2935 ) );
NAND3_X1 _u10_u20_U751  ( .A1(_u10_u20_n2927 ), .A2(_u10_u20_n2937 ), .A3(_u10_u20_n2220 ), .ZN(_u10_u20_n2936 ) );
NAND2_X1 _u10_u20_U750  ( .A1(_u10_u20_n2935 ), .A2(_u10_u20_n2936 ), .ZN(_u10_u20_n2932 ) );
INV_X1 _u10_u20_U749  ( .A(_u10_u20_n1937 ), .ZN(_u10_u20_n2350 ) );
NAND2_X1 _u10_u20_U748  ( .A1(_u10_u20_n1913 ), .A2(_u10_u20_n2350 ), .ZN(_u10_u20_n2934 ) );
NAND2_X1 _u10_u20_U747  ( .A1(_u10_u20_n2386 ), .A2(_u10_u20_n2934 ), .ZN(_u10_u20_n2933 ) );
NAND3_X1 _u10_u20_U746  ( .A1(_u10_u20_n2931 ), .A2(_u10_u20_n2932 ), .A3(_u10_u20_n2933 ), .ZN(_u10_u20_n2921 ) );
OR2_X1 _u10_u20_U745  ( .A1(_u10_u20_n2213 ), .A2(_u10_u20_n2386 ), .ZN(_u10_u20_n2930 ) );
NAND2_X1 _u10_u20_U744  ( .A1(_u10_u20_n2049 ), .A2(_u10_u20_n2930 ), .ZN(_u10_u20_n2228 ) );
AND2_X1 _u10_u20_U743  ( .A1(_u10_u20_n2228 ), .A2(_u10_u20_n2699 ), .ZN(_u10_u20_n2929 ) );
NOR2_X1 _u10_u20_U742  ( .A1(_u10_u20_n2929 ), .A2(_u10_u20_n2495 ), .ZN(_u10_u20_n2922 ) );
NOR2_X1 _u10_u20_U741  ( .A1(_u10_u20_n2633 ), .A2(_u10_u20_n2877 ), .ZN(_u10_u20_n2928 ) );
NOR2_X1 _u10_u20_U740  ( .A1(_u10_u20_n2928 ), .A2(_u10_u20_n2886 ), .ZN(_u10_u20_n2923 ) );
NOR2_X1 _u10_u20_U739  ( .A1(_u10_u20_n2927 ), .A2(_u10_u20_n2531 ), .ZN(_u10_u20_n2926 ) );
NOR2_X1 _u10_u20_U738  ( .A1(_u10_u20_n2926 ), .A2(_u10_u20_n2687 ), .ZN(_u10_u20_n2925 ) );
NOR2_X1 _u10_u20_U737  ( .A1(_u10_u20_n2925 ), .A2(_u10_u20_n1849 ), .ZN(_u10_u20_n2924 ) );
NOR4_X1 _u10_u20_U736  ( .A1(_u10_u20_n2921 ), .A2(_u10_u20_n2922 ), .A3(_u10_u20_n2923 ), .A4(_u10_u20_n2924 ), .ZN(_u10_u20_n2920 ) );
NAND4_X1 _u10_u20_U735  ( .A1(_u10_u20_n2917 ), .A2(_u10_u20_n2918 ), .A3(_u10_u20_n2919 ), .A4(_u10_u20_n2920 ), .ZN(_u10_u20_n2312 ) );
NOR2_X1 _u10_u20_U734  ( .A1(_u10_u20_n2600 ), .A2(_u10_u20_n2686 ), .ZN(_u10_u20_n2401 ) );
NAND2_X1 _u10_u20_U733  ( .A1(_u10_u20_n2401 ), .A2(_u10_u20_n2549 ), .ZN(_u10_u20_n2547 ) );
INV_X1 _u10_u20_U732  ( .A(_u10_u20_n2547 ), .ZN(_u10_u20_n2794 ) );
NAND3_X1 _u10_u20_U731  ( .A1(_u10_u20_n2364 ), .A2(_u10_u20_n2667 ), .A3(_u10_u20_n2794 ), .ZN(_u10_u20_n2535 ) );
INV_X1 _u10_u20_U730  ( .A(_u10_u20_n2535 ), .ZN(_u10_u20_n2586 ) );
NAND2_X1 _u10_u20_U729  ( .A1(_u10_u20_n2586 ), .A2(_u10_u20_n2571 ), .ZN(_u10_u20_n2916 ) );
NAND2_X1 _u10_u20_U728  ( .A1(_u10_u20_n2837 ), .A2(_u10_u20_n2916 ), .ZN(_u10_u20_n2436 ) );
NAND2_X1 _u10_u20_U727  ( .A1(_u10_u20_n2915 ), .A2(_u10_u20_n2571 ), .ZN(_u10_u20_n2914 ) );
NAND2_X1 _u10_u20_U726  ( .A1(_u10_u20_n2166 ), .A2(_u10_u20_n2914 ), .ZN(_u10_u20_n2017 ) );
NOR2_X1 _u10_u20_U725  ( .A1(_u10_u20_n2485 ), .A2(_u10_u20_n1841 ), .ZN(_u10_u20_n2913 ) );
OR4_X1 _u10_u20_U724  ( .A1(_u10_u20_n2436 ), .A2(_u10_u20_n2017 ), .A3(_u10_u20_n2913 ), .A4(_u10_u20_n2442 ), .ZN(_u10_u20_n2912 ) );
NAND2_X1 _u10_u20_U723  ( .A1(_u10_u20_n2709 ), .A2(_u10_u20_n2912 ), .ZN(_u10_u20_n2888 ) );
NAND3_X1 _u10_u20_U722  ( .A1(_u10_u20_n2078 ), .A2(_u10_u20_n2031 ), .A3(1'b0), .ZN(_u10_u20_n2580 ) );
INV_X1 _u10_u20_U721  ( .A(_u10_u20_n2580 ), .ZN(_u10_u20_n2680 ) );
AND2_X1 _u10_u20_U720  ( .A1(_u10_u20_n2680 ), .A2(_u10_u20_n2668 ), .ZN(_u10_u20_n1950 ) );
NAND2_X1 _u10_u20_U719  ( .A1(_u10_u20_n1950 ), .A2(_u10_u20_n2089 ), .ZN(_u10_u20_n2095 ) );
INV_X1 _u10_u20_U718  ( .A(_u10_u20_n2095 ), .ZN(_u10_u20_n2542 ) );
NAND2_X1 _u10_u20_U717  ( .A1(_u10_u20_n2542 ), .A2(_u10_u20_n2446 ), .ZN(_u10_u20_n1887 ) );
NOR2_X1 _u10_u20_U716  ( .A1(_u10_u20_n1887 ), .A2(_u10_u20_n2911 ), .ZN(_u10_u20_n2114 ) );
INV_X1 _u10_u20_U715  ( .A(_u10_u20_n2114 ), .ZN(_u10_u20_n1940 ) );
NAND3_X1 _u10_u20_U714  ( .A1(_u10_u20_n2535 ), .A2(_u10_u20_n1940 ), .A3(_u10_u20_n2910 ), .ZN(_u10_u20_n2524 ) );
NAND2_X1 _u10_u20_U713  ( .A1(_u10_u20_n2524 ), .A2(_u10_u20_n2488 ), .ZN(_u10_u20_n2889 ) );
NAND2_X1 _u10_u20_U712  ( .A1(_u10_u20_n2220 ), .A2(_u10_u20_n1940 ), .ZN(_u10_u20_n2763 ) );
NOR2_X1 _u10_u20_U711  ( .A1(_u10_u20_n2763 ), .A2(_u10_u20_n2586 ), .ZN(_u10_u20_n2808 ) );
NOR2_X1 _u10_u20_U710  ( .A1(_u10_u20_n2808 ), .A2(_u10_u20_n2350 ), .ZN(_u10_u20_n2908 ) );
NOR2_X1 _u10_u20_U709  ( .A1(_u10_u20_n2544 ), .A2(_u10_u20_n1950 ), .ZN(_u10_u20_n2899 ) );
NOR2_X1 _u10_u20_U708  ( .A1(_u10_u20_n2899 ), .A2(_u10_u20_n2159 ), .ZN(_u10_u20_n2909 ) );
NOR2_X1 _u10_u20_U707  ( .A1(_u10_u20_n2908 ), .A2(_u10_u20_n2909 ), .ZN(_u10_u20_n2890 ) );
NOR3_X1 _u10_u20_U706  ( .A1(_u10_u20_n2547 ), .A2(_u10_u20_n1846 ), .A3(_u10_u20_n2907 ), .ZN(_u10_u20_n2892 ) );
NOR3_X1 _u10_u20_U705  ( .A1(_u10_u20_n2240 ), .A2(_u10_u20_n2377 ), .A3(_u10_u20_n1911 ), .ZN(_u10_u20_n2906 ) );
NOR2_X1 _u10_u20_U704  ( .A1(_u10_u20_n2906 ), .A2(_u10_u20_n2535 ), .ZN(_u10_u20_n2893 ) );
NAND2_X1 _u10_u20_U703  ( .A1(_u10_u20_n2554 ), .A2(_u10_u20_n2446 ), .ZN(_u10_u20_n2903 ) );
AND3_X1 _u10_u20_U702  ( .A1(_u10_u20_n2210 ), .A2(_u10_u20_n2905 ), .A3(_u10_u20_n1887 ), .ZN(_u10_u20_n2904 ) );
NAND4_X1 _u10_u20_U701  ( .A1(_u10_u20_n2902 ), .A2(_u10_u20_n2498 ), .A3(_u10_u20_n2903 ), .A4(_u10_u20_n2904 ), .ZN(_u10_u20_n2788 ) );
INV_X1 _u10_u20_U700  ( .A(_u10_u20_n2788 ), .ZN(_u10_u20_n2901 ) );
NOR2_X1 _u10_u20_U699  ( .A1(_u10_u20_n2901 ), .A2(_u10_u20_n1888 ), .ZN(_u10_u20_n2894 ) );
NOR2_X1 _u10_u20_U698  ( .A1(_u10_u20_n2401 ), .A2(_u10_u20_n2553 ), .ZN(_u10_u20_n2900 ) );
NOR2_X1 _u10_u20_U697  ( .A1(_u10_u20_n2900 ), .A2(_u10_u20_n1954 ), .ZN(_u10_u20_n2897 ) );
NOR2_X1 _u10_u20_U696  ( .A1(1'b0), .A2(_u10_u20_n2899 ), .ZN(_u10_u20_n2898 ) );
NOR2_X1 _u10_u20_U695  ( .A1(_u10_u20_n2897 ), .A2(_u10_u20_n2898 ), .ZN(_u10_u20_n2896 ) );
NOR2_X1 _u10_u20_U694  ( .A1(_u10_u20_n2896 ), .A2(_u10_u20_n1843 ), .ZN(_u10_u20_n2895 ) );
NOR4_X1 _u10_u20_U693  ( .A1(_u10_u20_n2892 ), .A2(_u10_u20_n2893 ), .A3(_u10_u20_n2894 ), .A4(_u10_u20_n2895 ), .ZN(_u10_u20_n2891 ) );
NAND4_X1 _u10_u20_U692  ( .A1(_u10_u20_n2888 ), .A2(_u10_u20_n2889 ), .A3(_u10_u20_n2890 ), .A4(_u10_u20_n2891 ), .ZN(_u10_u20_n2610 ) );
NOR4_X1 _u10_u20_U691  ( .A1(_u10_u20_n2670 ), .A2(_u10_u20_n2312 ), .A3(_u10_u20_n2610 ), .A4(_u10_u20_n2887 ), .ZN(_u10_u20_n2724 ) );
NOR2_X1 _u10_u20_U690  ( .A1(_u10_u20_n2883 ), .A2(_u10_u20_n2535 ), .ZN(_u10_u20_n2861 ) );
NOR2_X1 _u10_u20_U689  ( .A1(_u10_u20_n1855 ), .A2(_u10_u20_n1869 ), .ZN(_u10_u20_n2862 ) );
NOR2_X1 _u10_u20_U688  ( .A1(_u10_u20_n2886 ), .A2(_u10_u20_n2695 ), .ZN(_u10_u20_n2863 ) );
NAND2_X1 _u10_u20_U687  ( .A1(_u10_u20_n2813 ), .A2(_u10_u20_n2885 ), .ZN(_u10_u20_n2864 ) );
NAND2_X1 _u10_u20_U686  ( .A1(_u10_u20_n2114 ), .A2(_u10_u20_n2884 ), .ZN(_u10_u20_n2865 ) );
NAND2_X1 _u10_u20_U685  ( .A1(1'b0), .A2(_u10_u20_n2667 ), .ZN(_u10_u20_n2112 ) );
NOR3_X1 _u10_u20_U684  ( .A1(_u10_u20_n2883 ), .A2(_u10_u20_n2112 ), .A3(_u10_u20_n2719 ), .ZN(_u10_u20_n2878 ) );
INV_X1 _u10_u20_U683  ( .A(_u10_u20_n2112 ), .ZN(_u10_u20_n1856 ) );
NAND2_X1 _u10_u20_U682  ( .A1(_u10_u20_n2364 ), .A2(_u10_u20_n1856 ), .ZN(_u10_u20_n2882 ) );
NAND2_X1 _u10_u20_U681  ( .A1(_u10_u20_n2882 ), .A2(_u10_u20_n1869 ), .ZN(_u10_u20_n2050 ) );
INV_X1 _u10_u20_U680  ( .A(_u10_u20_n2050 ), .ZN(_u10_u20_n1939 ) );
NOR2_X1 _u10_u20_U679  ( .A1(_u10_u20_n1939 ), .A2(_u10_u20_n1841 ), .ZN(_u10_u20_n2881 ) );
NOR2_X1 _u10_u20_U678  ( .A1(_u10_u20_n2881 ), .A2(_u10_u20_n2840 ), .ZN(_u10_u20_n2880 ) );
NOR2_X1 _u10_u20_U677  ( .A1(_u10_u20_n2880 ), .A2(_u10_u20_n1836 ), .ZN(_u10_u20_n2879 ) );
NOR2_X1 _u10_u20_U676  ( .A1(_u10_u20_n2878 ), .A2(_u10_u20_n2879 ), .ZN(_u10_u20_n2866 ) );
NOR2_X1 _u10_u20_U675  ( .A1(_u10_u20_n2081 ), .A2(_u10_u20_n2877 ), .ZN(_u10_u20_n1840 ) );
NAND2_X1 _u10_u20_U674  ( .A1(_u10_u20_n1840 ), .A2(_u10_u20_n2115 ), .ZN(_u10_u20_n1873 ) );
NAND2_X1 _u10_u20_U673  ( .A1(_u10_u20_n2695 ), .A2(_u10_u20_n1940 ), .ZN(_u10_u20_n1874 ) );
NOR3_X1 _u10_u20_U672  ( .A1(_u10_u20_n2050 ), .A2(_u10_u20_n1873 ), .A3(_u10_u20_n1874 ), .ZN(_u10_u20_n2876 ) );
NOR2_X1 _u10_u20_U671  ( .A1(_u10_u20_n2876 ), .A2(_u10_u20_n1913 ), .ZN(_u10_u20_n2868 ) );
NAND2_X1 _u10_u20_U670  ( .A1(_u10_u20_n2875 ), .A2(_u10_u20_n2466 ), .ZN(_u10_u20_n2872 ) );
INV_X1 _u10_u20_U669  ( .A(_u10_u20_n1979 ), .ZN(_u10_u20_n2746 ) );
NAND2_X1 _u10_u20_U668  ( .A1(_u10_u20_n2874 ), .A2(_u10_u20_n2746 ), .ZN(_u10_u20_n1935 ) );
NAND3_X1 _u10_u20_U667  ( .A1(_u10_u20_n1935 ), .A2(_u10_u20_n1936 ), .A3(_u10_u20_n2467 ), .ZN(_u10_u20_n2873 ) );
NAND2_X1 _u10_u20_U666  ( .A1(_u10_u20_n2872 ), .A2(_u10_u20_n2873 ), .ZN(_u10_u20_n2264 ) );
AND2_X1 _u10_u20_U665  ( .A1(_u10_u20_n2264 ), .A2(_u10_u20_n2461 ), .ZN(_u10_u20_n2869 ) );
AND2_X1 _u10_u20_U664  ( .A1(_u10_u20_n1966 ), .A2(_u10_u20_n2761 ), .ZN(_u10_u20_n2870 ) );
NOR2_X1 _u10_u20_U663  ( .A1(_u10_u20_n2159 ), .A2(_u10_u20_n2163 ), .ZN(_u10_u20_n2871 ) );
NOR4_X1 _u10_u20_U662  ( .A1(_u10_u20_n2868 ), .A2(_u10_u20_n2869 ), .A3(_u10_u20_n2870 ), .A4(_u10_u20_n2871 ), .ZN(_u10_u20_n2867 ) );
NAND4_X1 _u10_u20_U661  ( .A1(_u10_u20_n2864 ), .A2(_u10_u20_n2865 ), .A3(_u10_u20_n2866 ), .A4(_u10_u20_n2867 ), .ZN(_u10_u20_n1992 ) );
NOR4_X1 _u10_u20_U660  ( .A1(_u10_u20_n2861 ), .A2(_u10_u20_n2862 ), .A3(_u10_u20_n2863 ), .A4(_u10_u20_n1992 ), .ZN(_u10_u20_n2725 ) );
NAND2_X1 _u10_u20_U659  ( .A1(_u10_u20_n2364 ), .A2(_u10_u20_n1846 ), .ZN(_u10_u20_n2744 ) );
NAND4_X1 _u10_u20_U658  ( .A1(_u10_u20_n2765 ), .A2(_u10_u20_n1939 ), .A3(_u10_u20_n2744 ), .A4(_u10_u20_n2535 ), .ZN(_u10_u20_n2860 ) );
NAND2_X1 _u10_u20_U657  ( .A1(_u10_u20_n2049 ), .A2(_u10_u20_n2860 ), .ZN(_u10_u20_n2856 ) );
NOR4_X1 _u10_u20_U656  ( .A1(1'b0), .A2(_u10_u20_n2858 ), .A3(_u10_u20_n2859 ), .A4(_u10_u20_n2051 ), .ZN(_u10_u20_n2857 ) );
NAND4_X1 _u10_u20_U655  ( .A1(_u10_u20_n2228 ), .A2(_u10_u20_n2855 ), .A3(_u10_u20_n2856 ), .A4(_u10_u20_n2857 ), .ZN(_u10_u20_n2854 ) );
NAND2_X1 _u10_u20_U654  ( .A1(_u10_u20_n2043 ), .A2(_u10_u20_n2854 ), .ZN(_u10_u20_n2821 ) );
INV_X1 _u10_u20_U653  ( .A(_u10_u20_n2071 ), .ZN(_u10_u20_n2279 ) );
INV_X1 _u10_u20_U652  ( .A(_u10_u20_n2599 ), .ZN(_u10_u20_n2357 ) );
OR2_X1 _u10_u20_U651  ( .A1(_u10_u20_n2744 ), .A2(_u10_u20_n2853 ), .ZN(_u10_u20_n2844 ) );
NAND2_X1 _u10_u20_U650  ( .A1(_u10_u20_n2131 ), .A2(_u10_u20_n2852 ), .ZN(_u10_u20_n2851 ) );
NAND2_X1 _u10_u20_U649  ( .A1(_u10_u20_n2082 ), .A2(_u10_u20_n2851 ), .ZN(_u10_u20_n2848 ) );
NAND2_X1 _u10_u20_U648  ( .A1(_u10_u20_n2850 ), .A2(_u10_u20_n2600 ), .ZN(_u10_u20_n2849 ) );
NAND3_X1 _u10_u20_U647  ( .A1(_u10_u20_n2848 ), .A2(_u10_u20_n2077 ), .A3(_u10_u20_n2849 ), .ZN(_u10_u20_n2287 ) );
NAND2_X1 _u10_u20_U646  ( .A1(_u10_u20_n2082 ), .A2(_u10_u20_n2050 ), .ZN(_u10_u20_n2847 ) );
NAND2_X1 _u10_u20_U645  ( .A1(_u10_u20_n2846 ), .A2(_u10_u20_n2847 ), .ZN(_u10_u20_n2074 ) );
NOR3_X1 _u10_u20_U644  ( .A1(_u10_u20_n2287 ), .A2(_u10_u20_n2596 ), .A3(_u10_u20_n2074 ), .ZN(_u10_u20_n2845 ) );
NAND4_X1 _u10_u20_U643  ( .A1(_u10_u20_n2357 ), .A2(_u10_u20_n2837 ), .A3(_u10_u20_n2844 ), .A4(_u10_u20_n2845 ), .ZN(_u10_u20_n2843 ) );
NAND2_X1 _u10_u20_U642  ( .A1(_u10_u20_n2279 ), .A2(_u10_u20_n2843 ), .ZN(_u10_u20_n2822 ) );
NOR3_X1 _u10_u20_U641  ( .A1(_u10_u20_n1925 ), .A2(_u10_u20_n2842 ), .A3(_u10_u20_n2686 ), .ZN(_u10_u20_n2841 ) );
NOR3_X1 _u10_u20_U640  ( .A1(_u10_u20_n2840 ), .A2(_u10_u20_n2599 ), .A3(_u10_u20_n2841 ), .ZN(_u10_u20_n2839 ) );
AND4_X1 _u10_u20_U639  ( .A1(_u10_u20_n2836 ), .A2(_u10_u20_n2837 ), .A3(_u10_u20_n2838 ), .A4(_u10_u20_n2839 ), .ZN(_u10_u20_n2454 ) );
NOR2_X1 _u10_u20_U638  ( .A1(_u10_u20_n2719 ), .A2(_u10_u20_n2835 ), .ZN(_u10_u20_n2773 ) );
NOR2_X1 _u10_u20_U637  ( .A1(_u10_u20_n2138 ), .A2(_u10_u20_n2773 ), .ZN(_u10_u20_n2814 ) );
NAND2_X1 _u10_u20_U636  ( .A1(_u10_u20_n2814 ), .A2(_u10_u20_n1869 ), .ZN(_u10_u20_n2834 ) );
NAND2_X1 _u10_u20_U635  ( .A1(_u10_u20_n2833 ), .A2(_u10_u20_n2834 ), .ZN(_u10_u20_n2832 ) );
NAND2_X1 _u10_u20_U634  ( .A1(_u10_u20_n2454 ), .A2(_u10_u20_n2832 ), .ZN(_u10_u20_n2831 ) );
NAND2_X1 _u10_u20_U633  ( .A1(_u10_u20_n2830 ), .A2(_u10_u20_n2831 ), .ZN(_u10_u20_n2823 ) );
INV_X1 _u10_u20_U632  ( .A(_u10_u20_n2025 ), .ZN(_u10_u20_n2470 ) );
NAND2_X1 _u10_u20_U631  ( .A1(_u10_u20_n1979 ), .A2(_u10_u20_n1936 ), .ZN(_u10_u20_n2829 ) );
AND2_X1 _u10_u20_U630  ( .A1(_u10_u20_n2828 ), .A2(_u10_u20_n2829 ), .ZN(_u10_u20_n2469 ) );
NAND2_X1 _u10_u20_U629  ( .A1(_u10_u20_n2469 ), .A2(_u10_u20_n2269 ), .ZN(_u10_u20_n2161 ) );
INV_X1 _u10_u20_U628  ( .A(_u10_u20_n2161 ), .ZN(_u10_u20_n2276 ) );
NOR2_X1 _u10_u20_U627  ( .A1(_u10_u20_n2274 ), .A2(_u10_u20_n2719 ), .ZN(_u10_u20_n2827 ) );
NOR3_X1 _u10_u20_U626  ( .A1(_u10_u20_n2827 ), .A2(_u10_u20_n2742 ), .A3(_u10_u20_n2680 ), .ZN(_u10_u20_n2826 ) );
NAND3_X1 _u10_u20_U625  ( .A1(_u10_u20_n2276 ), .A2(_u10_u20_n2108 ), .A3(_u10_u20_n2826 ), .ZN(_u10_u20_n2825 ) );
NAND2_X1 _u10_u20_U624  ( .A1(_u10_u20_n2470 ), .A2(_u10_u20_n2825 ), .ZN(_u10_u20_n2824 ) );
NAND4_X1 _u10_u20_U623  ( .A1(_u10_u20_n2821 ), .A2(_u10_u20_n2822 ), .A3(_u10_u20_n2823 ), .A4(_u10_u20_n2824 ), .ZN(_u10_u20_n2804 ) );
NAND2_X1 _u10_u20_U622  ( .A1(_u10_u20_n2131 ), .A2(_u10_u20_n2744 ), .ZN(_u10_u20_n2820 ) );
NAND2_X1 _u10_u20_U621  ( .A1(_u10_u20_n2571 ), .A2(_u10_u20_n2820 ), .ZN(_u10_u20_n2817 ) );
NOR2_X1 _u10_u20_U620  ( .A1(_u10_u20_n2819 ), .A2(_u10_u20_n2436 ), .ZN(_u10_u20_n2818 ) );
NAND4_X1 _u10_u20_U619  ( .A1(_u10_u20_n2437 ), .A2(_u10_u20_n2355 ), .A3(_u10_u20_n2817 ), .A4(_u10_u20_n2818 ), .ZN(_u10_u20_n2816 ) );
NAND2_X1 _u10_u20_U618  ( .A1(_u10_u20_n2815 ), .A2(_u10_u20_n2816 ), .ZN(_u10_u20_n2809 ) );
INV_X1 _u10_u20_U617  ( .A(_u10_u20_n2814 ), .ZN(_u10_u20_n2812 ) );
OR2_X1 _u10_u20_U616  ( .A1(_u10_u20_n1911 ), .A2(_u10_u20_n2813 ), .ZN(_u10_u20_n1884 ) );
NAND2_X1 _u10_u20_U615  ( .A1(_u10_u20_n2812 ), .A2(_u10_u20_n1884 ), .ZN(_u10_u20_n2810 ) );
NOR2_X1 _u10_u20_U614  ( .A1(_u10_u20_n1894 ), .A2(_u10_u20_n2461 ), .ZN(_u10_u20_n1948 ) );
OR2_X1 _u10_u20_U613  ( .A1(_u10_u20_n1847 ), .A2(_u10_u20_n1948 ), .ZN(_u10_u20_n2811 ) );
NAND3_X1 _u10_u20_U612  ( .A1(_u10_u20_n2809 ), .A2(_u10_u20_n2810 ), .A3(_u10_u20_n2811 ), .ZN(_u10_u20_n2805 ) );
NOR2_X1 _u10_u20_U611  ( .A1(_u10_u20_n2808 ), .A2(_u10_u20_n2775 ), .ZN(_u10_u20_n2806 ) );
AND2_X1 _u10_u20_U610  ( .A1(_u10_u20_n2721 ), .A2(_u10_u20_n1911 ), .ZN(_u10_u20_n2807 ) );
NOR4_X1 _u10_u20_U609  ( .A1(_u10_u20_n2804 ), .A2(_u10_u20_n2805 ), .A3(_u10_u20_n2806 ), .A4(_u10_u20_n2807 ), .ZN(_u10_u20_n2726 ) );
NAND2_X1 _u10_u20_U608  ( .A1(_u10_u20_n2803 ), .A2(_u10_u20_n2112 ), .ZN(_u10_u20_n2802 ) );
NAND2_X1 _u10_u20_U607  ( .A1(_u10_u20_n2364 ), .A2(_u10_u20_n2802 ), .ZN(_u10_u20_n2801 ) );
NAND2_X1 _u10_u20_U606  ( .A1(_u10_u20_n2800 ), .A2(_u10_u20_n2801 ), .ZN(_u10_u20_n2799 ) );
NAND2_X1 _u10_u20_U605  ( .A1(_u10_u20_n1937 ), .A2(_u10_u20_n2799 ), .ZN(_u10_u20_n2780 ) );
NAND2_X1 _u10_u20_U604  ( .A1(_u10_u20_n2775 ), .A2(_u10_u20_n2798 ), .ZN(_u10_u20_n2796 ) );
INV_X1 _u10_u20_U603  ( .A(_u10_u20_n2131 ), .ZN(_u10_u20_n2797 ) );
NAND2_X1 _u10_u20_U602  ( .A1(_u10_u20_n2796 ), .A2(_u10_u20_n2797 ), .ZN(_u10_u20_n2781 ) );
OR4_X1 _u10_u20_U601  ( .A1(_u10_u20_n2795 ), .A2(_u10_u20_n2303 ), .A3(_u10_u20_n2553 ), .A4(_u10_u20_n2554 ), .ZN(_u10_u20_n2792 ) );
NAND3_X1 _u10_u20_U600  ( .A1(_u10_u20_n1847 ), .A2(_u10_u20_n2097 ), .A3(_u10_u20_n2096 ), .ZN(_u10_u20_n2793 ) );
NOR4_X1 _u10_u20_U599  ( .A1(_u10_u20_n2792 ), .A2(_u10_u20_n2793 ), .A3(_u10_u20_n2542 ), .A4(_u10_u20_n2794 ), .ZN(_u10_u20_n2791 ) );
NOR2_X1 _u10_u20_U598  ( .A1(_u10_u20_n2791 ), .A2(_u10_u20_n2085 ), .ZN(_u10_u20_n2783 ) );
NAND2_X1 _u10_u20_U597  ( .A1(_u10_u20_n2114 ), .A2(_u10_u20_n2049 ), .ZN(_u10_u20_n2700 ) );
INV_X1 _u10_u20_U596  ( .A(_u10_u20_n2700 ), .ZN(_u10_u20_n2784 ) );
NAND4_X1 _u10_u20_U595  ( .A1(_u10_u20_n2001 ), .A2(_u10_u20_n2547 ), .A3(_u10_u20_n2368 ), .A4(_u10_u20_n1847 ), .ZN(_u10_u20_n2787 ) );
NOR4_X1 _u10_u20_U594  ( .A1(_u10_u20_n2787 ), .A2(_u10_u20_n2788 ), .A3(_u10_u20_n2789 ), .A4(_u10_u20_n2790 ), .ZN(_u10_u20_n2786 ) );
NOR2_X1 _u10_u20_U593  ( .A1(_u10_u20_n2786 ), .A2(_u10_u20_n2000 ), .ZN(_u10_u20_n2785 ) );
NOR3_X1 _u10_u20_U592  ( .A1(_u10_u20_n2783 ), .A2(_u10_u20_n2784 ), .A3(_u10_u20_n2785 ), .ZN(_u10_u20_n2782 ) );
NAND3_X1 _u10_u20_U591  ( .A1(_u10_u20_n2780 ), .A2(_u10_u20_n2781 ), .A3(_u10_u20_n2782 ), .ZN(_u10_u20_n2728 ) );
OR3_X1 _u10_u20_U590  ( .A1(_u10_u20_n2138 ), .A2(_u10_u20_n2633 ), .A3(_u10_u20_n2779 ), .ZN(_u10_u20_n2778 ) );
NAND2_X1 _u10_u20_U589  ( .A1(_u10_u20_n2777 ), .A2(_u10_u20_n2778 ), .ZN(_u10_u20_n2767 ) );
NAND3_X1 _u10_u20_U588  ( .A1(_u10_u20_n2775 ), .A2(_u10_u20_n2083 ), .A3(_u10_u20_n2776 ), .ZN(_u10_u20_n2774 ) );
NAND2_X1 _u10_u20_U587  ( .A1(_u10_u20_n2773 ), .A2(_u10_u20_n2774 ), .ZN(_u10_u20_n2768 ) );
NAND2_X1 _u10_u20_U586  ( .A1(_u10_u20_n2218 ), .A2(_u10_u20_n2772 ), .ZN(_u10_u20_n2769 ) );
NAND2_X1 _u10_u20_U585  ( .A1(_u10_u20_n2302 ), .A2(_u10_u20_n2467 ), .ZN(_u10_u20_n2771 ) );
NAND2_X1 _u10_u20_U584  ( .A1(_u10_u20_n2461 ), .A2(_u10_u20_n2771 ), .ZN(_u10_u20_n2770 ) );
NAND4_X1 _u10_u20_U583  ( .A1(_u10_u20_n2767 ), .A2(_u10_u20_n2768 ), .A3(_u10_u20_n2769 ), .A4(_u10_u20_n2770 ), .ZN(_u10_u20_n2729 ) );
NAND3_X1 _u10_u20_U582  ( .A1(_u10_u20_n2668 ), .A2(_u10_u20_n2600 ), .A3(_u10_u20_n2276 ), .ZN(_u10_u20_n2766 ) );
NAND2_X1 _u10_u20_U581  ( .A1(_u10_u20_n1894 ), .A2(_u10_u20_n2766 ), .ZN(_u10_u20_n2753 ) );
NAND3_X1 _u10_u20_U580  ( .A1(_u10_u20_n2456 ), .A2(_u10_u20_n2744 ), .A3(_u10_u20_n2765 ), .ZN(_u10_u20_n2764 ) );
NAND2_X1 _u10_u20_U579  ( .A1(_u10_u20_n2377 ), .A2(_u10_u20_n2764 ), .ZN(_u10_u20_n2754 ) );
NAND2_X1 _u10_u20_U578  ( .A1(_u10_u20_n2763 ), .A2(_u10_u20_n2007 ), .ZN(_u10_u20_n2755 ) );
NOR2_X1 _u10_u20_U577  ( .A1(_u10_u20_n2531 ), .A2(_u10_u20_n2744 ), .ZN(_u10_u20_n2760 ) );
INV_X1 _u10_u20_U576  ( .A(_u10_u20_n2762 ), .ZN(_u10_u20_n2189 ) );
NOR3_X1 _u10_u20_U575  ( .A1(_u10_u20_n2760 ), .A2(_u10_u20_n2761 ), .A3(_u10_u20_n2189 ), .ZN(_u10_u20_n2759 ) );
NOR2_X1 _u10_u20_U574  ( .A1(_u10_u20_n2759 ), .A2(_u10_u20_n1849 ), .ZN(_u10_u20_n2757 ) );
NOR2_X1 _u10_u20_U573  ( .A1(_u10_u20_n1817 ), .A2(_u10_u20_n2665 ), .ZN(_u10_u20_n2758 ) );
NOR2_X1 _u10_u20_U572  ( .A1(_u10_u20_n2757 ), .A2(_u10_u20_n2758 ), .ZN(_u10_u20_n2756 ) );
NAND4_X1 _u10_u20_U571  ( .A1(_u10_u20_n2753 ), .A2(_u10_u20_n2754 ), .A3(_u10_u20_n2755 ), .A4(_u10_u20_n2756 ), .ZN(_u10_u20_n2730 ) );
INV_X1 _u10_u20_U570  ( .A(_u10_u20_n2359 ), .ZN(_u10_u20_n1899 ) );
NAND4_X1 _u10_u20_U569  ( .A1(_u10_u20_n2078 ), .A2(_u10_u20_n2580 ), .A3(_u10_u20_n2748 ), .A4(_u10_u20_n2752 ), .ZN(_u10_u20_n2751 ) );
NAND2_X1 _u10_u20_U568  ( .A1(_u10_u20_n1899 ), .A2(_u10_u20_n2751 ), .ZN(_u10_u20_n2732 ) );
INV_X1 _u10_u20_U567  ( .A(_u10_u20_n2750 ), .ZN(_u10_u20_n2379 ) );
NAND3_X1 _u10_u20_U566  ( .A1(_u10_u20_n1856 ), .A2(_u10_u20_n2669 ), .A3(_u10_u20_n2364 ), .ZN(_u10_u20_n2749 ) );
AND2_X1 _u10_u20_U565  ( .A1(_u10_u20_n2748 ), .A2(_u10_u20_n2749 ), .ZN(_u10_u20_n2034 ) );
NAND2_X1 _u10_u20_U564  ( .A1(_u10_u20_n2105 ), .A2(_u10_u20_n2669 ), .ZN(_u10_u20_n2745 ) );
AND3_X1 _u10_u20_U563  ( .A1(_u10_u20_n2745 ), .A2(_u10_u20_n2746 ), .A3(_u10_u20_n2747 ), .ZN(_u10_u20_n2380 ) );
NOR2_X1 _u10_u20_U562  ( .A1(_u10_u20_n2274 ), .A2(_u10_u20_n2744 ), .ZN(_u10_u20_n2743 ) );
NOR4_X1 _u10_u20_U561  ( .A1(_u10_u20_n2742 ), .A2(_u10_u20_n2680 ), .A3(_u10_u20_n2743 ), .A4(_u10_u20_n2428 ), .ZN(_u10_u20_n2741 ) );
NAND4_X1 _u10_u20_U560  ( .A1(_u10_u20_n2379 ), .A2(_u10_u20_n2034 ), .A3(_u10_u20_n2380 ), .A4(_u10_u20_n2741 ), .ZN(_u10_u20_n2740 ) );
NAND2_X1 _u10_u20_U559  ( .A1(_u10_u20_n1967 ), .A2(_u10_u20_n2740 ), .ZN(_u10_u20_n2733 ) );
NAND3_X1 _u10_u20_U558  ( .A1(_u10_u20_n2739 ), .A2(_u10_u20_n2368 ), .A3(_u10_u20_n2255 ), .ZN(_u10_u20_n2738 ) );
NAND2_X1 _u10_u20_U557  ( .A1(_u10_u20_n2737 ), .A2(_u10_u20_n2738 ), .ZN(_u10_u20_n2734 ) );
NAND2_X1 _u10_u20_U556  ( .A1(_u10_u20_n2736 ), .A2(_u10_u20_n2524 ), .ZN(_u10_u20_n2735 ) );
NAND4_X1 _u10_u20_U555  ( .A1(_u10_u20_n2732 ), .A2(_u10_u20_n2733 ), .A3(_u10_u20_n2734 ), .A4(_u10_u20_n2735 ), .ZN(_u10_u20_n2731 ) );
NOR4_X1 _u10_u20_U554  ( .A1(_u10_u20_n2728 ), .A2(_u10_u20_n2729 ), .A3(_u10_u20_n2730 ), .A4(_u10_u20_n2731 ), .ZN(_u10_u20_n2727 ) );
NAND4_X1 _u10_u20_U553  ( .A1(_u10_u20_n2724 ), .A2(_u10_u20_n2725 ), .A3(_u10_u20_n2726 ), .A4(_u10_u20_n2727 ), .ZN(_u10_u20_n2723 ) );
MUX2_X1 _u10_u20_U552  ( .A(_u10_u20_n2723 ), .B(_u10_SYNOPSYS_UNCONNECTED_4 ), .S(_u10_u20_n1819 ), .Z(_u10_u20_n1809 ) );
NAND2_X1 _u10_u20_U551  ( .A1(_u10_u20_n2002 ), .A2(_u10_u20_n2722 ), .ZN(_u10_u20_n2713 ) );
NAND2_X1 _u10_u20_U550  ( .A1(_u10_u20_n2720 ), .A2(_u10_u20_n2721 ), .ZN(_u10_u20_n2714 ) );
NAND2_X1 _u10_u20_U549  ( .A1(_u10_u20_n2256 ), .A2(_u10_u20_n2719 ), .ZN(_u10_u20_n2715 ) );
NOR2_X1 _u10_u20_U548  ( .A1(_u10_u20_n2106 ), .A2(_u10_u20_n2037 ), .ZN(_u10_u20_n2717 ) );
AND2_X1 _u10_u20_U547  ( .A1(_u10_u20_n1966 ), .A2(_u10_u20_n2054 ), .ZN(_u10_u20_n2718 ) );
NOR2_X1 _u10_u20_U546  ( .A1(_u10_u20_n2717 ), .A2(_u10_u20_n2718 ), .ZN(_u10_u20_n2716 ) );
NAND4_X1 _u10_u20_U545  ( .A1(_u10_u20_n2713 ), .A2(_u10_u20_n2714 ), .A3(_u10_u20_n2715 ), .A4(_u10_u20_n2716 ), .ZN(_u10_u20_n2608 ) );
NAND2_X1 _u10_u20_U544  ( .A1(1'b0), .A2(_u10_u20_n2669 ), .ZN(_u10_u20_n2385 ) );
INV_X1 _u10_u20_U543  ( .A(_u10_u20_n2385 ), .ZN(_u10_u20_n1977 ) );
NAND2_X1 _u10_u20_U542  ( .A1(_u10_u20_n1977 ), .A2(_u10_u20_n2668 ), .ZN(_u10_u20_n2712 ) );
NAND2_X1 _u10_u20_U541  ( .A1(_u10_u20_n2712 ), .A2(_u10_u20_n2092 ), .ZN(_u10_u20_n1844 ) );
NAND2_X1 _u10_u20_U540  ( .A1(_u10_u20_n1894 ), .A2(_u10_u20_n1844 ), .ZN(_u10_u20_n2705 ) );
NAND2_X1 _u10_u20_U539  ( .A1(_u10_u20_n1894 ), .A2(_u10_u20_n2305 ), .ZN(_u10_u20_n2711 ) );
NAND2_X1 _u10_u20_U538  ( .A1(_u10_u20_n2711 ), .A2(_u10_u20_n2025 ), .ZN(_u10_u20_n1932 ) );
NAND2_X1 _u10_u20_U537  ( .A1(_u10_u20_n2710 ), .A2(_u10_u20_n1932 ), .ZN(_u10_u20_n2706 ) );
NAND2_X1 _u10_u20_U536  ( .A1(_u10_u20_n2708 ), .A2(_u10_u20_n2709 ), .ZN(_u10_u20_n2707 ) );
NAND3_X1 _u10_u20_U535  ( .A1(_u10_u20_n2705 ), .A2(_u10_u20_n2706 ), .A3(_u10_u20_n2707 ), .ZN(_u10_u20_n2701 ) );
NOR2_X1 _u10_u20_U534  ( .A1(_u10_u20_n1843 ), .A2(_u10_u20_n2545 ), .ZN(_u10_u20_n2702 ) );
NOR2_X1 _u10_u20_U533  ( .A1(_u10_u20_n2346 ), .A2(_u10_u20_n2700 ), .ZN(_u10_u20_n2703 ) );
NOR2_X1 _u10_u20_U532  ( .A1(_u10_u20_n2000 ), .A2(_u10_u20_n1887 ), .ZN(_u10_u20_n2704 ) );
NOR4_X1 _u10_u20_U531  ( .A1(_u10_u20_n2701 ), .A2(_u10_u20_n2702 ), .A3(_u10_u20_n2703 ), .A4(_u10_u20_n2704 ), .ZN(_u10_u20_n2671 ) );
NAND2_X1 _u10_u20_U530  ( .A1(_u10_u20_n2699 ), .A2(_u10_u20_n2700 ), .ZN(_u10_u20_n2698 ) );
NAND2_X1 _u10_u20_U529  ( .A1(_u10_u20_n2063 ), .A2(_u10_u20_n2698 ), .ZN(_u10_u20_n2682 ) );
NAND2_X1 _u10_u20_U528  ( .A1(_u10_u20_n2697 ), .A2(_u10_u20_n2103 ), .ZN(_u10_u20_n2696 ) );
NAND2_X1 _u10_u20_U527  ( .A1(_u10_u20_n2695 ), .A2(_u10_u20_n2696 ), .ZN(_u10_u20_n2694 ) );
NAND2_X1 _u10_u20_U526  ( .A1(_u10_u20_n1937 ), .A2(_u10_u20_n2694 ), .ZN(_u10_u20_n2683 ) );
INV_X1 _u10_u20_U525  ( .A(_u10_u20_n2693 ), .ZN(_u10_u20_n2691 ) );
NAND3_X1 _u10_u20_U524  ( .A1(_u10_u20_n2103 ), .A2(_u10_u20_n2502 ), .A3(1'b0), .ZN(_u10_u20_n2692 ) );
NAND2_X1 _u10_u20_U523  ( .A1(_u10_u20_n2691 ), .A2(_u10_u20_n2692 ), .ZN(_u10_u20_n2690 ) );
NAND2_X1 _u10_u20_U522  ( .A1(_u10_u20_n2236 ), .A2(_u10_u20_n2690 ), .ZN(_u10_u20_n2684 ) );
NAND3_X1 _u10_u20_U521  ( .A1(_u10_u20_n2688 ), .A2(_u10_u20_n1913 ), .A3(_u10_u20_n2689 ), .ZN(_u10_u20_n2335 ) );
NAND3_X1 _u10_u20_U520  ( .A1(_u10_u20_n2536 ), .A2(_u10_u20_n2103 ), .A3(1'b0), .ZN(_u10_u20_n2052 ) );
NOR2_X1 _u10_u20_U519  ( .A1(_u10_u20_n2052 ), .A2(_u10_u20_n2687 ), .ZN(_u10_u20_n1851 ) );
NAND2_X1 _u10_u20_U518  ( .A1(_u10_u20_n1851 ), .A2(_u10_u20_n2078 ), .ZN(_u10_u20_n2582 ) );
NOR2_X1 _u10_u20_U517  ( .A1(_u10_u20_n2686 ), .A2(_u10_u20_n2582 ), .ZN(_u10_u20_n2094 ) );
NAND3_X1 _u10_u20_U516  ( .A1(_u10_u20_n2251 ), .A2(_u10_u20_n2335 ), .A3(_u10_u20_n2094 ), .ZN(_u10_u20_n2685 ) );
NAND4_X1 _u10_u20_U515  ( .A1(_u10_u20_n2682 ), .A2(_u10_u20_n2683 ), .A3(_u10_u20_n2684 ), .A4(_u10_u20_n2685 ), .ZN(_u10_u20_n2673 ) );
INV_X1 _u10_u20_U514  ( .A(_u10_u20_n2291 ), .ZN(_u10_u20_n2057 ) );
AND2_X1 _u10_u20_U513  ( .A1(_u10_u20_n1851 ), .A2(_u10_u20_n2057 ), .ZN(_u10_u20_n2674 ) );
INV_X1 _u10_u20_U512  ( .A(_u10_u20_n1874 ), .ZN(_u10_u20_n2681 ) );
NOR2_X1 _u10_u20_U511  ( .A1(_u10_u20_n2007 ), .A2(_u10_u20_n1911 ), .ZN(_u10_u20_n2486 ) );
NOR2_X1 _u10_u20_U510  ( .A1(_u10_u20_n2681 ), .A2(_u10_u20_n2486 ), .ZN(_u10_u20_n2675 ) );
NOR2_X1 _u10_u20_U509  ( .A1(_u10_u20_n1977 ), .A2(_u10_u20_n2680 ), .ZN(_u10_u20_n2679 ) );
NOR2_X1 _u10_u20_U508  ( .A1(_u10_u20_n2679 ), .A2(_u10_u20_n2030 ), .ZN(_u10_u20_n2678 ) );
NOR2_X1 _u10_u20_U507  ( .A1(_u10_u20_n2678 ), .A2(_u10_u20_n2094 ), .ZN(_u10_u20_n2677 ) );
NOR2_X1 _u10_u20_U506  ( .A1(_u10_u20_n2677 ), .A2(_u10_u20_n2025 ), .ZN(_u10_u20_n2676 ) );
NOR4_X1 _u10_u20_U505  ( .A1(_u10_u20_n2673 ), .A2(_u10_u20_n2674 ), .A3(_u10_u20_n2675 ), .A4(_u10_u20_n2676 ), .ZN(_u10_u20_n2672 ) );
AND2_X1 _u10_u20_U504  ( .A1(_u10_u20_n2671 ), .A2(_u10_u20_n2672 ), .ZN(_u10_u20_n1990 ) );
INV_X1 _u10_u20_U503  ( .A(_u10_u20_n2670 ), .ZN(_u10_u20_n2660 ) );
NAND4_X1 _u10_u20_U502  ( .A1(_u10_u20_n2251 ), .A2(_u10_u20_n2669 ), .A3(_u10_u20_n2162 ), .A4(_u10_u20_n2169 ), .ZN(_u10_u20_n2664 ) );
AND3_X1 _u10_u20_U501  ( .A1(_u10_u20_n1977 ), .A2(_u10_u20_n2668 ), .A3(_u10_u20_n2089 ), .ZN(_u10_u20_n2555 ) );
NAND2_X1 _u10_u20_U500  ( .A1(_u10_u20_n2555 ), .A2(_u10_u20_n2667 ), .ZN(_u10_u20_n2666 ) );
NAND3_X1 _u10_u20_U499  ( .A1(_u10_u20_n2664 ), .A2(_u10_u20_n2665 ), .A3(_u10_u20_n2666 ), .ZN(_u10_u20_n1988 ) );
INV_X1 _u10_u20_U498  ( .A(_u10_u20_n1988 ), .ZN(_u10_u20_n2661 ) );
NAND2_X1 _u10_u20_U497  ( .A1(1'b0), .A2(_u10_u20_n2043 ), .ZN(_u10_u20_n2662 ) );
NAND2_X1 _u10_u20_U496  ( .A1(_u10_u20_n2169 ), .A2(1'b0), .ZN(_u10_u20_n2663 ) );
NAND4_X1 _u10_u20_U495  ( .A1(_u10_u20_n2660 ), .A2(_u10_u20_n2661 ), .A3(_u10_u20_n2662 ), .A4(_u10_u20_n2663 ), .ZN(_u10_u20_n2650 ) );
NAND2_X1 _u10_u20_U494  ( .A1(_u10_u20_n2659 ), .A2(1'b0), .ZN(_u10_u20_n2193 ) );
INV_X1 _u10_u20_U493  ( .A(_u10_u20_n2193 ), .ZN(_u10_u20_n2143 ) );
NAND2_X1 _u10_u20_U492  ( .A1(_u10_u20_n2143 ), .A2(_u10_u20_n2036 ), .ZN(_u10_u20_n2286 ) );
INV_X1 _u10_u20_U491  ( .A(_u10_u20_n2286 ), .ZN(_u10_u20_n2577 ) );
NAND2_X1 _u10_u20_U490  ( .A1(_u10_u20_n2577 ), .A2(_u10_u20_n2278 ), .ZN(_u10_u20_n2474 ) );
INV_X1 _u10_u20_U489  ( .A(_u10_u20_n2474 ), .ZN(_u10_u20_n2306 ) );
NAND2_X1 _u10_u20_U488  ( .A1(_u10_u20_n2306 ), .A2(_u10_u20_n2251 ), .ZN(_u10_u20_n2654 ) );
NAND2_X1 _u10_u20_U487  ( .A1(_u10_u20_n2649 ), .A2(_u10_u20_n2658 ), .ZN(_u10_u20_n2655 ) );
NAND2_X1 _u10_u20_U486  ( .A1(_u10_u20_n2657 ), .A2(_u10_u20_n2445 ), .ZN(_u10_u20_n2656 ) );
NAND3_X1 _u10_u20_U485  ( .A1(_u10_u20_n2654 ), .A2(_u10_u20_n2655 ), .A3(_u10_u20_n2656 ), .ZN(_u10_u20_n2651 ) );
NOR2_X1 _u10_u20_U484  ( .A1(_u10_u20_n2366 ), .A2(_u10_u20_n2376 ), .ZN(_u10_u20_n2652 ) );
AND2_X1 _u10_u20_U483  ( .A1(_u10_u20_n1966 ), .A2(_u10_u20_n2528 ), .ZN(_u10_u20_n2653 ) );
NOR4_X1 _u10_u20_U482  ( .A1(_u10_u20_n2650 ), .A2(_u10_u20_n2651 ), .A3(_u10_u20_n2652 ), .A4(_u10_u20_n2653 ), .ZN(_u10_u20_n2613 ) );
NAND2_X1 _u10_u20_U481  ( .A1(_u10_u20_n1891 ), .A2(1'b0), .ZN(_u10_u20_n2636 ) );
NAND2_X1 _u10_u20_U480  ( .A1(_u10_u20_n1868 ), .A2(_u10_u20_n2113 ), .ZN(_u10_u20_n2101 ) );
NOR4_X1 _u10_u20_U479  ( .A1(_u10_u20_n2649 ), .A2(_u10_u20_n2216 ), .A3(_u10_u20_n2101 ), .A4(_u10_u20_n2634 ), .ZN(_u10_u20_n2648 ) );
NOR2_X1 _u10_u20_U478  ( .A1(_u10_u20_n2648 ), .A2(_u10_u20_n2254 ), .ZN(_u10_u20_n2638 ) );
NOR2_X1 _u10_u20_U477  ( .A1(_u10_u20_n2106 ), .A2(_u10_u20_n2643 ), .ZN(_u10_u20_n2645 ) );
NAND2_X1 _u10_u20_U476  ( .A1(1'b0), .A2(_u10_u20_n2049 ), .ZN(_u10_u20_n2647 ) );
NAND2_X1 _u10_u20_U475  ( .A1(_u10_u20_n2646 ), .A2(_u10_u20_n2647 ), .ZN(_u10_u20_n2348 ) );
NOR2_X1 _u10_u20_U474  ( .A1(_u10_u20_n2645 ), .A2(_u10_u20_n2348 ), .ZN(_u10_u20_n2644 ) );
NOR2_X1 _u10_u20_U473  ( .A1(_u10_u20_n2644 ), .A2(_u10_u20_n2495 ), .ZN(_u10_u20_n2639 ) );
NOR2_X1 _u10_u20_U472  ( .A1(_u10_u20_n2643 ), .A2(_u10_u20_n2203 ), .ZN(_u10_u20_n2642 ) );
NOR3_X1 _u10_u20_U471  ( .A1(_u10_u20_n2101 ), .A2(1'b0), .A3(_u10_u20_n2642 ), .ZN(_u10_u20_n2641 ) );
NOR2_X1 _u10_u20_U470  ( .A1(_u10_u20_n2641 ), .A2(_u10_u20_n2253 ), .ZN(_u10_u20_n2640 ) );
NOR3_X1 _u10_u20_U469  ( .A1(_u10_u20_n2638 ), .A2(_u10_u20_n2639 ), .A3(_u10_u20_n2640 ), .ZN(_u10_u20_n2637 ) );
NAND3_X1 _u10_u20_U468  ( .A1(_u10_u20_n2635 ), .A2(_u10_u20_n2636 ), .A3(_u10_u20_n2637 ), .ZN(_u10_u20_n2615 ) );
NOR3_X1 _u10_u20_U467  ( .A1(_u10_u20_n2174 ), .A2(_u10_u20_n2175 ), .A3(_u10_u20_n2179 ), .ZN(_u10_u20_n2631 ) );
NAND3_X1 _u10_u20_U466  ( .A1(_u10_u20_n2223 ), .A2(_u10_u20_n2236 ), .A3(_u10_u20_n2631 ), .ZN(_u10_u20_n2622 ) );
OR2_X1 _u10_u20_U465  ( .A1(_u10_u20_n1960 ), .A2(_u10_u20_n1959 ), .ZN(_u10_u20_n2625 ) );
NOR3_X1 _u10_u20_U464  ( .A1(_u10_u20_n2101 ), .A2(_u10_u20_n2633 ), .A3(_u10_u20_n2634 ), .ZN(_u10_u20_n2523 ) );
OR2_X1 _u10_u20_U463  ( .A1(_u10_u20_n2632 ), .A2(_u10_u20_n2523 ), .ZN(_u10_u20_n2627 ) );
INV_X1 _u10_u20_U462  ( .A(_u10_u20_n2631 ), .ZN(_u10_u20_n2628 ) );
NAND2_X1 _u10_u20_U461  ( .A1(_u10_u20_n2630 ), .A2(_u10_u20_n1922 ), .ZN(_u10_u20_n2629 ) );
NAND3_X1 _u10_u20_U460  ( .A1(_u10_u20_n2627 ), .A2(_u10_u20_n2628 ), .A3(_u10_u20_n2629 ), .ZN(_u10_u20_n2626 ) );
NAND2_X1 _u10_u20_U459  ( .A1(_u10_u20_n2625 ), .A2(_u10_u20_n2626 ), .ZN(_u10_u20_n2624 ) );
NAND3_X1 _u10_u20_U458  ( .A1(_u10_u20_n2622 ), .A2(_u10_u20_n2623 ), .A3(_u10_u20_n2624 ), .ZN(_u10_u20_n2616 ) );
AND2_X1 _u10_u20_U457  ( .A1(_u10_u20_n2621 ), .A2(_u10_u20_n2358 ), .ZN(_u10_u20_n2620 ) );
NOR2_X1 _u10_u20_U456  ( .A1(_u10_u20_n2523 ), .A2(_u10_u20_n2620 ), .ZN(_u10_u20_n2617 ) );
INV_X1 _u10_u20_U455  ( .A(_u10_u20_n2101 ), .ZN(_u10_u20_n2221 ) );
NOR2_X1 _u10_u20_U454  ( .A1(_u10_u20_n1911 ), .A2(_u10_u20_n2488 ), .ZN(_u10_u20_n2619 ) );
NOR2_X1 _u10_u20_U453  ( .A1(_u10_u20_n2221 ), .A2(_u10_u20_n2619 ), .ZN(_u10_u20_n2618 ) );
NOR4_X1 _u10_u20_U452  ( .A1(_u10_u20_n2615 ), .A2(_u10_u20_n2616 ), .A3(_u10_u20_n2617 ), .A4(_u10_u20_n2618 ), .ZN(_u10_u20_n2614 ) );
AND2_X1 _u10_u20_U451  ( .A1(_u10_u20_n2613 ), .A2(_u10_u20_n2614 ), .ZN(_u10_u20_n2314 ) );
NAND3_X1 _u10_u20_U450  ( .A1(_u10_u20_n2612 ), .A2(_u10_u20_n1990 ), .A3(_u10_u20_n2314 ), .ZN(_u10_u20_n2609 ) );
NOR4_X1 _u10_u20_U449  ( .A1(_u10_u20_n2608 ), .A2(_u10_u20_n2609 ), .A3(_u10_u20_n2610 ), .A4(_u10_u20_n2611 ), .ZN(_u10_u20_n2388 ) );
NAND2_X1 _u10_u20_U448  ( .A1(_u10_u20_n2346 ), .A2(_u10_u20_n2607 ), .ZN(_u10_u20_n2191 ) );
NAND2_X1 _u10_u20_U447  ( .A1(_u10_u20_n2143 ), .A2(_u10_u20_n2191 ), .ZN(_u10_u20_n2556 ) );
INV_X1 _u10_u20_U446  ( .A(_u10_u20_n2348 ), .ZN(_u10_u20_n2603 ) );
NAND3_X1 _u10_u20_U445  ( .A1(_u10_u20_n2535 ), .A2(_u10_u20_n2485 ), .A3(_u10_u20_n2456 ), .ZN(_u10_u20_n2606 ) );
NAND2_X1 _u10_u20_U444  ( .A1(_u10_u20_n2049 ), .A2(_u10_u20_n2606 ), .ZN(_u10_u20_n2604 ) );
NAND3_X1 _u10_u20_U443  ( .A1(_u10_u20_n2603 ), .A2(_u10_u20_n2604 ), .A3(_u10_u20_n2605 ), .ZN(_u10_u20_n2602 ) );
NAND2_X1 _u10_u20_U442  ( .A1(_u10_u20_n2043 ), .A2(_u10_u20_n2602 ), .ZN(_u10_u20_n2557 ) );
INV_X1 _u10_u20_U441  ( .A(_u10_u20_n2601 ), .ZN(_u10_u20_n2590 ) );
NAND2_X1 _u10_u20_U440  ( .A1(_u10_u20_n2599 ), .A2(_u10_u20_n2600 ), .ZN(_u10_u20_n2597 ) );
NAND2_X1 _u10_u20_U439  ( .A1(_u10_u20_n2082 ), .A2(_u10_u20_n2101 ), .ZN(_u10_u20_n2598 ) );
AND2_X1 _u10_u20_U438  ( .A1(_u10_u20_n2597 ), .A2(_u10_u20_n2598 ), .ZN(_u10_u20_n2281 ) );
NAND3_X1 _u10_u20_U437  ( .A1(_u10_u20_n1969 ), .A2(_u10_u20_n2582 ), .A3(_u10_u20_n2281 ), .ZN(_u10_u20_n2073 ) );
INV_X1 _u10_u20_U436  ( .A(_u10_u20_n2073 ), .ZN(_u10_u20_n2591 ) );
NOR2_X1 _u10_u20_U435  ( .A1(_u10_u20_n1816 ), .A2(_u10_u20_n2077 ), .ZN(_u10_u20_n2595 ) );
NOR2_X1 _u10_u20_U434  ( .A1(_u10_u20_n2595 ), .A2(_u10_u20_n2596 ), .ZN(_u10_u20_n2592 ) );
NAND3_X1 _u10_u20_U433  ( .A1(_u10_u20_n2107 ), .A2(_u10_u20_n2536 ), .A3(1'b0), .ZN(_u10_u20_n2438 ) );
INV_X1 _u10_u20_U432  ( .A(_u10_u20_n2438 ), .ZN(_u10_u20_n2427 ) );
NOR4_X1 _u10_u20_U431  ( .A1(1'b0), .A2(_u10_u20_n2594 ), .A3(_u10_u20_n2577 ), .A4(_u10_u20_n2427 ), .ZN(_u10_u20_n2593 ) );
NAND4_X1 _u10_u20_U430  ( .A1(_u10_u20_n2590 ), .A2(_u10_u20_n2591 ), .A3(_u10_u20_n2592 ), .A4(_u10_u20_n2593 ), .ZN(_u10_u20_n2589 ) );
NAND2_X1 _u10_u20_U429  ( .A1(_u10_u20_n2279 ), .A2(_u10_u20_n2589 ), .ZN(_u10_u20_n2558 ) );
NAND3_X1 _u10_u20_U428  ( .A1(_u10_u20_n2587 ), .A2(_u10_u20_n2115 ), .A3(_u10_u20_n2588 ), .ZN(_u10_u20_n2585 ) );
NOR4_X1 _u10_u20_U427  ( .A1(_u10_u20_n2585 ), .A2(_u10_u20_n2586 ), .A3(1'b0), .A4(_u10_u20_n2114 ), .ZN(_u10_u20_n2583 ) );
NOR2_X1 _u10_u20_U426  ( .A1(_u10_u20_n2583 ), .A2(_u10_u20_n2584 ), .ZN(_u10_u20_n2560 ) );
OR2_X1 _u10_u20_U425  ( .A1(_u10_u20_n2582 ), .A2(1'b0), .ZN(_u10_u20_n2581 ) );
NAND2_X1 _u10_u20_U424  ( .A1(_u10_u20_n2580 ), .A2(_u10_u20_n2581 ), .ZN(_u10_u20_n1974 ) );
INV_X1 _u10_u20_U423  ( .A(_u10_u20_n1974 ), .ZN(_u10_u20_n1901 ) );
AND4_X1 _u10_u20_U422  ( .A1(_u10_u20_n1901 ), .A2(_u10_u20_n2385 ), .A3(_u10_u20_n2578 ), .A4(_u10_u20_n2579 ), .ZN(_u10_u20_n2424 ) );
NOR2_X1 _u10_u20_U421  ( .A1(1'b0), .A2(_u10_u20_n2424 ), .ZN(_u10_u20_n2574 ) );
NOR3_X1 _u10_u20_U420  ( .A1(_u10_u20_n2427 ), .A2(1'b0), .A3(_u10_u20_n2577 ), .ZN(_u10_u20_n2576 ) );
NOR2_X1 _u10_u20_U419  ( .A1(_u10_u20_n2576 ), .A2(_u10_u20_n1976 ), .ZN(_u10_u20_n2575 ) );
NOR3_X1 _u10_u20_U418  ( .A1(_u10_u20_n2574 ), .A2(_u10_u20_n1979 ), .A3(_u10_u20_n2575 ), .ZN(_u10_u20_n2572 ) );
NOR2_X1 _u10_u20_U417  ( .A1(_u10_u20_n2572 ), .A2(_u10_u20_n2573 ), .ZN(_u10_u20_n2561 ) );
INV_X1 _u10_u20_U416  ( .A(_u10_u20_n2061 ), .ZN(_u10_u20_n2453 ) );
NOR2_X1 _u10_u20_U415  ( .A1(_u10_u20_n2453 ), .A2(_u10_u20_n1851 ), .ZN(_u10_u20_n2018 ) );
NAND2_X1 _u10_u20_U414  ( .A1(1'b0), .A2(_u10_u20_n2571 ), .ZN(_u10_u20_n2570 ) );
NAND2_X1 _u10_u20_U413  ( .A1(_u10_u20_n2018 ), .A2(_u10_u20_n2570 ), .ZN(_u10_u20_n1837 ) );
INV_X1 _u10_u20_U412  ( .A(_u10_u20_n1837 ), .ZN(_u10_u20_n2568 ) );
NAND2_X1 _u10_u20_U411  ( .A1(1'b0), .A2(_u10_u20_n2536 ), .ZN(_u10_u20_n2569 ) );
NAND2_X1 _u10_u20_U410  ( .A1(_u10_u20_n2568 ), .A2(_u10_u20_n2569 ), .ZN(_u10_u20_n2564 ) );
NOR2_X1 _u10_u20_U409  ( .A1(_u10_u20_n1841 ), .A2(_u10_u20_n1868 ), .ZN(_u10_u20_n2565 ) );
INV_X1 _u10_u20_U408  ( .A(_u10_u20_n2567 ), .ZN(_u10_u20_n2566 ) );
NOR4_X1 _u10_u20_U407  ( .A1(_u10_u20_n2564 ), .A2(_u10_u20_n2565 ), .A3(_u10_u20_n2143 ), .A4(_u10_u20_n2566 ), .ZN(_u10_u20_n2563 ) );
NOR2_X1 _u10_u20_U406  ( .A1(_u10_u20_n2563 ), .A2(_u10_u20_n2014 ), .ZN(_u10_u20_n2562 ) );
NOR3_X1 _u10_u20_U405  ( .A1(_u10_u20_n2560 ), .A2(_u10_u20_n2561 ), .A3(_u10_u20_n2562 ), .ZN(_u10_u20_n2559 ) );
NAND4_X1 _u10_u20_U404  ( .A1(_u10_u20_n2556 ), .A2(_u10_u20_n2557 ), .A3(_u10_u20_n2558 ), .A4(_u10_u20_n2559 ), .ZN(_u10_u20_n2511 ) );
INV_X1 _u10_u20_U403  ( .A(_u10_u20_n2085 ), .ZN(_u10_u20_n2293 ) );
NOR2_X1 _u10_u20_U402  ( .A1(_u10_u20_n2554 ), .A2(_u10_u20_n2555 ), .ZN(_u10_u20_n2444 ) );
NAND2_X1 _u10_u20_U401  ( .A1(_u10_u20_n2553 ), .A2(_u10_u20_n2549 ), .ZN(_u10_u20_n2552 ) );
AND2_X1 _u10_u20_U400  ( .A1(_u10_u20_n2444 ), .A2(_u10_u20_n2552 ), .ZN(_u10_u20_n2295 ) );
NAND2_X1 _u10_u20_U399  ( .A1(_u10_u20_n2551 ), .A2(_u10_u20_n2549 ), .ZN(_u10_u20_n2538 ) );
AND2_X1 _u10_u20_U398  ( .A1(_u10_u20_n2427 ), .A2(_u10_u20_n2108 ), .ZN(_u10_u20_n2460 ) );
NOR4_X1 _u10_u20_U397  ( .A1(_u10_u20_n2460 ), .A2(_u10_u20_n2306 ), .A3(_u10_u20_n2094 ), .A4(_u10_u20_n2550 ), .ZN(_u10_u20_n2409 ) );
INV_X1 _u10_u20_U396  ( .A(_u10_u20_n2409 ), .ZN(_u10_u20_n2407 ) );
NAND2_X1 _u10_u20_U395  ( .A1(_u10_u20_n2549 ), .A2(_u10_u20_n2407 ), .ZN(_u10_u20_n2546 ) );
NAND3_X1 _u10_u20_U394  ( .A1(_u10_u20_n2546 ), .A2(_u10_u20_n2547 ), .A3(_u10_u20_n2548 ), .ZN(_u10_u20_n2501 ) );
INV_X1 _u10_u20_U393  ( .A(_u10_u20_n2501 ), .ZN(_u10_u20_n2539 ) );
NOR2_X1 _u10_u20_U392  ( .A1(1'b0), .A2(_u10_u20_n2545 ), .ZN(_u10_u20_n2541 ) );
AND2_X1 _u10_u20_U391  ( .A1(_u10_u20_n2544 ), .A2(_u10_u20_n2089 ), .ZN(_u10_u20_n2543 ) );
NOR3_X1 _u10_u20_U390  ( .A1(_u10_u20_n2541 ), .A2(_u10_u20_n2542 ), .A3(_u10_u20_n2543 ), .ZN(_u10_u20_n2540 ) );
NAND4_X1 _u10_u20_U389  ( .A1(_u10_u20_n2295 ), .A2(_u10_u20_n2538 ), .A3(_u10_u20_n2539 ), .A4(_u10_u20_n2540 ), .ZN(_u10_u20_n2537 ) );
NAND2_X1 _u10_u20_U388  ( .A1(_u10_u20_n2293 ), .A2(_u10_u20_n2537 ), .ZN(_u10_u20_n2515 ) );
NAND2_X1 _u10_u20_U387  ( .A1(_u10_u20_n2536 ), .A2(_u10_u20_n2508 ), .ZN(_u10_u20_n2526 ) );
NAND2_X1 _u10_u20_U386  ( .A1(_u10_u20_n2535 ), .A2(_u10_u20_n1940 ), .ZN(_u10_u20_n2532 ) );
NOR4_X1 _u10_u20_U385  ( .A1(_u10_u20_n2532 ), .A2(_u10_u20_n2533 ), .A3(1'b0), .A4(_u10_u20_n2534 ), .ZN(_u10_u20_n2530 ) );
NOR2_X1 _u10_u20_U384  ( .A1(_u10_u20_n2530 ), .A2(_u10_u20_n2531 ), .ZN(_u10_u20_n2529 ) );
NOR4_X1 _u10_u20_U383  ( .A1(_u10_u20_n2528 ), .A2(_u10_u20_n2143 ), .A3(_u10_u20_n2189 ), .A4(_u10_u20_n2529 ), .ZN(_u10_u20_n2527 ) );
NAND4_X1 _u10_u20_U382  ( .A1(_u10_u20_n2019 ), .A2(_u10_u20_n2526 ), .A3(_u10_u20_n2018 ), .A4(_u10_u20_n2527 ), .ZN(_u10_u20_n2525 ) );
NAND2_X1 _u10_u20_U381  ( .A1(_u10_u20_n2183 ), .A2(_u10_u20_n2525 ), .ZN(_u10_u20_n2516 ) );
INV_X1 _u10_u20_U380  ( .A(_u10_u20_n2524 ), .ZN(_u10_u20_n2396 ) );
NAND2_X1 _u10_u20_U379  ( .A1(_u10_u20_n2396 ), .A2(_u10_u20_n2523 ), .ZN(_u10_u20_n2522 ) );
NAND2_X1 _u10_u20_U378  ( .A1(_u10_u20_n1866 ), .A2(_u10_u20_n2522 ), .ZN(_u10_u20_n2519 ) );
AND2_X1 _u10_u20_U377  ( .A1(_u10_u20_n2493 ), .A2(_u10_u20_n1961 ), .ZN(_u10_u20_n2429 ) );
NAND2_X1 _u10_u20_U376  ( .A1(_u10_u20_n2429 ), .A2(_u10_u20_n2175 ), .ZN(_u10_u20_n2510 ) );
NAND2_X1 _u10_u20_U375  ( .A1(_u10_u20_n2510 ), .A2(_u10_u20_n1864 ), .ZN(_u10_u20_n2521 ) );
NAND3_X1 _u10_u20_U374  ( .A1(_u10_u20_n2519 ), .A2(_u10_u20_n2520 ), .A3(_u10_u20_n2521 ), .ZN(_u10_u20_n2518 ) );
NAND2_X1 _u10_u20_U373  ( .A1(_u10_u20_n1861 ), .A2(_u10_u20_n2518 ), .ZN(_u10_u20_n2517 ) );
NAND3_X1 _u10_u20_U372  ( .A1(_u10_u20_n2515 ), .A2(_u10_u20_n2516 ), .A3(_u10_u20_n2517 ), .ZN(_u10_u20_n2512 ) );
NOR2_X1 _u10_u20_U371  ( .A1(_u10_u20_n1913 ), .A2(_u10_u20_n1940 ), .ZN(_u10_u20_n2513 ) );
NOR2_X1 _u10_u20_U370  ( .A1(_u10_u20_n2113 ), .A2(_u10_u20_n2350 ), .ZN(_u10_u20_n2514 ) );
NOR4_X1 _u10_u20_U369  ( .A1(_u10_u20_n2511 ), .A2(_u10_u20_n2512 ), .A3(_u10_u20_n2513 ), .A4(_u10_u20_n2514 ), .ZN(_u10_u20_n2389 ) );
NAND2_X1 _u10_u20_U368  ( .A1(_u10_u20_n2509 ), .A2(_u10_u20_n2510 ), .ZN(_u10_u20_n2477 ) );
NAND2_X1 _u10_u20_U367  ( .A1(_u10_u20_n2507 ), .A2(_u10_u20_n2508 ), .ZN(_u10_u20_n2504 ) );
NAND2_X1 _u10_u20_U366  ( .A1(1'b0), .A2(_u10_u20_n2506 ), .ZN(_u10_u20_n2505 ) );
NAND2_X1 _u10_u20_U365  ( .A1(_u10_u20_n2504 ), .A2(_u10_u20_n2505 ), .ZN(_u10_u20_n2503 ) );
NAND2_X1 _u10_u20_U364  ( .A1(_u10_u20_n2502 ), .A2(_u10_u20_n2503 ), .ZN(_u10_u20_n2478 ) );
NAND2_X1 _u10_u20_U363  ( .A1(_u10_u20_n2501 ), .A2(_u10_u20_n2446 ), .ZN(_u10_u20_n2497 ) );
INV_X1 _u10_u20_U362  ( .A(_u10_u20_n2500 ), .ZN(_u10_u20_n2499 ) );
NAND3_X1 _u10_u20_U361  ( .A1(_u10_u20_n2497 ), .A2(_u10_u20_n2498 ), .A3(_u10_u20_n2499 ), .ZN(_u10_u20_n2496 ) );
NAND2_X1 _u10_u20_U360  ( .A1(_u10_u20_n2445 ), .A2(_u10_u20_n2496 ), .ZN(_u10_u20_n2479 ) );
NOR2_X1 _u10_u20_U359  ( .A1(_u10_u20_n2429 ), .A2(_u10_u20_n2495 ), .ZN(_u10_u20_n2491 ) );
INV_X1 _u10_u20_U358  ( .A(_u10_u20_n2191 ), .ZN(_u10_u20_n2494 ) );
NOR2_X1 _u10_u20_U357  ( .A1(_u10_u20_n2493 ), .A2(_u10_u20_n2494 ), .ZN(_u10_u20_n2492 ) );
NOR2_X1 _u10_u20_U356  ( .A1(_u10_u20_n2491 ), .A2(_u10_u20_n2492 ), .ZN(_u10_u20_n2489 ) );
NOR2_X1 _u10_u20_U355  ( .A1(_u10_u20_n2489 ), .A2(_u10_u20_n2490 ), .ZN(_u10_u20_n2481 ) );
NAND2_X1 _u10_u20_U354  ( .A1(_u10_u20_n2253 ), .A2(_u10_u20_n1859 ), .ZN(_u10_u20_n2398 ) );
NOR2_X1 _u10_u20_U353  ( .A1(_u10_u20_n2488 ), .A2(_u10_u20_n2398 ), .ZN(_u10_u20_n2487 ) );
NOR2_X1 _u10_u20_U352  ( .A1(_u10_u20_n2220 ), .A2(_u10_u20_n2487 ), .ZN(_u10_u20_n2482 ) );
AND2_X1 _u10_u20_U351  ( .A1(_u10_u20_n2350 ), .A2(_u10_u20_n2486 ), .ZN(_u10_u20_n2484 ) );
NOR2_X1 _u10_u20_U350  ( .A1(_u10_u20_n2484 ), .A2(_u10_u20_n2485 ), .ZN(_u10_u20_n2483 ) );
NOR3_X1 _u10_u20_U349  ( .A1(_u10_u20_n2481 ), .A2(_u10_u20_n2482 ), .A3(_u10_u20_n2483 ), .ZN(_u10_u20_n2480 ) );
NAND4_X1 _u10_u20_U348  ( .A1(_u10_u20_n2477 ), .A2(_u10_u20_n2478 ), .A3(_u10_u20_n2479 ), .A4(_u10_u20_n2480 ), .ZN(_u10_u20_n2447 ) );
NAND2_X1 _u10_u20_U347  ( .A1(_u10_u20_n2476 ), .A2(_u10_u20_n1936 ), .ZN(_u10_u20_n2472 ) );
NAND2_X1 _u10_u20_U346  ( .A1(_u10_u20_n2427 ), .A2(_u10_u20_n2278 ), .ZN(_u10_u20_n2473 ) );
NAND4_X1 _u10_u20_U345  ( .A1(_u10_u20_n2472 ), .A2(_u10_u20_n2473 ), .A3(_u10_u20_n2474 ), .A4(_u10_u20_n2475 ), .ZN(_u10_u20_n2471 ) );
NAND2_X1 _u10_u20_U344  ( .A1(_u10_u20_n2470 ), .A2(_u10_u20_n2471 ), .ZN(_u10_u20_n2457 ) );
NAND2_X1 _u10_u20_U343  ( .A1(_u10_u20_n2409 ), .A2(_u10_u20_n2469 ), .ZN(_u10_u20_n2468 ) );
NAND2_X1 _u10_u20_U342  ( .A1(_u10_u20_n2467 ), .A2(_u10_u20_n2468 ), .ZN(_u10_u20_n2463 ) );
NAND2_X1 _u10_u20_U341  ( .A1(_u10_u20_n1844 ), .A2(_u10_u20_n2466 ), .ZN(_u10_u20_n2465 ) );
NAND3_X1 _u10_u20_U340  ( .A1(_u10_u20_n2463 ), .A2(_u10_u20_n2464 ), .A3(_u10_u20_n2465 ), .ZN(_u10_u20_n2462 ) );
NAND2_X1 _u10_u20_U339  ( .A1(_u10_u20_n2461 ), .A2(_u10_u20_n2462 ), .ZN(_u10_u20_n2458 ) );
NAND2_X1 _u10_u20_U338  ( .A1(_u10_u20_n2460 ), .A2(_u10_u20_n2251 ), .ZN(_u10_u20_n2459 ) );
NAND3_X1 _u10_u20_U337  ( .A1(_u10_u20_n2457 ), .A2(_u10_u20_n2458 ), .A3(_u10_u20_n2459 ), .ZN(_u10_u20_n2448 ) );
NOR2_X1 _u10_u20_U336  ( .A1(_u10_u20_n2455 ), .A2(_u10_u20_n2456 ), .ZN(_u10_u20_n2449 ) );
NAND2_X1 _u10_u20_U335  ( .A1(_u10_u20_n2454 ), .A2(_u10_u20_n2438 ), .ZN(_u10_u20_n2452 ) );
NOR4_X1 _u10_u20_U334  ( .A1(_u10_u20_n2452 ), .A2(_u10_u20_n2453 ), .A3(_u10_u20_n2443 ), .A4(_u10_u20_n2143 ), .ZN(_u10_u20_n2451 ) );
NOR2_X1 _u10_u20_U333  ( .A1(_u10_u20_n2451 ), .A2(_u10_u20_n2356 ), .ZN(_u10_u20_n2450 ) );
NOR4_X1 _u10_u20_U332  ( .A1(_u10_u20_n2447 ), .A2(_u10_u20_n2448 ), .A3(_u10_u20_n2449 ), .A4(_u10_u20_n2450 ), .ZN(_u10_u20_n2390 ) );
NAND2_X1 _u10_u20_U331  ( .A1(_u10_u20_n2445 ), .A2(_u10_u20_n2446 ), .ZN(_u10_u20_n2155 ) );
INV_X1 _u10_u20_U330  ( .A(_u10_u20_n2155 ), .ZN(_u10_u20_n1892 ) );
INV_X1 _u10_u20_U329  ( .A(_u10_u20_n2444 ), .ZN(_u10_u20_n2088 ) );
NAND2_X1 _u10_u20_U328  ( .A1(_u10_u20_n1892 ), .A2(_u10_u20_n2088 ), .ZN(_u10_u20_n2337 ) );
NOR3_X1 _u10_u20_U327  ( .A1(_u10_u20_n2441 ), .A2(_u10_u20_n2442 ), .A3(_u10_u20_n2443 ), .ZN(_u10_u20_n2440 ) );
NAND4_X1 _u10_u20_U326  ( .A1(_u10_u20_n2193 ), .A2(_u10_u20_n2355 ), .A3(_u10_u20_n2439 ), .A4(_u10_u20_n2440 ), .ZN(_u10_u20_n2434 ) );
NAND3_X1 _u10_u20_U325  ( .A1(_u10_u20_n2437 ), .A2(_u10_u20_n2438 ), .A3(_u10_u20_n2059 ), .ZN(_u10_u20_n2435 ) );
NOR4_X1 _u10_u20_U324  ( .A1(_u10_u20_n2434 ), .A2(_u10_u20_n2435 ), .A3(_u10_u20_n1837 ), .A4(_u10_u20_n2436 ), .ZN(_u10_u20_n2433 ) );
NOR2_X1 _u10_u20_U323  ( .A1(_u10_u20_n2433 ), .A2(_u10_u20_n1836 ), .ZN(_u10_u20_n2415 ) );
INV_X1 _u10_u20_U322  ( .A(_u10_u20_n2432 ), .ZN(_u10_u20_n2178 ) );
NOR2_X1 _u10_u20_U321  ( .A1(_u10_u20_n1960 ), .A2(_u10_u20_n2431 ), .ZN(_u10_u20_n2430 ) );
NOR4_X1 _u10_u20_U320  ( .A1(_u10_u20_n2178 ), .A2(_u10_u20_n2429 ), .A3(_u10_u20_n2430 ), .A4(_u10_u20_n2179 ), .ZN(_u10_u20_n2416 ) );
NOR2_X1 _u10_u20_U319  ( .A1(_u10_u20_n2427 ), .A2(_u10_u20_n2428 ), .ZN(_u10_u20_n2426 ) );
NAND4_X1 _u10_u20_U318  ( .A1(_u10_u20_n2286 ), .A2(_u10_u20_n1969 ), .A3(_u10_u20_n2282 ), .A4(_u10_u20_n2426 ), .ZN(_u10_u20_n2425 ) );
NAND2_X1 _u10_u20_U317  ( .A1(_u10_u20_n2031 ), .A2(_u10_u20_n2425 ), .ZN(_u10_u20_n2422 ) );
NAND3_X1 _u10_u20_U316  ( .A1(_u10_u20_n2422 ), .A2(_u10_u20_n2423 ), .A3(_u10_u20_n2424 ), .ZN(_u10_u20_n2419 ) );
NOR4_X1 _u10_u20_U315  ( .A1(_u10_u20_n2419 ), .A2(_u10_u20_n1978 ), .A3(_u10_u20_n2420 ), .A4(_u10_u20_n2421 ), .ZN(_u10_u20_n2418 ) );
NOR2_X1 _u10_u20_U314  ( .A1(_u10_u20_n2418 ), .A2(_u10_u20_n2359 ), .ZN(_u10_u20_n2417 ) );
NOR3_X1 _u10_u20_U313  ( .A1(_u10_u20_n2415 ), .A2(_u10_u20_n2416 ), .A3(_u10_u20_n2417 ), .ZN(_u10_u20_n2414 ) );
NAND4_X1 _u10_u20_U312  ( .A1(_u10_u20_n2337 ), .A2(_u10_u20_n2412 ), .A3(_u10_u20_n2413 ), .A4(_u10_u20_n2414 ), .ZN(_u10_u20_n2392 ) );
NAND2_X1 _u10_u20_U311  ( .A1(_u10_u20_n2411 ), .A2(_u10_u20_n1936 ), .ZN(_u10_u20_n2410 ) );
NAND2_X1 _u10_u20_U310  ( .A1(_u10_u20_n2409 ), .A2(_u10_u20_n2410 ), .ZN(_u10_u20_n2408 ) );
NAND3_X1 _u10_u20_U309  ( .A1(_u10_u20_n2408 ), .A2(_u10_u20_n2305 ), .A3(_u10_u20_n1894 ), .ZN(_u10_u20_n2402 ) );
NAND3_X1 _u10_u20_U308  ( .A1(_u10_u20_n2329 ), .A2(_u10_u20_n2407 ), .A3(_u10_u20_n2255 ), .ZN(_u10_u20_n2403 ) );
NAND3_X1 _u10_u20_U307  ( .A1(_u10_u20_n1924 ), .A2(_u10_u20_n2405 ), .A3(_u10_u20_n2406 ), .ZN(_u10_u20_n2404 ) );
NAND3_X1 _u10_u20_U306  ( .A1(_u10_u20_n2402 ), .A2(_u10_u20_n2403 ), .A3(_u10_u20_n2404 ), .ZN(_u10_u20_n2393 ) );
INV_X1 _u10_u20_U305  ( .A(_u10_u20_n1932 ), .ZN(_u10_u20_n2399 ) );
NOR2_X1 _u10_u20_U304  ( .A1(_u10_u20_n2401 ), .A2(_u10_u20_n2161 ), .ZN(_u10_u20_n2400 ) );
NOR2_X1 _u10_u20_U303  ( .A1(_u10_u20_n2399 ), .A2(_u10_u20_n2400 ), .ZN(_u10_u20_n2394 ) );
NOR2_X1 _u10_u20_U302  ( .A1(_u10_u20_n2110 ), .A2(_u10_u20_n2398 ), .ZN(_u10_u20_n2397 ) );
NOR2_X1 _u10_u20_U301  ( .A1(_u10_u20_n2396 ), .A2(_u10_u20_n2397 ), .ZN(_u10_u20_n2395 ) );
NOR4_X1 _u10_u20_U300  ( .A1(_u10_u20_n2392 ), .A2(_u10_u20_n2393 ), .A3(_u10_u20_n2394 ), .A4(_u10_u20_n2395 ), .ZN(_u10_u20_n2391 ) );
NAND4_X1 _u10_u20_U299  ( .A1(_u10_u20_n2388 ), .A2(_u10_u20_n2389 ), .A3(_u10_u20_n2390 ), .A4(_u10_u20_n2391 ), .ZN(_u10_u20_n2387 ) );
MUX2_X1 _u10_u20_U298  ( .A(_u10_u20_n2387 ), .B(_u10_SYNOPSYS_UNCONNECTED_5 ), .S(_u10_u20_n1819 ), .Z(_u10_u20_n1810 ) );
NAND2_X1 _u10_u20_U297  ( .A1(_u10_u20_n2386 ), .A2(_u10_u20_n2007 ), .ZN(_u10_u20_n2369 ) );
AND2_X1 _u10_u20_U296  ( .A1(1'b0), .A2(_u10_u20_n2195 ), .ZN(_u10_u20_n2308 ) );
NAND2_X1 _u10_u20_U295  ( .A1(_u10_u20_n2308 ), .A2(_u10_u20_n2036 ), .ZN(_u10_u20_n2384 ) );
AND2_X1 _u10_u20_U294  ( .A1(_u10_u20_n2384 ), .A2(_u10_u20_n2385 ), .ZN(_u10_u20_n2275 ) );
AND4_X1 _u10_u20_U293  ( .A1(_u10_u20_n2275 ), .A2(_u10_u20_n2286 ), .A3(_u10_u20_n2383 ), .A4(_u10_u20_n2285 ), .ZN(_u10_u20_n2225 ) );
NAND3_X1 _u10_u20_U292  ( .A1(_u10_u20_n2195 ), .A2(_u10_u20_n2223 ), .A3(1'b0), .ZN(_u10_u20_n2021 ) );
INV_X1 _u10_u20_U291  ( .A(_u10_u20_n2021 ), .ZN(_u10_u20_n2167 ) );
NAND2_X1 _u10_u20_U290  ( .A1(_u10_u20_n2036 ), .A2(_u10_u20_n2167 ), .ZN(_u10_u20_n1970 ) );
AND3_X1 _u10_u20_U289  ( .A1(_u10_u20_n1970 ), .A2(_u10_u20_n2164 ), .A3(_u10_u20_n2382 ), .ZN(_u10_u20_n2381 ) );
NAND4_X1 _u10_u20_U288  ( .A1(_u10_u20_n2225 ), .A2(_u10_u20_n2379 ), .A3(_u10_u20_n2380 ), .A4(_u10_u20_n2381 ), .ZN(_u10_u20_n2378 ) );
NAND2_X1 _u10_u20_U287  ( .A1(_u10_u20_n1967 ), .A2(_u10_u20_n2378 ), .ZN(_u10_u20_n2370 ) );
NAND2_X1 _u10_u20_U286  ( .A1(_u10_u20_n2081 ), .A2(_u10_u20_n2377 ), .ZN(_u10_u20_n2371 ) );
NOR2_X1 _u10_u20_U285  ( .A1(_u10_u20_n2375 ), .A2(_u10_u20_n2376 ), .ZN(_u10_u20_n2373 ) );
NOR2_X1 _u10_u20_U284  ( .A1(_u10_u20_n2373 ), .A2(_u10_u20_n2374 ), .ZN(_u10_u20_n2372 ) );
NAND4_X1 _u10_u20_U283  ( .A1(_u10_u20_n2369 ), .A2(_u10_u20_n2370 ), .A3(_u10_u20_n2371 ), .A4(_u10_u20_n2372 ), .ZN(_u10_u20_n2309 ) );
NOR2_X1 _u10_u20_U282  ( .A1(_u10_u20_n2000 ), .A2(_u10_u20_n2368 ), .ZN(_u10_u20_n2360 ) );
NOR2_X1 _u10_u20_U281  ( .A1(_u10_u20_n2366 ), .A2(_u10_u20_n2367 ), .ZN(_u10_u20_n2361 ) );
NOR2_X1 _u10_u20_U280  ( .A1(_u10_u20_n1868 ), .A2(_u10_u20_n2365 ), .ZN(_u10_u20_n2362 ) );
NOR2_X1 _u10_u20_U279  ( .A1(_u10_u20_n2364 ), .A2(_u10_u20_n1859 ), .ZN(_u10_u20_n2363 ) );
NOR4_X1 _u10_u20_U278  ( .A1(_u10_u20_n2360 ), .A2(_u10_u20_n2361 ), .A3(_u10_u20_n2362 ), .A4(_u10_u20_n2363 ), .ZN(_u10_u20_n2316 ) );
NOR2_X1 _u10_u20_U277  ( .A1(_u10_u20_n2359 ), .A2(_u10_u20_n1970 ), .ZN(_u10_u20_n2351 ) );
NOR2_X1 _u10_u20_U276  ( .A1(_u10_u20_n2358 ), .A2(_u10_u20_n1840 ), .ZN(_u10_u20_n2352 ) );
NOR2_X1 _u10_u20_U275  ( .A1(_u10_u20_n2356 ), .A2(_u10_u20_n2357 ), .ZN(_u10_u20_n2353 ) );
NOR2_X1 _u10_u20_U274  ( .A1(_u10_u20_n1836 ), .A2(_u10_u20_n2355 ), .ZN(_u10_u20_n2354 ) );
NOR4_X1 _u10_u20_U273  ( .A1(_u10_u20_n2351 ), .A2(_u10_u20_n2352 ), .A3(_u10_u20_n2353 ), .A4(_u10_u20_n2354 ), .ZN(_u10_u20_n2317 ) );
NOR2_X1 _u10_u20_U272  ( .A1(_u10_u20_n1873 ), .A2(_u10_u20_n2101 ), .ZN(_u10_u20_n2349 ) );
NOR2_X1 _u10_u20_U271  ( .A1(_u10_u20_n2349 ), .A2(_u10_u20_n2350 ), .ZN(_u10_u20_n2338 ) );
NOR2_X1 _u10_u20_U270  ( .A1(_u10_u20_n2347 ), .A2(_u10_u20_n2348 ), .ZN(_u10_u20_n2345 ) );
NOR2_X1 _u10_u20_U269  ( .A1(_u10_u20_n2345 ), .A2(_u10_u20_n2346 ), .ZN(_u10_u20_n2339 ) );
NOR2_X1 _u10_u20_U268  ( .A1(_u10_u20_n2344 ), .A2(_u10_u20_n2142 ), .ZN(_u10_u20_n2340 ) );
NOR2_X1 _u10_u20_U267  ( .A1(_u10_u20_n2342 ), .A2(_u10_u20_n2343 ), .ZN(_u10_u20_n2341 ) );
NOR4_X1 _u10_u20_U266  ( .A1(_u10_u20_n2338 ), .A2(_u10_u20_n2339 ), .A3(_u10_u20_n2340 ), .A4(_u10_u20_n2341 ), .ZN(_u10_u20_n2318 ) );
INV_X1 _u10_u20_U265  ( .A(_u10_u20_n2337 ), .ZN(_u10_u20_n2320 ) );
NOR2_X1 _u10_u20_U264  ( .A1(_u10_u20_n1970 ), .A2(1'b0), .ZN(_u10_u20_n2027 ) );
INV_X1 _u10_u20_U263  ( .A(_u10_u20_n2027 ), .ZN(_u10_u20_n2331 ) );
NOR2_X1 _u10_u20_U262  ( .A1(_u10_u20_n2174 ), .A2(_u10_u20_n2216 ), .ZN(_u10_u20_n2333 ) );
AND2_X1 _u10_u20_U261  ( .A1(_u10_u20_n1928 ), .A2(_u10_u20_n2336 ), .ZN(_u10_u20_n2334 ) );
NOR4_X1 _u10_u20_U260  ( .A1(_u10_u20_n1937 ), .A2(_u10_u20_n2333 ), .A3(_u10_u20_n2334 ), .A4(_u10_u20_n2335 ), .ZN(_u10_u20_n2332 ) );
NOR3_X1 _u10_u20_U259  ( .A1(_u10_u20_n2331 ), .A2(_u10_u20_n2332 ), .A3(_u10_u20_n1915 ), .ZN(_u10_u20_n2321 ) );
NOR3_X1 _u10_u20_U258  ( .A1(_u10_u20_n2291 ), .A2(_u10_u20_n2330 ), .A3(_u10_u20_n2021 ), .ZN(_u10_u20_n2322 ) );
NOR2_X1 _u10_u20_U257  ( .A1(_u10_u20_n2329 ), .A2(_u10_u20_n2169 ), .ZN(_u10_u20_n2324 ) );
NOR2_X1 _u10_u20_U256  ( .A1(1'b0), .A2(_u10_u20_n2328 ), .ZN(_u10_u20_n2327 ) );
NOR2_X1 _u10_u20_U255  ( .A1(_u10_u20_n2326 ), .A2(_u10_u20_n2327 ), .ZN(_u10_u20_n2325 ) );
NOR3_X1 _u10_u20_U254  ( .A1(_u10_u20_n2324 ), .A2(1'b0), .A3(_u10_u20_n2325 ), .ZN(_u10_u20_n2323 ) );
NOR4_X1 _u10_u20_U253  ( .A1(_u10_u20_n2320 ), .A2(_u10_u20_n2321 ), .A3(_u10_u20_n2322 ), .A4(_u10_u20_n2323 ), .ZN(_u10_u20_n2319 ) );
AND4_X1 _u10_u20_U252  ( .A1(_u10_u20_n2316 ), .A2(_u10_u20_n2317 ), .A3(_u10_u20_n2318 ), .A4(_u10_u20_n2319 ), .ZN(_u10_u20_n1991 ) );
INV_X1 _u10_u20_U251  ( .A(_u10_u20_n2315 ), .ZN(_u10_u20_n2313 ) );
NAND3_X1 _u10_u20_U250  ( .A1(_u10_u20_n1991 ), .A2(_u10_u20_n2313 ), .A3(_u10_u20_n2314 ), .ZN(_u10_u20_n2310 ) );
NOR4_X1 _u10_u20_U249  ( .A1(_u10_u20_n2309 ), .A2(_u10_u20_n2310 ), .A3(_u10_u20_n2311 ), .A4(_u10_u20_n2312 ), .ZN(_u10_u20_n2117 ) );
NAND3_X1 _u10_u20_U248  ( .A1(_u10_u20_n2108 ), .A2(_u10_u20_n2107 ), .A3(_u10_u20_n2308 ), .ZN(_u10_u20_n2217 ) );
NOR3_X1 _u10_u20_U247  ( .A1(_u10_u20_n2306 ), .A2(_u10_u20_n2307 ), .A3(_u10_u20_n2027 ), .ZN(_u10_u20_n2277 ) );
NAND3_X1 _u10_u20_U246  ( .A1(_u10_u20_n2217 ), .A2(_u10_u20_n2305 ), .A3(_u10_u20_n2277 ), .ZN(_u10_u20_n2157 ) );
NAND2_X1 _u10_u20_U245  ( .A1(_u10_u20_n2089 ), .A2(_u10_u20_n2157 ), .ZN(_u10_u20_n2296 ) );
INV_X1 _u10_u20_U244  ( .A(_u10_u20_n2304 ), .ZN(_u10_u20_n2297 ) );
NOR2_X1 _u10_u20_U243  ( .A1(_u10_u20_n2302 ), .A2(_u10_u20_n2303 ), .ZN(_u10_u20_n2299 ) );
NOR3_X1 _u10_u20_U242  ( .A1(_u10_u20_n2299 ), .A2(_u10_u20_n2300 ), .A3(_u10_u20_n2301 ), .ZN(_u10_u20_n2298 ) );
NAND4_X1 _u10_u20_U241  ( .A1(_u10_u20_n2295 ), .A2(_u10_u20_n2296 ), .A3(_u10_u20_n2297 ), .A4(_u10_u20_n2298 ), .ZN(_u10_u20_n2294 ) );
NAND2_X1 _u10_u20_U240  ( .A1(_u10_u20_n2293 ), .A2(_u10_u20_n2294 ), .ZN(_u10_u20_n2257 ) );
NAND2_X1 _u10_u20_U239  ( .A1(_u10_u20_n2165 ), .A2(_u10_u20_n2166 ), .ZN(_u10_u20_n2288 ) );
NAND2_X1 _u10_u20_U238  ( .A1(_u10_u20_n2078 ), .A2(_u10_u20_n2279 ), .ZN(_u10_u20_n2292 ) );
NAND2_X1 _u10_u20_U237  ( .A1(_u10_u20_n2291 ), .A2(_u10_u20_n2292 ), .ZN(_u10_u20_n2290 ) );
NAND2_X1 _u10_u20_U236  ( .A1(_u10_u20_n2059 ), .A2(_u10_u20_n2290 ), .ZN(_u10_u20_n2289 ) );
NAND2_X1 _u10_u20_U235  ( .A1(_u10_u20_n2288 ), .A2(_u10_u20_n2289 ), .ZN(_u10_u20_n2201 ) );
NAND2_X1 _u10_u20_U234  ( .A1(1'b0), .A2(_u10_u20_n2201 ), .ZN(_u10_u20_n2258 ) );
INV_X1 _u10_u20_U233  ( .A(_u10_u20_n2287 ), .ZN(_u10_u20_n2283 ) );
AND4_X1 _u10_u20_U232  ( .A1(_u10_u20_n2285 ), .A2(_u10_u20_n2226 ), .A3(_u10_u20_n1970 ), .A4(_u10_u20_n2286 ), .ZN(_u10_u20_n2284 ) );
NAND4_X1 _u10_u20_U231  ( .A1(_u10_u20_n2281 ), .A2(_u10_u20_n2282 ), .A3(_u10_u20_n2283 ), .A4(_u10_u20_n2284 ), .ZN(_u10_u20_n2280 ) );
NAND2_X1 _u10_u20_U230  ( .A1(_u10_u20_n2279 ), .A2(_u10_u20_n2280 ), .ZN(_u10_u20_n2259 ) );
NAND4_X1 _u10_u20_U229  ( .A1(_u10_u20_n2275 ), .A2(_u10_u20_n2276 ), .A3(_u10_u20_n2277 ), .A4(_u10_u20_n2278 ), .ZN(_u10_u20_n2271 ) );
NAND2_X1 _u10_u20_U228  ( .A1(_u10_u20_n1933 ), .A2(_u10_u20_n2164 ), .ZN(_u10_u20_n2272 ) );
NOR2_X1 _u10_u20_U227  ( .A1(_u10_u20_n2274 ), .A2(_u10_u20_n2130 ), .ZN(_u10_u20_n2273 ) );
NOR4_X1 _u10_u20_U226  ( .A1(_u10_u20_n2271 ), .A2(_u10_u20_n2272 ), .A3(_u10_u20_n1978 ), .A4(_u10_u20_n2273 ), .ZN(_u10_u20_n2270 ) );
NOR2_X1 _u10_u20_U225  ( .A1(_u10_u20_n2270 ), .A2(_u10_u20_n2025 ), .ZN(_u10_u20_n2261 ) );
NAND3_X1 _u10_u20_U224  ( .A1(_u10_u20_n1933 ), .A2(_u10_u20_n1936 ), .A3(_u10_u20_n2269 ), .ZN(_u10_u20_n2268 ) );
NOR3_X1 _u10_u20_U223  ( .A1(_u10_u20_n2268 ), .A2(_u10_u20_n1844 ), .A3(_u10_u20_n2157 ), .ZN(_u10_u20_n2267 ) );
NOR2_X1 _u10_u20_U222  ( .A1(1'b0), .A2(_u10_u20_n2267 ), .ZN(_u10_u20_n2265 ) );
NOR3_X1 _u10_u20_U221  ( .A1(_u10_u20_n2264 ), .A2(_u10_u20_n2265 ), .A3(_u10_u20_n2266 ), .ZN(_u10_u20_n2263 ) );
NOR2_X1 _u10_u20_U220  ( .A1(_u10_u20_n2263 ), .A2(_u10_u20_n1843 ), .ZN(_u10_u20_n2262 ) );
NOR2_X1 _u10_u20_U219  ( .A1(_u10_u20_n2261 ), .A2(_u10_u20_n2262 ), .ZN(_u10_u20_n2260 ) );
NAND4_X1 _u10_u20_U218  ( .A1(_u10_u20_n2257 ), .A2(_u10_u20_n2258 ), .A3(_u10_u20_n2259 ), .A4(_u10_u20_n2260 ), .ZN(_u10_u20_n2230 ) );
INV_X1 _u10_u20_U217  ( .A(_u10_u20_n2217 ), .ZN(_u10_u20_n2242 ) );
NAND2_X1 _u10_u20_U216  ( .A1(_u10_u20_n2168 ), .A2(_u10_u20_n2169 ), .ZN(_u10_u20_n2244 ) );
NAND2_X1 _u10_u20_U215  ( .A1(_u10_u20_n2255 ), .A2(_u10_u20_n2256 ), .ZN(_u10_u20_n2245 ) );
NAND2_X1 _u10_u20_U214  ( .A1(_u10_u20_n2253 ), .A2(_u10_u20_n2254 ), .ZN(_u10_u20_n2252 ) );
NAND2_X1 _u10_u20_U213  ( .A1(_u10_u20_n2251 ), .A2(_u10_u20_n2252 ), .ZN(_u10_u20_n2246 ) );
NAND2_X1 _u10_u20_U212  ( .A1(_u10_u20_n2152 ), .A2(_u10_u20_n1928 ), .ZN(_u10_u20_n2250 ) );
NAND2_X1 _u10_u20_U211  ( .A1(_u10_u20_n2249 ), .A2(_u10_u20_n2250 ), .ZN(_u10_u20_n2248 ) );
NAND2_X1 _u10_u20_U210  ( .A1(_u10_u20_n2105 ), .A2(_u10_u20_n2248 ), .ZN(_u10_u20_n2247 ) );
NAND4_X1 _u10_u20_U209  ( .A1(_u10_u20_n2244 ), .A2(_u10_u20_n2245 ), .A3(_u10_u20_n2246 ), .A4(_u10_u20_n2247 ), .ZN(_u10_u20_n2243 ) );
NAND2_X1 _u10_u20_U208  ( .A1(_u10_u20_n2242 ), .A2(_u10_u20_n2243 ), .ZN(_u10_u20_n2237 ) );
NAND2_X1 _u10_u20_U207  ( .A1(1'b0), .A2(_u10_u20_n2241 ), .ZN(_u10_u20_n2238 ) );
NAND2_X1 _u10_u20_U206  ( .A1(_u10_u20_n2214 ), .A2(_u10_u20_n2240 ), .ZN(_u10_u20_n2239 ) );
NAND3_X1 _u10_u20_U205  ( .A1(_u10_u20_n2237 ), .A2(_u10_u20_n2238 ), .A3(_u10_u20_n2239 ), .ZN(_u10_u20_n2231 ) );
AND2_X1 _u10_u20_U204  ( .A1(_u10_u20_n2200 ), .A2(_u10_u20_n2236 ), .ZN(_u10_u20_n2232 ) );
NOR2_X1 _u10_u20_U203  ( .A1(_u10_u20_n2234 ), .A2(_u10_u20_n2235 ), .ZN(_u10_u20_n2233 ) );
NOR4_X1 _u10_u20_U202  ( .A1(_u10_u20_n2230 ), .A2(_u10_u20_n2231 ), .A3(_u10_u20_n2232 ), .A4(_u10_u20_n2233 ), .ZN(_u10_u20_n2118 ) );
NAND2_X1 _u10_u20_U201  ( .A1(_u10_u20_n2214 ), .A2(_u10_u20_n2049 ), .ZN(_u10_u20_n2229 ) );
NAND2_X1 _u10_u20_U200  ( .A1(_u10_u20_n2228 ), .A2(_u10_u20_n2229 ), .ZN(_u10_u20_n2227 ) );
NAND2_X1 _u10_u20_U199  ( .A1(_u10_u20_n2043 ), .A2(_u10_u20_n2227 ), .ZN(_u10_u20_n2204 ) );
NAND2_X1 _u10_u20_U198  ( .A1(_u10_u20_n2225 ), .A2(_u10_u20_n2226 ), .ZN(_u10_u20_n2224 ) );
NAND2_X1 _u10_u20_U197  ( .A1(_u10_u20_n1899 ), .A2(_u10_u20_n2224 ), .ZN(_u10_u20_n2205 ) );
NAND2_X1 _u10_u20_U196  ( .A1(_u10_u20_n2222 ), .A2(_u10_u20_n2223 ), .ZN(_u10_u20_n1870 ) );
NAND4_X1 _u10_u20_U195  ( .A1(_u10_u20_n2220 ), .A2(_u10_u20_n2131 ), .A3(_u10_u20_n2221 ), .A4(_u10_u20_n1870 ), .ZN(_u10_u20_n2219 ) );
NAND2_X1 _u10_u20_U194  ( .A1(_u10_u20_n2218 ), .A2(_u10_u20_n2219 ), .ZN(_u10_u20_n2206 ) );
NOR2_X1 _u10_u20_U193  ( .A1(_u10_u20_n1925 ), .A2(_u10_u20_n2217 ), .ZN(_u10_u20_n2215 ) );
NOR4_X1 _u10_u20_U192  ( .A1(_u10_u20_n2213 ), .A2(_u10_u20_n2214 ), .A3(_u10_u20_n2215 ), .A4(_u10_u20_n2216 ), .ZN(_u10_u20_n2211 ) );
NOR2_X1 _u10_u20_U191  ( .A1(_u10_u20_n2211 ), .A2(_u10_u20_n2212 ), .ZN(_u10_u20_n2208 ) );
NOR2_X1 _u10_u20_U190  ( .A1(_u10_u20_n1888 ), .A2(_u10_u20_n2210 ), .ZN(_u10_u20_n2209 ) );
NOR2_X1 _u10_u20_U189  ( .A1(_u10_u20_n2208 ), .A2(_u10_u20_n2209 ), .ZN(_u10_u20_n2207 ) );
NAND4_X1 _u10_u20_U188  ( .A1(_u10_u20_n2204 ), .A2(_u10_u20_n2205 ), .A3(_u10_u20_n2206 ), .A4(_u10_u20_n2207 ), .ZN(_u10_u20_n2170 ) );
OR2_X1 _u10_u20_U187  ( .A1(_u10_u20_n2202 ), .A2(_u10_u20_n2203 ), .ZN(_u10_u20_n2197 ) );
NAND2_X1 _u10_u20_U186  ( .A1(1'b0), .A2(_u10_u20_n2201 ), .ZN(_u10_u20_n2198 ) );
NAND2_X1 _u10_u20_U185  ( .A1(_u10_u20_n2063 ), .A2(_u10_u20_n2200 ), .ZN(_u10_u20_n2199 ) );
NAND3_X1 _u10_u20_U184  ( .A1(_u10_u20_n2197 ), .A2(_u10_u20_n2198 ), .A3(_u10_u20_n2199 ), .ZN(_u10_u20_n2196 ) );
NAND2_X1 _u10_u20_U183  ( .A1(_u10_u20_n2195 ), .A2(_u10_u20_n2196 ), .ZN(_u10_u20_n2180 ) );
NAND2_X1 _u10_u20_U182  ( .A1(_u10_u20_n2195 ), .A2(_u10_u20_n1918 ), .ZN(_u10_u20_n2192 ) );
NAND4_X1 _u10_u20_U181  ( .A1(_u10_u20_n2192 ), .A2(_u10_u20_n2021 ), .A3(_u10_u20_n2193 ), .A4(_u10_u20_n2194 ), .ZN(_u10_u20_n2188 ) );
NAND2_X1 _u10_u20_U180  ( .A1(_u10_u20_n2188 ), .A2(_u10_u20_n2191 ), .ZN(_u10_u20_n2181 ) );
NAND2_X1 _u10_u20_U179  ( .A1(1'b0), .A2(_u10_u20_n2190 ), .ZN(_u10_u20_n2185 ) );
NAND2_X1 _u10_u20_U178  ( .A1(_u10_u20_n2189 ), .A2(_u10_SYNOPSYS_UNCONNECTED_6 ), .ZN(_u10_u20_n2186 ) );
INV_X1 _u10_u20_U177  ( .A(_u10_u20_n2188 ), .ZN(_u10_u20_n2187 ) );
NAND3_X1 _u10_u20_U176  ( .A1(_u10_u20_n2185 ), .A2(_u10_u20_n2186 ), .A3(_u10_u20_n2187 ), .ZN(_u10_u20_n2184 ) );
NAND2_X1 _u10_u20_U175  ( .A1(_u10_u20_n2183 ), .A2(_u10_u20_n2184 ), .ZN(_u10_u20_n2182 ) );
NAND3_X1 _u10_u20_U174  ( .A1(_u10_u20_n2180 ), .A2(_u10_u20_n2181 ), .A3(_u10_u20_n2182 ), .ZN(_u10_u20_n2171 ) );
INV_X1 _u10_u20_U173  ( .A(_u10_u20_n2179 ), .ZN(_u10_u20_n1963 ) );
NOR2_X1 _u10_u20_U172  ( .A1(_u10_u20_n1963 ), .A2(_u10_u20_n2178 ), .ZN(_u10_u20_n2172 ) );
INV_X1 _u10_u20_U171  ( .A(_u10_u20_n2177 ), .ZN(_u10_u20_n2176 ) );
NOR3_X1 _u10_u20_U170  ( .A1(_u10_u20_n2174 ), .A2(_u10_u20_n2175 ), .A3(_u10_u20_n2176 ), .ZN(_u10_u20_n2173 ) );
NOR4_X1 _u10_u20_U169  ( .A1(_u10_u20_n2170 ), .A2(_u10_u20_n2171 ), .A3(_u10_u20_n2172 ), .A4(_u10_u20_n2173 ), .ZN(_u10_u20_n2119 ) );
NAND3_X1 _u10_u20_U168  ( .A1(_u10_u20_n2168 ), .A2(_u10_u20_n2169 ), .A3(1'b0), .ZN(_u10_u20_n2148 ) );
NAND3_X1 _u10_u20_U167  ( .A1(_u10_u20_n2165 ), .A2(_u10_u20_n2166 ), .A3(_u10_u20_n2167 ), .ZN(_u10_u20_n2149 ) );
NAND4_X1 _u10_u20_U166  ( .A1(_u10_u20_n2162 ), .A2(_u10_u20_n1933 ), .A3(_u10_u20_n2163 ), .A4(_u10_u20_n2164 ), .ZN(_u10_u20_n2160 ) );
NOR4_X1 _u10_u20_U165  ( .A1(_u10_u20_n2160 ), .A2(_u10_u20_n2157 ), .A3(_u10_u20_n1844 ), .A4(_u10_u20_n2161 ), .ZN(_u10_u20_n2158 ) );
NOR2_X1 _u10_u20_U164  ( .A1(_u10_u20_n2158 ), .A2(_u10_u20_n2159 ), .ZN(_u10_u20_n2153 ) );
INV_X1 _u10_u20_U163  ( .A(_u10_u20_n2157 ), .ZN(_u10_u20_n2129 ) );
NOR3_X1 _u10_u20_U162  ( .A1(_u10_u20_n2155 ), .A2(_u10_u20_n2129 ), .A3(_u10_u20_n2156 ), .ZN(_u10_u20_n2154 ) );
NOR2_X1 _u10_u20_U161  ( .A1(_u10_u20_n2153 ), .A2(_u10_u20_n2154 ), .ZN(_u10_u20_n2150 ) );
NAND3_X1 _u10_u20_U160  ( .A1(1'b0), .A2(_u10_u20_n1928 ), .A3(_u10_u20_n2152 ), .ZN(_u10_u20_n2151 ) );
NAND4_X1 _u10_u20_U159  ( .A1(_u10_u20_n2148 ), .A2(_u10_u20_n2149 ), .A3(_u10_u20_n2150 ), .A4(_u10_u20_n2151 ), .ZN(_u10_u20_n2121 ) );
NAND2_X1 _u10_u20_U158  ( .A1(_u10_u20_n2107 ), .A2(_u10_u20_n2147 ), .ZN(_u10_u20_n2146 ) );
NAND2_X1 _u10_u20_U157  ( .A1(_u10_u20_n2145 ), .A2(_u10_u20_n2146 ), .ZN(_u10_u20_n2144 ) );
NAND2_X1 _u10_u20_U156  ( .A1(_u10_u20_n2143 ), .A2(_u10_u20_n2144 ), .ZN(_u10_u20_n2134 ) );
NAND2_X1 _u10_u20_U155  ( .A1(_u10_u20_n2141 ), .A2(_u10_u20_n2142 ), .ZN(_u10_u20_n2140 ) );
NAND2_X1 _u10_u20_U154  ( .A1(_u10_u20_n2139 ), .A2(_u10_u20_n2140 ), .ZN(_u10_u20_n2135 ) );
OR2_X1 _u10_u20_U153  ( .A1(_u10_u20_n2110 ), .A2(_u10_u20_n1911 ), .ZN(_u10_u20_n2137 ) );
NAND2_X1 _u10_u20_U152  ( .A1(_u10_u20_n2137 ), .A2(_u10_u20_n2138 ), .ZN(_u10_u20_n2136 ) );
NAND3_X1 _u10_u20_U151  ( .A1(_u10_u20_n2134 ), .A2(_u10_u20_n2135 ), .A3(_u10_u20_n2136 ), .ZN(_u10_u20_n2122 ) );
NOR2_X1 _u10_u20_U150  ( .A1(_u10_u20_n2133 ), .A2(_u10_u20_n1891 ), .ZN(_u10_u20_n2132 ) );
NOR2_X1 _u10_u20_U149  ( .A1(_u10_u20_n2131 ), .A2(_u10_u20_n2132 ), .ZN(_u10_u20_n2123 ) );
NOR2_X1 _u10_u20_U148  ( .A1(_u10_u20_n2129 ), .A2(_u10_u20_n2130 ), .ZN(_u10_u20_n2127 ) );
NOR2_X1 _u10_u20_U147  ( .A1(_u10_u20_n2127 ), .A2(_u10_u20_n2128 ), .ZN(_u10_u20_n2125 ) );
NOR2_X1 _u10_u20_U146  ( .A1(_u10_u20_n2125 ), .A2(_u10_u20_n2126 ), .ZN(_u10_u20_n2124 ) );
NOR4_X1 _u10_u20_U145  ( .A1(_u10_u20_n2121 ), .A2(_u10_u20_n2122 ), .A3(_u10_u20_n2123 ), .A4(_u10_u20_n2124 ), .ZN(_u10_u20_n2120 ) );
NAND4_X1 _u10_u20_U144  ( .A1(_u10_u20_n2117 ), .A2(_u10_u20_n2118 ), .A3(_u10_u20_n2119 ), .A4(_u10_u20_n2120 ), .ZN(_u10_u20_n2116 ) );
MUX2_X1 _u10_u20_U143  ( .A(_u10_u20_n2116 ), .B(_u10_SYNOPSYS_UNCONNECTED_6 ), .S(_u10_u20_n1819 ), .Z(_u10_u20_n1811 ) );
INV_X1 _u10_u20_U142  ( .A(_u10_u20_n2115 ), .ZN(_u10_u20_n2006 ) );
NOR3_X1 _u10_u20_U141  ( .A1(_u10_u20_n2006 ), .A2(_u10_u20_n2114 ), .A3(_u10_u20_n2081 ), .ZN(_u10_u20_n1854 ) );
NAND2_X1 _u10_u20_U140  ( .A1(_u10_u20_n2112 ), .A2(_u10_u20_n2113 ), .ZN(_u10_u20_n1872 ) );
INV_X1 _u10_u20_U139  ( .A(_u10_u20_n1872 ), .ZN(_u10_u20_n1882 ) );
NAND4_X1 _u10_u20_U138  ( .A1(_u10_u20_n1854 ), .A2(_u10_u20_n1882 ), .A3(_u10_u20_n2111 ), .A4(_u10_u20_n1868 ), .ZN(_u10_u20_n2109 ) );
NAND2_X1 _u10_u20_U137  ( .A1(_u10_u20_n2109 ), .A2(_u10_u20_n2110 ), .ZN(_u10_u20_n2098 ) );
NAND2_X1 _u10_u20_U136  ( .A1(1'b0), .A2(_u10_u20_n1983 ), .ZN(_u10_u20_n2023 ) );
INV_X1 _u10_u20_U135  ( .A(_u10_u20_n2023 ), .ZN(_u10_u20_n2035 ) );
NAND3_X1 _u10_u20_U134  ( .A1(_u10_u20_n2035 ), .A2(_u10_u20_n2107 ), .A3(_u10_u20_n2108 ), .ZN(_u10_u20_n1916 ) );
INV_X1 _u10_u20_U133  ( .A(_u10_u20_n1916 ), .ZN(_u10_u20_n2093 ) );
NAND3_X1 _u10_u20_U132  ( .A1(_u10_u20_n2105 ), .A2(_u10_u20_n2106 ), .A3(_u10_u20_n2093 ), .ZN(_u10_u20_n2039 ) );
NAND2_X1 _u10_u20_U131  ( .A1(_u10_u20_n2039 ), .A2(_u10_u20_n1930 ), .ZN(_u10_u20_n2104 ) );
NAND2_X1 _u10_u20_U130  ( .A1(_u10_u20_n2103 ), .A2(_u10_u20_n2104 ), .ZN(_u10_u20_n1863 ) );
OR2_X1 _u10_u20_U129  ( .A1(_u10_u20_n1863 ), .A2(_u10_u20_n2102 ), .ZN(_u10_u20_n2099 ) );
NAND2_X1 _u10_u20_U128  ( .A1(_u10_u20_n1890 ), .A2(_u10_u20_n2101 ), .ZN(_u10_u20_n2100 ) );
NAND3_X1 _u10_u20_U127  ( .A1(_u10_u20_n2098 ), .A2(_u10_u20_n2099 ), .A3(_u10_u20_n2100 ), .ZN(_u10_u20_n2066 ) );
NAND4_X1 _u10_u20_U126  ( .A1(_u10_u20_n2095 ), .A2(_u10_u20_n2096 ), .A3(_u10_u20_n1896 ), .A4(_u10_u20_n2097 ), .ZN(_u10_u20_n2086 ) );
NOR4_X1 _u10_u20_U125  ( .A1(_u10_u20_n2093 ), .A2(_u10_u20_n2027 ), .A3(_u10_u20_n2094 ), .A4(_u10_u20_n2026 ), .ZN(_u10_u20_n1952 ) );
NOR2_X1 _u10_u20_U124  ( .A1(1'b0), .A2(_u10_u20_n1952 ), .ZN(_u10_u20_n1951 ) );
INV_X1 _u10_u20_U123  ( .A(_u10_u20_n1951 ), .ZN(_u10_u20_n2090 ) );
NAND4_X1 _u10_u20_U122  ( .A1(_u10_u20_n2089 ), .A2(_u10_u20_n2090 ), .A3(_u10_u20_n2091 ), .A4(_u10_u20_n2092 ), .ZN(_u10_u20_n1893 ) );
NOR4_X1 _u10_u20_U121  ( .A1(_u10_u20_n2086 ), .A2(_u10_u20_n1893 ), .A3(_u10_u20_n2087 ), .A4(_u10_u20_n2088 ), .ZN(_u10_u20_n2084 ) );
NOR2_X1 _u10_u20_U120  ( .A1(_u10_u20_n2084 ), .A2(_u10_u20_n2085 ), .ZN(_u10_u20_n2067 ) );
NOR2_X1 _u10_u20_U119  ( .A1(_u10_u20_n2083 ), .A2(_u10_u20_n1869 ), .ZN(_u10_u20_n2068 ) );
NAND2_X1 _u10_u20_U118  ( .A1(_u10_u20_n2081 ), .A2(_u10_u20_n2082 ), .ZN(_u10_u20_n2075 ) );
NAND2_X1 _u10_u20_U117  ( .A1(_u10_u20_n2035 ), .A2(_u10_u20_n2019 ), .ZN(_u10_u20_n2060 ) );
NAND2_X1 _u10_u20_U116  ( .A1(_u10_u20_n2080 ), .A2(_u10_u20_n2060 ), .ZN(_u10_u20_n2079 ) );
NAND2_X1 _u10_u20_U115  ( .A1(_u10_u20_n2078 ), .A2(_u10_u20_n2079 ), .ZN(_u10_u20_n2076 ) );
NAND4_X1 _u10_u20_U114  ( .A1(_u10_u20_n2075 ), .A2(_u10_u20_n2076 ), .A3(_u10_u20_n1970 ), .A4(_u10_u20_n2077 ), .ZN(_u10_u20_n2072 ) );
NOR4_X1 _u10_u20_U113  ( .A1(_u10_u20_n2072 ), .A2(_u10_u20_n2073 ), .A3(_u10_u20_n1975 ), .A4(_u10_u20_n2074 ), .ZN(_u10_u20_n2070 ) );
NOR2_X1 _u10_u20_U112  ( .A1(_u10_u20_n2070 ), .A2(_u10_u20_n2071 ), .ZN(_u10_u20_n2069 ) );
NOR4_X1 _u10_u20_U111  ( .A1(_u10_u20_n2066 ), .A2(_u10_u20_n2067 ), .A3(_u10_u20_n2068 ), .A4(_u10_u20_n2069 ), .ZN(_u10_u20_n1820 ) );
NAND2_X1 _u10_u20_U110  ( .A1(1'b0), .A2(_u10_u20_n1983 ), .ZN(_u10_u20_n2065 ) );
NAND4_X1 _u10_u20_U109  ( .A1(_u10_u20_n2065 ), .A2(_u10_u20_n2023 ), .A3(_u10_u20_n2021 ), .A4(_u10_u20_n2052 ), .ZN(_u10_u20_n2064 ) );
NAND2_X1 _u10_u20_U108  ( .A1(_u10_u20_n2063 ), .A2(_u10_u20_n2064 ), .ZN(_u10_u20_n2040 ) );
NAND4_X1 _u10_u20_U107  ( .A1(_u10_u20_n2059 ), .A2(_u10_u20_n2060 ), .A3(_u10_u20_n2061 ), .A4(_u10_u20_n2062 ), .ZN(_u10_u20_n2058 ) );
NAND2_X1 _u10_u20_U106  ( .A1(_u10_u20_n2057 ), .A2(_u10_u20_n2058 ), .ZN(_u10_u20_n2041 ) );
NOR4_X1 _u10_u20_U105  ( .A1(1'b0), .A2(_u10_u20_n2054 ), .A3(_u10_u20_n2055 ), .A4(_u10_u20_n2056 ), .ZN(_u10_u20_n2053 ) );
NAND4_X1 _u10_u20_U104  ( .A1(_u10_u20_n2021 ), .A2(_u10_u20_n2052 ), .A3(_u10_u20_n2023 ), .A4(_u10_u20_n2053 ), .ZN(_u10_u20_n1964 ) );
INV_X1 _u10_u20_U103  ( .A(_u10_u20_n1964 ), .ZN(_u10_u20_n2045 ) );
NAND2_X1 _u10_u20_U102  ( .A1(_u10_u20_n2051 ), .A2(_u10_SYNOPSYS_UNCONNECTED_7 ), .ZN(_u10_u20_n2046 ) );
NAND2_X1 _u10_u20_U101  ( .A1(_u10_u20_n2049 ), .A2(_u10_u20_n2050 ), .ZN(_u10_u20_n2047 ) );
NAND4_X1 _u10_u20_U100  ( .A1(_u10_u20_n2045 ), .A2(_u10_u20_n2046 ), .A3(_u10_u20_n2047 ), .A4(_u10_u20_n2048 ), .ZN(_u10_u20_n2044 ) );
NAND2_X1 _u10_u20_U99  ( .A1(_u10_u20_n2043 ), .A2(_u10_u20_n2044 ), .ZN(_u10_u20_n2042 ) );
NAND3_X1 _u10_u20_U98  ( .A1(_u10_u20_n2040 ), .A2(_u10_u20_n2041 ), .A3(_u10_u20_n2042 ), .ZN(_u10_u20_n2009 ) );
AND2_X1 _u10_u20_U97  ( .A1(_u10_u20_n2038 ), .A2(_u10_u20_n2039 ), .ZN(_u10_u20_n1929 ) );
NOR2_X1 _u10_u20_U96  ( .A1(_u10_u20_n1929 ), .A2(_u10_u20_n2037 ), .ZN(_u10_u20_n2010 ) );
NAND2_X1 _u10_u20_U95  ( .A1(_u10_u20_n2035 ), .A2(_u10_u20_n2036 ), .ZN(_u10_u20_n1902 ) );
NAND3_X1 _u10_u20_U94  ( .A1(_u10_u20_n1902 ), .A2(_u10_u20_n2033 ), .A3(_u10_u20_n2034 ), .ZN(_u10_u20_n1973 ) );
NOR2_X1 _u10_u20_U93  ( .A1(_u10_u20_n1978 ), .A2(_u10_u20_n1973 ), .ZN(_u10_u20_n2032 ) );
NOR2_X1 _u10_u20_U92  ( .A1(1'b0), .A2(_u10_u20_n2032 ), .ZN(_u10_u20_n2028 ) );
NOR2_X1 _u10_u20_U91  ( .A1(_u10_u20_n2030 ), .A2(_u10_u20_n2031 ), .ZN(_u10_u20_n2029 ) );
NOR4_X1 _u10_u20_U90  ( .A1(_u10_u20_n2026 ), .A2(_u10_u20_n2027 ), .A3(_u10_u20_n2028 ), .A4(_u10_u20_n2029 ), .ZN(_u10_u20_n2024 ) );
NOR2_X1 _u10_u20_U89  ( .A1(_u10_u20_n2024 ), .A2(_u10_u20_n2025 ), .ZN(_u10_u20_n2011 ) );
NAND3_X1 _u10_u20_U88  ( .A1(_u10_u20_n2021 ), .A2(_u10_u20_n2022 ), .A3(_u10_u20_n2023 ), .ZN(_u10_u20_n2020 ) );
AND2_X1 _u10_u20_U87  ( .A1(_u10_u20_n2019 ), .A2(_u10_u20_n2020 ), .ZN(_u10_u20_n1838 ) );
INV_X1 _u10_u20_U86  ( .A(_u10_u20_n2018 ), .ZN(_u10_u20_n2016 ) );
NOR4_X1 _u10_u20_U85  ( .A1(_u10_u20_n2015 ), .A2(_u10_u20_n1838 ), .A3(_u10_u20_n2016 ), .A4(_u10_u20_n2017 ), .ZN(_u10_u20_n2013 ) );
NOR2_X1 _u10_u20_U84  ( .A1(_u10_u20_n2013 ), .A2(_u10_u20_n2014 ), .ZN(_u10_u20_n2012 ) );
NOR4_X1 _u10_u20_U83  ( .A1(_u10_u20_n2009 ), .A2(_u10_u20_n2010 ), .A3(_u10_u20_n2011 ), .A4(_u10_u20_n2012 ), .ZN(_u10_u20_n1821 ) );
NAND2_X1 _u10_u20_U82  ( .A1(_u10_u20_n1924 ), .A2(_u10_u20_n2008 ), .ZN(_u10_u20_n1993 ) );
NAND2_X1 _u10_u20_U81  ( .A1(_u10_u20_n2006 ), .A2(_u10_u20_n2007 ), .ZN(_u10_u20_n1994 ) );
NAND2_X1 _u10_u20_U80  ( .A1(_u10_u20_n2004 ), .A2(_u10_u20_n2005 ), .ZN(_u10_u20_n1995 ) );
AND2_X1 _u10_u20_U79  ( .A1(_u10_u20_n2002 ), .A2(_u10_u20_n2003 ), .ZN(_u10_u20_n1998 ) );
NOR2_X1 _u10_u20_U78  ( .A1(_u10_u20_n2000 ), .A2(_u10_u20_n2001 ), .ZN(_u10_u20_n1999 ) );
NOR3_X1 _u10_u20_U77  ( .A1(_u10_u20_n1997 ), .A2(_u10_u20_n1998 ), .A3(_u10_u20_n1999 ), .ZN(_u10_u20_n1996 ) );
NAND4_X1 _u10_u20_U76  ( .A1(_u10_u20_n1993 ), .A2(_u10_u20_n1994 ), .A3(_u10_u20_n1995 ), .A4(_u10_u20_n1996 ), .ZN(_u10_u20_n1985 ) );
INV_X1 _u10_u20_U75  ( .A(_u10_u20_n1992 ), .ZN(_u10_u20_n1989 ) );
NAND3_X1 _u10_u20_U74  ( .A1(_u10_u20_n1989 ), .A2(_u10_u20_n1990 ), .A3(_u10_u20_n1991 ), .ZN(_u10_u20_n1986 ) );
NOR4_X1 _u10_u20_U73  ( .A1(_u10_u20_n1985 ), .A2(_u10_u20_n1986 ), .A3(_u10_u20_n1987 ), .A4(_u10_u20_n1988 ), .ZN(_u10_u20_n1822 ) );
INV_X1 _u10_u20_U72  ( .A(_u10_u20_n1984 ), .ZN(_u10_u20_n1980 ) );
NAND4_X1 _u10_u20_U71  ( .A1(_u10_u20_n1980 ), .A2(_u10_u20_n1981 ), .A3(_u10_u20_n1982 ), .A4(_u10_u20_n1983 ), .ZN(_u10_u20_n1941 ) );
NOR3_X1 _u10_u20_U70  ( .A1(_u10_u20_n1977 ), .A2(_u10_u20_n1978 ), .A3(_u10_u20_n1979 ), .ZN(_u10_u20_n1971 ) );
NOR4_X1 _u10_u20_U69  ( .A1(_u10_u20_n1973 ), .A2(_u10_u20_n1974 ), .A3(_u10_u20_n1975 ), .A4(_u10_u20_n1976 ), .ZN(_u10_u20_n1972 ) );
NAND4_X1 _u10_u20_U68  ( .A1(_u10_u20_n1969 ), .A2(_u10_u20_n1970 ), .A3(_u10_u20_n1971 ), .A4(_u10_u20_n1972 ), .ZN(_u10_u20_n1968 ) );
NAND2_X1 _u10_u20_U67  ( .A1(_u10_u20_n1967 ), .A2(_u10_u20_n1968 ), .ZN(_u10_u20_n1942 ) );
NAND3_X1 _u10_u20_U66  ( .A1(_u10_u20_n1964 ), .A2(_u10_u20_n1965 ), .A3(_u10_u20_n1966 ), .ZN(_u10_u20_n1943 ) );
AND4_X1 _u10_u20_U65  ( .A1(_u10_u20_n1961 ), .A2(_u10_u20_n1863 ), .A3(_u10_u20_n1962 ), .A4(_u10_u20_n1963 ), .ZN(_u10_u20_n1957 ) );
NOR2_X1 _u10_u20_U64  ( .A1(_u10_u20_n1959 ), .A2(_u10_u20_n1960 ), .ZN(_u10_u20_n1958 ) );
NOR2_X1 _u10_u20_U63  ( .A1(_u10_u20_n1957 ), .A2(_u10_u20_n1958 ), .ZN(_u10_u20_n1945 ) );
NOR2_X1 _u10_u20_U62  ( .A1(_u10_u20_n1955 ), .A2(_u10_u20_n1956 ), .ZN(_u10_u20_n1953 ) );
NOR4_X1 _u10_u20_U61  ( .A1(_u10_u20_n1952 ), .A2(_u10_u20_n1953 ), .A3(_u10_u20_n1846 ), .A4(_u10_u20_n1954 ), .ZN(_u10_u20_n1946 ) );
NOR2_X1 _u10_u20_U60  ( .A1(_u10_u20_n1950 ), .A2(_u10_u20_n1951 ), .ZN(_u10_u20_n1949 ) );
NOR2_X1 _u10_u20_U59  ( .A1(_u10_u20_n1948 ), .A2(_u10_u20_n1949 ), .ZN(_u10_u20_n1947 ) );
NOR3_X1 _u10_u20_U58  ( .A1(_u10_u20_n1945 ), .A2(_u10_u20_n1946 ), .A3(_u10_u20_n1947 ), .ZN(_u10_u20_n1944 ) );
NAND4_X1 _u10_u20_U57  ( .A1(_u10_u20_n1941 ), .A2(_u10_u20_n1942 ), .A3(_u10_u20_n1943 ), .A4(_u10_u20_n1944 ), .ZN(_u10_u20_n1824 ) );
NAND2_X1 _u10_u20_U56  ( .A1(_u10_u20_n1939 ), .A2(_u10_u20_n1940 ), .ZN(_u10_u20_n1938 ) );
NAND2_X1 _u10_u20_U55  ( .A1(_u10_u20_n1937 ), .A2(_u10_u20_n1938 ), .ZN(_u10_u20_n1903 ) );
NAND2_X1 _u10_u20_U54  ( .A1(_u10_u20_n1935 ), .A2(_u10_u20_n1936 ), .ZN(_u10_u20_n1934 ) );
NAND2_X1 _u10_u20_U53  ( .A1(_u10_u20_n1933 ), .A2(_u10_u20_n1934 ), .ZN(_u10_u20_n1931 ) );
NAND2_X1 _u10_u20_U52  ( .A1(_u10_u20_n1931 ), .A2(_u10_u20_n1932 ), .ZN(_u10_u20_n1904 ) );
NAND2_X1 _u10_u20_U51  ( .A1(_u10_u20_n1929 ), .A2(_u10_u20_n1930 ), .ZN(_u10_u20_n1927 ) );
NAND2_X1 _u10_u20_U50  ( .A1(_u10_u20_n1927 ), .A2(_u10_u20_n1928 ), .ZN(_u10_u20_n1905 ) );
NOR3_X1 _u10_u20_U49  ( .A1(_u10_u20_n1916 ), .A2(_u10_u20_n1925 ), .A3(_u10_u20_n1926 ), .ZN(_u10_u20_n1919 ) );
NOR2_X1 _u10_u20_U48  ( .A1(_u10_u20_n1923 ), .A2(_u10_u20_n1924 ), .ZN(_u10_u20_n1921 ) );
NOR2_X1 _u10_u20_U47  ( .A1(_u10_u20_n1921 ), .A2(_u10_u20_n1922 ), .ZN(_u10_u20_n1920 ) );
NOR2_X1 _u10_u20_U46  ( .A1(_u10_u20_n1919 ), .A2(_u10_u20_n1920 ), .ZN(_u10_u20_n1917 ) );
NOR2_X1 _u10_u20_U45  ( .A1(_u10_u20_n1917 ), .A2(_u10_u20_n1918 ), .ZN(_u10_u20_n1907 ) );
NOR2_X1 _u10_u20_U44  ( .A1(_u10_u20_n1915 ), .A2(_u10_u20_n1916 ), .ZN(_u10_u20_n1914 ) );
NOR2_X1 _u10_u20_U43  ( .A1(_u10_u20_n1914 ), .A2(1'b0), .ZN(_u10_u20_n1912 ) );
NOR2_X1 _u10_u20_U42  ( .A1(_u10_u20_n1912 ), .A2(_u10_u20_n1913 ), .ZN(_u10_u20_n1908 ) );
NOR2_X1 _u10_u20_U41  ( .A1(_u10_u20_n1891 ), .A2(_u10_u20_n1911 ), .ZN(_u10_u20_n1910 ) );
NOR2_X1 _u10_u20_U40  ( .A1(_u10_u20_n1910 ), .A2(_u10_u20_n1868 ), .ZN(_u10_u20_n1909 ) );
NOR3_X1 _u10_u20_U39  ( .A1(_u10_u20_n1907 ), .A2(_u10_u20_n1908 ), .A3(_u10_u20_n1909 ), .ZN(_u10_u20_n1906 ) );
NAND4_X1 _u10_u20_U38  ( .A1(_u10_u20_n1903 ), .A2(_u10_u20_n1904 ), .A3(_u10_u20_n1905 ), .A4(_u10_u20_n1906 ), .ZN(_u10_u20_n1825 ) );
NAND2_X1 _u10_u20_U37  ( .A1(_u10_u20_n1901 ), .A2(_u10_u20_n1902 ), .ZN(_u10_u20_n1900 ) );
NAND2_X1 _u10_u20_U36  ( .A1(_u10_u20_n1899 ), .A2(_u10_u20_n1900 ), .ZN(_u10_u20_n1875 ) );
OR2_X1 _u10_u20_U35  ( .A1(_u10_u20_n1847 ), .A2(_u10_u20_n1898 ), .ZN(_u10_u20_n1897 ) );
NAND2_X1 _u10_u20_U34  ( .A1(_u10_u20_n1896 ), .A2(_u10_u20_n1897 ), .ZN(_u10_u20_n1895 ) );
NAND2_X1 _u10_u20_U33  ( .A1(_u10_u20_n1894 ), .A2(_u10_u20_n1895 ), .ZN(_u10_u20_n1876 ) );
NAND2_X1 _u10_u20_U32  ( .A1(_u10_u20_n1892 ), .A2(_u10_u20_n1893 ), .ZN(_u10_u20_n1877 ) );
NOR3_X1 _u10_u20_U31  ( .A1(_u10_u20_n1884 ), .A2(_u10_u20_n1890 ), .A3(_u10_u20_n1891 ), .ZN(_u10_u20_n1889 ) );
NOR2_X1 _u10_u20_U30  ( .A1(_u10_u20_n1840 ), .A2(_u10_u20_n1889 ), .ZN(_u10_u20_n1879 ) );
NOR2_X1 _u10_u20_U29  ( .A1(_u10_u20_n1887 ), .A2(_u10_u20_n1888 ), .ZN(_u10_u20_n1880 ) );
NOR3_X1 _u10_u20_U28  ( .A1(_u10_u20_n1884 ), .A2(_u10_u20_n1885 ), .A3(_u10_u20_n1886 ), .ZN(_u10_u20_n1883 ) );
NOR2_X1 _u10_u20_U27  ( .A1(_u10_u20_n1882 ), .A2(_u10_u20_n1883 ), .ZN(_u10_u20_n1881 ) );
NOR3_X1 _u10_u20_U26  ( .A1(_u10_u20_n1879 ), .A2(_u10_u20_n1880 ), .A3(_u10_u20_n1881 ), .ZN(_u10_u20_n1878 ) );
NAND4_X1 _u10_u20_U25  ( .A1(_u10_u20_n1875 ), .A2(_u10_u20_n1876 ), .A3(_u10_u20_n1877 ), .A4(_u10_u20_n1878 ), .ZN(_u10_u20_n1826 ) );
NOR3_X1 _u10_u20_U24  ( .A1(_u10_u20_n1872 ), .A2(_u10_u20_n1873 ), .A3(_u10_u20_n1874 ), .ZN(_u10_u20_n1871 ) );
NAND4_X1 _u10_u20_U23  ( .A1(_u10_u20_n1868 ), .A2(_u10_u20_n1869 ), .A3(_u10_u20_n1870 ), .A4(_u10_u20_n1871 ), .ZN(_u10_u20_n1867 ) );
NAND2_X1 _u10_u20_U22  ( .A1(_u10_u20_n1866 ), .A2(_u10_u20_n1867 ), .ZN(_u10_u20_n1865 ) );
NAND3_X1 _u10_u20_U21  ( .A1(_u10_u20_n1863 ), .A2(_u10_u20_n1864 ), .A3(_u10_u20_n1865 ), .ZN(_u10_u20_n1862 ) );
NAND2_X1 _u10_u20_U20  ( .A1(_u10_u20_n1861 ), .A2(_u10_u20_n1862 ), .ZN(_u10_u20_n1828 ) );
NAND3_X1 _u10_u20_U19  ( .A1(_u10_u20_n1858 ), .A2(_u10_u20_n1859 ), .A3(_u10_u20_n1860 ), .ZN(_u10_u20_n1857 ) );
NAND2_X1 _u10_u20_U18  ( .A1(_u10_u20_n1856 ), .A2(_u10_u20_n1857 ), .ZN(_u10_u20_n1829 ) );
OR2_X1 _u10_u20_U17  ( .A1(_u10_u20_n1854 ), .A2(_u10_u20_n1855 ), .ZN(_u10_u20_n1830 ) );
NOR2_X1 _u10_u20_U16  ( .A1(_u10_u20_n1852 ), .A2(_u10_u20_n1853 ), .ZN(_u10_u20_n1850 ) );
NOR3_X1 _u10_u20_U15  ( .A1(_u10_u20_n1850 ), .A2(_u10_u20_n1851 ), .A3(_u10_u20_n1838 ), .ZN(_u10_u20_n1848 ) );
NOR2_X1 _u10_u20_U14  ( .A1(_u10_u20_n1848 ), .A2(_u10_u20_n1849 ), .ZN(_u10_u20_n1832 ) );
NOR2_X1 _u10_u20_U13  ( .A1(_u10_u20_n1846 ), .A2(_u10_u20_n1847 ), .ZN(_u10_u20_n1845 ) );
NOR3_X1 _u10_u20_U12  ( .A1(_u10_u20_n1844 ), .A2(1'b0), .A3(_u10_u20_n1845 ), .ZN(_u10_u20_n1842 ) );
NOR2_X1 _u10_u20_U11  ( .A1(_u10_u20_n1842 ), .A2(_u10_u20_n1843 ), .ZN(_u10_u20_n1833 ) );
NOR2_X1 _u10_u20_U10  ( .A1(_u10_u20_n1840 ), .A2(_u10_u20_n1841 ), .ZN(_u10_u20_n1839 ) );
NOR3_X1 _u10_u20_U9  ( .A1(_u10_u20_n1837 ), .A2(_u10_u20_n1838 ), .A3(_u10_u20_n1839 ), .ZN(_u10_u20_n1835 ) );
NOR2_X1 _u10_u20_U8  ( .A1(_u10_u20_n1835 ), .A2(_u10_u20_n1836 ), .ZN(_u10_u20_n1834 ) );
NOR3_X1 _u10_u20_U7  ( .A1(_u10_u20_n1832 ), .A2(_u10_u20_n1833 ), .A3(_u10_u20_n1834 ), .ZN(_u10_u20_n1831 ) );
NAND4_X1 _u10_u20_U6  ( .A1(_u10_u20_n1828 ), .A2(_u10_u20_n1829 ), .A3(_u10_u20_n1830 ), .A4(_u10_u20_n1831 ), .ZN(_u10_u20_n1827 ) );
NOR4_X1 _u10_u20_U5  ( .A1(_u10_u20_n1824 ), .A2(_u10_u20_n1825 ), .A3(_u10_u20_n1826 ), .A4(_u10_u20_n1827 ), .ZN(_u10_u20_n1823 ) );
NAND4_X1 _u10_u20_U4  ( .A1(_u10_u20_n1820 ), .A2(_u10_u20_n1821 ), .A3(_u10_u20_n1822 ), .A4(_u10_u20_n1823 ), .ZN(_u10_u20_n1818 ) );
MUX2_X1 _u10_u20_U3  ( .A(_u10_u20_n1818 ), .B(_u10_SYNOPSYS_UNCONNECTED_7 ),.S(_u10_u20_n1819 ), .Z(_u10_u20_n1812 ) );
DFFR_X1 _u10_u20_state_reg_1_  ( .D(_u10_u20_n1812 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_7 ), .QN(_u10_u20_n1814 ));
DFFR_X1 _u10_u20_state_reg_2_  ( .D(_u10_u20_n1811 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_6 ), .QN(_u10_u20_n1815 ));
DFFR_X1 _u10_u20_state_reg_3_  ( .D(_u10_u20_n1810 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_5 ), .QN(_u10_u20_n1816 ));
DFFR_X1 _u10_u20_state_reg_4_  ( .D(_u10_u20_n1809 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_4 ), .QN(_u10_u20_n1817 ));
DFFR_X1 _u10_u20_state_reg_0_  ( .D(_u10_u20_n1808 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_8 ), .QN(_u10_u20_n1813 ));
NOR2_X1 _u10_u3_U1606  ( .A1(_u10_SYNOPSYS_UNCONNECTED_11 ), .A2(_u10_u3_n1814 ), .ZN(_u10_u3_n3174 ) );
NOR3_X1 _u10_u3_U1605  ( .A1(_u10_SYNOPSYS_UNCONNECTED_10 ), .A2(_u10_u3_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_13 ), .ZN(_u10_u3_n3328 ) );
NAND2_X1 _u10_u3_U1604  ( .A1(_u10_u3_n3174 ), .A2(_u10_u3_n3328 ), .ZN(_u10_u3_n1843 ) );
INV_X1 _u10_u3_U1603  ( .A(_u10_u3_n1843 ), .ZN(_u10_u3_n2461 ) );
INV_X1 _u10_u3_U1602  ( .A(1'b0), .ZN(_u10_u3_n2466 ) );
INV_X1 _u10_u3_U1601  ( .A(1'b0), .ZN(_u10_u3_n2305 ) );
NAND2_X1 _u10_u3_U1600  ( .A1(_u10_u3_n2466 ), .A2(_u10_u3_n2305 ), .ZN(_u10_u3_n1954 ) );
INV_X1 _u10_u3_U1599  ( .A(_u10_u3_n1954 ), .ZN(_u10_u3_n2467 ) );
INV_X1 _u10_u3_U1598  ( .A(1'b0), .ZN(_u10_u3_n1936 ) );
NOR2_X1 _u10_u3_U1597  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u3_n2223 ) );
INV_X1 _u10_u3_U1596  ( .A(1'b0), .ZN(_u10_u3_n1922 ) );
NAND2_X1 _u10_u3_U1595  ( .A1(_u10_u3_n2223 ), .A2(_u10_u3_n1922 ), .ZN(_u10_u3_n2200 ) );
NOR2_X1 _u10_u3_U1594  ( .A1(_u10_u3_n2200 ), .A2(1'b0), .ZN(_u10_u3_n2502 ));
INV_X1 _u10_u3_U1593  ( .A(1'b0), .ZN(_u10_u3_n2978 ) );
INV_X1 _u10_u3_U1592  ( .A(1'b0), .ZN(_u10_u3_n3000 ) );
NAND2_X1 _u10_u3_U1591  ( .A1(_u10_u3_n2978 ), .A2(_u10_u3_n3000 ), .ZN(_u10_u3_n3356 ) );
INV_X1 _u10_u3_U1590  ( .A(1'b0), .ZN(_u10_u3_n2405 ) );
INV_X1 _u10_u3_U1589  ( .A(1'b0), .ZN(_u10_u3_n2972 ) );
NAND2_X1 _u10_u3_U1588  ( .A1(_u10_u3_n2405 ), .A2(_u10_u3_n2972 ), .ZN(_u10_u3_n2008 ) );
NOR2_X1 _u10_u3_U1587  ( .A1(_u10_u3_n3356 ), .A2(_u10_u3_n2008 ), .ZN(_u10_u3_n2195 ) );
NAND2_X1 _u10_u3_U1586  ( .A1(_u10_u3_n2502 ), .A2(_u10_u3_n2195 ), .ZN(_u10_u3_n2490 ) );
INV_X1 _u10_u3_U1585  ( .A(1'b0), .ZN(_u10_u3_n3040 ) );
INV_X1 _u10_u3_U1584  ( .A(1'b0), .ZN(_u10_u3_n3006 ) );
NAND2_X1 _u10_u3_U1583  ( .A1(_u10_u3_n3040 ), .A2(_u10_u3_n3006 ), .ZN(_u10_u3_n2508 ) );
NOR2_X1 _u10_u3_U1582  ( .A1(_u10_u3_n2508 ), .A2(1'b0), .ZN(_u10_u3_n2493 ));
INV_X1 _u10_u3_U1581  ( .A(1'b0), .ZN(_u10_u3_n2038 ) );
NAND2_X1 _u10_u3_U1580  ( .A1(_u10_u3_n2493 ), .A2(_u10_u3_n2038 ), .ZN(_u10_u3_n2174 ) );
NOR2_X1 _u10_u3_U1579  ( .A1(_u10_u3_n2490 ), .A2(_u10_u3_n2174 ), .ZN(_u10_u3_n2659 ) );
INV_X1 _u10_u3_U1578  ( .A(1'b0), .ZN(_u10_u3_n2175 ) );
NAND3_X1 _u10_u3_U1577  ( .A1(_u10_u3_n2659 ), .A2(_u10_u3_n2175 ), .A3(1'b0), .ZN(_u10_u3_n3189 ) );
NOR2_X1 _u10_u3_U1576  ( .A1(_u10_u3_n3189 ), .A2(1'b0), .ZN(_u10_u3_n2528 ));
INV_X1 _u10_u3_U1575  ( .A(1'b0), .ZN(_u10_u3_n2837 ) );
NAND2_X1 _u10_u3_U1574  ( .A1(_u10_u3_n2528 ), .A2(_u10_u3_n2837 ), .ZN(_u10_u3_n2567 ) );
INV_X1 _u10_u3_U1573  ( .A(1'b0), .ZN(_u10_u3_n2080 ) );
INV_X1 _u10_u3_U1572  ( .A(1'b0), .ZN(_u10_u3_n2166 ) );
NAND2_X1 _u10_u3_U1571  ( .A1(_u10_u3_n2080 ), .A2(_u10_u3_n2166 ), .ZN(_u10_u3_n2840 ) );
NOR2_X1 _u10_u3_U1570  ( .A1(_u10_u3_n2567 ), .A2(_u10_u3_n2840 ), .ZN(_u10_u3_n2443 ) );
INV_X1 _u10_u3_U1569  ( .A(1'b0), .ZN(_u10_u3_n2600 ) );
INV_X1 _u10_u3_U1568  ( .A(1'b0), .ZN(_u10_u3_n2836 ) );
NAND2_X1 _u10_u3_U1567  ( .A1(_u10_u3_n2600 ), .A2(_u10_u3_n2836 ), .ZN(_u10_u3_n2428 ) );
INV_X1 _u10_u3_U1566  ( .A(_u10_u3_n2428 ), .ZN(_u10_u3_n2078 ) );
NAND2_X1 _u10_u3_U1565  ( .A1(_u10_u3_n2443 ), .A2(_u10_u3_n2078 ), .ZN(_u10_u3_n2282 ) );
INV_X1 _u10_u3_U1564  ( .A(1'b0), .ZN(_u10_u3_n2874 ) );
INV_X1 _u10_u3_U1563  ( .A(1'b0), .ZN(_u10_u3_n2031 ) );
NAND2_X1 _u10_u3_U1562  ( .A1(_u10_u3_n2874 ), .A2(_u10_u3_n2031 ), .ZN(_u10_u3_n1976 ) );
NOR2_X1 _u10_u3_U1561  ( .A1(_u10_u3_n2282 ), .A2(_u10_u3_n1976 ), .ZN(_u10_u3_n2411 ) );
NAND3_X1 _u10_u3_U1560  ( .A1(_u10_u3_n2467 ), .A2(_u10_u3_n1936 ), .A3(_u10_u3_n2411 ), .ZN(_u10_u3_n2464 ) );
NAND3_X1 _u10_u3_U1559  ( .A1(_u10_u3_n2166 ), .A2(_u10_u3_n2837 ), .A3(1'b0), .ZN(_u10_u3_n3276 ) );
INV_X1 _u10_u3_U1558  ( .A(_u10_u3_n3276 ), .ZN(_u10_u3_n2442 ) );
NAND3_X1 _u10_u3_U1557  ( .A1(_u10_u3_n2836 ), .A2(_u10_u3_n2080 ), .A3(_u10_u3_n2442 ), .ZN(_u10_u3_n2838 ) );
INV_X1 _u10_u3_U1556  ( .A(_u10_u3_n2838 ), .ZN(_u10_u3_n2850 ) );
NOR2_X1 _u10_u3_U1555  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u3_n2953 ) );
NAND2_X1 _u10_u3_U1554  ( .A1(_u10_u3_n2850 ), .A2(_u10_u3_n2953 ), .ZN(_u10_u3_n2947 ) );
INV_X1 _u10_u3_U1553  ( .A(_u10_u3_n2947 ), .ZN(_u10_u3_n2420 ) );
NAND2_X1 _u10_u3_U1552  ( .A1(_u10_u3_n1936 ), .A2(_u10_u3_n2874 ), .ZN(_u10_u3_n2030 ) );
INV_X1 _u10_u3_U1551  ( .A(_u10_u3_n2030 ), .ZN(_u10_u3_n2162 ) );
NAND2_X1 _u10_u3_U1550  ( .A1(_u10_u3_n2420 ), .A2(_u10_u3_n2162 ), .ZN(_u10_u3_n2828 ) );
INV_X1 _u10_u3_U1549  ( .A(_u10_u3_n2828 ), .ZN(_u10_u3_n2551 ) );
NAND2_X1 _u10_u3_U1548  ( .A1(_u10_u3_n2551 ), .A2(_u10_u3_n2467 ), .ZN(_u10_u3_n3416 ) );
NAND2_X1 _u10_u3_U1547  ( .A1(_u10_u3_n2464 ), .A2(_u10_u3_n3416 ), .ZN(_u10_u3_n2266 ) );
INV_X1 _u10_u3_U1546  ( .A(_u10_u3_n2266 ), .ZN(_u10_u3_n3410 ) );
NAND2_X1 _u10_u3_U1545  ( .A1(1'b0), .A2(_u10_u3_n2305 ), .ZN(_u10_u3_n3411 ) );
INV_X1 _u10_u3_U1544  ( .A(_u10_u3_n3356 ), .ZN(_u10_u3_n1983 ) );
NAND3_X1 _u10_u3_U1543  ( .A1(_u10_u3_n1983 ), .A2(_u10_u3_n2405 ), .A3(1'b0), .ZN(_u10_u3_n2022 ) );
INV_X1 _u10_u3_U1542  ( .A(_u10_u3_n2022 ), .ZN(_u10_u3_n2056 ) );
INV_X1 _u10_u3_U1541  ( .A(_u10_u3_n2840 ), .ZN(_u10_u3_n2059 ) );
INV_X1 _u10_u3_U1540  ( .A(1'b0), .ZN(_u10_u3_n1965 ) );
NAND2_X1 _u10_u3_U1539  ( .A1(_u10_u3_n2837 ), .A2(_u10_u3_n1965 ), .ZN(_u10_u3_n1852 ) );
INV_X1 _u10_u3_U1538  ( .A(_u10_u3_n1852 ), .ZN(_u10_u3_n3190 ) );
INV_X1 _u10_u3_U1537  ( .A(1'b0), .ZN(_u10_u3_n1853 ) );
NAND2_X1 _u10_u3_U1536  ( .A1(_u10_u3_n3190 ), .A2(_u10_u3_n1853 ), .ZN(_u10_u3_n2687 ) );
INV_X1 _u10_u3_U1535  ( .A(_u10_u3_n2687 ), .ZN(_u10_u3_n2019 ) );
NAND2_X1 _u10_u3_U1534  ( .A1(_u10_u3_n2059 ), .A2(_u10_u3_n2019 ), .ZN(_u10_u3_n2330 ) );
NOR2_X1 _u10_u3_U1533  ( .A1(_u10_u3_n2428 ), .A2(_u10_u3_n2330 ), .ZN(_u10_u3_n2036 ) );
NAND2_X1 _u10_u3_U1532  ( .A1(_u10_u3_n2056 ), .A2(_u10_u3_n2036 ), .ZN(_u10_u3_n3379 ) );
NOR2_X1 _u10_u3_U1531  ( .A1(_u10_u3_n3379 ), .A2(_u10_u3_n2030 ), .ZN(_u10_u3_n2026 ) );
INV_X1 _u10_u3_U1530  ( .A(1'b0), .ZN(_u10_u3_n2431 ) );
NOR2_X1 _u10_u3_U1529  ( .A1(_u10_u3_n2431 ), .A2(1'b0), .ZN(_u10_u3_n3062 ));
NAND2_X1 _u10_u3_U1528  ( .A1(_u10_u3_n3062 ), .A2(_u10_u3_n2195 ), .ZN(_u10_u3_n3407 ) );
NOR3_X1 _u10_u3_U1527  ( .A1(_u10_u3_n2687 ), .A2(1'b0), .A3(_u10_u3_n3407 ),.ZN(_u10_u3_n3275 ) );
NAND3_X1 _u10_u3_U1526  ( .A1(_u10_u3_n2836 ), .A2(_u10_u3_n2080 ), .A3(_u10_u3_n3275 ), .ZN(_u10_u3_n3297 ) );
INV_X1 _u10_u3_U1525  ( .A(_u10_u3_n3297 ), .ZN(_u10_u3_n3172 ) );
NAND2_X1 _u10_u3_U1524  ( .A1(_u10_u3_n3172 ), .A2(_u10_u3_n2600 ), .ZN(_u10_u3_n2226 ) );
NOR2_X1 _u10_u3_U1523  ( .A1(_u10_u3_n2226 ), .A2(1'b0), .ZN(_u10_u3_n2307 ));
INV_X1 _u10_u3_U1522  ( .A(_u10_u3_n2490 ), .ZN(_u10_u3_n2536 ) );
NAND3_X1 _u10_u3_U1521  ( .A1(_u10_u3_n2536 ), .A2(_u10_u3_n3040 ), .A3(1'b0), .ZN(_u10_u3_n3226 ) );
NOR2_X1 _u10_u3_U1520  ( .A1(_u10_u3_n3226 ), .A2(_u10_u3_n2330 ), .ZN(_u10_u3_n2441 ) );
NAND2_X1 _u10_u3_U1519  ( .A1(_u10_u3_n2441 ), .A2(_u10_u3_n2953 ), .ZN(_u10_u3_n2579 ) );
NOR2_X1 _u10_u3_U1518  ( .A1(_u10_u3_n2579 ), .A2(_u10_u3_n2030 ), .ZN(_u10_u3_n2550 ) );
NOR3_X1 _u10_u3_U1517  ( .A1(_u10_u3_n2026 ), .A2(_u10_u3_n2307 ), .A3(_u10_u3_n2550 ), .ZN(_u10_u3_n3394 ) );
NAND2_X1 _u10_u3_U1516  ( .A1(1'b0), .A2(_u10_u3_n2978 ), .ZN(_u10_u3_n3115 ) );
NOR2_X1 _u10_u3_U1515  ( .A1(_u10_u3_n3115 ), .A2(_u10_u3_n2330 ), .ZN(_u10_u3_n3126 ) );
NAND2_X1 _u10_u3_U1514  ( .A1(_u10_u3_n2162 ), .A2(_u10_u3_n2031 ), .ZN(_u10_u3_n2686 ) );
NOR2_X1 _u10_u3_U1513  ( .A1(_u10_u3_n2686 ), .A2(_u10_u3_n2428 ), .ZN(_u10_u3_n2108 ) );
NAND2_X1 _u10_u3_U1512  ( .A1(_u10_u3_n3126 ), .A2(_u10_u3_n2108 ), .ZN(_u10_u3_n3415 ) );
NAND2_X1 _u10_u3_U1511  ( .A1(_u10_u3_n3394 ), .A2(_u10_u3_n3415 ), .ZN(_u10_u3_n3089 ) );
NAND2_X1 _u10_u3_U1510  ( .A1(_u10_u3_n3089 ), .A2(_u10_u3_n2305 ), .ZN(_u10_u3_n3414 ) );
NAND2_X1 _u10_u3_U1509  ( .A1(_u10_u3_n2466 ), .A2(_u10_u3_n3414 ), .ZN(_u10_u3_n3118 ) );
NAND2_X1 _u10_u3_U1508  ( .A1(_u10_u3_n2078 ), .A2(_u10_u3_n2080 ), .ZN(_u10_u3_n2596 ) );
NAND2_X1 _u10_u3_U1507  ( .A1(1'b0), .A2(_u10_u3_n2493 ), .ZN(_u10_u3_n1961 ) );
NOR3_X1 _u10_u3_U1506  ( .A1(_u10_u3_n2490 ), .A2(1'b0), .A3(_u10_u3_n1961 ),.ZN(_u10_u3_n2054 ) );
NAND2_X1 _u10_u3_U1505  ( .A1(_u10_u3_n2054 ), .A2(_u10_u3_n3190 ), .ZN(_u10_u3_n2061 ) );
OR2_X1 _u10_u3_U1504  ( .A1(_u10_u3_n2596 ), .A2(_u10_u3_n2061 ), .ZN(_u10_u3_n1969 ) );
NOR3_X1 _u10_u3_U1503  ( .A1(_u10_u3_n1976 ), .A2(1'b0), .A3(_u10_u3_n1969 ),.ZN(_u10_u3_n2710 ) );
NAND2_X1 _u10_u3_U1502  ( .A1(_u10_u3_n2710 ), .A2(_u10_u3_n2467 ), .ZN(_u10_u3_n2545 ) );
INV_X1 _u10_u3_U1501  ( .A(_u10_u3_n2545 ), .ZN(_u10_u3_n2087 ) );
NOR2_X1 _u10_u3_U1500  ( .A1(_u10_u3_n3118 ), .A2(_u10_u3_n2087 ), .ZN(_u10_u3_n3145 ) );
NOR2_X1 _u10_u3_U1499  ( .A1(_u10_u3_n2030 ), .A2(1'b0), .ZN(_u10_u3_n2668 ));
NAND2_X1 _u10_u3_U1498  ( .A1(1'b0), .A2(_u10_u3_n2668 ), .ZN(_u10_u3_n2163 ) );
INV_X1 _u10_u3_U1497  ( .A(_u10_u3_n2163 ), .ZN(_u10_u3_n2875 ) );
INV_X1 _u10_u3_U1496  ( .A(_u10_u3_n1976 ), .ZN(_u10_u3_n2747 ) );
NAND3_X1 _u10_u3_U1495  ( .A1(_u10_u3_n2747 ), .A2(_u10_u3_n2600 ), .A3(1'b0), .ZN(_u10_u3_n3393 ) );
NOR3_X1 _u10_u3_U1494  ( .A1(1'b0), .A2(1'b0), .A3(_u10_u3_n3393 ), .ZN(_u10_u3_n3180 ) );
INV_X1 _u10_u3_U1493  ( .A(1'b0), .ZN(_u10_u3_n2113 ) );
INV_X1 _u10_u3_U1492  ( .A(1'b0), .ZN(_u10_u3_n3066 ) );
NAND2_X1 _u10_u3_U1491  ( .A1(_u10_u3_n2175 ), .A2(_u10_u3_n3066 ), .ZN(_u10_u3_n2216 ) );
INV_X1 _u10_u3_U1490  ( .A(_u10_u3_n2659 ), .ZN(_u10_u3_n2643 ) );
NOR2_X1 _u10_u3_U1489  ( .A1(_u10_u3_n2216 ), .A2(_u10_u3_n2643 ), .ZN(_u10_u3_n2049 ) );
AND2_X1 _u10_u3_U1488  ( .A1(_u10_u3_n2049 ), .A2(_u10_u3_n1853 ), .ZN(_u10_u3_n3223 ) );
NAND2_X1 _u10_u3_U1487  ( .A1(_u10_u3_n3223 ), .A2(_u10_u3_n1965 ), .ZN(_u10_u3_n2531 ) );
NOR2_X1 _u10_u3_U1486  ( .A1(_u10_u3_n2531 ), .A2(1'b0), .ZN(_u10_u3_n2884 ));
NAND2_X1 _u10_u3_U1485  ( .A1(_u10_u3_n2884 ), .A2(_u10_u3_n2166 ), .ZN(_u10_u3_n1841 ) );
NOR2_X1 _u10_u3_U1484  ( .A1(_u10_u3_n1841 ), .A2(1'b0), .ZN(_u10_u3_n3129 ));
NAND2_X1 _u10_u3_U1483  ( .A1(_u10_u3_n3129 ), .A2(_u10_u3_n2836 ), .ZN(_u10_u3_n2842 ) );
INV_X1 _u10_u3_U1482  ( .A(_u10_u3_n2842 ), .ZN(_u10_u3_n2833 ) );
NAND2_X1 _u10_u3_U1481  ( .A1(_u10_u3_n2833 ), .A2(_u10_u3_n2600 ), .ZN(_u10_u3_n2853 ) );
INV_X1 _u10_u3_U1480  ( .A(_u10_u3_n2853 ), .ZN(_u10_u3_n2082 ) );
NAND2_X1 _u10_u3_U1479  ( .A1(_u10_u3_n2082 ), .A2(_u10_u3_n2031 ), .ZN(_u10_u3_n2274 ) );
INV_X1 _u10_u3_U1478  ( .A(_u10_u3_n2274 ), .ZN(_u10_u3_n2669 ) );
NAND3_X1 _u10_u3_U1477  ( .A1(_u10_u3_n2668 ), .A2(_u10_u3_n2113 ), .A3(_u10_u3_n2669 ), .ZN(_u10_u3_n1858 ) );
INV_X1 _u10_u3_U1476  ( .A(_u10_u3_n1858 ), .ZN(_u10_u3_n3067 ) );
NAND2_X1 _u10_u3_U1475  ( .A1(_u10_u3_n3067 ), .A2(1'b0), .ZN(_u10_u3_n2092 ) );
INV_X1 _u10_u3_U1474  ( .A(_u10_u3_n2092 ), .ZN(_u10_u3_n3294 ) );
INV_X1 _u10_u3_U1473  ( .A(1'b0), .ZN(_u10_u3_n2446 ) );
INV_X1 _u10_u3_U1472  ( .A(1'b0), .ZN(_u10_u3_n2996 ) );
NAND2_X1 _u10_u3_U1471  ( .A1(_u10_u3_n3067 ), .A2(_u10_u3_n2996 ), .ZN(_u10_u3_n1847 ) );
NOR3_X1 _u10_u3_U1470  ( .A1(_u10_u3_n2446 ), .A2(1'b0), .A3(_u10_u3_n1847 ),.ZN(_u10_u3_n3413 ) );
NOR4_X1 _u10_u3_U1469  ( .A1(_u10_u3_n2875 ), .A2(_u10_u3_n3180 ), .A3(_u10_u3_n3294 ), .A4(_u10_u3_n3413 ), .ZN(_u10_u3_n3412 ) );
NAND4_X1 _u10_u3_U1468  ( .A1(_u10_u3_n3410 ), .A2(_u10_u3_n3411 ), .A3(_u10_u3_n3145 ), .A4(_u10_u3_n3412 ), .ZN(_u10_u3_n3409 ) );
NAND2_X1 _u10_u3_U1467  ( .A1(_u10_u3_n2461 ), .A2(_u10_u3_n3409 ), .ZN(_u10_u3_n3380 ) );
NOR2_X1 _u10_u3_U1466  ( .A1(_u10_u3_n1817 ), .A2(_u10_u3_n1816 ), .ZN(_u10_u3_n3368 ) );
AND2_X1 _u10_u3_U1465  ( .A1(_u10_u3_n3368 ), .A2(_u10_u3_n1813 ), .ZN(_u10_u3_n3320 ) );
NOR2_X1 _u10_u3_U1464  ( .A1(_u10_SYNOPSYS_UNCONNECTED_12 ), .A2(_u10_u3_n1815 ), .ZN(_u10_u3_n3236 ) );
NAND2_X1 _u10_u3_U1463  ( .A1(_u10_u3_n3320 ), .A2(_u10_u3_n3236 ), .ZN(_u10_u3_n2607 ) );
INV_X1 _u10_u3_U1462  ( .A(_u10_u3_n2607 ), .ZN(_u10_u3_n1966 ) );
INV_X1 _u10_u3_U1461  ( .A(_u10_u3_n2200 ), .ZN(_u10_u3_n3216 ) );
NAND2_X1 _u10_u3_U1460  ( .A1(1'b0), .A2(_u10_u3_n3216 ), .ZN(_u10_u3_n2367 ) );
INV_X1 _u10_u3_U1459  ( .A(_u10_u3_n2367 ), .ZN(_u10_u3_n3183 ) );
NAND2_X1 _u10_u3_U1458  ( .A1(_u10_u3_n3183 ), .A2(_u10_u3_n2195 ), .ZN(_u10_u3_n2194 ) );
INV_X1 _u10_u3_U1457  ( .A(_u10_u3_n2194 ), .ZN(_u10_u3_n2055 ) );
NAND2_X1 _u10_u3_U1456  ( .A1(_u10_u3_n2055 ), .A2(_u10_u3_n1853 ), .ZN(_u10_u3_n3401 ) );
INV_X1 _u10_u3_U1455  ( .A(_u10_u3_n2531 ), .ZN(_u10_u3_n2190 ) );
INV_X1 _u10_u3_U1454  ( .A(1'b0), .ZN(_u10_u3_n3001 ) );
NAND2_X1 _u10_u3_U1453  ( .A1(_u10_u3_n3001 ), .A2(_u10_u3_n2466 ), .ZN(_u10_u3_n2156 ) );
NOR2_X1 _u10_u3_U1452  ( .A1(_u10_u3_n2166 ), .A2(_u10_u3_n2596 ), .ZN(_u10_u3_n2594 ) );
NAND2_X1 _u10_u3_U1451  ( .A1(_u10_u3_n2594 ), .A2(_u10_u3_n2031 ), .ZN(_u10_u3_n2752 ) );
INV_X1 _u10_u3_U1450  ( .A(_u10_u3_n2752 ), .ZN(_u10_u3_n2421 ) );
NAND2_X1 _u10_u3_U1449  ( .A1(_u10_u3_n2421 ), .A2(_u10_u3_n2874 ), .ZN(_u10_u3_n2033 ) );
INV_X1 _u10_u3_U1448  ( .A(_u10_u3_n2033 ), .ZN(_u10_u3_n2742 ) );
NAND3_X1 _u10_u3_U1447  ( .A1(_u10_u3_n2305 ), .A2(_u10_u3_n1936 ), .A3(_u10_u3_n2742 ), .ZN(_u10_u3_n1896 ) );
OR3_X1 _u10_u3_U1446  ( .A1(_u10_u3_n2156 ), .A2(1'b0), .A3(_u10_u3_n1896 ),.ZN(_u10_u3_n2905 ) );
NAND2_X1 _u10_u3_U1445  ( .A1(_u10_u3_n2113 ), .A2(_u10_u3_n2996 ), .ZN(_u10_u3_n2719 ) );
NOR2_X1 _u10_u3_U1444  ( .A1(_u10_u3_n2719 ), .A2(1'b0), .ZN(_u10_u3_n2941 ));
INV_X1 _u10_u3_U1443  ( .A(_u10_u3_n2941 ), .ZN(_u10_u3_n2911 ) );
NOR2_X1 _u10_u3_U1442  ( .A1(_u10_u3_n2905 ), .A2(_u10_u3_n2911 ), .ZN(_u10_u3_n3222 ) );
INV_X1 _u10_u3_U1441  ( .A(_u10_u3_n3222 ), .ZN(_u10_u3_n2695 ) );
INV_X1 _u10_u3_U1440  ( .A(_u10_u3_n2156 ), .ZN(_u10_u3_n2089 ) );
NAND3_X1 _u10_u3_U1439  ( .A1(_u10_u3_n2089 ), .A2(_u10_u3_n2446 ), .A3(_u10_u3_n3180 ), .ZN(_u10_u3_n2902 ) );
NOR2_X1 _u10_u3_U1438  ( .A1(_u10_u3_n2902 ), .A2(_u10_u3_n2911 ), .ZN(_u10_u3_n2533 ) );
INV_X1 _u10_u3_U1437  ( .A(_u10_u3_n2533 ), .ZN(_u10_u3_n2485 ) );
NAND2_X1 _u10_u3_U1436  ( .A1(_u10_u3_n2695 ), .A2(_u10_u3_n2485 ), .ZN(_u10_u3_n2721 ) );
NAND2_X1 _u10_u3_U1435  ( .A1(1'b0), .A2(_u10_u3_n2113 ), .ZN(_u10_u3_n1868 ) );
INV_X1 _u10_u3_U1434  ( .A(_u10_u3_n1868 ), .ZN(_u10_u3_n2534 ) );
NOR2_X1 _u10_u3_U1433  ( .A1(_u10_u3_n2721 ), .A2(_u10_u3_n2534 ), .ZN(_u10_u3_n3231 ) );
NAND2_X1 _u10_u3_U1432  ( .A1(_u10_u3_n2467 ), .A2(_u10_u3_n3001 ), .ZN(_u10_u3_n2303 ) );
INV_X1 _u10_u3_U1431  ( .A(_u10_u3_n2303 ), .ZN(_u10_u3_n2549 ) );
INV_X1 _u10_u3_U1430  ( .A(1'b0), .ZN(_u10_u3_n2803 ) );
NAND2_X1 _u10_u3_U1429  ( .A1(_u10_u3_n2803 ), .A2(_u10_u3_n2446 ), .ZN(_u10_u3_n1846 ) );
INV_X1 _u10_u3_U1428  ( .A(_u10_u3_n1846 ), .ZN(_u10_u3_n2667 ) );
NAND3_X1 _u10_u3_U1427  ( .A1(_u10_u3_n2549 ), .A2(_u10_u3_n2667 ), .A3(1'b0), .ZN(_u10_u3_n2739 ) );
INV_X1 _u10_u3_U1426  ( .A(_u10_u3_n2739 ), .ZN(_u10_u3_n3272 ) );
INV_X1 _u10_u3_U1425  ( .A(_u10_u3_n2719 ), .ZN(_u10_u3_n2364 ) );
NAND2_X1 _u10_u3_U1424  ( .A1(_u10_u3_n3272 ), .A2(_u10_u3_n2364 ), .ZN(_u10_u3_n2852 ) );
INV_X1 _u10_u3_U1423  ( .A(_u10_u3_n2852 ), .ZN(_u10_u3_n2214 ) );
NAND2_X1 _u10_u3_U1422  ( .A1(_u10_u3_n2875 ), .A2(_u10_u3_n2089 ), .ZN(_u10_u3_n2097 ) );
INV_X1 _u10_u3_U1421  ( .A(_u10_u3_n2097 ), .ZN(_u10_u3_n2300 ) );
NAND2_X1 _u10_u3_U1420  ( .A1(_u10_u3_n2300 ), .A2(_u10_u3_n2446 ), .ZN(_u10_u3_n2001 ) );
NOR2_X1 _u10_u3_U1419  ( .A1(_u10_u3_n2001 ), .A2(_u10_u3_n2911 ), .ZN(_u10_u3_n2877 ) );
NOR2_X1 _u10_u3_U1418  ( .A1(_u10_u3_n2214 ), .A2(_u10_u3_n2877 ), .ZN(_u10_u3_n2940 ) );
NAND2_X1 _u10_u3_U1417  ( .A1(_u10_u3_n3231 ), .A2(_u10_u3_n2940 ), .ZN(_u10_u3_n3408 ) );
NAND2_X1 _u10_u3_U1416  ( .A1(_u10_u3_n2190 ), .A2(_u10_u3_n3408 ), .ZN(_u10_u3_n3402 ) );
NOR2_X1 _u10_u3_U1415  ( .A1(_u10_u3_n2446 ), .A2(_u10_u3_n2911 ), .ZN(_u10_u3_n3059 ) );
NAND2_X1 _u10_u3_U1414  ( .A1(_u10_u3_n3059 ), .A2(_u10_u3_n2190 ), .ZN(_u10_u3_n3404 ) );
AND3_X1 _u10_u3_U1413  ( .A1(_u10_u3_n3407 ), .A2(_u10_u3_n3226 ), .A3(_u10_u3_n3115 ), .ZN(_u10_u3_n3058 ) );
NAND2_X1 _u10_u3_U1412  ( .A1(_u10_u3_n3058 ), .A2(_u10_u3_n2022 ), .ZN(_u10_u3_n3406 ) );
NAND2_X1 _u10_u3_U1411  ( .A1(_u10_u3_n1853 ), .A2(_u10_u3_n3406 ), .ZN(_u10_u3_n3405 ) );
AND3_X1 _u10_u3_U1410  ( .A1(_u10_u3_n3404 ), .A2(_u10_u3_n1965 ), .A3(_u10_u3_n3405 ), .ZN(_u10_u3_n3063 ) );
NAND2_X1 _u10_u3_U1409  ( .A1(_u10_u3_n2667 ), .A2(_u10_u3_n3001 ), .ZN(_u10_u3_n1898 ) );
INV_X1 _u10_u3_U1408  ( .A(_u10_u3_n1898 ), .ZN(_u10_u3_n2835 ) );
NAND3_X1 _u10_u3_U1407  ( .A1(_u10_u3_n2364 ), .A2(_u10_u3_n2835 ), .A3(1'b0), .ZN(_u10_u3_n1869 ) );
NOR2_X1 _u10_u3_U1406  ( .A1(_u10_u3_n1869 ), .A2(_u10_u3_n2531 ), .ZN(_u10_u3_n2761 ) );
NOR3_X1 _u10_u3_U1405  ( .A1(_u10_u3_n2761 ), .A2(_u10_u3_n2528 ), .A3(_u10_u3_n2054 ), .ZN(_u10_u3_n3403 ) );
NAND4_X1 _u10_u3_U1404  ( .A1(_u10_u3_n3401 ), .A2(_u10_u3_n3402 ), .A3(_u10_u3_n3063 ), .A4(_u10_u3_n3403 ), .ZN(_u10_u3_n3400 ) );
NAND2_X1 _u10_u3_U1403  ( .A1(_u10_u3_n1966 ), .A2(_u10_u3_n3400 ), .ZN(_u10_u3_n3381 ) );
AND2_X1 _u10_u3_U1402  ( .A1(_u10_u3_n3368 ), .A2(_u10_SYNOPSYS_UNCONNECTED_13 ), .ZN(_u10_u3_n3319 ) );
NAND2_X1 _u10_u3_U1401  ( .A1(_u10_u3_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_12 ), .ZN(_u10_u3_n1849 ) );
INV_X1 _u10_u3_U1400  ( .A(_u10_u3_n1849 ), .ZN(_u10_u3_n2183 ) );
NAND2_X1 _u10_u3_U1399  ( .A1(_u10_u3_n2884 ), .A2(_u10_u3_n2183 ), .ZN(_u10_u3_n2883 ) );
INV_X1 _u10_u3_U1398  ( .A(_u10_u3_n2883 ), .ZN(_u10_u3_n1890 ) );
INV_X1 _u10_u3_U1397  ( .A(_u10_u3_n2940 ), .ZN(_u10_u3_n3278 ) );
NAND2_X1 _u10_u3_U1396  ( .A1(_u10_u3_n1890 ), .A2(_u10_u3_n3278 ), .ZN(_u10_u3_n3382 ) );
NAND2_X1 _u10_u3_U1395  ( .A1(_u10_u3_n3059 ), .A2(_u10_u3_n2669 ), .ZN(_u10_u3_n3399 ) );
NAND2_X1 _u10_u3_U1394  ( .A1(_u10_u3_n2031 ), .A2(_u10_u3_n3399 ), .ZN(_u10_u3_n3398 ) );
NAND2_X1 _u10_u3_U1393  ( .A1(_u10_u3_n2162 ), .A2(_u10_u3_n3398 ), .ZN(_u10_u3_n3395 ) );
NAND3_X1 _u10_u3_U1392  ( .A1(_u10_u3_n2747 ), .A2(_u10_u3_n2078 ), .A3(_u10_u3_n3126 ), .ZN(_u10_u3_n3396 ) );
NAND2_X1 _u10_u3_U1391  ( .A1(_u10_u3_n2055 ), .A2(_u10_u3_n2036 ), .ZN(_u10_u3_n2285 ) );
NOR2_X1 _u10_u3_U1390  ( .A1(_u10_u3_n2285 ), .A2(_u10_u3_n2030 ), .ZN(_u10_u3_n3349 ) );
INV_X1 _u10_u3_U1389  ( .A(_u10_u3_n3349 ), .ZN(_u10_u3_n1933 ) );
INV_X1 _u10_u3_U1388  ( .A(_u10_u3_n2710 ), .ZN(_u10_u3_n3397 ) );
NAND4_X1 _u10_u3_U1387  ( .A1(_u10_u3_n3395 ), .A2(_u10_u3_n3396 ), .A3(_u10_u3_n1933 ), .A4(_u10_u3_n3397 ), .ZN(_u10_u3_n3389 ) );
NAND2_X1 _u10_u3_U1386  ( .A1(_u10_u3_n1936 ), .A2(_u10_u3_n2828 ), .ZN(_u10_u3_n3141 ) );
INV_X1 _u10_u3_U1385  ( .A(_u10_u3_n3141 ), .ZN(_u10_u3_n2302 ) );
NAND2_X1 _u10_u3_U1384  ( .A1(_u10_u3_n3394 ), .A2(_u10_u3_n2302 ), .ZN(_u10_u3_n3390 ) );
NOR2_X1 _u10_u3_U1383  ( .A1(_u10_u3_n1869 ), .A2(_u10_u3_n2274 ), .ZN(_u10_u3_n3378 ) );
INV_X1 _u10_u3_U1382  ( .A(_u10_u3_n3378 ), .ZN(_u10_u3_n2748 ) );
NOR2_X1 _u10_u3_U1381  ( .A1(1'b0), .A2(_u10_u3_n2748 ), .ZN(_u10_u3_n3391 ));
NAND2_X1 _u10_u3_U1380  ( .A1(_u10_u3_n2534 ), .A2(_u10_u3_n2669 ), .ZN(_u10_u3_n2383 ) );
INV_X1 _u10_u3_U1379  ( .A(_u10_u3_n2383 ), .ZN(_u10_u3_n1978 ) );
NAND2_X1 _u10_u3_U1378  ( .A1(_u10_u3_n1978 ), .A2(_u10_u3_n2874 ), .ZN(_u10_u3_n3392 ) );
INV_X1 _u10_u3_U1377  ( .A(_u10_u3_n2411 ), .ZN(_u10_u3_n2164 ) );
NAND4_X1 _u10_u3_U1376  ( .A1(_u10_u3_n3392 ), .A2(_u10_u3_n3393 ), .A3(_u10_u3_n2033 ), .A4(_u10_u3_n2164 ), .ZN(_u10_u3_n2476 ) );
NOR4_X1 _u10_u3_U1375  ( .A1(_u10_u3_n3389 ), .A2(_u10_u3_n3390 ), .A3(_u10_u3_n3391 ), .A4(_u10_u3_n2476 ), .ZN(_u10_u3_n3388 ) );
NAND2_X1 _u10_u3_U1374  ( .A1(_u10_u3_n3236 ), .A2(_u10_u3_n3328 ), .ZN(_u10_u3_n2025 ) );
NOR2_X1 _u10_u3_U1373  ( .A1(_u10_u3_n3388 ), .A2(_u10_u3_n2025 ), .ZN(_u10_u3_n3384 ) );
NOR2_X1 _u10_u3_U1372  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u3_n2152 ) );
NAND2_X1 _u10_u3_U1371  ( .A1(_u10_u3_n2152 ), .A2(_u10_u3_n2175 ), .ZN(_u10_u3_n2722 ) );
INV_X1 _u10_u3_U1370  ( .A(_u10_u3_n2722 ), .ZN(_u10_u3_n2588 ) );
NAND2_X1 _u10_u3_U1369  ( .A1(_u10_u3_n2549 ), .A2(_u10_u3_n3349 ), .ZN(_u10_u3_n2091 ) );
NOR2_X1 _u10_u3_U1368  ( .A1(_u10_u3_n2091 ), .A2(_u10_u3_n1846 ), .ZN(_u10_u3_n2128 ) );
NAND3_X1 _u10_u3_U1367  ( .A1(_u10_u3_n3066 ), .A2(_u10_u3_n2113 ), .A3(_u10_u3_n2128 ), .ZN(_u10_u3_n2342 ) );
INV_X1 _u10_u3_U1366  ( .A(_u10_u3_n2342 ), .ZN(_u10_u3_n3316 ) );
NAND2_X1 _u10_u3_U1365  ( .A1(_u10_u3_n2588 ), .A2(_u10_u3_n3316 ), .ZN(_u10_u3_n2142 ) );
NOR2_X1 _u10_u3_U1364  ( .A1(_u10_u3_n1954 ), .A2(_u10_u3_n1898 ), .ZN(_u10_u3_n2255 ) );
NAND2_X1 _u10_u3_U1363  ( .A1(_u10_u3_n2255 ), .A2(_u10_u3_n2996 ), .ZN(_u10_u3_n1915 ) );
INV_X1 _u10_u3_U1362  ( .A(_u10_u3_n1915 ), .ZN(_u10_u3_n2251 ) );
NAND2_X1 _u10_u3_U1361  ( .A1(_u10_u3_n2251 ), .A2(_u10_u3_n2113 ), .ZN(_u10_u3_n1925 ) );
INV_X1 _u10_u3_U1360  ( .A(_u10_u3_n2026 ), .ZN(_u10_u3_n3340 ) );
NOR3_X1 _u10_u3_U1359  ( .A1(_u10_u3_n1925 ), .A2(_u10_u3_n2216 ), .A3(_u10_u3_n3340 ), .ZN(_u10_u3_n2003 ) );
INV_X1 _u10_u3_U1358  ( .A(1'b0), .ZN(_u10_u3_n1930 ) );
NAND2_X1 _u10_u3_U1357  ( .A1(_u10_u3_n2003 ), .A2(_u10_u3_n1930 ), .ZN(_u10_u3_n3387 ) );
AND2_X1 _u10_u3_U1356  ( .A1(_u10_u3_n2142 ), .A2(_u10_u3_n3387 ), .ZN(_u10_u3_n3366 ) );
NOR3_X1 _u10_u3_U1355  ( .A1(_u10_u3_n1813 ), .A2(_u10_u3_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_9 ), .ZN(_u10_u3_n3360 ) );
NOR2_X1 _u10_u3_U1354  ( .A1(_u10_SYNOPSYS_UNCONNECTED_11 ), .A2(_u10_SYNOPSYS_UNCONNECTED_12 ), .ZN(_u10_u3_n3136 ) );
NAND2_X1 _u10_u3_U1353  ( .A1(_u10_u3_n3360 ), .A2(_u10_u3_n3136 ), .ZN(_u10_u3_n2344 ) );
NOR2_X1 _u10_u3_U1352  ( .A1(_u10_u3_n3366 ), .A2(_u10_u3_n2344 ), .ZN(_u10_u3_n3385 ) );
NOR3_X1 _u10_u3_U1351  ( .A1(_u10_SYNOPSYS_UNCONNECTED_9 ), .A2(_u10_u3_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_13 ), .ZN(_u10_u3_n3342 ) );
NAND2_X1 _u10_u3_U1350  ( .A1(_u10_u3_n3342 ), .A2(_u10_u3_n3136 ), .ZN(_u10_u3_n2584 ) );
NOR2_X1 _u10_u3_U1349  ( .A1(_u10_u3_n2584 ), .A2(1'b0), .ZN(_u10_u3_n2139 ));
INV_X1 _u10_u3_U1348  ( .A(_u10_u3_n2216 ), .ZN(_u10_u3_n2106 ) );
AND2_X1 _u10_u3_U1347  ( .A1(_u10_u3_n2152 ), .A2(_u10_u3_n2106 ), .ZN(_u10_u3_n2336 ) );
NAND2_X1 _u10_u3_U1346  ( .A1(_u10_u3_n2139 ), .A2(_u10_u3_n2336 ), .ZN(_u10_u3_n2365 ) );
INV_X1 _u10_u3_U1345  ( .A(_u10_u3_n2365 ), .ZN(_u10_u3_n2004 ) );
AND2_X1 _u10_u3_U1344  ( .A1(_u10_u3_n2877 ), .A2(_u10_u3_n2004 ), .ZN(_u10_u3_n3386 ) );
NOR3_X1 _u10_u3_U1343  ( .A1(_u10_u3_n3384 ), .A2(_u10_u3_n3385 ), .A3(_u10_u3_n3386 ), .ZN(_u10_u3_n3383 ) );
NAND4_X1 _u10_u3_U1342  ( .A1(_u10_u3_n3380 ), .A2(_u10_u3_n3381 ), .A3(_u10_u3_n3382 ), .A4(_u10_u3_n3383 ), .ZN(_u10_u3_n3191 ) );
NAND2_X1 _u10_u3_U1341  ( .A1(_u10_u3_n2285 ), .A2(_u10_u3_n3379 ), .ZN(_u10_u3_n1975 ) );
NOR3_X1 _u10_u3_U1340  ( .A1(_u10_u3_n3378 ), .A2(1'b0), .A3(_u10_u3_n1975 ),.ZN(_u10_u3_n3122 ) );
AND4_X1 _u10_u3_U1339  ( .A1(_u10_u3_n2752 ), .A2(_u10_u3_n2383 ), .A3(_u10_u3_n1969 ), .A4(_u10_u3_n3122 ), .ZN(_u10_u3_n3377 ) );
NOR2_X1 _u10_u3_U1338  ( .A1(_u10_u3_n1814 ), .A2(_u10_u3_n1815 ), .ZN(_u10_u3_n3147 ) );
NAND2_X1 _u10_u3_U1337  ( .A1(_u10_u3_n3328 ), .A2(_u10_u3_n3147 ), .ZN(_u10_u3_n2359 ) );
NOR2_X1 _u10_u3_U1336  ( .A1(_u10_u3_n3377 ), .A2(_u10_u3_n2359 ), .ZN(_u10_u3_n3362 ) );
INV_X1 _u10_u3_U1335  ( .A(_u10_u3_n2008 ), .ZN(_u10_u3_n3097 ) );
NOR3_X1 _u10_u3_U1334  ( .A1(_u10_SYNOPSYS_UNCONNECTED_9 ), .A2(_u10_u3_n1813 ), .A3(_u10_SYNOPSYS_UNCONNECTED_10 ), .ZN(_u10_u3_n3269 ) );
NAND2_X1 _u10_u3_U1333  ( .A1(_u10_u3_n3269 ), .A2(_u10_u3_n3136 ), .ZN(_u10_u3_n3109 ) );
INV_X1 _u10_u3_U1332  ( .A(_u10_u3_n3109 ), .ZN(_u10_u3_n2999 ) );
INV_X1 _u10_u3_U1331  ( .A(_u10_u3_n2508 ), .ZN(_u10_u3_n2103 ) );
NAND2_X1 _u10_u3_U1330  ( .A1(_u10_u3_n2336 ), .A2(_u10_u3_n2103 ), .ZN(_u10_u3_n2249 ) );
NOR2_X1 _u10_u3_U1329  ( .A1(_u10_u3_n2249 ), .A2(1'b0), .ZN(_u10_u3_n1866 ));
NAND2_X1 _u10_u3_U1328  ( .A1(_u10_u3_n1866 ), .A2(_u10_u3_n1922 ), .ZN(_u10_u3_n2632 ) );
INV_X1 _u10_u3_U1327  ( .A(_u10_u3_n2223 ), .ZN(_u10_u3_n1918 ) );
NOR2_X1 _u10_u3_U1326  ( .A1(_u10_u3_n2632 ), .A2(_u10_u3_n1918 ), .ZN(_u10_u3_n1981 ) );
NAND3_X1 _u10_u3_U1325  ( .A1(_u10_u3_n3097 ), .A2(_u10_u3_n2999 ), .A3(_u10_u3_n1981 ), .ZN(_u10_u3_n3034 ) );
NOR3_X1 _u10_u3_U1324  ( .A1(_u10_SYNOPSYS_UNCONNECTED_10 ), .A2(_u10_SYNOPSYS_UNCONNECTED_9 ), .A3(_u10_SYNOPSYS_UNCONNECTED_13 ),.ZN(_u10_u3_n3302 ) );
NAND2_X1 _u10_u3_U1323  ( .A1(_u10_u3_n3302 ), .A2(_u10_u3_n3174 ), .ZN(_u10_u3_n3162 ) );
INV_X1 _u10_u3_U1322  ( .A(_u10_u3_n3162 ), .ZN(_u10_u3_n2979 ) );
NAND2_X1 _u10_u3_U1321  ( .A1(_u10_u3_n2979 ), .A2(_u10_u3_n2972 ), .ZN(_u10_u3_n1984 ) );
AND2_X1 _u10_u3_U1320  ( .A1(_u10_u3_n3302 ), .A2(_u10_u3_n3136 ), .ZN(_u10_u3_n2977 ) );
NAND3_X1 _u10_u3_U1319  ( .A1(_u10_u3_n2977 ), .A2(_u10_u3_n3000 ), .A3(_u10_u3_n3097 ), .ZN(_u10_u3_n3376 ) );
NAND2_X1 _u10_u3_U1318  ( .A1(_u10_u3_n1984 ), .A2(_u10_u3_n3376 ), .ZN(_u10_u3_n3375 ) );
NAND2_X1 _u10_u3_U1317  ( .A1(_u10_u3_n1981 ), .A2(_u10_u3_n3375 ), .ZN(_u10_u3_n2798 ) );
NAND2_X1 _u10_u3_U1316  ( .A1(_u10_u3_n3034 ), .A2(_u10_u3_n2798 ), .ZN(_u10_u3_n2007 ) );
NAND2_X1 _u10_u3_U1315  ( .A1(_u10_u3_n3269 ), .A2(_u10_u3_n3147 ), .ZN(_u10_u3_n2102 ) );
NOR2_X1 _u10_u3_U1314  ( .A1(_u10_u3_n2249 ), .A2(_u10_u3_n2102 ), .ZN(_u10_u3_n3323 ) );
INV_X1 _u10_u3_U1313  ( .A(_u10_u3_n3323 ), .ZN(_u10_u3_n3374 ) );
INV_X1 _u10_u3_U1312  ( .A(_u10_u3_n2344 ), .ZN(_u10_u3_n2002 ) );
NAND2_X1 _u10_u3_U1311  ( .A1(_u10_u3_n2336 ), .A2(_u10_u3_n2002 ), .ZN(_u10_u3_n3225 ) );
NAND2_X1 _u10_u3_U1310  ( .A1(_u10_u3_n3374 ), .A2(_u10_u3_n3225 ), .ZN(_u10_u3_n2488 ) );
NAND2_X1 _u10_u3_U1309  ( .A1(_u10_u3_n3342 ), .A2(_u10_u3_n3236 ), .ZN(_u10_u3_n2253 ) );
NOR2_X1 _u10_u3_U1308  ( .A1(_u10_u3_n2253 ), .A2(1'b0), .ZN(_u10_u3_n1885 ));
NAND2_X1 _u10_u3_U1307  ( .A1(_u10_u3_n3360 ), .A2(_u10_u3_n3174 ), .ZN(_u10_u3_n2254 ) );
INV_X1 _u10_u3_U1306  ( .A(_u10_u3_n2254 ), .ZN(_u10_u3_n2986 ) );
NAND2_X1 _u10_u3_U1305  ( .A1(_u10_u3_n2106 ), .A2(_u10_u3_n2986 ), .ZN(_u10_u3_n1913 ) );
INV_X1 _u10_u3_U1304  ( .A(_u10_u3_n1913 ), .ZN(_u10_u3_n2377 ) );
OR4_X1 _u10_u3_U1303  ( .A1(_u10_u3_n2007 ), .A2(_u10_u3_n2488 ), .A3(_u10_u3_n1885 ), .A4(_u10_u3_n2377 ), .ZN(_u10_u3_n3373 ) );
NAND2_X1 _u10_u3_U1302  ( .A1(_u10_u3_n2534 ), .A2(_u10_u3_n3373 ), .ZN(_u10_u3_n3370 ) );
NAND2_X1 _u10_u3_U1301  ( .A1(_u10_u3_n3342 ), .A2(_u10_u3_n3174 ), .ZN(_u10_u3_n2037 ) );
NAND2_X1 _u10_u3_U1300  ( .A1(_u10_u3_n2037 ), .A2(_u10_u3_n2254 ), .ZN(_u10_u3_n3372 ) );
NAND2_X1 _u10_u3_U1299  ( .A1(_u10_u3_n2003 ), .A2(_u10_u3_n3372 ), .ZN(_u10_u3_n3371 ) );
NAND2_X1 _u10_u3_U1298  ( .A1(_u10_u3_n3370 ), .A2(_u10_u3_n3371 ), .ZN(_u10_u3_n3363 ) );
NOR2_X1 _u10_u3_U1297  ( .A1(_u10_u3_n2490 ), .A2(_u10_u3_n1961 ), .ZN(_u10_u3_n3369 ) );
NAND2_X1 _u10_u3_U1296  ( .A1(_u10_u3_n2534 ), .A2(_u10_u3_n2049 ), .ZN(_u10_u3_n2646 ) );
INV_X1 _u10_u3_U1295  ( .A(_u10_u3_n2646 ), .ZN(_u10_u3_n3055 ) );
NOR2_X1 _u10_u3_U1294  ( .A1(_u10_u3_n3369 ), .A2(_u10_u3_n3055 ), .ZN(_u10_u3_n3367 ) );
NAND2_X1 _u10_u3_U1293  ( .A1(_u10_u3_n3368 ), .A2(_u10_u3_n3147 ), .ZN(_u10_u3_n2495 ) );
NOR2_X1 _u10_u3_U1292  ( .A1(_u10_u3_n3367 ), .A2(_u10_u3_n2495 ), .ZN(_u10_u3_n3364 ) );
INV_X1 _u10_u3_U1291  ( .A(_u10_u3_n2139 ), .ZN(_u10_u3_n3254 ) );
NOR2_X1 _u10_u3_U1290  ( .A1(_u10_u3_n3366 ), .A2(_u10_u3_n3254 ), .ZN(_u10_u3_n3365 ) );
NOR4_X1 _u10_u3_U1289  ( .A1(_u10_u3_n3362 ), .A2(_u10_u3_n3363 ), .A3(_u10_u3_n3364 ), .A4(_u10_u3_n3365 ), .ZN(_u10_u3_n3305 ) );
NAND2_X1 _u10_u3_U1288  ( .A1(_u10_u3_n3302 ), .A2(_u10_u3_n3147 ), .ZN(_u10_u3_n2980 ) );
NAND2_X1 _u10_u3_U1287  ( .A1(_u10_u3_n2102 ), .A2(_u10_u3_n2980 ), .ZN(_u10_u3_n2177 ) );
NAND2_X1 _u10_u3_U1286  ( .A1(_u10_u3_n2003 ), .A2(_u10_u3_n2493 ), .ZN(_u10_u3_n1962 ) );
NAND2_X1 _u10_u3_U1285  ( .A1(_u10_u3_n1961 ), .A2(_u10_u3_n1962 ), .ZN(_u10_u3_n3361 ) );
NAND2_X1 _u10_u3_U1284  ( .A1(_u10_u3_n2177 ), .A2(_u10_u3_n3361 ), .ZN(_u10_u3_n3357 ) );
NAND2_X1 _u10_u3_U1283  ( .A1(_u10_u3_n3236 ), .A2(_u10_u3_n3360 ), .ZN(_u10_u3_n1859 ) );
INV_X1 _u10_u3_U1282  ( .A(_u10_u3_n1859 ), .ZN(_u10_u3_n2256 ) );
NAND3_X1 _u10_u3_U1281  ( .A1(_u10_u3_n2256 ), .A2(_u10_u3_n2113 ), .A3(_u10_u3_n2128 ), .ZN(_u10_u3_n3358 ) );
NOR2_X1 _u10_u3_U1280  ( .A1(_u10_u3_n2877 ), .A2(_u10_u3_n3222 ), .ZN(_u10_u3_n3347 ) );
NAND2_X1 _u10_u3_U1279  ( .A1(_u10_u3_n3347 ), .A2(_u10_u3_n1869 ), .ZN(_u10_u3_n2005 ) );
NAND2_X1 _u10_u3_U1278  ( .A1(_u10_u3_n2488 ), .A2(_u10_u3_n2005 ), .ZN(_u10_u3_n3359 ) );
NAND3_X1 _u10_u3_U1277  ( .A1(_u10_u3_n3357 ), .A2(_u10_u3_n3358 ), .A3(_u10_u3_n3359 ), .ZN(_u10_u3_n3352 ) );
NAND2_X1 _u10_u3_U1276  ( .A1(_u10_u3_n3320 ), .A2(_u10_u3_n3136 ), .ZN(_u10_u3_n2356 ) );
INV_X1 _u10_u3_U1275  ( .A(_u10_u3_n2356 ), .ZN(_u10_u3_n2830 ) );
NAND2_X1 _u10_u3_U1274  ( .A1(_u10_u3_n2830 ), .A2(_u10_u3_n2836 ), .ZN(_u10_u3_n2291 ) );
NOR3_X1 _u10_u3_U1273  ( .A1(_u10_u3_n2291 ), .A2(_u10_u3_n2330 ), .A3(_u10_u3_n2022 ), .ZN(_u10_u3_n3353 ) );
INV_X1 _u10_u3_U1272  ( .A(_u10_u3_n1925 ), .ZN(_u10_u3_n2105 ) );
AND2_X1 _u10_u3_U1271  ( .A1(_u10_u3_n2108 ), .A2(_u10_u3_n2105 ), .ZN(_u10_u3_n2915 ) );
INV_X1 _u10_u3_U1270  ( .A(_u10_u3_n2330 ), .ZN(_u10_u3_n2107 ) );
NAND2_X1 _u10_u3_U1269  ( .A1(_u10_u3_n2915 ), .A2(_u10_u3_n2107 ), .ZN(_u10_u3_n2203 ) );
INV_X1 _u10_u3_U1268  ( .A(_u10_u3_n2203 ), .ZN(_u10_u3_n1982 ) );
NAND2_X1 _u10_u3_U1267  ( .A1(_u10_u3_n1982 ), .A2(_u10_u3_n2536 ), .ZN(_u10_u3_n2587 ) );
INV_X1 _u10_u3_U1266  ( .A(_u10_u3_n2587 ), .ZN(_u10_u3_n2697 ) );
NAND3_X1 _u10_u3_U1265  ( .A1(_u10_u3_n2697 ), .A2(_u10_u3_n2493 ), .A3(_u10_u3_n2377 ), .ZN(_u10_u3_n2412 ) );
INV_X1 _u10_u3_U1264  ( .A(_u10_u3_n2412 ), .ZN(_u10_u3_n3354 ) );
NAND2_X1 _u10_u3_U1263  ( .A1(_u10_u3_n3174 ), .A2(_u10_u3_n3269 ), .ZN(_u10_u3_n2375 ) );
INV_X1 _u10_u3_U1262  ( .A(_u10_u3_n2375 ), .ZN(_u10_u3_n2507 ) );
NAND2_X1 _u10_u3_U1261  ( .A1(_u10_u3_n1981 ), .A2(_u10_u3_n2507 ), .ZN(_u10_u3_n2621 ) );
NOR4_X1 _u10_u3_U1260  ( .A1(1'b0), .A2(_u10_u3_n3356 ), .A3(_u10_u3_n2203 ),.A4(_u10_u3_n2621 ), .ZN(_u10_u3_n3355 ) );
NOR4_X1 _u10_u3_U1259  ( .A1(_u10_u3_n3352 ), .A2(_u10_u3_n3353 ), .A3(_u10_u3_n3354 ), .A4(_u10_u3_n3355 ), .ZN(_u10_u3_n3306 ) );
NOR2_X1 _u10_u3_U1258  ( .A1(_u10_u3_n2842 ), .A2(_u10_u3_n2356 ), .ZN(_u10_u3_n1891 ) );
INV_X1 _u10_u3_U1257  ( .A(_u10_u3_n1869 ), .ZN(_u10_u3_n2885 ) );
NAND2_X1 _u10_u3_U1256  ( .A1(_u10_u3_n1891 ), .A2(_u10_u3_n2885 ), .ZN(_u10_u3_n3330 ) );
NAND2_X1 _u10_u3_U1255  ( .A1(_u10_u3_n2761 ), .A2(_u10_u3_n2837 ), .ZN(_u10_u3_n3351 ) );
NAND3_X1 _u10_u3_U1254  ( .A1(_u10_u3_n2884 ), .A2(_u10_u3_n2080 ), .A3(_u10_u3_n2915 ), .ZN(_u10_u3_n2762 ) );
NAND2_X1 _u10_u3_U1253  ( .A1(_u10_u3_n2055 ), .A2(_u10_u3_n2019 ), .ZN(_u10_u3_n3259 ) );
NAND4_X1 _u10_u3_U1252  ( .A1(_u10_u3_n3351 ), .A2(_u10_u3_n2762 ), .A3(_u10_u3_n2061 ), .A4(_u10_u3_n3259 ), .ZN(_u10_u3_n3350 ) );
NAND2_X1 _u10_u3_U1251  ( .A1(_u10_u3_n2183 ), .A2(_u10_u3_n3350 ), .ZN(_u10_u3_n3331 ) );
NAND2_X1 _u10_u3_U1250  ( .A1(_u10_u3_n3349 ), .A2(_u10_u3_n2305 ), .ZN(_u10_u3_n3348 ) );
NAND2_X1 _u10_u3_U1249  ( .A1(_u10_u3_n1896 ), .A2(_u10_u3_n3348 ), .ZN(_u10_u3_n3176 ) );
NAND2_X1 _u10_u3_U1248  ( .A1(_u10_u3_n2461 ), .A2(_u10_u3_n3176 ), .ZN(_u10_u3_n3332 ) );
INV_X1 _u10_u3_U1247  ( .A(_u10_u3_n2495 ), .ZN(_u10_u3_n2063 ) );
NAND2_X1 _u10_u3_U1246  ( .A1(_u10_u3_n2049 ), .A2(_u10_u3_n2063 ), .ZN(_u10_u3_n2886 ) );
NOR2_X1 _u10_u3_U1245  ( .A1(_u10_u3_n3347 ), .A2(_u10_u3_n2886 ), .ZN(_u10_u3_n3334 ) );
NAND2_X1 _u10_u3_U1244  ( .A1(1'b0), .A2(_u10_u3_n2835 ), .ZN(_u10_u3_n3344 ) );
NAND2_X1 _u10_u3_U1243  ( .A1(_u10_u3_n2001 ), .A2(_u10_u3_n2905 ), .ZN(_u10_u3_n3346 ) );
NAND2_X1 _u10_u3_U1242  ( .A1(_u10_u3_n3346 ), .A2(_u10_u3_n2803 ), .ZN(_u10_u3_n3345 ) );
NAND2_X1 _u10_u3_U1241  ( .A1(_u10_u3_n2087 ), .A2(_u10_u3_n2835 ), .ZN(_u10_u3_n2413 ) );
INV_X1 _u10_u3_U1240  ( .A(_u10_u3_n2128 ), .ZN(_u10_u3_n2235 ) );
NAND4_X1 _u10_u3_U1239  ( .A1(_u10_u3_n3344 ), .A2(_u10_u3_n3345 ), .A3(_u10_u3_n2413 ), .A4(_u10_u3_n2235 ), .ZN(_u10_u3_n3329 ) );
NOR2_X1 _u10_u3_U1238  ( .A1(_u10_u3_n1915 ), .A2(_u10_u3_n3340 ), .ZN(_u10_u3_n3343 ) );
NOR3_X1 _u10_u3_U1237  ( .A1(_u10_u3_n3329 ), .A2(1'b0), .A3(_u10_u3_n3343 ),.ZN(_u10_u3_n3341 ) );
NAND2_X1 _u10_u3_U1236  ( .A1(_u10_u3_n3342 ), .A2(_u10_u3_n3147 ), .ZN(_u10_u3_n2688 ) );
NOR2_X1 _u10_u3_U1235  ( .A1(_u10_u3_n3341 ), .A2(_u10_u3_n2688 ), .ZN(_u10_u3_n3335 ) );
NOR2_X1 _u10_u3_U1234  ( .A1(_u10_u3_n2256 ), .A2(_u10_u3_n1885 ), .ZN(_u10_u3_n2689 ) );
NOR2_X1 _u10_u3_U1233  ( .A1(1'b0), .A2(_u10_u3_n2413 ), .ZN(_u10_u3_n3338 ));
NOR2_X1 _u10_u3_U1232  ( .A1(_u10_u3_n1925 ), .A2(_u10_u3_n3340 ), .ZN(_u10_u3_n3339 ) );
NOR3_X1 _u10_u3_U1231  ( .A1(_u10_u3_n2005 ), .A2(_u10_u3_n3338 ), .A3(_u10_u3_n3339 ), .ZN(_u10_u3_n3337 ) );
NOR2_X1 _u10_u3_U1230  ( .A1(_u10_u3_n2689 ), .A2(_u10_u3_n3337 ), .ZN(_u10_u3_n3336 ) );
NOR3_X1 _u10_u3_U1229  ( .A1(_u10_u3_n3334 ), .A2(_u10_u3_n3335 ), .A3(_u10_u3_n3336 ), .ZN(_u10_u3_n3333 ) );
NAND4_X1 _u10_u3_U1228  ( .A1(_u10_u3_n3330 ), .A2(_u10_u3_n3331 ), .A3(_u10_u3_n3332 ), .A4(_u10_u3_n3333 ), .ZN(_u10_u3_n3308 ) );
NAND3_X1 _u10_u3_U1227  ( .A1(_u10_SYNOPSYS_UNCONNECTED_13 ), .A2(_u10_SYNOPSYS_UNCONNECTED_10 ), .A3(_u10_u3_n3147 ), .ZN(_u10_u3_n2126 ) );
INV_X1 _u10_u3_U1226  ( .A(_u10_u3_n2126 ), .ZN(_u10_u3_n2329 ) );
NAND2_X1 _u10_u3_U1225  ( .A1(_u10_u3_n2329 ), .A2(_u10_u3_n3329 ), .ZN(_u10_u3_n3324 ) );
NAND2_X1 _u10_u3_U1224  ( .A1(_u10_u3_n3328 ), .A2(_u10_u3_n3136 ), .ZN(_u10_u3_n2000 ) );
INV_X1 _u10_u3_U1223  ( .A(_u10_u3_n2000 ), .ZN(_u10_u3_n2445 ) );
NAND3_X1 _u10_u3_U1222  ( .A1(_u10_u3_n2446 ), .A2(_u10_u3_n3001 ), .A3(_u10_u3_n2087 ), .ZN(_u10_u3_n3327 ) );
NAND2_X1 _u10_u3_U1221  ( .A1(_u10_u3_n3327 ), .A2(_u10_u3_n2905 ), .ZN(_u10_u3_n2500 ) );
NAND2_X1 _u10_u3_U1220  ( .A1(_u10_u3_n2445 ), .A2(_u10_u3_n2500 ), .ZN(_u10_u3_n3325 ) );
NAND2_X1 _u10_u3_U1219  ( .A1(1'b0), .A2(_u10_u3_n2979 ), .ZN(_u10_u3_n3326 ) );
NAND3_X1 _u10_u3_U1218  ( .A1(_u10_u3_n3324 ), .A2(_u10_u3_n3325 ), .A3(_u10_u3_n3326 ), .ZN(_u10_u3_n3309 ) );
AND2_X1 _u10_u3_U1217  ( .A1(_u10_u3_n2877 ), .A2(_u10_u3_n3223 ), .ZN(_u10_u3_n2858 ) );
NAND2_X1 _u10_u3_U1216  ( .A1(_u10_u3_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_11 ), .ZN(_u10_u3_n2346 ) );
INV_X1 _u10_u3_U1215  ( .A(_u10_u3_n2346 ), .ZN(_u10_u3_n2043 ) );
NAND2_X1 _u10_u3_U1214  ( .A1(_u10_u3_n2858 ), .A2(_u10_u3_n2043 ), .ZN(_u10_u3_n3321 ) );
NAND2_X1 _u10_u3_U1213  ( .A1(_u10_u3_n1982 ), .A2(_u10_u3_n2195 ), .ZN(_u10_u3_n3268 ) );
INV_X1 _u10_u3_U1212  ( .A(_u10_u3_n3268 ), .ZN(_u10_u3_n2222 ) );
NAND3_X1 _u10_u3_U1211  ( .A1(_u10_u3_n3323 ), .A2(_u10_u3_n3216 ), .A3(_u10_u3_n2222 ), .ZN(_u10_u3_n3322 ) );
NAND2_X1 _u10_u3_U1210  ( .A1(_u10_u3_n3321 ), .A2(_u10_u3_n3322 ), .ZN(_u10_u3_n2374 ) );
NAND2_X1 _u10_u3_U1209  ( .A1(_u10_u3_n3320 ), .A2(_u10_u3_n3174 ), .ZN(_u10_u3_n2014 ) );
NOR2_X1 _u10_u3_U1208  ( .A1(_u10_u3_n1841 ), .A2(_u10_u3_n2014 ), .ZN(_u10_u3_n2813 ) );
NAND2_X1 _u10_u3_U1207  ( .A1(_u10_u3_n2813 ), .A2(_u10_u3_n2534 ), .ZN(_u10_u3_n3310 ) );
NAND2_X1 _u10_u3_U1206  ( .A1(_u10_u3_n3319 ), .A2(_u10_u3_n3136 ), .ZN(_u10_u3_n1836 ) );
INV_X1 _u10_u3_U1205  ( .A(_u10_u3_n1836 ), .ZN(_u10_u3_n2815 ) );
NAND2_X1 _u10_u3_U1204  ( .A1(_u10_u3_n2534 ), .A2(_u10_u3_n3129 ), .ZN(_u10_u3_n2439 ) );
NAND2_X1 _u10_u3_U1203  ( .A1(_u10_u3_n2055 ), .A2(_u10_u3_n2107 ), .ZN(_u10_u3_n2062 ) );
NAND2_X1 _u10_u3_U1202  ( .A1(_u10_u3_n2439 ), .A2(_u10_u3_n2062 ), .ZN(_u10_u3_n3318 ) );
NAND2_X1 _u10_u3_U1201  ( .A1(_u10_u3_n2815 ), .A2(_u10_u3_n3318 ), .ZN(_u10_u3_n3311 ) );
NAND2_X1 _u10_u3_U1200  ( .A1(_u10_u3_n2986 ), .A2(_u10_u3_n2175 ), .ZN(_u10_u3_n3317 ) );
NAND2_X1 _u10_u3_U1199  ( .A1(_u10_u3_n2253 ), .A2(_u10_u3_n3317 ), .ZN(_u10_u3_n3157 ) );
NAND2_X1 _u10_u3_U1198  ( .A1(_u10_u3_n3316 ), .A2(_u10_u3_n3157 ), .ZN(_u10_u3_n3312 ) );
NOR2_X1 _u10_u3_U1197  ( .A1(_u10_u3_n2495 ), .A2(_u10_u3_n2194 ), .ZN(_u10_u3_n3314 ) );
NOR2_X1 _u10_u3_U1196  ( .A1(_u10_u3_n2375 ), .A2(_u10_u3_n2367 ), .ZN(_u10_u3_n3315 ) );
NOR2_X1 _u10_u3_U1195  ( .A1(_u10_u3_n3314 ), .A2(_u10_u3_n3315 ), .ZN(_u10_u3_n3313 ) );
NAND4_X1 _u10_u3_U1194  ( .A1(_u10_u3_n3310 ), .A2(_u10_u3_n3311 ), .A3(_u10_u3_n3312 ), .A4(_u10_u3_n3313 ), .ZN(_u10_u3_n2315 ) );
NOR4_X1 _u10_u3_U1193  ( .A1(_u10_u3_n3308 ), .A2(_u10_u3_n3309 ), .A3(_u10_u3_n2374 ), .A4(_u10_u3_n2315 ), .ZN(_u10_u3_n3307 ) );
NAND3_X1 _u10_u3_U1192  ( .A1(_u10_u3_n3305 ), .A2(_u10_u3_n3306 ), .A3(_u10_u3_n3307 ), .ZN(_u10_u3_n1987 ) );
AND2_X1 _u10_u3_U1191  ( .A1(1'b0), .A2(_u10_u3_n2977 ), .ZN(_u10_u3_n3240 ));
NAND2_X1 _u10_u3_U1190  ( .A1(_u10_u3_n1891 ), .A2(_u10_u3_n2534 ), .ZN(_u10_u3_n3303 ) );
NAND4_X1 _u10_u3_U1189  ( .A1(_u10_u3_n1982 ), .A2(_u10_u3_n2659 ), .A3(_u10_u3_n2256 ), .A4(_u10_u3_n2175 ), .ZN(_u10_u3_n3304 ) );
AND2_X1 _u10_u3_U1188  ( .A1(_u10_u3_n3303 ), .A2(_u10_u3_n3304 ), .ZN(_u10_u3_n2612 ) );
NAND2_X1 _u10_u3_U1187  ( .A1(_u10_u3_n3302 ), .A2(_u10_u3_n3236 ), .ZN(_u10_u3_n2985 ) );
OR2_X1 _u10_u3_U1186  ( .A1(_u10_u3_n2431 ), .A2(_u10_u3_n2985 ), .ZN(_u10_u3_n3299 ) );
OR2_X1 _u10_u3_U1185  ( .A1(_u10_u3_n2282 ), .A2(_u10_u3_n2359 ), .ZN(_u10_u3_n3300 ) );
NAND2_X1 _u10_u3_U1184  ( .A1(_u10_u3_n1890 ), .A2(_u10_u3_n2534 ), .ZN(_u10_u3_n3301 ) );
NAND4_X1 _u10_u3_U1183  ( .A1(_u10_u3_n2612 ), .A2(_u10_u3_n3299 ), .A3(_u10_u3_n3300 ), .A4(_u10_u3_n3301 ), .ZN(_u10_u3_n3279 ) );
INV_X1 _u10_u3_U1182  ( .A(_u10_u3_n2464 ), .ZN(_u10_u3_n3295 ) );
NAND2_X1 _u10_u3_U1181  ( .A1(_u10_u3_n3295 ), .A2(_u10_u3_n2835 ), .ZN(_u10_u3_n2623 ) );
INV_X1 _u10_u3_U1180  ( .A(_u10_u3_n2623 ), .ZN(_u10_u3_n3185 ) );
INV_X1 _u10_u3_U1179  ( .A(_u10_u3_n2688 ), .ZN(_u10_u3_n2169 ) );
NAND2_X1 _u10_u3_U1178  ( .A1(_u10_u3_n3185 ), .A2(_u10_u3_n2169 ), .ZN(_u10_u3_n3286 ) );
NAND2_X1 _u10_u3_U1177  ( .A1(_u10_u3_n2833 ), .A2(_u10_u3_n3278 ), .ZN(_u10_u3_n3298 ) );
NAND3_X1 _u10_u3_U1176  ( .A1(_u10_u3_n3297 ), .A2(_u10_u3_n2838 ), .A3(_u10_u3_n3298 ), .ZN(_u10_u3_n3296 ) );
NAND2_X1 _u10_u3_U1175  ( .A1(_u10_u3_n2830 ), .A2(_u10_u3_n3296 ), .ZN(_u10_u3_n3287 ) );
NAND2_X1 _u10_u3_U1174  ( .A1(_u10_u3_n3295 ), .A2(_u10_u3_n3001 ), .ZN(_u10_u3_n3292 ) );
NAND2_X1 _u10_u3_U1173  ( .A1(_u10_u3_n3294 ), .A2(_u10_u3_n2089 ), .ZN(_u10_u3_n3293 ) );
AND2_X1 _u10_u3_U1172  ( .A1(_u10_u3_n3292 ), .A2(_u10_u3_n3293 ), .ZN(_u10_u3_n2548 ) );
NAND2_X1 _u10_u3_U1171  ( .A1(_u10_u3_n2548 ), .A2(_u10_u3_n2091 ), .ZN(_u10_u3_n2304 ) );
NAND2_X1 _u10_u3_U1170  ( .A1(_u10_u3_n2304 ), .A2(_u10_u3_n2446 ), .ZN(_u10_u3_n3290 ) );
NAND2_X1 _u10_u3_U1169  ( .A1(_u10_u3_n2549 ), .A2(_u10_u3_n2446 ), .ZN(_u10_u3_n2790 ) );
NOR2_X1 _u10_u3_U1168  ( .A1(_u10_u3_n1936 ), .A2(_u10_u3_n2790 ), .ZN(_u10_u3_n2789 ) );
INV_X1 _u10_u3_U1167  ( .A(_u10_u3_n2789 ), .ZN(_u10_u3_n3291 ) );
OR2_X1 _u10_u3_U1166  ( .A1(_u10_u3_n2828 ), .A2(_u10_u3_n2790 ), .ZN(_u10_u3_n2498 ) );
NAND4_X1 _u10_u3_U1165  ( .A1(_u10_u3_n3290 ), .A2(_u10_u3_n3291 ), .A3(_u10_u3_n2498 ), .A4(_u10_u3_n2001 ), .ZN(_u10_u3_n3289 ) );
NAND2_X1 _u10_u3_U1164  ( .A1(_u10_u3_n2445 ), .A2(_u10_u3_n3289 ), .ZN(_u10_u3_n3288 ) );
NAND3_X1 _u10_u3_U1163  ( .A1(_u10_u3_n3286 ), .A2(_u10_u3_n3287 ), .A3(_u10_u3_n3288 ), .ZN(_u10_u3_n3280 ) );
NOR2_X1 _u10_u3_U1162  ( .A1(_u10_u3_n2940 ), .A2(_u10_u3_n1913 ), .ZN(_u10_u3_n3281 ) );
INV_X1 _u10_u3_U1161  ( .A(1'b0), .ZN(_u10_u3_n1864 ) );
NAND2_X1 _u10_u3_U1160  ( .A1(1'b0), .A2(_u10_u3_n2588 ), .ZN(_u10_u3_n2141 ) );
INV_X1 _u10_u3_U1159  ( .A(_u10_u3_n2141 ), .ZN(_u10_u3_n3159 ) );
NAND3_X1 _u10_u3_U1158  ( .A1(_u10_u3_n2103 ), .A2(_u10_u3_n1864 ), .A3(_u10_u3_n3159 ), .ZN(_u10_u3_n2520 ) );
INV_X1 _u10_u3_U1157  ( .A(_u10_u3_n2520 ), .ZN(_u10_u3_n2630 ) );
INV_X1 _u10_u3_U1156  ( .A(_u10_u3_n2307 ), .ZN(_u10_u3_n2382 ) );
NOR4_X1 _u10_u3_U1155  ( .A1(_u10_u3_n2382 ), .A2(_u10_u3_n2722 ), .A3(_u10_u3_n1925 ), .A4(_u10_u3_n2508 ), .ZN(_u10_u3_n3260 ) );
NOR2_X1 _u10_u3_U1154  ( .A1(_u10_u3_n2498 ), .A2(_u10_u3_n2911 ), .ZN(_u10_u3_n2633 ) );
NOR2_X1 _u10_u3_U1153  ( .A1(_u10_u3_n2633 ), .A2(_u10_u3_n3278 ), .ZN(_u10_u3_n3285 ) );
INV_X1 _u10_u3_U1152  ( .A(_u10_u3_n1866 ), .ZN(_u10_u3_n1926 ) );
NOR2_X1 _u10_u3_U1151  ( .A1(_u10_u3_n3285 ), .A2(_u10_u3_n1926 ), .ZN(_u10_u3_n3284 ) );
NOR4_X1 _u10_u3_U1150  ( .A1(1'b0), .A2(_u10_u3_n2630 ), .A3(_u10_u3_n3260 ),.A4(_u10_u3_n3284 ), .ZN(_u10_u3_n3283 ) );
NOR2_X1 _u10_u3_U1149  ( .A1(_u10_u3_n3283 ), .A2(_u10_u3_n2980 ), .ZN(_u10_u3_n3282 ) );
NOR4_X1 _u10_u3_U1148  ( .A1(_u10_u3_n3279 ), .A2(_u10_u3_n3280 ), .A3(_u10_u3_n3281 ), .A4(_u10_u3_n3282 ), .ZN(_u10_u3_n3241 ) );
NAND2_X1 _u10_u3_U1147  ( .A1(_u10_u3_n1836 ), .A2(_u10_u3_n2291 ), .ZN(_u10_u3_n2147 ) );
NAND2_X1 _u10_u3_U1146  ( .A1(_u10_u3_n2443 ), .A2(_u10_u3_n2147 ), .ZN(_u10_u3_n3261 ) );
INV_X1 _u10_u3_U1145  ( .A(_u10_u3_n1841 ), .ZN(_u10_u3_n2571 ) );
NAND2_X1 _u10_u3_U1144  ( .A1(_u10_u3_n2571 ), .A2(_u10_u3_n3278 ), .ZN(_u10_u3_n3277 ) );
NAND2_X1 _u10_u3_U1143  ( .A1(_u10_u3_n3276 ), .A2(_u10_u3_n3277 ), .ZN(_u10_u3_n2819 ) );
OR2_X1 _u10_u3_U1142  ( .A1(_u10_u3_n2819 ), .A2(_u10_u3_n3275 ), .ZN(_u10_u3_n3273 ) );
NAND2_X1 _u10_u3_U1141  ( .A1(_u10_u3_n2815 ), .A2(_u10_u3_n2080 ), .ZN(_u10_u3_n3274 ) );
NAND2_X1 _u10_u3_U1140  ( .A1(_u10_u3_n2014 ), .A2(_u10_u3_n3274 ), .ZN(_u10_u3_n2165 ) );
NAND2_X1 _u10_u3_U1139  ( .A1(_u10_u3_n3273 ), .A2(_u10_u3_n2165 ), .ZN(_u10_u3_n3262 ) );
NAND2_X1 _u10_u3_U1138  ( .A1(_u10_u3_n2688 ), .A2(_u10_u3_n2126 ), .ZN(_u10_u3_n1956 ) );
INV_X1 _u10_u3_U1137  ( .A(_u10_u3_n1956 ), .ZN(_u10_u3_n1860 ) );
NOR2_X1 _u10_u3_U1136  ( .A1(1'b0), .A2(_u10_u3_n2498 ), .ZN(_u10_u3_n3271 ));
NOR2_X1 _u10_u3_U1135  ( .A1(_u10_u3_n3271 ), .A2(_u10_u3_n3272 ), .ZN(_u10_u3_n3270 ) );
NOR2_X1 _u10_u3_U1134  ( .A1(_u10_u3_n1860 ), .A2(_u10_u3_n3270 ), .ZN(_u10_u3_n3264 ) );
INV_X1 _u10_u3_U1133  ( .A(_u10_u3_n2632 ), .ZN(_u10_u3_n3202 ) );
NAND2_X1 _u10_u3_U1132  ( .A1(_u10_u3_n3236 ), .A2(_u10_u3_n3269 ), .ZN(_u10_u3_n3036 ) );
INV_X1 _u10_u3_U1131  ( .A(_u10_u3_n3036 ), .ZN(_u10_u3_n1960 ) );
NAND2_X1 _u10_u3_U1130  ( .A1(_u10_u3_n3202 ), .A2(_u10_u3_n1960 ), .ZN(_u10_u3_n3079 ) );
NOR3_X1 _u10_u3_U1129  ( .A1(_u10_u3_n3079 ), .A2(1'b0), .A3(_u10_u3_n3268 ),.ZN(_u10_u3_n3265 ) );
INV_X1 _u10_u3_U1128  ( .A(_u10_u3_n2014 ), .ZN(_u10_u3_n2709 ) );
NAND2_X1 _u10_u3_U1127  ( .A1(_u10_u3_n2709 ), .A2(_u10_u3_n2166 ), .ZN(_u10_u3_n2145 ) );
INV_X1 _u10_u3_U1126  ( .A(_u10_u3_n2145 ), .ZN(_u10_u3_n3258 ) );
NOR2_X1 _u10_u3_U1125  ( .A1(_u10_u3_n3258 ), .A2(_u10_u3_n2183 ), .ZN(_u10_u3_n3267 ) );
NOR2_X1 _u10_u3_U1124  ( .A1(_u10_u3_n3267 ), .A2(_u10_u3_n2567 ), .ZN(_u10_u3_n3266 ) );
NOR3_X1 _u10_u3_U1123  ( .A1(_u10_u3_n3264 ), .A2(_u10_u3_n3265 ), .A3(_u10_u3_n3266 ), .ZN(_u10_u3_n3263 ) );
NAND3_X1 _u10_u3_U1122  ( .A1(_u10_u3_n3261 ), .A2(_u10_u3_n3262 ), .A3(_u10_u3_n3263 ), .ZN(_u10_u3_n3243 ) );
INV_X1 _u10_u3_U1121  ( .A(_u10_u3_n2102 ), .ZN(_u10_u3_n2509 ) );
NAND2_X1 _u10_u3_U1120  ( .A1(_u10_u3_n3260 ), .A2(_u10_u3_n2509 ), .ZN(_u10_u3_n3247 ) );
INV_X1 _u10_u3_U1119  ( .A(_u10_u3_n3259 ), .ZN(_u10_u3_n2015 ) );
NAND2_X1 _u10_u3_U1118  ( .A1(_u10_u3_n2015 ), .A2(_u10_u3_n3258 ), .ZN(_u10_u3_n3248 ) );
NAND2_X1 _u10_u3_U1117  ( .A1(_u10_u3_n2251 ), .A2(_u10_u3_n2169 ), .ZN(_u10_u3_n3255 ) );
OR2_X1 _u10_u3_U1116  ( .A1(_u10_u3_n3157 ), .A2(_u10_u3_n2256 ), .ZN(_u10_u3_n3257 ) );
NAND2_X1 _u10_u3_U1115  ( .A1(_u10_u3_n2105 ), .A2(_u10_u3_n3257 ), .ZN(_u10_u3_n3256 ) );
AND2_X1 _u10_u3_U1114  ( .A1(_u10_u3_n3255 ), .A2(_u10_u3_n3256 ), .ZN(_u10_u3_n3212 ) );
INV_X1 _u10_u3_U1113  ( .A(_u10_u3_n2037 ), .ZN(_u10_u3_n2987 ) );
NAND2_X1 _u10_u3_U1112  ( .A1(_u10_u3_n2987 ), .A2(_u10_u3_n2038 ), .ZN(_u10_u3_n2212 ) );
NOR2_X1 _u10_u3_U1111  ( .A1(_u10_u3_n2212 ), .A2(1'b0), .ZN(_u10_u3_n2658 ));
INV_X1 _u10_u3_U1110  ( .A(_u10_u3_n2658 ), .ZN(_u10_u3_n2343 ) );
NAND2_X1 _u10_u3_U1109  ( .A1(_u10_u3_n2344 ), .A2(_u10_u3_n3254 ), .ZN(_u10_u3_n1928 ) );
NAND2_X1 _u10_u3_U1108  ( .A1(_u10_u3_n2588 ), .A2(_u10_u3_n1928 ), .ZN(_u10_u3_n3253 ) );
NAND2_X1 _u10_u3_U1107  ( .A1(_u10_u3_n2343 ), .A2(_u10_u3_n3253 ), .ZN(_u10_u3_n3252 ) );
NAND2_X1 _u10_u3_U1106  ( .A1(_u10_u3_n2105 ), .A2(_u10_u3_n3252 ), .ZN(_u10_u3_n3251 ) );
NAND2_X1 _u10_u3_U1105  ( .A1(_u10_u3_n3212 ), .A2(_u10_u3_n3251 ), .ZN(_u10_u3_n3250 ) );
NAND2_X1 _u10_u3_U1104  ( .A1(_u10_u3_n2307 ), .A2(_u10_u3_n3250 ), .ZN(_u10_u3_n3249 ) );
NAND3_X1 _u10_u3_U1103  ( .A1(_u10_u3_n3247 ), .A2(_u10_u3_n3248 ), .A3(_u10_u3_n3249 ), .ZN(_u10_u3_n3244 ) );
AND2_X1 _u10_u3_U1102  ( .A1(_u10_u3_n2915 ), .A2(_u10_u3_n2059 ), .ZN(_u10_u3_n2957 ) );
AND3_X1 _u10_u3_U1101  ( .A1(_u10_u3_n3223 ), .A2(_u10_u3_n2837 ), .A3(_u10_u3_n2957 ), .ZN(_u10_u3_n2051 ) );
NOR2_X1 _u10_u3_U1100  ( .A1(_u10_u3_n2528 ), .A2(_u10_u3_n2051 ), .ZN(_u10_u3_n2605 ) );
NOR2_X1 _u10_u3_U1099  ( .A1(_u10_u3_n2605 ), .A2(_u10_u3_n2346 ), .ZN(_u10_u3_n3245 ) );
NOR2_X1 _u10_u3_U1098  ( .A1(_u10_u3_n2291 ), .A2(_u10_u3_n2062 ), .ZN(_u10_u3_n3246 ) );
NOR4_X1 _u10_u3_U1097  ( .A1(_u10_u3_n3243 ), .A2(_u10_u3_n3244 ), .A3(_u10_u3_n3245 ), .A4(_u10_u3_n3246 ), .ZN(_u10_u3_n3242 ) );
NAND2_X1 _u10_u3_U1096  ( .A1(_u10_u3_n3241 ), .A2(_u10_u3_n3242 ), .ZN(_u10_u3_n2311 ) );
OR3_X1 _u10_u3_U1095  ( .A1(_u10_u3_n1987 ), .A2(_u10_u3_n3240 ), .A3(_u10_u3_n2311 ), .ZN(_u10_u3_n3192 ) );
INV_X1 _u10_u3_U1094  ( .A(_u10_u3_n2886 ), .ZN(_u10_u3_n2720 ) );
NOR2_X1 _u10_u3_U1093  ( .A1(_u10_u3_n2004 ), .A2(_u10_u3_n2720 ), .ZN(_u10_u3_n2455 ) );
INV_X1 _u10_u3_U1092  ( .A(_u10_u3_n2488 ), .ZN(_u10_u3_n2938 ) );
AND3_X1 _u10_u3_U1091  ( .A1(_u10_u3_n2455 ), .A2(_u10_u3_n1859 ), .A3(_u10_u3_n2938 ), .ZN(_u10_u3_n3239 ) );
INV_X1 _u10_u3_U1090  ( .A(_u10_u3_n2633 ), .ZN(_u10_u3_n2937 ) );
NOR2_X1 _u10_u3_U1089  ( .A1(_u10_u3_n3239 ), .A2(_u10_u3_n2937 ), .ZN(_u10_u3_n3227 ) );
NOR2_X1 _u10_u3_U1088  ( .A1(_u10_u3_n1976 ), .A2(_u10_u3_n1969 ), .ZN(_u10_u3_n3237 ) );
NOR2_X1 _u10_u3_U1087  ( .A1(1'b0), .A2(_u10_u3_n2947 ), .ZN(_u10_u3_n3238 ));
NOR3_X1 _u10_u3_U1086  ( .A1(_u10_u3_n2476 ), .A2(_u10_u3_n3237 ), .A3(_u10_u3_n3238 ), .ZN(_u10_u3_n3235 ) );
NOR3_X1 _u10_u3_U1085  ( .A1(_u10_u3_n1813 ), .A2(_u10_u3_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_10 ), .ZN(_u10_u3_n3135 ) );
NAND2_X1 _u10_u3_U1084  ( .A1(_u10_u3_n3135 ), .A2(_u10_u3_n3236 ), .ZN(_u10_u3_n2573 ) );
NOR2_X1 _u10_u3_U1083  ( .A1(_u10_u3_n3235 ), .A2(_u10_u3_n2573 ), .ZN(_u10_u3_n3228 ) );
NOR2_X1 _u10_u3_U1082  ( .A1(_u10_u3_n2216 ), .A2(_u10_u3_n1868 ), .ZN(_u10_u3_n3233 ) );
INV_X1 _u10_u3_U1081  ( .A(_u10_u3_n2550 ), .ZN(_u10_u3_n2475 ) );
NOR3_X1 _u10_u3_U1080  ( .A1(_u10_u3_n2475 ), .A2(1'b0), .A3(_u10_u3_n1925 ),.ZN(_u10_u3_n3234 ) );
NOR3_X1 _u10_u3_U1079  ( .A1(_u10_u3_n3233 ), .A2(1'b0), .A3(_u10_u3_n3234 ),.ZN(_u10_u3_n3232 ) );
NOR2_X1 _u10_u3_U1078  ( .A1(_u10_u3_n3232 ), .A2(_u10_u3_n2037 ), .ZN(_u10_u3_n3229 ) );
NOR2_X1 _u10_u3_U1077  ( .A1(_u10_u3_n3231 ), .A2(_u10_u3_n2365 ), .ZN(_u10_u3_n3230 ) );
NOR4_X1 _u10_u3_U1076  ( .A1(_u10_u3_n3227 ), .A2(_u10_u3_n3228 ), .A3(_u10_u3_n3229 ), .A4(_u10_u3_n3230 ), .ZN(_u10_u3_n3205 ) );
NOR3_X1 _u10_u3_U1075  ( .A1(_u10_u3_n3226 ), .A2(_u10_u3_n2687 ), .A3(_u10_u3_n2145 ), .ZN(_u10_u3_n3217 ) );
NOR3_X1 _u10_u3_U1074  ( .A1(_u10_u3_n3225 ), .A2(1'b0), .A3(_u10_u3_n2587 ),.ZN(_u10_u3_n3218 ) );
NOR2_X1 _u10_u3_U1073  ( .A1(_u10_u3_n3159 ), .A2(1'b0), .ZN(_u10_u3_n3224 ));
NOR2_X1 _u10_u3_U1072  ( .A1(_u10_u3_n3224 ), .A2(_u10_u3_n2584 ), .ZN(_u10_u3_n3219 ) );
NAND2_X1 _u10_u3_U1071  ( .A1(_u10_u3_n3222 ), .A2(_u10_u3_n3223 ), .ZN(_u10_u3_n2048 ) );
INV_X1 _u10_u3_U1070  ( .A(_u10_u3_n2048 ), .ZN(_u10_u3_n2859 ) );
NOR2_X1 _u10_u3_U1069  ( .A1(_u10_u3_n2859 ), .A2(_u10_u3_n2054 ), .ZN(_u10_u3_n3221 ) );
NOR2_X1 _u10_u3_U1068  ( .A1(_u10_u3_n3221 ), .A2(_u10_u3_n2346 ), .ZN(_u10_u3_n3220 ) );
NOR4_X1 _u10_u3_U1067  ( .A1(_u10_u3_n3217 ), .A2(_u10_u3_n3218 ), .A3(_u10_u3_n3219 ), .A4(_u10_u3_n3220 ), .ZN(_u10_u3_n3206 ) );
NAND2_X1 _u10_u3_U1066  ( .A1(_u10_u3_n2377 ), .A2(_u10_u3_n2721 ), .ZN(_u10_u3_n3213 ) );
AND4_X1 _u10_u3_U1065  ( .A1(1'b0), .A2(_u10_u3_n2502 ), .A3(_u10_u3_n2972 ),.A4(_u10_u3_n3040 ), .ZN(_u10_u3_n2406 ) );
NAND2_X1 _u10_u3_U1064  ( .A1(_u10_u3_n2406 ), .A2(_u10_u3_n2979 ), .ZN(_u10_u3_n3214 ) );
NAND2_X1 _u10_u3_U1063  ( .A1(_u10_u3_n2630 ), .A2(_u10_u3_n3216 ), .ZN(_u10_u3_n2376 ) );
INV_X1 _u10_u3_U1062  ( .A(_u10_u3_n2376 ), .ZN(_u10_u3_n3108 ) );
NAND2_X1 _u10_u3_U1061  ( .A1(_u10_u3_n3108 ), .A2(_u10_u3_n2507 ), .ZN(_u10_u3_n3215 ) );
NOR2_X1 _u10_u3_U1060  ( .A1(_u10_u3_n2937 ), .A2(1'b0), .ZN(_u10_u3_n2649 ));
INV_X1 _u10_u3_U1059  ( .A(_u10_u3_n2253 ), .ZN(_u10_u3_n2971 ) );
NAND2_X1 _u10_u3_U1058  ( .A1(_u10_u3_n2649 ), .A2(_u10_u3_n2971 ), .ZN(_u10_u3_n2918 ) );
NAND4_X1 _u10_u3_U1057  ( .A1(_u10_u3_n3213 ), .A2(_u10_u3_n3214 ), .A3(_u10_u3_n3215 ), .A4(_u10_u3_n2918 ), .ZN(_u10_u3_n3208 ) );
NOR2_X1 _u10_u3_U1056  ( .A1(_u10_u3_n2000 ), .A2(_u10_u3_n2902 ), .ZN(_u10_u3_n3209 ) );
NOR2_X1 _u10_u3_U1055  ( .A1(_u10_u3_n3212 ), .A2(_u10_u3_n2475 ), .ZN(_u10_u3_n3210 ) );
INV_X1 _u10_u3_U1054  ( .A(_u10_u3_n2441 ), .ZN(_u10_u3_n3128 ) );
NOR2_X1 _u10_u3_U1053  ( .A1(_u10_u3_n2356 ), .A2(_u10_u3_n3128 ), .ZN(_u10_u3_n3211 ) );
NOR4_X1 _u10_u3_U1052  ( .A1(_u10_u3_n3208 ), .A2(_u10_u3_n3209 ), .A3(_u10_u3_n3210 ), .A4(_u10_u3_n3211 ), .ZN(_u10_u3_n3207 ) );
NAND3_X1 _u10_u3_U1051  ( .A1(_u10_u3_n3205 ), .A2(_u10_u3_n3206 ), .A3(_u10_u3_n3207 ), .ZN(_u10_u3_n2611 ) );
NOR2_X1 _u10_u3_U1050  ( .A1(_u10_u3_n2212 ), .A2(_u10_u3_n2216 ), .ZN(_u10_u3_n1937 ) );
NOR2_X1 _u10_u3_U1049  ( .A1(_u10_u3_n2533 ), .A2(_u10_u3_n2214 ), .ZN(_u10_u3_n2765 ) );
INV_X1 _u10_u3_U1048  ( .A(_u10_u3_n2005 ), .ZN(_u10_u3_n2111 ) );
AND2_X1 _u10_u3_U1047  ( .A1(_u10_u3_n2765 ), .A2(_u10_u3_n2111 ), .ZN(_u10_u3_n3201 ) );
INV_X1 _u10_u3_U1046  ( .A(_u10_u3_n3059 ), .ZN(_u10_u3_n3076 ) );
NAND2_X1 _u10_u3_U1045  ( .A1(_u10_u3_n3201 ), .A2(_u10_u3_n3076 ), .ZN(_u10_u3_n3204 ) );
NAND2_X1 _u10_u3_U1044  ( .A1(_u10_u3_n1937 ), .A2(_u10_u3_n3204 ), .ZN(_u10_u3_n3193 ) );
NAND2_X1 _u10_u3_U1043  ( .A1(_u10_u3_n2254 ), .A2(_u10_u3_n2212 ), .ZN(_u10_u3_n3203 ) );
NAND3_X1 _u10_u3_U1042  ( .A1(_u10_u3_n3203 ), .A2(_u10_u3_n2175 ), .A3(_u10_u3_n2649 ), .ZN(_u10_u3_n3194 ) );
NOR2_X1 _u10_u3_U1041  ( .A1(_u10_u3_n2985 ), .A2(1'b0), .ZN(_u10_u3_n1959 ));
NAND2_X1 _u10_u3_U1040  ( .A1(_u10_u3_n1959 ), .A2(_u10_u3_n3202 ), .ZN(_u10_u3_n2202 ) );
NAND4_X1 _u10_u3_U1039  ( .A1(_u10_u3_n3079 ), .A2(_u10_u3_n2621 ), .A3(_u10_u3_n2202 ), .A4(_u10_u3_n2798 ), .ZN(_u10_u3_n3200 ) );
NAND2_X1 _u10_u3_U1038  ( .A1(_u10_u3_n3201 ), .A2(_u10_u3_n2937 ), .ZN(_u10_u3_n2772 ) );
NAND2_X1 _u10_u3_U1037  ( .A1(_u10_u3_n3200 ), .A2(_u10_u3_n2772 ), .ZN(_u10_u3_n3195 ) );
NAND2_X1 _u10_u3_U1036  ( .A1(_u10_u3_n2765 ), .A2(_u10_u3_n1869 ), .ZN(_u10_u3_n3199 ) );
NAND2_X1 _u10_u3_U1035  ( .A1(_u10_u3_n2049 ), .A2(_u10_u3_n3199 ), .ZN(_u10_u3_n3057 ) );
NOR2_X1 _u10_u3_U1034  ( .A1(_u10_u3_n2495 ), .A2(_u10_u3_n3057 ), .ZN(_u10_u3_n3197 ) );
NOR2_X1 _u10_u3_U1033  ( .A1(_u10_u3_n2883 ), .A2(_u10_u3_n2485 ), .ZN(_u10_u3_n3198 ) );
NOR2_X1 _u10_u3_U1032  ( .A1(_u10_u3_n3197 ), .A2(_u10_u3_n3198 ), .ZN(_u10_u3_n3196 ) );
NAND4_X1 _u10_u3_U1031  ( .A1(_u10_u3_n3193 ), .A2(_u10_u3_n3194 ), .A3(_u10_u3_n3195 ), .A4(_u10_u3_n3196 ), .ZN(_u10_u3_n2887 ) );
NOR4_X1 _u10_u3_U1030  ( .A1(_u10_u3_n3191 ), .A2(_u10_u3_n3192 ), .A3(_u10_u3_n2611 ), .A4(_u10_u3_n2887 ), .ZN(_u10_u3_n3015 ) );
NAND3_X1 _u10_u3_U1029  ( .A1(_u10_u3_n3190 ), .A2(_u10_u3_n2049 ), .A3(_u10_u3_n2957 ), .ZN(_u10_u3_n2699 ) );
OR2_X1 _u10_u3_U1028  ( .A1(_u10_u3_n2699 ), .A2(_u10_u3_n1813 ), .ZN(_u10_u3_n3187 ) );
NAND3_X1 _u10_u3_U1027  ( .A1(_u10_u3_n2978 ), .A2(_u10_u3_n2405 ), .A3(1'b0), .ZN(_u10_u3_n3188 ) );
NAND4_X1 _u10_u3_U1026  ( .A1(_u10_u3_n3058 ), .A2(_u10_u3_n3187 ), .A3(_u10_u3_n3188 ), .A4(_u10_u3_n3189 ), .ZN(_u10_u3_n3186 ) );
NAND2_X1 _u10_u3_U1025  ( .A1(_u10_u3_n2063 ), .A2(_u10_u3_n3186 ), .ZN(_u10_u3_n3163 ) );
NAND2_X1 _u10_u3_U1024  ( .A1(_u10_u3_n3185 ), .A2(_u10_u3_n2329 ), .ZN(_u10_u3_n3164 ) );
NAND2_X1 _u10_u3_U1023  ( .A1(_u10_u3_n2689 ), .A2(_u10_u3_n2365 ), .ZN(_u10_u3_n2736 ) );
NOR2_X1 _u10_u3_U1022  ( .A1(_u10_u3_n2736 ), .A2(_u10_u3_n2488 ), .ZN(_u10_u3_n1855 ) );
INV_X1 _u10_u3_U1021  ( .A(_u10_u3_n1855 ), .ZN(_u10_u3_n3184 ) );
NOR2_X1 _u10_u3_U1020  ( .A1(_u10_u3_n2274 ), .A2(_u10_u3_n2359 ), .ZN(_u10_u3_n2952 ) );
NOR2_X1 _u10_u3_U1019  ( .A1(_u10_u3_n3184 ), .A2(_u10_u3_n2952 ), .ZN(_u10_u3_n2776 ) );
OR2_X1 _u10_u3_U1018  ( .A1(_u10_u3_n2852 ), .A2(_u10_u3_n2776 ), .ZN(_u10_u3_n3165 ) );
NAND2_X1 _u10_u3_U1017  ( .A1(_u10_u3_n3126 ), .A2(_u10_u3_n2915 ), .ZN(_u10_u3_n3065 ) );
NOR3_X1 _u10_u3_U1016  ( .A1(_u10_u3_n3065 ), .A2(1'b0), .A3(_u10_u3_n2632 ),.ZN(_u10_u3_n3182 ) );
NOR3_X1 _u10_u3_U1015  ( .A1(_u10_u3_n3182 ), .A2(_u10_u3_n3183 ), .A3(_u10_u3_n3108 ), .ZN(_u10_u3_n3181 ) );
NOR2_X1 _u10_u3_U1014  ( .A1(_u10_u3_n3181 ), .A2(_u10_u3_n3162 ), .ZN(_u10_u3_n3167 ) );
INV_X1 _u10_u3_U1013  ( .A(_u10_u3_n3180 ), .ZN(_u10_u3_n3140 ) );
NAND3_X1 _u10_u3_U1012  ( .A1(_u10_u3_n3140 ), .A2(_u10_u3_n2163 ), .A3(_u10_u3_n2092 ), .ZN(_u10_u3_n3175 ) );
NOR4_X1 _u10_u3_U1011  ( .A1(_u10_u3_n2411 ), .A2(_u10_u3_n2710 ), .A3(_u10_u3_n3141 ), .A4(_u10_u3_n3089 ), .ZN(_u10_u3_n3179 ) );
NOR2_X1 _u10_u3_U1010  ( .A1(1'b0), .A2(_u10_u3_n3179 ), .ZN(_u10_u3_n3177 ));
NOR2_X1 _u10_u3_U1009  ( .A1(_u10_u3_n1898 ), .A2(_u10_u3_n1847 ), .ZN(_u10_u3_n3178 ) );
NOR4_X1 _u10_u3_U1008  ( .A1(_u10_u3_n3175 ), .A2(_u10_u3_n3176 ), .A3(_u10_u3_n3177 ), .A4(_u10_u3_n3178 ), .ZN(_u10_u3_n3173 ) );
NAND2_X1 _u10_u3_U1007  ( .A1(_u10_u3_n3135 ), .A2(_u10_u3_n3174 ), .ZN(_u10_u3_n2159 ) );
NOR2_X1 _u10_u3_U1006  ( .A1(_u10_u3_n3173 ), .A2(_u10_u3_n2159 ), .ZN(_u10_u3_n3168 ) );
OR3_X1 _u10_u3_U1005  ( .A1(_u10_u3_n3172 ), .A2(1'b0), .A3(_u10_u3_n3126 ),.ZN(_u10_u3_n3171 ) );
NAND2_X1 _u10_u3_U1004  ( .A1(_u10_u3_n2600 ), .A2(_u10_u3_n3171 ), .ZN(_u10_u3_n3153 ) );
AND3_X1 _u10_u3_U1003  ( .A1(_u10_u3_n3153 ), .A2(_u10_u3_n2947 ), .A3(_u10_u3_n2579 ), .ZN(_u10_u3_n3170 ) );
NOR2_X1 _u10_u3_U1002  ( .A1(_u10_u3_n3170 ), .A2(_u10_u3_n2359 ), .ZN(_u10_u3_n3169 ) );
NOR3_X1 _u10_u3_U1001  ( .A1(_u10_u3_n3167 ), .A2(_u10_u3_n3168 ), .A3(_u10_u3_n3169 ), .ZN(_u10_u3_n3166 ) );
NAND4_X1 _u10_u3_U1000  ( .A1(_u10_u3_n3163 ), .A2(_u10_u3_n3164 ), .A3(_u10_u3_n3165 ), .A4(_u10_u3_n3166 ), .ZN(_u10_u3_n3130 ) );
NAND2_X1 _u10_u3_U999  ( .A1(_u10_u3_n2375 ), .A2(_u10_u3_n3162 ), .ZN(_u10_u3_n1923 ) );
NAND2_X1 _u10_u3_U998  ( .A1(_u10_u3_n3062 ), .A2(_u10_u3_n1923 ), .ZN(_u10_u3_n3154 ) );
NAND2_X1 _u10_u3_U997  ( .A1(_u10_u3_n2103 ), .A2(_u10_u3_n2509 ), .ZN(_u10_u3_n3161 ) );
NAND2_X1 _u10_u3_U996  ( .A1(_u10_u3_n2344 ), .A2(_u10_u3_n3161 ), .ZN(_u10_u3_n3160 ) );
NAND2_X1 _u10_u3_U995  ( .A1(_u10_u3_n3159 ), .A2(_u10_u3_n3160 ), .ZN(_u10_u3_n2635 ) );
AND3_X1 _u10_u3_U994  ( .A1(_u10_u3_n2549 ), .A2(_u10_u3_n2108 ), .A3(_u10_u3_n3126 ), .ZN(_u10_u3_n3093 ) );
NAND2_X1 _u10_u3_U993  ( .A1(_u10_u3_n3093 ), .A2(_u10_u3_n2941 ), .ZN(_u10_u3_n3158 ) );
NAND3_X1 _u10_u3_U992  ( .A1(_u10_u3_n3076 ), .A2(_u10_u3_n3066 ), .A3(_u10_u3_n3158 ), .ZN(_u10_u3_n3156 ) );
NAND2_X1 _u10_u3_U991  ( .A1(_u10_u3_n3156 ), .A2(_u10_u3_n3157 ), .ZN(_u10_u3_n3155 ) );
NAND3_X1 _u10_u3_U990  ( .A1(_u10_u3_n3154 ), .A2(_u10_u3_n2635 ), .A3(_u10_u3_n3155 ), .ZN(_u10_u3_n3131 ) );
INV_X1 _u10_u3_U989  ( .A(_u10_u3_n2594 ), .ZN(_u10_u3_n2846 ) );
NAND3_X1 _u10_u3_U988  ( .A1(_u10_u3_n2162 ), .A2(_u10_u3_n2082 ), .A3(_u10_u3_n2105 ), .ZN(_u10_u3_n2077 ) );
NAND4_X1 _u10_u3_U987  ( .A1(_u10_u3_n3153 ), .A2(_u10_u3_n1969 ), .A3(_u10_u3_n2846 ), .A4(_u10_u3_n2077 ), .ZN(_u10_u3_n3148 ) );
NAND2_X1 _u10_u3_U986  ( .A1(_u10_u3_n2838 ), .A2(_u10_u3_n3128 ), .ZN(_u10_u3_n3152 ) );
NAND2_X1 _u10_u3_U985  ( .A1(_u10_u3_n3152 ), .A2(_u10_u3_n2600 ), .ZN(_u10_u3_n3151 ) );
NAND2_X1 _u10_u3_U984  ( .A1(_u10_u3_n2282 ), .A2(_u10_u3_n3151 ), .ZN(_u10_u3_n2601 ) );
NOR4_X1 _u10_u3_U983  ( .A1(_u10_u3_n2885 ), .A2(_u10_u3_n2534 ), .A3(_u10_u3_n2214 ), .A4(_u10_u3_n3059 ), .ZN(_u10_u3_n3150 ) );
NOR2_X1 _u10_u3_U982  ( .A1(_u10_u3_n3150 ), .A2(_u10_u3_n2853 ), .ZN(_u10_u3_n3149 ) );
NOR4_X1 _u10_u3_U981  ( .A1(_u10_u3_n3148 ), .A2(_u10_u3_n2601 ), .A3(_u10_u3_n3149 ), .A4(_u10_u3_n1975 ), .ZN(_u10_u3_n3146 ) );
NAND3_X1 _u10_u3_U980  ( .A1(_u10_SYNOPSYS_UNCONNECTED_13 ), .A2(_u10_SYNOPSYS_UNCONNECTED_9 ), .A3(_u10_u3_n3147 ), .ZN(_u10_u3_n2071 ) );
NOR2_X1 _u10_u3_U979  ( .A1(_u10_u3_n3146 ), .A2(_u10_u3_n2071 ), .ZN(_u10_u3_n3132 ) );
NOR2_X1 _u10_u3_U978  ( .A1(1'b0), .A2(_u10_u3_n1847 ), .ZN(_u10_u3_n3143 ));
INV_X1 _u10_u3_U977  ( .A(_u10_u3_n3145 ), .ZN(_u10_u3_n3144 ) );
NOR2_X1 _u10_u3_U976  ( .A1(_u10_u3_n3143 ), .A2(_u10_u3_n3144 ), .ZN(_u10_u3_n3142 ) );
NOR2_X1 _u10_u3_U975  ( .A1(1'b0), .A2(_u10_u3_n3142 ), .ZN(_u10_u3_n3137 ));
NAND2_X1 _u10_u3_U974  ( .A1(_u10_u3_n2549 ), .A2(_u10_u3_n3141 ), .ZN(_u10_u3_n3138 ) );
NAND2_X1 _u10_u3_U973  ( .A1(_u10_u3_n1896 ), .A2(_u10_u3_n3140 ), .ZN(_u10_u3_n2544 ) );
NAND2_X1 _u10_u3_U972  ( .A1(_u10_u3_n2089 ), .A2(_u10_u3_n2544 ), .ZN(_u10_u3_n3139 ) );
NAND2_X1 _u10_u3_U971  ( .A1(_u10_u3_n3138 ), .A2(_u10_u3_n3139 ), .ZN(_u10_u3_n2795 ) );
NOR4_X1 _u10_u3_U970  ( .A1(_u10_u3_n2300 ), .A2(_u10_u3_n3137 ), .A3(_u10_u3_n2304 ), .A4(_u10_u3_n2795 ), .ZN(_u10_u3_n3134 ) );
NAND2_X1 _u10_u3_U969  ( .A1(_u10_u3_n3135 ), .A2(_u10_u3_n3136 ), .ZN(_u10_u3_n2085 ) );
NOR2_X1 _u10_u3_U968  ( .A1(_u10_u3_n3134 ), .A2(_u10_u3_n2085 ), .ZN(_u10_u3_n3133 ) );
NOR4_X1 _u10_u3_U967  ( .A1(_u10_u3_n3130 ), .A2(_u10_u3_n3131 ), .A3(_u10_u3_n3132 ), .A4(_u10_u3_n3133 ), .ZN(_u10_u3_n3016 ) );
INV_X1 _u10_u3_U966  ( .A(_u10_u3_n2686 ), .ZN(_u10_u3_n2278 ) );
NAND4_X1 _u10_u3_U965  ( .A1(_u10_u3_n2105 ), .A2(_u10_u3_n2278 ), .A3(_u10_u3_n3129 ), .A4(_u10_u3_n2600 ), .ZN(_u10_u3_n2437 ) );
NAND2_X1 _u10_u3_U964  ( .A1(_u10_u3_n3128 ), .A2(_u10_u3_n2437 ), .ZN(_u10_u3_n3127 ) );
NAND2_X1 _u10_u3_U963  ( .A1(_u10_u3_n2815 ), .A2(_u10_u3_n3127 ), .ZN(_u10_u3_n3098 ) );
INV_X1 _u10_u3_U962  ( .A(_u10_u3_n2573 ), .ZN(_u10_u3_n1967 ) );
NAND2_X1 _u10_u3_U961  ( .A1(_u10_u3_n3126 ), .A2(_u10_u3_n2078 ), .ZN(_u10_u3_n3123 ) );
NAND2_X1 _u10_u3_U960  ( .A1(_u10_u3_n3076 ), .A2(_u10_u3_n1925 ), .ZN(_u10_u3_n3125 ) );
NAND2_X1 _u10_u3_U959  ( .A1(_u10_u3_n2669 ), .A2(_u10_u3_n3125 ), .ZN(_u10_u3_n3124 ) );
NAND4_X1 _u10_u3_U958  ( .A1(_u10_u3_n3122 ), .A2(_u10_u3_n3123 ), .A3(_u10_u3_n3124 ), .A4(_u10_u3_n2579 ), .ZN(_u10_u3_n3121 ) );
NAND2_X1 _u10_u3_U957  ( .A1(_u10_u3_n3121 ), .A2(_u10_u3_n2874 ), .ZN(_u10_u3_n3120 ) );
NAND2_X1 _u10_u3_U956  ( .A1(_u10_u3_n2382 ), .A2(_u10_u3_n3120 ), .ZN(_u10_u3_n3119 ) );
NAND2_X1 _u10_u3_U955  ( .A1(_u10_u3_n1967 ), .A2(_u10_u3_n3119 ), .ZN(_u10_u3_n3099 ) );
NAND2_X1 _u10_u3_U954  ( .A1(_u10_u3_n3118 ), .A2(_u10_u3_n3001 ), .ZN(_u10_u3_n3117 ) );
NAND2_X1 _u10_u3_U953  ( .A1(_u10_u3_n2446 ), .A2(_u10_u3_n3117 ), .ZN(_u10_u3_n3116 ) );
NAND2_X1 _u10_u3_U952  ( .A1(_u10_u3_n2445 ), .A2(_u10_u3_n3116 ), .ZN(_u10_u3_n3100 ) );
OR2_X1 _u10_u3_U951  ( .A1(_u10_u3_n3115 ), .A2(_u10_u3_n2687 ), .ZN(_u10_u3_n3114 ) );
AND3_X1 _u10_u3_U950  ( .A1(_u10_u3_n2061 ), .A2(_u10_u3_n2166 ), .A3(_u10_u3_n3114 ), .ZN(_u10_u3_n3045 ) );
NOR2_X1 _u10_u3_U949  ( .A1(1'b0), .A2(_u10_u3_n3045 ), .ZN(_u10_u3_n3113 ));
NOR2_X1 _u10_u3_U948  ( .A1(_u10_u3_n3113 ), .A2(1'b0), .ZN(_u10_u3_n3112 ));
NOR2_X1 _u10_u3_U947  ( .A1(_u10_u3_n3112 ), .A2(_u10_u3_n2356 ), .ZN(_u10_u3_n3102 ) );
NAND2_X1 _u10_u3_U946  ( .A1(_u10_u3_n2571 ), .A2(_u10_u3_n2165 ), .ZN(_u10_u3_n3078 ) );
NAND2_X1 _u10_u3_U945  ( .A1(_u10_u3_n2365 ), .A2(_u10_u3_n3078 ), .ZN(_u10_u3_n2241 ) );
NOR2_X1 _u10_u3_U944  ( .A1(_u10_u3_n2377 ), .A2(_u10_u3_n2241 ), .ZN(_u10_u3_n3111 ) );
NOR2_X1 _u10_u3_U943  ( .A1(_u10_u3_n3111 ), .A2(_u10_u3_n1869 ), .ZN(_u10_u3_n3103 ) );
NOR2_X1 _u10_u3_U942  ( .A1(_u10_u3_n2999 ), .A2(_u10_u3_n2977 ), .ZN(_u10_u3_n3061 ) );
NOR2_X1 _u10_u3_U941  ( .A1(_u10_u3_n3061 ), .A2(_u10_u3_n2367 ), .ZN(_u10_u3_n3106 ) );
NAND2_X1 _u10_u3_U940  ( .A1(_u10_u3_n2977 ), .A2(_u10_u3_n3000 ), .ZN(_u10_u3_n3110 ) );
NAND2_X1 _u10_u3_U939  ( .A1(_u10_u3_n3109 ), .A2(_u10_u3_n3110 ), .ZN(_u10_u3_n1924 ) );
AND2_X1 _u10_u3_U938  ( .A1(_u10_u3_n1924 ), .A2(_u10_u3_n3108 ), .ZN(_u10_u3_n3107 ) );
NOR2_X1 _u10_u3_U937  ( .A1(_u10_u3_n3106 ), .A2(_u10_u3_n3107 ), .ZN(_u10_u3_n3105 ) );
NOR2_X1 _u10_u3_U936  ( .A1(_u10_u3_n3105 ), .A2(_u10_u3_n2008 ), .ZN(_u10_u3_n3104 ) );
NOR3_X1 _u10_u3_U935  ( .A1(_u10_u3_n3102 ), .A2(_u10_u3_n3103 ), .A3(_u10_u3_n3104 ), .ZN(_u10_u3_n3101 ) );
NAND4_X1 _u10_u3_U934  ( .A1(_u10_u3_n3098 ), .A2(_u10_u3_n3099 ), .A3(_u10_u3_n3100 ), .A4(_u10_u3_n3101 ), .ZN(_u10_u3_n3071 ) );
NOR2_X1 _u10_u3_U933  ( .A1(_u10_u3_n1926 ), .A2(_u10_u3_n2980 ), .ZN(_u10_u3_n2218 ) );
INV_X1 _u10_u3_U932  ( .A(_u10_u3_n2721 ), .ZN(_u10_u3_n2910 ) );
NAND2_X1 _u10_u3_U931  ( .A1(_u10_u3_n2910 ), .A2(_u10_u3_n1869 ), .ZN(_u10_u3_n2779 ) );
NAND2_X1 _u10_u3_U930  ( .A1(_u10_u3_n2218 ), .A2(_u10_u3_n2779 ), .ZN(_u10_u3_n3081 ) );
NAND2_X1 _u10_u3_U929  ( .A1(_u10_u3_n1922 ), .A2(_u10_u3_n1864 ), .ZN(_u10_u3_n2179 ) );
NOR3_X1 _u10_u3_U928  ( .A1(_u10_u3_n1961 ), .A2(_u10_u3_n1918 ), .A3(_u10_u3_n2179 ), .ZN(_u10_u3_n2693 ) );
NAND2_X1 _u10_u3_U927  ( .A1(_u10_u3_n3097 ), .A2(_u10_u3_n1924 ), .ZN(_u10_u3_n3096 ) );
NAND2_X1 _u10_u3_U926  ( .A1(_u10_u3_n1984 ), .A2(_u10_u3_n3096 ), .ZN(_u10_u3_n2506 ) );
INV_X1 _u10_u3_U925  ( .A(_u10_u3_n2506 ), .ZN(_u10_u3_n2366 ) );
NAND2_X1 _u10_u3_U924  ( .A1(_u10_u3_n2366 ), .A2(_u10_u3_n2375 ), .ZN(_u10_u3_n2236 ) );
NAND2_X1 _u10_u3_U923  ( .A1(_u10_u3_n2693 ), .A2(_u10_u3_n2236 ), .ZN(_u10_u3_n3082 ) );
NAND2_X1 _u10_u3_U922  ( .A1(1'b0), .A2(_u10_u3_n2126 ), .ZN(_u10_u3_n3095 ));
NAND2_X1 _u10_u3_U921  ( .A1(_u10_u3_n1956 ), .A2(_u10_u3_n3095 ), .ZN(_u10_u3_n2907 ) );
OR2_X1 _u10_u3_U920  ( .A1(_u10_u3_n2902 ), .A2(_u10_u3_n2907 ), .ZN(_u10_u3_n3085 ) );
NAND2_X1 _u10_u3_U919  ( .A1(_u10_u3_n2256 ), .A2(_u10_u3_n2113 ), .ZN(_u10_u3_n3094 ) );
NAND2_X1 _u10_u3_U918  ( .A1(_u10_u3_n2688 ), .A2(_u10_u3_n3094 ), .ZN(_u10_u3_n3092 ) );
NAND2_X1 _u10_u3_U917  ( .A1(_u10_u3_n3093 ), .A2(_u10_u3_n3092 ), .ZN(_u10_u3_n3086 ) );
INV_X1 _u10_u3_U916  ( .A(_u10_u3_n2159 ), .ZN(_u10_u3_n1894 ) );
NAND2_X1 _u10_u3_U915  ( .A1(_u10_u3_n3067 ), .A2(_u10_u3_n1894 ), .ZN(_u10_u3_n3091 ) );
INV_X1 _u10_u3_U914  ( .A(_u10_u3_n3092 ), .ZN(_u10_u3_n2234 ) );
NAND3_X1 _u10_u3_U913  ( .A1(_u10_u3_n3091 ), .A2(_u10_u3_n2126 ), .A3(_u10_u3_n2234 ), .ZN(_u10_u3_n3090 ) );
NAND2_X1 _u10_u3_U912  ( .A1(1'b0), .A2(_u10_u3_n3090 ), .ZN(_u10_u3_n3087 ));
NAND3_X1 _u10_u3_U911  ( .A1(_u10_u3_n2329 ), .A2(_u10_u3_n3089 ), .A3(_u10_u3_n2549 ), .ZN(_u10_u3_n3088 ) );
NAND4_X1 _u10_u3_U910  ( .A1(_u10_u3_n3085 ), .A2(_u10_u3_n3086 ), .A3(_u10_u3_n3087 ), .A4(_u10_u3_n3088 ), .ZN(_u10_u3_n3084 ) );
NAND2_X1 _u10_u3_U909  ( .A1(_u10_u3_n3084 ), .A2(_u10_u3_n2803 ), .ZN(_u10_u3_n3083 ) );
NAND3_X1 _u10_u3_U908  ( .A1(_u10_u3_n3081 ), .A2(_u10_u3_n3082 ), .A3(_u10_u3_n3083 ), .ZN(_u10_u3_n3072 ) );
INV_X1 _u10_u3_U907  ( .A(_u10_u3_n2689 ), .ZN(_u10_u3_n1955 ) );
NOR3_X1 _u10_u3_U906  ( .A1(_u10_u3_n1955 ), .A2(_u10_u3_n2813 ), .A3(_u10_u3_n2488 ), .ZN(_u10_u3_n3080 ) );
NOR2_X1 _u10_u3_U905  ( .A1(_u10_u3_n3080 ), .A2(_u10_u3_n2485 ), .ZN(_u10_u3_n3073 ) );
NAND3_X1 _u10_u3_U904  ( .A1(_u10_u3_n2621 ), .A2(_u10_u3_n2202 ), .A3(_u10_u3_n3079 ), .ZN(_u10_u3_n2110 ) );
NOR2_X1 _u10_u3_U903  ( .A1(_u10_u3_n2110 ), .A2(_u10_u3_n2218 ), .ZN(_u10_u3_n2775 ) );
INV_X1 _u10_u3_U902  ( .A(_u10_u3_n2775 ), .ZN(_u10_u3_n3024 ) );
INV_X1 _u10_u3_U901  ( .A(_u10_u3_n3078 ), .ZN(_u10_u3_n2133 ) );
INV_X1 _u10_u3_U900  ( .A(_u10_u3_n2007 ), .ZN(_u10_u3_n2358 ) );
NAND2_X1 _u10_u3_U899  ( .A1(_u10_u3_n2358 ), .A2(_u10_u3_n2886 ), .ZN(_u10_u3_n2240 ) );
INV_X1 _u10_u3_U898  ( .A(_u10_u3_n2240 ), .ZN(_u10_u3_n2083 ) );
NOR3_X1 _u10_u3_U897  ( .A1(_u10_u3_n2952 ), .A2(_u10_u3_n2004 ), .A3(_u10_u3_n1891 ), .ZN(_u10_u3_n3077 ) );
NAND3_X1 _u10_u3_U896  ( .A1(_u10_u3_n2083 ), .A2(_u10_u3_n2938 ), .A3(_u10_u3_n3077 ), .ZN(_u10_u3_n1886 ) );
NOR3_X1 _u10_u3_U895  ( .A1(_u10_u3_n3024 ), .A2(_u10_u3_n2133 ), .A3(_u10_u3_n1886 ), .ZN(_u10_u3_n3075 ) );
NOR2_X1 _u10_u3_U894  ( .A1(_u10_u3_n3075 ), .A2(_u10_u3_n3076 ), .ZN(_u10_u3_n3074 ) );
NOR4_X1 _u10_u3_U893  ( .A1(_u10_u3_n3071 ), .A2(_u10_u3_n3072 ), .A3(_u10_u3_n3073 ), .A4(_u10_u3_n3074 ), .ZN(_u10_u3_n3017 ) );
INV_X1 _u10_u3_U892  ( .A(_u10_u3_n3065 ), .ZN(_u10_u3_n3043 ) );
NAND2_X1 _u10_u3_U891  ( .A1(_u10_u3_n3043 ), .A2(_u10_u3_n2106 ), .ZN(_u10_u3_n3070 ) );
NAND2_X1 _u10_u3_U890  ( .A1(_u10_u3_n3070 ), .A2(_u10_u3_n2038 ), .ZN(_u10_u3_n3068 ) );
NAND2_X1 _u10_u3_U889  ( .A1(_u10_u3_n2344 ), .A2(_u10_u3_n2584 ), .ZN(_u10_u3_n3069 ) );
NAND3_X1 _u10_u3_U888  ( .A1(_u10_u3_n3068 ), .A2(_u10_u3_n1930 ), .A3(_u10_u3_n3069 ), .ZN(_u10_u3_n3047 ) );
NAND2_X1 _u10_u3_U887  ( .A1(_u10_u3_n2835 ), .A2(_u10_u3_n2466 ), .ZN(_u10_u3_n2130 ) );
INV_X1 _u10_u3_U886  ( .A(_u10_u3_n2130 ), .ZN(_u10_u3_n2168 ) );
NAND3_X1 _u10_u3_U885  ( .A1(_u10_u3_n3067 ), .A2(_u10_u3_n2329 ), .A3(_u10_u3_n2168 ), .ZN(_u10_u3_n2665 ) );
NAND3_X1 _u10_u3_U884  ( .A1(_u10_u3_n3065 ), .A2(_u10_u3_n3066 ), .A3(_u10_u3_n2342 ), .ZN(_u10_u3_n3064 ) );
NAND3_X1 _u10_u3_U883  ( .A1(_u10_u3_n3064 ), .A2(_u10_u3_n2175 ), .A3(_u10_u3_n2987 ), .ZN(_u10_u3_n3048 ) );
NOR3_X1 _u10_u3_U882  ( .A1(_u10_u3_n1849 ), .A2(1'b0), .A3(_u10_u3_n3063 ),.ZN(_u10_u3_n3050 ) );
NOR3_X1 _u10_u3_U881  ( .A1(_u10_u3_n2406 ), .A2(1'b0), .A3(_u10_u3_n3062 ),.ZN(_u10_u3_n3060 ) );
NOR3_X1 _u10_u3_U880  ( .A1(_u10_u3_n3060 ), .A2(1'b0), .A3(_u10_u3_n3061 ),.ZN(_u10_u3_n3051 ) );
NAND2_X1 _u10_u3_U879  ( .A1(_u10_u3_n3059 ), .A2(_u10_u3_n2049 ), .ZN(_u10_u3_n3056 ) );
NAND3_X1 _u10_u3_U878  ( .A1(_u10_u3_n3056 ), .A2(_u10_u3_n3057 ), .A3(_u10_u3_n3058 ), .ZN(_u10_u3_n3054 ) );
NOR4_X1 _u10_u3_U877  ( .A1(_u10_u3_n3054 ), .A2(_u10_u3_n3055 ), .A3(_u10_u3_n2055 ), .A4(_u10_u3_n2056 ), .ZN(_u10_u3_n3053 ) );
NOR3_X1 _u10_u3_U876  ( .A1(_u10_u3_n2346 ), .A2(1'b0), .A3(_u10_u3_n3053 ),.ZN(_u10_u3_n3052 ) );
NOR3_X1 _u10_u3_U875  ( .A1(_u10_u3_n3050 ), .A2(_u10_u3_n3051 ), .A3(_u10_u3_n3052 ), .ZN(_u10_u3_n3049 ) );
NAND4_X1 _u10_u3_U874  ( .A1(_u10_u3_n3047 ), .A2(_u10_u3_n2665 ), .A3(_u10_u3_n3048 ), .A4(_u10_u3_n3049 ), .ZN(_u10_u3_n3019 ) );
NAND2_X1 _u10_u3_U873  ( .A1(_u10_u3_n2056 ), .A2(_u10_u3_n2019 ), .ZN(_u10_u3_n3046 ) );
NAND2_X1 _u10_u3_U872  ( .A1(_u10_u3_n3045 ), .A2(_u10_u3_n3046 ), .ZN(_u10_u3_n3044 ) );
NAND2_X1 _u10_u3_U871  ( .A1(_u10_u3_n3044 ), .A2(_u10_u3_n2165 ), .ZN(_u10_u3_n3028 ) );
OR2_X1 _u10_u3_U870  ( .A1(_u10_u3_n2179 ), .A2(_u10_u3_n1961 ), .ZN(_u10_u3_n3037 ) );
NAND2_X1 _u10_u3_U869  ( .A1(_u10_u3_n3043 ), .A2(_u10_u3_n2336 ), .ZN(_u10_u3_n3042 ) );
NAND2_X1 _u10_u3_U868  ( .A1(_u10_u3_n3042 ), .A2(_u10_u3_n3006 ), .ZN(_u10_u3_n3041 ) );
NAND2_X1 _u10_u3_U867  ( .A1(_u10_u3_n3040 ), .A2(_u10_u3_n3041 ), .ZN(_u10_u3_n3026 ) );
NAND4_X1 _u10_u3_U866  ( .A1(_u10_u3_n3026 ), .A2(_u10_u3_n2520 ), .A3(_u10_u3_n1962 ), .A4(_u10_u3_n1864 ), .ZN(_u10_u3_n3039 ) );
NAND2_X1 _u10_u3_U865  ( .A1(_u10_u3_n3039 ), .A2(_u10_u3_n1922 ), .ZN(_u10_u3_n3038 ) );
NAND2_X1 _u10_u3_U864  ( .A1(_u10_u3_n3037 ), .A2(_u10_u3_n3038 ), .ZN(_u10_u3_n3035 ) );
NAND2_X1 _u10_u3_U863  ( .A1(_u10_u3_n2985 ), .A2(_u10_u3_n3036 ), .ZN(_u10_u3_n2432 ) );
NAND2_X1 _u10_u3_U862  ( .A1(_u10_u3_n3035 ), .A2(_u10_u3_n2432 ), .ZN(_u10_u3_n3029 ) );
INV_X1 _u10_u3_U861  ( .A(_u10_u3_n3034 ), .ZN(_u10_u3_n2777 ) );
INV_X1 _u10_u3_U860  ( .A(_u10_u3_n2772 ), .ZN(_u10_u3_n3032 ) );
NAND2_X1 _u10_u3_U859  ( .A1(_u10_u3_n1982 ), .A2(_u10_u3_n2978 ), .ZN(_u10_u3_n3033 ) );
NAND2_X1 _u10_u3_U858  ( .A1(_u10_u3_n3032 ), .A2(_u10_u3_n3033 ), .ZN(_u10_u3_n3031 ) );
NAND2_X1 _u10_u3_U857  ( .A1(_u10_u3_n2777 ), .A2(_u10_u3_n3031 ), .ZN(_u10_u3_n3030 ) );
NAND3_X1 _u10_u3_U856  ( .A1(_u10_u3_n3028 ), .A2(_u10_u3_n3029 ), .A3(_u10_u3_n3030 ), .ZN(_u10_u3_n3020 ) );
NOR3_X1 _u10_u3_U855  ( .A1(_u10_u3_n2179 ), .A2(1'b0), .A3(_u10_u3_n2375 ),.ZN(_u10_u3_n3027 ) );
NOR2_X1 _u10_u3_U854  ( .A1(_u10_u3_n3027 ), .A2(_u10_u3_n2177 ), .ZN(_u10_u3_n3025 ) );
NOR2_X1 _u10_u3_U853  ( .A1(_u10_u3_n3025 ), .A2(_u10_u3_n3026 ), .ZN(_u10_u3_n3021 ) );
NOR2_X1 _u10_u3_U852  ( .A1(_u10_u3_n2256 ), .A2(_u10_u3_n3024 ), .ZN(_u10_u3_n3023 ) );
NOR2_X1 _u10_u3_U851  ( .A1(_u10_u3_n3023 ), .A2(_u10_u3_n1868 ), .ZN(_u10_u3_n3022 ) );
NOR4_X1 _u10_u3_U850  ( .A1(_u10_u3_n3019 ), .A2(_u10_u3_n3020 ), .A3(_u10_u3_n3021 ), .A4(_u10_u3_n3022 ), .ZN(_u10_u3_n3018 ) );
NAND4_X1 _u10_u3_U849  ( .A1(_u10_u3_n3015 ), .A2(_u10_u3_n3016 ), .A3(_u10_u3_n3017 ), .A4(_u10_u3_n3018 ), .ZN(_u10_u3_n2958 ) );
NOR2_X1 _u10_u3_U848  ( .A1(1'b0), .A2(_u10_u3_n2573 ), .ZN(_u10_u3_n3011 ));
NOR2_X1 _u10_u3_U847  ( .A1(1'b0), .A2(_u10_u3_n2359 ), .ZN(_u10_u3_n3012 ));
NOR2_X1 _u10_u3_U846  ( .A1(1'b0), .A2(_u10_u3_n1859 ), .ZN(_u10_u3_n3013 ));
NOR2_X1 _u10_u3_U845  ( .A1(1'b0), .A2(_u10_u3_n1836 ), .ZN(_u10_u3_n3014 ));
NOR4_X1 _u10_u3_U844  ( .A1(_u10_u3_n3011 ), .A2(_u10_u3_n3012 ), .A3(_u10_u3_n3013 ), .A4(_u10_u3_n3014 ), .ZN(_u10_u3_n2959 ) );
NOR2_X1 _u10_u3_U843  ( .A1(1'b0), .A2(_u10_u3_n2025 ), .ZN(_u10_u3_n3007 ));
NOR2_X1 _u10_u3_U842  ( .A1(1'b0), .A2(_u10_u3_n2085 ), .ZN(_u10_u3_n3008 ));
NOR2_X1 _u10_u3_U841  ( .A1(1'b0), .A2(_u10_u3_n2607 ), .ZN(_u10_u3_n3009 ));
NOR2_X1 _u10_u3_U840  ( .A1(1'b0), .A2(_u10_u3_n2071 ), .ZN(_u10_u3_n3010 ));
NOR4_X1 _u10_u3_U839  ( .A1(_u10_u3_n3007 ), .A2(_u10_u3_n3008 ), .A3(_u10_u3_n3009 ), .A4(_u10_u3_n3010 ), .ZN(_u10_u3_n2960 ) );
NAND2_X1 _u10_u3_U838  ( .A1(_u10_u3_n1894 ), .A2(_u10_u3_n2466 ), .ZN(_u10_u3_n3002 ) );
NAND2_X1 _u10_u3_U837  ( .A1(_u10_u3_n2830 ), .A2(_u10_u3_n2600 ), .ZN(_u10_u3_n3003 ) );
NAND2_X1 _u10_u3_U836  ( .A1(_u10_u3_n1960 ), .A2(_u10_u3_n2431 ), .ZN(_u10_u3_n3004 ) );
NAND2_X1 _u10_u3_U835  ( .A1(_u10_u3_n2002 ), .A2(_u10_u3_n3006 ), .ZN(_u10_u3_n3005 ) );
NAND4_X1 _u10_u3_U834  ( .A1(_u10_u3_n3002 ), .A2(_u10_u3_n3003 ), .A3(_u10_u3_n3004 ), .A4(_u10_u3_n3005 ), .ZN(_u10_u3_n2992 ) );
NAND2_X1 _u10_u3_U833  ( .A1(_u10_u3_n2461 ), .A2(_u10_u3_n3001 ), .ZN(_u10_u3_n2997 ) );
NAND2_X1 _u10_u3_U832  ( .A1(_u10_u3_n2999 ), .A2(_u10_u3_n3000 ), .ZN(_u10_u3_n2998 ) );
NAND2_X1 _u10_u3_U831  ( .A1(_u10_u3_n2997 ), .A2(_u10_u3_n2998 ), .ZN(_u10_u3_n2993 ) );
NOR2_X1 _u10_u3_U830  ( .A1(_u10_SYNOPSYS_UNCONNECTED_9 ), .A2(_u10_u3_n2996 ), .ZN(_u10_u3_n2995 ) );
NOR2_X1 _u10_u3_U829  ( .A1(_u10_u3_n2995 ), .A2(_u10_u3_n2126 ), .ZN(_u10_u3_n2994 ) );
NOR4_X1 _u10_u3_U828  ( .A1(_u10_u3_n2992 ), .A2(_u10_u3_n2993 ), .A3(next_ch), .A4(_u10_u3_n2994 ), .ZN(_u10_u3_n2961 ) );
NAND2_X1 _u10_u3_U827  ( .A1(_u10_u3_n2445 ), .A2(_u10_u3_n2803 ), .ZN(_u10_u3_n2988 ) );
OR2_X1 _u10_u3_U826  ( .A1(_u10_u3_n2584 ), .A2(1'b0), .ZN(_u10_u3_n2989 ));
NAND2_X1 _u10_u3_U825  ( .A1(_u10_u3_n2709 ), .A2(_u10_u3_n2080 ), .ZN(_u10_u3_n2990 ) );
NAND2_X1 _u10_u3_U824  ( .A1(_u10_u3_n2183 ), .A2(_u10_u3_n2166 ), .ZN(_u10_u3_n2991 ) );
NAND4_X1 _u10_u3_U823  ( .A1(_u10_u3_n2988 ), .A2(_u10_u3_n2989 ), .A3(_u10_u3_n2990 ), .A4(_u10_u3_n2991 ), .ZN(_u10_u3_n2963 ) );
NAND2_X1 _u10_u3_U822  ( .A1(_u10_u3_n2987 ), .A2(_u10_u3_n1930 ), .ZN(_u10_u3_n2981 ) );
NAND2_X1 _u10_u3_U821  ( .A1(_u10_u3_n2986 ), .A2(_u10_u3_n2038 ), .ZN(_u10_u3_n2982 ) );
OR2_X1 _u10_u3_U820  ( .A1(_u10_u3_n2985 ), .A2(1'b0), .ZN(_u10_u3_n2983 ));
NAND2_X1 _u10_u3_U819  ( .A1(_u10_u3_n2169 ), .A2(_u10_u3_n2113 ), .ZN(_u10_u3_n2984 ) );
NAND4_X1 _u10_u3_U818  ( .A1(_u10_u3_n2981 ), .A2(_u10_u3_n2982 ), .A3(_u10_u3_n2983 ), .A4(_u10_u3_n2984 ), .ZN(_u10_u3_n2964 ) );
NAND2_X1 _u10_u3_U817  ( .A1(_u10_u3_n2509 ), .A2(_u10_u3_n1864 ), .ZN(_u10_u3_n2973 ) );
INV_X1 _u10_u3_U816  ( .A(_u10_u3_n2980 ), .ZN(_u10_u3_n1861 ) );
NAND2_X1 _u10_u3_U815  ( .A1(_u10_u3_n1861 ), .A2(_u10_u3_n1922 ), .ZN(_u10_u3_n2974 ) );
NAND2_X1 _u10_u3_U814  ( .A1(_u10_u3_n2979 ), .A2(_u10_u3_n2405 ), .ZN(_u10_u3_n2975 ) );
NAND2_X1 _u10_u3_U813  ( .A1(_u10_u3_n2977 ), .A2(_u10_u3_n2978 ), .ZN(_u10_u3_n2976 ) );
NAND4_X1 _u10_u3_U812  ( .A1(_u10_u3_n2973 ), .A2(_u10_u3_n2974 ), .A3(_u10_u3_n2975 ), .A4(_u10_u3_n2976 ), .ZN(_u10_u3_n2965 ) );
NAND2_X1 _u10_u3_U811  ( .A1(_u10_u3_n2507 ), .A2(_u10_u3_n2972 ), .ZN(_u10_u3_n2967 ) );
NAND2_X1 _u10_u3_U810  ( .A1(_u10_u3_n2043 ), .A2(_u10_u3_n1965 ), .ZN(_u10_u3_n2968 ) );
NAND2_X1 _u10_u3_U809  ( .A1(_u10_u3_n2063 ), .A2(_u10_u3_n1853 ), .ZN(_u10_u3_n2969 ) );
NAND2_X1 _u10_u3_U808  ( .A1(_u10_u3_n2971 ), .A2(_u10_u3_n2175 ), .ZN(_u10_u3_n2970 ) );
NAND4_X1 _u10_u3_U807  ( .A1(_u10_u3_n2967 ), .A2(_u10_u3_n2968 ), .A3(_u10_u3_n2969 ), .A4(_u10_u3_n2970 ), .ZN(_u10_u3_n2966 ) );
NOR4_X1 _u10_u3_U806  ( .A1(_u10_u3_n2963 ), .A2(_u10_u3_n2964 ), .A3(_u10_u3_n2965 ), .A4(_u10_u3_n2966 ), .ZN(_u10_u3_n2962 ) );
AND4_X1 _u10_u3_U805  ( .A1(_u10_u3_n2959 ), .A2(_u10_u3_n2960 ), .A3(_u10_u3_n2961 ), .A4(_u10_u3_n2962 ), .ZN(_u10_u3_n1819 ) );
MUX2_X1 _u10_u3_U804  ( .A(_u10_u3_n2958 ), .B(_u10_SYNOPSYS_UNCONNECTED_13 ), .S(_u10_u3_n1819 ), .Z(_u10_u3_n1808 ) );
NOR2_X1 _u10_u3_U803  ( .A1(_u10_u3_n2531 ), .A2(_u10_u3_n2607 ), .ZN(_u10_u3_n1911 ) );
NAND2_X1 _u10_u3_U802  ( .A1(_u10_u3_n1911 ), .A2(_u10_u3_n2957 ), .ZN(_u10_u3_n2954 ) );
NAND2_X1 _u10_u3_U801  ( .A1(_u10_u3_n1853 ), .A2(_u10_u3_n1965 ), .ZN(_u10_u3_n2956 ) );
NAND2_X1 _u10_u3_U800  ( .A1(_u10_u3_n1966 ), .A2(_u10_u3_n2956 ), .ZN(_u10_u3_n2955 ) );
NAND2_X1 _u10_u3_U799  ( .A1(_u10_u3_n2954 ), .A2(_u10_u3_n2955 ), .ZN(_u10_u3_n2670 ) );
NOR3_X1 _u10_u3_U798  ( .A1(_u10_u3_n1852 ), .A2(1'b0), .A3(_u10_u3_n1853 ),.ZN(_u10_u3_n2708 ) );
NAND2_X1 _u10_u3_U797  ( .A1(_u10_u3_n2708 ), .A2(_u10_u3_n2080 ), .ZN(_u10_u3_n2355 ) );
NOR2_X1 _u10_u3_U796  ( .A1(_u10_u3_n2355 ), .A2(1'b0), .ZN(_u10_u3_n2599 ));
NAND2_X1 _u10_u3_U795  ( .A1(_u10_u3_n2953 ), .A2(_u10_u3_n2599 ), .ZN(_u10_u3_n2423 ) );
OR2_X1 _u10_u3_U794  ( .A1(_u10_u3_n2423 ), .A2(_u10_u3_n2359 ), .ZN(_u10_u3_n2949 ) );
NAND3_X1 _u10_u3_U793  ( .A1(_u10_u3_n2105 ), .A2(_u10_u3_n1936 ), .A3(_u10_u3_n2952 ), .ZN(_u10_u3_n2950 ) );
NAND3_X1 _u10_u3_U792  ( .A1(_u10_u3_n2549 ), .A2(_u10_u3_n1936 ), .A3(1'b0),.ZN(_u10_u3_n2096 ) );
INV_X1 _u10_u3_U791  ( .A(_u10_u3_n2096 ), .ZN(_u10_u3_n2301 ) );
NAND2_X1 _u10_u3_U790  ( .A1(_u10_u3_n2301 ), .A2(_u10_u3_n2446 ), .ZN(_u10_u3_n2368 ) );
INV_X1 _u10_u3_U789  ( .A(_u10_u3_n2368 ), .ZN(_u10_u3_n2326 ) );
NAND2_X1 _u10_u3_U788  ( .A1(_u10_u3_n2326 ), .A2(_u10_u3_n2941 ), .ZN(_u10_u3_n2800 ) );
INV_X1 _u10_u3_U787  ( .A(_u10_u3_n2800 ), .ZN(_u10_u3_n2081 ) );
NAND2_X1 _u10_u3_U786  ( .A1(_u10_u3_n2081 ), .A2(_u10_u3_n2049 ), .ZN(_u10_u3_n2855 ) );
INV_X1 _u10_u3_U785  ( .A(_u10_u3_n2855 ), .ZN(_u10_u3_n2347 ) );
NAND2_X1 _u10_u3_U784  ( .A1(_u10_u3_n2347 ), .A2(_u10_u3_n2063 ), .ZN(_u10_u3_n2951 ) );
NAND3_X1 _u10_u3_U783  ( .A1(_u10_u3_n2949 ), .A2(_u10_u3_n2950 ), .A3(_u10_u3_n2951 ), .ZN(_u10_u3_n1997 ) );
INV_X1 _u10_u3_U782  ( .A(_u10_u3_n1997 ), .ZN(_u10_u3_n2917 ) );
AND2_X1 _u10_u3_U781  ( .A1(_u10_u3_n2709 ), .A2(_u10_u3_n2708 ), .ZN(_u10_u3_n2942 ) );
INV_X1 _u10_u3_U780  ( .A(_u10_u3_n2907 ), .ZN(_u10_u3_n2737 ) );
NAND2_X1 _u10_u3_U779  ( .A1(_u10_u3_n2737 ), .A2(_u10_u3_n2803 ), .ZN(_u10_u3_n1888 ) );
NOR2_X1 _u10_u3_U778  ( .A1(_u10_u3_n2001 ), .A2(_u10_u3_n1888 ), .ZN(_u10_u3_n2943 ) );
NAND4_X1 _u10_u3_U777  ( .A1(1'b0), .A2(_u10_u3_n2078 ), .A3(_u10_u3_n2059 ),.A4(_u10_u3_n2031 ), .ZN(_u10_u3_n2578 ) );
NOR3_X1 _u10_u3_U776  ( .A1(_u10_u3_n2719 ), .A2(_u10_u3_n2130 ), .A3(_u10_u3_n2305 ), .ZN(_u10_u3_n2386 ) );
NAND2_X1 _u10_u3_U775  ( .A1(_u10_u3_n2386 ), .A2(_u10_u3_n2669 ), .ZN(_u10_u3_n2948 ) );
NAND3_X1 _u10_u3_U774  ( .A1(_u10_u3_n2578 ), .A2(_u10_u3_n2947 ), .A3(_u10_u3_n2948 ), .ZN(_u10_u3_n2750 ) );
NOR2_X1 _u10_u3_U773  ( .A1(_u10_u3_n2274 ), .A2(_u10_u3_n2852 ), .ZN(_u10_u3_n2946 ) );
NOR3_X1 _u10_u3_U772  ( .A1(_u10_u3_n2750 ), .A2(1'b0), .A3(_u10_u3_n2946 ),.ZN(_u10_u3_n2945 ) );
NOR2_X1 _u10_u3_U771  ( .A1(_u10_u3_n2945 ), .A2(_u10_u3_n2359 ), .ZN(_u10_u3_n2944 ) );
NOR3_X1 _u10_u3_U770  ( .A1(_u10_u3_n2942 ), .A2(_u10_u3_n2943 ), .A3(_u10_u3_n2944 ), .ZN(_u10_u3_n2919 ) );
NOR2_X1 _u10_u3_U769  ( .A1(_u10_u3_n2423 ), .A2(1'b0), .ZN(_u10_u3_n1979 ));
NAND3_X1 _u10_u3_U768  ( .A1(_u10_u3_n2549 ), .A2(_u10_u3_n1936 ), .A3(_u10_u3_n1979 ), .ZN(_u10_u3_n2328 ) );
INV_X1 _u10_u3_U767  ( .A(_u10_u3_n2328 ), .ZN(_u10_u3_n2554 ) );
NAND3_X1 _u10_u3_U766  ( .A1(_u10_u3_n2941 ), .A2(_u10_u3_n2446 ), .A3(_u10_u3_n2554 ), .ZN(_u10_u3_n2115 ) );
NOR2_X1 _u10_u3_U765  ( .A1(_u10_u3_n2578 ), .A2(_u10_u3_n2030 ), .ZN(_u10_u3_n2553 ) );
INV_X1 _u10_u3_U764  ( .A(_u10_u3_n2553 ), .ZN(_u10_u3_n2269 ) );
NOR2_X1 _u10_u3_U763  ( .A1(_u10_u3_n2269 ), .A2(_u10_u3_n2790 ), .ZN(_u10_u3_n2657 ) );
INV_X1 _u10_u3_U762  ( .A(_u10_u3_n2657 ), .ZN(_u10_u3_n2210 ) );
NOR2_X1 _u10_u3_U761  ( .A1(_u10_u3_n2210 ), .A2(_u10_u3_n2911 ), .ZN(_u10_u3_n2213 ) );
INV_X1 _u10_u3_U760  ( .A(_u10_u3_n2213 ), .ZN(_u10_u3_n2456 ) );
NAND2_X1 _u10_u3_U759  ( .A1(_u10_u3_n2115 ), .A2(_u10_u3_n2456 ), .ZN(_u10_u3_n2634 ) );
INV_X1 _u10_u3_U758  ( .A(_u10_u3_n2634 ), .ZN(_u10_u3_n2220 ) );
NOR2_X1 _u10_u3_U757  ( .A1(_u10_u3_n2081 ), .A2(_u10_u3_n2386 ), .ZN(_u10_u3_n2131 ) );
NAND2_X1 _u10_u3_U756  ( .A1(_u10_u3_n2940 ), .A2(_u10_u3_n2131 ), .ZN(_u10_u3_n2138 ) );
INV_X1 _u10_u3_U755  ( .A(_u10_u3_n2138 ), .ZN(_u10_u3_n2927 ) );
NAND2_X1 _u10_u3_U754  ( .A1(_u10_u3_n2220 ), .A2(_u10_u3_n2927 ), .ZN(_u10_u3_n2939 ) );
NAND2_X1 _u10_u3_U753  ( .A1(_u10_u3_n1885 ), .A2(_u10_u3_n2939 ), .ZN(_u10_u3_n2931 ) );
NAND3_X1 _u10_u3_U752  ( .A1(_u10_u3_n1859 ), .A2(_u10_u3_n2365 ), .A3(_u10_u3_n2938 ), .ZN(_u10_u3_n2935 ) );
NAND3_X1 _u10_u3_U751  ( .A1(_u10_u3_n2927 ), .A2(_u10_u3_n2937 ), .A3(_u10_u3_n2220 ), .ZN(_u10_u3_n2936 ) );
NAND2_X1 _u10_u3_U750  ( .A1(_u10_u3_n2935 ), .A2(_u10_u3_n2936 ), .ZN(_u10_u3_n2932 ) );
INV_X1 _u10_u3_U749  ( .A(_u10_u3_n1937 ), .ZN(_u10_u3_n2350 ) );
NAND2_X1 _u10_u3_U748  ( .A1(_u10_u3_n1913 ), .A2(_u10_u3_n2350 ), .ZN(_u10_u3_n2934 ) );
NAND2_X1 _u10_u3_U747  ( .A1(_u10_u3_n2386 ), .A2(_u10_u3_n2934 ), .ZN(_u10_u3_n2933 ) );
NAND3_X1 _u10_u3_U746  ( .A1(_u10_u3_n2931 ), .A2(_u10_u3_n2932 ), .A3(_u10_u3_n2933 ), .ZN(_u10_u3_n2921 ) );
OR2_X1 _u10_u3_U745  ( .A1(_u10_u3_n2213 ), .A2(_u10_u3_n2386 ), .ZN(_u10_u3_n2930 ) );
NAND2_X1 _u10_u3_U744  ( .A1(_u10_u3_n2049 ), .A2(_u10_u3_n2930 ), .ZN(_u10_u3_n2228 ) );
AND2_X1 _u10_u3_U743  ( .A1(_u10_u3_n2228 ), .A2(_u10_u3_n2699 ), .ZN(_u10_u3_n2929 ) );
NOR2_X1 _u10_u3_U742  ( .A1(_u10_u3_n2929 ), .A2(_u10_u3_n2495 ), .ZN(_u10_u3_n2922 ) );
NOR2_X1 _u10_u3_U741  ( .A1(_u10_u3_n2633 ), .A2(_u10_u3_n2877 ), .ZN(_u10_u3_n2928 ) );
NOR2_X1 _u10_u3_U740  ( .A1(_u10_u3_n2928 ), .A2(_u10_u3_n2886 ), .ZN(_u10_u3_n2923 ) );
NOR2_X1 _u10_u3_U739  ( .A1(_u10_u3_n2927 ), .A2(_u10_u3_n2531 ), .ZN(_u10_u3_n2926 ) );
NOR2_X1 _u10_u3_U738  ( .A1(_u10_u3_n2926 ), .A2(_u10_u3_n2687 ), .ZN(_u10_u3_n2925 ) );
NOR2_X1 _u10_u3_U737  ( .A1(_u10_u3_n2925 ), .A2(_u10_u3_n1849 ), .ZN(_u10_u3_n2924 ) );
NOR4_X1 _u10_u3_U736  ( .A1(_u10_u3_n2921 ), .A2(_u10_u3_n2922 ), .A3(_u10_u3_n2923 ), .A4(_u10_u3_n2924 ), .ZN(_u10_u3_n2920 ) );
NAND4_X1 _u10_u3_U735  ( .A1(_u10_u3_n2917 ), .A2(_u10_u3_n2918 ), .A3(_u10_u3_n2919 ), .A4(_u10_u3_n2920 ), .ZN(_u10_u3_n2312 ) );
NOR2_X1 _u10_u3_U734  ( .A1(_u10_u3_n2600 ), .A2(_u10_u3_n2686 ), .ZN(_u10_u3_n2401 ) );
NAND2_X1 _u10_u3_U733  ( .A1(_u10_u3_n2401 ), .A2(_u10_u3_n2549 ), .ZN(_u10_u3_n2547 ) );
INV_X1 _u10_u3_U732  ( .A(_u10_u3_n2547 ), .ZN(_u10_u3_n2794 ) );
NAND3_X1 _u10_u3_U731  ( .A1(_u10_u3_n2364 ), .A2(_u10_u3_n2667 ), .A3(_u10_u3_n2794 ), .ZN(_u10_u3_n2535 ) );
INV_X1 _u10_u3_U730  ( .A(_u10_u3_n2535 ), .ZN(_u10_u3_n2586 ) );
NAND2_X1 _u10_u3_U729  ( .A1(_u10_u3_n2586 ), .A2(_u10_u3_n2571 ), .ZN(_u10_u3_n2916 ) );
NAND2_X1 _u10_u3_U728  ( .A1(_u10_u3_n2837 ), .A2(_u10_u3_n2916 ), .ZN(_u10_u3_n2436 ) );
NAND2_X1 _u10_u3_U727  ( .A1(_u10_u3_n2915 ), .A2(_u10_u3_n2571 ), .ZN(_u10_u3_n2914 ) );
NAND2_X1 _u10_u3_U726  ( .A1(_u10_u3_n2166 ), .A2(_u10_u3_n2914 ), .ZN(_u10_u3_n2017 ) );
NOR2_X1 _u10_u3_U725  ( .A1(_u10_u3_n2485 ), .A2(_u10_u3_n1841 ), .ZN(_u10_u3_n2913 ) );
OR4_X1 _u10_u3_U724  ( .A1(_u10_u3_n2436 ), .A2(_u10_u3_n2017 ), .A3(_u10_u3_n2913 ), .A4(_u10_u3_n2442 ), .ZN(_u10_u3_n2912 ) );
NAND2_X1 _u10_u3_U723  ( .A1(_u10_u3_n2709 ), .A2(_u10_u3_n2912 ), .ZN(_u10_u3_n2888 ) );
NAND3_X1 _u10_u3_U722  ( .A1(_u10_u3_n2078 ), .A2(_u10_u3_n2031 ), .A3(1'b0),.ZN(_u10_u3_n2580 ) );
INV_X1 _u10_u3_U721  ( .A(_u10_u3_n2580 ), .ZN(_u10_u3_n2680 ) );
AND2_X1 _u10_u3_U720  ( .A1(_u10_u3_n2680 ), .A2(_u10_u3_n2668 ), .ZN(_u10_u3_n1950 ) );
NAND2_X1 _u10_u3_U719  ( .A1(_u10_u3_n1950 ), .A2(_u10_u3_n2089 ), .ZN(_u10_u3_n2095 ) );
INV_X1 _u10_u3_U718  ( .A(_u10_u3_n2095 ), .ZN(_u10_u3_n2542 ) );
NAND2_X1 _u10_u3_U717  ( .A1(_u10_u3_n2542 ), .A2(_u10_u3_n2446 ), .ZN(_u10_u3_n1887 ) );
NOR2_X1 _u10_u3_U716  ( .A1(_u10_u3_n1887 ), .A2(_u10_u3_n2911 ), .ZN(_u10_u3_n2114 ) );
INV_X1 _u10_u3_U715  ( .A(_u10_u3_n2114 ), .ZN(_u10_u3_n1940 ) );
NAND3_X1 _u10_u3_U714  ( .A1(_u10_u3_n2535 ), .A2(_u10_u3_n1940 ), .A3(_u10_u3_n2910 ), .ZN(_u10_u3_n2524 ) );
NAND2_X1 _u10_u3_U713  ( .A1(_u10_u3_n2524 ), .A2(_u10_u3_n2488 ), .ZN(_u10_u3_n2889 ) );
NAND2_X1 _u10_u3_U712  ( .A1(_u10_u3_n2220 ), .A2(_u10_u3_n1940 ), .ZN(_u10_u3_n2763 ) );
NOR2_X1 _u10_u3_U711  ( .A1(_u10_u3_n2763 ), .A2(_u10_u3_n2586 ), .ZN(_u10_u3_n2808 ) );
NOR2_X1 _u10_u3_U710  ( .A1(_u10_u3_n2808 ), .A2(_u10_u3_n2350 ), .ZN(_u10_u3_n2908 ) );
NOR2_X1 _u10_u3_U709  ( .A1(_u10_u3_n2544 ), .A2(_u10_u3_n1950 ), .ZN(_u10_u3_n2899 ) );
NOR2_X1 _u10_u3_U708  ( .A1(_u10_u3_n2899 ), .A2(_u10_u3_n2159 ), .ZN(_u10_u3_n2909 ) );
NOR2_X1 _u10_u3_U707  ( .A1(_u10_u3_n2908 ), .A2(_u10_u3_n2909 ), .ZN(_u10_u3_n2890 ) );
NOR3_X1 _u10_u3_U706  ( .A1(_u10_u3_n2547 ), .A2(_u10_u3_n1846 ), .A3(_u10_u3_n2907 ), .ZN(_u10_u3_n2892 ) );
NOR3_X1 _u10_u3_U705  ( .A1(_u10_u3_n2240 ), .A2(_u10_u3_n2377 ), .A3(_u10_u3_n1911 ), .ZN(_u10_u3_n2906 ) );
NOR2_X1 _u10_u3_U704  ( .A1(_u10_u3_n2906 ), .A2(_u10_u3_n2535 ), .ZN(_u10_u3_n2893 ) );
NAND2_X1 _u10_u3_U703  ( .A1(_u10_u3_n2554 ), .A2(_u10_u3_n2446 ), .ZN(_u10_u3_n2903 ) );
AND3_X1 _u10_u3_U702  ( .A1(_u10_u3_n2210 ), .A2(_u10_u3_n2905 ), .A3(_u10_u3_n1887 ), .ZN(_u10_u3_n2904 ) );
NAND4_X1 _u10_u3_U701  ( .A1(_u10_u3_n2902 ), .A2(_u10_u3_n2498 ), .A3(_u10_u3_n2903 ), .A4(_u10_u3_n2904 ), .ZN(_u10_u3_n2788 ) );
INV_X1 _u10_u3_U700  ( .A(_u10_u3_n2788 ), .ZN(_u10_u3_n2901 ) );
NOR2_X1 _u10_u3_U699  ( .A1(_u10_u3_n2901 ), .A2(_u10_u3_n1888 ), .ZN(_u10_u3_n2894 ) );
NOR2_X1 _u10_u3_U698  ( .A1(_u10_u3_n2401 ), .A2(_u10_u3_n2553 ), .ZN(_u10_u3_n2900 ) );
NOR2_X1 _u10_u3_U697  ( .A1(_u10_u3_n2900 ), .A2(_u10_u3_n1954 ), .ZN(_u10_u3_n2897 ) );
NOR2_X1 _u10_u3_U696  ( .A1(1'b0), .A2(_u10_u3_n2899 ), .ZN(_u10_u3_n2898 ));
NOR2_X1 _u10_u3_U695  ( .A1(_u10_u3_n2897 ), .A2(_u10_u3_n2898 ), .ZN(_u10_u3_n2896 ) );
NOR2_X1 _u10_u3_U694  ( .A1(_u10_u3_n2896 ), .A2(_u10_u3_n1843 ), .ZN(_u10_u3_n2895 ) );
NOR4_X1 _u10_u3_U693  ( .A1(_u10_u3_n2892 ), .A2(_u10_u3_n2893 ), .A3(_u10_u3_n2894 ), .A4(_u10_u3_n2895 ), .ZN(_u10_u3_n2891 ) );
NAND4_X1 _u10_u3_U692  ( .A1(_u10_u3_n2888 ), .A2(_u10_u3_n2889 ), .A3(_u10_u3_n2890 ), .A4(_u10_u3_n2891 ), .ZN(_u10_u3_n2610 ) );
NOR4_X1 _u10_u3_U691  ( .A1(_u10_u3_n2670 ), .A2(_u10_u3_n2312 ), .A3(_u10_u3_n2610 ), .A4(_u10_u3_n2887 ), .ZN(_u10_u3_n2724 ) );
NOR2_X1 _u10_u3_U690  ( .A1(_u10_u3_n2883 ), .A2(_u10_u3_n2535 ), .ZN(_u10_u3_n2861 ) );
NOR2_X1 _u10_u3_U689  ( .A1(_u10_u3_n1855 ), .A2(_u10_u3_n1869 ), .ZN(_u10_u3_n2862 ) );
NOR2_X1 _u10_u3_U688  ( .A1(_u10_u3_n2886 ), .A2(_u10_u3_n2695 ), .ZN(_u10_u3_n2863 ) );
NAND2_X1 _u10_u3_U687  ( .A1(_u10_u3_n2813 ), .A2(_u10_u3_n2885 ), .ZN(_u10_u3_n2864 ) );
NAND2_X1 _u10_u3_U686  ( .A1(_u10_u3_n2114 ), .A2(_u10_u3_n2884 ), .ZN(_u10_u3_n2865 ) );
NAND2_X1 _u10_u3_U685  ( .A1(1'b0), .A2(_u10_u3_n2667 ), .ZN(_u10_u3_n2112 ));
NOR3_X1 _u10_u3_U684  ( .A1(_u10_u3_n2883 ), .A2(_u10_u3_n2112 ), .A3(_u10_u3_n2719 ), .ZN(_u10_u3_n2878 ) );
INV_X1 _u10_u3_U683  ( .A(_u10_u3_n2112 ), .ZN(_u10_u3_n1856 ) );
NAND2_X1 _u10_u3_U682  ( .A1(_u10_u3_n2364 ), .A2(_u10_u3_n1856 ), .ZN(_u10_u3_n2882 ) );
NAND2_X1 _u10_u3_U681  ( .A1(_u10_u3_n2882 ), .A2(_u10_u3_n1869 ), .ZN(_u10_u3_n2050 ) );
INV_X1 _u10_u3_U680  ( .A(_u10_u3_n2050 ), .ZN(_u10_u3_n1939 ) );
NOR2_X1 _u10_u3_U679  ( .A1(_u10_u3_n1939 ), .A2(_u10_u3_n1841 ), .ZN(_u10_u3_n2881 ) );
NOR2_X1 _u10_u3_U678  ( .A1(_u10_u3_n2881 ), .A2(_u10_u3_n2840 ), .ZN(_u10_u3_n2880 ) );
NOR2_X1 _u10_u3_U677  ( .A1(_u10_u3_n2880 ), .A2(_u10_u3_n1836 ), .ZN(_u10_u3_n2879 ) );
NOR2_X1 _u10_u3_U676  ( .A1(_u10_u3_n2878 ), .A2(_u10_u3_n2879 ), .ZN(_u10_u3_n2866 ) );
NOR2_X1 _u10_u3_U675  ( .A1(_u10_u3_n2081 ), .A2(_u10_u3_n2877 ), .ZN(_u10_u3_n1840 ) );
NAND2_X1 _u10_u3_U674  ( .A1(_u10_u3_n1840 ), .A2(_u10_u3_n2115 ), .ZN(_u10_u3_n1873 ) );
NAND2_X1 _u10_u3_U673  ( .A1(_u10_u3_n2695 ), .A2(_u10_u3_n1940 ), .ZN(_u10_u3_n1874 ) );
NOR3_X1 _u10_u3_U672  ( .A1(_u10_u3_n2050 ), .A2(_u10_u3_n1873 ), .A3(_u10_u3_n1874 ), .ZN(_u10_u3_n2876 ) );
NOR2_X1 _u10_u3_U671  ( .A1(_u10_u3_n2876 ), .A2(_u10_u3_n1913 ), .ZN(_u10_u3_n2868 ) );
NAND2_X1 _u10_u3_U670  ( .A1(_u10_u3_n2875 ), .A2(_u10_u3_n2466 ), .ZN(_u10_u3_n2872 ) );
INV_X1 _u10_u3_U669  ( .A(_u10_u3_n1979 ), .ZN(_u10_u3_n2746 ) );
NAND2_X1 _u10_u3_U668  ( .A1(_u10_u3_n2874 ), .A2(_u10_u3_n2746 ), .ZN(_u10_u3_n1935 ) );
NAND3_X1 _u10_u3_U667  ( .A1(_u10_u3_n1935 ), .A2(_u10_u3_n1936 ), .A3(_u10_u3_n2467 ), .ZN(_u10_u3_n2873 ) );
NAND2_X1 _u10_u3_U666  ( .A1(_u10_u3_n2872 ), .A2(_u10_u3_n2873 ), .ZN(_u10_u3_n2264 ) );
AND2_X1 _u10_u3_U665  ( .A1(_u10_u3_n2264 ), .A2(_u10_u3_n2461 ), .ZN(_u10_u3_n2869 ) );
AND2_X1 _u10_u3_U664  ( .A1(_u10_u3_n1966 ), .A2(_u10_u3_n2761 ), .ZN(_u10_u3_n2870 ) );
NOR2_X1 _u10_u3_U663  ( .A1(_u10_u3_n2159 ), .A2(_u10_u3_n2163 ), .ZN(_u10_u3_n2871 ) );
NOR4_X1 _u10_u3_U662  ( .A1(_u10_u3_n2868 ), .A2(_u10_u3_n2869 ), .A3(_u10_u3_n2870 ), .A4(_u10_u3_n2871 ), .ZN(_u10_u3_n2867 ) );
NAND4_X1 _u10_u3_U661  ( .A1(_u10_u3_n2864 ), .A2(_u10_u3_n2865 ), .A3(_u10_u3_n2866 ), .A4(_u10_u3_n2867 ), .ZN(_u10_u3_n1992 ) );
NOR4_X1 _u10_u3_U660  ( .A1(_u10_u3_n2861 ), .A2(_u10_u3_n2862 ), .A3(_u10_u3_n2863 ), .A4(_u10_u3_n1992 ), .ZN(_u10_u3_n2725 ) );
NAND2_X1 _u10_u3_U659  ( .A1(_u10_u3_n2364 ), .A2(_u10_u3_n1846 ), .ZN(_u10_u3_n2744 ) );
NAND4_X1 _u10_u3_U658  ( .A1(_u10_u3_n2765 ), .A2(_u10_u3_n1939 ), .A3(_u10_u3_n2744 ), .A4(_u10_u3_n2535 ), .ZN(_u10_u3_n2860 ) );
NAND2_X1 _u10_u3_U657  ( .A1(_u10_u3_n2049 ), .A2(_u10_u3_n2860 ), .ZN(_u10_u3_n2856 ) );
NOR4_X1 _u10_u3_U656  ( .A1(1'b0), .A2(_u10_u3_n2858 ), .A3(_u10_u3_n2859 ),.A4(_u10_u3_n2051 ), .ZN(_u10_u3_n2857 ) );
NAND4_X1 _u10_u3_U655  ( .A1(_u10_u3_n2228 ), .A2(_u10_u3_n2855 ), .A3(_u10_u3_n2856 ), .A4(_u10_u3_n2857 ), .ZN(_u10_u3_n2854 ) );
NAND2_X1 _u10_u3_U654  ( .A1(_u10_u3_n2043 ), .A2(_u10_u3_n2854 ), .ZN(_u10_u3_n2821 ) );
INV_X1 _u10_u3_U653  ( .A(_u10_u3_n2071 ), .ZN(_u10_u3_n2279 ) );
INV_X1 _u10_u3_U652  ( .A(_u10_u3_n2599 ), .ZN(_u10_u3_n2357 ) );
OR2_X1 _u10_u3_U651  ( .A1(_u10_u3_n2744 ), .A2(_u10_u3_n2853 ), .ZN(_u10_u3_n2844 ) );
NAND2_X1 _u10_u3_U650  ( .A1(_u10_u3_n2131 ), .A2(_u10_u3_n2852 ), .ZN(_u10_u3_n2851 ) );
NAND2_X1 _u10_u3_U649  ( .A1(_u10_u3_n2082 ), .A2(_u10_u3_n2851 ), .ZN(_u10_u3_n2848 ) );
NAND2_X1 _u10_u3_U648  ( .A1(_u10_u3_n2850 ), .A2(_u10_u3_n2600 ), .ZN(_u10_u3_n2849 ) );
NAND3_X1 _u10_u3_U647  ( .A1(_u10_u3_n2848 ), .A2(_u10_u3_n2077 ), .A3(_u10_u3_n2849 ), .ZN(_u10_u3_n2287 ) );
NAND2_X1 _u10_u3_U646  ( .A1(_u10_u3_n2082 ), .A2(_u10_u3_n2050 ), .ZN(_u10_u3_n2847 ) );
NAND2_X1 _u10_u3_U645  ( .A1(_u10_u3_n2846 ), .A2(_u10_u3_n2847 ), .ZN(_u10_u3_n2074 ) );
NOR3_X1 _u10_u3_U644  ( .A1(_u10_u3_n2287 ), .A2(_u10_u3_n2596 ), .A3(_u10_u3_n2074 ), .ZN(_u10_u3_n2845 ) );
NAND4_X1 _u10_u3_U643  ( .A1(_u10_u3_n2357 ), .A2(_u10_u3_n2837 ), .A3(_u10_u3_n2844 ), .A4(_u10_u3_n2845 ), .ZN(_u10_u3_n2843 ) );
NAND2_X1 _u10_u3_U642  ( .A1(_u10_u3_n2279 ), .A2(_u10_u3_n2843 ), .ZN(_u10_u3_n2822 ) );
NOR3_X1 _u10_u3_U641  ( .A1(_u10_u3_n1925 ), .A2(_u10_u3_n2842 ), .A3(_u10_u3_n2686 ), .ZN(_u10_u3_n2841 ) );
NOR3_X1 _u10_u3_U640  ( .A1(_u10_u3_n2840 ), .A2(_u10_u3_n2599 ), .A3(_u10_u3_n2841 ), .ZN(_u10_u3_n2839 ) );
AND4_X1 _u10_u3_U639  ( .A1(_u10_u3_n2836 ), .A2(_u10_u3_n2837 ), .A3(_u10_u3_n2838 ), .A4(_u10_u3_n2839 ), .ZN(_u10_u3_n2454 ) );
NOR2_X1 _u10_u3_U638  ( .A1(_u10_u3_n2719 ), .A2(_u10_u3_n2835 ), .ZN(_u10_u3_n2773 ) );
NOR2_X1 _u10_u3_U637  ( .A1(_u10_u3_n2138 ), .A2(_u10_u3_n2773 ), .ZN(_u10_u3_n2814 ) );
NAND2_X1 _u10_u3_U636  ( .A1(_u10_u3_n2814 ), .A2(_u10_u3_n1869 ), .ZN(_u10_u3_n2834 ) );
NAND2_X1 _u10_u3_U635  ( .A1(_u10_u3_n2833 ), .A2(_u10_u3_n2834 ), .ZN(_u10_u3_n2832 ) );
NAND2_X1 _u10_u3_U634  ( .A1(_u10_u3_n2454 ), .A2(_u10_u3_n2832 ), .ZN(_u10_u3_n2831 ) );
NAND2_X1 _u10_u3_U633  ( .A1(_u10_u3_n2830 ), .A2(_u10_u3_n2831 ), .ZN(_u10_u3_n2823 ) );
INV_X1 _u10_u3_U632  ( .A(_u10_u3_n2025 ), .ZN(_u10_u3_n2470 ) );
NAND2_X1 _u10_u3_U631  ( .A1(_u10_u3_n1979 ), .A2(_u10_u3_n1936 ), .ZN(_u10_u3_n2829 ) );
AND2_X1 _u10_u3_U630  ( .A1(_u10_u3_n2828 ), .A2(_u10_u3_n2829 ), .ZN(_u10_u3_n2469 ) );
NAND2_X1 _u10_u3_U629  ( .A1(_u10_u3_n2469 ), .A2(_u10_u3_n2269 ), .ZN(_u10_u3_n2161 ) );
INV_X1 _u10_u3_U628  ( .A(_u10_u3_n2161 ), .ZN(_u10_u3_n2276 ) );
NOR2_X1 _u10_u3_U627  ( .A1(_u10_u3_n2274 ), .A2(_u10_u3_n2719 ), .ZN(_u10_u3_n2827 ) );
NOR3_X1 _u10_u3_U626  ( .A1(_u10_u3_n2827 ), .A2(_u10_u3_n2742 ), .A3(_u10_u3_n2680 ), .ZN(_u10_u3_n2826 ) );
NAND3_X1 _u10_u3_U625  ( .A1(_u10_u3_n2276 ), .A2(_u10_u3_n2108 ), .A3(_u10_u3_n2826 ), .ZN(_u10_u3_n2825 ) );
NAND2_X1 _u10_u3_U624  ( .A1(_u10_u3_n2470 ), .A2(_u10_u3_n2825 ), .ZN(_u10_u3_n2824 ) );
NAND4_X1 _u10_u3_U623  ( .A1(_u10_u3_n2821 ), .A2(_u10_u3_n2822 ), .A3(_u10_u3_n2823 ), .A4(_u10_u3_n2824 ), .ZN(_u10_u3_n2804 ) );
NAND2_X1 _u10_u3_U622  ( .A1(_u10_u3_n2131 ), .A2(_u10_u3_n2744 ), .ZN(_u10_u3_n2820 ) );
NAND2_X1 _u10_u3_U621  ( .A1(_u10_u3_n2571 ), .A2(_u10_u3_n2820 ), .ZN(_u10_u3_n2817 ) );
NOR2_X1 _u10_u3_U620  ( .A1(_u10_u3_n2819 ), .A2(_u10_u3_n2436 ), .ZN(_u10_u3_n2818 ) );
NAND4_X1 _u10_u3_U619  ( .A1(_u10_u3_n2437 ), .A2(_u10_u3_n2355 ), .A3(_u10_u3_n2817 ), .A4(_u10_u3_n2818 ), .ZN(_u10_u3_n2816 ) );
NAND2_X1 _u10_u3_U618  ( .A1(_u10_u3_n2815 ), .A2(_u10_u3_n2816 ), .ZN(_u10_u3_n2809 ) );
INV_X1 _u10_u3_U617  ( .A(_u10_u3_n2814 ), .ZN(_u10_u3_n2812 ) );
OR2_X1 _u10_u3_U616  ( .A1(_u10_u3_n1911 ), .A2(_u10_u3_n2813 ), .ZN(_u10_u3_n1884 ) );
NAND2_X1 _u10_u3_U615  ( .A1(_u10_u3_n2812 ), .A2(_u10_u3_n1884 ), .ZN(_u10_u3_n2810 ) );
NOR2_X1 _u10_u3_U614  ( .A1(_u10_u3_n1894 ), .A2(_u10_u3_n2461 ), .ZN(_u10_u3_n1948 ) );
OR2_X1 _u10_u3_U613  ( .A1(_u10_u3_n1847 ), .A2(_u10_u3_n1948 ), .ZN(_u10_u3_n2811 ) );
NAND3_X1 _u10_u3_U612  ( .A1(_u10_u3_n2809 ), .A2(_u10_u3_n2810 ), .A3(_u10_u3_n2811 ), .ZN(_u10_u3_n2805 ) );
NOR2_X1 _u10_u3_U611  ( .A1(_u10_u3_n2808 ), .A2(_u10_u3_n2775 ), .ZN(_u10_u3_n2806 ) );
AND2_X1 _u10_u3_U610  ( .A1(_u10_u3_n2721 ), .A2(_u10_u3_n1911 ), .ZN(_u10_u3_n2807 ) );
NOR4_X1 _u10_u3_U609  ( .A1(_u10_u3_n2804 ), .A2(_u10_u3_n2805 ), .A3(_u10_u3_n2806 ), .A4(_u10_u3_n2807 ), .ZN(_u10_u3_n2726 ) );
NAND2_X1 _u10_u3_U608  ( .A1(_u10_u3_n2803 ), .A2(_u10_u3_n2112 ), .ZN(_u10_u3_n2802 ) );
NAND2_X1 _u10_u3_U607  ( .A1(_u10_u3_n2364 ), .A2(_u10_u3_n2802 ), .ZN(_u10_u3_n2801 ) );
NAND2_X1 _u10_u3_U606  ( .A1(_u10_u3_n2800 ), .A2(_u10_u3_n2801 ), .ZN(_u10_u3_n2799 ) );
NAND2_X1 _u10_u3_U605  ( .A1(_u10_u3_n1937 ), .A2(_u10_u3_n2799 ), .ZN(_u10_u3_n2780 ) );
NAND2_X1 _u10_u3_U604  ( .A1(_u10_u3_n2775 ), .A2(_u10_u3_n2798 ), .ZN(_u10_u3_n2796 ) );
INV_X1 _u10_u3_U603  ( .A(_u10_u3_n2131 ), .ZN(_u10_u3_n2797 ) );
NAND2_X1 _u10_u3_U602  ( .A1(_u10_u3_n2796 ), .A2(_u10_u3_n2797 ), .ZN(_u10_u3_n2781 ) );
OR4_X1 _u10_u3_U601  ( .A1(_u10_u3_n2795 ), .A2(_u10_u3_n2303 ), .A3(_u10_u3_n2553 ), .A4(_u10_u3_n2554 ), .ZN(_u10_u3_n2792 ) );
NAND3_X1 _u10_u3_U600  ( .A1(_u10_u3_n1847 ), .A2(_u10_u3_n2097 ), .A3(_u10_u3_n2096 ), .ZN(_u10_u3_n2793 ) );
NOR4_X1 _u10_u3_U599  ( .A1(_u10_u3_n2792 ), .A2(_u10_u3_n2793 ), .A3(_u10_u3_n2542 ), .A4(_u10_u3_n2794 ), .ZN(_u10_u3_n2791 ) );
NOR2_X1 _u10_u3_U598  ( .A1(_u10_u3_n2791 ), .A2(_u10_u3_n2085 ), .ZN(_u10_u3_n2783 ) );
NAND2_X1 _u10_u3_U597  ( .A1(_u10_u3_n2114 ), .A2(_u10_u3_n2049 ), .ZN(_u10_u3_n2700 ) );
INV_X1 _u10_u3_U596  ( .A(_u10_u3_n2700 ), .ZN(_u10_u3_n2784 ) );
NAND4_X1 _u10_u3_U595  ( .A1(_u10_u3_n2001 ), .A2(_u10_u3_n2547 ), .A3(_u10_u3_n2368 ), .A4(_u10_u3_n1847 ), .ZN(_u10_u3_n2787 ) );
NOR4_X1 _u10_u3_U594  ( .A1(_u10_u3_n2787 ), .A2(_u10_u3_n2788 ), .A3(_u10_u3_n2789 ), .A4(_u10_u3_n2790 ), .ZN(_u10_u3_n2786 ) );
NOR2_X1 _u10_u3_U593  ( .A1(_u10_u3_n2786 ), .A2(_u10_u3_n2000 ), .ZN(_u10_u3_n2785 ) );
NOR3_X1 _u10_u3_U592  ( .A1(_u10_u3_n2783 ), .A2(_u10_u3_n2784 ), .A3(_u10_u3_n2785 ), .ZN(_u10_u3_n2782 ) );
NAND3_X1 _u10_u3_U591  ( .A1(_u10_u3_n2780 ), .A2(_u10_u3_n2781 ), .A3(_u10_u3_n2782 ), .ZN(_u10_u3_n2728 ) );
OR3_X1 _u10_u3_U590  ( .A1(_u10_u3_n2138 ), .A2(_u10_u3_n2633 ), .A3(_u10_u3_n2779 ), .ZN(_u10_u3_n2778 ) );
NAND2_X1 _u10_u3_U589  ( .A1(_u10_u3_n2777 ), .A2(_u10_u3_n2778 ), .ZN(_u10_u3_n2767 ) );
NAND3_X1 _u10_u3_U588  ( .A1(_u10_u3_n2775 ), .A2(_u10_u3_n2083 ), .A3(_u10_u3_n2776 ), .ZN(_u10_u3_n2774 ) );
NAND2_X1 _u10_u3_U587  ( .A1(_u10_u3_n2773 ), .A2(_u10_u3_n2774 ), .ZN(_u10_u3_n2768 ) );
NAND2_X1 _u10_u3_U586  ( .A1(_u10_u3_n2218 ), .A2(_u10_u3_n2772 ), .ZN(_u10_u3_n2769 ) );
NAND2_X1 _u10_u3_U585  ( .A1(_u10_u3_n2302 ), .A2(_u10_u3_n2467 ), .ZN(_u10_u3_n2771 ) );
NAND2_X1 _u10_u3_U584  ( .A1(_u10_u3_n2461 ), .A2(_u10_u3_n2771 ), .ZN(_u10_u3_n2770 ) );
NAND4_X1 _u10_u3_U583  ( .A1(_u10_u3_n2767 ), .A2(_u10_u3_n2768 ), .A3(_u10_u3_n2769 ), .A4(_u10_u3_n2770 ), .ZN(_u10_u3_n2729 ) );
NAND3_X1 _u10_u3_U582  ( .A1(_u10_u3_n2668 ), .A2(_u10_u3_n2600 ), .A3(_u10_u3_n2276 ), .ZN(_u10_u3_n2766 ) );
NAND2_X1 _u10_u3_U581  ( .A1(_u10_u3_n1894 ), .A2(_u10_u3_n2766 ), .ZN(_u10_u3_n2753 ) );
NAND3_X1 _u10_u3_U580  ( .A1(_u10_u3_n2456 ), .A2(_u10_u3_n2744 ), .A3(_u10_u3_n2765 ), .ZN(_u10_u3_n2764 ) );
NAND2_X1 _u10_u3_U579  ( .A1(_u10_u3_n2377 ), .A2(_u10_u3_n2764 ), .ZN(_u10_u3_n2754 ) );
NAND2_X1 _u10_u3_U578  ( .A1(_u10_u3_n2763 ), .A2(_u10_u3_n2007 ), .ZN(_u10_u3_n2755 ) );
NOR2_X1 _u10_u3_U577  ( .A1(_u10_u3_n2531 ), .A2(_u10_u3_n2744 ), .ZN(_u10_u3_n2760 ) );
INV_X1 _u10_u3_U576  ( .A(_u10_u3_n2762 ), .ZN(_u10_u3_n2189 ) );
NOR3_X1 _u10_u3_U575  ( .A1(_u10_u3_n2760 ), .A2(_u10_u3_n2761 ), .A3(_u10_u3_n2189 ), .ZN(_u10_u3_n2759 ) );
NOR2_X1 _u10_u3_U574  ( .A1(_u10_u3_n2759 ), .A2(_u10_u3_n1849 ), .ZN(_u10_u3_n2757 ) );
NOR2_X1 _u10_u3_U573  ( .A1(_u10_u3_n1817 ), .A2(_u10_u3_n2665 ), .ZN(_u10_u3_n2758 ) );
NOR2_X1 _u10_u3_U572  ( .A1(_u10_u3_n2757 ), .A2(_u10_u3_n2758 ), .ZN(_u10_u3_n2756 ) );
NAND4_X1 _u10_u3_U571  ( .A1(_u10_u3_n2753 ), .A2(_u10_u3_n2754 ), .A3(_u10_u3_n2755 ), .A4(_u10_u3_n2756 ), .ZN(_u10_u3_n2730 ) );
INV_X1 _u10_u3_U570  ( .A(_u10_u3_n2359 ), .ZN(_u10_u3_n1899 ) );
NAND4_X1 _u10_u3_U569  ( .A1(_u10_u3_n2078 ), .A2(_u10_u3_n2580 ), .A3(_u10_u3_n2748 ), .A4(_u10_u3_n2752 ), .ZN(_u10_u3_n2751 ) );
NAND2_X1 _u10_u3_U568  ( .A1(_u10_u3_n1899 ), .A2(_u10_u3_n2751 ), .ZN(_u10_u3_n2732 ) );
INV_X1 _u10_u3_U567  ( .A(_u10_u3_n2750 ), .ZN(_u10_u3_n2379 ) );
NAND3_X1 _u10_u3_U566  ( .A1(_u10_u3_n1856 ), .A2(_u10_u3_n2669 ), .A3(_u10_u3_n2364 ), .ZN(_u10_u3_n2749 ) );
AND2_X1 _u10_u3_U565  ( .A1(_u10_u3_n2748 ), .A2(_u10_u3_n2749 ), .ZN(_u10_u3_n2034 ) );
NAND2_X1 _u10_u3_U564  ( .A1(_u10_u3_n2105 ), .A2(_u10_u3_n2669 ), .ZN(_u10_u3_n2745 ) );
AND3_X1 _u10_u3_U563  ( .A1(_u10_u3_n2745 ), .A2(_u10_u3_n2746 ), .A3(_u10_u3_n2747 ), .ZN(_u10_u3_n2380 ) );
NOR2_X1 _u10_u3_U562  ( .A1(_u10_u3_n2274 ), .A2(_u10_u3_n2744 ), .ZN(_u10_u3_n2743 ) );
NOR4_X1 _u10_u3_U561  ( .A1(_u10_u3_n2742 ), .A2(_u10_u3_n2680 ), .A3(_u10_u3_n2743 ), .A4(_u10_u3_n2428 ), .ZN(_u10_u3_n2741 ) );
NAND4_X1 _u10_u3_U560  ( .A1(_u10_u3_n2379 ), .A2(_u10_u3_n2034 ), .A3(_u10_u3_n2380 ), .A4(_u10_u3_n2741 ), .ZN(_u10_u3_n2740 ) );
NAND2_X1 _u10_u3_U559  ( .A1(_u10_u3_n1967 ), .A2(_u10_u3_n2740 ), .ZN(_u10_u3_n2733 ) );
NAND3_X1 _u10_u3_U558  ( .A1(_u10_u3_n2739 ), .A2(_u10_u3_n2368 ), .A3(_u10_u3_n2255 ), .ZN(_u10_u3_n2738 ) );
NAND2_X1 _u10_u3_U557  ( .A1(_u10_u3_n2737 ), .A2(_u10_u3_n2738 ), .ZN(_u10_u3_n2734 ) );
NAND2_X1 _u10_u3_U556  ( .A1(_u10_u3_n2736 ), .A2(_u10_u3_n2524 ), .ZN(_u10_u3_n2735 ) );
NAND4_X1 _u10_u3_U555  ( .A1(_u10_u3_n2732 ), .A2(_u10_u3_n2733 ), .A3(_u10_u3_n2734 ), .A4(_u10_u3_n2735 ), .ZN(_u10_u3_n2731 ) );
NOR4_X1 _u10_u3_U554  ( .A1(_u10_u3_n2728 ), .A2(_u10_u3_n2729 ), .A3(_u10_u3_n2730 ), .A4(_u10_u3_n2731 ), .ZN(_u10_u3_n2727 ) );
NAND4_X1 _u10_u3_U553  ( .A1(_u10_u3_n2724 ), .A2(_u10_u3_n2725 ), .A3(_u10_u3_n2726 ), .A4(_u10_u3_n2727 ), .ZN(_u10_u3_n2723 ) );
MUX2_X1 _u10_u3_U552  ( .A(_u10_u3_n2723 ), .B(_u10_SYNOPSYS_UNCONNECTED_9 ),.S(_u10_u3_n1819 ), .Z(_u10_u3_n1809 ) );
NAND2_X1 _u10_u3_U551  ( .A1(_u10_u3_n2002 ), .A2(_u10_u3_n2722 ), .ZN(_u10_u3_n2713 ) );
NAND2_X1 _u10_u3_U550  ( .A1(_u10_u3_n2720 ), .A2(_u10_u3_n2721 ), .ZN(_u10_u3_n2714 ) );
NAND2_X1 _u10_u3_U549  ( .A1(_u10_u3_n2256 ), .A2(_u10_u3_n2719 ), .ZN(_u10_u3_n2715 ) );
NOR2_X1 _u10_u3_U548  ( .A1(_u10_u3_n2106 ), .A2(_u10_u3_n2037 ), .ZN(_u10_u3_n2717 ) );
AND2_X1 _u10_u3_U547  ( .A1(_u10_u3_n1966 ), .A2(_u10_u3_n2054 ), .ZN(_u10_u3_n2718 ) );
NOR2_X1 _u10_u3_U546  ( .A1(_u10_u3_n2717 ), .A2(_u10_u3_n2718 ), .ZN(_u10_u3_n2716 ) );
NAND4_X1 _u10_u3_U545  ( .A1(_u10_u3_n2713 ), .A2(_u10_u3_n2714 ), .A3(_u10_u3_n2715 ), .A4(_u10_u3_n2716 ), .ZN(_u10_u3_n2608 ) );
NAND2_X1 _u10_u3_U544  ( .A1(1'b0), .A2(_u10_u3_n2669 ), .ZN(_u10_u3_n2385 ));
INV_X1 _u10_u3_U543  ( .A(_u10_u3_n2385 ), .ZN(_u10_u3_n1977 ) );
NAND2_X1 _u10_u3_U542  ( .A1(_u10_u3_n1977 ), .A2(_u10_u3_n2668 ), .ZN(_u10_u3_n2712 ) );
NAND2_X1 _u10_u3_U541  ( .A1(_u10_u3_n2712 ), .A2(_u10_u3_n2092 ), .ZN(_u10_u3_n1844 ) );
NAND2_X1 _u10_u3_U540  ( .A1(_u10_u3_n1894 ), .A2(_u10_u3_n1844 ), .ZN(_u10_u3_n2705 ) );
NAND2_X1 _u10_u3_U539  ( .A1(_u10_u3_n1894 ), .A2(_u10_u3_n2305 ), .ZN(_u10_u3_n2711 ) );
NAND2_X1 _u10_u3_U538  ( .A1(_u10_u3_n2711 ), .A2(_u10_u3_n2025 ), .ZN(_u10_u3_n1932 ) );
NAND2_X1 _u10_u3_U537  ( .A1(_u10_u3_n2710 ), .A2(_u10_u3_n1932 ), .ZN(_u10_u3_n2706 ) );
NAND2_X1 _u10_u3_U536  ( .A1(_u10_u3_n2708 ), .A2(_u10_u3_n2709 ), .ZN(_u10_u3_n2707 ) );
NAND3_X1 _u10_u3_U535  ( .A1(_u10_u3_n2705 ), .A2(_u10_u3_n2706 ), .A3(_u10_u3_n2707 ), .ZN(_u10_u3_n2701 ) );
NOR2_X1 _u10_u3_U534  ( .A1(_u10_u3_n1843 ), .A2(_u10_u3_n2545 ), .ZN(_u10_u3_n2702 ) );
NOR2_X1 _u10_u3_U533  ( .A1(_u10_u3_n2346 ), .A2(_u10_u3_n2700 ), .ZN(_u10_u3_n2703 ) );
NOR2_X1 _u10_u3_U532  ( .A1(_u10_u3_n2000 ), .A2(_u10_u3_n1887 ), .ZN(_u10_u3_n2704 ) );
NOR4_X1 _u10_u3_U531  ( .A1(_u10_u3_n2701 ), .A2(_u10_u3_n2702 ), .A3(_u10_u3_n2703 ), .A4(_u10_u3_n2704 ), .ZN(_u10_u3_n2671 ) );
NAND2_X1 _u10_u3_U530  ( .A1(_u10_u3_n2699 ), .A2(_u10_u3_n2700 ), .ZN(_u10_u3_n2698 ) );
NAND2_X1 _u10_u3_U529  ( .A1(_u10_u3_n2063 ), .A2(_u10_u3_n2698 ), .ZN(_u10_u3_n2682 ) );
NAND2_X1 _u10_u3_U528  ( .A1(_u10_u3_n2697 ), .A2(_u10_u3_n2103 ), .ZN(_u10_u3_n2696 ) );
NAND2_X1 _u10_u3_U527  ( .A1(_u10_u3_n2695 ), .A2(_u10_u3_n2696 ), .ZN(_u10_u3_n2694 ) );
NAND2_X1 _u10_u3_U526  ( .A1(_u10_u3_n1937 ), .A2(_u10_u3_n2694 ), .ZN(_u10_u3_n2683 ) );
INV_X1 _u10_u3_U525  ( .A(_u10_u3_n2693 ), .ZN(_u10_u3_n2691 ) );
NAND3_X1 _u10_u3_U524  ( .A1(_u10_u3_n2103 ), .A2(_u10_u3_n2502 ), .A3(1'b0),.ZN(_u10_u3_n2692 ) );
NAND2_X1 _u10_u3_U523  ( .A1(_u10_u3_n2691 ), .A2(_u10_u3_n2692 ), .ZN(_u10_u3_n2690 ) );
NAND2_X1 _u10_u3_U522  ( .A1(_u10_u3_n2236 ), .A2(_u10_u3_n2690 ), .ZN(_u10_u3_n2684 ) );
NAND3_X1 _u10_u3_U521  ( .A1(_u10_u3_n2688 ), .A2(_u10_u3_n1913 ), .A3(_u10_u3_n2689 ), .ZN(_u10_u3_n2335 ) );
NAND3_X1 _u10_u3_U520  ( .A1(_u10_u3_n2536 ), .A2(_u10_u3_n2103 ), .A3(1'b0),.ZN(_u10_u3_n2052 ) );
NOR2_X1 _u10_u3_U519  ( .A1(_u10_u3_n2052 ), .A2(_u10_u3_n2687 ), .ZN(_u10_u3_n1851 ) );
NAND2_X1 _u10_u3_U518  ( .A1(_u10_u3_n1851 ), .A2(_u10_u3_n2078 ), .ZN(_u10_u3_n2582 ) );
NOR2_X1 _u10_u3_U517  ( .A1(_u10_u3_n2686 ), .A2(_u10_u3_n2582 ), .ZN(_u10_u3_n2094 ) );
NAND3_X1 _u10_u3_U516  ( .A1(_u10_u3_n2251 ), .A2(_u10_u3_n2335 ), .A3(_u10_u3_n2094 ), .ZN(_u10_u3_n2685 ) );
NAND4_X1 _u10_u3_U515  ( .A1(_u10_u3_n2682 ), .A2(_u10_u3_n2683 ), .A3(_u10_u3_n2684 ), .A4(_u10_u3_n2685 ), .ZN(_u10_u3_n2673 ) );
INV_X1 _u10_u3_U514  ( .A(_u10_u3_n2291 ), .ZN(_u10_u3_n2057 ) );
AND2_X1 _u10_u3_U513  ( .A1(_u10_u3_n1851 ), .A2(_u10_u3_n2057 ), .ZN(_u10_u3_n2674 ) );
INV_X1 _u10_u3_U512  ( .A(_u10_u3_n1874 ), .ZN(_u10_u3_n2681 ) );
NOR2_X1 _u10_u3_U511  ( .A1(_u10_u3_n2007 ), .A2(_u10_u3_n1911 ), .ZN(_u10_u3_n2486 ) );
NOR2_X1 _u10_u3_U510  ( .A1(_u10_u3_n2681 ), .A2(_u10_u3_n2486 ), .ZN(_u10_u3_n2675 ) );
NOR2_X1 _u10_u3_U509  ( .A1(_u10_u3_n1977 ), .A2(_u10_u3_n2680 ), .ZN(_u10_u3_n2679 ) );
NOR2_X1 _u10_u3_U508  ( .A1(_u10_u3_n2679 ), .A2(_u10_u3_n2030 ), .ZN(_u10_u3_n2678 ) );
NOR2_X1 _u10_u3_U507  ( .A1(_u10_u3_n2678 ), .A2(_u10_u3_n2094 ), .ZN(_u10_u3_n2677 ) );
NOR2_X1 _u10_u3_U506  ( .A1(_u10_u3_n2677 ), .A2(_u10_u3_n2025 ), .ZN(_u10_u3_n2676 ) );
NOR4_X1 _u10_u3_U505  ( .A1(_u10_u3_n2673 ), .A2(_u10_u3_n2674 ), .A3(_u10_u3_n2675 ), .A4(_u10_u3_n2676 ), .ZN(_u10_u3_n2672 ) );
AND2_X1 _u10_u3_U504  ( .A1(_u10_u3_n2671 ), .A2(_u10_u3_n2672 ), .ZN(_u10_u3_n1990 ) );
INV_X1 _u10_u3_U503  ( .A(_u10_u3_n2670 ), .ZN(_u10_u3_n2660 ) );
NAND4_X1 _u10_u3_U502  ( .A1(_u10_u3_n2251 ), .A2(_u10_u3_n2669 ), .A3(_u10_u3_n2162 ), .A4(_u10_u3_n2169 ), .ZN(_u10_u3_n2664 ) );
AND3_X1 _u10_u3_U501  ( .A1(_u10_u3_n1977 ), .A2(_u10_u3_n2668 ), .A3(_u10_u3_n2089 ), .ZN(_u10_u3_n2555 ) );
NAND2_X1 _u10_u3_U500  ( .A1(_u10_u3_n2555 ), .A2(_u10_u3_n2667 ), .ZN(_u10_u3_n2666 ) );
NAND3_X1 _u10_u3_U499  ( .A1(_u10_u3_n2664 ), .A2(_u10_u3_n2665 ), .A3(_u10_u3_n2666 ), .ZN(_u10_u3_n1988 ) );
INV_X1 _u10_u3_U498  ( .A(_u10_u3_n1988 ), .ZN(_u10_u3_n2661 ) );
NAND2_X1 _u10_u3_U497  ( .A1(1'b0), .A2(_u10_u3_n2043 ), .ZN(_u10_u3_n2662 ));
NAND2_X1 _u10_u3_U496  ( .A1(_u10_u3_n2169 ), .A2(1'b0), .ZN(_u10_u3_n2663 ));
NAND4_X1 _u10_u3_U495  ( .A1(_u10_u3_n2660 ), .A2(_u10_u3_n2661 ), .A3(_u10_u3_n2662 ), .A4(_u10_u3_n2663 ), .ZN(_u10_u3_n2650 ) );
NAND2_X1 _u10_u3_U494  ( .A1(_u10_u3_n2659 ), .A2(1'b0), .ZN(_u10_u3_n2193 ));
INV_X1 _u10_u3_U493  ( .A(_u10_u3_n2193 ), .ZN(_u10_u3_n2143 ) );
NAND2_X1 _u10_u3_U492  ( .A1(_u10_u3_n2143 ), .A2(_u10_u3_n2036 ), .ZN(_u10_u3_n2286 ) );
INV_X1 _u10_u3_U491  ( .A(_u10_u3_n2286 ), .ZN(_u10_u3_n2577 ) );
NAND2_X1 _u10_u3_U490  ( .A1(_u10_u3_n2577 ), .A2(_u10_u3_n2278 ), .ZN(_u10_u3_n2474 ) );
INV_X1 _u10_u3_U489  ( .A(_u10_u3_n2474 ), .ZN(_u10_u3_n2306 ) );
NAND2_X1 _u10_u3_U488  ( .A1(_u10_u3_n2306 ), .A2(_u10_u3_n2251 ), .ZN(_u10_u3_n2654 ) );
NAND2_X1 _u10_u3_U487  ( .A1(_u10_u3_n2649 ), .A2(_u10_u3_n2658 ), .ZN(_u10_u3_n2655 ) );
NAND2_X1 _u10_u3_U486  ( .A1(_u10_u3_n2657 ), .A2(_u10_u3_n2445 ), .ZN(_u10_u3_n2656 ) );
NAND3_X1 _u10_u3_U485  ( .A1(_u10_u3_n2654 ), .A2(_u10_u3_n2655 ), .A3(_u10_u3_n2656 ), .ZN(_u10_u3_n2651 ) );
NOR2_X1 _u10_u3_U484  ( .A1(_u10_u3_n2366 ), .A2(_u10_u3_n2376 ), .ZN(_u10_u3_n2652 ) );
AND2_X1 _u10_u3_U483  ( .A1(_u10_u3_n1966 ), .A2(_u10_u3_n2528 ), .ZN(_u10_u3_n2653 ) );
NOR4_X1 _u10_u3_U482  ( .A1(_u10_u3_n2650 ), .A2(_u10_u3_n2651 ), .A3(_u10_u3_n2652 ), .A4(_u10_u3_n2653 ), .ZN(_u10_u3_n2613 ) );
NAND2_X1 _u10_u3_U481  ( .A1(_u10_u3_n1891 ), .A2(1'b0), .ZN(_u10_u3_n2636 ));
NAND2_X1 _u10_u3_U480  ( .A1(_u10_u3_n1868 ), .A2(_u10_u3_n2113 ), .ZN(_u10_u3_n2101 ) );
NOR4_X1 _u10_u3_U479  ( .A1(_u10_u3_n2649 ), .A2(_u10_u3_n2216 ), .A3(_u10_u3_n2101 ), .A4(_u10_u3_n2634 ), .ZN(_u10_u3_n2648 ) );
NOR2_X1 _u10_u3_U478  ( .A1(_u10_u3_n2648 ), .A2(_u10_u3_n2254 ), .ZN(_u10_u3_n2638 ) );
NOR2_X1 _u10_u3_U477  ( .A1(_u10_u3_n2106 ), .A2(_u10_u3_n2643 ), .ZN(_u10_u3_n2645 ) );
NAND2_X1 _u10_u3_U476  ( .A1(1'b0), .A2(_u10_u3_n2049 ), .ZN(_u10_u3_n2647 ));
NAND2_X1 _u10_u3_U475  ( .A1(_u10_u3_n2646 ), .A2(_u10_u3_n2647 ), .ZN(_u10_u3_n2348 ) );
NOR2_X1 _u10_u3_U474  ( .A1(_u10_u3_n2645 ), .A2(_u10_u3_n2348 ), .ZN(_u10_u3_n2644 ) );
NOR2_X1 _u10_u3_U473  ( .A1(_u10_u3_n2644 ), .A2(_u10_u3_n2495 ), .ZN(_u10_u3_n2639 ) );
NOR2_X1 _u10_u3_U472  ( .A1(_u10_u3_n2643 ), .A2(_u10_u3_n2203 ), .ZN(_u10_u3_n2642 ) );
NOR3_X1 _u10_u3_U471  ( .A1(_u10_u3_n2101 ), .A2(1'b0), .A3(_u10_u3_n2642 ),.ZN(_u10_u3_n2641 ) );
NOR2_X1 _u10_u3_U470  ( .A1(_u10_u3_n2641 ), .A2(_u10_u3_n2253 ), .ZN(_u10_u3_n2640 ) );
NOR3_X1 _u10_u3_U469  ( .A1(_u10_u3_n2638 ), .A2(_u10_u3_n2639 ), .A3(_u10_u3_n2640 ), .ZN(_u10_u3_n2637 ) );
NAND3_X1 _u10_u3_U468  ( .A1(_u10_u3_n2635 ), .A2(_u10_u3_n2636 ), .A3(_u10_u3_n2637 ), .ZN(_u10_u3_n2615 ) );
NOR3_X1 _u10_u3_U467  ( .A1(_u10_u3_n2174 ), .A2(_u10_u3_n2175 ), .A3(_u10_u3_n2179 ), .ZN(_u10_u3_n2631 ) );
NAND3_X1 _u10_u3_U466  ( .A1(_u10_u3_n2223 ), .A2(_u10_u3_n2236 ), .A3(_u10_u3_n2631 ), .ZN(_u10_u3_n2622 ) );
OR2_X1 _u10_u3_U465  ( .A1(_u10_u3_n1960 ), .A2(_u10_u3_n1959 ), .ZN(_u10_u3_n2625 ) );
NOR3_X1 _u10_u3_U464  ( .A1(_u10_u3_n2101 ), .A2(_u10_u3_n2633 ), .A3(_u10_u3_n2634 ), .ZN(_u10_u3_n2523 ) );
OR2_X1 _u10_u3_U463  ( .A1(_u10_u3_n2632 ), .A2(_u10_u3_n2523 ), .ZN(_u10_u3_n2627 ) );
INV_X1 _u10_u3_U462  ( .A(_u10_u3_n2631 ), .ZN(_u10_u3_n2628 ) );
NAND2_X1 _u10_u3_U461  ( .A1(_u10_u3_n2630 ), .A2(_u10_u3_n1922 ), .ZN(_u10_u3_n2629 ) );
NAND3_X1 _u10_u3_U460  ( .A1(_u10_u3_n2627 ), .A2(_u10_u3_n2628 ), .A3(_u10_u3_n2629 ), .ZN(_u10_u3_n2626 ) );
NAND2_X1 _u10_u3_U459  ( .A1(_u10_u3_n2625 ), .A2(_u10_u3_n2626 ), .ZN(_u10_u3_n2624 ) );
NAND3_X1 _u10_u3_U458  ( .A1(_u10_u3_n2622 ), .A2(_u10_u3_n2623 ), .A3(_u10_u3_n2624 ), .ZN(_u10_u3_n2616 ) );
AND2_X1 _u10_u3_U457  ( .A1(_u10_u3_n2621 ), .A2(_u10_u3_n2358 ), .ZN(_u10_u3_n2620 ) );
NOR2_X1 _u10_u3_U456  ( .A1(_u10_u3_n2523 ), .A2(_u10_u3_n2620 ), .ZN(_u10_u3_n2617 ) );
INV_X1 _u10_u3_U455  ( .A(_u10_u3_n2101 ), .ZN(_u10_u3_n2221 ) );
NOR2_X1 _u10_u3_U454  ( .A1(_u10_u3_n1911 ), .A2(_u10_u3_n2488 ), .ZN(_u10_u3_n2619 ) );
NOR2_X1 _u10_u3_U453  ( .A1(_u10_u3_n2221 ), .A2(_u10_u3_n2619 ), .ZN(_u10_u3_n2618 ) );
NOR4_X1 _u10_u3_U452  ( .A1(_u10_u3_n2615 ), .A2(_u10_u3_n2616 ), .A3(_u10_u3_n2617 ), .A4(_u10_u3_n2618 ), .ZN(_u10_u3_n2614 ) );
AND2_X1 _u10_u3_U451  ( .A1(_u10_u3_n2613 ), .A2(_u10_u3_n2614 ), .ZN(_u10_u3_n2314 ) );
NAND3_X1 _u10_u3_U450  ( .A1(_u10_u3_n2612 ), .A2(_u10_u3_n1990 ), .A3(_u10_u3_n2314 ), .ZN(_u10_u3_n2609 ) );
NOR4_X1 _u10_u3_U449  ( .A1(_u10_u3_n2608 ), .A2(_u10_u3_n2609 ), .A3(_u10_u3_n2610 ), .A4(_u10_u3_n2611 ), .ZN(_u10_u3_n2388 ) );
NAND2_X1 _u10_u3_U448  ( .A1(_u10_u3_n2346 ), .A2(_u10_u3_n2607 ), .ZN(_u10_u3_n2191 ) );
NAND2_X1 _u10_u3_U447  ( .A1(_u10_u3_n2143 ), .A2(_u10_u3_n2191 ), .ZN(_u10_u3_n2556 ) );
INV_X1 _u10_u3_U446  ( .A(_u10_u3_n2348 ), .ZN(_u10_u3_n2603 ) );
NAND3_X1 _u10_u3_U445  ( .A1(_u10_u3_n2535 ), .A2(_u10_u3_n2485 ), .A3(_u10_u3_n2456 ), .ZN(_u10_u3_n2606 ) );
NAND2_X1 _u10_u3_U444  ( .A1(_u10_u3_n2049 ), .A2(_u10_u3_n2606 ), .ZN(_u10_u3_n2604 ) );
NAND3_X1 _u10_u3_U443  ( .A1(_u10_u3_n2603 ), .A2(_u10_u3_n2604 ), .A3(_u10_u3_n2605 ), .ZN(_u10_u3_n2602 ) );
NAND2_X1 _u10_u3_U442  ( .A1(_u10_u3_n2043 ), .A2(_u10_u3_n2602 ), .ZN(_u10_u3_n2557 ) );
INV_X1 _u10_u3_U441  ( .A(_u10_u3_n2601 ), .ZN(_u10_u3_n2590 ) );
NAND2_X1 _u10_u3_U440  ( .A1(_u10_u3_n2599 ), .A2(_u10_u3_n2600 ), .ZN(_u10_u3_n2597 ) );
NAND2_X1 _u10_u3_U439  ( .A1(_u10_u3_n2082 ), .A2(_u10_u3_n2101 ), .ZN(_u10_u3_n2598 ) );
AND2_X1 _u10_u3_U438  ( .A1(_u10_u3_n2597 ), .A2(_u10_u3_n2598 ), .ZN(_u10_u3_n2281 ) );
NAND3_X1 _u10_u3_U437  ( .A1(_u10_u3_n1969 ), .A2(_u10_u3_n2582 ), .A3(_u10_u3_n2281 ), .ZN(_u10_u3_n2073 ) );
INV_X1 _u10_u3_U436  ( .A(_u10_u3_n2073 ), .ZN(_u10_u3_n2591 ) );
NOR2_X1 _u10_u3_U435  ( .A1(_u10_u3_n1816 ), .A2(_u10_u3_n2077 ), .ZN(_u10_u3_n2595 ) );
NOR2_X1 _u10_u3_U434  ( .A1(_u10_u3_n2595 ), .A2(_u10_u3_n2596 ), .ZN(_u10_u3_n2592 ) );
NAND3_X1 _u10_u3_U433  ( .A1(_u10_u3_n2107 ), .A2(_u10_u3_n2536 ), .A3(1'b0),.ZN(_u10_u3_n2438 ) );
INV_X1 _u10_u3_U432  ( .A(_u10_u3_n2438 ), .ZN(_u10_u3_n2427 ) );
NOR4_X1 _u10_u3_U431  ( .A1(1'b0), .A2(_u10_u3_n2594 ), .A3(_u10_u3_n2577 ),.A4(_u10_u3_n2427 ), .ZN(_u10_u3_n2593 ) );
NAND4_X1 _u10_u3_U430  ( .A1(_u10_u3_n2590 ), .A2(_u10_u3_n2591 ), .A3(_u10_u3_n2592 ), .A4(_u10_u3_n2593 ), .ZN(_u10_u3_n2589 ) );
NAND2_X1 _u10_u3_U429  ( .A1(_u10_u3_n2279 ), .A2(_u10_u3_n2589 ), .ZN(_u10_u3_n2558 ) );
NAND3_X1 _u10_u3_U428  ( .A1(_u10_u3_n2587 ), .A2(_u10_u3_n2115 ), .A3(_u10_u3_n2588 ), .ZN(_u10_u3_n2585 ) );
NOR4_X1 _u10_u3_U427  ( .A1(_u10_u3_n2585 ), .A2(_u10_u3_n2586 ), .A3(1'b0),.A4(_u10_u3_n2114 ), .ZN(_u10_u3_n2583 ) );
NOR2_X1 _u10_u3_U426  ( .A1(_u10_u3_n2583 ), .A2(_u10_u3_n2584 ), .ZN(_u10_u3_n2560 ) );
OR2_X1 _u10_u3_U425  ( .A1(_u10_u3_n2582 ), .A2(1'b0), .ZN(_u10_u3_n2581 ));
NAND2_X1 _u10_u3_U424  ( .A1(_u10_u3_n2580 ), .A2(_u10_u3_n2581 ), .ZN(_u10_u3_n1974 ) );
INV_X1 _u10_u3_U423  ( .A(_u10_u3_n1974 ), .ZN(_u10_u3_n1901 ) );
AND4_X1 _u10_u3_U422  ( .A1(_u10_u3_n1901 ), .A2(_u10_u3_n2385 ), .A3(_u10_u3_n2578 ), .A4(_u10_u3_n2579 ), .ZN(_u10_u3_n2424 ) );
NOR2_X1 _u10_u3_U421  ( .A1(1'b0), .A2(_u10_u3_n2424 ), .ZN(_u10_u3_n2574 ));
NOR3_X1 _u10_u3_U420  ( .A1(_u10_u3_n2427 ), .A2(1'b0), .A3(_u10_u3_n2577 ),.ZN(_u10_u3_n2576 ) );
NOR2_X1 _u10_u3_U419  ( .A1(_u10_u3_n2576 ), .A2(_u10_u3_n1976 ), .ZN(_u10_u3_n2575 ) );
NOR3_X1 _u10_u3_U418  ( .A1(_u10_u3_n2574 ), .A2(_u10_u3_n1979 ), .A3(_u10_u3_n2575 ), .ZN(_u10_u3_n2572 ) );
NOR2_X1 _u10_u3_U417  ( .A1(_u10_u3_n2572 ), .A2(_u10_u3_n2573 ), .ZN(_u10_u3_n2561 ) );
INV_X1 _u10_u3_U416  ( .A(_u10_u3_n2061 ), .ZN(_u10_u3_n2453 ) );
NOR2_X1 _u10_u3_U415  ( .A1(_u10_u3_n2453 ), .A2(_u10_u3_n1851 ), .ZN(_u10_u3_n2018 ) );
NAND2_X1 _u10_u3_U414  ( .A1(1'b0), .A2(_u10_u3_n2571 ), .ZN(_u10_u3_n2570 ));
NAND2_X1 _u10_u3_U413  ( .A1(_u10_u3_n2018 ), .A2(_u10_u3_n2570 ), .ZN(_u10_u3_n1837 ) );
INV_X1 _u10_u3_U412  ( .A(_u10_u3_n1837 ), .ZN(_u10_u3_n2568 ) );
NAND2_X1 _u10_u3_U411  ( .A1(1'b0), .A2(_u10_u3_n2536 ), .ZN(_u10_u3_n2569 ));
NAND2_X1 _u10_u3_U410  ( .A1(_u10_u3_n2568 ), .A2(_u10_u3_n2569 ), .ZN(_u10_u3_n2564 ) );
NOR2_X1 _u10_u3_U409  ( .A1(_u10_u3_n1841 ), .A2(_u10_u3_n1868 ), .ZN(_u10_u3_n2565 ) );
INV_X1 _u10_u3_U408  ( .A(_u10_u3_n2567 ), .ZN(_u10_u3_n2566 ) );
NOR4_X1 _u10_u3_U407  ( .A1(_u10_u3_n2564 ), .A2(_u10_u3_n2565 ), .A3(_u10_u3_n2143 ), .A4(_u10_u3_n2566 ), .ZN(_u10_u3_n2563 ) );
NOR2_X1 _u10_u3_U406  ( .A1(_u10_u3_n2563 ), .A2(_u10_u3_n2014 ), .ZN(_u10_u3_n2562 ) );
NOR3_X1 _u10_u3_U405  ( .A1(_u10_u3_n2560 ), .A2(_u10_u3_n2561 ), .A3(_u10_u3_n2562 ), .ZN(_u10_u3_n2559 ) );
NAND4_X1 _u10_u3_U404  ( .A1(_u10_u3_n2556 ), .A2(_u10_u3_n2557 ), .A3(_u10_u3_n2558 ), .A4(_u10_u3_n2559 ), .ZN(_u10_u3_n2511 ) );
INV_X1 _u10_u3_U403  ( .A(_u10_u3_n2085 ), .ZN(_u10_u3_n2293 ) );
NOR2_X1 _u10_u3_U402  ( .A1(_u10_u3_n2554 ), .A2(_u10_u3_n2555 ), .ZN(_u10_u3_n2444 ) );
NAND2_X1 _u10_u3_U401  ( .A1(_u10_u3_n2553 ), .A2(_u10_u3_n2549 ), .ZN(_u10_u3_n2552 ) );
AND2_X1 _u10_u3_U400  ( .A1(_u10_u3_n2444 ), .A2(_u10_u3_n2552 ), .ZN(_u10_u3_n2295 ) );
NAND2_X1 _u10_u3_U399  ( .A1(_u10_u3_n2551 ), .A2(_u10_u3_n2549 ), .ZN(_u10_u3_n2538 ) );
AND2_X1 _u10_u3_U398  ( .A1(_u10_u3_n2427 ), .A2(_u10_u3_n2108 ), .ZN(_u10_u3_n2460 ) );
NOR4_X1 _u10_u3_U397  ( .A1(_u10_u3_n2460 ), .A2(_u10_u3_n2306 ), .A3(_u10_u3_n2094 ), .A4(_u10_u3_n2550 ), .ZN(_u10_u3_n2409 ) );
INV_X1 _u10_u3_U396  ( .A(_u10_u3_n2409 ), .ZN(_u10_u3_n2407 ) );
NAND2_X1 _u10_u3_U395  ( .A1(_u10_u3_n2549 ), .A2(_u10_u3_n2407 ), .ZN(_u10_u3_n2546 ) );
NAND3_X1 _u10_u3_U394  ( .A1(_u10_u3_n2546 ), .A2(_u10_u3_n2547 ), .A3(_u10_u3_n2548 ), .ZN(_u10_u3_n2501 ) );
INV_X1 _u10_u3_U393  ( .A(_u10_u3_n2501 ), .ZN(_u10_u3_n2539 ) );
NOR2_X1 _u10_u3_U392  ( .A1(1'b0), .A2(_u10_u3_n2545 ), .ZN(_u10_u3_n2541 ));
AND2_X1 _u10_u3_U391  ( .A1(_u10_u3_n2544 ), .A2(_u10_u3_n2089 ), .ZN(_u10_u3_n2543 ) );
NOR3_X1 _u10_u3_U390  ( .A1(_u10_u3_n2541 ), .A2(_u10_u3_n2542 ), .A3(_u10_u3_n2543 ), .ZN(_u10_u3_n2540 ) );
NAND4_X1 _u10_u3_U389  ( .A1(_u10_u3_n2295 ), .A2(_u10_u3_n2538 ), .A3(_u10_u3_n2539 ), .A4(_u10_u3_n2540 ), .ZN(_u10_u3_n2537 ) );
NAND2_X1 _u10_u3_U388  ( .A1(_u10_u3_n2293 ), .A2(_u10_u3_n2537 ), .ZN(_u10_u3_n2515 ) );
NAND2_X1 _u10_u3_U387  ( .A1(_u10_u3_n2536 ), .A2(_u10_u3_n2508 ), .ZN(_u10_u3_n2526 ) );
NAND2_X1 _u10_u3_U386  ( .A1(_u10_u3_n2535 ), .A2(_u10_u3_n1940 ), .ZN(_u10_u3_n2532 ) );
NOR4_X1 _u10_u3_U385  ( .A1(_u10_u3_n2532 ), .A2(_u10_u3_n2533 ), .A3(1'b0),.A4(_u10_u3_n2534 ), .ZN(_u10_u3_n2530 ) );
NOR2_X1 _u10_u3_U384  ( .A1(_u10_u3_n2530 ), .A2(_u10_u3_n2531 ), .ZN(_u10_u3_n2529 ) );
NOR4_X1 _u10_u3_U383  ( .A1(_u10_u3_n2528 ), .A2(_u10_u3_n2143 ), .A3(_u10_u3_n2189 ), .A4(_u10_u3_n2529 ), .ZN(_u10_u3_n2527 ) );
NAND4_X1 _u10_u3_U382  ( .A1(_u10_u3_n2019 ), .A2(_u10_u3_n2526 ), .A3(_u10_u3_n2018 ), .A4(_u10_u3_n2527 ), .ZN(_u10_u3_n2525 ) );
NAND2_X1 _u10_u3_U381  ( .A1(_u10_u3_n2183 ), .A2(_u10_u3_n2525 ), .ZN(_u10_u3_n2516 ) );
INV_X1 _u10_u3_U380  ( .A(_u10_u3_n2524 ), .ZN(_u10_u3_n2396 ) );
NAND2_X1 _u10_u3_U379  ( .A1(_u10_u3_n2396 ), .A2(_u10_u3_n2523 ), .ZN(_u10_u3_n2522 ) );
NAND2_X1 _u10_u3_U378  ( .A1(_u10_u3_n1866 ), .A2(_u10_u3_n2522 ), .ZN(_u10_u3_n2519 ) );
AND2_X1 _u10_u3_U377  ( .A1(_u10_u3_n2493 ), .A2(_u10_u3_n1961 ), .ZN(_u10_u3_n2429 ) );
NAND2_X1 _u10_u3_U376  ( .A1(_u10_u3_n2429 ), .A2(_u10_u3_n2175 ), .ZN(_u10_u3_n2510 ) );
NAND2_X1 _u10_u3_U375  ( .A1(_u10_u3_n2510 ), .A2(_u10_u3_n1864 ), .ZN(_u10_u3_n2521 ) );
NAND3_X1 _u10_u3_U374  ( .A1(_u10_u3_n2519 ), .A2(_u10_u3_n2520 ), .A3(_u10_u3_n2521 ), .ZN(_u10_u3_n2518 ) );
NAND2_X1 _u10_u3_U373  ( .A1(_u10_u3_n1861 ), .A2(_u10_u3_n2518 ), .ZN(_u10_u3_n2517 ) );
NAND3_X1 _u10_u3_U372  ( .A1(_u10_u3_n2515 ), .A2(_u10_u3_n2516 ), .A3(_u10_u3_n2517 ), .ZN(_u10_u3_n2512 ) );
NOR2_X1 _u10_u3_U371  ( .A1(_u10_u3_n1913 ), .A2(_u10_u3_n1940 ), .ZN(_u10_u3_n2513 ) );
NOR2_X1 _u10_u3_U370  ( .A1(_u10_u3_n2113 ), .A2(_u10_u3_n2350 ), .ZN(_u10_u3_n2514 ) );
NOR4_X1 _u10_u3_U369  ( .A1(_u10_u3_n2511 ), .A2(_u10_u3_n2512 ), .A3(_u10_u3_n2513 ), .A4(_u10_u3_n2514 ), .ZN(_u10_u3_n2389 ) );
NAND2_X1 _u10_u3_U368  ( .A1(_u10_u3_n2509 ), .A2(_u10_u3_n2510 ), .ZN(_u10_u3_n2477 ) );
NAND2_X1 _u10_u3_U367  ( .A1(_u10_u3_n2507 ), .A2(_u10_u3_n2508 ), .ZN(_u10_u3_n2504 ) );
NAND2_X1 _u10_u3_U366  ( .A1(1'b0), .A2(_u10_u3_n2506 ), .ZN(_u10_u3_n2505 ));
NAND2_X1 _u10_u3_U365  ( .A1(_u10_u3_n2504 ), .A2(_u10_u3_n2505 ), .ZN(_u10_u3_n2503 ) );
NAND2_X1 _u10_u3_U364  ( .A1(_u10_u3_n2502 ), .A2(_u10_u3_n2503 ), .ZN(_u10_u3_n2478 ) );
NAND2_X1 _u10_u3_U363  ( .A1(_u10_u3_n2501 ), .A2(_u10_u3_n2446 ), .ZN(_u10_u3_n2497 ) );
INV_X1 _u10_u3_U362  ( .A(_u10_u3_n2500 ), .ZN(_u10_u3_n2499 ) );
NAND3_X1 _u10_u3_U361  ( .A1(_u10_u3_n2497 ), .A2(_u10_u3_n2498 ), .A3(_u10_u3_n2499 ), .ZN(_u10_u3_n2496 ) );
NAND2_X1 _u10_u3_U360  ( .A1(_u10_u3_n2445 ), .A2(_u10_u3_n2496 ), .ZN(_u10_u3_n2479 ) );
NOR2_X1 _u10_u3_U359  ( .A1(_u10_u3_n2429 ), .A2(_u10_u3_n2495 ), .ZN(_u10_u3_n2491 ) );
INV_X1 _u10_u3_U358  ( .A(_u10_u3_n2191 ), .ZN(_u10_u3_n2494 ) );
NOR2_X1 _u10_u3_U357  ( .A1(_u10_u3_n2493 ), .A2(_u10_u3_n2494 ), .ZN(_u10_u3_n2492 ) );
NOR2_X1 _u10_u3_U356  ( .A1(_u10_u3_n2491 ), .A2(_u10_u3_n2492 ), .ZN(_u10_u3_n2489 ) );
NOR2_X1 _u10_u3_U355  ( .A1(_u10_u3_n2489 ), .A2(_u10_u3_n2490 ), .ZN(_u10_u3_n2481 ) );
NAND2_X1 _u10_u3_U354  ( .A1(_u10_u3_n2253 ), .A2(_u10_u3_n1859 ), .ZN(_u10_u3_n2398 ) );
NOR2_X1 _u10_u3_U353  ( .A1(_u10_u3_n2488 ), .A2(_u10_u3_n2398 ), .ZN(_u10_u3_n2487 ) );
NOR2_X1 _u10_u3_U352  ( .A1(_u10_u3_n2220 ), .A2(_u10_u3_n2487 ), .ZN(_u10_u3_n2482 ) );
AND2_X1 _u10_u3_U351  ( .A1(_u10_u3_n2350 ), .A2(_u10_u3_n2486 ), .ZN(_u10_u3_n2484 ) );
NOR2_X1 _u10_u3_U350  ( .A1(_u10_u3_n2484 ), .A2(_u10_u3_n2485 ), .ZN(_u10_u3_n2483 ) );
NOR3_X1 _u10_u3_U349  ( .A1(_u10_u3_n2481 ), .A2(_u10_u3_n2482 ), .A3(_u10_u3_n2483 ), .ZN(_u10_u3_n2480 ) );
NAND4_X1 _u10_u3_U348  ( .A1(_u10_u3_n2477 ), .A2(_u10_u3_n2478 ), .A3(_u10_u3_n2479 ), .A4(_u10_u3_n2480 ), .ZN(_u10_u3_n2447 ) );
NAND2_X1 _u10_u3_U347  ( .A1(_u10_u3_n2476 ), .A2(_u10_u3_n1936 ), .ZN(_u10_u3_n2472 ) );
NAND2_X1 _u10_u3_U346  ( .A1(_u10_u3_n2427 ), .A2(_u10_u3_n2278 ), .ZN(_u10_u3_n2473 ) );
NAND4_X1 _u10_u3_U345  ( .A1(_u10_u3_n2472 ), .A2(_u10_u3_n2473 ), .A3(_u10_u3_n2474 ), .A4(_u10_u3_n2475 ), .ZN(_u10_u3_n2471 ) );
NAND2_X1 _u10_u3_U344  ( .A1(_u10_u3_n2470 ), .A2(_u10_u3_n2471 ), .ZN(_u10_u3_n2457 ) );
NAND2_X1 _u10_u3_U343  ( .A1(_u10_u3_n2409 ), .A2(_u10_u3_n2469 ), .ZN(_u10_u3_n2468 ) );
NAND2_X1 _u10_u3_U342  ( .A1(_u10_u3_n2467 ), .A2(_u10_u3_n2468 ), .ZN(_u10_u3_n2463 ) );
NAND2_X1 _u10_u3_U341  ( .A1(_u10_u3_n1844 ), .A2(_u10_u3_n2466 ), .ZN(_u10_u3_n2465 ) );
NAND3_X1 _u10_u3_U340  ( .A1(_u10_u3_n2463 ), .A2(_u10_u3_n2464 ), .A3(_u10_u3_n2465 ), .ZN(_u10_u3_n2462 ) );
NAND2_X1 _u10_u3_U339  ( .A1(_u10_u3_n2461 ), .A2(_u10_u3_n2462 ), .ZN(_u10_u3_n2458 ) );
NAND2_X1 _u10_u3_U338  ( .A1(_u10_u3_n2460 ), .A2(_u10_u3_n2251 ), .ZN(_u10_u3_n2459 ) );
NAND3_X1 _u10_u3_U337  ( .A1(_u10_u3_n2457 ), .A2(_u10_u3_n2458 ), .A3(_u10_u3_n2459 ), .ZN(_u10_u3_n2448 ) );
NOR2_X1 _u10_u3_U336  ( .A1(_u10_u3_n2455 ), .A2(_u10_u3_n2456 ), .ZN(_u10_u3_n2449 ) );
NAND2_X1 _u10_u3_U335  ( .A1(_u10_u3_n2454 ), .A2(_u10_u3_n2438 ), .ZN(_u10_u3_n2452 ) );
NOR4_X1 _u10_u3_U334  ( .A1(_u10_u3_n2452 ), .A2(_u10_u3_n2453 ), .A3(_u10_u3_n2443 ), .A4(_u10_u3_n2143 ), .ZN(_u10_u3_n2451 ) );
NOR2_X1 _u10_u3_U333  ( .A1(_u10_u3_n2451 ), .A2(_u10_u3_n2356 ), .ZN(_u10_u3_n2450 ) );
NOR4_X1 _u10_u3_U332  ( .A1(_u10_u3_n2447 ), .A2(_u10_u3_n2448 ), .A3(_u10_u3_n2449 ), .A4(_u10_u3_n2450 ), .ZN(_u10_u3_n2390 ) );
NAND2_X1 _u10_u3_U331  ( .A1(_u10_u3_n2445 ), .A2(_u10_u3_n2446 ), .ZN(_u10_u3_n2155 ) );
INV_X1 _u10_u3_U330  ( .A(_u10_u3_n2155 ), .ZN(_u10_u3_n1892 ) );
INV_X1 _u10_u3_U329  ( .A(_u10_u3_n2444 ), .ZN(_u10_u3_n2088 ) );
NAND2_X1 _u10_u3_U328  ( .A1(_u10_u3_n1892 ), .A2(_u10_u3_n2088 ), .ZN(_u10_u3_n2337 ) );
NOR3_X1 _u10_u3_U327  ( .A1(_u10_u3_n2441 ), .A2(_u10_u3_n2442 ), .A3(_u10_u3_n2443 ), .ZN(_u10_u3_n2440 ) );
NAND4_X1 _u10_u3_U326  ( .A1(_u10_u3_n2193 ), .A2(_u10_u3_n2355 ), .A3(_u10_u3_n2439 ), .A4(_u10_u3_n2440 ), .ZN(_u10_u3_n2434 ) );
NAND3_X1 _u10_u3_U325  ( .A1(_u10_u3_n2437 ), .A2(_u10_u3_n2438 ), .A3(_u10_u3_n2059 ), .ZN(_u10_u3_n2435 ) );
NOR4_X1 _u10_u3_U324  ( .A1(_u10_u3_n2434 ), .A2(_u10_u3_n2435 ), .A3(_u10_u3_n1837 ), .A4(_u10_u3_n2436 ), .ZN(_u10_u3_n2433 ) );
NOR2_X1 _u10_u3_U323  ( .A1(_u10_u3_n2433 ), .A2(_u10_u3_n1836 ), .ZN(_u10_u3_n2415 ) );
INV_X1 _u10_u3_U322  ( .A(_u10_u3_n2432 ), .ZN(_u10_u3_n2178 ) );
NOR2_X1 _u10_u3_U321  ( .A1(_u10_u3_n1960 ), .A2(_u10_u3_n2431 ), .ZN(_u10_u3_n2430 ) );
NOR4_X1 _u10_u3_U320  ( .A1(_u10_u3_n2178 ), .A2(_u10_u3_n2429 ), .A3(_u10_u3_n2430 ), .A4(_u10_u3_n2179 ), .ZN(_u10_u3_n2416 ) );
NOR2_X1 _u10_u3_U319  ( .A1(_u10_u3_n2427 ), .A2(_u10_u3_n2428 ), .ZN(_u10_u3_n2426 ) );
NAND4_X1 _u10_u3_U318  ( .A1(_u10_u3_n2286 ), .A2(_u10_u3_n1969 ), .A3(_u10_u3_n2282 ), .A4(_u10_u3_n2426 ), .ZN(_u10_u3_n2425 ) );
NAND2_X1 _u10_u3_U317  ( .A1(_u10_u3_n2031 ), .A2(_u10_u3_n2425 ), .ZN(_u10_u3_n2422 ) );
NAND3_X1 _u10_u3_U316  ( .A1(_u10_u3_n2422 ), .A2(_u10_u3_n2423 ), .A3(_u10_u3_n2424 ), .ZN(_u10_u3_n2419 ) );
NOR4_X1 _u10_u3_U315  ( .A1(_u10_u3_n2419 ), .A2(_u10_u3_n1978 ), .A3(_u10_u3_n2420 ), .A4(_u10_u3_n2421 ), .ZN(_u10_u3_n2418 ) );
NOR2_X1 _u10_u3_U314  ( .A1(_u10_u3_n2418 ), .A2(_u10_u3_n2359 ), .ZN(_u10_u3_n2417 ) );
NOR3_X1 _u10_u3_U313  ( .A1(_u10_u3_n2415 ), .A2(_u10_u3_n2416 ), .A3(_u10_u3_n2417 ), .ZN(_u10_u3_n2414 ) );
NAND4_X1 _u10_u3_U312  ( .A1(_u10_u3_n2337 ), .A2(_u10_u3_n2412 ), .A3(_u10_u3_n2413 ), .A4(_u10_u3_n2414 ), .ZN(_u10_u3_n2392 ) );
NAND2_X1 _u10_u3_U311  ( .A1(_u10_u3_n2411 ), .A2(_u10_u3_n1936 ), .ZN(_u10_u3_n2410 ) );
NAND2_X1 _u10_u3_U310  ( .A1(_u10_u3_n2409 ), .A2(_u10_u3_n2410 ), .ZN(_u10_u3_n2408 ) );
NAND3_X1 _u10_u3_U309  ( .A1(_u10_u3_n2408 ), .A2(_u10_u3_n2305 ), .A3(_u10_u3_n1894 ), .ZN(_u10_u3_n2402 ) );
NAND3_X1 _u10_u3_U308  ( .A1(_u10_u3_n2329 ), .A2(_u10_u3_n2407 ), .A3(_u10_u3_n2255 ), .ZN(_u10_u3_n2403 ) );
NAND3_X1 _u10_u3_U307  ( .A1(_u10_u3_n1924 ), .A2(_u10_u3_n2405 ), .A3(_u10_u3_n2406 ), .ZN(_u10_u3_n2404 ) );
NAND3_X1 _u10_u3_U306  ( .A1(_u10_u3_n2402 ), .A2(_u10_u3_n2403 ), .A3(_u10_u3_n2404 ), .ZN(_u10_u3_n2393 ) );
INV_X1 _u10_u3_U305  ( .A(_u10_u3_n1932 ), .ZN(_u10_u3_n2399 ) );
NOR2_X1 _u10_u3_U304  ( .A1(_u10_u3_n2401 ), .A2(_u10_u3_n2161 ), .ZN(_u10_u3_n2400 ) );
NOR2_X1 _u10_u3_U303  ( .A1(_u10_u3_n2399 ), .A2(_u10_u3_n2400 ), .ZN(_u10_u3_n2394 ) );
NOR2_X1 _u10_u3_U302  ( .A1(_u10_u3_n2110 ), .A2(_u10_u3_n2398 ), .ZN(_u10_u3_n2397 ) );
NOR2_X1 _u10_u3_U301  ( .A1(_u10_u3_n2396 ), .A2(_u10_u3_n2397 ), .ZN(_u10_u3_n2395 ) );
NOR4_X1 _u10_u3_U300  ( .A1(_u10_u3_n2392 ), .A2(_u10_u3_n2393 ), .A3(_u10_u3_n2394 ), .A4(_u10_u3_n2395 ), .ZN(_u10_u3_n2391 ) );
NAND4_X1 _u10_u3_U299  ( .A1(_u10_u3_n2388 ), .A2(_u10_u3_n2389 ), .A3(_u10_u3_n2390 ), .A4(_u10_u3_n2391 ), .ZN(_u10_u3_n2387 ) );
MUX2_X1 _u10_u3_U298  ( .A(_u10_u3_n2387 ), .B(_u10_SYNOPSYS_UNCONNECTED_10 ), .S(_u10_u3_n1819 ), .Z(_u10_u3_n1810 ) );
NAND2_X1 _u10_u3_U297  ( .A1(_u10_u3_n2386 ), .A2(_u10_u3_n2007 ), .ZN(_u10_u3_n2369 ) );
AND2_X1 _u10_u3_U296  ( .A1(1'b0), .A2(_u10_u3_n2195 ), .ZN(_u10_u3_n2308 ));
NAND2_X1 _u10_u3_U295  ( .A1(_u10_u3_n2308 ), .A2(_u10_u3_n2036 ), .ZN(_u10_u3_n2384 ) );
AND2_X1 _u10_u3_U294  ( .A1(_u10_u3_n2384 ), .A2(_u10_u3_n2385 ), .ZN(_u10_u3_n2275 ) );
AND4_X1 _u10_u3_U293  ( .A1(_u10_u3_n2275 ), .A2(_u10_u3_n2286 ), .A3(_u10_u3_n2383 ), .A4(_u10_u3_n2285 ), .ZN(_u10_u3_n2225 ) );
NAND3_X1 _u10_u3_U292  ( .A1(_u10_u3_n2195 ), .A2(_u10_u3_n2223 ), .A3(1'b0),.ZN(_u10_u3_n2021 ) );
INV_X1 _u10_u3_U291  ( .A(_u10_u3_n2021 ), .ZN(_u10_u3_n2167 ) );
NAND2_X1 _u10_u3_U290  ( .A1(_u10_u3_n2036 ), .A2(_u10_u3_n2167 ), .ZN(_u10_u3_n1970 ) );
AND3_X1 _u10_u3_U289  ( .A1(_u10_u3_n1970 ), .A2(_u10_u3_n2164 ), .A3(_u10_u3_n2382 ), .ZN(_u10_u3_n2381 ) );
NAND4_X1 _u10_u3_U288  ( .A1(_u10_u3_n2225 ), .A2(_u10_u3_n2379 ), .A3(_u10_u3_n2380 ), .A4(_u10_u3_n2381 ), .ZN(_u10_u3_n2378 ) );
NAND2_X1 _u10_u3_U287  ( .A1(_u10_u3_n1967 ), .A2(_u10_u3_n2378 ), .ZN(_u10_u3_n2370 ) );
NAND2_X1 _u10_u3_U286  ( .A1(_u10_u3_n2081 ), .A2(_u10_u3_n2377 ), .ZN(_u10_u3_n2371 ) );
NOR2_X1 _u10_u3_U285  ( .A1(_u10_u3_n2375 ), .A2(_u10_u3_n2376 ), .ZN(_u10_u3_n2373 ) );
NOR2_X1 _u10_u3_U284  ( .A1(_u10_u3_n2373 ), .A2(_u10_u3_n2374 ), .ZN(_u10_u3_n2372 ) );
NAND4_X1 _u10_u3_U283  ( .A1(_u10_u3_n2369 ), .A2(_u10_u3_n2370 ), .A3(_u10_u3_n2371 ), .A4(_u10_u3_n2372 ), .ZN(_u10_u3_n2309 ) );
NOR2_X1 _u10_u3_U282  ( .A1(_u10_u3_n2000 ), .A2(_u10_u3_n2368 ), .ZN(_u10_u3_n2360 ) );
NOR2_X1 _u10_u3_U281  ( .A1(_u10_u3_n2366 ), .A2(_u10_u3_n2367 ), .ZN(_u10_u3_n2361 ) );
NOR2_X1 _u10_u3_U280  ( .A1(_u10_u3_n1868 ), .A2(_u10_u3_n2365 ), .ZN(_u10_u3_n2362 ) );
NOR2_X1 _u10_u3_U279  ( .A1(_u10_u3_n2364 ), .A2(_u10_u3_n1859 ), .ZN(_u10_u3_n2363 ) );
NOR4_X1 _u10_u3_U278  ( .A1(_u10_u3_n2360 ), .A2(_u10_u3_n2361 ), .A3(_u10_u3_n2362 ), .A4(_u10_u3_n2363 ), .ZN(_u10_u3_n2316 ) );
NOR2_X1 _u10_u3_U277  ( .A1(_u10_u3_n2359 ), .A2(_u10_u3_n1970 ), .ZN(_u10_u3_n2351 ) );
NOR2_X1 _u10_u3_U276  ( .A1(_u10_u3_n2358 ), .A2(_u10_u3_n1840 ), .ZN(_u10_u3_n2352 ) );
NOR2_X1 _u10_u3_U275  ( .A1(_u10_u3_n2356 ), .A2(_u10_u3_n2357 ), .ZN(_u10_u3_n2353 ) );
NOR2_X1 _u10_u3_U274  ( .A1(_u10_u3_n1836 ), .A2(_u10_u3_n2355 ), .ZN(_u10_u3_n2354 ) );
NOR4_X1 _u10_u3_U273  ( .A1(_u10_u3_n2351 ), .A2(_u10_u3_n2352 ), .A3(_u10_u3_n2353 ), .A4(_u10_u3_n2354 ), .ZN(_u10_u3_n2317 ) );
NOR2_X1 _u10_u3_U272  ( .A1(_u10_u3_n1873 ), .A2(_u10_u3_n2101 ), .ZN(_u10_u3_n2349 ) );
NOR2_X1 _u10_u3_U271  ( .A1(_u10_u3_n2349 ), .A2(_u10_u3_n2350 ), .ZN(_u10_u3_n2338 ) );
NOR2_X1 _u10_u3_U270  ( .A1(_u10_u3_n2347 ), .A2(_u10_u3_n2348 ), .ZN(_u10_u3_n2345 ) );
NOR2_X1 _u10_u3_U269  ( .A1(_u10_u3_n2345 ), .A2(_u10_u3_n2346 ), .ZN(_u10_u3_n2339 ) );
NOR2_X1 _u10_u3_U268  ( .A1(_u10_u3_n2344 ), .A2(_u10_u3_n2142 ), .ZN(_u10_u3_n2340 ) );
NOR2_X1 _u10_u3_U267  ( .A1(_u10_u3_n2342 ), .A2(_u10_u3_n2343 ), .ZN(_u10_u3_n2341 ) );
NOR4_X1 _u10_u3_U266  ( .A1(_u10_u3_n2338 ), .A2(_u10_u3_n2339 ), .A3(_u10_u3_n2340 ), .A4(_u10_u3_n2341 ), .ZN(_u10_u3_n2318 ) );
INV_X1 _u10_u3_U265  ( .A(_u10_u3_n2337 ), .ZN(_u10_u3_n2320 ) );
NOR2_X1 _u10_u3_U264  ( .A1(_u10_u3_n1970 ), .A2(1'b0), .ZN(_u10_u3_n2027 ));
INV_X1 _u10_u3_U263  ( .A(_u10_u3_n2027 ), .ZN(_u10_u3_n2331 ) );
NOR2_X1 _u10_u3_U262  ( .A1(_u10_u3_n2174 ), .A2(_u10_u3_n2216 ), .ZN(_u10_u3_n2333 ) );
AND2_X1 _u10_u3_U261  ( .A1(_u10_u3_n1928 ), .A2(_u10_u3_n2336 ), .ZN(_u10_u3_n2334 ) );
NOR4_X1 _u10_u3_U260  ( .A1(_u10_u3_n1937 ), .A2(_u10_u3_n2333 ), .A3(_u10_u3_n2334 ), .A4(_u10_u3_n2335 ), .ZN(_u10_u3_n2332 ) );
NOR3_X1 _u10_u3_U259  ( .A1(_u10_u3_n2331 ), .A2(_u10_u3_n2332 ), .A3(_u10_u3_n1915 ), .ZN(_u10_u3_n2321 ) );
NOR3_X1 _u10_u3_U258  ( .A1(_u10_u3_n2291 ), .A2(_u10_u3_n2330 ), .A3(_u10_u3_n2021 ), .ZN(_u10_u3_n2322 ) );
NOR2_X1 _u10_u3_U257  ( .A1(_u10_u3_n2329 ), .A2(_u10_u3_n2169 ), .ZN(_u10_u3_n2324 ) );
NOR2_X1 _u10_u3_U256  ( .A1(1'b0), .A2(_u10_u3_n2328 ), .ZN(_u10_u3_n2327 ));
NOR2_X1 _u10_u3_U255  ( .A1(_u10_u3_n2326 ), .A2(_u10_u3_n2327 ), .ZN(_u10_u3_n2325 ) );
NOR3_X1 _u10_u3_U254  ( .A1(_u10_u3_n2324 ), .A2(1'b0), .A3(_u10_u3_n2325 ),.ZN(_u10_u3_n2323 ) );
NOR4_X1 _u10_u3_U253  ( .A1(_u10_u3_n2320 ), .A2(_u10_u3_n2321 ), .A3(_u10_u3_n2322 ), .A4(_u10_u3_n2323 ), .ZN(_u10_u3_n2319 ) );
AND4_X1 _u10_u3_U252  ( .A1(_u10_u3_n2316 ), .A2(_u10_u3_n2317 ), .A3(_u10_u3_n2318 ), .A4(_u10_u3_n2319 ), .ZN(_u10_u3_n1991 ) );
INV_X1 _u10_u3_U251  ( .A(_u10_u3_n2315 ), .ZN(_u10_u3_n2313 ) );
NAND3_X1 _u10_u3_U250  ( .A1(_u10_u3_n1991 ), .A2(_u10_u3_n2313 ), .A3(_u10_u3_n2314 ), .ZN(_u10_u3_n2310 ) );
NOR4_X1 _u10_u3_U249  ( .A1(_u10_u3_n2309 ), .A2(_u10_u3_n2310 ), .A3(_u10_u3_n2311 ), .A4(_u10_u3_n2312 ), .ZN(_u10_u3_n2117 ) );
NAND3_X1 _u10_u3_U248  ( .A1(_u10_u3_n2108 ), .A2(_u10_u3_n2107 ), .A3(_u10_u3_n2308 ), .ZN(_u10_u3_n2217 ) );
NOR3_X1 _u10_u3_U247  ( .A1(_u10_u3_n2306 ), .A2(_u10_u3_n2307 ), .A3(_u10_u3_n2027 ), .ZN(_u10_u3_n2277 ) );
NAND3_X1 _u10_u3_U246  ( .A1(_u10_u3_n2217 ), .A2(_u10_u3_n2305 ), .A3(_u10_u3_n2277 ), .ZN(_u10_u3_n2157 ) );
NAND2_X1 _u10_u3_U245  ( .A1(_u10_u3_n2089 ), .A2(_u10_u3_n2157 ), .ZN(_u10_u3_n2296 ) );
INV_X1 _u10_u3_U244  ( .A(_u10_u3_n2304 ), .ZN(_u10_u3_n2297 ) );
NOR2_X1 _u10_u3_U243  ( .A1(_u10_u3_n2302 ), .A2(_u10_u3_n2303 ), .ZN(_u10_u3_n2299 ) );
NOR3_X1 _u10_u3_U242  ( .A1(_u10_u3_n2299 ), .A2(_u10_u3_n2300 ), .A3(_u10_u3_n2301 ), .ZN(_u10_u3_n2298 ) );
NAND4_X1 _u10_u3_U241  ( .A1(_u10_u3_n2295 ), .A2(_u10_u3_n2296 ), .A3(_u10_u3_n2297 ), .A4(_u10_u3_n2298 ), .ZN(_u10_u3_n2294 ) );
NAND2_X1 _u10_u3_U240  ( .A1(_u10_u3_n2293 ), .A2(_u10_u3_n2294 ), .ZN(_u10_u3_n2257 ) );
NAND2_X1 _u10_u3_U239  ( .A1(_u10_u3_n2165 ), .A2(_u10_u3_n2166 ), .ZN(_u10_u3_n2288 ) );
NAND2_X1 _u10_u3_U238  ( .A1(_u10_u3_n2078 ), .A2(_u10_u3_n2279 ), .ZN(_u10_u3_n2292 ) );
NAND2_X1 _u10_u3_U237  ( .A1(_u10_u3_n2291 ), .A2(_u10_u3_n2292 ), .ZN(_u10_u3_n2290 ) );
NAND2_X1 _u10_u3_U236  ( .A1(_u10_u3_n2059 ), .A2(_u10_u3_n2290 ), .ZN(_u10_u3_n2289 ) );
NAND2_X1 _u10_u3_U235  ( .A1(_u10_u3_n2288 ), .A2(_u10_u3_n2289 ), .ZN(_u10_u3_n2201 ) );
NAND2_X1 _u10_u3_U234  ( .A1(1'b0), .A2(_u10_u3_n2201 ), .ZN(_u10_u3_n2258 ));
INV_X1 _u10_u3_U233  ( .A(_u10_u3_n2287 ), .ZN(_u10_u3_n2283 ) );
AND4_X1 _u10_u3_U232  ( .A1(_u10_u3_n2285 ), .A2(_u10_u3_n2226 ), .A3(_u10_u3_n1970 ), .A4(_u10_u3_n2286 ), .ZN(_u10_u3_n2284 ) );
NAND4_X1 _u10_u3_U231  ( .A1(_u10_u3_n2281 ), .A2(_u10_u3_n2282 ), .A3(_u10_u3_n2283 ), .A4(_u10_u3_n2284 ), .ZN(_u10_u3_n2280 ) );
NAND2_X1 _u10_u3_U230  ( .A1(_u10_u3_n2279 ), .A2(_u10_u3_n2280 ), .ZN(_u10_u3_n2259 ) );
NAND4_X1 _u10_u3_U229  ( .A1(_u10_u3_n2275 ), .A2(_u10_u3_n2276 ), .A3(_u10_u3_n2277 ), .A4(_u10_u3_n2278 ), .ZN(_u10_u3_n2271 ) );
NAND2_X1 _u10_u3_U228  ( .A1(_u10_u3_n1933 ), .A2(_u10_u3_n2164 ), .ZN(_u10_u3_n2272 ) );
NOR2_X1 _u10_u3_U227  ( .A1(_u10_u3_n2274 ), .A2(_u10_u3_n2130 ), .ZN(_u10_u3_n2273 ) );
NOR4_X1 _u10_u3_U226  ( .A1(_u10_u3_n2271 ), .A2(_u10_u3_n2272 ), .A3(_u10_u3_n1978 ), .A4(_u10_u3_n2273 ), .ZN(_u10_u3_n2270 ) );
NOR2_X1 _u10_u3_U225  ( .A1(_u10_u3_n2270 ), .A2(_u10_u3_n2025 ), .ZN(_u10_u3_n2261 ) );
NAND3_X1 _u10_u3_U224  ( .A1(_u10_u3_n1933 ), .A2(_u10_u3_n1936 ), .A3(_u10_u3_n2269 ), .ZN(_u10_u3_n2268 ) );
NOR3_X1 _u10_u3_U223  ( .A1(_u10_u3_n2268 ), .A2(_u10_u3_n1844 ), .A3(_u10_u3_n2157 ), .ZN(_u10_u3_n2267 ) );
NOR2_X1 _u10_u3_U222  ( .A1(1'b0), .A2(_u10_u3_n2267 ), .ZN(_u10_u3_n2265 ));
NOR3_X1 _u10_u3_U221  ( .A1(_u10_u3_n2264 ), .A2(_u10_u3_n2265 ), .A3(_u10_u3_n2266 ), .ZN(_u10_u3_n2263 ) );
NOR2_X1 _u10_u3_U220  ( .A1(_u10_u3_n2263 ), .A2(_u10_u3_n1843 ), .ZN(_u10_u3_n2262 ) );
NOR2_X1 _u10_u3_U219  ( .A1(_u10_u3_n2261 ), .A2(_u10_u3_n2262 ), .ZN(_u10_u3_n2260 ) );
NAND4_X1 _u10_u3_U218  ( .A1(_u10_u3_n2257 ), .A2(_u10_u3_n2258 ), .A3(_u10_u3_n2259 ), .A4(_u10_u3_n2260 ), .ZN(_u10_u3_n2230 ) );
INV_X1 _u10_u3_U217  ( .A(_u10_u3_n2217 ), .ZN(_u10_u3_n2242 ) );
NAND2_X1 _u10_u3_U216  ( .A1(_u10_u3_n2168 ), .A2(_u10_u3_n2169 ), .ZN(_u10_u3_n2244 ) );
NAND2_X1 _u10_u3_U215  ( .A1(_u10_u3_n2255 ), .A2(_u10_u3_n2256 ), .ZN(_u10_u3_n2245 ) );
NAND2_X1 _u10_u3_U214  ( .A1(_u10_u3_n2253 ), .A2(_u10_u3_n2254 ), .ZN(_u10_u3_n2252 ) );
NAND2_X1 _u10_u3_U213  ( .A1(_u10_u3_n2251 ), .A2(_u10_u3_n2252 ), .ZN(_u10_u3_n2246 ) );
NAND2_X1 _u10_u3_U212  ( .A1(_u10_u3_n2152 ), .A2(_u10_u3_n1928 ), .ZN(_u10_u3_n2250 ) );
NAND2_X1 _u10_u3_U211  ( .A1(_u10_u3_n2249 ), .A2(_u10_u3_n2250 ), .ZN(_u10_u3_n2248 ) );
NAND2_X1 _u10_u3_U210  ( .A1(_u10_u3_n2105 ), .A2(_u10_u3_n2248 ), .ZN(_u10_u3_n2247 ) );
NAND4_X1 _u10_u3_U209  ( .A1(_u10_u3_n2244 ), .A2(_u10_u3_n2245 ), .A3(_u10_u3_n2246 ), .A4(_u10_u3_n2247 ), .ZN(_u10_u3_n2243 ) );
NAND2_X1 _u10_u3_U208  ( .A1(_u10_u3_n2242 ), .A2(_u10_u3_n2243 ), .ZN(_u10_u3_n2237 ) );
NAND2_X1 _u10_u3_U207  ( .A1(1'b0), .A2(_u10_u3_n2241 ), .ZN(_u10_u3_n2238 ));
NAND2_X1 _u10_u3_U206  ( .A1(_u10_u3_n2214 ), .A2(_u10_u3_n2240 ), .ZN(_u10_u3_n2239 ) );
NAND3_X1 _u10_u3_U205  ( .A1(_u10_u3_n2237 ), .A2(_u10_u3_n2238 ), .A3(_u10_u3_n2239 ), .ZN(_u10_u3_n2231 ) );
AND2_X1 _u10_u3_U204  ( .A1(_u10_u3_n2200 ), .A2(_u10_u3_n2236 ), .ZN(_u10_u3_n2232 ) );
NOR2_X1 _u10_u3_U203  ( .A1(_u10_u3_n2234 ), .A2(_u10_u3_n2235 ), .ZN(_u10_u3_n2233 ) );
NOR4_X1 _u10_u3_U202  ( .A1(_u10_u3_n2230 ), .A2(_u10_u3_n2231 ), .A3(_u10_u3_n2232 ), .A4(_u10_u3_n2233 ), .ZN(_u10_u3_n2118 ) );
NAND2_X1 _u10_u3_U201  ( .A1(_u10_u3_n2214 ), .A2(_u10_u3_n2049 ), .ZN(_u10_u3_n2229 ) );
NAND2_X1 _u10_u3_U200  ( .A1(_u10_u3_n2228 ), .A2(_u10_u3_n2229 ), .ZN(_u10_u3_n2227 ) );
NAND2_X1 _u10_u3_U199  ( .A1(_u10_u3_n2043 ), .A2(_u10_u3_n2227 ), .ZN(_u10_u3_n2204 ) );
NAND2_X1 _u10_u3_U198  ( .A1(_u10_u3_n2225 ), .A2(_u10_u3_n2226 ), .ZN(_u10_u3_n2224 ) );
NAND2_X1 _u10_u3_U197  ( .A1(_u10_u3_n1899 ), .A2(_u10_u3_n2224 ), .ZN(_u10_u3_n2205 ) );
NAND2_X1 _u10_u3_U196  ( .A1(_u10_u3_n2222 ), .A2(_u10_u3_n2223 ), .ZN(_u10_u3_n1870 ) );
NAND4_X1 _u10_u3_U195  ( .A1(_u10_u3_n2220 ), .A2(_u10_u3_n2131 ), .A3(_u10_u3_n2221 ), .A4(_u10_u3_n1870 ), .ZN(_u10_u3_n2219 ) );
NAND2_X1 _u10_u3_U194  ( .A1(_u10_u3_n2218 ), .A2(_u10_u3_n2219 ), .ZN(_u10_u3_n2206 ) );
NOR2_X1 _u10_u3_U193  ( .A1(_u10_u3_n1925 ), .A2(_u10_u3_n2217 ), .ZN(_u10_u3_n2215 ) );
NOR4_X1 _u10_u3_U192  ( .A1(_u10_u3_n2213 ), .A2(_u10_u3_n2214 ), .A3(_u10_u3_n2215 ), .A4(_u10_u3_n2216 ), .ZN(_u10_u3_n2211 ) );
NOR2_X1 _u10_u3_U191  ( .A1(_u10_u3_n2211 ), .A2(_u10_u3_n2212 ), .ZN(_u10_u3_n2208 ) );
NOR2_X1 _u10_u3_U190  ( .A1(_u10_u3_n1888 ), .A2(_u10_u3_n2210 ), .ZN(_u10_u3_n2209 ) );
NOR2_X1 _u10_u3_U189  ( .A1(_u10_u3_n2208 ), .A2(_u10_u3_n2209 ), .ZN(_u10_u3_n2207 ) );
NAND4_X1 _u10_u3_U188  ( .A1(_u10_u3_n2204 ), .A2(_u10_u3_n2205 ), .A3(_u10_u3_n2206 ), .A4(_u10_u3_n2207 ), .ZN(_u10_u3_n2170 ) );
OR2_X1 _u10_u3_U187  ( .A1(_u10_u3_n2202 ), .A2(_u10_u3_n2203 ), .ZN(_u10_u3_n2197 ) );
NAND2_X1 _u10_u3_U186  ( .A1(1'b0), .A2(_u10_u3_n2201 ), .ZN(_u10_u3_n2198 ));
NAND2_X1 _u10_u3_U185  ( .A1(_u10_u3_n2063 ), .A2(_u10_u3_n2200 ), .ZN(_u10_u3_n2199 ) );
NAND3_X1 _u10_u3_U184  ( .A1(_u10_u3_n2197 ), .A2(_u10_u3_n2198 ), .A3(_u10_u3_n2199 ), .ZN(_u10_u3_n2196 ) );
NAND2_X1 _u10_u3_U183  ( .A1(_u10_u3_n2195 ), .A2(_u10_u3_n2196 ), .ZN(_u10_u3_n2180 ) );
NAND2_X1 _u10_u3_U182  ( .A1(_u10_u3_n2195 ), .A2(_u10_u3_n1918 ), .ZN(_u10_u3_n2192 ) );
NAND4_X1 _u10_u3_U181  ( .A1(_u10_u3_n2192 ), .A2(_u10_u3_n2021 ), .A3(_u10_u3_n2193 ), .A4(_u10_u3_n2194 ), .ZN(_u10_u3_n2188 ) );
NAND2_X1 _u10_u3_U180  ( .A1(_u10_u3_n2188 ), .A2(_u10_u3_n2191 ), .ZN(_u10_u3_n2181 ) );
NAND2_X1 _u10_u3_U179  ( .A1(1'b0), .A2(_u10_u3_n2190 ), .ZN(_u10_u3_n2185 ));
NAND2_X1 _u10_u3_U178  ( .A1(_u10_u3_n2189 ), .A2(_u10_SYNOPSYS_UNCONNECTED_11 ), .ZN(_u10_u3_n2186 ) );
INV_X1 _u10_u3_U177  ( .A(_u10_u3_n2188 ), .ZN(_u10_u3_n2187 ) );
NAND3_X1 _u10_u3_U176  ( .A1(_u10_u3_n2185 ), .A2(_u10_u3_n2186 ), .A3(_u10_u3_n2187 ), .ZN(_u10_u3_n2184 ) );
NAND2_X1 _u10_u3_U175  ( .A1(_u10_u3_n2183 ), .A2(_u10_u3_n2184 ), .ZN(_u10_u3_n2182 ) );
NAND3_X1 _u10_u3_U174  ( .A1(_u10_u3_n2180 ), .A2(_u10_u3_n2181 ), .A3(_u10_u3_n2182 ), .ZN(_u10_u3_n2171 ) );
INV_X1 _u10_u3_U173  ( .A(_u10_u3_n2179 ), .ZN(_u10_u3_n1963 ) );
NOR2_X1 _u10_u3_U172  ( .A1(_u10_u3_n1963 ), .A2(_u10_u3_n2178 ), .ZN(_u10_u3_n2172 ) );
INV_X1 _u10_u3_U171  ( .A(_u10_u3_n2177 ), .ZN(_u10_u3_n2176 ) );
NOR3_X1 _u10_u3_U170  ( .A1(_u10_u3_n2174 ), .A2(_u10_u3_n2175 ), .A3(_u10_u3_n2176 ), .ZN(_u10_u3_n2173 ) );
NOR4_X1 _u10_u3_U169  ( .A1(_u10_u3_n2170 ), .A2(_u10_u3_n2171 ), .A3(_u10_u3_n2172 ), .A4(_u10_u3_n2173 ), .ZN(_u10_u3_n2119 ) );
NAND3_X1 _u10_u3_U168  ( .A1(_u10_u3_n2168 ), .A2(_u10_u3_n2169 ), .A3(1'b0),.ZN(_u10_u3_n2148 ) );
NAND3_X1 _u10_u3_U167  ( .A1(_u10_u3_n2165 ), .A2(_u10_u3_n2166 ), .A3(_u10_u3_n2167 ), .ZN(_u10_u3_n2149 ) );
NAND4_X1 _u10_u3_U166  ( .A1(_u10_u3_n2162 ), .A2(_u10_u3_n1933 ), .A3(_u10_u3_n2163 ), .A4(_u10_u3_n2164 ), .ZN(_u10_u3_n2160 ) );
NOR4_X1 _u10_u3_U165  ( .A1(_u10_u3_n2160 ), .A2(_u10_u3_n2157 ), .A3(_u10_u3_n1844 ), .A4(_u10_u3_n2161 ), .ZN(_u10_u3_n2158 ) );
NOR2_X1 _u10_u3_U164  ( .A1(_u10_u3_n2158 ), .A2(_u10_u3_n2159 ), .ZN(_u10_u3_n2153 ) );
INV_X1 _u10_u3_U163  ( .A(_u10_u3_n2157 ), .ZN(_u10_u3_n2129 ) );
NOR3_X1 _u10_u3_U162  ( .A1(_u10_u3_n2155 ), .A2(_u10_u3_n2129 ), .A3(_u10_u3_n2156 ), .ZN(_u10_u3_n2154 ) );
NOR2_X1 _u10_u3_U161  ( .A1(_u10_u3_n2153 ), .A2(_u10_u3_n2154 ), .ZN(_u10_u3_n2150 ) );
NAND3_X1 _u10_u3_U160  ( .A1(1'b0), .A2(_u10_u3_n1928 ), .A3(_u10_u3_n2152 ),.ZN(_u10_u3_n2151 ) );
NAND4_X1 _u10_u3_U159  ( .A1(_u10_u3_n2148 ), .A2(_u10_u3_n2149 ), .A3(_u10_u3_n2150 ), .A4(_u10_u3_n2151 ), .ZN(_u10_u3_n2121 ) );
NAND2_X1 _u10_u3_U158  ( .A1(_u10_u3_n2107 ), .A2(_u10_u3_n2147 ), .ZN(_u10_u3_n2146 ) );
NAND2_X1 _u10_u3_U157  ( .A1(_u10_u3_n2145 ), .A2(_u10_u3_n2146 ), .ZN(_u10_u3_n2144 ) );
NAND2_X1 _u10_u3_U156  ( .A1(_u10_u3_n2143 ), .A2(_u10_u3_n2144 ), .ZN(_u10_u3_n2134 ) );
NAND2_X1 _u10_u3_U155  ( .A1(_u10_u3_n2141 ), .A2(_u10_u3_n2142 ), .ZN(_u10_u3_n2140 ) );
NAND2_X1 _u10_u3_U154  ( .A1(_u10_u3_n2139 ), .A2(_u10_u3_n2140 ), .ZN(_u10_u3_n2135 ) );
OR2_X1 _u10_u3_U153  ( .A1(_u10_u3_n2110 ), .A2(_u10_u3_n1911 ), .ZN(_u10_u3_n2137 ) );
NAND2_X1 _u10_u3_U152  ( .A1(_u10_u3_n2137 ), .A2(_u10_u3_n2138 ), .ZN(_u10_u3_n2136 ) );
NAND3_X1 _u10_u3_U151  ( .A1(_u10_u3_n2134 ), .A2(_u10_u3_n2135 ), .A3(_u10_u3_n2136 ), .ZN(_u10_u3_n2122 ) );
NOR2_X1 _u10_u3_U150  ( .A1(_u10_u3_n2133 ), .A2(_u10_u3_n1891 ), .ZN(_u10_u3_n2132 ) );
NOR2_X1 _u10_u3_U149  ( .A1(_u10_u3_n2131 ), .A2(_u10_u3_n2132 ), .ZN(_u10_u3_n2123 ) );
NOR2_X1 _u10_u3_U148  ( .A1(_u10_u3_n2129 ), .A2(_u10_u3_n2130 ), .ZN(_u10_u3_n2127 ) );
NOR2_X1 _u10_u3_U147  ( .A1(_u10_u3_n2127 ), .A2(_u10_u3_n2128 ), .ZN(_u10_u3_n2125 ) );
NOR2_X1 _u10_u3_U146  ( .A1(_u10_u3_n2125 ), .A2(_u10_u3_n2126 ), .ZN(_u10_u3_n2124 ) );
NOR4_X1 _u10_u3_U145  ( .A1(_u10_u3_n2121 ), .A2(_u10_u3_n2122 ), .A3(_u10_u3_n2123 ), .A4(_u10_u3_n2124 ), .ZN(_u10_u3_n2120 ) );
NAND4_X1 _u10_u3_U144  ( .A1(_u10_u3_n2117 ), .A2(_u10_u3_n2118 ), .A3(_u10_u3_n2119 ), .A4(_u10_u3_n2120 ), .ZN(_u10_u3_n2116 ) );
MUX2_X1 _u10_u3_U143  ( .A(_u10_u3_n2116 ), .B(_u10_SYNOPSYS_UNCONNECTED_11 ), .S(_u10_u3_n1819 ), .Z(_u10_u3_n1811 ) );
INV_X1 _u10_u3_U142  ( .A(_u10_u3_n2115 ), .ZN(_u10_u3_n2006 ) );
NOR3_X1 _u10_u3_U141  ( .A1(_u10_u3_n2006 ), .A2(_u10_u3_n2114 ), .A3(_u10_u3_n2081 ), .ZN(_u10_u3_n1854 ) );
NAND2_X1 _u10_u3_U140  ( .A1(_u10_u3_n2112 ), .A2(_u10_u3_n2113 ), .ZN(_u10_u3_n1872 ) );
INV_X1 _u10_u3_U139  ( .A(_u10_u3_n1872 ), .ZN(_u10_u3_n1882 ) );
NAND4_X1 _u10_u3_U138  ( .A1(_u10_u3_n1854 ), .A2(_u10_u3_n1882 ), .A3(_u10_u3_n2111 ), .A4(_u10_u3_n1868 ), .ZN(_u10_u3_n2109 ) );
NAND2_X1 _u10_u3_U137  ( .A1(_u10_u3_n2109 ), .A2(_u10_u3_n2110 ), .ZN(_u10_u3_n2098 ) );
NAND2_X1 _u10_u3_U136  ( .A1(1'b0), .A2(_u10_u3_n1983 ), .ZN(_u10_u3_n2023 ));
INV_X1 _u10_u3_U135  ( .A(_u10_u3_n2023 ), .ZN(_u10_u3_n2035 ) );
NAND3_X1 _u10_u3_U134  ( .A1(_u10_u3_n2035 ), .A2(_u10_u3_n2107 ), .A3(_u10_u3_n2108 ), .ZN(_u10_u3_n1916 ) );
INV_X1 _u10_u3_U133  ( .A(_u10_u3_n1916 ), .ZN(_u10_u3_n2093 ) );
NAND3_X1 _u10_u3_U132  ( .A1(_u10_u3_n2105 ), .A2(_u10_u3_n2106 ), .A3(_u10_u3_n2093 ), .ZN(_u10_u3_n2039 ) );
NAND2_X1 _u10_u3_U131  ( .A1(_u10_u3_n2039 ), .A2(_u10_u3_n1930 ), .ZN(_u10_u3_n2104 ) );
NAND2_X1 _u10_u3_U130  ( .A1(_u10_u3_n2103 ), .A2(_u10_u3_n2104 ), .ZN(_u10_u3_n1863 ) );
OR2_X1 _u10_u3_U129  ( .A1(_u10_u3_n1863 ), .A2(_u10_u3_n2102 ), .ZN(_u10_u3_n2099 ) );
NAND2_X1 _u10_u3_U128  ( .A1(_u10_u3_n1890 ), .A2(_u10_u3_n2101 ), .ZN(_u10_u3_n2100 ) );
NAND3_X1 _u10_u3_U127  ( .A1(_u10_u3_n2098 ), .A2(_u10_u3_n2099 ), .A3(_u10_u3_n2100 ), .ZN(_u10_u3_n2066 ) );
NAND4_X1 _u10_u3_U126  ( .A1(_u10_u3_n2095 ), .A2(_u10_u3_n2096 ), .A3(_u10_u3_n1896 ), .A4(_u10_u3_n2097 ), .ZN(_u10_u3_n2086 ) );
NOR4_X1 _u10_u3_U125  ( .A1(_u10_u3_n2093 ), .A2(_u10_u3_n2027 ), .A3(_u10_u3_n2094 ), .A4(_u10_u3_n2026 ), .ZN(_u10_u3_n1952 ) );
NOR2_X1 _u10_u3_U124  ( .A1(1'b0), .A2(_u10_u3_n1952 ), .ZN(_u10_u3_n1951 ));
INV_X1 _u10_u3_U123  ( .A(_u10_u3_n1951 ), .ZN(_u10_u3_n2090 ) );
NAND4_X1 _u10_u3_U122  ( .A1(_u10_u3_n2089 ), .A2(_u10_u3_n2090 ), .A3(_u10_u3_n2091 ), .A4(_u10_u3_n2092 ), .ZN(_u10_u3_n1893 ) );
NOR4_X1 _u10_u3_U121  ( .A1(_u10_u3_n2086 ), .A2(_u10_u3_n1893 ), .A3(_u10_u3_n2087 ), .A4(_u10_u3_n2088 ), .ZN(_u10_u3_n2084 ) );
NOR2_X1 _u10_u3_U120  ( .A1(_u10_u3_n2084 ), .A2(_u10_u3_n2085 ), .ZN(_u10_u3_n2067 ) );
NOR2_X1 _u10_u3_U119  ( .A1(_u10_u3_n2083 ), .A2(_u10_u3_n1869 ), .ZN(_u10_u3_n2068 ) );
NAND2_X1 _u10_u3_U118  ( .A1(_u10_u3_n2081 ), .A2(_u10_u3_n2082 ), .ZN(_u10_u3_n2075 ) );
NAND2_X1 _u10_u3_U117  ( .A1(_u10_u3_n2035 ), .A2(_u10_u3_n2019 ), .ZN(_u10_u3_n2060 ) );
NAND2_X1 _u10_u3_U116  ( .A1(_u10_u3_n2080 ), .A2(_u10_u3_n2060 ), .ZN(_u10_u3_n2079 ) );
NAND2_X1 _u10_u3_U115  ( .A1(_u10_u3_n2078 ), .A2(_u10_u3_n2079 ), .ZN(_u10_u3_n2076 ) );
NAND4_X1 _u10_u3_U114  ( .A1(_u10_u3_n2075 ), .A2(_u10_u3_n2076 ), .A3(_u10_u3_n1970 ), .A4(_u10_u3_n2077 ), .ZN(_u10_u3_n2072 ) );
NOR4_X1 _u10_u3_U113  ( .A1(_u10_u3_n2072 ), .A2(_u10_u3_n2073 ), .A3(_u10_u3_n1975 ), .A4(_u10_u3_n2074 ), .ZN(_u10_u3_n2070 ) );
NOR2_X1 _u10_u3_U112  ( .A1(_u10_u3_n2070 ), .A2(_u10_u3_n2071 ), .ZN(_u10_u3_n2069 ) );
NOR4_X1 _u10_u3_U111  ( .A1(_u10_u3_n2066 ), .A2(_u10_u3_n2067 ), .A3(_u10_u3_n2068 ), .A4(_u10_u3_n2069 ), .ZN(_u10_u3_n1820 ) );
NAND2_X1 _u10_u3_U110  ( .A1(1'b0), .A2(_u10_u3_n1983 ), .ZN(_u10_u3_n2065 ));
NAND4_X1 _u10_u3_U109  ( .A1(_u10_u3_n2065 ), .A2(_u10_u3_n2023 ), .A3(_u10_u3_n2021 ), .A4(_u10_u3_n2052 ), .ZN(_u10_u3_n2064 ) );
NAND2_X1 _u10_u3_U108  ( .A1(_u10_u3_n2063 ), .A2(_u10_u3_n2064 ), .ZN(_u10_u3_n2040 ) );
NAND4_X1 _u10_u3_U107  ( .A1(_u10_u3_n2059 ), .A2(_u10_u3_n2060 ), .A3(_u10_u3_n2061 ), .A4(_u10_u3_n2062 ), .ZN(_u10_u3_n2058 ) );
NAND2_X1 _u10_u3_U106  ( .A1(_u10_u3_n2057 ), .A2(_u10_u3_n2058 ), .ZN(_u10_u3_n2041 ) );
NOR4_X1 _u10_u3_U105  ( .A1(1'b0), .A2(_u10_u3_n2054 ), .A3(_u10_u3_n2055 ),.A4(_u10_u3_n2056 ), .ZN(_u10_u3_n2053 ) );
NAND4_X1 _u10_u3_U104  ( .A1(_u10_u3_n2021 ), .A2(_u10_u3_n2052 ), .A3(_u10_u3_n2023 ), .A4(_u10_u3_n2053 ), .ZN(_u10_u3_n1964 ) );
INV_X1 _u10_u3_U103  ( .A(_u10_u3_n1964 ), .ZN(_u10_u3_n2045 ) );
NAND2_X1 _u10_u3_U102  ( .A1(_u10_u3_n2051 ), .A2(_u10_SYNOPSYS_UNCONNECTED_12 ), .ZN(_u10_u3_n2046 ) );
NAND2_X1 _u10_u3_U101  ( .A1(_u10_u3_n2049 ), .A2(_u10_u3_n2050 ), .ZN(_u10_u3_n2047 ) );
NAND4_X1 _u10_u3_U100  ( .A1(_u10_u3_n2045 ), .A2(_u10_u3_n2046 ), .A3(_u10_u3_n2047 ), .A4(_u10_u3_n2048 ), .ZN(_u10_u3_n2044 ) );
NAND2_X1 _u10_u3_U99  ( .A1(_u10_u3_n2043 ), .A2(_u10_u3_n2044 ), .ZN(_u10_u3_n2042 ) );
NAND3_X1 _u10_u3_U98  ( .A1(_u10_u3_n2040 ), .A2(_u10_u3_n2041 ), .A3(_u10_u3_n2042 ), .ZN(_u10_u3_n2009 ) );
AND2_X1 _u10_u3_U97  ( .A1(_u10_u3_n2038 ), .A2(_u10_u3_n2039 ), .ZN(_u10_u3_n1929 ) );
NOR2_X1 _u10_u3_U96  ( .A1(_u10_u3_n1929 ), .A2(_u10_u3_n2037 ), .ZN(_u10_u3_n2010 ) );
NAND2_X1 _u10_u3_U95  ( .A1(_u10_u3_n2035 ), .A2(_u10_u3_n2036 ), .ZN(_u10_u3_n1902 ) );
NAND3_X1 _u10_u3_U94  ( .A1(_u10_u3_n1902 ), .A2(_u10_u3_n2033 ), .A3(_u10_u3_n2034 ), .ZN(_u10_u3_n1973 ) );
NOR2_X1 _u10_u3_U93  ( .A1(_u10_u3_n1978 ), .A2(_u10_u3_n1973 ), .ZN(_u10_u3_n2032 ) );
NOR2_X1 _u10_u3_U92  ( .A1(1'b0), .A2(_u10_u3_n2032 ), .ZN(_u10_u3_n2028 ));
NOR2_X1 _u10_u3_U91  ( .A1(_u10_u3_n2030 ), .A2(_u10_u3_n2031 ), .ZN(_u10_u3_n2029 ) );
NOR4_X1 _u10_u3_U90  ( .A1(_u10_u3_n2026 ), .A2(_u10_u3_n2027 ), .A3(_u10_u3_n2028 ), .A4(_u10_u3_n2029 ), .ZN(_u10_u3_n2024 ) );
NOR2_X1 _u10_u3_U89  ( .A1(_u10_u3_n2024 ), .A2(_u10_u3_n2025 ), .ZN(_u10_u3_n2011 ) );
NAND3_X1 _u10_u3_U88  ( .A1(_u10_u3_n2021 ), .A2(_u10_u3_n2022 ), .A3(_u10_u3_n2023 ), .ZN(_u10_u3_n2020 ) );
AND2_X1 _u10_u3_U87  ( .A1(_u10_u3_n2019 ), .A2(_u10_u3_n2020 ), .ZN(_u10_u3_n1838 ) );
INV_X1 _u10_u3_U86  ( .A(_u10_u3_n2018 ), .ZN(_u10_u3_n2016 ) );
NOR4_X1 _u10_u3_U85  ( .A1(_u10_u3_n2015 ), .A2(_u10_u3_n1838 ), .A3(_u10_u3_n2016 ), .A4(_u10_u3_n2017 ), .ZN(_u10_u3_n2013 ) );
NOR2_X1 _u10_u3_U84  ( .A1(_u10_u3_n2013 ), .A2(_u10_u3_n2014 ), .ZN(_u10_u3_n2012 ) );
NOR4_X1 _u10_u3_U83  ( .A1(_u10_u3_n2009 ), .A2(_u10_u3_n2010 ), .A3(_u10_u3_n2011 ), .A4(_u10_u3_n2012 ), .ZN(_u10_u3_n1821 ) );
NAND2_X1 _u10_u3_U82  ( .A1(_u10_u3_n1924 ), .A2(_u10_u3_n2008 ), .ZN(_u10_u3_n1993 ) );
NAND2_X1 _u10_u3_U81  ( .A1(_u10_u3_n2006 ), .A2(_u10_u3_n2007 ), .ZN(_u10_u3_n1994 ) );
NAND2_X1 _u10_u3_U80  ( .A1(_u10_u3_n2004 ), .A2(_u10_u3_n2005 ), .ZN(_u10_u3_n1995 ) );
AND2_X1 _u10_u3_U79  ( .A1(_u10_u3_n2002 ), .A2(_u10_u3_n2003 ), .ZN(_u10_u3_n1998 ) );
NOR2_X1 _u10_u3_U78  ( .A1(_u10_u3_n2000 ), .A2(_u10_u3_n2001 ), .ZN(_u10_u3_n1999 ) );
NOR3_X1 _u10_u3_U77  ( .A1(_u10_u3_n1997 ), .A2(_u10_u3_n1998 ), .A3(_u10_u3_n1999 ), .ZN(_u10_u3_n1996 ) );
NAND4_X1 _u10_u3_U76  ( .A1(_u10_u3_n1993 ), .A2(_u10_u3_n1994 ), .A3(_u10_u3_n1995 ), .A4(_u10_u3_n1996 ), .ZN(_u10_u3_n1985 ) );
INV_X1 _u10_u3_U75  ( .A(_u10_u3_n1992 ), .ZN(_u10_u3_n1989 ) );
NAND3_X1 _u10_u3_U74  ( .A1(_u10_u3_n1989 ), .A2(_u10_u3_n1990 ), .A3(_u10_u3_n1991 ), .ZN(_u10_u3_n1986 ) );
NOR4_X1 _u10_u3_U73  ( .A1(_u10_u3_n1985 ), .A2(_u10_u3_n1986 ), .A3(_u10_u3_n1987 ), .A4(_u10_u3_n1988 ), .ZN(_u10_u3_n1822 ) );
INV_X1 _u10_u3_U72  ( .A(_u10_u3_n1984 ), .ZN(_u10_u3_n1980 ) );
NAND4_X1 _u10_u3_U71  ( .A1(_u10_u3_n1980 ), .A2(_u10_u3_n1981 ), .A3(_u10_u3_n1982 ), .A4(_u10_u3_n1983 ), .ZN(_u10_u3_n1941 ) );
NOR3_X1 _u10_u3_U70  ( .A1(_u10_u3_n1977 ), .A2(_u10_u3_n1978 ), .A3(_u10_u3_n1979 ), .ZN(_u10_u3_n1971 ) );
NOR4_X1 _u10_u3_U69  ( .A1(_u10_u3_n1973 ), .A2(_u10_u3_n1974 ), .A3(_u10_u3_n1975 ), .A4(_u10_u3_n1976 ), .ZN(_u10_u3_n1972 ) );
NAND4_X1 _u10_u3_U68  ( .A1(_u10_u3_n1969 ), .A2(_u10_u3_n1970 ), .A3(_u10_u3_n1971 ), .A4(_u10_u3_n1972 ), .ZN(_u10_u3_n1968 ) );
NAND2_X1 _u10_u3_U67  ( .A1(_u10_u3_n1967 ), .A2(_u10_u3_n1968 ), .ZN(_u10_u3_n1942 ) );
NAND3_X1 _u10_u3_U66  ( .A1(_u10_u3_n1964 ), .A2(_u10_u3_n1965 ), .A3(_u10_u3_n1966 ), .ZN(_u10_u3_n1943 ) );
AND4_X1 _u10_u3_U65  ( .A1(_u10_u3_n1961 ), .A2(_u10_u3_n1863 ), .A3(_u10_u3_n1962 ), .A4(_u10_u3_n1963 ), .ZN(_u10_u3_n1957 ) );
NOR2_X1 _u10_u3_U64  ( .A1(_u10_u3_n1959 ), .A2(_u10_u3_n1960 ), .ZN(_u10_u3_n1958 ) );
NOR2_X1 _u10_u3_U63  ( .A1(_u10_u3_n1957 ), .A2(_u10_u3_n1958 ), .ZN(_u10_u3_n1945 ) );
NOR2_X1 _u10_u3_U62  ( .A1(_u10_u3_n1955 ), .A2(_u10_u3_n1956 ), .ZN(_u10_u3_n1953 ) );
NOR4_X1 _u10_u3_U61  ( .A1(_u10_u3_n1952 ), .A2(_u10_u3_n1953 ), .A3(_u10_u3_n1846 ), .A4(_u10_u3_n1954 ), .ZN(_u10_u3_n1946 ) );
NOR2_X1 _u10_u3_U60  ( .A1(_u10_u3_n1950 ), .A2(_u10_u3_n1951 ), .ZN(_u10_u3_n1949 ) );
NOR2_X1 _u10_u3_U59  ( .A1(_u10_u3_n1948 ), .A2(_u10_u3_n1949 ), .ZN(_u10_u3_n1947 ) );
NOR3_X1 _u10_u3_U58  ( .A1(_u10_u3_n1945 ), .A2(_u10_u3_n1946 ), .A3(_u10_u3_n1947 ), .ZN(_u10_u3_n1944 ) );
NAND4_X1 _u10_u3_U57  ( .A1(_u10_u3_n1941 ), .A2(_u10_u3_n1942 ), .A3(_u10_u3_n1943 ), .A4(_u10_u3_n1944 ), .ZN(_u10_u3_n1824 ) );
NAND2_X1 _u10_u3_U56  ( .A1(_u10_u3_n1939 ), .A2(_u10_u3_n1940 ), .ZN(_u10_u3_n1938 ) );
NAND2_X1 _u10_u3_U55  ( .A1(_u10_u3_n1937 ), .A2(_u10_u3_n1938 ), .ZN(_u10_u3_n1903 ) );
NAND2_X1 _u10_u3_U54  ( .A1(_u10_u3_n1935 ), .A2(_u10_u3_n1936 ), .ZN(_u10_u3_n1934 ) );
NAND2_X1 _u10_u3_U53  ( .A1(_u10_u3_n1933 ), .A2(_u10_u3_n1934 ), .ZN(_u10_u3_n1931 ) );
NAND2_X1 _u10_u3_U52  ( .A1(_u10_u3_n1931 ), .A2(_u10_u3_n1932 ), .ZN(_u10_u3_n1904 ) );
NAND2_X1 _u10_u3_U51  ( .A1(_u10_u3_n1929 ), .A2(_u10_u3_n1930 ), .ZN(_u10_u3_n1927 ) );
NAND2_X1 _u10_u3_U50  ( .A1(_u10_u3_n1927 ), .A2(_u10_u3_n1928 ), .ZN(_u10_u3_n1905 ) );
NOR3_X1 _u10_u3_U49  ( .A1(_u10_u3_n1916 ), .A2(_u10_u3_n1925 ), .A3(_u10_u3_n1926 ), .ZN(_u10_u3_n1919 ) );
NOR2_X1 _u10_u3_U48  ( .A1(_u10_u3_n1923 ), .A2(_u10_u3_n1924 ), .ZN(_u10_u3_n1921 ) );
NOR2_X1 _u10_u3_U47  ( .A1(_u10_u3_n1921 ), .A2(_u10_u3_n1922 ), .ZN(_u10_u3_n1920 ) );
NOR2_X1 _u10_u3_U46  ( .A1(_u10_u3_n1919 ), .A2(_u10_u3_n1920 ), .ZN(_u10_u3_n1917 ) );
NOR2_X1 _u10_u3_U45  ( .A1(_u10_u3_n1917 ), .A2(_u10_u3_n1918 ), .ZN(_u10_u3_n1907 ) );
NOR2_X1 _u10_u3_U44  ( .A1(_u10_u3_n1915 ), .A2(_u10_u3_n1916 ), .ZN(_u10_u3_n1914 ) );
NOR2_X1 _u10_u3_U43  ( .A1(_u10_u3_n1914 ), .A2(1'b0), .ZN(_u10_u3_n1912 ));
NOR2_X1 _u10_u3_U42  ( .A1(_u10_u3_n1912 ), .A2(_u10_u3_n1913 ), .ZN(_u10_u3_n1908 ) );
NOR2_X1 _u10_u3_U41  ( .A1(_u10_u3_n1891 ), .A2(_u10_u3_n1911 ), .ZN(_u10_u3_n1910 ) );
NOR2_X1 _u10_u3_U40  ( .A1(_u10_u3_n1910 ), .A2(_u10_u3_n1868 ), .ZN(_u10_u3_n1909 ) );
NOR3_X1 _u10_u3_U39  ( .A1(_u10_u3_n1907 ), .A2(_u10_u3_n1908 ), .A3(_u10_u3_n1909 ), .ZN(_u10_u3_n1906 ) );
NAND4_X1 _u10_u3_U38  ( .A1(_u10_u3_n1903 ), .A2(_u10_u3_n1904 ), .A3(_u10_u3_n1905 ), .A4(_u10_u3_n1906 ), .ZN(_u10_u3_n1825 ) );
NAND2_X1 _u10_u3_U37  ( .A1(_u10_u3_n1901 ), .A2(_u10_u3_n1902 ), .ZN(_u10_u3_n1900 ) );
NAND2_X1 _u10_u3_U36  ( .A1(_u10_u3_n1899 ), .A2(_u10_u3_n1900 ), .ZN(_u10_u3_n1875 ) );
OR2_X1 _u10_u3_U35  ( .A1(_u10_u3_n1847 ), .A2(_u10_u3_n1898 ), .ZN(_u10_u3_n1897 ) );
NAND2_X1 _u10_u3_U34  ( .A1(_u10_u3_n1896 ), .A2(_u10_u3_n1897 ), .ZN(_u10_u3_n1895 ) );
NAND2_X1 _u10_u3_U33  ( .A1(_u10_u3_n1894 ), .A2(_u10_u3_n1895 ), .ZN(_u10_u3_n1876 ) );
NAND2_X1 _u10_u3_U32  ( .A1(_u10_u3_n1892 ), .A2(_u10_u3_n1893 ), .ZN(_u10_u3_n1877 ) );
NOR3_X1 _u10_u3_U31  ( .A1(_u10_u3_n1884 ), .A2(_u10_u3_n1890 ), .A3(_u10_u3_n1891 ), .ZN(_u10_u3_n1889 ) );
NOR2_X1 _u10_u3_U30  ( .A1(_u10_u3_n1840 ), .A2(_u10_u3_n1889 ), .ZN(_u10_u3_n1879 ) );
NOR2_X1 _u10_u3_U29  ( .A1(_u10_u3_n1887 ), .A2(_u10_u3_n1888 ), .ZN(_u10_u3_n1880 ) );
NOR3_X1 _u10_u3_U28  ( .A1(_u10_u3_n1884 ), .A2(_u10_u3_n1885 ), .A3(_u10_u3_n1886 ), .ZN(_u10_u3_n1883 ) );
NOR2_X1 _u10_u3_U27  ( .A1(_u10_u3_n1882 ), .A2(_u10_u3_n1883 ), .ZN(_u10_u3_n1881 ) );
NOR3_X1 _u10_u3_U26  ( .A1(_u10_u3_n1879 ), .A2(_u10_u3_n1880 ), .A3(_u10_u3_n1881 ), .ZN(_u10_u3_n1878 ) );
NAND4_X1 _u10_u3_U25  ( .A1(_u10_u3_n1875 ), .A2(_u10_u3_n1876 ), .A3(_u10_u3_n1877 ), .A4(_u10_u3_n1878 ), .ZN(_u10_u3_n1826 ) );
NOR3_X1 _u10_u3_U24  ( .A1(_u10_u3_n1872 ), .A2(_u10_u3_n1873 ), .A3(_u10_u3_n1874 ), .ZN(_u10_u3_n1871 ) );
NAND4_X1 _u10_u3_U23  ( .A1(_u10_u3_n1868 ), .A2(_u10_u3_n1869 ), .A3(_u10_u3_n1870 ), .A4(_u10_u3_n1871 ), .ZN(_u10_u3_n1867 ) );
NAND2_X1 _u10_u3_U22  ( .A1(_u10_u3_n1866 ), .A2(_u10_u3_n1867 ), .ZN(_u10_u3_n1865 ) );
NAND3_X1 _u10_u3_U21  ( .A1(_u10_u3_n1863 ), .A2(_u10_u3_n1864 ), .A3(_u10_u3_n1865 ), .ZN(_u10_u3_n1862 ) );
NAND2_X1 _u10_u3_U20  ( .A1(_u10_u3_n1861 ), .A2(_u10_u3_n1862 ), .ZN(_u10_u3_n1828 ) );
NAND3_X1 _u10_u3_U19  ( .A1(_u10_u3_n1858 ), .A2(_u10_u3_n1859 ), .A3(_u10_u3_n1860 ), .ZN(_u10_u3_n1857 ) );
NAND2_X1 _u10_u3_U18  ( .A1(_u10_u3_n1856 ), .A2(_u10_u3_n1857 ), .ZN(_u10_u3_n1829 ) );
OR2_X1 _u10_u3_U17  ( .A1(_u10_u3_n1854 ), .A2(_u10_u3_n1855 ), .ZN(_u10_u3_n1830 ) );
NOR2_X1 _u10_u3_U16  ( .A1(_u10_u3_n1852 ), .A2(_u10_u3_n1853 ), .ZN(_u10_u3_n1850 ) );
NOR3_X1 _u10_u3_U15  ( .A1(_u10_u3_n1850 ), .A2(_u10_u3_n1851 ), .A3(_u10_u3_n1838 ), .ZN(_u10_u3_n1848 ) );
NOR2_X1 _u10_u3_U14  ( .A1(_u10_u3_n1848 ), .A2(_u10_u3_n1849 ), .ZN(_u10_u3_n1832 ) );
NOR2_X1 _u10_u3_U13  ( .A1(_u10_u3_n1846 ), .A2(_u10_u3_n1847 ), .ZN(_u10_u3_n1845 ) );
NOR3_X1 _u10_u3_U12  ( .A1(_u10_u3_n1844 ), .A2(1'b0), .A3(_u10_u3_n1845 ),.ZN(_u10_u3_n1842 ) );
NOR2_X1 _u10_u3_U11  ( .A1(_u10_u3_n1842 ), .A2(_u10_u3_n1843 ), .ZN(_u10_u3_n1833 ) );
NOR2_X1 _u10_u3_U10  ( .A1(_u10_u3_n1840 ), .A2(_u10_u3_n1841 ), .ZN(_u10_u3_n1839 ) );
NOR3_X1 _u10_u3_U9  ( .A1(_u10_u3_n1837 ), .A2(_u10_u3_n1838 ), .A3(_u10_u3_n1839 ), .ZN(_u10_u3_n1835 ) );
NOR2_X1 _u10_u3_U8  ( .A1(_u10_u3_n1835 ), .A2(_u10_u3_n1836 ), .ZN(_u10_u3_n1834 ) );
NOR3_X1 _u10_u3_U7  ( .A1(_u10_u3_n1832 ), .A2(_u10_u3_n1833 ), .A3(_u10_u3_n1834 ), .ZN(_u10_u3_n1831 ) );
NAND4_X1 _u10_u3_U6  ( .A1(_u10_u3_n1828 ), .A2(_u10_u3_n1829 ), .A3(_u10_u3_n1830 ), .A4(_u10_u3_n1831 ), .ZN(_u10_u3_n1827 ) );
NOR4_X1 _u10_u3_U5  ( .A1(_u10_u3_n1824 ), .A2(_u10_u3_n1825 ), .A3(_u10_u3_n1826 ), .A4(_u10_u3_n1827 ), .ZN(_u10_u3_n1823 ) );
NAND4_X1 _u10_u3_U4  ( .A1(_u10_u3_n1820 ), .A2(_u10_u3_n1821 ), .A3(_u10_u3_n1822 ), .A4(_u10_u3_n1823 ), .ZN(_u10_u3_n1818 ) );
MUX2_X1 _u10_u3_U3  ( .A(_u10_u3_n1818 ), .B(_u10_SYNOPSYS_UNCONNECTED_12 ),.S(_u10_u3_n1819 ), .Z(_u10_u3_n1812 ) );
DFFR_X1 _u10_u3_state_reg_1_  ( .D(_u10_u3_n1812 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_12 ), .QN(_u10_u3_n1814 ));
DFFR_X1 _u10_u3_state_reg_2_  ( .D(_u10_u3_n1811 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_11 ), .QN(_u10_u3_n1815 ));
DFFR_X1 _u10_u3_state_reg_3_  ( .D(_u10_u3_n1810 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_10 ), .QN(_u10_u3_n1816 ));
DFFR_X1 _u10_u3_state_reg_4_  ( .D(_u10_u3_n1809 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_9 ), .QN(_u10_u3_n1817 ));
DFFR_X1 _u10_u3_state_reg_0_  ( .D(_u10_u3_n1808 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_13 ), .QN(_u10_u3_n1813 ));
NOR2_X1 _u10_u4_U1606  ( .A1(_u10_SYNOPSYS_UNCONNECTED_16 ), .A2(_u10_u4_n1814 ), .ZN(_u10_u4_n3174 ) );
NOR3_X1 _u10_u4_U1605  ( .A1(_u10_SYNOPSYS_UNCONNECTED_15 ), .A2(_u10_u4_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_18 ), .ZN(_u10_u4_n3328 ) );
NAND2_X1 _u10_u4_U1604  ( .A1(_u10_u4_n3174 ), .A2(_u10_u4_n3328 ), .ZN(_u10_u4_n1843 ) );
INV_X1 _u10_u4_U1603  ( .A(_u10_u4_n1843 ), .ZN(_u10_u4_n2461 ) );
INV_X1 _u10_u4_U1602  ( .A(1'b0), .ZN(_u10_u4_n2466 ) );
INV_X1 _u10_u4_U1601  ( .A(1'b0), .ZN(_u10_u4_n2305 ) );
NAND2_X1 _u10_u4_U1600  ( .A1(_u10_u4_n2466 ), .A2(_u10_u4_n2305 ), .ZN(_u10_u4_n1954 ) );
INV_X1 _u10_u4_U1599  ( .A(_u10_u4_n1954 ), .ZN(_u10_u4_n2467 ) );
INV_X1 _u10_u4_U1598  ( .A(1'b0), .ZN(_u10_u4_n1936 ) );
NOR2_X1 _u10_u4_U1597  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u4_n2223 ) );
INV_X1 _u10_u4_U1596  ( .A(1'b0), .ZN(_u10_u4_n1922 ) );
NAND2_X1 _u10_u4_U1595  ( .A1(_u10_u4_n2223 ), .A2(_u10_u4_n1922 ), .ZN(_u10_u4_n2200 ) );
NOR2_X1 _u10_u4_U1594  ( .A1(_u10_u4_n2200 ), .A2(1'b0), .ZN(_u10_u4_n2502 ));
INV_X1 _u10_u4_U1593  ( .A(1'b0), .ZN(_u10_u4_n2978 ) );
INV_X1 _u10_u4_U1592  ( .A(1'b0), .ZN(_u10_u4_n3000 ) );
NAND2_X1 _u10_u4_U1591  ( .A1(_u10_u4_n2978 ), .A2(_u10_u4_n3000 ), .ZN(_u10_u4_n3356 ) );
INV_X1 _u10_u4_U1590  ( .A(1'b0), .ZN(_u10_u4_n2405 ) );
INV_X1 _u10_u4_U1589  ( .A(1'b0), .ZN(_u10_u4_n2972 ) );
NAND2_X1 _u10_u4_U1588  ( .A1(_u10_u4_n2405 ), .A2(_u10_u4_n2972 ), .ZN(_u10_u4_n2008 ) );
NOR2_X1 _u10_u4_U1587  ( .A1(_u10_u4_n3356 ), .A2(_u10_u4_n2008 ), .ZN(_u10_u4_n2195 ) );
NAND2_X1 _u10_u4_U1586  ( .A1(_u10_u4_n2502 ), .A2(_u10_u4_n2195 ), .ZN(_u10_u4_n2490 ) );
INV_X1 _u10_u4_U1585  ( .A(1'b0), .ZN(_u10_u4_n3040 ) );
INV_X1 _u10_u4_U1584  ( .A(1'b0), .ZN(_u10_u4_n3006 ) );
NAND2_X1 _u10_u4_U1583  ( .A1(_u10_u4_n3040 ), .A2(_u10_u4_n3006 ), .ZN(_u10_u4_n2508 ) );
NOR2_X1 _u10_u4_U1582  ( .A1(_u10_u4_n2508 ), .A2(1'b0), .ZN(_u10_u4_n2493 ));
INV_X1 _u10_u4_U1581  ( .A(1'b0), .ZN(_u10_u4_n2038 ) );
NAND2_X1 _u10_u4_U1580  ( .A1(_u10_u4_n2493 ), .A2(_u10_u4_n2038 ), .ZN(_u10_u4_n2174 ) );
NOR2_X1 _u10_u4_U1579  ( .A1(_u10_u4_n2490 ), .A2(_u10_u4_n2174 ), .ZN(_u10_u4_n2659 ) );
INV_X1 _u10_u4_U1578  ( .A(1'b0), .ZN(_u10_u4_n2175 ) );
NAND3_X1 _u10_u4_U1577  ( .A1(_u10_u4_n2659 ), .A2(_u10_u4_n2175 ), .A3(1'b0), .ZN(_u10_u4_n3189 ) );
NOR2_X1 _u10_u4_U1576  ( .A1(_u10_u4_n3189 ), .A2(1'b0), .ZN(_u10_u4_n2528 ));
INV_X1 _u10_u4_U1575  ( .A(1'b0), .ZN(_u10_u4_n2837 ) );
NAND2_X1 _u10_u4_U1574  ( .A1(_u10_u4_n2528 ), .A2(_u10_u4_n2837 ), .ZN(_u10_u4_n2567 ) );
INV_X1 _u10_u4_U1573  ( .A(1'b0), .ZN(_u10_u4_n2080 ) );
INV_X1 _u10_u4_U1572  ( .A(1'b0), .ZN(_u10_u4_n2166 ) );
NAND2_X1 _u10_u4_U1571  ( .A1(_u10_u4_n2080 ), .A2(_u10_u4_n2166 ), .ZN(_u10_u4_n2840 ) );
NOR2_X1 _u10_u4_U1570  ( .A1(_u10_u4_n2567 ), .A2(_u10_u4_n2840 ), .ZN(_u10_u4_n2443 ) );
INV_X1 _u10_u4_U1569  ( .A(1'b0), .ZN(_u10_u4_n2600 ) );
INV_X1 _u10_u4_U1568  ( .A(1'b0), .ZN(_u10_u4_n2836 ) );
NAND2_X1 _u10_u4_U1567  ( .A1(_u10_u4_n2600 ), .A2(_u10_u4_n2836 ), .ZN(_u10_u4_n2428 ) );
INV_X1 _u10_u4_U1566  ( .A(_u10_u4_n2428 ), .ZN(_u10_u4_n2078 ) );
NAND2_X1 _u10_u4_U1565  ( .A1(_u10_u4_n2443 ), .A2(_u10_u4_n2078 ), .ZN(_u10_u4_n2282 ) );
INV_X1 _u10_u4_U1564  ( .A(1'b0), .ZN(_u10_u4_n2874 ) );
INV_X1 _u10_u4_U1563  ( .A(1'b0), .ZN(_u10_u4_n2031 ) );
NAND2_X1 _u10_u4_U1562  ( .A1(_u10_u4_n2874 ), .A2(_u10_u4_n2031 ), .ZN(_u10_u4_n1976 ) );
NOR2_X1 _u10_u4_U1561  ( .A1(_u10_u4_n2282 ), .A2(_u10_u4_n1976 ), .ZN(_u10_u4_n2411 ) );
NAND3_X1 _u10_u4_U1560  ( .A1(_u10_u4_n2467 ), .A2(_u10_u4_n1936 ), .A3(_u10_u4_n2411 ), .ZN(_u10_u4_n2464 ) );
NAND3_X1 _u10_u4_U1559  ( .A1(_u10_u4_n2166 ), .A2(_u10_u4_n2837 ), .A3(1'b0), .ZN(_u10_u4_n3276 ) );
INV_X1 _u10_u4_U1558  ( .A(_u10_u4_n3276 ), .ZN(_u10_u4_n2442 ) );
NAND3_X1 _u10_u4_U1557  ( .A1(_u10_u4_n2836 ), .A2(_u10_u4_n2080 ), .A3(_u10_u4_n2442 ), .ZN(_u10_u4_n2838 ) );
INV_X1 _u10_u4_U1556  ( .A(_u10_u4_n2838 ), .ZN(_u10_u4_n2850 ) );
NOR2_X1 _u10_u4_U1555  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u4_n2953 ) );
NAND2_X1 _u10_u4_U1554  ( .A1(_u10_u4_n2850 ), .A2(_u10_u4_n2953 ), .ZN(_u10_u4_n2947 ) );
INV_X1 _u10_u4_U1553  ( .A(_u10_u4_n2947 ), .ZN(_u10_u4_n2420 ) );
NAND2_X1 _u10_u4_U1552  ( .A1(_u10_u4_n1936 ), .A2(_u10_u4_n2874 ), .ZN(_u10_u4_n2030 ) );
INV_X1 _u10_u4_U1551  ( .A(_u10_u4_n2030 ), .ZN(_u10_u4_n2162 ) );
NAND2_X1 _u10_u4_U1550  ( .A1(_u10_u4_n2420 ), .A2(_u10_u4_n2162 ), .ZN(_u10_u4_n2828 ) );
INV_X1 _u10_u4_U1549  ( .A(_u10_u4_n2828 ), .ZN(_u10_u4_n2551 ) );
NAND2_X1 _u10_u4_U1548  ( .A1(_u10_u4_n2551 ), .A2(_u10_u4_n2467 ), .ZN(_u10_u4_n3416 ) );
NAND2_X1 _u10_u4_U1547  ( .A1(_u10_u4_n2464 ), .A2(_u10_u4_n3416 ), .ZN(_u10_u4_n2266 ) );
INV_X1 _u10_u4_U1546  ( .A(_u10_u4_n2266 ), .ZN(_u10_u4_n3410 ) );
NAND2_X1 _u10_u4_U1545  ( .A1(1'b0), .A2(_u10_u4_n2305 ), .ZN(_u10_u4_n3411 ) );
INV_X1 _u10_u4_U1544  ( .A(_u10_u4_n3356 ), .ZN(_u10_u4_n1983 ) );
NAND3_X1 _u10_u4_U1543  ( .A1(_u10_u4_n1983 ), .A2(_u10_u4_n2405 ), .A3(1'b0), .ZN(_u10_u4_n2022 ) );
INV_X1 _u10_u4_U1542  ( .A(_u10_u4_n2022 ), .ZN(_u10_u4_n2056 ) );
INV_X1 _u10_u4_U1541  ( .A(_u10_u4_n2840 ), .ZN(_u10_u4_n2059 ) );
INV_X1 _u10_u4_U1540  ( .A(1'b0), .ZN(_u10_u4_n1965 ) );
NAND2_X1 _u10_u4_U1539  ( .A1(_u10_u4_n2837 ), .A2(_u10_u4_n1965 ), .ZN(_u10_u4_n1852 ) );
INV_X1 _u10_u4_U1538  ( .A(_u10_u4_n1852 ), .ZN(_u10_u4_n3190 ) );
INV_X1 _u10_u4_U1537  ( .A(1'b0), .ZN(_u10_u4_n1853 ) );
NAND2_X1 _u10_u4_U1536  ( .A1(_u10_u4_n3190 ), .A2(_u10_u4_n1853 ), .ZN(_u10_u4_n2687 ) );
INV_X1 _u10_u4_U1535  ( .A(_u10_u4_n2687 ), .ZN(_u10_u4_n2019 ) );
NAND2_X1 _u10_u4_U1534  ( .A1(_u10_u4_n2059 ), .A2(_u10_u4_n2019 ), .ZN(_u10_u4_n2330 ) );
NOR2_X1 _u10_u4_U1533  ( .A1(_u10_u4_n2428 ), .A2(_u10_u4_n2330 ), .ZN(_u10_u4_n2036 ) );
NAND2_X1 _u10_u4_U1532  ( .A1(_u10_u4_n2056 ), .A2(_u10_u4_n2036 ), .ZN(_u10_u4_n3379 ) );
NOR2_X1 _u10_u4_U1531  ( .A1(_u10_u4_n3379 ), .A2(_u10_u4_n2030 ), .ZN(_u10_u4_n2026 ) );
INV_X1 _u10_u4_U1530  ( .A(1'b0), .ZN(_u10_u4_n2431 ) );
NOR2_X1 _u10_u4_U1529  ( .A1(_u10_u4_n2431 ), .A2(1'b0), .ZN(_u10_u4_n3062 ));
NAND2_X1 _u10_u4_U1528  ( .A1(_u10_u4_n3062 ), .A2(_u10_u4_n2195 ), .ZN(_u10_u4_n3407 ) );
NOR3_X1 _u10_u4_U1527  ( .A1(_u10_u4_n2687 ), .A2(1'b0), .A3(_u10_u4_n3407 ),.ZN(_u10_u4_n3275 ) );
NAND3_X1 _u10_u4_U1526  ( .A1(_u10_u4_n2836 ), .A2(_u10_u4_n2080 ), .A3(_u10_u4_n3275 ), .ZN(_u10_u4_n3297 ) );
INV_X1 _u10_u4_U1525  ( .A(_u10_u4_n3297 ), .ZN(_u10_u4_n3172 ) );
NAND2_X1 _u10_u4_U1524  ( .A1(_u10_u4_n3172 ), .A2(_u10_u4_n2600 ), .ZN(_u10_u4_n2226 ) );
NOR2_X1 _u10_u4_U1523  ( .A1(_u10_u4_n2226 ), .A2(1'b0), .ZN(_u10_u4_n2307 ));
INV_X1 _u10_u4_U1522  ( .A(_u10_u4_n2490 ), .ZN(_u10_u4_n2536 ) );
NAND3_X1 _u10_u4_U1521  ( .A1(_u10_u4_n2536 ), .A2(_u10_u4_n3040 ), .A3(1'b0), .ZN(_u10_u4_n3226 ) );
NOR2_X1 _u10_u4_U1520  ( .A1(_u10_u4_n3226 ), .A2(_u10_u4_n2330 ), .ZN(_u10_u4_n2441 ) );
NAND2_X1 _u10_u4_U1519  ( .A1(_u10_u4_n2441 ), .A2(_u10_u4_n2953 ), .ZN(_u10_u4_n2579 ) );
NOR2_X1 _u10_u4_U1518  ( .A1(_u10_u4_n2579 ), .A2(_u10_u4_n2030 ), .ZN(_u10_u4_n2550 ) );
NOR3_X1 _u10_u4_U1517  ( .A1(_u10_u4_n2026 ), .A2(_u10_u4_n2307 ), .A3(_u10_u4_n2550 ), .ZN(_u10_u4_n3394 ) );
NAND2_X1 _u10_u4_U1516  ( .A1(1'b0), .A2(_u10_u4_n2978 ), .ZN(_u10_u4_n3115 ) );
NOR2_X1 _u10_u4_U1515  ( .A1(_u10_u4_n3115 ), .A2(_u10_u4_n2330 ), .ZN(_u10_u4_n3126 ) );
NAND2_X1 _u10_u4_U1514  ( .A1(_u10_u4_n2162 ), .A2(_u10_u4_n2031 ), .ZN(_u10_u4_n2686 ) );
NOR2_X1 _u10_u4_U1513  ( .A1(_u10_u4_n2686 ), .A2(_u10_u4_n2428 ), .ZN(_u10_u4_n2108 ) );
NAND2_X1 _u10_u4_U1512  ( .A1(_u10_u4_n3126 ), .A2(_u10_u4_n2108 ), .ZN(_u10_u4_n3415 ) );
NAND2_X1 _u10_u4_U1511  ( .A1(_u10_u4_n3394 ), .A2(_u10_u4_n3415 ), .ZN(_u10_u4_n3089 ) );
NAND2_X1 _u10_u4_U1510  ( .A1(_u10_u4_n3089 ), .A2(_u10_u4_n2305 ), .ZN(_u10_u4_n3414 ) );
NAND2_X1 _u10_u4_U1509  ( .A1(_u10_u4_n2466 ), .A2(_u10_u4_n3414 ), .ZN(_u10_u4_n3118 ) );
NAND2_X1 _u10_u4_U1508  ( .A1(_u10_u4_n2078 ), .A2(_u10_u4_n2080 ), .ZN(_u10_u4_n2596 ) );
NAND2_X1 _u10_u4_U1507  ( .A1(1'b0), .A2(_u10_u4_n2493 ), .ZN(_u10_u4_n1961 ) );
NOR3_X1 _u10_u4_U1506  ( .A1(_u10_u4_n2490 ), .A2(1'b0), .A3(_u10_u4_n1961 ),.ZN(_u10_u4_n2054 ) );
NAND2_X1 _u10_u4_U1505  ( .A1(_u10_u4_n2054 ), .A2(_u10_u4_n3190 ), .ZN(_u10_u4_n2061 ) );
OR2_X1 _u10_u4_U1504  ( .A1(_u10_u4_n2596 ), .A2(_u10_u4_n2061 ), .ZN(_u10_u4_n1969 ) );
NOR3_X1 _u10_u4_U1503  ( .A1(_u10_u4_n1976 ), .A2(1'b0), .A3(_u10_u4_n1969 ),.ZN(_u10_u4_n2710 ) );
NAND2_X1 _u10_u4_U1502  ( .A1(_u10_u4_n2710 ), .A2(_u10_u4_n2467 ), .ZN(_u10_u4_n2545 ) );
INV_X1 _u10_u4_U1501  ( .A(_u10_u4_n2545 ), .ZN(_u10_u4_n2087 ) );
NOR2_X1 _u10_u4_U1500  ( .A1(_u10_u4_n3118 ), .A2(_u10_u4_n2087 ), .ZN(_u10_u4_n3145 ) );
NOR2_X1 _u10_u4_U1499  ( .A1(_u10_u4_n2030 ), .A2(1'b0), .ZN(_u10_u4_n2668 ));
NAND2_X1 _u10_u4_U1498  ( .A1(1'b0), .A2(_u10_u4_n2668 ), .ZN(_u10_u4_n2163 ) );
INV_X1 _u10_u4_U1497  ( .A(_u10_u4_n2163 ), .ZN(_u10_u4_n2875 ) );
INV_X1 _u10_u4_U1496  ( .A(_u10_u4_n1976 ), .ZN(_u10_u4_n2747 ) );
NAND3_X1 _u10_u4_U1495  ( .A1(_u10_u4_n2747 ), .A2(_u10_u4_n2600 ), .A3(1'b0), .ZN(_u10_u4_n3393 ) );
NOR3_X1 _u10_u4_U1494  ( .A1(1'b0), .A2(1'b0), .A3(_u10_u4_n3393 ), .ZN(_u10_u4_n3180 ) );
INV_X1 _u10_u4_U1493  ( .A(1'b0), .ZN(_u10_u4_n2113 ) );
INV_X1 _u10_u4_U1492  ( .A(1'b0), .ZN(_u10_u4_n3066 ) );
NAND2_X1 _u10_u4_U1491  ( .A1(_u10_u4_n2175 ), .A2(_u10_u4_n3066 ), .ZN(_u10_u4_n2216 ) );
INV_X1 _u10_u4_U1490  ( .A(_u10_u4_n2659 ), .ZN(_u10_u4_n2643 ) );
NOR2_X1 _u10_u4_U1489  ( .A1(_u10_u4_n2216 ), .A2(_u10_u4_n2643 ), .ZN(_u10_u4_n2049 ) );
AND2_X1 _u10_u4_U1488  ( .A1(_u10_u4_n2049 ), .A2(_u10_u4_n1853 ), .ZN(_u10_u4_n3223 ) );
NAND2_X1 _u10_u4_U1487  ( .A1(_u10_u4_n3223 ), .A2(_u10_u4_n1965 ), .ZN(_u10_u4_n2531 ) );
NOR2_X1 _u10_u4_U1486  ( .A1(_u10_u4_n2531 ), .A2(1'b0), .ZN(_u10_u4_n2884 ));
NAND2_X1 _u10_u4_U1485  ( .A1(_u10_u4_n2884 ), .A2(_u10_u4_n2166 ), .ZN(_u10_u4_n1841 ) );
NOR2_X1 _u10_u4_U1484  ( .A1(_u10_u4_n1841 ), .A2(1'b0), .ZN(_u10_u4_n3129 ));
NAND2_X1 _u10_u4_U1483  ( .A1(_u10_u4_n3129 ), .A2(_u10_u4_n2836 ), .ZN(_u10_u4_n2842 ) );
INV_X1 _u10_u4_U1482  ( .A(_u10_u4_n2842 ), .ZN(_u10_u4_n2833 ) );
NAND2_X1 _u10_u4_U1481  ( .A1(_u10_u4_n2833 ), .A2(_u10_u4_n2600 ), .ZN(_u10_u4_n2853 ) );
INV_X1 _u10_u4_U1480  ( .A(_u10_u4_n2853 ), .ZN(_u10_u4_n2082 ) );
NAND2_X1 _u10_u4_U1479  ( .A1(_u10_u4_n2082 ), .A2(_u10_u4_n2031 ), .ZN(_u10_u4_n2274 ) );
INV_X1 _u10_u4_U1478  ( .A(_u10_u4_n2274 ), .ZN(_u10_u4_n2669 ) );
NAND3_X1 _u10_u4_U1477  ( .A1(_u10_u4_n2668 ), .A2(_u10_u4_n2113 ), .A3(_u10_u4_n2669 ), .ZN(_u10_u4_n1858 ) );
INV_X1 _u10_u4_U1476  ( .A(_u10_u4_n1858 ), .ZN(_u10_u4_n3067 ) );
NAND2_X1 _u10_u4_U1475  ( .A1(_u10_u4_n3067 ), .A2(1'b0), .ZN(_u10_u4_n2092 ) );
INV_X1 _u10_u4_U1474  ( .A(_u10_u4_n2092 ), .ZN(_u10_u4_n3294 ) );
INV_X1 _u10_u4_U1473  ( .A(1'b0), .ZN(_u10_u4_n2446 ) );
INV_X1 _u10_u4_U1472  ( .A(1'b0), .ZN(_u10_u4_n2996 ) );
NAND2_X1 _u10_u4_U1471  ( .A1(_u10_u4_n3067 ), .A2(_u10_u4_n2996 ), .ZN(_u10_u4_n1847 ) );
NOR3_X1 _u10_u4_U1470  ( .A1(_u10_u4_n2446 ), .A2(1'b0), .A3(_u10_u4_n1847 ),.ZN(_u10_u4_n3413 ) );
NOR4_X1 _u10_u4_U1469  ( .A1(_u10_u4_n2875 ), .A2(_u10_u4_n3180 ), .A3(_u10_u4_n3294 ), .A4(_u10_u4_n3413 ), .ZN(_u10_u4_n3412 ) );
NAND4_X1 _u10_u4_U1468  ( .A1(_u10_u4_n3410 ), .A2(_u10_u4_n3411 ), .A3(_u10_u4_n3145 ), .A4(_u10_u4_n3412 ), .ZN(_u10_u4_n3409 ) );
NAND2_X1 _u10_u4_U1467  ( .A1(_u10_u4_n2461 ), .A2(_u10_u4_n3409 ), .ZN(_u10_u4_n3380 ) );
NOR2_X1 _u10_u4_U1466  ( .A1(_u10_u4_n1817 ), .A2(_u10_u4_n1816 ), .ZN(_u10_u4_n3368 ) );
AND2_X1 _u10_u4_U1465  ( .A1(_u10_u4_n3368 ), .A2(_u10_u4_n1813 ), .ZN(_u10_u4_n3320 ) );
NOR2_X1 _u10_u4_U1464  ( .A1(_u10_SYNOPSYS_UNCONNECTED_17 ), .A2(_u10_u4_n1815 ), .ZN(_u10_u4_n3236 ) );
NAND2_X1 _u10_u4_U1463  ( .A1(_u10_u4_n3320 ), .A2(_u10_u4_n3236 ), .ZN(_u10_u4_n2607 ) );
INV_X1 _u10_u4_U1462  ( .A(_u10_u4_n2607 ), .ZN(_u10_u4_n1966 ) );
INV_X1 _u10_u4_U1461  ( .A(_u10_u4_n2200 ), .ZN(_u10_u4_n3216 ) );
NAND2_X1 _u10_u4_U1460  ( .A1(1'b0), .A2(_u10_u4_n3216 ), .ZN(_u10_u4_n2367 ) );
INV_X1 _u10_u4_U1459  ( .A(_u10_u4_n2367 ), .ZN(_u10_u4_n3183 ) );
NAND2_X1 _u10_u4_U1458  ( .A1(_u10_u4_n3183 ), .A2(_u10_u4_n2195 ), .ZN(_u10_u4_n2194 ) );
INV_X1 _u10_u4_U1457  ( .A(_u10_u4_n2194 ), .ZN(_u10_u4_n2055 ) );
NAND2_X1 _u10_u4_U1456  ( .A1(_u10_u4_n2055 ), .A2(_u10_u4_n1853 ), .ZN(_u10_u4_n3401 ) );
INV_X1 _u10_u4_U1455  ( .A(_u10_u4_n2531 ), .ZN(_u10_u4_n2190 ) );
INV_X1 _u10_u4_U1454  ( .A(1'b0), .ZN(_u10_u4_n3001 ) );
NAND2_X1 _u10_u4_U1453  ( .A1(_u10_u4_n3001 ), .A2(_u10_u4_n2466 ), .ZN(_u10_u4_n2156 ) );
NOR2_X1 _u10_u4_U1452  ( .A1(_u10_u4_n2166 ), .A2(_u10_u4_n2596 ), .ZN(_u10_u4_n2594 ) );
NAND2_X1 _u10_u4_U1451  ( .A1(_u10_u4_n2594 ), .A2(_u10_u4_n2031 ), .ZN(_u10_u4_n2752 ) );
INV_X1 _u10_u4_U1450  ( .A(_u10_u4_n2752 ), .ZN(_u10_u4_n2421 ) );
NAND2_X1 _u10_u4_U1449  ( .A1(_u10_u4_n2421 ), .A2(_u10_u4_n2874 ), .ZN(_u10_u4_n2033 ) );
INV_X1 _u10_u4_U1448  ( .A(_u10_u4_n2033 ), .ZN(_u10_u4_n2742 ) );
NAND3_X1 _u10_u4_U1447  ( .A1(_u10_u4_n2305 ), .A2(_u10_u4_n1936 ), .A3(_u10_u4_n2742 ), .ZN(_u10_u4_n1896 ) );
OR3_X1 _u10_u4_U1446  ( .A1(_u10_u4_n2156 ), .A2(1'b0), .A3(_u10_u4_n1896 ),.ZN(_u10_u4_n2905 ) );
NAND2_X1 _u10_u4_U1445  ( .A1(_u10_u4_n2113 ), .A2(_u10_u4_n2996 ), .ZN(_u10_u4_n2719 ) );
NOR2_X1 _u10_u4_U1444  ( .A1(_u10_u4_n2719 ), .A2(1'b0), .ZN(_u10_u4_n2941 ));
INV_X1 _u10_u4_U1443  ( .A(_u10_u4_n2941 ), .ZN(_u10_u4_n2911 ) );
NOR2_X1 _u10_u4_U1442  ( .A1(_u10_u4_n2905 ), .A2(_u10_u4_n2911 ), .ZN(_u10_u4_n3222 ) );
INV_X1 _u10_u4_U1441  ( .A(_u10_u4_n3222 ), .ZN(_u10_u4_n2695 ) );
INV_X1 _u10_u4_U1440  ( .A(_u10_u4_n2156 ), .ZN(_u10_u4_n2089 ) );
NAND3_X1 _u10_u4_U1439  ( .A1(_u10_u4_n2089 ), .A2(_u10_u4_n2446 ), .A3(_u10_u4_n3180 ), .ZN(_u10_u4_n2902 ) );
NOR2_X1 _u10_u4_U1438  ( .A1(_u10_u4_n2902 ), .A2(_u10_u4_n2911 ), .ZN(_u10_u4_n2533 ) );
INV_X1 _u10_u4_U1437  ( .A(_u10_u4_n2533 ), .ZN(_u10_u4_n2485 ) );
NAND2_X1 _u10_u4_U1436  ( .A1(_u10_u4_n2695 ), .A2(_u10_u4_n2485 ), .ZN(_u10_u4_n2721 ) );
NAND2_X1 _u10_u4_U1435  ( .A1(1'b0), .A2(_u10_u4_n2113 ), .ZN(_u10_u4_n1868 ) );
INV_X1 _u10_u4_U1434  ( .A(_u10_u4_n1868 ), .ZN(_u10_u4_n2534 ) );
NOR2_X1 _u10_u4_U1433  ( .A1(_u10_u4_n2721 ), .A2(_u10_u4_n2534 ), .ZN(_u10_u4_n3231 ) );
NAND2_X1 _u10_u4_U1432  ( .A1(_u10_u4_n2467 ), .A2(_u10_u4_n3001 ), .ZN(_u10_u4_n2303 ) );
INV_X1 _u10_u4_U1431  ( .A(_u10_u4_n2303 ), .ZN(_u10_u4_n2549 ) );
INV_X1 _u10_u4_U1430  ( .A(1'b0), .ZN(_u10_u4_n2803 ) );
NAND2_X1 _u10_u4_U1429  ( .A1(_u10_u4_n2803 ), .A2(_u10_u4_n2446 ), .ZN(_u10_u4_n1846 ) );
INV_X1 _u10_u4_U1428  ( .A(_u10_u4_n1846 ), .ZN(_u10_u4_n2667 ) );
NAND3_X1 _u10_u4_U1427  ( .A1(_u10_u4_n2549 ), .A2(_u10_u4_n2667 ), .A3(1'b0), .ZN(_u10_u4_n2739 ) );
INV_X1 _u10_u4_U1426  ( .A(_u10_u4_n2739 ), .ZN(_u10_u4_n3272 ) );
INV_X1 _u10_u4_U1425  ( .A(_u10_u4_n2719 ), .ZN(_u10_u4_n2364 ) );
NAND2_X1 _u10_u4_U1424  ( .A1(_u10_u4_n3272 ), .A2(_u10_u4_n2364 ), .ZN(_u10_u4_n2852 ) );
INV_X1 _u10_u4_U1423  ( .A(_u10_u4_n2852 ), .ZN(_u10_u4_n2214 ) );
NAND2_X1 _u10_u4_U1422  ( .A1(_u10_u4_n2875 ), .A2(_u10_u4_n2089 ), .ZN(_u10_u4_n2097 ) );
INV_X1 _u10_u4_U1421  ( .A(_u10_u4_n2097 ), .ZN(_u10_u4_n2300 ) );
NAND2_X1 _u10_u4_U1420  ( .A1(_u10_u4_n2300 ), .A2(_u10_u4_n2446 ), .ZN(_u10_u4_n2001 ) );
NOR2_X1 _u10_u4_U1419  ( .A1(_u10_u4_n2001 ), .A2(_u10_u4_n2911 ), .ZN(_u10_u4_n2877 ) );
NOR2_X1 _u10_u4_U1418  ( .A1(_u10_u4_n2214 ), .A2(_u10_u4_n2877 ), .ZN(_u10_u4_n2940 ) );
NAND2_X1 _u10_u4_U1417  ( .A1(_u10_u4_n3231 ), .A2(_u10_u4_n2940 ), .ZN(_u10_u4_n3408 ) );
NAND2_X1 _u10_u4_U1416  ( .A1(_u10_u4_n2190 ), .A2(_u10_u4_n3408 ), .ZN(_u10_u4_n3402 ) );
NOR2_X1 _u10_u4_U1415  ( .A1(_u10_u4_n2446 ), .A2(_u10_u4_n2911 ), .ZN(_u10_u4_n3059 ) );
NAND2_X1 _u10_u4_U1414  ( .A1(_u10_u4_n3059 ), .A2(_u10_u4_n2190 ), .ZN(_u10_u4_n3404 ) );
AND3_X1 _u10_u4_U1413  ( .A1(_u10_u4_n3407 ), .A2(_u10_u4_n3226 ), .A3(_u10_u4_n3115 ), .ZN(_u10_u4_n3058 ) );
NAND2_X1 _u10_u4_U1412  ( .A1(_u10_u4_n3058 ), .A2(_u10_u4_n2022 ), .ZN(_u10_u4_n3406 ) );
NAND2_X1 _u10_u4_U1411  ( .A1(_u10_u4_n1853 ), .A2(_u10_u4_n3406 ), .ZN(_u10_u4_n3405 ) );
AND3_X1 _u10_u4_U1410  ( .A1(_u10_u4_n3404 ), .A2(_u10_u4_n1965 ), .A3(_u10_u4_n3405 ), .ZN(_u10_u4_n3063 ) );
NAND2_X1 _u10_u4_U1409  ( .A1(_u10_u4_n2667 ), .A2(_u10_u4_n3001 ), .ZN(_u10_u4_n1898 ) );
INV_X1 _u10_u4_U1408  ( .A(_u10_u4_n1898 ), .ZN(_u10_u4_n2835 ) );
NAND3_X1 _u10_u4_U1407  ( .A1(_u10_u4_n2364 ), .A2(_u10_u4_n2835 ), .A3(1'b0), .ZN(_u10_u4_n1869 ) );
NOR2_X1 _u10_u4_U1406  ( .A1(_u10_u4_n1869 ), .A2(_u10_u4_n2531 ), .ZN(_u10_u4_n2761 ) );
NOR3_X1 _u10_u4_U1405  ( .A1(_u10_u4_n2761 ), .A2(_u10_u4_n2528 ), .A3(_u10_u4_n2054 ), .ZN(_u10_u4_n3403 ) );
NAND4_X1 _u10_u4_U1404  ( .A1(_u10_u4_n3401 ), .A2(_u10_u4_n3402 ), .A3(_u10_u4_n3063 ), .A4(_u10_u4_n3403 ), .ZN(_u10_u4_n3400 ) );
NAND2_X1 _u10_u4_U1403  ( .A1(_u10_u4_n1966 ), .A2(_u10_u4_n3400 ), .ZN(_u10_u4_n3381 ) );
AND2_X1 _u10_u4_U1402  ( .A1(_u10_u4_n3368 ), .A2(_u10_SYNOPSYS_UNCONNECTED_18 ), .ZN(_u10_u4_n3319 ) );
NAND2_X1 _u10_u4_U1401  ( .A1(_u10_u4_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_17 ), .ZN(_u10_u4_n1849 ) );
INV_X1 _u10_u4_U1400  ( .A(_u10_u4_n1849 ), .ZN(_u10_u4_n2183 ) );
NAND2_X1 _u10_u4_U1399  ( .A1(_u10_u4_n2884 ), .A2(_u10_u4_n2183 ), .ZN(_u10_u4_n2883 ) );
INV_X1 _u10_u4_U1398  ( .A(_u10_u4_n2883 ), .ZN(_u10_u4_n1890 ) );
INV_X1 _u10_u4_U1397  ( .A(_u10_u4_n2940 ), .ZN(_u10_u4_n3278 ) );
NAND2_X1 _u10_u4_U1396  ( .A1(_u10_u4_n1890 ), .A2(_u10_u4_n3278 ), .ZN(_u10_u4_n3382 ) );
NAND2_X1 _u10_u4_U1395  ( .A1(_u10_u4_n3059 ), .A2(_u10_u4_n2669 ), .ZN(_u10_u4_n3399 ) );
NAND2_X1 _u10_u4_U1394  ( .A1(_u10_u4_n2031 ), .A2(_u10_u4_n3399 ), .ZN(_u10_u4_n3398 ) );
NAND2_X1 _u10_u4_U1393  ( .A1(_u10_u4_n2162 ), .A2(_u10_u4_n3398 ), .ZN(_u10_u4_n3395 ) );
NAND3_X1 _u10_u4_U1392  ( .A1(_u10_u4_n2747 ), .A2(_u10_u4_n2078 ), .A3(_u10_u4_n3126 ), .ZN(_u10_u4_n3396 ) );
NAND2_X1 _u10_u4_U1391  ( .A1(_u10_u4_n2055 ), .A2(_u10_u4_n2036 ), .ZN(_u10_u4_n2285 ) );
NOR2_X1 _u10_u4_U1390  ( .A1(_u10_u4_n2285 ), .A2(_u10_u4_n2030 ), .ZN(_u10_u4_n3349 ) );
INV_X1 _u10_u4_U1389  ( .A(_u10_u4_n3349 ), .ZN(_u10_u4_n1933 ) );
INV_X1 _u10_u4_U1388  ( .A(_u10_u4_n2710 ), .ZN(_u10_u4_n3397 ) );
NAND4_X1 _u10_u4_U1387  ( .A1(_u10_u4_n3395 ), .A2(_u10_u4_n3396 ), .A3(_u10_u4_n1933 ), .A4(_u10_u4_n3397 ), .ZN(_u10_u4_n3389 ) );
NAND2_X1 _u10_u4_U1386  ( .A1(_u10_u4_n1936 ), .A2(_u10_u4_n2828 ), .ZN(_u10_u4_n3141 ) );
INV_X1 _u10_u4_U1385  ( .A(_u10_u4_n3141 ), .ZN(_u10_u4_n2302 ) );
NAND2_X1 _u10_u4_U1384  ( .A1(_u10_u4_n3394 ), .A2(_u10_u4_n2302 ), .ZN(_u10_u4_n3390 ) );
NOR2_X1 _u10_u4_U1383  ( .A1(_u10_u4_n1869 ), .A2(_u10_u4_n2274 ), .ZN(_u10_u4_n3378 ) );
INV_X1 _u10_u4_U1382  ( .A(_u10_u4_n3378 ), .ZN(_u10_u4_n2748 ) );
NOR2_X1 _u10_u4_U1381  ( .A1(1'b0), .A2(_u10_u4_n2748 ), .ZN(_u10_u4_n3391 ));
NAND2_X1 _u10_u4_U1380  ( .A1(_u10_u4_n2534 ), .A2(_u10_u4_n2669 ), .ZN(_u10_u4_n2383 ) );
INV_X1 _u10_u4_U1379  ( .A(_u10_u4_n2383 ), .ZN(_u10_u4_n1978 ) );
NAND2_X1 _u10_u4_U1378  ( .A1(_u10_u4_n1978 ), .A2(_u10_u4_n2874 ), .ZN(_u10_u4_n3392 ) );
INV_X1 _u10_u4_U1377  ( .A(_u10_u4_n2411 ), .ZN(_u10_u4_n2164 ) );
NAND4_X1 _u10_u4_U1376  ( .A1(_u10_u4_n3392 ), .A2(_u10_u4_n3393 ), .A3(_u10_u4_n2033 ), .A4(_u10_u4_n2164 ), .ZN(_u10_u4_n2476 ) );
NOR4_X1 _u10_u4_U1375  ( .A1(_u10_u4_n3389 ), .A2(_u10_u4_n3390 ), .A3(_u10_u4_n3391 ), .A4(_u10_u4_n2476 ), .ZN(_u10_u4_n3388 ) );
NAND2_X1 _u10_u4_U1374  ( .A1(_u10_u4_n3236 ), .A2(_u10_u4_n3328 ), .ZN(_u10_u4_n2025 ) );
NOR2_X1 _u10_u4_U1373  ( .A1(_u10_u4_n3388 ), .A2(_u10_u4_n2025 ), .ZN(_u10_u4_n3384 ) );
NOR2_X1 _u10_u4_U1372  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u4_n2152 ) );
NAND2_X1 _u10_u4_U1371  ( .A1(_u10_u4_n2152 ), .A2(_u10_u4_n2175 ), .ZN(_u10_u4_n2722 ) );
INV_X1 _u10_u4_U1370  ( .A(_u10_u4_n2722 ), .ZN(_u10_u4_n2588 ) );
NAND2_X1 _u10_u4_U1369  ( .A1(_u10_u4_n2549 ), .A2(_u10_u4_n3349 ), .ZN(_u10_u4_n2091 ) );
NOR2_X1 _u10_u4_U1368  ( .A1(_u10_u4_n2091 ), .A2(_u10_u4_n1846 ), .ZN(_u10_u4_n2128 ) );
NAND3_X1 _u10_u4_U1367  ( .A1(_u10_u4_n3066 ), .A2(_u10_u4_n2113 ), .A3(_u10_u4_n2128 ), .ZN(_u10_u4_n2342 ) );
INV_X1 _u10_u4_U1366  ( .A(_u10_u4_n2342 ), .ZN(_u10_u4_n3316 ) );
NAND2_X1 _u10_u4_U1365  ( .A1(_u10_u4_n2588 ), .A2(_u10_u4_n3316 ), .ZN(_u10_u4_n2142 ) );
NOR2_X1 _u10_u4_U1364  ( .A1(_u10_u4_n1954 ), .A2(_u10_u4_n1898 ), .ZN(_u10_u4_n2255 ) );
NAND2_X1 _u10_u4_U1363  ( .A1(_u10_u4_n2255 ), .A2(_u10_u4_n2996 ), .ZN(_u10_u4_n1915 ) );
INV_X1 _u10_u4_U1362  ( .A(_u10_u4_n1915 ), .ZN(_u10_u4_n2251 ) );
NAND2_X1 _u10_u4_U1361  ( .A1(_u10_u4_n2251 ), .A2(_u10_u4_n2113 ), .ZN(_u10_u4_n1925 ) );
INV_X1 _u10_u4_U1360  ( .A(_u10_u4_n2026 ), .ZN(_u10_u4_n3340 ) );
NOR3_X1 _u10_u4_U1359  ( .A1(_u10_u4_n1925 ), .A2(_u10_u4_n2216 ), .A3(_u10_u4_n3340 ), .ZN(_u10_u4_n2003 ) );
INV_X1 _u10_u4_U1358  ( .A(1'b0), .ZN(_u10_u4_n1930 ) );
NAND2_X1 _u10_u4_U1357  ( .A1(_u10_u4_n2003 ), .A2(_u10_u4_n1930 ), .ZN(_u10_u4_n3387 ) );
AND2_X1 _u10_u4_U1356  ( .A1(_u10_u4_n2142 ), .A2(_u10_u4_n3387 ), .ZN(_u10_u4_n3366 ) );
NOR3_X1 _u10_u4_U1355  ( .A1(_u10_u4_n1813 ), .A2(_u10_u4_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_14 ), .ZN(_u10_u4_n3360 ) );
NOR2_X1 _u10_u4_U1354  ( .A1(_u10_SYNOPSYS_UNCONNECTED_16 ), .A2(_u10_SYNOPSYS_UNCONNECTED_17 ), .ZN(_u10_u4_n3136 ) );
NAND2_X1 _u10_u4_U1353  ( .A1(_u10_u4_n3360 ), .A2(_u10_u4_n3136 ), .ZN(_u10_u4_n2344 ) );
NOR2_X1 _u10_u4_U1352  ( .A1(_u10_u4_n3366 ), .A2(_u10_u4_n2344 ), .ZN(_u10_u4_n3385 ) );
NOR3_X1 _u10_u4_U1351  ( .A1(_u10_SYNOPSYS_UNCONNECTED_14 ), .A2(_u10_u4_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_18 ), .ZN(_u10_u4_n3342 ) );
NAND2_X1 _u10_u4_U1350  ( .A1(_u10_u4_n3342 ), .A2(_u10_u4_n3136 ), .ZN(_u10_u4_n2584 ) );
NOR2_X1 _u10_u4_U1349  ( .A1(_u10_u4_n2584 ), .A2(1'b0), .ZN(_u10_u4_n2139 ));
INV_X1 _u10_u4_U1348  ( .A(_u10_u4_n2216 ), .ZN(_u10_u4_n2106 ) );
AND2_X1 _u10_u4_U1347  ( .A1(_u10_u4_n2152 ), .A2(_u10_u4_n2106 ), .ZN(_u10_u4_n2336 ) );
NAND2_X1 _u10_u4_U1346  ( .A1(_u10_u4_n2139 ), .A2(_u10_u4_n2336 ), .ZN(_u10_u4_n2365 ) );
INV_X1 _u10_u4_U1345  ( .A(_u10_u4_n2365 ), .ZN(_u10_u4_n2004 ) );
AND2_X1 _u10_u4_U1344  ( .A1(_u10_u4_n2877 ), .A2(_u10_u4_n2004 ), .ZN(_u10_u4_n3386 ) );
NOR3_X1 _u10_u4_U1343  ( .A1(_u10_u4_n3384 ), .A2(_u10_u4_n3385 ), .A3(_u10_u4_n3386 ), .ZN(_u10_u4_n3383 ) );
NAND4_X1 _u10_u4_U1342  ( .A1(_u10_u4_n3380 ), .A2(_u10_u4_n3381 ), .A3(_u10_u4_n3382 ), .A4(_u10_u4_n3383 ), .ZN(_u10_u4_n3191 ) );
NAND2_X1 _u10_u4_U1341  ( .A1(_u10_u4_n2285 ), .A2(_u10_u4_n3379 ), .ZN(_u10_u4_n1975 ) );
NOR3_X1 _u10_u4_U1340  ( .A1(_u10_u4_n3378 ), .A2(1'b0), .A3(_u10_u4_n1975 ),.ZN(_u10_u4_n3122 ) );
AND4_X1 _u10_u4_U1339  ( .A1(_u10_u4_n2752 ), .A2(_u10_u4_n2383 ), .A3(_u10_u4_n1969 ), .A4(_u10_u4_n3122 ), .ZN(_u10_u4_n3377 ) );
NOR2_X1 _u10_u4_U1338  ( .A1(_u10_u4_n1814 ), .A2(_u10_u4_n1815 ), .ZN(_u10_u4_n3147 ) );
NAND2_X1 _u10_u4_U1337  ( .A1(_u10_u4_n3328 ), .A2(_u10_u4_n3147 ), .ZN(_u10_u4_n2359 ) );
NOR2_X1 _u10_u4_U1336  ( .A1(_u10_u4_n3377 ), .A2(_u10_u4_n2359 ), .ZN(_u10_u4_n3362 ) );
INV_X1 _u10_u4_U1335  ( .A(_u10_u4_n2008 ), .ZN(_u10_u4_n3097 ) );
NOR3_X1 _u10_u4_U1334  ( .A1(_u10_SYNOPSYS_UNCONNECTED_14 ), .A2(_u10_u4_n1813 ), .A3(_u10_SYNOPSYS_UNCONNECTED_15 ), .ZN(_u10_u4_n3269 ) );
NAND2_X1 _u10_u4_U1333  ( .A1(_u10_u4_n3269 ), .A2(_u10_u4_n3136 ), .ZN(_u10_u4_n3109 ) );
INV_X1 _u10_u4_U1332  ( .A(_u10_u4_n3109 ), .ZN(_u10_u4_n2999 ) );
INV_X1 _u10_u4_U1331  ( .A(_u10_u4_n2508 ), .ZN(_u10_u4_n2103 ) );
NAND2_X1 _u10_u4_U1330  ( .A1(_u10_u4_n2336 ), .A2(_u10_u4_n2103 ), .ZN(_u10_u4_n2249 ) );
NOR2_X1 _u10_u4_U1329  ( .A1(_u10_u4_n2249 ), .A2(1'b0), .ZN(_u10_u4_n1866 ));
NAND2_X1 _u10_u4_U1328  ( .A1(_u10_u4_n1866 ), .A2(_u10_u4_n1922 ), .ZN(_u10_u4_n2632 ) );
INV_X1 _u10_u4_U1327  ( .A(_u10_u4_n2223 ), .ZN(_u10_u4_n1918 ) );
NOR2_X1 _u10_u4_U1326  ( .A1(_u10_u4_n2632 ), .A2(_u10_u4_n1918 ), .ZN(_u10_u4_n1981 ) );
NAND3_X1 _u10_u4_U1325  ( .A1(_u10_u4_n3097 ), .A2(_u10_u4_n2999 ), .A3(_u10_u4_n1981 ), .ZN(_u10_u4_n3034 ) );
NOR3_X1 _u10_u4_U1324  ( .A1(_u10_SYNOPSYS_UNCONNECTED_15 ), .A2(_u10_SYNOPSYS_UNCONNECTED_14 ), .A3(_u10_SYNOPSYS_UNCONNECTED_18 ),.ZN(_u10_u4_n3302 ) );
NAND2_X1 _u10_u4_U1323  ( .A1(_u10_u4_n3302 ), .A2(_u10_u4_n3174 ), .ZN(_u10_u4_n3162 ) );
INV_X1 _u10_u4_U1322  ( .A(_u10_u4_n3162 ), .ZN(_u10_u4_n2979 ) );
NAND2_X1 _u10_u4_U1321  ( .A1(_u10_u4_n2979 ), .A2(_u10_u4_n2972 ), .ZN(_u10_u4_n1984 ) );
AND2_X1 _u10_u4_U1320  ( .A1(_u10_u4_n3302 ), .A2(_u10_u4_n3136 ), .ZN(_u10_u4_n2977 ) );
NAND3_X1 _u10_u4_U1319  ( .A1(_u10_u4_n2977 ), .A2(_u10_u4_n3000 ), .A3(_u10_u4_n3097 ), .ZN(_u10_u4_n3376 ) );
NAND2_X1 _u10_u4_U1318  ( .A1(_u10_u4_n1984 ), .A2(_u10_u4_n3376 ), .ZN(_u10_u4_n3375 ) );
NAND2_X1 _u10_u4_U1317  ( .A1(_u10_u4_n1981 ), .A2(_u10_u4_n3375 ), .ZN(_u10_u4_n2798 ) );
NAND2_X1 _u10_u4_U1316  ( .A1(_u10_u4_n3034 ), .A2(_u10_u4_n2798 ), .ZN(_u10_u4_n2007 ) );
NAND2_X1 _u10_u4_U1315  ( .A1(_u10_u4_n3269 ), .A2(_u10_u4_n3147 ), .ZN(_u10_u4_n2102 ) );
NOR2_X1 _u10_u4_U1314  ( .A1(_u10_u4_n2249 ), .A2(_u10_u4_n2102 ), .ZN(_u10_u4_n3323 ) );
INV_X1 _u10_u4_U1313  ( .A(_u10_u4_n3323 ), .ZN(_u10_u4_n3374 ) );
INV_X1 _u10_u4_U1312  ( .A(_u10_u4_n2344 ), .ZN(_u10_u4_n2002 ) );
NAND2_X1 _u10_u4_U1311  ( .A1(_u10_u4_n2336 ), .A2(_u10_u4_n2002 ), .ZN(_u10_u4_n3225 ) );
NAND2_X1 _u10_u4_U1310  ( .A1(_u10_u4_n3374 ), .A2(_u10_u4_n3225 ), .ZN(_u10_u4_n2488 ) );
NAND2_X1 _u10_u4_U1309  ( .A1(_u10_u4_n3342 ), .A2(_u10_u4_n3236 ), .ZN(_u10_u4_n2253 ) );
NOR2_X1 _u10_u4_U1308  ( .A1(_u10_u4_n2253 ), .A2(1'b0), .ZN(_u10_u4_n1885 ));
NAND2_X1 _u10_u4_U1307  ( .A1(_u10_u4_n3360 ), .A2(_u10_u4_n3174 ), .ZN(_u10_u4_n2254 ) );
INV_X1 _u10_u4_U1306  ( .A(_u10_u4_n2254 ), .ZN(_u10_u4_n2986 ) );
NAND2_X1 _u10_u4_U1305  ( .A1(_u10_u4_n2106 ), .A2(_u10_u4_n2986 ), .ZN(_u10_u4_n1913 ) );
INV_X1 _u10_u4_U1304  ( .A(_u10_u4_n1913 ), .ZN(_u10_u4_n2377 ) );
OR4_X1 _u10_u4_U1303  ( .A1(_u10_u4_n2007 ), .A2(_u10_u4_n2488 ), .A3(_u10_u4_n1885 ), .A4(_u10_u4_n2377 ), .ZN(_u10_u4_n3373 ) );
NAND2_X1 _u10_u4_U1302  ( .A1(_u10_u4_n2534 ), .A2(_u10_u4_n3373 ), .ZN(_u10_u4_n3370 ) );
NAND2_X1 _u10_u4_U1301  ( .A1(_u10_u4_n3342 ), .A2(_u10_u4_n3174 ), .ZN(_u10_u4_n2037 ) );
NAND2_X1 _u10_u4_U1300  ( .A1(_u10_u4_n2037 ), .A2(_u10_u4_n2254 ), .ZN(_u10_u4_n3372 ) );
NAND2_X1 _u10_u4_U1299  ( .A1(_u10_u4_n2003 ), .A2(_u10_u4_n3372 ), .ZN(_u10_u4_n3371 ) );
NAND2_X1 _u10_u4_U1298  ( .A1(_u10_u4_n3370 ), .A2(_u10_u4_n3371 ), .ZN(_u10_u4_n3363 ) );
NOR2_X1 _u10_u4_U1297  ( .A1(_u10_u4_n2490 ), .A2(_u10_u4_n1961 ), .ZN(_u10_u4_n3369 ) );
NAND2_X1 _u10_u4_U1296  ( .A1(_u10_u4_n2534 ), .A2(_u10_u4_n2049 ), .ZN(_u10_u4_n2646 ) );
INV_X1 _u10_u4_U1295  ( .A(_u10_u4_n2646 ), .ZN(_u10_u4_n3055 ) );
NOR2_X1 _u10_u4_U1294  ( .A1(_u10_u4_n3369 ), .A2(_u10_u4_n3055 ), .ZN(_u10_u4_n3367 ) );
NAND2_X1 _u10_u4_U1293  ( .A1(_u10_u4_n3368 ), .A2(_u10_u4_n3147 ), .ZN(_u10_u4_n2495 ) );
NOR2_X1 _u10_u4_U1292  ( .A1(_u10_u4_n3367 ), .A2(_u10_u4_n2495 ), .ZN(_u10_u4_n3364 ) );
INV_X1 _u10_u4_U1291  ( .A(_u10_u4_n2139 ), .ZN(_u10_u4_n3254 ) );
NOR2_X1 _u10_u4_U1290  ( .A1(_u10_u4_n3366 ), .A2(_u10_u4_n3254 ), .ZN(_u10_u4_n3365 ) );
NOR4_X1 _u10_u4_U1289  ( .A1(_u10_u4_n3362 ), .A2(_u10_u4_n3363 ), .A3(_u10_u4_n3364 ), .A4(_u10_u4_n3365 ), .ZN(_u10_u4_n3305 ) );
NAND2_X1 _u10_u4_U1288  ( .A1(_u10_u4_n3302 ), .A2(_u10_u4_n3147 ), .ZN(_u10_u4_n2980 ) );
NAND2_X1 _u10_u4_U1287  ( .A1(_u10_u4_n2102 ), .A2(_u10_u4_n2980 ), .ZN(_u10_u4_n2177 ) );
NAND2_X1 _u10_u4_U1286  ( .A1(_u10_u4_n2003 ), .A2(_u10_u4_n2493 ), .ZN(_u10_u4_n1962 ) );
NAND2_X1 _u10_u4_U1285  ( .A1(_u10_u4_n1961 ), .A2(_u10_u4_n1962 ), .ZN(_u10_u4_n3361 ) );
NAND2_X1 _u10_u4_U1284  ( .A1(_u10_u4_n2177 ), .A2(_u10_u4_n3361 ), .ZN(_u10_u4_n3357 ) );
NAND2_X1 _u10_u4_U1283  ( .A1(_u10_u4_n3236 ), .A2(_u10_u4_n3360 ), .ZN(_u10_u4_n1859 ) );
INV_X1 _u10_u4_U1282  ( .A(_u10_u4_n1859 ), .ZN(_u10_u4_n2256 ) );
NAND3_X1 _u10_u4_U1281  ( .A1(_u10_u4_n2256 ), .A2(_u10_u4_n2113 ), .A3(_u10_u4_n2128 ), .ZN(_u10_u4_n3358 ) );
NOR2_X1 _u10_u4_U1280  ( .A1(_u10_u4_n2877 ), .A2(_u10_u4_n3222 ), .ZN(_u10_u4_n3347 ) );
NAND2_X1 _u10_u4_U1279  ( .A1(_u10_u4_n3347 ), .A2(_u10_u4_n1869 ), .ZN(_u10_u4_n2005 ) );
NAND2_X1 _u10_u4_U1278  ( .A1(_u10_u4_n2488 ), .A2(_u10_u4_n2005 ), .ZN(_u10_u4_n3359 ) );
NAND3_X1 _u10_u4_U1277  ( .A1(_u10_u4_n3357 ), .A2(_u10_u4_n3358 ), .A3(_u10_u4_n3359 ), .ZN(_u10_u4_n3352 ) );
NAND2_X1 _u10_u4_U1276  ( .A1(_u10_u4_n3320 ), .A2(_u10_u4_n3136 ), .ZN(_u10_u4_n2356 ) );
INV_X1 _u10_u4_U1275  ( .A(_u10_u4_n2356 ), .ZN(_u10_u4_n2830 ) );
NAND2_X1 _u10_u4_U1274  ( .A1(_u10_u4_n2830 ), .A2(_u10_u4_n2836 ), .ZN(_u10_u4_n2291 ) );
NOR3_X1 _u10_u4_U1273  ( .A1(_u10_u4_n2291 ), .A2(_u10_u4_n2330 ), .A3(_u10_u4_n2022 ), .ZN(_u10_u4_n3353 ) );
INV_X1 _u10_u4_U1272  ( .A(_u10_u4_n1925 ), .ZN(_u10_u4_n2105 ) );
AND2_X1 _u10_u4_U1271  ( .A1(_u10_u4_n2108 ), .A2(_u10_u4_n2105 ), .ZN(_u10_u4_n2915 ) );
INV_X1 _u10_u4_U1270  ( .A(_u10_u4_n2330 ), .ZN(_u10_u4_n2107 ) );
NAND2_X1 _u10_u4_U1269  ( .A1(_u10_u4_n2915 ), .A2(_u10_u4_n2107 ), .ZN(_u10_u4_n2203 ) );
INV_X1 _u10_u4_U1268  ( .A(_u10_u4_n2203 ), .ZN(_u10_u4_n1982 ) );
NAND2_X1 _u10_u4_U1267  ( .A1(_u10_u4_n1982 ), .A2(_u10_u4_n2536 ), .ZN(_u10_u4_n2587 ) );
INV_X1 _u10_u4_U1266  ( .A(_u10_u4_n2587 ), .ZN(_u10_u4_n2697 ) );
NAND3_X1 _u10_u4_U1265  ( .A1(_u10_u4_n2697 ), .A2(_u10_u4_n2493 ), .A3(_u10_u4_n2377 ), .ZN(_u10_u4_n2412 ) );
INV_X1 _u10_u4_U1264  ( .A(_u10_u4_n2412 ), .ZN(_u10_u4_n3354 ) );
NAND2_X1 _u10_u4_U1263  ( .A1(_u10_u4_n3174 ), .A2(_u10_u4_n3269 ), .ZN(_u10_u4_n2375 ) );
INV_X1 _u10_u4_U1262  ( .A(_u10_u4_n2375 ), .ZN(_u10_u4_n2507 ) );
NAND2_X1 _u10_u4_U1261  ( .A1(_u10_u4_n1981 ), .A2(_u10_u4_n2507 ), .ZN(_u10_u4_n2621 ) );
NOR4_X1 _u10_u4_U1260  ( .A1(1'b0), .A2(_u10_u4_n3356 ), .A3(_u10_u4_n2203 ),.A4(_u10_u4_n2621 ), .ZN(_u10_u4_n3355 ) );
NOR4_X1 _u10_u4_U1259  ( .A1(_u10_u4_n3352 ), .A2(_u10_u4_n3353 ), .A3(_u10_u4_n3354 ), .A4(_u10_u4_n3355 ), .ZN(_u10_u4_n3306 ) );
NOR2_X1 _u10_u4_U1258  ( .A1(_u10_u4_n2842 ), .A2(_u10_u4_n2356 ), .ZN(_u10_u4_n1891 ) );
INV_X1 _u10_u4_U1257  ( .A(_u10_u4_n1869 ), .ZN(_u10_u4_n2885 ) );
NAND2_X1 _u10_u4_U1256  ( .A1(_u10_u4_n1891 ), .A2(_u10_u4_n2885 ), .ZN(_u10_u4_n3330 ) );
NAND2_X1 _u10_u4_U1255  ( .A1(_u10_u4_n2761 ), .A2(_u10_u4_n2837 ), .ZN(_u10_u4_n3351 ) );
NAND3_X1 _u10_u4_U1254  ( .A1(_u10_u4_n2884 ), .A2(_u10_u4_n2080 ), .A3(_u10_u4_n2915 ), .ZN(_u10_u4_n2762 ) );
NAND2_X1 _u10_u4_U1253  ( .A1(_u10_u4_n2055 ), .A2(_u10_u4_n2019 ), .ZN(_u10_u4_n3259 ) );
NAND4_X1 _u10_u4_U1252  ( .A1(_u10_u4_n3351 ), .A2(_u10_u4_n2762 ), .A3(_u10_u4_n2061 ), .A4(_u10_u4_n3259 ), .ZN(_u10_u4_n3350 ) );
NAND2_X1 _u10_u4_U1251  ( .A1(_u10_u4_n2183 ), .A2(_u10_u4_n3350 ), .ZN(_u10_u4_n3331 ) );
NAND2_X1 _u10_u4_U1250  ( .A1(_u10_u4_n3349 ), .A2(_u10_u4_n2305 ), .ZN(_u10_u4_n3348 ) );
NAND2_X1 _u10_u4_U1249  ( .A1(_u10_u4_n1896 ), .A2(_u10_u4_n3348 ), .ZN(_u10_u4_n3176 ) );
NAND2_X1 _u10_u4_U1248  ( .A1(_u10_u4_n2461 ), .A2(_u10_u4_n3176 ), .ZN(_u10_u4_n3332 ) );
INV_X1 _u10_u4_U1247  ( .A(_u10_u4_n2495 ), .ZN(_u10_u4_n2063 ) );
NAND2_X1 _u10_u4_U1246  ( .A1(_u10_u4_n2049 ), .A2(_u10_u4_n2063 ), .ZN(_u10_u4_n2886 ) );
NOR2_X1 _u10_u4_U1245  ( .A1(_u10_u4_n3347 ), .A2(_u10_u4_n2886 ), .ZN(_u10_u4_n3334 ) );
NAND2_X1 _u10_u4_U1244  ( .A1(1'b0), .A2(_u10_u4_n2835 ), .ZN(_u10_u4_n3344 ) );
NAND2_X1 _u10_u4_U1243  ( .A1(_u10_u4_n2001 ), .A2(_u10_u4_n2905 ), .ZN(_u10_u4_n3346 ) );
NAND2_X1 _u10_u4_U1242  ( .A1(_u10_u4_n3346 ), .A2(_u10_u4_n2803 ), .ZN(_u10_u4_n3345 ) );
NAND2_X1 _u10_u4_U1241  ( .A1(_u10_u4_n2087 ), .A2(_u10_u4_n2835 ), .ZN(_u10_u4_n2413 ) );
INV_X1 _u10_u4_U1240  ( .A(_u10_u4_n2128 ), .ZN(_u10_u4_n2235 ) );
NAND4_X1 _u10_u4_U1239  ( .A1(_u10_u4_n3344 ), .A2(_u10_u4_n3345 ), .A3(_u10_u4_n2413 ), .A4(_u10_u4_n2235 ), .ZN(_u10_u4_n3329 ) );
NOR2_X1 _u10_u4_U1238  ( .A1(_u10_u4_n1915 ), .A2(_u10_u4_n3340 ), .ZN(_u10_u4_n3343 ) );
NOR3_X1 _u10_u4_U1237  ( .A1(_u10_u4_n3329 ), .A2(1'b0), .A3(_u10_u4_n3343 ),.ZN(_u10_u4_n3341 ) );
NAND2_X1 _u10_u4_U1236  ( .A1(_u10_u4_n3342 ), .A2(_u10_u4_n3147 ), .ZN(_u10_u4_n2688 ) );
NOR2_X1 _u10_u4_U1235  ( .A1(_u10_u4_n3341 ), .A2(_u10_u4_n2688 ), .ZN(_u10_u4_n3335 ) );
NOR2_X1 _u10_u4_U1234  ( .A1(_u10_u4_n2256 ), .A2(_u10_u4_n1885 ), .ZN(_u10_u4_n2689 ) );
NOR2_X1 _u10_u4_U1233  ( .A1(1'b0), .A2(_u10_u4_n2413 ), .ZN(_u10_u4_n3338 ));
NOR2_X1 _u10_u4_U1232  ( .A1(_u10_u4_n1925 ), .A2(_u10_u4_n3340 ), .ZN(_u10_u4_n3339 ) );
NOR3_X1 _u10_u4_U1231  ( .A1(_u10_u4_n2005 ), .A2(_u10_u4_n3338 ), .A3(_u10_u4_n3339 ), .ZN(_u10_u4_n3337 ) );
NOR2_X1 _u10_u4_U1230  ( .A1(_u10_u4_n2689 ), .A2(_u10_u4_n3337 ), .ZN(_u10_u4_n3336 ) );
NOR3_X1 _u10_u4_U1229  ( .A1(_u10_u4_n3334 ), .A2(_u10_u4_n3335 ), .A3(_u10_u4_n3336 ), .ZN(_u10_u4_n3333 ) );
NAND4_X1 _u10_u4_U1228  ( .A1(_u10_u4_n3330 ), .A2(_u10_u4_n3331 ), .A3(_u10_u4_n3332 ), .A4(_u10_u4_n3333 ), .ZN(_u10_u4_n3308 ) );
NAND3_X1 _u10_u4_U1227  ( .A1(_u10_SYNOPSYS_UNCONNECTED_18 ), .A2(_u10_SYNOPSYS_UNCONNECTED_15 ), .A3(_u10_u4_n3147 ), .ZN(_u10_u4_n2126 ) );
INV_X1 _u10_u4_U1226  ( .A(_u10_u4_n2126 ), .ZN(_u10_u4_n2329 ) );
NAND2_X1 _u10_u4_U1225  ( .A1(_u10_u4_n2329 ), .A2(_u10_u4_n3329 ), .ZN(_u10_u4_n3324 ) );
NAND2_X1 _u10_u4_U1224  ( .A1(_u10_u4_n3328 ), .A2(_u10_u4_n3136 ), .ZN(_u10_u4_n2000 ) );
INV_X1 _u10_u4_U1223  ( .A(_u10_u4_n2000 ), .ZN(_u10_u4_n2445 ) );
NAND3_X1 _u10_u4_U1222  ( .A1(_u10_u4_n2446 ), .A2(_u10_u4_n3001 ), .A3(_u10_u4_n2087 ), .ZN(_u10_u4_n3327 ) );
NAND2_X1 _u10_u4_U1221  ( .A1(_u10_u4_n3327 ), .A2(_u10_u4_n2905 ), .ZN(_u10_u4_n2500 ) );
NAND2_X1 _u10_u4_U1220  ( .A1(_u10_u4_n2445 ), .A2(_u10_u4_n2500 ), .ZN(_u10_u4_n3325 ) );
NAND2_X1 _u10_u4_U1219  ( .A1(1'b0), .A2(_u10_u4_n2979 ), .ZN(_u10_u4_n3326 ) );
NAND3_X1 _u10_u4_U1218  ( .A1(_u10_u4_n3324 ), .A2(_u10_u4_n3325 ), .A3(_u10_u4_n3326 ), .ZN(_u10_u4_n3309 ) );
AND2_X1 _u10_u4_U1217  ( .A1(_u10_u4_n2877 ), .A2(_u10_u4_n3223 ), .ZN(_u10_u4_n2858 ) );
NAND2_X1 _u10_u4_U1216  ( .A1(_u10_u4_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_16 ), .ZN(_u10_u4_n2346 ) );
INV_X1 _u10_u4_U1215  ( .A(_u10_u4_n2346 ), .ZN(_u10_u4_n2043 ) );
NAND2_X1 _u10_u4_U1214  ( .A1(_u10_u4_n2858 ), .A2(_u10_u4_n2043 ), .ZN(_u10_u4_n3321 ) );
NAND2_X1 _u10_u4_U1213  ( .A1(_u10_u4_n1982 ), .A2(_u10_u4_n2195 ), .ZN(_u10_u4_n3268 ) );
INV_X1 _u10_u4_U1212  ( .A(_u10_u4_n3268 ), .ZN(_u10_u4_n2222 ) );
NAND3_X1 _u10_u4_U1211  ( .A1(_u10_u4_n3323 ), .A2(_u10_u4_n3216 ), .A3(_u10_u4_n2222 ), .ZN(_u10_u4_n3322 ) );
NAND2_X1 _u10_u4_U1210  ( .A1(_u10_u4_n3321 ), .A2(_u10_u4_n3322 ), .ZN(_u10_u4_n2374 ) );
NAND2_X1 _u10_u4_U1209  ( .A1(_u10_u4_n3320 ), .A2(_u10_u4_n3174 ), .ZN(_u10_u4_n2014 ) );
NOR2_X1 _u10_u4_U1208  ( .A1(_u10_u4_n1841 ), .A2(_u10_u4_n2014 ), .ZN(_u10_u4_n2813 ) );
NAND2_X1 _u10_u4_U1207  ( .A1(_u10_u4_n2813 ), .A2(_u10_u4_n2534 ), .ZN(_u10_u4_n3310 ) );
NAND2_X1 _u10_u4_U1206  ( .A1(_u10_u4_n3319 ), .A2(_u10_u4_n3136 ), .ZN(_u10_u4_n1836 ) );
INV_X1 _u10_u4_U1205  ( .A(_u10_u4_n1836 ), .ZN(_u10_u4_n2815 ) );
NAND2_X1 _u10_u4_U1204  ( .A1(_u10_u4_n2534 ), .A2(_u10_u4_n3129 ), .ZN(_u10_u4_n2439 ) );
NAND2_X1 _u10_u4_U1203  ( .A1(_u10_u4_n2055 ), .A2(_u10_u4_n2107 ), .ZN(_u10_u4_n2062 ) );
NAND2_X1 _u10_u4_U1202  ( .A1(_u10_u4_n2439 ), .A2(_u10_u4_n2062 ), .ZN(_u10_u4_n3318 ) );
NAND2_X1 _u10_u4_U1201  ( .A1(_u10_u4_n2815 ), .A2(_u10_u4_n3318 ), .ZN(_u10_u4_n3311 ) );
NAND2_X1 _u10_u4_U1200  ( .A1(_u10_u4_n2986 ), .A2(_u10_u4_n2175 ), .ZN(_u10_u4_n3317 ) );
NAND2_X1 _u10_u4_U1199  ( .A1(_u10_u4_n2253 ), .A2(_u10_u4_n3317 ), .ZN(_u10_u4_n3157 ) );
NAND2_X1 _u10_u4_U1198  ( .A1(_u10_u4_n3316 ), .A2(_u10_u4_n3157 ), .ZN(_u10_u4_n3312 ) );
NOR2_X1 _u10_u4_U1197  ( .A1(_u10_u4_n2495 ), .A2(_u10_u4_n2194 ), .ZN(_u10_u4_n3314 ) );
NOR2_X1 _u10_u4_U1196  ( .A1(_u10_u4_n2375 ), .A2(_u10_u4_n2367 ), .ZN(_u10_u4_n3315 ) );
NOR2_X1 _u10_u4_U1195  ( .A1(_u10_u4_n3314 ), .A2(_u10_u4_n3315 ), .ZN(_u10_u4_n3313 ) );
NAND4_X1 _u10_u4_U1194  ( .A1(_u10_u4_n3310 ), .A2(_u10_u4_n3311 ), .A3(_u10_u4_n3312 ), .A4(_u10_u4_n3313 ), .ZN(_u10_u4_n2315 ) );
NOR4_X1 _u10_u4_U1193  ( .A1(_u10_u4_n3308 ), .A2(_u10_u4_n3309 ), .A3(_u10_u4_n2374 ), .A4(_u10_u4_n2315 ), .ZN(_u10_u4_n3307 ) );
NAND3_X1 _u10_u4_U1192  ( .A1(_u10_u4_n3305 ), .A2(_u10_u4_n3306 ), .A3(_u10_u4_n3307 ), .ZN(_u10_u4_n1987 ) );
AND2_X1 _u10_u4_U1191  ( .A1(1'b0), .A2(_u10_u4_n2977 ), .ZN(_u10_u4_n3240 ));
NAND2_X1 _u10_u4_U1190  ( .A1(_u10_u4_n1891 ), .A2(_u10_u4_n2534 ), .ZN(_u10_u4_n3303 ) );
NAND4_X1 _u10_u4_U1189  ( .A1(_u10_u4_n1982 ), .A2(_u10_u4_n2659 ), .A3(_u10_u4_n2256 ), .A4(_u10_u4_n2175 ), .ZN(_u10_u4_n3304 ) );
AND2_X1 _u10_u4_U1188  ( .A1(_u10_u4_n3303 ), .A2(_u10_u4_n3304 ), .ZN(_u10_u4_n2612 ) );
NAND2_X1 _u10_u4_U1187  ( .A1(_u10_u4_n3302 ), .A2(_u10_u4_n3236 ), .ZN(_u10_u4_n2985 ) );
OR2_X1 _u10_u4_U1186  ( .A1(_u10_u4_n2431 ), .A2(_u10_u4_n2985 ), .ZN(_u10_u4_n3299 ) );
OR2_X1 _u10_u4_U1185  ( .A1(_u10_u4_n2282 ), .A2(_u10_u4_n2359 ), .ZN(_u10_u4_n3300 ) );
NAND2_X1 _u10_u4_U1184  ( .A1(_u10_u4_n1890 ), .A2(_u10_u4_n2534 ), .ZN(_u10_u4_n3301 ) );
NAND4_X1 _u10_u4_U1183  ( .A1(_u10_u4_n2612 ), .A2(_u10_u4_n3299 ), .A3(_u10_u4_n3300 ), .A4(_u10_u4_n3301 ), .ZN(_u10_u4_n3279 ) );
INV_X1 _u10_u4_U1182  ( .A(_u10_u4_n2464 ), .ZN(_u10_u4_n3295 ) );
NAND2_X1 _u10_u4_U1181  ( .A1(_u10_u4_n3295 ), .A2(_u10_u4_n2835 ), .ZN(_u10_u4_n2623 ) );
INV_X1 _u10_u4_U1180  ( .A(_u10_u4_n2623 ), .ZN(_u10_u4_n3185 ) );
INV_X1 _u10_u4_U1179  ( .A(_u10_u4_n2688 ), .ZN(_u10_u4_n2169 ) );
NAND2_X1 _u10_u4_U1178  ( .A1(_u10_u4_n3185 ), .A2(_u10_u4_n2169 ), .ZN(_u10_u4_n3286 ) );
NAND2_X1 _u10_u4_U1177  ( .A1(_u10_u4_n2833 ), .A2(_u10_u4_n3278 ), .ZN(_u10_u4_n3298 ) );
NAND3_X1 _u10_u4_U1176  ( .A1(_u10_u4_n3297 ), .A2(_u10_u4_n2838 ), .A3(_u10_u4_n3298 ), .ZN(_u10_u4_n3296 ) );
NAND2_X1 _u10_u4_U1175  ( .A1(_u10_u4_n2830 ), .A2(_u10_u4_n3296 ), .ZN(_u10_u4_n3287 ) );
NAND2_X1 _u10_u4_U1174  ( .A1(_u10_u4_n3295 ), .A2(_u10_u4_n3001 ), .ZN(_u10_u4_n3292 ) );
NAND2_X1 _u10_u4_U1173  ( .A1(_u10_u4_n3294 ), .A2(_u10_u4_n2089 ), .ZN(_u10_u4_n3293 ) );
AND2_X1 _u10_u4_U1172  ( .A1(_u10_u4_n3292 ), .A2(_u10_u4_n3293 ), .ZN(_u10_u4_n2548 ) );
NAND2_X1 _u10_u4_U1171  ( .A1(_u10_u4_n2548 ), .A2(_u10_u4_n2091 ), .ZN(_u10_u4_n2304 ) );
NAND2_X1 _u10_u4_U1170  ( .A1(_u10_u4_n2304 ), .A2(_u10_u4_n2446 ), .ZN(_u10_u4_n3290 ) );
NAND2_X1 _u10_u4_U1169  ( .A1(_u10_u4_n2549 ), .A2(_u10_u4_n2446 ), .ZN(_u10_u4_n2790 ) );
NOR2_X1 _u10_u4_U1168  ( .A1(_u10_u4_n1936 ), .A2(_u10_u4_n2790 ), .ZN(_u10_u4_n2789 ) );
INV_X1 _u10_u4_U1167  ( .A(_u10_u4_n2789 ), .ZN(_u10_u4_n3291 ) );
OR2_X1 _u10_u4_U1166  ( .A1(_u10_u4_n2828 ), .A2(_u10_u4_n2790 ), .ZN(_u10_u4_n2498 ) );
NAND4_X1 _u10_u4_U1165  ( .A1(_u10_u4_n3290 ), .A2(_u10_u4_n3291 ), .A3(_u10_u4_n2498 ), .A4(_u10_u4_n2001 ), .ZN(_u10_u4_n3289 ) );
NAND2_X1 _u10_u4_U1164  ( .A1(_u10_u4_n2445 ), .A2(_u10_u4_n3289 ), .ZN(_u10_u4_n3288 ) );
NAND3_X1 _u10_u4_U1163  ( .A1(_u10_u4_n3286 ), .A2(_u10_u4_n3287 ), .A3(_u10_u4_n3288 ), .ZN(_u10_u4_n3280 ) );
NOR2_X1 _u10_u4_U1162  ( .A1(_u10_u4_n2940 ), .A2(_u10_u4_n1913 ), .ZN(_u10_u4_n3281 ) );
INV_X1 _u10_u4_U1161  ( .A(1'b0), .ZN(_u10_u4_n1864 ) );
NAND2_X1 _u10_u4_U1160  ( .A1(1'b0), .A2(_u10_u4_n2588 ), .ZN(_u10_u4_n2141 ) );
INV_X1 _u10_u4_U1159  ( .A(_u10_u4_n2141 ), .ZN(_u10_u4_n3159 ) );
NAND3_X1 _u10_u4_U1158  ( .A1(_u10_u4_n2103 ), .A2(_u10_u4_n1864 ), .A3(_u10_u4_n3159 ), .ZN(_u10_u4_n2520 ) );
INV_X1 _u10_u4_U1157  ( .A(_u10_u4_n2520 ), .ZN(_u10_u4_n2630 ) );
INV_X1 _u10_u4_U1156  ( .A(_u10_u4_n2307 ), .ZN(_u10_u4_n2382 ) );
NOR4_X1 _u10_u4_U1155  ( .A1(_u10_u4_n2382 ), .A2(_u10_u4_n2722 ), .A3(_u10_u4_n1925 ), .A4(_u10_u4_n2508 ), .ZN(_u10_u4_n3260 ) );
NOR2_X1 _u10_u4_U1154  ( .A1(_u10_u4_n2498 ), .A2(_u10_u4_n2911 ), .ZN(_u10_u4_n2633 ) );
NOR2_X1 _u10_u4_U1153  ( .A1(_u10_u4_n2633 ), .A2(_u10_u4_n3278 ), .ZN(_u10_u4_n3285 ) );
INV_X1 _u10_u4_U1152  ( .A(_u10_u4_n1866 ), .ZN(_u10_u4_n1926 ) );
NOR2_X1 _u10_u4_U1151  ( .A1(_u10_u4_n3285 ), .A2(_u10_u4_n1926 ), .ZN(_u10_u4_n3284 ) );
NOR4_X1 _u10_u4_U1150  ( .A1(1'b0), .A2(_u10_u4_n2630 ), .A3(_u10_u4_n3260 ),.A4(_u10_u4_n3284 ), .ZN(_u10_u4_n3283 ) );
NOR2_X1 _u10_u4_U1149  ( .A1(_u10_u4_n3283 ), .A2(_u10_u4_n2980 ), .ZN(_u10_u4_n3282 ) );
NOR4_X1 _u10_u4_U1148  ( .A1(_u10_u4_n3279 ), .A2(_u10_u4_n3280 ), .A3(_u10_u4_n3281 ), .A4(_u10_u4_n3282 ), .ZN(_u10_u4_n3241 ) );
NAND2_X1 _u10_u4_U1147  ( .A1(_u10_u4_n1836 ), .A2(_u10_u4_n2291 ), .ZN(_u10_u4_n2147 ) );
NAND2_X1 _u10_u4_U1146  ( .A1(_u10_u4_n2443 ), .A2(_u10_u4_n2147 ), .ZN(_u10_u4_n3261 ) );
INV_X1 _u10_u4_U1145  ( .A(_u10_u4_n1841 ), .ZN(_u10_u4_n2571 ) );
NAND2_X1 _u10_u4_U1144  ( .A1(_u10_u4_n2571 ), .A2(_u10_u4_n3278 ), .ZN(_u10_u4_n3277 ) );
NAND2_X1 _u10_u4_U1143  ( .A1(_u10_u4_n3276 ), .A2(_u10_u4_n3277 ), .ZN(_u10_u4_n2819 ) );
OR2_X1 _u10_u4_U1142  ( .A1(_u10_u4_n2819 ), .A2(_u10_u4_n3275 ), .ZN(_u10_u4_n3273 ) );
NAND2_X1 _u10_u4_U1141  ( .A1(_u10_u4_n2815 ), .A2(_u10_u4_n2080 ), .ZN(_u10_u4_n3274 ) );
NAND2_X1 _u10_u4_U1140  ( .A1(_u10_u4_n2014 ), .A2(_u10_u4_n3274 ), .ZN(_u10_u4_n2165 ) );
NAND2_X1 _u10_u4_U1139  ( .A1(_u10_u4_n3273 ), .A2(_u10_u4_n2165 ), .ZN(_u10_u4_n3262 ) );
NAND2_X1 _u10_u4_U1138  ( .A1(_u10_u4_n2688 ), .A2(_u10_u4_n2126 ), .ZN(_u10_u4_n1956 ) );
INV_X1 _u10_u4_U1137  ( .A(_u10_u4_n1956 ), .ZN(_u10_u4_n1860 ) );
NOR2_X1 _u10_u4_U1136  ( .A1(1'b0), .A2(_u10_u4_n2498 ), .ZN(_u10_u4_n3271 ));
NOR2_X1 _u10_u4_U1135  ( .A1(_u10_u4_n3271 ), .A2(_u10_u4_n3272 ), .ZN(_u10_u4_n3270 ) );
NOR2_X1 _u10_u4_U1134  ( .A1(_u10_u4_n1860 ), .A2(_u10_u4_n3270 ), .ZN(_u10_u4_n3264 ) );
INV_X1 _u10_u4_U1133  ( .A(_u10_u4_n2632 ), .ZN(_u10_u4_n3202 ) );
NAND2_X1 _u10_u4_U1132  ( .A1(_u10_u4_n3236 ), .A2(_u10_u4_n3269 ), .ZN(_u10_u4_n3036 ) );
INV_X1 _u10_u4_U1131  ( .A(_u10_u4_n3036 ), .ZN(_u10_u4_n1960 ) );
NAND2_X1 _u10_u4_U1130  ( .A1(_u10_u4_n3202 ), .A2(_u10_u4_n1960 ), .ZN(_u10_u4_n3079 ) );
NOR3_X1 _u10_u4_U1129  ( .A1(_u10_u4_n3079 ), .A2(1'b0), .A3(_u10_u4_n3268 ),.ZN(_u10_u4_n3265 ) );
INV_X1 _u10_u4_U1128  ( .A(_u10_u4_n2014 ), .ZN(_u10_u4_n2709 ) );
NAND2_X1 _u10_u4_U1127  ( .A1(_u10_u4_n2709 ), .A2(_u10_u4_n2166 ), .ZN(_u10_u4_n2145 ) );
INV_X1 _u10_u4_U1126  ( .A(_u10_u4_n2145 ), .ZN(_u10_u4_n3258 ) );
NOR2_X1 _u10_u4_U1125  ( .A1(_u10_u4_n3258 ), .A2(_u10_u4_n2183 ), .ZN(_u10_u4_n3267 ) );
NOR2_X1 _u10_u4_U1124  ( .A1(_u10_u4_n3267 ), .A2(_u10_u4_n2567 ), .ZN(_u10_u4_n3266 ) );
NOR3_X1 _u10_u4_U1123  ( .A1(_u10_u4_n3264 ), .A2(_u10_u4_n3265 ), .A3(_u10_u4_n3266 ), .ZN(_u10_u4_n3263 ) );
NAND3_X1 _u10_u4_U1122  ( .A1(_u10_u4_n3261 ), .A2(_u10_u4_n3262 ), .A3(_u10_u4_n3263 ), .ZN(_u10_u4_n3243 ) );
INV_X1 _u10_u4_U1121  ( .A(_u10_u4_n2102 ), .ZN(_u10_u4_n2509 ) );
NAND2_X1 _u10_u4_U1120  ( .A1(_u10_u4_n3260 ), .A2(_u10_u4_n2509 ), .ZN(_u10_u4_n3247 ) );
INV_X1 _u10_u4_U1119  ( .A(_u10_u4_n3259 ), .ZN(_u10_u4_n2015 ) );
NAND2_X1 _u10_u4_U1118  ( .A1(_u10_u4_n2015 ), .A2(_u10_u4_n3258 ), .ZN(_u10_u4_n3248 ) );
NAND2_X1 _u10_u4_U1117  ( .A1(_u10_u4_n2251 ), .A2(_u10_u4_n2169 ), .ZN(_u10_u4_n3255 ) );
OR2_X1 _u10_u4_U1116  ( .A1(_u10_u4_n3157 ), .A2(_u10_u4_n2256 ), .ZN(_u10_u4_n3257 ) );
NAND2_X1 _u10_u4_U1115  ( .A1(_u10_u4_n2105 ), .A2(_u10_u4_n3257 ), .ZN(_u10_u4_n3256 ) );
AND2_X1 _u10_u4_U1114  ( .A1(_u10_u4_n3255 ), .A2(_u10_u4_n3256 ), .ZN(_u10_u4_n3212 ) );
INV_X1 _u10_u4_U1113  ( .A(_u10_u4_n2037 ), .ZN(_u10_u4_n2987 ) );
NAND2_X1 _u10_u4_U1112  ( .A1(_u10_u4_n2987 ), .A2(_u10_u4_n2038 ), .ZN(_u10_u4_n2212 ) );
NOR2_X1 _u10_u4_U1111  ( .A1(_u10_u4_n2212 ), .A2(1'b0), .ZN(_u10_u4_n2658 ));
INV_X1 _u10_u4_U1110  ( .A(_u10_u4_n2658 ), .ZN(_u10_u4_n2343 ) );
NAND2_X1 _u10_u4_U1109  ( .A1(_u10_u4_n2344 ), .A2(_u10_u4_n3254 ), .ZN(_u10_u4_n1928 ) );
NAND2_X1 _u10_u4_U1108  ( .A1(_u10_u4_n2588 ), .A2(_u10_u4_n1928 ), .ZN(_u10_u4_n3253 ) );
NAND2_X1 _u10_u4_U1107  ( .A1(_u10_u4_n2343 ), .A2(_u10_u4_n3253 ), .ZN(_u10_u4_n3252 ) );
NAND2_X1 _u10_u4_U1106  ( .A1(_u10_u4_n2105 ), .A2(_u10_u4_n3252 ), .ZN(_u10_u4_n3251 ) );
NAND2_X1 _u10_u4_U1105  ( .A1(_u10_u4_n3212 ), .A2(_u10_u4_n3251 ), .ZN(_u10_u4_n3250 ) );
NAND2_X1 _u10_u4_U1104  ( .A1(_u10_u4_n2307 ), .A2(_u10_u4_n3250 ), .ZN(_u10_u4_n3249 ) );
NAND3_X1 _u10_u4_U1103  ( .A1(_u10_u4_n3247 ), .A2(_u10_u4_n3248 ), .A3(_u10_u4_n3249 ), .ZN(_u10_u4_n3244 ) );
AND2_X1 _u10_u4_U1102  ( .A1(_u10_u4_n2915 ), .A2(_u10_u4_n2059 ), .ZN(_u10_u4_n2957 ) );
AND3_X1 _u10_u4_U1101  ( .A1(_u10_u4_n3223 ), .A2(_u10_u4_n2837 ), .A3(_u10_u4_n2957 ), .ZN(_u10_u4_n2051 ) );
NOR2_X1 _u10_u4_U1100  ( .A1(_u10_u4_n2528 ), .A2(_u10_u4_n2051 ), .ZN(_u10_u4_n2605 ) );
NOR2_X1 _u10_u4_U1099  ( .A1(_u10_u4_n2605 ), .A2(_u10_u4_n2346 ), .ZN(_u10_u4_n3245 ) );
NOR2_X1 _u10_u4_U1098  ( .A1(_u10_u4_n2291 ), .A2(_u10_u4_n2062 ), .ZN(_u10_u4_n3246 ) );
NOR4_X1 _u10_u4_U1097  ( .A1(_u10_u4_n3243 ), .A2(_u10_u4_n3244 ), .A3(_u10_u4_n3245 ), .A4(_u10_u4_n3246 ), .ZN(_u10_u4_n3242 ) );
NAND2_X1 _u10_u4_U1096  ( .A1(_u10_u4_n3241 ), .A2(_u10_u4_n3242 ), .ZN(_u10_u4_n2311 ) );
OR3_X1 _u10_u4_U1095  ( .A1(_u10_u4_n1987 ), .A2(_u10_u4_n3240 ), .A3(_u10_u4_n2311 ), .ZN(_u10_u4_n3192 ) );
INV_X1 _u10_u4_U1094  ( .A(_u10_u4_n2886 ), .ZN(_u10_u4_n2720 ) );
NOR2_X1 _u10_u4_U1093  ( .A1(_u10_u4_n2004 ), .A2(_u10_u4_n2720 ), .ZN(_u10_u4_n2455 ) );
INV_X1 _u10_u4_U1092  ( .A(_u10_u4_n2488 ), .ZN(_u10_u4_n2938 ) );
AND3_X1 _u10_u4_U1091  ( .A1(_u10_u4_n2455 ), .A2(_u10_u4_n1859 ), .A3(_u10_u4_n2938 ), .ZN(_u10_u4_n3239 ) );
INV_X1 _u10_u4_U1090  ( .A(_u10_u4_n2633 ), .ZN(_u10_u4_n2937 ) );
NOR2_X1 _u10_u4_U1089  ( .A1(_u10_u4_n3239 ), .A2(_u10_u4_n2937 ), .ZN(_u10_u4_n3227 ) );
NOR2_X1 _u10_u4_U1088  ( .A1(_u10_u4_n1976 ), .A2(_u10_u4_n1969 ), .ZN(_u10_u4_n3237 ) );
NOR2_X1 _u10_u4_U1087  ( .A1(1'b0), .A2(_u10_u4_n2947 ), .ZN(_u10_u4_n3238 ));
NOR3_X1 _u10_u4_U1086  ( .A1(_u10_u4_n2476 ), .A2(_u10_u4_n3237 ), .A3(_u10_u4_n3238 ), .ZN(_u10_u4_n3235 ) );
NOR3_X1 _u10_u4_U1085  ( .A1(_u10_u4_n1813 ), .A2(_u10_u4_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_15 ), .ZN(_u10_u4_n3135 ) );
NAND2_X1 _u10_u4_U1084  ( .A1(_u10_u4_n3135 ), .A2(_u10_u4_n3236 ), .ZN(_u10_u4_n2573 ) );
NOR2_X1 _u10_u4_U1083  ( .A1(_u10_u4_n3235 ), .A2(_u10_u4_n2573 ), .ZN(_u10_u4_n3228 ) );
NOR2_X1 _u10_u4_U1082  ( .A1(_u10_u4_n2216 ), .A2(_u10_u4_n1868 ), .ZN(_u10_u4_n3233 ) );
INV_X1 _u10_u4_U1081  ( .A(_u10_u4_n2550 ), .ZN(_u10_u4_n2475 ) );
NOR3_X1 _u10_u4_U1080  ( .A1(_u10_u4_n2475 ), .A2(1'b0), .A3(_u10_u4_n1925 ),.ZN(_u10_u4_n3234 ) );
NOR3_X1 _u10_u4_U1079  ( .A1(_u10_u4_n3233 ), .A2(1'b0), .A3(_u10_u4_n3234 ),.ZN(_u10_u4_n3232 ) );
NOR2_X1 _u10_u4_U1078  ( .A1(_u10_u4_n3232 ), .A2(_u10_u4_n2037 ), .ZN(_u10_u4_n3229 ) );
NOR2_X1 _u10_u4_U1077  ( .A1(_u10_u4_n3231 ), .A2(_u10_u4_n2365 ), .ZN(_u10_u4_n3230 ) );
NOR4_X1 _u10_u4_U1076  ( .A1(_u10_u4_n3227 ), .A2(_u10_u4_n3228 ), .A3(_u10_u4_n3229 ), .A4(_u10_u4_n3230 ), .ZN(_u10_u4_n3205 ) );
NOR3_X1 _u10_u4_U1075  ( .A1(_u10_u4_n3226 ), .A2(_u10_u4_n2687 ), .A3(_u10_u4_n2145 ), .ZN(_u10_u4_n3217 ) );
NOR3_X1 _u10_u4_U1074  ( .A1(_u10_u4_n3225 ), .A2(1'b0), .A3(_u10_u4_n2587 ),.ZN(_u10_u4_n3218 ) );
NOR2_X1 _u10_u4_U1073  ( .A1(_u10_u4_n3159 ), .A2(1'b0), .ZN(_u10_u4_n3224 ));
NOR2_X1 _u10_u4_U1072  ( .A1(_u10_u4_n3224 ), .A2(_u10_u4_n2584 ), .ZN(_u10_u4_n3219 ) );
NAND2_X1 _u10_u4_U1071  ( .A1(_u10_u4_n3222 ), .A2(_u10_u4_n3223 ), .ZN(_u10_u4_n2048 ) );
INV_X1 _u10_u4_U1070  ( .A(_u10_u4_n2048 ), .ZN(_u10_u4_n2859 ) );
NOR2_X1 _u10_u4_U1069  ( .A1(_u10_u4_n2859 ), .A2(_u10_u4_n2054 ), .ZN(_u10_u4_n3221 ) );
NOR2_X1 _u10_u4_U1068  ( .A1(_u10_u4_n3221 ), .A2(_u10_u4_n2346 ), .ZN(_u10_u4_n3220 ) );
NOR4_X1 _u10_u4_U1067  ( .A1(_u10_u4_n3217 ), .A2(_u10_u4_n3218 ), .A3(_u10_u4_n3219 ), .A4(_u10_u4_n3220 ), .ZN(_u10_u4_n3206 ) );
NAND2_X1 _u10_u4_U1066  ( .A1(_u10_u4_n2377 ), .A2(_u10_u4_n2721 ), .ZN(_u10_u4_n3213 ) );
AND4_X1 _u10_u4_U1065  ( .A1(1'b0), .A2(_u10_u4_n2502 ), .A3(_u10_u4_n2972 ),.A4(_u10_u4_n3040 ), .ZN(_u10_u4_n2406 ) );
NAND2_X1 _u10_u4_U1064  ( .A1(_u10_u4_n2406 ), .A2(_u10_u4_n2979 ), .ZN(_u10_u4_n3214 ) );
NAND2_X1 _u10_u4_U1063  ( .A1(_u10_u4_n2630 ), .A2(_u10_u4_n3216 ), .ZN(_u10_u4_n2376 ) );
INV_X1 _u10_u4_U1062  ( .A(_u10_u4_n2376 ), .ZN(_u10_u4_n3108 ) );
NAND2_X1 _u10_u4_U1061  ( .A1(_u10_u4_n3108 ), .A2(_u10_u4_n2507 ), .ZN(_u10_u4_n3215 ) );
NOR2_X1 _u10_u4_U1060  ( .A1(_u10_u4_n2937 ), .A2(1'b0), .ZN(_u10_u4_n2649 ));
INV_X1 _u10_u4_U1059  ( .A(_u10_u4_n2253 ), .ZN(_u10_u4_n2971 ) );
NAND2_X1 _u10_u4_U1058  ( .A1(_u10_u4_n2649 ), .A2(_u10_u4_n2971 ), .ZN(_u10_u4_n2918 ) );
NAND4_X1 _u10_u4_U1057  ( .A1(_u10_u4_n3213 ), .A2(_u10_u4_n3214 ), .A3(_u10_u4_n3215 ), .A4(_u10_u4_n2918 ), .ZN(_u10_u4_n3208 ) );
NOR2_X1 _u10_u4_U1056  ( .A1(_u10_u4_n2000 ), .A2(_u10_u4_n2902 ), .ZN(_u10_u4_n3209 ) );
NOR2_X1 _u10_u4_U1055  ( .A1(_u10_u4_n3212 ), .A2(_u10_u4_n2475 ), .ZN(_u10_u4_n3210 ) );
INV_X1 _u10_u4_U1054  ( .A(_u10_u4_n2441 ), .ZN(_u10_u4_n3128 ) );
NOR2_X1 _u10_u4_U1053  ( .A1(_u10_u4_n2356 ), .A2(_u10_u4_n3128 ), .ZN(_u10_u4_n3211 ) );
NOR4_X1 _u10_u4_U1052  ( .A1(_u10_u4_n3208 ), .A2(_u10_u4_n3209 ), .A3(_u10_u4_n3210 ), .A4(_u10_u4_n3211 ), .ZN(_u10_u4_n3207 ) );
NAND3_X1 _u10_u4_U1051  ( .A1(_u10_u4_n3205 ), .A2(_u10_u4_n3206 ), .A3(_u10_u4_n3207 ), .ZN(_u10_u4_n2611 ) );
NOR2_X1 _u10_u4_U1050  ( .A1(_u10_u4_n2212 ), .A2(_u10_u4_n2216 ), .ZN(_u10_u4_n1937 ) );
NOR2_X1 _u10_u4_U1049  ( .A1(_u10_u4_n2533 ), .A2(_u10_u4_n2214 ), .ZN(_u10_u4_n2765 ) );
INV_X1 _u10_u4_U1048  ( .A(_u10_u4_n2005 ), .ZN(_u10_u4_n2111 ) );
AND2_X1 _u10_u4_U1047  ( .A1(_u10_u4_n2765 ), .A2(_u10_u4_n2111 ), .ZN(_u10_u4_n3201 ) );
INV_X1 _u10_u4_U1046  ( .A(_u10_u4_n3059 ), .ZN(_u10_u4_n3076 ) );
NAND2_X1 _u10_u4_U1045  ( .A1(_u10_u4_n3201 ), .A2(_u10_u4_n3076 ), .ZN(_u10_u4_n3204 ) );
NAND2_X1 _u10_u4_U1044  ( .A1(_u10_u4_n1937 ), .A2(_u10_u4_n3204 ), .ZN(_u10_u4_n3193 ) );
NAND2_X1 _u10_u4_U1043  ( .A1(_u10_u4_n2254 ), .A2(_u10_u4_n2212 ), .ZN(_u10_u4_n3203 ) );
NAND3_X1 _u10_u4_U1042  ( .A1(_u10_u4_n3203 ), .A2(_u10_u4_n2175 ), .A3(_u10_u4_n2649 ), .ZN(_u10_u4_n3194 ) );
NOR2_X1 _u10_u4_U1041  ( .A1(_u10_u4_n2985 ), .A2(1'b0), .ZN(_u10_u4_n1959 ));
NAND2_X1 _u10_u4_U1040  ( .A1(_u10_u4_n1959 ), .A2(_u10_u4_n3202 ), .ZN(_u10_u4_n2202 ) );
NAND4_X1 _u10_u4_U1039  ( .A1(_u10_u4_n3079 ), .A2(_u10_u4_n2621 ), .A3(_u10_u4_n2202 ), .A4(_u10_u4_n2798 ), .ZN(_u10_u4_n3200 ) );
NAND2_X1 _u10_u4_U1038  ( .A1(_u10_u4_n3201 ), .A2(_u10_u4_n2937 ), .ZN(_u10_u4_n2772 ) );
NAND2_X1 _u10_u4_U1037  ( .A1(_u10_u4_n3200 ), .A2(_u10_u4_n2772 ), .ZN(_u10_u4_n3195 ) );
NAND2_X1 _u10_u4_U1036  ( .A1(_u10_u4_n2765 ), .A2(_u10_u4_n1869 ), .ZN(_u10_u4_n3199 ) );
NAND2_X1 _u10_u4_U1035  ( .A1(_u10_u4_n2049 ), .A2(_u10_u4_n3199 ), .ZN(_u10_u4_n3057 ) );
NOR2_X1 _u10_u4_U1034  ( .A1(_u10_u4_n2495 ), .A2(_u10_u4_n3057 ), .ZN(_u10_u4_n3197 ) );
NOR2_X1 _u10_u4_U1033  ( .A1(_u10_u4_n2883 ), .A2(_u10_u4_n2485 ), .ZN(_u10_u4_n3198 ) );
NOR2_X1 _u10_u4_U1032  ( .A1(_u10_u4_n3197 ), .A2(_u10_u4_n3198 ), .ZN(_u10_u4_n3196 ) );
NAND4_X1 _u10_u4_U1031  ( .A1(_u10_u4_n3193 ), .A2(_u10_u4_n3194 ), .A3(_u10_u4_n3195 ), .A4(_u10_u4_n3196 ), .ZN(_u10_u4_n2887 ) );
NOR4_X1 _u10_u4_U1030  ( .A1(_u10_u4_n3191 ), .A2(_u10_u4_n3192 ), .A3(_u10_u4_n2611 ), .A4(_u10_u4_n2887 ), .ZN(_u10_u4_n3015 ) );
NAND3_X1 _u10_u4_U1029  ( .A1(_u10_u4_n3190 ), .A2(_u10_u4_n2049 ), .A3(_u10_u4_n2957 ), .ZN(_u10_u4_n2699 ) );
OR2_X1 _u10_u4_U1028  ( .A1(_u10_u4_n2699 ), .A2(_u10_u4_n1813 ), .ZN(_u10_u4_n3187 ) );
NAND3_X1 _u10_u4_U1027  ( .A1(_u10_u4_n2978 ), .A2(_u10_u4_n2405 ), .A3(1'b0), .ZN(_u10_u4_n3188 ) );
NAND4_X1 _u10_u4_U1026  ( .A1(_u10_u4_n3058 ), .A2(_u10_u4_n3187 ), .A3(_u10_u4_n3188 ), .A4(_u10_u4_n3189 ), .ZN(_u10_u4_n3186 ) );
NAND2_X1 _u10_u4_U1025  ( .A1(_u10_u4_n2063 ), .A2(_u10_u4_n3186 ), .ZN(_u10_u4_n3163 ) );
NAND2_X1 _u10_u4_U1024  ( .A1(_u10_u4_n3185 ), .A2(_u10_u4_n2329 ), .ZN(_u10_u4_n3164 ) );
NAND2_X1 _u10_u4_U1023  ( .A1(_u10_u4_n2689 ), .A2(_u10_u4_n2365 ), .ZN(_u10_u4_n2736 ) );
NOR2_X1 _u10_u4_U1022  ( .A1(_u10_u4_n2736 ), .A2(_u10_u4_n2488 ), .ZN(_u10_u4_n1855 ) );
INV_X1 _u10_u4_U1021  ( .A(_u10_u4_n1855 ), .ZN(_u10_u4_n3184 ) );
NOR2_X1 _u10_u4_U1020  ( .A1(_u10_u4_n2274 ), .A2(_u10_u4_n2359 ), .ZN(_u10_u4_n2952 ) );
NOR2_X1 _u10_u4_U1019  ( .A1(_u10_u4_n3184 ), .A2(_u10_u4_n2952 ), .ZN(_u10_u4_n2776 ) );
OR2_X1 _u10_u4_U1018  ( .A1(_u10_u4_n2852 ), .A2(_u10_u4_n2776 ), .ZN(_u10_u4_n3165 ) );
NAND2_X1 _u10_u4_U1017  ( .A1(_u10_u4_n3126 ), .A2(_u10_u4_n2915 ), .ZN(_u10_u4_n3065 ) );
NOR3_X1 _u10_u4_U1016  ( .A1(_u10_u4_n3065 ), .A2(1'b0), .A3(_u10_u4_n2632 ),.ZN(_u10_u4_n3182 ) );
NOR3_X1 _u10_u4_U1015  ( .A1(_u10_u4_n3182 ), .A2(_u10_u4_n3183 ), .A3(_u10_u4_n3108 ), .ZN(_u10_u4_n3181 ) );
NOR2_X1 _u10_u4_U1014  ( .A1(_u10_u4_n3181 ), .A2(_u10_u4_n3162 ), .ZN(_u10_u4_n3167 ) );
INV_X1 _u10_u4_U1013  ( .A(_u10_u4_n3180 ), .ZN(_u10_u4_n3140 ) );
NAND3_X1 _u10_u4_U1012  ( .A1(_u10_u4_n3140 ), .A2(_u10_u4_n2163 ), .A3(_u10_u4_n2092 ), .ZN(_u10_u4_n3175 ) );
NOR4_X1 _u10_u4_U1011  ( .A1(_u10_u4_n2411 ), .A2(_u10_u4_n2710 ), .A3(_u10_u4_n3141 ), .A4(_u10_u4_n3089 ), .ZN(_u10_u4_n3179 ) );
NOR2_X1 _u10_u4_U1010  ( .A1(1'b0), .A2(_u10_u4_n3179 ), .ZN(_u10_u4_n3177 ));
NOR2_X1 _u10_u4_U1009  ( .A1(_u10_u4_n1898 ), .A2(_u10_u4_n1847 ), .ZN(_u10_u4_n3178 ) );
NOR4_X1 _u10_u4_U1008  ( .A1(_u10_u4_n3175 ), .A2(_u10_u4_n3176 ), .A3(_u10_u4_n3177 ), .A4(_u10_u4_n3178 ), .ZN(_u10_u4_n3173 ) );
NAND2_X1 _u10_u4_U1007  ( .A1(_u10_u4_n3135 ), .A2(_u10_u4_n3174 ), .ZN(_u10_u4_n2159 ) );
NOR2_X1 _u10_u4_U1006  ( .A1(_u10_u4_n3173 ), .A2(_u10_u4_n2159 ), .ZN(_u10_u4_n3168 ) );
OR3_X1 _u10_u4_U1005  ( .A1(_u10_u4_n3172 ), .A2(1'b0), .A3(_u10_u4_n3126 ),.ZN(_u10_u4_n3171 ) );
NAND2_X1 _u10_u4_U1004  ( .A1(_u10_u4_n2600 ), .A2(_u10_u4_n3171 ), .ZN(_u10_u4_n3153 ) );
AND3_X1 _u10_u4_U1003  ( .A1(_u10_u4_n3153 ), .A2(_u10_u4_n2947 ), .A3(_u10_u4_n2579 ), .ZN(_u10_u4_n3170 ) );
NOR2_X1 _u10_u4_U1002  ( .A1(_u10_u4_n3170 ), .A2(_u10_u4_n2359 ), .ZN(_u10_u4_n3169 ) );
NOR3_X1 _u10_u4_U1001  ( .A1(_u10_u4_n3167 ), .A2(_u10_u4_n3168 ), .A3(_u10_u4_n3169 ), .ZN(_u10_u4_n3166 ) );
NAND4_X1 _u10_u4_U1000  ( .A1(_u10_u4_n3163 ), .A2(_u10_u4_n3164 ), .A3(_u10_u4_n3165 ), .A4(_u10_u4_n3166 ), .ZN(_u10_u4_n3130 ) );
NAND2_X1 _u10_u4_U999  ( .A1(_u10_u4_n2375 ), .A2(_u10_u4_n3162 ), .ZN(_u10_u4_n1923 ) );
NAND2_X1 _u10_u4_U998  ( .A1(_u10_u4_n3062 ), .A2(_u10_u4_n1923 ), .ZN(_u10_u4_n3154 ) );
NAND2_X1 _u10_u4_U997  ( .A1(_u10_u4_n2103 ), .A2(_u10_u4_n2509 ), .ZN(_u10_u4_n3161 ) );
NAND2_X1 _u10_u4_U996  ( .A1(_u10_u4_n2344 ), .A2(_u10_u4_n3161 ), .ZN(_u10_u4_n3160 ) );
NAND2_X1 _u10_u4_U995  ( .A1(_u10_u4_n3159 ), .A2(_u10_u4_n3160 ), .ZN(_u10_u4_n2635 ) );
AND3_X1 _u10_u4_U994  ( .A1(_u10_u4_n2549 ), .A2(_u10_u4_n2108 ), .A3(_u10_u4_n3126 ), .ZN(_u10_u4_n3093 ) );
NAND2_X1 _u10_u4_U993  ( .A1(_u10_u4_n3093 ), .A2(_u10_u4_n2941 ), .ZN(_u10_u4_n3158 ) );
NAND3_X1 _u10_u4_U992  ( .A1(_u10_u4_n3076 ), .A2(_u10_u4_n3066 ), .A3(_u10_u4_n3158 ), .ZN(_u10_u4_n3156 ) );
NAND2_X1 _u10_u4_U991  ( .A1(_u10_u4_n3156 ), .A2(_u10_u4_n3157 ), .ZN(_u10_u4_n3155 ) );
NAND3_X1 _u10_u4_U990  ( .A1(_u10_u4_n3154 ), .A2(_u10_u4_n2635 ), .A3(_u10_u4_n3155 ), .ZN(_u10_u4_n3131 ) );
INV_X1 _u10_u4_U989  ( .A(_u10_u4_n2594 ), .ZN(_u10_u4_n2846 ) );
NAND3_X1 _u10_u4_U988  ( .A1(_u10_u4_n2162 ), .A2(_u10_u4_n2082 ), .A3(_u10_u4_n2105 ), .ZN(_u10_u4_n2077 ) );
NAND4_X1 _u10_u4_U987  ( .A1(_u10_u4_n3153 ), .A2(_u10_u4_n1969 ), .A3(_u10_u4_n2846 ), .A4(_u10_u4_n2077 ), .ZN(_u10_u4_n3148 ) );
NAND2_X1 _u10_u4_U986  ( .A1(_u10_u4_n2838 ), .A2(_u10_u4_n3128 ), .ZN(_u10_u4_n3152 ) );
NAND2_X1 _u10_u4_U985  ( .A1(_u10_u4_n3152 ), .A2(_u10_u4_n2600 ), .ZN(_u10_u4_n3151 ) );
NAND2_X1 _u10_u4_U984  ( .A1(_u10_u4_n2282 ), .A2(_u10_u4_n3151 ), .ZN(_u10_u4_n2601 ) );
NOR4_X1 _u10_u4_U983  ( .A1(_u10_u4_n2885 ), .A2(_u10_u4_n2534 ), .A3(_u10_u4_n2214 ), .A4(_u10_u4_n3059 ), .ZN(_u10_u4_n3150 ) );
NOR2_X1 _u10_u4_U982  ( .A1(_u10_u4_n3150 ), .A2(_u10_u4_n2853 ), .ZN(_u10_u4_n3149 ) );
NOR4_X1 _u10_u4_U981  ( .A1(_u10_u4_n3148 ), .A2(_u10_u4_n2601 ), .A3(_u10_u4_n3149 ), .A4(_u10_u4_n1975 ), .ZN(_u10_u4_n3146 ) );
NAND3_X1 _u10_u4_U980  ( .A1(_u10_SYNOPSYS_UNCONNECTED_18 ), .A2(_u10_SYNOPSYS_UNCONNECTED_14 ), .A3(_u10_u4_n3147 ), .ZN(_u10_u4_n2071 ) );
NOR2_X1 _u10_u4_U979  ( .A1(_u10_u4_n3146 ), .A2(_u10_u4_n2071 ), .ZN(_u10_u4_n3132 ) );
NOR2_X1 _u10_u4_U978  ( .A1(1'b0), .A2(_u10_u4_n1847 ), .ZN(_u10_u4_n3143 ));
INV_X1 _u10_u4_U977  ( .A(_u10_u4_n3145 ), .ZN(_u10_u4_n3144 ) );
NOR2_X1 _u10_u4_U976  ( .A1(_u10_u4_n3143 ), .A2(_u10_u4_n3144 ), .ZN(_u10_u4_n3142 ) );
NOR2_X1 _u10_u4_U975  ( .A1(1'b0), .A2(_u10_u4_n3142 ), .ZN(_u10_u4_n3137 ));
NAND2_X1 _u10_u4_U974  ( .A1(_u10_u4_n2549 ), .A2(_u10_u4_n3141 ), .ZN(_u10_u4_n3138 ) );
NAND2_X1 _u10_u4_U973  ( .A1(_u10_u4_n1896 ), .A2(_u10_u4_n3140 ), .ZN(_u10_u4_n2544 ) );
NAND2_X1 _u10_u4_U972  ( .A1(_u10_u4_n2089 ), .A2(_u10_u4_n2544 ), .ZN(_u10_u4_n3139 ) );
NAND2_X1 _u10_u4_U971  ( .A1(_u10_u4_n3138 ), .A2(_u10_u4_n3139 ), .ZN(_u10_u4_n2795 ) );
NOR4_X1 _u10_u4_U970  ( .A1(_u10_u4_n2300 ), .A2(_u10_u4_n3137 ), .A3(_u10_u4_n2304 ), .A4(_u10_u4_n2795 ), .ZN(_u10_u4_n3134 ) );
NAND2_X1 _u10_u4_U969  ( .A1(_u10_u4_n3135 ), .A2(_u10_u4_n3136 ), .ZN(_u10_u4_n2085 ) );
NOR2_X1 _u10_u4_U968  ( .A1(_u10_u4_n3134 ), .A2(_u10_u4_n2085 ), .ZN(_u10_u4_n3133 ) );
NOR4_X1 _u10_u4_U967  ( .A1(_u10_u4_n3130 ), .A2(_u10_u4_n3131 ), .A3(_u10_u4_n3132 ), .A4(_u10_u4_n3133 ), .ZN(_u10_u4_n3016 ) );
INV_X1 _u10_u4_U966  ( .A(_u10_u4_n2686 ), .ZN(_u10_u4_n2278 ) );
NAND4_X1 _u10_u4_U965  ( .A1(_u10_u4_n2105 ), .A2(_u10_u4_n2278 ), .A3(_u10_u4_n3129 ), .A4(_u10_u4_n2600 ), .ZN(_u10_u4_n2437 ) );
NAND2_X1 _u10_u4_U964  ( .A1(_u10_u4_n3128 ), .A2(_u10_u4_n2437 ), .ZN(_u10_u4_n3127 ) );
NAND2_X1 _u10_u4_U963  ( .A1(_u10_u4_n2815 ), .A2(_u10_u4_n3127 ), .ZN(_u10_u4_n3098 ) );
INV_X1 _u10_u4_U962  ( .A(_u10_u4_n2573 ), .ZN(_u10_u4_n1967 ) );
NAND2_X1 _u10_u4_U961  ( .A1(_u10_u4_n3126 ), .A2(_u10_u4_n2078 ), .ZN(_u10_u4_n3123 ) );
NAND2_X1 _u10_u4_U960  ( .A1(_u10_u4_n3076 ), .A2(_u10_u4_n1925 ), .ZN(_u10_u4_n3125 ) );
NAND2_X1 _u10_u4_U959  ( .A1(_u10_u4_n2669 ), .A2(_u10_u4_n3125 ), .ZN(_u10_u4_n3124 ) );
NAND4_X1 _u10_u4_U958  ( .A1(_u10_u4_n3122 ), .A2(_u10_u4_n3123 ), .A3(_u10_u4_n3124 ), .A4(_u10_u4_n2579 ), .ZN(_u10_u4_n3121 ) );
NAND2_X1 _u10_u4_U957  ( .A1(_u10_u4_n3121 ), .A2(_u10_u4_n2874 ), .ZN(_u10_u4_n3120 ) );
NAND2_X1 _u10_u4_U956  ( .A1(_u10_u4_n2382 ), .A2(_u10_u4_n3120 ), .ZN(_u10_u4_n3119 ) );
NAND2_X1 _u10_u4_U955  ( .A1(_u10_u4_n1967 ), .A2(_u10_u4_n3119 ), .ZN(_u10_u4_n3099 ) );
NAND2_X1 _u10_u4_U954  ( .A1(_u10_u4_n3118 ), .A2(_u10_u4_n3001 ), .ZN(_u10_u4_n3117 ) );
NAND2_X1 _u10_u4_U953  ( .A1(_u10_u4_n2446 ), .A2(_u10_u4_n3117 ), .ZN(_u10_u4_n3116 ) );
NAND2_X1 _u10_u4_U952  ( .A1(_u10_u4_n2445 ), .A2(_u10_u4_n3116 ), .ZN(_u10_u4_n3100 ) );
OR2_X1 _u10_u4_U951  ( .A1(_u10_u4_n3115 ), .A2(_u10_u4_n2687 ), .ZN(_u10_u4_n3114 ) );
AND3_X1 _u10_u4_U950  ( .A1(_u10_u4_n2061 ), .A2(_u10_u4_n2166 ), .A3(_u10_u4_n3114 ), .ZN(_u10_u4_n3045 ) );
NOR2_X1 _u10_u4_U949  ( .A1(1'b0), .A2(_u10_u4_n3045 ), .ZN(_u10_u4_n3113 ));
NOR2_X1 _u10_u4_U948  ( .A1(_u10_u4_n3113 ), .A2(1'b0), .ZN(_u10_u4_n3112 ));
NOR2_X1 _u10_u4_U947  ( .A1(_u10_u4_n3112 ), .A2(_u10_u4_n2356 ), .ZN(_u10_u4_n3102 ) );
NAND2_X1 _u10_u4_U946  ( .A1(_u10_u4_n2571 ), .A2(_u10_u4_n2165 ), .ZN(_u10_u4_n3078 ) );
NAND2_X1 _u10_u4_U945  ( .A1(_u10_u4_n2365 ), .A2(_u10_u4_n3078 ), .ZN(_u10_u4_n2241 ) );
NOR2_X1 _u10_u4_U944  ( .A1(_u10_u4_n2377 ), .A2(_u10_u4_n2241 ), .ZN(_u10_u4_n3111 ) );
NOR2_X1 _u10_u4_U943  ( .A1(_u10_u4_n3111 ), .A2(_u10_u4_n1869 ), .ZN(_u10_u4_n3103 ) );
NOR2_X1 _u10_u4_U942  ( .A1(_u10_u4_n2999 ), .A2(_u10_u4_n2977 ), .ZN(_u10_u4_n3061 ) );
NOR2_X1 _u10_u4_U941  ( .A1(_u10_u4_n3061 ), .A2(_u10_u4_n2367 ), .ZN(_u10_u4_n3106 ) );
NAND2_X1 _u10_u4_U940  ( .A1(_u10_u4_n2977 ), .A2(_u10_u4_n3000 ), .ZN(_u10_u4_n3110 ) );
NAND2_X1 _u10_u4_U939  ( .A1(_u10_u4_n3109 ), .A2(_u10_u4_n3110 ), .ZN(_u10_u4_n1924 ) );
AND2_X1 _u10_u4_U938  ( .A1(_u10_u4_n1924 ), .A2(_u10_u4_n3108 ), .ZN(_u10_u4_n3107 ) );
NOR2_X1 _u10_u4_U937  ( .A1(_u10_u4_n3106 ), .A2(_u10_u4_n3107 ), .ZN(_u10_u4_n3105 ) );
NOR2_X1 _u10_u4_U936  ( .A1(_u10_u4_n3105 ), .A2(_u10_u4_n2008 ), .ZN(_u10_u4_n3104 ) );
NOR3_X1 _u10_u4_U935  ( .A1(_u10_u4_n3102 ), .A2(_u10_u4_n3103 ), .A3(_u10_u4_n3104 ), .ZN(_u10_u4_n3101 ) );
NAND4_X1 _u10_u4_U934  ( .A1(_u10_u4_n3098 ), .A2(_u10_u4_n3099 ), .A3(_u10_u4_n3100 ), .A4(_u10_u4_n3101 ), .ZN(_u10_u4_n3071 ) );
NOR2_X1 _u10_u4_U933  ( .A1(_u10_u4_n1926 ), .A2(_u10_u4_n2980 ), .ZN(_u10_u4_n2218 ) );
INV_X1 _u10_u4_U932  ( .A(_u10_u4_n2721 ), .ZN(_u10_u4_n2910 ) );
NAND2_X1 _u10_u4_U931  ( .A1(_u10_u4_n2910 ), .A2(_u10_u4_n1869 ), .ZN(_u10_u4_n2779 ) );
NAND2_X1 _u10_u4_U930  ( .A1(_u10_u4_n2218 ), .A2(_u10_u4_n2779 ), .ZN(_u10_u4_n3081 ) );
NAND2_X1 _u10_u4_U929  ( .A1(_u10_u4_n1922 ), .A2(_u10_u4_n1864 ), .ZN(_u10_u4_n2179 ) );
NOR3_X1 _u10_u4_U928  ( .A1(_u10_u4_n1961 ), .A2(_u10_u4_n1918 ), .A3(_u10_u4_n2179 ), .ZN(_u10_u4_n2693 ) );
NAND2_X1 _u10_u4_U927  ( .A1(_u10_u4_n3097 ), .A2(_u10_u4_n1924 ), .ZN(_u10_u4_n3096 ) );
NAND2_X1 _u10_u4_U926  ( .A1(_u10_u4_n1984 ), .A2(_u10_u4_n3096 ), .ZN(_u10_u4_n2506 ) );
INV_X1 _u10_u4_U925  ( .A(_u10_u4_n2506 ), .ZN(_u10_u4_n2366 ) );
NAND2_X1 _u10_u4_U924  ( .A1(_u10_u4_n2366 ), .A2(_u10_u4_n2375 ), .ZN(_u10_u4_n2236 ) );
NAND2_X1 _u10_u4_U923  ( .A1(_u10_u4_n2693 ), .A2(_u10_u4_n2236 ), .ZN(_u10_u4_n3082 ) );
NAND2_X1 _u10_u4_U922  ( .A1(1'b0), .A2(_u10_u4_n2126 ), .ZN(_u10_u4_n3095 ));
NAND2_X1 _u10_u4_U921  ( .A1(_u10_u4_n1956 ), .A2(_u10_u4_n3095 ), .ZN(_u10_u4_n2907 ) );
OR2_X1 _u10_u4_U920  ( .A1(_u10_u4_n2902 ), .A2(_u10_u4_n2907 ), .ZN(_u10_u4_n3085 ) );
NAND2_X1 _u10_u4_U919  ( .A1(_u10_u4_n2256 ), .A2(_u10_u4_n2113 ), .ZN(_u10_u4_n3094 ) );
NAND2_X1 _u10_u4_U918  ( .A1(_u10_u4_n2688 ), .A2(_u10_u4_n3094 ), .ZN(_u10_u4_n3092 ) );
NAND2_X1 _u10_u4_U917  ( .A1(_u10_u4_n3093 ), .A2(_u10_u4_n3092 ), .ZN(_u10_u4_n3086 ) );
INV_X1 _u10_u4_U916  ( .A(_u10_u4_n2159 ), .ZN(_u10_u4_n1894 ) );
NAND2_X1 _u10_u4_U915  ( .A1(_u10_u4_n3067 ), .A2(_u10_u4_n1894 ), .ZN(_u10_u4_n3091 ) );
INV_X1 _u10_u4_U914  ( .A(_u10_u4_n3092 ), .ZN(_u10_u4_n2234 ) );
NAND3_X1 _u10_u4_U913  ( .A1(_u10_u4_n3091 ), .A2(_u10_u4_n2126 ), .A3(_u10_u4_n2234 ), .ZN(_u10_u4_n3090 ) );
NAND2_X1 _u10_u4_U912  ( .A1(1'b0), .A2(_u10_u4_n3090 ), .ZN(_u10_u4_n3087 ));
NAND3_X1 _u10_u4_U911  ( .A1(_u10_u4_n2329 ), .A2(_u10_u4_n3089 ), .A3(_u10_u4_n2549 ), .ZN(_u10_u4_n3088 ) );
NAND4_X1 _u10_u4_U910  ( .A1(_u10_u4_n3085 ), .A2(_u10_u4_n3086 ), .A3(_u10_u4_n3087 ), .A4(_u10_u4_n3088 ), .ZN(_u10_u4_n3084 ) );
NAND2_X1 _u10_u4_U909  ( .A1(_u10_u4_n3084 ), .A2(_u10_u4_n2803 ), .ZN(_u10_u4_n3083 ) );
NAND3_X1 _u10_u4_U908  ( .A1(_u10_u4_n3081 ), .A2(_u10_u4_n3082 ), .A3(_u10_u4_n3083 ), .ZN(_u10_u4_n3072 ) );
INV_X1 _u10_u4_U907  ( .A(_u10_u4_n2689 ), .ZN(_u10_u4_n1955 ) );
NOR3_X1 _u10_u4_U906  ( .A1(_u10_u4_n1955 ), .A2(_u10_u4_n2813 ), .A3(_u10_u4_n2488 ), .ZN(_u10_u4_n3080 ) );
NOR2_X1 _u10_u4_U905  ( .A1(_u10_u4_n3080 ), .A2(_u10_u4_n2485 ), .ZN(_u10_u4_n3073 ) );
NAND3_X1 _u10_u4_U904  ( .A1(_u10_u4_n2621 ), .A2(_u10_u4_n2202 ), .A3(_u10_u4_n3079 ), .ZN(_u10_u4_n2110 ) );
NOR2_X1 _u10_u4_U903  ( .A1(_u10_u4_n2110 ), .A2(_u10_u4_n2218 ), .ZN(_u10_u4_n2775 ) );
INV_X1 _u10_u4_U902  ( .A(_u10_u4_n2775 ), .ZN(_u10_u4_n3024 ) );
INV_X1 _u10_u4_U901  ( .A(_u10_u4_n3078 ), .ZN(_u10_u4_n2133 ) );
INV_X1 _u10_u4_U900  ( .A(_u10_u4_n2007 ), .ZN(_u10_u4_n2358 ) );
NAND2_X1 _u10_u4_U899  ( .A1(_u10_u4_n2358 ), .A2(_u10_u4_n2886 ), .ZN(_u10_u4_n2240 ) );
INV_X1 _u10_u4_U898  ( .A(_u10_u4_n2240 ), .ZN(_u10_u4_n2083 ) );
NOR3_X1 _u10_u4_U897  ( .A1(_u10_u4_n2952 ), .A2(_u10_u4_n2004 ), .A3(_u10_u4_n1891 ), .ZN(_u10_u4_n3077 ) );
NAND3_X1 _u10_u4_U896  ( .A1(_u10_u4_n2083 ), .A2(_u10_u4_n2938 ), .A3(_u10_u4_n3077 ), .ZN(_u10_u4_n1886 ) );
NOR3_X1 _u10_u4_U895  ( .A1(_u10_u4_n3024 ), .A2(_u10_u4_n2133 ), .A3(_u10_u4_n1886 ), .ZN(_u10_u4_n3075 ) );
NOR2_X1 _u10_u4_U894  ( .A1(_u10_u4_n3075 ), .A2(_u10_u4_n3076 ), .ZN(_u10_u4_n3074 ) );
NOR4_X1 _u10_u4_U893  ( .A1(_u10_u4_n3071 ), .A2(_u10_u4_n3072 ), .A3(_u10_u4_n3073 ), .A4(_u10_u4_n3074 ), .ZN(_u10_u4_n3017 ) );
INV_X1 _u10_u4_U892  ( .A(_u10_u4_n3065 ), .ZN(_u10_u4_n3043 ) );
NAND2_X1 _u10_u4_U891  ( .A1(_u10_u4_n3043 ), .A2(_u10_u4_n2106 ), .ZN(_u10_u4_n3070 ) );
NAND2_X1 _u10_u4_U890  ( .A1(_u10_u4_n3070 ), .A2(_u10_u4_n2038 ), .ZN(_u10_u4_n3068 ) );
NAND2_X1 _u10_u4_U889  ( .A1(_u10_u4_n2344 ), .A2(_u10_u4_n2584 ), .ZN(_u10_u4_n3069 ) );
NAND3_X1 _u10_u4_U888  ( .A1(_u10_u4_n3068 ), .A2(_u10_u4_n1930 ), .A3(_u10_u4_n3069 ), .ZN(_u10_u4_n3047 ) );
NAND2_X1 _u10_u4_U887  ( .A1(_u10_u4_n2835 ), .A2(_u10_u4_n2466 ), .ZN(_u10_u4_n2130 ) );
INV_X1 _u10_u4_U886  ( .A(_u10_u4_n2130 ), .ZN(_u10_u4_n2168 ) );
NAND3_X1 _u10_u4_U885  ( .A1(_u10_u4_n3067 ), .A2(_u10_u4_n2329 ), .A3(_u10_u4_n2168 ), .ZN(_u10_u4_n2665 ) );
NAND3_X1 _u10_u4_U884  ( .A1(_u10_u4_n3065 ), .A2(_u10_u4_n3066 ), .A3(_u10_u4_n2342 ), .ZN(_u10_u4_n3064 ) );
NAND3_X1 _u10_u4_U883  ( .A1(_u10_u4_n3064 ), .A2(_u10_u4_n2175 ), .A3(_u10_u4_n2987 ), .ZN(_u10_u4_n3048 ) );
NOR3_X1 _u10_u4_U882  ( .A1(_u10_u4_n1849 ), .A2(1'b0), .A3(_u10_u4_n3063 ),.ZN(_u10_u4_n3050 ) );
NOR3_X1 _u10_u4_U881  ( .A1(_u10_u4_n2406 ), .A2(1'b0), .A3(_u10_u4_n3062 ),.ZN(_u10_u4_n3060 ) );
NOR3_X1 _u10_u4_U880  ( .A1(_u10_u4_n3060 ), .A2(1'b0), .A3(_u10_u4_n3061 ),.ZN(_u10_u4_n3051 ) );
NAND2_X1 _u10_u4_U879  ( .A1(_u10_u4_n3059 ), .A2(_u10_u4_n2049 ), .ZN(_u10_u4_n3056 ) );
NAND3_X1 _u10_u4_U878  ( .A1(_u10_u4_n3056 ), .A2(_u10_u4_n3057 ), .A3(_u10_u4_n3058 ), .ZN(_u10_u4_n3054 ) );
NOR4_X1 _u10_u4_U877  ( .A1(_u10_u4_n3054 ), .A2(_u10_u4_n3055 ), .A3(_u10_u4_n2055 ), .A4(_u10_u4_n2056 ), .ZN(_u10_u4_n3053 ) );
NOR3_X1 _u10_u4_U876  ( .A1(_u10_u4_n2346 ), .A2(1'b0), .A3(_u10_u4_n3053 ),.ZN(_u10_u4_n3052 ) );
NOR3_X1 _u10_u4_U875  ( .A1(_u10_u4_n3050 ), .A2(_u10_u4_n3051 ), .A3(_u10_u4_n3052 ), .ZN(_u10_u4_n3049 ) );
NAND4_X1 _u10_u4_U874  ( .A1(_u10_u4_n3047 ), .A2(_u10_u4_n2665 ), .A3(_u10_u4_n3048 ), .A4(_u10_u4_n3049 ), .ZN(_u10_u4_n3019 ) );
NAND2_X1 _u10_u4_U873  ( .A1(_u10_u4_n2056 ), .A2(_u10_u4_n2019 ), .ZN(_u10_u4_n3046 ) );
NAND2_X1 _u10_u4_U872  ( .A1(_u10_u4_n3045 ), .A2(_u10_u4_n3046 ), .ZN(_u10_u4_n3044 ) );
NAND2_X1 _u10_u4_U871  ( .A1(_u10_u4_n3044 ), .A2(_u10_u4_n2165 ), .ZN(_u10_u4_n3028 ) );
OR2_X1 _u10_u4_U870  ( .A1(_u10_u4_n2179 ), .A2(_u10_u4_n1961 ), .ZN(_u10_u4_n3037 ) );
NAND2_X1 _u10_u4_U869  ( .A1(_u10_u4_n3043 ), .A2(_u10_u4_n2336 ), .ZN(_u10_u4_n3042 ) );
NAND2_X1 _u10_u4_U868  ( .A1(_u10_u4_n3042 ), .A2(_u10_u4_n3006 ), .ZN(_u10_u4_n3041 ) );
NAND2_X1 _u10_u4_U867  ( .A1(_u10_u4_n3040 ), .A2(_u10_u4_n3041 ), .ZN(_u10_u4_n3026 ) );
NAND4_X1 _u10_u4_U866  ( .A1(_u10_u4_n3026 ), .A2(_u10_u4_n2520 ), .A3(_u10_u4_n1962 ), .A4(_u10_u4_n1864 ), .ZN(_u10_u4_n3039 ) );
NAND2_X1 _u10_u4_U865  ( .A1(_u10_u4_n3039 ), .A2(_u10_u4_n1922 ), .ZN(_u10_u4_n3038 ) );
NAND2_X1 _u10_u4_U864  ( .A1(_u10_u4_n3037 ), .A2(_u10_u4_n3038 ), .ZN(_u10_u4_n3035 ) );
NAND2_X1 _u10_u4_U863  ( .A1(_u10_u4_n2985 ), .A2(_u10_u4_n3036 ), .ZN(_u10_u4_n2432 ) );
NAND2_X1 _u10_u4_U862  ( .A1(_u10_u4_n3035 ), .A2(_u10_u4_n2432 ), .ZN(_u10_u4_n3029 ) );
INV_X1 _u10_u4_U861  ( .A(_u10_u4_n3034 ), .ZN(_u10_u4_n2777 ) );
INV_X1 _u10_u4_U860  ( .A(_u10_u4_n2772 ), .ZN(_u10_u4_n3032 ) );
NAND2_X1 _u10_u4_U859  ( .A1(_u10_u4_n1982 ), .A2(_u10_u4_n2978 ), .ZN(_u10_u4_n3033 ) );
NAND2_X1 _u10_u4_U858  ( .A1(_u10_u4_n3032 ), .A2(_u10_u4_n3033 ), .ZN(_u10_u4_n3031 ) );
NAND2_X1 _u10_u4_U857  ( .A1(_u10_u4_n2777 ), .A2(_u10_u4_n3031 ), .ZN(_u10_u4_n3030 ) );
NAND3_X1 _u10_u4_U856  ( .A1(_u10_u4_n3028 ), .A2(_u10_u4_n3029 ), .A3(_u10_u4_n3030 ), .ZN(_u10_u4_n3020 ) );
NOR3_X1 _u10_u4_U855  ( .A1(_u10_u4_n2179 ), .A2(1'b0), .A3(_u10_u4_n2375 ),.ZN(_u10_u4_n3027 ) );
NOR2_X1 _u10_u4_U854  ( .A1(_u10_u4_n3027 ), .A2(_u10_u4_n2177 ), .ZN(_u10_u4_n3025 ) );
NOR2_X1 _u10_u4_U853  ( .A1(_u10_u4_n3025 ), .A2(_u10_u4_n3026 ), .ZN(_u10_u4_n3021 ) );
NOR2_X1 _u10_u4_U852  ( .A1(_u10_u4_n2256 ), .A2(_u10_u4_n3024 ), .ZN(_u10_u4_n3023 ) );
NOR2_X1 _u10_u4_U851  ( .A1(_u10_u4_n3023 ), .A2(_u10_u4_n1868 ), .ZN(_u10_u4_n3022 ) );
NOR4_X1 _u10_u4_U850  ( .A1(_u10_u4_n3019 ), .A2(_u10_u4_n3020 ), .A3(_u10_u4_n3021 ), .A4(_u10_u4_n3022 ), .ZN(_u10_u4_n3018 ) );
NAND4_X1 _u10_u4_U849  ( .A1(_u10_u4_n3015 ), .A2(_u10_u4_n3016 ), .A3(_u10_u4_n3017 ), .A4(_u10_u4_n3018 ), .ZN(_u10_u4_n2958 ) );
NOR2_X1 _u10_u4_U848  ( .A1(1'b0), .A2(_u10_u4_n2573 ), .ZN(_u10_u4_n3011 ));
NOR2_X1 _u10_u4_U847  ( .A1(1'b0), .A2(_u10_u4_n2359 ), .ZN(_u10_u4_n3012 ));
NOR2_X1 _u10_u4_U846  ( .A1(1'b0), .A2(_u10_u4_n1859 ), .ZN(_u10_u4_n3013 ));
NOR2_X1 _u10_u4_U845  ( .A1(1'b0), .A2(_u10_u4_n1836 ), .ZN(_u10_u4_n3014 ));
NOR4_X1 _u10_u4_U844  ( .A1(_u10_u4_n3011 ), .A2(_u10_u4_n3012 ), .A3(_u10_u4_n3013 ), .A4(_u10_u4_n3014 ), .ZN(_u10_u4_n2959 ) );
NOR2_X1 _u10_u4_U843  ( .A1(1'b0), .A2(_u10_u4_n2025 ), .ZN(_u10_u4_n3007 ));
NOR2_X1 _u10_u4_U842  ( .A1(1'b0), .A2(_u10_u4_n2085 ), .ZN(_u10_u4_n3008 ));
NOR2_X1 _u10_u4_U841  ( .A1(1'b0), .A2(_u10_u4_n2607 ), .ZN(_u10_u4_n3009 ));
NOR2_X1 _u10_u4_U840  ( .A1(1'b0), .A2(_u10_u4_n2071 ), .ZN(_u10_u4_n3010 ));
NOR4_X1 _u10_u4_U839  ( .A1(_u10_u4_n3007 ), .A2(_u10_u4_n3008 ), .A3(_u10_u4_n3009 ), .A4(_u10_u4_n3010 ), .ZN(_u10_u4_n2960 ) );
NAND2_X1 _u10_u4_U838  ( .A1(_u10_u4_n1894 ), .A2(_u10_u4_n2466 ), .ZN(_u10_u4_n3002 ) );
NAND2_X1 _u10_u4_U837  ( .A1(_u10_u4_n2830 ), .A2(_u10_u4_n2600 ), .ZN(_u10_u4_n3003 ) );
NAND2_X1 _u10_u4_U836  ( .A1(_u10_u4_n1960 ), .A2(_u10_u4_n2431 ), .ZN(_u10_u4_n3004 ) );
NAND2_X1 _u10_u4_U835  ( .A1(_u10_u4_n2002 ), .A2(_u10_u4_n3006 ), .ZN(_u10_u4_n3005 ) );
NAND4_X1 _u10_u4_U834  ( .A1(_u10_u4_n3002 ), .A2(_u10_u4_n3003 ), .A3(_u10_u4_n3004 ), .A4(_u10_u4_n3005 ), .ZN(_u10_u4_n2992 ) );
NAND2_X1 _u10_u4_U833  ( .A1(_u10_u4_n2461 ), .A2(_u10_u4_n3001 ), .ZN(_u10_u4_n2997 ) );
NAND2_X1 _u10_u4_U832  ( .A1(_u10_u4_n2999 ), .A2(_u10_u4_n3000 ), .ZN(_u10_u4_n2998 ) );
NAND2_X1 _u10_u4_U831  ( .A1(_u10_u4_n2997 ), .A2(_u10_u4_n2998 ), .ZN(_u10_u4_n2993 ) );
NOR2_X1 _u10_u4_U830  ( .A1(_u10_SYNOPSYS_UNCONNECTED_14 ), .A2(_u10_u4_n2996 ), .ZN(_u10_u4_n2995 ) );
NOR2_X1 _u10_u4_U829  ( .A1(_u10_u4_n2995 ), .A2(_u10_u4_n2126 ), .ZN(_u10_u4_n2994 ) );
NOR4_X1 _u10_u4_U828  ( .A1(_u10_u4_n2992 ), .A2(_u10_u4_n2993 ), .A3(next_ch), .A4(_u10_u4_n2994 ), .ZN(_u10_u4_n2961 ) );
NAND2_X1 _u10_u4_U827  ( .A1(_u10_u4_n2445 ), .A2(_u10_u4_n2803 ), .ZN(_u10_u4_n2988 ) );
OR2_X1 _u10_u4_U826  ( .A1(_u10_u4_n2584 ), .A2(1'b0), .ZN(_u10_u4_n2989 ));
NAND2_X1 _u10_u4_U825  ( .A1(_u10_u4_n2709 ), .A2(_u10_u4_n2080 ), .ZN(_u10_u4_n2990 ) );
NAND2_X1 _u10_u4_U824  ( .A1(_u10_u4_n2183 ), .A2(_u10_u4_n2166 ), .ZN(_u10_u4_n2991 ) );
NAND4_X1 _u10_u4_U823  ( .A1(_u10_u4_n2988 ), .A2(_u10_u4_n2989 ), .A3(_u10_u4_n2990 ), .A4(_u10_u4_n2991 ), .ZN(_u10_u4_n2963 ) );
NAND2_X1 _u10_u4_U822  ( .A1(_u10_u4_n2987 ), .A2(_u10_u4_n1930 ), .ZN(_u10_u4_n2981 ) );
NAND2_X1 _u10_u4_U821  ( .A1(_u10_u4_n2986 ), .A2(_u10_u4_n2038 ), .ZN(_u10_u4_n2982 ) );
OR2_X1 _u10_u4_U820  ( .A1(_u10_u4_n2985 ), .A2(1'b0), .ZN(_u10_u4_n2983 ));
NAND2_X1 _u10_u4_U819  ( .A1(_u10_u4_n2169 ), .A2(_u10_u4_n2113 ), .ZN(_u10_u4_n2984 ) );
NAND4_X1 _u10_u4_U818  ( .A1(_u10_u4_n2981 ), .A2(_u10_u4_n2982 ), .A3(_u10_u4_n2983 ), .A4(_u10_u4_n2984 ), .ZN(_u10_u4_n2964 ) );
NAND2_X1 _u10_u4_U817  ( .A1(_u10_u4_n2509 ), .A2(_u10_u4_n1864 ), .ZN(_u10_u4_n2973 ) );
INV_X1 _u10_u4_U816  ( .A(_u10_u4_n2980 ), .ZN(_u10_u4_n1861 ) );
NAND2_X1 _u10_u4_U815  ( .A1(_u10_u4_n1861 ), .A2(_u10_u4_n1922 ), .ZN(_u10_u4_n2974 ) );
NAND2_X1 _u10_u4_U814  ( .A1(_u10_u4_n2979 ), .A2(_u10_u4_n2405 ), .ZN(_u10_u4_n2975 ) );
NAND2_X1 _u10_u4_U813  ( .A1(_u10_u4_n2977 ), .A2(_u10_u4_n2978 ), .ZN(_u10_u4_n2976 ) );
NAND4_X1 _u10_u4_U812  ( .A1(_u10_u4_n2973 ), .A2(_u10_u4_n2974 ), .A3(_u10_u4_n2975 ), .A4(_u10_u4_n2976 ), .ZN(_u10_u4_n2965 ) );
NAND2_X1 _u10_u4_U811  ( .A1(_u10_u4_n2507 ), .A2(_u10_u4_n2972 ), .ZN(_u10_u4_n2967 ) );
NAND2_X1 _u10_u4_U810  ( .A1(_u10_u4_n2043 ), .A2(_u10_u4_n1965 ), .ZN(_u10_u4_n2968 ) );
NAND2_X1 _u10_u4_U809  ( .A1(_u10_u4_n2063 ), .A2(_u10_u4_n1853 ), .ZN(_u10_u4_n2969 ) );
NAND2_X1 _u10_u4_U808  ( .A1(_u10_u4_n2971 ), .A2(_u10_u4_n2175 ), .ZN(_u10_u4_n2970 ) );
NAND4_X1 _u10_u4_U807  ( .A1(_u10_u4_n2967 ), .A2(_u10_u4_n2968 ), .A3(_u10_u4_n2969 ), .A4(_u10_u4_n2970 ), .ZN(_u10_u4_n2966 ) );
NOR4_X1 _u10_u4_U806  ( .A1(_u10_u4_n2963 ), .A2(_u10_u4_n2964 ), .A3(_u10_u4_n2965 ), .A4(_u10_u4_n2966 ), .ZN(_u10_u4_n2962 ) );
AND4_X1 _u10_u4_U805  ( .A1(_u10_u4_n2959 ), .A2(_u10_u4_n2960 ), .A3(_u10_u4_n2961 ), .A4(_u10_u4_n2962 ), .ZN(_u10_u4_n1819 ) );
MUX2_X1 _u10_u4_U804  ( .A(_u10_u4_n2958 ), .B(_u10_SYNOPSYS_UNCONNECTED_18 ), .S(_u10_u4_n1819 ), .Z(_u10_u4_n1808 ) );
NOR2_X1 _u10_u4_U803  ( .A1(_u10_u4_n2531 ), .A2(_u10_u4_n2607 ), .ZN(_u10_u4_n1911 ) );
NAND2_X1 _u10_u4_U802  ( .A1(_u10_u4_n1911 ), .A2(_u10_u4_n2957 ), .ZN(_u10_u4_n2954 ) );
NAND2_X1 _u10_u4_U801  ( .A1(_u10_u4_n1853 ), .A2(_u10_u4_n1965 ), .ZN(_u10_u4_n2956 ) );
NAND2_X1 _u10_u4_U800  ( .A1(_u10_u4_n1966 ), .A2(_u10_u4_n2956 ), .ZN(_u10_u4_n2955 ) );
NAND2_X1 _u10_u4_U799  ( .A1(_u10_u4_n2954 ), .A2(_u10_u4_n2955 ), .ZN(_u10_u4_n2670 ) );
NOR3_X1 _u10_u4_U798  ( .A1(_u10_u4_n1852 ), .A2(1'b0), .A3(_u10_u4_n1853 ),.ZN(_u10_u4_n2708 ) );
NAND2_X1 _u10_u4_U797  ( .A1(_u10_u4_n2708 ), .A2(_u10_u4_n2080 ), .ZN(_u10_u4_n2355 ) );
NOR2_X1 _u10_u4_U796  ( .A1(_u10_u4_n2355 ), .A2(1'b0), .ZN(_u10_u4_n2599 ));
NAND2_X1 _u10_u4_U795  ( .A1(_u10_u4_n2953 ), .A2(_u10_u4_n2599 ), .ZN(_u10_u4_n2423 ) );
OR2_X1 _u10_u4_U794  ( .A1(_u10_u4_n2423 ), .A2(_u10_u4_n2359 ), .ZN(_u10_u4_n2949 ) );
NAND3_X1 _u10_u4_U793  ( .A1(_u10_u4_n2105 ), .A2(_u10_u4_n1936 ), .A3(_u10_u4_n2952 ), .ZN(_u10_u4_n2950 ) );
NAND3_X1 _u10_u4_U792  ( .A1(_u10_u4_n2549 ), .A2(_u10_u4_n1936 ), .A3(1'b0),.ZN(_u10_u4_n2096 ) );
INV_X1 _u10_u4_U791  ( .A(_u10_u4_n2096 ), .ZN(_u10_u4_n2301 ) );
NAND2_X1 _u10_u4_U790  ( .A1(_u10_u4_n2301 ), .A2(_u10_u4_n2446 ), .ZN(_u10_u4_n2368 ) );
INV_X1 _u10_u4_U789  ( .A(_u10_u4_n2368 ), .ZN(_u10_u4_n2326 ) );
NAND2_X1 _u10_u4_U788  ( .A1(_u10_u4_n2326 ), .A2(_u10_u4_n2941 ), .ZN(_u10_u4_n2800 ) );
INV_X1 _u10_u4_U787  ( .A(_u10_u4_n2800 ), .ZN(_u10_u4_n2081 ) );
NAND2_X1 _u10_u4_U786  ( .A1(_u10_u4_n2081 ), .A2(_u10_u4_n2049 ), .ZN(_u10_u4_n2855 ) );
INV_X1 _u10_u4_U785  ( .A(_u10_u4_n2855 ), .ZN(_u10_u4_n2347 ) );
NAND2_X1 _u10_u4_U784  ( .A1(_u10_u4_n2347 ), .A2(_u10_u4_n2063 ), .ZN(_u10_u4_n2951 ) );
NAND3_X1 _u10_u4_U783  ( .A1(_u10_u4_n2949 ), .A2(_u10_u4_n2950 ), .A3(_u10_u4_n2951 ), .ZN(_u10_u4_n1997 ) );
INV_X1 _u10_u4_U782  ( .A(_u10_u4_n1997 ), .ZN(_u10_u4_n2917 ) );
AND2_X1 _u10_u4_U781  ( .A1(_u10_u4_n2709 ), .A2(_u10_u4_n2708 ), .ZN(_u10_u4_n2942 ) );
INV_X1 _u10_u4_U780  ( .A(_u10_u4_n2907 ), .ZN(_u10_u4_n2737 ) );
NAND2_X1 _u10_u4_U779  ( .A1(_u10_u4_n2737 ), .A2(_u10_u4_n2803 ), .ZN(_u10_u4_n1888 ) );
NOR2_X1 _u10_u4_U778  ( .A1(_u10_u4_n2001 ), .A2(_u10_u4_n1888 ), .ZN(_u10_u4_n2943 ) );
NAND4_X1 _u10_u4_U777  ( .A1(1'b0), .A2(_u10_u4_n2078 ), .A3(_u10_u4_n2059 ),.A4(_u10_u4_n2031 ), .ZN(_u10_u4_n2578 ) );
NOR3_X1 _u10_u4_U776  ( .A1(_u10_u4_n2719 ), .A2(_u10_u4_n2130 ), .A3(_u10_u4_n2305 ), .ZN(_u10_u4_n2386 ) );
NAND2_X1 _u10_u4_U775  ( .A1(_u10_u4_n2386 ), .A2(_u10_u4_n2669 ), .ZN(_u10_u4_n2948 ) );
NAND3_X1 _u10_u4_U774  ( .A1(_u10_u4_n2578 ), .A2(_u10_u4_n2947 ), .A3(_u10_u4_n2948 ), .ZN(_u10_u4_n2750 ) );
NOR2_X1 _u10_u4_U773  ( .A1(_u10_u4_n2274 ), .A2(_u10_u4_n2852 ), .ZN(_u10_u4_n2946 ) );
NOR3_X1 _u10_u4_U772  ( .A1(_u10_u4_n2750 ), .A2(1'b0), .A3(_u10_u4_n2946 ),.ZN(_u10_u4_n2945 ) );
NOR2_X1 _u10_u4_U771  ( .A1(_u10_u4_n2945 ), .A2(_u10_u4_n2359 ), .ZN(_u10_u4_n2944 ) );
NOR3_X1 _u10_u4_U770  ( .A1(_u10_u4_n2942 ), .A2(_u10_u4_n2943 ), .A3(_u10_u4_n2944 ), .ZN(_u10_u4_n2919 ) );
NOR2_X1 _u10_u4_U769  ( .A1(_u10_u4_n2423 ), .A2(1'b0), .ZN(_u10_u4_n1979 ));
NAND3_X1 _u10_u4_U768  ( .A1(_u10_u4_n2549 ), .A2(_u10_u4_n1936 ), .A3(_u10_u4_n1979 ), .ZN(_u10_u4_n2328 ) );
INV_X1 _u10_u4_U767  ( .A(_u10_u4_n2328 ), .ZN(_u10_u4_n2554 ) );
NAND3_X1 _u10_u4_U766  ( .A1(_u10_u4_n2941 ), .A2(_u10_u4_n2446 ), .A3(_u10_u4_n2554 ), .ZN(_u10_u4_n2115 ) );
NOR2_X1 _u10_u4_U765  ( .A1(_u10_u4_n2578 ), .A2(_u10_u4_n2030 ), .ZN(_u10_u4_n2553 ) );
INV_X1 _u10_u4_U764  ( .A(_u10_u4_n2553 ), .ZN(_u10_u4_n2269 ) );
NOR2_X1 _u10_u4_U763  ( .A1(_u10_u4_n2269 ), .A2(_u10_u4_n2790 ), .ZN(_u10_u4_n2657 ) );
INV_X1 _u10_u4_U762  ( .A(_u10_u4_n2657 ), .ZN(_u10_u4_n2210 ) );
NOR2_X1 _u10_u4_U761  ( .A1(_u10_u4_n2210 ), .A2(_u10_u4_n2911 ), .ZN(_u10_u4_n2213 ) );
INV_X1 _u10_u4_U760  ( .A(_u10_u4_n2213 ), .ZN(_u10_u4_n2456 ) );
NAND2_X1 _u10_u4_U759  ( .A1(_u10_u4_n2115 ), .A2(_u10_u4_n2456 ), .ZN(_u10_u4_n2634 ) );
INV_X1 _u10_u4_U758  ( .A(_u10_u4_n2634 ), .ZN(_u10_u4_n2220 ) );
NOR2_X1 _u10_u4_U757  ( .A1(_u10_u4_n2081 ), .A2(_u10_u4_n2386 ), .ZN(_u10_u4_n2131 ) );
NAND2_X1 _u10_u4_U756  ( .A1(_u10_u4_n2940 ), .A2(_u10_u4_n2131 ), .ZN(_u10_u4_n2138 ) );
INV_X1 _u10_u4_U755  ( .A(_u10_u4_n2138 ), .ZN(_u10_u4_n2927 ) );
NAND2_X1 _u10_u4_U754  ( .A1(_u10_u4_n2220 ), .A2(_u10_u4_n2927 ), .ZN(_u10_u4_n2939 ) );
NAND2_X1 _u10_u4_U753  ( .A1(_u10_u4_n1885 ), .A2(_u10_u4_n2939 ), .ZN(_u10_u4_n2931 ) );
NAND3_X1 _u10_u4_U752  ( .A1(_u10_u4_n1859 ), .A2(_u10_u4_n2365 ), .A3(_u10_u4_n2938 ), .ZN(_u10_u4_n2935 ) );
NAND3_X1 _u10_u4_U751  ( .A1(_u10_u4_n2927 ), .A2(_u10_u4_n2937 ), .A3(_u10_u4_n2220 ), .ZN(_u10_u4_n2936 ) );
NAND2_X1 _u10_u4_U750  ( .A1(_u10_u4_n2935 ), .A2(_u10_u4_n2936 ), .ZN(_u10_u4_n2932 ) );
INV_X1 _u10_u4_U749  ( .A(_u10_u4_n1937 ), .ZN(_u10_u4_n2350 ) );
NAND2_X1 _u10_u4_U748  ( .A1(_u10_u4_n1913 ), .A2(_u10_u4_n2350 ), .ZN(_u10_u4_n2934 ) );
NAND2_X1 _u10_u4_U747  ( .A1(_u10_u4_n2386 ), .A2(_u10_u4_n2934 ), .ZN(_u10_u4_n2933 ) );
NAND3_X1 _u10_u4_U746  ( .A1(_u10_u4_n2931 ), .A2(_u10_u4_n2932 ), .A3(_u10_u4_n2933 ), .ZN(_u10_u4_n2921 ) );
OR2_X1 _u10_u4_U745  ( .A1(_u10_u4_n2213 ), .A2(_u10_u4_n2386 ), .ZN(_u10_u4_n2930 ) );
NAND2_X1 _u10_u4_U744  ( .A1(_u10_u4_n2049 ), .A2(_u10_u4_n2930 ), .ZN(_u10_u4_n2228 ) );
AND2_X1 _u10_u4_U743  ( .A1(_u10_u4_n2228 ), .A2(_u10_u4_n2699 ), .ZN(_u10_u4_n2929 ) );
NOR2_X1 _u10_u4_U742  ( .A1(_u10_u4_n2929 ), .A2(_u10_u4_n2495 ), .ZN(_u10_u4_n2922 ) );
NOR2_X1 _u10_u4_U741  ( .A1(_u10_u4_n2633 ), .A2(_u10_u4_n2877 ), .ZN(_u10_u4_n2928 ) );
NOR2_X1 _u10_u4_U740  ( .A1(_u10_u4_n2928 ), .A2(_u10_u4_n2886 ), .ZN(_u10_u4_n2923 ) );
NOR2_X1 _u10_u4_U739  ( .A1(_u10_u4_n2927 ), .A2(_u10_u4_n2531 ), .ZN(_u10_u4_n2926 ) );
NOR2_X1 _u10_u4_U738  ( .A1(_u10_u4_n2926 ), .A2(_u10_u4_n2687 ), .ZN(_u10_u4_n2925 ) );
NOR2_X1 _u10_u4_U737  ( .A1(_u10_u4_n2925 ), .A2(_u10_u4_n1849 ), .ZN(_u10_u4_n2924 ) );
NOR4_X1 _u10_u4_U736  ( .A1(_u10_u4_n2921 ), .A2(_u10_u4_n2922 ), .A3(_u10_u4_n2923 ), .A4(_u10_u4_n2924 ), .ZN(_u10_u4_n2920 ) );
NAND4_X1 _u10_u4_U735  ( .A1(_u10_u4_n2917 ), .A2(_u10_u4_n2918 ), .A3(_u10_u4_n2919 ), .A4(_u10_u4_n2920 ), .ZN(_u10_u4_n2312 ) );
NOR2_X1 _u10_u4_U734  ( .A1(_u10_u4_n2600 ), .A2(_u10_u4_n2686 ), .ZN(_u10_u4_n2401 ) );
NAND2_X1 _u10_u4_U733  ( .A1(_u10_u4_n2401 ), .A2(_u10_u4_n2549 ), .ZN(_u10_u4_n2547 ) );
INV_X1 _u10_u4_U732  ( .A(_u10_u4_n2547 ), .ZN(_u10_u4_n2794 ) );
NAND3_X1 _u10_u4_U731  ( .A1(_u10_u4_n2364 ), .A2(_u10_u4_n2667 ), .A3(_u10_u4_n2794 ), .ZN(_u10_u4_n2535 ) );
INV_X1 _u10_u4_U730  ( .A(_u10_u4_n2535 ), .ZN(_u10_u4_n2586 ) );
NAND2_X1 _u10_u4_U729  ( .A1(_u10_u4_n2586 ), .A2(_u10_u4_n2571 ), .ZN(_u10_u4_n2916 ) );
NAND2_X1 _u10_u4_U728  ( .A1(_u10_u4_n2837 ), .A2(_u10_u4_n2916 ), .ZN(_u10_u4_n2436 ) );
NAND2_X1 _u10_u4_U727  ( .A1(_u10_u4_n2915 ), .A2(_u10_u4_n2571 ), .ZN(_u10_u4_n2914 ) );
NAND2_X1 _u10_u4_U726  ( .A1(_u10_u4_n2166 ), .A2(_u10_u4_n2914 ), .ZN(_u10_u4_n2017 ) );
NOR2_X1 _u10_u4_U725  ( .A1(_u10_u4_n2485 ), .A2(_u10_u4_n1841 ), .ZN(_u10_u4_n2913 ) );
OR4_X1 _u10_u4_U724  ( .A1(_u10_u4_n2436 ), .A2(_u10_u4_n2017 ), .A3(_u10_u4_n2913 ), .A4(_u10_u4_n2442 ), .ZN(_u10_u4_n2912 ) );
NAND2_X1 _u10_u4_U723  ( .A1(_u10_u4_n2709 ), .A2(_u10_u4_n2912 ), .ZN(_u10_u4_n2888 ) );
NAND3_X1 _u10_u4_U722  ( .A1(_u10_u4_n2078 ), .A2(_u10_u4_n2031 ), .A3(1'b0),.ZN(_u10_u4_n2580 ) );
INV_X1 _u10_u4_U721  ( .A(_u10_u4_n2580 ), .ZN(_u10_u4_n2680 ) );
AND2_X1 _u10_u4_U720  ( .A1(_u10_u4_n2680 ), .A2(_u10_u4_n2668 ), .ZN(_u10_u4_n1950 ) );
NAND2_X1 _u10_u4_U719  ( .A1(_u10_u4_n1950 ), .A2(_u10_u4_n2089 ), .ZN(_u10_u4_n2095 ) );
INV_X1 _u10_u4_U718  ( .A(_u10_u4_n2095 ), .ZN(_u10_u4_n2542 ) );
NAND2_X1 _u10_u4_U717  ( .A1(_u10_u4_n2542 ), .A2(_u10_u4_n2446 ), .ZN(_u10_u4_n1887 ) );
NOR2_X1 _u10_u4_U716  ( .A1(_u10_u4_n1887 ), .A2(_u10_u4_n2911 ), .ZN(_u10_u4_n2114 ) );
INV_X1 _u10_u4_U715  ( .A(_u10_u4_n2114 ), .ZN(_u10_u4_n1940 ) );
NAND3_X1 _u10_u4_U714  ( .A1(_u10_u4_n2535 ), .A2(_u10_u4_n1940 ), .A3(_u10_u4_n2910 ), .ZN(_u10_u4_n2524 ) );
NAND2_X1 _u10_u4_U713  ( .A1(_u10_u4_n2524 ), .A2(_u10_u4_n2488 ), .ZN(_u10_u4_n2889 ) );
NAND2_X1 _u10_u4_U712  ( .A1(_u10_u4_n2220 ), .A2(_u10_u4_n1940 ), .ZN(_u10_u4_n2763 ) );
NOR2_X1 _u10_u4_U711  ( .A1(_u10_u4_n2763 ), .A2(_u10_u4_n2586 ), .ZN(_u10_u4_n2808 ) );
NOR2_X1 _u10_u4_U710  ( .A1(_u10_u4_n2808 ), .A2(_u10_u4_n2350 ), .ZN(_u10_u4_n2908 ) );
NOR2_X1 _u10_u4_U709  ( .A1(_u10_u4_n2544 ), .A2(_u10_u4_n1950 ), .ZN(_u10_u4_n2899 ) );
NOR2_X1 _u10_u4_U708  ( .A1(_u10_u4_n2899 ), .A2(_u10_u4_n2159 ), .ZN(_u10_u4_n2909 ) );
NOR2_X1 _u10_u4_U707  ( .A1(_u10_u4_n2908 ), .A2(_u10_u4_n2909 ), .ZN(_u10_u4_n2890 ) );
NOR3_X1 _u10_u4_U706  ( .A1(_u10_u4_n2547 ), .A2(_u10_u4_n1846 ), .A3(_u10_u4_n2907 ), .ZN(_u10_u4_n2892 ) );
NOR3_X1 _u10_u4_U705  ( .A1(_u10_u4_n2240 ), .A2(_u10_u4_n2377 ), .A3(_u10_u4_n1911 ), .ZN(_u10_u4_n2906 ) );
NOR2_X1 _u10_u4_U704  ( .A1(_u10_u4_n2906 ), .A2(_u10_u4_n2535 ), .ZN(_u10_u4_n2893 ) );
NAND2_X1 _u10_u4_U703  ( .A1(_u10_u4_n2554 ), .A2(_u10_u4_n2446 ), .ZN(_u10_u4_n2903 ) );
AND3_X1 _u10_u4_U702  ( .A1(_u10_u4_n2210 ), .A2(_u10_u4_n2905 ), .A3(_u10_u4_n1887 ), .ZN(_u10_u4_n2904 ) );
NAND4_X1 _u10_u4_U701  ( .A1(_u10_u4_n2902 ), .A2(_u10_u4_n2498 ), .A3(_u10_u4_n2903 ), .A4(_u10_u4_n2904 ), .ZN(_u10_u4_n2788 ) );
INV_X1 _u10_u4_U700  ( .A(_u10_u4_n2788 ), .ZN(_u10_u4_n2901 ) );
NOR2_X1 _u10_u4_U699  ( .A1(_u10_u4_n2901 ), .A2(_u10_u4_n1888 ), .ZN(_u10_u4_n2894 ) );
NOR2_X1 _u10_u4_U698  ( .A1(_u10_u4_n2401 ), .A2(_u10_u4_n2553 ), .ZN(_u10_u4_n2900 ) );
NOR2_X1 _u10_u4_U697  ( .A1(_u10_u4_n2900 ), .A2(_u10_u4_n1954 ), .ZN(_u10_u4_n2897 ) );
NOR2_X1 _u10_u4_U696  ( .A1(1'b0), .A2(_u10_u4_n2899 ), .ZN(_u10_u4_n2898 ));
NOR2_X1 _u10_u4_U695  ( .A1(_u10_u4_n2897 ), .A2(_u10_u4_n2898 ), .ZN(_u10_u4_n2896 ) );
NOR2_X1 _u10_u4_U694  ( .A1(_u10_u4_n2896 ), .A2(_u10_u4_n1843 ), .ZN(_u10_u4_n2895 ) );
NOR4_X1 _u10_u4_U693  ( .A1(_u10_u4_n2892 ), .A2(_u10_u4_n2893 ), .A3(_u10_u4_n2894 ), .A4(_u10_u4_n2895 ), .ZN(_u10_u4_n2891 ) );
NAND4_X1 _u10_u4_U692  ( .A1(_u10_u4_n2888 ), .A2(_u10_u4_n2889 ), .A3(_u10_u4_n2890 ), .A4(_u10_u4_n2891 ), .ZN(_u10_u4_n2610 ) );
NOR4_X1 _u10_u4_U691  ( .A1(_u10_u4_n2670 ), .A2(_u10_u4_n2312 ), .A3(_u10_u4_n2610 ), .A4(_u10_u4_n2887 ), .ZN(_u10_u4_n2724 ) );
NOR2_X1 _u10_u4_U690  ( .A1(_u10_u4_n2883 ), .A2(_u10_u4_n2535 ), .ZN(_u10_u4_n2861 ) );
NOR2_X1 _u10_u4_U689  ( .A1(_u10_u4_n1855 ), .A2(_u10_u4_n1869 ), .ZN(_u10_u4_n2862 ) );
NOR2_X1 _u10_u4_U688  ( .A1(_u10_u4_n2886 ), .A2(_u10_u4_n2695 ), .ZN(_u10_u4_n2863 ) );
NAND2_X1 _u10_u4_U687  ( .A1(_u10_u4_n2813 ), .A2(_u10_u4_n2885 ), .ZN(_u10_u4_n2864 ) );
NAND2_X1 _u10_u4_U686  ( .A1(_u10_u4_n2114 ), .A2(_u10_u4_n2884 ), .ZN(_u10_u4_n2865 ) );
NAND2_X1 _u10_u4_U685  ( .A1(1'b0), .A2(_u10_u4_n2667 ), .ZN(_u10_u4_n2112 ));
NOR3_X1 _u10_u4_U684  ( .A1(_u10_u4_n2883 ), .A2(_u10_u4_n2112 ), .A3(_u10_u4_n2719 ), .ZN(_u10_u4_n2878 ) );
INV_X1 _u10_u4_U683  ( .A(_u10_u4_n2112 ), .ZN(_u10_u4_n1856 ) );
NAND2_X1 _u10_u4_U682  ( .A1(_u10_u4_n2364 ), .A2(_u10_u4_n1856 ), .ZN(_u10_u4_n2882 ) );
NAND2_X1 _u10_u4_U681  ( .A1(_u10_u4_n2882 ), .A2(_u10_u4_n1869 ), .ZN(_u10_u4_n2050 ) );
INV_X1 _u10_u4_U680  ( .A(_u10_u4_n2050 ), .ZN(_u10_u4_n1939 ) );
NOR2_X1 _u10_u4_U679  ( .A1(_u10_u4_n1939 ), .A2(_u10_u4_n1841 ), .ZN(_u10_u4_n2881 ) );
NOR2_X1 _u10_u4_U678  ( .A1(_u10_u4_n2881 ), .A2(_u10_u4_n2840 ), .ZN(_u10_u4_n2880 ) );
NOR2_X1 _u10_u4_U677  ( .A1(_u10_u4_n2880 ), .A2(_u10_u4_n1836 ), .ZN(_u10_u4_n2879 ) );
NOR2_X1 _u10_u4_U676  ( .A1(_u10_u4_n2878 ), .A2(_u10_u4_n2879 ), .ZN(_u10_u4_n2866 ) );
NOR2_X1 _u10_u4_U675  ( .A1(_u10_u4_n2081 ), .A2(_u10_u4_n2877 ), .ZN(_u10_u4_n1840 ) );
NAND2_X1 _u10_u4_U674  ( .A1(_u10_u4_n1840 ), .A2(_u10_u4_n2115 ), .ZN(_u10_u4_n1873 ) );
NAND2_X1 _u10_u4_U673  ( .A1(_u10_u4_n2695 ), .A2(_u10_u4_n1940 ), .ZN(_u10_u4_n1874 ) );
NOR3_X1 _u10_u4_U672  ( .A1(_u10_u4_n2050 ), .A2(_u10_u4_n1873 ), .A3(_u10_u4_n1874 ), .ZN(_u10_u4_n2876 ) );
NOR2_X1 _u10_u4_U671  ( .A1(_u10_u4_n2876 ), .A2(_u10_u4_n1913 ), .ZN(_u10_u4_n2868 ) );
NAND2_X1 _u10_u4_U670  ( .A1(_u10_u4_n2875 ), .A2(_u10_u4_n2466 ), .ZN(_u10_u4_n2872 ) );
INV_X1 _u10_u4_U669  ( .A(_u10_u4_n1979 ), .ZN(_u10_u4_n2746 ) );
NAND2_X1 _u10_u4_U668  ( .A1(_u10_u4_n2874 ), .A2(_u10_u4_n2746 ), .ZN(_u10_u4_n1935 ) );
NAND3_X1 _u10_u4_U667  ( .A1(_u10_u4_n1935 ), .A2(_u10_u4_n1936 ), .A3(_u10_u4_n2467 ), .ZN(_u10_u4_n2873 ) );
NAND2_X1 _u10_u4_U666  ( .A1(_u10_u4_n2872 ), .A2(_u10_u4_n2873 ), .ZN(_u10_u4_n2264 ) );
AND2_X1 _u10_u4_U665  ( .A1(_u10_u4_n2264 ), .A2(_u10_u4_n2461 ), .ZN(_u10_u4_n2869 ) );
AND2_X1 _u10_u4_U664  ( .A1(_u10_u4_n1966 ), .A2(_u10_u4_n2761 ), .ZN(_u10_u4_n2870 ) );
NOR2_X1 _u10_u4_U663  ( .A1(_u10_u4_n2159 ), .A2(_u10_u4_n2163 ), .ZN(_u10_u4_n2871 ) );
NOR4_X1 _u10_u4_U662  ( .A1(_u10_u4_n2868 ), .A2(_u10_u4_n2869 ), .A3(_u10_u4_n2870 ), .A4(_u10_u4_n2871 ), .ZN(_u10_u4_n2867 ) );
NAND4_X1 _u10_u4_U661  ( .A1(_u10_u4_n2864 ), .A2(_u10_u4_n2865 ), .A3(_u10_u4_n2866 ), .A4(_u10_u4_n2867 ), .ZN(_u10_u4_n1992 ) );
NOR4_X1 _u10_u4_U660  ( .A1(_u10_u4_n2861 ), .A2(_u10_u4_n2862 ), .A3(_u10_u4_n2863 ), .A4(_u10_u4_n1992 ), .ZN(_u10_u4_n2725 ) );
NAND2_X1 _u10_u4_U659  ( .A1(_u10_u4_n2364 ), .A2(_u10_u4_n1846 ), .ZN(_u10_u4_n2744 ) );
NAND4_X1 _u10_u4_U658  ( .A1(_u10_u4_n2765 ), .A2(_u10_u4_n1939 ), .A3(_u10_u4_n2744 ), .A4(_u10_u4_n2535 ), .ZN(_u10_u4_n2860 ) );
NAND2_X1 _u10_u4_U657  ( .A1(_u10_u4_n2049 ), .A2(_u10_u4_n2860 ), .ZN(_u10_u4_n2856 ) );
NOR4_X1 _u10_u4_U656  ( .A1(1'b0), .A2(_u10_u4_n2858 ), .A3(_u10_u4_n2859 ),.A4(_u10_u4_n2051 ), .ZN(_u10_u4_n2857 ) );
NAND4_X1 _u10_u4_U655  ( .A1(_u10_u4_n2228 ), .A2(_u10_u4_n2855 ), .A3(_u10_u4_n2856 ), .A4(_u10_u4_n2857 ), .ZN(_u10_u4_n2854 ) );
NAND2_X1 _u10_u4_U654  ( .A1(_u10_u4_n2043 ), .A2(_u10_u4_n2854 ), .ZN(_u10_u4_n2821 ) );
INV_X1 _u10_u4_U653  ( .A(_u10_u4_n2071 ), .ZN(_u10_u4_n2279 ) );
INV_X1 _u10_u4_U652  ( .A(_u10_u4_n2599 ), .ZN(_u10_u4_n2357 ) );
OR2_X1 _u10_u4_U651  ( .A1(_u10_u4_n2744 ), .A2(_u10_u4_n2853 ), .ZN(_u10_u4_n2844 ) );
NAND2_X1 _u10_u4_U650  ( .A1(_u10_u4_n2131 ), .A2(_u10_u4_n2852 ), .ZN(_u10_u4_n2851 ) );
NAND2_X1 _u10_u4_U649  ( .A1(_u10_u4_n2082 ), .A2(_u10_u4_n2851 ), .ZN(_u10_u4_n2848 ) );
NAND2_X1 _u10_u4_U648  ( .A1(_u10_u4_n2850 ), .A2(_u10_u4_n2600 ), .ZN(_u10_u4_n2849 ) );
NAND3_X1 _u10_u4_U647  ( .A1(_u10_u4_n2848 ), .A2(_u10_u4_n2077 ), .A3(_u10_u4_n2849 ), .ZN(_u10_u4_n2287 ) );
NAND2_X1 _u10_u4_U646  ( .A1(_u10_u4_n2082 ), .A2(_u10_u4_n2050 ), .ZN(_u10_u4_n2847 ) );
NAND2_X1 _u10_u4_U645  ( .A1(_u10_u4_n2846 ), .A2(_u10_u4_n2847 ), .ZN(_u10_u4_n2074 ) );
NOR3_X1 _u10_u4_U644  ( .A1(_u10_u4_n2287 ), .A2(_u10_u4_n2596 ), .A3(_u10_u4_n2074 ), .ZN(_u10_u4_n2845 ) );
NAND4_X1 _u10_u4_U643  ( .A1(_u10_u4_n2357 ), .A2(_u10_u4_n2837 ), .A3(_u10_u4_n2844 ), .A4(_u10_u4_n2845 ), .ZN(_u10_u4_n2843 ) );
NAND2_X1 _u10_u4_U642  ( .A1(_u10_u4_n2279 ), .A2(_u10_u4_n2843 ), .ZN(_u10_u4_n2822 ) );
NOR3_X1 _u10_u4_U641  ( .A1(_u10_u4_n1925 ), .A2(_u10_u4_n2842 ), .A3(_u10_u4_n2686 ), .ZN(_u10_u4_n2841 ) );
NOR3_X1 _u10_u4_U640  ( .A1(_u10_u4_n2840 ), .A2(_u10_u4_n2599 ), .A3(_u10_u4_n2841 ), .ZN(_u10_u4_n2839 ) );
AND4_X1 _u10_u4_U639  ( .A1(_u10_u4_n2836 ), .A2(_u10_u4_n2837 ), .A3(_u10_u4_n2838 ), .A4(_u10_u4_n2839 ), .ZN(_u10_u4_n2454 ) );
NOR2_X1 _u10_u4_U638  ( .A1(_u10_u4_n2719 ), .A2(_u10_u4_n2835 ), .ZN(_u10_u4_n2773 ) );
NOR2_X1 _u10_u4_U637  ( .A1(_u10_u4_n2138 ), .A2(_u10_u4_n2773 ), .ZN(_u10_u4_n2814 ) );
NAND2_X1 _u10_u4_U636  ( .A1(_u10_u4_n2814 ), .A2(_u10_u4_n1869 ), .ZN(_u10_u4_n2834 ) );
NAND2_X1 _u10_u4_U635  ( .A1(_u10_u4_n2833 ), .A2(_u10_u4_n2834 ), .ZN(_u10_u4_n2832 ) );
NAND2_X1 _u10_u4_U634  ( .A1(_u10_u4_n2454 ), .A2(_u10_u4_n2832 ), .ZN(_u10_u4_n2831 ) );
NAND2_X1 _u10_u4_U633  ( .A1(_u10_u4_n2830 ), .A2(_u10_u4_n2831 ), .ZN(_u10_u4_n2823 ) );
INV_X1 _u10_u4_U632  ( .A(_u10_u4_n2025 ), .ZN(_u10_u4_n2470 ) );
NAND2_X1 _u10_u4_U631  ( .A1(_u10_u4_n1979 ), .A2(_u10_u4_n1936 ), .ZN(_u10_u4_n2829 ) );
AND2_X1 _u10_u4_U630  ( .A1(_u10_u4_n2828 ), .A2(_u10_u4_n2829 ), .ZN(_u10_u4_n2469 ) );
NAND2_X1 _u10_u4_U629  ( .A1(_u10_u4_n2469 ), .A2(_u10_u4_n2269 ), .ZN(_u10_u4_n2161 ) );
INV_X1 _u10_u4_U628  ( .A(_u10_u4_n2161 ), .ZN(_u10_u4_n2276 ) );
NOR2_X1 _u10_u4_U627  ( .A1(_u10_u4_n2274 ), .A2(_u10_u4_n2719 ), .ZN(_u10_u4_n2827 ) );
NOR3_X1 _u10_u4_U626  ( .A1(_u10_u4_n2827 ), .A2(_u10_u4_n2742 ), .A3(_u10_u4_n2680 ), .ZN(_u10_u4_n2826 ) );
NAND3_X1 _u10_u4_U625  ( .A1(_u10_u4_n2276 ), .A2(_u10_u4_n2108 ), .A3(_u10_u4_n2826 ), .ZN(_u10_u4_n2825 ) );
NAND2_X1 _u10_u4_U624  ( .A1(_u10_u4_n2470 ), .A2(_u10_u4_n2825 ), .ZN(_u10_u4_n2824 ) );
NAND4_X1 _u10_u4_U623  ( .A1(_u10_u4_n2821 ), .A2(_u10_u4_n2822 ), .A3(_u10_u4_n2823 ), .A4(_u10_u4_n2824 ), .ZN(_u10_u4_n2804 ) );
NAND2_X1 _u10_u4_U622  ( .A1(_u10_u4_n2131 ), .A2(_u10_u4_n2744 ), .ZN(_u10_u4_n2820 ) );
NAND2_X1 _u10_u4_U621  ( .A1(_u10_u4_n2571 ), .A2(_u10_u4_n2820 ), .ZN(_u10_u4_n2817 ) );
NOR2_X1 _u10_u4_U620  ( .A1(_u10_u4_n2819 ), .A2(_u10_u4_n2436 ), .ZN(_u10_u4_n2818 ) );
NAND4_X1 _u10_u4_U619  ( .A1(_u10_u4_n2437 ), .A2(_u10_u4_n2355 ), .A3(_u10_u4_n2817 ), .A4(_u10_u4_n2818 ), .ZN(_u10_u4_n2816 ) );
NAND2_X1 _u10_u4_U618  ( .A1(_u10_u4_n2815 ), .A2(_u10_u4_n2816 ), .ZN(_u10_u4_n2809 ) );
INV_X1 _u10_u4_U617  ( .A(_u10_u4_n2814 ), .ZN(_u10_u4_n2812 ) );
OR2_X1 _u10_u4_U616  ( .A1(_u10_u4_n1911 ), .A2(_u10_u4_n2813 ), .ZN(_u10_u4_n1884 ) );
NAND2_X1 _u10_u4_U615  ( .A1(_u10_u4_n2812 ), .A2(_u10_u4_n1884 ), .ZN(_u10_u4_n2810 ) );
NOR2_X1 _u10_u4_U614  ( .A1(_u10_u4_n1894 ), .A2(_u10_u4_n2461 ), .ZN(_u10_u4_n1948 ) );
OR2_X1 _u10_u4_U613  ( .A1(_u10_u4_n1847 ), .A2(_u10_u4_n1948 ), .ZN(_u10_u4_n2811 ) );
NAND3_X1 _u10_u4_U612  ( .A1(_u10_u4_n2809 ), .A2(_u10_u4_n2810 ), .A3(_u10_u4_n2811 ), .ZN(_u10_u4_n2805 ) );
NOR2_X1 _u10_u4_U611  ( .A1(_u10_u4_n2808 ), .A2(_u10_u4_n2775 ), .ZN(_u10_u4_n2806 ) );
AND2_X1 _u10_u4_U610  ( .A1(_u10_u4_n2721 ), .A2(_u10_u4_n1911 ), .ZN(_u10_u4_n2807 ) );
NOR4_X1 _u10_u4_U609  ( .A1(_u10_u4_n2804 ), .A2(_u10_u4_n2805 ), .A3(_u10_u4_n2806 ), .A4(_u10_u4_n2807 ), .ZN(_u10_u4_n2726 ) );
NAND2_X1 _u10_u4_U608  ( .A1(_u10_u4_n2803 ), .A2(_u10_u4_n2112 ), .ZN(_u10_u4_n2802 ) );
NAND2_X1 _u10_u4_U607  ( .A1(_u10_u4_n2364 ), .A2(_u10_u4_n2802 ), .ZN(_u10_u4_n2801 ) );
NAND2_X1 _u10_u4_U606  ( .A1(_u10_u4_n2800 ), .A2(_u10_u4_n2801 ), .ZN(_u10_u4_n2799 ) );
NAND2_X1 _u10_u4_U605  ( .A1(_u10_u4_n1937 ), .A2(_u10_u4_n2799 ), .ZN(_u10_u4_n2780 ) );
NAND2_X1 _u10_u4_U604  ( .A1(_u10_u4_n2775 ), .A2(_u10_u4_n2798 ), .ZN(_u10_u4_n2796 ) );
INV_X1 _u10_u4_U603  ( .A(_u10_u4_n2131 ), .ZN(_u10_u4_n2797 ) );
NAND2_X1 _u10_u4_U602  ( .A1(_u10_u4_n2796 ), .A2(_u10_u4_n2797 ), .ZN(_u10_u4_n2781 ) );
OR4_X1 _u10_u4_U601  ( .A1(_u10_u4_n2795 ), .A2(_u10_u4_n2303 ), .A3(_u10_u4_n2553 ), .A4(_u10_u4_n2554 ), .ZN(_u10_u4_n2792 ) );
NAND3_X1 _u10_u4_U600  ( .A1(_u10_u4_n1847 ), .A2(_u10_u4_n2097 ), .A3(_u10_u4_n2096 ), .ZN(_u10_u4_n2793 ) );
NOR4_X1 _u10_u4_U599  ( .A1(_u10_u4_n2792 ), .A2(_u10_u4_n2793 ), .A3(_u10_u4_n2542 ), .A4(_u10_u4_n2794 ), .ZN(_u10_u4_n2791 ) );
NOR2_X1 _u10_u4_U598  ( .A1(_u10_u4_n2791 ), .A2(_u10_u4_n2085 ), .ZN(_u10_u4_n2783 ) );
NAND2_X1 _u10_u4_U597  ( .A1(_u10_u4_n2114 ), .A2(_u10_u4_n2049 ), .ZN(_u10_u4_n2700 ) );
INV_X1 _u10_u4_U596  ( .A(_u10_u4_n2700 ), .ZN(_u10_u4_n2784 ) );
NAND4_X1 _u10_u4_U595  ( .A1(_u10_u4_n2001 ), .A2(_u10_u4_n2547 ), .A3(_u10_u4_n2368 ), .A4(_u10_u4_n1847 ), .ZN(_u10_u4_n2787 ) );
NOR4_X1 _u10_u4_U594  ( .A1(_u10_u4_n2787 ), .A2(_u10_u4_n2788 ), .A3(_u10_u4_n2789 ), .A4(_u10_u4_n2790 ), .ZN(_u10_u4_n2786 ) );
NOR2_X1 _u10_u4_U593  ( .A1(_u10_u4_n2786 ), .A2(_u10_u4_n2000 ), .ZN(_u10_u4_n2785 ) );
NOR3_X1 _u10_u4_U592  ( .A1(_u10_u4_n2783 ), .A2(_u10_u4_n2784 ), .A3(_u10_u4_n2785 ), .ZN(_u10_u4_n2782 ) );
NAND3_X1 _u10_u4_U591  ( .A1(_u10_u4_n2780 ), .A2(_u10_u4_n2781 ), .A3(_u10_u4_n2782 ), .ZN(_u10_u4_n2728 ) );
OR3_X1 _u10_u4_U590  ( .A1(_u10_u4_n2138 ), .A2(_u10_u4_n2633 ), .A3(_u10_u4_n2779 ), .ZN(_u10_u4_n2778 ) );
NAND2_X1 _u10_u4_U589  ( .A1(_u10_u4_n2777 ), .A2(_u10_u4_n2778 ), .ZN(_u10_u4_n2767 ) );
NAND3_X1 _u10_u4_U588  ( .A1(_u10_u4_n2775 ), .A2(_u10_u4_n2083 ), .A3(_u10_u4_n2776 ), .ZN(_u10_u4_n2774 ) );
NAND2_X1 _u10_u4_U587  ( .A1(_u10_u4_n2773 ), .A2(_u10_u4_n2774 ), .ZN(_u10_u4_n2768 ) );
NAND2_X1 _u10_u4_U586  ( .A1(_u10_u4_n2218 ), .A2(_u10_u4_n2772 ), .ZN(_u10_u4_n2769 ) );
NAND2_X1 _u10_u4_U585  ( .A1(_u10_u4_n2302 ), .A2(_u10_u4_n2467 ), .ZN(_u10_u4_n2771 ) );
NAND2_X1 _u10_u4_U584  ( .A1(_u10_u4_n2461 ), .A2(_u10_u4_n2771 ), .ZN(_u10_u4_n2770 ) );
NAND4_X1 _u10_u4_U583  ( .A1(_u10_u4_n2767 ), .A2(_u10_u4_n2768 ), .A3(_u10_u4_n2769 ), .A4(_u10_u4_n2770 ), .ZN(_u10_u4_n2729 ) );
NAND3_X1 _u10_u4_U582  ( .A1(_u10_u4_n2668 ), .A2(_u10_u4_n2600 ), .A3(_u10_u4_n2276 ), .ZN(_u10_u4_n2766 ) );
NAND2_X1 _u10_u4_U581  ( .A1(_u10_u4_n1894 ), .A2(_u10_u4_n2766 ), .ZN(_u10_u4_n2753 ) );
NAND3_X1 _u10_u4_U580  ( .A1(_u10_u4_n2456 ), .A2(_u10_u4_n2744 ), .A3(_u10_u4_n2765 ), .ZN(_u10_u4_n2764 ) );
NAND2_X1 _u10_u4_U579  ( .A1(_u10_u4_n2377 ), .A2(_u10_u4_n2764 ), .ZN(_u10_u4_n2754 ) );
NAND2_X1 _u10_u4_U578  ( .A1(_u10_u4_n2763 ), .A2(_u10_u4_n2007 ), .ZN(_u10_u4_n2755 ) );
NOR2_X1 _u10_u4_U577  ( .A1(_u10_u4_n2531 ), .A2(_u10_u4_n2744 ), .ZN(_u10_u4_n2760 ) );
INV_X1 _u10_u4_U576  ( .A(_u10_u4_n2762 ), .ZN(_u10_u4_n2189 ) );
NOR3_X1 _u10_u4_U575  ( .A1(_u10_u4_n2760 ), .A2(_u10_u4_n2761 ), .A3(_u10_u4_n2189 ), .ZN(_u10_u4_n2759 ) );
NOR2_X1 _u10_u4_U574  ( .A1(_u10_u4_n2759 ), .A2(_u10_u4_n1849 ), .ZN(_u10_u4_n2757 ) );
NOR2_X1 _u10_u4_U573  ( .A1(_u10_u4_n1817 ), .A2(_u10_u4_n2665 ), .ZN(_u10_u4_n2758 ) );
NOR2_X1 _u10_u4_U572  ( .A1(_u10_u4_n2757 ), .A2(_u10_u4_n2758 ), .ZN(_u10_u4_n2756 ) );
NAND4_X1 _u10_u4_U571  ( .A1(_u10_u4_n2753 ), .A2(_u10_u4_n2754 ), .A3(_u10_u4_n2755 ), .A4(_u10_u4_n2756 ), .ZN(_u10_u4_n2730 ) );
INV_X1 _u10_u4_U570  ( .A(_u10_u4_n2359 ), .ZN(_u10_u4_n1899 ) );
NAND4_X1 _u10_u4_U569  ( .A1(_u10_u4_n2078 ), .A2(_u10_u4_n2580 ), .A3(_u10_u4_n2748 ), .A4(_u10_u4_n2752 ), .ZN(_u10_u4_n2751 ) );
NAND2_X1 _u10_u4_U568  ( .A1(_u10_u4_n1899 ), .A2(_u10_u4_n2751 ), .ZN(_u10_u4_n2732 ) );
INV_X1 _u10_u4_U567  ( .A(_u10_u4_n2750 ), .ZN(_u10_u4_n2379 ) );
NAND3_X1 _u10_u4_U566  ( .A1(_u10_u4_n1856 ), .A2(_u10_u4_n2669 ), .A3(_u10_u4_n2364 ), .ZN(_u10_u4_n2749 ) );
AND2_X1 _u10_u4_U565  ( .A1(_u10_u4_n2748 ), .A2(_u10_u4_n2749 ), .ZN(_u10_u4_n2034 ) );
NAND2_X1 _u10_u4_U564  ( .A1(_u10_u4_n2105 ), .A2(_u10_u4_n2669 ), .ZN(_u10_u4_n2745 ) );
AND3_X1 _u10_u4_U563  ( .A1(_u10_u4_n2745 ), .A2(_u10_u4_n2746 ), .A3(_u10_u4_n2747 ), .ZN(_u10_u4_n2380 ) );
NOR2_X1 _u10_u4_U562  ( .A1(_u10_u4_n2274 ), .A2(_u10_u4_n2744 ), .ZN(_u10_u4_n2743 ) );
NOR4_X1 _u10_u4_U561  ( .A1(_u10_u4_n2742 ), .A2(_u10_u4_n2680 ), .A3(_u10_u4_n2743 ), .A4(_u10_u4_n2428 ), .ZN(_u10_u4_n2741 ) );
NAND4_X1 _u10_u4_U560  ( .A1(_u10_u4_n2379 ), .A2(_u10_u4_n2034 ), .A3(_u10_u4_n2380 ), .A4(_u10_u4_n2741 ), .ZN(_u10_u4_n2740 ) );
NAND2_X1 _u10_u4_U559  ( .A1(_u10_u4_n1967 ), .A2(_u10_u4_n2740 ), .ZN(_u10_u4_n2733 ) );
NAND3_X1 _u10_u4_U558  ( .A1(_u10_u4_n2739 ), .A2(_u10_u4_n2368 ), .A3(_u10_u4_n2255 ), .ZN(_u10_u4_n2738 ) );
NAND2_X1 _u10_u4_U557  ( .A1(_u10_u4_n2737 ), .A2(_u10_u4_n2738 ), .ZN(_u10_u4_n2734 ) );
NAND2_X1 _u10_u4_U556  ( .A1(_u10_u4_n2736 ), .A2(_u10_u4_n2524 ), .ZN(_u10_u4_n2735 ) );
NAND4_X1 _u10_u4_U555  ( .A1(_u10_u4_n2732 ), .A2(_u10_u4_n2733 ), .A3(_u10_u4_n2734 ), .A4(_u10_u4_n2735 ), .ZN(_u10_u4_n2731 ) );
NOR4_X1 _u10_u4_U554  ( .A1(_u10_u4_n2728 ), .A2(_u10_u4_n2729 ), .A3(_u10_u4_n2730 ), .A4(_u10_u4_n2731 ), .ZN(_u10_u4_n2727 ) );
NAND4_X1 _u10_u4_U553  ( .A1(_u10_u4_n2724 ), .A2(_u10_u4_n2725 ), .A3(_u10_u4_n2726 ), .A4(_u10_u4_n2727 ), .ZN(_u10_u4_n2723 ) );
MUX2_X1 _u10_u4_U552  ( .A(_u10_u4_n2723 ), .B(_u10_SYNOPSYS_UNCONNECTED_14 ), .S(_u10_u4_n1819 ), .Z(_u10_u4_n1809 ) );
NAND2_X1 _u10_u4_U551  ( .A1(_u10_u4_n2002 ), .A2(_u10_u4_n2722 ), .ZN(_u10_u4_n2713 ) );
NAND2_X1 _u10_u4_U550  ( .A1(_u10_u4_n2720 ), .A2(_u10_u4_n2721 ), .ZN(_u10_u4_n2714 ) );
NAND2_X1 _u10_u4_U549  ( .A1(_u10_u4_n2256 ), .A2(_u10_u4_n2719 ), .ZN(_u10_u4_n2715 ) );
NOR2_X1 _u10_u4_U548  ( .A1(_u10_u4_n2106 ), .A2(_u10_u4_n2037 ), .ZN(_u10_u4_n2717 ) );
AND2_X1 _u10_u4_U547  ( .A1(_u10_u4_n1966 ), .A2(_u10_u4_n2054 ), .ZN(_u10_u4_n2718 ) );
NOR2_X1 _u10_u4_U546  ( .A1(_u10_u4_n2717 ), .A2(_u10_u4_n2718 ), .ZN(_u10_u4_n2716 ) );
NAND4_X1 _u10_u4_U545  ( .A1(_u10_u4_n2713 ), .A2(_u10_u4_n2714 ), .A3(_u10_u4_n2715 ), .A4(_u10_u4_n2716 ), .ZN(_u10_u4_n2608 ) );
NAND2_X1 _u10_u4_U544  ( .A1(1'b0), .A2(_u10_u4_n2669 ), .ZN(_u10_u4_n2385 ));
INV_X1 _u10_u4_U543  ( .A(_u10_u4_n2385 ), .ZN(_u10_u4_n1977 ) );
NAND2_X1 _u10_u4_U542  ( .A1(_u10_u4_n1977 ), .A2(_u10_u4_n2668 ), .ZN(_u10_u4_n2712 ) );
NAND2_X1 _u10_u4_U541  ( .A1(_u10_u4_n2712 ), .A2(_u10_u4_n2092 ), .ZN(_u10_u4_n1844 ) );
NAND2_X1 _u10_u4_U540  ( .A1(_u10_u4_n1894 ), .A2(_u10_u4_n1844 ), .ZN(_u10_u4_n2705 ) );
NAND2_X1 _u10_u4_U539  ( .A1(_u10_u4_n1894 ), .A2(_u10_u4_n2305 ), .ZN(_u10_u4_n2711 ) );
NAND2_X1 _u10_u4_U538  ( .A1(_u10_u4_n2711 ), .A2(_u10_u4_n2025 ), .ZN(_u10_u4_n1932 ) );
NAND2_X1 _u10_u4_U537  ( .A1(_u10_u4_n2710 ), .A2(_u10_u4_n1932 ), .ZN(_u10_u4_n2706 ) );
NAND2_X1 _u10_u4_U536  ( .A1(_u10_u4_n2708 ), .A2(_u10_u4_n2709 ), .ZN(_u10_u4_n2707 ) );
NAND3_X1 _u10_u4_U535  ( .A1(_u10_u4_n2705 ), .A2(_u10_u4_n2706 ), .A3(_u10_u4_n2707 ), .ZN(_u10_u4_n2701 ) );
NOR2_X1 _u10_u4_U534  ( .A1(_u10_u4_n1843 ), .A2(_u10_u4_n2545 ), .ZN(_u10_u4_n2702 ) );
NOR2_X1 _u10_u4_U533  ( .A1(_u10_u4_n2346 ), .A2(_u10_u4_n2700 ), .ZN(_u10_u4_n2703 ) );
NOR2_X1 _u10_u4_U532  ( .A1(_u10_u4_n2000 ), .A2(_u10_u4_n1887 ), .ZN(_u10_u4_n2704 ) );
NOR4_X1 _u10_u4_U531  ( .A1(_u10_u4_n2701 ), .A2(_u10_u4_n2702 ), .A3(_u10_u4_n2703 ), .A4(_u10_u4_n2704 ), .ZN(_u10_u4_n2671 ) );
NAND2_X1 _u10_u4_U530  ( .A1(_u10_u4_n2699 ), .A2(_u10_u4_n2700 ), .ZN(_u10_u4_n2698 ) );
NAND2_X1 _u10_u4_U529  ( .A1(_u10_u4_n2063 ), .A2(_u10_u4_n2698 ), .ZN(_u10_u4_n2682 ) );
NAND2_X1 _u10_u4_U528  ( .A1(_u10_u4_n2697 ), .A2(_u10_u4_n2103 ), .ZN(_u10_u4_n2696 ) );
NAND2_X1 _u10_u4_U527  ( .A1(_u10_u4_n2695 ), .A2(_u10_u4_n2696 ), .ZN(_u10_u4_n2694 ) );
NAND2_X1 _u10_u4_U526  ( .A1(_u10_u4_n1937 ), .A2(_u10_u4_n2694 ), .ZN(_u10_u4_n2683 ) );
INV_X1 _u10_u4_U525  ( .A(_u10_u4_n2693 ), .ZN(_u10_u4_n2691 ) );
NAND3_X1 _u10_u4_U524  ( .A1(_u10_u4_n2103 ), .A2(_u10_u4_n2502 ), .A3(1'b0),.ZN(_u10_u4_n2692 ) );
NAND2_X1 _u10_u4_U523  ( .A1(_u10_u4_n2691 ), .A2(_u10_u4_n2692 ), .ZN(_u10_u4_n2690 ) );
NAND2_X1 _u10_u4_U522  ( .A1(_u10_u4_n2236 ), .A2(_u10_u4_n2690 ), .ZN(_u10_u4_n2684 ) );
NAND3_X1 _u10_u4_U521  ( .A1(_u10_u4_n2688 ), .A2(_u10_u4_n1913 ), .A3(_u10_u4_n2689 ), .ZN(_u10_u4_n2335 ) );
NAND3_X1 _u10_u4_U520  ( .A1(_u10_u4_n2536 ), .A2(_u10_u4_n2103 ), .A3(1'b0),.ZN(_u10_u4_n2052 ) );
NOR2_X1 _u10_u4_U519  ( .A1(_u10_u4_n2052 ), .A2(_u10_u4_n2687 ), .ZN(_u10_u4_n1851 ) );
NAND2_X1 _u10_u4_U518  ( .A1(_u10_u4_n1851 ), .A2(_u10_u4_n2078 ), .ZN(_u10_u4_n2582 ) );
NOR2_X1 _u10_u4_U517  ( .A1(_u10_u4_n2686 ), .A2(_u10_u4_n2582 ), .ZN(_u10_u4_n2094 ) );
NAND3_X1 _u10_u4_U516  ( .A1(_u10_u4_n2251 ), .A2(_u10_u4_n2335 ), .A3(_u10_u4_n2094 ), .ZN(_u10_u4_n2685 ) );
NAND4_X1 _u10_u4_U515  ( .A1(_u10_u4_n2682 ), .A2(_u10_u4_n2683 ), .A3(_u10_u4_n2684 ), .A4(_u10_u4_n2685 ), .ZN(_u10_u4_n2673 ) );
INV_X1 _u10_u4_U514  ( .A(_u10_u4_n2291 ), .ZN(_u10_u4_n2057 ) );
AND2_X1 _u10_u4_U513  ( .A1(_u10_u4_n1851 ), .A2(_u10_u4_n2057 ), .ZN(_u10_u4_n2674 ) );
INV_X1 _u10_u4_U512  ( .A(_u10_u4_n1874 ), .ZN(_u10_u4_n2681 ) );
NOR2_X1 _u10_u4_U511  ( .A1(_u10_u4_n2007 ), .A2(_u10_u4_n1911 ), .ZN(_u10_u4_n2486 ) );
NOR2_X1 _u10_u4_U510  ( .A1(_u10_u4_n2681 ), .A2(_u10_u4_n2486 ), .ZN(_u10_u4_n2675 ) );
NOR2_X1 _u10_u4_U509  ( .A1(_u10_u4_n1977 ), .A2(_u10_u4_n2680 ), .ZN(_u10_u4_n2679 ) );
NOR2_X1 _u10_u4_U508  ( .A1(_u10_u4_n2679 ), .A2(_u10_u4_n2030 ), .ZN(_u10_u4_n2678 ) );
NOR2_X1 _u10_u4_U507  ( .A1(_u10_u4_n2678 ), .A2(_u10_u4_n2094 ), .ZN(_u10_u4_n2677 ) );
NOR2_X1 _u10_u4_U506  ( .A1(_u10_u4_n2677 ), .A2(_u10_u4_n2025 ), .ZN(_u10_u4_n2676 ) );
NOR4_X1 _u10_u4_U505  ( .A1(_u10_u4_n2673 ), .A2(_u10_u4_n2674 ), .A3(_u10_u4_n2675 ), .A4(_u10_u4_n2676 ), .ZN(_u10_u4_n2672 ) );
AND2_X1 _u10_u4_U504  ( .A1(_u10_u4_n2671 ), .A2(_u10_u4_n2672 ), .ZN(_u10_u4_n1990 ) );
INV_X1 _u10_u4_U503  ( .A(_u10_u4_n2670 ), .ZN(_u10_u4_n2660 ) );
NAND4_X1 _u10_u4_U502  ( .A1(_u10_u4_n2251 ), .A2(_u10_u4_n2669 ), .A3(_u10_u4_n2162 ), .A4(_u10_u4_n2169 ), .ZN(_u10_u4_n2664 ) );
AND3_X1 _u10_u4_U501  ( .A1(_u10_u4_n1977 ), .A2(_u10_u4_n2668 ), .A3(_u10_u4_n2089 ), .ZN(_u10_u4_n2555 ) );
NAND2_X1 _u10_u4_U500  ( .A1(_u10_u4_n2555 ), .A2(_u10_u4_n2667 ), .ZN(_u10_u4_n2666 ) );
NAND3_X1 _u10_u4_U499  ( .A1(_u10_u4_n2664 ), .A2(_u10_u4_n2665 ), .A3(_u10_u4_n2666 ), .ZN(_u10_u4_n1988 ) );
INV_X1 _u10_u4_U498  ( .A(_u10_u4_n1988 ), .ZN(_u10_u4_n2661 ) );
NAND2_X1 _u10_u4_U497  ( .A1(1'b0), .A2(_u10_u4_n2043 ), .ZN(_u10_u4_n2662 ));
NAND2_X1 _u10_u4_U496  ( .A1(_u10_u4_n2169 ), .A2(1'b0), .ZN(_u10_u4_n2663 ));
NAND4_X1 _u10_u4_U495  ( .A1(_u10_u4_n2660 ), .A2(_u10_u4_n2661 ), .A3(_u10_u4_n2662 ), .A4(_u10_u4_n2663 ), .ZN(_u10_u4_n2650 ) );
NAND2_X1 _u10_u4_U494  ( .A1(_u10_u4_n2659 ), .A2(1'b0), .ZN(_u10_u4_n2193 ));
INV_X1 _u10_u4_U493  ( .A(_u10_u4_n2193 ), .ZN(_u10_u4_n2143 ) );
NAND2_X1 _u10_u4_U492  ( .A1(_u10_u4_n2143 ), .A2(_u10_u4_n2036 ), .ZN(_u10_u4_n2286 ) );
INV_X1 _u10_u4_U491  ( .A(_u10_u4_n2286 ), .ZN(_u10_u4_n2577 ) );
NAND2_X1 _u10_u4_U490  ( .A1(_u10_u4_n2577 ), .A2(_u10_u4_n2278 ), .ZN(_u10_u4_n2474 ) );
INV_X1 _u10_u4_U489  ( .A(_u10_u4_n2474 ), .ZN(_u10_u4_n2306 ) );
NAND2_X1 _u10_u4_U488  ( .A1(_u10_u4_n2306 ), .A2(_u10_u4_n2251 ), .ZN(_u10_u4_n2654 ) );
NAND2_X1 _u10_u4_U487  ( .A1(_u10_u4_n2649 ), .A2(_u10_u4_n2658 ), .ZN(_u10_u4_n2655 ) );
NAND2_X1 _u10_u4_U486  ( .A1(_u10_u4_n2657 ), .A2(_u10_u4_n2445 ), .ZN(_u10_u4_n2656 ) );
NAND3_X1 _u10_u4_U485  ( .A1(_u10_u4_n2654 ), .A2(_u10_u4_n2655 ), .A3(_u10_u4_n2656 ), .ZN(_u10_u4_n2651 ) );
NOR2_X1 _u10_u4_U484  ( .A1(_u10_u4_n2366 ), .A2(_u10_u4_n2376 ), .ZN(_u10_u4_n2652 ) );
AND2_X1 _u10_u4_U483  ( .A1(_u10_u4_n1966 ), .A2(_u10_u4_n2528 ), .ZN(_u10_u4_n2653 ) );
NOR4_X1 _u10_u4_U482  ( .A1(_u10_u4_n2650 ), .A2(_u10_u4_n2651 ), .A3(_u10_u4_n2652 ), .A4(_u10_u4_n2653 ), .ZN(_u10_u4_n2613 ) );
NAND2_X1 _u10_u4_U481  ( .A1(_u10_u4_n1891 ), .A2(1'b0), .ZN(_u10_u4_n2636 ));
NAND2_X1 _u10_u4_U480  ( .A1(_u10_u4_n1868 ), .A2(_u10_u4_n2113 ), .ZN(_u10_u4_n2101 ) );
NOR4_X1 _u10_u4_U479  ( .A1(_u10_u4_n2649 ), .A2(_u10_u4_n2216 ), .A3(_u10_u4_n2101 ), .A4(_u10_u4_n2634 ), .ZN(_u10_u4_n2648 ) );
NOR2_X1 _u10_u4_U478  ( .A1(_u10_u4_n2648 ), .A2(_u10_u4_n2254 ), .ZN(_u10_u4_n2638 ) );
NOR2_X1 _u10_u4_U477  ( .A1(_u10_u4_n2106 ), .A2(_u10_u4_n2643 ), .ZN(_u10_u4_n2645 ) );
NAND2_X1 _u10_u4_U476  ( .A1(1'b0), .A2(_u10_u4_n2049 ), .ZN(_u10_u4_n2647 ));
NAND2_X1 _u10_u4_U475  ( .A1(_u10_u4_n2646 ), .A2(_u10_u4_n2647 ), .ZN(_u10_u4_n2348 ) );
NOR2_X1 _u10_u4_U474  ( .A1(_u10_u4_n2645 ), .A2(_u10_u4_n2348 ), .ZN(_u10_u4_n2644 ) );
NOR2_X1 _u10_u4_U473  ( .A1(_u10_u4_n2644 ), .A2(_u10_u4_n2495 ), .ZN(_u10_u4_n2639 ) );
NOR2_X1 _u10_u4_U472  ( .A1(_u10_u4_n2643 ), .A2(_u10_u4_n2203 ), .ZN(_u10_u4_n2642 ) );
NOR3_X1 _u10_u4_U471  ( .A1(_u10_u4_n2101 ), .A2(1'b0), .A3(_u10_u4_n2642 ),.ZN(_u10_u4_n2641 ) );
NOR2_X1 _u10_u4_U470  ( .A1(_u10_u4_n2641 ), .A2(_u10_u4_n2253 ), .ZN(_u10_u4_n2640 ) );
NOR3_X1 _u10_u4_U469  ( .A1(_u10_u4_n2638 ), .A2(_u10_u4_n2639 ), .A3(_u10_u4_n2640 ), .ZN(_u10_u4_n2637 ) );
NAND3_X1 _u10_u4_U468  ( .A1(_u10_u4_n2635 ), .A2(_u10_u4_n2636 ), .A3(_u10_u4_n2637 ), .ZN(_u10_u4_n2615 ) );
NOR3_X1 _u10_u4_U467  ( .A1(_u10_u4_n2174 ), .A2(_u10_u4_n2175 ), .A3(_u10_u4_n2179 ), .ZN(_u10_u4_n2631 ) );
NAND3_X1 _u10_u4_U466  ( .A1(_u10_u4_n2223 ), .A2(_u10_u4_n2236 ), .A3(_u10_u4_n2631 ), .ZN(_u10_u4_n2622 ) );
OR2_X1 _u10_u4_U465  ( .A1(_u10_u4_n1960 ), .A2(_u10_u4_n1959 ), .ZN(_u10_u4_n2625 ) );
NOR3_X1 _u10_u4_U464  ( .A1(_u10_u4_n2101 ), .A2(_u10_u4_n2633 ), .A3(_u10_u4_n2634 ), .ZN(_u10_u4_n2523 ) );
OR2_X1 _u10_u4_U463  ( .A1(_u10_u4_n2632 ), .A2(_u10_u4_n2523 ), .ZN(_u10_u4_n2627 ) );
INV_X1 _u10_u4_U462  ( .A(_u10_u4_n2631 ), .ZN(_u10_u4_n2628 ) );
NAND2_X1 _u10_u4_U461  ( .A1(_u10_u4_n2630 ), .A2(_u10_u4_n1922 ), .ZN(_u10_u4_n2629 ) );
NAND3_X1 _u10_u4_U460  ( .A1(_u10_u4_n2627 ), .A2(_u10_u4_n2628 ), .A3(_u10_u4_n2629 ), .ZN(_u10_u4_n2626 ) );
NAND2_X1 _u10_u4_U459  ( .A1(_u10_u4_n2625 ), .A2(_u10_u4_n2626 ), .ZN(_u10_u4_n2624 ) );
NAND3_X1 _u10_u4_U458  ( .A1(_u10_u4_n2622 ), .A2(_u10_u4_n2623 ), .A3(_u10_u4_n2624 ), .ZN(_u10_u4_n2616 ) );
AND2_X1 _u10_u4_U457  ( .A1(_u10_u4_n2621 ), .A2(_u10_u4_n2358 ), .ZN(_u10_u4_n2620 ) );
NOR2_X1 _u10_u4_U456  ( .A1(_u10_u4_n2523 ), .A2(_u10_u4_n2620 ), .ZN(_u10_u4_n2617 ) );
INV_X1 _u10_u4_U455  ( .A(_u10_u4_n2101 ), .ZN(_u10_u4_n2221 ) );
NOR2_X1 _u10_u4_U454  ( .A1(_u10_u4_n1911 ), .A2(_u10_u4_n2488 ), .ZN(_u10_u4_n2619 ) );
NOR2_X1 _u10_u4_U453  ( .A1(_u10_u4_n2221 ), .A2(_u10_u4_n2619 ), .ZN(_u10_u4_n2618 ) );
NOR4_X1 _u10_u4_U452  ( .A1(_u10_u4_n2615 ), .A2(_u10_u4_n2616 ), .A3(_u10_u4_n2617 ), .A4(_u10_u4_n2618 ), .ZN(_u10_u4_n2614 ) );
AND2_X1 _u10_u4_U451  ( .A1(_u10_u4_n2613 ), .A2(_u10_u4_n2614 ), .ZN(_u10_u4_n2314 ) );
NAND3_X1 _u10_u4_U450  ( .A1(_u10_u4_n2612 ), .A2(_u10_u4_n1990 ), .A3(_u10_u4_n2314 ), .ZN(_u10_u4_n2609 ) );
NOR4_X1 _u10_u4_U449  ( .A1(_u10_u4_n2608 ), .A2(_u10_u4_n2609 ), .A3(_u10_u4_n2610 ), .A4(_u10_u4_n2611 ), .ZN(_u10_u4_n2388 ) );
NAND2_X1 _u10_u4_U448  ( .A1(_u10_u4_n2346 ), .A2(_u10_u4_n2607 ), .ZN(_u10_u4_n2191 ) );
NAND2_X1 _u10_u4_U447  ( .A1(_u10_u4_n2143 ), .A2(_u10_u4_n2191 ), .ZN(_u10_u4_n2556 ) );
INV_X1 _u10_u4_U446  ( .A(_u10_u4_n2348 ), .ZN(_u10_u4_n2603 ) );
NAND3_X1 _u10_u4_U445  ( .A1(_u10_u4_n2535 ), .A2(_u10_u4_n2485 ), .A3(_u10_u4_n2456 ), .ZN(_u10_u4_n2606 ) );
NAND2_X1 _u10_u4_U444  ( .A1(_u10_u4_n2049 ), .A2(_u10_u4_n2606 ), .ZN(_u10_u4_n2604 ) );
NAND3_X1 _u10_u4_U443  ( .A1(_u10_u4_n2603 ), .A2(_u10_u4_n2604 ), .A3(_u10_u4_n2605 ), .ZN(_u10_u4_n2602 ) );
NAND2_X1 _u10_u4_U442  ( .A1(_u10_u4_n2043 ), .A2(_u10_u4_n2602 ), .ZN(_u10_u4_n2557 ) );
INV_X1 _u10_u4_U441  ( .A(_u10_u4_n2601 ), .ZN(_u10_u4_n2590 ) );
NAND2_X1 _u10_u4_U440  ( .A1(_u10_u4_n2599 ), .A2(_u10_u4_n2600 ), .ZN(_u10_u4_n2597 ) );
NAND2_X1 _u10_u4_U439  ( .A1(_u10_u4_n2082 ), .A2(_u10_u4_n2101 ), .ZN(_u10_u4_n2598 ) );
AND2_X1 _u10_u4_U438  ( .A1(_u10_u4_n2597 ), .A2(_u10_u4_n2598 ), .ZN(_u10_u4_n2281 ) );
NAND3_X1 _u10_u4_U437  ( .A1(_u10_u4_n1969 ), .A2(_u10_u4_n2582 ), .A3(_u10_u4_n2281 ), .ZN(_u10_u4_n2073 ) );
INV_X1 _u10_u4_U436  ( .A(_u10_u4_n2073 ), .ZN(_u10_u4_n2591 ) );
NOR2_X1 _u10_u4_U435  ( .A1(_u10_u4_n1816 ), .A2(_u10_u4_n2077 ), .ZN(_u10_u4_n2595 ) );
NOR2_X1 _u10_u4_U434  ( .A1(_u10_u4_n2595 ), .A2(_u10_u4_n2596 ), .ZN(_u10_u4_n2592 ) );
NAND3_X1 _u10_u4_U433  ( .A1(_u10_u4_n2107 ), .A2(_u10_u4_n2536 ), .A3(1'b0),.ZN(_u10_u4_n2438 ) );
INV_X1 _u10_u4_U432  ( .A(_u10_u4_n2438 ), .ZN(_u10_u4_n2427 ) );
NOR4_X1 _u10_u4_U431  ( .A1(1'b0), .A2(_u10_u4_n2594 ), .A3(_u10_u4_n2577 ),.A4(_u10_u4_n2427 ), .ZN(_u10_u4_n2593 ) );
NAND4_X1 _u10_u4_U430  ( .A1(_u10_u4_n2590 ), .A2(_u10_u4_n2591 ), .A3(_u10_u4_n2592 ), .A4(_u10_u4_n2593 ), .ZN(_u10_u4_n2589 ) );
NAND2_X1 _u10_u4_U429  ( .A1(_u10_u4_n2279 ), .A2(_u10_u4_n2589 ), .ZN(_u10_u4_n2558 ) );
NAND3_X1 _u10_u4_U428  ( .A1(_u10_u4_n2587 ), .A2(_u10_u4_n2115 ), .A3(_u10_u4_n2588 ), .ZN(_u10_u4_n2585 ) );
NOR4_X1 _u10_u4_U427  ( .A1(_u10_u4_n2585 ), .A2(_u10_u4_n2586 ), .A3(1'b0),.A4(_u10_u4_n2114 ), .ZN(_u10_u4_n2583 ) );
NOR2_X1 _u10_u4_U426  ( .A1(_u10_u4_n2583 ), .A2(_u10_u4_n2584 ), .ZN(_u10_u4_n2560 ) );
OR2_X1 _u10_u4_U425  ( .A1(_u10_u4_n2582 ), .A2(1'b0), .ZN(_u10_u4_n2581 ));
NAND2_X1 _u10_u4_U424  ( .A1(_u10_u4_n2580 ), .A2(_u10_u4_n2581 ), .ZN(_u10_u4_n1974 ) );
INV_X1 _u10_u4_U423  ( .A(_u10_u4_n1974 ), .ZN(_u10_u4_n1901 ) );
AND4_X1 _u10_u4_U422  ( .A1(_u10_u4_n1901 ), .A2(_u10_u4_n2385 ), .A3(_u10_u4_n2578 ), .A4(_u10_u4_n2579 ), .ZN(_u10_u4_n2424 ) );
NOR2_X1 _u10_u4_U421  ( .A1(1'b0), .A2(_u10_u4_n2424 ), .ZN(_u10_u4_n2574 ));
NOR3_X1 _u10_u4_U420  ( .A1(_u10_u4_n2427 ), .A2(1'b0), .A3(_u10_u4_n2577 ),.ZN(_u10_u4_n2576 ) );
NOR2_X1 _u10_u4_U419  ( .A1(_u10_u4_n2576 ), .A2(_u10_u4_n1976 ), .ZN(_u10_u4_n2575 ) );
NOR3_X1 _u10_u4_U418  ( .A1(_u10_u4_n2574 ), .A2(_u10_u4_n1979 ), .A3(_u10_u4_n2575 ), .ZN(_u10_u4_n2572 ) );
NOR2_X1 _u10_u4_U417  ( .A1(_u10_u4_n2572 ), .A2(_u10_u4_n2573 ), .ZN(_u10_u4_n2561 ) );
INV_X1 _u10_u4_U416  ( .A(_u10_u4_n2061 ), .ZN(_u10_u4_n2453 ) );
NOR2_X1 _u10_u4_U415  ( .A1(_u10_u4_n2453 ), .A2(_u10_u4_n1851 ), .ZN(_u10_u4_n2018 ) );
NAND2_X1 _u10_u4_U414  ( .A1(1'b0), .A2(_u10_u4_n2571 ), .ZN(_u10_u4_n2570 ));
NAND2_X1 _u10_u4_U413  ( .A1(_u10_u4_n2018 ), .A2(_u10_u4_n2570 ), .ZN(_u10_u4_n1837 ) );
INV_X1 _u10_u4_U412  ( .A(_u10_u4_n1837 ), .ZN(_u10_u4_n2568 ) );
NAND2_X1 _u10_u4_U411  ( .A1(1'b0), .A2(_u10_u4_n2536 ), .ZN(_u10_u4_n2569 ));
NAND2_X1 _u10_u4_U410  ( .A1(_u10_u4_n2568 ), .A2(_u10_u4_n2569 ), .ZN(_u10_u4_n2564 ) );
NOR2_X1 _u10_u4_U409  ( .A1(_u10_u4_n1841 ), .A2(_u10_u4_n1868 ), .ZN(_u10_u4_n2565 ) );
INV_X1 _u10_u4_U408  ( .A(_u10_u4_n2567 ), .ZN(_u10_u4_n2566 ) );
NOR4_X1 _u10_u4_U407  ( .A1(_u10_u4_n2564 ), .A2(_u10_u4_n2565 ), .A3(_u10_u4_n2143 ), .A4(_u10_u4_n2566 ), .ZN(_u10_u4_n2563 ) );
NOR2_X1 _u10_u4_U406  ( .A1(_u10_u4_n2563 ), .A2(_u10_u4_n2014 ), .ZN(_u10_u4_n2562 ) );
NOR3_X1 _u10_u4_U405  ( .A1(_u10_u4_n2560 ), .A2(_u10_u4_n2561 ), .A3(_u10_u4_n2562 ), .ZN(_u10_u4_n2559 ) );
NAND4_X1 _u10_u4_U404  ( .A1(_u10_u4_n2556 ), .A2(_u10_u4_n2557 ), .A3(_u10_u4_n2558 ), .A4(_u10_u4_n2559 ), .ZN(_u10_u4_n2511 ) );
INV_X1 _u10_u4_U403  ( .A(_u10_u4_n2085 ), .ZN(_u10_u4_n2293 ) );
NOR2_X1 _u10_u4_U402  ( .A1(_u10_u4_n2554 ), .A2(_u10_u4_n2555 ), .ZN(_u10_u4_n2444 ) );
NAND2_X1 _u10_u4_U401  ( .A1(_u10_u4_n2553 ), .A2(_u10_u4_n2549 ), .ZN(_u10_u4_n2552 ) );
AND2_X1 _u10_u4_U400  ( .A1(_u10_u4_n2444 ), .A2(_u10_u4_n2552 ), .ZN(_u10_u4_n2295 ) );
NAND2_X1 _u10_u4_U399  ( .A1(_u10_u4_n2551 ), .A2(_u10_u4_n2549 ), .ZN(_u10_u4_n2538 ) );
AND2_X1 _u10_u4_U398  ( .A1(_u10_u4_n2427 ), .A2(_u10_u4_n2108 ), .ZN(_u10_u4_n2460 ) );
NOR4_X1 _u10_u4_U397  ( .A1(_u10_u4_n2460 ), .A2(_u10_u4_n2306 ), .A3(_u10_u4_n2094 ), .A4(_u10_u4_n2550 ), .ZN(_u10_u4_n2409 ) );
INV_X1 _u10_u4_U396  ( .A(_u10_u4_n2409 ), .ZN(_u10_u4_n2407 ) );
NAND2_X1 _u10_u4_U395  ( .A1(_u10_u4_n2549 ), .A2(_u10_u4_n2407 ), .ZN(_u10_u4_n2546 ) );
NAND3_X1 _u10_u4_U394  ( .A1(_u10_u4_n2546 ), .A2(_u10_u4_n2547 ), .A3(_u10_u4_n2548 ), .ZN(_u10_u4_n2501 ) );
INV_X1 _u10_u4_U393  ( .A(_u10_u4_n2501 ), .ZN(_u10_u4_n2539 ) );
NOR2_X1 _u10_u4_U392  ( .A1(1'b0), .A2(_u10_u4_n2545 ), .ZN(_u10_u4_n2541 ));
AND2_X1 _u10_u4_U391  ( .A1(_u10_u4_n2544 ), .A2(_u10_u4_n2089 ), .ZN(_u10_u4_n2543 ) );
NOR3_X1 _u10_u4_U390  ( .A1(_u10_u4_n2541 ), .A2(_u10_u4_n2542 ), .A3(_u10_u4_n2543 ), .ZN(_u10_u4_n2540 ) );
NAND4_X1 _u10_u4_U389  ( .A1(_u10_u4_n2295 ), .A2(_u10_u4_n2538 ), .A3(_u10_u4_n2539 ), .A4(_u10_u4_n2540 ), .ZN(_u10_u4_n2537 ) );
NAND2_X1 _u10_u4_U388  ( .A1(_u10_u4_n2293 ), .A2(_u10_u4_n2537 ), .ZN(_u10_u4_n2515 ) );
NAND2_X1 _u10_u4_U387  ( .A1(_u10_u4_n2536 ), .A2(_u10_u4_n2508 ), .ZN(_u10_u4_n2526 ) );
NAND2_X1 _u10_u4_U386  ( .A1(_u10_u4_n2535 ), .A2(_u10_u4_n1940 ), .ZN(_u10_u4_n2532 ) );
NOR4_X1 _u10_u4_U385  ( .A1(_u10_u4_n2532 ), .A2(_u10_u4_n2533 ), .A3(1'b0),.A4(_u10_u4_n2534 ), .ZN(_u10_u4_n2530 ) );
NOR2_X1 _u10_u4_U384  ( .A1(_u10_u4_n2530 ), .A2(_u10_u4_n2531 ), .ZN(_u10_u4_n2529 ) );
NOR4_X1 _u10_u4_U383  ( .A1(_u10_u4_n2528 ), .A2(_u10_u4_n2143 ), .A3(_u10_u4_n2189 ), .A4(_u10_u4_n2529 ), .ZN(_u10_u4_n2527 ) );
NAND4_X1 _u10_u4_U382  ( .A1(_u10_u4_n2019 ), .A2(_u10_u4_n2526 ), .A3(_u10_u4_n2018 ), .A4(_u10_u4_n2527 ), .ZN(_u10_u4_n2525 ) );
NAND2_X1 _u10_u4_U381  ( .A1(_u10_u4_n2183 ), .A2(_u10_u4_n2525 ), .ZN(_u10_u4_n2516 ) );
INV_X1 _u10_u4_U380  ( .A(_u10_u4_n2524 ), .ZN(_u10_u4_n2396 ) );
NAND2_X1 _u10_u4_U379  ( .A1(_u10_u4_n2396 ), .A2(_u10_u4_n2523 ), .ZN(_u10_u4_n2522 ) );
NAND2_X1 _u10_u4_U378  ( .A1(_u10_u4_n1866 ), .A2(_u10_u4_n2522 ), .ZN(_u10_u4_n2519 ) );
AND2_X1 _u10_u4_U377  ( .A1(_u10_u4_n2493 ), .A2(_u10_u4_n1961 ), .ZN(_u10_u4_n2429 ) );
NAND2_X1 _u10_u4_U376  ( .A1(_u10_u4_n2429 ), .A2(_u10_u4_n2175 ), .ZN(_u10_u4_n2510 ) );
NAND2_X1 _u10_u4_U375  ( .A1(_u10_u4_n2510 ), .A2(_u10_u4_n1864 ), .ZN(_u10_u4_n2521 ) );
NAND3_X1 _u10_u4_U374  ( .A1(_u10_u4_n2519 ), .A2(_u10_u4_n2520 ), .A3(_u10_u4_n2521 ), .ZN(_u10_u4_n2518 ) );
NAND2_X1 _u10_u4_U373  ( .A1(_u10_u4_n1861 ), .A2(_u10_u4_n2518 ), .ZN(_u10_u4_n2517 ) );
NAND3_X1 _u10_u4_U372  ( .A1(_u10_u4_n2515 ), .A2(_u10_u4_n2516 ), .A3(_u10_u4_n2517 ), .ZN(_u10_u4_n2512 ) );
NOR2_X1 _u10_u4_U371  ( .A1(_u10_u4_n1913 ), .A2(_u10_u4_n1940 ), .ZN(_u10_u4_n2513 ) );
NOR2_X1 _u10_u4_U370  ( .A1(_u10_u4_n2113 ), .A2(_u10_u4_n2350 ), .ZN(_u10_u4_n2514 ) );
NOR4_X1 _u10_u4_U369  ( .A1(_u10_u4_n2511 ), .A2(_u10_u4_n2512 ), .A3(_u10_u4_n2513 ), .A4(_u10_u4_n2514 ), .ZN(_u10_u4_n2389 ) );
NAND2_X1 _u10_u4_U368  ( .A1(_u10_u4_n2509 ), .A2(_u10_u4_n2510 ), .ZN(_u10_u4_n2477 ) );
NAND2_X1 _u10_u4_U367  ( .A1(_u10_u4_n2507 ), .A2(_u10_u4_n2508 ), .ZN(_u10_u4_n2504 ) );
NAND2_X1 _u10_u4_U366  ( .A1(1'b0), .A2(_u10_u4_n2506 ), .ZN(_u10_u4_n2505 ));
NAND2_X1 _u10_u4_U365  ( .A1(_u10_u4_n2504 ), .A2(_u10_u4_n2505 ), .ZN(_u10_u4_n2503 ) );
NAND2_X1 _u10_u4_U364  ( .A1(_u10_u4_n2502 ), .A2(_u10_u4_n2503 ), .ZN(_u10_u4_n2478 ) );
NAND2_X1 _u10_u4_U363  ( .A1(_u10_u4_n2501 ), .A2(_u10_u4_n2446 ), .ZN(_u10_u4_n2497 ) );
INV_X1 _u10_u4_U362  ( .A(_u10_u4_n2500 ), .ZN(_u10_u4_n2499 ) );
NAND3_X1 _u10_u4_U361  ( .A1(_u10_u4_n2497 ), .A2(_u10_u4_n2498 ), .A3(_u10_u4_n2499 ), .ZN(_u10_u4_n2496 ) );
NAND2_X1 _u10_u4_U360  ( .A1(_u10_u4_n2445 ), .A2(_u10_u4_n2496 ), .ZN(_u10_u4_n2479 ) );
NOR2_X1 _u10_u4_U359  ( .A1(_u10_u4_n2429 ), .A2(_u10_u4_n2495 ), .ZN(_u10_u4_n2491 ) );
INV_X1 _u10_u4_U358  ( .A(_u10_u4_n2191 ), .ZN(_u10_u4_n2494 ) );
NOR2_X1 _u10_u4_U357  ( .A1(_u10_u4_n2493 ), .A2(_u10_u4_n2494 ), .ZN(_u10_u4_n2492 ) );
NOR2_X1 _u10_u4_U356  ( .A1(_u10_u4_n2491 ), .A2(_u10_u4_n2492 ), .ZN(_u10_u4_n2489 ) );
NOR2_X1 _u10_u4_U355  ( .A1(_u10_u4_n2489 ), .A2(_u10_u4_n2490 ), .ZN(_u10_u4_n2481 ) );
NAND2_X1 _u10_u4_U354  ( .A1(_u10_u4_n2253 ), .A2(_u10_u4_n1859 ), .ZN(_u10_u4_n2398 ) );
NOR2_X1 _u10_u4_U353  ( .A1(_u10_u4_n2488 ), .A2(_u10_u4_n2398 ), .ZN(_u10_u4_n2487 ) );
NOR2_X1 _u10_u4_U352  ( .A1(_u10_u4_n2220 ), .A2(_u10_u4_n2487 ), .ZN(_u10_u4_n2482 ) );
AND2_X1 _u10_u4_U351  ( .A1(_u10_u4_n2350 ), .A2(_u10_u4_n2486 ), .ZN(_u10_u4_n2484 ) );
NOR2_X1 _u10_u4_U350  ( .A1(_u10_u4_n2484 ), .A2(_u10_u4_n2485 ), .ZN(_u10_u4_n2483 ) );
NOR3_X1 _u10_u4_U349  ( .A1(_u10_u4_n2481 ), .A2(_u10_u4_n2482 ), .A3(_u10_u4_n2483 ), .ZN(_u10_u4_n2480 ) );
NAND4_X1 _u10_u4_U348  ( .A1(_u10_u4_n2477 ), .A2(_u10_u4_n2478 ), .A3(_u10_u4_n2479 ), .A4(_u10_u4_n2480 ), .ZN(_u10_u4_n2447 ) );
NAND2_X1 _u10_u4_U347  ( .A1(_u10_u4_n2476 ), .A2(_u10_u4_n1936 ), .ZN(_u10_u4_n2472 ) );
NAND2_X1 _u10_u4_U346  ( .A1(_u10_u4_n2427 ), .A2(_u10_u4_n2278 ), .ZN(_u10_u4_n2473 ) );
NAND4_X1 _u10_u4_U345  ( .A1(_u10_u4_n2472 ), .A2(_u10_u4_n2473 ), .A3(_u10_u4_n2474 ), .A4(_u10_u4_n2475 ), .ZN(_u10_u4_n2471 ) );
NAND2_X1 _u10_u4_U344  ( .A1(_u10_u4_n2470 ), .A2(_u10_u4_n2471 ), .ZN(_u10_u4_n2457 ) );
NAND2_X1 _u10_u4_U343  ( .A1(_u10_u4_n2409 ), .A2(_u10_u4_n2469 ), .ZN(_u10_u4_n2468 ) );
NAND2_X1 _u10_u4_U342  ( .A1(_u10_u4_n2467 ), .A2(_u10_u4_n2468 ), .ZN(_u10_u4_n2463 ) );
NAND2_X1 _u10_u4_U341  ( .A1(_u10_u4_n1844 ), .A2(_u10_u4_n2466 ), .ZN(_u10_u4_n2465 ) );
NAND3_X1 _u10_u4_U340  ( .A1(_u10_u4_n2463 ), .A2(_u10_u4_n2464 ), .A3(_u10_u4_n2465 ), .ZN(_u10_u4_n2462 ) );
NAND2_X1 _u10_u4_U339  ( .A1(_u10_u4_n2461 ), .A2(_u10_u4_n2462 ), .ZN(_u10_u4_n2458 ) );
NAND2_X1 _u10_u4_U338  ( .A1(_u10_u4_n2460 ), .A2(_u10_u4_n2251 ), .ZN(_u10_u4_n2459 ) );
NAND3_X1 _u10_u4_U337  ( .A1(_u10_u4_n2457 ), .A2(_u10_u4_n2458 ), .A3(_u10_u4_n2459 ), .ZN(_u10_u4_n2448 ) );
NOR2_X1 _u10_u4_U336  ( .A1(_u10_u4_n2455 ), .A2(_u10_u4_n2456 ), .ZN(_u10_u4_n2449 ) );
NAND2_X1 _u10_u4_U335  ( .A1(_u10_u4_n2454 ), .A2(_u10_u4_n2438 ), .ZN(_u10_u4_n2452 ) );
NOR4_X1 _u10_u4_U334  ( .A1(_u10_u4_n2452 ), .A2(_u10_u4_n2453 ), .A3(_u10_u4_n2443 ), .A4(_u10_u4_n2143 ), .ZN(_u10_u4_n2451 ) );
NOR2_X1 _u10_u4_U333  ( .A1(_u10_u4_n2451 ), .A2(_u10_u4_n2356 ), .ZN(_u10_u4_n2450 ) );
NOR4_X1 _u10_u4_U332  ( .A1(_u10_u4_n2447 ), .A2(_u10_u4_n2448 ), .A3(_u10_u4_n2449 ), .A4(_u10_u4_n2450 ), .ZN(_u10_u4_n2390 ) );
NAND2_X1 _u10_u4_U331  ( .A1(_u10_u4_n2445 ), .A2(_u10_u4_n2446 ), .ZN(_u10_u4_n2155 ) );
INV_X1 _u10_u4_U330  ( .A(_u10_u4_n2155 ), .ZN(_u10_u4_n1892 ) );
INV_X1 _u10_u4_U329  ( .A(_u10_u4_n2444 ), .ZN(_u10_u4_n2088 ) );
NAND2_X1 _u10_u4_U328  ( .A1(_u10_u4_n1892 ), .A2(_u10_u4_n2088 ), .ZN(_u10_u4_n2337 ) );
NOR3_X1 _u10_u4_U327  ( .A1(_u10_u4_n2441 ), .A2(_u10_u4_n2442 ), .A3(_u10_u4_n2443 ), .ZN(_u10_u4_n2440 ) );
NAND4_X1 _u10_u4_U326  ( .A1(_u10_u4_n2193 ), .A2(_u10_u4_n2355 ), .A3(_u10_u4_n2439 ), .A4(_u10_u4_n2440 ), .ZN(_u10_u4_n2434 ) );
NAND3_X1 _u10_u4_U325  ( .A1(_u10_u4_n2437 ), .A2(_u10_u4_n2438 ), .A3(_u10_u4_n2059 ), .ZN(_u10_u4_n2435 ) );
NOR4_X1 _u10_u4_U324  ( .A1(_u10_u4_n2434 ), .A2(_u10_u4_n2435 ), .A3(_u10_u4_n1837 ), .A4(_u10_u4_n2436 ), .ZN(_u10_u4_n2433 ) );
NOR2_X1 _u10_u4_U323  ( .A1(_u10_u4_n2433 ), .A2(_u10_u4_n1836 ), .ZN(_u10_u4_n2415 ) );
INV_X1 _u10_u4_U322  ( .A(_u10_u4_n2432 ), .ZN(_u10_u4_n2178 ) );
NOR2_X1 _u10_u4_U321  ( .A1(_u10_u4_n1960 ), .A2(_u10_u4_n2431 ), .ZN(_u10_u4_n2430 ) );
NOR4_X1 _u10_u4_U320  ( .A1(_u10_u4_n2178 ), .A2(_u10_u4_n2429 ), .A3(_u10_u4_n2430 ), .A4(_u10_u4_n2179 ), .ZN(_u10_u4_n2416 ) );
NOR2_X1 _u10_u4_U319  ( .A1(_u10_u4_n2427 ), .A2(_u10_u4_n2428 ), .ZN(_u10_u4_n2426 ) );
NAND4_X1 _u10_u4_U318  ( .A1(_u10_u4_n2286 ), .A2(_u10_u4_n1969 ), .A3(_u10_u4_n2282 ), .A4(_u10_u4_n2426 ), .ZN(_u10_u4_n2425 ) );
NAND2_X1 _u10_u4_U317  ( .A1(_u10_u4_n2031 ), .A2(_u10_u4_n2425 ), .ZN(_u10_u4_n2422 ) );
NAND3_X1 _u10_u4_U316  ( .A1(_u10_u4_n2422 ), .A2(_u10_u4_n2423 ), .A3(_u10_u4_n2424 ), .ZN(_u10_u4_n2419 ) );
NOR4_X1 _u10_u4_U315  ( .A1(_u10_u4_n2419 ), .A2(_u10_u4_n1978 ), .A3(_u10_u4_n2420 ), .A4(_u10_u4_n2421 ), .ZN(_u10_u4_n2418 ) );
NOR2_X1 _u10_u4_U314  ( .A1(_u10_u4_n2418 ), .A2(_u10_u4_n2359 ), .ZN(_u10_u4_n2417 ) );
NOR3_X1 _u10_u4_U313  ( .A1(_u10_u4_n2415 ), .A2(_u10_u4_n2416 ), .A3(_u10_u4_n2417 ), .ZN(_u10_u4_n2414 ) );
NAND4_X1 _u10_u4_U312  ( .A1(_u10_u4_n2337 ), .A2(_u10_u4_n2412 ), .A3(_u10_u4_n2413 ), .A4(_u10_u4_n2414 ), .ZN(_u10_u4_n2392 ) );
NAND2_X1 _u10_u4_U311  ( .A1(_u10_u4_n2411 ), .A2(_u10_u4_n1936 ), .ZN(_u10_u4_n2410 ) );
NAND2_X1 _u10_u4_U310  ( .A1(_u10_u4_n2409 ), .A2(_u10_u4_n2410 ), .ZN(_u10_u4_n2408 ) );
NAND3_X1 _u10_u4_U309  ( .A1(_u10_u4_n2408 ), .A2(_u10_u4_n2305 ), .A3(_u10_u4_n1894 ), .ZN(_u10_u4_n2402 ) );
NAND3_X1 _u10_u4_U308  ( .A1(_u10_u4_n2329 ), .A2(_u10_u4_n2407 ), .A3(_u10_u4_n2255 ), .ZN(_u10_u4_n2403 ) );
NAND3_X1 _u10_u4_U307  ( .A1(_u10_u4_n1924 ), .A2(_u10_u4_n2405 ), .A3(_u10_u4_n2406 ), .ZN(_u10_u4_n2404 ) );
NAND3_X1 _u10_u4_U306  ( .A1(_u10_u4_n2402 ), .A2(_u10_u4_n2403 ), .A3(_u10_u4_n2404 ), .ZN(_u10_u4_n2393 ) );
INV_X1 _u10_u4_U305  ( .A(_u10_u4_n1932 ), .ZN(_u10_u4_n2399 ) );
NOR2_X1 _u10_u4_U304  ( .A1(_u10_u4_n2401 ), .A2(_u10_u4_n2161 ), .ZN(_u10_u4_n2400 ) );
NOR2_X1 _u10_u4_U303  ( .A1(_u10_u4_n2399 ), .A2(_u10_u4_n2400 ), .ZN(_u10_u4_n2394 ) );
NOR2_X1 _u10_u4_U302  ( .A1(_u10_u4_n2110 ), .A2(_u10_u4_n2398 ), .ZN(_u10_u4_n2397 ) );
NOR2_X1 _u10_u4_U301  ( .A1(_u10_u4_n2396 ), .A2(_u10_u4_n2397 ), .ZN(_u10_u4_n2395 ) );
NOR4_X1 _u10_u4_U300  ( .A1(_u10_u4_n2392 ), .A2(_u10_u4_n2393 ), .A3(_u10_u4_n2394 ), .A4(_u10_u4_n2395 ), .ZN(_u10_u4_n2391 ) );
NAND4_X1 _u10_u4_U299  ( .A1(_u10_u4_n2388 ), .A2(_u10_u4_n2389 ), .A3(_u10_u4_n2390 ), .A4(_u10_u4_n2391 ), .ZN(_u10_u4_n2387 ) );
MUX2_X1 _u10_u4_U298  ( .A(_u10_u4_n2387 ), .B(_u10_SYNOPSYS_UNCONNECTED_15 ), .S(_u10_u4_n1819 ), .Z(_u10_u4_n1810 ) );
NAND2_X1 _u10_u4_U297  ( .A1(_u10_u4_n2386 ), .A2(_u10_u4_n2007 ), .ZN(_u10_u4_n2369 ) );
AND2_X1 _u10_u4_U296  ( .A1(1'b0), .A2(_u10_u4_n2195 ), .ZN(_u10_u4_n2308 ));
NAND2_X1 _u10_u4_U295  ( .A1(_u10_u4_n2308 ), .A2(_u10_u4_n2036 ), .ZN(_u10_u4_n2384 ) );
AND2_X1 _u10_u4_U294  ( .A1(_u10_u4_n2384 ), .A2(_u10_u4_n2385 ), .ZN(_u10_u4_n2275 ) );
AND4_X1 _u10_u4_U293  ( .A1(_u10_u4_n2275 ), .A2(_u10_u4_n2286 ), .A3(_u10_u4_n2383 ), .A4(_u10_u4_n2285 ), .ZN(_u10_u4_n2225 ) );
NAND3_X1 _u10_u4_U292  ( .A1(_u10_u4_n2195 ), .A2(_u10_u4_n2223 ), .A3(1'b0),.ZN(_u10_u4_n2021 ) );
INV_X1 _u10_u4_U291  ( .A(_u10_u4_n2021 ), .ZN(_u10_u4_n2167 ) );
NAND2_X1 _u10_u4_U290  ( .A1(_u10_u4_n2036 ), .A2(_u10_u4_n2167 ), .ZN(_u10_u4_n1970 ) );
AND3_X1 _u10_u4_U289  ( .A1(_u10_u4_n1970 ), .A2(_u10_u4_n2164 ), .A3(_u10_u4_n2382 ), .ZN(_u10_u4_n2381 ) );
NAND4_X1 _u10_u4_U288  ( .A1(_u10_u4_n2225 ), .A2(_u10_u4_n2379 ), .A3(_u10_u4_n2380 ), .A4(_u10_u4_n2381 ), .ZN(_u10_u4_n2378 ) );
NAND2_X1 _u10_u4_U287  ( .A1(_u10_u4_n1967 ), .A2(_u10_u4_n2378 ), .ZN(_u10_u4_n2370 ) );
NAND2_X1 _u10_u4_U286  ( .A1(_u10_u4_n2081 ), .A2(_u10_u4_n2377 ), .ZN(_u10_u4_n2371 ) );
NOR2_X1 _u10_u4_U285  ( .A1(_u10_u4_n2375 ), .A2(_u10_u4_n2376 ), .ZN(_u10_u4_n2373 ) );
NOR2_X1 _u10_u4_U284  ( .A1(_u10_u4_n2373 ), .A2(_u10_u4_n2374 ), .ZN(_u10_u4_n2372 ) );
NAND4_X1 _u10_u4_U283  ( .A1(_u10_u4_n2369 ), .A2(_u10_u4_n2370 ), .A3(_u10_u4_n2371 ), .A4(_u10_u4_n2372 ), .ZN(_u10_u4_n2309 ) );
NOR2_X1 _u10_u4_U282  ( .A1(_u10_u4_n2000 ), .A2(_u10_u4_n2368 ), .ZN(_u10_u4_n2360 ) );
NOR2_X1 _u10_u4_U281  ( .A1(_u10_u4_n2366 ), .A2(_u10_u4_n2367 ), .ZN(_u10_u4_n2361 ) );
NOR2_X1 _u10_u4_U280  ( .A1(_u10_u4_n1868 ), .A2(_u10_u4_n2365 ), .ZN(_u10_u4_n2362 ) );
NOR2_X1 _u10_u4_U279  ( .A1(_u10_u4_n2364 ), .A2(_u10_u4_n1859 ), .ZN(_u10_u4_n2363 ) );
NOR4_X1 _u10_u4_U278  ( .A1(_u10_u4_n2360 ), .A2(_u10_u4_n2361 ), .A3(_u10_u4_n2362 ), .A4(_u10_u4_n2363 ), .ZN(_u10_u4_n2316 ) );
NOR2_X1 _u10_u4_U277  ( .A1(_u10_u4_n2359 ), .A2(_u10_u4_n1970 ), .ZN(_u10_u4_n2351 ) );
NOR2_X1 _u10_u4_U276  ( .A1(_u10_u4_n2358 ), .A2(_u10_u4_n1840 ), .ZN(_u10_u4_n2352 ) );
NOR2_X1 _u10_u4_U275  ( .A1(_u10_u4_n2356 ), .A2(_u10_u4_n2357 ), .ZN(_u10_u4_n2353 ) );
NOR2_X1 _u10_u4_U274  ( .A1(_u10_u4_n1836 ), .A2(_u10_u4_n2355 ), .ZN(_u10_u4_n2354 ) );
NOR4_X1 _u10_u4_U273  ( .A1(_u10_u4_n2351 ), .A2(_u10_u4_n2352 ), .A3(_u10_u4_n2353 ), .A4(_u10_u4_n2354 ), .ZN(_u10_u4_n2317 ) );
NOR2_X1 _u10_u4_U272  ( .A1(_u10_u4_n1873 ), .A2(_u10_u4_n2101 ), .ZN(_u10_u4_n2349 ) );
NOR2_X1 _u10_u4_U271  ( .A1(_u10_u4_n2349 ), .A2(_u10_u4_n2350 ), .ZN(_u10_u4_n2338 ) );
NOR2_X1 _u10_u4_U270  ( .A1(_u10_u4_n2347 ), .A2(_u10_u4_n2348 ), .ZN(_u10_u4_n2345 ) );
NOR2_X1 _u10_u4_U269  ( .A1(_u10_u4_n2345 ), .A2(_u10_u4_n2346 ), .ZN(_u10_u4_n2339 ) );
NOR2_X1 _u10_u4_U268  ( .A1(_u10_u4_n2344 ), .A2(_u10_u4_n2142 ), .ZN(_u10_u4_n2340 ) );
NOR2_X1 _u10_u4_U267  ( .A1(_u10_u4_n2342 ), .A2(_u10_u4_n2343 ), .ZN(_u10_u4_n2341 ) );
NOR4_X1 _u10_u4_U266  ( .A1(_u10_u4_n2338 ), .A2(_u10_u4_n2339 ), .A3(_u10_u4_n2340 ), .A4(_u10_u4_n2341 ), .ZN(_u10_u4_n2318 ) );
INV_X1 _u10_u4_U265  ( .A(_u10_u4_n2337 ), .ZN(_u10_u4_n2320 ) );
NOR2_X1 _u10_u4_U264  ( .A1(_u10_u4_n1970 ), .A2(1'b0), .ZN(_u10_u4_n2027 ));
INV_X1 _u10_u4_U263  ( .A(_u10_u4_n2027 ), .ZN(_u10_u4_n2331 ) );
NOR2_X1 _u10_u4_U262  ( .A1(_u10_u4_n2174 ), .A2(_u10_u4_n2216 ), .ZN(_u10_u4_n2333 ) );
AND2_X1 _u10_u4_U261  ( .A1(_u10_u4_n1928 ), .A2(_u10_u4_n2336 ), .ZN(_u10_u4_n2334 ) );
NOR4_X1 _u10_u4_U260  ( .A1(_u10_u4_n1937 ), .A2(_u10_u4_n2333 ), .A3(_u10_u4_n2334 ), .A4(_u10_u4_n2335 ), .ZN(_u10_u4_n2332 ) );
NOR3_X1 _u10_u4_U259  ( .A1(_u10_u4_n2331 ), .A2(_u10_u4_n2332 ), .A3(_u10_u4_n1915 ), .ZN(_u10_u4_n2321 ) );
NOR3_X1 _u10_u4_U258  ( .A1(_u10_u4_n2291 ), .A2(_u10_u4_n2330 ), .A3(_u10_u4_n2021 ), .ZN(_u10_u4_n2322 ) );
NOR2_X1 _u10_u4_U257  ( .A1(_u10_u4_n2329 ), .A2(_u10_u4_n2169 ), .ZN(_u10_u4_n2324 ) );
NOR2_X1 _u10_u4_U256  ( .A1(1'b0), .A2(_u10_u4_n2328 ), .ZN(_u10_u4_n2327 ));
NOR2_X1 _u10_u4_U255  ( .A1(_u10_u4_n2326 ), .A2(_u10_u4_n2327 ), .ZN(_u10_u4_n2325 ) );
NOR3_X1 _u10_u4_U254  ( .A1(_u10_u4_n2324 ), .A2(1'b0), .A3(_u10_u4_n2325 ),.ZN(_u10_u4_n2323 ) );
NOR4_X1 _u10_u4_U253  ( .A1(_u10_u4_n2320 ), .A2(_u10_u4_n2321 ), .A3(_u10_u4_n2322 ), .A4(_u10_u4_n2323 ), .ZN(_u10_u4_n2319 ) );
AND4_X1 _u10_u4_U252  ( .A1(_u10_u4_n2316 ), .A2(_u10_u4_n2317 ), .A3(_u10_u4_n2318 ), .A4(_u10_u4_n2319 ), .ZN(_u10_u4_n1991 ) );
INV_X1 _u10_u4_U251  ( .A(_u10_u4_n2315 ), .ZN(_u10_u4_n2313 ) );
NAND3_X1 _u10_u4_U250  ( .A1(_u10_u4_n1991 ), .A2(_u10_u4_n2313 ), .A3(_u10_u4_n2314 ), .ZN(_u10_u4_n2310 ) );
NOR4_X1 _u10_u4_U249  ( .A1(_u10_u4_n2309 ), .A2(_u10_u4_n2310 ), .A3(_u10_u4_n2311 ), .A4(_u10_u4_n2312 ), .ZN(_u10_u4_n2117 ) );
NAND3_X1 _u10_u4_U248  ( .A1(_u10_u4_n2108 ), .A2(_u10_u4_n2107 ), .A3(_u10_u4_n2308 ), .ZN(_u10_u4_n2217 ) );
NOR3_X1 _u10_u4_U247  ( .A1(_u10_u4_n2306 ), .A2(_u10_u4_n2307 ), .A3(_u10_u4_n2027 ), .ZN(_u10_u4_n2277 ) );
NAND3_X1 _u10_u4_U246  ( .A1(_u10_u4_n2217 ), .A2(_u10_u4_n2305 ), .A3(_u10_u4_n2277 ), .ZN(_u10_u4_n2157 ) );
NAND2_X1 _u10_u4_U245  ( .A1(_u10_u4_n2089 ), .A2(_u10_u4_n2157 ), .ZN(_u10_u4_n2296 ) );
INV_X1 _u10_u4_U244  ( .A(_u10_u4_n2304 ), .ZN(_u10_u4_n2297 ) );
NOR2_X1 _u10_u4_U243  ( .A1(_u10_u4_n2302 ), .A2(_u10_u4_n2303 ), .ZN(_u10_u4_n2299 ) );
NOR3_X1 _u10_u4_U242  ( .A1(_u10_u4_n2299 ), .A2(_u10_u4_n2300 ), .A3(_u10_u4_n2301 ), .ZN(_u10_u4_n2298 ) );
NAND4_X1 _u10_u4_U241  ( .A1(_u10_u4_n2295 ), .A2(_u10_u4_n2296 ), .A3(_u10_u4_n2297 ), .A4(_u10_u4_n2298 ), .ZN(_u10_u4_n2294 ) );
NAND2_X1 _u10_u4_U240  ( .A1(_u10_u4_n2293 ), .A2(_u10_u4_n2294 ), .ZN(_u10_u4_n2257 ) );
NAND2_X1 _u10_u4_U239  ( .A1(_u10_u4_n2165 ), .A2(_u10_u4_n2166 ), .ZN(_u10_u4_n2288 ) );
NAND2_X1 _u10_u4_U238  ( .A1(_u10_u4_n2078 ), .A2(_u10_u4_n2279 ), .ZN(_u10_u4_n2292 ) );
NAND2_X1 _u10_u4_U237  ( .A1(_u10_u4_n2291 ), .A2(_u10_u4_n2292 ), .ZN(_u10_u4_n2290 ) );
NAND2_X1 _u10_u4_U236  ( .A1(_u10_u4_n2059 ), .A2(_u10_u4_n2290 ), .ZN(_u10_u4_n2289 ) );
NAND2_X1 _u10_u4_U235  ( .A1(_u10_u4_n2288 ), .A2(_u10_u4_n2289 ), .ZN(_u10_u4_n2201 ) );
NAND2_X1 _u10_u4_U234  ( .A1(1'b0), .A2(_u10_u4_n2201 ), .ZN(_u10_u4_n2258 ));
INV_X1 _u10_u4_U233  ( .A(_u10_u4_n2287 ), .ZN(_u10_u4_n2283 ) );
AND4_X1 _u10_u4_U232  ( .A1(_u10_u4_n2285 ), .A2(_u10_u4_n2226 ), .A3(_u10_u4_n1970 ), .A4(_u10_u4_n2286 ), .ZN(_u10_u4_n2284 ) );
NAND4_X1 _u10_u4_U231  ( .A1(_u10_u4_n2281 ), .A2(_u10_u4_n2282 ), .A3(_u10_u4_n2283 ), .A4(_u10_u4_n2284 ), .ZN(_u10_u4_n2280 ) );
NAND2_X1 _u10_u4_U230  ( .A1(_u10_u4_n2279 ), .A2(_u10_u4_n2280 ), .ZN(_u10_u4_n2259 ) );
NAND4_X1 _u10_u4_U229  ( .A1(_u10_u4_n2275 ), .A2(_u10_u4_n2276 ), .A3(_u10_u4_n2277 ), .A4(_u10_u4_n2278 ), .ZN(_u10_u4_n2271 ) );
NAND2_X1 _u10_u4_U228  ( .A1(_u10_u4_n1933 ), .A2(_u10_u4_n2164 ), .ZN(_u10_u4_n2272 ) );
NOR2_X1 _u10_u4_U227  ( .A1(_u10_u4_n2274 ), .A2(_u10_u4_n2130 ), .ZN(_u10_u4_n2273 ) );
NOR4_X1 _u10_u4_U226  ( .A1(_u10_u4_n2271 ), .A2(_u10_u4_n2272 ), .A3(_u10_u4_n1978 ), .A4(_u10_u4_n2273 ), .ZN(_u10_u4_n2270 ) );
NOR2_X1 _u10_u4_U225  ( .A1(_u10_u4_n2270 ), .A2(_u10_u4_n2025 ), .ZN(_u10_u4_n2261 ) );
NAND3_X1 _u10_u4_U224  ( .A1(_u10_u4_n1933 ), .A2(_u10_u4_n1936 ), .A3(_u10_u4_n2269 ), .ZN(_u10_u4_n2268 ) );
NOR3_X1 _u10_u4_U223  ( .A1(_u10_u4_n2268 ), .A2(_u10_u4_n1844 ), .A3(_u10_u4_n2157 ), .ZN(_u10_u4_n2267 ) );
NOR2_X1 _u10_u4_U222  ( .A1(1'b0), .A2(_u10_u4_n2267 ), .ZN(_u10_u4_n2265 ));
NOR3_X1 _u10_u4_U221  ( .A1(_u10_u4_n2264 ), .A2(_u10_u4_n2265 ), .A3(_u10_u4_n2266 ), .ZN(_u10_u4_n2263 ) );
NOR2_X1 _u10_u4_U220  ( .A1(_u10_u4_n2263 ), .A2(_u10_u4_n1843 ), .ZN(_u10_u4_n2262 ) );
NOR2_X1 _u10_u4_U219  ( .A1(_u10_u4_n2261 ), .A2(_u10_u4_n2262 ), .ZN(_u10_u4_n2260 ) );
NAND4_X1 _u10_u4_U218  ( .A1(_u10_u4_n2257 ), .A2(_u10_u4_n2258 ), .A3(_u10_u4_n2259 ), .A4(_u10_u4_n2260 ), .ZN(_u10_u4_n2230 ) );
INV_X1 _u10_u4_U217  ( .A(_u10_u4_n2217 ), .ZN(_u10_u4_n2242 ) );
NAND2_X1 _u10_u4_U216  ( .A1(_u10_u4_n2168 ), .A2(_u10_u4_n2169 ), .ZN(_u10_u4_n2244 ) );
NAND2_X1 _u10_u4_U215  ( .A1(_u10_u4_n2255 ), .A2(_u10_u4_n2256 ), .ZN(_u10_u4_n2245 ) );
NAND2_X1 _u10_u4_U214  ( .A1(_u10_u4_n2253 ), .A2(_u10_u4_n2254 ), .ZN(_u10_u4_n2252 ) );
NAND2_X1 _u10_u4_U213  ( .A1(_u10_u4_n2251 ), .A2(_u10_u4_n2252 ), .ZN(_u10_u4_n2246 ) );
NAND2_X1 _u10_u4_U212  ( .A1(_u10_u4_n2152 ), .A2(_u10_u4_n1928 ), .ZN(_u10_u4_n2250 ) );
NAND2_X1 _u10_u4_U211  ( .A1(_u10_u4_n2249 ), .A2(_u10_u4_n2250 ), .ZN(_u10_u4_n2248 ) );
NAND2_X1 _u10_u4_U210  ( .A1(_u10_u4_n2105 ), .A2(_u10_u4_n2248 ), .ZN(_u10_u4_n2247 ) );
NAND4_X1 _u10_u4_U209  ( .A1(_u10_u4_n2244 ), .A2(_u10_u4_n2245 ), .A3(_u10_u4_n2246 ), .A4(_u10_u4_n2247 ), .ZN(_u10_u4_n2243 ) );
NAND2_X1 _u10_u4_U208  ( .A1(_u10_u4_n2242 ), .A2(_u10_u4_n2243 ), .ZN(_u10_u4_n2237 ) );
NAND2_X1 _u10_u4_U207  ( .A1(1'b0), .A2(_u10_u4_n2241 ), .ZN(_u10_u4_n2238 ));
NAND2_X1 _u10_u4_U206  ( .A1(_u10_u4_n2214 ), .A2(_u10_u4_n2240 ), .ZN(_u10_u4_n2239 ) );
NAND3_X1 _u10_u4_U205  ( .A1(_u10_u4_n2237 ), .A2(_u10_u4_n2238 ), .A3(_u10_u4_n2239 ), .ZN(_u10_u4_n2231 ) );
AND2_X1 _u10_u4_U204  ( .A1(_u10_u4_n2200 ), .A2(_u10_u4_n2236 ), .ZN(_u10_u4_n2232 ) );
NOR2_X1 _u10_u4_U203  ( .A1(_u10_u4_n2234 ), .A2(_u10_u4_n2235 ), .ZN(_u10_u4_n2233 ) );
NOR4_X1 _u10_u4_U202  ( .A1(_u10_u4_n2230 ), .A2(_u10_u4_n2231 ), .A3(_u10_u4_n2232 ), .A4(_u10_u4_n2233 ), .ZN(_u10_u4_n2118 ) );
NAND2_X1 _u10_u4_U201  ( .A1(_u10_u4_n2214 ), .A2(_u10_u4_n2049 ), .ZN(_u10_u4_n2229 ) );
NAND2_X1 _u10_u4_U200  ( .A1(_u10_u4_n2228 ), .A2(_u10_u4_n2229 ), .ZN(_u10_u4_n2227 ) );
NAND2_X1 _u10_u4_U199  ( .A1(_u10_u4_n2043 ), .A2(_u10_u4_n2227 ), .ZN(_u10_u4_n2204 ) );
NAND2_X1 _u10_u4_U198  ( .A1(_u10_u4_n2225 ), .A2(_u10_u4_n2226 ), .ZN(_u10_u4_n2224 ) );
NAND2_X1 _u10_u4_U197  ( .A1(_u10_u4_n1899 ), .A2(_u10_u4_n2224 ), .ZN(_u10_u4_n2205 ) );
NAND2_X1 _u10_u4_U196  ( .A1(_u10_u4_n2222 ), .A2(_u10_u4_n2223 ), .ZN(_u10_u4_n1870 ) );
NAND4_X1 _u10_u4_U195  ( .A1(_u10_u4_n2220 ), .A2(_u10_u4_n2131 ), .A3(_u10_u4_n2221 ), .A4(_u10_u4_n1870 ), .ZN(_u10_u4_n2219 ) );
NAND2_X1 _u10_u4_U194  ( .A1(_u10_u4_n2218 ), .A2(_u10_u4_n2219 ), .ZN(_u10_u4_n2206 ) );
NOR2_X1 _u10_u4_U193  ( .A1(_u10_u4_n1925 ), .A2(_u10_u4_n2217 ), .ZN(_u10_u4_n2215 ) );
NOR4_X1 _u10_u4_U192  ( .A1(_u10_u4_n2213 ), .A2(_u10_u4_n2214 ), .A3(_u10_u4_n2215 ), .A4(_u10_u4_n2216 ), .ZN(_u10_u4_n2211 ) );
NOR2_X1 _u10_u4_U191  ( .A1(_u10_u4_n2211 ), .A2(_u10_u4_n2212 ), .ZN(_u10_u4_n2208 ) );
NOR2_X1 _u10_u4_U190  ( .A1(_u10_u4_n1888 ), .A2(_u10_u4_n2210 ), .ZN(_u10_u4_n2209 ) );
NOR2_X1 _u10_u4_U189  ( .A1(_u10_u4_n2208 ), .A2(_u10_u4_n2209 ), .ZN(_u10_u4_n2207 ) );
NAND4_X1 _u10_u4_U188  ( .A1(_u10_u4_n2204 ), .A2(_u10_u4_n2205 ), .A3(_u10_u4_n2206 ), .A4(_u10_u4_n2207 ), .ZN(_u10_u4_n2170 ) );
OR2_X1 _u10_u4_U187  ( .A1(_u10_u4_n2202 ), .A2(_u10_u4_n2203 ), .ZN(_u10_u4_n2197 ) );
NAND2_X1 _u10_u4_U186  ( .A1(1'b0), .A2(_u10_u4_n2201 ), .ZN(_u10_u4_n2198 ));
NAND2_X1 _u10_u4_U185  ( .A1(_u10_u4_n2063 ), .A2(_u10_u4_n2200 ), .ZN(_u10_u4_n2199 ) );
NAND3_X1 _u10_u4_U184  ( .A1(_u10_u4_n2197 ), .A2(_u10_u4_n2198 ), .A3(_u10_u4_n2199 ), .ZN(_u10_u4_n2196 ) );
NAND2_X1 _u10_u4_U183  ( .A1(_u10_u4_n2195 ), .A2(_u10_u4_n2196 ), .ZN(_u10_u4_n2180 ) );
NAND2_X1 _u10_u4_U182  ( .A1(_u10_u4_n2195 ), .A2(_u10_u4_n1918 ), .ZN(_u10_u4_n2192 ) );
NAND4_X1 _u10_u4_U181  ( .A1(_u10_u4_n2192 ), .A2(_u10_u4_n2021 ), .A3(_u10_u4_n2193 ), .A4(_u10_u4_n2194 ), .ZN(_u10_u4_n2188 ) );
NAND2_X1 _u10_u4_U180  ( .A1(_u10_u4_n2188 ), .A2(_u10_u4_n2191 ), .ZN(_u10_u4_n2181 ) );
NAND2_X1 _u10_u4_U179  ( .A1(1'b0), .A2(_u10_u4_n2190 ), .ZN(_u10_u4_n2185 ));
NAND2_X1 _u10_u4_U178  ( .A1(_u10_u4_n2189 ), .A2(_u10_SYNOPSYS_UNCONNECTED_16 ), .ZN(_u10_u4_n2186 ) );
INV_X1 _u10_u4_U177  ( .A(_u10_u4_n2188 ), .ZN(_u10_u4_n2187 ) );
NAND3_X1 _u10_u4_U176  ( .A1(_u10_u4_n2185 ), .A2(_u10_u4_n2186 ), .A3(_u10_u4_n2187 ), .ZN(_u10_u4_n2184 ) );
NAND2_X1 _u10_u4_U175  ( .A1(_u10_u4_n2183 ), .A2(_u10_u4_n2184 ), .ZN(_u10_u4_n2182 ) );
NAND3_X1 _u10_u4_U174  ( .A1(_u10_u4_n2180 ), .A2(_u10_u4_n2181 ), .A3(_u10_u4_n2182 ), .ZN(_u10_u4_n2171 ) );
INV_X1 _u10_u4_U173  ( .A(_u10_u4_n2179 ), .ZN(_u10_u4_n1963 ) );
NOR2_X1 _u10_u4_U172  ( .A1(_u10_u4_n1963 ), .A2(_u10_u4_n2178 ), .ZN(_u10_u4_n2172 ) );
INV_X1 _u10_u4_U171  ( .A(_u10_u4_n2177 ), .ZN(_u10_u4_n2176 ) );
NOR3_X1 _u10_u4_U170  ( .A1(_u10_u4_n2174 ), .A2(_u10_u4_n2175 ), .A3(_u10_u4_n2176 ), .ZN(_u10_u4_n2173 ) );
NOR4_X1 _u10_u4_U169  ( .A1(_u10_u4_n2170 ), .A2(_u10_u4_n2171 ), .A3(_u10_u4_n2172 ), .A4(_u10_u4_n2173 ), .ZN(_u10_u4_n2119 ) );
NAND3_X1 _u10_u4_U168  ( .A1(_u10_u4_n2168 ), .A2(_u10_u4_n2169 ), .A3(1'b0),.ZN(_u10_u4_n2148 ) );
NAND3_X1 _u10_u4_U167  ( .A1(_u10_u4_n2165 ), .A2(_u10_u4_n2166 ), .A3(_u10_u4_n2167 ), .ZN(_u10_u4_n2149 ) );
NAND4_X1 _u10_u4_U166  ( .A1(_u10_u4_n2162 ), .A2(_u10_u4_n1933 ), .A3(_u10_u4_n2163 ), .A4(_u10_u4_n2164 ), .ZN(_u10_u4_n2160 ) );
NOR4_X1 _u10_u4_U165  ( .A1(_u10_u4_n2160 ), .A2(_u10_u4_n2157 ), .A3(_u10_u4_n1844 ), .A4(_u10_u4_n2161 ), .ZN(_u10_u4_n2158 ) );
NOR2_X1 _u10_u4_U164  ( .A1(_u10_u4_n2158 ), .A2(_u10_u4_n2159 ), .ZN(_u10_u4_n2153 ) );
INV_X1 _u10_u4_U163  ( .A(_u10_u4_n2157 ), .ZN(_u10_u4_n2129 ) );
NOR3_X1 _u10_u4_U162  ( .A1(_u10_u4_n2155 ), .A2(_u10_u4_n2129 ), .A3(_u10_u4_n2156 ), .ZN(_u10_u4_n2154 ) );
NOR2_X1 _u10_u4_U161  ( .A1(_u10_u4_n2153 ), .A2(_u10_u4_n2154 ), .ZN(_u10_u4_n2150 ) );
NAND3_X1 _u10_u4_U160  ( .A1(1'b0), .A2(_u10_u4_n1928 ), .A3(_u10_u4_n2152 ),.ZN(_u10_u4_n2151 ) );
NAND4_X1 _u10_u4_U159  ( .A1(_u10_u4_n2148 ), .A2(_u10_u4_n2149 ), .A3(_u10_u4_n2150 ), .A4(_u10_u4_n2151 ), .ZN(_u10_u4_n2121 ) );
NAND2_X1 _u10_u4_U158  ( .A1(_u10_u4_n2107 ), .A2(_u10_u4_n2147 ), .ZN(_u10_u4_n2146 ) );
NAND2_X1 _u10_u4_U157  ( .A1(_u10_u4_n2145 ), .A2(_u10_u4_n2146 ), .ZN(_u10_u4_n2144 ) );
NAND2_X1 _u10_u4_U156  ( .A1(_u10_u4_n2143 ), .A2(_u10_u4_n2144 ), .ZN(_u10_u4_n2134 ) );
NAND2_X1 _u10_u4_U155  ( .A1(_u10_u4_n2141 ), .A2(_u10_u4_n2142 ), .ZN(_u10_u4_n2140 ) );
NAND2_X1 _u10_u4_U154  ( .A1(_u10_u4_n2139 ), .A2(_u10_u4_n2140 ), .ZN(_u10_u4_n2135 ) );
OR2_X1 _u10_u4_U153  ( .A1(_u10_u4_n2110 ), .A2(_u10_u4_n1911 ), .ZN(_u10_u4_n2137 ) );
NAND2_X1 _u10_u4_U152  ( .A1(_u10_u4_n2137 ), .A2(_u10_u4_n2138 ), .ZN(_u10_u4_n2136 ) );
NAND3_X1 _u10_u4_U151  ( .A1(_u10_u4_n2134 ), .A2(_u10_u4_n2135 ), .A3(_u10_u4_n2136 ), .ZN(_u10_u4_n2122 ) );
NOR2_X1 _u10_u4_U150  ( .A1(_u10_u4_n2133 ), .A2(_u10_u4_n1891 ), .ZN(_u10_u4_n2132 ) );
NOR2_X1 _u10_u4_U149  ( .A1(_u10_u4_n2131 ), .A2(_u10_u4_n2132 ), .ZN(_u10_u4_n2123 ) );
NOR2_X1 _u10_u4_U148  ( .A1(_u10_u4_n2129 ), .A2(_u10_u4_n2130 ), .ZN(_u10_u4_n2127 ) );
NOR2_X1 _u10_u4_U147  ( .A1(_u10_u4_n2127 ), .A2(_u10_u4_n2128 ), .ZN(_u10_u4_n2125 ) );
NOR2_X1 _u10_u4_U146  ( .A1(_u10_u4_n2125 ), .A2(_u10_u4_n2126 ), .ZN(_u10_u4_n2124 ) );
NOR4_X1 _u10_u4_U145  ( .A1(_u10_u4_n2121 ), .A2(_u10_u4_n2122 ), .A3(_u10_u4_n2123 ), .A4(_u10_u4_n2124 ), .ZN(_u10_u4_n2120 ) );
NAND4_X1 _u10_u4_U144  ( .A1(_u10_u4_n2117 ), .A2(_u10_u4_n2118 ), .A3(_u10_u4_n2119 ), .A4(_u10_u4_n2120 ), .ZN(_u10_u4_n2116 ) );
MUX2_X1 _u10_u4_U143  ( .A(_u10_u4_n2116 ), .B(_u10_SYNOPSYS_UNCONNECTED_16 ), .S(_u10_u4_n1819 ), .Z(_u10_u4_n1811 ) );
INV_X1 _u10_u4_U142  ( .A(_u10_u4_n2115 ), .ZN(_u10_u4_n2006 ) );
NOR3_X1 _u10_u4_U141  ( .A1(_u10_u4_n2006 ), .A2(_u10_u4_n2114 ), .A3(_u10_u4_n2081 ), .ZN(_u10_u4_n1854 ) );
NAND2_X1 _u10_u4_U140  ( .A1(_u10_u4_n2112 ), .A2(_u10_u4_n2113 ), .ZN(_u10_u4_n1872 ) );
INV_X1 _u10_u4_U139  ( .A(_u10_u4_n1872 ), .ZN(_u10_u4_n1882 ) );
NAND4_X1 _u10_u4_U138  ( .A1(_u10_u4_n1854 ), .A2(_u10_u4_n1882 ), .A3(_u10_u4_n2111 ), .A4(_u10_u4_n1868 ), .ZN(_u10_u4_n2109 ) );
NAND2_X1 _u10_u4_U137  ( .A1(_u10_u4_n2109 ), .A2(_u10_u4_n2110 ), .ZN(_u10_u4_n2098 ) );
NAND2_X1 _u10_u4_U136  ( .A1(1'b0), .A2(_u10_u4_n1983 ), .ZN(_u10_u4_n2023 ));
INV_X1 _u10_u4_U135  ( .A(_u10_u4_n2023 ), .ZN(_u10_u4_n2035 ) );
NAND3_X1 _u10_u4_U134  ( .A1(_u10_u4_n2035 ), .A2(_u10_u4_n2107 ), .A3(_u10_u4_n2108 ), .ZN(_u10_u4_n1916 ) );
INV_X1 _u10_u4_U133  ( .A(_u10_u4_n1916 ), .ZN(_u10_u4_n2093 ) );
NAND3_X1 _u10_u4_U132  ( .A1(_u10_u4_n2105 ), .A2(_u10_u4_n2106 ), .A3(_u10_u4_n2093 ), .ZN(_u10_u4_n2039 ) );
NAND2_X1 _u10_u4_U131  ( .A1(_u10_u4_n2039 ), .A2(_u10_u4_n1930 ), .ZN(_u10_u4_n2104 ) );
NAND2_X1 _u10_u4_U130  ( .A1(_u10_u4_n2103 ), .A2(_u10_u4_n2104 ), .ZN(_u10_u4_n1863 ) );
OR2_X1 _u10_u4_U129  ( .A1(_u10_u4_n1863 ), .A2(_u10_u4_n2102 ), .ZN(_u10_u4_n2099 ) );
NAND2_X1 _u10_u4_U128  ( .A1(_u10_u4_n1890 ), .A2(_u10_u4_n2101 ), .ZN(_u10_u4_n2100 ) );
NAND3_X1 _u10_u4_U127  ( .A1(_u10_u4_n2098 ), .A2(_u10_u4_n2099 ), .A3(_u10_u4_n2100 ), .ZN(_u10_u4_n2066 ) );
NAND4_X1 _u10_u4_U126  ( .A1(_u10_u4_n2095 ), .A2(_u10_u4_n2096 ), .A3(_u10_u4_n1896 ), .A4(_u10_u4_n2097 ), .ZN(_u10_u4_n2086 ) );
NOR4_X1 _u10_u4_U125  ( .A1(_u10_u4_n2093 ), .A2(_u10_u4_n2027 ), .A3(_u10_u4_n2094 ), .A4(_u10_u4_n2026 ), .ZN(_u10_u4_n1952 ) );
NOR2_X1 _u10_u4_U124  ( .A1(1'b0), .A2(_u10_u4_n1952 ), .ZN(_u10_u4_n1951 ));
INV_X1 _u10_u4_U123  ( .A(_u10_u4_n1951 ), .ZN(_u10_u4_n2090 ) );
NAND4_X1 _u10_u4_U122  ( .A1(_u10_u4_n2089 ), .A2(_u10_u4_n2090 ), .A3(_u10_u4_n2091 ), .A4(_u10_u4_n2092 ), .ZN(_u10_u4_n1893 ) );
NOR4_X1 _u10_u4_U121  ( .A1(_u10_u4_n2086 ), .A2(_u10_u4_n1893 ), .A3(_u10_u4_n2087 ), .A4(_u10_u4_n2088 ), .ZN(_u10_u4_n2084 ) );
NOR2_X1 _u10_u4_U120  ( .A1(_u10_u4_n2084 ), .A2(_u10_u4_n2085 ), .ZN(_u10_u4_n2067 ) );
NOR2_X1 _u10_u4_U119  ( .A1(_u10_u4_n2083 ), .A2(_u10_u4_n1869 ), .ZN(_u10_u4_n2068 ) );
NAND2_X1 _u10_u4_U118  ( .A1(_u10_u4_n2081 ), .A2(_u10_u4_n2082 ), .ZN(_u10_u4_n2075 ) );
NAND2_X1 _u10_u4_U117  ( .A1(_u10_u4_n2035 ), .A2(_u10_u4_n2019 ), .ZN(_u10_u4_n2060 ) );
NAND2_X1 _u10_u4_U116  ( .A1(_u10_u4_n2080 ), .A2(_u10_u4_n2060 ), .ZN(_u10_u4_n2079 ) );
NAND2_X1 _u10_u4_U115  ( .A1(_u10_u4_n2078 ), .A2(_u10_u4_n2079 ), .ZN(_u10_u4_n2076 ) );
NAND4_X1 _u10_u4_U114  ( .A1(_u10_u4_n2075 ), .A2(_u10_u4_n2076 ), .A3(_u10_u4_n1970 ), .A4(_u10_u4_n2077 ), .ZN(_u10_u4_n2072 ) );
NOR4_X1 _u10_u4_U113  ( .A1(_u10_u4_n2072 ), .A2(_u10_u4_n2073 ), .A3(_u10_u4_n1975 ), .A4(_u10_u4_n2074 ), .ZN(_u10_u4_n2070 ) );
NOR2_X1 _u10_u4_U112  ( .A1(_u10_u4_n2070 ), .A2(_u10_u4_n2071 ), .ZN(_u10_u4_n2069 ) );
NOR4_X1 _u10_u4_U111  ( .A1(_u10_u4_n2066 ), .A2(_u10_u4_n2067 ), .A3(_u10_u4_n2068 ), .A4(_u10_u4_n2069 ), .ZN(_u10_u4_n1820 ) );
NAND2_X1 _u10_u4_U110  ( .A1(1'b0), .A2(_u10_u4_n1983 ), .ZN(_u10_u4_n2065 ));
NAND4_X1 _u10_u4_U109  ( .A1(_u10_u4_n2065 ), .A2(_u10_u4_n2023 ), .A3(_u10_u4_n2021 ), .A4(_u10_u4_n2052 ), .ZN(_u10_u4_n2064 ) );
NAND2_X1 _u10_u4_U108  ( .A1(_u10_u4_n2063 ), .A2(_u10_u4_n2064 ), .ZN(_u10_u4_n2040 ) );
NAND4_X1 _u10_u4_U107  ( .A1(_u10_u4_n2059 ), .A2(_u10_u4_n2060 ), .A3(_u10_u4_n2061 ), .A4(_u10_u4_n2062 ), .ZN(_u10_u4_n2058 ) );
NAND2_X1 _u10_u4_U106  ( .A1(_u10_u4_n2057 ), .A2(_u10_u4_n2058 ), .ZN(_u10_u4_n2041 ) );
NOR4_X1 _u10_u4_U105  ( .A1(1'b0), .A2(_u10_u4_n2054 ), .A3(_u10_u4_n2055 ),.A4(_u10_u4_n2056 ), .ZN(_u10_u4_n2053 ) );
NAND4_X1 _u10_u4_U104  ( .A1(_u10_u4_n2021 ), .A2(_u10_u4_n2052 ), .A3(_u10_u4_n2023 ), .A4(_u10_u4_n2053 ), .ZN(_u10_u4_n1964 ) );
INV_X1 _u10_u4_U103  ( .A(_u10_u4_n1964 ), .ZN(_u10_u4_n2045 ) );
NAND2_X1 _u10_u4_U102  ( .A1(_u10_u4_n2051 ), .A2(_u10_SYNOPSYS_UNCONNECTED_17 ), .ZN(_u10_u4_n2046 ) );
NAND2_X1 _u10_u4_U101  ( .A1(_u10_u4_n2049 ), .A2(_u10_u4_n2050 ), .ZN(_u10_u4_n2047 ) );
NAND4_X1 _u10_u4_U100  ( .A1(_u10_u4_n2045 ), .A2(_u10_u4_n2046 ), .A3(_u10_u4_n2047 ), .A4(_u10_u4_n2048 ), .ZN(_u10_u4_n2044 ) );
NAND2_X1 _u10_u4_U99  ( .A1(_u10_u4_n2043 ), .A2(_u10_u4_n2044 ), .ZN(_u10_u4_n2042 ) );
NAND3_X1 _u10_u4_U98  ( .A1(_u10_u4_n2040 ), .A2(_u10_u4_n2041 ), .A3(_u10_u4_n2042 ), .ZN(_u10_u4_n2009 ) );
AND2_X1 _u10_u4_U97  ( .A1(_u10_u4_n2038 ), .A2(_u10_u4_n2039 ), .ZN(_u10_u4_n1929 ) );
NOR2_X1 _u10_u4_U96  ( .A1(_u10_u4_n1929 ), .A2(_u10_u4_n2037 ), .ZN(_u10_u4_n2010 ) );
NAND2_X1 _u10_u4_U95  ( .A1(_u10_u4_n2035 ), .A2(_u10_u4_n2036 ), .ZN(_u10_u4_n1902 ) );
NAND3_X1 _u10_u4_U94  ( .A1(_u10_u4_n1902 ), .A2(_u10_u4_n2033 ), .A3(_u10_u4_n2034 ), .ZN(_u10_u4_n1973 ) );
NOR2_X1 _u10_u4_U93  ( .A1(_u10_u4_n1978 ), .A2(_u10_u4_n1973 ), .ZN(_u10_u4_n2032 ) );
NOR2_X1 _u10_u4_U92  ( .A1(1'b0), .A2(_u10_u4_n2032 ), .ZN(_u10_u4_n2028 ));
NOR2_X1 _u10_u4_U91  ( .A1(_u10_u4_n2030 ), .A2(_u10_u4_n2031 ), .ZN(_u10_u4_n2029 ) );
NOR4_X1 _u10_u4_U90  ( .A1(_u10_u4_n2026 ), .A2(_u10_u4_n2027 ), .A3(_u10_u4_n2028 ), .A4(_u10_u4_n2029 ), .ZN(_u10_u4_n2024 ) );
NOR2_X1 _u10_u4_U89  ( .A1(_u10_u4_n2024 ), .A2(_u10_u4_n2025 ), .ZN(_u10_u4_n2011 ) );
NAND3_X1 _u10_u4_U88  ( .A1(_u10_u4_n2021 ), .A2(_u10_u4_n2022 ), .A3(_u10_u4_n2023 ), .ZN(_u10_u4_n2020 ) );
AND2_X1 _u10_u4_U87  ( .A1(_u10_u4_n2019 ), .A2(_u10_u4_n2020 ), .ZN(_u10_u4_n1838 ) );
INV_X1 _u10_u4_U86  ( .A(_u10_u4_n2018 ), .ZN(_u10_u4_n2016 ) );
NOR4_X1 _u10_u4_U85  ( .A1(_u10_u4_n2015 ), .A2(_u10_u4_n1838 ), .A3(_u10_u4_n2016 ), .A4(_u10_u4_n2017 ), .ZN(_u10_u4_n2013 ) );
NOR2_X1 _u10_u4_U84  ( .A1(_u10_u4_n2013 ), .A2(_u10_u4_n2014 ), .ZN(_u10_u4_n2012 ) );
NOR4_X1 _u10_u4_U83  ( .A1(_u10_u4_n2009 ), .A2(_u10_u4_n2010 ), .A3(_u10_u4_n2011 ), .A4(_u10_u4_n2012 ), .ZN(_u10_u4_n1821 ) );
NAND2_X1 _u10_u4_U82  ( .A1(_u10_u4_n1924 ), .A2(_u10_u4_n2008 ), .ZN(_u10_u4_n1993 ) );
NAND2_X1 _u10_u4_U81  ( .A1(_u10_u4_n2006 ), .A2(_u10_u4_n2007 ), .ZN(_u10_u4_n1994 ) );
NAND2_X1 _u10_u4_U80  ( .A1(_u10_u4_n2004 ), .A2(_u10_u4_n2005 ), .ZN(_u10_u4_n1995 ) );
AND2_X1 _u10_u4_U79  ( .A1(_u10_u4_n2002 ), .A2(_u10_u4_n2003 ), .ZN(_u10_u4_n1998 ) );
NOR2_X1 _u10_u4_U78  ( .A1(_u10_u4_n2000 ), .A2(_u10_u4_n2001 ), .ZN(_u10_u4_n1999 ) );
NOR3_X1 _u10_u4_U77  ( .A1(_u10_u4_n1997 ), .A2(_u10_u4_n1998 ), .A3(_u10_u4_n1999 ), .ZN(_u10_u4_n1996 ) );
NAND4_X1 _u10_u4_U76  ( .A1(_u10_u4_n1993 ), .A2(_u10_u4_n1994 ), .A3(_u10_u4_n1995 ), .A4(_u10_u4_n1996 ), .ZN(_u10_u4_n1985 ) );
INV_X1 _u10_u4_U75  ( .A(_u10_u4_n1992 ), .ZN(_u10_u4_n1989 ) );
NAND3_X1 _u10_u4_U74  ( .A1(_u10_u4_n1989 ), .A2(_u10_u4_n1990 ), .A3(_u10_u4_n1991 ), .ZN(_u10_u4_n1986 ) );
NOR4_X1 _u10_u4_U73  ( .A1(_u10_u4_n1985 ), .A2(_u10_u4_n1986 ), .A3(_u10_u4_n1987 ), .A4(_u10_u4_n1988 ), .ZN(_u10_u4_n1822 ) );
INV_X1 _u10_u4_U72  ( .A(_u10_u4_n1984 ), .ZN(_u10_u4_n1980 ) );
NAND4_X1 _u10_u4_U71  ( .A1(_u10_u4_n1980 ), .A2(_u10_u4_n1981 ), .A3(_u10_u4_n1982 ), .A4(_u10_u4_n1983 ), .ZN(_u10_u4_n1941 ) );
NOR3_X1 _u10_u4_U70  ( .A1(_u10_u4_n1977 ), .A2(_u10_u4_n1978 ), .A3(_u10_u4_n1979 ), .ZN(_u10_u4_n1971 ) );
NOR4_X1 _u10_u4_U69  ( .A1(_u10_u4_n1973 ), .A2(_u10_u4_n1974 ), .A3(_u10_u4_n1975 ), .A4(_u10_u4_n1976 ), .ZN(_u10_u4_n1972 ) );
NAND4_X1 _u10_u4_U68  ( .A1(_u10_u4_n1969 ), .A2(_u10_u4_n1970 ), .A3(_u10_u4_n1971 ), .A4(_u10_u4_n1972 ), .ZN(_u10_u4_n1968 ) );
NAND2_X1 _u10_u4_U67  ( .A1(_u10_u4_n1967 ), .A2(_u10_u4_n1968 ), .ZN(_u10_u4_n1942 ) );
NAND3_X1 _u10_u4_U66  ( .A1(_u10_u4_n1964 ), .A2(_u10_u4_n1965 ), .A3(_u10_u4_n1966 ), .ZN(_u10_u4_n1943 ) );
AND4_X1 _u10_u4_U65  ( .A1(_u10_u4_n1961 ), .A2(_u10_u4_n1863 ), .A3(_u10_u4_n1962 ), .A4(_u10_u4_n1963 ), .ZN(_u10_u4_n1957 ) );
NOR2_X1 _u10_u4_U64  ( .A1(_u10_u4_n1959 ), .A2(_u10_u4_n1960 ), .ZN(_u10_u4_n1958 ) );
NOR2_X1 _u10_u4_U63  ( .A1(_u10_u4_n1957 ), .A2(_u10_u4_n1958 ), .ZN(_u10_u4_n1945 ) );
NOR2_X1 _u10_u4_U62  ( .A1(_u10_u4_n1955 ), .A2(_u10_u4_n1956 ), .ZN(_u10_u4_n1953 ) );
NOR4_X1 _u10_u4_U61  ( .A1(_u10_u4_n1952 ), .A2(_u10_u4_n1953 ), .A3(_u10_u4_n1846 ), .A4(_u10_u4_n1954 ), .ZN(_u10_u4_n1946 ) );
NOR2_X1 _u10_u4_U60  ( .A1(_u10_u4_n1950 ), .A2(_u10_u4_n1951 ), .ZN(_u10_u4_n1949 ) );
NOR2_X1 _u10_u4_U59  ( .A1(_u10_u4_n1948 ), .A2(_u10_u4_n1949 ), .ZN(_u10_u4_n1947 ) );
NOR3_X1 _u10_u4_U58  ( .A1(_u10_u4_n1945 ), .A2(_u10_u4_n1946 ), .A3(_u10_u4_n1947 ), .ZN(_u10_u4_n1944 ) );
NAND4_X1 _u10_u4_U57  ( .A1(_u10_u4_n1941 ), .A2(_u10_u4_n1942 ), .A3(_u10_u4_n1943 ), .A4(_u10_u4_n1944 ), .ZN(_u10_u4_n1824 ) );
NAND2_X1 _u10_u4_U56  ( .A1(_u10_u4_n1939 ), .A2(_u10_u4_n1940 ), .ZN(_u10_u4_n1938 ) );
NAND2_X1 _u10_u4_U55  ( .A1(_u10_u4_n1937 ), .A2(_u10_u4_n1938 ), .ZN(_u10_u4_n1903 ) );
NAND2_X1 _u10_u4_U54  ( .A1(_u10_u4_n1935 ), .A2(_u10_u4_n1936 ), .ZN(_u10_u4_n1934 ) );
NAND2_X1 _u10_u4_U53  ( .A1(_u10_u4_n1933 ), .A2(_u10_u4_n1934 ), .ZN(_u10_u4_n1931 ) );
NAND2_X1 _u10_u4_U52  ( .A1(_u10_u4_n1931 ), .A2(_u10_u4_n1932 ), .ZN(_u10_u4_n1904 ) );
NAND2_X1 _u10_u4_U51  ( .A1(_u10_u4_n1929 ), .A2(_u10_u4_n1930 ), .ZN(_u10_u4_n1927 ) );
NAND2_X1 _u10_u4_U50  ( .A1(_u10_u4_n1927 ), .A2(_u10_u4_n1928 ), .ZN(_u10_u4_n1905 ) );
NOR3_X1 _u10_u4_U49  ( .A1(_u10_u4_n1916 ), .A2(_u10_u4_n1925 ), .A3(_u10_u4_n1926 ), .ZN(_u10_u4_n1919 ) );
NOR2_X1 _u10_u4_U48  ( .A1(_u10_u4_n1923 ), .A2(_u10_u4_n1924 ), .ZN(_u10_u4_n1921 ) );
NOR2_X1 _u10_u4_U47  ( .A1(_u10_u4_n1921 ), .A2(_u10_u4_n1922 ), .ZN(_u10_u4_n1920 ) );
NOR2_X1 _u10_u4_U46  ( .A1(_u10_u4_n1919 ), .A2(_u10_u4_n1920 ), .ZN(_u10_u4_n1917 ) );
NOR2_X1 _u10_u4_U45  ( .A1(_u10_u4_n1917 ), .A2(_u10_u4_n1918 ), .ZN(_u10_u4_n1907 ) );
NOR2_X1 _u10_u4_U44  ( .A1(_u10_u4_n1915 ), .A2(_u10_u4_n1916 ), .ZN(_u10_u4_n1914 ) );
NOR2_X1 _u10_u4_U43  ( .A1(_u10_u4_n1914 ), .A2(1'b0), .ZN(_u10_u4_n1912 ));
NOR2_X1 _u10_u4_U42  ( .A1(_u10_u4_n1912 ), .A2(_u10_u4_n1913 ), .ZN(_u10_u4_n1908 ) );
NOR2_X1 _u10_u4_U41  ( .A1(_u10_u4_n1891 ), .A2(_u10_u4_n1911 ), .ZN(_u10_u4_n1910 ) );
NOR2_X1 _u10_u4_U40  ( .A1(_u10_u4_n1910 ), .A2(_u10_u4_n1868 ), .ZN(_u10_u4_n1909 ) );
NOR3_X1 _u10_u4_U39  ( .A1(_u10_u4_n1907 ), .A2(_u10_u4_n1908 ), .A3(_u10_u4_n1909 ), .ZN(_u10_u4_n1906 ) );
NAND4_X1 _u10_u4_U38  ( .A1(_u10_u4_n1903 ), .A2(_u10_u4_n1904 ), .A3(_u10_u4_n1905 ), .A4(_u10_u4_n1906 ), .ZN(_u10_u4_n1825 ) );
NAND2_X1 _u10_u4_U37  ( .A1(_u10_u4_n1901 ), .A2(_u10_u4_n1902 ), .ZN(_u10_u4_n1900 ) );
NAND2_X1 _u10_u4_U36  ( .A1(_u10_u4_n1899 ), .A2(_u10_u4_n1900 ), .ZN(_u10_u4_n1875 ) );
OR2_X1 _u10_u4_U35  ( .A1(_u10_u4_n1847 ), .A2(_u10_u4_n1898 ), .ZN(_u10_u4_n1897 ) );
NAND2_X1 _u10_u4_U34  ( .A1(_u10_u4_n1896 ), .A2(_u10_u4_n1897 ), .ZN(_u10_u4_n1895 ) );
NAND2_X1 _u10_u4_U33  ( .A1(_u10_u4_n1894 ), .A2(_u10_u4_n1895 ), .ZN(_u10_u4_n1876 ) );
NAND2_X1 _u10_u4_U32  ( .A1(_u10_u4_n1892 ), .A2(_u10_u4_n1893 ), .ZN(_u10_u4_n1877 ) );
NOR3_X1 _u10_u4_U31  ( .A1(_u10_u4_n1884 ), .A2(_u10_u4_n1890 ), .A3(_u10_u4_n1891 ), .ZN(_u10_u4_n1889 ) );
NOR2_X1 _u10_u4_U30  ( .A1(_u10_u4_n1840 ), .A2(_u10_u4_n1889 ), .ZN(_u10_u4_n1879 ) );
NOR2_X1 _u10_u4_U29  ( .A1(_u10_u4_n1887 ), .A2(_u10_u4_n1888 ), .ZN(_u10_u4_n1880 ) );
NOR3_X1 _u10_u4_U28  ( .A1(_u10_u4_n1884 ), .A2(_u10_u4_n1885 ), .A3(_u10_u4_n1886 ), .ZN(_u10_u4_n1883 ) );
NOR2_X1 _u10_u4_U27  ( .A1(_u10_u4_n1882 ), .A2(_u10_u4_n1883 ), .ZN(_u10_u4_n1881 ) );
NOR3_X1 _u10_u4_U26  ( .A1(_u10_u4_n1879 ), .A2(_u10_u4_n1880 ), .A3(_u10_u4_n1881 ), .ZN(_u10_u4_n1878 ) );
NAND4_X1 _u10_u4_U25  ( .A1(_u10_u4_n1875 ), .A2(_u10_u4_n1876 ), .A3(_u10_u4_n1877 ), .A4(_u10_u4_n1878 ), .ZN(_u10_u4_n1826 ) );
NOR3_X1 _u10_u4_U24  ( .A1(_u10_u4_n1872 ), .A2(_u10_u4_n1873 ), .A3(_u10_u4_n1874 ), .ZN(_u10_u4_n1871 ) );
NAND4_X1 _u10_u4_U23  ( .A1(_u10_u4_n1868 ), .A2(_u10_u4_n1869 ), .A3(_u10_u4_n1870 ), .A4(_u10_u4_n1871 ), .ZN(_u10_u4_n1867 ) );
NAND2_X1 _u10_u4_U22  ( .A1(_u10_u4_n1866 ), .A2(_u10_u4_n1867 ), .ZN(_u10_u4_n1865 ) );
NAND3_X1 _u10_u4_U21  ( .A1(_u10_u4_n1863 ), .A2(_u10_u4_n1864 ), .A3(_u10_u4_n1865 ), .ZN(_u10_u4_n1862 ) );
NAND2_X1 _u10_u4_U20  ( .A1(_u10_u4_n1861 ), .A2(_u10_u4_n1862 ), .ZN(_u10_u4_n1828 ) );
NAND3_X1 _u10_u4_U19  ( .A1(_u10_u4_n1858 ), .A2(_u10_u4_n1859 ), .A3(_u10_u4_n1860 ), .ZN(_u10_u4_n1857 ) );
NAND2_X1 _u10_u4_U18  ( .A1(_u10_u4_n1856 ), .A2(_u10_u4_n1857 ), .ZN(_u10_u4_n1829 ) );
OR2_X1 _u10_u4_U17  ( .A1(_u10_u4_n1854 ), .A2(_u10_u4_n1855 ), .ZN(_u10_u4_n1830 ) );
NOR2_X1 _u10_u4_U16  ( .A1(_u10_u4_n1852 ), .A2(_u10_u4_n1853 ), .ZN(_u10_u4_n1850 ) );
NOR3_X1 _u10_u4_U15  ( .A1(_u10_u4_n1850 ), .A2(_u10_u4_n1851 ), .A3(_u10_u4_n1838 ), .ZN(_u10_u4_n1848 ) );
NOR2_X1 _u10_u4_U14  ( .A1(_u10_u4_n1848 ), .A2(_u10_u4_n1849 ), .ZN(_u10_u4_n1832 ) );
NOR2_X1 _u10_u4_U13  ( .A1(_u10_u4_n1846 ), .A2(_u10_u4_n1847 ), .ZN(_u10_u4_n1845 ) );
NOR3_X1 _u10_u4_U12  ( .A1(_u10_u4_n1844 ), .A2(1'b0), .A3(_u10_u4_n1845 ),.ZN(_u10_u4_n1842 ) );
NOR2_X1 _u10_u4_U11  ( .A1(_u10_u4_n1842 ), .A2(_u10_u4_n1843 ), .ZN(_u10_u4_n1833 ) );
NOR2_X1 _u10_u4_U10  ( .A1(_u10_u4_n1840 ), .A2(_u10_u4_n1841 ), .ZN(_u10_u4_n1839 ) );
NOR3_X1 _u10_u4_U9  ( .A1(_u10_u4_n1837 ), .A2(_u10_u4_n1838 ), .A3(_u10_u4_n1839 ), .ZN(_u10_u4_n1835 ) );
NOR2_X1 _u10_u4_U8  ( .A1(_u10_u4_n1835 ), .A2(_u10_u4_n1836 ), .ZN(_u10_u4_n1834 ) );
NOR3_X1 _u10_u4_U7  ( .A1(_u10_u4_n1832 ), .A2(_u10_u4_n1833 ), .A3(_u10_u4_n1834 ), .ZN(_u10_u4_n1831 ) );
NAND4_X1 _u10_u4_U6  ( .A1(_u10_u4_n1828 ), .A2(_u10_u4_n1829 ), .A3(_u10_u4_n1830 ), .A4(_u10_u4_n1831 ), .ZN(_u10_u4_n1827 ) );
NOR4_X1 _u10_u4_U5  ( .A1(_u10_u4_n1824 ), .A2(_u10_u4_n1825 ), .A3(_u10_u4_n1826 ), .A4(_u10_u4_n1827 ), .ZN(_u10_u4_n1823 ) );
NAND4_X1 _u10_u4_U4  ( .A1(_u10_u4_n1820 ), .A2(_u10_u4_n1821 ), .A3(_u10_u4_n1822 ), .A4(_u10_u4_n1823 ), .ZN(_u10_u4_n1818 ) );
MUX2_X1 _u10_u4_U3  ( .A(_u10_u4_n1818 ), .B(_u10_SYNOPSYS_UNCONNECTED_17 ),.S(_u10_u4_n1819 ), .Z(_u10_u4_n1812 ) );
DFFR_X1 _u10_u4_state_reg_1_  ( .D(_u10_u4_n1812 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_17 ), .QN(_u10_u4_n1814 ));
DFFR_X1 _u10_u4_state_reg_2_  ( .D(_u10_u4_n1811 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_16 ), .QN(_u10_u4_n1815 ));
DFFR_X1 _u10_u4_state_reg_3_  ( .D(_u10_u4_n1810 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_15 ), .QN(_u10_u4_n1816 ));
DFFR_X1 _u10_u4_state_reg_4_  ( .D(_u10_u4_n1809 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_14 ), .QN(_u10_u4_n1817 ));
DFFR_X1 _u10_u4_state_reg_0_  ( .D(_u10_u4_n1808 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_18 ), .QN(_u10_u4_n1813 ));
NOR2_X1 _u10_u5_U1606  ( .A1(_u10_SYNOPSYS_UNCONNECTED_21 ), .A2(_u10_u5_n1814 ), .ZN(_u10_u5_n3174 ) );
NOR3_X1 _u10_u5_U1605  ( .A1(_u10_SYNOPSYS_UNCONNECTED_20 ), .A2(_u10_u5_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_23 ), .ZN(_u10_u5_n3328 ) );
NAND2_X1 _u10_u5_U1604  ( .A1(_u10_u5_n3174 ), .A2(_u10_u5_n3328 ), .ZN(_u10_u5_n1843 ) );
INV_X1 _u10_u5_U1603  ( .A(_u10_u5_n1843 ), .ZN(_u10_u5_n2461 ) );
INV_X1 _u10_u5_U1602  ( .A(1'b0), .ZN(_u10_u5_n2466 ) );
INV_X1 _u10_u5_U1601  ( .A(1'b0), .ZN(_u10_u5_n2305 ) );
NAND2_X1 _u10_u5_U1600  ( .A1(_u10_u5_n2466 ), .A2(_u10_u5_n2305 ), .ZN(_u10_u5_n1954 ) );
INV_X1 _u10_u5_U1599  ( .A(_u10_u5_n1954 ), .ZN(_u10_u5_n2467 ) );
INV_X1 _u10_u5_U1598  ( .A(1'b0), .ZN(_u10_u5_n1936 ) );
NOR2_X1 _u10_u5_U1597  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u5_n2223 ) );
INV_X1 _u10_u5_U1596  ( .A(1'b0), .ZN(_u10_u5_n1922 ) );
NAND2_X1 _u10_u5_U1595  ( .A1(_u10_u5_n2223 ), .A2(_u10_u5_n1922 ), .ZN(_u10_u5_n2200 ) );
NOR2_X1 _u10_u5_U1594  ( .A1(_u10_u5_n2200 ), .A2(1'b0), .ZN(_u10_u5_n2502 ));
INV_X1 _u10_u5_U1593  ( .A(1'b0), .ZN(_u10_u5_n2978 ) );
INV_X1 _u10_u5_U1592  ( .A(1'b0), .ZN(_u10_u5_n3000 ) );
NAND2_X1 _u10_u5_U1591  ( .A1(_u10_u5_n2978 ), .A2(_u10_u5_n3000 ), .ZN(_u10_u5_n3356 ) );
INV_X1 _u10_u5_U1590  ( .A(1'b0), .ZN(_u10_u5_n2405 ) );
INV_X1 _u10_u5_U1589  ( .A(1'b0), .ZN(_u10_u5_n2972 ) );
NAND2_X1 _u10_u5_U1588  ( .A1(_u10_u5_n2405 ), .A2(_u10_u5_n2972 ), .ZN(_u10_u5_n2008 ) );
NOR2_X1 _u10_u5_U1587  ( .A1(_u10_u5_n3356 ), .A2(_u10_u5_n2008 ), .ZN(_u10_u5_n2195 ) );
NAND2_X1 _u10_u5_U1586  ( .A1(_u10_u5_n2502 ), .A2(_u10_u5_n2195 ), .ZN(_u10_u5_n2490 ) );
INV_X1 _u10_u5_U1585  ( .A(1'b0), .ZN(_u10_u5_n3040 ) );
INV_X1 _u10_u5_U1584  ( .A(1'b0), .ZN(_u10_u5_n3006 ) );
NAND2_X1 _u10_u5_U1583  ( .A1(_u10_u5_n3040 ), .A2(_u10_u5_n3006 ), .ZN(_u10_u5_n2508 ) );
NOR2_X1 _u10_u5_U1582  ( .A1(_u10_u5_n2508 ), .A2(1'b0), .ZN(_u10_u5_n2493 ));
INV_X1 _u10_u5_U1581  ( .A(1'b0), .ZN(_u10_u5_n2038 ) );
NAND2_X1 _u10_u5_U1580  ( .A1(_u10_u5_n2493 ), .A2(_u10_u5_n2038 ), .ZN(_u10_u5_n2174 ) );
NOR2_X1 _u10_u5_U1579  ( .A1(_u10_u5_n2490 ), .A2(_u10_u5_n2174 ), .ZN(_u10_u5_n2659 ) );
INV_X1 _u10_u5_U1578  ( .A(1'b0), .ZN(_u10_u5_n2175 ) );
NAND3_X1 _u10_u5_U1577  ( .A1(_u10_u5_n2659 ), .A2(_u10_u5_n2175 ), .A3(1'b0), .ZN(_u10_u5_n3189 ) );
NOR2_X1 _u10_u5_U1576  ( .A1(_u10_u5_n3189 ), .A2(1'b0), .ZN(_u10_u5_n2528 ));
INV_X1 _u10_u5_U1575  ( .A(1'b0), .ZN(_u10_u5_n2837 ) );
NAND2_X1 _u10_u5_U1574  ( .A1(_u10_u5_n2528 ), .A2(_u10_u5_n2837 ), .ZN(_u10_u5_n2567 ) );
INV_X1 _u10_u5_U1573  ( .A(1'b0), .ZN(_u10_u5_n2080 ) );
INV_X1 _u10_u5_U1572  ( .A(1'b0), .ZN(_u10_u5_n2166 ) );
NAND2_X1 _u10_u5_U1571  ( .A1(_u10_u5_n2080 ), .A2(_u10_u5_n2166 ), .ZN(_u10_u5_n2840 ) );
NOR2_X1 _u10_u5_U1570  ( .A1(_u10_u5_n2567 ), .A2(_u10_u5_n2840 ), .ZN(_u10_u5_n2443 ) );
INV_X1 _u10_u5_U1569  ( .A(1'b0), .ZN(_u10_u5_n2600 ) );
INV_X1 _u10_u5_U1568  ( .A(1'b0), .ZN(_u10_u5_n2836 ) );
NAND2_X1 _u10_u5_U1567  ( .A1(_u10_u5_n2600 ), .A2(_u10_u5_n2836 ), .ZN(_u10_u5_n2428 ) );
INV_X1 _u10_u5_U1566  ( .A(_u10_u5_n2428 ), .ZN(_u10_u5_n2078 ) );
NAND2_X1 _u10_u5_U1565  ( .A1(_u10_u5_n2443 ), .A2(_u10_u5_n2078 ), .ZN(_u10_u5_n2282 ) );
INV_X1 _u10_u5_U1564  ( .A(1'b0), .ZN(_u10_u5_n2874 ) );
INV_X1 _u10_u5_U1563  ( .A(1'b0), .ZN(_u10_u5_n2031 ) );
NAND2_X1 _u10_u5_U1562  ( .A1(_u10_u5_n2874 ), .A2(_u10_u5_n2031 ), .ZN(_u10_u5_n1976 ) );
NOR2_X1 _u10_u5_U1561  ( .A1(_u10_u5_n2282 ), .A2(_u10_u5_n1976 ), .ZN(_u10_u5_n2411 ) );
NAND3_X1 _u10_u5_U1560  ( .A1(_u10_u5_n2467 ), .A2(_u10_u5_n1936 ), .A3(_u10_u5_n2411 ), .ZN(_u10_u5_n2464 ) );
NAND3_X1 _u10_u5_U1559  ( .A1(_u10_u5_n2166 ), .A2(_u10_u5_n2837 ), .A3(1'b0), .ZN(_u10_u5_n3276 ) );
INV_X1 _u10_u5_U1558  ( .A(_u10_u5_n3276 ), .ZN(_u10_u5_n2442 ) );
NAND3_X1 _u10_u5_U1557  ( .A1(_u10_u5_n2836 ), .A2(_u10_u5_n2080 ), .A3(_u10_u5_n2442 ), .ZN(_u10_u5_n2838 ) );
INV_X1 _u10_u5_U1556  ( .A(_u10_u5_n2838 ), .ZN(_u10_u5_n2850 ) );
NOR2_X1 _u10_u5_U1555  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u5_n2953 ) );
NAND2_X1 _u10_u5_U1554  ( .A1(_u10_u5_n2850 ), .A2(_u10_u5_n2953 ), .ZN(_u10_u5_n2947 ) );
INV_X1 _u10_u5_U1553  ( .A(_u10_u5_n2947 ), .ZN(_u10_u5_n2420 ) );
NAND2_X1 _u10_u5_U1552  ( .A1(_u10_u5_n1936 ), .A2(_u10_u5_n2874 ), .ZN(_u10_u5_n2030 ) );
INV_X1 _u10_u5_U1551  ( .A(_u10_u5_n2030 ), .ZN(_u10_u5_n2162 ) );
NAND2_X1 _u10_u5_U1550  ( .A1(_u10_u5_n2420 ), .A2(_u10_u5_n2162 ), .ZN(_u10_u5_n2828 ) );
INV_X1 _u10_u5_U1549  ( .A(_u10_u5_n2828 ), .ZN(_u10_u5_n2551 ) );
NAND2_X1 _u10_u5_U1548  ( .A1(_u10_u5_n2551 ), .A2(_u10_u5_n2467 ), .ZN(_u10_u5_n3416 ) );
NAND2_X1 _u10_u5_U1547  ( .A1(_u10_u5_n2464 ), .A2(_u10_u5_n3416 ), .ZN(_u10_u5_n2266 ) );
INV_X1 _u10_u5_U1546  ( .A(_u10_u5_n2266 ), .ZN(_u10_u5_n3410 ) );
NAND2_X1 _u10_u5_U1545  ( .A1(1'b0), .A2(_u10_u5_n2305 ), .ZN(_u10_u5_n3411 ) );
INV_X1 _u10_u5_U1544  ( .A(_u10_u5_n3356 ), .ZN(_u10_u5_n1983 ) );
NAND3_X1 _u10_u5_U1543  ( .A1(_u10_u5_n1983 ), .A2(_u10_u5_n2405 ), .A3(1'b0), .ZN(_u10_u5_n2022 ) );
INV_X1 _u10_u5_U1542  ( .A(_u10_u5_n2022 ), .ZN(_u10_u5_n2056 ) );
INV_X1 _u10_u5_U1541  ( .A(_u10_u5_n2840 ), .ZN(_u10_u5_n2059 ) );
INV_X1 _u10_u5_U1540  ( .A(1'b0), .ZN(_u10_u5_n1965 ) );
NAND2_X1 _u10_u5_U1539  ( .A1(_u10_u5_n2837 ), .A2(_u10_u5_n1965 ), .ZN(_u10_u5_n1852 ) );
INV_X1 _u10_u5_U1538  ( .A(_u10_u5_n1852 ), .ZN(_u10_u5_n3190 ) );
INV_X1 _u10_u5_U1537  ( .A(1'b0), .ZN(_u10_u5_n1853 ) );
NAND2_X1 _u10_u5_U1536  ( .A1(_u10_u5_n3190 ), .A2(_u10_u5_n1853 ), .ZN(_u10_u5_n2687 ) );
INV_X1 _u10_u5_U1535  ( .A(_u10_u5_n2687 ), .ZN(_u10_u5_n2019 ) );
NAND2_X1 _u10_u5_U1534  ( .A1(_u10_u5_n2059 ), .A2(_u10_u5_n2019 ), .ZN(_u10_u5_n2330 ) );
NOR2_X1 _u10_u5_U1533  ( .A1(_u10_u5_n2428 ), .A2(_u10_u5_n2330 ), .ZN(_u10_u5_n2036 ) );
NAND2_X1 _u10_u5_U1532  ( .A1(_u10_u5_n2056 ), .A2(_u10_u5_n2036 ), .ZN(_u10_u5_n3379 ) );
NOR2_X1 _u10_u5_U1531  ( .A1(_u10_u5_n3379 ), .A2(_u10_u5_n2030 ), .ZN(_u10_u5_n2026 ) );
INV_X1 _u10_u5_U1530  ( .A(1'b0), .ZN(_u10_u5_n2431 ) );
NOR2_X1 _u10_u5_U1529  ( .A1(_u10_u5_n2431 ), .A2(1'b0), .ZN(_u10_u5_n3062 ));
NAND2_X1 _u10_u5_U1528  ( .A1(_u10_u5_n3062 ), .A2(_u10_u5_n2195 ), .ZN(_u10_u5_n3407 ) );
NOR3_X1 _u10_u5_U1527  ( .A1(_u10_u5_n2687 ), .A2(1'b0), .A3(_u10_u5_n3407 ),.ZN(_u10_u5_n3275 ) );
NAND3_X1 _u10_u5_U1526  ( .A1(_u10_u5_n2836 ), .A2(_u10_u5_n2080 ), .A3(_u10_u5_n3275 ), .ZN(_u10_u5_n3297 ) );
INV_X1 _u10_u5_U1525  ( .A(_u10_u5_n3297 ), .ZN(_u10_u5_n3172 ) );
NAND2_X1 _u10_u5_U1524  ( .A1(_u10_u5_n3172 ), .A2(_u10_u5_n2600 ), .ZN(_u10_u5_n2226 ) );
NOR2_X1 _u10_u5_U1523  ( .A1(_u10_u5_n2226 ), .A2(1'b0), .ZN(_u10_u5_n2307 ));
INV_X1 _u10_u5_U1522  ( .A(_u10_u5_n2490 ), .ZN(_u10_u5_n2536 ) );
NAND3_X1 _u10_u5_U1521  ( .A1(_u10_u5_n2536 ), .A2(_u10_u5_n3040 ), .A3(1'b0), .ZN(_u10_u5_n3226 ) );
NOR2_X1 _u10_u5_U1520  ( .A1(_u10_u5_n3226 ), .A2(_u10_u5_n2330 ), .ZN(_u10_u5_n2441 ) );
NAND2_X1 _u10_u5_U1519  ( .A1(_u10_u5_n2441 ), .A2(_u10_u5_n2953 ), .ZN(_u10_u5_n2579 ) );
NOR2_X1 _u10_u5_U1518  ( .A1(_u10_u5_n2579 ), .A2(_u10_u5_n2030 ), .ZN(_u10_u5_n2550 ) );
NOR3_X1 _u10_u5_U1517  ( .A1(_u10_u5_n2026 ), .A2(_u10_u5_n2307 ), .A3(_u10_u5_n2550 ), .ZN(_u10_u5_n3394 ) );
NAND2_X1 _u10_u5_U1516  ( .A1(1'b0), .A2(_u10_u5_n2978 ), .ZN(_u10_u5_n3115 ) );
NOR2_X1 _u10_u5_U1515  ( .A1(_u10_u5_n3115 ), .A2(_u10_u5_n2330 ), .ZN(_u10_u5_n3126 ) );
NAND2_X1 _u10_u5_U1514  ( .A1(_u10_u5_n2162 ), .A2(_u10_u5_n2031 ), .ZN(_u10_u5_n2686 ) );
NOR2_X1 _u10_u5_U1513  ( .A1(_u10_u5_n2686 ), .A2(_u10_u5_n2428 ), .ZN(_u10_u5_n2108 ) );
NAND2_X1 _u10_u5_U1512  ( .A1(_u10_u5_n3126 ), .A2(_u10_u5_n2108 ), .ZN(_u10_u5_n3415 ) );
NAND2_X1 _u10_u5_U1511  ( .A1(_u10_u5_n3394 ), .A2(_u10_u5_n3415 ), .ZN(_u10_u5_n3089 ) );
NAND2_X1 _u10_u5_U1510  ( .A1(_u10_u5_n3089 ), .A2(_u10_u5_n2305 ), .ZN(_u10_u5_n3414 ) );
NAND2_X1 _u10_u5_U1509  ( .A1(_u10_u5_n2466 ), .A2(_u10_u5_n3414 ), .ZN(_u10_u5_n3118 ) );
NAND2_X1 _u10_u5_U1508  ( .A1(_u10_u5_n2078 ), .A2(_u10_u5_n2080 ), .ZN(_u10_u5_n2596 ) );
NAND2_X1 _u10_u5_U1507  ( .A1(1'b0), .A2(_u10_u5_n2493 ), .ZN(_u10_u5_n1961 ) );
NOR3_X1 _u10_u5_U1506  ( .A1(_u10_u5_n2490 ), .A2(1'b0), .A3(_u10_u5_n1961 ),.ZN(_u10_u5_n2054 ) );
NAND2_X1 _u10_u5_U1505  ( .A1(_u10_u5_n2054 ), .A2(_u10_u5_n3190 ), .ZN(_u10_u5_n2061 ) );
OR2_X1 _u10_u5_U1504  ( .A1(_u10_u5_n2596 ), .A2(_u10_u5_n2061 ), .ZN(_u10_u5_n1969 ) );
NOR3_X1 _u10_u5_U1503  ( .A1(_u10_u5_n1976 ), .A2(1'b0), .A3(_u10_u5_n1969 ),.ZN(_u10_u5_n2710 ) );
NAND2_X1 _u10_u5_U1502  ( .A1(_u10_u5_n2710 ), .A2(_u10_u5_n2467 ), .ZN(_u10_u5_n2545 ) );
INV_X1 _u10_u5_U1501  ( .A(_u10_u5_n2545 ), .ZN(_u10_u5_n2087 ) );
NOR2_X1 _u10_u5_U1500  ( .A1(_u10_u5_n3118 ), .A2(_u10_u5_n2087 ), .ZN(_u10_u5_n3145 ) );
NOR2_X1 _u10_u5_U1499  ( .A1(_u10_u5_n2030 ), .A2(1'b0), .ZN(_u10_u5_n2668 ));
NAND2_X1 _u10_u5_U1498  ( .A1(1'b0), .A2(_u10_u5_n2668 ), .ZN(_u10_u5_n2163 ) );
INV_X1 _u10_u5_U1497  ( .A(_u10_u5_n2163 ), .ZN(_u10_u5_n2875 ) );
INV_X1 _u10_u5_U1496  ( .A(_u10_u5_n1976 ), .ZN(_u10_u5_n2747 ) );
NAND3_X1 _u10_u5_U1495  ( .A1(_u10_u5_n2747 ), .A2(_u10_u5_n2600 ), .A3(1'b0), .ZN(_u10_u5_n3393 ) );
NOR3_X1 _u10_u5_U1494  ( .A1(1'b0), .A2(1'b0), .A3(_u10_u5_n3393 ), .ZN(_u10_u5_n3180 ) );
INV_X1 _u10_u5_U1493  ( .A(1'b0), .ZN(_u10_u5_n2113 ) );
INV_X1 _u10_u5_U1492  ( .A(1'b0), .ZN(_u10_u5_n3066 ) );
NAND2_X1 _u10_u5_U1491  ( .A1(_u10_u5_n2175 ), .A2(_u10_u5_n3066 ), .ZN(_u10_u5_n2216 ) );
INV_X1 _u10_u5_U1490  ( .A(_u10_u5_n2659 ), .ZN(_u10_u5_n2643 ) );
NOR2_X1 _u10_u5_U1489  ( .A1(_u10_u5_n2216 ), .A2(_u10_u5_n2643 ), .ZN(_u10_u5_n2049 ) );
AND2_X1 _u10_u5_U1488  ( .A1(_u10_u5_n2049 ), .A2(_u10_u5_n1853 ), .ZN(_u10_u5_n3223 ) );
NAND2_X1 _u10_u5_U1487  ( .A1(_u10_u5_n3223 ), .A2(_u10_u5_n1965 ), .ZN(_u10_u5_n2531 ) );
NOR2_X1 _u10_u5_U1486  ( .A1(_u10_u5_n2531 ), .A2(1'b0), .ZN(_u10_u5_n2884 ));
NAND2_X1 _u10_u5_U1485  ( .A1(_u10_u5_n2884 ), .A2(_u10_u5_n2166 ), .ZN(_u10_u5_n1841 ) );
NOR2_X1 _u10_u5_U1484  ( .A1(_u10_u5_n1841 ), .A2(1'b0), .ZN(_u10_u5_n3129 ));
NAND2_X1 _u10_u5_U1483  ( .A1(_u10_u5_n3129 ), .A2(_u10_u5_n2836 ), .ZN(_u10_u5_n2842 ) );
INV_X1 _u10_u5_U1482  ( .A(_u10_u5_n2842 ), .ZN(_u10_u5_n2833 ) );
NAND2_X1 _u10_u5_U1481  ( .A1(_u10_u5_n2833 ), .A2(_u10_u5_n2600 ), .ZN(_u10_u5_n2853 ) );
INV_X1 _u10_u5_U1480  ( .A(_u10_u5_n2853 ), .ZN(_u10_u5_n2082 ) );
NAND2_X1 _u10_u5_U1479  ( .A1(_u10_u5_n2082 ), .A2(_u10_u5_n2031 ), .ZN(_u10_u5_n2274 ) );
INV_X1 _u10_u5_U1478  ( .A(_u10_u5_n2274 ), .ZN(_u10_u5_n2669 ) );
NAND3_X1 _u10_u5_U1477  ( .A1(_u10_u5_n2668 ), .A2(_u10_u5_n2113 ), .A3(_u10_u5_n2669 ), .ZN(_u10_u5_n1858 ) );
INV_X1 _u10_u5_U1476  ( .A(_u10_u5_n1858 ), .ZN(_u10_u5_n3067 ) );
NAND2_X1 _u10_u5_U1475  ( .A1(_u10_u5_n3067 ), .A2(1'b0), .ZN(_u10_u5_n2092 ) );
INV_X1 _u10_u5_U1474  ( .A(_u10_u5_n2092 ), .ZN(_u10_u5_n3294 ) );
INV_X1 _u10_u5_U1473  ( .A(1'b0), .ZN(_u10_u5_n2446 ) );
INV_X1 _u10_u5_U1472  ( .A(1'b0), .ZN(_u10_u5_n2996 ) );
NAND2_X1 _u10_u5_U1471  ( .A1(_u10_u5_n3067 ), .A2(_u10_u5_n2996 ), .ZN(_u10_u5_n1847 ) );
NOR3_X1 _u10_u5_U1470  ( .A1(_u10_u5_n2446 ), .A2(1'b0), .A3(_u10_u5_n1847 ),.ZN(_u10_u5_n3413 ) );
NOR4_X1 _u10_u5_U1469  ( .A1(_u10_u5_n2875 ), .A2(_u10_u5_n3180 ), .A3(_u10_u5_n3294 ), .A4(_u10_u5_n3413 ), .ZN(_u10_u5_n3412 ) );
NAND4_X1 _u10_u5_U1468  ( .A1(_u10_u5_n3410 ), .A2(_u10_u5_n3411 ), .A3(_u10_u5_n3145 ), .A4(_u10_u5_n3412 ), .ZN(_u10_u5_n3409 ) );
NAND2_X1 _u10_u5_U1467  ( .A1(_u10_u5_n2461 ), .A2(_u10_u5_n3409 ), .ZN(_u10_u5_n3380 ) );
NOR2_X1 _u10_u5_U1466  ( .A1(_u10_u5_n1817 ), .A2(_u10_u5_n1816 ), .ZN(_u10_u5_n3368 ) );
AND2_X1 _u10_u5_U1465  ( .A1(_u10_u5_n3368 ), .A2(_u10_u5_n1813 ), .ZN(_u10_u5_n3320 ) );
NOR2_X1 _u10_u5_U1464  ( .A1(_u10_SYNOPSYS_UNCONNECTED_22 ), .A2(_u10_u5_n1815 ), .ZN(_u10_u5_n3236 ) );
NAND2_X1 _u10_u5_U1463  ( .A1(_u10_u5_n3320 ), .A2(_u10_u5_n3236 ), .ZN(_u10_u5_n2607 ) );
INV_X1 _u10_u5_U1462  ( .A(_u10_u5_n2607 ), .ZN(_u10_u5_n1966 ) );
INV_X1 _u10_u5_U1461  ( .A(_u10_u5_n2200 ), .ZN(_u10_u5_n3216 ) );
NAND2_X1 _u10_u5_U1460  ( .A1(1'b0), .A2(_u10_u5_n3216 ), .ZN(_u10_u5_n2367 ) );
INV_X1 _u10_u5_U1459  ( .A(_u10_u5_n2367 ), .ZN(_u10_u5_n3183 ) );
NAND2_X1 _u10_u5_U1458  ( .A1(_u10_u5_n3183 ), .A2(_u10_u5_n2195 ), .ZN(_u10_u5_n2194 ) );
INV_X1 _u10_u5_U1457  ( .A(_u10_u5_n2194 ), .ZN(_u10_u5_n2055 ) );
NAND2_X1 _u10_u5_U1456  ( .A1(_u10_u5_n2055 ), .A2(_u10_u5_n1853 ), .ZN(_u10_u5_n3401 ) );
INV_X1 _u10_u5_U1455  ( .A(_u10_u5_n2531 ), .ZN(_u10_u5_n2190 ) );
INV_X1 _u10_u5_U1454  ( .A(1'b0), .ZN(_u10_u5_n3001 ) );
NAND2_X1 _u10_u5_U1453  ( .A1(_u10_u5_n3001 ), .A2(_u10_u5_n2466 ), .ZN(_u10_u5_n2156 ) );
NOR2_X1 _u10_u5_U1452  ( .A1(_u10_u5_n2166 ), .A2(_u10_u5_n2596 ), .ZN(_u10_u5_n2594 ) );
NAND2_X1 _u10_u5_U1451  ( .A1(_u10_u5_n2594 ), .A2(_u10_u5_n2031 ), .ZN(_u10_u5_n2752 ) );
INV_X1 _u10_u5_U1450  ( .A(_u10_u5_n2752 ), .ZN(_u10_u5_n2421 ) );
NAND2_X1 _u10_u5_U1449  ( .A1(_u10_u5_n2421 ), .A2(_u10_u5_n2874 ), .ZN(_u10_u5_n2033 ) );
INV_X1 _u10_u5_U1448  ( .A(_u10_u5_n2033 ), .ZN(_u10_u5_n2742 ) );
NAND3_X1 _u10_u5_U1447  ( .A1(_u10_u5_n2305 ), .A2(_u10_u5_n1936 ), .A3(_u10_u5_n2742 ), .ZN(_u10_u5_n1896 ) );
OR3_X1 _u10_u5_U1446  ( .A1(_u10_u5_n2156 ), .A2(1'b0), .A3(_u10_u5_n1896 ),.ZN(_u10_u5_n2905 ) );
NAND2_X1 _u10_u5_U1445  ( .A1(_u10_u5_n2113 ), .A2(_u10_u5_n2996 ), .ZN(_u10_u5_n2719 ) );
NOR2_X1 _u10_u5_U1444  ( .A1(_u10_u5_n2719 ), .A2(1'b0), .ZN(_u10_u5_n2941 ));
INV_X1 _u10_u5_U1443  ( .A(_u10_u5_n2941 ), .ZN(_u10_u5_n2911 ) );
NOR2_X1 _u10_u5_U1442  ( .A1(_u10_u5_n2905 ), .A2(_u10_u5_n2911 ), .ZN(_u10_u5_n3222 ) );
INV_X1 _u10_u5_U1441  ( .A(_u10_u5_n3222 ), .ZN(_u10_u5_n2695 ) );
INV_X1 _u10_u5_U1440  ( .A(_u10_u5_n2156 ), .ZN(_u10_u5_n2089 ) );
NAND3_X1 _u10_u5_U1439  ( .A1(_u10_u5_n2089 ), .A2(_u10_u5_n2446 ), .A3(_u10_u5_n3180 ), .ZN(_u10_u5_n2902 ) );
NOR2_X1 _u10_u5_U1438  ( .A1(_u10_u5_n2902 ), .A2(_u10_u5_n2911 ), .ZN(_u10_u5_n2533 ) );
INV_X1 _u10_u5_U1437  ( .A(_u10_u5_n2533 ), .ZN(_u10_u5_n2485 ) );
NAND2_X1 _u10_u5_U1436  ( .A1(_u10_u5_n2695 ), .A2(_u10_u5_n2485 ), .ZN(_u10_u5_n2721 ) );
NAND2_X1 _u10_u5_U1435  ( .A1(1'b0), .A2(_u10_u5_n2113 ), .ZN(_u10_u5_n1868 ) );
INV_X1 _u10_u5_U1434  ( .A(_u10_u5_n1868 ), .ZN(_u10_u5_n2534 ) );
NOR2_X1 _u10_u5_U1433  ( .A1(_u10_u5_n2721 ), .A2(_u10_u5_n2534 ), .ZN(_u10_u5_n3231 ) );
NAND2_X1 _u10_u5_U1432  ( .A1(_u10_u5_n2467 ), .A2(_u10_u5_n3001 ), .ZN(_u10_u5_n2303 ) );
INV_X1 _u10_u5_U1431  ( .A(_u10_u5_n2303 ), .ZN(_u10_u5_n2549 ) );
INV_X1 _u10_u5_U1430  ( .A(1'b0), .ZN(_u10_u5_n2803 ) );
NAND2_X1 _u10_u5_U1429  ( .A1(_u10_u5_n2803 ), .A2(_u10_u5_n2446 ), .ZN(_u10_u5_n1846 ) );
INV_X1 _u10_u5_U1428  ( .A(_u10_u5_n1846 ), .ZN(_u10_u5_n2667 ) );
NAND3_X1 _u10_u5_U1427  ( .A1(_u10_u5_n2549 ), .A2(_u10_u5_n2667 ), .A3(1'b0), .ZN(_u10_u5_n2739 ) );
INV_X1 _u10_u5_U1426  ( .A(_u10_u5_n2739 ), .ZN(_u10_u5_n3272 ) );
INV_X1 _u10_u5_U1425  ( .A(_u10_u5_n2719 ), .ZN(_u10_u5_n2364 ) );
NAND2_X1 _u10_u5_U1424  ( .A1(_u10_u5_n3272 ), .A2(_u10_u5_n2364 ), .ZN(_u10_u5_n2852 ) );
INV_X1 _u10_u5_U1423  ( .A(_u10_u5_n2852 ), .ZN(_u10_u5_n2214 ) );
NAND2_X1 _u10_u5_U1422  ( .A1(_u10_u5_n2875 ), .A2(_u10_u5_n2089 ), .ZN(_u10_u5_n2097 ) );
INV_X1 _u10_u5_U1421  ( .A(_u10_u5_n2097 ), .ZN(_u10_u5_n2300 ) );
NAND2_X1 _u10_u5_U1420  ( .A1(_u10_u5_n2300 ), .A2(_u10_u5_n2446 ), .ZN(_u10_u5_n2001 ) );
NOR2_X1 _u10_u5_U1419  ( .A1(_u10_u5_n2001 ), .A2(_u10_u5_n2911 ), .ZN(_u10_u5_n2877 ) );
NOR2_X1 _u10_u5_U1418  ( .A1(_u10_u5_n2214 ), .A2(_u10_u5_n2877 ), .ZN(_u10_u5_n2940 ) );
NAND2_X1 _u10_u5_U1417  ( .A1(_u10_u5_n3231 ), .A2(_u10_u5_n2940 ), .ZN(_u10_u5_n3408 ) );
NAND2_X1 _u10_u5_U1416  ( .A1(_u10_u5_n2190 ), .A2(_u10_u5_n3408 ), .ZN(_u10_u5_n3402 ) );
NOR2_X1 _u10_u5_U1415  ( .A1(_u10_u5_n2446 ), .A2(_u10_u5_n2911 ), .ZN(_u10_u5_n3059 ) );
NAND2_X1 _u10_u5_U1414  ( .A1(_u10_u5_n3059 ), .A2(_u10_u5_n2190 ), .ZN(_u10_u5_n3404 ) );
AND3_X1 _u10_u5_U1413  ( .A1(_u10_u5_n3407 ), .A2(_u10_u5_n3226 ), .A3(_u10_u5_n3115 ), .ZN(_u10_u5_n3058 ) );
NAND2_X1 _u10_u5_U1412  ( .A1(_u10_u5_n3058 ), .A2(_u10_u5_n2022 ), .ZN(_u10_u5_n3406 ) );
NAND2_X1 _u10_u5_U1411  ( .A1(_u10_u5_n1853 ), .A2(_u10_u5_n3406 ), .ZN(_u10_u5_n3405 ) );
AND3_X1 _u10_u5_U1410  ( .A1(_u10_u5_n3404 ), .A2(_u10_u5_n1965 ), .A3(_u10_u5_n3405 ), .ZN(_u10_u5_n3063 ) );
NAND2_X1 _u10_u5_U1409  ( .A1(_u10_u5_n2667 ), .A2(_u10_u5_n3001 ), .ZN(_u10_u5_n1898 ) );
INV_X1 _u10_u5_U1408  ( .A(_u10_u5_n1898 ), .ZN(_u10_u5_n2835 ) );
NAND3_X1 _u10_u5_U1407  ( .A1(_u10_u5_n2364 ), .A2(_u10_u5_n2835 ), .A3(1'b0), .ZN(_u10_u5_n1869 ) );
NOR2_X1 _u10_u5_U1406  ( .A1(_u10_u5_n1869 ), .A2(_u10_u5_n2531 ), .ZN(_u10_u5_n2761 ) );
NOR3_X1 _u10_u5_U1405  ( .A1(_u10_u5_n2761 ), .A2(_u10_u5_n2528 ), .A3(_u10_u5_n2054 ), .ZN(_u10_u5_n3403 ) );
NAND4_X1 _u10_u5_U1404  ( .A1(_u10_u5_n3401 ), .A2(_u10_u5_n3402 ), .A3(_u10_u5_n3063 ), .A4(_u10_u5_n3403 ), .ZN(_u10_u5_n3400 ) );
NAND2_X1 _u10_u5_U1403  ( .A1(_u10_u5_n1966 ), .A2(_u10_u5_n3400 ), .ZN(_u10_u5_n3381 ) );
AND2_X1 _u10_u5_U1402  ( .A1(_u10_u5_n3368 ), .A2(_u10_SYNOPSYS_UNCONNECTED_23 ), .ZN(_u10_u5_n3319 ) );
NAND2_X1 _u10_u5_U1401  ( .A1(_u10_u5_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_22 ), .ZN(_u10_u5_n1849 ) );
INV_X1 _u10_u5_U1400  ( .A(_u10_u5_n1849 ), .ZN(_u10_u5_n2183 ) );
NAND2_X1 _u10_u5_U1399  ( .A1(_u10_u5_n2884 ), .A2(_u10_u5_n2183 ), .ZN(_u10_u5_n2883 ) );
INV_X1 _u10_u5_U1398  ( .A(_u10_u5_n2883 ), .ZN(_u10_u5_n1890 ) );
INV_X1 _u10_u5_U1397  ( .A(_u10_u5_n2940 ), .ZN(_u10_u5_n3278 ) );
NAND2_X1 _u10_u5_U1396  ( .A1(_u10_u5_n1890 ), .A2(_u10_u5_n3278 ), .ZN(_u10_u5_n3382 ) );
NAND2_X1 _u10_u5_U1395  ( .A1(_u10_u5_n3059 ), .A2(_u10_u5_n2669 ), .ZN(_u10_u5_n3399 ) );
NAND2_X1 _u10_u5_U1394  ( .A1(_u10_u5_n2031 ), .A2(_u10_u5_n3399 ), .ZN(_u10_u5_n3398 ) );
NAND2_X1 _u10_u5_U1393  ( .A1(_u10_u5_n2162 ), .A2(_u10_u5_n3398 ), .ZN(_u10_u5_n3395 ) );
NAND3_X1 _u10_u5_U1392  ( .A1(_u10_u5_n2747 ), .A2(_u10_u5_n2078 ), .A3(_u10_u5_n3126 ), .ZN(_u10_u5_n3396 ) );
NAND2_X1 _u10_u5_U1391  ( .A1(_u10_u5_n2055 ), .A2(_u10_u5_n2036 ), .ZN(_u10_u5_n2285 ) );
NOR2_X1 _u10_u5_U1390  ( .A1(_u10_u5_n2285 ), .A2(_u10_u5_n2030 ), .ZN(_u10_u5_n3349 ) );
INV_X1 _u10_u5_U1389  ( .A(_u10_u5_n3349 ), .ZN(_u10_u5_n1933 ) );
INV_X1 _u10_u5_U1388  ( .A(_u10_u5_n2710 ), .ZN(_u10_u5_n3397 ) );
NAND4_X1 _u10_u5_U1387  ( .A1(_u10_u5_n3395 ), .A2(_u10_u5_n3396 ), .A3(_u10_u5_n1933 ), .A4(_u10_u5_n3397 ), .ZN(_u10_u5_n3389 ) );
NAND2_X1 _u10_u5_U1386  ( .A1(_u10_u5_n1936 ), .A2(_u10_u5_n2828 ), .ZN(_u10_u5_n3141 ) );
INV_X1 _u10_u5_U1385  ( .A(_u10_u5_n3141 ), .ZN(_u10_u5_n2302 ) );
NAND2_X1 _u10_u5_U1384  ( .A1(_u10_u5_n3394 ), .A2(_u10_u5_n2302 ), .ZN(_u10_u5_n3390 ) );
NOR2_X1 _u10_u5_U1383  ( .A1(_u10_u5_n1869 ), .A2(_u10_u5_n2274 ), .ZN(_u10_u5_n3378 ) );
INV_X1 _u10_u5_U1382  ( .A(_u10_u5_n3378 ), .ZN(_u10_u5_n2748 ) );
NOR2_X1 _u10_u5_U1381  ( .A1(1'b0), .A2(_u10_u5_n2748 ), .ZN(_u10_u5_n3391 ));
NAND2_X1 _u10_u5_U1380  ( .A1(_u10_u5_n2534 ), .A2(_u10_u5_n2669 ), .ZN(_u10_u5_n2383 ) );
INV_X1 _u10_u5_U1379  ( .A(_u10_u5_n2383 ), .ZN(_u10_u5_n1978 ) );
NAND2_X1 _u10_u5_U1378  ( .A1(_u10_u5_n1978 ), .A2(_u10_u5_n2874 ), .ZN(_u10_u5_n3392 ) );
INV_X1 _u10_u5_U1377  ( .A(_u10_u5_n2411 ), .ZN(_u10_u5_n2164 ) );
NAND4_X1 _u10_u5_U1376  ( .A1(_u10_u5_n3392 ), .A2(_u10_u5_n3393 ), .A3(_u10_u5_n2033 ), .A4(_u10_u5_n2164 ), .ZN(_u10_u5_n2476 ) );
NOR4_X1 _u10_u5_U1375  ( .A1(_u10_u5_n3389 ), .A2(_u10_u5_n3390 ), .A3(_u10_u5_n3391 ), .A4(_u10_u5_n2476 ), .ZN(_u10_u5_n3388 ) );
NAND2_X1 _u10_u5_U1374  ( .A1(_u10_u5_n3236 ), .A2(_u10_u5_n3328 ), .ZN(_u10_u5_n2025 ) );
NOR2_X1 _u10_u5_U1373  ( .A1(_u10_u5_n3388 ), .A2(_u10_u5_n2025 ), .ZN(_u10_u5_n3384 ) );
NOR2_X1 _u10_u5_U1372  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u5_n2152 ) );
NAND2_X1 _u10_u5_U1371  ( .A1(_u10_u5_n2152 ), .A2(_u10_u5_n2175 ), .ZN(_u10_u5_n2722 ) );
INV_X1 _u10_u5_U1370  ( .A(_u10_u5_n2722 ), .ZN(_u10_u5_n2588 ) );
NAND2_X1 _u10_u5_U1369  ( .A1(_u10_u5_n2549 ), .A2(_u10_u5_n3349 ), .ZN(_u10_u5_n2091 ) );
NOR2_X1 _u10_u5_U1368  ( .A1(_u10_u5_n2091 ), .A2(_u10_u5_n1846 ), .ZN(_u10_u5_n2128 ) );
NAND3_X1 _u10_u5_U1367  ( .A1(_u10_u5_n3066 ), .A2(_u10_u5_n2113 ), .A3(_u10_u5_n2128 ), .ZN(_u10_u5_n2342 ) );
INV_X1 _u10_u5_U1366  ( .A(_u10_u5_n2342 ), .ZN(_u10_u5_n3316 ) );
NAND2_X1 _u10_u5_U1365  ( .A1(_u10_u5_n2588 ), .A2(_u10_u5_n3316 ), .ZN(_u10_u5_n2142 ) );
NOR2_X1 _u10_u5_U1364  ( .A1(_u10_u5_n1954 ), .A2(_u10_u5_n1898 ), .ZN(_u10_u5_n2255 ) );
NAND2_X1 _u10_u5_U1363  ( .A1(_u10_u5_n2255 ), .A2(_u10_u5_n2996 ), .ZN(_u10_u5_n1915 ) );
INV_X1 _u10_u5_U1362  ( .A(_u10_u5_n1915 ), .ZN(_u10_u5_n2251 ) );
NAND2_X1 _u10_u5_U1361  ( .A1(_u10_u5_n2251 ), .A2(_u10_u5_n2113 ), .ZN(_u10_u5_n1925 ) );
INV_X1 _u10_u5_U1360  ( .A(_u10_u5_n2026 ), .ZN(_u10_u5_n3340 ) );
NOR3_X1 _u10_u5_U1359  ( .A1(_u10_u5_n1925 ), .A2(_u10_u5_n2216 ), .A3(_u10_u5_n3340 ), .ZN(_u10_u5_n2003 ) );
INV_X1 _u10_u5_U1358  ( .A(1'b0), .ZN(_u10_u5_n1930 ) );
NAND2_X1 _u10_u5_U1357  ( .A1(_u10_u5_n2003 ), .A2(_u10_u5_n1930 ), .ZN(_u10_u5_n3387 ) );
AND2_X1 _u10_u5_U1356  ( .A1(_u10_u5_n2142 ), .A2(_u10_u5_n3387 ), .ZN(_u10_u5_n3366 ) );
NOR3_X1 _u10_u5_U1355  ( .A1(_u10_u5_n1813 ), .A2(_u10_u5_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_19 ), .ZN(_u10_u5_n3360 ) );
NOR2_X1 _u10_u5_U1354  ( .A1(_u10_SYNOPSYS_UNCONNECTED_21 ), .A2(_u10_SYNOPSYS_UNCONNECTED_22 ), .ZN(_u10_u5_n3136 ) );
NAND2_X1 _u10_u5_U1353  ( .A1(_u10_u5_n3360 ), .A2(_u10_u5_n3136 ), .ZN(_u10_u5_n2344 ) );
NOR2_X1 _u10_u5_U1352  ( .A1(_u10_u5_n3366 ), .A2(_u10_u5_n2344 ), .ZN(_u10_u5_n3385 ) );
NOR3_X1 _u10_u5_U1351  ( .A1(_u10_SYNOPSYS_UNCONNECTED_19 ), .A2(_u10_u5_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_23 ), .ZN(_u10_u5_n3342 ) );
NAND2_X1 _u10_u5_U1350  ( .A1(_u10_u5_n3342 ), .A2(_u10_u5_n3136 ), .ZN(_u10_u5_n2584 ) );
NOR2_X1 _u10_u5_U1349  ( .A1(_u10_u5_n2584 ), .A2(1'b0), .ZN(_u10_u5_n2139 ));
INV_X1 _u10_u5_U1348  ( .A(_u10_u5_n2216 ), .ZN(_u10_u5_n2106 ) );
AND2_X1 _u10_u5_U1347  ( .A1(_u10_u5_n2152 ), .A2(_u10_u5_n2106 ), .ZN(_u10_u5_n2336 ) );
NAND2_X1 _u10_u5_U1346  ( .A1(_u10_u5_n2139 ), .A2(_u10_u5_n2336 ), .ZN(_u10_u5_n2365 ) );
INV_X1 _u10_u5_U1345  ( .A(_u10_u5_n2365 ), .ZN(_u10_u5_n2004 ) );
AND2_X1 _u10_u5_U1344  ( .A1(_u10_u5_n2877 ), .A2(_u10_u5_n2004 ), .ZN(_u10_u5_n3386 ) );
NOR3_X1 _u10_u5_U1343  ( .A1(_u10_u5_n3384 ), .A2(_u10_u5_n3385 ), .A3(_u10_u5_n3386 ), .ZN(_u10_u5_n3383 ) );
NAND4_X1 _u10_u5_U1342  ( .A1(_u10_u5_n3380 ), .A2(_u10_u5_n3381 ), .A3(_u10_u5_n3382 ), .A4(_u10_u5_n3383 ), .ZN(_u10_u5_n3191 ) );
NAND2_X1 _u10_u5_U1341  ( .A1(_u10_u5_n2285 ), .A2(_u10_u5_n3379 ), .ZN(_u10_u5_n1975 ) );
NOR3_X1 _u10_u5_U1340  ( .A1(_u10_u5_n3378 ), .A2(1'b0), .A3(_u10_u5_n1975 ),.ZN(_u10_u5_n3122 ) );
AND4_X1 _u10_u5_U1339  ( .A1(_u10_u5_n2752 ), .A2(_u10_u5_n2383 ), .A3(_u10_u5_n1969 ), .A4(_u10_u5_n3122 ), .ZN(_u10_u5_n3377 ) );
NOR2_X1 _u10_u5_U1338  ( .A1(_u10_u5_n1814 ), .A2(_u10_u5_n1815 ), .ZN(_u10_u5_n3147 ) );
NAND2_X1 _u10_u5_U1337  ( .A1(_u10_u5_n3328 ), .A2(_u10_u5_n3147 ), .ZN(_u10_u5_n2359 ) );
NOR2_X1 _u10_u5_U1336  ( .A1(_u10_u5_n3377 ), .A2(_u10_u5_n2359 ), .ZN(_u10_u5_n3362 ) );
INV_X1 _u10_u5_U1335  ( .A(_u10_u5_n2008 ), .ZN(_u10_u5_n3097 ) );
NOR3_X1 _u10_u5_U1334  ( .A1(_u10_SYNOPSYS_UNCONNECTED_19 ), .A2(_u10_u5_n1813 ), .A3(_u10_SYNOPSYS_UNCONNECTED_20 ), .ZN(_u10_u5_n3269 ) );
NAND2_X1 _u10_u5_U1333  ( .A1(_u10_u5_n3269 ), .A2(_u10_u5_n3136 ), .ZN(_u10_u5_n3109 ) );
INV_X1 _u10_u5_U1332  ( .A(_u10_u5_n3109 ), .ZN(_u10_u5_n2999 ) );
INV_X1 _u10_u5_U1331  ( .A(_u10_u5_n2508 ), .ZN(_u10_u5_n2103 ) );
NAND2_X1 _u10_u5_U1330  ( .A1(_u10_u5_n2336 ), .A2(_u10_u5_n2103 ), .ZN(_u10_u5_n2249 ) );
NOR2_X1 _u10_u5_U1329  ( .A1(_u10_u5_n2249 ), .A2(1'b0), .ZN(_u10_u5_n1866 ));
NAND2_X1 _u10_u5_U1328  ( .A1(_u10_u5_n1866 ), .A2(_u10_u5_n1922 ), .ZN(_u10_u5_n2632 ) );
INV_X1 _u10_u5_U1327  ( .A(_u10_u5_n2223 ), .ZN(_u10_u5_n1918 ) );
NOR2_X1 _u10_u5_U1326  ( .A1(_u10_u5_n2632 ), .A2(_u10_u5_n1918 ), .ZN(_u10_u5_n1981 ) );
NAND3_X1 _u10_u5_U1325  ( .A1(_u10_u5_n3097 ), .A2(_u10_u5_n2999 ), .A3(_u10_u5_n1981 ), .ZN(_u10_u5_n3034 ) );
NOR3_X1 _u10_u5_U1324  ( .A1(_u10_SYNOPSYS_UNCONNECTED_20 ), .A2(_u10_SYNOPSYS_UNCONNECTED_19 ), .A3(_u10_SYNOPSYS_UNCONNECTED_23 ),.ZN(_u10_u5_n3302 ) );
NAND2_X1 _u10_u5_U1323  ( .A1(_u10_u5_n3302 ), .A2(_u10_u5_n3174 ), .ZN(_u10_u5_n3162 ) );
INV_X1 _u10_u5_U1322  ( .A(_u10_u5_n3162 ), .ZN(_u10_u5_n2979 ) );
NAND2_X1 _u10_u5_U1321  ( .A1(_u10_u5_n2979 ), .A2(_u10_u5_n2972 ), .ZN(_u10_u5_n1984 ) );
AND2_X1 _u10_u5_U1320  ( .A1(_u10_u5_n3302 ), .A2(_u10_u5_n3136 ), .ZN(_u10_u5_n2977 ) );
NAND3_X1 _u10_u5_U1319  ( .A1(_u10_u5_n2977 ), .A2(_u10_u5_n3000 ), .A3(_u10_u5_n3097 ), .ZN(_u10_u5_n3376 ) );
NAND2_X1 _u10_u5_U1318  ( .A1(_u10_u5_n1984 ), .A2(_u10_u5_n3376 ), .ZN(_u10_u5_n3375 ) );
NAND2_X1 _u10_u5_U1317  ( .A1(_u10_u5_n1981 ), .A2(_u10_u5_n3375 ), .ZN(_u10_u5_n2798 ) );
NAND2_X1 _u10_u5_U1316  ( .A1(_u10_u5_n3034 ), .A2(_u10_u5_n2798 ), .ZN(_u10_u5_n2007 ) );
NAND2_X1 _u10_u5_U1315  ( .A1(_u10_u5_n3269 ), .A2(_u10_u5_n3147 ), .ZN(_u10_u5_n2102 ) );
NOR2_X1 _u10_u5_U1314  ( .A1(_u10_u5_n2249 ), .A2(_u10_u5_n2102 ), .ZN(_u10_u5_n3323 ) );
INV_X1 _u10_u5_U1313  ( .A(_u10_u5_n3323 ), .ZN(_u10_u5_n3374 ) );
INV_X1 _u10_u5_U1312  ( .A(_u10_u5_n2344 ), .ZN(_u10_u5_n2002 ) );
NAND2_X1 _u10_u5_U1311  ( .A1(_u10_u5_n2336 ), .A2(_u10_u5_n2002 ), .ZN(_u10_u5_n3225 ) );
NAND2_X1 _u10_u5_U1310  ( .A1(_u10_u5_n3374 ), .A2(_u10_u5_n3225 ), .ZN(_u10_u5_n2488 ) );
NAND2_X1 _u10_u5_U1309  ( .A1(_u10_u5_n3342 ), .A2(_u10_u5_n3236 ), .ZN(_u10_u5_n2253 ) );
NOR2_X1 _u10_u5_U1308  ( .A1(_u10_u5_n2253 ), .A2(1'b0), .ZN(_u10_u5_n1885 ));
NAND2_X1 _u10_u5_U1307  ( .A1(_u10_u5_n3360 ), .A2(_u10_u5_n3174 ), .ZN(_u10_u5_n2254 ) );
INV_X1 _u10_u5_U1306  ( .A(_u10_u5_n2254 ), .ZN(_u10_u5_n2986 ) );
NAND2_X1 _u10_u5_U1305  ( .A1(_u10_u5_n2106 ), .A2(_u10_u5_n2986 ), .ZN(_u10_u5_n1913 ) );
INV_X1 _u10_u5_U1304  ( .A(_u10_u5_n1913 ), .ZN(_u10_u5_n2377 ) );
OR4_X1 _u10_u5_U1303  ( .A1(_u10_u5_n2007 ), .A2(_u10_u5_n2488 ), .A3(_u10_u5_n1885 ), .A4(_u10_u5_n2377 ), .ZN(_u10_u5_n3373 ) );
NAND2_X1 _u10_u5_U1302  ( .A1(_u10_u5_n2534 ), .A2(_u10_u5_n3373 ), .ZN(_u10_u5_n3370 ) );
NAND2_X1 _u10_u5_U1301  ( .A1(_u10_u5_n3342 ), .A2(_u10_u5_n3174 ), .ZN(_u10_u5_n2037 ) );
NAND2_X1 _u10_u5_U1300  ( .A1(_u10_u5_n2037 ), .A2(_u10_u5_n2254 ), .ZN(_u10_u5_n3372 ) );
NAND2_X1 _u10_u5_U1299  ( .A1(_u10_u5_n2003 ), .A2(_u10_u5_n3372 ), .ZN(_u10_u5_n3371 ) );
NAND2_X1 _u10_u5_U1298  ( .A1(_u10_u5_n3370 ), .A2(_u10_u5_n3371 ), .ZN(_u10_u5_n3363 ) );
NOR2_X1 _u10_u5_U1297  ( .A1(_u10_u5_n2490 ), .A2(_u10_u5_n1961 ), .ZN(_u10_u5_n3369 ) );
NAND2_X1 _u10_u5_U1296  ( .A1(_u10_u5_n2534 ), .A2(_u10_u5_n2049 ), .ZN(_u10_u5_n2646 ) );
INV_X1 _u10_u5_U1295  ( .A(_u10_u5_n2646 ), .ZN(_u10_u5_n3055 ) );
NOR2_X1 _u10_u5_U1294  ( .A1(_u10_u5_n3369 ), .A2(_u10_u5_n3055 ), .ZN(_u10_u5_n3367 ) );
NAND2_X1 _u10_u5_U1293  ( .A1(_u10_u5_n3368 ), .A2(_u10_u5_n3147 ), .ZN(_u10_u5_n2495 ) );
NOR2_X1 _u10_u5_U1292  ( .A1(_u10_u5_n3367 ), .A2(_u10_u5_n2495 ), .ZN(_u10_u5_n3364 ) );
INV_X1 _u10_u5_U1291  ( .A(_u10_u5_n2139 ), .ZN(_u10_u5_n3254 ) );
NOR2_X1 _u10_u5_U1290  ( .A1(_u10_u5_n3366 ), .A2(_u10_u5_n3254 ), .ZN(_u10_u5_n3365 ) );
NOR4_X1 _u10_u5_U1289  ( .A1(_u10_u5_n3362 ), .A2(_u10_u5_n3363 ), .A3(_u10_u5_n3364 ), .A4(_u10_u5_n3365 ), .ZN(_u10_u5_n3305 ) );
NAND2_X1 _u10_u5_U1288  ( .A1(_u10_u5_n3302 ), .A2(_u10_u5_n3147 ), .ZN(_u10_u5_n2980 ) );
NAND2_X1 _u10_u5_U1287  ( .A1(_u10_u5_n2102 ), .A2(_u10_u5_n2980 ), .ZN(_u10_u5_n2177 ) );
NAND2_X1 _u10_u5_U1286  ( .A1(_u10_u5_n2003 ), .A2(_u10_u5_n2493 ), .ZN(_u10_u5_n1962 ) );
NAND2_X1 _u10_u5_U1285  ( .A1(_u10_u5_n1961 ), .A2(_u10_u5_n1962 ), .ZN(_u10_u5_n3361 ) );
NAND2_X1 _u10_u5_U1284  ( .A1(_u10_u5_n2177 ), .A2(_u10_u5_n3361 ), .ZN(_u10_u5_n3357 ) );
NAND2_X1 _u10_u5_U1283  ( .A1(_u10_u5_n3236 ), .A2(_u10_u5_n3360 ), .ZN(_u10_u5_n1859 ) );
INV_X1 _u10_u5_U1282  ( .A(_u10_u5_n1859 ), .ZN(_u10_u5_n2256 ) );
NAND3_X1 _u10_u5_U1281  ( .A1(_u10_u5_n2256 ), .A2(_u10_u5_n2113 ), .A3(_u10_u5_n2128 ), .ZN(_u10_u5_n3358 ) );
NOR2_X1 _u10_u5_U1280  ( .A1(_u10_u5_n2877 ), .A2(_u10_u5_n3222 ), .ZN(_u10_u5_n3347 ) );
NAND2_X1 _u10_u5_U1279  ( .A1(_u10_u5_n3347 ), .A2(_u10_u5_n1869 ), .ZN(_u10_u5_n2005 ) );
NAND2_X1 _u10_u5_U1278  ( .A1(_u10_u5_n2488 ), .A2(_u10_u5_n2005 ), .ZN(_u10_u5_n3359 ) );
NAND3_X1 _u10_u5_U1277  ( .A1(_u10_u5_n3357 ), .A2(_u10_u5_n3358 ), .A3(_u10_u5_n3359 ), .ZN(_u10_u5_n3352 ) );
NAND2_X1 _u10_u5_U1276  ( .A1(_u10_u5_n3320 ), .A2(_u10_u5_n3136 ), .ZN(_u10_u5_n2356 ) );
INV_X1 _u10_u5_U1275  ( .A(_u10_u5_n2356 ), .ZN(_u10_u5_n2830 ) );
NAND2_X1 _u10_u5_U1274  ( .A1(_u10_u5_n2830 ), .A2(_u10_u5_n2836 ), .ZN(_u10_u5_n2291 ) );
NOR3_X1 _u10_u5_U1273  ( .A1(_u10_u5_n2291 ), .A2(_u10_u5_n2330 ), .A3(_u10_u5_n2022 ), .ZN(_u10_u5_n3353 ) );
INV_X1 _u10_u5_U1272  ( .A(_u10_u5_n1925 ), .ZN(_u10_u5_n2105 ) );
AND2_X1 _u10_u5_U1271  ( .A1(_u10_u5_n2108 ), .A2(_u10_u5_n2105 ), .ZN(_u10_u5_n2915 ) );
INV_X1 _u10_u5_U1270  ( .A(_u10_u5_n2330 ), .ZN(_u10_u5_n2107 ) );
NAND2_X1 _u10_u5_U1269  ( .A1(_u10_u5_n2915 ), .A2(_u10_u5_n2107 ), .ZN(_u10_u5_n2203 ) );
INV_X1 _u10_u5_U1268  ( .A(_u10_u5_n2203 ), .ZN(_u10_u5_n1982 ) );
NAND2_X1 _u10_u5_U1267  ( .A1(_u10_u5_n1982 ), .A2(_u10_u5_n2536 ), .ZN(_u10_u5_n2587 ) );
INV_X1 _u10_u5_U1266  ( .A(_u10_u5_n2587 ), .ZN(_u10_u5_n2697 ) );
NAND3_X1 _u10_u5_U1265  ( .A1(_u10_u5_n2697 ), .A2(_u10_u5_n2493 ), .A3(_u10_u5_n2377 ), .ZN(_u10_u5_n2412 ) );
INV_X1 _u10_u5_U1264  ( .A(_u10_u5_n2412 ), .ZN(_u10_u5_n3354 ) );
NAND2_X1 _u10_u5_U1263  ( .A1(_u10_u5_n3174 ), .A2(_u10_u5_n3269 ), .ZN(_u10_u5_n2375 ) );
INV_X1 _u10_u5_U1262  ( .A(_u10_u5_n2375 ), .ZN(_u10_u5_n2507 ) );
NAND2_X1 _u10_u5_U1261  ( .A1(_u10_u5_n1981 ), .A2(_u10_u5_n2507 ), .ZN(_u10_u5_n2621 ) );
NOR4_X1 _u10_u5_U1260  ( .A1(1'b0), .A2(_u10_u5_n3356 ), .A3(_u10_u5_n2203 ),.A4(_u10_u5_n2621 ), .ZN(_u10_u5_n3355 ) );
NOR4_X1 _u10_u5_U1259  ( .A1(_u10_u5_n3352 ), .A2(_u10_u5_n3353 ), .A3(_u10_u5_n3354 ), .A4(_u10_u5_n3355 ), .ZN(_u10_u5_n3306 ) );
NOR2_X1 _u10_u5_U1258  ( .A1(_u10_u5_n2842 ), .A2(_u10_u5_n2356 ), .ZN(_u10_u5_n1891 ) );
INV_X1 _u10_u5_U1257  ( .A(_u10_u5_n1869 ), .ZN(_u10_u5_n2885 ) );
NAND2_X1 _u10_u5_U1256  ( .A1(_u10_u5_n1891 ), .A2(_u10_u5_n2885 ), .ZN(_u10_u5_n3330 ) );
NAND2_X1 _u10_u5_U1255  ( .A1(_u10_u5_n2761 ), .A2(_u10_u5_n2837 ), .ZN(_u10_u5_n3351 ) );
NAND3_X1 _u10_u5_U1254  ( .A1(_u10_u5_n2884 ), .A2(_u10_u5_n2080 ), .A3(_u10_u5_n2915 ), .ZN(_u10_u5_n2762 ) );
NAND2_X1 _u10_u5_U1253  ( .A1(_u10_u5_n2055 ), .A2(_u10_u5_n2019 ), .ZN(_u10_u5_n3259 ) );
NAND4_X1 _u10_u5_U1252  ( .A1(_u10_u5_n3351 ), .A2(_u10_u5_n2762 ), .A3(_u10_u5_n2061 ), .A4(_u10_u5_n3259 ), .ZN(_u10_u5_n3350 ) );
NAND2_X1 _u10_u5_U1251  ( .A1(_u10_u5_n2183 ), .A2(_u10_u5_n3350 ), .ZN(_u10_u5_n3331 ) );
NAND2_X1 _u10_u5_U1250  ( .A1(_u10_u5_n3349 ), .A2(_u10_u5_n2305 ), .ZN(_u10_u5_n3348 ) );
NAND2_X1 _u10_u5_U1249  ( .A1(_u10_u5_n1896 ), .A2(_u10_u5_n3348 ), .ZN(_u10_u5_n3176 ) );
NAND2_X1 _u10_u5_U1248  ( .A1(_u10_u5_n2461 ), .A2(_u10_u5_n3176 ), .ZN(_u10_u5_n3332 ) );
INV_X1 _u10_u5_U1247  ( .A(_u10_u5_n2495 ), .ZN(_u10_u5_n2063 ) );
NAND2_X1 _u10_u5_U1246  ( .A1(_u10_u5_n2049 ), .A2(_u10_u5_n2063 ), .ZN(_u10_u5_n2886 ) );
NOR2_X1 _u10_u5_U1245  ( .A1(_u10_u5_n3347 ), .A2(_u10_u5_n2886 ), .ZN(_u10_u5_n3334 ) );
NAND2_X1 _u10_u5_U1244  ( .A1(1'b0), .A2(_u10_u5_n2835 ), .ZN(_u10_u5_n3344 ) );
NAND2_X1 _u10_u5_U1243  ( .A1(_u10_u5_n2001 ), .A2(_u10_u5_n2905 ), .ZN(_u10_u5_n3346 ) );
NAND2_X1 _u10_u5_U1242  ( .A1(_u10_u5_n3346 ), .A2(_u10_u5_n2803 ), .ZN(_u10_u5_n3345 ) );
NAND2_X1 _u10_u5_U1241  ( .A1(_u10_u5_n2087 ), .A2(_u10_u5_n2835 ), .ZN(_u10_u5_n2413 ) );
INV_X1 _u10_u5_U1240  ( .A(_u10_u5_n2128 ), .ZN(_u10_u5_n2235 ) );
NAND4_X1 _u10_u5_U1239  ( .A1(_u10_u5_n3344 ), .A2(_u10_u5_n3345 ), .A3(_u10_u5_n2413 ), .A4(_u10_u5_n2235 ), .ZN(_u10_u5_n3329 ) );
NOR2_X1 _u10_u5_U1238  ( .A1(_u10_u5_n1915 ), .A2(_u10_u5_n3340 ), .ZN(_u10_u5_n3343 ) );
NOR3_X1 _u10_u5_U1237  ( .A1(_u10_u5_n3329 ), .A2(1'b0), .A3(_u10_u5_n3343 ),.ZN(_u10_u5_n3341 ) );
NAND2_X1 _u10_u5_U1236  ( .A1(_u10_u5_n3342 ), .A2(_u10_u5_n3147 ), .ZN(_u10_u5_n2688 ) );
NOR2_X1 _u10_u5_U1235  ( .A1(_u10_u5_n3341 ), .A2(_u10_u5_n2688 ), .ZN(_u10_u5_n3335 ) );
NOR2_X1 _u10_u5_U1234  ( .A1(_u10_u5_n2256 ), .A2(_u10_u5_n1885 ), .ZN(_u10_u5_n2689 ) );
NOR2_X1 _u10_u5_U1233  ( .A1(1'b0), .A2(_u10_u5_n2413 ), .ZN(_u10_u5_n3338 ));
NOR2_X1 _u10_u5_U1232  ( .A1(_u10_u5_n1925 ), .A2(_u10_u5_n3340 ), .ZN(_u10_u5_n3339 ) );
NOR3_X1 _u10_u5_U1231  ( .A1(_u10_u5_n2005 ), .A2(_u10_u5_n3338 ), .A3(_u10_u5_n3339 ), .ZN(_u10_u5_n3337 ) );
NOR2_X1 _u10_u5_U1230  ( .A1(_u10_u5_n2689 ), .A2(_u10_u5_n3337 ), .ZN(_u10_u5_n3336 ) );
NOR3_X1 _u10_u5_U1229  ( .A1(_u10_u5_n3334 ), .A2(_u10_u5_n3335 ), .A3(_u10_u5_n3336 ), .ZN(_u10_u5_n3333 ) );
NAND4_X1 _u10_u5_U1228  ( .A1(_u10_u5_n3330 ), .A2(_u10_u5_n3331 ), .A3(_u10_u5_n3332 ), .A4(_u10_u5_n3333 ), .ZN(_u10_u5_n3308 ) );
NAND3_X1 _u10_u5_U1227  ( .A1(_u10_SYNOPSYS_UNCONNECTED_23 ), .A2(_u10_SYNOPSYS_UNCONNECTED_20 ), .A3(_u10_u5_n3147 ), .ZN(_u10_u5_n2126 ) );
INV_X1 _u10_u5_U1226  ( .A(_u10_u5_n2126 ), .ZN(_u10_u5_n2329 ) );
NAND2_X1 _u10_u5_U1225  ( .A1(_u10_u5_n2329 ), .A2(_u10_u5_n3329 ), .ZN(_u10_u5_n3324 ) );
NAND2_X1 _u10_u5_U1224  ( .A1(_u10_u5_n3328 ), .A2(_u10_u5_n3136 ), .ZN(_u10_u5_n2000 ) );
INV_X1 _u10_u5_U1223  ( .A(_u10_u5_n2000 ), .ZN(_u10_u5_n2445 ) );
NAND3_X1 _u10_u5_U1222  ( .A1(_u10_u5_n2446 ), .A2(_u10_u5_n3001 ), .A3(_u10_u5_n2087 ), .ZN(_u10_u5_n3327 ) );
NAND2_X1 _u10_u5_U1221  ( .A1(_u10_u5_n3327 ), .A2(_u10_u5_n2905 ), .ZN(_u10_u5_n2500 ) );
NAND2_X1 _u10_u5_U1220  ( .A1(_u10_u5_n2445 ), .A2(_u10_u5_n2500 ), .ZN(_u10_u5_n3325 ) );
NAND2_X1 _u10_u5_U1219  ( .A1(1'b0), .A2(_u10_u5_n2979 ), .ZN(_u10_u5_n3326 ) );
NAND3_X1 _u10_u5_U1218  ( .A1(_u10_u5_n3324 ), .A2(_u10_u5_n3325 ), .A3(_u10_u5_n3326 ), .ZN(_u10_u5_n3309 ) );
AND2_X1 _u10_u5_U1217  ( .A1(_u10_u5_n2877 ), .A2(_u10_u5_n3223 ), .ZN(_u10_u5_n2858 ) );
NAND2_X1 _u10_u5_U1216  ( .A1(_u10_u5_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_21 ), .ZN(_u10_u5_n2346 ) );
INV_X1 _u10_u5_U1215  ( .A(_u10_u5_n2346 ), .ZN(_u10_u5_n2043 ) );
NAND2_X1 _u10_u5_U1214  ( .A1(_u10_u5_n2858 ), .A2(_u10_u5_n2043 ), .ZN(_u10_u5_n3321 ) );
NAND2_X1 _u10_u5_U1213  ( .A1(_u10_u5_n1982 ), .A2(_u10_u5_n2195 ), .ZN(_u10_u5_n3268 ) );
INV_X1 _u10_u5_U1212  ( .A(_u10_u5_n3268 ), .ZN(_u10_u5_n2222 ) );
NAND3_X1 _u10_u5_U1211  ( .A1(_u10_u5_n3323 ), .A2(_u10_u5_n3216 ), .A3(_u10_u5_n2222 ), .ZN(_u10_u5_n3322 ) );
NAND2_X1 _u10_u5_U1210  ( .A1(_u10_u5_n3321 ), .A2(_u10_u5_n3322 ), .ZN(_u10_u5_n2374 ) );
NAND2_X1 _u10_u5_U1209  ( .A1(_u10_u5_n3320 ), .A2(_u10_u5_n3174 ), .ZN(_u10_u5_n2014 ) );
NOR2_X1 _u10_u5_U1208  ( .A1(_u10_u5_n1841 ), .A2(_u10_u5_n2014 ), .ZN(_u10_u5_n2813 ) );
NAND2_X1 _u10_u5_U1207  ( .A1(_u10_u5_n2813 ), .A2(_u10_u5_n2534 ), .ZN(_u10_u5_n3310 ) );
NAND2_X1 _u10_u5_U1206  ( .A1(_u10_u5_n3319 ), .A2(_u10_u5_n3136 ), .ZN(_u10_u5_n1836 ) );
INV_X1 _u10_u5_U1205  ( .A(_u10_u5_n1836 ), .ZN(_u10_u5_n2815 ) );
NAND2_X1 _u10_u5_U1204  ( .A1(_u10_u5_n2534 ), .A2(_u10_u5_n3129 ), .ZN(_u10_u5_n2439 ) );
NAND2_X1 _u10_u5_U1203  ( .A1(_u10_u5_n2055 ), .A2(_u10_u5_n2107 ), .ZN(_u10_u5_n2062 ) );
NAND2_X1 _u10_u5_U1202  ( .A1(_u10_u5_n2439 ), .A2(_u10_u5_n2062 ), .ZN(_u10_u5_n3318 ) );
NAND2_X1 _u10_u5_U1201  ( .A1(_u10_u5_n2815 ), .A2(_u10_u5_n3318 ), .ZN(_u10_u5_n3311 ) );
NAND2_X1 _u10_u5_U1200  ( .A1(_u10_u5_n2986 ), .A2(_u10_u5_n2175 ), .ZN(_u10_u5_n3317 ) );
NAND2_X1 _u10_u5_U1199  ( .A1(_u10_u5_n2253 ), .A2(_u10_u5_n3317 ), .ZN(_u10_u5_n3157 ) );
NAND2_X1 _u10_u5_U1198  ( .A1(_u10_u5_n3316 ), .A2(_u10_u5_n3157 ), .ZN(_u10_u5_n3312 ) );
NOR2_X1 _u10_u5_U1197  ( .A1(_u10_u5_n2495 ), .A2(_u10_u5_n2194 ), .ZN(_u10_u5_n3314 ) );
NOR2_X1 _u10_u5_U1196  ( .A1(_u10_u5_n2375 ), .A2(_u10_u5_n2367 ), .ZN(_u10_u5_n3315 ) );
NOR2_X1 _u10_u5_U1195  ( .A1(_u10_u5_n3314 ), .A2(_u10_u5_n3315 ), .ZN(_u10_u5_n3313 ) );
NAND4_X1 _u10_u5_U1194  ( .A1(_u10_u5_n3310 ), .A2(_u10_u5_n3311 ), .A3(_u10_u5_n3312 ), .A4(_u10_u5_n3313 ), .ZN(_u10_u5_n2315 ) );
NOR4_X1 _u10_u5_U1193  ( .A1(_u10_u5_n3308 ), .A2(_u10_u5_n3309 ), .A3(_u10_u5_n2374 ), .A4(_u10_u5_n2315 ), .ZN(_u10_u5_n3307 ) );
NAND3_X1 _u10_u5_U1192  ( .A1(_u10_u5_n3305 ), .A2(_u10_u5_n3306 ), .A3(_u10_u5_n3307 ), .ZN(_u10_u5_n1987 ) );
AND2_X1 _u10_u5_U1191  ( .A1(1'b0), .A2(_u10_u5_n2977 ), .ZN(_u10_u5_n3240 ));
NAND2_X1 _u10_u5_U1190  ( .A1(_u10_u5_n1891 ), .A2(_u10_u5_n2534 ), .ZN(_u10_u5_n3303 ) );
NAND4_X1 _u10_u5_U1189  ( .A1(_u10_u5_n1982 ), .A2(_u10_u5_n2659 ), .A3(_u10_u5_n2256 ), .A4(_u10_u5_n2175 ), .ZN(_u10_u5_n3304 ) );
AND2_X1 _u10_u5_U1188  ( .A1(_u10_u5_n3303 ), .A2(_u10_u5_n3304 ), .ZN(_u10_u5_n2612 ) );
NAND2_X1 _u10_u5_U1187  ( .A1(_u10_u5_n3302 ), .A2(_u10_u5_n3236 ), .ZN(_u10_u5_n2985 ) );
OR2_X1 _u10_u5_U1186  ( .A1(_u10_u5_n2431 ), .A2(_u10_u5_n2985 ), .ZN(_u10_u5_n3299 ) );
OR2_X1 _u10_u5_U1185  ( .A1(_u10_u5_n2282 ), .A2(_u10_u5_n2359 ), .ZN(_u10_u5_n3300 ) );
NAND2_X1 _u10_u5_U1184  ( .A1(_u10_u5_n1890 ), .A2(_u10_u5_n2534 ), .ZN(_u10_u5_n3301 ) );
NAND4_X1 _u10_u5_U1183  ( .A1(_u10_u5_n2612 ), .A2(_u10_u5_n3299 ), .A3(_u10_u5_n3300 ), .A4(_u10_u5_n3301 ), .ZN(_u10_u5_n3279 ) );
INV_X1 _u10_u5_U1182  ( .A(_u10_u5_n2464 ), .ZN(_u10_u5_n3295 ) );
NAND2_X1 _u10_u5_U1181  ( .A1(_u10_u5_n3295 ), .A2(_u10_u5_n2835 ), .ZN(_u10_u5_n2623 ) );
INV_X1 _u10_u5_U1180  ( .A(_u10_u5_n2623 ), .ZN(_u10_u5_n3185 ) );
INV_X1 _u10_u5_U1179  ( .A(_u10_u5_n2688 ), .ZN(_u10_u5_n2169 ) );
NAND2_X1 _u10_u5_U1178  ( .A1(_u10_u5_n3185 ), .A2(_u10_u5_n2169 ), .ZN(_u10_u5_n3286 ) );
NAND2_X1 _u10_u5_U1177  ( .A1(_u10_u5_n2833 ), .A2(_u10_u5_n3278 ), .ZN(_u10_u5_n3298 ) );
NAND3_X1 _u10_u5_U1176  ( .A1(_u10_u5_n3297 ), .A2(_u10_u5_n2838 ), .A3(_u10_u5_n3298 ), .ZN(_u10_u5_n3296 ) );
NAND2_X1 _u10_u5_U1175  ( .A1(_u10_u5_n2830 ), .A2(_u10_u5_n3296 ), .ZN(_u10_u5_n3287 ) );
NAND2_X1 _u10_u5_U1174  ( .A1(_u10_u5_n3295 ), .A2(_u10_u5_n3001 ), .ZN(_u10_u5_n3292 ) );
NAND2_X1 _u10_u5_U1173  ( .A1(_u10_u5_n3294 ), .A2(_u10_u5_n2089 ), .ZN(_u10_u5_n3293 ) );
AND2_X1 _u10_u5_U1172  ( .A1(_u10_u5_n3292 ), .A2(_u10_u5_n3293 ), .ZN(_u10_u5_n2548 ) );
NAND2_X1 _u10_u5_U1171  ( .A1(_u10_u5_n2548 ), .A2(_u10_u5_n2091 ), .ZN(_u10_u5_n2304 ) );
NAND2_X1 _u10_u5_U1170  ( .A1(_u10_u5_n2304 ), .A2(_u10_u5_n2446 ), .ZN(_u10_u5_n3290 ) );
NAND2_X1 _u10_u5_U1169  ( .A1(_u10_u5_n2549 ), .A2(_u10_u5_n2446 ), .ZN(_u10_u5_n2790 ) );
NOR2_X1 _u10_u5_U1168  ( .A1(_u10_u5_n1936 ), .A2(_u10_u5_n2790 ), .ZN(_u10_u5_n2789 ) );
INV_X1 _u10_u5_U1167  ( .A(_u10_u5_n2789 ), .ZN(_u10_u5_n3291 ) );
OR2_X1 _u10_u5_U1166  ( .A1(_u10_u5_n2828 ), .A2(_u10_u5_n2790 ), .ZN(_u10_u5_n2498 ) );
NAND4_X1 _u10_u5_U1165  ( .A1(_u10_u5_n3290 ), .A2(_u10_u5_n3291 ), .A3(_u10_u5_n2498 ), .A4(_u10_u5_n2001 ), .ZN(_u10_u5_n3289 ) );
NAND2_X1 _u10_u5_U1164  ( .A1(_u10_u5_n2445 ), .A2(_u10_u5_n3289 ), .ZN(_u10_u5_n3288 ) );
NAND3_X1 _u10_u5_U1163  ( .A1(_u10_u5_n3286 ), .A2(_u10_u5_n3287 ), .A3(_u10_u5_n3288 ), .ZN(_u10_u5_n3280 ) );
NOR2_X1 _u10_u5_U1162  ( .A1(_u10_u5_n2940 ), .A2(_u10_u5_n1913 ), .ZN(_u10_u5_n3281 ) );
INV_X1 _u10_u5_U1161  ( .A(1'b0), .ZN(_u10_u5_n1864 ) );
NAND2_X1 _u10_u5_U1160  ( .A1(1'b0), .A2(_u10_u5_n2588 ), .ZN(_u10_u5_n2141 ) );
INV_X1 _u10_u5_U1159  ( .A(_u10_u5_n2141 ), .ZN(_u10_u5_n3159 ) );
NAND3_X1 _u10_u5_U1158  ( .A1(_u10_u5_n2103 ), .A2(_u10_u5_n1864 ), .A3(_u10_u5_n3159 ), .ZN(_u10_u5_n2520 ) );
INV_X1 _u10_u5_U1157  ( .A(_u10_u5_n2520 ), .ZN(_u10_u5_n2630 ) );
INV_X1 _u10_u5_U1156  ( .A(_u10_u5_n2307 ), .ZN(_u10_u5_n2382 ) );
NOR4_X1 _u10_u5_U1155  ( .A1(_u10_u5_n2382 ), .A2(_u10_u5_n2722 ), .A3(_u10_u5_n1925 ), .A4(_u10_u5_n2508 ), .ZN(_u10_u5_n3260 ) );
NOR2_X1 _u10_u5_U1154  ( .A1(_u10_u5_n2498 ), .A2(_u10_u5_n2911 ), .ZN(_u10_u5_n2633 ) );
NOR2_X1 _u10_u5_U1153  ( .A1(_u10_u5_n2633 ), .A2(_u10_u5_n3278 ), .ZN(_u10_u5_n3285 ) );
INV_X1 _u10_u5_U1152  ( .A(_u10_u5_n1866 ), .ZN(_u10_u5_n1926 ) );
NOR2_X1 _u10_u5_U1151  ( .A1(_u10_u5_n3285 ), .A2(_u10_u5_n1926 ), .ZN(_u10_u5_n3284 ) );
NOR4_X1 _u10_u5_U1150  ( .A1(1'b0), .A2(_u10_u5_n2630 ), .A3(_u10_u5_n3260 ),.A4(_u10_u5_n3284 ), .ZN(_u10_u5_n3283 ) );
NOR2_X1 _u10_u5_U1149  ( .A1(_u10_u5_n3283 ), .A2(_u10_u5_n2980 ), .ZN(_u10_u5_n3282 ) );
NOR4_X1 _u10_u5_U1148  ( .A1(_u10_u5_n3279 ), .A2(_u10_u5_n3280 ), .A3(_u10_u5_n3281 ), .A4(_u10_u5_n3282 ), .ZN(_u10_u5_n3241 ) );
NAND2_X1 _u10_u5_U1147  ( .A1(_u10_u5_n1836 ), .A2(_u10_u5_n2291 ), .ZN(_u10_u5_n2147 ) );
NAND2_X1 _u10_u5_U1146  ( .A1(_u10_u5_n2443 ), .A2(_u10_u5_n2147 ), .ZN(_u10_u5_n3261 ) );
INV_X1 _u10_u5_U1145  ( .A(_u10_u5_n1841 ), .ZN(_u10_u5_n2571 ) );
NAND2_X1 _u10_u5_U1144  ( .A1(_u10_u5_n2571 ), .A2(_u10_u5_n3278 ), .ZN(_u10_u5_n3277 ) );
NAND2_X1 _u10_u5_U1143  ( .A1(_u10_u5_n3276 ), .A2(_u10_u5_n3277 ), .ZN(_u10_u5_n2819 ) );
OR2_X1 _u10_u5_U1142  ( .A1(_u10_u5_n2819 ), .A2(_u10_u5_n3275 ), .ZN(_u10_u5_n3273 ) );
NAND2_X1 _u10_u5_U1141  ( .A1(_u10_u5_n2815 ), .A2(_u10_u5_n2080 ), .ZN(_u10_u5_n3274 ) );
NAND2_X1 _u10_u5_U1140  ( .A1(_u10_u5_n2014 ), .A2(_u10_u5_n3274 ), .ZN(_u10_u5_n2165 ) );
NAND2_X1 _u10_u5_U1139  ( .A1(_u10_u5_n3273 ), .A2(_u10_u5_n2165 ), .ZN(_u10_u5_n3262 ) );
NAND2_X1 _u10_u5_U1138  ( .A1(_u10_u5_n2688 ), .A2(_u10_u5_n2126 ), .ZN(_u10_u5_n1956 ) );
INV_X1 _u10_u5_U1137  ( .A(_u10_u5_n1956 ), .ZN(_u10_u5_n1860 ) );
NOR2_X1 _u10_u5_U1136  ( .A1(1'b0), .A2(_u10_u5_n2498 ), .ZN(_u10_u5_n3271 ));
NOR2_X1 _u10_u5_U1135  ( .A1(_u10_u5_n3271 ), .A2(_u10_u5_n3272 ), .ZN(_u10_u5_n3270 ) );
NOR2_X1 _u10_u5_U1134  ( .A1(_u10_u5_n1860 ), .A2(_u10_u5_n3270 ), .ZN(_u10_u5_n3264 ) );
INV_X1 _u10_u5_U1133  ( .A(_u10_u5_n2632 ), .ZN(_u10_u5_n3202 ) );
NAND2_X1 _u10_u5_U1132  ( .A1(_u10_u5_n3236 ), .A2(_u10_u5_n3269 ), .ZN(_u10_u5_n3036 ) );
INV_X1 _u10_u5_U1131  ( .A(_u10_u5_n3036 ), .ZN(_u10_u5_n1960 ) );
NAND2_X1 _u10_u5_U1130  ( .A1(_u10_u5_n3202 ), .A2(_u10_u5_n1960 ), .ZN(_u10_u5_n3079 ) );
NOR3_X1 _u10_u5_U1129  ( .A1(_u10_u5_n3079 ), .A2(1'b0), .A3(_u10_u5_n3268 ),.ZN(_u10_u5_n3265 ) );
INV_X1 _u10_u5_U1128  ( .A(_u10_u5_n2014 ), .ZN(_u10_u5_n2709 ) );
NAND2_X1 _u10_u5_U1127  ( .A1(_u10_u5_n2709 ), .A2(_u10_u5_n2166 ), .ZN(_u10_u5_n2145 ) );
INV_X1 _u10_u5_U1126  ( .A(_u10_u5_n2145 ), .ZN(_u10_u5_n3258 ) );
NOR2_X1 _u10_u5_U1125  ( .A1(_u10_u5_n3258 ), .A2(_u10_u5_n2183 ), .ZN(_u10_u5_n3267 ) );
NOR2_X1 _u10_u5_U1124  ( .A1(_u10_u5_n3267 ), .A2(_u10_u5_n2567 ), .ZN(_u10_u5_n3266 ) );
NOR3_X1 _u10_u5_U1123  ( .A1(_u10_u5_n3264 ), .A2(_u10_u5_n3265 ), .A3(_u10_u5_n3266 ), .ZN(_u10_u5_n3263 ) );
NAND3_X1 _u10_u5_U1122  ( .A1(_u10_u5_n3261 ), .A2(_u10_u5_n3262 ), .A3(_u10_u5_n3263 ), .ZN(_u10_u5_n3243 ) );
INV_X1 _u10_u5_U1121  ( .A(_u10_u5_n2102 ), .ZN(_u10_u5_n2509 ) );
NAND2_X1 _u10_u5_U1120  ( .A1(_u10_u5_n3260 ), .A2(_u10_u5_n2509 ), .ZN(_u10_u5_n3247 ) );
INV_X1 _u10_u5_U1119  ( .A(_u10_u5_n3259 ), .ZN(_u10_u5_n2015 ) );
NAND2_X1 _u10_u5_U1118  ( .A1(_u10_u5_n2015 ), .A2(_u10_u5_n3258 ), .ZN(_u10_u5_n3248 ) );
NAND2_X1 _u10_u5_U1117  ( .A1(_u10_u5_n2251 ), .A2(_u10_u5_n2169 ), .ZN(_u10_u5_n3255 ) );
OR2_X1 _u10_u5_U1116  ( .A1(_u10_u5_n3157 ), .A2(_u10_u5_n2256 ), .ZN(_u10_u5_n3257 ) );
NAND2_X1 _u10_u5_U1115  ( .A1(_u10_u5_n2105 ), .A2(_u10_u5_n3257 ), .ZN(_u10_u5_n3256 ) );
AND2_X1 _u10_u5_U1114  ( .A1(_u10_u5_n3255 ), .A2(_u10_u5_n3256 ), .ZN(_u10_u5_n3212 ) );
INV_X1 _u10_u5_U1113  ( .A(_u10_u5_n2037 ), .ZN(_u10_u5_n2987 ) );
NAND2_X1 _u10_u5_U1112  ( .A1(_u10_u5_n2987 ), .A2(_u10_u5_n2038 ), .ZN(_u10_u5_n2212 ) );
NOR2_X1 _u10_u5_U1111  ( .A1(_u10_u5_n2212 ), .A2(1'b0), .ZN(_u10_u5_n2658 ));
INV_X1 _u10_u5_U1110  ( .A(_u10_u5_n2658 ), .ZN(_u10_u5_n2343 ) );
NAND2_X1 _u10_u5_U1109  ( .A1(_u10_u5_n2344 ), .A2(_u10_u5_n3254 ), .ZN(_u10_u5_n1928 ) );
NAND2_X1 _u10_u5_U1108  ( .A1(_u10_u5_n2588 ), .A2(_u10_u5_n1928 ), .ZN(_u10_u5_n3253 ) );
NAND2_X1 _u10_u5_U1107  ( .A1(_u10_u5_n2343 ), .A2(_u10_u5_n3253 ), .ZN(_u10_u5_n3252 ) );
NAND2_X1 _u10_u5_U1106  ( .A1(_u10_u5_n2105 ), .A2(_u10_u5_n3252 ), .ZN(_u10_u5_n3251 ) );
NAND2_X1 _u10_u5_U1105  ( .A1(_u10_u5_n3212 ), .A2(_u10_u5_n3251 ), .ZN(_u10_u5_n3250 ) );
NAND2_X1 _u10_u5_U1104  ( .A1(_u10_u5_n2307 ), .A2(_u10_u5_n3250 ), .ZN(_u10_u5_n3249 ) );
NAND3_X1 _u10_u5_U1103  ( .A1(_u10_u5_n3247 ), .A2(_u10_u5_n3248 ), .A3(_u10_u5_n3249 ), .ZN(_u10_u5_n3244 ) );
AND2_X1 _u10_u5_U1102  ( .A1(_u10_u5_n2915 ), .A2(_u10_u5_n2059 ), .ZN(_u10_u5_n2957 ) );
AND3_X1 _u10_u5_U1101  ( .A1(_u10_u5_n3223 ), .A2(_u10_u5_n2837 ), .A3(_u10_u5_n2957 ), .ZN(_u10_u5_n2051 ) );
NOR2_X1 _u10_u5_U1100  ( .A1(_u10_u5_n2528 ), .A2(_u10_u5_n2051 ), .ZN(_u10_u5_n2605 ) );
NOR2_X1 _u10_u5_U1099  ( .A1(_u10_u5_n2605 ), .A2(_u10_u5_n2346 ), .ZN(_u10_u5_n3245 ) );
NOR2_X1 _u10_u5_U1098  ( .A1(_u10_u5_n2291 ), .A2(_u10_u5_n2062 ), .ZN(_u10_u5_n3246 ) );
NOR4_X1 _u10_u5_U1097  ( .A1(_u10_u5_n3243 ), .A2(_u10_u5_n3244 ), .A3(_u10_u5_n3245 ), .A4(_u10_u5_n3246 ), .ZN(_u10_u5_n3242 ) );
NAND2_X1 _u10_u5_U1096  ( .A1(_u10_u5_n3241 ), .A2(_u10_u5_n3242 ), .ZN(_u10_u5_n2311 ) );
OR3_X1 _u10_u5_U1095  ( .A1(_u10_u5_n1987 ), .A2(_u10_u5_n3240 ), .A3(_u10_u5_n2311 ), .ZN(_u10_u5_n3192 ) );
INV_X1 _u10_u5_U1094  ( .A(_u10_u5_n2886 ), .ZN(_u10_u5_n2720 ) );
NOR2_X1 _u10_u5_U1093  ( .A1(_u10_u5_n2004 ), .A2(_u10_u5_n2720 ), .ZN(_u10_u5_n2455 ) );
INV_X1 _u10_u5_U1092  ( .A(_u10_u5_n2488 ), .ZN(_u10_u5_n2938 ) );
AND3_X1 _u10_u5_U1091  ( .A1(_u10_u5_n2455 ), .A2(_u10_u5_n1859 ), .A3(_u10_u5_n2938 ), .ZN(_u10_u5_n3239 ) );
INV_X1 _u10_u5_U1090  ( .A(_u10_u5_n2633 ), .ZN(_u10_u5_n2937 ) );
NOR2_X1 _u10_u5_U1089  ( .A1(_u10_u5_n3239 ), .A2(_u10_u5_n2937 ), .ZN(_u10_u5_n3227 ) );
NOR2_X1 _u10_u5_U1088  ( .A1(_u10_u5_n1976 ), .A2(_u10_u5_n1969 ), .ZN(_u10_u5_n3237 ) );
NOR2_X1 _u10_u5_U1087  ( .A1(1'b0), .A2(_u10_u5_n2947 ), .ZN(_u10_u5_n3238 ));
NOR3_X1 _u10_u5_U1086  ( .A1(_u10_u5_n2476 ), .A2(_u10_u5_n3237 ), .A3(_u10_u5_n3238 ), .ZN(_u10_u5_n3235 ) );
NOR3_X1 _u10_u5_U1085  ( .A1(_u10_u5_n1813 ), .A2(_u10_u5_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_20 ), .ZN(_u10_u5_n3135 ) );
NAND2_X1 _u10_u5_U1084  ( .A1(_u10_u5_n3135 ), .A2(_u10_u5_n3236 ), .ZN(_u10_u5_n2573 ) );
NOR2_X1 _u10_u5_U1083  ( .A1(_u10_u5_n3235 ), .A2(_u10_u5_n2573 ), .ZN(_u10_u5_n3228 ) );
NOR2_X1 _u10_u5_U1082  ( .A1(_u10_u5_n2216 ), .A2(_u10_u5_n1868 ), .ZN(_u10_u5_n3233 ) );
INV_X1 _u10_u5_U1081  ( .A(_u10_u5_n2550 ), .ZN(_u10_u5_n2475 ) );
NOR3_X1 _u10_u5_U1080  ( .A1(_u10_u5_n2475 ), .A2(1'b0), .A3(_u10_u5_n1925 ),.ZN(_u10_u5_n3234 ) );
NOR3_X1 _u10_u5_U1079  ( .A1(_u10_u5_n3233 ), .A2(1'b0), .A3(_u10_u5_n3234 ),.ZN(_u10_u5_n3232 ) );
NOR2_X1 _u10_u5_U1078  ( .A1(_u10_u5_n3232 ), .A2(_u10_u5_n2037 ), .ZN(_u10_u5_n3229 ) );
NOR2_X1 _u10_u5_U1077  ( .A1(_u10_u5_n3231 ), .A2(_u10_u5_n2365 ), .ZN(_u10_u5_n3230 ) );
NOR4_X1 _u10_u5_U1076  ( .A1(_u10_u5_n3227 ), .A2(_u10_u5_n3228 ), .A3(_u10_u5_n3229 ), .A4(_u10_u5_n3230 ), .ZN(_u10_u5_n3205 ) );
NOR3_X1 _u10_u5_U1075  ( .A1(_u10_u5_n3226 ), .A2(_u10_u5_n2687 ), .A3(_u10_u5_n2145 ), .ZN(_u10_u5_n3217 ) );
NOR3_X1 _u10_u5_U1074  ( .A1(_u10_u5_n3225 ), .A2(1'b0), .A3(_u10_u5_n2587 ),.ZN(_u10_u5_n3218 ) );
NOR2_X1 _u10_u5_U1073  ( .A1(_u10_u5_n3159 ), .A2(1'b0), .ZN(_u10_u5_n3224 ));
NOR2_X1 _u10_u5_U1072  ( .A1(_u10_u5_n3224 ), .A2(_u10_u5_n2584 ), .ZN(_u10_u5_n3219 ) );
NAND2_X1 _u10_u5_U1071  ( .A1(_u10_u5_n3222 ), .A2(_u10_u5_n3223 ), .ZN(_u10_u5_n2048 ) );
INV_X1 _u10_u5_U1070  ( .A(_u10_u5_n2048 ), .ZN(_u10_u5_n2859 ) );
NOR2_X1 _u10_u5_U1069  ( .A1(_u10_u5_n2859 ), .A2(_u10_u5_n2054 ), .ZN(_u10_u5_n3221 ) );
NOR2_X1 _u10_u5_U1068  ( .A1(_u10_u5_n3221 ), .A2(_u10_u5_n2346 ), .ZN(_u10_u5_n3220 ) );
NOR4_X1 _u10_u5_U1067  ( .A1(_u10_u5_n3217 ), .A2(_u10_u5_n3218 ), .A3(_u10_u5_n3219 ), .A4(_u10_u5_n3220 ), .ZN(_u10_u5_n3206 ) );
NAND2_X1 _u10_u5_U1066  ( .A1(_u10_u5_n2377 ), .A2(_u10_u5_n2721 ), .ZN(_u10_u5_n3213 ) );
AND4_X1 _u10_u5_U1065  ( .A1(1'b0), .A2(_u10_u5_n2502 ), .A3(_u10_u5_n2972 ),.A4(_u10_u5_n3040 ), .ZN(_u10_u5_n2406 ) );
NAND2_X1 _u10_u5_U1064  ( .A1(_u10_u5_n2406 ), .A2(_u10_u5_n2979 ), .ZN(_u10_u5_n3214 ) );
NAND2_X1 _u10_u5_U1063  ( .A1(_u10_u5_n2630 ), .A2(_u10_u5_n3216 ), .ZN(_u10_u5_n2376 ) );
INV_X1 _u10_u5_U1062  ( .A(_u10_u5_n2376 ), .ZN(_u10_u5_n3108 ) );
NAND2_X1 _u10_u5_U1061  ( .A1(_u10_u5_n3108 ), .A2(_u10_u5_n2507 ), .ZN(_u10_u5_n3215 ) );
NOR2_X1 _u10_u5_U1060  ( .A1(_u10_u5_n2937 ), .A2(1'b0), .ZN(_u10_u5_n2649 ));
INV_X1 _u10_u5_U1059  ( .A(_u10_u5_n2253 ), .ZN(_u10_u5_n2971 ) );
NAND2_X1 _u10_u5_U1058  ( .A1(_u10_u5_n2649 ), .A2(_u10_u5_n2971 ), .ZN(_u10_u5_n2918 ) );
NAND4_X1 _u10_u5_U1057  ( .A1(_u10_u5_n3213 ), .A2(_u10_u5_n3214 ), .A3(_u10_u5_n3215 ), .A4(_u10_u5_n2918 ), .ZN(_u10_u5_n3208 ) );
NOR2_X1 _u10_u5_U1056  ( .A1(_u10_u5_n2000 ), .A2(_u10_u5_n2902 ), .ZN(_u10_u5_n3209 ) );
NOR2_X1 _u10_u5_U1055  ( .A1(_u10_u5_n3212 ), .A2(_u10_u5_n2475 ), .ZN(_u10_u5_n3210 ) );
INV_X1 _u10_u5_U1054  ( .A(_u10_u5_n2441 ), .ZN(_u10_u5_n3128 ) );
NOR2_X1 _u10_u5_U1053  ( .A1(_u10_u5_n2356 ), .A2(_u10_u5_n3128 ), .ZN(_u10_u5_n3211 ) );
NOR4_X1 _u10_u5_U1052  ( .A1(_u10_u5_n3208 ), .A2(_u10_u5_n3209 ), .A3(_u10_u5_n3210 ), .A4(_u10_u5_n3211 ), .ZN(_u10_u5_n3207 ) );
NAND3_X1 _u10_u5_U1051  ( .A1(_u10_u5_n3205 ), .A2(_u10_u5_n3206 ), .A3(_u10_u5_n3207 ), .ZN(_u10_u5_n2611 ) );
NOR2_X1 _u10_u5_U1050  ( .A1(_u10_u5_n2212 ), .A2(_u10_u5_n2216 ), .ZN(_u10_u5_n1937 ) );
NOR2_X1 _u10_u5_U1049  ( .A1(_u10_u5_n2533 ), .A2(_u10_u5_n2214 ), .ZN(_u10_u5_n2765 ) );
INV_X1 _u10_u5_U1048  ( .A(_u10_u5_n2005 ), .ZN(_u10_u5_n2111 ) );
AND2_X1 _u10_u5_U1047  ( .A1(_u10_u5_n2765 ), .A2(_u10_u5_n2111 ), .ZN(_u10_u5_n3201 ) );
INV_X1 _u10_u5_U1046  ( .A(_u10_u5_n3059 ), .ZN(_u10_u5_n3076 ) );
NAND2_X1 _u10_u5_U1045  ( .A1(_u10_u5_n3201 ), .A2(_u10_u5_n3076 ), .ZN(_u10_u5_n3204 ) );
NAND2_X1 _u10_u5_U1044  ( .A1(_u10_u5_n1937 ), .A2(_u10_u5_n3204 ), .ZN(_u10_u5_n3193 ) );
NAND2_X1 _u10_u5_U1043  ( .A1(_u10_u5_n2254 ), .A2(_u10_u5_n2212 ), .ZN(_u10_u5_n3203 ) );
NAND3_X1 _u10_u5_U1042  ( .A1(_u10_u5_n3203 ), .A2(_u10_u5_n2175 ), .A3(_u10_u5_n2649 ), .ZN(_u10_u5_n3194 ) );
NOR2_X1 _u10_u5_U1041  ( .A1(_u10_u5_n2985 ), .A2(1'b0), .ZN(_u10_u5_n1959 ));
NAND2_X1 _u10_u5_U1040  ( .A1(_u10_u5_n1959 ), .A2(_u10_u5_n3202 ), .ZN(_u10_u5_n2202 ) );
NAND4_X1 _u10_u5_U1039  ( .A1(_u10_u5_n3079 ), .A2(_u10_u5_n2621 ), .A3(_u10_u5_n2202 ), .A4(_u10_u5_n2798 ), .ZN(_u10_u5_n3200 ) );
NAND2_X1 _u10_u5_U1038  ( .A1(_u10_u5_n3201 ), .A2(_u10_u5_n2937 ), .ZN(_u10_u5_n2772 ) );
NAND2_X1 _u10_u5_U1037  ( .A1(_u10_u5_n3200 ), .A2(_u10_u5_n2772 ), .ZN(_u10_u5_n3195 ) );
NAND2_X1 _u10_u5_U1036  ( .A1(_u10_u5_n2765 ), .A2(_u10_u5_n1869 ), .ZN(_u10_u5_n3199 ) );
NAND2_X1 _u10_u5_U1035  ( .A1(_u10_u5_n2049 ), .A2(_u10_u5_n3199 ), .ZN(_u10_u5_n3057 ) );
NOR2_X1 _u10_u5_U1034  ( .A1(_u10_u5_n2495 ), .A2(_u10_u5_n3057 ), .ZN(_u10_u5_n3197 ) );
NOR2_X1 _u10_u5_U1033  ( .A1(_u10_u5_n2883 ), .A2(_u10_u5_n2485 ), .ZN(_u10_u5_n3198 ) );
NOR2_X1 _u10_u5_U1032  ( .A1(_u10_u5_n3197 ), .A2(_u10_u5_n3198 ), .ZN(_u10_u5_n3196 ) );
NAND4_X1 _u10_u5_U1031  ( .A1(_u10_u5_n3193 ), .A2(_u10_u5_n3194 ), .A3(_u10_u5_n3195 ), .A4(_u10_u5_n3196 ), .ZN(_u10_u5_n2887 ) );
NOR4_X1 _u10_u5_U1030  ( .A1(_u10_u5_n3191 ), .A2(_u10_u5_n3192 ), .A3(_u10_u5_n2611 ), .A4(_u10_u5_n2887 ), .ZN(_u10_u5_n3015 ) );
NAND3_X1 _u10_u5_U1029  ( .A1(_u10_u5_n3190 ), .A2(_u10_u5_n2049 ), .A3(_u10_u5_n2957 ), .ZN(_u10_u5_n2699 ) );
OR2_X1 _u10_u5_U1028  ( .A1(_u10_u5_n2699 ), .A2(_u10_u5_n1813 ), .ZN(_u10_u5_n3187 ) );
NAND3_X1 _u10_u5_U1027  ( .A1(_u10_u5_n2978 ), .A2(_u10_u5_n2405 ), .A3(1'b0), .ZN(_u10_u5_n3188 ) );
NAND4_X1 _u10_u5_U1026  ( .A1(_u10_u5_n3058 ), .A2(_u10_u5_n3187 ), .A3(_u10_u5_n3188 ), .A4(_u10_u5_n3189 ), .ZN(_u10_u5_n3186 ) );
NAND2_X1 _u10_u5_U1025  ( .A1(_u10_u5_n2063 ), .A2(_u10_u5_n3186 ), .ZN(_u10_u5_n3163 ) );
NAND2_X1 _u10_u5_U1024  ( .A1(_u10_u5_n3185 ), .A2(_u10_u5_n2329 ), .ZN(_u10_u5_n3164 ) );
NAND2_X1 _u10_u5_U1023  ( .A1(_u10_u5_n2689 ), .A2(_u10_u5_n2365 ), .ZN(_u10_u5_n2736 ) );
NOR2_X1 _u10_u5_U1022  ( .A1(_u10_u5_n2736 ), .A2(_u10_u5_n2488 ), .ZN(_u10_u5_n1855 ) );
INV_X1 _u10_u5_U1021  ( .A(_u10_u5_n1855 ), .ZN(_u10_u5_n3184 ) );
NOR2_X1 _u10_u5_U1020  ( .A1(_u10_u5_n2274 ), .A2(_u10_u5_n2359 ), .ZN(_u10_u5_n2952 ) );
NOR2_X1 _u10_u5_U1019  ( .A1(_u10_u5_n3184 ), .A2(_u10_u5_n2952 ), .ZN(_u10_u5_n2776 ) );
OR2_X1 _u10_u5_U1018  ( .A1(_u10_u5_n2852 ), .A2(_u10_u5_n2776 ), .ZN(_u10_u5_n3165 ) );
NAND2_X1 _u10_u5_U1017  ( .A1(_u10_u5_n3126 ), .A2(_u10_u5_n2915 ), .ZN(_u10_u5_n3065 ) );
NOR3_X1 _u10_u5_U1016  ( .A1(_u10_u5_n3065 ), .A2(1'b0), .A3(_u10_u5_n2632 ),.ZN(_u10_u5_n3182 ) );
NOR3_X1 _u10_u5_U1015  ( .A1(_u10_u5_n3182 ), .A2(_u10_u5_n3183 ), .A3(_u10_u5_n3108 ), .ZN(_u10_u5_n3181 ) );
NOR2_X1 _u10_u5_U1014  ( .A1(_u10_u5_n3181 ), .A2(_u10_u5_n3162 ), .ZN(_u10_u5_n3167 ) );
INV_X1 _u10_u5_U1013  ( .A(_u10_u5_n3180 ), .ZN(_u10_u5_n3140 ) );
NAND3_X1 _u10_u5_U1012  ( .A1(_u10_u5_n3140 ), .A2(_u10_u5_n2163 ), .A3(_u10_u5_n2092 ), .ZN(_u10_u5_n3175 ) );
NOR4_X1 _u10_u5_U1011  ( .A1(_u10_u5_n2411 ), .A2(_u10_u5_n2710 ), .A3(_u10_u5_n3141 ), .A4(_u10_u5_n3089 ), .ZN(_u10_u5_n3179 ) );
NOR2_X1 _u10_u5_U1010  ( .A1(1'b0), .A2(_u10_u5_n3179 ), .ZN(_u10_u5_n3177 ));
NOR2_X1 _u10_u5_U1009  ( .A1(_u10_u5_n1898 ), .A2(_u10_u5_n1847 ), .ZN(_u10_u5_n3178 ) );
NOR4_X1 _u10_u5_U1008  ( .A1(_u10_u5_n3175 ), .A2(_u10_u5_n3176 ), .A3(_u10_u5_n3177 ), .A4(_u10_u5_n3178 ), .ZN(_u10_u5_n3173 ) );
NAND2_X1 _u10_u5_U1007  ( .A1(_u10_u5_n3135 ), .A2(_u10_u5_n3174 ), .ZN(_u10_u5_n2159 ) );
NOR2_X1 _u10_u5_U1006  ( .A1(_u10_u5_n3173 ), .A2(_u10_u5_n2159 ), .ZN(_u10_u5_n3168 ) );
OR3_X1 _u10_u5_U1005  ( .A1(_u10_u5_n3172 ), .A2(1'b0), .A3(_u10_u5_n3126 ),.ZN(_u10_u5_n3171 ) );
NAND2_X1 _u10_u5_U1004  ( .A1(_u10_u5_n2600 ), .A2(_u10_u5_n3171 ), .ZN(_u10_u5_n3153 ) );
AND3_X1 _u10_u5_U1003  ( .A1(_u10_u5_n3153 ), .A2(_u10_u5_n2947 ), .A3(_u10_u5_n2579 ), .ZN(_u10_u5_n3170 ) );
NOR2_X1 _u10_u5_U1002  ( .A1(_u10_u5_n3170 ), .A2(_u10_u5_n2359 ), .ZN(_u10_u5_n3169 ) );
NOR3_X1 _u10_u5_U1001  ( .A1(_u10_u5_n3167 ), .A2(_u10_u5_n3168 ), .A3(_u10_u5_n3169 ), .ZN(_u10_u5_n3166 ) );
NAND4_X1 _u10_u5_U1000  ( .A1(_u10_u5_n3163 ), .A2(_u10_u5_n3164 ), .A3(_u10_u5_n3165 ), .A4(_u10_u5_n3166 ), .ZN(_u10_u5_n3130 ) );
NAND2_X1 _u10_u5_U999  ( .A1(_u10_u5_n2375 ), .A2(_u10_u5_n3162 ), .ZN(_u10_u5_n1923 ) );
NAND2_X1 _u10_u5_U998  ( .A1(_u10_u5_n3062 ), .A2(_u10_u5_n1923 ), .ZN(_u10_u5_n3154 ) );
NAND2_X1 _u10_u5_U997  ( .A1(_u10_u5_n2103 ), .A2(_u10_u5_n2509 ), .ZN(_u10_u5_n3161 ) );
NAND2_X1 _u10_u5_U996  ( .A1(_u10_u5_n2344 ), .A2(_u10_u5_n3161 ), .ZN(_u10_u5_n3160 ) );
NAND2_X1 _u10_u5_U995  ( .A1(_u10_u5_n3159 ), .A2(_u10_u5_n3160 ), .ZN(_u10_u5_n2635 ) );
AND3_X1 _u10_u5_U994  ( .A1(_u10_u5_n2549 ), .A2(_u10_u5_n2108 ), .A3(_u10_u5_n3126 ), .ZN(_u10_u5_n3093 ) );
NAND2_X1 _u10_u5_U993  ( .A1(_u10_u5_n3093 ), .A2(_u10_u5_n2941 ), .ZN(_u10_u5_n3158 ) );
NAND3_X1 _u10_u5_U992  ( .A1(_u10_u5_n3076 ), .A2(_u10_u5_n3066 ), .A3(_u10_u5_n3158 ), .ZN(_u10_u5_n3156 ) );
NAND2_X1 _u10_u5_U991  ( .A1(_u10_u5_n3156 ), .A2(_u10_u5_n3157 ), .ZN(_u10_u5_n3155 ) );
NAND3_X1 _u10_u5_U990  ( .A1(_u10_u5_n3154 ), .A2(_u10_u5_n2635 ), .A3(_u10_u5_n3155 ), .ZN(_u10_u5_n3131 ) );
INV_X1 _u10_u5_U989  ( .A(_u10_u5_n2594 ), .ZN(_u10_u5_n2846 ) );
NAND3_X1 _u10_u5_U988  ( .A1(_u10_u5_n2162 ), .A2(_u10_u5_n2082 ), .A3(_u10_u5_n2105 ), .ZN(_u10_u5_n2077 ) );
NAND4_X1 _u10_u5_U987  ( .A1(_u10_u5_n3153 ), .A2(_u10_u5_n1969 ), .A3(_u10_u5_n2846 ), .A4(_u10_u5_n2077 ), .ZN(_u10_u5_n3148 ) );
NAND2_X1 _u10_u5_U986  ( .A1(_u10_u5_n2838 ), .A2(_u10_u5_n3128 ), .ZN(_u10_u5_n3152 ) );
NAND2_X1 _u10_u5_U985  ( .A1(_u10_u5_n3152 ), .A2(_u10_u5_n2600 ), .ZN(_u10_u5_n3151 ) );
NAND2_X1 _u10_u5_U984  ( .A1(_u10_u5_n2282 ), .A2(_u10_u5_n3151 ), .ZN(_u10_u5_n2601 ) );
NOR4_X1 _u10_u5_U983  ( .A1(_u10_u5_n2885 ), .A2(_u10_u5_n2534 ), .A3(_u10_u5_n2214 ), .A4(_u10_u5_n3059 ), .ZN(_u10_u5_n3150 ) );
NOR2_X1 _u10_u5_U982  ( .A1(_u10_u5_n3150 ), .A2(_u10_u5_n2853 ), .ZN(_u10_u5_n3149 ) );
NOR4_X1 _u10_u5_U981  ( .A1(_u10_u5_n3148 ), .A2(_u10_u5_n2601 ), .A3(_u10_u5_n3149 ), .A4(_u10_u5_n1975 ), .ZN(_u10_u5_n3146 ) );
NAND3_X1 _u10_u5_U980  ( .A1(_u10_SYNOPSYS_UNCONNECTED_23 ), .A2(_u10_SYNOPSYS_UNCONNECTED_19 ), .A3(_u10_u5_n3147 ), .ZN(_u10_u5_n2071 ) );
NOR2_X1 _u10_u5_U979  ( .A1(_u10_u5_n3146 ), .A2(_u10_u5_n2071 ), .ZN(_u10_u5_n3132 ) );
NOR2_X1 _u10_u5_U978  ( .A1(1'b0), .A2(_u10_u5_n1847 ), .ZN(_u10_u5_n3143 ));
INV_X1 _u10_u5_U977  ( .A(_u10_u5_n3145 ), .ZN(_u10_u5_n3144 ) );
NOR2_X1 _u10_u5_U976  ( .A1(_u10_u5_n3143 ), .A2(_u10_u5_n3144 ), .ZN(_u10_u5_n3142 ) );
NOR2_X1 _u10_u5_U975  ( .A1(1'b0), .A2(_u10_u5_n3142 ), .ZN(_u10_u5_n3137 ));
NAND2_X1 _u10_u5_U974  ( .A1(_u10_u5_n2549 ), .A2(_u10_u5_n3141 ), .ZN(_u10_u5_n3138 ) );
NAND2_X1 _u10_u5_U973  ( .A1(_u10_u5_n1896 ), .A2(_u10_u5_n3140 ), .ZN(_u10_u5_n2544 ) );
NAND2_X1 _u10_u5_U972  ( .A1(_u10_u5_n2089 ), .A2(_u10_u5_n2544 ), .ZN(_u10_u5_n3139 ) );
NAND2_X1 _u10_u5_U971  ( .A1(_u10_u5_n3138 ), .A2(_u10_u5_n3139 ), .ZN(_u10_u5_n2795 ) );
NOR4_X1 _u10_u5_U970  ( .A1(_u10_u5_n2300 ), .A2(_u10_u5_n3137 ), .A3(_u10_u5_n2304 ), .A4(_u10_u5_n2795 ), .ZN(_u10_u5_n3134 ) );
NAND2_X1 _u10_u5_U969  ( .A1(_u10_u5_n3135 ), .A2(_u10_u5_n3136 ), .ZN(_u10_u5_n2085 ) );
NOR2_X1 _u10_u5_U968  ( .A1(_u10_u5_n3134 ), .A2(_u10_u5_n2085 ), .ZN(_u10_u5_n3133 ) );
NOR4_X1 _u10_u5_U967  ( .A1(_u10_u5_n3130 ), .A2(_u10_u5_n3131 ), .A3(_u10_u5_n3132 ), .A4(_u10_u5_n3133 ), .ZN(_u10_u5_n3016 ) );
INV_X1 _u10_u5_U966  ( .A(_u10_u5_n2686 ), .ZN(_u10_u5_n2278 ) );
NAND4_X1 _u10_u5_U965  ( .A1(_u10_u5_n2105 ), .A2(_u10_u5_n2278 ), .A3(_u10_u5_n3129 ), .A4(_u10_u5_n2600 ), .ZN(_u10_u5_n2437 ) );
NAND2_X1 _u10_u5_U964  ( .A1(_u10_u5_n3128 ), .A2(_u10_u5_n2437 ), .ZN(_u10_u5_n3127 ) );
NAND2_X1 _u10_u5_U963  ( .A1(_u10_u5_n2815 ), .A2(_u10_u5_n3127 ), .ZN(_u10_u5_n3098 ) );
INV_X1 _u10_u5_U962  ( .A(_u10_u5_n2573 ), .ZN(_u10_u5_n1967 ) );
NAND2_X1 _u10_u5_U961  ( .A1(_u10_u5_n3126 ), .A2(_u10_u5_n2078 ), .ZN(_u10_u5_n3123 ) );
NAND2_X1 _u10_u5_U960  ( .A1(_u10_u5_n3076 ), .A2(_u10_u5_n1925 ), .ZN(_u10_u5_n3125 ) );
NAND2_X1 _u10_u5_U959  ( .A1(_u10_u5_n2669 ), .A2(_u10_u5_n3125 ), .ZN(_u10_u5_n3124 ) );
NAND4_X1 _u10_u5_U958  ( .A1(_u10_u5_n3122 ), .A2(_u10_u5_n3123 ), .A3(_u10_u5_n3124 ), .A4(_u10_u5_n2579 ), .ZN(_u10_u5_n3121 ) );
NAND2_X1 _u10_u5_U957  ( .A1(_u10_u5_n3121 ), .A2(_u10_u5_n2874 ), .ZN(_u10_u5_n3120 ) );
NAND2_X1 _u10_u5_U956  ( .A1(_u10_u5_n2382 ), .A2(_u10_u5_n3120 ), .ZN(_u10_u5_n3119 ) );
NAND2_X1 _u10_u5_U955  ( .A1(_u10_u5_n1967 ), .A2(_u10_u5_n3119 ), .ZN(_u10_u5_n3099 ) );
NAND2_X1 _u10_u5_U954  ( .A1(_u10_u5_n3118 ), .A2(_u10_u5_n3001 ), .ZN(_u10_u5_n3117 ) );
NAND2_X1 _u10_u5_U953  ( .A1(_u10_u5_n2446 ), .A2(_u10_u5_n3117 ), .ZN(_u10_u5_n3116 ) );
NAND2_X1 _u10_u5_U952  ( .A1(_u10_u5_n2445 ), .A2(_u10_u5_n3116 ), .ZN(_u10_u5_n3100 ) );
OR2_X1 _u10_u5_U951  ( .A1(_u10_u5_n3115 ), .A2(_u10_u5_n2687 ), .ZN(_u10_u5_n3114 ) );
AND3_X1 _u10_u5_U950  ( .A1(_u10_u5_n2061 ), .A2(_u10_u5_n2166 ), .A3(_u10_u5_n3114 ), .ZN(_u10_u5_n3045 ) );
NOR2_X1 _u10_u5_U949  ( .A1(1'b0), .A2(_u10_u5_n3045 ), .ZN(_u10_u5_n3113 ));
NOR2_X1 _u10_u5_U948  ( .A1(_u10_u5_n3113 ), .A2(1'b0), .ZN(_u10_u5_n3112 ));
NOR2_X1 _u10_u5_U947  ( .A1(_u10_u5_n3112 ), .A2(_u10_u5_n2356 ), .ZN(_u10_u5_n3102 ) );
NAND2_X1 _u10_u5_U946  ( .A1(_u10_u5_n2571 ), .A2(_u10_u5_n2165 ), .ZN(_u10_u5_n3078 ) );
NAND2_X1 _u10_u5_U945  ( .A1(_u10_u5_n2365 ), .A2(_u10_u5_n3078 ), .ZN(_u10_u5_n2241 ) );
NOR2_X1 _u10_u5_U944  ( .A1(_u10_u5_n2377 ), .A2(_u10_u5_n2241 ), .ZN(_u10_u5_n3111 ) );
NOR2_X1 _u10_u5_U943  ( .A1(_u10_u5_n3111 ), .A2(_u10_u5_n1869 ), .ZN(_u10_u5_n3103 ) );
NOR2_X1 _u10_u5_U942  ( .A1(_u10_u5_n2999 ), .A2(_u10_u5_n2977 ), .ZN(_u10_u5_n3061 ) );
NOR2_X1 _u10_u5_U941  ( .A1(_u10_u5_n3061 ), .A2(_u10_u5_n2367 ), .ZN(_u10_u5_n3106 ) );
NAND2_X1 _u10_u5_U940  ( .A1(_u10_u5_n2977 ), .A2(_u10_u5_n3000 ), .ZN(_u10_u5_n3110 ) );
NAND2_X1 _u10_u5_U939  ( .A1(_u10_u5_n3109 ), .A2(_u10_u5_n3110 ), .ZN(_u10_u5_n1924 ) );
AND2_X1 _u10_u5_U938  ( .A1(_u10_u5_n1924 ), .A2(_u10_u5_n3108 ), .ZN(_u10_u5_n3107 ) );
NOR2_X1 _u10_u5_U937  ( .A1(_u10_u5_n3106 ), .A2(_u10_u5_n3107 ), .ZN(_u10_u5_n3105 ) );
NOR2_X1 _u10_u5_U936  ( .A1(_u10_u5_n3105 ), .A2(_u10_u5_n2008 ), .ZN(_u10_u5_n3104 ) );
NOR3_X1 _u10_u5_U935  ( .A1(_u10_u5_n3102 ), .A2(_u10_u5_n3103 ), .A3(_u10_u5_n3104 ), .ZN(_u10_u5_n3101 ) );
NAND4_X1 _u10_u5_U934  ( .A1(_u10_u5_n3098 ), .A2(_u10_u5_n3099 ), .A3(_u10_u5_n3100 ), .A4(_u10_u5_n3101 ), .ZN(_u10_u5_n3071 ) );
NOR2_X1 _u10_u5_U933  ( .A1(_u10_u5_n1926 ), .A2(_u10_u5_n2980 ), .ZN(_u10_u5_n2218 ) );
INV_X1 _u10_u5_U932  ( .A(_u10_u5_n2721 ), .ZN(_u10_u5_n2910 ) );
NAND2_X1 _u10_u5_U931  ( .A1(_u10_u5_n2910 ), .A2(_u10_u5_n1869 ), .ZN(_u10_u5_n2779 ) );
NAND2_X1 _u10_u5_U930  ( .A1(_u10_u5_n2218 ), .A2(_u10_u5_n2779 ), .ZN(_u10_u5_n3081 ) );
NAND2_X1 _u10_u5_U929  ( .A1(_u10_u5_n1922 ), .A2(_u10_u5_n1864 ), .ZN(_u10_u5_n2179 ) );
NOR3_X1 _u10_u5_U928  ( .A1(_u10_u5_n1961 ), .A2(_u10_u5_n1918 ), .A3(_u10_u5_n2179 ), .ZN(_u10_u5_n2693 ) );
NAND2_X1 _u10_u5_U927  ( .A1(_u10_u5_n3097 ), .A2(_u10_u5_n1924 ), .ZN(_u10_u5_n3096 ) );
NAND2_X1 _u10_u5_U926  ( .A1(_u10_u5_n1984 ), .A2(_u10_u5_n3096 ), .ZN(_u10_u5_n2506 ) );
INV_X1 _u10_u5_U925  ( .A(_u10_u5_n2506 ), .ZN(_u10_u5_n2366 ) );
NAND2_X1 _u10_u5_U924  ( .A1(_u10_u5_n2366 ), .A2(_u10_u5_n2375 ), .ZN(_u10_u5_n2236 ) );
NAND2_X1 _u10_u5_U923  ( .A1(_u10_u5_n2693 ), .A2(_u10_u5_n2236 ), .ZN(_u10_u5_n3082 ) );
NAND2_X1 _u10_u5_U922  ( .A1(1'b0), .A2(_u10_u5_n2126 ), .ZN(_u10_u5_n3095 ));
NAND2_X1 _u10_u5_U921  ( .A1(_u10_u5_n1956 ), .A2(_u10_u5_n3095 ), .ZN(_u10_u5_n2907 ) );
OR2_X1 _u10_u5_U920  ( .A1(_u10_u5_n2902 ), .A2(_u10_u5_n2907 ), .ZN(_u10_u5_n3085 ) );
NAND2_X1 _u10_u5_U919  ( .A1(_u10_u5_n2256 ), .A2(_u10_u5_n2113 ), .ZN(_u10_u5_n3094 ) );
NAND2_X1 _u10_u5_U918  ( .A1(_u10_u5_n2688 ), .A2(_u10_u5_n3094 ), .ZN(_u10_u5_n3092 ) );
NAND2_X1 _u10_u5_U917  ( .A1(_u10_u5_n3093 ), .A2(_u10_u5_n3092 ), .ZN(_u10_u5_n3086 ) );
INV_X1 _u10_u5_U916  ( .A(_u10_u5_n2159 ), .ZN(_u10_u5_n1894 ) );
NAND2_X1 _u10_u5_U915  ( .A1(_u10_u5_n3067 ), .A2(_u10_u5_n1894 ), .ZN(_u10_u5_n3091 ) );
INV_X1 _u10_u5_U914  ( .A(_u10_u5_n3092 ), .ZN(_u10_u5_n2234 ) );
NAND3_X1 _u10_u5_U913  ( .A1(_u10_u5_n3091 ), .A2(_u10_u5_n2126 ), .A3(_u10_u5_n2234 ), .ZN(_u10_u5_n3090 ) );
NAND2_X1 _u10_u5_U912  ( .A1(1'b0), .A2(_u10_u5_n3090 ), .ZN(_u10_u5_n3087 ));
NAND3_X1 _u10_u5_U911  ( .A1(_u10_u5_n2329 ), .A2(_u10_u5_n3089 ), .A3(_u10_u5_n2549 ), .ZN(_u10_u5_n3088 ) );
NAND4_X1 _u10_u5_U910  ( .A1(_u10_u5_n3085 ), .A2(_u10_u5_n3086 ), .A3(_u10_u5_n3087 ), .A4(_u10_u5_n3088 ), .ZN(_u10_u5_n3084 ) );
NAND2_X1 _u10_u5_U909  ( .A1(_u10_u5_n3084 ), .A2(_u10_u5_n2803 ), .ZN(_u10_u5_n3083 ) );
NAND3_X1 _u10_u5_U908  ( .A1(_u10_u5_n3081 ), .A2(_u10_u5_n3082 ), .A3(_u10_u5_n3083 ), .ZN(_u10_u5_n3072 ) );
INV_X1 _u10_u5_U907  ( .A(_u10_u5_n2689 ), .ZN(_u10_u5_n1955 ) );
NOR3_X1 _u10_u5_U906  ( .A1(_u10_u5_n1955 ), .A2(_u10_u5_n2813 ), .A3(_u10_u5_n2488 ), .ZN(_u10_u5_n3080 ) );
NOR2_X1 _u10_u5_U905  ( .A1(_u10_u5_n3080 ), .A2(_u10_u5_n2485 ), .ZN(_u10_u5_n3073 ) );
NAND3_X1 _u10_u5_U904  ( .A1(_u10_u5_n2621 ), .A2(_u10_u5_n2202 ), .A3(_u10_u5_n3079 ), .ZN(_u10_u5_n2110 ) );
NOR2_X1 _u10_u5_U903  ( .A1(_u10_u5_n2110 ), .A2(_u10_u5_n2218 ), .ZN(_u10_u5_n2775 ) );
INV_X1 _u10_u5_U902  ( .A(_u10_u5_n2775 ), .ZN(_u10_u5_n3024 ) );
INV_X1 _u10_u5_U901  ( .A(_u10_u5_n3078 ), .ZN(_u10_u5_n2133 ) );
INV_X1 _u10_u5_U900  ( .A(_u10_u5_n2007 ), .ZN(_u10_u5_n2358 ) );
NAND2_X1 _u10_u5_U899  ( .A1(_u10_u5_n2358 ), .A2(_u10_u5_n2886 ), .ZN(_u10_u5_n2240 ) );
INV_X1 _u10_u5_U898  ( .A(_u10_u5_n2240 ), .ZN(_u10_u5_n2083 ) );
NOR3_X1 _u10_u5_U897  ( .A1(_u10_u5_n2952 ), .A2(_u10_u5_n2004 ), .A3(_u10_u5_n1891 ), .ZN(_u10_u5_n3077 ) );
NAND3_X1 _u10_u5_U896  ( .A1(_u10_u5_n2083 ), .A2(_u10_u5_n2938 ), .A3(_u10_u5_n3077 ), .ZN(_u10_u5_n1886 ) );
NOR3_X1 _u10_u5_U895  ( .A1(_u10_u5_n3024 ), .A2(_u10_u5_n2133 ), .A3(_u10_u5_n1886 ), .ZN(_u10_u5_n3075 ) );
NOR2_X1 _u10_u5_U894  ( .A1(_u10_u5_n3075 ), .A2(_u10_u5_n3076 ), .ZN(_u10_u5_n3074 ) );
NOR4_X1 _u10_u5_U893  ( .A1(_u10_u5_n3071 ), .A2(_u10_u5_n3072 ), .A3(_u10_u5_n3073 ), .A4(_u10_u5_n3074 ), .ZN(_u10_u5_n3017 ) );
INV_X1 _u10_u5_U892  ( .A(_u10_u5_n3065 ), .ZN(_u10_u5_n3043 ) );
NAND2_X1 _u10_u5_U891  ( .A1(_u10_u5_n3043 ), .A2(_u10_u5_n2106 ), .ZN(_u10_u5_n3070 ) );
NAND2_X1 _u10_u5_U890  ( .A1(_u10_u5_n3070 ), .A2(_u10_u5_n2038 ), .ZN(_u10_u5_n3068 ) );
NAND2_X1 _u10_u5_U889  ( .A1(_u10_u5_n2344 ), .A2(_u10_u5_n2584 ), .ZN(_u10_u5_n3069 ) );
NAND3_X1 _u10_u5_U888  ( .A1(_u10_u5_n3068 ), .A2(_u10_u5_n1930 ), .A3(_u10_u5_n3069 ), .ZN(_u10_u5_n3047 ) );
NAND2_X1 _u10_u5_U887  ( .A1(_u10_u5_n2835 ), .A2(_u10_u5_n2466 ), .ZN(_u10_u5_n2130 ) );
INV_X1 _u10_u5_U886  ( .A(_u10_u5_n2130 ), .ZN(_u10_u5_n2168 ) );
NAND3_X1 _u10_u5_U885  ( .A1(_u10_u5_n3067 ), .A2(_u10_u5_n2329 ), .A3(_u10_u5_n2168 ), .ZN(_u10_u5_n2665 ) );
NAND3_X1 _u10_u5_U884  ( .A1(_u10_u5_n3065 ), .A2(_u10_u5_n3066 ), .A3(_u10_u5_n2342 ), .ZN(_u10_u5_n3064 ) );
NAND3_X1 _u10_u5_U883  ( .A1(_u10_u5_n3064 ), .A2(_u10_u5_n2175 ), .A3(_u10_u5_n2987 ), .ZN(_u10_u5_n3048 ) );
NOR3_X1 _u10_u5_U882  ( .A1(_u10_u5_n1849 ), .A2(1'b0), .A3(_u10_u5_n3063 ),.ZN(_u10_u5_n3050 ) );
NOR3_X1 _u10_u5_U881  ( .A1(_u10_u5_n2406 ), .A2(1'b0), .A3(_u10_u5_n3062 ),.ZN(_u10_u5_n3060 ) );
NOR3_X1 _u10_u5_U880  ( .A1(_u10_u5_n3060 ), .A2(1'b0), .A3(_u10_u5_n3061 ),.ZN(_u10_u5_n3051 ) );
NAND2_X1 _u10_u5_U879  ( .A1(_u10_u5_n3059 ), .A2(_u10_u5_n2049 ), .ZN(_u10_u5_n3056 ) );
NAND3_X1 _u10_u5_U878  ( .A1(_u10_u5_n3056 ), .A2(_u10_u5_n3057 ), .A3(_u10_u5_n3058 ), .ZN(_u10_u5_n3054 ) );
NOR4_X1 _u10_u5_U877  ( .A1(_u10_u5_n3054 ), .A2(_u10_u5_n3055 ), .A3(_u10_u5_n2055 ), .A4(_u10_u5_n2056 ), .ZN(_u10_u5_n3053 ) );
NOR3_X1 _u10_u5_U876  ( .A1(_u10_u5_n2346 ), .A2(1'b0), .A3(_u10_u5_n3053 ),.ZN(_u10_u5_n3052 ) );
NOR3_X1 _u10_u5_U875  ( .A1(_u10_u5_n3050 ), .A2(_u10_u5_n3051 ), .A3(_u10_u5_n3052 ), .ZN(_u10_u5_n3049 ) );
NAND4_X1 _u10_u5_U874  ( .A1(_u10_u5_n3047 ), .A2(_u10_u5_n2665 ), .A3(_u10_u5_n3048 ), .A4(_u10_u5_n3049 ), .ZN(_u10_u5_n3019 ) );
NAND2_X1 _u10_u5_U873  ( .A1(_u10_u5_n2056 ), .A2(_u10_u5_n2019 ), .ZN(_u10_u5_n3046 ) );
NAND2_X1 _u10_u5_U872  ( .A1(_u10_u5_n3045 ), .A2(_u10_u5_n3046 ), .ZN(_u10_u5_n3044 ) );
NAND2_X1 _u10_u5_U871  ( .A1(_u10_u5_n3044 ), .A2(_u10_u5_n2165 ), .ZN(_u10_u5_n3028 ) );
OR2_X1 _u10_u5_U870  ( .A1(_u10_u5_n2179 ), .A2(_u10_u5_n1961 ), .ZN(_u10_u5_n3037 ) );
NAND2_X1 _u10_u5_U869  ( .A1(_u10_u5_n3043 ), .A2(_u10_u5_n2336 ), .ZN(_u10_u5_n3042 ) );
NAND2_X1 _u10_u5_U868  ( .A1(_u10_u5_n3042 ), .A2(_u10_u5_n3006 ), .ZN(_u10_u5_n3041 ) );
NAND2_X1 _u10_u5_U867  ( .A1(_u10_u5_n3040 ), .A2(_u10_u5_n3041 ), .ZN(_u10_u5_n3026 ) );
NAND4_X1 _u10_u5_U866  ( .A1(_u10_u5_n3026 ), .A2(_u10_u5_n2520 ), .A3(_u10_u5_n1962 ), .A4(_u10_u5_n1864 ), .ZN(_u10_u5_n3039 ) );
NAND2_X1 _u10_u5_U865  ( .A1(_u10_u5_n3039 ), .A2(_u10_u5_n1922 ), .ZN(_u10_u5_n3038 ) );
NAND2_X1 _u10_u5_U864  ( .A1(_u10_u5_n3037 ), .A2(_u10_u5_n3038 ), .ZN(_u10_u5_n3035 ) );
NAND2_X1 _u10_u5_U863  ( .A1(_u10_u5_n2985 ), .A2(_u10_u5_n3036 ), .ZN(_u10_u5_n2432 ) );
NAND2_X1 _u10_u5_U862  ( .A1(_u10_u5_n3035 ), .A2(_u10_u5_n2432 ), .ZN(_u10_u5_n3029 ) );
INV_X1 _u10_u5_U861  ( .A(_u10_u5_n3034 ), .ZN(_u10_u5_n2777 ) );
INV_X1 _u10_u5_U860  ( .A(_u10_u5_n2772 ), .ZN(_u10_u5_n3032 ) );
NAND2_X1 _u10_u5_U859  ( .A1(_u10_u5_n1982 ), .A2(_u10_u5_n2978 ), .ZN(_u10_u5_n3033 ) );
NAND2_X1 _u10_u5_U858  ( .A1(_u10_u5_n3032 ), .A2(_u10_u5_n3033 ), .ZN(_u10_u5_n3031 ) );
NAND2_X1 _u10_u5_U857  ( .A1(_u10_u5_n2777 ), .A2(_u10_u5_n3031 ), .ZN(_u10_u5_n3030 ) );
NAND3_X1 _u10_u5_U856  ( .A1(_u10_u5_n3028 ), .A2(_u10_u5_n3029 ), .A3(_u10_u5_n3030 ), .ZN(_u10_u5_n3020 ) );
NOR3_X1 _u10_u5_U855  ( .A1(_u10_u5_n2179 ), .A2(1'b0), .A3(_u10_u5_n2375 ),.ZN(_u10_u5_n3027 ) );
NOR2_X1 _u10_u5_U854  ( .A1(_u10_u5_n3027 ), .A2(_u10_u5_n2177 ), .ZN(_u10_u5_n3025 ) );
NOR2_X1 _u10_u5_U853  ( .A1(_u10_u5_n3025 ), .A2(_u10_u5_n3026 ), .ZN(_u10_u5_n3021 ) );
NOR2_X1 _u10_u5_U852  ( .A1(_u10_u5_n2256 ), .A2(_u10_u5_n3024 ), .ZN(_u10_u5_n3023 ) );
NOR2_X1 _u10_u5_U851  ( .A1(_u10_u5_n3023 ), .A2(_u10_u5_n1868 ), .ZN(_u10_u5_n3022 ) );
NOR4_X1 _u10_u5_U850  ( .A1(_u10_u5_n3019 ), .A2(_u10_u5_n3020 ), .A3(_u10_u5_n3021 ), .A4(_u10_u5_n3022 ), .ZN(_u10_u5_n3018 ) );
NAND4_X1 _u10_u5_U849  ( .A1(_u10_u5_n3015 ), .A2(_u10_u5_n3016 ), .A3(_u10_u5_n3017 ), .A4(_u10_u5_n3018 ), .ZN(_u10_u5_n2958 ) );
NOR2_X1 _u10_u5_U848  ( .A1(1'b0), .A2(_u10_u5_n2573 ), .ZN(_u10_u5_n3011 ));
NOR2_X1 _u10_u5_U847  ( .A1(1'b0), .A2(_u10_u5_n2359 ), .ZN(_u10_u5_n3012 ));
NOR2_X1 _u10_u5_U846  ( .A1(1'b0), .A2(_u10_u5_n1859 ), .ZN(_u10_u5_n3013 ));
NOR2_X1 _u10_u5_U845  ( .A1(1'b0), .A2(_u10_u5_n1836 ), .ZN(_u10_u5_n3014 ));
NOR4_X1 _u10_u5_U844  ( .A1(_u10_u5_n3011 ), .A2(_u10_u5_n3012 ), .A3(_u10_u5_n3013 ), .A4(_u10_u5_n3014 ), .ZN(_u10_u5_n2959 ) );
NOR2_X1 _u10_u5_U843  ( .A1(1'b0), .A2(_u10_u5_n2025 ), .ZN(_u10_u5_n3007 ));
NOR2_X1 _u10_u5_U842  ( .A1(1'b0), .A2(_u10_u5_n2085 ), .ZN(_u10_u5_n3008 ));
NOR2_X1 _u10_u5_U841  ( .A1(1'b0), .A2(_u10_u5_n2607 ), .ZN(_u10_u5_n3009 ));
NOR2_X1 _u10_u5_U840  ( .A1(1'b0), .A2(_u10_u5_n2071 ), .ZN(_u10_u5_n3010 ));
NOR4_X1 _u10_u5_U839  ( .A1(_u10_u5_n3007 ), .A2(_u10_u5_n3008 ), .A3(_u10_u5_n3009 ), .A4(_u10_u5_n3010 ), .ZN(_u10_u5_n2960 ) );
NAND2_X1 _u10_u5_U838  ( .A1(_u10_u5_n1894 ), .A2(_u10_u5_n2466 ), .ZN(_u10_u5_n3002 ) );
NAND2_X1 _u10_u5_U837  ( .A1(_u10_u5_n2830 ), .A2(_u10_u5_n2600 ), .ZN(_u10_u5_n3003 ) );
NAND2_X1 _u10_u5_U836  ( .A1(_u10_u5_n1960 ), .A2(_u10_u5_n2431 ), .ZN(_u10_u5_n3004 ) );
NAND2_X1 _u10_u5_U835  ( .A1(_u10_u5_n2002 ), .A2(_u10_u5_n3006 ), .ZN(_u10_u5_n3005 ) );
NAND4_X1 _u10_u5_U834  ( .A1(_u10_u5_n3002 ), .A2(_u10_u5_n3003 ), .A3(_u10_u5_n3004 ), .A4(_u10_u5_n3005 ), .ZN(_u10_u5_n2992 ) );
NAND2_X1 _u10_u5_U833  ( .A1(_u10_u5_n2461 ), .A2(_u10_u5_n3001 ), .ZN(_u10_u5_n2997 ) );
NAND2_X1 _u10_u5_U832  ( .A1(_u10_u5_n2999 ), .A2(_u10_u5_n3000 ), .ZN(_u10_u5_n2998 ) );
NAND2_X1 _u10_u5_U831  ( .A1(_u10_u5_n2997 ), .A2(_u10_u5_n2998 ), .ZN(_u10_u5_n2993 ) );
NOR2_X1 _u10_u5_U830  ( .A1(_u10_SYNOPSYS_UNCONNECTED_19 ), .A2(_u10_u5_n2996 ), .ZN(_u10_u5_n2995 ) );
NOR2_X1 _u10_u5_U829  ( .A1(_u10_u5_n2995 ), .A2(_u10_u5_n2126 ), .ZN(_u10_u5_n2994 ) );
NOR4_X1 _u10_u5_U828  ( .A1(_u10_u5_n2992 ), .A2(_u10_u5_n2993 ), .A3(next_ch), .A4(_u10_u5_n2994 ), .ZN(_u10_u5_n2961 ) );
NAND2_X1 _u10_u5_U827  ( .A1(_u10_u5_n2445 ), .A2(_u10_u5_n2803 ), .ZN(_u10_u5_n2988 ) );
OR2_X1 _u10_u5_U826  ( .A1(_u10_u5_n2584 ), .A2(1'b0), .ZN(_u10_u5_n2989 ));
NAND2_X1 _u10_u5_U825  ( .A1(_u10_u5_n2709 ), .A2(_u10_u5_n2080 ), .ZN(_u10_u5_n2990 ) );
NAND2_X1 _u10_u5_U824  ( .A1(_u10_u5_n2183 ), .A2(_u10_u5_n2166 ), .ZN(_u10_u5_n2991 ) );
NAND4_X1 _u10_u5_U823  ( .A1(_u10_u5_n2988 ), .A2(_u10_u5_n2989 ), .A3(_u10_u5_n2990 ), .A4(_u10_u5_n2991 ), .ZN(_u10_u5_n2963 ) );
NAND2_X1 _u10_u5_U822  ( .A1(_u10_u5_n2987 ), .A2(_u10_u5_n1930 ), .ZN(_u10_u5_n2981 ) );
NAND2_X1 _u10_u5_U821  ( .A1(_u10_u5_n2986 ), .A2(_u10_u5_n2038 ), .ZN(_u10_u5_n2982 ) );
OR2_X1 _u10_u5_U820  ( .A1(_u10_u5_n2985 ), .A2(1'b0), .ZN(_u10_u5_n2983 ));
NAND2_X1 _u10_u5_U819  ( .A1(_u10_u5_n2169 ), .A2(_u10_u5_n2113 ), .ZN(_u10_u5_n2984 ) );
NAND4_X1 _u10_u5_U818  ( .A1(_u10_u5_n2981 ), .A2(_u10_u5_n2982 ), .A3(_u10_u5_n2983 ), .A4(_u10_u5_n2984 ), .ZN(_u10_u5_n2964 ) );
NAND2_X1 _u10_u5_U817  ( .A1(_u10_u5_n2509 ), .A2(_u10_u5_n1864 ), .ZN(_u10_u5_n2973 ) );
INV_X1 _u10_u5_U816  ( .A(_u10_u5_n2980 ), .ZN(_u10_u5_n1861 ) );
NAND2_X1 _u10_u5_U815  ( .A1(_u10_u5_n1861 ), .A2(_u10_u5_n1922 ), .ZN(_u10_u5_n2974 ) );
NAND2_X1 _u10_u5_U814  ( .A1(_u10_u5_n2979 ), .A2(_u10_u5_n2405 ), .ZN(_u10_u5_n2975 ) );
NAND2_X1 _u10_u5_U813  ( .A1(_u10_u5_n2977 ), .A2(_u10_u5_n2978 ), .ZN(_u10_u5_n2976 ) );
NAND4_X1 _u10_u5_U812  ( .A1(_u10_u5_n2973 ), .A2(_u10_u5_n2974 ), .A3(_u10_u5_n2975 ), .A4(_u10_u5_n2976 ), .ZN(_u10_u5_n2965 ) );
NAND2_X1 _u10_u5_U811  ( .A1(_u10_u5_n2507 ), .A2(_u10_u5_n2972 ), .ZN(_u10_u5_n2967 ) );
NAND2_X1 _u10_u5_U810  ( .A1(_u10_u5_n2043 ), .A2(_u10_u5_n1965 ), .ZN(_u10_u5_n2968 ) );
NAND2_X1 _u10_u5_U809  ( .A1(_u10_u5_n2063 ), .A2(_u10_u5_n1853 ), .ZN(_u10_u5_n2969 ) );
NAND2_X1 _u10_u5_U808  ( .A1(_u10_u5_n2971 ), .A2(_u10_u5_n2175 ), .ZN(_u10_u5_n2970 ) );
NAND4_X1 _u10_u5_U807  ( .A1(_u10_u5_n2967 ), .A2(_u10_u5_n2968 ), .A3(_u10_u5_n2969 ), .A4(_u10_u5_n2970 ), .ZN(_u10_u5_n2966 ) );
NOR4_X1 _u10_u5_U806  ( .A1(_u10_u5_n2963 ), .A2(_u10_u5_n2964 ), .A3(_u10_u5_n2965 ), .A4(_u10_u5_n2966 ), .ZN(_u10_u5_n2962 ) );
AND4_X1 _u10_u5_U805  ( .A1(_u10_u5_n2959 ), .A2(_u10_u5_n2960 ), .A3(_u10_u5_n2961 ), .A4(_u10_u5_n2962 ), .ZN(_u10_u5_n1819 ) );
MUX2_X1 _u10_u5_U804  ( .A(_u10_u5_n2958 ), .B(_u10_SYNOPSYS_UNCONNECTED_23 ), .S(_u10_u5_n1819 ), .Z(_u10_u5_n1808 ) );
NOR2_X1 _u10_u5_U803  ( .A1(_u10_u5_n2531 ), .A2(_u10_u5_n2607 ), .ZN(_u10_u5_n1911 ) );
NAND2_X1 _u10_u5_U802  ( .A1(_u10_u5_n1911 ), .A2(_u10_u5_n2957 ), .ZN(_u10_u5_n2954 ) );
NAND2_X1 _u10_u5_U801  ( .A1(_u10_u5_n1853 ), .A2(_u10_u5_n1965 ), .ZN(_u10_u5_n2956 ) );
NAND2_X1 _u10_u5_U800  ( .A1(_u10_u5_n1966 ), .A2(_u10_u5_n2956 ), .ZN(_u10_u5_n2955 ) );
NAND2_X1 _u10_u5_U799  ( .A1(_u10_u5_n2954 ), .A2(_u10_u5_n2955 ), .ZN(_u10_u5_n2670 ) );
NOR3_X1 _u10_u5_U798  ( .A1(_u10_u5_n1852 ), .A2(1'b0), .A3(_u10_u5_n1853 ),.ZN(_u10_u5_n2708 ) );
NAND2_X1 _u10_u5_U797  ( .A1(_u10_u5_n2708 ), .A2(_u10_u5_n2080 ), .ZN(_u10_u5_n2355 ) );
NOR2_X1 _u10_u5_U796  ( .A1(_u10_u5_n2355 ), .A2(1'b0), .ZN(_u10_u5_n2599 ));
NAND2_X1 _u10_u5_U795  ( .A1(_u10_u5_n2953 ), .A2(_u10_u5_n2599 ), .ZN(_u10_u5_n2423 ) );
OR2_X1 _u10_u5_U794  ( .A1(_u10_u5_n2423 ), .A2(_u10_u5_n2359 ), .ZN(_u10_u5_n2949 ) );
NAND3_X1 _u10_u5_U793  ( .A1(_u10_u5_n2105 ), .A2(_u10_u5_n1936 ), .A3(_u10_u5_n2952 ), .ZN(_u10_u5_n2950 ) );
NAND3_X1 _u10_u5_U792  ( .A1(_u10_u5_n2549 ), .A2(_u10_u5_n1936 ), .A3(1'b0),.ZN(_u10_u5_n2096 ) );
INV_X1 _u10_u5_U791  ( .A(_u10_u5_n2096 ), .ZN(_u10_u5_n2301 ) );
NAND2_X1 _u10_u5_U790  ( .A1(_u10_u5_n2301 ), .A2(_u10_u5_n2446 ), .ZN(_u10_u5_n2368 ) );
INV_X1 _u10_u5_U789  ( .A(_u10_u5_n2368 ), .ZN(_u10_u5_n2326 ) );
NAND2_X1 _u10_u5_U788  ( .A1(_u10_u5_n2326 ), .A2(_u10_u5_n2941 ), .ZN(_u10_u5_n2800 ) );
INV_X1 _u10_u5_U787  ( .A(_u10_u5_n2800 ), .ZN(_u10_u5_n2081 ) );
NAND2_X1 _u10_u5_U786  ( .A1(_u10_u5_n2081 ), .A2(_u10_u5_n2049 ), .ZN(_u10_u5_n2855 ) );
INV_X1 _u10_u5_U785  ( .A(_u10_u5_n2855 ), .ZN(_u10_u5_n2347 ) );
NAND2_X1 _u10_u5_U784  ( .A1(_u10_u5_n2347 ), .A2(_u10_u5_n2063 ), .ZN(_u10_u5_n2951 ) );
NAND3_X1 _u10_u5_U783  ( .A1(_u10_u5_n2949 ), .A2(_u10_u5_n2950 ), .A3(_u10_u5_n2951 ), .ZN(_u10_u5_n1997 ) );
INV_X1 _u10_u5_U782  ( .A(_u10_u5_n1997 ), .ZN(_u10_u5_n2917 ) );
AND2_X1 _u10_u5_U781  ( .A1(_u10_u5_n2709 ), .A2(_u10_u5_n2708 ), .ZN(_u10_u5_n2942 ) );
INV_X1 _u10_u5_U780  ( .A(_u10_u5_n2907 ), .ZN(_u10_u5_n2737 ) );
NAND2_X1 _u10_u5_U779  ( .A1(_u10_u5_n2737 ), .A2(_u10_u5_n2803 ), .ZN(_u10_u5_n1888 ) );
NOR2_X1 _u10_u5_U778  ( .A1(_u10_u5_n2001 ), .A2(_u10_u5_n1888 ), .ZN(_u10_u5_n2943 ) );
NAND4_X1 _u10_u5_U777  ( .A1(1'b0), .A2(_u10_u5_n2078 ), .A3(_u10_u5_n2059 ),.A4(_u10_u5_n2031 ), .ZN(_u10_u5_n2578 ) );
NOR3_X1 _u10_u5_U776  ( .A1(_u10_u5_n2719 ), .A2(_u10_u5_n2130 ), .A3(_u10_u5_n2305 ), .ZN(_u10_u5_n2386 ) );
NAND2_X1 _u10_u5_U775  ( .A1(_u10_u5_n2386 ), .A2(_u10_u5_n2669 ), .ZN(_u10_u5_n2948 ) );
NAND3_X1 _u10_u5_U774  ( .A1(_u10_u5_n2578 ), .A2(_u10_u5_n2947 ), .A3(_u10_u5_n2948 ), .ZN(_u10_u5_n2750 ) );
NOR2_X1 _u10_u5_U773  ( .A1(_u10_u5_n2274 ), .A2(_u10_u5_n2852 ), .ZN(_u10_u5_n2946 ) );
NOR3_X1 _u10_u5_U772  ( .A1(_u10_u5_n2750 ), .A2(1'b0), .A3(_u10_u5_n2946 ),.ZN(_u10_u5_n2945 ) );
NOR2_X1 _u10_u5_U771  ( .A1(_u10_u5_n2945 ), .A2(_u10_u5_n2359 ), .ZN(_u10_u5_n2944 ) );
NOR3_X1 _u10_u5_U770  ( .A1(_u10_u5_n2942 ), .A2(_u10_u5_n2943 ), .A3(_u10_u5_n2944 ), .ZN(_u10_u5_n2919 ) );
NOR2_X1 _u10_u5_U769  ( .A1(_u10_u5_n2423 ), .A2(1'b0), .ZN(_u10_u5_n1979 ));
NAND3_X1 _u10_u5_U768  ( .A1(_u10_u5_n2549 ), .A2(_u10_u5_n1936 ), .A3(_u10_u5_n1979 ), .ZN(_u10_u5_n2328 ) );
INV_X1 _u10_u5_U767  ( .A(_u10_u5_n2328 ), .ZN(_u10_u5_n2554 ) );
NAND3_X1 _u10_u5_U766  ( .A1(_u10_u5_n2941 ), .A2(_u10_u5_n2446 ), .A3(_u10_u5_n2554 ), .ZN(_u10_u5_n2115 ) );
NOR2_X1 _u10_u5_U765  ( .A1(_u10_u5_n2578 ), .A2(_u10_u5_n2030 ), .ZN(_u10_u5_n2553 ) );
INV_X1 _u10_u5_U764  ( .A(_u10_u5_n2553 ), .ZN(_u10_u5_n2269 ) );
NOR2_X1 _u10_u5_U763  ( .A1(_u10_u5_n2269 ), .A2(_u10_u5_n2790 ), .ZN(_u10_u5_n2657 ) );
INV_X1 _u10_u5_U762  ( .A(_u10_u5_n2657 ), .ZN(_u10_u5_n2210 ) );
NOR2_X1 _u10_u5_U761  ( .A1(_u10_u5_n2210 ), .A2(_u10_u5_n2911 ), .ZN(_u10_u5_n2213 ) );
INV_X1 _u10_u5_U760  ( .A(_u10_u5_n2213 ), .ZN(_u10_u5_n2456 ) );
NAND2_X1 _u10_u5_U759  ( .A1(_u10_u5_n2115 ), .A2(_u10_u5_n2456 ), .ZN(_u10_u5_n2634 ) );
INV_X1 _u10_u5_U758  ( .A(_u10_u5_n2634 ), .ZN(_u10_u5_n2220 ) );
NOR2_X1 _u10_u5_U757  ( .A1(_u10_u5_n2081 ), .A2(_u10_u5_n2386 ), .ZN(_u10_u5_n2131 ) );
NAND2_X1 _u10_u5_U756  ( .A1(_u10_u5_n2940 ), .A2(_u10_u5_n2131 ), .ZN(_u10_u5_n2138 ) );
INV_X1 _u10_u5_U755  ( .A(_u10_u5_n2138 ), .ZN(_u10_u5_n2927 ) );
NAND2_X1 _u10_u5_U754  ( .A1(_u10_u5_n2220 ), .A2(_u10_u5_n2927 ), .ZN(_u10_u5_n2939 ) );
NAND2_X1 _u10_u5_U753  ( .A1(_u10_u5_n1885 ), .A2(_u10_u5_n2939 ), .ZN(_u10_u5_n2931 ) );
NAND3_X1 _u10_u5_U752  ( .A1(_u10_u5_n1859 ), .A2(_u10_u5_n2365 ), .A3(_u10_u5_n2938 ), .ZN(_u10_u5_n2935 ) );
NAND3_X1 _u10_u5_U751  ( .A1(_u10_u5_n2927 ), .A2(_u10_u5_n2937 ), .A3(_u10_u5_n2220 ), .ZN(_u10_u5_n2936 ) );
NAND2_X1 _u10_u5_U750  ( .A1(_u10_u5_n2935 ), .A2(_u10_u5_n2936 ), .ZN(_u10_u5_n2932 ) );
INV_X1 _u10_u5_U749  ( .A(_u10_u5_n1937 ), .ZN(_u10_u5_n2350 ) );
NAND2_X1 _u10_u5_U748  ( .A1(_u10_u5_n1913 ), .A2(_u10_u5_n2350 ), .ZN(_u10_u5_n2934 ) );
NAND2_X1 _u10_u5_U747  ( .A1(_u10_u5_n2386 ), .A2(_u10_u5_n2934 ), .ZN(_u10_u5_n2933 ) );
NAND3_X1 _u10_u5_U746  ( .A1(_u10_u5_n2931 ), .A2(_u10_u5_n2932 ), .A3(_u10_u5_n2933 ), .ZN(_u10_u5_n2921 ) );
OR2_X1 _u10_u5_U745  ( .A1(_u10_u5_n2213 ), .A2(_u10_u5_n2386 ), .ZN(_u10_u5_n2930 ) );
NAND2_X1 _u10_u5_U744  ( .A1(_u10_u5_n2049 ), .A2(_u10_u5_n2930 ), .ZN(_u10_u5_n2228 ) );
AND2_X1 _u10_u5_U743  ( .A1(_u10_u5_n2228 ), .A2(_u10_u5_n2699 ), .ZN(_u10_u5_n2929 ) );
NOR2_X1 _u10_u5_U742  ( .A1(_u10_u5_n2929 ), .A2(_u10_u5_n2495 ), .ZN(_u10_u5_n2922 ) );
NOR2_X1 _u10_u5_U741  ( .A1(_u10_u5_n2633 ), .A2(_u10_u5_n2877 ), .ZN(_u10_u5_n2928 ) );
NOR2_X1 _u10_u5_U740  ( .A1(_u10_u5_n2928 ), .A2(_u10_u5_n2886 ), .ZN(_u10_u5_n2923 ) );
NOR2_X1 _u10_u5_U739  ( .A1(_u10_u5_n2927 ), .A2(_u10_u5_n2531 ), .ZN(_u10_u5_n2926 ) );
NOR2_X1 _u10_u5_U738  ( .A1(_u10_u5_n2926 ), .A2(_u10_u5_n2687 ), .ZN(_u10_u5_n2925 ) );
NOR2_X1 _u10_u5_U737  ( .A1(_u10_u5_n2925 ), .A2(_u10_u5_n1849 ), .ZN(_u10_u5_n2924 ) );
NOR4_X1 _u10_u5_U736  ( .A1(_u10_u5_n2921 ), .A2(_u10_u5_n2922 ), .A3(_u10_u5_n2923 ), .A4(_u10_u5_n2924 ), .ZN(_u10_u5_n2920 ) );
NAND4_X1 _u10_u5_U735  ( .A1(_u10_u5_n2917 ), .A2(_u10_u5_n2918 ), .A3(_u10_u5_n2919 ), .A4(_u10_u5_n2920 ), .ZN(_u10_u5_n2312 ) );
NOR2_X1 _u10_u5_U734  ( .A1(_u10_u5_n2600 ), .A2(_u10_u5_n2686 ), .ZN(_u10_u5_n2401 ) );
NAND2_X1 _u10_u5_U733  ( .A1(_u10_u5_n2401 ), .A2(_u10_u5_n2549 ), .ZN(_u10_u5_n2547 ) );
INV_X1 _u10_u5_U732  ( .A(_u10_u5_n2547 ), .ZN(_u10_u5_n2794 ) );
NAND3_X1 _u10_u5_U731  ( .A1(_u10_u5_n2364 ), .A2(_u10_u5_n2667 ), .A3(_u10_u5_n2794 ), .ZN(_u10_u5_n2535 ) );
INV_X1 _u10_u5_U730  ( .A(_u10_u5_n2535 ), .ZN(_u10_u5_n2586 ) );
NAND2_X1 _u10_u5_U729  ( .A1(_u10_u5_n2586 ), .A2(_u10_u5_n2571 ), .ZN(_u10_u5_n2916 ) );
NAND2_X1 _u10_u5_U728  ( .A1(_u10_u5_n2837 ), .A2(_u10_u5_n2916 ), .ZN(_u10_u5_n2436 ) );
NAND2_X1 _u10_u5_U727  ( .A1(_u10_u5_n2915 ), .A2(_u10_u5_n2571 ), .ZN(_u10_u5_n2914 ) );
NAND2_X1 _u10_u5_U726  ( .A1(_u10_u5_n2166 ), .A2(_u10_u5_n2914 ), .ZN(_u10_u5_n2017 ) );
NOR2_X1 _u10_u5_U725  ( .A1(_u10_u5_n2485 ), .A2(_u10_u5_n1841 ), .ZN(_u10_u5_n2913 ) );
OR4_X1 _u10_u5_U724  ( .A1(_u10_u5_n2436 ), .A2(_u10_u5_n2017 ), .A3(_u10_u5_n2913 ), .A4(_u10_u5_n2442 ), .ZN(_u10_u5_n2912 ) );
NAND2_X1 _u10_u5_U723  ( .A1(_u10_u5_n2709 ), .A2(_u10_u5_n2912 ), .ZN(_u10_u5_n2888 ) );
NAND3_X1 _u10_u5_U722  ( .A1(_u10_u5_n2078 ), .A2(_u10_u5_n2031 ), .A3(1'b0),.ZN(_u10_u5_n2580 ) );
INV_X1 _u10_u5_U721  ( .A(_u10_u5_n2580 ), .ZN(_u10_u5_n2680 ) );
AND2_X1 _u10_u5_U720  ( .A1(_u10_u5_n2680 ), .A2(_u10_u5_n2668 ), .ZN(_u10_u5_n1950 ) );
NAND2_X1 _u10_u5_U719  ( .A1(_u10_u5_n1950 ), .A2(_u10_u5_n2089 ), .ZN(_u10_u5_n2095 ) );
INV_X1 _u10_u5_U718  ( .A(_u10_u5_n2095 ), .ZN(_u10_u5_n2542 ) );
NAND2_X1 _u10_u5_U717  ( .A1(_u10_u5_n2542 ), .A2(_u10_u5_n2446 ), .ZN(_u10_u5_n1887 ) );
NOR2_X1 _u10_u5_U716  ( .A1(_u10_u5_n1887 ), .A2(_u10_u5_n2911 ), .ZN(_u10_u5_n2114 ) );
INV_X1 _u10_u5_U715  ( .A(_u10_u5_n2114 ), .ZN(_u10_u5_n1940 ) );
NAND3_X1 _u10_u5_U714  ( .A1(_u10_u5_n2535 ), .A2(_u10_u5_n1940 ), .A3(_u10_u5_n2910 ), .ZN(_u10_u5_n2524 ) );
NAND2_X1 _u10_u5_U713  ( .A1(_u10_u5_n2524 ), .A2(_u10_u5_n2488 ), .ZN(_u10_u5_n2889 ) );
NAND2_X1 _u10_u5_U712  ( .A1(_u10_u5_n2220 ), .A2(_u10_u5_n1940 ), .ZN(_u10_u5_n2763 ) );
NOR2_X1 _u10_u5_U711  ( .A1(_u10_u5_n2763 ), .A2(_u10_u5_n2586 ), .ZN(_u10_u5_n2808 ) );
NOR2_X1 _u10_u5_U710  ( .A1(_u10_u5_n2808 ), .A2(_u10_u5_n2350 ), .ZN(_u10_u5_n2908 ) );
NOR2_X1 _u10_u5_U709  ( .A1(_u10_u5_n2544 ), .A2(_u10_u5_n1950 ), .ZN(_u10_u5_n2899 ) );
NOR2_X1 _u10_u5_U708  ( .A1(_u10_u5_n2899 ), .A2(_u10_u5_n2159 ), .ZN(_u10_u5_n2909 ) );
NOR2_X1 _u10_u5_U707  ( .A1(_u10_u5_n2908 ), .A2(_u10_u5_n2909 ), .ZN(_u10_u5_n2890 ) );
NOR3_X1 _u10_u5_U706  ( .A1(_u10_u5_n2547 ), .A2(_u10_u5_n1846 ), .A3(_u10_u5_n2907 ), .ZN(_u10_u5_n2892 ) );
NOR3_X1 _u10_u5_U705  ( .A1(_u10_u5_n2240 ), .A2(_u10_u5_n2377 ), .A3(_u10_u5_n1911 ), .ZN(_u10_u5_n2906 ) );
NOR2_X1 _u10_u5_U704  ( .A1(_u10_u5_n2906 ), .A2(_u10_u5_n2535 ), .ZN(_u10_u5_n2893 ) );
NAND2_X1 _u10_u5_U703  ( .A1(_u10_u5_n2554 ), .A2(_u10_u5_n2446 ), .ZN(_u10_u5_n2903 ) );
AND3_X1 _u10_u5_U702  ( .A1(_u10_u5_n2210 ), .A2(_u10_u5_n2905 ), .A3(_u10_u5_n1887 ), .ZN(_u10_u5_n2904 ) );
NAND4_X1 _u10_u5_U701  ( .A1(_u10_u5_n2902 ), .A2(_u10_u5_n2498 ), .A3(_u10_u5_n2903 ), .A4(_u10_u5_n2904 ), .ZN(_u10_u5_n2788 ) );
INV_X1 _u10_u5_U700  ( .A(_u10_u5_n2788 ), .ZN(_u10_u5_n2901 ) );
NOR2_X1 _u10_u5_U699  ( .A1(_u10_u5_n2901 ), .A2(_u10_u5_n1888 ), .ZN(_u10_u5_n2894 ) );
NOR2_X1 _u10_u5_U698  ( .A1(_u10_u5_n2401 ), .A2(_u10_u5_n2553 ), .ZN(_u10_u5_n2900 ) );
NOR2_X1 _u10_u5_U697  ( .A1(_u10_u5_n2900 ), .A2(_u10_u5_n1954 ), .ZN(_u10_u5_n2897 ) );
NOR2_X1 _u10_u5_U696  ( .A1(1'b0), .A2(_u10_u5_n2899 ), .ZN(_u10_u5_n2898 ));
NOR2_X1 _u10_u5_U695  ( .A1(_u10_u5_n2897 ), .A2(_u10_u5_n2898 ), .ZN(_u10_u5_n2896 ) );
NOR2_X1 _u10_u5_U694  ( .A1(_u10_u5_n2896 ), .A2(_u10_u5_n1843 ), .ZN(_u10_u5_n2895 ) );
NOR4_X1 _u10_u5_U693  ( .A1(_u10_u5_n2892 ), .A2(_u10_u5_n2893 ), .A3(_u10_u5_n2894 ), .A4(_u10_u5_n2895 ), .ZN(_u10_u5_n2891 ) );
NAND4_X1 _u10_u5_U692  ( .A1(_u10_u5_n2888 ), .A2(_u10_u5_n2889 ), .A3(_u10_u5_n2890 ), .A4(_u10_u5_n2891 ), .ZN(_u10_u5_n2610 ) );
NOR4_X1 _u10_u5_U691  ( .A1(_u10_u5_n2670 ), .A2(_u10_u5_n2312 ), .A3(_u10_u5_n2610 ), .A4(_u10_u5_n2887 ), .ZN(_u10_u5_n2724 ) );
NOR2_X1 _u10_u5_U690  ( .A1(_u10_u5_n2883 ), .A2(_u10_u5_n2535 ), .ZN(_u10_u5_n2861 ) );
NOR2_X1 _u10_u5_U689  ( .A1(_u10_u5_n1855 ), .A2(_u10_u5_n1869 ), .ZN(_u10_u5_n2862 ) );
NOR2_X1 _u10_u5_U688  ( .A1(_u10_u5_n2886 ), .A2(_u10_u5_n2695 ), .ZN(_u10_u5_n2863 ) );
NAND2_X1 _u10_u5_U687  ( .A1(_u10_u5_n2813 ), .A2(_u10_u5_n2885 ), .ZN(_u10_u5_n2864 ) );
NAND2_X1 _u10_u5_U686  ( .A1(_u10_u5_n2114 ), .A2(_u10_u5_n2884 ), .ZN(_u10_u5_n2865 ) );
NAND2_X1 _u10_u5_U685  ( .A1(1'b0), .A2(_u10_u5_n2667 ), .ZN(_u10_u5_n2112 ));
NOR3_X1 _u10_u5_U684  ( .A1(_u10_u5_n2883 ), .A2(_u10_u5_n2112 ), .A3(_u10_u5_n2719 ), .ZN(_u10_u5_n2878 ) );
INV_X1 _u10_u5_U683  ( .A(_u10_u5_n2112 ), .ZN(_u10_u5_n1856 ) );
NAND2_X1 _u10_u5_U682  ( .A1(_u10_u5_n2364 ), .A2(_u10_u5_n1856 ), .ZN(_u10_u5_n2882 ) );
NAND2_X1 _u10_u5_U681  ( .A1(_u10_u5_n2882 ), .A2(_u10_u5_n1869 ), .ZN(_u10_u5_n2050 ) );
INV_X1 _u10_u5_U680  ( .A(_u10_u5_n2050 ), .ZN(_u10_u5_n1939 ) );
NOR2_X1 _u10_u5_U679  ( .A1(_u10_u5_n1939 ), .A2(_u10_u5_n1841 ), .ZN(_u10_u5_n2881 ) );
NOR2_X1 _u10_u5_U678  ( .A1(_u10_u5_n2881 ), .A2(_u10_u5_n2840 ), .ZN(_u10_u5_n2880 ) );
NOR2_X1 _u10_u5_U677  ( .A1(_u10_u5_n2880 ), .A2(_u10_u5_n1836 ), .ZN(_u10_u5_n2879 ) );
NOR2_X1 _u10_u5_U676  ( .A1(_u10_u5_n2878 ), .A2(_u10_u5_n2879 ), .ZN(_u10_u5_n2866 ) );
NOR2_X1 _u10_u5_U675  ( .A1(_u10_u5_n2081 ), .A2(_u10_u5_n2877 ), .ZN(_u10_u5_n1840 ) );
NAND2_X1 _u10_u5_U674  ( .A1(_u10_u5_n1840 ), .A2(_u10_u5_n2115 ), .ZN(_u10_u5_n1873 ) );
NAND2_X1 _u10_u5_U673  ( .A1(_u10_u5_n2695 ), .A2(_u10_u5_n1940 ), .ZN(_u10_u5_n1874 ) );
NOR3_X1 _u10_u5_U672  ( .A1(_u10_u5_n2050 ), .A2(_u10_u5_n1873 ), .A3(_u10_u5_n1874 ), .ZN(_u10_u5_n2876 ) );
NOR2_X1 _u10_u5_U671  ( .A1(_u10_u5_n2876 ), .A2(_u10_u5_n1913 ), .ZN(_u10_u5_n2868 ) );
NAND2_X1 _u10_u5_U670  ( .A1(_u10_u5_n2875 ), .A2(_u10_u5_n2466 ), .ZN(_u10_u5_n2872 ) );
INV_X1 _u10_u5_U669  ( .A(_u10_u5_n1979 ), .ZN(_u10_u5_n2746 ) );
NAND2_X1 _u10_u5_U668  ( .A1(_u10_u5_n2874 ), .A2(_u10_u5_n2746 ), .ZN(_u10_u5_n1935 ) );
NAND3_X1 _u10_u5_U667  ( .A1(_u10_u5_n1935 ), .A2(_u10_u5_n1936 ), .A3(_u10_u5_n2467 ), .ZN(_u10_u5_n2873 ) );
NAND2_X1 _u10_u5_U666  ( .A1(_u10_u5_n2872 ), .A2(_u10_u5_n2873 ), .ZN(_u10_u5_n2264 ) );
AND2_X1 _u10_u5_U665  ( .A1(_u10_u5_n2264 ), .A2(_u10_u5_n2461 ), .ZN(_u10_u5_n2869 ) );
AND2_X1 _u10_u5_U664  ( .A1(_u10_u5_n1966 ), .A2(_u10_u5_n2761 ), .ZN(_u10_u5_n2870 ) );
NOR2_X1 _u10_u5_U663  ( .A1(_u10_u5_n2159 ), .A2(_u10_u5_n2163 ), .ZN(_u10_u5_n2871 ) );
NOR4_X1 _u10_u5_U662  ( .A1(_u10_u5_n2868 ), .A2(_u10_u5_n2869 ), .A3(_u10_u5_n2870 ), .A4(_u10_u5_n2871 ), .ZN(_u10_u5_n2867 ) );
NAND4_X1 _u10_u5_U661  ( .A1(_u10_u5_n2864 ), .A2(_u10_u5_n2865 ), .A3(_u10_u5_n2866 ), .A4(_u10_u5_n2867 ), .ZN(_u10_u5_n1992 ) );
NOR4_X1 _u10_u5_U660  ( .A1(_u10_u5_n2861 ), .A2(_u10_u5_n2862 ), .A3(_u10_u5_n2863 ), .A4(_u10_u5_n1992 ), .ZN(_u10_u5_n2725 ) );
NAND2_X1 _u10_u5_U659  ( .A1(_u10_u5_n2364 ), .A2(_u10_u5_n1846 ), .ZN(_u10_u5_n2744 ) );
NAND4_X1 _u10_u5_U658  ( .A1(_u10_u5_n2765 ), .A2(_u10_u5_n1939 ), .A3(_u10_u5_n2744 ), .A4(_u10_u5_n2535 ), .ZN(_u10_u5_n2860 ) );
NAND2_X1 _u10_u5_U657  ( .A1(_u10_u5_n2049 ), .A2(_u10_u5_n2860 ), .ZN(_u10_u5_n2856 ) );
NOR4_X1 _u10_u5_U656  ( .A1(1'b0), .A2(_u10_u5_n2858 ), .A3(_u10_u5_n2859 ),.A4(_u10_u5_n2051 ), .ZN(_u10_u5_n2857 ) );
NAND4_X1 _u10_u5_U655  ( .A1(_u10_u5_n2228 ), .A2(_u10_u5_n2855 ), .A3(_u10_u5_n2856 ), .A4(_u10_u5_n2857 ), .ZN(_u10_u5_n2854 ) );
NAND2_X1 _u10_u5_U654  ( .A1(_u10_u5_n2043 ), .A2(_u10_u5_n2854 ), .ZN(_u10_u5_n2821 ) );
INV_X1 _u10_u5_U653  ( .A(_u10_u5_n2071 ), .ZN(_u10_u5_n2279 ) );
INV_X1 _u10_u5_U652  ( .A(_u10_u5_n2599 ), .ZN(_u10_u5_n2357 ) );
OR2_X1 _u10_u5_U651  ( .A1(_u10_u5_n2744 ), .A2(_u10_u5_n2853 ), .ZN(_u10_u5_n2844 ) );
NAND2_X1 _u10_u5_U650  ( .A1(_u10_u5_n2131 ), .A2(_u10_u5_n2852 ), .ZN(_u10_u5_n2851 ) );
NAND2_X1 _u10_u5_U649  ( .A1(_u10_u5_n2082 ), .A2(_u10_u5_n2851 ), .ZN(_u10_u5_n2848 ) );
NAND2_X1 _u10_u5_U648  ( .A1(_u10_u5_n2850 ), .A2(_u10_u5_n2600 ), .ZN(_u10_u5_n2849 ) );
NAND3_X1 _u10_u5_U647  ( .A1(_u10_u5_n2848 ), .A2(_u10_u5_n2077 ), .A3(_u10_u5_n2849 ), .ZN(_u10_u5_n2287 ) );
NAND2_X1 _u10_u5_U646  ( .A1(_u10_u5_n2082 ), .A2(_u10_u5_n2050 ), .ZN(_u10_u5_n2847 ) );
NAND2_X1 _u10_u5_U645  ( .A1(_u10_u5_n2846 ), .A2(_u10_u5_n2847 ), .ZN(_u10_u5_n2074 ) );
NOR3_X1 _u10_u5_U644  ( .A1(_u10_u5_n2287 ), .A2(_u10_u5_n2596 ), .A3(_u10_u5_n2074 ), .ZN(_u10_u5_n2845 ) );
NAND4_X1 _u10_u5_U643  ( .A1(_u10_u5_n2357 ), .A2(_u10_u5_n2837 ), .A3(_u10_u5_n2844 ), .A4(_u10_u5_n2845 ), .ZN(_u10_u5_n2843 ) );
NAND2_X1 _u10_u5_U642  ( .A1(_u10_u5_n2279 ), .A2(_u10_u5_n2843 ), .ZN(_u10_u5_n2822 ) );
NOR3_X1 _u10_u5_U641  ( .A1(_u10_u5_n1925 ), .A2(_u10_u5_n2842 ), .A3(_u10_u5_n2686 ), .ZN(_u10_u5_n2841 ) );
NOR3_X1 _u10_u5_U640  ( .A1(_u10_u5_n2840 ), .A2(_u10_u5_n2599 ), .A3(_u10_u5_n2841 ), .ZN(_u10_u5_n2839 ) );
AND4_X1 _u10_u5_U639  ( .A1(_u10_u5_n2836 ), .A2(_u10_u5_n2837 ), .A3(_u10_u5_n2838 ), .A4(_u10_u5_n2839 ), .ZN(_u10_u5_n2454 ) );
NOR2_X1 _u10_u5_U638  ( .A1(_u10_u5_n2719 ), .A2(_u10_u5_n2835 ), .ZN(_u10_u5_n2773 ) );
NOR2_X1 _u10_u5_U637  ( .A1(_u10_u5_n2138 ), .A2(_u10_u5_n2773 ), .ZN(_u10_u5_n2814 ) );
NAND2_X1 _u10_u5_U636  ( .A1(_u10_u5_n2814 ), .A2(_u10_u5_n1869 ), .ZN(_u10_u5_n2834 ) );
NAND2_X1 _u10_u5_U635  ( .A1(_u10_u5_n2833 ), .A2(_u10_u5_n2834 ), .ZN(_u10_u5_n2832 ) );
NAND2_X1 _u10_u5_U634  ( .A1(_u10_u5_n2454 ), .A2(_u10_u5_n2832 ), .ZN(_u10_u5_n2831 ) );
NAND2_X1 _u10_u5_U633  ( .A1(_u10_u5_n2830 ), .A2(_u10_u5_n2831 ), .ZN(_u10_u5_n2823 ) );
INV_X1 _u10_u5_U632  ( .A(_u10_u5_n2025 ), .ZN(_u10_u5_n2470 ) );
NAND2_X1 _u10_u5_U631  ( .A1(_u10_u5_n1979 ), .A2(_u10_u5_n1936 ), .ZN(_u10_u5_n2829 ) );
AND2_X1 _u10_u5_U630  ( .A1(_u10_u5_n2828 ), .A2(_u10_u5_n2829 ), .ZN(_u10_u5_n2469 ) );
NAND2_X1 _u10_u5_U629  ( .A1(_u10_u5_n2469 ), .A2(_u10_u5_n2269 ), .ZN(_u10_u5_n2161 ) );
INV_X1 _u10_u5_U628  ( .A(_u10_u5_n2161 ), .ZN(_u10_u5_n2276 ) );
NOR2_X1 _u10_u5_U627  ( .A1(_u10_u5_n2274 ), .A2(_u10_u5_n2719 ), .ZN(_u10_u5_n2827 ) );
NOR3_X1 _u10_u5_U626  ( .A1(_u10_u5_n2827 ), .A2(_u10_u5_n2742 ), .A3(_u10_u5_n2680 ), .ZN(_u10_u5_n2826 ) );
NAND3_X1 _u10_u5_U625  ( .A1(_u10_u5_n2276 ), .A2(_u10_u5_n2108 ), .A3(_u10_u5_n2826 ), .ZN(_u10_u5_n2825 ) );
NAND2_X1 _u10_u5_U624  ( .A1(_u10_u5_n2470 ), .A2(_u10_u5_n2825 ), .ZN(_u10_u5_n2824 ) );
NAND4_X1 _u10_u5_U623  ( .A1(_u10_u5_n2821 ), .A2(_u10_u5_n2822 ), .A3(_u10_u5_n2823 ), .A4(_u10_u5_n2824 ), .ZN(_u10_u5_n2804 ) );
NAND2_X1 _u10_u5_U622  ( .A1(_u10_u5_n2131 ), .A2(_u10_u5_n2744 ), .ZN(_u10_u5_n2820 ) );
NAND2_X1 _u10_u5_U621  ( .A1(_u10_u5_n2571 ), .A2(_u10_u5_n2820 ), .ZN(_u10_u5_n2817 ) );
NOR2_X1 _u10_u5_U620  ( .A1(_u10_u5_n2819 ), .A2(_u10_u5_n2436 ), .ZN(_u10_u5_n2818 ) );
NAND4_X1 _u10_u5_U619  ( .A1(_u10_u5_n2437 ), .A2(_u10_u5_n2355 ), .A3(_u10_u5_n2817 ), .A4(_u10_u5_n2818 ), .ZN(_u10_u5_n2816 ) );
NAND2_X1 _u10_u5_U618  ( .A1(_u10_u5_n2815 ), .A2(_u10_u5_n2816 ), .ZN(_u10_u5_n2809 ) );
INV_X1 _u10_u5_U617  ( .A(_u10_u5_n2814 ), .ZN(_u10_u5_n2812 ) );
OR2_X1 _u10_u5_U616  ( .A1(_u10_u5_n1911 ), .A2(_u10_u5_n2813 ), .ZN(_u10_u5_n1884 ) );
NAND2_X1 _u10_u5_U615  ( .A1(_u10_u5_n2812 ), .A2(_u10_u5_n1884 ), .ZN(_u10_u5_n2810 ) );
NOR2_X1 _u10_u5_U614  ( .A1(_u10_u5_n1894 ), .A2(_u10_u5_n2461 ), .ZN(_u10_u5_n1948 ) );
OR2_X1 _u10_u5_U613  ( .A1(_u10_u5_n1847 ), .A2(_u10_u5_n1948 ), .ZN(_u10_u5_n2811 ) );
NAND3_X1 _u10_u5_U612  ( .A1(_u10_u5_n2809 ), .A2(_u10_u5_n2810 ), .A3(_u10_u5_n2811 ), .ZN(_u10_u5_n2805 ) );
NOR2_X1 _u10_u5_U611  ( .A1(_u10_u5_n2808 ), .A2(_u10_u5_n2775 ), .ZN(_u10_u5_n2806 ) );
AND2_X1 _u10_u5_U610  ( .A1(_u10_u5_n2721 ), .A2(_u10_u5_n1911 ), .ZN(_u10_u5_n2807 ) );
NOR4_X1 _u10_u5_U609  ( .A1(_u10_u5_n2804 ), .A2(_u10_u5_n2805 ), .A3(_u10_u5_n2806 ), .A4(_u10_u5_n2807 ), .ZN(_u10_u5_n2726 ) );
NAND2_X1 _u10_u5_U608  ( .A1(_u10_u5_n2803 ), .A2(_u10_u5_n2112 ), .ZN(_u10_u5_n2802 ) );
NAND2_X1 _u10_u5_U607  ( .A1(_u10_u5_n2364 ), .A2(_u10_u5_n2802 ), .ZN(_u10_u5_n2801 ) );
NAND2_X1 _u10_u5_U606  ( .A1(_u10_u5_n2800 ), .A2(_u10_u5_n2801 ), .ZN(_u10_u5_n2799 ) );
NAND2_X1 _u10_u5_U605  ( .A1(_u10_u5_n1937 ), .A2(_u10_u5_n2799 ), .ZN(_u10_u5_n2780 ) );
NAND2_X1 _u10_u5_U604  ( .A1(_u10_u5_n2775 ), .A2(_u10_u5_n2798 ), .ZN(_u10_u5_n2796 ) );
INV_X1 _u10_u5_U603  ( .A(_u10_u5_n2131 ), .ZN(_u10_u5_n2797 ) );
NAND2_X1 _u10_u5_U602  ( .A1(_u10_u5_n2796 ), .A2(_u10_u5_n2797 ), .ZN(_u10_u5_n2781 ) );
OR4_X1 _u10_u5_U601  ( .A1(_u10_u5_n2795 ), .A2(_u10_u5_n2303 ), .A3(_u10_u5_n2553 ), .A4(_u10_u5_n2554 ), .ZN(_u10_u5_n2792 ) );
NAND3_X1 _u10_u5_U600  ( .A1(_u10_u5_n1847 ), .A2(_u10_u5_n2097 ), .A3(_u10_u5_n2096 ), .ZN(_u10_u5_n2793 ) );
NOR4_X1 _u10_u5_U599  ( .A1(_u10_u5_n2792 ), .A2(_u10_u5_n2793 ), .A3(_u10_u5_n2542 ), .A4(_u10_u5_n2794 ), .ZN(_u10_u5_n2791 ) );
NOR2_X1 _u10_u5_U598  ( .A1(_u10_u5_n2791 ), .A2(_u10_u5_n2085 ), .ZN(_u10_u5_n2783 ) );
NAND2_X1 _u10_u5_U597  ( .A1(_u10_u5_n2114 ), .A2(_u10_u5_n2049 ), .ZN(_u10_u5_n2700 ) );
INV_X1 _u10_u5_U596  ( .A(_u10_u5_n2700 ), .ZN(_u10_u5_n2784 ) );
NAND4_X1 _u10_u5_U595  ( .A1(_u10_u5_n2001 ), .A2(_u10_u5_n2547 ), .A3(_u10_u5_n2368 ), .A4(_u10_u5_n1847 ), .ZN(_u10_u5_n2787 ) );
NOR4_X1 _u10_u5_U594  ( .A1(_u10_u5_n2787 ), .A2(_u10_u5_n2788 ), .A3(_u10_u5_n2789 ), .A4(_u10_u5_n2790 ), .ZN(_u10_u5_n2786 ) );
NOR2_X1 _u10_u5_U593  ( .A1(_u10_u5_n2786 ), .A2(_u10_u5_n2000 ), .ZN(_u10_u5_n2785 ) );
NOR3_X1 _u10_u5_U592  ( .A1(_u10_u5_n2783 ), .A2(_u10_u5_n2784 ), .A3(_u10_u5_n2785 ), .ZN(_u10_u5_n2782 ) );
NAND3_X1 _u10_u5_U591  ( .A1(_u10_u5_n2780 ), .A2(_u10_u5_n2781 ), .A3(_u10_u5_n2782 ), .ZN(_u10_u5_n2728 ) );
OR3_X1 _u10_u5_U590  ( .A1(_u10_u5_n2138 ), .A2(_u10_u5_n2633 ), .A3(_u10_u5_n2779 ), .ZN(_u10_u5_n2778 ) );
NAND2_X1 _u10_u5_U589  ( .A1(_u10_u5_n2777 ), .A2(_u10_u5_n2778 ), .ZN(_u10_u5_n2767 ) );
NAND3_X1 _u10_u5_U588  ( .A1(_u10_u5_n2775 ), .A2(_u10_u5_n2083 ), .A3(_u10_u5_n2776 ), .ZN(_u10_u5_n2774 ) );
NAND2_X1 _u10_u5_U587  ( .A1(_u10_u5_n2773 ), .A2(_u10_u5_n2774 ), .ZN(_u10_u5_n2768 ) );
NAND2_X1 _u10_u5_U586  ( .A1(_u10_u5_n2218 ), .A2(_u10_u5_n2772 ), .ZN(_u10_u5_n2769 ) );
NAND2_X1 _u10_u5_U585  ( .A1(_u10_u5_n2302 ), .A2(_u10_u5_n2467 ), .ZN(_u10_u5_n2771 ) );
NAND2_X1 _u10_u5_U584  ( .A1(_u10_u5_n2461 ), .A2(_u10_u5_n2771 ), .ZN(_u10_u5_n2770 ) );
NAND4_X1 _u10_u5_U583  ( .A1(_u10_u5_n2767 ), .A2(_u10_u5_n2768 ), .A3(_u10_u5_n2769 ), .A4(_u10_u5_n2770 ), .ZN(_u10_u5_n2729 ) );
NAND3_X1 _u10_u5_U582  ( .A1(_u10_u5_n2668 ), .A2(_u10_u5_n2600 ), .A3(_u10_u5_n2276 ), .ZN(_u10_u5_n2766 ) );
NAND2_X1 _u10_u5_U581  ( .A1(_u10_u5_n1894 ), .A2(_u10_u5_n2766 ), .ZN(_u10_u5_n2753 ) );
NAND3_X1 _u10_u5_U580  ( .A1(_u10_u5_n2456 ), .A2(_u10_u5_n2744 ), .A3(_u10_u5_n2765 ), .ZN(_u10_u5_n2764 ) );
NAND2_X1 _u10_u5_U579  ( .A1(_u10_u5_n2377 ), .A2(_u10_u5_n2764 ), .ZN(_u10_u5_n2754 ) );
NAND2_X1 _u10_u5_U578  ( .A1(_u10_u5_n2763 ), .A2(_u10_u5_n2007 ), .ZN(_u10_u5_n2755 ) );
NOR2_X1 _u10_u5_U577  ( .A1(_u10_u5_n2531 ), .A2(_u10_u5_n2744 ), .ZN(_u10_u5_n2760 ) );
INV_X1 _u10_u5_U576  ( .A(_u10_u5_n2762 ), .ZN(_u10_u5_n2189 ) );
NOR3_X1 _u10_u5_U575  ( .A1(_u10_u5_n2760 ), .A2(_u10_u5_n2761 ), .A3(_u10_u5_n2189 ), .ZN(_u10_u5_n2759 ) );
NOR2_X1 _u10_u5_U574  ( .A1(_u10_u5_n2759 ), .A2(_u10_u5_n1849 ), .ZN(_u10_u5_n2757 ) );
NOR2_X1 _u10_u5_U573  ( .A1(_u10_u5_n1817 ), .A2(_u10_u5_n2665 ), .ZN(_u10_u5_n2758 ) );
NOR2_X1 _u10_u5_U572  ( .A1(_u10_u5_n2757 ), .A2(_u10_u5_n2758 ), .ZN(_u10_u5_n2756 ) );
NAND4_X1 _u10_u5_U571  ( .A1(_u10_u5_n2753 ), .A2(_u10_u5_n2754 ), .A3(_u10_u5_n2755 ), .A4(_u10_u5_n2756 ), .ZN(_u10_u5_n2730 ) );
INV_X1 _u10_u5_U570  ( .A(_u10_u5_n2359 ), .ZN(_u10_u5_n1899 ) );
NAND4_X1 _u10_u5_U569  ( .A1(_u10_u5_n2078 ), .A2(_u10_u5_n2580 ), .A3(_u10_u5_n2748 ), .A4(_u10_u5_n2752 ), .ZN(_u10_u5_n2751 ) );
NAND2_X1 _u10_u5_U568  ( .A1(_u10_u5_n1899 ), .A2(_u10_u5_n2751 ), .ZN(_u10_u5_n2732 ) );
INV_X1 _u10_u5_U567  ( .A(_u10_u5_n2750 ), .ZN(_u10_u5_n2379 ) );
NAND3_X1 _u10_u5_U566  ( .A1(_u10_u5_n1856 ), .A2(_u10_u5_n2669 ), .A3(_u10_u5_n2364 ), .ZN(_u10_u5_n2749 ) );
AND2_X1 _u10_u5_U565  ( .A1(_u10_u5_n2748 ), .A2(_u10_u5_n2749 ), .ZN(_u10_u5_n2034 ) );
NAND2_X1 _u10_u5_U564  ( .A1(_u10_u5_n2105 ), .A2(_u10_u5_n2669 ), .ZN(_u10_u5_n2745 ) );
AND3_X1 _u10_u5_U563  ( .A1(_u10_u5_n2745 ), .A2(_u10_u5_n2746 ), .A3(_u10_u5_n2747 ), .ZN(_u10_u5_n2380 ) );
NOR2_X1 _u10_u5_U562  ( .A1(_u10_u5_n2274 ), .A2(_u10_u5_n2744 ), .ZN(_u10_u5_n2743 ) );
NOR4_X1 _u10_u5_U561  ( .A1(_u10_u5_n2742 ), .A2(_u10_u5_n2680 ), .A3(_u10_u5_n2743 ), .A4(_u10_u5_n2428 ), .ZN(_u10_u5_n2741 ) );
NAND4_X1 _u10_u5_U560  ( .A1(_u10_u5_n2379 ), .A2(_u10_u5_n2034 ), .A3(_u10_u5_n2380 ), .A4(_u10_u5_n2741 ), .ZN(_u10_u5_n2740 ) );
NAND2_X1 _u10_u5_U559  ( .A1(_u10_u5_n1967 ), .A2(_u10_u5_n2740 ), .ZN(_u10_u5_n2733 ) );
NAND3_X1 _u10_u5_U558  ( .A1(_u10_u5_n2739 ), .A2(_u10_u5_n2368 ), .A3(_u10_u5_n2255 ), .ZN(_u10_u5_n2738 ) );
NAND2_X1 _u10_u5_U557  ( .A1(_u10_u5_n2737 ), .A2(_u10_u5_n2738 ), .ZN(_u10_u5_n2734 ) );
NAND2_X1 _u10_u5_U556  ( .A1(_u10_u5_n2736 ), .A2(_u10_u5_n2524 ), .ZN(_u10_u5_n2735 ) );
NAND4_X1 _u10_u5_U555  ( .A1(_u10_u5_n2732 ), .A2(_u10_u5_n2733 ), .A3(_u10_u5_n2734 ), .A4(_u10_u5_n2735 ), .ZN(_u10_u5_n2731 ) );
NOR4_X1 _u10_u5_U554  ( .A1(_u10_u5_n2728 ), .A2(_u10_u5_n2729 ), .A3(_u10_u5_n2730 ), .A4(_u10_u5_n2731 ), .ZN(_u10_u5_n2727 ) );
NAND4_X1 _u10_u5_U553  ( .A1(_u10_u5_n2724 ), .A2(_u10_u5_n2725 ), .A3(_u10_u5_n2726 ), .A4(_u10_u5_n2727 ), .ZN(_u10_u5_n2723 ) );
MUX2_X1 _u10_u5_U552  ( .A(_u10_u5_n2723 ), .B(_u10_SYNOPSYS_UNCONNECTED_19 ), .S(_u10_u5_n1819 ), .Z(_u10_u5_n1809 ) );
NAND2_X1 _u10_u5_U551  ( .A1(_u10_u5_n2002 ), .A2(_u10_u5_n2722 ), .ZN(_u10_u5_n2713 ) );
NAND2_X1 _u10_u5_U550  ( .A1(_u10_u5_n2720 ), .A2(_u10_u5_n2721 ), .ZN(_u10_u5_n2714 ) );
NAND2_X1 _u10_u5_U549  ( .A1(_u10_u5_n2256 ), .A2(_u10_u5_n2719 ), .ZN(_u10_u5_n2715 ) );
NOR2_X1 _u10_u5_U548  ( .A1(_u10_u5_n2106 ), .A2(_u10_u5_n2037 ), .ZN(_u10_u5_n2717 ) );
AND2_X1 _u10_u5_U547  ( .A1(_u10_u5_n1966 ), .A2(_u10_u5_n2054 ), .ZN(_u10_u5_n2718 ) );
NOR2_X1 _u10_u5_U546  ( .A1(_u10_u5_n2717 ), .A2(_u10_u5_n2718 ), .ZN(_u10_u5_n2716 ) );
NAND4_X1 _u10_u5_U545  ( .A1(_u10_u5_n2713 ), .A2(_u10_u5_n2714 ), .A3(_u10_u5_n2715 ), .A4(_u10_u5_n2716 ), .ZN(_u10_u5_n2608 ) );
NAND2_X1 _u10_u5_U544  ( .A1(1'b0), .A2(_u10_u5_n2669 ), .ZN(_u10_u5_n2385 ));
INV_X1 _u10_u5_U543  ( .A(_u10_u5_n2385 ), .ZN(_u10_u5_n1977 ) );
NAND2_X1 _u10_u5_U542  ( .A1(_u10_u5_n1977 ), .A2(_u10_u5_n2668 ), .ZN(_u10_u5_n2712 ) );
NAND2_X1 _u10_u5_U541  ( .A1(_u10_u5_n2712 ), .A2(_u10_u5_n2092 ), .ZN(_u10_u5_n1844 ) );
NAND2_X1 _u10_u5_U540  ( .A1(_u10_u5_n1894 ), .A2(_u10_u5_n1844 ), .ZN(_u10_u5_n2705 ) );
NAND2_X1 _u10_u5_U539  ( .A1(_u10_u5_n1894 ), .A2(_u10_u5_n2305 ), .ZN(_u10_u5_n2711 ) );
NAND2_X1 _u10_u5_U538  ( .A1(_u10_u5_n2711 ), .A2(_u10_u5_n2025 ), .ZN(_u10_u5_n1932 ) );
NAND2_X1 _u10_u5_U537  ( .A1(_u10_u5_n2710 ), .A2(_u10_u5_n1932 ), .ZN(_u10_u5_n2706 ) );
NAND2_X1 _u10_u5_U536  ( .A1(_u10_u5_n2708 ), .A2(_u10_u5_n2709 ), .ZN(_u10_u5_n2707 ) );
NAND3_X1 _u10_u5_U535  ( .A1(_u10_u5_n2705 ), .A2(_u10_u5_n2706 ), .A3(_u10_u5_n2707 ), .ZN(_u10_u5_n2701 ) );
NOR2_X1 _u10_u5_U534  ( .A1(_u10_u5_n1843 ), .A2(_u10_u5_n2545 ), .ZN(_u10_u5_n2702 ) );
NOR2_X1 _u10_u5_U533  ( .A1(_u10_u5_n2346 ), .A2(_u10_u5_n2700 ), .ZN(_u10_u5_n2703 ) );
NOR2_X1 _u10_u5_U532  ( .A1(_u10_u5_n2000 ), .A2(_u10_u5_n1887 ), .ZN(_u10_u5_n2704 ) );
NOR4_X1 _u10_u5_U531  ( .A1(_u10_u5_n2701 ), .A2(_u10_u5_n2702 ), .A3(_u10_u5_n2703 ), .A4(_u10_u5_n2704 ), .ZN(_u10_u5_n2671 ) );
NAND2_X1 _u10_u5_U530  ( .A1(_u10_u5_n2699 ), .A2(_u10_u5_n2700 ), .ZN(_u10_u5_n2698 ) );
NAND2_X1 _u10_u5_U529  ( .A1(_u10_u5_n2063 ), .A2(_u10_u5_n2698 ), .ZN(_u10_u5_n2682 ) );
NAND2_X1 _u10_u5_U528  ( .A1(_u10_u5_n2697 ), .A2(_u10_u5_n2103 ), .ZN(_u10_u5_n2696 ) );
NAND2_X1 _u10_u5_U527  ( .A1(_u10_u5_n2695 ), .A2(_u10_u5_n2696 ), .ZN(_u10_u5_n2694 ) );
NAND2_X1 _u10_u5_U526  ( .A1(_u10_u5_n1937 ), .A2(_u10_u5_n2694 ), .ZN(_u10_u5_n2683 ) );
INV_X1 _u10_u5_U525  ( .A(_u10_u5_n2693 ), .ZN(_u10_u5_n2691 ) );
NAND3_X1 _u10_u5_U524  ( .A1(_u10_u5_n2103 ), .A2(_u10_u5_n2502 ), .A3(1'b0),.ZN(_u10_u5_n2692 ) );
NAND2_X1 _u10_u5_U523  ( .A1(_u10_u5_n2691 ), .A2(_u10_u5_n2692 ), .ZN(_u10_u5_n2690 ) );
NAND2_X1 _u10_u5_U522  ( .A1(_u10_u5_n2236 ), .A2(_u10_u5_n2690 ), .ZN(_u10_u5_n2684 ) );
NAND3_X1 _u10_u5_U521  ( .A1(_u10_u5_n2688 ), .A2(_u10_u5_n1913 ), .A3(_u10_u5_n2689 ), .ZN(_u10_u5_n2335 ) );
NAND3_X1 _u10_u5_U520  ( .A1(_u10_u5_n2536 ), .A2(_u10_u5_n2103 ), .A3(1'b0),.ZN(_u10_u5_n2052 ) );
NOR2_X1 _u10_u5_U519  ( .A1(_u10_u5_n2052 ), .A2(_u10_u5_n2687 ), .ZN(_u10_u5_n1851 ) );
NAND2_X1 _u10_u5_U518  ( .A1(_u10_u5_n1851 ), .A2(_u10_u5_n2078 ), .ZN(_u10_u5_n2582 ) );
NOR2_X1 _u10_u5_U517  ( .A1(_u10_u5_n2686 ), .A2(_u10_u5_n2582 ), .ZN(_u10_u5_n2094 ) );
NAND3_X1 _u10_u5_U516  ( .A1(_u10_u5_n2251 ), .A2(_u10_u5_n2335 ), .A3(_u10_u5_n2094 ), .ZN(_u10_u5_n2685 ) );
NAND4_X1 _u10_u5_U515  ( .A1(_u10_u5_n2682 ), .A2(_u10_u5_n2683 ), .A3(_u10_u5_n2684 ), .A4(_u10_u5_n2685 ), .ZN(_u10_u5_n2673 ) );
INV_X1 _u10_u5_U514  ( .A(_u10_u5_n2291 ), .ZN(_u10_u5_n2057 ) );
AND2_X1 _u10_u5_U513  ( .A1(_u10_u5_n1851 ), .A2(_u10_u5_n2057 ), .ZN(_u10_u5_n2674 ) );
INV_X1 _u10_u5_U512  ( .A(_u10_u5_n1874 ), .ZN(_u10_u5_n2681 ) );
NOR2_X1 _u10_u5_U511  ( .A1(_u10_u5_n2007 ), .A2(_u10_u5_n1911 ), .ZN(_u10_u5_n2486 ) );
NOR2_X1 _u10_u5_U510  ( .A1(_u10_u5_n2681 ), .A2(_u10_u5_n2486 ), .ZN(_u10_u5_n2675 ) );
NOR2_X1 _u10_u5_U509  ( .A1(_u10_u5_n1977 ), .A2(_u10_u5_n2680 ), .ZN(_u10_u5_n2679 ) );
NOR2_X1 _u10_u5_U508  ( .A1(_u10_u5_n2679 ), .A2(_u10_u5_n2030 ), .ZN(_u10_u5_n2678 ) );
NOR2_X1 _u10_u5_U507  ( .A1(_u10_u5_n2678 ), .A2(_u10_u5_n2094 ), .ZN(_u10_u5_n2677 ) );
NOR2_X1 _u10_u5_U506  ( .A1(_u10_u5_n2677 ), .A2(_u10_u5_n2025 ), .ZN(_u10_u5_n2676 ) );
NOR4_X1 _u10_u5_U505  ( .A1(_u10_u5_n2673 ), .A2(_u10_u5_n2674 ), .A3(_u10_u5_n2675 ), .A4(_u10_u5_n2676 ), .ZN(_u10_u5_n2672 ) );
AND2_X1 _u10_u5_U504  ( .A1(_u10_u5_n2671 ), .A2(_u10_u5_n2672 ), .ZN(_u10_u5_n1990 ) );
INV_X1 _u10_u5_U503  ( .A(_u10_u5_n2670 ), .ZN(_u10_u5_n2660 ) );
NAND4_X1 _u10_u5_U502  ( .A1(_u10_u5_n2251 ), .A2(_u10_u5_n2669 ), .A3(_u10_u5_n2162 ), .A4(_u10_u5_n2169 ), .ZN(_u10_u5_n2664 ) );
AND3_X1 _u10_u5_U501  ( .A1(_u10_u5_n1977 ), .A2(_u10_u5_n2668 ), .A3(_u10_u5_n2089 ), .ZN(_u10_u5_n2555 ) );
NAND2_X1 _u10_u5_U500  ( .A1(_u10_u5_n2555 ), .A2(_u10_u5_n2667 ), .ZN(_u10_u5_n2666 ) );
NAND3_X1 _u10_u5_U499  ( .A1(_u10_u5_n2664 ), .A2(_u10_u5_n2665 ), .A3(_u10_u5_n2666 ), .ZN(_u10_u5_n1988 ) );
INV_X1 _u10_u5_U498  ( .A(_u10_u5_n1988 ), .ZN(_u10_u5_n2661 ) );
NAND2_X1 _u10_u5_U497  ( .A1(1'b0), .A2(_u10_u5_n2043 ), .ZN(_u10_u5_n2662 ));
NAND2_X1 _u10_u5_U496  ( .A1(_u10_u5_n2169 ), .A2(1'b0), .ZN(_u10_u5_n2663 ));
NAND4_X1 _u10_u5_U495  ( .A1(_u10_u5_n2660 ), .A2(_u10_u5_n2661 ), .A3(_u10_u5_n2662 ), .A4(_u10_u5_n2663 ), .ZN(_u10_u5_n2650 ) );
NAND2_X1 _u10_u5_U494  ( .A1(_u10_u5_n2659 ), .A2(1'b0), .ZN(_u10_u5_n2193 ));
INV_X1 _u10_u5_U493  ( .A(_u10_u5_n2193 ), .ZN(_u10_u5_n2143 ) );
NAND2_X1 _u10_u5_U492  ( .A1(_u10_u5_n2143 ), .A2(_u10_u5_n2036 ), .ZN(_u10_u5_n2286 ) );
INV_X1 _u10_u5_U491  ( .A(_u10_u5_n2286 ), .ZN(_u10_u5_n2577 ) );
NAND2_X1 _u10_u5_U490  ( .A1(_u10_u5_n2577 ), .A2(_u10_u5_n2278 ), .ZN(_u10_u5_n2474 ) );
INV_X1 _u10_u5_U489  ( .A(_u10_u5_n2474 ), .ZN(_u10_u5_n2306 ) );
NAND2_X1 _u10_u5_U488  ( .A1(_u10_u5_n2306 ), .A2(_u10_u5_n2251 ), .ZN(_u10_u5_n2654 ) );
NAND2_X1 _u10_u5_U487  ( .A1(_u10_u5_n2649 ), .A2(_u10_u5_n2658 ), .ZN(_u10_u5_n2655 ) );
NAND2_X1 _u10_u5_U486  ( .A1(_u10_u5_n2657 ), .A2(_u10_u5_n2445 ), .ZN(_u10_u5_n2656 ) );
NAND3_X1 _u10_u5_U485  ( .A1(_u10_u5_n2654 ), .A2(_u10_u5_n2655 ), .A3(_u10_u5_n2656 ), .ZN(_u10_u5_n2651 ) );
NOR2_X1 _u10_u5_U484  ( .A1(_u10_u5_n2366 ), .A2(_u10_u5_n2376 ), .ZN(_u10_u5_n2652 ) );
AND2_X1 _u10_u5_U483  ( .A1(_u10_u5_n1966 ), .A2(_u10_u5_n2528 ), .ZN(_u10_u5_n2653 ) );
NOR4_X1 _u10_u5_U482  ( .A1(_u10_u5_n2650 ), .A2(_u10_u5_n2651 ), .A3(_u10_u5_n2652 ), .A4(_u10_u5_n2653 ), .ZN(_u10_u5_n2613 ) );
NAND2_X1 _u10_u5_U481  ( .A1(_u10_u5_n1891 ), .A2(1'b0), .ZN(_u10_u5_n2636 ));
NAND2_X1 _u10_u5_U480  ( .A1(_u10_u5_n1868 ), .A2(_u10_u5_n2113 ), .ZN(_u10_u5_n2101 ) );
NOR4_X1 _u10_u5_U479  ( .A1(_u10_u5_n2649 ), .A2(_u10_u5_n2216 ), .A3(_u10_u5_n2101 ), .A4(_u10_u5_n2634 ), .ZN(_u10_u5_n2648 ) );
NOR2_X1 _u10_u5_U478  ( .A1(_u10_u5_n2648 ), .A2(_u10_u5_n2254 ), .ZN(_u10_u5_n2638 ) );
NOR2_X1 _u10_u5_U477  ( .A1(_u10_u5_n2106 ), .A2(_u10_u5_n2643 ), .ZN(_u10_u5_n2645 ) );
NAND2_X1 _u10_u5_U476  ( .A1(1'b0), .A2(_u10_u5_n2049 ), .ZN(_u10_u5_n2647 ));
NAND2_X1 _u10_u5_U475  ( .A1(_u10_u5_n2646 ), .A2(_u10_u5_n2647 ), .ZN(_u10_u5_n2348 ) );
NOR2_X1 _u10_u5_U474  ( .A1(_u10_u5_n2645 ), .A2(_u10_u5_n2348 ), .ZN(_u10_u5_n2644 ) );
NOR2_X1 _u10_u5_U473  ( .A1(_u10_u5_n2644 ), .A2(_u10_u5_n2495 ), .ZN(_u10_u5_n2639 ) );
NOR2_X1 _u10_u5_U472  ( .A1(_u10_u5_n2643 ), .A2(_u10_u5_n2203 ), .ZN(_u10_u5_n2642 ) );
NOR3_X1 _u10_u5_U471  ( .A1(_u10_u5_n2101 ), .A2(1'b0), .A3(_u10_u5_n2642 ),.ZN(_u10_u5_n2641 ) );
NOR2_X1 _u10_u5_U470  ( .A1(_u10_u5_n2641 ), .A2(_u10_u5_n2253 ), .ZN(_u10_u5_n2640 ) );
NOR3_X1 _u10_u5_U469  ( .A1(_u10_u5_n2638 ), .A2(_u10_u5_n2639 ), .A3(_u10_u5_n2640 ), .ZN(_u10_u5_n2637 ) );
NAND3_X1 _u10_u5_U468  ( .A1(_u10_u5_n2635 ), .A2(_u10_u5_n2636 ), .A3(_u10_u5_n2637 ), .ZN(_u10_u5_n2615 ) );
NOR3_X1 _u10_u5_U467  ( .A1(_u10_u5_n2174 ), .A2(_u10_u5_n2175 ), .A3(_u10_u5_n2179 ), .ZN(_u10_u5_n2631 ) );
NAND3_X1 _u10_u5_U466  ( .A1(_u10_u5_n2223 ), .A2(_u10_u5_n2236 ), .A3(_u10_u5_n2631 ), .ZN(_u10_u5_n2622 ) );
OR2_X1 _u10_u5_U465  ( .A1(_u10_u5_n1960 ), .A2(_u10_u5_n1959 ), .ZN(_u10_u5_n2625 ) );
NOR3_X1 _u10_u5_U464  ( .A1(_u10_u5_n2101 ), .A2(_u10_u5_n2633 ), .A3(_u10_u5_n2634 ), .ZN(_u10_u5_n2523 ) );
OR2_X1 _u10_u5_U463  ( .A1(_u10_u5_n2632 ), .A2(_u10_u5_n2523 ), .ZN(_u10_u5_n2627 ) );
INV_X1 _u10_u5_U462  ( .A(_u10_u5_n2631 ), .ZN(_u10_u5_n2628 ) );
NAND2_X1 _u10_u5_U461  ( .A1(_u10_u5_n2630 ), .A2(_u10_u5_n1922 ), .ZN(_u10_u5_n2629 ) );
NAND3_X1 _u10_u5_U460  ( .A1(_u10_u5_n2627 ), .A2(_u10_u5_n2628 ), .A3(_u10_u5_n2629 ), .ZN(_u10_u5_n2626 ) );
NAND2_X1 _u10_u5_U459  ( .A1(_u10_u5_n2625 ), .A2(_u10_u5_n2626 ), .ZN(_u10_u5_n2624 ) );
NAND3_X1 _u10_u5_U458  ( .A1(_u10_u5_n2622 ), .A2(_u10_u5_n2623 ), .A3(_u10_u5_n2624 ), .ZN(_u10_u5_n2616 ) );
AND2_X1 _u10_u5_U457  ( .A1(_u10_u5_n2621 ), .A2(_u10_u5_n2358 ), .ZN(_u10_u5_n2620 ) );
NOR2_X1 _u10_u5_U456  ( .A1(_u10_u5_n2523 ), .A2(_u10_u5_n2620 ), .ZN(_u10_u5_n2617 ) );
INV_X1 _u10_u5_U455  ( .A(_u10_u5_n2101 ), .ZN(_u10_u5_n2221 ) );
NOR2_X1 _u10_u5_U454  ( .A1(_u10_u5_n1911 ), .A2(_u10_u5_n2488 ), .ZN(_u10_u5_n2619 ) );
NOR2_X1 _u10_u5_U453  ( .A1(_u10_u5_n2221 ), .A2(_u10_u5_n2619 ), .ZN(_u10_u5_n2618 ) );
NOR4_X1 _u10_u5_U452  ( .A1(_u10_u5_n2615 ), .A2(_u10_u5_n2616 ), .A3(_u10_u5_n2617 ), .A4(_u10_u5_n2618 ), .ZN(_u10_u5_n2614 ) );
AND2_X1 _u10_u5_U451  ( .A1(_u10_u5_n2613 ), .A2(_u10_u5_n2614 ), .ZN(_u10_u5_n2314 ) );
NAND3_X1 _u10_u5_U450  ( .A1(_u10_u5_n2612 ), .A2(_u10_u5_n1990 ), .A3(_u10_u5_n2314 ), .ZN(_u10_u5_n2609 ) );
NOR4_X1 _u10_u5_U449  ( .A1(_u10_u5_n2608 ), .A2(_u10_u5_n2609 ), .A3(_u10_u5_n2610 ), .A4(_u10_u5_n2611 ), .ZN(_u10_u5_n2388 ) );
NAND2_X1 _u10_u5_U448  ( .A1(_u10_u5_n2346 ), .A2(_u10_u5_n2607 ), .ZN(_u10_u5_n2191 ) );
NAND2_X1 _u10_u5_U447  ( .A1(_u10_u5_n2143 ), .A2(_u10_u5_n2191 ), .ZN(_u10_u5_n2556 ) );
INV_X1 _u10_u5_U446  ( .A(_u10_u5_n2348 ), .ZN(_u10_u5_n2603 ) );
NAND3_X1 _u10_u5_U445  ( .A1(_u10_u5_n2535 ), .A2(_u10_u5_n2485 ), .A3(_u10_u5_n2456 ), .ZN(_u10_u5_n2606 ) );
NAND2_X1 _u10_u5_U444  ( .A1(_u10_u5_n2049 ), .A2(_u10_u5_n2606 ), .ZN(_u10_u5_n2604 ) );
NAND3_X1 _u10_u5_U443  ( .A1(_u10_u5_n2603 ), .A2(_u10_u5_n2604 ), .A3(_u10_u5_n2605 ), .ZN(_u10_u5_n2602 ) );
NAND2_X1 _u10_u5_U442  ( .A1(_u10_u5_n2043 ), .A2(_u10_u5_n2602 ), .ZN(_u10_u5_n2557 ) );
INV_X1 _u10_u5_U441  ( .A(_u10_u5_n2601 ), .ZN(_u10_u5_n2590 ) );
NAND2_X1 _u10_u5_U440  ( .A1(_u10_u5_n2599 ), .A2(_u10_u5_n2600 ), .ZN(_u10_u5_n2597 ) );
NAND2_X1 _u10_u5_U439  ( .A1(_u10_u5_n2082 ), .A2(_u10_u5_n2101 ), .ZN(_u10_u5_n2598 ) );
AND2_X1 _u10_u5_U438  ( .A1(_u10_u5_n2597 ), .A2(_u10_u5_n2598 ), .ZN(_u10_u5_n2281 ) );
NAND3_X1 _u10_u5_U437  ( .A1(_u10_u5_n1969 ), .A2(_u10_u5_n2582 ), .A3(_u10_u5_n2281 ), .ZN(_u10_u5_n2073 ) );
INV_X1 _u10_u5_U436  ( .A(_u10_u5_n2073 ), .ZN(_u10_u5_n2591 ) );
NOR2_X1 _u10_u5_U435  ( .A1(_u10_u5_n1816 ), .A2(_u10_u5_n2077 ), .ZN(_u10_u5_n2595 ) );
NOR2_X1 _u10_u5_U434  ( .A1(_u10_u5_n2595 ), .A2(_u10_u5_n2596 ), .ZN(_u10_u5_n2592 ) );
NAND3_X1 _u10_u5_U433  ( .A1(_u10_u5_n2107 ), .A2(_u10_u5_n2536 ), .A3(1'b0),.ZN(_u10_u5_n2438 ) );
INV_X1 _u10_u5_U432  ( .A(_u10_u5_n2438 ), .ZN(_u10_u5_n2427 ) );
NOR4_X1 _u10_u5_U431  ( .A1(1'b0), .A2(_u10_u5_n2594 ), .A3(_u10_u5_n2577 ),.A4(_u10_u5_n2427 ), .ZN(_u10_u5_n2593 ) );
NAND4_X1 _u10_u5_U430  ( .A1(_u10_u5_n2590 ), .A2(_u10_u5_n2591 ), .A3(_u10_u5_n2592 ), .A4(_u10_u5_n2593 ), .ZN(_u10_u5_n2589 ) );
NAND2_X1 _u10_u5_U429  ( .A1(_u10_u5_n2279 ), .A2(_u10_u5_n2589 ), .ZN(_u10_u5_n2558 ) );
NAND3_X1 _u10_u5_U428  ( .A1(_u10_u5_n2587 ), .A2(_u10_u5_n2115 ), .A3(_u10_u5_n2588 ), .ZN(_u10_u5_n2585 ) );
NOR4_X1 _u10_u5_U427  ( .A1(_u10_u5_n2585 ), .A2(_u10_u5_n2586 ), .A3(1'b0),.A4(_u10_u5_n2114 ), .ZN(_u10_u5_n2583 ) );
NOR2_X1 _u10_u5_U426  ( .A1(_u10_u5_n2583 ), .A2(_u10_u5_n2584 ), .ZN(_u10_u5_n2560 ) );
OR2_X1 _u10_u5_U425  ( .A1(_u10_u5_n2582 ), .A2(1'b0), .ZN(_u10_u5_n2581 ));
NAND2_X1 _u10_u5_U424  ( .A1(_u10_u5_n2580 ), .A2(_u10_u5_n2581 ), .ZN(_u10_u5_n1974 ) );
INV_X1 _u10_u5_U423  ( .A(_u10_u5_n1974 ), .ZN(_u10_u5_n1901 ) );
AND4_X1 _u10_u5_U422  ( .A1(_u10_u5_n1901 ), .A2(_u10_u5_n2385 ), .A3(_u10_u5_n2578 ), .A4(_u10_u5_n2579 ), .ZN(_u10_u5_n2424 ) );
NOR2_X1 _u10_u5_U421  ( .A1(1'b0), .A2(_u10_u5_n2424 ), .ZN(_u10_u5_n2574 ));
NOR3_X1 _u10_u5_U420  ( .A1(_u10_u5_n2427 ), .A2(1'b0), .A3(_u10_u5_n2577 ),.ZN(_u10_u5_n2576 ) );
NOR2_X1 _u10_u5_U419  ( .A1(_u10_u5_n2576 ), .A2(_u10_u5_n1976 ), .ZN(_u10_u5_n2575 ) );
NOR3_X1 _u10_u5_U418  ( .A1(_u10_u5_n2574 ), .A2(_u10_u5_n1979 ), .A3(_u10_u5_n2575 ), .ZN(_u10_u5_n2572 ) );
NOR2_X1 _u10_u5_U417  ( .A1(_u10_u5_n2572 ), .A2(_u10_u5_n2573 ), .ZN(_u10_u5_n2561 ) );
INV_X1 _u10_u5_U416  ( .A(_u10_u5_n2061 ), .ZN(_u10_u5_n2453 ) );
NOR2_X1 _u10_u5_U415  ( .A1(_u10_u5_n2453 ), .A2(_u10_u5_n1851 ), .ZN(_u10_u5_n2018 ) );
NAND2_X1 _u10_u5_U414  ( .A1(1'b0), .A2(_u10_u5_n2571 ), .ZN(_u10_u5_n2570 ));
NAND2_X1 _u10_u5_U413  ( .A1(_u10_u5_n2018 ), .A2(_u10_u5_n2570 ), .ZN(_u10_u5_n1837 ) );
INV_X1 _u10_u5_U412  ( .A(_u10_u5_n1837 ), .ZN(_u10_u5_n2568 ) );
NAND2_X1 _u10_u5_U411  ( .A1(1'b0), .A2(_u10_u5_n2536 ), .ZN(_u10_u5_n2569 ));
NAND2_X1 _u10_u5_U410  ( .A1(_u10_u5_n2568 ), .A2(_u10_u5_n2569 ), .ZN(_u10_u5_n2564 ) );
NOR2_X1 _u10_u5_U409  ( .A1(_u10_u5_n1841 ), .A2(_u10_u5_n1868 ), .ZN(_u10_u5_n2565 ) );
INV_X1 _u10_u5_U408  ( .A(_u10_u5_n2567 ), .ZN(_u10_u5_n2566 ) );
NOR4_X1 _u10_u5_U407  ( .A1(_u10_u5_n2564 ), .A2(_u10_u5_n2565 ), .A3(_u10_u5_n2143 ), .A4(_u10_u5_n2566 ), .ZN(_u10_u5_n2563 ) );
NOR2_X1 _u10_u5_U406  ( .A1(_u10_u5_n2563 ), .A2(_u10_u5_n2014 ), .ZN(_u10_u5_n2562 ) );
NOR3_X1 _u10_u5_U405  ( .A1(_u10_u5_n2560 ), .A2(_u10_u5_n2561 ), .A3(_u10_u5_n2562 ), .ZN(_u10_u5_n2559 ) );
NAND4_X1 _u10_u5_U404  ( .A1(_u10_u5_n2556 ), .A2(_u10_u5_n2557 ), .A3(_u10_u5_n2558 ), .A4(_u10_u5_n2559 ), .ZN(_u10_u5_n2511 ) );
INV_X1 _u10_u5_U403  ( .A(_u10_u5_n2085 ), .ZN(_u10_u5_n2293 ) );
NOR2_X1 _u10_u5_U402  ( .A1(_u10_u5_n2554 ), .A2(_u10_u5_n2555 ), .ZN(_u10_u5_n2444 ) );
NAND2_X1 _u10_u5_U401  ( .A1(_u10_u5_n2553 ), .A2(_u10_u5_n2549 ), .ZN(_u10_u5_n2552 ) );
AND2_X1 _u10_u5_U400  ( .A1(_u10_u5_n2444 ), .A2(_u10_u5_n2552 ), .ZN(_u10_u5_n2295 ) );
NAND2_X1 _u10_u5_U399  ( .A1(_u10_u5_n2551 ), .A2(_u10_u5_n2549 ), .ZN(_u10_u5_n2538 ) );
AND2_X1 _u10_u5_U398  ( .A1(_u10_u5_n2427 ), .A2(_u10_u5_n2108 ), .ZN(_u10_u5_n2460 ) );
NOR4_X1 _u10_u5_U397  ( .A1(_u10_u5_n2460 ), .A2(_u10_u5_n2306 ), .A3(_u10_u5_n2094 ), .A4(_u10_u5_n2550 ), .ZN(_u10_u5_n2409 ) );
INV_X1 _u10_u5_U396  ( .A(_u10_u5_n2409 ), .ZN(_u10_u5_n2407 ) );
NAND2_X1 _u10_u5_U395  ( .A1(_u10_u5_n2549 ), .A2(_u10_u5_n2407 ), .ZN(_u10_u5_n2546 ) );
NAND3_X1 _u10_u5_U394  ( .A1(_u10_u5_n2546 ), .A2(_u10_u5_n2547 ), .A3(_u10_u5_n2548 ), .ZN(_u10_u5_n2501 ) );
INV_X1 _u10_u5_U393  ( .A(_u10_u5_n2501 ), .ZN(_u10_u5_n2539 ) );
NOR2_X1 _u10_u5_U392  ( .A1(1'b0), .A2(_u10_u5_n2545 ), .ZN(_u10_u5_n2541 ));
AND2_X1 _u10_u5_U391  ( .A1(_u10_u5_n2544 ), .A2(_u10_u5_n2089 ), .ZN(_u10_u5_n2543 ) );
NOR3_X1 _u10_u5_U390  ( .A1(_u10_u5_n2541 ), .A2(_u10_u5_n2542 ), .A3(_u10_u5_n2543 ), .ZN(_u10_u5_n2540 ) );
NAND4_X1 _u10_u5_U389  ( .A1(_u10_u5_n2295 ), .A2(_u10_u5_n2538 ), .A3(_u10_u5_n2539 ), .A4(_u10_u5_n2540 ), .ZN(_u10_u5_n2537 ) );
NAND2_X1 _u10_u5_U388  ( .A1(_u10_u5_n2293 ), .A2(_u10_u5_n2537 ), .ZN(_u10_u5_n2515 ) );
NAND2_X1 _u10_u5_U387  ( .A1(_u10_u5_n2536 ), .A2(_u10_u5_n2508 ), .ZN(_u10_u5_n2526 ) );
NAND2_X1 _u10_u5_U386  ( .A1(_u10_u5_n2535 ), .A2(_u10_u5_n1940 ), .ZN(_u10_u5_n2532 ) );
NOR4_X1 _u10_u5_U385  ( .A1(_u10_u5_n2532 ), .A2(_u10_u5_n2533 ), .A3(1'b0),.A4(_u10_u5_n2534 ), .ZN(_u10_u5_n2530 ) );
NOR2_X1 _u10_u5_U384  ( .A1(_u10_u5_n2530 ), .A2(_u10_u5_n2531 ), .ZN(_u10_u5_n2529 ) );
NOR4_X1 _u10_u5_U383  ( .A1(_u10_u5_n2528 ), .A2(_u10_u5_n2143 ), .A3(_u10_u5_n2189 ), .A4(_u10_u5_n2529 ), .ZN(_u10_u5_n2527 ) );
NAND4_X1 _u10_u5_U382  ( .A1(_u10_u5_n2019 ), .A2(_u10_u5_n2526 ), .A3(_u10_u5_n2018 ), .A4(_u10_u5_n2527 ), .ZN(_u10_u5_n2525 ) );
NAND2_X1 _u10_u5_U381  ( .A1(_u10_u5_n2183 ), .A2(_u10_u5_n2525 ), .ZN(_u10_u5_n2516 ) );
INV_X1 _u10_u5_U380  ( .A(_u10_u5_n2524 ), .ZN(_u10_u5_n2396 ) );
NAND2_X1 _u10_u5_U379  ( .A1(_u10_u5_n2396 ), .A2(_u10_u5_n2523 ), .ZN(_u10_u5_n2522 ) );
NAND2_X1 _u10_u5_U378  ( .A1(_u10_u5_n1866 ), .A2(_u10_u5_n2522 ), .ZN(_u10_u5_n2519 ) );
AND2_X1 _u10_u5_U377  ( .A1(_u10_u5_n2493 ), .A2(_u10_u5_n1961 ), .ZN(_u10_u5_n2429 ) );
NAND2_X1 _u10_u5_U376  ( .A1(_u10_u5_n2429 ), .A2(_u10_u5_n2175 ), .ZN(_u10_u5_n2510 ) );
NAND2_X1 _u10_u5_U375  ( .A1(_u10_u5_n2510 ), .A2(_u10_u5_n1864 ), .ZN(_u10_u5_n2521 ) );
NAND3_X1 _u10_u5_U374  ( .A1(_u10_u5_n2519 ), .A2(_u10_u5_n2520 ), .A3(_u10_u5_n2521 ), .ZN(_u10_u5_n2518 ) );
NAND2_X1 _u10_u5_U373  ( .A1(_u10_u5_n1861 ), .A2(_u10_u5_n2518 ), .ZN(_u10_u5_n2517 ) );
NAND3_X1 _u10_u5_U372  ( .A1(_u10_u5_n2515 ), .A2(_u10_u5_n2516 ), .A3(_u10_u5_n2517 ), .ZN(_u10_u5_n2512 ) );
NOR2_X1 _u10_u5_U371  ( .A1(_u10_u5_n1913 ), .A2(_u10_u5_n1940 ), .ZN(_u10_u5_n2513 ) );
NOR2_X1 _u10_u5_U370  ( .A1(_u10_u5_n2113 ), .A2(_u10_u5_n2350 ), .ZN(_u10_u5_n2514 ) );
NOR4_X1 _u10_u5_U369  ( .A1(_u10_u5_n2511 ), .A2(_u10_u5_n2512 ), .A3(_u10_u5_n2513 ), .A4(_u10_u5_n2514 ), .ZN(_u10_u5_n2389 ) );
NAND2_X1 _u10_u5_U368  ( .A1(_u10_u5_n2509 ), .A2(_u10_u5_n2510 ), .ZN(_u10_u5_n2477 ) );
NAND2_X1 _u10_u5_U367  ( .A1(_u10_u5_n2507 ), .A2(_u10_u5_n2508 ), .ZN(_u10_u5_n2504 ) );
NAND2_X1 _u10_u5_U366  ( .A1(1'b0), .A2(_u10_u5_n2506 ), .ZN(_u10_u5_n2505 ));
NAND2_X1 _u10_u5_U365  ( .A1(_u10_u5_n2504 ), .A2(_u10_u5_n2505 ), .ZN(_u10_u5_n2503 ) );
NAND2_X1 _u10_u5_U364  ( .A1(_u10_u5_n2502 ), .A2(_u10_u5_n2503 ), .ZN(_u10_u5_n2478 ) );
NAND2_X1 _u10_u5_U363  ( .A1(_u10_u5_n2501 ), .A2(_u10_u5_n2446 ), .ZN(_u10_u5_n2497 ) );
INV_X1 _u10_u5_U362  ( .A(_u10_u5_n2500 ), .ZN(_u10_u5_n2499 ) );
NAND3_X1 _u10_u5_U361  ( .A1(_u10_u5_n2497 ), .A2(_u10_u5_n2498 ), .A3(_u10_u5_n2499 ), .ZN(_u10_u5_n2496 ) );
NAND2_X1 _u10_u5_U360  ( .A1(_u10_u5_n2445 ), .A2(_u10_u5_n2496 ), .ZN(_u10_u5_n2479 ) );
NOR2_X1 _u10_u5_U359  ( .A1(_u10_u5_n2429 ), .A2(_u10_u5_n2495 ), .ZN(_u10_u5_n2491 ) );
INV_X1 _u10_u5_U358  ( .A(_u10_u5_n2191 ), .ZN(_u10_u5_n2494 ) );
NOR2_X1 _u10_u5_U357  ( .A1(_u10_u5_n2493 ), .A2(_u10_u5_n2494 ), .ZN(_u10_u5_n2492 ) );
NOR2_X1 _u10_u5_U356  ( .A1(_u10_u5_n2491 ), .A2(_u10_u5_n2492 ), .ZN(_u10_u5_n2489 ) );
NOR2_X1 _u10_u5_U355  ( .A1(_u10_u5_n2489 ), .A2(_u10_u5_n2490 ), .ZN(_u10_u5_n2481 ) );
NAND2_X1 _u10_u5_U354  ( .A1(_u10_u5_n2253 ), .A2(_u10_u5_n1859 ), .ZN(_u10_u5_n2398 ) );
NOR2_X1 _u10_u5_U353  ( .A1(_u10_u5_n2488 ), .A2(_u10_u5_n2398 ), .ZN(_u10_u5_n2487 ) );
NOR2_X1 _u10_u5_U352  ( .A1(_u10_u5_n2220 ), .A2(_u10_u5_n2487 ), .ZN(_u10_u5_n2482 ) );
AND2_X1 _u10_u5_U351  ( .A1(_u10_u5_n2350 ), .A2(_u10_u5_n2486 ), .ZN(_u10_u5_n2484 ) );
NOR2_X1 _u10_u5_U350  ( .A1(_u10_u5_n2484 ), .A2(_u10_u5_n2485 ), .ZN(_u10_u5_n2483 ) );
NOR3_X1 _u10_u5_U349  ( .A1(_u10_u5_n2481 ), .A2(_u10_u5_n2482 ), .A3(_u10_u5_n2483 ), .ZN(_u10_u5_n2480 ) );
NAND4_X1 _u10_u5_U348  ( .A1(_u10_u5_n2477 ), .A2(_u10_u5_n2478 ), .A3(_u10_u5_n2479 ), .A4(_u10_u5_n2480 ), .ZN(_u10_u5_n2447 ) );
NAND2_X1 _u10_u5_U347  ( .A1(_u10_u5_n2476 ), .A2(_u10_u5_n1936 ), .ZN(_u10_u5_n2472 ) );
NAND2_X1 _u10_u5_U346  ( .A1(_u10_u5_n2427 ), .A2(_u10_u5_n2278 ), .ZN(_u10_u5_n2473 ) );
NAND4_X1 _u10_u5_U345  ( .A1(_u10_u5_n2472 ), .A2(_u10_u5_n2473 ), .A3(_u10_u5_n2474 ), .A4(_u10_u5_n2475 ), .ZN(_u10_u5_n2471 ) );
NAND2_X1 _u10_u5_U344  ( .A1(_u10_u5_n2470 ), .A2(_u10_u5_n2471 ), .ZN(_u10_u5_n2457 ) );
NAND2_X1 _u10_u5_U343  ( .A1(_u10_u5_n2409 ), .A2(_u10_u5_n2469 ), .ZN(_u10_u5_n2468 ) );
NAND2_X1 _u10_u5_U342  ( .A1(_u10_u5_n2467 ), .A2(_u10_u5_n2468 ), .ZN(_u10_u5_n2463 ) );
NAND2_X1 _u10_u5_U341  ( .A1(_u10_u5_n1844 ), .A2(_u10_u5_n2466 ), .ZN(_u10_u5_n2465 ) );
NAND3_X1 _u10_u5_U340  ( .A1(_u10_u5_n2463 ), .A2(_u10_u5_n2464 ), .A3(_u10_u5_n2465 ), .ZN(_u10_u5_n2462 ) );
NAND2_X1 _u10_u5_U339  ( .A1(_u10_u5_n2461 ), .A2(_u10_u5_n2462 ), .ZN(_u10_u5_n2458 ) );
NAND2_X1 _u10_u5_U338  ( .A1(_u10_u5_n2460 ), .A2(_u10_u5_n2251 ), .ZN(_u10_u5_n2459 ) );
NAND3_X1 _u10_u5_U337  ( .A1(_u10_u5_n2457 ), .A2(_u10_u5_n2458 ), .A3(_u10_u5_n2459 ), .ZN(_u10_u5_n2448 ) );
NOR2_X1 _u10_u5_U336  ( .A1(_u10_u5_n2455 ), .A2(_u10_u5_n2456 ), .ZN(_u10_u5_n2449 ) );
NAND2_X1 _u10_u5_U335  ( .A1(_u10_u5_n2454 ), .A2(_u10_u5_n2438 ), .ZN(_u10_u5_n2452 ) );
NOR4_X1 _u10_u5_U334  ( .A1(_u10_u5_n2452 ), .A2(_u10_u5_n2453 ), .A3(_u10_u5_n2443 ), .A4(_u10_u5_n2143 ), .ZN(_u10_u5_n2451 ) );
NOR2_X1 _u10_u5_U333  ( .A1(_u10_u5_n2451 ), .A2(_u10_u5_n2356 ), .ZN(_u10_u5_n2450 ) );
NOR4_X1 _u10_u5_U332  ( .A1(_u10_u5_n2447 ), .A2(_u10_u5_n2448 ), .A3(_u10_u5_n2449 ), .A4(_u10_u5_n2450 ), .ZN(_u10_u5_n2390 ) );
NAND2_X1 _u10_u5_U331  ( .A1(_u10_u5_n2445 ), .A2(_u10_u5_n2446 ), .ZN(_u10_u5_n2155 ) );
INV_X1 _u10_u5_U330  ( .A(_u10_u5_n2155 ), .ZN(_u10_u5_n1892 ) );
INV_X1 _u10_u5_U329  ( .A(_u10_u5_n2444 ), .ZN(_u10_u5_n2088 ) );
NAND2_X1 _u10_u5_U328  ( .A1(_u10_u5_n1892 ), .A2(_u10_u5_n2088 ), .ZN(_u10_u5_n2337 ) );
NOR3_X1 _u10_u5_U327  ( .A1(_u10_u5_n2441 ), .A2(_u10_u5_n2442 ), .A3(_u10_u5_n2443 ), .ZN(_u10_u5_n2440 ) );
NAND4_X1 _u10_u5_U326  ( .A1(_u10_u5_n2193 ), .A2(_u10_u5_n2355 ), .A3(_u10_u5_n2439 ), .A4(_u10_u5_n2440 ), .ZN(_u10_u5_n2434 ) );
NAND3_X1 _u10_u5_U325  ( .A1(_u10_u5_n2437 ), .A2(_u10_u5_n2438 ), .A3(_u10_u5_n2059 ), .ZN(_u10_u5_n2435 ) );
NOR4_X1 _u10_u5_U324  ( .A1(_u10_u5_n2434 ), .A2(_u10_u5_n2435 ), .A3(_u10_u5_n1837 ), .A4(_u10_u5_n2436 ), .ZN(_u10_u5_n2433 ) );
NOR2_X1 _u10_u5_U323  ( .A1(_u10_u5_n2433 ), .A2(_u10_u5_n1836 ), .ZN(_u10_u5_n2415 ) );
INV_X1 _u10_u5_U322  ( .A(_u10_u5_n2432 ), .ZN(_u10_u5_n2178 ) );
NOR2_X1 _u10_u5_U321  ( .A1(_u10_u5_n1960 ), .A2(_u10_u5_n2431 ), .ZN(_u10_u5_n2430 ) );
NOR4_X1 _u10_u5_U320  ( .A1(_u10_u5_n2178 ), .A2(_u10_u5_n2429 ), .A3(_u10_u5_n2430 ), .A4(_u10_u5_n2179 ), .ZN(_u10_u5_n2416 ) );
NOR2_X1 _u10_u5_U319  ( .A1(_u10_u5_n2427 ), .A2(_u10_u5_n2428 ), .ZN(_u10_u5_n2426 ) );
NAND4_X1 _u10_u5_U318  ( .A1(_u10_u5_n2286 ), .A2(_u10_u5_n1969 ), .A3(_u10_u5_n2282 ), .A4(_u10_u5_n2426 ), .ZN(_u10_u5_n2425 ) );
NAND2_X1 _u10_u5_U317  ( .A1(_u10_u5_n2031 ), .A2(_u10_u5_n2425 ), .ZN(_u10_u5_n2422 ) );
NAND3_X1 _u10_u5_U316  ( .A1(_u10_u5_n2422 ), .A2(_u10_u5_n2423 ), .A3(_u10_u5_n2424 ), .ZN(_u10_u5_n2419 ) );
NOR4_X1 _u10_u5_U315  ( .A1(_u10_u5_n2419 ), .A2(_u10_u5_n1978 ), .A3(_u10_u5_n2420 ), .A4(_u10_u5_n2421 ), .ZN(_u10_u5_n2418 ) );
NOR2_X1 _u10_u5_U314  ( .A1(_u10_u5_n2418 ), .A2(_u10_u5_n2359 ), .ZN(_u10_u5_n2417 ) );
NOR3_X1 _u10_u5_U313  ( .A1(_u10_u5_n2415 ), .A2(_u10_u5_n2416 ), .A3(_u10_u5_n2417 ), .ZN(_u10_u5_n2414 ) );
NAND4_X1 _u10_u5_U312  ( .A1(_u10_u5_n2337 ), .A2(_u10_u5_n2412 ), .A3(_u10_u5_n2413 ), .A4(_u10_u5_n2414 ), .ZN(_u10_u5_n2392 ) );
NAND2_X1 _u10_u5_U311  ( .A1(_u10_u5_n2411 ), .A2(_u10_u5_n1936 ), .ZN(_u10_u5_n2410 ) );
NAND2_X1 _u10_u5_U310  ( .A1(_u10_u5_n2409 ), .A2(_u10_u5_n2410 ), .ZN(_u10_u5_n2408 ) );
NAND3_X1 _u10_u5_U309  ( .A1(_u10_u5_n2408 ), .A2(_u10_u5_n2305 ), .A3(_u10_u5_n1894 ), .ZN(_u10_u5_n2402 ) );
NAND3_X1 _u10_u5_U308  ( .A1(_u10_u5_n2329 ), .A2(_u10_u5_n2407 ), .A3(_u10_u5_n2255 ), .ZN(_u10_u5_n2403 ) );
NAND3_X1 _u10_u5_U307  ( .A1(_u10_u5_n1924 ), .A2(_u10_u5_n2405 ), .A3(_u10_u5_n2406 ), .ZN(_u10_u5_n2404 ) );
NAND3_X1 _u10_u5_U306  ( .A1(_u10_u5_n2402 ), .A2(_u10_u5_n2403 ), .A3(_u10_u5_n2404 ), .ZN(_u10_u5_n2393 ) );
INV_X1 _u10_u5_U305  ( .A(_u10_u5_n1932 ), .ZN(_u10_u5_n2399 ) );
NOR2_X1 _u10_u5_U304  ( .A1(_u10_u5_n2401 ), .A2(_u10_u5_n2161 ), .ZN(_u10_u5_n2400 ) );
NOR2_X1 _u10_u5_U303  ( .A1(_u10_u5_n2399 ), .A2(_u10_u5_n2400 ), .ZN(_u10_u5_n2394 ) );
NOR2_X1 _u10_u5_U302  ( .A1(_u10_u5_n2110 ), .A2(_u10_u5_n2398 ), .ZN(_u10_u5_n2397 ) );
NOR2_X1 _u10_u5_U301  ( .A1(_u10_u5_n2396 ), .A2(_u10_u5_n2397 ), .ZN(_u10_u5_n2395 ) );
NOR4_X1 _u10_u5_U300  ( .A1(_u10_u5_n2392 ), .A2(_u10_u5_n2393 ), .A3(_u10_u5_n2394 ), .A4(_u10_u5_n2395 ), .ZN(_u10_u5_n2391 ) );
NAND4_X1 _u10_u5_U299  ( .A1(_u10_u5_n2388 ), .A2(_u10_u5_n2389 ), .A3(_u10_u5_n2390 ), .A4(_u10_u5_n2391 ), .ZN(_u10_u5_n2387 ) );
MUX2_X1 _u10_u5_U298  ( .A(_u10_u5_n2387 ), .B(_u10_SYNOPSYS_UNCONNECTED_20 ), .S(_u10_u5_n1819 ), .Z(_u10_u5_n1810 ) );
NAND2_X1 _u10_u5_U297  ( .A1(_u10_u5_n2386 ), .A2(_u10_u5_n2007 ), .ZN(_u10_u5_n2369 ) );
AND2_X1 _u10_u5_U296  ( .A1(1'b0), .A2(_u10_u5_n2195 ), .ZN(_u10_u5_n2308 ));
NAND2_X1 _u10_u5_U295  ( .A1(_u10_u5_n2308 ), .A2(_u10_u5_n2036 ), .ZN(_u10_u5_n2384 ) );
AND2_X1 _u10_u5_U294  ( .A1(_u10_u5_n2384 ), .A2(_u10_u5_n2385 ), .ZN(_u10_u5_n2275 ) );
AND4_X1 _u10_u5_U293  ( .A1(_u10_u5_n2275 ), .A2(_u10_u5_n2286 ), .A3(_u10_u5_n2383 ), .A4(_u10_u5_n2285 ), .ZN(_u10_u5_n2225 ) );
NAND3_X1 _u10_u5_U292  ( .A1(_u10_u5_n2195 ), .A2(_u10_u5_n2223 ), .A3(1'b0),.ZN(_u10_u5_n2021 ) );
INV_X1 _u10_u5_U291  ( .A(_u10_u5_n2021 ), .ZN(_u10_u5_n2167 ) );
NAND2_X1 _u10_u5_U290  ( .A1(_u10_u5_n2036 ), .A2(_u10_u5_n2167 ), .ZN(_u10_u5_n1970 ) );
AND3_X1 _u10_u5_U289  ( .A1(_u10_u5_n1970 ), .A2(_u10_u5_n2164 ), .A3(_u10_u5_n2382 ), .ZN(_u10_u5_n2381 ) );
NAND4_X1 _u10_u5_U288  ( .A1(_u10_u5_n2225 ), .A2(_u10_u5_n2379 ), .A3(_u10_u5_n2380 ), .A4(_u10_u5_n2381 ), .ZN(_u10_u5_n2378 ) );
NAND2_X1 _u10_u5_U287  ( .A1(_u10_u5_n1967 ), .A2(_u10_u5_n2378 ), .ZN(_u10_u5_n2370 ) );
NAND2_X1 _u10_u5_U286  ( .A1(_u10_u5_n2081 ), .A2(_u10_u5_n2377 ), .ZN(_u10_u5_n2371 ) );
NOR2_X1 _u10_u5_U285  ( .A1(_u10_u5_n2375 ), .A2(_u10_u5_n2376 ), .ZN(_u10_u5_n2373 ) );
NOR2_X1 _u10_u5_U284  ( .A1(_u10_u5_n2373 ), .A2(_u10_u5_n2374 ), .ZN(_u10_u5_n2372 ) );
NAND4_X1 _u10_u5_U283  ( .A1(_u10_u5_n2369 ), .A2(_u10_u5_n2370 ), .A3(_u10_u5_n2371 ), .A4(_u10_u5_n2372 ), .ZN(_u10_u5_n2309 ) );
NOR2_X1 _u10_u5_U282  ( .A1(_u10_u5_n2000 ), .A2(_u10_u5_n2368 ), .ZN(_u10_u5_n2360 ) );
NOR2_X1 _u10_u5_U281  ( .A1(_u10_u5_n2366 ), .A2(_u10_u5_n2367 ), .ZN(_u10_u5_n2361 ) );
NOR2_X1 _u10_u5_U280  ( .A1(_u10_u5_n1868 ), .A2(_u10_u5_n2365 ), .ZN(_u10_u5_n2362 ) );
NOR2_X1 _u10_u5_U279  ( .A1(_u10_u5_n2364 ), .A2(_u10_u5_n1859 ), .ZN(_u10_u5_n2363 ) );
NOR4_X1 _u10_u5_U278  ( .A1(_u10_u5_n2360 ), .A2(_u10_u5_n2361 ), .A3(_u10_u5_n2362 ), .A4(_u10_u5_n2363 ), .ZN(_u10_u5_n2316 ) );
NOR2_X1 _u10_u5_U277  ( .A1(_u10_u5_n2359 ), .A2(_u10_u5_n1970 ), .ZN(_u10_u5_n2351 ) );
NOR2_X1 _u10_u5_U276  ( .A1(_u10_u5_n2358 ), .A2(_u10_u5_n1840 ), .ZN(_u10_u5_n2352 ) );
NOR2_X1 _u10_u5_U275  ( .A1(_u10_u5_n2356 ), .A2(_u10_u5_n2357 ), .ZN(_u10_u5_n2353 ) );
NOR2_X1 _u10_u5_U274  ( .A1(_u10_u5_n1836 ), .A2(_u10_u5_n2355 ), .ZN(_u10_u5_n2354 ) );
NOR4_X1 _u10_u5_U273  ( .A1(_u10_u5_n2351 ), .A2(_u10_u5_n2352 ), .A3(_u10_u5_n2353 ), .A4(_u10_u5_n2354 ), .ZN(_u10_u5_n2317 ) );
NOR2_X1 _u10_u5_U272  ( .A1(_u10_u5_n1873 ), .A2(_u10_u5_n2101 ), .ZN(_u10_u5_n2349 ) );
NOR2_X1 _u10_u5_U271  ( .A1(_u10_u5_n2349 ), .A2(_u10_u5_n2350 ), .ZN(_u10_u5_n2338 ) );
NOR2_X1 _u10_u5_U270  ( .A1(_u10_u5_n2347 ), .A2(_u10_u5_n2348 ), .ZN(_u10_u5_n2345 ) );
NOR2_X1 _u10_u5_U269  ( .A1(_u10_u5_n2345 ), .A2(_u10_u5_n2346 ), .ZN(_u10_u5_n2339 ) );
NOR2_X1 _u10_u5_U268  ( .A1(_u10_u5_n2344 ), .A2(_u10_u5_n2142 ), .ZN(_u10_u5_n2340 ) );
NOR2_X1 _u10_u5_U267  ( .A1(_u10_u5_n2342 ), .A2(_u10_u5_n2343 ), .ZN(_u10_u5_n2341 ) );
NOR4_X1 _u10_u5_U266  ( .A1(_u10_u5_n2338 ), .A2(_u10_u5_n2339 ), .A3(_u10_u5_n2340 ), .A4(_u10_u5_n2341 ), .ZN(_u10_u5_n2318 ) );
INV_X1 _u10_u5_U265  ( .A(_u10_u5_n2337 ), .ZN(_u10_u5_n2320 ) );
NOR2_X1 _u10_u5_U264  ( .A1(_u10_u5_n1970 ), .A2(1'b0), .ZN(_u10_u5_n2027 ));
INV_X1 _u10_u5_U263  ( .A(_u10_u5_n2027 ), .ZN(_u10_u5_n2331 ) );
NOR2_X1 _u10_u5_U262  ( .A1(_u10_u5_n2174 ), .A2(_u10_u5_n2216 ), .ZN(_u10_u5_n2333 ) );
AND2_X1 _u10_u5_U261  ( .A1(_u10_u5_n1928 ), .A2(_u10_u5_n2336 ), .ZN(_u10_u5_n2334 ) );
NOR4_X1 _u10_u5_U260  ( .A1(_u10_u5_n1937 ), .A2(_u10_u5_n2333 ), .A3(_u10_u5_n2334 ), .A4(_u10_u5_n2335 ), .ZN(_u10_u5_n2332 ) );
NOR3_X1 _u10_u5_U259  ( .A1(_u10_u5_n2331 ), .A2(_u10_u5_n2332 ), .A3(_u10_u5_n1915 ), .ZN(_u10_u5_n2321 ) );
NOR3_X1 _u10_u5_U258  ( .A1(_u10_u5_n2291 ), .A2(_u10_u5_n2330 ), .A3(_u10_u5_n2021 ), .ZN(_u10_u5_n2322 ) );
NOR2_X1 _u10_u5_U257  ( .A1(_u10_u5_n2329 ), .A2(_u10_u5_n2169 ), .ZN(_u10_u5_n2324 ) );
NOR2_X1 _u10_u5_U256  ( .A1(1'b0), .A2(_u10_u5_n2328 ), .ZN(_u10_u5_n2327 ));
NOR2_X1 _u10_u5_U255  ( .A1(_u10_u5_n2326 ), .A2(_u10_u5_n2327 ), .ZN(_u10_u5_n2325 ) );
NOR3_X1 _u10_u5_U254  ( .A1(_u10_u5_n2324 ), .A2(1'b0), .A3(_u10_u5_n2325 ),.ZN(_u10_u5_n2323 ) );
NOR4_X1 _u10_u5_U253  ( .A1(_u10_u5_n2320 ), .A2(_u10_u5_n2321 ), .A3(_u10_u5_n2322 ), .A4(_u10_u5_n2323 ), .ZN(_u10_u5_n2319 ) );
AND4_X1 _u10_u5_U252  ( .A1(_u10_u5_n2316 ), .A2(_u10_u5_n2317 ), .A3(_u10_u5_n2318 ), .A4(_u10_u5_n2319 ), .ZN(_u10_u5_n1991 ) );
INV_X1 _u10_u5_U251  ( .A(_u10_u5_n2315 ), .ZN(_u10_u5_n2313 ) );
NAND3_X1 _u10_u5_U250  ( .A1(_u10_u5_n1991 ), .A2(_u10_u5_n2313 ), .A3(_u10_u5_n2314 ), .ZN(_u10_u5_n2310 ) );
NOR4_X1 _u10_u5_U249  ( .A1(_u10_u5_n2309 ), .A2(_u10_u5_n2310 ), .A3(_u10_u5_n2311 ), .A4(_u10_u5_n2312 ), .ZN(_u10_u5_n2117 ) );
NAND3_X1 _u10_u5_U248  ( .A1(_u10_u5_n2108 ), .A2(_u10_u5_n2107 ), .A3(_u10_u5_n2308 ), .ZN(_u10_u5_n2217 ) );
NOR3_X1 _u10_u5_U247  ( .A1(_u10_u5_n2306 ), .A2(_u10_u5_n2307 ), .A3(_u10_u5_n2027 ), .ZN(_u10_u5_n2277 ) );
NAND3_X1 _u10_u5_U246  ( .A1(_u10_u5_n2217 ), .A2(_u10_u5_n2305 ), .A3(_u10_u5_n2277 ), .ZN(_u10_u5_n2157 ) );
NAND2_X1 _u10_u5_U245  ( .A1(_u10_u5_n2089 ), .A2(_u10_u5_n2157 ), .ZN(_u10_u5_n2296 ) );
INV_X1 _u10_u5_U244  ( .A(_u10_u5_n2304 ), .ZN(_u10_u5_n2297 ) );
NOR2_X1 _u10_u5_U243  ( .A1(_u10_u5_n2302 ), .A2(_u10_u5_n2303 ), .ZN(_u10_u5_n2299 ) );
NOR3_X1 _u10_u5_U242  ( .A1(_u10_u5_n2299 ), .A2(_u10_u5_n2300 ), .A3(_u10_u5_n2301 ), .ZN(_u10_u5_n2298 ) );
NAND4_X1 _u10_u5_U241  ( .A1(_u10_u5_n2295 ), .A2(_u10_u5_n2296 ), .A3(_u10_u5_n2297 ), .A4(_u10_u5_n2298 ), .ZN(_u10_u5_n2294 ) );
NAND2_X1 _u10_u5_U240  ( .A1(_u10_u5_n2293 ), .A2(_u10_u5_n2294 ), .ZN(_u10_u5_n2257 ) );
NAND2_X1 _u10_u5_U239  ( .A1(_u10_u5_n2165 ), .A2(_u10_u5_n2166 ), .ZN(_u10_u5_n2288 ) );
NAND2_X1 _u10_u5_U238  ( .A1(_u10_u5_n2078 ), .A2(_u10_u5_n2279 ), .ZN(_u10_u5_n2292 ) );
NAND2_X1 _u10_u5_U237  ( .A1(_u10_u5_n2291 ), .A2(_u10_u5_n2292 ), .ZN(_u10_u5_n2290 ) );
NAND2_X1 _u10_u5_U236  ( .A1(_u10_u5_n2059 ), .A2(_u10_u5_n2290 ), .ZN(_u10_u5_n2289 ) );
NAND2_X1 _u10_u5_U235  ( .A1(_u10_u5_n2288 ), .A2(_u10_u5_n2289 ), .ZN(_u10_u5_n2201 ) );
NAND2_X1 _u10_u5_U234  ( .A1(1'b0), .A2(_u10_u5_n2201 ), .ZN(_u10_u5_n2258 ));
INV_X1 _u10_u5_U233  ( .A(_u10_u5_n2287 ), .ZN(_u10_u5_n2283 ) );
AND4_X1 _u10_u5_U232  ( .A1(_u10_u5_n2285 ), .A2(_u10_u5_n2226 ), .A3(_u10_u5_n1970 ), .A4(_u10_u5_n2286 ), .ZN(_u10_u5_n2284 ) );
NAND4_X1 _u10_u5_U231  ( .A1(_u10_u5_n2281 ), .A2(_u10_u5_n2282 ), .A3(_u10_u5_n2283 ), .A4(_u10_u5_n2284 ), .ZN(_u10_u5_n2280 ) );
NAND2_X1 _u10_u5_U230  ( .A1(_u10_u5_n2279 ), .A2(_u10_u5_n2280 ), .ZN(_u10_u5_n2259 ) );
NAND4_X1 _u10_u5_U229  ( .A1(_u10_u5_n2275 ), .A2(_u10_u5_n2276 ), .A3(_u10_u5_n2277 ), .A4(_u10_u5_n2278 ), .ZN(_u10_u5_n2271 ) );
NAND2_X1 _u10_u5_U228  ( .A1(_u10_u5_n1933 ), .A2(_u10_u5_n2164 ), .ZN(_u10_u5_n2272 ) );
NOR2_X1 _u10_u5_U227  ( .A1(_u10_u5_n2274 ), .A2(_u10_u5_n2130 ), .ZN(_u10_u5_n2273 ) );
NOR4_X1 _u10_u5_U226  ( .A1(_u10_u5_n2271 ), .A2(_u10_u5_n2272 ), .A3(_u10_u5_n1978 ), .A4(_u10_u5_n2273 ), .ZN(_u10_u5_n2270 ) );
NOR2_X1 _u10_u5_U225  ( .A1(_u10_u5_n2270 ), .A2(_u10_u5_n2025 ), .ZN(_u10_u5_n2261 ) );
NAND3_X1 _u10_u5_U224  ( .A1(_u10_u5_n1933 ), .A2(_u10_u5_n1936 ), .A3(_u10_u5_n2269 ), .ZN(_u10_u5_n2268 ) );
NOR3_X1 _u10_u5_U223  ( .A1(_u10_u5_n2268 ), .A2(_u10_u5_n1844 ), .A3(_u10_u5_n2157 ), .ZN(_u10_u5_n2267 ) );
NOR2_X1 _u10_u5_U222  ( .A1(1'b0), .A2(_u10_u5_n2267 ), .ZN(_u10_u5_n2265 ));
NOR3_X1 _u10_u5_U221  ( .A1(_u10_u5_n2264 ), .A2(_u10_u5_n2265 ), .A3(_u10_u5_n2266 ), .ZN(_u10_u5_n2263 ) );
NOR2_X1 _u10_u5_U220  ( .A1(_u10_u5_n2263 ), .A2(_u10_u5_n1843 ), .ZN(_u10_u5_n2262 ) );
NOR2_X1 _u10_u5_U219  ( .A1(_u10_u5_n2261 ), .A2(_u10_u5_n2262 ), .ZN(_u10_u5_n2260 ) );
NAND4_X1 _u10_u5_U218  ( .A1(_u10_u5_n2257 ), .A2(_u10_u5_n2258 ), .A3(_u10_u5_n2259 ), .A4(_u10_u5_n2260 ), .ZN(_u10_u5_n2230 ) );
INV_X1 _u10_u5_U217  ( .A(_u10_u5_n2217 ), .ZN(_u10_u5_n2242 ) );
NAND2_X1 _u10_u5_U216  ( .A1(_u10_u5_n2168 ), .A2(_u10_u5_n2169 ), .ZN(_u10_u5_n2244 ) );
NAND2_X1 _u10_u5_U215  ( .A1(_u10_u5_n2255 ), .A2(_u10_u5_n2256 ), .ZN(_u10_u5_n2245 ) );
NAND2_X1 _u10_u5_U214  ( .A1(_u10_u5_n2253 ), .A2(_u10_u5_n2254 ), .ZN(_u10_u5_n2252 ) );
NAND2_X1 _u10_u5_U213  ( .A1(_u10_u5_n2251 ), .A2(_u10_u5_n2252 ), .ZN(_u10_u5_n2246 ) );
NAND2_X1 _u10_u5_U212  ( .A1(_u10_u5_n2152 ), .A2(_u10_u5_n1928 ), .ZN(_u10_u5_n2250 ) );
NAND2_X1 _u10_u5_U211  ( .A1(_u10_u5_n2249 ), .A2(_u10_u5_n2250 ), .ZN(_u10_u5_n2248 ) );
NAND2_X1 _u10_u5_U210  ( .A1(_u10_u5_n2105 ), .A2(_u10_u5_n2248 ), .ZN(_u10_u5_n2247 ) );
NAND4_X1 _u10_u5_U209  ( .A1(_u10_u5_n2244 ), .A2(_u10_u5_n2245 ), .A3(_u10_u5_n2246 ), .A4(_u10_u5_n2247 ), .ZN(_u10_u5_n2243 ) );
NAND2_X1 _u10_u5_U208  ( .A1(_u10_u5_n2242 ), .A2(_u10_u5_n2243 ), .ZN(_u10_u5_n2237 ) );
NAND2_X1 _u10_u5_U207  ( .A1(1'b0), .A2(_u10_u5_n2241 ), .ZN(_u10_u5_n2238 ));
NAND2_X1 _u10_u5_U206  ( .A1(_u10_u5_n2214 ), .A2(_u10_u5_n2240 ), .ZN(_u10_u5_n2239 ) );
NAND3_X1 _u10_u5_U205  ( .A1(_u10_u5_n2237 ), .A2(_u10_u5_n2238 ), .A3(_u10_u5_n2239 ), .ZN(_u10_u5_n2231 ) );
AND2_X1 _u10_u5_U204  ( .A1(_u10_u5_n2200 ), .A2(_u10_u5_n2236 ), .ZN(_u10_u5_n2232 ) );
NOR2_X1 _u10_u5_U203  ( .A1(_u10_u5_n2234 ), .A2(_u10_u5_n2235 ), .ZN(_u10_u5_n2233 ) );
NOR4_X1 _u10_u5_U202  ( .A1(_u10_u5_n2230 ), .A2(_u10_u5_n2231 ), .A3(_u10_u5_n2232 ), .A4(_u10_u5_n2233 ), .ZN(_u10_u5_n2118 ) );
NAND2_X1 _u10_u5_U201  ( .A1(_u10_u5_n2214 ), .A2(_u10_u5_n2049 ), .ZN(_u10_u5_n2229 ) );
NAND2_X1 _u10_u5_U200  ( .A1(_u10_u5_n2228 ), .A2(_u10_u5_n2229 ), .ZN(_u10_u5_n2227 ) );
NAND2_X1 _u10_u5_U199  ( .A1(_u10_u5_n2043 ), .A2(_u10_u5_n2227 ), .ZN(_u10_u5_n2204 ) );
NAND2_X1 _u10_u5_U198  ( .A1(_u10_u5_n2225 ), .A2(_u10_u5_n2226 ), .ZN(_u10_u5_n2224 ) );
NAND2_X1 _u10_u5_U197  ( .A1(_u10_u5_n1899 ), .A2(_u10_u5_n2224 ), .ZN(_u10_u5_n2205 ) );
NAND2_X1 _u10_u5_U196  ( .A1(_u10_u5_n2222 ), .A2(_u10_u5_n2223 ), .ZN(_u10_u5_n1870 ) );
NAND4_X1 _u10_u5_U195  ( .A1(_u10_u5_n2220 ), .A2(_u10_u5_n2131 ), .A3(_u10_u5_n2221 ), .A4(_u10_u5_n1870 ), .ZN(_u10_u5_n2219 ) );
NAND2_X1 _u10_u5_U194  ( .A1(_u10_u5_n2218 ), .A2(_u10_u5_n2219 ), .ZN(_u10_u5_n2206 ) );
NOR2_X1 _u10_u5_U193  ( .A1(_u10_u5_n1925 ), .A2(_u10_u5_n2217 ), .ZN(_u10_u5_n2215 ) );
NOR4_X1 _u10_u5_U192  ( .A1(_u10_u5_n2213 ), .A2(_u10_u5_n2214 ), .A3(_u10_u5_n2215 ), .A4(_u10_u5_n2216 ), .ZN(_u10_u5_n2211 ) );
NOR2_X1 _u10_u5_U191  ( .A1(_u10_u5_n2211 ), .A2(_u10_u5_n2212 ), .ZN(_u10_u5_n2208 ) );
NOR2_X1 _u10_u5_U190  ( .A1(_u10_u5_n1888 ), .A2(_u10_u5_n2210 ), .ZN(_u10_u5_n2209 ) );
NOR2_X1 _u10_u5_U189  ( .A1(_u10_u5_n2208 ), .A2(_u10_u5_n2209 ), .ZN(_u10_u5_n2207 ) );
NAND4_X1 _u10_u5_U188  ( .A1(_u10_u5_n2204 ), .A2(_u10_u5_n2205 ), .A3(_u10_u5_n2206 ), .A4(_u10_u5_n2207 ), .ZN(_u10_u5_n2170 ) );
OR2_X1 _u10_u5_U187  ( .A1(_u10_u5_n2202 ), .A2(_u10_u5_n2203 ), .ZN(_u10_u5_n2197 ) );
NAND2_X1 _u10_u5_U186  ( .A1(1'b0), .A2(_u10_u5_n2201 ), .ZN(_u10_u5_n2198 ));
NAND2_X1 _u10_u5_U185  ( .A1(_u10_u5_n2063 ), .A2(_u10_u5_n2200 ), .ZN(_u10_u5_n2199 ) );
NAND3_X1 _u10_u5_U184  ( .A1(_u10_u5_n2197 ), .A2(_u10_u5_n2198 ), .A3(_u10_u5_n2199 ), .ZN(_u10_u5_n2196 ) );
NAND2_X1 _u10_u5_U183  ( .A1(_u10_u5_n2195 ), .A2(_u10_u5_n2196 ), .ZN(_u10_u5_n2180 ) );
NAND2_X1 _u10_u5_U182  ( .A1(_u10_u5_n2195 ), .A2(_u10_u5_n1918 ), .ZN(_u10_u5_n2192 ) );
NAND4_X1 _u10_u5_U181  ( .A1(_u10_u5_n2192 ), .A2(_u10_u5_n2021 ), .A3(_u10_u5_n2193 ), .A4(_u10_u5_n2194 ), .ZN(_u10_u5_n2188 ) );
NAND2_X1 _u10_u5_U180  ( .A1(_u10_u5_n2188 ), .A2(_u10_u5_n2191 ), .ZN(_u10_u5_n2181 ) );
NAND2_X1 _u10_u5_U179  ( .A1(1'b0), .A2(_u10_u5_n2190 ), .ZN(_u10_u5_n2185 ));
NAND2_X1 _u10_u5_U178  ( .A1(_u10_u5_n2189 ), .A2(_u10_SYNOPSYS_UNCONNECTED_21 ), .ZN(_u10_u5_n2186 ) );
INV_X1 _u10_u5_U177  ( .A(_u10_u5_n2188 ), .ZN(_u10_u5_n2187 ) );
NAND3_X1 _u10_u5_U176  ( .A1(_u10_u5_n2185 ), .A2(_u10_u5_n2186 ), .A3(_u10_u5_n2187 ), .ZN(_u10_u5_n2184 ) );
NAND2_X1 _u10_u5_U175  ( .A1(_u10_u5_n2183 ), .A2(_u10_u5_n2184 ), .ZN(_u10_u5_n2182 ) );
NAND3_X1 _u10_u5_U174  ( .A1(_u10_u5_n2180 ), .A2(_u10_u5_n2181 ), .A3(_u10_u5_n2182 ), .ZN(_u10_u5_n2171 ) );
INV_X1 _u10_u5_U173  ( .A(_u10_u5_n2179 ), .ZN(_u10_u5_n1963 ) );
NOR2_X1 _u10_u5_U172  ( .A1(_u10_u5_n1963 ), .A2(_u10_u5_n2178 ), .ZN(_u10_u5_n2172 ) );
INV_X1 _u10_u5_U171  ( .A(_u10_u5_n2177 ), .ZN(_u10_u5_n2176 ) );
NOR3_X1 _u10_u5_U170  ( .A1(_u10_u5_n2174 ), .A2(_u10_u5_n2175 ), .A3(_u10_u5_n2176 ), .ZN(_u10_u5_n2173 ) );
NOR4_X1 _u10_u5_U169  ( .A1(_u10_u5_n2170 ), .A2(_u10_u5_n2171 ), .A3(_u10_u5_n2172 ), .A4(_u10_u5_n2173 ), .ZN(_u10_u5_n2119 ) );
NAND3_X1 _u10_u5_U168  ( .A1(_u10_u5_n2168 ), .A2(_u10_u5_n2169 ), .A3(1'b0),.ZN(_u10_u5_n2148 ) );
NAND3_X1 _u10_u5_U167  ( .A1(_u10_u5_n2165 ), .A2(_u10_u5_n2166 ), .A3(_u10_u5_n2167 ), .ZN(_u10_u5_n2149 ) );
NAND4_X1 _u10_u5_U166  ( .A1(_u10_u5_n2162 ), .A2(_u10_u5_n1933 ), .A3(_u10_u5_n2163 ), .A4(_u10_u5_n2164 ), .ZN(_u10_u5_n2160 ) );
NOR4_X1 _u10_u5_U165  ( .A1(_u10_u5_n2160 ), .A2(_u10_u5_n2157 ), .A3(_u10_u5_n1844 ), .A4(_u10_u5_n2161 ), .ZN(_u10_u5_n2158 ) );
NOR2_X1 _u10_u5_U164  ( .A1(_u10_u5_n2158 ), .A2(_u10_u5_n2159 ), .ZN(_u10_u5_n2153 ) );
INV_X1 _u10_u5_U163  ( .A(_u10_u5_n2157 ), .ZN(_u10_u5_n2129 ) );
NOR3_X1 _u10_u5_U162  ( .A1(_u10_u5_n2155 ), .A2(_u10_u5_n2129 ), .A3(_u10_u5_n2156 ), .ZN(_u10_u5_n2154 ) );
NOR2_X1 _u10_u5_U161  ( .A1(_u10_u5_n2153 ), .A2(_u10_u5_n2154 ), .ZN(_u10_u5_n2150 ) );
NAND3_X1 _u10_u5_U160  ( .A1(1'b0), .A2(_u10_u5_n1928 ), .A3(_u10_u5_n2152 ),.ZN(_u10_u5_n2151 ) );
NAND4_X1 _u10_u5_U159  ( .A1(_u10_u5_n2148 ), .A2(_u10_u5_n2149 ), .A3(_u10_u5_n2150 ), .A4(_u10_u5_n2151 ), .ZN(_u10_u5_n2121 ) );
NAND2_X1 _u10_u5_U158  ( .A1(_u10_u5_n2107 ), .A2(_u10_u5_n2147 ), .ZN(_u10_u5_n2146 ) );
NAND2_X1 _u10_u5_U157  ( .A1(_u10_u5_n2145 ), .A2(_u10_u5_n2146 ), .ZN(_u10_u5_n2144 ) );
NAND2_X1 _u10_u5_U156  ( .A1(_u10_u5_n2143 ), .A2(_u10_u5_n2144 ), .ZN(_u10_u5_n2134 ) );
NAND2_X1 _u10_u5_U155  ( .A1(_u10_u5_n2141 ), .A2(_u10_u5_n2142 ), .ZN(_u10_u5_n2140 ) );
NAND2_X1 _u10_u5_U154  ( .A1(_u10_u5_n2139 ), .A2(_u10_u5_n2140 ), .ZN(_u10_u5_n2135 ) );
OR2_X1 _u10_u5_U153  ( .A1(_u10_u5_n2110 ), .A2(_u10_u5_n1911 ), .ZN(_u10_u5_n2137 ) );
NAND2_X1 _u10_u5_U152  ( .A1(_u10_u5_n2137 ), .A2(_u10_u5_n2138 ), .ZN(_u10_u5_n2136 ) );
NAND3_X1 _u10_u5_U151  ( .A1(_u10_u5_n2134 ), .A2(_u10_u5_n2135 ), .A3(_u10_u5_n2136 ), .ZN(_u10_u5_n2122 ) );
NOR2_X1 _u10_u5_U150  ( .A1(_u10_u5_n2133 ), .A2(_u10_u5_n1891 ), .ZN(_u10_u5_n2132 ) );
NOR2_X1 _u10_u5_U149  ( .A1(_u10_u5_n2131 ), .A2(_u10_u5_n2132 ), .ZN(_u10_u5_n2123 ) );
NOR2_X1 _u10_u5_U148  ( .A1(_u10_u5_n2129 ), .A2(_u10_u5_n2130 ), .ZN(_u10_u5_n2127 ) );
NOR2_X1 _u10_u5_U147  ( .A1(_u10_u5_n2127 ), .A2(_u10_u5_n2128 ), .ZN(_u10_u5_n2125 ) );
NOR2_X1 _u10_u5_U146  ( .A1(_u10_u5_n2125 ), .A2(_u10_u5_n2126 ), .ZN(_u10_u5_n2124 ) );
NOR4_X1 _u10_u5_U145  ( .A1(_u10_u5_n2121 ), .A2(_u10_u5_n2122 ), .A3(_u10_u5_n2123 ), .A4(_u10_u5_n2124 ), .ZN(_u10_u5_n2120 ) );
NAND4_X1 _u10_u5_U144  ( .A1(_u10_u5_n2117 ), .A2(_u10_u5_n2118 ), .A3(_u10_u5_n2119 ), .A4(_u10_u5_n2120 ), .ZN(_u10_u5_n2116 ) );
MUX2_X1 _u10_u5_U143  ( .A(_u10_u5_n2116 ), .B(_u10_SYNOPSYS_UNCONNECTED_21 ), .S(_u10_u5_n1819 ), .Z(_u10_u5_n1811 ) );
INV_X1 _u10_u5_U142  ( .A(_u10_u5_n2115 ), .ZN(_u10_u5_n2006 ) );
NOR3_X1 _u10_u5_U141  ( .A1(_u10_u5_n2006 ), .A2(_u10_u5_n2114 ), .A3(_u10_u5_n2081 ), .ZN(_u10_u5_n1854 ) );
NAND2_X1 _u10_u5_U140  ( .A1(_u10_u5_n2112 ), .A2(_u10_u5_n2113 ), .ZN(_u10_u5_n1872 ) );
INV_X1 _u10_u5_U139  ( .A(_u10_u5_n1872 ), .ZN(_u10_u5_n1882 ) );
NAND4_X1 _u10_u5_U138  ( .A1(_u10_u5_n1854 ), .A2(_u10_u5_n1882 ), .A3(_u10_u5_n2111 ), .A4(_u10_u5_n1868 ), .ZN(_u10_u5_n2109 ) );
NAND2_X1 _u10_u5_U137  ( .A1(_u10_u5_n2109 ), .A2(_u10_u5_n2110 ), .ZN(_u10_u5_n2098 ) );
NAND2_X1 _u10_u5_U136  ( .A1(1'b0), .A2(_u10_u5_n1983 ), .ZN(_u10_u5_n2023 ));
INV_X1 _u10_u5_U135  ( .A(_u10_u5_n2023 ), .ZN(_u10_u5_n2035 ) );
NAND3_X1 _u10_u5_U134  ( .A1(_u10_u5_n2035 ), .A2(_u10_u5_n2107 ), .A3(_u10_u5_n2108 ), .ZN(_u10_u5_n1916 ) );
INV_X1 _u10_u5_U133  ( .A(_u10_u5_n1916 ), .ZN(_u10_u5_n2093 ) );
NAND3_X1 _u10_u5_U132  ( .A1(_u10_u5_n2105 ), .A2(_u10_u5_n2106 ), .A3(_u10_u5_n2093 ), .ZN(_u10_u5_n2039 ) );
NAND2_X1 _u10_u5_U131  ( .A1(_u10_u5_n2039 ), .A2(_u10_u5_n1930 ), .ZN(_u10_u5_n2104 ) );
NAND2_X1 _u10_u5_U130  ( .A1(_u10_u5_n2103 ), .A2(_u10_u5_n2104 ), .ZN(_u10_u5_n1863 ) );
OR2_X1 _u10_u5_U129  ( .A1(_u10_u5_n1863 ), .A2(_u10_u5_n2102 ), .ZN(_u10_u5_n2099 ) );
NAND2_X1 _u10_u5_U128  ( .A1(_u10_u5_n1890 ), .A2(_u10_u5_n2101 ), .ZN(_u10_u5_n2100 ) );
NAND3_X1 _u10_u5_U127  ( .A1(_u10_u5_n2098 ), .A2(_u10_u5_n2099 ), .A3(_u10_u5_n2100 ), .ZN(_u10_u5_n2066 ) );
NAND4_X1 _u10_u5_U126  ( .A1(_u10_u5_n2095 ), .A2(_u10_u5_n2096 ), .A3(_u10_u5_n1896 ), .A4(_u10_u5_n2097 ), .ZN(_u10_u5_n2086 ) );
NOR4_X1 _u10_u5_U125  ( .A1(_u10_u5_n2093 ), .A2(_u10_u5_n2027 ), .A3(_u10_u5_n2094 ), .A4(_u10_u5_n2026 ), .ZN(_u10_u5_n1952 ) );
NOR2_X1 _u10_u5_U124  ( .A1(1'b0), .A2(_u10_u5_n1952 ), .ZN(_u10_u5_n1951 ));
INV_X1 _u10_u5_U123  ( .A(_u10_u5_n1951 ), .ZN(_u10_u5_n2090 ) );
NAND4_X1 _u10_u5_U122  ( .A1(_u10_u5_n2089 ), .A2(_u10_u5_n2090 ), .A3(_u10_u5_n2091 ), .A4(_u10_u5_n2092 ), .ZN(_u10_u5_n1893 ) );
NOR4_X1 _u10_u5_U121  ( .A1(_u10_u5_n2086 ), .A2(_u10_u5_n1893 ), .A3(_u10_u5_n2087 ), .A4(_u10_u5_n2088 ), .ZN(_u10_u5_n2084 ) );
NOR2_X1 _u10_u5_U120  ( .A1(_u10_u5_n2084 ), .A2(_u10_u5_n2085 ), .ZN(_u10_u5_n2067 ) );
NOR2_X1 _u10_u5_U119  ( .A1(_u10_u5_n2083 ), .A2(_u10_u5_n1869 ), .ZN(_u10_u5_n2068 ) );
NAND2_X1 _u10_u5_U118  ( .A1(_u10_u5_n2081 ), .A2(_u10_u5_n2082 ), .ZN(_u10_u5_n2075 ) );
NAND2_X1 _u10_u5_U117  ( .A1(_u10_u5_n2035 ), .A2(_u10_u5_n2019 ), .ZN(_u10_u5_n2060 ) );
NAND2_X1 _u10_u5_U116  ( .A1(_u10_u5_n2080 ), .A2(_u10_u5_n2060 ), .ZN(_u10_u5_n2079 ) );
NAND2_X1 _u10_u5_U115  ( .A1(_u10_u5_n2078 ), .A2(_u10_u5_n2079 ), .ZN(_u10_u5_n2076 ) );
NAND4_X1 _u10_u5_U114  ( .A1(_u10_u5_n2075 ), .A2(_u10_u5_n2076 ), .A3(_u10_u5_n1970 ), .A4(_u10_u5_n2077 ), .ZN(_u10_u5_n2072 ) );
NOR4_X1 _u10_u5_U113  ( .A1(_u10_u5_n2072 ), .A2(_u10_u5_n2073 ), .A3(_u10_u5_n1975 ), .A4(_u10_u5_n2074 ), .ZN(_u10_u5_n2070 ) );
NOR2_X1 _u10_u5_U112  ( .A1(_u10_u5_n2070 ), .A2(_u10_u5_n2071 ), .ZN(_u10_u5_n2069 ) );
NOR4_X1 _u10_u5_U111  ( .A1(_u10_u5_n2066 ), .A2(_u10_u5_n2067 ), .A3(_u10_u5_n2068 ), .A4(_u10_u5_n2069 ), .ZN(_u10_u5_n1820 ) );
NAND2_X1 _u10_u5_U110  ( .A1(1'b0), .A2(_u10_u5_n1983 ), .ZN(_u10_u5_n2065 ));
NAND4_X1 _u10_u5_U109  ( .A1(_u10_u5_n2065 ), .A2(_u10_u5_n2023 ), .A3(_u10_u5_n2021 ), .A4(_u10_u5_n2052 ), .ZN(_u10_u5_n2064 ) );
NAND2_X1 _u10_u5_U108  ( .A1(_u10_u5_n2063 ), .A2(_u10_u5_n2064 ), .ZN(_u10_u5_n2040 ) );
NAND4_X1 _u10_u5_U107  ( .A1(_u10_u5_n2059 ), .A2(_u10_u5_n2060 ), .A3(_u10_u5_n2061 ), .A4(_u10_u5_n2062 ), .ZN(_u10_u5_n2058 ) );
NAND2_X1 _u10_u5_U106  ( .A1(_u10_u5_n2057 ), .A2(_u10_u5_n2058 ), .ZN(_u10_u5_n2041 ) );
NOR4_X1 _u10_u5_U105  ( .A1(1'b0), .A2(_u10_u5_n2054 ), .A3(_u10_u5_n2055 ),.A4(_u10_u5_n2056 ), .ZN(_u10_u5_n2053 ) );
NAND4_X1 _u10_u5_U104  ( .A1(_u10_u5_n2021 ), .A2(_u10_u5_n2052 ), .A3(_u10_u5_n2023 ), .A4(_u10_u5_n2053 ), .ZN(_u10_u5_n1964 ) );
INV_X1 _u10_u5_U103  ( .A(_u10_u5_n1964 ), .ZN(_u10_u5_n2045 ) );
NAND2_X1 _u10_u5_U102  ( .A1(_u10_u5_n2051 ), .A2(_u10_SYNOPSYS_UNCONNECTED_22 ), .ZN(_u10_u5_n2046 ) );
NAND2_X1 _u10_u5_U101  ( .A1(_u10_u5_n2049 ), .A2(_u10_u5_n2050 ), .ZN(_u10_u5_n2047 ) );
NAND4_X1 _u10_u5_U100  ( .A1(_u10_u5_n2045 ), .A2(_u10_u5_n2046 ), .A3(_u10_u5_n2047 ), .A4(_u10_u5_n2048 ), .ZN(_u10_u5_n2044 ) );
NAND2_X1 _u10_u5_U99  ( .A1(_u10_u5_n2043 ), .A2(_u10_u5_n2044 ), .ZN(_u10_u5_n2042 ) );
NAND3_X1 _u10_u5_U98  ( .A1(_u10_u5_n2040 ), .A2(_u10_u5_n2041 ), .A3(_u10_u5_n2042 ), .ZN(_u10_u5_n2009 ) );
AND2_X1 _u10_u5_U97  ( .A1(_u10_u5_n2038 ), .A2(_u10_u5_n2039 ), .ZN(_u10_u5_n1929 ) );
NOR2_X1 _u10_u5_U96  ( .A1(_u10_u5_n1929 ), .A2(_u10_u5_n2037 ), .ZN(_u10_u5_n2010 ) );
NAND2_X1 _u10_u5_U95  ( .A1(_u10_u5_n2035 ), .A2(_u10_u5_n2036 ), .ZN(_u10_u5_n1902 ) );
NAND3_X1 _u10_u5_U94  ( .A1(_u10_u5_n1902 ), .A2(_u10_u5_n2033 ), .A3(_u10_u5_n2034 ), .ZN(_u10_u5_n1973 ) );
NOR2_X1 _u10_u5_U93  ( .A1(_u10_u5_n1978 ), .A2(_u10_u5_n1973 ), .ZN(_u10_u5_n2032 ) );
NOR2_X1 _u10_u5_U92  ( .A1(1'b0), .A2(_u10_u5_n2032 ), .ZN(_u10_u5_n2028 ));
NOR2_X1 _u10_u5_U91  ( .A1(_u10_u5_n2030 ), .A2(_u10_u5_n2031 ), .ZN(_u10_u5_n2029 ) );
NOR4_X1 _u10_u5_U90  ( .A1(_u10_u5_n2026 ), .A2(_u10_u5_n2027 ), .A3(_u10_u5_n2028 ), .A4(_u10_u5_n2029 ), .ZN(_u10_u5_n2024 ) );
NOR2_X1 _u10_u5_U89  ( .A1(_u10_u5_n2024 ), .A2(_u10_u5_n2025 ), .ZN(_u10_u5_n2011 ) );
NAND3_X1 _u10_u5_U88  ( .A1(_u10_u5_n2021 ), .A2(_u10_u5_n2022 ), .A3(_u10_u5_n2023 ), .ZN(_u10_u5_n2020 ) );
AND2_X1 _u10_u5_U87  ( .A1(_u10_u5_n2019 ), .A2(_u10_u5_n2020 ), .ZN(_u10_u5_n1838 ) );
INV_X1 _u10_u5_U86  ( .A(_u10_u5_n2018 ), .ZN(_u10_u5_n2016 ) );
NOR4_X1 _u10_u5_U85  ( .A1(_u10_u5_n2015 ), .A2(_u10_u5_n1838 ), .A3(_u10_u5_n2016 ), .A4(_u10_u5_n2017 ), .ZN(_u10_u5_n2013 ) );
NOR2_X1 _u10_u5_U84  ( .A1(_u10_u5_n2013 ), .A2(_u10_u5_n2014 ), .ZN(_u10_u5_n2012 ) );
NOR4_X1 _u10_u5_U83  ( .A1(_u10_u5_n2009 ), .A2(_u10_u5_n2010 ), .A3(_u10_u5_n2011 ), .A4(_u10_u5_n2012 ), .ZN(_u10_u5_n1821 ) );
NAND2_X1 _u10_u5_U82  ( .A1(_u10_u5_n1924 ), .A2(_u10_u5_n2008 ), .ZN(_u10_u5_n1993 ) );
NAND2_X1 _u10_u5_U81  ( .A1(_u10_u5_n2006 ), .A2(_u10_u5_n2007 ), .ZN(_u10_u5_n1994 ) );
NAND2_X1 _u10_u5_U80  ( .A1(_u10_u5_n2004 ), .A2(_u10_u5_n2005 ), .ZN(_u10_u5_n1995 ) );
AND2_X1 _u10_u5_U79  ( .A1(_u10_u5_n2002 ), .A2(_u10_u5_n2003 ), .ZN(_u10_u5_n1998 ) );
NOR2_X1 _u10_u5_U78  ( .A1(_u10_u5_n2000 ), .A2(_u10_u5_n2001 ), .ZN(_u10_u5_n1999 ) );
NOR3_X1 _u10_u5_U77  ( .A1(_u10_u5_n1997 ), .A2(_u10_u5_n1998 ), .A3(_u10_u5_n1999 ), .ZN(_u10_u5_n1996 ) );
NAND4_X1 _u10_u5_U76  ( .A1(_u10_u5_n1993 ), .A2(_u10_u5_n1994 ), .A3(_u10_u5_n1995 ), .A4(_u10_u5_n1996 ), .ZN(_u10_u5_n1985 ) );
INV_X1 _u10_u5_U75  ( .A(_u10_u5_n1992 ), .ZN(_u10_u5_n1989 ) );
NAND3_X1 _u10_u5_U74  ( .A1(_u10_u5_n1989 ), .A2(_u10_u5_n1990 ), .A3(_u10_u5_n1991 ), .ZN(_u10_u5_n1986 ) );
NOR4_X1 _u10_u5_U73  ( .A1(_u10_u5_n1985 ), .A2(_u10_u5_n1986 ), .A3(_u10_u5_n1987 ), .A4(_u10_u5_n1988 ), .ZN(_u10_u5_n1822 ) );
INV_X1 _u10_u5_U72  ( .A(_u10_u5_n1984 ), .ZN(_u10_u5_n1980 ) );
NAND4_X1 _u10_u5_U71  ( .A1(_u10_u5_n1980 ), .A2(_u10_u5_n1981 ), .A3(_u10_u5_n1982 ), .A4(_u10_u5_n1983 ), .ZN(_u10_u5_n1941 ) );
NOR3_X1 _u10_u5_U70  ( .A1(_u10_u5_n1977 ), .A2(_u10_u5_n1978 ), .A3(_u10_u5_n1979 ), .ZN(_u10_u5_n1971 ) );
NOR4_X1 _u10_u5_U69  ( .A1(_u10_u5_n1973 ), .A2(_u10_u5_n1974 ), .A3(_u10_u5_n1975 ), .A4(_u10_u5_n1976 ), .ZN(_u10_u5_n1972 ) );
NAND4_X1 _u10_u5_U68  ( .A1(_u10_u5_n1969 ), .A2(_u10_u5_n1970 ), .A3(_u10_u5_n1971 ), .A4(_u10_u5_n1972 ), .ZN(_u10_u5_n1968 ) );
NAND2_X1 _u10_u5_U67  ( .A1(_u10_u5_n1967 ), .A2(_u10_u5_n1968 ), .ZN(_u10_u5_n1942 ) );
NAND3_X1 _u10_u5_U66  ( .A1(_u10_u5_n1964 ), .A2(_u10_u5_n1965 ), .A3(_u10_u5_n1966 ), .ZN(_u10_u5_n1943 ) );
AND4_X1 _u10_u5_U65  ( .A1(_u10_u5_n1961 ), .A2(_u10_u5_n1863 ), .A3(_u10_u5_n1962 ), .A4(_u10_u5_n1963 ), .ZN(_u10_u5_n1957 ) );
NOR2_X1 _u10_u5_U64  ( .A1(_u10_u5_n1959 ), .A2(_u10_u5_n1960 ), .ZN(_u10_u5_n1958 ) );
NOR2_X1 _u10_u5_U63  ( .A1(_u10_u5_n1957 ), .A2(_u10_u5_n1958 ), .ZN(_u10_u5_n1945 ) );
NOR2_X1 _u10_u5_U62  ( .A1(_u10_u5_n1955 ), .A2(_u10_u5_n1956 ), .ZN(_u10_u5_n1953 ) );
NOR4_X1 _u10_u5_U61  ( .A1(_u10_u5_n1952 ), .A2(_u10_u5_n1953 ), .A3(_u10_u5_n1846 ), .A4(_u10_u5_n1954 ), .ZN(_u10_u5_n1946 ) );
NOR2_X1 _u10_u5_U60  ( .A1(_u10_u5_n1950 ), .A2(_u10_u5_n1951 ), .ZN(_u10_u5_n1949 ) );
NOR2_X1 _u10_u5_U59  ( .A1(_u10_u5_n1948 ), .A2(_u10_u5_n1949 ), .ZN(_u10_u5_n1947 ) );
NOR3_X1 _u10_u5_U58  ( .A1(_u10_u5_n1945 ), .A2(_u10_u5_n1946 ), .A3(_u10_u5_n1947 ), .ZN(_u10_u5_n1944 ) );
NAND4_X1 _u10_u5_U57  ( .A1(_u10_u5_n1941 ), .A2(_u10_u5_n1942 ), .A3(_u10_u5_n1943 ), .A4(_u10_u5_n1944 ), .ZN(_u10_u5_n1824 ) );
NAND2_X1 _u10_u5_U56  ( .A1(_u10_u5_n1939 ), .A2(_u10_u5_n1940 ), .ZN(_u10_u5_n1938 ) );
NAND2_X1 _u10_u5_U55  ( .A1(_u10_u5_n1937 ), .A2(_u10_u5_n1938 ), .ZN(_u10_u5_n1903 ) );
NAND2_X1 _u10_u5_U54  ( .A1(_u10_u5_n1935 ), .A2(_u10_u5_n1936 ), .ZN(_u10_u5_n1934 ) );
NAND2_X1 _u10_u5_U53  ( .A1(_u10_u5_n1933 ), .A2(_u10_u5_n1934 ), .ZN(_u10_u5_n1931 ) );
NAND2_X1 _u10_u5_U52  ( .A1(_u10_u5_n1931 ), .A2(_u10_u5_n1932 ), .ZN(_u10_u5_n1904 ) );
NAND2_X1 _u10_u5_U51  ( .A1(_u10_u5_n1929 ), .A2(_u10_u5_n1930 ), .ZN(_u10_u5_n1927 ) );
NAND2_X1 _u10_u5_U50  ( .A1(_u10_u5_n1927 ), .A2(_u10_u5_n1928 ), .ZN(_u10_u5_n1905 ) );
NOR3_X1 _u10_u5_U49  ( .A1(_u10_u5_n1916 ), .A2(_u10_u5_n1925 ), .A3(_u10_u5_n1926 ), .ZN(_u10_u5_n1919 ) );
NOR2_X1 _u10_u5_U48  ( .A1(_u10_u5_n1923 ), .A2(_u10_u5_n1924 ), .ZN(_u10_u5_n1921 ) );
NOR2_X1 _u10_u5_U47  ( .A1(_u10_u5_n1921 ), .A2(_u10_u5_n1922 ), .ZN(_u10_u5_n1920 ) );
NOR2_X1 _u10_u5_U46  ( .A1(_u10_u5_n1919 ), .A2(_u10_u5_n1920 ), .ZN(_u10_u5_n1917 ) );
NOR2_X1 _u10_u5_U45  ( .A1(_u10_u5_n1917 ), .A2(_u10_u5_n1918 ), .ZN(_u10_u5_n1907 ) );
NOR2_X1 _u10_u5_U44  ( .A1(_u10_u5_n1915 ), .A2(_u10_u5_n1916 ), .ZN(_u10_u5_n1914 ) );
NOR2_X1 _u10_u5_U43  ( .A1(_u10_u5_n1914 ), .A2(1'b0), .ZN(_u10_u5_n1912 ));
NOR2_X1 _u10_u5_U42  ( .A1(_u10_u5_n1912 ), .A2(_u10_u5_n1913 ), .ZN(_u10_u5_n1908 ) );
NOR2_X1 _u10_u5_U41  ( .A1(_u10_u5_n1891 ), .A2(_u10_u5_n1911 ), .ZN(_u10_u5_n1910 ) );
NOR2_X1 _u10_u5_U40  ( .A1(_u10_u5_n1910 ), .A2(_u10_u5_n1868 ), .ZN(_u10_u5_n1909 ) );
NOR3_X1 _u10_u5_U39  ( .A1(_u10_u5_n1907 ), .A2(_u10_u5_n1908 ), .A3(_u10_u5_n1909 ), .ZN(_u10_u5_n1906 ) );
NAND4_X1 _u10_u5_U38  ( .A1(_u10_u5_n1903 ), .A2(_u10_u5_n1904 ), .A3(_u10_u5_n1905 ), .A4(_u10_u5_n1906 ), .ZN(_u10_u5_n1825 ) );
NAND2_X1 _u10_u5_U37  ( .A1(_u10_u5_n1901 ), .A2(_u10_u5_n1902 ), .ZN(_u10_u5_n1900 ) );
NAND2_X1 _u10_u5_U36  ( .A1(_u10_u5_n1899 ), .A2(_u10_u5_n1900 ), .ZN(_u10_u5_n1875 ) );
OR2_X1 _u10_u5_U35  ( .A1(_u10_u5_n1847 ), .A2(_u10_u5_n1898 ), .ZN(_u10_u5_n1897 ) );
NAND2_X1 _u10_u5_U34  ( .A1(_u10_u5_n1896 ), .A2(_u10_u5_n1897 ), .ZN(_u10_u5_n1895 ) );
NAND2_X1 _u10_u5_U33  ( .A1(_u10_u5_n1894 ), .A2(_u10_u5_n1895 ), .ZN(_u10_u5_n1876 ) );
NAND2_X1 _u10_u5_U32  ( .A1(_u10_u5_n1892 ), .A2(_u10_u5_n1893 ), .ZN(_u10_u5_n1877 ) );
NOR3_X1 _u10_u5_U31  ( .A1(_u10_u5_n1884 ), .A2(_u10_u5_n1890 ), .A3(_u10_u5_n1891 ), .ZN(_u10_u5_n1889 ) );
NOR2_X1 _u10_u5_U30  ( .A1(_u10_u5_n1840 ), .A2(_u10_u5_n1889 ), .ZN(_u10_u5_n1879 ) );
NOR2_X1 _u10_u5_U29  ( .A1(_u10_u5_n1887 ), .A2(_u10_u5_n1888 ), .ZN(_u10_u5_n1880 ) );
NOR3_X1 _u10_u5_U28  ( .A1(_u10_u5_n1884 ), .A2(_u10_u5_n1885 ), .A3(_u10_u5_n1886 ), .ZN(_u10_u5_n1883 ) );
NOR2_X1 _u10_u5_U27  ( .A1(_u10_u5_n1882 ), .A2(_u10_u5_n1883 ), .ZN(_u10_u5_n1881 ) );
NOR3_X1 _u10_u5_U26  ( .A1(_u10_u5_n1879 ), .A2(_u10_u5_n1880 ), .A3(_u10_u5_n1881 ), .ZN(_u10_u5_n1878 ) );
NAND4_X1 _u10_u5_U25  ( .A1(_u10_u5_n1875 ), .A2(_u10_u5_n1876 ), .A3(_u10_u5_n1877 ), .A4(_u10_u5_n1878 ), .ZN(_u10_u5_n1826 ) );
NOR3_X1 _u10_u5_U24  ( .A1(_u10_u5_n1872 ), .A2(_u10_u5_n1873 ), .A3(_u10_u5_n1874 ), .ZN(_u10_u5_n1871 ) );
NAND4_X1 _u10_u5_U23  ( .A1(_u10_u5_n1868 ), .A2(_u10_u5_n1869 ), .A3(_u10_u5_n1870 ), .A4(_u10_u5_n1871 ), .ZN(_u10_u5_n1867 ) );
NAND2_X1 _u10_u5_U22  ( .A1(_u10_u5_n1866 ), .A2(_u10_u5_n1867 ), .ZN(_u10_u5_n1865 ) );
NAND3_X1 _u10_u5_U21  ( .A1(_u10_u5_n1863 ), .A2(_u10_u5_n1864 ), .A3(_u10_u5_n1865 ), .ZN(_u10_u5_n1862 ) );
NAND2_X1 _u10_u5_U20  ( .A1(_u10_u5_n1861 ), .A2(_u10_u5_n1862 ), .ZN(_u10_u5_n1828 ) );
NAND3_X1 _u10_u5_U19  ( .A1(_u10_u5_n1858 ), .A2(_u10_u5_n1859 ), .A3(_u10_u5_n1860 ), .ZN(_u10_u5_n1857 ) );
NAND2_X1 _u10_u5_U18  ( .A1(_u10_u5_n1856 ), .A2(_u10_u5_n1857 ), .ZN(_u10_u5_n1829 ) );
OR2_X1 _u10_u5_U17  ( .A1(_u10_u5_n1854 ), .A2(_u10_u5_n1855 ), .ZN(_u10_u5_n1830 ) );
NOR2_X1 _u10_u5_U16  ( .A1(_u10_u5_n1852 ), .A2(_u10_u5_n1853 ), .ZN(_u10_u5_n1850 ) );
NOR3_X1 _u10_u5_U15  ( .A1(_u10_u5_n1850 ), .A2(_u10_u5_n1851 ), .A3(_u10_u5_n1838 ), .ZN(_u10_u5_n1848 ) );
NOR2_X1 _u10_u5_U14  ( .A1(_u10_u5_n1848 ), .A2(_u10_u5_n1849 ), .ZN(_u10_u5_n1832 ) );
NOR2_X1 _u10_u5_U13  ( .A1(_u10_u5_n1846 ), .A2(_u10_u5_n1847 ), .ZN(_u10_u5_n1845 ) );
NOR3_X1 _u10_u5_U12  ( .A1(_u10_u5_n1844 ), .A2(1'b0), .A3(_u10_u5_n1845 ),.ZN(_u10_u5_n1842 ) );
NOR2_X1 _u10_u5_U11  ( .A1(_u10_u5_n1842 ), .A2(_u10_u5_n1843 ), .ZN(_u10_u5_n1833 ) );
NOR2_X1 _u10_u5_U10  ( .A1(_u10_u5_n1840 ), .A2(_u10_u5_n1841 ), .ZN(_u10_u5_n1839 ) );
NOR3_X1 _u10_u5_U9  ( .A1(_u10_u5_n1837 ), .A2(_u10_u5_n1838 ), .A3(_u10_u5_n1839 ), .ZN(_u10_u5_n1835 ) );
NOR2_X1 _u10_u5_U8  ( .A1(_u10_u5_n1835 ), .A2(_u10_u5_n1836 ), .ZN(_u10_u5_n1834 ) );
NOR3_X1 _u10_u5_U7  ( .A1(_u10_u5_n1832 ), .A2(_u10_u5_n1833 ), .A3(_u10_u5_n1834 ), .ZN(_u10_u5_n1831 ) );
NAND4_X1 _u10_u5_U6  ( .A1(_u10_u5_n1828 ), .A2(_u10_u5_n1829 ), .A3(_u10_u5_n1830 ), .A4(_u10_u5_n1831 ), .ZN(_u10_u5_n1827 ) );
NOR4_X1 _u10_u5_U5  ( .A1(_u10_u5_n1824 ), .A2(_u10_u5_n1825 ), .A3(_u10_u5_n1826 ), .A4(_u10_u5_n1827 ), .ZN(_u10_u5_n1823 ) );
NAND4_X1 _u10_u5_U4  ( .A1(_u10_u5_n1820 ), .A2(_u10_u5_n1821 ), .A3(_u10_u5_n1822 ), .A4(_u10_u5_n1823 ), .ZN(_u10_u5_n1818 ) );
MUX2_X1 _u10_u5_U3  ( .A(_u10_u5_n1818 ), .B(_u10_SYNOPSYS_UNCONNECTED_22 ),.S(_u10_u5_n1819 ), .Z(_u10_u5_n1812 ) );
DFFR_X1 _u10_u5_state_reg_1_  ( .D(_u10_u5_n1812 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_22 ), .QN(_u10_u5_n1814 ));
DFFR_X1 _u10_u5_state_reg_2_  ( .D(_u10_u5_n1811 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_21 ), .QN(_u10_u5_n1815 ));
DFFR_X1 _u10_u5_state_reg_3_  ( .D(_u10_u5_n1810 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_20 ), .QN(_u10_u5_n1816 ));
DFFR_X1 _u10_u5_state_reg_4_  ( .D(_u10_u5_n1809 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_19 ), .QN(_u10_u5_n1817 ));
DFFR_X1 _u10_u5_state_reg_0_  ( .D(_u10_u5_n1808 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_23 ), .QN(_u10_u5_n1813 ));
NOR2_X1 _u10_u6_U1606  ( .A1(_u10_SYNOPSYS_UNCONNECTED_26 ), .A2(_u10_u6_n1814 ), .ZN(_u10_u6_n3174 ) );
NOR3_X1 _u10_u6_U1605  ( .A1(_u10_SYNOPSYS_UNCONNECTED_25 ), .A2(_u10_u6_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_28 ), .ZN(_u10_u6_n3328 ) );
NAND2_X1 _u10_u6_U1604  ( .A1(_u10_u6_n3174 ), .A2(_u10_u6_n3328 ), .ZN(_u10_u6_n1843 ) );
INV_X1 _u10_u6_U1603  ( .A(_u10_u6_n1843 ), .ZN(_u10_u6_n2461 ) );
INV_X1 _u10_u6_U1602  ( .A(1'b0), .ZN(_u10_u6_n2466 ) );
INV_X1 _u10_u6_U1601  ( .A(1'b0), .ZN(_u10_u6_n2305 ) );
NAND2_X1 _u10_u6_U1600  ( .A1(_u10_u6_n2466 ), .A2(_u10_u6_n2305 ), .ZN(_u10_u6_n1954 ) );
INV_X1 _u10_u6_U1599  ( .A(_u10_u6_n1954 ), .ZN(_u10_u6_n2467 ) );
INV_X1 _u10_u6_U1598  ( .A(1'b0), .ZN(_u10_u6_n1936 ) );
NOR2_X1 _u10_u6_U1597  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u6_n2223 ) );
INV_X1 _u10_u6_U1596  ( .A(1'b0), .ZN(_u10_u6_n1922 ) );
NAND2_X1 _u10_u6_U1595  ( .A1(_u10_u6_n2223 ), .A2(_u10_u6_n1922 ), .ZN(_u10_u6_n2200 ) );
NOR2_X1 _u10_u6_U1594  ( .A1(_u10_u6_n2200 ), .A2(1'b0), .ZN(_u10_u6_n2502 ));
INV_X1 _u10_u6_U1593  ( .A(1'b0), .ZN(_u10_u6_n2978 ) );
INV_X1 _u10_u6_U1592  ( .A(1'b0), .ZN(_u10_u6_n3000 ) );
NAND2_X1 _u10_u6_U1591  ( .A1(_u10_u6_n2978 ), .A2(_u10_u6_n3000 ), .ZN(_u10_u6_n3356 ) );
INV_X1 _u10_u6_U1590  ( .A(1'b0), .ZN(_u10_u6_n2405 ) );
INV_X1 _u10_u6_U1589  ( .A(1'b0), .ZN(_u10_u6_n2972 ) );
NAND2_X1 _u10_u6_U1588  ( .A1(_u10_u6_n2405 ), .A2(_u10_u6_n2972 ), .ZN(_u10_u6_n2008 ) );
NOR2_X1 _u10_u6_U1587  ( .A1(_u10_u6_n3356 ), .A2(_u10_u6_n2008 ), .ZN(_u10_u6_n2195 ) );
NAND2_X1 _u10_u6_U1586  ( .A1(_u10_u6_n2502 ), .A2(_u10_u6_n2195 ), .ZN(_u10_u6_n2490 ) );
INV_X1 _u10_u6_U1585  ( .A(1'b0), .ZN(_u10_u6_n3040 ) );
INV_X1 _u10_u6_U1584  ( .A(1'b0), .ZN(_u10_u6_n3006 ) );
NAND2_X1 _u10_u6_U1583  ( .A1(_u10_u6_n3040 ), .A2(_u10_u6_n3006 ), .ZN(_u10_u6_n2508 ) );
NOR2_X1 _u10_u6_U1582  ( .A1(_u10_u6_n2508 ), .A2(1'b0), .ZN(_u10_u6_n2493 ));
INV_X1 _u10_u6_U1581  ( .A(1'b0), .ZN(_u10_u6_n2038 ) );
NAND2_X1 _u10_u6_U1580  ( .A1(_u10_u6_n2493 ), .A2(_u10_u6_n2038 ), .ZN(_u10_u6_n2174 ) );
NOR2_X1 _u10_u6_U1579  ( .A1(_u10_u6_n2490 ), .A2(_u10_u6_n2174 ), .ZN(_u10_u6_n2659 ) );
INV_X1 _u10_u6_U1578  ( .A(1'b0), .ZN(_u10_u6_n2175 ) );
NAND3_X1 _u10_u6_U1577  ( .A1(_u10_u6_n2659 ), .A2(_u10_u6_n2175 ), .A3(1'b0), .ZN(_u10_u6_n3189 ) );
NOR2_X1 _u10_u6_U1576  ( .A1(_u10_u6_n3189 ), .A2(1'b0), .ZN(_u10_u6_n2528 ));
INV_X1 _u10_u6_U1575  ( .A(1'b0), .ZN(_u10_u6_n2837 ) );
NAND2_X1 _u10_u6_U1574  ( .A1(_u10_u6_n2528 ), .A2(_u10_u6_n2837 ), .ZN(_u10_u6_n2567 ) );
INV_X1 _u10_u6_U1573  ( .A(1'b0), .ZN(_u10_u6_n2080 ) );
INV_X1 _u10_u6_U1572  ( .A(1'b0), .ZN(_u10_u6_n2166 ) );
NAND2_X1 _u10_u6_U1571  ( .A1(_u10_u6_n2080 ), .A2(_u10_u6_n2166 ), .ZN(_u10_u6_n2840 ) );
NOR2_X1 _u10_u6_U1570  ( .A1(_u10_u6_n2567 ), .A2(_u10_u6_n2840 ), .ZN(_u10_u6_n2443 ) );
INV_X1 _u10_u6_U1569  ( .A(1'b0), .ZN(_u10_u6_n2600 ) );
INV_X1 _u10_u6_U1568  ( .A(1'b0), .ZN(_u10_u6_n2836 ) );
NAND2_X1 _u10_u6_U1567  ( .A1(_u10_u6_n2600 ), .A2(_u10_u6_n2836 ), .ZN(_u10_u6_n2428 ) );
INV_X1 _u10_u6_U1566  ( .A(_u10_u6_n2428 ), .ZN(_u10_u6_n2078 ) );
NAND2_X1 _u10_u6_U1565  ( .A1(_u10_u6_n2443 ), .A2(_u10_u6_n2078 ), .ZN(_u10_u6_n2282 ) );
INV_X1 _u10_u6_U1564  ( .A(1'b0), .ZN(_u10_u6_n2874 ) );
INV_X1 _u10_u6_U1563  ( .A(1'b0), .ZN(_u10_u6_n2031 ) );
NAND2_X1 _u10_u6_U1562  ( .A1(_u10_u6_n2874 ), .A2(_u10_u6_n2031 ), .ZN(_u10_u6_n1976 ) );
NOR2_X1 _u10_u6_U1561  ( .A1(_u10_u6_n2282 ), .A2(_u10_u6_n1976 ), .ZN(_u10_u6_n2411 ) );
NAND3_X1 _u10_u6_U1560  ( .A1(_u10_u6_n2467 ), .A2(_u10_u6_n1936 ), .A3(_u10_u6_n2411 ), .ZN(_u10_u6_n2464 ) );
NAND3_X1 _u10_u6_U1559  ( .A1(_u10_u6_n2166 ), .A2(_u10_u6_n2837 ), .A3(1'b0), .ZN(_u10_u6_n3276 ) );
INV_X1 _u10_u6_U1558  ( .A(_u10_u6_n3276 ), .ZN(_u10_u6_n2442 ) );
NAND3_X1 _u10_u6_U1557  ( .A1(_u10_u6_n2836 ), .A2(_u10_u6_n2080 ), .A3(_u10_u6_n2442 ), .ZN(_u10_u6_n2838 ) );
INV_X1 _u10_u6_U1556  ( .A(_u10_u6_n2838 ), .ZN(_u10_u6_n2850 ) );
NOR2_X1 _u10_u6_U1555  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u6_n2953 ) );
NAND2_X1 _u10_u6_U1554  ( .A1(_u10_u6_n2850 ), .A2(_u10_u6_n2953 ), .ZN(_u10_u6_n2947 ) );
INV_X1 _u10_u6_U1553  ( .A(_u10_u6_n2947 ), .ZN(_u10_u6_n2420 ) );
NAND2_X1 _u10_u6_U1552  ( .A1(_u10_u6_n1936 ), .A2(_u10_u6_n2874 ), .ZN(_u10_u6_n2030 ) );
INV_X1 _u10_u6_U1551  ( .A(_u10_u6_n2030 ), .ZN(_u10_u6_n2162 ) );
NAND2_X1 _u10_u6_U1550  ( .A1(_u10_u6_n2420 ), .A2(_u10_u6_n2162 ), .ZN(_u10_u6_n2828 ) );
INV_X1 _u10_u6_U1549  ( .A(_u10_u6_n2828 ), .ZN(_u10_u6_n2551 ) );
NAND2_X1 _u10_u6_U1548  ( .A1(_u10_u6_n2551 ), .A2(_u10_u6_n2467 ), .ZN(_u10_u6_n3416 ) );
NAND2_X1 _u10_u6_U1547  ( .A1(_u10_u6_n2464 ), .A2(_u10_u6_n3416 ), .ZN(_u10_u6_n2266 ) );
INV_X1 _u10_u6_U1546  ( .A(_u10_u6_n2266 ), .ZN(_u10_u6_n3410 ) );
NAND2_X1 _u10_u6_U1545  ( .A1(1'b0), .A2(_u10_u6_n2305 ), .ZN(_u10_u6_n3411 ) );
INV_X1 _u10_u6_U1544  ( .A(_u10_u6_n3356 ), .ZN(_u10_u6_n1983 ) );
NAND3_X1 _u10_u6_U1543  ( .A1(_u10_u6_n1983 ), .A2(_u10_u6_n2405 ), .A3(1'b0), .ZN(_u10_u6_n2022 ) );
INV_X1 _u10_u6_U1542  ( .A(_u10_u6_n2022 ), .ZN(_u10_u6_n2056 ) );
INV_X1 _u10_u6_U1541  ( .A(_u10_u6_n2840 ), .ZN(_u10_u6_n2059 ) );
INV_X1 _u10_u6_U1540  ( .A(1'b0), .ZN(_u10_u6_n1965 ) );
NAND2_X1 _u10_u6_U1539  ( .A1(_u10_u6_n2837 ), .A2(_u10_u6_n1965 ), .ZN(_u10_u6_n1852 ) );
INV_X1 _u10_u6_U1538  ( .A(_u10_u6_n1852 ), .ZN(_u10_u6_n3190 ) );
INV_X1 _u10_u6_U1537  ( .A(1'b0), .ZN(_u10_u6_n1853 ) );
NAND2_X1 _u10_u6_U1536  ( .A1(_u10_u6_n3190 ), .A2(_u10_u6_n1853 ), .ZN(_u10_u6_n2687 ) );
INV_X1 _u10_u6_U1535  ( .A(_u10_u6_n2687 ), .ZN(_u10_u6_n2019 ) );
NAND2_X1 _u10_u6_U1534  ( .A1(_u10_u6_n2059 ), .A2(_u10_u6_n2019 ), .ZN(_u10_u6_n2330 ) );
NOR2_X1 _u10_u6_U1533  ( .A1(_u10_u6_n2428 ), .A2(_u10_u6_n2330 ), .ZN(_u10_u6_n2036 ) );
NAND2_X1 _u10_u6_U1532  ( .A1(_u10_u6_n2056 ), .A2(_u10_u6_n2036 ), .ZN(_u10_u6_n3379 ) );
NOR2_X1 _u10_u6_U1531  ( .A1(_u10_u6_n3379 ), .A2(_u10_u6_n2030 ), .ZN(_u10_u6_n2026 ) );
INV_X1 _u10_u6_U1530  ( .A(1'b0), .ZN(_u10_u6_n2431 ) );
NOR2_X1 _u10_u6_U1529  ( .A1(_u10_u6_n2431 ), .A2(1'b0), .ZN(_u10_u6_n3062 ));
NAND2_X1 _u10_u6_U1528  ( .A1(_u10_u6_n3062 ), .A2(_u10_u6_n2195 ), .ZN(_u10_u6_n3407 ) );
NOR3_X1 _u10_u6_U1527  ( .A1(_u10_u6_n2687 ), .A2(1'b0), .A3(_u10_u6_n3407 ),.ZN(_u10_u6_n3275 ) );
NAND3_X1 _u10_u6_U1526  ( .A1(_u10_u6_n2836 ), .A2(_u10_u6_n2080 ), .A3(_u10_u6_n3275 ), .ZN(_u10_u6_n3297 ) );
INV_X1 _u10_u6_U1525  ( .A(_u10_u6_n3297 ), .ZN(_u10_u6_n3172 ) );
NAND2_X1 _u10_u6_U1524  ( .A1(_u10_u6_n3172 ), .A2(_u10_u6_n2600 ), .ZN(_u10_u6_n2226 ) );
NOR2_X1 _u10_u6_U1523  ( .A1(_u10_u6_n2226 ), .A2(1'b0), .ZN(_u10_u6_n2307 ));
INV_X1 _u10_u6_U1522  ( .A(_u10_u6_n2490 ), .ZN(_u10_u6_n2536 ) );
NAND3_X1 _u10_u6_U1521  ( .A1(_u10_u6_n2536 ), .A2(_u10_u6_n3040 ), .A3(1'b0), .ZN(_u10_u6_n3226 ) );
NOR2_X1 _u10_u6_U1520  ( .A1(_u10_u6_n3226 ), .A2(_u10_u6_n2330 ), .ZN(_u10_u6_n2441 ) );
NAND2_X1 _u10_u6_U1519  ( .A1(_u10_u6_n2441 ), .A2(_u10_u6_n2953 ), .ZN(_u10_u6_n2579 ) );
NOR2_X1 _u10_u6_U1518  ( .A1(_u10_u6_n2579 ), .A2(_u10_u6_n2030 ), .ZN(_u10_u6_n2550 ) );
NOR3_X1 _u10_u6_U1517  ( .A1(_u10_u6_n2026 ), .A2(_u10_u6_n2307 ), .A3(_u10_u6_n2550 ), .ZN(_u10_u6_n3394 ) );
NAND2_X1 _u10_u6_U1516  ( .A1(1'b0), .A2(_u10_u6_n2978 ), .ZN(_u10_u6_n3115 ) );
NOR2_X1 _u10_u6_U1515  ( .A1(_u10_u6_n3115 ), .A2(_u10_u6_n2330 ), .ZN(_u10_u6_n3126 ) );
NAND2_X1 _u10_u6_U1514  ( .A1(_u10_u6_n2162 ), .A2(_u10_u6_n2031 ), .ZN(_u10_u6_n2686 ) );
NOR2_X1 _u10_u6_U1513  ( .A1(_u10_u6_n2686 ), .A2(_u10_u6_n2428 ), .ZN(_u10_u6_n2108 ) );
NAND2_X1 _u10_u6_U1512  ( .A1(_u10_u6_n3126 ), .A2(_u10_u6_n2108 ), .ZN(_u10_u6_n3415 ) );
NAND2_X1 _u10_u6_U1511  ( .A1(_u10_u6_n3394 ), .A2(_u10_u6_n3415 ), .ZN(_u10_u6_n3089 ) );
NAND2_X1 _u10_u6_U1510  ( .A1(_u10_u6_n3089 ), .A2(_u10_u6_n2305 ), .ZN(_u10_u6_n3414 ) );
NAND2_X1 _u10_u6_U1509  ( .A1(_u10_u6_n2466 ), .A2(_u10_u6_n3414 ), .ZN(_u10_u6_n3118 ) );
NAND2_X1 _u10_u6_U1508  ( .A1(_u10_u6_n2078 ), .A2(_u10_u6_n2080 ), .ZN(_u10_u6_n2596 ) );
NAND2_X1 _u10_u6_U1507  ( .A1(1'b0), .A2(_u10_u6_n2493 ), .ZN(_u10_u6_n1961 ) );
NOR3_X1 _u10_u6_U1506  ( .A1(_u10_u6_n2490 ), .A2(1'b0), .A3(_u10_u6_n1961 ),.ZN(_u10_u6_n2054 ) );
NAND2_X1 _u10_u6_U1505  ( .A1(_u10_u6_n2054 ), .A2(_u10_u6_n3190 ), .ZN(_u10_u6_n2061 ) );
OR2_X1 _u10_u6_U1504  ( .A1(_u10_u6_n2596 ), .A2(_u10_u6_n2061 ), .ZN(_u10_u6_n1969 ) );
NOR3_X1 _u10_u6_U1503  ( .A1(_u10_u6_n1976 ), .A2(1'b0), .A3(_u10_u6_n1969 ),.ZN(_u10_u6_n2710 ) );
NAND2_X1 _u10_u6_U1502  ( .A1(_u10_u6_n2710 ), .A2(_u10_u6_n2467 ), .ZN(_u10_u6_n2545 ) );
INV_X1 _u10_u6_U1501  ( .A(_u10_u6_n2545 ), .ZN(_u10_u6_n2087 ) );
NOR2_X1 _u10_u6_U1500  ( .A1(_u10_u6_n3118 ), .A2(_u10_u6_n2087 ), .ZN(_u10_u6_n3145 ) );
NOR2_X1 _u10_u6_U1499  ( .A1(_u10_u6_n2030 ), .A2(1'b0), .ZN(_u10_u6_n2668 ));
NAND2_X1 _u10_u6_U1498  ( .A1(1'b0), .A2(_u10_u6_n2668 ), .ZN(_u10_u6_n2163 ) );
INV_X1 _u10_u6_U1497  ( .A(_u10_u6_n2163 ), .ZN(_u10_u6_n2875 ) );
INV_X1 _u10_u6_U1496  ( .A(_u10_u6_n1976 ), .ZN(_u10_u6_n2747 ) );
NAND3_X1 _u10_u6_U1495  ( .A1(_u10_u6_n2747 ), .A2(_u10_u6_n2600 ), .A3(1'b0), .ZN(_u10_u6_n3393 ) );
NOR3_X1 _u10_u6_U1494  ( .A1(1'b0), .A2(1'b0), .A3(_u10_u6_n3393 ), .ZN(_u10_u6_n3180 ) );
INV_X1 _u10_u6_U1493  ( .A(1'b0), .ZN(_u10_u6_n2113 ) );
INV_X1 _u10_u6_U1492  ( .A(1'b0), .ZN(_u10_u6_n3066 ) );
NAND2_X1 _u10_u6_U1491  ( .A1(_u10_u6_n2175 ), .A2(_u10_u6_n3066 ), .ZN(_u10_u6_n2216 ) );
INV_X1 _u10_u6_U1490  ( .A(_u10_u6_n2659 ), .ZN(_u10_u6_n2643 ) );
NOR2_X1 _u10_u6_U1489  ( .A1(_u10_u6_n2216 ), .A2(_u10_u6_n2643 ), .ZN(_u10_u6_n2049 ) );
AND2_X1 _u10_u6_U1488  ( .A1(_u10_u6_n2049 ), .A2(_u10_u6_n1853 ), .ZN(_u10_u6_n3223 ) );
NAND2_X1 _u10_u6_U1487  ( .A1(_u10_u6_n3223 ), .A2(_u10_u6_n1965 ), .ZN(_u10_u6_n2531 ) );
NOR2_X1 _u10_u6_U1486  ( .A1(_u10_u6_n2531 ), .A2(1'b0), .ZN(_u10_u6_n2884 ));
NAND2_X1 _u10_u6_U1485  ( .A1(_u10_u6_n2884 ), .A2(_u10_u6_n2166 ), .ZN(_u10_u6_n1841 ) );
NOR2_X1 _u10_u6_U1484  ( .A1(_u10_u6_n1841 ), .A2(1'b0), .ZN(_u10_u6_n3129 ));
NAND2_X1 _u10_u6_U1483  ( .A1(_u10_u6_n3129 ), .A2(_u10_u6_n2836 ), .ZN(_u10_u6_n2842 ) );
INV_X1 _u10_u6_U1482  ( .A(_u10_u6_n2842 ), .ZN(_u10_u6_n2833 ) );
NAND2_X1 _u10_u6_U1481  ( .A1(_u10_u6_n2833 ), .A2(_u10_u6_n2600 ), .ZN(_u10_u6_n2853 ) );
INV_X1 _u10_u6_U1480  ( .A(_u10_u6_n2853 ), .ZN(_u10_u6_n2082 ) );
NAND2_X1 _u10_u6_U1479  ( .A1(_u10_u6_n2082 ), .A2(_u10_u6_n2031 ), .ZN(_u10_u6_n2274 ) );
INV_X1 _u10_u6_U1478  ( .A(_u10_u6_n2274 ), .ZN(_u10_u6_n2669 ) );
NAND3_X1 _u10_u6_U1477  ( .A1(_u10_u6_n2668 ), .A2(_u10_u6_n2113 ), .A3(_u10_u6_n2669 ), .ZN(_u10_u6_n1858 ) );
INV_X1 _u10_u6_U1476  ( .A(_u10_u6_n1858 ), .ZN(_u10_u6_n3067 ) );
NAND2_X1 _u10_u6_U1475  ( .A1(_u10_u6_n3067 ), .A2(1'b0), .ZN(_u10_u6_n2092 ) );
INV_X1 _u10_u6_U1474  ( .A(_u10_u6_n2092 ), .ZN(_u10_u6_n3294 ) );
INV_X1 _u10_u6_U1473  ( .A(1'b0), .ZN(_u10_u6_n2446 ) );
INV_X1 _u10_u6_U1472  ( .A(1'b0), .ZN(_u10_u6_n2996 ) );
NAND2_X1 _u10_u6_U1471  ( .A1(_u10_u6_n3067 ), .A2(_u10_u6_n2996 ), .ZN(_u10_u6_n1847 ) );
NOR3_X1 _u10_u6_U1470  ( .A1(_u10_u6_n2446 ), .A2(1'b0), .A3(_u10_u6_n1847 ),.ZN(_u10_u6_n3413 ) );
NOR4_X1 _u10_u6_U1469  ( .A1(_u10_u6_n2875 ), .A2(_u10_u6_n3180 ), .A3(_u10_u6_n3294 ), .A4(_u10_u6_n3413 ), .ZN(_u10_u6_n3412 ) );
NAND4_X1 _u10_u6_U1468  ( .A1(_u10_u6_n3410 ), .A2(_u10_u6_n3411 ), .A3(_u10_u6_n3145 ), .A4(_u10_u6_n3412 ), .ZN(_u10_u6_n3409 ) );
NAND2_X1 _u10_u6_U1467  ( .A1(_u10_u6_n2461 ), .A2(_u10_u6_n3409 ), .ZN(_u10_u6_n3380 ) );
NOR2_X1 _u10_u6_U1466  ( .A1(_u10_u6_n1817 ), .A2(_u10_u6_n1816 ), .ZN(_u10_u6_n3368 ) );
AND2_X1 _u10_u6_U1465  ( .A1(_u10_u6_n3368 ), .A2(_u10_u6_n1813 ), .ZN(_u10_u6_n3320 ) );
NOR2_X1 _u10_u6_U1464  ( .A1(_u10_SYNOPSYS_UNCONNECTED_27 ), .A2(_u10_u6_n1815 ), .ZN(_u10_u6_n3236 ) );
NAND2_X1 _u10_u6_U1463  ( .A1(_u10_u6_n3320 ), .A2(_u10_u6_n3236 ), .ZN(_u10_u6_n2607 ) );
INV_X1 _u10_u6_U1462  ( .A(_u10_u6_n2607 ), .ZN(_u10_u6_n1966 ) );
INV_X1 _u10_u6_U1461  ( .A(_u10_u6_n2200 ), .ZN(_u10_u6_n3216 ) );
NAND2_X1 _u10_u6_U1460  ( .A1(1'b0), .A2(_u10_u6_n3216 ), .ZN(_u10_u6_n2367 ) );
INV_X1 _u10_u6_U1459  ( .A(_u10_u6_n2367 ), .ZN(_u10_u6_n3183 ) );
NAND2_X1 _u10_u6_U1458  ( .A1(_u10_u6_n3183 ), .A2(_u10_u6_n2195 ), .ZN(_u10_u6_n2194 ) );
INV_X1 _u10_u6_U1457  ( .A(_u10_u6_n2194 ), .ZN(_u10_u6_n2055 ) );
NAND2_X1 _u10_u6_U1456  ( .A1(_u10_u6_n2055 ), .A2(_u10_u6_n1853 ), .ZN(_u10_u6_n3401 ) );
INV_X1 _u10_u6_U1455  ( .A(_u10_u6_n2531 ), .ZN(_u10_u6_n2190 ) );
INV_X1 _u10_u6_U1454  ( .A(1'b0), .ZN(_u10_u6_n3001 ) );
NAND2_X1 _u10_u6_U1453  ( .A1(_u10_u6_n3001 ), .A2(_u10_u6_n2466 ), .ZN(_u10_u6_n2156 ) );
NOR2_X1 _u10_u6_U1452  ( .A1(_u10_u6_n2166 ), .A2(_u10_u6_n2596 ), .ZN(_u10_u6_n2594 ) );
NAND2_X1 _u10_u6_U1451  ( .A1(_u10_u6_n2594 ), .A2(_u10_u6_n2031 ), .ZN(_u10_u6_n2752 ) );
INV_X1 _u10_u6_U1450  ( .A(_u10_u6_n2752 ), .ZN(_u10_u6_n2421 ) );
NAND2_X1 _u10_u6_U1449  ( .A1(_u10_u6_n2421 ), .A2(_u10_u6_n2874 ), .ZN(_u10_u6_n2033 ) );
INV_X1 _u10_u6_U1448  ( .A(_u10_u6_n2033 ), .ZN(_u10_u6_n2742 ) );
NAND3_X1 _u10_u6_U1447  ( .A1(_u10_u6_n2305 ), .A2(_u10_u6_n1936 ), .A3(_u10_u6_n2742 ), .ZN(_u10_u6_n1896 ) );
OR3_X1 _u10_u6_U1446  ( .A1(_u10_u6_n2156 ), .A2(1'b0), .A3(_u10_u6_n1896 ),.ZN(_u10_u6_n2905 ) );
NAND2_X1 _u10_u6_U1445  ( .A1(_u10_u6_n2113 ), .A2(_u10_u6_n2996 ), .ZN(_u10_u6_n2719 ) );
NOR2_X1 _u10_u6_U1444  ( .A1(_u10_u6_n2719 ), .A2(1'b0), .ZN(_u10_u6_n2941 ));
INV_X1 _u10_u6_U1443  ( .A(_u10_u6_n2941 ), .ZN(_u10_u6_n2911 ) );
NOR2_X1 _u10_u6_U1442  ( .A1(_u10_u6_n2905 ), .A2(_u10_u6_n2911 ), .ZN(_u10_u6_n3222 ) );
INV_X1 _u10_u6_U1441  ( .A(_u10_u6_n3222 ), .ZN(_u10_u6_n2695 ) );
INV_X1 _u10_u6_U1440  ( .A(_u10_u6_n2156 ), .ZN(_u10_u6_n2089 ) );
NAND3_X1 _u10_u6_U1439  ( .A1(_u10_u6_n2089 ), .A2(_u10_u6_n2446 ), .A3(_u10_u6_n3180 ), .ZN(_u10_u6_n2902 ) );
NOR2_X1 _u10_u6_U1438  ( .A1(_u10_u6_n2902 ), .A2(_u10_u6_n2911 ), .ZN(_u10_u6_n2533 ) );
INV_X1 _u10_u6_U1437  ( .A(_u10_u6_n2533 ), .ZN(_u10_u6_n2485 ) );
NAND2_X1 _u10_u6_U1436  ( .A1(_u10_u6_n2695 ), .A2(_u10_u6_n2485 ), .ZN(_u10_u6_n2721 ) );
NAND2_X1 _u10_u6_U1435  ( .A1(1'b0), .A2(_u10_u6_n2113 ), .ZN(_u10_u6_n1868 ) );
INV_X1 _u10_u6_U1434  ( .A(_u10_u6_n1868 ), .ZN(_u10_u6_n2534 ) );
NOR2_X1 _u10_u6_U1433  ( .A1(_u10_u6_n2721 ), .A2(_u10_u6_n2534 ), .ZN(_u10_u6_n3231 ) );
NAND2_X1 _u10_u6_U1432  ( .A1(_u10_u6_n2467 ), .A2(_u10_u6_n3001 ), .ZN(_u10_u6_n2303 ) );
INV_X1 _u10_u6_U1431  ( .A(_u10_u6_n2303 ), .ZN(_u10_u6_n2549 ) );
INV_X1 _u10_u6_U1430  ( .A(1'b0), .ZN(_u10_u6_n2803 ) );
NAND2_X1 _u10_u6_U1429  ( .A1(_u10_u6_n2803 ), .A2(_u10_u6_n2446 ), .ZN(_u10_u6_n1846 ) );
INV_X1 _u10_u6_U1428  ( .A(_u10_u6_n1846 ), .ZN(_u10_u6_n2667 ) );
NAND3_X1 _u10_u6_U1427  ( .A1(_u10_u6_n2549 ), .A2(_u10_u6_n2667 ), .A3(1'b0), .ZN(_u10_u6_n2739 ) );
INV_X1 _u10_u6_U1426  ( .A(_u10_u6_n2739 ), .ZN(_u10_u6_n3272 ) );
INV_X1 _u10_u6_U1425  ( .A(_u10_u6_n2719 ), .ZN(_u10_u6_n2364 ) );
NAND2_X1 _u10_u6_U1424  ( .A1(_u10_u6_n3272 ), .A2(_u10_u6_n2364 ), .ZN(_u10_u6_n2852 ) );
INV_X1 _u10_u6_U1423  ( .A(_u10_u6_n2852 ), .ZN(_u10_u6_n2214 ) );
NAND2_X1 _u10_u6_U1422  ( .A1(_u10_u6_n2875 ), .A2(_u10_u6_n2089 ), .ZN(_u10_u6_n2097 ) );
INV_X1 _u10_u6_U1421  ( .A(_u10_u6_n2097 ), .ZN(_u10_u6_n2300 ) );
NAND2_X1 _u10_u6_U1420  ( .A1(_u10_u6_n2300 ), .A2(_u10_u6_n2446 ), .ZN(_u10_u6_n2001 ) );
NOR2_X1 _u10_u6_U1419  ( .A1(_u10_u6_n2001 ), .A2(_u10_u6_n2911 ), .ZN(_u10_u6_n2877 ) );
NOR2_X1 _u10_u6_U1418  ( .A1(_u10_u6_n2214 ), .A2(_u10_u6_n2877 ), .ZN(_u10_u6_n2940 ) );
NAND2_X1 _u10_u6_U1417  ( .A1(_u10_u6_n3231 ), .A2(_u10_u6_n2940 ), .ZN(_u10_u6_n3408 ) );
NAND2_X1 _u10_u6_U1416  ( .A1(_u10_u6_n2190 ), .A2(_u10_u6_n3408 ), .ZN(_u10_u6_n3402 ) );
NOR2_X1 _u10_u6_U1415  ( .A1(_u10_u6_n2446 ), .A2(_u10_u6_n2911 ), .ZN(_u10_u6_n3059 ) );
NAND2_X1 _u10_u6_U1414  ( .A1(_u10_u6_n3059 ), .A2(_u10_u6_n2190 ), .ZN(_u10_u6_n3404 ) );
AND3_X1 _u10_u6_U1413  ( .A1(_u10_u6_n3407 ), .A2(_u10_u6_n3226 ), .A3(_u10_u6_n3115 ), .ZN(_u10_u6_n3058 ) );
NAND2_X1 _u10_u6_U1412  ( .A1(_u10_u6_n3058 ), .A2(_u10_u6_n2022 ), .ZN(_u10_u6_n3406 ) );
NAND2_X1 _u10_u6_U1411  ( .A1(_u10_u6_n1853 ), .A2(_u10_u6_n3406 ), .ZN(_u10_u6_n3405 ) );
AND3_X1 _u10_u6_U1410  ( .A1(_u10_u6_n3404 ), .A2(_u10_u6_n1965 ), .A3(_u10_u6_n3405 ), .ZN(_u10_u6_n3063 ) );
NAND2_X1 _u10_u6_U1409  ( .A1(_u10_u6_n2667 ), .A2(_u10_u6_n3001 ), .ZN(_u10_u6_n1898 ) );
INV_X1 _u10_u6_U1408  ( .A(_u10_u6_n1898 ), .ZN(_u10_u6_n2835 ) );
NAND3_X1 _u10_u6_U1407  ( .A1(_u10_u6_n2364 ), .A2(_u10_u6_n2835 ), .A3(1'b0), .ZN(_u10_u6_n1869 ) );
NOR2_X1 _u10_u6_U1406  ( .A1(_u10_u6_n1869 ), .A2(_u10_u6_n2531 ), .ZN(_u10_u6_n2761 ) );
NOR3_X1 _u10_u6_U1405  ( .A1(_u10_u6_n2761 ), .A2(_u10_u6_n2528 ), .A3(_u10_u6_n2054 ), .ZN(_u10_u6_n3403 ) );
NAND4_X1 _u10_u6_U1404  ( .A1(_u10_u6_n3401 ), .A2(_u10_u6_n3402 ), .A3(_u10_u6_n3063 ), .A4(_u10_u6_n3403 ), .ZN(_u10_u6_n3400 ) );
NAND2_X1 _u10_u6_U1403  ( .A1(_u10_u6_n1966 ), .A2(_u10_u6_n3400 ), .ZN(_u10_u6_n3381 ) );
AND2_X1 _u10_u6_U1402  ( .A1(_u10_u6_n3368 ), .A2(_u10_SYNOPSYS_UNCONNECTED_28 ), .ZN(_u10_u6_n3319 ) );
NAND2_X1 _u10_u6_U1401  ( .A1(_u10_u6_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_27 ), .ZN(_u10_u6_n1849 ) );
INV_X1 _u10_u6_U1400  ( .A(_u10_u6_n1849 ), .ZN(_u10_u6_n2183 ) );
NAND2_X1 _u10_u6_U1399  ( .A1(_u10_u6_n2884 ), .A2(_u10_u6_n2183 ), .ZN(_u10_u6_n2883 ) );
INV_X1 _u10_u6_U1398  ( .A(_u10_u6_n2883 ), .ZN(_u10_u6_n1890 ) );
INV_X1 _u10_u6_U1397  ( .A(_u10_u6_n2940 ), .ZN(_u10_u6_n3278 ) );
NAND2_X1 _u10_u6_U1396  ( .A1(_u10_u6_n1890 ), .A2(_u10_u6_n3278 ), .ZN(_u10_u6_n3382 ) );
NAND2_X1 _u10_u6_U1395  ( .A1(_u10_u6_n3059 ), .A2(_u10_u6_n2669 ), .ZN(_u10_u6_n3399 ) );
NAND2_X1 _u10_u6_U1394  ( .A1(_u10_u6_n2031 ), .A2(_u10_u6_n3399 ), .ZN(_u10_u6_n3398 ) );
NAND2_X1 _u10_u6_U1393  ( .A1(_u10_u6_n2162 ), .A2(_u10_u6_n3398 ), .ZN(_u10_u6_n3395 ) );
NAND3_X1 _u10_u6_U1392  ( .A1(_u10_u6_n2747 ), .A2(_u10_u6_n2078 ), .A3(_u10_u6_n3126 ), .ZN(_u10_u6_n3396 ) );
NAND2_X1 _u10_u6_U1391  ( .A1(_u10_u6_n2055 ), .A2(_u10_u6_n2036 ), .ZN(_u10_u6_n2285 ) );
NOR2_X1 _u10_u6_U1390  ( .A1(_u10_u6_n2285 ), .A2(_u10_u6_n2030 ), .ZN(_u10_u6_n3349 ) );
INV_X1 _u10_u6_U1389  ( .A(_u10_u6_n3349 ), .ZN(_u10_u6_n1933 ) );
INV_X1 _u10_u6_U1388  ( .A(_u10_u6_n2710 ), .ZN(_u10_u6_n3397 ) );
NAND4_X1 _u10_u6_U1387  ( .A1(_u10_u6_n3395 ), .A2(_u10_u6_n3396 ), .A3(_u10_u6_n1933 ), .A4(_u10_u6_n3397 ), .ZN(_u10_u6_n3389 ) );
NAND2_X1 _u10_u6_U1386  ( .A1(_u10_u6_n1936 ), .A2(_u10_u6_n2828 ), .ZN(_u10_u6_n3141 ) );
INV_X1 _u10_u6_U1385  ( .A(_u10_u6_n3141 ), .ZN(_u10_u6_n2302 ) );
NAND2_X1 _u10_u6_U1384  ( .A1(_u10_u6_n3394 ), .A2(_u10_u6_n2302 ), .ZN(_u10_u6_n3390 ) );
NOR2_X1 _u10_u6_U1383  ( .A1(_u10_u6_n1869 ), .A2(_u10_u6_n2274 ), .ZN(_u10_u6_n3378 ) );
INV_X1 _u10_u6_U1382  ( .A(_u10_u6_n3378 ), .ZN(_u10_u6_n2748 ) );
NOR2_X1 _u10_u6_U1381  ( .A1(1'b0), .A2(_u10_u6_n2748 ), .ZN(_u10_u6_n3391 ));
NAND2_X1 _u10_u6_U1380  ( .A1(_u10_u6_n2534 ), .A2(_u10_u6_n2669 ), .ZN(_u10_u6_n2383 ) );
INV_X1 _u10_u6_U1379  ( .A(_u10_u6_n2383 ), .ZN(_u10_u6_n1978 ) );
NAND2_X1 _u10_u6_U1378  ( .A1(_u10_u6_n1978 ), .A2(_u10_u6_n2874 ), .ZN(_u10_u6_n3392 ) );
INV_X1 _u10_u6_U1377  ( .A(_u10_u6_n2411 ), .ZN(_u10_u6_n2164 ) );
NAND4_X1 _u10_u6_U1376  ( .A1(_u10_u6_n3392 ), .A2(_u10_u6_n3393 ), .A3(_u10_u6_n2033 ), .A4(_u10_u6_n2164 ), .ZN(_u10_u6_n2476 ) );
NOR4_X1 _u10_u6_U1375  ( .A1(_u10_u6_n3389 ), .A2(_u10_u6_n3390 ), .A3(_u10_u6_n3391 ), .A4(_u10_u6_n2476 ), .ZN(_u10_u6_n3388 ) );
NAND2_X1 _u10_u6_U1374  ( .A1(_u10_u6_n3236 ), .A2(_u10_u6_n3328 ), .ZN(_u10_u6_n2025 ) );
NOR2_X1 _u10_u6_U1373  ( .A1(_u10_u6_n3388 ), .A2(_u10_u6_n2025 ), .ZN(_u10_u6_n3384 ) );
NOR2_X1 _u10_u6_U1372  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u6_n2152 ) );
NAND2_X1 _u10_u6_U1371  ( .A1(_u10_u6_n2152 ), .A2(_u10_u6_n2175 ), .ZN(_u10_u6_n2722 ) );
INV_X1 _u10_u6_U1370  ( .A(_u10_u6_n2722 ), .ZN(_u10_u6_n2588 ) );
NAND2_X1 _u10_u6_U1369  ( .A1(_u10_u6_n2549 ), .A2(_u10_u6_n3349 ), .ZN(_u10_u6_n2091 ) );
NOR2_X1 _u10_u6_U1368  ( .A1(_u10_u6_n2091 ), .A2(_u10_u6_n1846 ), .ZN(_u10_u6_n2128 ) );
NAND3_X1 _u10_u6_U1367  ( .A1(_u10_u6_n3066 ), .A2(_u10_u6_n2113 ), .A3(_u10_u6_n2128 ), .ZN(_u10_u6_n2342 ) );
INV_X1 _u10_u6_U1366  ( .A(_u10_u6_n2342 ), .ZN(_u10_u6_n3316 ) );
NAND2_X1 _u10_u6_U1365  ( .A1(_u10_u6_n2588 ), .A2(_u10_u6_n3316 ), .ZN(_u10_u6_n2142 ) );
NOR2_X1 _u10_u6_U1364  ( .A1(_u10_u6_n1954 ), .A2(_u10_u6_n1898 ), .ZN(_u10_u6_n2255 ) );
NAND2_X1 _u10_u6_U1363  ( .A1(_u10_u6_n2255 ), .A2(_u10_u6_n2996 ), .ZN(_u10_u6_n1915 ) );
INV_X1 _u10_u6_U1362  ( .A(_u10_u6_n1915 ), .ZN(_u10_u6_n2251 ) );
NAND2_X1 _u10_u6_U1361  ( .A1(_u10_u6_n2251 ), .A2(_u10_u6_n2113 ), .ZN(_u10_u6_n1925 ) );
INV_X1 _u10_u6_U1360  ( .A(_u10_u6_n2026 ), .ZN(_u10_u6_n3340 ) );
NOR3_X1 _u10_u6_U1359  ( .A1(_u10_u6_n1925 ), .A2(_u10_u6_n2216 ), .A3(_u10_u6_n3340 ), .ZN(_u10_u6_n2003 ) );
INV_X1 _u10_u6_U1358  ( .A(1'b0), .ZN(_u10_u6_n1930 ) );
NAND2_X1 _u10_u6_U1357  ( .A1(_u10_u6_n2003 ), .A2(_u10_u6_n1930 ), .ZN(_u10_u6_n3387 ) );
AND2_X1 _u10_u6_U1356  ( .A1(_u10_u6_n2142 ), .A2(_u10_u6_n3387 ), .ZN(_u10_u6_n3366 ) );
NOR3_X1 _u10_u6_U1355  ( .A1(_u10_u6_n1813 ), .A2(_u10_u6_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_24 ), .ZN(_u10_u6_n3360 ) );
NOR2_X1 _u10_u6_U1354  ( .A1(_u10_SYNOPSYS_UNCONNECTED_26 ), .A2(_u10_SYNOPSYS_UNCONNECTED_27 ), .ZN(_u10_u6_n3136 ) );
NAND2_X1 _u10_u6_U1353  ( .A1(_u10_u6_n3360 ), .A2(_u10_u6_n3136 ), .ZN(_u10_u6_n2344 ) );
NOR2_X1 _u10_u6_U1352  ( .A1(_u10_u6_n3366 ), .A2(_u10_u6_n2344 ), .ZN(_u10_u6_n3385 ) );
NOR3_X1 _u10_u6_U1351  ( .A1(_u10_SYNOPSYS_UNCONNECTED_24 ), .A2(_u10_u6_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_28 ), .ZN(_u10_u6_n3342 ) );
NAND2_X1 _u10_u6_U1350  ( .A1(_u10_u6_n3342 ), .A2(_u10_u6_n3136 ), .ZN(_u10_u6_n2584 ) );
NOR2_X1 _u10_u6_U1349  ( .A1(_u10_u6_n2584 ), .A2(1'b0), .ZN(_u10_u6_n2139 ));
INV_X1 _u10_u6_U1348  ( .A(_u10_u6_n2216 ), .ZN(_u10_u6_n2106 ) );
AND2_X1 _u10_u6_U1347  ( .A1(_u10_u6_n2152 ), .A2(_u10_u6_n2106 ), .ZN(_u10_u6_n2336 ) );
NAND2_X1 _u10_u6_U1346  ( .A1(_u10_u6_n2139 ), .A2(_u10_u6_n2336 ), .ZN(_u10_u6_n2365 ) );
INV_X1 _u10_u6_U1345  ( .A(_u10_u6_n2365 ), .ZN(_u10_u6_n2004 ) );
AND2_X1 _u10_u6_U1344  ( .A1(_u10_u6_n2877 ), .A2(_u10_u6_n2004 ), .ZN(_u10_u6_n3386 ) );
NOR3_X1 _u10_u6_U1343  ( .A1(_u10_u6_n3384 ), .A2(_u10_u6_n3385 ), .A3(_u10_u6_n3386 ), .ZN(_u10_u6_n3383 ) );
NAND4_X1 _u10_u6_U1342  ( .A1(_u10_u6_n3380 ), .A2(_u10_u6_n3381 ), .A3(_u10_u6_n3382 ), .A4(_u10_u6_n3383 ), .ZN(_u10_u6_n3191 ) );
NAND2_X1 _u10_u6_U1341  ( .A1(_u10_u6_n2285 ), .A2(_u10_u6_n3379 ), .ZN(_u10_u6_n1975 ) );
NOR3_X1 _u10_u6_U1340  ( .A1(_u10_u6_n3378 ), .A2(1'b0), .A3(_u10_u6_n1975 ),.ZN(_u10_u6_n3122 ) );
AND4_X1 _u10_u6_U1339  ( .A1(_u10_u6_n2752 ), .A2(_u10_u6_n2383 ), .A3(_u10_u6_n1969 ), .A4(_u10_u6_n3122 ), .ZN(_u10_u6_n3377 ) );
NOR2_X1 _u10_u6_U1338  ( .A1(_u10_u6_n1814 ), .A2(_u10_u6_n1815 ), .ZN(_u10_u6_n3147 ) );
NAND2_X1 _u10_u6_U1337  ( .A1(_u10_u6_n3328 ), .A2(_u10_u6_n3147 ), .ZN(_u10_u6_n2359 ) );
NOR2_X1 _u10_u6_U1336  ( .A1(_u10_u6_n3377 ), .A2(_u10_u6_n2359 ), .ZN(_u10_u6_n3362 ) );
INV_X1 _u10_u6_U1335  ( .A(_u10_u6_n2008 ), .ZN(_u10_u6_n3097 ) );
NOR3_X1 _u10_u6_U1334  ( .A1(_u10_SYNOPSYS_UNCONNECTED_24 ), .A2(_u10_u6_n1813 ), .A3(_u10_SYNOPSYS_UNCONNECTED_25 ), .ZN(_u10_u6_n3269 ) );
NAND2_X1 _u10_u6_U1333  ( .A1(_u10_u6_n3269 ), .A2(_u10_u6_n3136 ), .ZN(_u10_u6_n3109 ) );
INV_X1 _u10_u6_U1332  ( .A(_u10_u6_n3109 ), .ZN(_u10_u6_n2999 ) );
INV_X1 _u10_u6_U1331  ( .A(_u10_u6_n2508 ), .ZN(_u10_u6_n2103 ) );
NAND2_X1 _u10_u6_U1330  ( .A1(_u10_u6_n2336 ), .A2(_u10_u6_n2103 ), .ZN(_u10_u6_n2249 ) );
NOR2_X1 _u10_u6_U1329  ( .A1(_u10_u6_n2249 ), .A2(1'b0), .ZN(_u10_u6_n1866 ));
NAND2_X1 _u10_u6_U1328  ( .A1(_u10_u6_n1866 ), .A2(_u10_u6_n1922 ), .ZN(_u10_u6_n2632 ) );
INV_X1 _u10_u6_U1327  ( .A(_u10_u6_n2223 ), .ZN(_u10_u6_n1918 ) );
NOR2_X1 _u10_u6_U1326  ( .A1(_u10_u6_n2632 ), .A2(_u10_u6_n1918 ), .ZN(_u10_u6_n1981 ) );
NAND3_X1 _u10_u6_U1325  ( .A1(_u10_u6_n3097 ), .A2(_u10_u6_n2999 ), .A3(_u10_u6_n1981 ), .ZN(_u10_u6_n3034 ) );
NOR3_X1 _u10_u6_U1324  ( .A1(_u10_SYNOPSYS_UNCONNECTED_25 ), .A2(_u10_SYNOPSYS_UNCONNECTED_24 ), .A3(_u10_SYNOPSYS_UNCONNECTED_28 ),.ZN(_u10_u6_n3302 ) );
NAND2_X1 _u10_u6_U1323  ( .A1(_u10_u6_n3302 ), .A2(_u10_u6_n3174 ), .ZN(_u10_u6_n3162 ) );
INV_X1 _u10_u6_U1322  ( .A(_u10_u6_n3162 ), .ZN(_u10_u6_n2979 ) );
NAND2_X1 _u10_u6_U1321  ( .A1(_u10_u6_n2979 ), .A2(_u10_u6_n2972 ), .ZN(_u10_u6_n1984 ) );
AND2_X1 _u10_u6_U1320  ( .A1(_u10_u6_n3302 ), .A2(_u10_u6_n3136 ), .ZN(_u10_u6_n2977 ) );
NAND3_X1 _u10_u6_U1319  ( .A1(_u10_u6_n2977 ), .A2(_u10_u6_n3000 ), .A3(_u10_u6_n3097 ), .ZN(_u10_u6_n3376 ) );
NAND2_X1 _u10_u6_U1318  ( .A1(_u10_u6_n1984 ), .A2(_u10_u6_n3376 ), .ZN(_u10_u6_n3375 ) );
NAND2_X1 _u10_u6_U1317  ( .A1(_u10_u6_n1981 ), .A2(_u10_u6_n3375 ), .ZN(_u10_u6_n2798 ) );
NAND2_X1 _u10_u6_U1316  ( .A1(_u10_u6_n3034 ), .A2(_u10_u6_n2798 ), .ZN(_u10_u6_n2007 ) );
NAND2_X1 _u10_u6_U1315  ( .A1(_u10_u6_n3269 ), .A2(_u10_u6_n3147 ), .ZN(_u10_u6_n2102 ) );
NOR2_X1 _u10_u6_U1314  ( .A1(_u10_u6_n2249 ), .A2(_u10_u6_n2102 ), .ZN(_u10_u6_n3323 ) );
INV_X1 _u10_u6_U1313  ( .A(_u10_u6_n3323 ), .ZN(_u10_u6_n3374 ) );
INV_X1 _u10_u6_U1312  ( .A(_u10_u6_n2344 ), .ZN(_u10_u6_n2002 ) );
NAND2_X1 _u10_u6_U1311  ( .A1(_u10_u6_n2336 ), .A2(_u10_u6_n2002 ), .ZN(_u10_u6_n3225 ) );
NAND2_X1 _u10_u6_U1310  ( .A1(_u10_u6_n3374 ), .A2(_u10_u6_n3225 ), .ZN(_u10_u6_n2488 ) );
NAND2_X1 _u10_u6_U1309  ( .A1(_u10_u6_n3342 ), .A2(_u10_u6_n3236 ), .ZN(_u10_u6_n2253 ) );
NOR2_X1 _u10_u6_U1308  ( .A1(_u10_u6_n2253 ), .A2(1'b0), .ZN(_u10_u6_n1885 ));
NAND2_X1 _u10_u6_U1307  ( .A1(_u10_u6_n3360 ), .A2(_u10_u6_n3174 ), .ZN(_u10_u6_n2254 ) );
INV_X1 _u10_u6_U1306  ( .A(_u10_u6_n2254 ), .ZN(_u10_u6_n2986 ) );
NAND2_X1 _u10_u6_U1305  ( .A1(_u10_u6_n2106 ), .A2(_u10_u6_n2986 ), .ZN(_u10_u6_n1913 ) );
INV_X1 _u10_u6_U1304  ( .A(_u10_u6_n1913 ), .ZN(_u10_u6_n2377 ) );
OR4_X1 _u10_u6_U1303  ( .A1(_u10_u6_n2007 ), .A2(_u10_u6_n2488 ), .A3(_u10_u6_n1885 ), .A4(_u10_u6_n2377 ), .ZN(_u10_u6_n3373 ) );
NAND2_X1 _u10_u6_U1302  ( .A1(_u10_u6_n2534 ), .A2(_u10_u6_n3373 ), .ZN(_u10_u6_n3370 ) );
NAND2_X1 _u10_u6_U1301  ( .A1(_u10_u6_n3342 ), .A2(_u10_u6_n3174 ), .ZN(_u10_u6_n2037 ) );
NAND2_X1 _u10_u6_U1300  ( .A1(_u10_u6_n2037 ), .A2(_u10_u6_n2254 ), .ZN(_u10_u6_n3372 ) );
NAND2_X1 _u10_u6_U1299  ( .A1(_u10_u6_n2003 ), .A2(_u10_u6_n3372 ), .ZN(_u10_u6_n3371 ) );
NAND2_X1 _u10_u6_U1298  ( .A1(_u10_u6_n3370 ), .A2(_u10_u6_n3371 ), .ZN(_u10_u6_n3363 ) );
NOR2_X1 _u10_u6_U1297  ( .A1(_u10_u6_n2490 ), .A2(_u10_u6_n1961 ), .ZN(_u10_u6_n3369 ) );
NAND2_X1 _u10_u6_U1296  ( .A1(_u10_u6_n2534 ), .A2(_u10_u6_n2049 ), .ZN(_u10_u6_n2646 ) );
INV_X1 _u10_u6_U1295  ( .A(_u10_u6_n2646 ), .ZN(_u10_u6_n3055 ) );
NOR2_X1 _u10_u6_U1294  ( .A1(_u10_u6_n3369 ), .A2(_u10_u6_n3055 ), .ZN(_u10_u6_n3367 ) );
NAND2_X1 _u10_u6_U1293  ( .A1(_u10_u6_n3368 ), .A2(_u10_u6_n3147 ), .ZN(_u10_u6_n2495 ) );
NOR2_X1 _u10_u6_U1292  ( .A1(_u10_u6_n3367 ), .A2(_u10_u6_n2495 ), .ZN(_u10_u6_n3364 ) );
INV_X1 _u10_u6_U1291  ( .A(_u10_u6_n2139 ), .ZN(_u10_u6_n3254 ) );
NOR2_X1 _u10_u6_U1290  ( .A1(_u10_u6_n3366 ), .A2(_u10_u6_n3254 ), .ZN(_u10_u6_n3365 ) );
NOR4_X1 _u10_u6_U1289  ( .A1(_u10_u6_n3362 ), .A2(_u10_u6_n3363 ), .A3(_u10_u6_n3364 ), .A4(_u10_u6_n3365 ), .ZN(_u10_u6_n3305 ) );
NAND2_X1 _u10_u6_U1288  ( .A1(_u10_u6_n3302 ), .A2(_u10_u6_n3147 ), .ZN(_u10_u6_n2980 ) );
NAND2_X1 _u10_u6_U1287  ( .A1(_u10_u6_n2102 ), .A2(_u10_u6_n2980 ), .ZN(_u10_u6_n2177 ) );
NAND2_X1 _u10_u6_U1286  ( .A1(_u10_u6_n2003 ), .A2(_u10_u6_n2493 ), .ZN(_u10_u6_n1962 ) );
NAND2_X1 _u10_u6_U1285  ( .A1(_u10_u6_n1961 ), .A2(_u10_u6_n1962 ), .ZN(_u10_u6_n3361 ) );
NAND2_X1 _u10_u6_U1284  ( .A1(_u10_u6_n2177 ), .A2(_u10_u6_n3361 ), .ZN(_u10_u6_n3357 ) );
NAND2_X1 _u10_u6_U1283  ( .A1(_u10_u6_n3236 ), .A2(_u10_u6_n3360 ), .ZN(_u10_u6_n1859 ) );
INV_X1 _u10_u6_U1282  ( .A(_u10_u6_n1859 ), .ZN(_u10_u6_n2256 ) );
NAND3_X1 _u10_u6_U1281  ( .A1(_u10_u6_n2256 ), .A2(_u10_u6_n2113 ), .A3(_u10_u6_n2128 ), .ZN(_u10_u6_n3358 ) );
NOR2_X1 _u10_u6_U1280  ( .A1(_u10_u6_n2877 ), .A2(_u10_u6_n3222 ), .ZN(_u10_u6_n3347 ) );
NAND2_X1 _u10_u6_U1279  ( .A1(_u10_u6_n3347 ), .A2(_u10_u6_n1869 ), .ZN(_u10_u6_n2005 ) );
NAND2_X1 _u10_u6_U1278  ( .A1(_u10_u6_n2488 ), .A2(_u10_u6_n2005 ), .ZN(_u10_u6_n3359 ) );
NAND3_X1 _u10_u6_U1277  ( .A1(_u10_u6_n3357 ), .A2(_u10_u6_n3358 ), .A3(_u10_u6_n3359 ), .ZN(_u10_u6_n3352 ) );
NAND2_X1 _u10_u6_U1276  ( .A1(_u10_u6_n3320 ), .A2(_u10_u6_n3136 ), .ZN(_u10_u6_n2356 ) );
INV_X1 _u10_u6_U1275  ( .A(_u10_u6_n2356 ), .ZN(_u10_u6_n2830 ) );
NAND2_X1 _u10_u6_U1274  ( .A1(_u10_u6_n2830 ), .A2(_u10_u6_n2836 ), .ZN(_u10_u6_n2291 ) );
NOR3_X1 _u10_u6_U1273  ( .A1(_u10_u6_n2291 ), .A2(_u10_u6_n2330 ), .A3(_u10_u6_n2022 ), .ZN(_u10_u6_n3353 ) );
INV_X1 _u10_u6_U1272  ( .A(_u10_u6_n1925 ), .ZN(_u10_u6_n2105 ) );
AND2_X1 _u10_u6_U1271  ( .A1(_u10_u6_n2108 ), .A2(_u10_u6_n2105 ), .ZN(_u10_u6_n2915 ) );
INV_X1 _u10_u6_U1270  ( .A(_u10_u6_n2330 ), .ZN(_u10_u6_n2107 ) );
NAND2_X1 _u10_u6_U1269  ( .A1(_u10_u6_n2915 ), .A2(_u10_u6_n2107 ), .ZN(_u10_u6_n2203 ) );
INV_X1 _u10_u6_U1268  ( .A(_u10_u6_n2203 ), .ZN(_u10_u6_n1982 ) );
NAND2_X1 _u10_u6_U1267  ( .A1(_u10_u6_n1982 ), .A2(_u10_u6_n2536 ), .ZN(_u10_u6_n2587 ) );
INV_X1 _u10_u6_U1266  ( .A(_u10_u6_n2587 ), .ZN(_u10_u6_n2697 ) );
NAND3_X1 _u10_u6_U1265  ( .A1(_u10_u6_n2697 ), .A2(_u10_u6_n2493 ), .A3(_u10_u6_n2377 ), .ZN(_u10_u6_n2412 ) );
INV_X1 _u10_u6_U1264  ( .A(_u10_u6_n2412 ), .ZN(_u10_u6_n3354 ) );
NAND2_X1 _u10_u6_U1263  ( .A1(_u10_u6_n3174 ), .A2(_u10_u6_n3269 ), .ZN(_u10_u6_n2375 ) );
INV_X1 _u10_u6_U1262  ( .A(_u10_u6_n2375 ), .ZN(_u10_u6_n2507 ) );
NAND2_X1 _u10_u6_U1261  ( .A1(_u10_u6_n1981 ), .A2(_u10_u6_n2507 ), .ZN(_u10_u6_n2621 ) );
NOR4_X1 _u10_u6_U1260  ( .A1(1'b0), .A2(_u10_u6_n3356 ), .A3(_u10_u6_n2203 ),.A4(_u10_u6_n2621 ), .ZN(_u10_u6_n3355 ) );
NOR4_X1 _u10_u6_U1259  ( .A1(_u10_u6_n3352 ), .A2(_u10_u6_n3353 ), .A3(_u10_u6_n3354 ), .A4(_u10_u6_n3355 ), .ZN(_u10_u6_n3306 ) );
NOR2_X1 _u10_u6_U1258  ( .A1(_u10_u6_n2842 ), .A2(_u10_u6_n2356 ), .ZN(_u10_u6_n1891 ) );
INV_X1 _u10_u6_U1257  ( .A(_u10_u6_n1869 ), .ZN(_u10_u6_n2885 ) );
NAND2_X1 _u10_u6_U1256  ( .A1(_u10_u6_n1891 ), .A2(_u10_u6_n2885 ), .ZN(_u10_u6_n3330 ) );
NAND2_X1 _u10_u6_U1255  ( .A1(_u10_u6_n2761 ), .A2(_u10_u6_n2837 ), .ZN(_u10_u6_n3351 ) );
NAND3_X1 _u10_u6_U1254  ( .A1(_u10_u6_n2884 ), .A2(_u10_u6_n2080 ), .A3(_u10_u6_n2915 ), .ZN(_u10_u6_n2762 ) );
NAND2_X1 _u10_u6_U1253  ( .A1(_u10_u6_n2055 ), .A2(_u10_u6_n2019 ), .ZN(_u10_u6_n3259 ) );
NAND4_X1 _u10_u6_U1252  ( .A1(_u10_u6_n3351 ), .A2(_u10_u6_n2762 ), .A3(_u10_u6_n2061 ), .A4(_u10_u6_n3259 ), .ZN(_u10_u6_n3350 ) );
NAND2_X1 _u10_u6_U1251  ( .A1(_u10_u6_n2183 ), .A2(_u10_u6_n3350 ), .ZN(_u10_u6_n3331 ) );
NAND2_X1 _u10_u6_U1250  ( .A1(_u10_u6_n3349 ), .A2(_u10_u6_n2305 ), .ZN(_u10_u6_n3348 ) );
NAND2_X1 _u10_u6_U1249  ( .A1(_u10_u6_n1896 ), .A2(_u10_u6_n3348 ), .ZN(_u10_u6_n3176 ) );
NAND2_X1 _u10_u6_U1248  ( .A1(_u10_u6_n2461 ), .A2(_u10_u6_n3176 ), .ZN(_u10_u6_n3332 ) );
INV_X1 _u10_u6_U1247  ( .A(_u10_u6_n2495 ), .ZN(_u10_u6_n2063 ) );
NAND2_X1 _u10_u6_U1246  ( .A1(_u10_u6_n2049 ), .A2(_u10_u6_n2063 ), .ZN(_u10_u6_n2886 ) );
NOR2_X1 _u10_u6_U1245  ( .A1(_u10_u6_n3347 ), .A2(_u10_u6_n2886 ), .ZN(_u10_u6_n3334 ) );
NAND2_X1 _u10_u6_U1244  ( .A1(1'b0), .A2(_u10_u6_n2835 ), .ZN(_u10_u6_n3344 ) );
NAND2_X1 _u10_u6_U1243  ( .A1(_u10_u6_n2001 ), .A2(_u10_u6_n2905 ), .ZN(_u10_u6_n3346 ) );
NAND2_X1 _u10_u6_U1242  ( .A1(_u10_u6_n3346 ), .A2(_u10_u6_n2803 ), .ZN(_u10_u6_n3345 ) );
NAND2_X1 _u10_u6_U1241  ( .A1(_u10_u6_n2087 ), .A2(_u10_u6_n2835 ), .ZN(_u10_u6_n2413 ) );
INV_X1 _u10_u6_U1240  ( .A(_u10_u6_n2128 ), .ZN(_u10_u6_n2235 ) );
NAND4_X1 _u10_u6_U1239  ( .A1(_u10_u6_n3344 ), .A2(_u10_u6_n3345 ), .A3(_u10_u6_n2413 ), .A4(_u10_u6_n2235 ), .ZN(_u10_u6_n3329 ) );
NOR2_X1 _u10_u6_U1238  ( .A1(_u10_u6_n1915 ), .A2(_u10_u6_n3340 ), .ZN(_u10_u6_n3343 ) );
NOR3_X1 _u10_u6_U1237  ( .A1(_u10_u6_n3329 ), .A2(1'b0), .A3(_u10_u6_n3343 ),.ZN(_u10_u6_n3341 ) );
NAND2_X1 _u10_u6_U1236  ( .A1(_u10_u6_n3342 ), .A2(_u10_u6_n3147 ), .ZN(_u10_u6_n2688 ) );
NOR2_X1 _u10_u6_U1235  ( .A1(_u10_u6_n3341 ), .A2(_u10_u6_n2688 ), .ZN(_u10_u6_n3335 ) );
NOR2_X1 _u10_u6_U1234  ( .A1(_u10_u6_n2256 ), .A2(_u10_u6_n1885 ), .ZN(_u10_u6_n2689 ) );
NOR2_X1 _u10_u6_U1233  ( .A1(1'b0), .A2(_u10_u6_n2413 ), .ZN(_u10_u6_n3338 ));
NOR2_X1 _u10_u6_U1232  ( .A1(_u10_u6_n1925 ), .A2(_u10_u6_n3340 ), .ZN(_u10_u6_n3339 ) );
NOR3_X1 _u10_u6_U1231  ( .A1(_u10_u6_n2005 ), .A2(_u10_u6_n3338 ), .A3(_u10_u6_n3339 ), .ZN(_u10_u6_n3337 ) );
NOR2_X1 _u10_u6_U1230  ( .A1(_u10_u6_n2689 ), .A2(_u10_u6_n3337 ), .ZN(_u10_u6_n3336 ) );
NOR3_X1 _u10_u6_U1229  ( .A1(_u10_u6_n3334 ), .A2(_u10_u6_n3335 ), .A3(_u10_u6_n3336 ), .ZN(_u10_u6_n3333 ) );
NAND4_X1 _u10_u6_U1228  ( .A1(_u10_u6_n3330 ), .A2(_u10_u6_n3331 ), .A3(_u10_u6_n3332 ), .A4(_u10_u6_n3333 ), .ZN(_u10_u6_n3308 ) );
NAND3_X1 _u10_u6_U1227  ( .A1(_u10_SYNOPSYS_UNCONNECTED_28 ), .A2(_u10_SYNOPSYS_UNCONNECTED_25 ), .A3(_u10_u6_n3147 ), .ZN(_u10_u6_n2126 ) );
INV_X1 _u10_u6_U1226  ( .A(_u10_u6_n2126 ), .ZN(_u10_u6_n2329 ) );
NAND2_X1 _u10_u6_U1225  ( .A1(_u10_u6_n2329 ), .A2(_u10_u6_n3329 ), .ZN(_u10_u6_n3324 ) );
NAND2_X1 _u10_u6_U1224  ( .A1(_u10_u6_n3328 ), .A2(_u10_u6_n3136 ), .ZN(_u10_u6_n2000 ) );
INV_X1 _u10_u6_U1223  ( .A(_u10_u6_n2000 ), .ZN(_u10_u6_n2445 ) );
NAND3_X1 _u10_u6_U1222  ( .A1(_u10_u6_n2446 ), .A2(_u10_u6_n3001 ), .A3(_u10_u6_n2087 ), .ZN(_u10_u6_n3327 ) );
NAND2_X1 _u10_u6_U1221  ( .A1(_u10_u6_n3327 ), .A2(_u10_u6_n2905 ), .ZN(_u10_u6_n2500 ) );
NAND2_X1 _u10_u6_U1220  ( .A1(_u10_u6_n2445 ), .A2(_u10_u6_n2500 ), .ZN(_u10_u6_n3325 ) );
NAND2_X1 _u10_u6_U1219  ( .A1(1'b0), .A2(_u10_u6_n2979 ), .ZN(_u10_u6_n3326 ) );
NAND3_X1 _u10_u6_U1218  ( .A1(_u10_u6_n3324 ), .A2(_u10_u6_n3325 ), .A3(_u10_u6_n3326 ), .ZN(_u10_u6_n3309 ) );
AND2_X1 _u10_u6_U1217  ( .A1(_u10_u6_n2877 ), .A2(_u10_u6_n3223 ), .ZN(_u10_u6_n2858 ) );
NAND2_X1 _u10_u6_U1216  ( .A1(_u10_u6_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_26 ), .ZN(_u10_u6_n2346 ) );
INV_X1 _u10_u6_U1215  ( .A(_u10_u6_n2346 ), .ZN(_u10_u6_n2043 ) );
NAND2_X1 _u10_u6_U1214  ( .A1(_u10_u6_n2858 ), .A2(_u10_u6_n2043 ), .ZN(_u10_u6_n3321 ) );
NAND2_X1 _u10_u6_U1213  ( .A1(_u10_u6_n1982 ), .A2(_u10_u6_n2195 ), .ZN(_u10_u6_n3268 ) );
INV_X1 _u10_u6_U1212  ( .A(_u10_u6_n3268 ), .ZN(_u10_u6_n2222 ) );
NAND3_X1 _u10_u6_U1211  ( .A1(_u10_u6_n3323 ), .A2(_u10_u6_n3216 ), .A3(_u10_u6_n2222 ), .ZN(_u10_u6_n3322 ) );
NAND2_X1 _u10_u6_U1210  ( .A1(_u10_u6_n3321 ), .A2(_u10_u6_n3322 ), .ZN(_u10_u6_n2374 ) );
NAND2_X1 _u10_u6_U1209  ( .A1(_u10_u6_n3320 ), .A2(_u10_u6_n3174 ), .ZN(_u10_u6_n2014 ) );
NOR2_X1 _u10_u6_U1208  ( .A1(_u10_u6_n1841 ), .A2(_u10_u6_n2014 ), .ZN(_u10_u6_n2813 ) );
NAND2_X1 _u10_u6_U1207  ( .A1(_u10_u6_n2813 ), .A2(_u10_u6_n2534 ), .ZN(_u10_u6_n3310 ) );
NAND2_X1 _u10_u6_U1206  ( .A1(_u10_u6_n3319 ), .A2(_u10_u6_n3136 ), .ZN(_u10_u6_n1836 ) );
INV_X1 _u10_u6_U1205  ( .A(_u10_u6_n1836 ), .ZN(_u10_u6_n2815 ) );
NAND2_X1 _u10_u6_U1204  ( .A1(_u10_u6_n2534 ), .A2(_u10_u6_n3129 ), .ZN(_u10_u6_n2439 ) );
NAND2_X1 _u10_u6_U1203  ( .A1(_u10_u6_n2055 ), .A2(_u10_u6_n2107 ), .ZN(_u10_u6_n2062 ) );
NAND2_X1 _u10_u6_U1202  ( .A1(_u10_u6_n2439 ), .A2(_u10_u6_n2062 ), .ZN(_u10_u6_n3318 ) );
NAND2_X1 _u10_u6_U1201  ( .A1(_u10_u6_n2815 ), .A2(_u10_u6_n3318 ), .ZN(_u10_u6_n3311 ) );
NAND2_X1 _u10_u6_U1200  ( .A1(_u10_u6_n2986 ), .A2(_u10_u6_n2175 ), .ZN(_u10_u6_n3317 ) );
NAND2_X1 _u10_u6_U1199  ( .A1(_u10_u6_n2253 ), .A2(_u10_u6_n3317 ), .ZN(_u10_u6_n3157 ) );
NAND2_X1 _u10_u6_U1198  ( .A1(_u10_u6_n3316 ), .A2(_u10_u6_n3157 ), .ZN(_u10_u6_n3312 ) );
NOR2_X1 _u10_u6_U1197  ( .A1(_u10_u6_n2495 ), .A2(_u10_u6_n2194 ), .ZN(_u10_u6_n3314 ) );
NOR2_X1 _u10_u6_U1196  ( .A1(_u10_u6_n2375 ), .A2(_u10_u6_n2367 ), .ZN(_u10_u6_n3315 ) );
NOR2_X1 _u10_u6_U1195  ( .A1(_u10_u6_n3314 ), .A2(_u10_u6_n3315 ), .ZN(_u10_u6_n3313 ) );
NAND4_X1 _u10_u6_U1194  ( .A1(_u10_u6_n3310 ), .A2(_u10_u6_n3311 ), .A3(_u10_u6_n3312 ), .A4(_u10_u6_n3313 ), .ZN(_u10_u6_n2315 ) );
NOR4_X1 _u10_u6_U1193  ( .A1(_u10_u6_n3308 ), .A2(_u10_u6_n3309 ), .A3(_u10_u6_n2374 ), .A4(_u10_u6_n2315 ), .ZN(_u10_u6_n3307 ) );
NAND3_X1 _u10_u6_U1192  ( .A1(_u10_u6_n3305 ), .A2(_u10_u6_n3306 ), .A3(_u10_u6_n3307 ), .ZN(_u10_u6_n1987 ) );
AND2_X1 _u10_u6_U1191  ( .A1(1'b0), .A2(_u10_u6_n2977 ), .ZN(_u10_u6_n3240 ));
NAND2_X1 _u10_u6_U1190  ( .A1(_u10_u6_n1891 ), .A2(_u10_u6_n2534 ), .ZN(_u10_u6_n3303 ) );
NAND4_X1 _u10_u6_U1189  ( .A1(_u10_u6_n1982 ), .A2(_u10_u6_n2659 ), .A3(_u10_u6_n2256 ), .A4(_u10_u6_n2175 ), .ZN(_u10_u6_n3304 ) );
AND2_X1 _u10_u6_U1188  ( .A1(_u10_u6_n3303 ), .A2(_u10_u6_n3304 ), .ZN(_u10_u6_n2612 ) );
NAND2_X1 _u10_u6_U1187  ( .A1(_u10_u6_n3302 ), .A2(_u10_u6_n3236 ), .ZN(_u10_u6_n2985 ) );
OR2_X1 _u10_u6_U1186  ( .A1(_u10_u6_n2431 ), .A2(_u10_u6_n2985 ), .ZN(_u10_u6_n3299 ) );
OR2_X1 _u10_u6_U1185  ( .A1(_u10_u6_n2282 ), .A2(_u10_u6_n2359 ), .ZN(_u10_u6_n3300 ) );
NAND2_X1 _u10_u6_U1184  ( .A1(_u10_u6_n1890 ), .A2(_u10_u6_n2534 ), .ZN(_u10_u6_n3301 ) );
NAND4_X1 _u10_u6_U1183  ( .A1(_u10_u6_n2612 ), .A2(_u10_u6_n3299 ), .A3(_u10_u6_n3300 ), .A4(_u10_u6_n3301 ), .ZN(_u10_u6_n3279 ) );
INV_X1 _u10_u6_U1182  ( .A(_u10_u6_n2464 ), .ZN(_u10_u6_n3295 ) );
NAND2_X1 _u10_u6_U1181  ( .A1(_u10_u6_n3295 ), .A2(_u10_u6_n2835 ), .ZN(_u10_u6_n2623 ) );
INV_X1 _u10_u6_U1180  ( .A(_u10_u6_n2623 ), .ZN(_u10_u6_n3185 ) );
INV_X1 _u10_u6_U1179  ( .A(_u10_u6_n2688 ), .ZN(_u10_u6_n2169 ) );
NAND2_X1 _u10_u6_U1178  ( .A1(_u10_u6_n3185 ), .A2(_u10_u6_n2169 ), .ZN(_u10_u6_n3286 ) );
NAND2_X1 _u10_u6_U1177  ( .A1(_u10_u6_n2833 ), .A2(_u10_u6_n3278 ), .ZN(_u10_u6_n3298 ) );
NAND3_X1 _u10_u6_U1176  ( .A1(_u10_u6_n3297 ), .A2(_u10_u6_n2838 ), .A3(_u10_u6_n3298 ), .ZN(_u10_u6_n3296 ) );
NAND2_X1 _u10_u6_U1175  ( .A1(_u10_u6_n2830 ), .A2(_u10_u6_n3296 ), .ZN(_u10_u6_n3287 ) );
NAND2_X1 _u10_u6_U1174  ( .A1(_u10_u6_n3295 ), .A2(_u10_u6_n3001 ), .ZN(_u10_u6_n3292 ) );
NAND2_X1 _u10_u6_U1173  ( .A1(_u10_u6_n3294 ), .A2(_u10_u6_n2089 ), .ZN(_u10_u6_n3293 ) );
AND2_X1 _u10_u6_U1172  ( .A1(_u10_u6_n3292 ), .A2(_u10_u6_n3293 ), .ZN(_u10_u6_n2548 ) );
NAND2_X1 _u10_u6_U1171  ( .A1(_u10_u6_n2548 ), .A2(_u10_u6_n2091 ), .ZN(_u10_u6_n2304 ) );
NAND2_X1 _u10_u6_U1170  ( .A1(_u10_u6_n2304 ), .A2(_u10_u6_n2446 ), .ZN(_u10_u6_n3290 ) );
NAND2_X1 _u10_u6_U1169  ( .A1(_u10_u6_n2549 ), .A2(_u10_u6_n2446 ), .ZN(_u10_u6_n2790 ) );
NOR2_X1 _u10_u6_U1168  ( .A1(_u10_u6_n1936 ), .A2(_u10_u6_n2790 ), .ZN(_u10_u6_n2789 ) );
INV_X1 _u10_u6_U1167  ( .A(_u10_u6_n2789 ), .ZN(_u10_u6_n3291 ) );
OR2_X1 _u10_u6_U1166  ( .A1(_u10_u6_n2828 ), .A2(_u10_u6_n2790 ), .ZN(_u10_u6_n2498 ) );
NAND4_X1 _u10_u6_U1165  ( .A1(_u10_u6_n3290 ), .A2(_u10_u6_n3291 ), .A3(_u10_u6_n2498 ), .A4(_u10_u6_n2001 ), .ZN(_u10_u6_n3289 ) );
NAND2_X1 _u10_u6_U1164  ( .A1(_u10_u6_n2445 ), .A2(_u10_u6_n3289 ), .ZN(_u10_u6_n3288 ) );
NAND3_X1 _u10_u6_U1163  ( .A1(_u10_u6_n3286 ), .A2(_u10_u6_n3287 ), .A3(_u10_u6_n3288 ), .ZN(_u10_u6_n3280 ) );
NOR2_X1 _u10_u6_U1162  ( .A1(_u10_u6_n2940 ), .A2(_u10_u6_n1913 ), .ZN(_u10_u6_n3281 ) );
INV_X1 _u10_u6_U1161  ( .A(1'b0), .ZN(_u10_u6_n1864 ) );
NAND2_X1 _u10_u6_U1160  ( .A1(1'b0), .A2(_u10_u6_n2588 ), .ZN(_u10_u6_n2141 ) );
INV_X1 _u10_u6_U1159  ( .A(_u10_u6_n2141 ), .ZN(_u10_u6_n3159 ) );
NAND3_X1 _u10_u6_U1158  ( .A1(_u10_u6_n2103 ), .A2(_u10_u6_n1864 ), .A3(_u10_u6_n3159 ), .ZN(_u10_u6_n2520 ) );
INV_X1 _u10_u6_U1157  ( .A(_u10_u6_n2520 ), .ZN(_u10_u6_n2630 ) );
INV_X1 _u10_u6_U1156  ( .A(_u10_u6_n2307 ), .ZN(_u10_u6_n2382 ) );
NOR4_X1 _u10_u6_U1155  ( .A1(_u10_u6_n2382 ), .A2(_u10_u6_n2722 ), .A3(_u10_u6_n1925 ), .A4(_u10_u6_n2508 ), .ZN(_u10_u6_n3260 ) );
NOR2_X1 _u10_u6_U1154  ( .A1(_u10_u6_n2498 ), .A2(_u10_u6_n2911 ), .ZN(_u10_u6_n2633 ) );
NOR2_X1 _u10_u6_U1153  ( .A1(_u10_u6_n2633 ), .A2(_u10_u6_n3278 ), .ZN(_u10_u6_n3285 ) );
INV_X1 _u10_u6_U1152  ( .A(_u10_u6_n1866 ), .ZN(_u10_u6_n1926 ) );
NOR2_X1 _u10_u6_U1151  ( .A1(_u10_u6_n3285 ), .A2(_u10_u6_n1926 ), .ZN(_u10_u6_n3284 ) );
NOR4_X1 _u10_u6_U1150  ( .A1(1'b0), .A2(_u10_u6_n2630 ), .A3(_u10_u6_n3260 ),.A4(_u10_u6_n3284 ), .ZN(_u10_u6_n3283 ) );
NOR2_X1 _u10_u6_U1149  ( .A1(_u10_u6_n3283 ), .A2(_u10_u6_n2980 ), .ZN(_u10_u6_n3282 ) );
NOR4_X1 _u10_u6_U1148  ( .A1(_u10_u6_n3279 ), .A2(_u10_u6_n3280 ), .A3(_u10_u6_n3281 ), .A4(_u10_u6_n3282 ), .ZN(_u10_u6_n3241 ) );
NAND2_X1 _u10_u6_U1147  ( .A1(_u10_u6_n1836 ), .A2(_u10_u6_n2291 ), .ZN(_u10_u6_n2147 ) );
NAND2_X1 _u10_u6_U1146  ( .A1(_u10_u6_n2443 ), .A2(_u10_u6_n2147 ), .ZN(_u10_u6_n3261 ) );
INV_X1 _u10_u6_U1145  ( .A(_u10_u6_n1841 ), .ZN(_u10_u6_n2571 ) );
NAND2_X1 _u10_u6_U1144  ( .A1(_u10_u6_n2571 ), .A2(_u10_u6_n3278 ), .ZN(_u10_u6_n3277 ) );
NAND2_X1 _u10_u6_U1143  ( .A1(_u10_u6_n3276 ), .A2(_u10_u6_n3277 ), .ZN(_u10_u6_n2819 ) );
OR2_X1 _u10_u6_U1142  ( .A1(_u10_u6_n2819 ), .A2(_u10_u6_n3275 ), .ZN(_u10_u6_n3273 ) );
NAND2_X1 _u10_u6_U1141  ( .A1(_u10_u6_n2815 ), .A2(_u10_u6_n2080 ), .ZN(_u10_u6_n3274 ) );
NAND2_X1 _u10_u6_U1140  ( .A1(_u10_u6_n2014 ), .A2(_u10_u6_n3274 ), .ZN(_u10_u6_n2165 ) );
NAND2_X1 _u10_u6_U1139  ( .A1(_u10_u6_n3273 ), .A2(_u10_u6_n2165 ), .ZN(_u10_u6_n3262 ) );
NAND2_X1 _u10_u6_U1138  ( .A1(_u10_u6_n2688 ), .A2(_u10_u6_n2126 ), .ZN(_u10_u6_n1956 ) );
INV_X1 _u10_u6_U1137  ( .A(_u10_u6_n1956 ), .ZN(_u10_u6_n1860 ) );
NOR2_X1 _u10_u6_U1136  ( .A1(1'b0), .A2(_u10_u6_n2498 ), .ZN(_u10_u6_n3271 ));
NOR2_X1 _u10_u6_U1135  ( .A1(_u10_u6_n3271 ), .A2(_u10_u6_n3272 ), .ZN(_u10_u6_n3270 ) );
NOR2_X1 _u10_u6_U1134  ( .A1(_u10_u6_n1860 ), .A2(_u10_u6_n3270 ), .ZN(_u10_u6_n3264 ) );
INV_X1 _u10_u6_U1133  ( .A(_u10_u6_n2632 ), .ZN(_u10_u6_n3202 ) );
NAND2_X1 _u10_u6_U1132  ( .A1(_u10_u6_n3236 ), .A2(_u10_u6_n3269 ), .ZN(_u10_u6_n3036 ) );
INV_X1 _u10_u6_U1131  ( .A(_u10_u6_n3036 ), .ZN(_u10_u6_n1960 ) );
NAND2_X1 _u10_u6_U1130  ( .A1(_u10_u6_n3202 ), .A2(_u10_u6_n1960 ), .ZN(_u10_u6_n3079 ) );
NOR3_X1 _u10_u6_U1129  ( .A1(_u10_u6_n3079 ), .A2(1'b0), .A3(_u10_u6_n3268 ),.ZN(_u10_u6_n3265 ) );
INV_X1 _u10_u6_U1128  ( .A(_u10_u6_n2014 ), .ZN(_u10_u6_n2709 ) );
NAND2_X1 _u10_u6_U1127  ( .A1(_u10_u6_n2709 ), .A2(_u10_u6_n2166 ), .ZN(_u10_u6_n2145 ) );
INV_X1 _u10_u6_U1126  ( .A(_u10_u6_n2145 ), .ZN(_u10_u6_n3258 ) );
NOR2_X1 _u10_u6_U1125  ( .A1(_u10_u6_n3258 ), .A2(_u10_u6_n2183 ), .ZN(_u10_u6_n3267 ) );
NOR2_X1 _u10_u6_U1124  ( .A1(_u10_u6_n3267 ), .A2(_u10_u6_n2567 ), .ZN(_u10_u6_n3266 ) );
NOR3_X1 _u10_u6_U1123  ( .A1(_u10_u6_n3264 ), .A2(_u10_u6_n3265 ), .A3(_u10_u6_n3266 ), .ZN(_u10_u6_n3263 ) );
NAND3_X1 _u10_u6_U1122  ( .A1(_u10_u6_n3261 ), .A2(_u10_u6_n3262 ), .A3(_u10_u6_n3263 ), .ZN(_u10_u6_n3243 ) );
INV_X1 _u10_u6_U1121  ( .A(_u10_u6_n2102 ), .ZN(_u10_u6_n2509 ) );
NAND2_X1 _u10_u6_U1120  ( .A1(_u10_u6_n3260 ), .A2(_u10_u6_n2509 ), .ZN(_u10_u6_n3247 ) );
INV_X1 _u10_u6_U1119  ( .A(_u10_u6_n3259 ), .ZN(_u10_u6_n2015 ) );
NAND2_X1 _u10_u6_U1118  ( .A1(_u10_u6_n2015 ), .A2(_u10_u6_n3258 ), .ZN(_u10_u6_n3248 ) );
NAND2_X1 _u10_u6_U1117  ( .A1(_u10_u6_n2251 ), .A2(_u10_u6_n2169 ), .ZN(_u10_u6_n3255 ) );
OR2_X1 _u10_u6_U1116  ( .A1(_u10_u6_n3157 ), .A2(_u10_u6_n2256 ), .ZN(_u10_u6_n3257 ) );
NAND2_X1 _u10_u6_U1115  ( .A1(_u10_u6_n2105 ), .A2(_u10_u6_n3257 ), .ZN(_u10_u6_n3256 ) );
AND2_X1 _u10_u6_U1114  ( .A1(_u10_u6_n3255 ), .A2(_u10_u6_n3256 ), .ZN(_u10_u6_n3212 ) );
INV_X1 _u10_u6_U1113  ( .A(_u10_u6_n2037 ), .ZN(_u10_u6_n2987 ) );
NAND2_X1 _u10_u6_U1112  ( .A1(_u10_u6_n2987 ), .A2(_u10_u6_n2038 ), .ZN(_u10_u6_n2212 ) );
NOR2_X1 _u10_u6_U1111  ( .A1(_u10_u6_n2212 ), .A2(1'b0), .ZN(_u10_u6_n2658 ));
INV_X1 _u10_u6_U1110  ( .A(_u10_u6_n2658 ), .ZN(_u10_u6_n2343 ) );
NAND2_X1 _u10_u6_U1109  ( .A1(_u10_u6_n2344 ), .A2(_u10_u6_n3254 ), .ZN(_u10_u6_n1928 ) );
NAND2_X1 _u10_u6_U1108  ( .A1(_u10_u6_n2588 ), .A2(_u10_u6_n1928 ), .ZN(_u10_u6_n3253 ) );
NAND2_X1 _u10_u6_U1107  ( .A1(_u10_u6_n2343 ), .A2(_u10_u6_n3253 ), .ZN(_u10_u6_n3252 ) );
NAND2_X1 _u10_u6_U1106  ( .A1(_u10_u6_n2105 ), .A2(_u10_u6_n3252 ), .ZN(_u10_u6_n3251 ) );
NAND2_X1 _u10_u6_U1105  ( .A1(_u10_u6_n3212 ), .A2(_u10_u6_n3251 ), .ZN(_u10_u6_n3250 ) );
NAND2_X1 _u10_u6_U1104  ( .A1(_u10_u6_n2307 ), .A2(_u10_u6_n3250 ), .ZN(_u10_u6_n3249 ) );
NAND3_X1 _u10_u6_U1103  ( .A1(_u10_u6_n3247 ), .A2(_u10_u6_n3248 ), .A3(_u10_u6_n3249 ), .ZN(_u10_u6_n3244 ) );
AND2_X1 _u10_u6_U1102  ( .A1(_u10_u6_n2915 ), .A2(_u10_u6_n2059 ), .ZN(_u10_u6_n2957 ) );
AND3_X1 _u10_u6_U1101  ( .A1(_u10_u6_n3223 ), .A2(_u10_u6_n2837 ), .A3(_u10_u6_n2957 ), .ZN(_u10_u6_n2051 ) );
NOR2_X1 _u10_u6_U1100  ( .A1(_u10_u6_n2528 ), .A2(_u10_u6_n2051 ), .ZN(_u10_u6_n2605 ) );
NOR2_X1 _u10_u6_U1099  ( .A1(_u10_u6_n2605 ), .A2(_u10_u6_n2346 ), .ZN(_u10_u6_n3245 ) );
NOR2_X1 _u10_u6_U1098  ( .A1(_u10_u6_n2291 ), .A2(_u10_u6_n2062 ), .ZN(_u10_u6_n3246 ) );
NOR4_X1 _u10_u6_U1097  ( .A1(_u10_u6_n3243 ), .A2(_u10_u6_n3244 ), .A3(_u10_u6_n3245 ), .A4(_u10_u6_n3246 ), .ZN(_u10_u6_n3242 ) );
NAND2_X1 _u10_u6_U1096  ( .A1(_u10_u6_n3241 ), .A2(_u10_u6_n3242 ), .ZN(_u10_u6_n2311 ) );
OR3_X1 _u10_u6_U1095  ( .A1(_u10_u6_n1987 ), .A2(_u10_u6_n3240 ), .A3(_u10_u6_n2311 ), .ZN(_u10_u6_n3192 ) );
INV_X1 _u10_u6_U1094  ( .A(_u10_u6_n2886 ), .ZN(_u10_u6_n2720 ) );
NOR2_X1 _u10_u6_U1093  ( .A1(_u10_u6_n2004 ), .A2(_u10_u6_n2720 ), .ZN(_u10_u6_n2455 ) );
INV_X1 _u10_u6_U1092  ( .A(_u10_u6_n2488 ), .ZN(_u10_u6_n2938 ) );
AND3_X1 _u10_u6_U1091  ( .A1(_u10_u6_n2455 ), .A2(_u10_u6_n1859 ), .A3(_u10_u6_n2938 ), .ZN(_u10_u6_n3239 ) );
INV_X1 _u10_u6_U1090  ( .A(_u10_u6_n2633 ), .ZN(_u10_u6_n2937 ) );
NOR2_X1 _u10_u6_U1089  ( .A1(_u10_u6_n3239 ), .A2(_u10_u6_n2937 ), .ZN(_u10_u6_n3227 ) );
NOR2_X1 _u10_u6_U1088  ( .A1(_u10_u6_n1976 ), .A2(_u10_u6_n1969 ), .ZN(_u10_u6_n3237 ) );
NOR2_X1 _u10_u6_U1087  ( .A1(1'b0), .A2(_u10_u6_n2947 ), .ZN(_u10_u6_n3238 ));
NOR3_X1 _u10_u6_U1086  ( .A1(_u10_u6_n2476 ), .A2(_u10_u6_n3237 ), .A3(_u10_u6_n3238 ), .ZN(_u10_u6_n3235 ) );
NOR3_X1 _u10_u6_U1085  ( .A1(_u10_u6_n1813 ), .A2(_u10_u6_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_25 ), .ZN(_u10_u6_n3135 ) );
NAND2_X1 _u10_u6_U1084  ( .A1(_u10_u6_n3135 ), .A2(_u10_u6_n3236 ), .ZN(_u10_u6_n2573 ) );
NOR2_X1 _u10_u6_U1083  ( .A1(_u10_u6_n3235 ), .A2(_u10_u6_n2573 ), .ZN(_u10_u6_n3228 ) );
NOR2_X1 _u10_u6_U1082  ( .A1(_u10_u6_n2216 ), .A2(_u10_u6_n1868 ), .ZN(_u10_u6_n3233 ) );
INV_X1 _u10_u6_U1081  ( .A(_u10_u6_n2550 ), .ZN(_u10_u6_n2475 ) );
NOR3_X1 _u10_u6_U1080  ( .A1(_u10_u6_n2475 ), .A2(1'b0), .A3(_u10_u6_n1925 ),.ZN(_u10_u6_n3234 ) );
NOR3_X1 _u10_u6_U1079  ( .A1(_u10_u6_n3233 ), .A2(1'b0), .A3(_u10_u6_n3234 ),.ZN(_u10_u6_n3232 ) );
NOR2_X1 _u10_u6_U1078  ( .A1(_u10_u6_n3232 ), .A2(_u10_u6_n2037 ), .ZN(_u10_u6_n3229 ) );
NOR2_X1 _u10_u6_U1077  ( .A1(_u10_u6_n3231 ), .A2(_u10_u6_n2365 ), .ZN(_u10_u6_n3230 ) );
NOR4_X1 _u10_u6_U1076  ( .A1(_u10_u6_n3227 ), .A2(_u10_u6_n3228 ), .A3(_u10_u6_n3229 ), .A4(_u10_u6_n3230 ), .ZN(_u10_u6_n3205 ) );
NOR3_X1 _u10_u6_U1075  ( .A1(_u10_u6_n3226 ), .A2(_u10_u6_n2687 ), .A3(_u10_u6_n2145 ), .ZN(_u10_u6_n3217 ) );
NOR3_X1 _u10_u6_U1074  ( .A1(_u10_u6_n3225 ), .A2(1'b0), .A3(_u10_u6_n2587 ),.ZN(_u10_u6_n3218 ) );
NOR2_X1 _u10_u6_U1073  ( .A1(_u10_u6_n3159 ), .A2(1'b0), .ZN(_u10_u6_n3224 ));
NOR2_X1 _u10_u6_U1072  ( .A1(_u10_u6_n3224 ), .A2(_u10_u6_n2584 ), .ZN(_u10_u6_n3219 ) );
NAND2_X1 _u10_u6_U1071  ( .A1(_u10_u6_n3222 ), .A2(_u10_u6_n3223 ), .ZN(_u10_u6_n2048 ) );
INV_X1 _u10_u6_U1070  ( .A(_u10_u6_n2048 ), .ZN(_u10_u6_n2859 ) );
NOR2_X1 _u10_u6_U1069  ( .A1(_u10_u6_n2859 ), .A2(_u10_u6_n2054 ), .ZN(_u10_u6_n3221 ) );
NOR2_X1 _u10_u6_U1068  ( .A1(_u10_u6_n3221 ), .A2(_u10_u6_n2346 ), .ZN(_u10_u6_n3220 ) );
NOR4_X1 _u10_u6_U1067  ( .A1(_u10_u6_n3217 ), .A2(_u10_u6_n3218 ), .A3(_u10_u6_n3219 ), .A4(_u10_u6_n3220 ), .ZN(_u10_u6_n3206 ) );
NAND2_X1 _u10_u6_U1066  ( .A1(_u10_u6_n2377 ), .A2(_u10_u6_n2721 ), .ZN(_u10_u6_n3213 ) );
AND4_X1 _u10_u6_U1065  ( .A1(1'b0), .A2(_u10_u6_n2502 ), .A3(_u10_u6_n2972 ),.A4(_u10_u6_n3040 ), .ZN(_u10_u6_n2406 ) );
NAND2_X1 _u10_u6_U1064  ( .A1(_u10_u6_n2406 ), .A2(_u10_u6_n2979 ), .ZN(_u10_u6_n3214 ) );
NAND2_X1 _u10_u6_U1063  ( .A1(_u10_u6_n2630 ), .A2(_u10_u6_n3216 ), .ZN(_u10_u6_n2376 ) );
INV_X1 _u10_u6_U1062  ( .A(_u10_u6_n2376 ), .ZN(_u10_u6_n3108 ) );
NAND2_X1 _u10_u6_U1061  ( .A1(_u10_u6_n3108 ), .A2(_u10_u6_n2507 ), .ZN(_u10_u6_n3215 ) );
NOR2_X1 _u10_u6_U1060  ( .A1(_u10_u6_n2937 ), .A2(1'b0), .ZN(_u10_u6_n2649 ));
INV_X1 _u10_u6_U1059  ( .A(_u10_u6_n2253 ), .ZN(_u10_u6_n2971 ) );
NAND2_X1 _u10_u6_U1058  ( .A1(_u10_u6_n2649 ), .A2(_u10_u6_n2971 ), .ZN(_u10_u6_n2918 ) );
NAND4_X1 _u10_u6_U1057  ( .A1(_u10_u6_n3213 ), .A2(_u10_u6_n3214 ), .A3(_u10_u6_n3215 ), .A4(_u10_u6_n2918 ), .ZN(_u10_u6_n3208 ) );
NOR2_X1 _u10_u6_U1056  ( .A1(_u10_u6_n2000 ), .A2(_u10_u6_n2902 ), .ZN(_u10_u6_n3209 ) );
NOR2_X1 _u10_u6_U1055  ( .A1(_u10_u6_n3212 ), .A2(_u10_u6_n2475 ), .ZN(_u10_u6_n3210 ) );
INV_X1 _u10_u6_U1054  ( .A(_u10_u6_n2441 ), .ZN(_u10_u6_n3128 ) );
NOR2_X1 _u10_u6_U1053  ( .A1(_u10_u6_n2356 ), .A2(_u10_u6_n3128 ), .ZN(_u10_u6_n3211 ) );
NOR4_X1 _u10_u6_U1052  ( .A1(_u10_u6_n3208 ), .A2(_u10_u6_n3209 ), .A3(_u10_u6_n3210 ), .A4(_u10_u6_n3211 ), .ZN(_u10_u6_n3207 ) );
NAND3_X1 _u10_u6_U1051  ( .A1(_u10_u6_n3205 ), .A2(_u10_u6_n3206 ), .A3(_u10_u6_n3207 ), .ZN(_u10_u6_n2611 ) );
NOR2_X1 _u10_u6_U1050  ( .A1(_u10_u6_n2212 ), .A2(_u10_u6_n2216 ), .ZN(_u10_u6_n1937 ) );
NOR2_X1 _u10_u6_U1049  ( .A1(_u10_u6_n2533 ), .A2(_u10_u6_n2214 ), .ZN(_u10_u6_n2765 ) );
INV_X1 _u10_u6_U1048  ( .A(_u10_u6_n2005 ), .ZN(_u10_u6_n2111 ) );
AND2_X1 _u10_u6_U1047  ( .A1(_u10_u6_n2765 ), .A2(_u10_u6_n2111 ), .ZN(_u10_u6_n3201 ) );
INV_X1 _u10_u6_U1046  ( .A(_u10_u6_n3059 ), .ZN(_u10_u6_n3076 ) );
NAND2_X1 _u10_u6_U1045  ( .A1(_u10_u6_n3201 ), .A2(_u10_u6_n3076 ), .ZN(_u10_u6_n3204 ) );
NAND2_X1 _u10_u6_U1044  ( .A1(_u10_u6_n1937 ), .A2(_u10_u6_n3204 ), .ZN(_u10_u6_n3193 ) );
NAND2_X1 _u10_u6_U1043  ( .A1(_u10_u6_n2254 ), .A2(_u10_u6_n2212 ), .ZN(_u10_u6_n3203 ) );
NAND3_X1 _u10_u6_U1042  ( .A1(_u10_u6_n3203 ), .A2(_u10_u6_n2175 ), .A3(_u10_u6_n2649 ), .ZN(_u10_u6_n3194 ) );
NOR2_X1 _u10_u6_U1041  ( .A1(_u10_u6_n2985 ), .A2(1'b0), .ZN(_u10_u6_n1959 ));
NAND2_X1 _u10_u6_U1040  ( .A1(_u10_u6_n1959 ), .A2(_u10_u6_n3202 ), .ZN(_u10_u6_n2202 ) );
NAND4_X1 _u10_u6_U1039  ( .A1(_u10_u6_n3079 ), .A2(_u10_u6_n2621 ), .A3(_u10_u6_n2202 ), .A4(_u10_u6_n2798 ), .ZN(_u10_u6_n3200 ) );
NAND2_X1 _u10_u6_U1038  ( .A1(_u10_u6_n3201 ), .A2(_u10_u6_n2937 ), .ZN(_u10_u6_n2772 ) );
NAND2_X1 _u10_u6_U1037  ( .A1(_u10_u6_n3200 ), .A2(_u10_u6_n2772 ), .ZN(_u10_u6_n3195 ) );
NAND2_X1 _u10_u6_U1036  ( .A1(_u10_u6_n2765 ), .A2(_u10_u6_n1869 ), .ZN(_u10_u6_n3199 ) );
NAND2_X1 _u10_u6_U1035  ( .A1(_u10_u6_n2049 ), .A2(_u10_u6_n3199 ), .ZN(_u10_u6_n3057 ) );
NOR2_X1 _u10_u6_U1034  ( .A1(_u10_u6_n2495 ), .A2(_u10_u6_n3057 ), .ZN(_u10_u6_n3197 ) );
NOR2_X1 _u10_u6_U1033  ( .A1(_u10_u6_n2883 ), .A2(_u10_u6_n2485 ), .ZN(_u10_u6_n3198 ) );
NOR2_X1 _u10_u6_U1032  ( .A1(_u10_u6_n3197 ), .A2(_u10_u6_n3198 ), .ZN(_u10_u6_n3196 ) );
NAND4_X1 _u10_u6_U1031  ( .A1(_u10_u6_n3193 ), .A2(_u10_u6_n3194 ), .A3(_u10_u6_n3195 ), .A4(_u10_u6_n3196 ), .ZN(_u10_u6_n2887 ) );
NOR4_X1 _u10_u6_U1030  ( .A1(_u10_u6_n3191 ), .A2(_u10_u6_n3192 ), .A3(_u10_u6_n2611 ), .A4(_u10_u6_n2887 ), .ZN(_u10_u6_n3015 ) );
NAND3_X1 _u10_u6_U1029  ( .A1(_u10_u6_n3190 ), .A2(_u10_u6_n2049 ), .A3(_u10_u6_n2957 ), .ZN(_u10_u6_n2699 ) );
OR2_X1 _u10_u6_U1028  ( .A1(_u10_u6_n2699 ), .A2(_u10_u6_n1813 ), .ZN(_u10_u6_n3187 ) );
NAND3_X1 _u10_u6_U1027  ( .A1(_u10_u6_n2978 ), .A2(_u10_u6_n2405 ), .A3(1'b0), .ZN(_u10_u6_n3188 ) );
NAND4_X1 _u10_u6_U1026  ( .A1(_u10_u6_n3058 ), .A2(_u10_u6_n3187 ), .A3(_u10_u6_n3188 ), .A4(_u10_u6_n3189 ), .ZN(_u10_u6_n3186 ) );
NAND2_X1 _u10_u6_U1025  ( .A1(_u10_u6_n2063 ), .A2(_u10_u6_n3186 ), .ZN(_u10_u6_n3163 ) );
NAND2_X1 _u10_u6_U1024  ( .A1(_u10_u6_n3185 ), .A2(_u10_u6_n2329 ), .ZN(_u10_u6_n3164 ) );
NAND2_X1 _u10_u6_U1023  ( .A1(_u10_u6_n2689 ), .A2(_u10_u6_n2365 ), .ZN(_u10_u6_n2736 ) );
NOR2_X1 _u10_u6_U1022  ( .A1(_u10_u6_n2736 ), .A2(_u10_u6_n2488 ), .ZN(_u10_u6_n1855 ) );
INV_X1 _u10_u6_U1021  ( .A(_u10_u6_n1855 ), .ZN(_u10_u6_n3184 ) );
NOR2_X1 _u10_u6_U1020  ( .A1(_u10_u6_n2274 ), .A2(_u10_u6_n2359 ), .ZN(_u10_u6_n2952 ) );
NOR2_X1 _u10_u6_U1019  ( .A1(_u10_u6_n3184 ), .A2(_u10_u6_n2952 ), .ZN(_u10_u6_n2776 ) );
OR2_X1 _u10_u6_U1018  ( .A1(_u10_u6_n2852 ), .A2(_u10_u6_n2776 ), .ZN(_u10_u6_n3165 ) );
NAND2_X1 _u10_u6_U1017  ( .A1(_u10_u6_n3126 ), .A2(_u10_u6_n2915 ), .ZN(_u10_u6_n3065 ) );
NOR3_X1 _u10_u6_U1016  ( .A1(_u10_u6_n3065 ), .A2(1'b0), .A3(_u10_u6_n2632 ),.ZN(_u10_u6_n3182 ) );
NOR3_X1 _u10_u6_U1015  ( .A1(_u10_u6_n3182 ), .A2(_u10_u6_n3183 ), .A3(_u10_u6_n3108 ), .ZN(_u10_u6_n3181 ) );
NOR2_X1 _u10_u6_U1014  ( .A1(_u10_u6_n3181 ), .A2(_u10_u6_n3162 ), .ZN(_u10_u6_n3167 ) );
INV_X1 _u10_u6_U1013  ( .A(_u10_u6_n3180 ), .ZN(_u10_u6_n3140 ) );
NAND3_X1 _u10_u6_U1012  ( .A1(_u10_u6_n3140 ), .A2(_u10_u6_n2163 ), .A3(_u10_u6_n2092 ), .ZN(_u10_u6_n3175 ) );
NOR4_X1 _u10_u6_U1011  ( .A1(_u10_u6_n2411 ), .A2(_u10_u6_n2710 ), .A3(_u10_u6_n3141 ), .A4(_u10_u6_n3089 ), .ZN(_u10_u6_n3179 ) );
NOR2_X1 _u10_u6_U1010  ( .A1(1'b0), .A2(_u10_u6_n3179 ), .ZN(_u10_u6_n3177 ));
NOR2_X1 _u10_u6_U1009  ( .A1(_u10_u6_n1898 ), .A2(_u10_u6_n1847 ), .ZN(_u10_u6_n3178 ) );
NOR4_X1 _u10_u6_U1008  ( .A1(_u10_u6_n3175 ), .A2(_u10_u6_n3176 ), .A3(_u10_u6_n3177 ), .A4(_u10_u6_n3178 ), .ZN(_u10_u6_n3173 ) );
NAND2_X1 _u10_u6_U1007  ( .A1(_u10_u6_n3135 ), .A2(_u10_u6_n3174 ), .ZN(_u10_u6_n2159 ) );
NOR2_X1 _u10_u6_U1006  ( .A1(_u10_u6_n3173 ), .A2(_u10_u6_n2159 ), .ZN(_u10_u6_n3168 ) );
OR3_X1 _u10_u6_U1005  ( .A1(_u10_u6_n3172 ), .A2(1'b0), .A3(_u10_u6_n3126 ),.ZN(_u10_u6_n3171 ) );
NAND2_X1 _u10_u6_U1004  ( .A1(_u10_u6_n2600 ), .A2(_u10_u6_n3171 ), .ZN(_u10_u6_n3153 ) );
AND3_X1 _u10_u6_U1003  ( .A1(_u10_u6_n3153 ), .A2(_u10_u6_n2947 ), .A3(_u10_u6_n2579 ), .ZN(_u10_u6_n3170 ) );
NOR2_X1 _u10_u6_U1002  ( .A1(_u10_u6_n3170 ), .A2(_u10_u6_n2359 ), .ZN(_u10_u6_n3169 ) );
NOR3_X1 _u10_u6_U1001  ( .A1(_u10_u6_n3167 ), .A2(_u10_u6_n3168 ), .A3(_u10_u6_n3169 ), .ZN(_u10_u6_n3166 ) );
NAND4_X1 _u10_u6_U1000  ( .A1(_u10_u6_n3163 ), .A2(_u10_u6_n3164 ), .A3(_u10_u6_n3165 ), .A4(_u10_u6_n3166 ), .ZN(_u10_u6_n3130 ) );
NAND2_X1 _u10_u6_U999  ( .A1(_u10_u6_n2375 ), .A2(_u10_u6_n3162 ), .ZN(_u10_u6_n1923 ) );
NAND2_X1 _u10_u6_U998  ( .A1(_u10_u6_n3062 ), .A2(_u10_u6_n1923 ), .ZN(_u10_u6_n3154 ) );
NAND2_X1 _u10_u6_U997  ( .A1(_u10_u6_n2103 ), .A2(_u10_u6_n2509 ), .ZN(_u10_u6_n3161 ) );
NAND2_X1 _u10_u6_U996  ( .A1(_u10_u6_n2344 ), .A2(_u10_u6_n3161 ), .ZN(_u10_u6_n3160 ) );
NAND2_X1 _u10_u6_U995  ( .A1(_u10_u6_n3159 ), .A2(_u10_u6_n3160 ), .ZN(_u10_u6_n2635 ) );
AND3_X1 _u10_u6_U994  ( .A1(_u10_u6_n2549 ), .A2(_u10_u6_n2108 ), .A3(_u10_u6_n3126 ), .ZN(_u10_u6_n3093 ) );
NAND2_X1 _u10_u6_U993  ( .A1(_u10_u6_n3093 ), .A2(_u10_u6_n2941 ), .ZN(_u10_u6_n3158 ) );
NAND3_X1 _u10_u6_U992  ( .A1(_u10_u6_n3076 ), .A2(_u10_u6_n3066 ), .A3(_u10_u6_n3158 ), .ZN(_u10_u6_n3156 ) );
NAND2_X1 _u10_u6_U991  ( .A1(_u10_u6_n3156 ), .A2(_u10_u6_n3157 ), .ZN(_u10_u6_n3155 ) );
NAND3_X1 _u10_u6_U990  ( .A1(_u10_u6_n3154 ), .A2(_u10_u6_n2635 ), .A3(_u10_u6_n3155 ), .ZN(_u10_u6_n3131 ) );
INV_X1 _u10_u6_U989  ( .A(_u10_u6_n2594 ), .ZN(_u10_u6_n2846 ) );
NAND3_X1 _u10_u6_U988  ( .A1(_u10_u6_n2162 ), .A2(_u10_u6_n2082 ), .A3(_u10_u6_n2105 ), .ZN(_u10_u6_n2077 ) );
NAND4_X1 _u10_u6_U987  ( .A1(_u10_u6_n3153 ), .A2(_u10_u6_n1969 ), .A3(_u10_u6_n2846 ), .A4(_u10_u6_n2077 ), .ZN(_u10_u6_n3148 ) );
NAND2_X1 _u10_u6_U986  ( .A1(_u10_u6_n2838 ), .A2(_u10_u6_n3128 ), .ZN(_u10_u6_n3152 ) );
NAND2_X1 _u10_u6_U985  ( .A1(_u10_u6_n3152 ), .A2(_u10_u6_n2600 ), .ZN(_u10_u6_n3151 ) );
NAND2_X1 _u10_u6_U984  ( .A1(_u10_u6_n2282 ), .A2(_u10_u6_n3151 ), .ZN(_u10_u6_n2601 ) );
NOR4_X1 _u10_u6_U983  ( .A1(_u10_u6_n2885 ), .A2(_u10_u6_n2534 ), .A3(_u10_u6_n2214 ), .A4(_u10_u6_n3059 ), .ZN(_u10_u6_n3150 ) );
NOR2_X1 _u10_u6_U982  ( .A1(_u10_u6_n3150 ), .A2(_u10_u6_n2853 ), .ZN(_u10_u6_n3149 ) );
NOR4_X1 _u10_u6_U981  ( .A1(_u10_u6_n3148 ), .A2(_u10_u6_n2601 ), .A3(_u10_u6_n3149 ), .A4(_u10_u6_n1975 ), .ZN(_u10_u6_n3146 ) );
NAND3_X1 _u10_u6_U980  ( .A1(_u10_SYNOPSYS_UNCONNECTED_28 ), .A2(_u10_SYNOPSYS_UNCONNECTED_24 ), .A3(_u10_u6_n3147 ), .ZN(_u10_u6_n2071 ) );
NOR2_X1 _u10_u6_U979  ( .A1(_u10_u6_n3146 ), .A2(_u10_u6_n2071 ), .ZN(_u10_u6_n3132 ) );
NOR2_X1 _u10_u6_U978  ( .A1(1'b0), .A2(_u10_u6_n1847 ), .ZN(_u10_u6_n3143 ));
INV_X1 _u10_u6_U977  ( .A(_u10_u6_n3145 ), .ZN(_u10_u6_n3144 ) );
NOR2_X1 _u10_u6_U976  ( .A1(_u10_u6_n3143 ), .A2(_u10_u6_n3144 ), .ZN(_u10_u6_n3142 ) );
NOR2_X1 _u10_u6_U975  ( .A1(1'b0), .A2(_u10_u6_n3142 ), .ZN(_u10_u6_n3137 ));
NAND2_X1 _u10_u6_U974  ( .A1(_u10_u6_n2549 ), .A2(_u10_u6_n3141 ), .ZN(_u10_u6_n3138 ) );
NAND2_X1 _u10_u6_U973  ( .A1(_u10_u6_n1896 ), .A2(_u10_u6_n3140 ), .ZN(_u10_u6_n2544 ) );
NAND2_X1 _u10_u6_U972  ( .A1(_u10_u6_n2089 ), .A2(_u10_u6_n2544 ), .ZN(_u10_u6_n3139 ) );
NAND2_X1 _u10_u6_U971  ( .A1(_u10_u6_n3138 ), .A2(_u10_u6_n3139 ), .ZN(_u10_u6_n2795 ) );
NOR4_X1 _u10_u6_U970  ( .A1(_u10_u6_n2300 ), .A2(_u10_u6_n3137 ), .A3(_u10_u6_n2304 ), .A4(_u10_u6_n2795 ), .ZN(_u10_u6_n3134 ) );
NAND2_X1 _u10_u6_U969  ( .A1(_u10_u6_n3135 ), .A2(_u10_u6_n3136 ), .ZN(_u10_u6_n2085 ) );
NOR2_X1 _u10_u6_U968  ( .A1(_u10_u6_n3134 ), .A2(_u10_u6_n2085 ), .ZN(_u10_u6_n3133 ) );
NOR4_X1 _u10_u6_U967  ( .A1(_u10_u6_n3130 ), .A2(_u10_u6_n3131 ), .A3(_u10_u6_n3132 ), .A4(_u10_u6_n3133 ), .ZN(_u10_u6_n3016 ) );
INV_X1 _u10_u6_U966  ( .A(_u10_u6_n2686 ), .ZN(_u10_u6_n2278 ) );
NAND4_X1 _u10_u6_U965  ( .A1(_u10_u6_n2105 ), .A2(_u10_u6_n2278 ), .A3(_u10_u6_n3129 ), .A4(_u10_u6_n2600 ), .ZN(_u10_u6_n2437 ) );
NAND2_X1 _u10_u6_U964  ( .A1(_u10_u6_n3128 ), .A2(_u10_u6_n2437 ), .ZN(_u10_u6_n3127 ) );
NAND2_X1 _u10_u6_U963  ( .A1(_u10_u6_n2815 ), .A2(_u10_u6_n3127 ), .ZN(_u10_u6_n3098 ) );
INV_X1 _u10_u6_U962  ( .A(_u10_u6_n2573 ), .ZN(_u10_u6_n1967 ) );
NAND2_X1 _u10_u6_U961  ( .A1(_u10_u6_n3126 ), .A2(_u10_u6_n2078 ), .ZN(_u10_u6_n3123 ) );
NAND2_X1 _u10_u6_U960  ( .A1(_u10_u6_n3076 ), .A2(_u10_u6_n1925 ), .ZN(_u10_u6_n3125 ) );
NAND2_X1 _u10_u6_U959  ( .A1(_u10_u6_n2669 ), .A2(_u10_u6_n3125 ), .ZN(_u10_u6_n3124 ) );
NAND4_X1 _u10_u6_U958  ( .A1(_u10_u6_n3122 ), .A2(_u10_u6_n3123 ), .A3(_u10_u6_n3124 ), .A4(_u10_u6_n2579 ), .ZN(_u10_u6_n3121 ) );
NAND2_X1 _u10_u6_U957  ( .A1(_u10_u6_n3121 ), .A2(_u10_u6_n2874 ), .ZN(_u10_u6_n3120 ) );
NAND2_X1 _u10_u6_U956  ( .A1(_u10_u6_n2382 ), .A2(_u10_u6_n3120 ), .ZN(_u10_u6_n3119 ) );
NAND2_X1 _u10_u6_U955  ( .A1(_u10_u6_n1967 ), .A2(_u10_u6_n3119 ), .ZN(_u10_u6_n3099 ) );
NAND2_X1 _u10_u6_U954  ( .A1(_u10_u6_n3118 ), .A2(_u10_u6_n3001 ), .ZN(_u10_u6_n3117 ) );
NAND2_X1 _u10_u6_U953  ( .A1(_u10_u6_n2446 ), .A2(_u10_u6_n3117 ), .ZN(_u10_u6_n3116 ) );
NAND2_X1 _u10_u6_U952  ( .A1(_u10_u6_n2445 ), .A2(_u10_u6_n3116 ), .ZN(_u10_u6_n3100 ) );
OR2_X1 _u10_u6_U951  ( .A1(_u10_u6_n3115 ), .A2(_u10_u6_n2687 ), .ZN(_u10_u6_n3114 ) );
AND3_X1 _u10_u6_U950  ( .A1(_u10_u6_n2061 ), .A2(_u10_u6_n2166 ), .A3(_u10_u6_n3114 ), .ZN(_u10_u6_n3045 ) );
NOR2_X1 _u10_u6_U949  ( .A1(1'b0), .A2(_u10_u6_n3045 ), .ZN(_u10_u6_n3113 ));
NOR2_X1 _u10_u6_U948  ( .A1(_u10_u6_n3113 ), .A2(1'b0), .ZN(_u10_u6_n3112 ));
NOR2_X1 _u10_u6_U947  ( .A1(_u10_u6_n3112 ), .A2(_u10_u6_n2356 ), .ZN(_u10_u6_n3102 ) );
NAND2_X1 _u10_u6_U946  ( .A1(_u10_u6_n2571 ), .A2(_u10_u6_n2165 ), .ZN(_u10_u6_n3078 ) );
NAND2_X1 _u10_u6_U945  ( .A1(_u10_u6_n2365 ), .A2(_u10_u6_n3078 ), .ZN(_u10_u6_n2241 ) );
NOR2_X1 _u10_u6_U944  ( .A1(_u10_u6_n2377 ), .A2(_u10_u6_n2241 ), .ZN(_u10_u6_n3111 ) );
NOR2_X1 _u10_u6_U943  ( .A1(_u10_u6_n3111 ), .A2(_u10_u6_n1869 ), .ZN(_u10_u6_n3103 ) );
NOR2_X1 _u10_u6_U942  ( .A1(_u10_u6_n2999 ), .A2(_u10_u6_n2977 ), .ZN(_u10_u6_n3061 ) );
NOR2_X1 _u10_u6_U941  ( .A1(_u10_u6_n3061 ), .A2(_u10_u6_n2367 ), .ZN(_u10_u6_n3106 ) );
NAND2_X1 _u10_u6_U940  ( .A1(_u10_u6_n2977 ), .A2(_u10_u6_n3000 ), .ZN(_u10_u6_n3110 ) );
NAND2_X1 _u10_u6_U939  ( .A1(_u10_u6_n3109 ), .A2(_u10_u6_n3110 ), .ZN(_u10_u6_n1924 ) );
AND2_X1 _u10_u6_U938  ( .A1(_u10_u6_n1924 ), .A2(_u10_u6_n3108 ), .ZN(_u10_u6_n3107 ) );
NOR2_X1 _u10_u6_U937  ( .A1(_u10_u6_n3106 ), .A2(_u10_u6_n3107 ), .ZN(_u10_u6_n3105 ) );
NOR2_X1 _u10_u6_U936  ( .A1(_u10_u6_n3105 ), .A2(_u10_u6_n2008 ), .ZN(_u10_u6_n3104 ) );
NOR3_X1 _u10_u6_U935  ( .A1(_u10_u6_n3102 ), .A2(_u10_u6_n3103 ), .A3(_u10_u6_n3104 ), .ZN(_u10_u6_n3101 ) );
NAND4_X1 _u10_u6_U934  ( .A1(_u10_u6_n3098 ), .A2(_u10_u6_n3099 ), .A3(_u10_u6_n3100 ), .A4(_u10_u6_n3101 ), .ZN(_u10_u6_n3071 ) );
NOR2_X1 _u10_u6_U933  ( .A1(_u10_u6_n1926 ), .A2(_u10_u6_n2980 ), .ZN(_u10_u6_n2218 ) );
INV_X1 _u10_u6_U932  ( .A(_u10_u6_n2721 ), .ZN(_u10_u6_n2910 ) );
NAND2_X1 _u10_u6_U931  ( .A1(_u10_u6_n2910 ), .A2(_u10_u6_n1869 ), .ZN(_u10_u6_n2779 ) );
NAND2_X1 _u10_u6_U930  ( .A1(_u10_u6_n2218 ), .A2(_u10_u6_n2779 ), .ZN(_u10_u6_n3081 ) );
NAND2_X1 _u10_u6_U929  ( .A1(_u10_u6_n1922 ), .A2(_u10_u6_n1864 ), .ZN(_u10_u6_n2179 ) );
NOR3_X1 _u10_u6_U928  ( .A1(_u10_u6_n1961 ), .A2(_u10_u6_n1918 ), .A3(_u10_u6_n2179 ), .ZN(_u10_u6_n2693 ) );
NAND2_X1 _u10_u6_U927  ( .A1(_u10_u6_n3097 ), .A2(_u10_u6_n1924 ), .ZN(_u10_u6_n3096 ) );
NAND2_X1 _u10_u6_U926  ( .A1(_u10_u6_n1984 ), .A2(_u10_u6_n3096 ), .ZN(_u10_u6_n2506 ) );
INV_X1 _u10_u6_U925  ( .A(_u10_u6_n2506 ), .ZN(_u10_u6_n2366 ) );
NAND2_X1 _u10_u6_U924  ( .A1(_u10_u6_n2366 ), .A2(_u10_u6_n2375 ), .ZN(_u10_u6_n2236 ) );
NAND2_X1 _u10_u6_U923  ( .A1(_u10_u6_n2693 ), .A2(_u10_u6_n2236 ), .ZN(_u10_u6_n3082 ) );
NAND2_X1 _u10_u6_U922  ( .A1(1'b0), .A2(_u10_u6_n2126 ), .ZN(_u10_u6_n3095 ));
NAND2_X1 _u10_u6_U921  ( .A1(_u10_u6_n1956 ), .A2(_u10_u6_n3095 ), .ZN(_u10_u6_n2907 ) );
OR2_X1 _u10_u6_U920  ( .A1(_u10_u6_n2902 ), .A2(_u10_u6_n2907 ), .ZN(_u10_u6_n3085 ) );
NAND2_X1 _u10_u6_U919  ( .A1(_u10_u6_n2256 ), .A2(_u10_u6_n2113 ), .ZN(_u10_u6_n3094 ) );
NAND2_X1 _u10_u6_U918  ( .A1(_u10_u6_n2688 ), .A2(_u10_u6_n3094 ), .ZN(_u10_u6_n3092 ) );
NAND2_X1 _u10_u6_U917  ( .A1(_u10_u6_n3093 ), .A2(_u10_u6_n3092 ), .ZN(_u10_u6_n3086 ) );
INV_X1 _u10_u6_U916  ( .A(_u10_u6_n2159 ), .ZN(_u10_u6_n1894 ) );
NAND2_X1 _u10_u6_U915  ( .A1(_u10_u6_n3067 ), .A2(_u10_u6_n1894 ), .ZN(_u10_u6_n3091 ) );
INV_X1 _u10_u6_U914  ( .A(_u10_u6_n3092 ), .ZN(_u10_u6_n2234 ) );
NAND3_X1 _u10_u6_U913  ( .A1(_u10_u6_n3091 ), .A2(_u10_u6_n2126 ), .A3(_u10_u6_n2234 ), .ZN(_u10_u6_n3090 ) );
NAND2_X1 _u10_u6_U912  ( .A1(1'b0), .A2(_u10_u6_n3090 ), .ZN(_u10_u6_n3087 ));
NAND3_X1 _u10_u6_U911  ( .A1(_u10_u6_n2329 ), .A2(_u10_u6_n3089 ), .A3(_u10_u6_n2549 ), .ZN(_u10_u6_n3088 ) );
NAND4_X1 _u10_u6_U910  ( .A1(_u10_u6_n3085 ), .A2(_u10_u6_n3086 ), .A3(_u10_u6_n3087 ), .A4(_u10_u6_n3088 ), .ZN(_u10_u6_n3084 ) );
NAND2_X1 _u10_u6_U909  ( .A1(_u10_u6_n3084 ), .A2(_u10_u6_n2803 ), .ZN(_u10_u6_n3083 ) );
NAND3_X1 _u10_u6_U908  ( .A1(_u10_u6_n3081 ), .A2(_u10_u6_n3082 ), .A3(_u10_u6_n3083 ), .ZN(_u10_u6_n3072 ) );
INV_X1 _u10_u6_U907  ( .A(_u10_u6_n2689 ), .ZN(_u10_u6_n1955 ) );
NOR3_X1 _u10_u6_U906  ( .A1(_u10_u6_n1955 ), .A2(_u10_u6_n2813 ), .A3(_u10_u6_n2488 ), .ZN(_u10_u6_n3080 ) );
NOR2_X1 _u10_u6_U905  ( .A1(_u10_u6_n3080 ), .A2(_u10_u6_n2485 ), .ZN(_u10_u6_n3073 ) );
NAND3_X1 _u10_u6_U904  ( .A1(_u10_u6_n2621 ), .A2(_u10_u6_n2202 ), .A3(_u10_u6_n3079 ), .ZN(_u10_u6_n2110 ) );
NOR2_X1 _u10_u6_U903  ( .A1(_u10_u6_n2110 ), .A2(_u10_u6_n2218 ), .ZN(_u10_u6_n2775 ) );
INV_X1 _u10_u6_U902  ( .A(_u10_u6_n2775 ), .ZN(_u10_u6_n3024 ) );
INV_X1 _u10_u6_U901  ( .A(_u10_u6_n3078 ), .ZN(_u10_u6_n2133 ) );
INV_X1 _u10_u6_U900  ( .A(_u10_u6_n2007 ), .ZN(_u10_u6_n2358 ) );
NAND2_X1 _u10_u6_U899  ( .A1(_u10_u6_n2358 ), .A2(_u10_u6_n2886 ), .ZN(_u10_u6_n2240 ) );
INV_X1 _u10_u6_U898  ( .A(_u10_u6_n2240 ), .ZN(_u10_u6_n2083 ) );
NOR3_X1 _u10_u6_U897  ( .A1(_u10_u6_n2952 ), .A2(_u10_u6_n2004 ), .A3(_u10_u6_n1891 ), .ZN(_u10_u6_n3077 ) );
NAND3_X1 _u10_u6_U896  ( .A1(_u10_u6_n2083 ), .A2(_u10_u6_n2938 ), .A3(_u10_u6_n3077 ), .ZN(_u10_u6_n1886 ) );
NOR3_X1 _u10_u6_U895  ( .A1(_u10_u6_n3024 ), .A2(_u10_u6_n2133 ), .A3(_u10_u6_n1886 ), .ZN(_u10_u6_n3075 ) );
NOR2_X1 _u10_u6_U894  ( .A1(_u10_u6_n3075 ), .A2(_u10_u6_n3076 ), .ZN(_u10_u6_n3074 ) );
NOR4_X1 _u10_u6_U893  ( .A1(_u10_u6_n3071 ), .A2(_u10_u6_n3072 ), .A3(_u10_u6_n3073 ), .A4(_u10_u6_n3074 ), .ZN(_u10_u6_n3017 ) );
INV_X1 _u10_u6_U892  ( .A(_u10_u6_n3065 ), .ZN(_u10_u6_n3043 ) );
NAND2_X1 _u10_u6_U891  ( .A1(_u10_u6_n3043 ), .A2(_u10_u6_n2106 ), .ZN(_u10_u6_n3070 ) );
NAND2_X1 _u10_u6_U890  ( .A1(_u10_u6_n3070 ), .A2(_u10_u6_n2038 ), .ZN(_u10_u6_n3068 ) );
NAND2_X1 _u10_u6_U889  ( .A1(_u10_u6_n2344 ), .A2(_u10_u6_n2584 ), .ZN(_u10_u6_n3069 ) );
NAND3_X1 _u10_u6_U888  ( .A1(_u10_u6_n3068 ), .A2(_u10_u6_n1930 ), .A3(_u10_u6_n3069 ), .ZN(_u10_u6_n3047 ) );
NAND2_X1 _u10_u6_U887  ( .A1(_u10_u6_n2835 ), .A2(_u10_u6_n2466 ), .ZN(_u10_u6_n2130 ) );
INV_X1 _u10_u6_U886  ( .A(_u10_u6_n2130 ), .ZN(_u10_u6_n2168 ) );
NAND3_X1 _u10_u6_U885  ( .A1(_u10_u6_n3067 ), .A2(_u10_u6_n2329 ), .A3(_u10_u6_n2168 ), .ZN(_u10_u6_n2665 ) );
NAND3_X1 _u10_u6_U884  ( .A1(_u10_u6_n3065 ), .A2(_u10_u6_n3066 ), .A3(_u10_u6_n2342 ), .ZN(_u10_u6_n3064 ) );
NAND3_X1 _u10_u6_U883  ( .A1(_u10_u6_n3064 ), .A2(_u10_u6_n2175 ), .A3(_u10_u6_n2987 ), .ZN(_u10_u6_n3048 ) );
NOR3_X1 _u10_u6_U882  ( .A1(_u10_u6_n1849 ), .A2(1'b0), .A3(_u10_u6_n3063 ),.ZN(_u10_u6_n3050 ) );
NOR3_X1 _u10_u6_U881  ( .A1(_u10_u6_n2406 ), .A2(1'b0), .A3(_u10_u6_n3062 ),.ZN(_u10_u6_n3060 ) );
NOR3_X1 _u10_u6_U880  ( .A1(_u10_u6_n3060 ), .A2(1'b0), .A3(_u10_u6_n3061 ),.ZN(_u10_u6_n3051 ) );
NAND2_X1 _u10_u6_U879  ( .A1(_u10_u6_n3059 ), .A2(_u10_u6_n2049 ), .ZN(_u10_u6_n3056 ) );
NAND3_X1 _u10_u6_U878  ( .A1(_u10_u6_n3056 ), .A2(_u10_u6_n3057 ), .A3(_u10_u6_n3058 ), .ZN(_u10_u6_n3054 ) );
NOR4_X1 _u10_u6_U877  ( .A1(_u10_u6_n3054 ), .A2(_u10_u6_n3055 ), .A3(_u10_u6_n2055 ), .A4(_u10_u6_n2056 ), .ZN(_u10_u6_n3053 ) );
NOR3_X1 _u10_u6_U876  ( .A1(_u10_u6_n2346 ), .A2(1'b0), .A3(_u10_u6_n3053 ),.ZN(_u10_u6_n3052 ) );
NOR3_X1 _u10_u6_U875  ( .A1(_u10_u6_n3050 ), .A2(_u10_u6_n3051 ), .A3(_u10_u6_n3052 ), .ZN(_u10_u6_n3049 ) );
NAND4_X1 _u10_u6_U874  ( .A1(_u10_u6_n3047 ), .A2(_u10_u6_n2665 ), .A3(_u10_u6_n3048 ), .A4(_u10_u6_n3049 ), .ZN(_u10_u6_n3019 ) );
NAND2_X1 _u10_u6_U873  ( .A1(_u10_u6_n2056 ), .A2(_u10_u6_n2019 ), .ZN(_u10_u6_n3046 ) );
NAND2_X1 _u10_u6_U872  ( .A1(_u10_u6_n3045 ), .A2(_u10_u6_n3046 ), .ZN(_u10_u6_n3044 ) );
NAND2_X1 _u10_u6_U871  ( .A1(_u10_u6_n3044 ), .A2(_u10_u6_n2165 ), .ZN(_u10_u6_n3028 ) );
OR2_X1 _u10_u6_U870  ( .A1(_u10_u6_n2179 ), .A2(_u10_u6_n1961 ), .ZN(_u10_u6_n3037 ) );
NAND2_X1 _u10_u6_U869  ( .A1(_u10_u6_n3043 ), .A2(_u10_u6_n2336 ), .ZN(_u10_u6_n3042 ) );
NAND2_X1 _u10_u6_U868  ( .A1(_u10_u6_n3042 ), .A2(_u10_u6_n3006 ), .ZN(_u10_u6_n3041 ) );
NAND2_X1 _u10_u6_U867  ( .A1(_u10_u6_n3040 ), .A2(_u10_u6_n3041 ), .ZN(_u10_u6_n3026 ) );
NAND4_X1 _u10_u6_U866  ( .A1(_u10_u6_n3026 ), .A2(_u10_u6_n2520 ), .A3(_u10_u6_n1962 ), .A4(_u10_u6_n1864 ), .ZN(_u10_u6_n3039 ) );
NAND2_X1 _u10_u6_U865  ( .A1(_u10_u6_n3039 ), .A2(_u10_u6_n1922 ), .ZN(_u10_u6_n3038 ) );
NAND2_X1 _u10_u6_U864  ( .A1(_u10_u6_n3037 ), .A2(_u10_u6_n3038 ), .ZN(_u10_u6_n3035 ) );
NAND2_X1 _u10_u6_U863  ( .A1(_u10_u6_n2985 ), .A2(_u10_u6_n3036 ), .ZN(_u10_u6_n2432 ) );
NAND2_X1 _u10_u6_U862  ( .A1(_u10_u6_n3035 ), .A2(_u10_u6_n2432 ), .ZN(_u10_u6_n3029 ) );
INV_X1 _u10_u6_U861  ( .A(_u10_u6_n3034 ), .ZN(_u10_u6_n2777 ) );
INV_X1 _u10_u6_U860  ( .A(_u10_u6_n2772 ), .ZN(_u10_u6_n3032 ) );
NAND2_X1 _u10_u6_U859  ( .A1(_u10_u6_n1982 ), .A2(_u10_u6_n2978 ), .ZN(_u10_u6_n3033 ) );
NAND2_X1 _u10_u6_U858  ( .A1(_u10_u6_n3032 ), .A2(_u10_u6_n3033 ), .ZN(_u10_u6_n3031 ) );
NAND2_X1 _u10_u6_U857  ( .A1(_u10_u6_n2777 ), .A2(_u10_u6_n3031 ), .ZN(_u10_u6_n3030 ) );
NAND3_X1 _u10_u6_U856  ( .A1(_u10_u6_n3028 ), .A2(_u10_u6_n3029 ), .A3(_u10_u6_n3030 ), .ZN(_u10_u6_n3020 ) );
NOR3_X1 _u10_u6_U855  ( .A1(_u10_u6_n2179 ), .A2(1'b0), .A3(_u10_u6_n2375 ),.ZN(_u10_u6_n3027 ) );
NOR2_X1 _u10_u6_U854  ( .A1(_u10_u6_n3027 ), .A2(_u10_u6_n2177 ), .ZN(_u10_u6_n3025 ) );
NOR2_X1 _u10_u6_U853  ( .A1(_u10_u6_n3025 ), .A2(_u10_u6_n3026 ), .ZN(_u10_u6_n3021 ) );
NOR2_X1 _u10_u6_U852  ( .A1(_u10_u6_n2256 ), .A2(_u10_u6_n3024 ), .ZN(_u10_u6_n3023 ) );
NOR2_X1 _u10_u6_U851  ( .A1(_u10_u6_n3023 ), .A2(_u10_u6_n1868 ), .ZN(_u10_u6_n3022 ) );
NOR4_X1 _u10_u6_U850  ( .A1(_u10_u6_n3019 ), .A2(_u10_u6_n3020 ), .A3(_u10_u6_n3021 ), .A4(_u10_u6_n3022 ), .ZN(_u10_u6_n3018 ) );
NAND4_X1 _u10_u6_U849  ( .A1(_u10_u6_n3015 ), .A2(_u10_u6_n3016 ), .A3(_u10_u6_n3017 ), .A4(_u10_u6_n3018 ), .ZN(_u10_u6_n2958 ) );
NOR2_X1 _u10_u6_U848  ( .A1(1'b0), .A2(_u10_u6_n2573 ), .ZN(_u10_u6_n3011 ));
NOR2_X1 _u10_u6_U847  ( .A1(1'b0), .A2(_u10_u6_n2359 ), .ZN(_u10_u6_n3012 ));
NOR2_X1 _u10_u6_U846  ( .A1(1'b0), .A2(_u10_u6_n1859 ), .ZN(_u10_u6_n3013 ));
NOR2_X1 _u10_u6_U845  ( .A1(1'b0), .A2(_u10_u6_n1836 ), .ZN(_u10_u6_n3014 ));
NOR4_X1 _u10_u6_U844  ( .A1(_u10_u6_n3011 ), .A2(_u10_u6_n3012 ), .A3(_u10_u6_n3013 ), .A4(_u10_u6_n3014 ), .ZN(_u10_u6_n2959 ) );
NOR2_X1 _u10_u6_U843  ( .A1(1'b0), .A2(_u10_u6_n2025 ), .ZN(_u10_u6_n3007 ));
NOR2_X1 _u10_u6_U842  ( .A1(1'b0), .A2(_u10_u6_n2085 ), .ZN(_u10_u6_n3008 ));
NOR2_X1 _u10_u6_U841  ( .A1(1'b0), .A2(_u10_u6_n2607 ), .ZN(_u10_u6_n3009 ));
NOR2_X1 _u10_u6_U840  ( .A1(1'b0), .A2(_u10_u6_n2071 ), .ZN(_u10_u6_n3010 ));
NOR4_X1 _u10_u6_U839  ( .A1(_u10_u6_n3007 ), .A2(_u10_u6_n3008 ), .A3(_u10_u6_n3009 ), .A4(_u10_u6_n3010 ), .ZN(_u10_u6_n2960 ) );
NAND2_X1 _u10_u6_U838  ( .A1(_u10_u6_n1894 ), .A2(_u10_u6_n2466 ), .ZN(_u10_u6_n3002 ) );
NAND2_X1 _u10_u6_U837  ( .A1(_u10_u6_n2830 ), .A2(_u10_u6_n2600 ), .ZN(_u10_u6_n3003 ) );
NAND2_X1 _u10_u6_U836  ( .A1(_u10_u6_n1960 ), .A2(_u10_u6_n2431 ), .ZN(_u10_u6_n3004 ) );
NAND2_X1 _u10_u6_U835  ( .A1(_u10_u6_n2002 ), .A2(_u10_u6_n3006 ), .ZN(_u10_u6_n3005 ) );
NAND4_X1 _u10_u6_U834  ( .A1(_u10_u6_n3002 ), .A2(_u10_u6_n3003 ), .A3(_u10_u6_n3004 ), .A4(_u10_u6_n3005 ), .ZN(_u10_u6_n2992 ) );
NAND2_X1 _u10_u6_U833  ( .A1(_u10_u6_n2461 ), .A2(_u10_u6_n3001 ), .ZN(_u10_u6_n2997 ) );
NAND2_X1 _u10_u6_U832  ( .A1(_u10_u6_n2999 ), .A2(_u10_u6_n3000 ), .ZN(_u10_u6_n2998 ) );
NAND2_X1 _u10_u6_U831  ( .A1(_u10_u6_n2997 ), .A2(_u10_u6_n2998 ), .ZN(_u10_u6_n2993 ) );
NOR2_X1 _u10_u6_U830  ( .A1(_u10_SYNOPSYS_UNCONNECTED_24 ), .A2(_u10_u6_n2996 ), .ZN(_u10_u6_n2995 ) );
NOR2_X1 _u10_u6_U829  ( .A1(_u10_u6_n2995 ), .A2(_u10_u6_n2126 ), .ZN(_u10_u6_n2994 ) );
NOR4_X1 _u10_u6_U828  ( .A1(_u10_u6_n2992 ), .A2(_u10_u6_n2993 ), .A3(next_ch), .A4(_u10_u6_n2994 ), .ZN(_u10_u6_n2961 ) );
NAND2_X1 _u10_u6_U827  ( .A1(_u10_u6_n2445 ), .A2(_u10_u6_n2803 ), .ZN(_u10_u6_n2988 ) );
OR2_X1 _u10_u6_U826  ( .A1(_u10_u6_n2584 ), .A2(1'b0), .ZN(_u10_u6_n2989 ));
NAND2_X1 _u10_u6_U825  ( .A1(_u10_u6_n2709 ), .A2(_u10_u6_n2080 ), .ZN(_u10_u6_n2990 ) );
NAND2_X1 _u10_u6_U824  ( .A1(_u10_u6_n2183 ), .A2(_u10_u6_n2166 ), .ZN(_u10_u6_n2991 ) );
NAND4_X1 _u10_u6_U823  ( .A1(_u10_u6_n2988 ), .A2(_u10_u6_n2989 ), .A3(_u10_u6_n2990 ), .A4(_u10_u6_n2991 ), .ZN(_u10_u6_n2963 ) );
NAND2_X1 _u10_u6_U822  ( .A1(_u10_u6_n2987 ), .A2(_u10_u6_n1930 ), .ZN(_u10_u6_n2981 ) );
NAND2_X1 _u10_u6_U821  ( .A1(_u10_u6_n2986 ), .A2(_u10_u6_n2038 ), .ZN(_u10_u6_n2982 ) );
OR2_X1 _u10_u6_U820  ( .A1(_u10_u6_n2985 ), .A2(1'b0), .ZN(_u10_u6_n2983 ));
NAND2_X1 _u10_u6_U819  ( .A1(_u10_u6_n2169 ), .A2(_u10_u6_n2113 ), .ZN(_u10_u6_n2984 ) );
NAND4_X1 _u10_u6_U818  ( .A1(_u10_u6_n2981 ), .A2(_u10_u6_n2982 ), .A3(_u10_u6_n2983 ), .A4(_u10_u6_n2984 ), .ZN(_u10_u6_n2964 ) );
NAND2_X1 _u10_u6_U817  ( .A1(_u10_u6_n2509 ), .A2(_u10_u6_n1864 ), .ZN(_u10_u6_n2973 ) );
INV_X1 _u10_u6_U816  ( .A(_u10_u6_n2980 ), .ZN(_u10_u6_n1861 ) );
NAND2_X1 _u10_u6_U815  ( .A1(_u10_u6_n1861 ), .A2(_u10_u6_n1922 ), .ZN(_u10_u6_n2974 ) );
NAND2_X1 _u10_u6_U814  ( .A1(_u10_u6_n2979 ), .A2(_u10_u6_n2405 ), .ZN(_u10_u6_n2975 ) );
NAND2_X1 _u10_u6_U813  ( .A1(_u10_u6_n2977 ), .A2(_u10_u6_n2978 ), .ZN(_u10_u6_n2976 ) );
NAND4_X1 _u10_u6_U812  ( .A1(_u10_u6_n2973 ), .A2(_u10_u6_n2974 ), .A3(_u10_u6_n2975 ), .A4(_u10_u6_n2976 ), .ZN(_u10_u6_n2965 ) );
NAND2_X1 _u10_u6_U811  ( .A1(_u10_u6_n2507 ), .A2(_u10_u6_n2972 ), .ZN(_u10_u6_n2967 ) );
NAND2_X1 _u10_u6_U810  ( .A1(_u10_u6_n2043 ), .A2(_u10_u6_n1965 ), .ZN(_u10_u6_n2968 ) );
NAND2_X1 _u10_u6_U809  ( .A1(_u10_u6_n2063 ), .A2(_u10_u6_n1853 ), .ZN(_u10_u6_n2969 ) );
NAND2_X1 _u10_u6_U808  ( .A1(_u10_u6_n2971 ), .A2(_u10_u6_n2175 ), .ZN(_u10_u6_n2970 ) );
NAND4_X1 _u10_u6_U807  ( .A1(_u10_u6_n2967 ), .A2(_u10_u6_n2968 ), .A3(_u10_u6_n2969 ), .A4(_u10_u6_n2970 ), .ZN(_u10_u6_n2966 ) );
NOR4_X1 _u10_u6_U806  ( .A1(_u10_u6_n2963 ), .A2(_u10_u6_n2964 ), .A3(_u10_u6_n2965 ), .A4(_u10_u6_n2966 ), .ZN(_u10_u6_n2962 ) );
AND4_X1 _u10_u6_U805  ( .A1(_u10_u6_n2959 ), .A2(_u10_u6_n2960 ), .A3(_u10_u6_n2961 ), .A4(_u10_u6_n2962 ), .ZN(_u10_u6_n1819 ) );
MUX2_X1 _u10_u6_U804  ( .A(_u10_u6_n2958 ), .B(_u10_SYNOPSYS_UNCONNECTED_28 ), .S(_u10_u6_n1819 ), .Z(_u10_u6_n1808 ) );
NOR2_X1 _u10_u6_U803  ( .A1(_u10_u6_n2531 ), .A2(_u10_u6_n2607 ), .ZN(_u10_u6_n1911 ) );
NAND2_X1 _u10_u6_U802  ( .A1(_u10_u6_n1911 ), .A2(_u10_u6_n2957 ), .ZN(_u10_u6_n2954 ) );
NAND2_X1 _u10_u6_U801  ( .A1(_u10_u6_n1853 ), .A2(_u10_u6_n1965 ), .ZN(_u10_u6_n2956 ) );
NAND2_X1 _u10_u6_U800  ( .A1(_u10_u6_n1966 ), .A2(_u10_u6_n2956 ), .ZN(_u10_u6_n2955 ) );
NAND2_X1 _u10_u6_U799  ( .A1(_u10_u6_n2954 ), .A2(_u10_u6_n2955 ), .ZN(_u10_u6_n2670 ) );
NOR3_X1 _u10_u6_U798  ( .A1(_u10_u6_n1852 ), .A2(1'b0), .A3(_u10_u6_n1853 ),.ZN(_u10_u6_n2708 ) );
NAND2_X1 _u10_u6_U797  ( .A1(_u10_u6_n2708 ), .A2(_u10_u6_n2080 ), .ZN(_u10_u6_n2355 ) );
NOR2_X1 _u10_u6_U796  ( .A1(_u10_u6_n2355 ), .A2(1'b0), .ZN(_u10_u6_n2599 ));
NAND2_X1 _u10_u6_U795  ( .A1(_u10_u6_n2953 ), .A2(_u10_u6_n2599 ), .ZN(_u10_u6_n2423 ) );
OR2_X1 _u10_u6_U794  ( .A1(_u10_u6_n2423 ), .A2(_u10_u6_n2359 ), .ZN(_u10_u6_n2949 ) );
NAND3_X1 _u10_u6_U793  ( .A1(_u10_u6_n2105 ), .A2(_u10_u6_n1936 ), .A3(_u10_u6_n2952 ), .ZN(_u10_u6_n2950 ) );
NAND3_X1 _u10_u6_U792  ( .A1(_u10_u6_n2549 ), .A2(_u10_u6_n1936 ), .A3(1'b0),.ZN(_u10_u6_n2096 ) );
INV_X1 _u10_u6_U791  ( .A(_u10_u6_n2096 ), .ZN(_u10_u6_n2301 ) );
NAND2_X1 _u10_u6_U790  ( .A1(_u10_u6_n2301 ), .A2(_u10_u6_n2446 ), .ZN(_u10_u6_n2368 ) );
INV_X1 _u10_u6_U789  ( .A(_u10_u6_n2368 ), .ZN(_u10_u6_n2326 ) );
NAND2_X1 _u10_u6_U788  ( .A1(_u10_u6_n2326 ), .A2(_u10_u6_n2941 ), .ZN(_u10_u6_n2800 ) );
INV_X1 _u10_u6_U787  ( .A(_u10_u6_n2800 ), .ZN(_u10_u6_n2081 ) );
NAND2_X1 _u10_u6_U786  ( .A1(_u10_u6_n2081 ), .A2(_u10_u6_n2049 ), .ZN(_u10_u6_n2855 ) );
INV_X1 _u10_u6_U785  ( .A(_u10_u6_n2855 ), .ZN(_u10_u6_n2347 ) );
NAND2_X1 _u10_u6_U784  ( .A1(_u10_u6_n2347 ), .A2(_u10_u6_n2063 ), .ZN(_u10_u6_n2951 ) );
NAND3_X1 _u10_u6_U783  ( .A1(_u10_u6_n2949 ), .A2(_u10_u6_n2950 ), .A3(_u10_u6_n2951 ), .ZN(_u10_u6_n1997 ) );
INV_X1 _u10_u6_U782  ( .A(_u10_u6_n1997 ), .ZN(_u10_u6_n2917 ) );
AND2_X1 _u10_u6_U781  ( .A1(_u10_u6_n2709 ), .A2(_u10_u6_n2708 ), .ZN(_u10_u6_n2942 ) );
INV_X1 _u10_u6_U780  ( .A(_u10_u6_n2907 ), .ZN(_u10_u6_n2737 ) );
NAND2_X1 _u10_u6_U779  ( .A1(_u10_u6_n2737 ), .A2(_u10_u6_n2803 ), .ZN(_u10_u6_n1888 ) );
NOR2_X1 _u10_u6_U778  ( .A1(_u10_u6_n2001 ), .A2(_u10_u6_n1888 ), .ZN(_u10_u6_n2943 ) );
NAND4_X1 _u10_u6_U777  ( .A1(1'b0), .A2(_u10_u6_n2078 ), .A3(_u10_u6_n2059 ),.A4(_u10_u6_n2031 ), .ZN(_u10_u6_n2578 ) );
NOR3_X1 _u10_u6_U776  ( .A1(_u10_u6_n2719 ), .A2(_u10_u6_n2130 ), .A3(_u10_u6_n2305 ), .ZN(_u10_u6_n2386 ) );
NAND2_X1 _u10_u6_U775  ( .A1(_u10_u6_n2386 ), .A2(_u10_u6_n2669 ), .ZN(_u10_u6_n2948 ) );
NAND3_X1 _u10_u6_U774  ( .A1(_u10_u6_n2578 ), .A2(_u10_u6_n2947 ), .A3(_u10_u6_n2948 ), .ZN(_u10_u6_n2750 ) );
NOR2_X1 _u10_u6_U773  ( .A1(_u10_u6_n2274 ), .A2(_u10_u6_n2852 ), .ZN(_u10_u6_n2946 ) );
NOR3_X1 _u10_u6_U772  ( .A1(_u10_u6_n2750 ), .A2(1'b0), .A3(_u10_u6_n2946 ),.ZN(_u10_u6_n2945 ) );
NOR2_X1 _u10_u6_U771  ( .A1(_u10_u6_n2945 ), .A2(_u10_u6_n2359 ), .ZN(_u10_u6_n2944 ) );
NOR3_X1 _u10_u6_U770  ( .A1(_u10_u6_n2942 ), .A2(_u10_u6_n2943 ), .A3(_u10_u6_n2944 ), .ZN(_u10_u6_n2919 ) );
NOR2_X1 _u10_u6_U769  ( .A1(_u10_u6_n2423 ), .A2(1'b0), .ZN(_u10_u6_n1979 ));
NAND3_X1 _u10_u6_U768  ( .A1(_u10_u6_n2549 ), .A2(_u10_u6_n1936 ), .A3(_u10_u6_n1979 ), .ZN(_u10_u6_n2328 ) );
INV_X1 _u10_u6_U767  ( .A(_u10_u6_n2328 ), .ZN(_u10_u6_n2554 ) );
NAND3_X1 _u10_u6_U766  ( .A1(_u10_u6_n2941 ), .A2(_u10_u6_n2446 ), .A3(_u10_u6_n2554 ), .ZN(_u10_u6_n2115 ) );
NOR2_X1 _u10_u6_U765  ( .A1(_u10_u6_n2578 ), .A2(_u10_u6_n2030 ), .ZN(_u10_u6_n2553 ) );
INV_X1 _u10_u6_U764  ( .A(_u10_u6_n2553 ), .ZN(_u10_u6_n2269 ) );
NOR2_X1 _u10_u6_U763  ( .A1(_u10_u6_n2269 ), .A2(_u10_u6_n2790 ), .ZN(_u10_u6_n2657 ) );
INV_X1 _u10_u6_U762  ( .A(_u10_u6_n2657 ), .ZN(_u10_u6_n2210 ) );
NOR2_X1 _u10_u6_U761  ( .A1(_u10_u6_n2210 ), .A2(_u10_u6_n2911 ), .ZN(_u10_u6_n2213 ) );
INV_X1 _u10_u6_U760  ( .A(_u10_u6_n2213 ), .ZN(_u10_u6_n2456 ) );
NAND2_X1 _u10_u6_U759  ( .A1(_u10_u6_n2115 ), .A2(_u10_u6_n2456 ), .ZN(_u10_u6_n2634 ) );
INV_X1 _u10_u6_U758  ( .A(_u10_u6_n2634 ), .ZN(_u10_u6_n2220 ) );
NOR2_X1 _u10_u6_U757  ( .A1(_u10_u6_n2081 ), .A2(_u10_u6_n2386 ), .ZN(_u10_u6_n2131 ) );
NAND2_X1 _u10_u6_U756  ( .A1(_u10_u6_n2940 ), .A2(_u10_u6_n2131 ), .ZN(_u10_u6_n2138 ) );
INV_X1 _u10_u6_U755  ( .A(_u10_u6_n2138 ), .ZN(_u10_u6_n2927 ) );
NAND2_X1 _u10_u6_U754  ( .A1(_u10_u6_n2220 ), .A2(_u10_u6_n2927 ), .ZN(_u10_u6_n2939 ) );
NAND2_X1 _u10_u6_U753  ( .A1(_u10_u6_n1885 ), .A2(_u10_u6_n2939 ), .ZN(_u10_u6_n2931 ) );
NAND3_X1 _u10_u6_U752  ( .A1(_u10_u6_n1859 ), .A2(_u10_u6_n2365 ), .A3(_u10_u6_n2938 ), .ZN(_u10_u6_n2935 ) );
NAND3_X1 _u10_u6_U751  ( .A1(_u10_u6_n2927 ), .A2(_u10_u6_n2937 ), .A3(_u10_u6_n2220 ), .ZN(_u10_u6_n2936 ) );
NAND2_X1 _u10_u6_U750  ( .A1(_u10_u6_n2935 ), .A2(_u10_u6_n2936 ), .ZN(_u10_u6_n2932 ) );
INV_X1 _u10_u6_U749  ( .A(_u10_u6_n1937 ), .ZN(_u10_u6_n2350 ) );
NAND2_X1 _u10_u6_U748  ( .A1(_u10_u6_n1913 ), .A2(_u10_u6_n2350 ), .ZN(_u10_u6_n2934 ) );
NAND2_X1 _u10_u6_U747  ( .A1(_u10_u6_n2386 ), .A2(_u10_u6_n2934 ), .ZN(_u10_u6_n2933 ) );
NAND3_X1 _u10_u6_U746  ( .A1(_u10_u6_n2931 ), .A2(_u10_u6_n2932 ), .A3(_u10_u6_n2933 ), .ZN(_u10_u6_n2921 ) );
OR2_X1 _u10_u6_U745  ( .A1(_u10_u6_n2213 ), .A2(_u10_u6_n2386 ), .ZN(_u10_u6_n2930 ) );
NAND2_X1 _u10_u6_U744  ( .A1(_u10_u6_n2049 ), .A2(_u10_u6_n2930 ), .ZN(_u10_u6_n2228 ) );
AND2_X1 _u10_u6_U743  ( .A1(_u10_u6_n2228 ), .A2(_u10_u6_n2699 ), .ZN(_u10_u6_n2929 ) );
NOR2_X1 _u10_u6_U742  ( .A1(_u10_u6_n2929 ), .A2(_u10_u6_n2495 ), .ZN(_u10_u6_n2922 ) );
NOR2_X1 _u10_u6_U741  ( .A1(_u10_u6_n2633 ), .A2(_u10_u6_n2877 ), .ZN(_u10_u6_n2928 ) );
NOR2_X1 _u10_u6_U740  ( .A1(_u10_u6_n2928 ), .A2(_u10_u6_n2886 ), .ZN(_u10_u6_n2923 ) );
NOR2_X1 _u10_u6_U739  ( .A1(_u10_u6_n2927 ), .A2(_u10_u6_n2531 ), .ZN(_u10_u6_n2926 ) );
NOR2_X1 _u10_u6_U738  ( .A1(_u10_u6_n2926 ), .A2(_u10_u6_n2687 ), .ZN(_u10_u6_n2925 ) );
NOR2_X1 _u10_u6_U737  ( .A1(_u10_u6_n2925 ), .A2(_u10_u6_n1849 ), .ZN(_u10_u6_n2924 ) );
NOR4_X1 _u10_u6_U736  ( .A1(_u10_u6_n2921 ), .A2(_u10_u6_n2922 ), .A3(_u10_u6_n2923 ), .A4(_u10_u6_n2924 ), .ZN(_u10_u6_n2920 ) );
NAND4_X1 _u10_u6_U735  ( .A1(_u10_u6_n2917 ), .A2(_u10_u6_n2918 ), .A3(_u10_u6_n2919 ), .A4(_u10_u6_n2920 ), .ZN(_u10_u6_n2312 ) );
NOR2_X1 _u10_u6_U734  ( .A1(_u10_u6_n2600 ), .A2(_u10_u6_n2686 ), .ZN(_u10_u6_n2401 ) );
NAND2_X1 _u10_u6_U733  ( .A1(_u10_u6_n2401 ), .A2(_u10_u6_n2549 ), .ZN(_u10_u6_n2547 ) );
INV_X1 _u10_u6_U732  ( .A(_u10_u6_n2547 ), .ZN(_u10_u6_n2794 ) );
NAND3_X1 _u10_u6_U731  ( .A1(_u10_u6_n2364 ), .A2(_u10_u6_n2667 ), .A3(_u10_u6_n2794 ), .ZN(_u10_u6_n2535 ) );
INV_X1 _u10_u6_U730  ( .A(_u10_u6_n2535 ), .ZN(_u10_u6_n2586 ) );
NAND2_X1 _u10_u6_U729  ( .A1(_u10_u6_n2586 ), .A2(_u10_u6_n2571 ), .ZN(_u10_u6_n2916 ) );
NAND2_X1 _u10_u6_U728  ( .A1(_u10_u6_n2837 ), .A2(_u10_u6_n2916 ), .ZN(_u10_u6_n2436 ) );
NAND2_X1 _u10_u6_U727  ( .A1(_u10_u6_n2915 ), .A2(_u10_u6_n2571 ), .ZN(_u10_u6_n2914 ) );
NAND2_X1 _u10_u6_U726  ( .A1(_u10_u6_n2166 ), .A2(_u10_u6_n2914 ), .ZN(_u10_u6_n2017 ) );
NOR2_X1 _u10_u6_U725  ( .A1(_u10_u6_n2485 ), .A2(_u10_u6_n1841 ), .ZN(_u10_u6_n2913 ) );
OR4_X1 _u10_u6_U724  ( .A1(_u10_u6_n2436 ), .A2(_u10_u6_n2017 ), .A3(_u10_u6_n2913 ), .A4(_u10_u6_n2442 ), .ZN(_u10_u6_n2912 ) );
NAND2_X1 _u10_u6_U723  ( .A1(_u10_u6_n2709 ), .A2(_u10_u6_n2912 ), .ZN(_u10_u6_n2888 ) );
NAND3_X1 _u10_u6_U722  ( .A1(_u10_u6_n2078 ), .A2(_u10_u6_n2031 ), .A3(1'b0),.ZN(_u10_u6_n2580 ) );
INV_X1 _u10_u6_U721  ( .A(_u10_u6_n2580 ), .ZN(_u10_u6_n2680 ) );
AND2_X1 _u10_u6_U720  ( .A1(_u10_u6_n2680 ), .A2(_u10_u6_n2668 ), .ZN(_u10_u6_n1950 ) );
NAND2_X1 _u10_u6_U719  ( .A1(_u10_u6_n1950 ), .A2(_u10_u6_n2089 ), .ZN(_u10_u6_n2095 ) );
INV_X1 _u10_u6_U718  ( .A(_u10_u6_n2095 ), .ZN(_u10_u6_n2542 ) );
NAND2_X1 _u10_u6_U717  ( .A1(_u10_u6_n2542 ), .A2(_u10_u6_n2446 ), .ZN(_u10_u6_n1887 ) );
NOR2_X1 _u10_u6_U716  ( .A1(_u10_u6_n1887 ), .A2(_u10_u6_n2911 ), .ZN(_u10_u6_n2114 ) );
INV_X1 _u10_u6_U715  ( .A(_u10_u6_n2114 ), .ZN(_u10_u6_n1940 ) );
NAND3_X1 _u10_u6_U714  ( .A1(_u10_u6_n2535 ), .A2(_u10_u6_n1940 ), .A3(_u10_u6_n2910 ), .ZN(_u10_u6_n2524 ) );
NAND2_X1 _u10_u6_U713  ( .A1(_u10_u6_n2524 ), .A2(_u10_u6_n2488 ), .ZN(_u10_u6_n2889 ) );
NAND2_X1 _u10_u6_U712  ( .A1(_u10_u6_n2220 ), .A2(_u10_u6_n1940 ), .ZN(_u10_u6_n2763 ) );
NOR2_X1 _u10_u6_U711  ( .A1(_u10_u6_n2763 ), .A2(_u10_u6_n2586 ), .ZN(_u10_u6_n2808 ) );
NOR2_X1 _u10_u6_U710  ( .A1(_u10_u6_n2808 ), .A2(_u10_u6_n2350 ), .ZN(_u10_u6_n2908 ) );
NOR2_X1 _u10_u6_U709  ( .A1(_u10_u6_n2544 ), .A2(_u10_u6_n1950 ), .ZN(_u10_u6_n2899 ) );
NOR2_X1 _u10_u6_U708  ( .A1(_u10_u6_n2899 ), .A2(_u10_u6_n2159 ), .ZN(_u10_u6_n2909 ) );
NOR2_X1 _u10_u6_U707  ( .A1(_u10_u6_n2908 ), .A2(_u10_u6_n2909 ), .ZN(_u10_u6_n2890 ) );
NOR3_X1 _u10_u6_U706  ( .A1(_u10_u6_n2547 ), .A2(_u10_u6_n1846 ), .A3(_u10_u6_n2907 ), .ZN(_u10_u6_n2892 ) );
NOR3_X1 _u10_u6_U705  ( .A1(_u10_u6_n2240 ), .A2(_u10_u6_n2377 ), .A3(_u10_u6_n1911 ), .ZN(_u10_u6_n2906 ) );
NOR2_X1 _u10_u6_U704  ( .A1(_u10_u6_n2906 ), .A2(_u10_u6_n2535 ), .ZN(_u10_u6_n2893 ) );
NAND2_X1 _u10_u6_U703  ( .A1(_u10_u6_n2554 ), .A2(_u10_u6_n2446 ), .ZN(_u10_u6_n2903 ) );
AND3_X1 _u10_u6_U702  ( .A1(_u10_u6_n2210 ), .A2(_u10_u6_n2905 ), .A3(_u10_u6_n1887 ), .ZN(_u10_u6_n2904 ) );
NAND4_X1 _u10_u6_U701  ( .A1(_u10_u6_n2902 ), .A2(_u10_u6_n2498 ), .A3(_u10_u6_n2903 ), .A4(_u10_u6_n2904 ), .ZN(_u10_u6_n2788 ) );
INV_X1 _u10_u6_U700  ( .A(_u10_u6_n2788 ), .ZN(_u10_u6_n2901 ) );
NOR2_X1 _u10_u6_U699  ( .A1(_u10_u6_n2901 ), .A2(_u10_u6_n1888 ), .ZN(_u10_u6_n2894 ) );
NOR2_X1 _u10_u6_U698  ( .A1(_u10_u6_n2401 ), .A2(_u10_u6_n2553 ), .ZN(_u10_u6_n2900 ) );
NOR2_X1 _u10_u6_U697  ( .A1(_u10_u6_n2900 ), .A2(_u10_u6_n1954 ), .ZN(_u10_u6_n2897 ) );
NOR2_X1 _u10_u6_U696  ( .A1(1'b0), .A2(_u10_u6_n2899 ), .ZN(_u10_u6_n2898 ));
NOR2_X1 _u10_u6_U695  ( .A1(_u10_u6_n2897 ), .A2(_u10_u6_n2898 ), .ZN(_u10_u6_n2896 ) );
NOR2_X1 _u10_u6_U694  ( .A1(_u10_u6_n2896 ), .A2(_u10_u6_n1843 ), .ZN(_u10_u6_n2895 ) );
NOR4_X1 _u10_u6_U693  ( .A1(_u10_u6_n2892 ), .A2(_u10_u6_n2893 ), .A3(_u10_u6_n2894 ), .A4(_u10_u6_n2895 ), .ZN(_u10_u6_n2891 ) );
NAND4_X1 _u10_u6_U692  ( .A1(_u10_u6_n2888 ), .A2(_u10_u6_n2889 ), .A3(_u10_u6_n2890 ), .A4(_u10_u6_n2891 ), .ZN(_u10_u6_n2610 ) );
NOR4_X1 _u10_u6_U691  ( .A1(_u10_u6_n2670 ), .A2(_u10_u6_n2312 ), .A3(_u10_u6_n2610 ), .A4(_u10_u6_n2887 ), .ZN(_u10_u6_n2724 ) );
NOR2_X1 _u10_u6_U690  ( .A1(_u10_u6_n2883 ), .A2(_u10_u6_n2535 ), .ZN(_u10_u6_n2861 ) );
NOR2_X1 _u10_u6_U689  ( .A1(_u10_u6_n1855 ), .A2(_u10_u6_n1869 ), .ZN(_u10_u6_n2862 ) );
NOR2_X1 _u10_u6_U688  ( .A1(_u10_u6_n2886 ), .A2(_u10_u6_n2695 ), .ZN(_u10_u6_n2863 ) );
NAND2_X1 _u10_u6_U687  ( .A1(_u10_u6_n2813 ), .A2(_u10_u6_n2885 ), .ZN(_u10_u6_n2864 ) );
NAND2_X1 _u10_u6_U686  ( .A1(_u10_u6_n2114 ), .A2(_u10_u6_n2884 ), .ZN(_u10_u6_n2865 ) );
NAND2_X1 _u10_u6_U685  ( .A1(1'b0), .A2(_u10_u6_n2667 ), .ZN(_u10_u6_n2112 ));
NOR3_X1 _u10_u6_U684  ( .A1(_u10_u6_n2883 ), .A2(_u10_u6_n2112 ), .A3(_u10_u6_n2719 ), .ZN(_u10_u6_n2878 ) );
INV_X1 _u10_u6_U683  ( .A(_u10_u6_n2112 ), .ZN(_u10_u6_n1856 ) );
NAND2_X1 _u10_u6_U682  ( .A1(_u10_u6_n2364 ), .A2(_u10_u6_n1856 ), .ZN(_u10_u6_n2882 ) );
NAND2_X1 _u10_u6_U681  ( .A1(_u10_u6_n2882 ), .A2(_u10_u6_n1869 ), .ZN(_u10_u6_n2050 ) );
INV_X1 _u10_u6_U680  ( .A(_u10_u6_n2050 ), .ZN(_u10_u6_n1939 ) );
NOR2_X1 _u10_u6_U679  ( .A1(_u10_u6_n1939 ), .A2(_u10_u6_n1841 ), .ZN(_u10_u6_n2881 ) );
NOR2_X1 _u10_u6_U678  ( .A1(_u10_u6_n2881 ), .A2(_u10_u6_n2840 ), .ZN(_u10_u6_n2880 ) );
NOR2_X1 _u10_u6_U677  ( .A1(_u10_u6_n2880 ), .A2(_u10_u6_n1836 ), .ZN(_u10_u6_n2879 ) );
NOR2_X1 _u10_u6_U676  ( .A1(_u10_u6_n2878 ), .A2(_u10_u6_n2879 ), .ZN(_u10_u6_n2866 ) );
NOR2_X1 _u10_u6_U675  ( .A1(_u10_u6_n2081 ), .A2(_u10_u6_n2877 ), .ZN(_u10_u6_n1840 ) );
NAND2_X1 _u10_u6_U674  ( .A1(_u10_u6_n1840 ), .A2(_u10_u6_n2115 ), .ZN(_u10_u6_n1873 ) );
NAND2_X1 _u10_u6_U673  ( .A1(_u10_u6_n2695 ), .A2(_u10_u6_n1940 ), .ZN(_u10_u6_n1874 ) );
NOR3_X1 _u10_u6_U672  ( .A1(_u10_u6_n2050 ), .A2(_u10_u6_n1873 ), .A3(_u10_u6_n1874 ), .ZN(_u10_u6_n2876 ) );
NOR2_X1 _u10_u6_U671  ( .A1(_u10_u6_n2876 ), .A2(_u10_u6_n1913 ), .ZN(_u10_u6_n2868 ) );
NAND2_X1 _u10_u6_U670  ( .A1(_u10_u6_n2875 ), .A2(_u10_u6_n2466 ), .ZN(_u10_u6_n2872 ) );
INV_X1 _u10_u6_U669  ( .A(_u10_u6_n1979 ), .ZN(_u10_u6_n2746 ) );
NAND2_X1 _u10_u6_U668  ( .A1(_u10_u6_n2874 ), .A2(_u10_u6_n2746 ), .ZN(_u10_u6_n1935 ) );
NAND3_X1 _u10_u6_U667  ( .A1(_u10_u6_n1935 ), .A2(_u10_u6_n1936 ), .A3(_u10_u6_n2467 ), .ZN(_u10_u6_n2873 ) );
NAND2_X1 _u10_u6_U666  ( .A1(_u10_u6_n2872 ), .A2(_u10_u6_n2873 ), .ZN(_u10_u6_n2264 ) );
AND2_X1 _u10_u6_U665  ( .A1(_u10_u6_n2264 ), .A2(_u10_u6_n2461 ), .ZN(_u10_u6_n2869 ) );
AND2_X1 _u10_u6_U664  ( .A1(_u10_u6_n1966 ), .A2(_u10_u6_n2761 ), .ZN(_u10_u6_n2870 ) );
NOR2_X1 _u10_u6_U663  ( .A1(_u10_u6_n2159 ), .A2(_u10_u6_n2163 ), .ZN(_u10_u6_n2871 ) );
NOR4_X1 _u10_u6_U662  ( .A1(_u10_u6_n2868 ), .A2(_u10_u6_n2869 ), .A3(_u10_u6_n2870 ), .A4(_u10_u6_n2871 ), .ZN(_u10_u6_n2867 ) );
NAND4_X1 _u10_u6_U661  ( .A1(_u10_u6_n2864 ), .A2(_u10_u6_n2865 ), .A3(_u10_u6_n2866 ), .A4(_u10_u6_n2867 ), .ZN(_u10_u6_n1992 ) );
NOR4_X1 _u10_u6_U660  ( .A1(_u10_u6_n2861 ), .A2(_u10_u6_n2862 ), .A3(_u10_u6_n2863 ), .A4(_u10_u6_n1992 ), .ZN(_u10_u6_n2725 ) );
NAND2_X1 _u10_u6_U659  ( .A1(_u10_u6_n2364 ), .A2(_u10_u6_n1846 ), .ZN(_u10_u6_n2744 ) );
NAND4_X1 _u10_u6_U658  ( .A1(_u10_u6_n2765 ), .A2(_u10_u6_n1939 ), .A3(_u10_u6_n2744 ), .A4(_u10_u6_n2535 ), .ZN(_u10_u6_n2860 ) );
NAND2_X1 _u10_u6_U657  ( .A1(_u10_u6_n2049 ), .A2(_u10_u6_n2860 ), .ZN(_u10_u6_n2856 ) );
NOR4_X1 _u10_u6_U656  ( .A1(1'b0), .A2(_u10_u6_n2858 ), .A3(_u10_u6_n2859 ),.A4(_u10_u6_n2051 ), .ZN(_u10_u6_n2857 ) );
NAND4_X1 _u10_u6_U655  ( .A1(_u10_u6_n2228 ), .A2(_u10_u6_n2855 ), .A3(_u10_u6_n2856 ), .A4(_u10_u6_n2857 ), .ZN(_u10_u6_n2854 ) );
NAND2_X1 _u10_u6_U654  ( .A1(_u10_u6_n2043 ), .A2(_u10_u6_n2854 ), .ZN(_u10_u6_n2821 ) );
INV_X1 _u10_u6_U653  ( .A(_u10_u6_n2071 ), .ZN(_u10_u6_n2279 ) );
INV_X1 _u10_u6_U652  ( .A(_u10_u6_n2599 ), .ZN(_u10_u6_n2357 ) );
OR2_X1 _u10_u6_U651  ( .A1(_u10_u6_n2744 ), .A2(_u10_u6_n2853 ), .ZN(_u10_u6_n2844 ) );
NAND2_X1 _u10_u6_U650  ( .A1(_u10_u6_n2131 ), .A2(_u10_u6_n2852 ), .ZN(_u10_u6_n2851 ) );
NAND2_X1 _u10_u6_U649  ( .A1(_u10_u6_n2082 ), .A2(_u10_u6_n2851 ), .ZN(_u10_u6_n2848 ) );
NAND2_X1 _u10_u6_U648  ( .A1(_u10_u6_n2850 ), .A2(_u10_u6_n2600 ), .ZN(_u10_u6_n2849 ) );
NAND3_X1 _u10_u6_U647  ( .A1(_u10_u6_n2848 ), .A2(_u10_u6_n2077 ), .A3(_u10_u6_n2849 ), .ZN(_u10_u6_n2287 ) );
NAND2_X1 _u10_u6_U646  ( .A1(_u10_u6_n2082 ), .A2(_u10_u6_n2050 ), .ZN(_u10_u6_n2847 ) );
NAND2_X1 _u10_u6_U645  ( .A1(_u10_u6_n2846 ), .A2(_u10_u6_n2847 ), .ZN(_u10_u6_n2074 ) );
NOR3_X1 _u10_u6_U644  ( .A1(_u10_u6_n2287 ), .A2(_u10_u6_n2596 ), .A3(_u10_u6_n2074 ), .ZN(_u10_u6_n2845 ) );
NAND4_X1 _u10_u6_U643  ( .A1(_u10_u6_n2357 ), .A2(_u10_u6_n2837 ), .A3(_u10_u6_n2844 ), .A4(_u10_u6_n2845 ), .ZN(_u10_u6_n2843 ) );
NAND2_X1 _u10_u6_U642  ( .A1(_u10_u6_n2279 ), .A2(_u10_u6_n2843 ), .ZN(_u10_u6_n2822 ) );
NOR3_X1 _u10_u6_U641  ( .A1(_u10_u6_n1925 ), .A2(_u10_u6_n2842 ), .A3(_u10_u6_n2686 ), .ZN(_u10_u6_n2841 ) );
NOR3_X1 _u10_u6_U640  ( .A1(_u10_u6_n2840 ), .A2(_u10_u6_n2599 ), .A3(_u10_u6_n2841 ), .ZN(_u10_u6_n2839 ) );
AND4_X1 _u10_u6_U639  ( .A1(_u10_u6_n2836 ), .A2(_u10_u6_n2837 ), .A3(_u10_u6_n2838 ), .A4(_u10_u6_n2839 ), .ZN(_u10_u6_n2454 ) );
NOR2_X1 _u10_u6_U638  ( .A1(_u10_u6_n2719 ), .A2(_u10_u6_n2835 ), .ZN(_u10_u6_n2773 ) );
NOR2_X1 _u10_u6_U637  ( .A1(_u10_u6_n2138 ), .A2(_u10_u6_n2773 ), .ZN(_u10_u6_n2814 ) );
NAND2_X1 _u10_u6_U636  ( .A1(_u10_u6_n2814 ), .A2(_u10_u6_n1869 ), .ZN(_u10_u6_n2834 ) );
NAND2_X1 _u10_u6_U635  ( .A1(_u10_u6_n2833 ), .A2(_u10_u6_n2834 ), .ZN(_u10_u6_n2832 ) );
NAND2_X1 _u10_u6_U634  ( .A1(_u10_u6_n2454 ), .A2(_u10_u6_n2832 ), .ZN(_u10_u6_n2831 ) );
NAND2_X1 _u10_u6_U633  ( .A1(_u10_u6_n2830 ), .A2(_u10_u6_n2831 ), .ZN(_u10_u6_n2823 ) );
INV_X1 _u10_u6_U632  ( .A(_u10_u6_n2025 ), .ZN(_u10_u6_n2470 ) );
NAND2_X1 _u10_u6_U631  ( .A1(_u10_u6_n1979 ), .A2(_u10_u6_n1936 ), .ZN(_u10_u6_n2829 ) );
AND2_X1 _u10_u6_U630  ( .A1(_u10_u6_n2828 ), .A2(_u10_u6_n2829 ), .ZN(_u10_u6_n2469 ) );
NAND2_X1 _u10_u6_U629  ( .A1(_u10_u6_n2469 ), .A2(_u10_u6_n2269 ), .ZN(_u10_u6_n2161 ) );
INV_X1 _u10_u6_U628  ( .A(_u10_u6_n2161 ), .ZN(_u10_u6_n2276 ) );
NOR2_X1 _u10_u6_U627  ( .A1(_u10_u6_n2274 ), .A2(_u10_u6_n2719 ), .ZN(_u10_u6_n2827 ) );
NOR3_X1 _u10_u6_U626  ( .A1(_u10_u6_n2827 ), .A2(_u10_u6_n2742 ), .A3(_u10_u6_n2680 ), .ZN(_u10_u6_n2826 ) );
NAND3_X1 _u10_u6_U625  ( .A1(_u10_u6_n2276 ), .A2(_u10_u6_n2108 ), .A3(_u10_u6_n2826 ), .ZN(_u10_u6_n2825 ) );
NAND2_X1 _u10_u6_U624  ( .A1(_u10_u6_n2470 ), .A2(_u10_u6_n2825 ), .ZN(_u10_u6_n2824 ) );
NAND4_X1 _u10_u6_U623  ( .A1(_u10_u6_n2821 ), .A2(_u10_u6_n2822 ), .A3(_u10_u6_n2823 ), .A4(_u10_u6_n2824 ), .ZN(_u10_u6_n2804 ) );
NAND2_X1 _u10_u6_U622  ( .A1(_u10_u6_n2131 ), .A2(_u10_u6_n2744 ), .ZN(_u10_u6_n2820 ) );
NAND2_X1 _u10_u6_U621  ( .A1(_u10_u6_n2571 ), .A2(_u10_u6_n2820 ), .ZN(_u10_u6_n2817 ) );
NOR2_X1 _u10_u6_U620  ( .A1(_u10_u6_n2819 ), .A2(_u10_u6_n2436 ), .ZN(_u10_u6_n2818 ) );
NAND4_X1 _u10_u6_U619  ( .A1(_u10_u6_n2437 ), .A2(_u10_u6_n2355 ), .A3(_u10_u6_n2817 ), .A4(_u10_u6_n2818 ), .ZN(_u10_u6_n2816 ) );
NAND2_X1 _u10_u6_U618  ( .A1(_u10_u6_n2815 ), .A2(_u10_u6_n2816 ), .ZN(_u10_u6_n2809 ) );
INV_X1 _u10_u6_U617  ( .A(_u10_u6_n2814 ), .ZN(_u10_u6_n2812 ) );
OR2_X1 _u10_u6_U616  ( .A1(_u10_u6_n1911 ), .A2(_u10_u6_n2813 ), .ZN(_u10_u6_n1884 ) );
NAND2_X1 _u10_u6_U615  ( .A1(_u10_u6_n2812 ), .A2(_u10_u6_n1884 ), .ZN(_u10_u6_n2810 ) );
NOR2_X1 _u10_u6_U614  ( .A1(_u10_u6_n1894 ), .A2(_u10_u6_n2461 ), .ZN(_u10_u6_n1948 ) );
OR2_X1 _u10_u6_U613  ( .A1(_u10_u6_n1847 ), .A2(_u10_u6_n1948 ), .ZN(_u10_u6_n2811 ) );
NAND3_X1 _u10_u6_U612  ( .A1(_u10_u6_n2809 ), .A2(_u10_u6_n2810 ), .A3(_u10_u6_n2811 ), .ZN(_u10_u6_n2805 ) );
NOR2_X1 _u10_u6_U611  ( .A1(_u10_u6_n2808 ), .A2(_u10_u6_n2775 ), .ZN(_u10_u6_n2806 ) );
AND2_X1 _u10_u6_U610  ( .A1(_u10_u6_n2721 ), .A2(_u10_u6_n1911 ), .ZN(_u10_u6_n2807 ) );
NOR4_X1 _u10_u6_U609  ( .A1(_u10_u6_n2804 ), .A2(_u10_u6_n2805 ), .A3(_u10_u6_n2806 ), .A4(_u10_u6_n2807 ), .ZN(_u10_u6_n2726 ) );
NAND2_X1 _u10_u6_U608  ( .A1(_u10_u6_n2803 ), .A2(_u10_u6_n2112 ), .ZN(_u10_u6_n2802 ) );
NAND2_X1 _u10_u6_U607  ( .A1(_u10_u6_n2364 ), .A2(_u10_u6_n2802 ), .ZN(_u10_u6_n2801 ) );
NAND2_X1 _u10_u6_U606  ( .A1(_u10_u6_n2800 ), .A2(_u10_u6_n2801 ), .ZN(_u10_u6_n2799 ) );
NAND2_X1 _u10_u6_U605  ( .A1(_u10_u6_n1937 ), .A2(_u10_u6_n2799 ), .ZN(_u10_u6_n2780 ) );
NAND2_X1 _u10_u6_U604  ( .A1(_u10_u6_n2775 ), .A2(_u10_u6_n2798 ), .ZN(_u10_u6_n2796 ) );
INV_X1 _u10_u6_U603  ( .A(_u10_u6_n2131 ), .ZN(_u10_u6_n2797 ) );
NAND2_X1 _u10_u6_U602  ( .A1(_u10_u6_n2796 ), .A2(_u10_u6_n2797 ), .ZN(_u10_u6_n2781 ) );
OR4_X1 _u10_u6_U601  ( .A1(_u10_u6_n2795 ), .A2(_u10_u6_n2303 ), .A3(_u10_u6_n2553 ), .A4(_u10_u6_n2554 ), .ZN(_u10_u6_n2792 ) );
NAND3_X1 _u10_u6_U600  ( .A1(_u10_u6_n1847 ), .A2(_u10_u6_n2097 ), .A3(_u10_u6_n2096 ), .ZN(_u10_u6_n2793 ) );
NOR4_X1 _u10_u6_U599  ( .A1(_u10_u6_n2792 ), .A2(_u10_u6_n2793 ), .A3(_u10_u6_n2542 ), .A4(_u10_u6_n2794 ), .ZN(_u10_u6_n2791 ) );
NOR2_X1 _u10_u6_U598  ( .A1(_u10_u6_n2791 ), .A2(_u10_u6_n2085 ), .ZN(_u10_u6_n2783 ) );
NAND2_X1 _u10_u6_U597  ( .A1(_u10_u6_n2114 ), .A2(_u10_u6_n2049 ), .ZN(_u10_u6_n2700 ) );
INV_X1 _u10_u6_U596  ( .A(_u10_u6_n2700 ), .ZN(_u10_u6_n2784 ) );
NAND4_X1 _u10_u6_U595  ( .A1(_u10_u6_n2001 ), .A2(_u10_u6_n2547 ), .A3(_u10_u6_n2368 ), .A4(_u10_u6_n1847 ), .ZN(_u10_u6_n2787 ) );
NOR4_X1 _u10_u6_U594  ( .A1(_u10_u6_n2787 ), .A2(_u10_u6_n2788 ), .A3(_u10_u6_n2789 ), .A4(_u10_u6_n2790 ), .ZN(_u10_u6_n2786 ) );
NOR2_X1 _u10_u6_U593  ( .A1(_u10_u6_n2786 ), .A2(_u10_u6_n2000 ), .ZN(_u10_u6_n2785 ) );
NOR3_X1 _u10_u6_U592  ( .A1(_u10_u6_n2783 ), .A2(_u10_u6_n2784 ), .A3(_u10_u6_n2785 ), .ZN(_u10_u6_n2782 ) );
NAND3_X1 _u10_u6_U591  ( .A1(_u10_u6_n2780 ), .A2(_u10_u6_n2781 ), .A3(_u10_u6_n2782 ), .ZN(_u10_u6_n2728 ) );
OR3_X1 _u10_u6_U590  ( .A1(_u10_u6_n2138 ), .A2(_u10_u6_n2633 ), .A3(_u10_u6_n2779 ), .ZN(_u10_u6_n2778 ) );
NAND2_X1 _u10_u6_U589  ( .A1(_u10_u6_n2777 ), .A2(_u10_u6_n2778 ), .ZN(_u10_u6_n2767 ) );
NAND3_X1 _u10_u6_U588  ( .A1(_u10_u6_n2775 ), .A2(_u10_u6_n2083 ), .A3(_u10_u6_n2776 ), .ZN(_u10_u6_n2774 ) );
NAND2_X1 _u10_u6_U587  ( .A1(_u10_u6_n2773 ), .A2(_u10_u6_n2774 ), .ZN(_u10_u6_n2768 ) );
NAND2_X1 _u10_u6_U586  ( .A1(_u10_u6_n2218 ), .A2(_u10_u6_n2772 ), .ZN(_u10_u6_n2769 ) );
NAND2_X1 _u10_u6_U585  ( .A1(_u10_u6_n2302 ), .A2(_u10_u6_n2467 ), .ZN(_u10_u6_n2771 ) );
NAND2_X1 _u10_u6_U584  ( .A1(_u10_u6_n2461 ), .A2(_u10_u6_n2771 ), .ZN(_u10_u6_n2770 ) );
NAND4_X1 _u10_u6_U583  ( .A1(_u10_u6_n2767 ), .A2(_u10_u6_n2768 ), .A3(_u10_u6_n2769 ), .A4(_u10_u6_n2770 ), .ZN(_u10_u6_n2729 ) );
NAND3_X1 _u10_u6_U582  ( .A1(_u10_u6_n2668 ), .A2(_u10_u6_n2600 ), .A3(_u10_u6_n2276 ), .ZN(_u10_u6_n2766 ) );
NAND2_X1 _u10_u6_U581  ( .A1(_u10_u6_n1894 ), .A2(_u10_u6_n2766 ), .ZN(_u10_u6_n2753 ) );
NAND3_X1 _u10_u6_U580  ( .A1(_u10_u6_n2456 ), .A2(_u10_u6_n2744 ), .A3(_u10_u6_n2765 ), .ZN(_u10_u6_n2764 ) );
NAND2_X1 _u10_u6_U579  ( .A1(_u10_u6_n2377 ), .A2(_u10_u6_n2764 ), .ZN(_u10_u6_n2754 ) );
NAND2_X1 _u10_u6_U578  ( .A1(_u10_u6_n2763 ), .A2(_u10_u6_n2007 ), .ZN(_u10_u6_n2755 ) );
NOR2_X1 _u10_u6_U577  ( .A1(_u10_u6_n2531 ), .A2(_u10_u6_n2744 ), .ZN(_u10_u6_n2760 ) );
INV_X1 _u10_u6_U576  ( .A(_u10_u6_n2762 ), .ZN(_u10_u6_n2189 ) );
NOR3_X1 _u10_u6_U575  ( .A1(_u10_u6_n2760 ), .A2(_u10_u6_n2761 ), .A3(_u10_u6_n2189 ), .ZN(_u10_u6_n2759 ) );
NOR2_X1 _u10_u6_U574  ( .A1(_u10_u6_n2759 ), .A2(_u10_u6_n1849 ), .ZN(_u10_u6_n2757 ) );
NOR2_X1 _u10_u6_U573  ( .A1(_u10_u6_n1817 ), .A2(_u10_u6_n2665 ), .ZN(_u10_u6_n2758 ) );
NOR2_X1 _u10_u6_U572  ( .A1(_u10_u6_n2757 ), .A2(_u10_u6_n2758 ), .ZN(_u10_u6_n2756 ) );
NAND4_X1 _u10_u6_U571  ( .A1(_u10_u6_n2753 ), .A2(_u10_u6_n2754 ), .A3(_u10_u6_n2755 ), .A4(_u10_u6_n2756 ), .ZN(_u10_u6_n2730 ) );
INV_X1 _u10_u6_U570  ( .A(_u10_u6_n2359 ), .ZN(_u10_u6_n1899 ) );
NAND4_X1 _u10_u6_U569  ( .A1(_u10_u6_n2078 ), .A2(_u10_u6_n2580 ), .A3(_u10_u6_n2748 ), .A4(_u10_u6_n2752 ), .ZN(_u10_u6_n2751 ) );
NAND2_X1 _u10_u6_U568  ( .A1(_u10_u6_n1899 ), .A2(_u10_u6_n2751 ), .ZN(_u10_u6_n2732 ) );
INV_X1 _u10_u6_U567  ( .A(_u10_u6_n2750 ), .ZN(_u10_u6_n2379 ) );
NAND3_X1 _u10_u6_U566  ( .A1(_u10_u6_n1856 ), .A2(_u10_u6_n2669 ), .A3(_u10_u6_n2364 ), .ZN(_u10_u6_n2749 ) );
AND2_X1 _u10_u6_U565  ( .A1(_u10_u6_n2748 ), .A2(_u10_u6_n2749 ), .ZN(_u10_u6_n2034 ) );
NAND2_X1 _u10_u6_U564  ( .A1(_u10_u6_n2105 ), .A2(_u10_u6_n2669 ), .ZN(_u10_u6_n2745 ) );
AND3_X1 _u10_u6_U563  ( .A1(_u10_u6_n2745 ), .A2(_u10_u6_n2746 ), .A3(_u10_u6_n2747 ), .ZN(_u10_u6_n2380 ) );
NOR2_X1 _u10_u6_U562  ( .A1(_u10_u6_n2274 ), .A2(_u10_u6_n2744 ), .ZN(_u10_u6_n2743 ) );
NOR4_X1 _u10_u6_U561  ( .A1(_u10_u6_n2742 ), .A2(_u10_u6_n2680 ), .A3(_u10_u6_n2743 ), .A4(_u10_u6_n2428 ), .ZN(_u10_u6_n2741 ) );
NAND4_X1 _u10_u6_U560  ( .A1(_u10_u6_n2379 ), .A2(_u10_u6_n2034 ), .A3(_u10_u6_n2380 ), .A4(_u10_u6_n2741 ), .ZN(_u10_u6_n2740 ) );
NAND2_X1 _u10_u6_U559  ( .A1(_u10_u6_n1967 ), .A2(_u10_u6_n2740 ), .ZN(_u10_u6_n2733 ) );
NAND3_X1 _u10_u6_U558  ( .A1(_u10_u6_n2739 ), .A2(_u10_u6_n2368 ), .A3(_u10_u6_n2255 ), .ZN(_u10_u6_n2738 ) );
NAND2_X1 _u10_u6_U557  ( .A1(_u10_u6_n2737 ), .A2(_u10_u6_n2738 ), .ZN(_u10_u6_n2734 ) );
NAND2_X1 _u10_u6_U556  ( .A1(_u10_u6_n2736 ), .A2(_u10_u6_n2524 ), .ZN(_u10_u6_n2735 ) );
NAND4_X1 _u10_u6_U555  ( .A1(_u10_u6_n2732 ), .A2(_u10_u6_n2733 ), .A3(_u10_u6_n2734 ), .A4(_u10_u6_n2735 ), .ZN(_u10_u6_n2731 ) );
NOR4_X1 _u10_u6_U554  ( .A1(_u10_u6_n2728 ), .A2(_u10_u6_n2729 ), .A3(_u10_u6_n2730 ), .A4(_u10_u6_n2731 ), .ZN(_u10_u6_n2727 ) );
NAND4_X1 _u10_u6_U553  ( .A1(_u10_u6_n2724 ), .A2(_u10_u6_n2725 ), .A3(_u10_u6_n2726 ), .A4(_u10_u6_n2727 ), .ZN(_u10_u6_n2723 ) );
MUX2_X1 _u10_u6_U552  ( .A(_u10_u6_n2723 ), .B(_u10_SYNOPSYS_UNCONNECTED_24 ), .S(_u10_u6_n1819 ), .Z(_u10_u6_n1809 ) );
NAND2_X1 _u10_u6_U551  ( .A1(_u10_u6_n2002 ), .A2(_u10_u6_n2722 ), .ZN(_u10_u6_n2713 ) );
NAND2_X1 _u10_u6_U550  ( .A1(_u10_u6_n2720 ), .A2(_u10_u6_n2721 ), .ZN(_u10_u6_n2714 ) );
NAND2_X1 _u10_u6_U549  ( .A1(_u10_u6_n2256 ), .A2(_u10_u6_n2719 ), .ZN(_u10_u6_n2715 ) );
NOR2_X1 _u10_u6_U548  ( .A1(_u10_u6_n2106 ), .A2(_u10_u6_n2037 ), .ZN(_u10_u6_n2717 ) );
AND2_X1 _u10_u6_U547  ( .A1(_u10_u6_n1966 ), .A2(_u10_u6_n2054 ), .ZN(_u10_u6_n2718 ) );
NOR2_X1 _u10_u6_U546  ( .A1(_u10_u6_n2717 ), .A2(_u10_u6_n2718 ), .ZN(_u10_u6_n2716 ) );
NAND4_X1 _u10_u6_U545  ( .A1(_u10_u6_n2713 ), .A2(_u10_u6_n2714 ), .A3(_u10_u6_n2715 ), .A4(_u10_u6_n2716 ), .ZN(_u10_u6_n2608 ) );
NAND2_X1 _u10_u6_U544  ( .A1(1'b0), .A2(_u10_u6_n2669 ), .ZN(_u10_u6_n2385 ));
INV_X1 _u10_u6_U543  ( .A(_u10_u6_n2385 ), .ZN(_u10_u6_n1977 ) );
NAND2_X1 _u10_u6_U542  ( .A1(_u10_u6_n1977 ), .A2(_u10_u6_n2668 ), .ZN(_u10_u6_n2712 ) );
NAND2_X1 _u10_u6_U541  ( .A1(_u10_u6_n2712 ), .A2(_u10_u6_n2092 ), .ZN(_u10_u6_n1844 ) );
NAND2_X1 _u10_u6_U540  ( .A1(_u10_u6_n1894 ), .A2(_u10_u6_n1844 ), .ZN(_u10_u6_n2705 ) );
NAND2_X1 _u10_u6_U539  ( .A1(_u10_u6_n1894 ), .A2(_u10_u6_n2305 ), .ZN(_u10_u6_n2711 ) );
NAND2_X1 _u10_u6_U538  ( .A1(_u10_u6_n2711 ), .A2(_u10_u6_n2025 ), .ZN(_u10_u6_n1932 ) );
NAND2_X1 _u10_u6_U537  ( .A1(_u10_u6_n2710 ), .A2(_u10_u6_n1932 ), .ZN(_u10_u6_n2706 ) );
NAND2_X1 _u10_u6_U536  ( .A1(_u10_u6_n2708 ), .A2(_u10_u6_n2709 ), .ZN(_u10_u6_n2707 ) );
NAND3_X1 _u10_u6_U535  ( .A1(_u10_u6_n2705 ), .A2(_u10_u6_n2706 ), .A3(_u10_u6_n2707 ), .ZN(_u10_u6_n2701 ) );
NOR2_X1 _u10_u6_U534  ( .A1(_u10_u6_n1843 ), .A2(_u10_u6_n2545 ), .ZN(_u10_u6_n2702 ) );
NOR2_X1 _u10_u6_U533  ( .A1(_u10_u6_n2346 ), .A2(_u10_u6_n2700 ), .ZN(_u10_u6_n2703 ) );
NOR2_X1 _u10_u6_U532  ( .A1(_u10_u6_n2000 ), .A2(_u10_u6_n1887 ), .ZN(_u10_u6_n2704 ) );
NOR4_X1 _u10_u6_U531  ( .A1(_u10_u6_n2701 ), .A2(_u10_u6_n2702 ), .A3(_u10_u6_n2703 ), .A4(_u10_u6_n2704 ), .ZN(_u10_u6_n2671 ) );
NAND2_X1 _u10_u6_U530  ( .A1(_u10_u6_n2699 ), .A2(_u10_u6_n2700 ), .ZN(_u10_u6_n2698 ) );
NAND2_X1 _u10_u6_U529  ( .A1(_u10_u6_n2063 ), .A2(_u10_u6_n2698 ), .ZN(_u10_u6_n2682 ) );
NAND2_X1 _u10_u6_U528  ( .A1(_u10_u6_n2697 ), .A2(_u10_u6_n2103 ), .ZN(_u10_u6_n2696 ) );
NAND2_X1 _u10_u6_U527  ( .A1(_u10_u6_n2695 ), .A2(_u10_u6_n2696 ), .ZN(_u10_u6_n2694 ) );
NAND2_X1 _u10_u6_U526  ( .A1(_u10_u6_n1937 ), .A2(_u10_u6_n2694 ), .ZN(_u10_u6_n2683 ) );
INV_X1 _u10_u6_U525  ( .A(_u10_u6_n2693 ), .ZN(_u10_u6_n2691 ) );
NAND3_X1 _u10_u6_U524  ( .A1(_u10_u6_n2103 ), .A2(_u10_u6_n2502 ), .A3(1'b0),.ZN(_u10_u6_n2692 ) );
NAND2_X1 _u10_u6_U523  ( .A1(_u10_u6_n2691 ), .A2(_u10_u6_n2692 ), .ZN(_u10_u6_n2690 ) );
NAND2_X1 _u10_u6_U522  ( .A1(_u10_u6_n2236 ), .A2(_u10_u6_n2690 ), .ZN(_u10_u6_n2684 ) );
NAND3_X1 _u10_u6_U521  ( .A1(_u10_u6_n2688 ), .A2(_u10_u6_n1913 ), .A3(_u10_u6_n2689 ), .ZN(_u10_u6_n2335 ) );
NAND3_X1 _u10_u6_U520  ( .A1(_u10_u6_n2536 ), .A2(_u10_u6_n2103 ), .A3(1'b0),.ZN(_u10_u6_n2052 ) );
NOR2_X1 _u10_u6_U519  ( .A1(_u10_u6_n2052 ), .A2(_u10_u6_n2687 ), .ZN(_u10_u6_n1851 ) );
NAND2_X1 _u10_u6_U518  ( .A1(_u10_u6_n1851 ), .A2(_u10_u6_n2078 ), .ZN(_u10_u6_n2582 ) );
NOR2_X1 _u10_u6_U517  ( .A1(_u10_u6_n2686 ), .A2(_u10_u6_n2582 ), .ZN(_u10_u6_n2094 ) );
NAND3_X1 _u10_u6_U516  ( .A1(_u10_u6_n2251 ), .A2(_u10_u6_n2335 ), .A3(_u10_u6_n2094 ), .ZN(_u10_u6_n2685 ) );
NAND4_X1 _u10_u6_U515  ( .A1(_u10_u6_n2682 ), .A2(_u10_u6_n2683 ), .A3(_u10_u6_n2684 ), .A4(_u10_u6_n2685 ), .ZN(_u10_u6_n2673 ) );
INV_X1 _u10_u6_U514  ( .A(_u10_u6_n2291 ), .ZN(_u10_u6_n2057 ) );
AND2_X1 _u10_u6_U513  ( .A1(_u10_u6_n1851 ), .A2(_u10_u6_n2057 ), .ZN(_u10_u6_n2674 ) );
INV_X1 _u10_u6_U512  ( .A(_u10_u6_n1874 ), .ZN(_u10_u6_n2681 ) );
NOR2_X1 _u10_u6_U511  ( .A1(_u10_u6_n2007 ), .A2(_u10_u6_n1911 ), .ZN(_u10_u6_n2486 ) );
NOR2_X1 _u10_u6_U510  ( .A1(_u10_u6_n2681 ), .A2(_u10_u6_n2486 ), .ZN(_u10_u6_n2675 ) );
NOR2_X1 _u10_u6_U509  ( .A1(_u10_u6_n1977 ), .A2(_u10_u6_n2680 ), .ZN(_u10_u6_n2679 ) );
NOR2_X1 _u10_u6_U508  ( .A1(_u10_u6_n2679 ), .A2(_u10_u6_n2030 ), .ZN(_u10_u6_n2678 ) );
NOR2_X1 _u10_u6_U507  ( .A1(_u10_u6_n2678 ), .A2(_u10_u6_n2094 ), .ZN(_u10_u6_n2677 ) );
NOR2_X1 _u10_u6_U506  ( .A1(_u10_u6_n2677 ), .A2(_u10_u6_n2025 ), .ZN(_u10_u6_n2676 ) );
NOR4_X1 _u10_u6_U505  ( .A1(_u10_u6_n2673 ), .A2(_u10_u6_n2674 ), .A3(_u10_u6_n2675 ), .A4(_u10_u6_n2676 ), .ZN(_u10_u6_n2672 ) );
AND2_X1 _u10_u6_U504  ( .A1(_u10_u6_n2671 ), .A2(_u10_u6_n2672 ), .ZN(_u10_u6_n1990 ) );
INV_X1 _u10_u6_U503  ( .A(_u10_u6_n2670 ), .ZN(_u10_u6_n2660 ) );
NAND4_X1 _u10_u6_U502  ( .A1(_u10_u6_n2251 ), .A2(_u10_u6_n2669 ), .A3(_u10_u6_n2162 ), .A4(_u10_u6_n2169 ), .ZN(_u10_u6_n2664 ) );
AND3_X1 _u10_u6_U501  ( .A1(_u10_u6_n1977 ), .A2(_u10_u6_n2668 ), .A3(_u10_u6_n2089 ), .ZN(_u10_u6_n2555 ) );
NAND2_X1 _u10_u6_U500  ( .A1(_u10_u6_n2555 ), .A2(_u10_u6_n2667 ), .ZN(_u10_u6_n2666 ) );
NAND3_X1 _u10_u6_U499  ( .A1(_u10_u6_n2664 ), .A2(_u10_u6_n2665 ), .A3(_u10_u6_n2666 ), .ZN(_u10_u6_n1988 ) );
INV_X1 _u10_u6_U498  ( .A(_u10_u6_n1988 ), .ZN(_u10_u6_n2661 ) );
NAND2_X1 _u10_u6_U497  ( .A1(1'b0), .A2(_u10_u6_n2043 ), .ZN(_u10_u6_n2662 ));
NAND2_X1 _u10_u6_U496  ( .A1(_u10_u6_n2169 ), .A2(1'b0), .ZN(_u10_u6_n2663 ));
NAND4_X1 _u10_u6_U495  ( .A1(_u10_u6_n2660 ), .A2(_u10_u6_n2661 ), .A3(_u10_u6_n2662 ), .A4(_u10_u6_n2663 ), .ZN(_u10_u6_n2650 ) );
NAND2_X1 _u10_u6_U494  ( .A1(_u10_u6_n2659 ), .A2(1'b0), .ZN(_u10_u6_n2193 ));
INV_X1 _u10_u6_U493  ( .A(_u10_u6_n2193 ), .ZN(_u10_u6_n2143 ) );
NAND2_X1 _u10_u6_U492  ( .A1(_u10_u6_n2143 ), .A2(_u10_u6_n2036 ), .ZN(_u10_u6_n2286 ) );
INV_X1 _u10_u6_U491  ( .A(_u10_u6_n2286 ), .ZN(_u10_u6_n2577 ) );
NAND2_X1 _u10_u6_U490  ( .A1(_u10_u6_n2577 ), .A2(_u10_u6_n2278 ), .ZN(_u10_u6_n2474 ) );
INV_X1 _u10_u6_U489  ( .A(_u10_u6_n2474 ), .ZN(_u10_u6_n2306 ) );
NAND2_X1 _u10_u6_U488  ( .A1(_u10_u6_n2306 ), .A2(_u10_u6_n2251 ), .ZN(_u10_u6_n2654 ) );
NAND2_X1 _u10_u6_U487  ( .A1(_u10_u6_n2649 ), .A2(_u10_u6_n2658 ), .ZN(_u10_u6_n2655 ) );
NAND2_X1 _u10_u6_U486  ( .A1(_u10_u6_n2657 ), .A2(_u10_u6_n2445 ), .ZN(_u10_u6_n2656 ) );
NAND3_X1 _u10_u6_U485  ( .A1(_u10_u6_n2654 ), .A2(_u10_u6_n2655 ), .A3(_u10_u6_n2656 ), .ZN(_u10_u6_n2651 ) );
NOR2_X1 _u10_u6_U484  ( .A1(_u10_u6_n2366 ), .A2(_u10_u6_n2376 ), .ZN(_u10_u6_n2652 ) );
AND2_X1 _u10_u6_U483  ( .A1(_u10_u6_n1966 ), .A2(_u10_u6_n2528 ), .ZN(_u10_u6_n2653 ) );
NOR4_X1 _u10_u6_U482  ( .A1(_u10_u6_n2650 ), .A2(_u10_u6_n2651 ), .A3(_u10_u6_n2652 ), .A4(_u10_u6_n2653 ), .ZN(_u10_u6_n2613 ) );
NAND2_X1 _u10_u6_U481  ( .A1(_u10_u6_n1891 ), .A2(1'b0), .ZN(_u10_u6_n2636 ));
NAND2_X1 _u10_u6_U480  ( .A1(_u10_u6_n1868 ), .A2(_u10_u6_n2113 ), .ZN(_u10_u6_n2101 ) );
NOR4_X1 _u10_u6_U479  ( .A1(_u10_u6_n2649 ), .A2(_u10_u6_n2216 ), .A3(_u10_u6_n2101 ), .A4(_u10_u6_n2634 ), .ZN(_u10_u6_n2648 ) );
NOR2_X1 _u10_u6_U478  ( .A1(_u10_u6_n2648 ), .A2(_u10_u6_n2254 ), .ZN(_u10_u6_n2638 ) );
NOR2_X1 _u10_u6_U477  ( .A1(_u10_u6_n2106 ), .A2(_u10_u6_n2643 ), .ZN(_u10_u6_n2645 ) );
NAND2_X1 _u10_u6_U476  ( .A1(1'b0), .A2(_u10_u6_n2049 ), .ZN(_u10_u6_n2647 ));
NAND2_X1 _u10_u6_U475  ( .A1(_u10_u6_n2646 ), .A2(_u10_u6_n2647 ), .ZN(_u10_u6_n2348 ) );
NOR2_X1 _u10_u6_U474  ( .A1(_u10_u6_n2645 ), .A2(_u10_u6_n2348 ), .ZN(_u10_u6_n2644 ) );
NOR2_X1 _u10_u6_U473  ( .A1(_u10_u6_n2644 ), .A2(_u10_u6_n2495 ), .ZN(_u10_u6_n2639 ) );
NOR2_X1 _u10_u6_U472  ( .A1(_u10_u6_n2643 ), .A2(_u10_u6_n2203 ), .ZN(_u10_u6_n2642 ) );
NOR3_X1 _u10_u6_U471  ( .A1(_u10_u6_n2101 ), .A2(1'b0), .A3(_u10_u6_n2642 ),.ZN(_u10_u6_n2641 ) );
NOR2_X1 _u10_u6_U470  ( .A1(_u10_u6_n2641 ), .A2(_u10_u6_n2253 ), .ZN(_u10_u6_n2640 ) );
NOR3_X1 _u10_u6_U469  ( .A1(_u10_u6_n2638 ), .A2(_u10_u6_n2639 ), .A3(_u10_u6_n2640 ), .ZN(_u10_u6_n2637 ) );
NAND3_X1 _u10_u6_U468  ( .A1(_u10_u6_n2635 ), .A2(_u10_u6_n2636 ), .A3(_u10_u6_n2637 ), .ZN(_u10_u6_n2615 ) );
NOR3_X1 _u10_u6_U467  ( .A1(_u10_u6_n2174 ), .A2(_u10_u6_n2175 ), .A3(_u10_u6_n2179 ), .ZN(_u10_u6_n2631 ) );
NAND3_X1 _u10_u6_U466  ( .A1(_u10_u6_n2223 ), .A2(_u10_u6_n2236 ), .A3(_u10_u6_n2631 ), .ZN(_u10_u6_n2622 ) );
OR2_X1 _u10_u6_U465  ( .A1(_u10_u6_n1960 ), .A2(_u10_u6_n1959 ), .ZN(_u10_u6_n2625 ) );
NOR3_X1 _u10_u6_U464  ( .A1(_u10_u6_n2101 ), .A2(_u10_u6_n2633 ), .A3(_u10_u6_n2634 ), .ZN(_u10_u6_n2523 ) );
OR2_X1 _u10_u6_U463  ( .A1(_u10_u6_n2632 ), .A2(_u10_u6_n2523 ), .ZN(_u10_u6_n2627 ) );
INV_X1 _u10_u6_U462  ( .A(_u10_u6_n2631 ), .ZN(_u10_u6_n2628 ) );
NAND2_X1 _u10_u6_U461  ( .A1(_u10_u6_n2630 ), .A2(_u10_u6_n1922 ), .ZN(_u10_u6_n2629 ) );
NAND3_X1 _u10_u6_U460  ( .A1(_u10_u6_n2627 ), .A2(_u10_u6_n2628 ), .A3(_u10_u6_n2629 ), .ZN(_u10_u6_n2626 ) );
NAND2_X1 _u10_u6_U459  ( .A1(_u10_u6_n2625 ), .A2(_u10_u6_n2626 ), .ZN(_u10_u6_n2624 ) );
NAND3_X1 _u10_u6_U458  ( .A1(_u10_u6_n2622 ), .A2(_u10_u6_n2623 ), .A3(_u10_u6_n2624 ), .ZN(_u10_u6_n2616 ) );
AND2_X1 _u10_u6_U457  ( .A1(_u10_u6_n2621 ), .A2(_u10_u6_n2358 ), .ZN(_u10_u6_n2620 ) );
NOR2_X1 _u10_u6_U456  ( .A1(_u10_u6_n2523 ), .A2(_u10_u6_n2620 ), .ZN(_u10_u6_n2617 ) );
INV_X1 _u10_u6_U455  ( .A(_u10_u6_n2101 ), .ZN(_u10_u6_n2221 ) );
NOR2_X1 _u10_u6_U454  ( .A1(_u10_u6_n1911 ), .A2(_u10_u6_n2488 ), .ZN(_u10_u6_n2619 ) );
NOR2_X1 _u10_u6_U453  ( .A1(_u10_u6_n2221 ), .A2(_u10_u6_n2619 ), .ZN(_u10_u6_n2618 ) );
NOR4_X1 _u10_u6_U452  ( .A1(_u10_u6_n2615 ), .A2(_u10_u6_n2616 ), .A3(_u10_u6_n2617 ), .A4(_u10_u6_n2618 ), .ZN(_u10_u6_n2614 ) );
AND2_X1 _u10_u6_U451  ( .A1(_u10_u6_n2613 ), .A2(_u10_u6_n2614 ), .ZN(_u10_u6_n2314 ) );
NAND3_X1 _u10_u6_U450  ( .A1(_u10_u6_n2612 ), .A2(_u10_u6_n1990 ), .A3(_u10_u6_n2314 ), .ZN(_u10_u6_n2609 ) );
NOR4_X1 _u10_u6_U449  ( .A1(_u10_u6_n2608 ), .A2(_u10_u6_n2609 ), .A3(_u10_u6_n2610 ), .A4(_u10_u6_n2611 ), .ZN(_u10_u6_n2388 ) );
NAND2_X1 _u10_u6_U448  ( .A1(_u10_u6_n2346 ), .A2(_u10_u6_n2607 ), .ZN(_u10_u6_n2191 ) );
NAND2_X1 _u10_u6_U447  ( .A1(_u10_u6_n2143 ), .A2(_u10_u6_n2191 ), .ZN(_u10_u6_n2556 ) );
INV_X1 _u10_u6_U446  ( .A(_u10_u6_n2348 ), .ZN(_u10_u6_n2603 ) );
NAND3_X1 _u10_u6_U445  ( .A1(_u10_u6_n2535 ), .A2(_u10_u6_n2485 ), .A3(_u10_u6_n2456 ), .ZN(_u10_u6_n2606 ) );
NAND2_X1 _u10_u6_U444  ( .A1(_u10_u6_n2049 ), .A2(_u10_u6_n2606 ), .ZN(_u10_u6_n2604 ) );
NAND3_X1 _u10_u6_U443  ( .A1(_u10_u6_n2603 ), .A2(_u10_u6_n2604 ), .A3(_u10_u6_n2605 ), .ZN(_u10_u6_n2602 ) );
NAND2_X1 _u10_u6_U442  ( .A1(_u10_u6_n2043 ), .A2(_u10_u6_n2602 ), .ZN(_u10_u6_n2557 ) );
INV_X1 _u10_u6_U441  ( .A(_u10_u6_n2601 ), .ZN(_u10_u6_n2590 ) );
NAND2_X1 _u10_u6_U440  ( .A1(_u10_u6_n2599 ), .A2(_u10_u6_n2600 ), .ZN(_u10_u6_n2597 ) );
NAND2_X1 _u10_u6_U439  ( .A1(_u10_u6_n2082 ), .A2(_u10_u6_n2101 ), .ZN(_u10_u6_n2598 ) );
AND2_X1 _u10_u6_U438  ( .A1(_u10_u6_n2597 ), .A2(_u10_u6_n2598 ), .ZN(_u10_u6_n2281 ) );
NAND3_X1 _u10_u6_U437  ( .A1(_u10_u6_n1969 ), .A2(_u10_u6_n2582 ), .A3(_u10_u6_n2281 ), .ZN(_u10_u6_n2073 ) );
INV_X1 _u10_u6_U436  ( .A(_u10_u6_n2073 ), .ZN(_u10_u6_n2591 ) );
NOR2_X1 _u10_u6_U435  ( .A1(_u10_u6_n1816 ), .A2(_u10_u6_n2077 ), .ZN(_u10_u6_n2595 ) );
NOR2_X1 _u10_u6_U434  ( .A1(_u10_u6_n2595 ), .A2(_u10_u6_n2596 ), .ZN(_u10_u6_n2592 ) );
NAND3_X1 _u10_u6_U433  ( .A1(_u10_u6_n2107 ), .A2(_u10_u6_n2536 ), .A3(1'b0),.ZN(_u10_u6_n2438 ) );
INV_X1 _u10_u6_U432  ( .A(_u10_u6_n2438 ), .ZN(_u10_u6_n2427 ) );
NOR4_X1 _u10_u6_U431  ( .A1(1'b0), .A2(_u10_u6_n2594 ), .A3(_u10_u6_n2577 ),.A4(_u10_u6_n2427 ), .ZN(_u10_u6_n2593 ) );
NAND4_X1 _u10_u6_U430  ( .A1(_u10_u6_n2590 ), .A2(_u10_u6_n2591 ), .A3(_u10_u6_n2592 ), .A4(_u10_u6_n2593 ), .ZN(_u10_u6_n2589 ) );
NAND2_X1 _u10_u6_U429  ( .A1(_u10_u6_n2279 ), .A2(_u10_u6_n2589 ), .ZN(_u10_u6_n2558 ) );
NAND3_X1 _u10_u6_U428  ( .A1(_u10_u6_n2587 ), .A2(_u10_u6_n2115 ), .A3(_u10_u6_n2588 ), .ZN(_u10_u6_n2585 ) );
NOR4_X1 _u10_u6_U427  ( .A1(_u10_u6_n2585 ), .A2(_u10_u6_n2586 ), .A3(1'b0),.A4(_u10_u6_n2114 ), .ZN(_u10_u6_n2583 ) );
NOR2_X1 _u10_u6_U426  ( .A1(_u10_u6_n2583 ), .A2(_u10_u6_n2584 ), .ZN(_u10_u6_n2560 ) );
OR2_X1 _u10_u6_U425  ( .A1(_u10_u6_n2582 ), .A2(1'b0), .ZN(_u10_u6_n2581 ));
NAND2_X1 _u10_u6_U424  ( .A1(_u10_u6_n2580 ), .A2(_u10_u6_n2581 ), .ZN(_u10_u6_n1974 ) );
INV_X1 _u10_u6_U423  ( .A(_u10_u6_n1974 ), .ZN(_u10_u6_n1901 ) );
AND4_X1 _u10_u6_U422  ( .A1(_u10_u6_n1901 ), .A2(_u10_u6_n2385 ), .A3(_u10_u6_n2578 ), .A4(_u10_u6_n2579 ), .ZN(_u10_u6_n2424 ) );
NOR2_X1 _u10_u6_U421  ( .A1(1'b0), .A2(_u10_u6_n2424 ), .ZN(_u10_u6_n2574 ));
NOR3_X1 _u10_u6_U420  ( .A1(_u10_u6_n2427 ), .A2(1'b0), .A3(_u10_u6_n2577 ),.ZN(_u10_u6_n2576 ) );
NOR2_X1 _u10_u6_U419  ( .A1(_u10_u6_n2576 ), .A2(_u10_u6_n1976 ), .ZN(_u10_u6_n2575 ) );
NOR3_X1 _u10_u6_U418  ( .A1(_u10_u6_n2574 ), .A2(_u10_u6_n1979 ), .A3(_u10_u6_n2575 ), .ZN(_u10_u6_n2572 ) );
NOR2_X1 _u10_u6_U417  ( .A1(_u10_u6_n2572 ), .A2(_u10_u6_n2573 ), .ZN(_u10_u6_n2561 ) );
INV_X1 _u10_u6_U416  ( .A(_u10_u6_n2061 ), .ZN(_u10_u6_n2453 ) );
NOR2_X1 _u10_u6_U415  ( .A1(_u10_u6_n2453 ), .A2(_u10_u6_n1851 ), .ZN(_u10_u6_n2018 ) );
NAND2_X1 _u10_u6_U414  ( .A1(1'b0), .A2(_u10_u6_n2571 ), .ZN(_u10_u6_n2570 ));
NAND2_X1 _u10_u6_U413  ( .A1(_u10_u6_n2018 ), .A2(_u10_u6_n2570 ), .ZN(_u10_u6_n1837 ) );
INV_X1 _u10_u6_U412  ( .A(_u10_u6_n1837 ), .ZN(_u10_u6_n2568 ) );
NAND2_X1 _u10_u6_U411  ( .A1(1'b0), .A2(_u10_u6_n2536 ), .ZN(_u10_u6_n2569 ));
NAND2_X1 _u10_u6_U410  ( .A1(_u10_u6_n2568 ), .A2(_u10_u6_n2569 ), .ZN(_u10_u6_n2564 ) );
NOR2_X1 _u10_u6_U409  ( .A1(_u10_u6_n1841 ), .A2(_u10_u6_n1868 ), .ZN(_u10_u6_n2565 ) );
INV_X1 _u10_u6_U408  ( .A(_u10_u6_n2567 ), .ZN(_u10_u6_n2566 ) );
NOR4_X1 _u10_u6_U407  ( .A1(_u10_u6_n2564 ), .A2(_u10_u6_n2565 ), .A3(_u10_u6_n2143 ), .A4(_u10_u6_n2566 ), .ZN(_u10_u6_n2563 ) );
NOR2_X1 _u10_u6_U406  ( .A1(_u10_u6_n2563 ), .A2(_u10_u6_n2014 ), .ZN(_u10_u6_n2562 ) );
NOR3_X1 _u10_u6_U405  ( .A1(_u10_u6_n2560 ), .A2(_u10_u6_n2561 ), .A3(_u10_u6_n2562 ), .ZN(_u10_u6_n2559 ) );
NAND4_X1 _u10_u6_U404  ( .A1(_u10_u6_n2556 ), .A2(_u10_u6_n2557 ), .A3(_u10_u6_n2558 ), .A4(_u10_u6_n2559 ), .ZN(_u10_u6_n2511 ) );
INV_X1 _u10_u6_U403  ( .A(_u10_u6_n2085 ), .ZN(_u10_u6_n2293 ) );
NOR2_X1 _u10_u6_U402  ( .A1(_u10_u6_n2554 ), .A2(_u10_u6_n2555 ), .ZN(_u10_u6_n2444 ) );
NAND2_X1 _u10_u6_U401  ( .A1(_u10_u6_n2553 ), .A2(_u10_u6_n2549 ), .ZN(_u10_u6_n2552 ) );
AND2_X1 _u10_u6_U400  ( .A1(_u10_u6_n2444 ), .A2(_u10_u6_n2552 ), .ZN(_u10_u6_n2295 ) );
NAND2_X1 _u10_u6_U399  ( .A1(_u10_u6_n2551 ), .A2(_u10_u6_n2549 ), .ZN(_u10_u6_n2538 ) );
AND2_X1 _u10_u6_U398  ( .A1(_u10_u6_n2427 ), .A2(_u10_u6_n2108 ), .ZN(_u10_u6_n2460 ) );
NOR4_X1 _u10_u6_U397  ( .A1(_u10_u6_n2460 ), .A2(_u10_u6_n2306 ), .A3(_u10_u6_n2094 ), .A4(_u10_u6_n2550 ), .ZN(_u10_u6_n2409 ) );
INV_X1 _u10_u6_U396  ( .A(_u10_u6_n2409 ), .ZN(_u10_u6_n2407 ) );
NAND2_X1 _u10_u6_U395  ( .A1(_u10_u6_n2549 ), .A2(_u10_u6_n2407 ), .ZN(_u10_u6_n2546 ) );
NAND3_X1 _u10_u6_U394  ( .A1(_u10_u6_n2546 ), .A2(_u10_u6_n2547 ), .A3(_u10_u6_n2548 ), .ZN(_u10_u6_n2501 ) );
INV_X1 _u10_u6_U393  ( .A(_u10_u6_n2501 ), .ZN(_u10_u6_n2539 ) );
NOR2_X1 _u10_u6_U392  ( .A1(1'b0), .A2(_u10_u6_n2545 ), .ZN(_u10_u6_n2541 ));
AND2_X1 _u10_u6_U391  ( .A1(_u10_u6_n2544 ), .A2(_u10_u6_n2089 ), .ZN(_u10_u6_n2543 ) );
NOR3_X1 _u10_u6_U390  ( .A1(_u10_u6_n2541 ), .A2(_u10_u6_n2542 ), .A3(_u10_u6_n2543 ), .ZN(_u10_u6_n2540 ) );
NAND4_X1 _u10_u6_U389  ( .A1(_u10_u6_n2295 ), .A2(_u10_u6_n2538 ), .A3(_u10_u6_n2539 ), .A4(_u10_u6_n2540 ), .ZN(_u10_u6_n2537 ) );
NAND2_X1 _u10_u6_U388  ( .A1(_u10_u6_n2293 ), .A2(_u10_u6_n2537 ), .ZN(_u10_u6_n2515 ) );
NAND2_X1 _u10_u6_U387  ( .A1(_u10_u6_n2536 ), .A2(_u10_u6_n2508 ), .ZN(_u10_u6_n2526 ) );
NAND2_X1 _u10_u6_U386  ( .A1(_u10_u6_n2535 ), .A2(_u10_u6_n1940 ), .ZN(_u10_u6_n2532 ) );
NOR4_X1 _u10_u6_U385  ( .A1(_u10_u6_n2532 ), .A2(_u10_u6_n2533 ), .A3(1'b0),.A4(_u10_u6_n2534 ), .ZN(_u10_u6_n2530 ) );
NOR2_X1 _u10_u6_U384  ( .A1(_u10_u6_n2530 ), .A2(_u10_u6_n2531 ), .ZN(_u10_u6_n2529 ) );
NOR4_X1 _u10_u6_U383  ( .A1(_u10_u6_n2528 ), .A2(_u10_u6_n2143 ), .A3(_u10_u6_n2189 ), .A4(_u10_u6_n2529 ), .ZN(_u10_u6_n2527 ) );
NAND4_X1 _u10_u6_U382  ( .A1(_u10_u6_n2019 ), .A2(_u10_u6_n2526 ), .A3(_u10_u6_n2018 ), .A4(_u10_u6_n2527 ), .ZN(_u10_u6_n2525 ) );
NAND2_X1 _u10_u6_U381  ( .A1(_u10_u6_n2183 ), .A2(_u10_u6_n2525 ), .ZN(_u10_u6_n2516 ) );
INV_X1 _u10_u6_U380  ( .A(_u10_u6_n2524 ), .ZN(_u10_u6_n2396 ) );
NAND2_X1 _u10_u6_U379  ( .A1(_u10_u6_n2396 ), .A2(_u10_u6_n2523 ), .ZN(_u10_u6_n2522 ) );
NAND2_X1 _u10_u6_U378  ( .A1(_u10_u6_n1866 ), .A2(_u10_u6_n2522 ), .ZN(_u10_u6_n2519 ) );
AND2_X1 _u10_u6_U377  ( .A1(_u10_u6_n2493 ), .A2(_u10_u6_n1961 ), .ZN(_u10_u6_n2429 ) );
NAND2_X1 _u10_u6_U376  ( .A1(_u10_u6_n2429 ), .A2(_u10_u6_n2175 ), .ZN(_u10_u6_n2510 ) );
NAND2_X1 _u10_u6_U375  ( .A1(_u10_u6_n2510 ), .A2(_u10_u6_n1864 ), .ZN(_u10_u6_n2521 ) );
NAND3_X1 _u10_u6_U374  ( .A1(_u10_u6_n2519 ), .A2(_u10_u6_n2520 ), .A3(_u10_u6_n2521 ), .ZN(_u10_u6_n2518 ) );
NAND2_X1 _u10_u6_U373  ( .A1(_u10_u6_n1861 ), .A2(_u10_u6_n2518 ), .ZN(_u10_u6_n2517 ) );
NAND3_X1 _u10_u6_U372  ( .A1(_u10_u6_n2515 ), .A2(_u10_u6_n2516 ), .A3(_u10_u6_n2517 ), .ZN(_u10_u6_n2512 ) );
NOR2_X1 _u10_u6_U371  ( .A1(_u10_u6_n1913 ), .A2(_u10_u6_n1940 ), .ZN(_u10_u6_n2513 ) );
NOR2_X1 _u10_u6_U370  ( .A1(_u10_u6_n2113 ), .A2(_u10_u6_n2350 ), .ZN(_u10_u6_n2514 ) );
NOR4_X1 _u10_u6_U369  ( .A1(_u10_u6_n2511 ), .A2(_u10_u6_n2512 ), .A3(_u10_u6_n2513 ), .A4(_u10_u6_n2514 ), .ZN(_u10_u6_n2389 ) );
NAND2_X1 _u10_u6_U368  ( .A1(_u10_u6_n2509 ), .A2(_u10_u6_n2510 ), .ZN(_u10_u6_n2477 ) );
NAND2_X1 _u10_u6_U367  ( .A1(_u10_u6_n2507 ), .A2(_u10_u6_n2508 ), .ZN(_u10_u6_n2504 ) );
NAND2_X1 _u10_u6_U366  ( .A1(1'b0), .A2(_u10_u6_n2506 ), .ZN(_u10_u6_n2505 ));
NAND2_X1 _u10_u6_U365  ( .A1(_u10_u6_n2504 ), .A2(_u10_u6_n2505 ), .ZN(_u10_u6_n2503 ) );
NAND2_X1 _u10_u6_U364  ( .A1(_u10_u6_n2502 ), .A2(_u10_u6_n2503 ), .ZN(_u10_u6_n2478 ) );
NAND2_X1 _u10_u6_U363  ( .A1(_u10_u6_n2501 ), .A2(_u10_u6_n2446 ), .ZN(_u10_u6_n2497 ) );
INV_X1 _u10_u6_U362  ( .A(_u10_u6_n2500 ), .ZN(_u10_u6_n2499 ) );
NAND3_X1 _u10_u6_U361  ( .A1(_u10_u6_n2497 ), .A2(_u10_u6_n2498 ), .A3(_u10_u6_n2499 ), .ZN(_u10_u6_n2496 ) );
NAND2_X1 _u10_u6_U360  ( .A1(_u10_u6_n2445 ), .A2(_u10_u6_n2496 ), .ZN(_u10_u6_n2479 ) );
NOR2_X1 _u10_u6_U359  ( .A1(_u10_u6_n2429 ), .A2(_u10_u6_n2495 ), .ZN(_u10_u6_n2491 ) );
INV_X1 _u10_u6_U358  ( .A(_u10_u6_n2191 ), .ZN(_u10_u6_n2494 ) );
NOR2_X1 _u10_u6_U357  ( .A1(_u10_u6_n2493 ), .A2(_u10_u6_n2494 ), .ZN(_u10_u6_n2492 ) );
NOR2_X1 _u10_u6_U356  ( .A1(_u10_u6_n2491 ), .A2(_u10_u6_n2492 ), .ZN(_u10_u6_n2489 ) );
NOR2_X1 _u10_u6_U355  ( .A1(_u10_u6_n2489 ), .A2(_u10_u6_n2490 ), .ZN(_u10_u6_n2481 ) );
NAND2_X1 _u10_u6_U354  ( .A1(_u10_u6_n2253 ), .A2(_u10_u6_n1859 ), .ZN(_u10_u6_n2398 ) );
NOR2_X1 _u10_u6_U353  ( .A1(_u10_u6_n2488 ), .A2(_u10_u6_n2398 ), .ZN(_u10_u6_n2487 ) );
NOR2_X1 _u10_u6_U352  ( .A1(_u10_u6_n2220 ), .A2(_u10_u6_n2487 ), .ZN(_u10_u6_n2482 ) );
AND2_X1 _u10_u6_U351  ( .A1(_u10_u6_n2350 ), .A2(_u10_u6_n2486 ), .ZN(_u10_u6_n2484 ) );
NOR2_X1 _u10_u6_U350  ( .A1(_u10_u6_n2484 ), .A2(_u10_u6_n2485 ), .ZN(_u10_u6_n2483 ) );
NOR3_X1 _u10_u6_U349  ( .A1(_u10_u6_n2481 ), .A2(_u10_u6_n2482 ), .A3(_u10_u6_n2483 ), .ZN(_u10_u6_n2480 ) );
NAND4_X1 _u10_u6_U348  ( .A1(_u10_u6_n2477 ), .A2(_u10_u6_n2478 ), .A3(_u10_u6_n2479 ), .A4(_u10_u6_n2480 ), .ZN(_u10_u6_n2447 ) );
NAND2_X1 _u10_u6_U347  ( .A1(_u10_u6_n2476 ), .A2(_u10_u6_n1936 ), .ZN(_u10_u6_n2472 ) );
NAND2_X1 _u10_u6_U346  ( .A1(_u10_u6_n2427 ), .A2(_u10_u6_n2278 ), .ZN(_u10_u6_n2473 ) );
NAND4_X1 _u10_u6_U345  ( .A1(_u10_u6_n2472 ), .A2(_u10_u6_n2473 ), .A3(_u10_u6_n2474 ), .A4(_u10_u6_n2475 ), .ZN(_u10_u6_n2471 ) );
NAND2_X1 _u10_u6_U344  ( .A1(_u10_u6_n2470 ), .A2(_u10_u6_n2471 ), .ZN(_u10_u6_n2457 ) );
NAND2_X1 _u10_u6_U343  ( .A1(_u10_u6_n2409 ), .A2(_u10_u6_n2469 ), .ZN(_u10_u6_n2468 ) );
NAND2_X1 _u10_u6_U342  ( .A1(_u10_u6_n2467 ), .A2(_u10_u6_n2468 ), .ZN(_u10_u6_n2463 ) );
NAND2_X1 _u10_u6_U341  ( .A1(_u10_u6_n1844 ), .A2(_u10_u6_n2466 ), .ZN(_u10_u6_n2465 ) );
NAND3_X1 _u10_u6_U340  ( .A1(_u10_u6_n2463 ), .A2(_u10_u6_n2464 ), .A3(_u10_u6_n2465 ), .ZN(_u10_u6_n2462 ) );
NAND2_X1 _u10_u6_U339  ( .A1(_u10_u6_n2461 ), .A2(_u10_u6_n2462 ), .ZN(_u10_u6_n2458 ) );
NAND2_X1 _u10_u6_U338  ( .A1(_u10_u6_n2460 ), .A2(_u10_u6_n2251 ), .ZN(_u10_u6_n2459 ) );
NAND3_X1 _u10_u6_U337  ( .A1(_u10_u6_n2457 ), .A2(_u10_u6_n2458 ), .A3(_u10_u6_n2459 ), .ZN(_u10_u6_n2448 ) );
NOR2_X1 _u10_u6_U336  ( .A1(_u10_u6_n2455 ), .A2(_u10_u6_n2456 ), .ZN(_u10_u6_n2449 ) );
NAND2_X1 _u10_u6_U335  ( .A1(_u10_u6_n2454 ), .A2(_u10_u6_n2438 ), .ZN(_u10_u6_n2452 ) );
NOR4_X1 _u10_u6_U334  ( .A1(_u10_u6_n2452 ), .A2(_u10_u6_n2453 ), .A3(_u10_u6_n2443 ), .A4(_u10_u6_n2143 ), .ZN(_u10_u6_n2451 ) );
NOR2_X1 _u10_u6_U333  ( .A1(_u10_u6_n2451 ), .A2(_u10_u6_n2356 ), .ZN(_u10_u6_n2450 ) );
NOR4_X1 _u10_u6_U332  ( .A1(_u10_u6_n2447 ), .A2(_u10_u6_n2448 ), .A3(_u10_u6_n2449 ), .A4(_u10_u6_n2450 ), .ZN(_u10_u6_n2390 ) );
NAND2_X1 _u10_u6_U331  ( .A1(_u10_u6_n2445 ), .A2(_u10_u6_n2446 ), .ZN(_u10_u6_n2155 ) );
INV_X1 _u10_u6_U330  ( .A(_u10_u6_n2155 ), .ZN(_u10_u6_n1892 ) );
INV_X1 _u10_u6_U329  ( .A(_u10_u6_n2444 ), .ZN(_u10_u6_n2088 ) );
NAND2_X1 _u10_u6_U328  ( .A1(_u10_u6_n1892 ), .A2(_u10_u6_n2088 ), .ZN(_u10_u6_n2337 ) );
NOR3_X1 _u10_u6_U327  ( .A1(_u10_u6_n2441 ), .A2(_u10_u6_n2442 ), .A3(_u10_u6_n2443 ), .ZN(_u10_u6_n2440 ) );
NAND4_X1 _u10_u6_U326  ( .A1(_u10_u6_n2193 ), .A2(_u10_u6_n2355 ), .A3(_u10_u6_n2439 ), .A4(_u10_u6_n2440 ), .ZN(_u10_u6_n2434 ) );
NAND3_X1 _u10_u6_U325  ( .A1(_u10_u6_n2437 ), .A2(_u10_u6_n2438 ), .A3(_u10_u6_n2059 ), .ZN(_u10_u6_n2435 ) );
NOR4_X1 _u10_u6_U324  ( .A1(_u10_u6_n2434 ), .A2(_u10_u6_n2435 ), .A3(_u10_u6_n1837 ), .A4(_u10_u6_n2436 ), .ZN(_u10_u6_n2433 ) );
NOR2_X1 _u10_u6_U323  ( .A1(_u10_u6_n2433 ), .A2(_u10_u6_n1836 ), .ZN(_u10_u6_n2415 ) );
INV_X1 _u10_u6_U322  ( .A(_u10_u6_n2432 ), .ZN(_u10_u6_n2178 ) );
NOR2_X1 _u10_u6_U321  ( .A1(_u10_u6_n1960 ), .A2(_u10_u6_n2431 ), .ZN(_u10_u6_n2430 ) );
NOR4_X1 _u10_u6_U320  ( .A1(_u10_u6_n2178 ), .A2(_u10_u6_n2429 ), .A3(_u10_u6_n2430 ), .A4(_u10_u6_n2179 ), .ZN(_u10_u6_n2416 ) );
NOR2_X1 _u10_u6_U319  ( .A1(_u10_u6_n2427 ), .A2(_u10_u6_n2428 ), .ZN(_u10_u6_n2426 ) );
NAND4_X1 _u10_u6_U318  ( .A1(_u10_u6_n2286 ), .A2(_u10_u6_n1969 ), .A3(_u10_u6_n2282 ), .A4(_u10_u6_n2426 ), .ZN(_u10_u6_n2425 ) );
NAND2_X1 _u10_u6_U317  ( .A1(_u10_u6_n2031 ), .A2(_u10_u6_n2425 ), .ZN(_u10_u6_n2422 ) );
NAND3_X1 _u10_u6_U316  ( .A1(_u10_u6_n2422 ), .A2(_u10_u6_n2423 ), .A3(_u10_u6_n2424 ), .ZN(_u10_u6_n2419 ) );
NOR4_X1 _u10_u6_U315  ( .A1(_u10_u6_n2419 ), .A2(_u10_u6_n1978 ), .A3(_u10_u6_n2420 ), .A4(_u10_u6_n2421 ), .ZN(_u10_u6_n2418 ) );
NOR2_X1 _u10_u6_U314  ( .A1(_u10_u6_n2418 ), .A2(_u10_u6_n2359 ), .ZN(_u10_u6_n2417 ) );
NOR3_X1 _u10_u6_U313  ( .A1(_u10_u6_n2415 ), .A2(_u10_u6_n2416 ), .A3(_u10_u6_n2417 ), .ZN(_u10_u6_n2414 ) );
NAND4_X1 _u10_u6_U312  ( .A1(_u10_u6_n2337 ), .A2(_u10_u6_n2412 ), .A3(_u10_u6_n2413 ), .A4(_u10_u6_n2414 ), .ZN(_u10_u6_n2392 ) );
NAND2_X1 _u10_u6_U311  ( .A1(_u10_u6_n2411 ), .A2(_u10_u6_n1936 ), .ZN(_u10_u6_n2410 ) );
NAND2_X1 _u10_u6_U310  ( .A1(_u10_u6_n2409 ), .A2(_u10_u6_n2410 ), .ZN(_u10_u6_n2408 ) );
NAND3_X1 _u10_u6_U309  ( .A1(_u10_u6_n2408 ), .A2(_u10_u6_n2305 ), .A3(_u10_u6_n1894 ), .ZN(_u10_u6_n2402 ) );
NAND3_X1 _u10_u6_U308  ( .A1(_u10_u6_n2329 ), .A2(_u10_u6_n2407 ), .A3(_u10_u6_n2255 ), .ZN(_u10_u6_n2403 ) );
NAND3_X1 _u10_u6_U307  ( .A1(_u10_u6_n1924 ), .A2(_u10_u6_n2405 ), .A3(_u10_u6_n2406 ), .ZN(_u10_u6_n2404 ) );
NAND3_X1 _u10_u6_U306  ( .A1(_u10_u6_n2402 ), .A2(_u10_u6_n2403 ), .A3(_u10_u6_n2404 ), .ZN(_u10_u6_n2393 ) );
INV_X1 _u10_u6_U305  ( .A(_u10_u6_n1932 ), .ZN(_u10_u6_n2399 ) );
NOR2_X1 _u10_u6_U304  ( .A1(_u10_u6_n2401 ), .A2(_u10_u6_n2161 ), .ZN(_u10_u6_n2400 ) );
NOR2_X1 _u10_u6_U303  ( .A1(_u10_u6_n2399 ), .A2(_u10_u6_n2400 ), .ZN(_u10_u6_n2394 ) );
NOR2_X1 _u10_u6_U302  ( .A1(_u10_u6_n2110 ), .A2(_u10_u6_n2398 ), .ZN(_u10_u6_n2397 ) );
NOR2_X1 _u10_u6_U301  ( .A1(_u10_u6_n2396 ), .A2(_u10_u6_n2397 ), .ZN(_u10_u6_n2395 ) );
NOR4_X1 _u10_u6_U300  ( .A1(_u10_u6_n2392 ), .A2(_u10_u6_n2393 ), .A3(_u10_u6_n2394 ), .A4(_u10_u6_n2395 ), .ZN(_u10_u6_n2391 ) );
NAND4_X1 _u10_u6_U299  ( .A1(_u10_u6_n2388 ), .A2(_u10_u6_n2389 ), .A3(_u10_u6_n2390 ), .A4(_u10_u6_n2391 ), .ZN(_u10_u6_n2387 ) );
MUX2_X1 _u10_u6_U298  ( .A(_u10_u6_n2387 ), .B(_u10_SYNOPSYS_UNCONNECTED_25 ), .S(_u10_u6_n1819 ), .Z(_u10_u6_n1810 ) );
NAND2_X1 _u10_u6_U297  ( .A1(_u10_u6_n2386 ), .A2(_u10_u6_n2007 ), .ZN(_u10_u6_n2369 ) );
AND2_X1 _u10_u6_U296  ( .A1(1'b0), .A2(_u10_u6_n2195 ), .ZN(_u10_u6_n2308 ));
NAND2_X1 _u10_u6_U295  ( .A1(_u10_u6_n2308 ), .A2(_u10_u6_n2036 ), .ZN(_u10_u6_n2384 ) );
AND2_X1 _u10_u6_U294  ( .A1(_u10_u6_n2384 ), .A2(_u10_u6_n2385 ), .ZN(_u10_u6_n2275 ) );
AND4_X1 _u10_u6_U293  ( .A1(_u10_u6_n2275 ), .A2(_u10_u6_n2286 ), .A3(_u10_u6_n2383 ), .A4(_u10_u6_n2285 ), .ZN(_u10_u6_n2225 ) );
NAND3_X1 _u10_u6_U292  ( .A1(_u10_u6_n2195 ), .A2(_u10_u6_n2223 ), .A3(1'b0),.ZN(_u10_u6_n2021 ) );
INV_X1 _u10_u6_U291  ( .A(_u10_u6_n2021 ), .ZN(_u10_u6_n2167 ) );
NAND2_X1 _u10_u6_U290  ( .A1(_u10_u6_n2036 ), .A2(_u10_u6_n2167 ), .ZN(_u10_u6_n1970 ) );
AND3_X1 _u10_u6_U289  ( .A1(_u10_u6_n1970 ), .A2(_u10_u6_n2164 ), .A3(_u10_u6_n2382 ), .ZN(_u10_u6_n2381 ) );
NAND4_X1 _u10_u6_U288  ( .A1(_u10_u6_n2225 ), .A2(_u10_u6_n2379 ), .A3(_u10_u6_n2380 ), .A4(_u10_u6_n2381 ), .ZN(_u10_u6_n2378 ) );
NAND2_X1 _u10_u6_U287  ( .A1(_u10_u6_n1967 ), .A2(_u10_u6_n2378 ), .ZN(_u10_u6_n2370 ) );
NAND2_X1 _u10_u6_U286  ( .A1(_u10_u6_n2081 ), .A2(_u10_u6_n2377 ), .ZN(_u10_u6_n2371 ) );
NOR2_X1 _u10_u6_U285  ( .A1(_u10_u6_n2375 ), .A2(_u10_u6_n2376 ), .ZN(_u10_u6_n2373 ) );
NOR2_X1 _u10_u6_U284  ( .A1(_u10_u6_n2373 ), .A2(_u10_u6_n2374 ), .ZN(_u10_u6_n2372 ) );
NAND4_X1 _u10_u6_U283  ( .A1(_u10_u6_n2369 ), .A2(_u10_u6_n2370 ), .A3(_u10_u6_n2371 ), .A4(_u10_u6_n2372 ), .ZN(_u10_u6_n2309 ) );
NOR2_X1 _u10_u6_U282  ( .A1(_u10_u6_n2000 ), .A2(_u10_u6_n2368 ), .ZN(_u10_u6_n2360 ) );
NOR2_X1 _u10_u6_U281  ( .A1(_u10_u6_n2366 ), .A2(_u10_u6_n2367 ), .ZN(_u10_u6_n2361 ) );
NOR2_X1 _u10_u6_U280  ( .A1(_u10_u6_n1868 ), .A2(_u10_u6_n2365 ), .ZN(_u10_u6_n2362 ) );
NOR2_X1 _u10_u6_U279  ( .A1(_u10_u6_n2364 ), .A2(_u10_u6_n1859 ), .ZN(_u10_u6_n2363 ) );
NOR4_X1 _u10_u6_U278  ( .A1(_u10_u6_n2360 ), .A2(_u10_u6_n2361 ), .A3(_u10_u6_n2362 ), .A4(_u10_u6_n2363 ), .ZN(_u10_u6_n2316 ) );
NOR2_X1 _u10_u6_U277  ( .A1(_u10_u6_n2359 ), .A2(_u10_u6_n1970 ), .ZN(_u10_u6_n2351 ) );
NOR2_X1 _u10_u6_U276  ( .A1(_u10_u6_n2358 ), .A2(_u10_u6_n1840 ), .ZN(_u10_u6_n2352 ) );
NOR2_X1 _u10_u6_U275  ( .A1(_u10_u6_n2356 ), .A2(_u10_u6_n2357 ), .ZN(_u10_u6_n2353 ) );
NOR2_X1 _u10_u6_U274  ( .A1(_u10_u6_n1836 ), .A2(_u10_u6_n2355 ), .ZN(_u10_u6_n2354 ) );
NOR4_X1 _u10_u6_U273  ( .A1(_u10_u6_n2351 ), .A2(_u10_u6_n2352 ), .A3(_u10_u6_n2353 ), .A4(_u10_u6_n2354 ), .ZN(_u10_u6_n2317 ) );
NOR2_X1 _u10_u6_U272  ( .A1(_u10_u6_n1873 ), .A2(_u10_u6_n2101 ), .ZN(_u10_u6_n2349 ) );
NOR2_X1 _u10_u6_U271  ( .A1(_u10_u6_n2349 ), .A2(_u10_u6_n2350 ), .ZN(_u10_u6_n2338 ) );
NOR2_X1 _u10_u6_U270  ( .A1(_u10_u6_n2347 ), .A2(_u10_u6_n2348 ), .ZN(_u10_u6_n2345 ) );
NOR2_X1 _u10_u6_U269  ( .A1(_u10_u6_n2345 ), .A2(_u10_u6_n2346 ), .ZN(_u10_u6_n2339 ) );
NOR2_X1 _u10_u6_U268  ( .A1(_u10_u6_n2344 ), .A2(_u10_u6_n2142 ), .ZN(_u10_u6_n2340 ) );
NOR2_X1 _u10_u6_U267  ( .A1(_u10_u6_n2342 ), .A2(_u10_u6_n2343 ), .ZN(_u10_u6_n2341 ) );
NOR4_X1 _u10_u6_U266  ( .A1(_u10_u6_n2338 ), .A2(_u10_u6_n2339 ), .A3(_u10_u6_n2340 ), .A4(_u10_u6_n2341 ), .ZN(_u10_u6_n2318 ) );
INV_X1 _u10_u6_U265  ( .A(_u10_u6_n2337 ), .ZN(_u10_u6_n2320 ) );
NOR2_X1 _u10_u6_U264  ( .A1(_u10_u6_n1970 ), .A2(1'b0), .ZN(_u10_u6_n2027 ));
INV_X1 _u10_u6_U263  ( .A(_u10_u6_n2027 ), .ZN(_u10_u6_n2331 ) );
NOR2_X1 _u10_u6_U262  ( .A1(_u10_u6_n2174 ), .A2(_u10_u6_n2216 ), .ZN(_u10_u6_n2333 ) );
AND2_X1 _u10_u6_U261  ( .A1(_u10_u6_n1928 ), .A2(_u10_u6_n2336 ), .ZN(_u10_u6_n2334 ) );
NOR4_X1 _u10_u6_U260  ( .A1(_u10_u6_n1937 ), .A2(_u10_u6_n2333 ), .A3(_u10_u6_n2334 ), .A4(_u10_u6_n2335 ), .ZN(_u10_u6_n2332 ) );
NOR3_X1 _u10_u6_U259  ( .A1(_u10_u6_n2331 ), .A2(_u10_u6_n2332 ), .A3(_u10_u6_n1915 ), .ZN(_u10_u6_n2321 ) );
NOR3_X1 _u10_u6_U258  ( .A1(_u10_u6_n2291 ), .A2(_u10_u6_n2330 ), .A3(_u10_u6_n2021 ), .ZN(_u10_u6_n2322 ) );
NOR2_X1 _u10_u6_U257  ( .A1(_u10_u6_n2329 ), .A2(_u10_u6_n2169 ), .ZN(_u10_u6_n2324 ) );
NOR2_X1 _u10_u6_U256  ( .A1(1'b0), .A2(_u10_u6_n2328 ), .ZN(_u10_u6_n2327 ));
NOR2_X1 _u10_u6_U255  ( .A1(_u10_u6_n2326 ), .A2(_u10_u6_n2327 ), .ZN(_u10_u6_n2325 ) );
NOR3_X1 _u10_u6_U254  ( .A1(_u10_u6_n2324 ), .A2(1'b0), .A3(_u10_u6_n2325 ),.ZN(_u10_u6_n2323 ) );
NOR4_X1 _u10_u6_U253  ( .A1(_u10_u6_n2320 ), .A2(_u10_u6_n2321 ), .A3(_u10_u6_n2322 ), .A4(_u10_u6_n2323 ), .ZN(_u10_u6_n2319 ) );
AND4_X1 _u10_u6_U252  ( .A1(_u10_u6_n2316 ), .A2(_u10_u6_n2317 ), .A3(_u10_u6_n2318 ), .A4(_u10_u6_n2319 ), .ZN(_u10_u6_n1991 ) );
INV_X1 _u10_u6_U251  ( .A(_u10_u6_n2315 ), .ZN(_u10_u6_n2313 ) );
NAND3_X1 _u10_u6_U250  ( .A1(_u10_u6_n1991 ), .A2(_u10_u6_n2313 ), .A3(_u10_u6_n2314 ), .ZN(_u10_u6_n2310 ) );
NOR4_X1 _u10_u6_U249  ( .A1(_u10_u6_n2309 ), .A2(_u10_u6_n2310 ), .A3(_u10_u6_n2311 ), .A4(_u10_u6_n2312 ), .ZN(_u10_u6_n2117 ) );
NAND3_X1 _u10_u6_U248  ( .A1(_u10_u6_n2108 ), .A2(_u10_u6_n2107 ), .A3(_u10_u6_n2308 ), .ZN(_u10_u6_n2217 ) );
NOR3_X1 _u10_u6_U247  ( .A1(_u10_u6_n2306 ), .A2(_u10_u6_n2307 ), .A3(_u10_u6_n2027 ), .ZN(_u10_u6_n2277 ) );
NAND3_X1 _u10_u6_U246  ( .A1(_u10_u6_n2217 ), .A2(_u10_u6_n2305 ), .A3(_u10_u6_n2277 ), .ZN(_u10_u6_n2157 ) );
NAND2_X1 _u10_u6_U245  ( .A1(_u10_u6_n2089 ), .A2(_u10_u6_n2157 ), .ZN(_u10_u6_n2296 ) );
INV_X1 _u10_u6_U244  ( .A(_u10_u6_n2304 ), .ZN(_u10_u6_n2297 ) );
NOR2_X1 _u10_u6_U243  ( .A1(_u10_u6_n2302 ), .A2(_u10_u6_n2303 ), .ZN(_u10_u6_n2299 ) );
NOR3_X1 _u10_u6_U242  ( .A1(_u10_u6_n2299 ), .A2(_u10_u6_n2300 ), .A3(_u10_u6_n2301 ), .ZN(_u10_u6_n2298 ) );
NAND4_X1 _u10_u6_U241  ( .A1(_u10_u6_n2295 ), .A2(_u10_u6_n2296 ), .A3(_u10_u6_n2297 ), .A4(_u10_u6_n2298 ), .ZN(_u10_u6_n2294 ) );
NAND2_X1 _u10_u6_U240  ( .A1(_u10_u6_n2293 ), .A2(_u10_u6_n2294 ), .ZN(_u10_u6_n2257 ) );
NAND2_X1 _u10_u6_U239  ( .A1(_u10_u6_n2165 ), .A2(_u10_u6_n2166 ), .ZN(_u10_u6_n2288 ) );
NAND2_X1 _u10_u6_U238  ( .A1(_u10_u6_n2078 ), .A2(_u10_u6_n2279 ), .ZN(_u10_u6_n2292 ) );
NAND2_X1 _u10_u6_U237  ( .A1(_u10_u6_n2291 ), .A2(_u10_u6_n2292 ), .ZN(_u10_u6_n2290 ) );
NAND2_X1 _u10_u6_U236  ( .A1(_u10_u6_n2059 ), .A2(_u10_u6_n2290 ), .ZN(_u10_u6_n2289 ) );
NAND2_X1 _u10_u6_U235  ( .A1(_u10_u6_n2288 ), .A2(_u10_u6_n2289 ), .ZN(_u10_u6_n2201 ) );
NAND2_X1 _u10_u6_U234  ( .A1(1'b0), .A2(_u10_u6_n2201 ), .ZN(_u10_u6_n2258 ));
INV_X1 _u10_u6_U233  ( .A(_u10_u6_n2287 ), .ZN(_u10_u6_n2283 ) );
AND4_X1 _u10_u6_U232  ( .A1(_u10_u6_n2285 ), .A2(_u10_u6_n2226 ), .A3(_u10_u6_n1970 ), .A4(_u10_u6_n2286 ), .ZN(_u10_u6_n2284 ) );
NAND4_X1 _u10_u6_U231  ( .A1(_u10_u6_n2281 ), .A2(_u10_u6_n2282 ), .A3(_u10_u6_n2283 ), .A4(_u10_u6_n2284 ), .ZN(_u10_u6_n2280 ) );
NAND2_X1 _u10_u6_U230  ( .A1(_u10_u6_n2279 ), .A2(_u10_u6_n2280 ), .ZN(_u10_u6_n2259 ) );
NAND4_X1 _u10_u6_U229  ( .A1(_u10_u6_n2275 ), .A2(_u10_u6_n2276 ), .A3(_u10_u6_n2277 ), .A4(_u10_u6_n2278 ), .ZN(_u10_u6_n2271 ) );
NAND2_X1 _u10_u6_U228  ( .A1(_u10_u6_n1933 ), .A2(_u10_u6_n2164 ), .ZN(_u10_u6_n2272 ) );
NOR2_X1 _u10_u6_U227  ( .A1(_u10_u6_n2274 ), .A2(_u10_u6_n2130 ), .ZN(_u10_u6_n2273 ) );
NOR4_X1 _u10_u6_U226  ( .A1(_u10_u6_n2271 ), .A2(_u10_u6_n2272 ), .A3(_u10_u6_n1978 ), .A4(_u10_u6_n2273 ), .ZN(_u10_u6_n2270 ) );
NOR2_X1 _u10_u6_U225  ( .A1(_u10_u6_n2270 ), .A2(_u10_u6_n2025 ), .ZN(_u10_u6_n2261 ) );
NAND3_X1 _u10_u6_U224  ( .A1(_u10_u6_n1933 ), .A2(_u10_u6_n1936 ), .A3(_u10_u6_n2269 ), .ZN(_u10_u6_n2268 ) );
NOR3_X1 _u10_u6_U223  ( .A1(_u10_u6_n2268 ), .A2(_u10_u6_n1844 ), .A3(_u10_u6_n2157 ), .ZN(_u10_u6_n2267 ) );
NOR2_X1 _u10_u6_U222  ( .A1(1'b0), .A2(_u10_u6_n2267 ), .ZN(_u10_u6_n2265 ));
NOR3_X1 _u10_u6_U221  ( .A1(_u10_u6_n2264 ), .A2(_u10_u6_n2265 ), .A3(_u10_u6_n2266 ), .ZN(_u10_u6_n2263 ) );
NOR2_X1 _u10_u6_U220  ( .A1(_u10_u6_n2263 ), .A2(_u10_u6_n1843 ), .ZN(_u10_u6_n2262 ) );
NOR2_X1 _u10_u6_U219  ( .A1(_u10_u6_n2261 ), .A2(_u10_u6_n2262 ), .ZN(_u10_u6_n2260 ) );
NAND4_X1 _u10_u6_U218  ( .A1(_u10_u6_n2257 ), .A2(_u10_u6_n2258 ), .A3(_u10_u6_n2259 ), .A4(_u10_u6_n2260 ), .ZN(_u10_u6_n2230 ) );
INV_X1 _u10_u6_U217  ( .A(_u10_u6_n2217 ), .ZN(_u10_u6_n2242 ) );
NAND2_X1 _u10_u6_U216  ( .A1(_u10_u6_n2168 ), .A2(_u10_u6_n2169 ), .ZN(_u10_u6_n2244 ) );
NAND2_X1 _u10_u6_U215  ( .A1(_u10_u6_n2255 ), .A2(_u10_u6_n2256 ), .ZN(_u10_u6_n2245 ) );
NAND2_X1 _u10_u6_U214  ( .A1(_u10_u6_n2253 ), .A2(_u10_u6_n2254 ), .ZN(_u10_u6_n2252 ) );
NAND2_X1 _u10_u6_U213  ( .A1(_u10_u6_n2251 ), .A2(_u10_u6_n2252 ), .ZN(_u10_u6_n2246 ) );
NAND2_X1 _u10_u6_U212  ( .A1(_u10_u6_n2152 ), .A2(_u10_u6_n1928 ), .ZN(_u10_u6_n2250 ) );
NAND2_X1 _u10_u6_U211  ( .A1(_u10_u6_n2249 ), .A2(_u10_u6_n2250 ), .ZN(_u10_u6_n2248 ) );
NAND2_X1 _u10_u6_U210  ( .A1(_u10_u6_n2105 ), .A2(_u10_u6_n2248 ), .ZN(_u10_u6_n2247 ) );
NAND4_X1 _u10_u6_U209  ( .A1(_u10_u6_n2244 ), .A2(_u10_u6_n2245 ), .A3(_u10_u6_n2246 ), .A4(_u10_u6_n2247 ), .ZN(_u10_u6_n2243 ) );
NAND2_X1 _u10_u6_U208  ( .A1(_u10_u6_n2242 ), .A2(_u10_u6_n2243 ), .ZN(_u10_u6_n2237 ) );
NAND2_X1 _u10_u6_U207  ( .A1(1'b0), .A2(_u10_u6_n2241 ), .ZN(_u10_u6_n2238 ));
NAND2_X1 _u10_u6_U206  ( .A1(_u10_u6_n2214 ), .A2(_u10_u6_n2240 ), .ZN(_u10_u6_n2239 ) );
NAND3_X1 _u10_u6_U205  ( .A1(_u10_u6_n2237 ), .A2(_u10_u6_n2238 ), .A3(_u10_u6_n2239 ), .ZN(_u10_u6_n2231 ) );
AND2_X1 _u10_u6_U204  ( .A1(_u10_u6_n2200 ), .A2(_u10_u6_n2236 ), .ZN(_u10_u6_n2232 ) );
NOR2_X1 _u10_u6_U203  ( .A1(_u10_u6_n2234 ), .A2(_u10_u6_n2235 ), .ZN(_u10_u6_n2233 ) );
NOR4_X1 _u10_u6_U202  ( .A1(_u10_u6_n2230 ), .A2(_u10_u6_n2231 ), .A3(_u10_u6_n2232 ), .A4(_u10_u6_n2233 ), .ZN(_u10_u6_n2118 ) );
NAND2_X1 _u10_u6_U201  ( .A1(_u10_u6_n2214 ), .A2(_u10_u6_n2049 ), .ZN(_u10_u6_n2229 ) );
NAND2_X1 _u10_u6_U200  ( .A1(_u10_u6_n2228 ), .A2(_u10_u6_n2229 ), .ZN(_u10_u6_n2227 ) );
NAND2_X1 _u10_u6_U199  ( .A1(_u10_u6_n2043 ), .A2(_u10_u6_n2227 ), .ZN(_u10_u6_n2204 ) );
NAND2_X1 _u10_u6_U198  ( .A1(_u10_u6_n2225 ), .A2(_u10_u6_n2226 ), .ZN(_u10_u6_n2224 ) );
NAND2_X1 _u10_u6_U197  ( .A1(_u10_u6_n1899 ), .A2(_u10_u6_n2224 ), .ZN(_u10_u6_n2205 ) );
NAND2_X1 _u10_u6_U196  ( .A1(_u10_u6_n2222 ), .A2(_u10_u6_n2223 ), .ZN(_u10_u6_n1870 ) );
NAND4_X1 _u10_u6_U195  ( .A1(_u10_u6_n2220 ), .A2(_u10_u6_n2131 ), .A3(_u10_u6_n2221 ), .A4(_u10_u6_n1870 ), .ZN(_u10_u6_n2219 ) );
NAND2_X1 _u10_u6_U194  ( .A1(_u10_u6_n2218 ), .A2(_u10_u6_n2219 ), .ZN(_u10_u6_n2206 ) );
NOR2_X1 _u10_u6_U193  ( .A1(_u10_u6_n1925 ), .A2(_u10_u6_n2217 ), .ZN(_u10_u6_n2215 ) );
NOR4_X1 _u10_u6_U192  ( .A1(_u10_u6_n2213 ), .A2(_u10_u6_n2214 ), .A3(_u10_u6_n2215 ), .A4(_u10_u6_n2216 ), .ZN(_u10_u6_n2211 ) );
NOR2_X1 _u10_u6_U191  ( .A1(_u10_u6_n2211 ), .A2(_u10_u6_n2212 ), .ZN(_u10_u6_n2208 ) );
NOR2_X1 _u10_u6_U190  ( .A1(_u10_u6_n1888 ), .A2(_u10_u6_n2210 ), .ZN(_u10_u6_n2209 ) );
NOR2_X1 _u10_u6_U189  ( .A1(_u10_u6_n2208 ), .A2(_u10_u6_n2209 ), .ZN(_u10_u6_n2207 ) );
NAND4_X1 _u10_u6_U188  ( .A1(_u10_u6_n2204 ), .A2(_u10_u6_n2205 ), .A3(_u10_u6_n2206 ), .A4(_u10_u6_n2207 ), .ZN(_u10_u6_n2170 ) );
OR2_X1 _u10_u6_U187  ( .A1(_u10_u6_n2202 ), .A2(_u10_u6_n2203 ), .ZN(_u10_u6_n2197 ) );
NAND2_X1 _u10_u6_U186  ( .A1(1'b0), .A2(_u10_u6_n2201 ), .ZN(_u10_u6_n2198 ));
NAND2_X1 _u10_u6_U185  ( .A1(_u10_u6_n2063 ), .A2(_u10_u6_n2200 ), .ZN(_u10_u6_n2199 ) );
NAND3_X1 _u10_u6_U184  ( .A1(_u10_u6_n2197 ), .A2(_u10_u6_n2198 ), .A3(_u10_u6_n2199 ), .ZN(_u10_u6_n2196 ) );
NAND2_X1 _u10_u6_U183  ( .A1(_u10_u6_n2195 ), .A2(_u10_u6_n2196 ), .ZN(_u10_u6_n2180 ) );
NAND2_X1 _u10_u6_U182  ( .A1(_u10_u6_n2195 ), .A2(_u10_u6_n1918 ), .ZN(_u10_u6_n2192 ) );
NAND4_X1 _u10_u6_U181  ( .A1(_u10_u6_n2192 ), .A2(_u10_u6_n2021 ), .A3(_u10_u6_n2193 ), .A4(_u10_u6_n2194 ), .ZN(_u10_u6_n2188 ) );
NAND2_X1 _u10_u6_U180  ( .A1(_u10_u6_n2188 ), .A2(_u10_u6_n2191 ), .ZN(_u10_u6_n2181 ) );
NAND2_X1 _u10_u6_U179  ( .A1(1'b0), .A2(_u10_u6_n2190 ), .ZN(_u10_u6_n2185 ));
NAND2_X1 _u10_u6_U178  ( .A1(_u10_u6_n2189 ), .A2(_u10_SYNOPSYS_UNCONNECTED_26 ), .ZN(_u10_u6_n2186 ) );
INV_X1 _u10_u6_U177  ( .A(_u10_u6_n2188 ), .ZN(_u10_u6_n2187 ) );
NAND3_X1 _u10_u6_U176  ( .A1(_u10_u6_n2185 ), .A2(_u10_u6_n2186 ), .A3(_u10_u6_n2187 ), .ZN(_u10_u6_n2184 ) );
NAND2_X1 _u10_u6_U175  ( .A1(_u10_u6_n2183 ), .A2(_u10_u6_n2184 ), .ZN(_u10_u6_n2182 ) );
NAND3_X1 _u10_u6_U174  ( .A1(_u10_u6_n2180 ), .A2(_u10_u6_n2181 ), .A3(_u10_u6_n2182 ), .ZN(_u10_u6_n2171 ) );
INV_X1 _u10_u6_U173  ( .A(_u10_u6_n2179 ), .ZN(_u10_u6_n1963 ) );
NOR2_X1 _u10_u6_U172  ( .A1(_u10_u6_n1963 ), .A2(_u10_u6_n2178 ), .ZN(_u10_u6_n2172 ) );
INV_X1 _u10_u6_U171  ( .A(_u10_u6_n2177 ), .ZN(_u10_u6_n2176 ) );
NOR3_X1 _u10_u6_U170  ( .A1(_u10_u6_n2174 ), .A2(_u10_u6_n2175 ), .A3(_u10_u6_n2176 ), .ZN(_u10_u6_n2173 ) );
NOR4_X1 _u10_u6_U169  ( .A1(_u10_u6_n2170 ), .A2(_u10_u6_n2171 ), .A3(_u10_u6_n2172 ), .A4(_u10_u6_n2173 ), .ZN(_u10_u6_n2119 ) );
NAND3_X1 _u10_u6_U168  ( .A1(_u10_u6_n2168 ), .A2(_u10_u6_n2169 ), .A3(1'b0),.ZN(_u10_u6_n2148 ) );
NAND3_X1 _u10_u6_U167  ( .A1(_u10_u6_n2165 ), .A2(_u10_u6_n2166 ), .A3(_u10_u6_n2167 ), .ZN(_u10_u6_n2149 ) );
NAND4_X1 _u10_u6_U166  ( .A1(_u10_u6_n2162 ), .A2(_u10_u6_n1933 ), .A3(_u10_u6_n2163 ), .A4(_u10_u6_n2164 ), .ZN(_u10_u6_n2160 ) );
NOR4_X1 _u10_u6_U165  ( .A1(_u10_u6_n2160 ), .A2(_u10_u6_n2157 ), .A3(_u10_u6_n1844 ), .A4(_u10_u6_n2161 ), .ZN(_u10_u6_n2158 ) );
NOR2_X1 _u10_u6_U164  ( .A1(_u10_u6_n2158 ), .A2(_u10_u6_n2159 ), .ZN(_u10_u6_n2153 ) );
INV_X1 _u10_u6_U163  ( .A(_u10_u6_n2157 ), .ZN(_u10_u6_n2129 ) );
NOR3_X1 _u10_u6_U162  ( .A1(_u10_u6_n2155 ), .A2(_u10_u6_n2129 ), .A3(_u10_u6_n2156 ), .ZN(_u10_u6_n2154 ) );
NOR2_X1 _u10_u6_U161  ( .A1(_u10_u6_n2153 ), .A2(_u10_u6_n2154 ), .ZN(_u10_u6_n2150 ) );
NAND3_X1 _u10_u6_U160  ( .A1(1'b0), .A2(_u10_u6_n1928 ), .A3(_u10_u6_n2152 ),.ZN(_u10_u6_n2151 ) );
NAND4_X1 _u10_u6_U159  ( .A1(_u10_u6_n2148 ), .A2(_u10_u6_n2149 ), .A3(_u10_u6_n2150 ), .A4(_u10_u6_n2151 ), .ZN(_u10_u6_n2121 ) );
NAND2_X1 _u10_u6_U158  ( .A1(_u10_u6_n2107 ), .A2(_u10_u6_n2147 ), .ZN(_u10_u6_n2146 ) );
NAND2_X1 _u10_u6_U157  ( .A1(_u10_u6_n2145 ), .A2(_u10_u6_n2146 ), .ZN(_u10_u6_n2144 ) );
NAND2_X1 _u10_u6_U156  ( .A1(_u10_u6_n2143 ), .A2(_u10_u6_n2144 ), .ZN(_u10_u6_n2134 ) );
NAND2_X1 _u10_u6_U155  ( .A1(_u10_u6_n2141 ), .A2(_u10_u6_n2142 ), .ZN(_u10_u6_n2140 ) );
NAND2_X1 _u10_u6_U154  ( .A1(_u10_u6_n2139 ), .A2(_u10_u6_n2140 ), .ZN(_u10_u6_n2135 ) );
OR2_X1 _u10_u6_U153  ( .A1(_u10_u6_n2110 ), .A2(_u10_u6_n1911 ), .ZN(_u10_u6_n2137 ) );
NAND2_X1 _u10_u6_U152  ( .A1(_u10_u6_n2137 ), .A2(_u10_u6_n2138 ), .ZN(_u10_u6_n2136 ) );
NAND3_X1 _u10_u6_U151  ( .A1(_u10_u6_n2134 ), .A2(_u10_u6_n2135 ), .A3(_u10_u6_n2136 ), .ZN(_u10_u6_n2122 ) );
NOR2_X1 _u10_u6_U150  ( .A1(_u10_u6_n2133 ), .A2(_u10_u6_n1891 ), .ZN(_u10_u6_n2132 ) );
NOR2_X1 _u10_u6_U149  ( .A1(_u10_u6_n2131 ), .A2(_u10_u6_n2132 ), .ZN(_u10_u6_n2123 ) );
NOR2_X1 _u10_u6_U148  ( .A1(_u10_u6_n2129 ), .A2(_u10_u6_n2130 ), .ZN(_u10_u6_n2127 ) );
NOR2_X1 _u10_u6_U147  ( .A1(_u10_u6_n2127 ), .A2(_u10_u6_n2128 ), .ZN(_u10_u6_n2125 ) );
NOR2_X1 _u10_u6_U146  ( .A1(_u10_u6_n2125 ), .A2(_u10_u6_n2126 ), .ZN(_u10_u6_n2124 ) );
NOR4_X1 _u10_u6_U145  ( .A1(_u10_u6_n2121 ), .A2(_u10_u6_n2122 ), .A3(_u10_u6_n2123 ), .A4(_u10_u6_n2124 ), .ZN(_u10_u6_n2120 ) );
NAND4_X1 _u10_u6_U144  ( .A1(_u10_u6_n2117 ), .A2(_u10_u6_n2118 ), .A3(_u10_u6_n2119 ), .A4(_u10_u6_n2120 ), .ZN(_u10_u6_n2116 ) );
MUX2_X1 _u10_u6_U143  ( .A(_u10_u6_n2116 ), .B(_u10_SYNOPSYS_UNCONNECTED_26 ), .S(_u10_u6_n1819 ), .Z(_u10_u6_n1811 ) );
INV_X1 _u10_u6_U142  ( .A(_u10_u6_n2115 ), .ZN(_u10_u6_n2006 ) );
NOR3_X1 _u10_u6_U141  ( .A1(_u10_u6_n2006 ), .A2(_u10_u6_n2114 ), .A3(_u10_u6_n2081 ), .ZN(_u10_u6_n1854 ) );
NAND2_X1 _u10_u6_U140  ( .A1(_u10_u6_n2112 ), .A2(_u10_u6_n2113 ), .ZN(_u10_u6_n1872 ) );
INV_X1 _u10_u6_U139  ( .A(_u10_u6_n1872 ), .ZN(_u10_u6_n1882 ) );
NAND4_X1 _u10_u6_U138  ( .A1(_u10_u6_n1854 ), .A2(_u10_u6_n1882 ), .A3(_u10_u6_n2111 ), .A4(_u10_u6_n1868 ), .ZN(_u10_u6_n2109 ) );
NAND2_X1 _u10_u6_U137  ( .A1(_u10_u6_n2109 ), .A2(_u10_u6_n2110 ), .ZN(_u10_u6_n2098 ) );
NAND2_X1 _u10_u6_U136  ( .A1(1'b0), .A2(_u10_u6_n1983 ), .ZN(_u10_u6_n2023 ));
INV_X1 _u10_u6_U135  ( .A(_u10_u6_n2023 ), .ZN(_u10_u6_n2035 ) );
NAND3_X1 _u10_u6_U134  ( .A1(_u10_u6_n2035 ), .A2(_u10_u6_n2107 ), .A3(_u10_u6_n2108 ), .ZN(_u10_u6_n1916 ) );
INV_X1 _u10_u6_U133  ( .A(_u10_u6_n1916 ), .ZN(_u10_u6_n2093 ) );
NAND3_X1 _u10_u6_U132  ( .A1(_u10_u6_n2105 ), .A2(_u10_u6_n2106 ), .A3(_u10_u6_n2093 ), .ZN(_u10_u6_n2039 ) );
NAND2_X1 _u10_u6_U131  ( .A1(_u10_u6_n2039 ), .A2(_u10_u6_n1930 ), .ZN(_u10_u6_n2104 ) );
NAND2_X1 _u10_u6_U130  ( .A1(_u10_u6_n2103 ), .A2(_u10_u6_n2104 ), .ZN(_u10_u6_n1863 ) );
OR2_X1 _u10_u6_U129  ( .A1(_u10_u6_n1863 ), .A2(_u10_u6_n2102 ), .ZN(_u10_u6_n2099 ) );
NAND2_X1 _u10_u6_U128  ( .A1(_u10_u6_n1890 ), .A2(_u10_u6_n2101 ), .ZN(_u10_u6_n2100 ) );
NAND3_X1 _u10_u6_U127  ( .A1(_u10_u6_n2098 ), .A2(_u10_u6_n2099 ), .A3(_u10_u6_n2100 ), .ZN(_u10_u6_n2066 ) );
NAND4_X1 _u10_u6_U126  ( .A1(_u10_u6_n2095 ), .A2(_u10_u6_n2096 ), .A3(_u10_u6_n1896 ), .A4(_u10_u6_n2097 ), .ZN(_u10_u6_n2086 ) );
NOR4_X1 _u10_u6_U125  ( .A1(_u10_u6_n2093 ), .A2(_u10_u6_n2027 ), .A3(_u10_u6_n2094 ), .A4(_u10_u6_n2026 ), .ZN(_u10_u6_n1952 ) );
NOR2_X1 _u10_u6_U124  ( .A1(1'b0), .A2(_u10_u6_n1952 ), .ZN(_u10_u6_n1951 ));
INV_X1 _u10_u6_U123  ( .A(_u10_u6_n1951 ), .ZN(_u10_u6_n2090 ) );
NAND4_X1 _u10_u6_U122  ( .A1(_u10_u6_n2089 ), .A2(_u10_u6_n2090 ), .A3(_u10_u6_n2091 ), .A4(_u10_u6_n2092 ), .ZN(_u10_u6_n1893 ) );
NOR4_X1 _u10_u6_U121  ( .A1(_u10_u6_n2086 ), .A2(_u10_u6_n1893 ), .A3(_u10_u6_n2087 ), .A4(_u10_u6_n2088 ), .ZN(_u10_u6_n2084 ) );
NOR2_X1 _u10_u6_U120  ( .A1(_u10_u6_n2084 ), .A2(_u10_u6_n2085 ), .ZN(_u10_u6_n2067 ) );
NOR2_X1 _u10_u6_U119  ( .A1(_u10_u6_n2083 ), .A2(_u10_u6_n1869 ), .ZN(_u10_u6_n2068 ) );
NAND2_X1 _u10_u6_U118  ( .A1(_u10_u6_n2081 ), .A2(_u10_u6_n2082 ), .ZN(_u10_u6_n2075 ) );
NAND2_X1 _u10_u6_U117  ( .A1(_u10_u6_n2035 ), .A2(_u10_u6_n2019 ), .ZN(_u10_u6_n2060 ) );
NAND2_X1 _u10_u6_U116  ( .A1(_u10_u6_n2080 ), .A2(_u10_u6_n2060 ), .ZN(_u10_u6_n2079 ) );
NAND2_X1 _u10_u6_U115  ( .A1(_u10_u6_n2078 ), .A2(_u10_u6_n2079 ), .ZN(_u10_u6_n2076 ) );
NAND4_X1 _u10_u6_U114  ( .A1(_u10_u6_n2075 ), .A2(_u10_u6_n2076 ), .A3(_u10_u6_n1970 ), .A4(_u10_u6_n2077 ), .ZN(_u10_u6_n2072 ) );
NOR4_X1 _u10_u6_U113  ( .A1(_u10_u6_n2072 ), .A2(_u10_u6_n2073 ), .A3(_u10_u6_n1975 ), .A4(_u10_u6_n2074 ), .ZN(_u10_u6_n2070 ) );
NOR2_X1 _u10_u6_U112  ( .A1(_u10_u6_n2070 ), .A2(_u10_u6_n2071 ), .ZN(_u10_u6_n2069 ) );
NOR4_X1 _u10_u6_U111  ( .A1(_u10_u6_n2066 ), .A2(_u10_u6_n2067 ), .A3(_u10_u6_n2068 ), .A4(_u10_u6_n2069 ), .ZN(_u10_u6_n1820 ) );
NAND2_X1 _u10_u6_U110  ( .A1(1'b0), .A2(_u10_u6_n1983 ), .ZN(_u10_u6_n2065 ));
NAND4_X1 _u10_u6_U109  ( .A1(_u10_u6_n2065 ), .A2(_u10_u6_n2023 ), .A3(_u10_u6_n2021 ), .A4(_u10_u6_n2052 ), .ZN(_u10_u6_n2064 ) );
NAND2_X1 _u10_u6_U108  ( .A1(_u10_u6_n2063 ), .A2(_u10_u6_n2064 ), .ZN(_u10_u6_n2040 ) );
NAND4_X1 _u10_u6_U107  ( .A1(_u10_u6_n2059 ), .A2(_u10_u6_n2060 ), .A3(_u10_u6_n2061 ), .A4(_u10_u6_n2062 ), .ZN(_u10_u6_n2058 ) );
NAND2_X1 _u10_u6_U106  ( .A1(_u10_u6_n2057 ), .A2(_u10_u6_n2058 ), .ZN(_u10_u6_n2041 ) );
NOR4_X1 _u10_u6_U105  ( .A1(1'b0), .A2(_u10_u6_n2054 ), .A3(_u10_u6_n2055 ),.A4(_u10_u6_n2056 ), .ZN(_u10_u6_n2053 ) );
NAND4_X1 _u10_u6_U104  ( .A1(_u10_u6_n2021 ), .A2(_u10_u6_n2052 ), .A3(_u10_u6_n2023 ), .A4(_u10_u6_n2053 ), .ZN(_u10_u6_n1964 ) );
INV_X1 _u10_u6_U103  ( .A(_u10_u6_n1964 ), .ZN(_u10_u6_n2045 ) );
NAND2_X1 _u10_u6_U102  ( .A1(_u10_u6_n2051 ), .A2(_u10_SYNOPSYS_UNCONNECTED_27 ), .ZN(_u10_u6_n2046 ) );
NAND2_X1 _u10_u6_U101  ( .A1(_u10_u6_n2049 ), .A2(_u10_u6_n2050 ), .ZN(_u10_u6_n2047 ) );
NAND4_X1 _u10_u6_U100  ( .A1(_u10_u6_n2045 ), .A2(_u10_u6_n2046 ), .A3(_u10_u6_n2047 ), .A4(_u10_u6_n2048 ), .ZN(_u10_u6_n2044 ) );
NAND2_X1 _u10_u6_U99  ( .A1(_u10_u6_n2043 ), .A2(_u10_u6_n2044 ), .ZN(_u10_u6_n2042 ) );
NAND3_X1 _u10_u6_U98  ( .A1(_u10_u6_n2040 ), .A2(_u10_u6_n2041 ), .A3(_u10_u6_n2042 ), .ZN(_u10_u6_n2009 ) );
AND2_X1 _u10_u6_U97  ( .A1(_u10_u6_n2038 ), .A2(_u10_u6_n2039 ), .ZN(_u10_u6_n1929 ) );
NOR2_X1 _u10_u6_U96  ( .A1(_u10_u6_n1929 ), .A2(_u10_u6_n2037 ), .ZN(_u10_u6_n2010 ) );
NAND2_X1 _u10_u6_U95  ( .A1(_u10_u6_n2035 ), .A2(_u10_u6_n2036 ), .ZN(_u10_u6_n1902 ) );
NAND3_X1 _u10_u6_U94  ( .A1(_u10_u6_n1902 ), .A2(_u10_u6_n2033 ), .A3(_u10_u6_n2034 ), .ZN(_u10_u6_n1973 ) );
NOR2_X1 _u10_u6_U93  ( .A1(_u10_u6_n1978 ), .A2(_u10_u6_n1973 ), .ZN(_u10_u6_n2032 ) );
NOR2_X1 _u10_u6_U92  ( .A1(1'b0), .A2(_u10_u6_n2032 ), .ZN(_u10_u6_n2028 ));
NOR2_X1 _u10_u6_U91  ( .A1(_u10_u6_n2030 ), .A2(_u10_u6_n2031 ), .ZN(_u10_u6_n2029 ) );
NOR4_X1 _u10_u6_U90  ( .A1(_u10_u6_n2026 ), .A2(_u10_u6_n2027 ), .A3(_u10_u6_n2028 ), .A4(_u10_u6_n2029 ), .ZN(_u10_u6_n2024 ) );
NOR2_X1 _u10_u6_U89  ( .A1(_u10_u6_n2024 ), .A2(_u10_u6_n2025 ), .ZN(_u10_u6_n2011 ) );
NAND3_X1 _u10_u6_U88  ( .A1(_u10_u6_n2021 ), .A2(_u10_u6_n2022 ), .A3(_u10_u6_n2023 ), .ZN(_u10_u6_n2020 ) );
AND2_X1 _u10_u6_U87  ( .A1(_u10_u6_n2019 ), .A2(_u10_u6_n2020 ), .ZN(_u10_u6_n1838 ) );
INV_X1 _u10_u6_U86  ( .A(_u10_u6_n2018 ), .ZN(_u10_u6_n2016 ) );
NOR4_X1 _u10_u6_U85  ( .A1(_u10_u6_n2015 ), .A2(_u10_u6_n1838 ), .A3(_u10_u6_n2016 ), .A4(_u10_u6_n2017 ), .ZN(_u10_u6_n2013 ) );
NOR2_X1 _u10_u6_U84  ( .A1(_u10_u6_n2013 ), .A2(_u10_u6_n2014 ), .ZN(_u10_u6_n2012 ) );
NOR4_X1 _u10_u6_U83  ( .A1(_u10_u6_n2009 ), .A2(_u10_u6_n2010 ), .A3(_u10_u6_n2011 ), .A4(_u10_u6_n2012 ), .ZN(_u10_u6_n1821 ) );
NAND2_X1 _u10_u6_U82  ( .A1(_u10_u6_n1924 ), .A2(_u10_u6_n2008 ), .ZN(_u10_u6_n1993 ) );
NAND2_X1 _u10_u6_U81  ( .A1(_u10_u6_n2006 ), .A2(_u10_u6_n2007 ), .ZN(_u10_u6_n1994 ) );
NAND2_X1 _u10_u6_U80  ( .A1(_u10_u6_n2004 ), .A2(_u10_u6_n2005 ), .ZN(_u10_u6_n1995 ) );
AND2_X1 _u10_u6_U79  ( .A1(_u10_u6_n2002 ), .A2(_u10_u6_n2003 ), .ZN(_u10_u6_n1998 ) );
NOR2_X1 _u10_u6_U78  ( .A1(_u10_u6_n2000 ), .A2(_u10_u6_n2001 ), .ZN(_u10_u6_n1999 ) );
NOR3_X1 _u10_u6_U77  ( .A1(_u10_u6_n1997 ), .A2(_u10_u6_n1998 ), .A3(_u10_u6_n1999 ), .ZN(_u10_u6_n1996 ) );
NAND4_X1 _u10_u6_U76  ( .A1(_u10_u6_n1993 ), .A2(_u10_u6_n1994 ), .A3(_u10_u6_n1995 ), .A4(_u10_u6_n1996 ), .ZN(_u10_u6_n1985 ) );
INV_X1 _u10_u6_U75  ( .A(_u10_u6_n1992 ), .ZN(_u10_u6_n1989 ) );
NAND3_X1 _u10_u6_U74  ( .A1(_u10_u6_n1989 ), .A2(_u10_u6_n1990 ), .A3(_u10_u6_n1991 ), .ZN(_u10_u6_n1986 ) );
NOR4_X1 _u10_u6_U73  ( .A1(_u10_u6_n1985 ), .A2(_u10_u6_n1986 ), .A3(_u10_u6_n1987 ), .A4(_u10_u6_n1988 ), .ZN(_u10_u6_n1822 ) );
INV_X1 _u10_u6_U72  ( .A(_u10_u6_n1984 ), .ZN(_u10_u6_n1980 ) );
NAND4_X1 _u10_u6_U71  ( .A1(_u10_u6_n1980 ), .A2(_u10_u6_n1981 ), .A3(_u10_u6_n1982 ), .A4(_u10_u6_n1983 ), .ZN(_u10_u6_n1941 ) );
NOR3_X1 _u10_u6_U70  ( .A1(_u10_u6_n1977 ), .A2(_u10_u6_n1978 ), .A3(_u10_u6_n1979 ), .ZN(_u10_u6_n1971 ) );
NOR4_X1 _u10_u6_U69  ( .A1(_u10_u6_n1973 ), .A2(_u10_u6_n1974 ), .A3(_u10_u6_n1975 ), .A4(_u10_u6_n1976 ), .ZN(_u10_u6_n1972 ) );
NAND4_X1 _u10_u6_U68  ( .A1(_u10_u6_n1969 ), .A2(_u10_u6_n1970 ), .A3(_u10_u6_n1971 ), .A4(_u10_u6_n1972 ), .ZN(_u10_u6_n1968 ) );
NAND2_X1 _u10_u6_U67  ( .A1(_u10_u6_n1967 ), .A2(_u10_u6_n1968 ), .ZN(_u10_u6_n1942 ) );
NAND3_X1 _u10_u6_U66  ( .A1(_u10_u6_n1964 ), .A2(_u10_u6_n1965 ), .A3(_u10_u6_n1966 ), .ZN(_u10_u6_n1943 ) );
AND4_X1 _u10_u6_U65  ( .A1(_u10_u6_n1961 ), .A2(_u10_u6_n1863 ), .A3(_u10_u6_n1962 ), .A4(_u10_u6_n1963 ), .ZN(_u10_u6_n1957 ) );
NOR2_X1 _u10_u6_U64  ( .A1(_u10_u6_n1959 ), .A2(_u10_u6_n1960 ), .ZN(_u10_u6_n1958 ) );
NOR2_X1 _u10_u6_U63  ( .A1(_u10_u6_n1957 ), .A2(_u10_u6_n1958 ), .ZN(_u10_u6_n1945 ) );
NOR2_X1 _u10_u6_U62  ( .A1(_u10_u6_n1955 ), .A2(_u10_u6_n1956 ), .ZN(_u10_u6_n1953 ) );
NOR4_X1 _u10_u6_U61  ( .A1(_u10_u6_n1952 ), .A2(_u10_u6_n1953 ), .A3(_u10_u6_n1846 ), .A4(_u10_u6_n1954 ), .ZN(_u10_u6_n1946 ) );
NOR2_X1 _u10_u6_U60  ( .A1(_u10_u6_n1950 ), .A2(_u10_u6_n1951 ), .ZN(_u10_u6_n1949 ) );
NOR2_X1 _u10_u6_U59  ( .A1(_u10_u6_n1948 ), .A2(_u10_u6_n1949 ), .ZN(_u10_u6_n1947 ) );
NOR3_X1 _u10_u6_U58  ( .A1(_u10_u6_n1945 ), .A2(_u10_u6_n1946 ), .A3(_u10_u6_n1947 ), .ZN(_u10_u6_n1944 ) );
NAND4_X1 _u10_u6_U57  ( .A1(_u10_u6_n1941 ), .A2(_u10_u6_n1942 ), .A3(_u10_u6_n1943 ), .A4(_u10_u6_n1944 ), .ZN(_u10_u6_n1824 ) );
NAND2_X1 _u10_u6_U56  ( .A1(_u10_u6_n1939 ), .A2(_u10_u6_n1940 ), .ZN(_u10_u6_n1938 ) );
NAND2_X1 _u10_u6_U55  ( .A1(_u10_u6_n1937 ), .A2(_u10_u6_n1938 ), .ZN(_u10_u6_n1903 ) );
NAND2_X1 _u10_u6_U54  ( .A1(_u10_u6_n1935 ), .A2(_u10_u6_n1936 ), .ZN(_u10_u6_n1934 ) );
NAND2_X1 _u10_u6_U53  ( .A1(_u10_u6_n1933 ), .A2(_u10_u6_n1934 ), .ZN(_u10_u6_n1931 ) );
NAND2_X1 _u10_u6_U52  ( .A1(_u10_u6_n1931 ), .A2(_u10_u6_n1932 ), .ZN(_u10_u6_n1904 ) );
NAND2_X1 _u10_u6_U51  ( .A1(_u10_u6_n1929 ), .A2(_u10_u6_n1930 ), .ZN(_u10_u6_n1927 ) );
NAND2_X1 _u10_u6_U50  ( .A1(_u10_u6_n1927 ), .A2(_u10_u6_n1928 ), .ZN(_u10_u6_n1905 ) );
NOR3_X1 _u10_u6_U49  ( .A1(_u10_u6_n1916 ), .A2(_u10_u6_n1925 ), .A3(_u10_u6_n1926 ), .ZN(_u10_u6_n1919 ) );
NOR2_X1 _u10_u6_U48  ( .A1(_u10_u6_n1923 ), .A2(_u10_u6_n1924 ), .ZN(_u10_u6_n1921 ) );
NOR2_X1 _u10_u6_U47  ( .A1(_u10_u6_n1921 ), .A2(_u10_u6_n1922 ), .ZN(_u10_u6_n1920 ) );
NOR2_X1 _u10_u6_U46  ( .A1(_u10_u6_n1919 ), .A2(_u10_u6_n1920 ), .ZN(_u10_u6_n1917 ) );
NOR2_X1 _u10_u6_U45  ( .A1(_u10_u6_n1917 ), .A2(_u10_u6_n1918 ), .ZN(_u10_u6_n1907 ) );
NOR2_X1 _u10_u6_U44  ( .A1(_u10_u6_n1915 ), .A2(_u10_u6_n1916 ), .ZN(_u10_u6_n1914 ) );
NOR2_X1 _u10_u6_U43  ( .A1(_u10_u6_n1914 ), .A2(1'b0), .ZN(_u10_u6_n1912 ));
NOR2_X1 _u10_u6_U42  ( .A1(_u10_u6_n1912 ), .A2(_u10_u6_n1913 ), .ZN(_u10_u6_n1908 ) );
NOR2_X1 _u10_u6_U41  ( .A1(_u10_u6_n1891 ), .A2(_u10_u6_n1911 ), .ZN(_u10_u6_n1910 ) );
NOR2_X1 _u10_u6_U40  ( .A1(_u10_u6_n1910 ), .A2(_u10_u6_n1868 ), .ZN(_u10_u6_n1909 ) );
NOR3_X1 _u10_u6_U39  ( .A1(_u10_u6_n1907 ), .A2(_u10_u6_n1908 ), .A3(_u10_u6_n1909 ), .ZN(_u10_u6_n1906 ) );
NAND4_X1 _u10_u6_U38  ( .A1(_u10_u6_n1903 ), .A2(_u10_u6_n1904 ), .A3(_u10_u6_n1905 ), .A4(_u10_u6_n1906 ), .ZN(_u10_u6_n1825 ) );
NAND2_X1 _u10_u6_U37  ( .A1(_u10_u6_n1901 ), .A2(_u10_u6_n1902 ), .ZN(_u10_u6_n1900 ) );
NAND2_X1 _u10_u6_U36  ( .A1(_u10_u6_n1899 ), .A2(_u10_u6_n1900 ), .ZN(_u10_u6_n1875 ) );
OR2_X1 _u10_u6_U35  ( .A1(_u10_u6_n1847 ), .A2(_u10_u6_n1898 ), .ZN(_u10_u6_n1897 ) );
NAND2_X1 _u10_u6_U34  ( .A1(_u10_u6_n1896 ), .A2(_u10_u6_n1897 ), .ZN(_u10_u6_n1895 ) );
NAND2_X1 _u10_u6_U33  ( .A1(_u10_u6_n1894 ), .A2(_u10_u6_n1895 ), .ZN(_u10_u6_n1876 ) );
NAND2_X1 _u10_u6_U32  ( .A1(_u10_u6_n1892 ), .A2(_u10_u6_n1893 ), .ZN(_u10_u6_n1877 ) );
NOR3_X1 _u10_u6_U31  ( .A1(_u10_u6_n1884 ), .A2(_u10_u6_n1890 ), .A3(_u10_u6_n1891 ), .ZN(_u10_u6_n1889 ) );
NOR2_X1 _u10_u6_U30  ( .A1(_u10_u6_n1840 ), .A2(_u10_u6_n1889 ), .ZN(_u10_u6_n1879 ) );
NOR2_X1 _u10_u6_U29  ( .A1(_u10_u6_n1887 ), .A2(_u10_u6_n1888 ), .ZN(_u10_u6_n1880 ) );
NOR3_X1 _u10_u6_U28  ( .A1(_u10_u6_n1884 ), .A2(_u10_u6_n1885 ), .A3(_u10_u6_n1886 ), .ZN(_u10_u6_n1883 ) );
NOR2_X1 _u10_u6_U27  ( .A1(_u10_u6_n1882 ), .A2(_u10_u6_n1883 ), .ZN(_u10_u6_n1881 ) );
NOR3_X1 _u10_u6_U26  ( .A1(_u10_u6_n1879 ), .A2(_u10_u6_n1880 ), .A3(_u10_u6_n1881 ), .ZN(_u10_u6_n1878 ) );
NAND4_X1 _u10_u6_U25  ( .A1(_u10_u6_n1875 ), .A2(_u10_u6_n1876 ), .A3(_u10_u6_n1877 ), .A4(_u10_u6_n1878 ), .ZN(_u10_u6_n1826 ) );
NOR3_X1 _u10_u6_U24  ( .A1(_u10_u6_n1872 ), .A2(_u10_u6_n1873 ), .A3(_u10_u6_n1874 ), .ZN(_u10_u6_n1871 ) );
NAND4_X1 _u10_u6_U23  ( .A1(_u10_u6_n1868 ), .A2(_u10_u6_n1869 ), .A3(_u10_u6_n1870 ), .A4(_u10_u6_n1871 ), .ZN(_u10_u6_n1867 ) );
NAND2_X1 _u10_u6_U22  ( .A1(_u10_u6_n1866 ), .A2(_u10_u6_n1867 ), .ZN(_u10_u6_n1865 ) );
NAND3_X1 _u10_u6_U21  ( .A1(_u10_u6_n1863 ), .A2(_u10_u6_n1864 ), .A3(_u10_u6_n1865 ), .ZN(_u10_u6_n1862 ) );
NAND2_X1 _u10_u6_U20  ( .A1(_u10_u6_n1861 ), .A2(_u10_u6_n1862 ), .ZN(_u10_u6_n1828 ) );
NAND3_X1 _u10_u6_U19  ( .A1(_u10_u6_n1858 ), .A2(_u10_u6_n1859 ), .A3(_u10_u6_n1860 ), .ZN(_u10_u6_n1857 ) );
NAND2_X1 _u10_u6_U18  ( .A1(_u10_u6_n1856 ), .A2(_u10_u6_n1857 ), .ZN(_u10_u6_n1829 ) );
OR2_X1 _u10_u6_U17  ( .A1(_u10_u6_n1854 ), .A2(_u10_u6_n1855 ), .ZN(_u10_u6_n1830 ) );
NOR2_X1 _u10_u6_U16  ( .A1(_u10_u6_n1852 ), .A2(_u10_u6_n1853 ), .ZN(_u10_u6_n1850 ) );
NOR3_X1 _u10_u6_U15  ( .A1(_u10_u6_n1850 ), .A2(_u10_u6_n1851 ), .A3(_u10_u6_n1838 ), .ZN(_u10_u6_n1848 ) );
NOR2_X1 _u10_u6_U14  ( .A1(_u10_u6_n1848 ), .A2(_u10_u6_n1849 ), .ZN(_u10_u6_n1832 ) );
NOR2_X1 _u10_u6_U13  ( .A1(_u10_u6_n1846 ), .A2(_u10_u6_n1847 ), .ZN(_u10_u6_n1845 ) );
NOR3_X1 _u10_u6_U12  ( .A1(_u10_u6_n1844 ), .A2(1'b0), .A3(_u10_u6_n1845 ),.ZN(_u10_u6_n1842 ) );
NOR2_X1 _u10_u6_U11  ( .A1(_u10_u6_n1842 ), .A2(_u10_u6_n1843 ), .ZN(_u10_u6_n1833 ) );
NOR2_X1 _u10_u6_U10  ( .A1(_u10_u6_n1840 ), .A2(_u10_u6_n1841 ), .ZN(_u10_u6_n1839 ) );
NOR3_X1 _u10_u6_U9  ( .A1(_u10_u6_n1837 ), .A2(_u10_u6_n1838 ), .A3(_u10_u6_n1839 ), .ZN(_u10_u6_n1835 ) );
NOR2_X1 _u10_u6_U8  ( .A1(_u10_u6_n1835 ), .A2(_u10_u6_n1836 ), .ZN(_u10_u6_n1834 ) );
NOR3_X1 _u10_u6_U7  ( .A1(_u10_u6_n1832 ), .A2(_u10_u6_n1833 ), .A3(_u10_u6_n1834 ), .ZN(_u10_u6_n1831 ) );
NAND4_X1 _u10_u6_U6  ( .A1(_u10_u6_n1828 ), .A2(_u10_u6_n1829 ), .A3(_u10_u6_n1830 ), .A4(_u10_u6_n1831 ), .ZN(_u10_u6_n1827 ) );
NOR4_X1 _u10_u6_U5  ( .A1(_u10_u6_n1824 ), .A2(_u10_u6_n1825 ), .A3(_u10_u6_n1826 ), .A4(_u10_u6_n1827 ), .ZN(_u10_u6_n1823 ) );
NAND4_X1 _u10_u6_U4  ( .A1(_u10_u6_n1820 ), .A2(_u10_u6_n1821 ), .A3(_u10_u6_n1822 ), .A4(_u10_u6_n1823 ), .ZN(_u10_u6_n1818 ) );
MUX2_X1 _u10_u6_U3  ( .A(_u10_u6_n1818 ), .B(_u10_SYNOPSYS_UNCONNECTED_27 ),.S(_u10_u6_n1819 ), .Z(_u10_u6_n1812 ) );
DFFR_X1 _u10_u6_state_reg_1_  ( .D(_u10_u6_n1812 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_27 ), .QN(_u10_u6_n1814 ));
DFFR_X1 _u10_u6_state_reg_2_  ( .D(_u10_u6_n1811 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_26 ), .QN(_u10_u6_n1815 ));
DFFR_X1 _u10_u6_state_reg_3_  ( .D(_u10_u6_n1810 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_25 ), .QN(_u10_u6_n1816 ));
DFFR_X1 _u10_u6_state_reg_4_  ( .D(_u10_u6_n1809 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_24 ), .QN(_u10_u6_n1817 ));
DFFR_X1 _u10_u6_state_reg_0_  ( .D(_u10_u6_n1808 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_28 ), .QN(_u10_u6_n1813 ));
NOR2_X1 _u10_u7_U1606  ( .A1(_u10_SYNOPSYS_UNCONNECTED_31 ), .A2(_u10_u7_n1814 ), .ZN(_u10_u7_n3174 ) );
NOR3_X1 _u10_u7_U1605  ( .A1(_u10_SYNOPSYS_UNCONNECTED_30 ), .A2(_u10_u7_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_33 ), .ZN(_u10_u7_n3328 ) );
NAND2_X1 _u10_u7_U1604  ( .A1(_u10_u7_n3174 ), .A2(_u10_u7_n3328 ), .ZN(_u10_u7_n1843 ) );
INV_X1 _u10_u7_U1603  ( .A(_u10_u7_n1843 ), .ZN(_u10_u7_n2461 ) );
INV_X1 _u10_u7_U1602  ( .A(1'b0), .ZN(_u10_u7_n2466 ) );
INV_X1 _u10_u7_U1601  ( .A(1'b0), .ZN(_u10_u7_n2305 ) );
NAND2_X1 _u10_u7_U1600  ( .A1(_u10_u7_n2466 ), .A2(_u10_u7_n2305 ), .ZN(_u10_u7_n1954 ) );
INV_X1 _u10_u7_U1599  ( .A(_u10_u7_n1954 ), .ZN(_u10_u7_n2467 ) );
INV_X1 _u10_u7_U1598  ( .A(1'b0), .ZN(_u10_u7_n1936 ) );
NOR2_X1 _u10_u7_U1597  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u7_n2223 ) );
INV_X1 _u10_u7_U1596  ( .A(1'b0), .ZN(_u10_u7_n1922 ) );
NAND2_X1 _u10_u7_U1595  ( .A1(_u10_u7_n2223 ), .A2(_u10_u7_n1922 ), .ZN(_u10_u7_n2200 ) );
NOR2_X1 _u10_u7_U1594  ( .A1(_u10_u7_n2200 ), .A2(1'b0), .ZN(_u10_u7_n2502 ));
INV_X1 _u10_u7_U1593  ( .A(1'b0), .ZN(_u10_u7_n2978 ) );
INV_X1 _u10_u7_U1592  ( .A(1'b0), .ZN(_u10_u7_n3000 ) );
NAND2_X1 _u10_u7_U1591  ( .A1(_u10_u7_n2978 ), .A2(_u10_u7_n3000 ), .ZN(_u10_u7_n3356 ) );
INV_X1 _u10_u7_U1590  ( .A(1'b0), .ZN(_u10_u7_n2405 ) );
INV_X1 _u10_u7_U1589  ( .A(1'b0), .ZN(_u10_u7_n2972 ) );
NAND2_X1 _u10_u7_U1588  ( .A1(_u10_u7_n2405 ), .A2(_u10_u7_n2972 ), .ZN(_u10_u7_n2008 ) );
NOR2_X1 _u10_u7_U1587  ( .A1(_u10_u7_n3356 ), .A2(_u10_u7_n2008 ), .ZN(_u10_u7_n2195 ) );
NAND2_X1 _u10_u7_U1586  ( .A1(_u10_u7_n2502 ), .A2(_u10_u7_n2195 ), .ZN(_u10_u7_n2490 ) );
INV_X1 _u10_u7_U1585  ( .A(1'b0), .ZN(_u10_u7_n3040 ) );
INV_X1 _u10_u7_U1584  ( .A(1'b0), .ZN(_u10_u7_n3006 ) );
NAND2_X1 _u10_u7_U1583  ( .A1(_u10_u7_n3040 ), .A2(_u10_u7_n3006 ), .ZN(_u10_u7_n2508 ) );
NOR2_X1 _u10_u7_U1582  ( .A1(_u10_u7_n2508 ), .A2(1'b0), .ZN(_u10_u7_n2493 ));
INV_X1 _u10_u7_U1581  ( .A(1'b0), .ZN(_u10_u7_n2038 ) );
NAND2_X1 _u10_u7_U1580  ( .A1(_u10_u7_n2493 ), .A2(_u10_u7_n2038 ), .ZN(_u10_u7_n2174 ) );
NOR2_X1 _u10_u7_U1579  ( .A1(_u10_u7_n2490 ), .A2(_u10_u7_n2174 ), .ZN(_u10_u7_n2659 ) );
INV_X1 _u10_u7_U1578  ( .A(1'b0), .ZN(_u10_u7_n2175 ) );
NAND3_X1 _u10_u7_U1577  ( .A1(_u10_u7_n2659 ), .A2(_u10_u7_n2175 ), .A3(1'b0), .ZN(_u10_u7_n3189 ) );
NOR2_X1 _u10_u7_U1576  ( .A1(_u10_u7_n3189 ), .A2(1'b0), .ZN(_u10_u7_n2528 ));
INV_X1 _u10_u7_U1575  ( .A(1'b0), .ZN(_u10_u7_n2837 ) );
NAND2_X1 _u10_u7_U1574  ( .A1(_u10_u7_n2528 ), .A2(_u10_u7_n2837 ), .ZN(_u10_u7_n2567 ) );
INV_X1 _u10_u7_U1573  ( .A(1'b0), .ZN(_u10_u7_n2080 ) );
INV_X1 _u10_u7_U1572  ( .A(1'b0), .ZN(_u10_u7_n2166 ) );
NAND2_X1 _u10_u7_U1571  ( .A1(_u10_u7_n2080 ), .A2(_u10_u7_n2166 ), .ZN(_u10_u7_n2840 ) );
NOR2_X1 _u10_u7_U1570  ( .A1(_u10_u7_n2567 ), .A2(_u10_u7_n2840 ), .ZN(_u10_u7_n2443 ) );
INV_X1 _u10_u7_U1569  ( .A(1'b0), .ZN(_u10_u7_n2600 ) );
INV_X1 _u10_u7_U1568  ( .A(1'b0), .ZN(_u10_u7_n2836 ) );
NAND2_X1 _u10_u7_U1567  ( .A1(_u10_u7_n2600 ), .A2(_u10_u7_n2836 ), .ZN(_u10_u7_n2428 ) );
INV_X1 _u10_u7_U1566  ( .A(_u10_u7_n2428 ), .ZN(_u10_u7_n2078 ) );
NAND2_X1 _u10_u7_U1565  ( .A1(_u10_u7_n2443 ), .A2(_u10_u7_n2078 ), .ZN(_u10_u7_n2282 ) );
INV_X1 _u10_u7_U1564  ( .A(1'b0), .ZN(_u10_u7_n2874 ) );
INV_X1 _u10_u7_U1563  ( .A(1'b0), .ZN(_u10_u7_n2031 ) );
NAND2_X1 _u10_u7_U1562  ( .A1(_u10_u7_n2874 ), .A2(_u10_u7_n2031 ), .ZN(_u10_u7_n1976 ) );
NOR2_X1 _u10_u7_U1561  ( .A1(_u10_u7_n2282 ), .A2(_u10_u7_n1976 ), .ZN(_u10_u7_n2411 ) );
NAND3_X1 _u10_u7_U1560  ( .A1(_u10_u7_n2467 ), .A2(_u10_u7_n1936 ), .A3(_u10_u7_n2411 ), .ZN(_u10_u7_n2464 ) );
NAND3_X1 _u10_u7_U1559  ( .A1(_u10_u7_n2166 ), .A2(_u10_u7_n2837 ), .A3(1'b0), .ZN(_u10_u7_n3276 ) );
INV_X1 _u10_u7_U1558  ( .A(_u10_u7_n3276 ), .ZN(_u10_u7_n2442 ) );
NAND3_X1 _u10_u7_U1557  ( .A1(_u10_u7_n2836 ), .A2(_u10_u7_n2080 ), .A3(_u10_u7_n2442 ), .ZN(_u10_u7_n2838 ) );
INV_X1 _u10_u7_U1556  ( .A(_u10_u7_n2838 ), .ZN(_u10_u7_n2850 ) );
NOR2_X1 _u10_u7_U1555  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u7_n2953 ) );
NAND2_X1 _u10_u7_U1554  ( .A1(_u10_u7_n2850 ), .A2(_u10_u7_n2953 ), .ZN(_u10_u7_n2947 ) );
INV_X1 _u10_u7_U1553  ( .A(_u10_u7_n2947 ), .ZN(_u10_u7_n2420 ) );
NAND2_X1 _u10_u7_U1552  ( .A1(_u10_u7_n1936 ), .A2(_u10_u7_n2874 ), .ZN(_u10_u7_n2030 ) );
INV_X1 _u10_u7_U1551  ( .A(_u10_u7_n2030 ), .ZN(_u10_u7_n2162 ) );
NAND2_X1 _u10_u7_U1550  ( .A1(_u10_u7_n2420 ), .A2(_u10_u7_n2162 ), .ZN(_u10_u7_n2828 ) );
INV_X1 _u10_u7_U1549  ( .A(_u10_u7_n2828 ), .ZN(_u10_u7_n2551 ) );
NAND2_X1 _u10_u7_U1548  ( .A1(_u10_u7_n2551 ), .A2(_u10_u7_n2467 ), .ZN(_u10_u7_n3416 ) );
NAND2_X1 _u10_u7_U1547  ( .A1(_u10_u7_n2464 ), .A2(_u10_u7_n3416 ), .ZN(_u10_u7_n2266 ) );
INV_X1 _u10_u7_U1546  ( .A(_u10_u7_n2266 ), .ZN(_u10_u7_n3410 ) );
NAND2_X1 _u10_u7_U1545  ( .A1(1'b0), .A2(_u10_u7_n2305 ), .ZN(_u10_u7_n3411 ) );
INV_X1 _u10_u7_U1544  ( .A(_u10_u7_n3356 ), .ZN(_u10_u7_n1983 ) );
NAND3_X1 _u10_u7_U1543  ( .A1(_u10_u7_n1983 ), .A2(_u10_u7_n2405 ), .A3(1'b0), .ZN(_u10_u7_n2022 ) );
INV_X1 _u10_u7_U1542  ( .A(_u10_u7_n2022 ), .ZN(_u10_u7_n2056 ) );
INV_X1 _u10_u7_U1541  ( .A(_u10_u7_n2840 ), .ZN(_u10_u7_n2059 ) );
INV_X1 _u10_u7_U1540  ( .A(1'b0), .ZN(_u10_u7_n1965 ) );
NAND2_X1 _u10_u7_U1539  ( .A1(_u10_u7_n2837 ), .A2(_u10_u7_n1965 ), .ZN(_u10_u7_n1852 ) );
INV_X1 _u10_u7_U1538  ( .A(_u10_u7_n1852 ), .ZN(_u10_u7_n3190 ) );
INV_X1 _u10_u7_U1537  ( .A(1'b0), .ZN(_u10_u7_n1853 ) );
NAND2_X1 _u10_u7_U1536  ( .A1(_u10_u7_n3190 ), .A2(_u10_u7_n1853 ), .ZN(_u10_u7_n2687 ) );
INV_X1 _u10_u7_U1535  ( .A(_u10_u7_n2687 ), .ZN(_u10_u7_n2019 ) );
NAND2_X1 _u10_u7_U1534  ( .A1(_u10_u7_n2059 ), .A2(_u10_u7_n2019 ), .ZN(_u10_u7_n2330 ) );
NOR2_X1 _u10_u7_U1533  ( .A1(_u10_u7_n2428 ), .A2(_u10_u7_n2330 ), .ZN(_u10_u7_n2036 ) );
NAND2_X1 _u10_u7_U1532  ( .A1(_u10_u7_n2056 ), .A2(_u10_u7_n2036 ), .ZN(_u10_u7_n3379 ) );
NOR2_X1 _u10_u7_U1531  ( .A1(_u10_u7_n3379 ), .A2(_u10_u7_n2030 ), .ZN(_u10_u7_n2026 ) );
INV_X1 _u10_u7_U1530  ( .A(1'b0), .ZN(_u10_u7_n2431 ) );
NOR2_X1 _u10_u7_U1529  ( .A1(_u10_u7_n2431 ), .A2(1'b0), .ZN(_u10_u7_n3062 ));
NAND2_X1 _u10_u7_U1528  ( .A1(_u10_u7_n3062 ), .A2(_u10_u7_n2195 ), .ZN(_u10_u7_n3407 ) );
NOR3_X1 _u10_u7_U1527  ( .A1(_u10_u7_n2687 ), .A2(1'b0), .A3(_u10_u7_n3407 ),.ZN(_u10_u7_n3275 ) );
NAND3_X1 _u10_u7_U1526  ( .A1(_u10_u7_n2836 ), .A2(_u10_u7_n2080 ), .A3(_u10_u7_n3275 ), .ZN(_u10_u7_n3297 ) );
INV_X1 _u10_u7_U1525  ( .A(_u10_u7_n3297 ), .ZN(_u10_u7_n3172 ) );
NAND2_X1 _u10_u7_U1524  ( .A1(_u10_u7_n3172 ), .A2(_u10_u7_n2600 ), .ZN(_u10_u7_n2226 ) );
NOR2_X1 _u10_u7_U1523  ( .A1(_u10_u7_n2226 ), .A2(1'b0), .ZN(_u10_u7_n2307 ));
INV_X1 _u10_u7_U1522  ( .A(_u10_u7_n2490 ), .ZN(_u10_u7_n2536 ) );
NAND3_X1 _u10_u7_U1521  ( .A1(_u10_u7_n2536 ), .A2(_u10_u7_n3040 ), .A3(1'b0), .ZN(_u10_u7_n3226 ) );
NOR2_X1 _u10_u7_U1520  ( .A1(_u10_u7_n3226 ), .A2(_u10_u7_n2330 ), .ZN(_u10_u7_n2441 ) );
NAND2_X1 _u10_u7_U1519  ( .A1(_u10_u7_n2441 ), .A2(_u10_u7_n2953 ), .ZN(_u10_u7_n2579 ) );
NOR2_X1 _u10_u7_U1518  ( .A1(_u10_u7_n2579 ), .A2(_u10_u7_n2030 ), .ZN(_u10_u7_n2550 ) );
NOR3_X1 _u10_u7_U1517  ( .A1(_u10_u7_n2026 ), .A2(_u10_u7_n2307 ), .A3(_u10_u7_n2550 ), .ZN(_u10_u7_n3394 ) );
NAND2_X1 _u10_u7_U1516  ( .A1(1'b0), .A2(_u10_u7_n2978 ), .ZN(_u10_u7_n3115 ) );
NOR2_X1 _u10_u7_U1515  ( .A1(_u10_u7_n3115 ), .A2(_u10_u7_n2330 ), .ZN(_u10_u7_n3126 ) );
NAND2_X1 _u10_u7_U1514  ( .A1(_u10_u7_n2162 ), .A2(_u10_u7_n2031 ), .ZN(_u10_u7_n2686 ) );
NOR2_X1 _u10_u7_U1513  ( .A1(_u10_u7_n2686 ), .A2(_u10_u7_n2428 ), .ZN(_u10_u7_n2108 ) );
NAND2_X1 _u10_u7_U1512  ( .A1(_u10_u7_n3126 ), .A2(_u10_u7_n2108 ), .ZN(_u10_u7_n3415 ) );
NAND2_X1 _u10_u7_U1511  ( .A1(_u10_u7_n3394 ), .A2(_u10_u7_n3415 ), .ZN(_u10_u7_n3089 ) );
NAND2_X1 _u10_u7_U1510  ( .A1(_u10_u7_n3089 ), .A2(_u10_u7_n2305 ), .ZN(_u10_u7_n3414 ) );
NAND2_X1 _u10_u7_U1509  ( .A1(_u10_u7_n2466 ), .A2(_u10_u7_n3414 ), .ZN(_u10_u7_n3118 ) );
NAND2_X1 _u10_u7_U1508  ( .A1(_u10_u7_n2078 ), .A2(_u10_u7_n2080 ), .ZN(_u10_u7_n2596 ) );
NAND2_X1 _u10_u7_U1507  ( .A1(1'b0), .A2(_u10_u7_n2493 ), .ZN(_u10_u7_n1961 ) );
NOR3_X1 _u10_u7_U1506  ( .A1(_u10_u7_n2490 ), .A2(1'b0), .A3(_u10_u7_n1961 ),.ZN(_u10_u7_n2054 ) );
NAND2_X1 _u10_u7_U1505  ( .A1(_u10_u7_n2054 ), .A2(_u10_u7_n3190 ), .ZN(_u10_u7_n2061 ) );
OR2_X1 _u10_u7_U1504  ( .A1(_u10_u7_n2596 ), .A2(_u10_u7_n2061 ), .ZN(_u10_u7_n1969 ) );
NOR3_X1 _u10_u7_U1503  ( .A1(_u10_u7_n1976 ), .A2(1'b0), .A3(_u10_u7_n1969 ),.ZN(_u10_u7_n2710 ) );
NAND2_X1 _u10_u7_U1502  ( .A1(_u10_u7_n2710 ), .A2(_u10_u7_n2467 ), .ZN(_u10_u7_n2545 ) );
INV_X1 _u10_u7_U1501  ( .A(_u10_u7_n2545 ), .ZN(_u10_u7_n2087 ) );
NOR2_X1 _u10_u7_U1500  ( .A1(_u10_u7_n3118 ), .A2(_u10_u7_n2087 ), .ZN(_u10_u7_n3145 ) );
NOR2_X1 _u10_u7_U1499  ( .A1(_u10_u7_n2030 ), .A2(1'b0), .ZN(_u10_u7_n2668 ));
NAND2_X1 _u10_u7_U1498  ( .A1(1'b0), .A2(_u10_u7_n2668 ), .ZN(_u10_u7_n2163 ) );
INV_X1 _u10_u7_U1497  ( .A(_u10_u7_n2163 ), .ZN(_u10_u7_n2875 ) );
INV_X1 _u10_u7_U1496  ( .A(_u10_u7_n1976 ), .ZN(_u10_u7_n2747 ) );
NAND3_X1 _u10_u7_U1495  ( .A1(_u10_u7_n2747 ), .A2(_u10_u7_n2600 ), .A3(1'b0), .ZN(_u10_u7_n3393 ) );
NOR3_X1 _u10_u7_U1494  ( .A1(1'b0), .A2(1'b0), .A3(_u10_u7_n3393 ), .ZN(_u10_u7_n3180 ) );
INV_X1 _u10_u7_U1493  ( .A(1'b0), .ZN(_u10_u7_n2113 ) );
INV_X1 _u10_u7_U1492  ( .A(1'b0), .ZN(_u10_u7_n3066 ) );
NAND2_X1 _u10_u7_U1491  ( .A1(_u10_u7_n2175 ), .A2(_u10_u7_n3066 ), .ZN(_u10_u7_n2216 ) );
INV_X1 _u10_u7_U1490  ( .A(_u10_u7_n2659 ), .ZN(_u10_u7_n2643 ) );
NOR2_X1 _u10_u7_U1489  ( .A1(_u10_u7_n2216 ), .A2(_u10_u7_n2643 ), .ZN(_u10_u7_n2049 ) );
AND2_X1 _u10_u7_U1488  ( .A1(_u10_u7_n2049 ), .A2(_u10_u7_n1853 ), .ZN(_u10_u7_n3223 ) );
NAND2_X1 _u10_u7_U1487  ( .A1(_u10_u7_n3223 ), .A2(_u10_u7_n1965 ), .ZN(_u10_u7_n2531 ) );
NOR2_X1 _u10_u7_U1486  ( .A1(_u10_u7_n2531 ), .A2(1'b0), .ZN(_u10_u7_n2884 ));
NAND2_X1 _u10_u7_U1485  ( .A1(_u10_u7_n2884 ), .A2(_u10_u7_n2166 ), .ZN(_u10_u7_n1841 ) );
NOR2_X1 _u10_u7_U1484  ( .A1(_u10_u7_n1841 ), .A2(1'b0), .ZN(_u10_u7_n3129 ));
NAND2_X1 _u10_u7_U1483  ( .A1(_u10_u7_n3129 ), .A2(_u10_u7_n2836 ), .ZN(_u10_u7_n2842 ) );
INV_X1 _u10_u7_U1482  ( .A(_u10_u7_n2842 ), .ZN(_u10_u7_n2833 ) );
NAND2_X1 _u10_u7_U1481  ( .A1(_u10_u7_n2833 ), .A2(_u10_u7_n2600 ), .ZN(_u10_u7_n2853 ) );
INV_X1 _u10_u7_U1480  ( .A(_u10_u7_n2853 ), .ZN(_u10_u7_n2082 ) );
NAND2_X1 _u10_u7_U1479  ( .A1(_u10_u7_n2082 ), .A2(_u10_u7_n2031 ), .ZN(_u10_u7_n2274 ) );
INV_X1 _u10_u7_U1478  ( .A(_u10_u7_n2274 ), .ZN(_u10_u7_n2669 ) );
NAND3_X1 _u10_u7_U1477  ( .A1(_u10_u7_n2668 ), .A2(_u10_u7_n2113 ), .A3(_u10_u7_n2669 ), .ZN(_u10_u7_n1858 ) );
INV_X1 _u10_u7_U1476  ( .A(_u10_u7_n1858 ), .ZN(_u10_u7_n3067 ) );
NAND2_X1 _u10_u7_U1475  ( .A1(_u10_u7_n3067 ), .A2(1'b0), .ZN(_u10_u7_n2092 ) );
INV_X1 _u10_u7_U1474  ( .A(_u10_u7_n2092 ), .ZN(_u10_u7_n3294 ) );
INV_X1 _u10_u7_U1473  ( .A(1'b0), .ZN(_u10_u7_n2446 ) );
INV_X1 _u10_u7_U1472  ( .A(1'b0), .ZN(_u10_u7_n2996 ) );
NAND2_X1 _u10_u7_U1471  ( .A1(_u10_u7_n3067 ), .A2(_u10_u7_n2996 ), .ZN(_u10_u7_n1847 ) );
NOR3_X1 _u10_u7_U1470  ( .A1(_u10_u7_n2446 ), .A2(1'b0), .A3(_u10_u7_n1847 ),.ZN(_u10_u7_n3413 ) );
NOR4_X1 _u10_u7_U1469  ( .A1(_u10_u7_n2875 ), .A2(_u10_u7_n3180 ), .A3(_u10_u7_n3294 ), .A4(_u10_u7_n3413 ), .ZN(_u10_u7_n3412 ) );
NAND4_X1 _u10_u7_U1468  ( .A1(_u10_u7_n3410 ), .A2(_u10_u7_n3411 ), .A3(_u10_u7_n3145 ), .A4(_u10_u7_n3412 ), .ZN(_u10_u7_n3409 ) );
NAND2_X1 _u10_u7_U1467  ( .A1(_u10_u7_n2461 ), .A2(_u10_u7_n3409 ), .ZN(_u10_u7_n3380 ) );
NOR2_X1 _u10_u7_U1466  ( .A1(_u10_u7_n1817 ), .A2(_u10_u7_n1816 ), .ZN(_u10_u7_n3368 ) );
AND2_X1 _u10_u7_U1465  ( .A1(_u10_u7_n3368 ), .A2(_u10_u7_n1813 ), .ZN(_u10_u7_n3320 ) );
NOR2_X1 _u10_u7_U1464  ( .A1(_u10_SYNOPSYS_UNCONNECTED_32 ), .A2(_u10_u7_n1815 ), .ZN(_u10_u7_n3236 ) );
NAND2_X1 _u10_u7_U1463  ( .A1(_u10_u7_n3320 ), .A2(_u10_u7_n3236 ), .ZN(_u10_u7_n2607 ) );
INV_X1 _u10_u7_U1462  ( .A(_u10_u7_n2607 ), .ZN(_u10_u7_n1966 ) );
INV_X1 _u10_u7_U1461  ( .A(_u10_u7_n2200 ), .ZN(_u10_u7_n3216 ) );
NAND2_X1 _u10_u7_U1460  ( .A1(1'b0), .A2(_u10_u7_n3216 ), .ZN(_u10_u7_n2367 ) );
INV_X1 _u10_u7_U1459  ( .A(_u10_u7_n2367 ), .ZN(_u10_u7_n3183 ) );
NAND2_X1 _u10_u7_U1458  ( .A1(_u10_u7_n3183 ), .A2(_u10_u7_n2195 ), .ZN(_u10_u7_n2194 ) );
INV_X1 _u10_u7_U1457  ( .A(_u10_u7_n2194 ), .ZN(_u10_u7_n2055 ) );
NAND2_X1 _u10_u7_U1456  ( .A1(_u10_u7_n2055 ), .A2(_u10_u7_n1853 ), .ZN(_u10_u7_n3401 ) );
INV_X1 _u10_u7_U1455  ( .A(_u10_u7_n2531 ), .ZN(_u10_u7_n2190 ) );
INV_X1 _u10_u7_U1454  ( .A(1'b0), .ZN(_u10_u7_n3001 ) );
NAND2_X1 _u10_u7_U1453  ( .A1(_u10_u7_n3001 ), .A2(_u10_u7_n2466 ), .ZN(_u10_u7_n2156 ) );
NOR2_X1 _u10_u7_U1452  ( .A1(_u10_u7_n2166 ), .A2(_u10_u7_n2596 ), .ZN(_u10_u7_n2594 ) );
NAND2_X1 _u10_u7_U1451  ( .A1(_u10_u7_n2594 ), .A2(_u10_u7_n2031 ), .ZN(_u10_u7_n2752 ) );
INV_X1 _u10_u7_U1450  ( .A(_u10_u7_n2752 ), .ZN(_u10_u7_n2421 ) );
NAND2_X1 _u10_u7_U1449  ( .A1(_u10_u7_n2421 ), .A2(_u10_u7_n2874 ), .ZN(_u10_u7_n2033 ) );
INV_X1 _u10_u7_U1448  ( .A(_u10_u7_n2033 ), .ZN(_u10_u7_n2742 ) );
NAND3_X1 _u10_u7_U1447  ( .A1(_u10_u7_n2305 ), .A2(_u10_u7_n1936 ), .A3(_u10_u7_n2742 ), .ZN(_u10_u7_n1896 ) );
OR3_X1 _u10_u7_U1446  ( .A1(_u10_u7_n2156 ), .A2(1'b0), .A3(_u10_u7_n1896 ),.ZN(_u10_u7_n2905 ) );
NAND2_X1 _u10_u7_U1445  ( .A1(_u10_u7_n2113 ), .A2(_u10_u7_n2996 ), .ZN(_u10_u7_n2719 ) );
NOR2_X1 _u10_u7_U1444  ( .A1(_u10_u7_n2719 ), .A2(1'b0), .ZN(_u10_u7_n2941 ));
INV_X1 _u10_u7_U1443  ( .A(_u10_u7_n2941 ), .ZN(_u10_u7_n2911 ) );
NOR2_X1 _u10_u7_U1442  ( .A1(_u10_u7_n2905 ), .A2(_u10_u7_n2911 ), .ZN(_u10_u7_n3222 ) );
INV_X1 _u10_u7_U1441  ( .A(_u10_u7_n3222 ), .ZN(_u10_u7_n2695 ) );
INV_X1 _u10_u7_U1440  ( .A(_u10_u7_n2156 ), .ZN(_u10_u7_n2089 ) );
NAND3_X1 _u10_u7_U1439  ( .A1(_u10_u7_n2089 ), .A2(_u10_u7_n2446 ), .A3(_u10_u7_n3180 ), .ZN(_u10_u7_n2902 ) );
NOR2_X1 _u10_u7_U1438  ( .A1(_u10_u7_n2902 ), .A2(_u10_u7_n2911 ), .ZN(_u10_u7_n2533 ) );
INV_X1 _u10_u7_U1437  ( .A(_u10_u7_n2533 ), .ZN(_u10_u7_n2485 ) );
NAND2_X1 _u10_u7_U1436  ( .A1(_u10_u7_n2695 ), .A2(_u10_u7_n2485 ), .ZN(_u10_u7_n2721 ) );
NAND2_X1 _u10_u7_U1435  ( .A1(1'b0), .A2(_u10_u7_n2113 ), .ZN(_u10_u7_n1868 ) );
INV_X1 _u10_u7_U1434  ( .A(_u10_u7_n1868 ), .ZN(_u10_u7_n2534 ) );
NOR2_X1 _u10_u7_U1433  ( .A1(_u10_u7_n2721 ), .A2(_u10_u7_n2534 ), .ZN(_u10_u7_n3231 ) );
NAND2_X1 _u10_u7_U1432  ( .A1(_u10_u7_n2467 ), .A2(_u10_u7_n3001 ), .ZN(_u10_u7_n2303 ) );
INV_X1 _u10_u7_U1431  ( .A(_u10_u7_n2303 ), .ZN(_u10_u7_n2549 ) );
INV_X1 _u10_u7_U1430  ( .A(1'b0), .ZN(_u10_u7_n2803 ) );
NAND2_X1 _u10_u7_U1429  ( .A1(_u10_u7_n2803 ), .A2(_u10_u7_n2446 ), .ZN(_u10_u7_n1846 ) );
INV_X1 _u10_u7_U1428  ( .A(_u10_u7_n1846 ), .ZN(_u10_u7_n2667 ) );
NAND3_X1 _u10_u7_U1427  ( .A1(_u10_u7_n2549 ), .A2(_u10_u7_n2667 ), .A3(1'b0), .ZN(_u10_u7_n2739 ) );
INV_X1 _u10_u7_U1426  ( .A(_u10_u7_n2739 ), .ZN(_u10_u7_n3272 ) );
INV_X1 _u10_u7_U1425  ( .A(_u10_u7_n2719 ), .ZN(_u10_u7_n2364 ) );
NAND2_X1 _u10_u7_U1424  ( .A1(_u10_u7_n3272 ), .A2(_u10_u7_n2364 ), .ZN(_u10_u7_n2852 ) );
INV_X1 _u10_u7_U1423  ( .A(_u10_u7_n2852 ), .ZN(_u10_u7_n2214 ) );
NAND2_X1 _u10_u7_U1422  ( .A1(_u10_u7_n2875 ), .A2(_u10_u7_n2089 ), .ZN(_u10_u7_n2097 ) );
INV_X1 _u10_u7_U1421  ( .A(_u10_u7_n2097 ), .ZN(_u10_u7_n2300 ) );
NAND2_X1 _u10_u7_U1420  ( .A1(_u10_u7_n2300 ), .A2(_u10_u7_n2446 ), .ZN(_u10_u7_n2001 ) );
NOR2_X1 _u10_u7_U1419  ( .A1(_u10_u7_n2001 ), .A2(_u10_u7_n2911 ), .ZN(_u10_u7_n2877 ) );
NOR2_X1 _u10_u7_U1418  ( .A1(_u10_u7_n2214 ), .A2(_u10_u7_n2877 ), .ZN(_u10_u7_n2940 ) );
NAND2_X1 _u10_u7_U1417  ( .A1(_u10_u7_n3231 ), .A2(_u10_u7_n2940 ), .ZN(_u10_u7_n3408 ) );
NAND2_X1 _u10_u7_U1416  ( .A1(_u10_u7_n2190 ), .A2(_u10_u7_n3408 ), .ZN(_u10_u7_n3402 ) );
NOR2_X1 _u10_u7_U1415  ( .A1(_u10_u7_n2446 ), .A2(_u10_u7_n2911 ), .ZN(_u10_u7_n3059 ) );
NAND2_X1 _u10_u7_U1414  ( .A1(_u10_u7_n3059 ), .A2(_u10_u7_n2190 ), .ZN(_u10_u7_n3404 ) );
AND3_X1 _u10_u7_U1413  ( .A1(_u10_u7_n3407 ), .A2(_u10_u7_n3226 ), .A3(_u10_u7_n3115 ), .ZN(_u10_u7_n3058 ) );
NAND2_X1 _u10_u7_U1412  ( .A1(_u10_u7_n3058 ), .A2(_u10_u7_n2022 ), .ZN(_u10_u7_n3406 ) );
NAND2_X1 _u10_u7_U1411  ( .A1(_u10_u7_n1853 ), .A2(_u10_u7_n3406 ), .ZN(_u10_u7_n3405 ) );
AND3_X1 _u10_u7_U1410  ( .A1(_u10_u7_n3404 ), .A2(_u10_u7_n1965 ), .A3(_u10_u7_n3405 ), .ZN(_u10_u7_n3063 ) );
NAND2_X1 _u10_u7_U1409  ( .A1(_u10_u7_n2667 ), .A2(_u10_u7_n3001 ), .ZN(_u10_u7_n1898 ) );
INV_X1 _u10_u7_U1408  ( .A(_u10_u7_n1898 ), .ZN(_u10_u7_n2835 ) );
NAND3_X1 _u10_u7_U1407  ( .A1(_u10_u7_n2364 ), .A2(_u10_u7_n2835 ), .A3(1'b0), .ZN(_u10_u7_n1869 ) );
NOR2_X1 _u10_u7_U1406  ( .A1(_u10_u7_n1869 ), .A2(_u10_u7_n2531 ), .ZN(_u10_u7_n2761 ) );
NOR3_X1 _u10_u7_U1405  ( .A1(_u10_u7_n2761 ), .A2(_u10_u7_n2528 ), .A3(_u10_u7_n2054 ), .ZN(_u10_u7_n3403 ) );
NAND4_X1 _u10_u7_U1404  ( .A1(_u10_u7_n3401 ), .A2(_u10_u7_n3402 ), .A3(_u10_u7_n3063 ), .A4(_u10_u7_n3403 ), .ZN(_u10_u7_n3400 ) );
NAND2_X1 _u10_u7_U1403  ( .A1(_u10_u7_n1966 ), .A2(_u10_u7_n3400 ), .ZN(_u10_u7_n3381 ) );
AND2_X1 _u10_u7_U1402  ( .A1(_u10_u7_n3368 ), .A2(_u10_SYNOPSYS_UNCONNECTED_33 ), .ZN(_u10_u7_n3319 ) );
NAND2_X1 _u10_u7_U1401  ( .A1(_u10_u7_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_32 ), .ZN(_u10_u7_n1849 ) );
INV_X1 _u10_u7_U1400  ( .A(_u10_u7_n1849 ), .ZN(_u10_u7_n2183 ) );
NAND2_X1 _u10_u7_U1399  ( .A1(_u10_u7_n2884 ), .A2(_u10_u7_n2183 ), .ZN(_u10_u7_n2883 ) );
INV_X1 _u10_u7_U1398  ( .A(_u10_u7_n2883 ), .ZN(_u10_u7_n1890 ) );
INV_X1 _u10_u7_U1397  ( .A(_u10_u7_n2940 ), .ZN(_u10_u7_n3278 ) );
NAND2_X1 _u10_u7_U1396  ( .A1(_u10_u7_n1890 ), .A2(_u10_u7_n3278 ), .ZN(_u10_u7_n3382 ) );
NAND2_X1 _u10_u7_U1395  ( .A1(_u10_u7_n3059 ), .A2(_u10_u7_n2669 ), .ZN(_u10_u7_n3399 ) );
NAND2_X1 _u10_u7_U1394  ( .A1(_u10_u7_n2031 ), .A2(_u10_u7_n3399 ), .ZN(_u10_u7_n3398 ) );
NAND2_X1 _u10_u7_U1393  ( .A1(_u10_u7_n2162 ), .A2(_u10_u7_n3398 ), .ZN(_u10_u7_n3395 ) );
NAND3_X1 _u10_u7_U1392  ( .A1(_u10_u7_n2747 ), .A2(_u10_u7_n2078 ), .A3(_u10_u7_n3126 ), .ZN(_u10_u7_n3396 ) );
NAND2_X1 _u10_u7_U1391  ( .A1(_u10_u7_n2055 ), .A2(_u10_u7_n2036 ), .ZN(_u10_u7_n2285 ) );
NOR2_X1 _u10_u7_U1390  ( .A1(_u10_u7_n2285 ), .A2(_u10_u7_n2030 ), .ZN(_u10_u7_n3349 ) );
INV_X1 _u10_u7_U1389  ( .A(_u10_u7_n3349 ), .ZN(_u10_u7_n1933 ) );
INV_X1 _u10_u7_U1388  ( .A(_u10_u7_n2710 ), .ZN(_u10_u7_n3397 ) );
NAND4_X1 _u10_u7_U1387  ( .A1(_u10_u7_n3395 ), .A2(_u10_u7_n3396 ), .A3(_u10_u7_n1933 ), .A4(_u10_u7_n3397 ), .ZN(_u10_u7_n3389 ) );
NAND2_X1 _u10_u7_U1386  ( .A1(_u10_u7_n1936 ), .A2(_u10_u7_n2828 ), .ZN(_u10_u7_n3141 ) );
INV_X1 _u10_u7_U1385  ( .A(_u10_u7_n3141 ), .ZN(_u10_u7_n2302 ) );
NAND2_X1 _u10_u7_U1384  ( .A1(_u10_u7_n3394 ), .A2(_u10_u7_n2302 ), .ZN(_u10_u7_n3390 ) );
NOR2_X1 _u10_u7_U1383  ( .A1(_u10_u7_n1869 ), .A2(_u10_u7_n2274 ), .ZN(_u10_u7_n3378 ) );
INV_X1 _u10_u7_U1382  ( .A(_u10_u7_n3378 ), .ZN(_u10_u7_n2748 ) );
NOR2_X1 _u10_u7_U1381  ( .A1(1'b0), .A2(_u10_u7_n2748 ), .ZN(_u10_u7_n3391 ));
NAND2_X1 _u10_u7_U1380  ( .A1(_u10_u7_n2534 ), .A2(_u10_u7_n2669 ), .ZN(_u10_u7_n2383 ) );
INV_X1 _u10_u7_U1379  ( .A(_u10_u7_n2383 ), .ZN(_u10_u7_n1978 ) );
NAND2_X1 _u10_u7_U1378  ( .A1(_u10_u7_n1978 ), .A2(_u10_u7_n2874 ), .ZN(_u10_u7_n3392 ) );
INV_X1 _u10_u7_U1377  ( .A(_u10_u7_n2411 ), .ZN(_u10_u7_n2164 ) );
NAND4_X1 _u10_u7_U1376  ( .A1(_u10_u7_n3392 ), .A2(_u10_u7_n3393 ), .A3(_u10_u7_n2033 ), .A4(_u10_u7_n2164 ), .ZN(_u10_u7_n2476 ) );
NOR4_X1 _u10_u7_U1375  ( .A1(_u10_u7_n3389 ), .A2(_u10_u7_n3390 ), .A3(_u10_u7_n3391 ), .A4(_u10_u7_n2476 ), .ZN(_u10_u7_n3388 ) );
NAND2_X1 _u10_u7_U1374  ( .A1(_u10_u7_n3236 ), .A2(_u10_u7_n3328 ), .ZN(_u10_u7_n2025 ) );
NOR2_X1 _u10_u7_U1373  ( .A1(_u10_u7_n3388 ), .A2(_u10_u7_n2025 ), .ZN(_u10_u7_n3384 ) );
NOR2_X1 _u10_u7_U1372  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u7_n2152 ) );
NAND2_X1 _u10_u7_U1371  ( .A1(_u10_u7_n2152 ), .A2(_u10_u7_n2175 ), .ZN(_u10_u7_n2722 ) );
INV_X1 _u10_u7_U1370  ( .A(_u10_u7_n2722 ), .ZN(_u10_u7_n2588 ) );
NAND2_X1 _u10_u7_U1369  ( .A1(_u10_u7_n2549 ), .A2(_u10_u7_n3349 ), .ZN(_u10_u7_n2091 ) );
NOR2_X1 _u10_u7_U1368  ( .A1(_u10_u7_n2091 ), .A2(_u10_u7_n1846 ), .ZN(_u10_u7_n2128 ) );
NAND3_X1 _u10_u7_U1367  ( .A1(_u10_u7_n3066 ), .A2(_u10_u7_n2113 ), .A3(_u10_u7_n2128 ), .ZN(_u10_u7_n2342 ) );
INV_X1 _u10_u7_U1366  ( .A(_u10_u7_n2342 ), .ZN(_u10_u7_n3316 ) );
NAND2_X1 _u10_u7_U1365  ( .A1(_u10_u7_n2588 ), .A2(_u10_u7_n3316 ), .ZN(_u10_u7_n2142 ) );
NOR2_X1 _u10_u7_U1364  ( .A1(_u10_u7_n1954 ), .A2(_u10_u7_n1898 ), .ZN(_u10_u7_n2255 ) );
NAND2_X1 _u10_u7_U1363  ( .A1(_u10_u7_n2255 ), .A2(_u10_u7_n2996 ), .ZN(_u10_u7_n1915 ) );
INV_X1 _u10_u7_U1362  ( .A(_u10_u7_n1915 ), .ZN(_u10_u7_n2251 ) );
NAND2_X1 _u10_u7_U1361  ( .A1(_u10_u7_n2251 ), .A2(_u10_u7_n2113 ), .ZN(_u10_u7_n1925 ) );
INV_X1 _u10_u7_U1360  ( .A(_u10_u7_n2026 ), .ZN(_u10_u7_n3340 ) );
NOR3_X1 _u10_u7_U1359  ( .A1(_u10_u7_n1925 ), .A2(_u10_u7_n2216 ), .A3(_u10_u7_n3340 ), .ZN(_u10_u7_n2003 ) );
INV_X1 _u10_u7_U1358  ( .A(1'b0), .ZN(_u10_u7_n1930 ) );
NAND2_X1 _u10_u7_U1357  ( .A1(_u10_u7_n2003 ), .A2(_u10_u7_n1930 ), .ZN(_u10_u7_n3387 ) );
AND2_X1 _u10_u7_U1356  ( .A1(_u10_u7_n2142 ), .A2(_u10_u7_n3387 ), .ZN(_u10_u7_n3366 ) );
NOR3_X1 _u10_u7_U1355  ( .A1(_u10_u7_n1813 ), .A2(_u10_u7_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_29 ), .ZN(_u10_u7_n3360 ) );
NOR2_X1 _u10_u7_U1354  ( .A1(_u10_SYNOPSYS_UNCONNECTED_31 ), .A2(_u10_SYNOPSYS_UNCONNECTED_32 ), .ZN(_u10_u7_n3136 ) );
NAND2_X1 _u10_u7_U1353  ( .A1(_u10_u7_n3360 ), .A2(_u10_u7_n3136 ), .ZN(_u10_u7_n2344 ) );
NOR2_X1 _u10_u7_U1352  ( .A1(_u10_u7_n3366 ), .A2(_u10_u7_n2344 ), .ZN(_u10_u7_n3385 ) );
NOR3_X1 _u10_u7_U1351  ( .A1(_u10_SYNOPSYS_UNCONNECTED_29 ), .A2(_u10_u7_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_33 ), .ZN(_u10_u7_n3342 ) );
NAND2_X1 _u10_u7_U1350  ( .A1(_u10_u7_n3342 ), .A2(_u10_u7_n3136 ), .ZN(_u10_u7_n2584 ) );
NOR2_X1 _u10_u7_U1349  ( .A1(_u10_u7_n2584 ), .A2(1'b0), .ZN(_u10_u7_n2139 ));
INV_X1 _u10_u7_U1348  ( .A(_u10_u7_n2216 ), .ZN(_u10_u7_n2106 ) );
AND2_X1 _u10_u7_U1347  ( .A1(_u10_u7_n2152 ), .A2(_u10_u7_n2106 ), .ZN(_u10_u7_n2336 ) );
NAND2_X1 _u10_u7_U1346  ( .A1(_u10_u7_n2139 ), .A2(_u10_u7_n2336 ), .ZN(_u10_u7_n2365 ) );
INV_X1 _u10_u7_U1345  ( .A(_u10_u7_n2365 ), .ZN(_u10_u7_n2004 ) );
AND2_X1 _u10_u7_U1344  ( .A1(_u10_u7_n2877 ), .A2(_u10_u7_n2004 ), .ZN(_u10_u7_n3386 ) );
NOR3_X1 _u10_u7_U1343  ( .A1(_u10_u7_n3384 ), .A2(_u10_u7_n3385 ), .A3(_u10_u7_n3386 ), .ZN(_u10_u7_n3383 ) );
NAND4_X1 _u10_u7_U1342  ( .A1(_u10_u7_n3380 ), .A2(_u10_u7_n3381 ), .A3(_u10_u7_n3382 ), .A4(_u10_u7_n3383 ), .ZN(_u10_u7_n3191 ) );
NAND2_X1 _u10_u7_U1341  ( .A1(_u10_u7_n2285 ), .A2(_u10_u7_n3379 ), .ZN(_u10_u7_n1975 ) );
NOR3_X1 _u10_u7_U1340  ( .A1(_u10_u7_n3378 ), .A2(1'b0), .A3(_u10_u7_n1975 ),.ZN(_u10_u7_n3122 ) );
AND4_X1 _u10_u7_U1339  ( .A1(_u10_u7_n2752 ), .A2(_u10_u7_n2383 ), .A3(_u10_u7_n1969 ), .A4(_u10_u7_n3122 ), .ZN(_u10_u7_n3377 ) );
NOR2_X1 _u10_u7_U1338  ( .A1(_u10_u7_n1814 ), .A2(_u10_u7_n1815 ), .ZN(_u10_u7_n3147 ) );
NAND2_X1 _u10_u7_U1337  ( .A1(_u10_u7_n3328 ), .A2(_u10_u7_n3147 ), .ZN(_u10_u7_n2359 ) );
NOR2_X1 _u10_u7_U1336  ( .A1(_u10_u7_n3377 ), .A2(_u10_u7_n2359 ), .ZN(_u10_u7_n3362 ) );
INV_X1 _u10_u7_U1335  ( .A(_u10_u7_n2008 ), .ZN(_u10_u7_n3097 ) );
NOR3_X1 _u10_u7_U1334  ( .A1(_u10_SYNOPSYS_UNCONNECTED_29 ), .A2(_u10_u7_n1813 ), .A3(_u10_SYNOPSYS_UNCONNECTED_30 ), .ZN(_u10_u7_n3269 ) );
NAND2_X1 _u10_u7_U1333  ( .A1(_u10_u7_n3269 ), .A2(_u10_u7_n3136 ), .ZN(_u10_u7_n3109 ) );
INV_X1 _u10_u7_U1332  ( .A(_u10_u7_n3109 ), .ZN(_u10_u7_n2999 ) );
INV_X1 _u10_u7_U1331  ( .A(_u10_u7_n2508 ), .ZN(_u10_u7_n2103 ) );
NAND2_X1 _u10_u7_U1330  ( .A1(_u10_u7_n2336 ), .A2(_u10_u7_n2103 ), .ZN(_u10_u7_n2249 ) );
NOR2_X1 _u10_u7_U1329  ( .A1(_u10_u7_n2249 ), .A2(1'b0), .ZN(_u10_u7_n1866 ));
NAND2_X1 _u10_u7_U1328  ( .A1(_u10_u7_n1866 ), .A2(_u10_u7_n1922 ), .ZN(_u10_u7_n2632 ) );
INV_X1 _u10_u7_U1327  ( .A(_u10_u7_n2223 ), .ZN(_u10_u7_n1918 ) );
NOR2_X1 _u10_u7_U1326  ( .A1(_u10_u7_n2632 ), .A2(_u10_u7_n1918 ), .ZN(_u10_u7_n1981 ) );
NAND3_X1 _u10_u7_U1325  ( .A1(_u10_u7_n3097 ), .A2(_u10_u7_n2999 ), .A3(_u10_u7_n1981 ), .ZN(_u10_u7_n3034 ) );
NOR3_X1 _u10_u7_U1324  ( .A1(_u10_SYNOPSYS_UNCONNECTED_30 ), .A2(_u10_SYNOPSYS_UNCONNECTED_29 ), .A3(_u10_SYNOPSYS_UNCONNECTED_33 ),.ZN(_u10_u7_n3302 ) );
NAND2_X1 _u10_u7_U1323  ( .A1(_u10_u7_n3302 ), .A2(_u10_u7_n3174 ), .ZN(_u10_u7_n3162 ) );
INV_X1 _u10_u7_U1322  ( .A(_u10_u7_n3162 ), .ZN(_u10_u7_n2979 ) );
NAND2_X1 _u10_u7_U1321  ( .A1(_u10_u7_n2979 ), .A2(_u10_u7_n2972 ), .ZN(_u10_u7_n1984 ) );
AND2_X1 _u10_u7_U1320  ( .A1(_u10_u7_n3302 ), .A2(_u10_u7_n3136 ), .ZN(_u10_u7_n2977 ) );
NAND3_X1 _u10_u7_U1319  ( .A1(_u10_u7_n2977 ), .A2(_u10_u7_n3000 ), .A3(_u10_u7_n3097 ), .ZN(_u10_u7_n3376 ) );
NAND2_X1 _u10_u7_U1318  ( .A1(_u10_u7_n1984 ), .A2(_u10_u7_n3376 ), .ZN(_u10_u7_n3375 ) );
NAND2_X1 _u10_u7_U1317  ( .A1(_u10_u7_n1981 ), .A2(_u10_u7_n3375 ), .ZN(_u10_u7_n2798 ) );
NAND2_X1 _u10_u7_U1316  ( .A1(_u10_u7_n3034 ), .A2(_u10_u7_n2798 ), .ZN(_u10_u7_n2007 ) );
NAND2_X1 _u10_u7_U1315  ( .A1(_u10_u7_n3269 ), .A2(_u10_u7_n3147 ), .ZN(_u10_u7_n2102 ) );
NOR2_X1 _u10_u7_U1314  ( .A1(_u10_u7_n2249 ), .A2(_u10_u7_n2102 ), .ZN(_u10_u7_n3323 ) );
INV_X1 _u10_u7_U1313  ( .A(_u10_u7_n3323 ), .ZN(_u10_u7_n3374 ) );
INV_X1 _u10_u7_U1312  ( .A(_u10_u7_n2344 ), .ZN(_u10_u7_n2002 ) );
NAND2_X1 _u10_u7_U1311  ( .A1(_u10_u7_n2336 ), .A2(_u10_u7_n2002 ), .ZN(_u10_u7_n3225 ) );
NAND2_X1 _u10_u7_U1310  ( .A1(_u10_u7_n3374 ), .A2(_u10_u7_n3225 ), .ZN(_u10_u7_n2488 ) );
NAND2_X1 _u10_u7_U1309  ( .A1(_u10_u7_n3342 ), .A2(_u10_u7_n3236 ), .ZN(_u10_u7_n2253 ) );
NOR2_X1 _u10_u7_U1308  ( .A1(_u10_u7_n2253 ), .A2(1'b0), .ZN(_u10_u7_n1885 ));
NAND2_X1 _u10_u7_U1307  ( .A1(_u10_u7_n3360 ), .A2(_u10_u7_n3174 ), .ZN(_u10_u7_n2254 ) );
INV_X1 _u10_u7_U1306  ( .A(_u10_u7_n2254 ), .ZN(_u10_u7_n2986 ) );
NAND2_X1 _u10_u7_U1305  ( .A1(_u10_u7_n2106 ), .A2(_u10_u7_n2986 ), .ZN(_u10_u7_n1913 ) );
INV_X1 _u10_u7_U1304  ( .A(_u10_u7_n1913 ), .ZN(_u10_u7_n2377 ) );
OR4_X1 _u10_u7_U1303  ( .A1(_u10_u7_n2007 ), .A2(_u10_u7_n2488 ), .A3(_u10_u7_n1885 ), .A4(_u10_u7_n2377 ), .ZN(_u10_u7_n3373 ) );
NAND2_X1 _u10_u7_U1302  ( .A1(_u10_u7_n2534 ), .A2(_u10_u7_n3373 ), .ZN(_u10_u7_n3370 ) );
NAND2_X1 _u10_u7_U1301  ( .A1(_u10_u7_n3342 ), .A2(_u10_u7_n3174 ), .ZN(_u10_u7_n2037 ) );
NAND2_X1 _u10_u7_U1300  ( .A1(_u10_u7_n2037 ), .A2(_u10_u7_n2254 ), .ZN(_u10_u7_n3372 ) );
NAND2_X1 _u10_u7_U1299  ( .A1(_u10_u7_n2003 ), .A2(_u10_u7_n3372 ), .ZN(_u10_u7_n3371 ) );
NAND2_X1 _u10_u7_U1298  ( .A1(_u10_u7_n3370 ), .A2(_u10_u7_n3371 ), .ZN(_u10_u7_n3363 ) );
NOR2_X1 _u10_u7_U1297  ( .A1(_u10_u7_n2490 ), .A2(_u10_u7_n1961 ), .ZN(_u10_u7_n3369 ) );
NAND2_X1 _u10_u7_U1296  ( .A1(_u10_u7_n2534 ), .A2(_u10_u7_n2049 ), .ZN(_u10_u7_n2646 ) );
INV_X1 _u10_u7_U1295  ( .A(_u10_u7_n2646 ), .ZN(_u10_u7_n3055 ) );
NOR2_X1 _u10_u7_U1294  ( .A1(_u10_u7_n3369 ), .A2(_u10_u7_n3055 ), .ZN(_u10_u7_n3367 ) );
NAND2_X1 _u10_u7_U1293  ( .A1(_u10_u7_n3368 ), .A2(_u10_u7_n3147 ), .ZN(_u10_u7_n2495 ) );
NOR2_X1 _u10_u7_U1292  ( .A1(_u10_u7_n3367 ), .A2(_u10_u7_n2495 ), .ZN(_u10_u7_n3364 ) );
INV_X1 _u10_u7_U1291  ( .A(_u10_u7_n2139 ), .ZN(_u10_u7_n3254 ) );
NOR2_X1 _u10_u7_U1290  ( .A1(_u10_u7_n3366 ), .A2(_u10_u7_n3254 ), .ZN(_u10_u7_n3365 ) );
NOR4_X1 _u10_u7_U1289  ( .A1(_u10_u7_n3362 ), .A2(_u10_u7_n3363 ), .A3(_u10_u7_n3364 ), .A4(_u10_u7_n3365 ), .ZN(_u10_u7_n3305 ) );
NAND2_X1 _u10_u7_U1288  ( .A1(_u10_u7_n3302 ), .A2(_u10_u7_n3147 ), .ZN(_u10_u7_n2980 ) );
NAND2_X1 _u10_u7_U1287  ( .A1(_u10_u7_n2102 ), .A2(_u10_u7_n2980 ), .ZN(_u10_u7_n2177 ) );
NAND2_X1 _u10_u7_U1286  ( .A1(_u10_u7_n2003 ), .A2(_u10_u7_n2493 ), .ZN(_u10_u7_n1962 ) );
NAND2_X1 _u10_u7_U1285  ( .A1(_u10_u7_n1961 ), .A2(_u10_u7_n1962 ), .ZN(_u10_u7_n3361 ) );
NAND2_X1 _u10_u7_U1284  ( .A1(_u10_u7_n2177 ), .A2(_u10_u7_n3361 ), .ZN(_u10_u7_n3357 ) );
NAND2_X1 _u10_u7_U1283  ( .A1(_u10_u7_n3236 ), .A2(_u10_u7_n3360 ), .ZN(_u10_u7_n1859 ) );
INV_X1 _u10_u7_U1282  ( .A(_u10_u7_n1859 ), .ZN(_u10_u7_n2256 ) );
NAND3_X1 _u10_u7_U1281  ( .A1(_u10_u7_n2256 ), .A2(_u10_u7_n2113 ), .A3(_u10_u7_n2128 ), .ZN(_u10_u7_n3358 ) );
NOR2_X1 _u10_u7_U1280  ( .A1(_u10_u7_n2877 ), .A2(_u10_u7_n3222 ), .ZN(_u10_u7_n3347 ) );
NAND2_X1 _u10_u7_U1279  ( .A1(_u10_u7_n3347 ), .A2(_u10_u7_n1869 ), .ZN(_u10_u7_n2005 ) );
NAND2_X1 _u10_u7_U1278  ( .A1(_u10_u7_n2488 ), .A2(_u10_u7_n2005 ), .ZN(_u10_u7_n3359 ) );
NAND3_X1 _u10_u7_U1277  ( .A1(_u10_u7_n3357 ), .A2(_u10_u7_n3358 ), .A3(_u10_u7_n3359 ), .ZN(_u10_u7_n3352 ) );
NAND2_X1 _u10_u7_U1276  ( .A1(_u10_u7_n3320 ), .A2(_u10_u7_n3136 ), .ZN(_u10_u7_n2356 ) );
INV_X1 _u10_u7_U1275  ( .A(_u10_u7_n2356 ), .ZN(_u10_u7_n2830 ) );
NAND2_X1 _u10_u7_U1274  ( .A1(_u10_u7_n2830 ), .A2(_u10_u7_n2836 ), .ZN(_u10_u7_n2291 ) );
NOR3_X1 _u10_u7_U1273  ( .A1(_u10_u7_n2291 ), .A2(_u10_u7_n2330 ), .A3(_u10_u7_n2022 ), .ZN(_u10_u7_n3353 ) );
INV_X1 _u10_u7_U1272  ( .A(_u10_u7_n1925 ), .ZN(_u10_u7_n2105 ) );
AND2_X1 _u10_u7_U1271  ( .A1(_u10_u7_n2108 ), .A2(_u10_u7_n2105 ), .ZN(_u10_u7_n2915 ) );
INV_X1 _u10_u7_U1270  ( .A(_u10_u7_n2330 ), .ZN(_u10_u7_n2107 ) );
NAND2_X1 _u10_u7_U1269  ( .A1(_u10_u7_n2915 ), .A2(_u10_u7_n2107 ), .ZN(_u10_u7_n2203 ) );
INV_X1 _u10_u7_U1268  ( .A(_u10_u7_n2203 ), .ZN(_u10_u7_n1982 ) );
NAND2_X1 _u10_u7_U1267  ( .A1(_u10_u7_n1982 ), .A2(_u10_u7_n2536 ), .ZN(_u10_u7_n2587 ) );
INV_X1 _u10_u7_U1266  ( .A(_u10_u7_n2587 ), .ZN(_u10_u7_n2697 ) );
NAND3_X1 _u10_u7_U1265  ( .A1(_u10_u7_n2697 ), .A2(_u10_u7_n2493 ), .A3(_u10_u7_n2377 ), .ZN(_u10_u7_n2412 ) );
INV_X1 _u10_u7_U1264  ( .A(_u10_u7_n2412 ), .ZN(_u10_u7_n3354 ) );
NAND2_X1 _u10_u7_U1263  ( .A1(_u10_u7_n3174 ), .A2(_u10_u7_n3269 ), .ZN(_u10_u7_n2375 ) );
INV_X1 _u10_u7_U1262  ( .A(_u10_u7_n2375 ), .ZN(_u10_u7_n2507 ) );
NAND2_X1 _u10_u7_U1261  ( .A1(_u10_u7_n1981 ), .A2(_u10_u7_n2507 ), .ZN(_u10_u7_n2621 ) );
NOR4_X1 _u10_u7_U1260  ( .A1(1'b0), .A2(_u10_u7_n3356 ), .A3(_u10_u7_n2203 ),.A4(_u10_u7_n2621 ), .ZN(_u10_u7_n3355 ) );
NOR4_X1 _u10_u7_U1259  ( .A1(_u10_u7_n3352 ), .A2(_u10_u7_n3353 ), .A3(_u10_u7_n3354 ), .A4(_u10_u7_n3355 ), .ZN(_u10_u7_n3306 ) );
NOR2_X1 _u10_u7_U1258  ( .A1(_u10_u7_n2842 ), .A2(_u10_u7_n2356 ), .ZN(_u10_u7_n1891 ) );
INV_X1 _u10_u7_U1257  ( .A(_u10_u7_n1869 ), .ZN(_u10_u7_n2885 ) );
NAND2_X1 _u10_u7_U1256  ( .A1(_u10_u7_n1891 ), .A2(_u10_u7_n2885 ), .ZN(_u10_u7_n3330 ) );
NAND2_X1 _u10_u7_U1255  ( .A1(_u10_u7_n2761 ), .A2(_u10_u7_n2837 ), .ZN(_u10_u7_n3351 ) );
NAND3_X1 _u10_u7_U1254  ( .A1(_u10_u7_n2884 ), .A2(_u10_u7_n2080 ), .A3(_u10_u7_n2915 ), .ZN(_u10_u7_n2762 ) );
NAND2_X1 _u10_u7_U1253  ( .A1(_u10_u7_n2055 ), .A2(_u10_u7_n2019 ), .ZN(_u10_u7_n3259 ) );
NAND4_X1 _u10_u7_U1252  ( .A1(_u10_u7_n3351 ), .A2(_u10_u7_n2762 ), .A3(_u10_u7_n2061 ), .A4(_u10_u7_n3259 ), .ZN(_u10_u7_n3350 ) );
NAND2_X1 _u10_u7_U1251  ( .A1(_u10_u7_n2183 ), .A2(_u10_u7_n3350 ), .ZN(_u10_u7_n3331 ) );
NAND2_X1 _u10_u7_U1250  ( .A1(_u10_u7_n3349 ), .A2(_u10_u7_n2305 ), .ZN(_u10_u7_n3348 ) );
NAND2_X1 _u10_u7_U1249  ( .A1(_u10_u7_n1896 ), .A2(_u10_u7_n3348 ), .ZN(_u10_u7_n3176 ) );
NAND2_X1 _u10_u7_U1248  ( .A1(_u10_u7_n2461 ), .A2(_u10_u7_n3176 ), .ZN(_u10_u7_n3332 ) );
INV_X1 _u10_u7_U1247  ( .A(_u10_u7_n2495 ), .ZN(_u10_u7_n2063 ) );
NAND2_X1 _u10_u7_U1246  ( .A1(_u10_u7_n2049 ), .A2(_u10_u7_n2063 ), .ZN(_u10_u7_n2886 ) );
NOR2_X1 _u10_u7_U1245  ( .A1(_u10_u7_n3347 ), .A2(_u10_u7_n2886 ), .ZN(_u10_u7_n3334 ) );
NAND2_X1 _u10_u7_U1244  ( .A1(1'b0), .A2(_u10_u7_n2835 ), .ZN(_u10_u7_n3344 ) );
NAND2_X1 _u10_u7_U1243  ( .A1(_u10_u7_n2001 ), .A2(_u10_u7_n2905 ), .ZN(_u10_u7_n3346 ) );
NAND2_X1 _u10_u7_U1242  ( .A1(_u10_u7_n3346 ), .A2(_u10_u7_n2803 ), .ZN(_u10_u7_n3345 ) );
NAND2_X1 _u10_u7_U1241  ( .A1(_u10_u7_n2087 ), .A2(_u10_u7_n2835 ), .ZN(_u10_u7_n2413 ) );
INV_X1 _u10_u7_U1240  ( .A(_u10_u7_n2128 ), .ZN(_u10_u7_n2235 ) );
NAND4_X1 _u10_u7_U1239  ( .A1(_u10_u7_n3344 ), .A2(_u10_u7_n3345 ), .A3(_u10_u7_n2413 ), .A4(_u10_u7_n2235 ), .ZN(_u10_u7_n3329 ) );
NOR2_X1 _u10_u7_U1238  ( .A1(_u10_u7_n1915 ), .A2(_u10_u7_n3340 ), .ZN(_u10_u7_n3343 ) );
NOR3_X1 _u10_u7_U1237  ( .A1(_u10_u7_n3329 ), .A2(1'b0), .A3(_u10_u7_n3343 ),.ZN(_u10_u7_n3341 ) );
NAND2_X1 _u10_u7_U1236  ( .A1(_u10_u7_n3342 ), .A2(_u10_u7_n3147 ), .ZN(_u10_u7_n2688 ) );
NOR2_X1 _u10_u7_U1235  ( .A1(_u10_u7_n3341 ), .A2(_u10_u7_n2688 ), .ZN(_u10_u7_n3335 ) );
NOR2_X1 _u10_u7_U1234  ( .A1(_u10_u7_n2256 ), .A2(_u10_u7_n1885 ), .ZN(_u10_u7_n2689 ) );
NOR2_X1 _u10_u7_U1233  ( .A1(1'b0), .A2(_u10_u7_n2413 ), .ZN(_u10_u7_n3338 ));
NOR2_X1 _u10_u7_U1232  ( .A1(_u10_u7_n1925 ), .A2(_u10_u7_n3340 ), .ZN(_u10_u7_n3339 ) );
NOR3_X1 _u10_u7_U1231  ( .A1(_u10_u7_n2005 ), .A2(_u10_u7_n3338 ), .A3(_u10_u7_n3339 ), .ZN(_u10_u7_n3337 ) );
NOR2_X1 _u10_u7_U1230  ( .A1(_u10_u7_n2689 ), .A2(_u10_u7_n3337 ), .ZN(_u10_u7_n3336 ) );
NOR3_X1 _u10_u7_U1229  ( .A1(_u10_u7_n3334 ), .A2(_u10_u7_n3335 ), .A3(_u10_u7_n3336 ), .ZN(_u10_u7_n3333 ) );
NAND4_X1 _u10_u7_U1228  ( .A1(_u10_u7_n3330 ), .A2(_u10_u7_n3331 ), .A3(_u10_u7_n3332 ), .A4(_u10_u7_n3333 ), .ZN(_u10_u7_n3308 ) );
NAND3_X1 _u10_u7_U1227  ( .A1(_u10_SYNOPSYS_UNCONNECTED_33 ), .A2(_u10_SYNOPSYS_UNCONNECTED_30 ), .A3(_u10_u7_n3147 ), .ZN(_u10_u7_n2126 ) );
INV_X1 _u10_u7_U1226  ( .A(_u10_u7_n2126 ), .ZN(_u10_u7_n2329 ) );
NAND2_X1 _u10_u7_U1225  ( .A1(_u10_u7_n2329 ), .A2(_u10_u7_n3329 ), .ZN(_u10_u7_n3324 ) );
NAND2_X1 _u10_u7_U1224  ( .A1(_u10_u7_n3328 ), .A2(_u10_u7_n3136 ), .ZN(_u10_u7_n2000 ) );
INV_X1 _u10_u7_U1223  ( .A(_u10_u7_n2000 ), .ZN(_u10_u7_n2445 ) );
NAND3_X1 _u10_u7_U1222  ( .A1(_u10_u7_n2446 ), .A2(_u10_u7_n3001 ), .A3(_u10_u7_n2087 ), .ZN(_u10_u7_n3327 ) );
NAND2_X1 _u10_u7_U1221  ( .A1(_u10_u7_n3327 ), .A2(_u10_u7_n2905 ), .ZN(_u10_u7_n2500 ) );
NAND2_X1 _u10_u7_U1220  ( .A1(_u10_u7_n2445 ), .A2(_u10_u7_n2500 ), .ZN(_u10_u7_n3325 ) );
NAND2_X1 _u10_u7_U1219  ( .A1(1'b0), .A2(_u10_u7_n2979 ), .ZN(_u10_u7_n3326 ) );
NAND3_X1 _u10_u7_U1218  ( .A1(_u10_u7_n3324 ), .A2(_u10_u7_n3325 ), .A3(_u10_u7_n3326 ), .ZN(_u10_u7_n3309 ) );
AND2_X1 _u10_u7_U1217  ( .A1(_u10_u7_n2877 ), .A2(_u10_u7_n3223 ), .ZN(_u10_u7_n2858 ) );
NAND2_X1 _u10_u7_U1216  ( .A1(_u10_u7_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_31 ), .ZN(_u10_u7_n2346 ) );
INV_X1 _u10_u7_U1215  ( .A(_u10_u7_n2346 ), .ZN(_u10_u7_n2043 ) );
NAND2_X1 _u10_u7_U1214  ( .A1(_u10_u7_n2858 ), .A2(_u10_u7_n2043 ), .ZN(_u10_u7_n3321 ) );
NAND2_X1 _u10_u7_U1213  ( .A1(_u10_u7_n1982 ), .A2(_u10_u7_n2195 ), .ZN(_u10_u7_n3268 ) );
INV_X1 _u10_u7_U1212  ( .A(_u10_u7_n3268 ), .ZN(_u10_u7_n2222 ) );
NAND3_X1 _u10_u7_U1211  ( .A1(_u10_u7_n3323 ), .A2(_u10_u7_n3216 ), .A3(_u10_u7_n2222 ), .ZN(_u10_u7_n3322 ) );
NAND2_X1 _u10_u7_U1210  ( .A1(_u10_u7_n3321 ), .A2(_u10_u7_n3322 ), .ZN(_u10_u7_n2374 ) );
NAND2_X1 _u10_u7_U1209  ( .A1(_u10_u7_n3320 ), .A2(_u10_u7_n3174 ), .ZN(_u10_u7_n2014 ) );
NOR2_X1 _u10_u7_U1208  ( .A1(_u10_u7_n1841 ), .A2(_u10_u7_n2014 ), .ZN(_u10_u7_n2813 ) );
NAND2_X1 _u10_u7_U1207  ( .A1(_u10_u7_n2813 ), .A2(_u10_u7_n2534 ), .ZN(_u10_u7_n3310 ) );
NAND2_X1 _u10_u7_U1206  ( .A1(_u10_u7_n3319 ), .A2(_u10_u7_n3136 ), .ZN(_u10_u7_n1836 ) );
INV_X1 _u10_u7_U1205  ( .A(_u10_u7_n1836 ), .ZN(_u10_u7_n2815 ) );
NAND2_X1 _u10_u7_U1204  ( .A1(_u10_u7_n2534 ), .A2(_u10_u7_n3129 ), .ZN(_u10_u7_n2439 ) );
NAND2_X1 _u10_u7_U1203  ( .A1(_u10_u7_n2055 ), .A2(_u10_u7_n2107 ), .ZN(_u10_u7_n2062 ) );
NAND2_X1 _u10_u7_U1202  ( .A1(_u10_u7_n2439 ), .A2(_u10_u7_n2062 ), .ZN(_u10_u7_n3318 ) );
NAND2_X1 _u10_u7_U1201  ( .A1(_u10_u7_n2815 ), .A2(_u10_u7_n3318 ), .ZN(_u10_u7_n3311 ) );
NAND2_X1 _u10_u7_U1200  ( .A1(_u10_u7_n2986 ), .A2(_u10_u7_n2175 ), .ZN(_u10_u7_n3317 ) );
NAND2_X1 _u10_u7_U1199  ( .A1(_u10_u7_n2253 ), .A2(_u10_u7_n3317 ), .ZN(_u10_u7_n3157 ) );
NAND2_X1 _u10_u7_U1198  ( .A1(_u10_u7_n3316 ), .A2(_u10_u7_n3157 ), .ZN(_u10_u7_n3312 ) );
NOR2_X1 _u10_u7_U1197  ( .A1(_u10_u7_n2495 ), .A2(_u10_u7_n2194 ), .ZN(_u10_u7_n3314 ) );
NOR2_X1 _u10_u7_U1196  ( .A1(_u10_u7_n2375 ), .A2(_u10_u7_n2367 ), .ZN(_u10_u7_n3315 ) );
NOR2_X1 _u10_u7_U1195  ( .A1(_u10_u7_n3314 ), .A2(_u10_u7_n3315 ), .ZN(_u10_u7_n3313 ) );
NAND4_X1 _u10_u7_U1194  ( .A1(_u10_u7_n3310 ), .A2(_u10_u7_n3311 ), .A3(_u10_u7_n3312 ), .A4(_u10_u7_n3313 ), .ZN(_u10_u7_n2315 ) );
NOR4_X1 _u10_u7_U1193  ( .A1(_u10_u7_n3308 ), .A2(_u10_u7_n3309 ), .A3(_u10_u7_n2374 ), .A4(_u10_u7_n2315 ), .ZN(_u10_u7_n3307 ) );
NAND3_X1 _u10_u7_U1192  ( .A1(_u10_u7_n3305 ), .A2(_u10_u7_n3306 ), .A3(_u10_u7_n3307 ), .ZN(_u10_u7_n1987 ) );
AND2_X1 _u10_u7_U1191  ( .A1(1'b0), .A2(_u10_u7_n2977 ), .ZN(_u10_u7_n3240 ));
NAND2_X1 _u10_u7_U1190  ( .A1(_u10_u7_n1891 ), .A2(_u10_u7_n2534 ), .ZN(_u10_u7_n3303 ) );
NAND4_X1 _u10_u7_U1189  ( .A1(_u10_u7_n1982 ), .A2(_u10_u7_n2659 ), .A3(_u10_u7_n2256 ), .A4(_u10_u7_n2175 ), .ZN(_u10_u7_n3304 ) );
AND2_X1 _u10_u7_U1188  ( .A1(_u10_u7_n3303 ), .A2(_u10_u7_n3304 ), .ZN(_u10_u7_n2612 ) );
NAND2_X1 _u10_u7_U1187  ( .A1(_u10_u7_n3302 ), .A2(_u10_u7_n3236 ), .ZN(_u10_u7_n2985 ) );
OR2_X1 _u10_u7_U1186  ( .A1(_u10_u7_n2431 ), .A2(_u10_u7_n2985 ), .ZN(_u10_u7_n3299 ) );
OR2_X1 _u10_u7_U1185  ( .A1(_u10_u7_n2282 ), .A2(_u10_u7_n2359 ), .ZN(_u10_u7_n3300 ) );
NAND2_X1 _u10_u7_U1184  ( .A1(_u10_u7_n1890 ), .A2(_u10_u7_n2534 ), .ZN(_u10_u7_n3301 ) );
NAND4_X1 _u10_u7_U1183  ( .A1(_u10_u7_n2612 ), .A2(_u10_u7_n3299 ), .A3(_u10_u7_n3300 ), .A4(_u10_u7_n3301 ), .ZN(_u10_u7_n3279 ) );
INV_X1 _u10_u7_U1182  ( .A(_u10_u7_n2464 ), .ZN(_u10_u7_n3295 ) );
NAND2_X1 _u10_u7_U1181  ( .A1(_u10_u7_n3295 ), .A2(_u10_u7_n2835 ), .ZN(_u10_u7_n2623 ) );
INV_X1 _u10_u7_U1180  ( .A(_u10_u7_n2623 ), .ZN(_u10_u7_n3185 ) );
INV_X1 _u10_u7_U1179  ( .A(_u10_u7_n2688 ), .ZN(_u10_u7_n2169 ) );
NAND2_X1 _u10_u7_U1178  ( .A1(_u10_u7_n3185 ), .A2(_u10_u7_n2169 ), .ZN(_u10_u7_n3286 ) );
NAND2_X1 _u10_u7_U1177  ( .A1(_u10_u7_n2833 ), .A2(_u10_u7_n3278 ), .ZN(_u10_u7_n3298 ) );
NAND3_X1 _u10_u7_U1176  ( .A1(_u10_u7_n3297 ), .A2(_u10_u7_n2838 ), .A3(_u10_u7_n3298 ), .ZN(_u10_u7_n3296 ) );
NAND2_X1 _u10_u7_U1175  ( .A1(_u10_u7_n2830 ), .A2(_u10_u7_n3296 ), .ZN(_u10_u7_n3287 ) );
NAND2_X1 _u10_u7_U1174  ( .A1(_u10_u7_n3295 ), .A2(_u10_u7_n3001 ), .ZN(_u10_u7_n3292 ) );
NAND2_X1 _u10_u7_U1173  ( .A1(_u10_u7_n3294 ), .A2(_u10_u7_n2089 ), .ZN(_u10_u7_n3293 ) );
AND2_X1 _u10_u7_U1172  ( .A1(_u10_u7_n3292 ), .A2(_u10_u7_n3293 ), .ZN(_u10_u7_n2548 ) );
NAND2_X1 _u10_u7_U1171  ( .A1(_u10_u7_n2548 ), .A2(_u10_u7_n2091 ), .ZN(_u10_u7_n2304 ) );
NAND2_X1 _u10_u7_U1170  ( .A1(_u10_u7_n2304 ), .A2(_u10_u7_n2446 ), .ZN(_u10_u7_n3290 ) );
NAND2_X1 _u10_u7_U1169  ( .A1(_u10_u7_n2549 ), .A2(_u10_u7_n2446 ), .ZN(_u10_u7_n2790 ) );
NOR2_X1 _u10_u7_U1168  ( .A1(_u10_u7_n1936 ), .A2(_u10_u7_n2790 ), .ZN(_u10_u7_n2789 ) );
INV_X1 _u10_u7_U1167  ( .A(_u10_u7_n2789 ), .ZN(_u10_u7_n3291 ) );
OR2_X1 _u10_u7_U1166  ( .A1(_u10_u7_n2828 ), .A2(_u10_u7_n2790 ), .ZN(_u10_u7_n2498 ) );
NAND4_X1 _u10_u7_U1165  ( .A1(_u10_u7_n3290 ), .A2(_u10_u7_n3291 ), .A3(_u10_u7_n2498 ), .A4(_u10_u7_n2001 ), .ZN(_u10_u7_n3289 ) );
NAND2_X1 _u10_u7_U1164  ( .A1(_u10_u7_n2445 ), .A2(_u10_u7_n3289 ), .ZN(_u10_u7_n3288 ) );
NAND3_X1 _u10_u7_U1163  ( .A1(_u10_u7_n3286 ), .A2(_u10_u7_n3287 ), .A3(_u10_u7_n3288 ), .ZN(_u10_u7_n3280 ) );
NOR2_X1 _u10_u7_U1162  ( .A1(_u10_u7_n2940 ), .A2(_u10_u7_n1913 ), .ZN(_u10_u7_n3281 ) );
INV_X1 _u10_u7_U1161  ( .A(1'b0), .ZN(_u10_u7_n1864 ) );
NAND2_X1 _u10_u7_U1160  ( .A1(1'b0), .A2(_u10_u7_n2588 ), .ZN(_u10_u7_n2141 ) );
INV_X1 _u10_u7_U1159  ( .A(_u10_u7_n2141 ), .ZN(_u10_u7_n3159 ) );
NAND3_X1 _u10_u7_U1158  ( .A1(_u10_u7_n2103 ), .A2(_u10_u7_n1864 ), .A3(_u10_u7_n3159 ), .ZN(_u10_u7_n2520 ) );
INV_X1 _u10_u7_U1157  ( .A(_u10_u7_n2520 ), .ZN(_u10_u7_n2630 ) );
INV_X1 _u10_u7_U1156  ( .A(_u10_u7_n2307 ), .ZN(_u10_u7_n2382 ) );
NOR4_X1 _u10_u7_U1155  ( .A1(_u10_u7_n2382 ), .A2(_u10_u7_n2722 ), .A3(_u10_u7_n1925 ), .A4(_u10_u7_n2508 ), .ZN(_u10_u7_n3260 ) );
NOR2_X1 _u10_u7_U1154  ( .A1(_u10_u7_n2498 ), .A2(_u10_u7_n2911 ), .ZN(_u10_u7_n2633 ) );
NOR2_X1 _u10_u7_U1153  ( .A1(_u10_u7_n2633 ), .A2(_u10_u7_n3278 ), .ZN(_u10_u7_n3285 ) );
INV_X1 _u10_u7_U1152  ( .A(_u10_u7_n1866 ), .ZN(_u10_u7_n1926 ) );
NOR2_X1 _u10_u7_U1151  ( .A1(_u10_u7_n3285 ), .A2(_u10_u7_n1926 ), .ZN(_u10_u7_n3284 ) );
NOR4_X1 _u10_u7_U1150  ( .A1(1'b0), .A2(_u10_u7_n2630 ), .A3(_u10_u7_n3260 ),.A4(_u10_u7_n3284 ), .ZN(_u10_u7_n3283 ) );
NOR2_X1 _u10_u7_U1149  ( .A1(_u10_u7_n3283 ), .A2(_u10_u7_n2980 ), .ZN(_u10_u7_n3282 ) );
NOR4_X1 _u10_u7_U1148  ( .A1(_u10_u7_n3279 ), .A2(_u10_u7_n3280 ), .A3(_u10_u7_n3281 ), .A4(_u10_u7_n3282 ), .ZN(_u10_u7_n3241 ) );
NAND2_X1 _u10_u7_U1147  ( .A1(_u10_u7_n1836 ), .A2(_u10_u7_n2291 ), .ZN(_u10_u7_n2147 ) );
NAND2_X1 _u10_u7_U1146  ( .A1(_u10_u7_n2443 ), .A2(_u10_u7_n2147 ), .ZN(_u10_u7_n3261 ) );
INV_X1 _u10_u7_U1145  ( .A(_u10_u7_n1841 ), .ZN(_u10_u7_n2571 ) );
NAND2_X1 _u10_u7_U1144  ( .A1(_u10_u7_n2571 ), .A2(_u10_u7_n3278 ), .ZN(_u10_u7_n3277 ) );
NAND2_X1 _u10_u7_U1143  ( .A1(_u10_u7_n3276 ), .A2(_u10_u7_n3277 ), .ZN(_u10_u7_n2819 ) );
OR2_X1 _u10_u7_U1142  ( .A1(_u10_u7_n2819 ), .A2(_u10_u7_n3275 ), .ZN(_u10_u7_n3273 ) );
NAND2_X1 _u10_u7_U1141  ( .A1(_u10_u7_n2815 ), .A2(_u10_u7_n2080 ), .ZN(_u10_u7_n3274 ) );
NAND2_X1 _u10_u7_U1140  ( .A1(_u10_u7_n2014 ), .A2(_u10_u7_n3274 ), .ZN(_u10_u7_n2165 ) );
NAND2_X1 _u10_u7_U1139  ( .A1(_u10_u7_n3273 ), .A2(_u10_u7_n2165 ), .ZN(_u10_u7_n3262 ) );
NAND2_X1 _u10_u7_U1138  ( .A1(_u10_u7_n2688 ), .A2(_u10_u7_n2126 ), .ZN(_u10_u7_n1956 ) );
INV_X1 _u10_u7_U1137  ( .A(_u10_u7_n1956 ), .ZN(_u10_u7_n1860 ) );
NOR2_X1 _u10_u7_U1136  ( .A1(1'b0), .A2(_u10_u7_n2498 ), .ZN(_u10_u7_n3271 ));
NOR2_X1 _u10_u7_U1135  ( .A1(_u10_u7_n3271 ), .A2(_u10_u7_n3272 ), .ZN(_u10_u7_n3270 ) );
NOR2_X1 _u10_u7_U1134  ( .A1(_u10_u7_n1860 ), .A2(_u10_u7_n3270 ), .ZN(_u10_u7_n3264 ) );
INV_X1 _u10_u7_U1133  ( .A(_u10_u7_n2632 ), .ZN(_u10_u7_n3202 ) );
NAND2_X1 _u10_u7_U1132  ( .A1(_u10_u7_n3236 ), .A2(_u10_u7_n3269 ), .ZN(_u10_u7_n3036 ) );
INV_X1 _u10_u7_U1131  ( .A(_u10_u7_n3036 ), .ZN(_u10_u7_n1960 ) );
NAND2_X1 _u10_u7_U1130  ( .A1(_u10_u7_n3202 ), .A2(_u10_u7_n1960 ), .ZN(_u10_u7_n3079 ) );
NOR3_X1 _u10_u7_U1129  ( .A1(_u10_u7_n3079 ), .A2(1'b0), .A3(_u10_u7_n3268 ),.ZN(_u10_u7_n3265 ) );
INV_X1 _u10_u7_U1128  ( .A(_u10_u7_n2014 ), .ZN(_u10_u7_n2709 ) );
NAND2_X1 _u10_u7_U1127  ( .A1(_u10_u7_n2709 ), .A2(_u10_u7_n2166 ), .ZN(_u10_u7_n2145 ) );
INV_X1 _u10_u7_U1126  ( .A(_u10_u7_n2145 ), .ZN(_u10_u7_n3258 ) );
NOR2_X1 _u10_u7_U1125  ( .A1(_u10_u7_n3258 ), .A2(_u10_u7_n2183 ), .ZN(_u10_u7_n3267 ) );
NOR2_X1 _u10_u7_U1124  ( .A1(_u10_u7_n3267 ), .A2(_u10_u7_n2567 ), .ZN(_u10_u7_n3266 ) );
NOR3_X1 _u10_u7_U1123  ( .A1(_u10_u7_n3264 ), .A2(_u10_u7_n3265 ), .A3(_u10_u7_n3266 ), .ZN(_u10_u7_n3263 ) );
NAND3_X1 _u10_u7_U1122  ( .A1(_u10_u7_n3261 ), .A2(_u10_u7_n3262 ), .A3(_u10_u7_n3263 ), .ZN(_u10_u7_n3243 ) );
INV_X1 _u10_u7_U1121  ( .A(_u10_u7_n2102 ), .ZN(_u10_u7_n2509 ) );
NAND2_X1 _u10_u7_U1120  ( .A1(_u10_u7_n3260 ), .A2(_u10_u7_n2509 ), .ZN(_u10_u7_n3247 ) );
INV_X1 _u10_u7_U1119  ( .A(_u10_u7_n3259 ), .ZN(_u10_u7_n2015 ) );
NAND2_X1 _u10_u7_U1118  ( .A1(_u10_u7_n2015 ), .A2(_u10_u7_n3258 ), .ZN(_u10_u7_n3248 ) );
NAND2_X1 _u10_u7_U1117  ( .A1(_u10_u7_n2251 ), .A2(_u10_u7_n2169 ), .ZN(_u10_u7_n3255 ) );
OR2_X1 _u10_u7_U1116  ( .A1(_u10_u7_n3157 ), .A2(_u10_u7_n2256 ), .ZN(_u10_u7_n3257 ) );
NAND2_X1 _u10_u7_U1115  ( .A1(_u10_u7_n2105 ), .A2(_u10_u7_n3257 ), .ZN(_u10_u7_n3256 ) );
AND2_X1 _u10_u7_U1114  ( .A1(_u10_u7_n3255 ), .A2(_u10_u7_n3256 ), .ZN(_u10_u7_n3212 ) );
INV_X1 _u10_u7_U1113  ( .A(_u10_u7_n2037 ), .ZN(_u10_u7_n2987 ) );
NAND2_X1 _u10_u7_U1112  ( .A1(_u10_u7_n2987 ), .A2(_u10_u7_n2038 ), .ZN(_u10_u7_n2212 ) );
NOR2_X1 _u10_u7_U1111  ( .A1(_u10_u7_n2212 ), .A2(1'b0), .ZN(_u10_u7_n2658 ));
INV_X1 _u10_u7_U1110  ( .A(_u10_u7_n2658 ), .ZN(_u10_u7_n2343 ) );
NAND2_X1 _u10_u7_U1109  ( .A1(_u10_u7_n2344 ), .A2(_u10_u7_n3254 ), .ZN(_u10_u7_n1928 ) );
NAND2_X1 _u10_u7_U1108  ( .A1(_u10_u7_n2588 ), .A2(_u10_u7_n1928 ), .ZN(_u10_u7_n3253 ) );
NAND2_X1 _u10_u7_U1107  ( .A1(_u10_u7_n2343 ), .A2(_u10_u7_n3253 ), .ZN(_u10_u7_n3252 ) );
NAND2_X1 _u10_u7_U1106  ( .A1(_u10_u7_n2105 ), .A2(_u10_u7_n3252 ), .ZN(_u10_u7_n3251 ) );
NAND2_X1 _u10_u7_U1105  ( .A1(_u10_u7_n3212 ), .A2(_u10_u7_n3251 ), .ZN(_u10_u7_n3250 ) );
NAND2_X1 _u10_u7_U1104  ( .A1(_u10_u7_n2307 ), .A2(_u10_u7_n3250 ), .ZN(_u10_u7_n3249 ) );
NAND3_X1 _u10_u7_U1103  ( .A1(_u10_u7_n3247 ), .A2(_u10_u7_n3248 ), .A3(_u10_u7_n3249 ), .ZN(_u10_u7_n3244 ) );
AND2_X1 _u10_u7_U1102  ( .A1(_u10_u7_n2915 ), .A2(_u10_u7_n2059 ), .ZN(_u10_u7_n2957 ) );
AND3_X1 _u10_u7_U1101  ( .A1(_u10_u7_n3223 ), .A2(_u10_u7_n2837 ), .A3(_u10_u7_n2957 ), .ZN(_u10_u7_n2051 ) );
NOR2_X1 _u10_u7_U1100  ( .A1(_u10_u7_n2528 ), .A2(_u10_u7_n2051 ), .ZN(_u10_u7_n2605 ) );
NOR2_X1 _u10_u7_U1099  ( .A1(_u10_u7_n2605 ), .A2(_u10_u7_n2346 ), .ZN(_u10_u7_n3245 ) );
NOR2_X1 _u10_u7_U1098  ( .A1(_u10_u7_n2291 ), .A2(_u10_u7_n2062 ), .ZN(_u10_u7_n3246 ) );
NOR4_X1 _u10_u7_U1097  ( .A1(_u10_u7_n3243 ), .A2(_u10_u7_n3244 ), .A3(_u10_u7_n3245 ), .A4(_u10_u7_n3246 ), .ZN(_u10_u7_n3242 ) );
NAND2_X1 _u10_u7_U1096  ( .A1(_u10_u7_n3241 ), .A2(_u10_u7_n3242 ), .ZN(_u10_u7_n2311 ) );
OR3_X1 _u10_u7_U1095  ( .A1(_u10_u7_n1987 ), .A2(_u10_u7_n3240 ), .A3(_u10_u7_n2311 ), .ZN(_u10_u7_n3192 ) );
INV_X1 _u10_u7_U1094  ( .A(_u10_u7_n2886 ), .ZN(_u10_u7_n2720 ) );
NOR2_X1 _u10_u7_U1093  ( .A1(_u10_u7_n2004 ), .A2(_u10_u7_n2720 ), .ZN(_u10_u7_n2455 ) );
INV_X1 _u10_u7_U1092  ( .A(_u10_u7_n2488 ), .ZN(_u10_u7_n2938 ) );
AND3_X1 _u10_u7_U1091  ( .A1(_u10_u7_n2455 ), .A2(_u10_u7_n1859 ), .A3(_u10_u7_n2938 ), .ZN(_u10_u7_n3239 ) );
INV_X1 _u10_u7_U1090  ( .A(_u10_u7_n2633 ), .ZN(_u10_u7_n2937 ) );
NOR2_X1 _u10_u7_U1089  ( .A1(_u10_u7_n3239 ), .A2(_u10_u7_n2937 ), .ZN(_u10_u7_n3227 ) );
NOR2_X1 _u10_u7_U1088  ( .A1(_u10_u7_n1976 ), .A2(_u10_u7_n1969 ), .ZN(_u10_u7_n3237 ) );
NOR2_X1 _u10_u7_U1087  ( .A1(1'b0), .A2(_u10_u7_n2947 ), .ZN(_u10_u7_n3238 ));
NOR3_X1 _u10_u7_U1086  ( .A1(_u10_u7_n2476 ), .A2(_u10_u7_n3237 ), .A3(_u10_u7_n3238 ), .ZN(_u10_u7_n3235 ) );
NOR3_X1 _u10_u7_U1085  ( .A1(_u10_u7_n1813 ), .A2(_u10_u7_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_30 ), .ZN(_u10_u7_n3135 ) );
NAND2_X1 _u10_u7_U1084  ( .A1(_u10_u7_n3135 ), .A2(_u10_u7_n3236 ), .ZN(_u10_u7_n2573 ) );
NOR2_X1 _u10_u7_U1083  ( .A1(_u10_u7_n3235 ), .A2(_u10_u7_n2573 ), .ZN(_u10_u7_n3228 ) );
NOR2_X1 _u10_u7_U1082  ( .A1(_u10_u7_n2216 ), .A2(_u10_u7_n1868 ), .ZN(_u10_u7_n3233 ) );
INV_X1 _u10_u7_U1081  ( .A(_u10_u7_n2550 ), .ZN(_u10_u7_n2475 ) );
NOR3_X1 _u10_u7_U1080  ( .A1(_u10_u7_n2475 ), .A2(1'b0), .A3(_u10_u7_n1925 ),.ZN(_u10_u7_n3234 ) );
NOR3_X1 _u10_u7_U1079  ( .A1(_u10_u7_n3233 ), .A2(1'b0), .A3(_u10_u7_n3234 ),.ZN(_u10_u7_n3232 ) );
NOR2_X1 _u10_u7_U1078  ( .A1(_u10_u7_n3232 ), .A2(_u10_u7_n2037 ), .ZN(_u10_u7_n3229 ) );
NOR2_X1 _u10_u7_U1077  ( .A1(_u10_u7_n3231 ), .A2(_u10_u7_n2365 ), .ZN(_u10_u7_n3230 ) );
NOR4_X1 _u10_u7_U1076  ( .A1(_u10_u7_n3227 ), .A2(_u10_u7_n3228 ), .A3(_u10_u7_n3229 ), .A4(_u10_u7_n3230 ), .ZN(_u10_u7_n3205 ) );
NOR3_X1 _u10_u7_U1075  ( .A1(_u10_u7_n3226 ), .A2(_u10_u7_n2687 ), .A3(_u10_u7_n2145 ), .ZN(_u10_u7_n3217 ) );
NOR3_X1 _u10_u7_U1074  ( .A1(_u10_u7_n3225 ), .A2(1'b0), .A3(_u10_u7_n2587 ),.ZN(_u10_u7_n3218 ) );
NOR2_X1 _u10_u7_U1073  ( .A1(_u10_u7_n3159 ), .A2(1'b0), .ZN(_u10_u7_n3224 ));
NOR2_X1 _u10_u7_U1072  ( .A1(_u10_u7_n3224 ), .A2(_u10_u7_n2584 ), .ZN(_u10_u7_n3219 ) );
NAND2_X1 _u10_u7_U1071  ( .A1(_u10_u7_n3222 ), .A2(_u10_u7_n3223 ), .ZN(_u10_u7_n2048 ) );
INV_X1 _u10_u7_U1070  ( .A(_u10_u7_n2048 ), .ZN(_u10_u7_n2859 ) );
NOR2_X1 _u10_u7_U1069  ( .A1(_u10_u7_n2859 ), .A2(_u10_u7_n2054 ), .ZN(_u10_u7_n3221 ) );
NOR2_X1 _u10_u7_U1068  ( .A1(_u10_u7_n3221 ), .A2(_u10_u7_n2346 ), .ZN(_u10_u7_n3220 ) );
NOR4_X1 _u10_u7_U1067  ( .A1(_u10_u7_n3217 ), .A2(_u10_u7_n3218 ), .A3(_u10_u7_n3219 ), .A4(_u10_u7_n3220 ), .ZN(_u10_u7_n3206 ) );
NAND2_X1 _u10_u7_U1066  ( .A1(_u10_u7_n2377 ), .A2(_u10_u7_n2721 ), .ZN(_u10_u7_n3213 ) );
AND4_X1 _u10_u7_U1065  ( .A1(1'b0), .A2(_u10_u7_n2502 ), .A3(_u10_u7_n2972 ),.A4(_u10_u7_n3040 ), .ZN(_u10_u7_n2406 ) );
NAND2_X1 _u10_u7_U1064  ( .A1(_u10_u7_n2406 ), .A2(_u10_u7_n2979 ), .ZN(_u10_u7_n3214 ) );
NAND2_X1 _u10_u7_U1063  ( .A1(_u10_u7_n2630 ), .A2(_u10_u7_n3216 ), .ZN(_u10_u7_n2376 ) );
INV_X1 _u10_u7_U1062  ( .A(_u10_u7_n2376 ), .ZN(_u10_u7_n3108 ) );
NAND2_X1 _u10_u7_U1061  ( .A1(_u10_u7_n3108 ), .A2(_u10_u7_n2507 ), .ZN(_u10_u7_n3215 ) );
NOR2_X1 _u10_u7_U1060  ( .A1(_u10_u7_n2937 ), .A2(1'b0), .ZN(_u10_u7_n2649 ));
INV_X1 _u10_u7_U1059  ( .A(_u10_u7_n2253 ), .ZN(_u10_u7_n2971 ) );
NAND2_X1 _u10_u7_U1058  ( .A1(_u10_u7_n2649 ), .A2(_u10_u7_n2971 ), .ZN(_u10_u7_n2918 ) );
NAND4_X1 _u10_u7_U1057  ( .A1(_u10_u7_n3213 ), .A2(_u10_u7_n3214 ), .A3(_u10_u7_n3215 ), .A4(_u10_u7_n2918 ), .ZN(_u10_u7_n3208 ) );
NOR2_X1 _u10_u7_U1056  ( .A1(_u10_u7_n2000 ), .A2(_u10_u7_n2902 ), .ZN(_u10_u7_n3209 ) );
NOR2_X1 _u10_u7_U1055  ( .A1(_u10_u7_n3212 ), .A2(_u10_u7_n2475 ), .ZN(_u10_u7_n3210 ) );
INV_X1 _u10_u7_U1054  ( .A(_u10_u7_n2441 ), .ZN(_u10_u7_n3128 ) );
NOR2_X1 _u10_u7_U1053  ( .A1(_u10_u7_n2356 ), .A2(_u10_u7_n3128 ), .ZN(_u10_u7_n3211 ) );
NOR4_X1 _u10_u7_U1052  ( .A1(_u10_u7_n3208 ), .A2(_u10_u7_n3209 ), .A3(_u10_u7_n3210 ), .A4(_u10_u7_n3211 ), .ZN(_u10_u7_n3207 ) );
NAND3_X1 _u10_u7_U1051  ( .A1(_u10_u7_n3205 ), .A2(_u10_u7_n3206 ), .A3(_u10_u7_n3207 ), .ZN(_u10_u7_n2611 ) );
NOR2_X1 _u10_u7_U1050  ( .A1(_u10_u7_n2212 ), .A2(_u10_u7_n2216 ), .ZN(_u10_u7_n1937 ) );
NOR2_X1 _u10_u7_U1049  ( .A1(_u10_u7_n2533 ), .A2(_u10_u7_n2214 ), .ZN(_u10_u7_n2765 ) );
INV_X1 _u10_u7_U1048  ( .A(_u10_u7_n2005 ), .ZN(_u10_u7_n2111 ) );
AND2_X1 _u10_u7_U1047  ( .A1(_u10_u7_n2765 ), .A2(_u10_u7_n2111 ), .ZN(_u10_u7_n3201 ) );
INV_X1 _u10_u7_U1046  ( .A(_u10_u7_n3059 ), .ZN(_u10_u7_n3076 ) );
NAND2_X1 _u10_u7_U1045  ( .A1(_u10_u7_n3201 ), .A2(_u10_u7_n3076 ), .ZN(_u10_u7_n3204 ) );
NAND2_X1 _u10_u7_U1044  ( .A1(_u10_u7_n1937 ), .A2(_u10_u7_n3204 ), .ZN(_u10_u7_n3193 ) );
NAND2_X1 _u10_u7_U1043  ( .A1(_u10_u7_n2254 ), .A2(_u10_u7_n2212 ), .ZN(_u10_u7_n3203 ) );
NAND3_X1 _u10_u7_U1042  ( .A1(_u10_u7_n3203 ), .A2(_u10_u7_n2175 ), .A3(_u10_u7_n2649 ), .ZN(_u10_u7_n3194 ) );
NOR2_X1 _u10_u7_U1041  ( .A1(_u10_u7_n2985 ), .A2(1'b0), .ZN(_u10_u7_n1959 ));
NAND2_X1 _u10_u7_U1040  ( .A1(_u10_u7_n1959 ), .A2(_u10_u7_n3202 ), .ZN(_u10_u7_n2202 ) );
NAND4_X1 _u10_u7_U1039  ( .A1(_u10_u7_n3079 ), .A2(_u10_u7_n2621 ), .A3(_u10_u7_n2202 ), .A4(_u10_u7_n2798 ), .ZN(_u10_u7_n3200 ) );
NAND2_X1 _u10_u7_U1038  ( .A1(_u10_u7_n3201 ), .A2(_u10_u7_n2937 ), .ZN(_u10_u7_n2772 ) );
NAND2_X1 _u10_u7_U1037  ( .A1(_u10_u7_n3200 ), .A2(_u10_u7_n2772 ), .ZN(_u10_u7_n3195 ) );
NAND2_X1 _u10_u7_U1036  ( .A1(_u10_u7_n2765 ), .A2(_u10_u7_n1869 ), .ZN(_u10_u7_n3199 ) );
NAND2_X1 _u10_u7_U1035  ( .A1(_u10_u7_n2049 ), .A2(_u10_u7_n3199 ), .ZN(_u10_u7_n3057 ) );
NOR2_X1 _u10_u7_U1034  ( .A1(_u10_u7_n2495 ), .A2(_u10_u7_n3057 ), .ZN(_u10_u7_n3197 ) );
NOR2_X1 _u10_u7_U1033  ( .A1(_u10_u7_n2883 ), .A2(_u10_u7_n2485 ), .ZN(_u10_u7_n3198 ) );
NOR2_X1 _u10_u7_U1032  ( .A1(_u10_u7_n3197 ), .A2(_u10_u7_n3198 ), .ZN(_u10_u7_n3196 ) );
NAND4_X1 _u10_u7_U1031  ( .A1(_u10_u7_n3193 ), .A2(_u10_u7_n3194 ), .A3(_u10_u7_n3195 ), .A4(_u10_u7_n3196 ), .ZN(_u10_u7_n2887 ) );
NOR4_X1 _u10_u7_U1030  ( .A1(_u10_u7_n3191 ), .A2(_u10_u7_n3192 ), .A3(_u10_u7_n2611 ), .A4(_u10_u7_n2887 ), .ZN(_u10_u7_n3015 ) );
NAND3_X1 _u10_u7_U1029  ( .A1(_u10_u7_n3190 ), .A2(_u10_u7_n2049 ), .A3(_u10_u7_n2957 ), .ZN(_u10_u7_n2699 ) );
OR2_X1 _u10_u7_U1028  ( .A1(_u10_u7_n2699 ), .A2(_u10_u7_n1813 ), .ZN(_u10_u7_n3187 ) );
NAND3_X1 _u10_u7_U1027  ( .A1(_u10_u7_n2978 ), .A2(_u10_u7_n2405 ), .A3(1'b0), .ZN(_u10_u7_n3188 ) );
NAND4_X1 _u10_u7_U1026  ( .A1(_u10_u7_n3058 ), .A2(_u10_u7_n3187 ), .A3(_u10_u7_n3188 ), .A4(_u10_u7_n3189 ), .ZN(_u10_u7_n3186 ) );
NAND2_X1 _u10_u7_U1025  ( .A1(_u10_u7_n2063 ), .A2(_u10_u7_n3186 ), .ZN(_u10_u7_n3163 ) );
NAND2_X1 _u10_u7_U1024  ( .A1(_u10_u7_n3185 ), .A2(_u10_u7_n2329 ), .ZN(_u10_u7_n3164 ) );
NAND2_X1 _u10_u7_U1023  ( .A1(_u10_u7_n2689 ), .A2(_u10_u7_n2365 ), .ZN(_u10_u7_n2736 ) );
NOR2_X1 _u10_u7_U1022  ( .A1(_u10_u7_n2736 ), .A2(_u10_u7_n2488 ), .ZN(_u10_u7_n1855 ) );
INV_X1 _u10_u7_U1021  ( .A(_u10_u7_n1855 ), .ZN(_u10_u7_n3184 ) );
NOR2_X1 _u10_u7_U1020  ( .A1(_u10_u7_n2274 ), .A2(_u10_u7_n2359 ), .ZN(_u10_u7_n2952 ) );
NOR2_X1 _u10_u7_U1019  ( .A1(_u10_u7_n3184 ), .A2(_u10_u7_n2952 ), .ZN(_u10_u7_n2776 ) );
OR2_X1 _u10_u7_U1018  ( .A1(_u10_u7_n2852 ), .A2(_u10_u7_n2776 ), .ZN(_u10_u7_n3165 ) );
NAND2_X1 _u10_u7_U1017  ( .A1(_u10_u7_n3126 ), .A2(_u10_u7_n2915 ), .ZN(_u10_u7_n3065 ) );
NOR3_X1 _u10_u7_U1016  ( .A1(_u10_u7_n3065 ), .A2(1'b0), .A3(_u10_u7_n2632 ),.ZN(_u10_u7_n3182 ) );
NOR3_X1 _u10_u7_U1015  ( .A1(_u10_u7_n3182 ), .A2(_u10_u7_n3183 ), .A3(_u10_u7_n3108 ), .ZN(_u10_u7_n3181 ) );
NOR2_X1 _u10_u7_U1014  ( .A1(_u10_u7_n3181 ), .A2(_u10_u7_n3162 ), .ZN(_u10_u7_n3167 ) );
INV_X1 _u10_u7_U1013  ( .A(_u10_u7_n3180 ), .ZN(_u10_u7_n3140 ) );
NAND3_X1 _u10_u7_U1012  ( .A1(_u10_u7_n3140 ), .A2(_u10_u7_n2163 ), .A3(_u10_u7_n2092 ), .ZN(_u10_u7_n3175 ) );
NOR4_X1 _u10_u7_U1011  ( .A1(_u10_u7_n2411 ), .A2(_u10_u7_n2710 ), .A3(_u10_u7_n3141 ), .A4(_u10_u7_n3089 ), .ZN(_u10_u7_n3179 ) );
NOR2_X1 _u10_u7_U1010  ( .A1(1'b0), .A2(_u10_u7_n3179 ), .ZN(_u10_u7_n3177 ));
NOR2_X1 _u10_u7_U1009  ( .A1(_u10_u7_n1898 ), .A2(_u10_u7_n1847 ), .ZN(_u10_u7_n3178 ) );
NOR4_X1 _u10_u7_U1008  ( .A1(_u10_u7_n3175 ), .A2(_u10_u7_n3176 ), .A3(_u10_u7_n3177 ), .A4(_u10_u7_n3178 ), .ZN(_u10_u7_n3173 ) );
NAND2_X1 _u10_u7_U1007  ( .A1(_u10_u7_n3135 ), .A2(_u10_u7_n3174 ), .ZN(_u10_u7_n2159 ) );
NOR2_X1 _u10_u7_U1006  ( .A1(_u10_u7_n3173 ), .A2(_u10_u7_n2159 ), .ZN(_u10_u7_n3168 ) );
OR3_X1 _u10_u7_U1005  ( .A1(_u10_u7_n3172 ), .A2(1'b0), .A3(_u10_u7_n3126 ),.ZN(_u10_u7_n3171 ) );
NAND2_X1 _u10_u7_U1004  ( .A1(_u10_u7_n2600 ), .A2(_u10_u7_n3171 ), .ZN(_u10_u7_n3153 ) );
AND3_X1 _u10_u7_U1003  ( .A1(_u10_u7_n3153 ), .A2(_u10_u7_n2947 ), .A3(_u10_u7_n2579 ), .ZN(_u10_u7_n3170 ) );
NOR2_X1 _u10_u7_U1002  ( .A1(_u10_u7_n3170 ), .A2(_u10_u7_n2359 ), .ZN(_u10_u7_n3169 ) );
NOR3_X1 _u10_u7_U1001  ( .A1(_u10_u7_n3167 ), .A2(_u10_u7_n3168 ), .A3(_u10_u7_n3169 ), .ZN(_u10_u7_n3166 ) );
NAND4_X1 _u10_u7_U1000  ( .A1(_u10_u7_n3163 ), .A2(_u10_u7_n3164 ), .A3(_u10_u7_n3165 ), .A4(_u10_u7_n3166 ), .ZN(_u10_u7_n3130 ) );
NAND2_X1 _u10_u7_U999  ( .A1(_u10_u7_n2375 ), .A2(_u10_u7_n3162 ), .ZN(_u10_u7_n1923 ) );
NAND2_X1 _u10_u7_U998  ( .A1(_u10_u7_n3062 ), .A2(_u10_u7_n1923 ), .ZN(_u10_u7_n3154 ) );
NAND2_X1 _u10_u7_U997  ( .A1(_u10_u7_n2103 ), .A2(_u10_u7_n2509 ), .ZN(_u10_u7_n3161 ) );
NAND2_X1 _u10_u7_U996  ( .A1(_u10_u7_n2344 ), .A2(_u10_u7_n3161 ), .ZN(_u10_u7_n3160 ) );
NAND2_X1 _u10_u7_U995  ( .A1(_u10_u7_n3159 ), .A2(_u10_u7_n3160 ), .ZN(_u10_u7_n2635 ) );
AND3_X1 _u10_u7_U994  ( .A1(_u10_u7_n2549 ), .A2(_u10_u7_n2108 ), .A3(_u10_u7_n3126 ), .ZN(_u10_u7_n3093 ) );
NAND2_X1 _u10_u7_U993  ( .A1(_u10_u7_n3093 ), .A2(_u10_u7_n2941 ), .ZN(_u10_u7_n3158 ) );
NAND3_X1 _u10_u7_U992  ( .A1(_u10_u7_n3076 ), .A2(_u10_u7_n3066 ), .A3(_u10_u7_n3158 ), .ZN(_u10_u7_n3156 ) );
NAND2_X1 _u10_u7_U991  ( .A1(_u10_u7_n3156 ), .A2(_u10_u7_n3157 ), .ZN(_u10_u7_n3155 ) );
NAND3_X1 _u10_u7_U990  ( .A1(_u10_u7_n3154 ), .A2(_u10_u7_n2635 ), .A3(_u10_u7_n3155 ), .ZN(_u10_u7_n3131 ) );
INV_X1 _u10_u7_U989  ( .A(_u10_u7_n2594 ), .ZN(_u10_u7_n2846 ) );
NAND3_X1 _u10_u7_U988  ( .A1(_u10_u7_n2162 ), .A2(_u10_u7_n2082 ), .A3(_u10_u7_n2105 ), .ZN(_u10_u7_n2077 ) );
NAND4_X1 _u10_u7_U987  ( .A1(_u10_u7_n3153 ), .A2(_u10_u7_n1969 ), .A3(_u10_u7_n2846 ), .A4(_u10_u7_n2077 ), .ZN(_u10_u7_n3148 ) );
NAND2_X1 _u10_u7_U986  ( .A1(_u10_u7_n2838 ), .A2(_u10_u7_n3128 ), .ZN(_u10_u7_n3152 ) );
NAND2_X1 _u10_u7_U985  ( .A1(_u10_u7_n3152 ), .A2(_u10_u7_n2600 ), .ZN(_u10_u7_n3151 ) );
NAND2_X1 _u10_u7_U984  ( .A1(_u10_u7_n2282 ), .A2(_u10_u7_n3151 ), .ZN(_u10_u7_n2601 ) );
NOR4_X1 _u10_u7_U983  ( .A1(_u10_u7_n2885 ), .A2(_u10_u7_n2534 ), .A3(_u10_u7_n2214 ), .A4(_u10_u7_n3059 ), .ZN(_u10_u7_n3150 ) );
NOR2_X1 _u10_u7_U982  ( .A1(_u10_u7_n3150 ), .A2(_u10_u7_n2853 ), .ZN(_u10_u7_n3149 ) );
NOR4_X1 _u10_u7_U981  ( .A1(_u10_u7_n3148 ), .A2(_u10_u7_n2601 ), .A3(_u10_u7_n3149 ), .A4(_u10_u7_n1975 ), .ZN(_u10_u7_n3146 ) );
NAND3_X1 _u10_u7_U980  ( .A1(_u10_SYNOPSYS_UNCONNECTED_33 ), .A2(_u10_SYNOPSYS_UNCONNECTED_29 ), .A3(_u10_u7_n3147 ), .ZN(_u10_u7_n2071 ) );
NOR2_X1 _u10_u7_U979  ( .A1(_u10_u7_n3146 ), .A2(_u10_u7_n2071 ), .ZN(_u10_u7_n3132 ) );
NOR2_X1 _u10_u7_U978  ( .A1(1'b0), .A2(_u10_u7_n1847 ), .ZN(_u10_u7_n3143 ));
INV_X1 _u10_u7_U977  ( .A(_u10_u7_n3145 ), .ZN(_u10_u7_n3144 ) );
NOR2_X1 _u10_u7_U976  ( .A1(_u10_u7_n3143 ), .A2(_u10_u7_n3144 ), .ZN(_u10_u7_n3142 ) );
NOR2_X1 _u10_u7_U975  ( .A1(1'b0), .A2(_u10_u7_n3142 ), .ZN(_u10_u7_n3137 ));
NAND2_X1 _u10_u7_U974  ( .A1(_u10_u7_n2549 ), .A2(_u10_u7_n3141 ), .ZN(_u10_u7_n3138 ) );
NAND2_X1 _u10_u7_U973  ( .A1(_u10_u7_n1896 ), .A2(_u10_u7_n3140 ), .ZN(_u10_u7_n2544 ) );
NAND2_X1 _u10_u7_U972  ( .A1(_u10_u7_n2089 ), .A2(_u10_u7_n2544 ), .ZN(_u10_u7_n3139 ) );
NAND2_X1 _u10_u7_U971  ( .A1(_u10_u7_n3138 ), .A2(_u10_u7_n3139 ), .ZN(_u10_u7_n2795 ) );
NOR4_X1 _u10_u7_U970  ( .A1(_u10_u7_n2300 ), .A2(_u10_u7_n3137 ), .A3(_u10_u7_n2304 ), .A4(_u10_u7_n2795 ), .ZN(_u10_u7_n3134 ) );
NAND2_X1 _u10_u7_U969  ( .A1(_u10_u7_n3135 ), .A2(_u10_u7_n3136 ), .ZN(_u10_u7_n2085 ) );
NOR2_X1 _u10_u7_U968  ( .A1(_u10_u7_n3134 ), .A2(_u10_u7_n2085 ), .ZN(_u10_u7_n3133 ) );
NOR4_X1 _u10_u7_U967  ( .A1(_u10_u7_n3130 ), .A2(_u10_u7_n3131 ), .A3(_u10_u7_n3132 ), .A4(_u10_u7_n3133 ), .ZN(_u10_u7_n3016 ) );
INV_X1 _u10_u7_U966  ( .A(_u10_u7_n2686 ), .ZN(_u10_u7_n2278 ) );
NAND4_X1 _u10_u7_U965  ( .A1(_u10_u7_n2105 ), .A2(_u10_u7_n2278 ), .A3(_u10_u7_n3129 ), .A4(_u10_u7_n2600 ), .ZN(_u10_u7_n2437 ) );
NAND2_X1 _u10_u7_U964  ( .A1(_u10_u7_n3128 ), .A2(_u10_u7_n2437 ), .ZN(_u10_u7_n3127 ) );
NAND2_X1 _u10_u7_U963  ( .A1(_u10_u7_n2815 ), .A2(_u10_u7_n3127 ), .ZN(_u10_u7_n3098 ) );
INV_X1 _u10_u7_U962  ( .A(_u10_u7_n2573 ), .ZN(_u10_u7_n1967 ) );
NAND2_X1 _u10_u7_U961  ( .A1(_u10_u7_n3126 ), .A2(_u10_u7_n2078 ), .ZN(_u10_u7_n3123 ) );
NAND2_X1 _u10_u7_U960  ( .A1(_u10_u7_n3076 ), .A2(_u10_u7_n1925 ), .ZN(_u10_u7_n3125 ) );
NAND2_X1 _u10_u7_U959  ( .A1(_u10_u7_n2669 ), .A2(_u10_u7_n3125 ), .ZN(_u10_u7_n3124 ) );
NAND4_X1 _u10_u7_U958  ( .A1(_u10_u7_n3122 ), .A2(_u10_u7_n3123 ), .A3(_u10_u7_n3124 ), .A4(_u10_u7_n2579 ), .ZN(_u10_u7_n3121 ) );
NAND2_X1 _u10_u7_U957  ( .A1(_u10_u7_n3121 ), .A2(_u10_u7_n2874 ), .ZN(_u10_u7_n3120 ) );
NAND2_X1 _u10_u7_U956  ( .A1(_u10_u7_n2382 ), .A2(_u10_u7_n3120 ), .ZN(_u10_u7_n3119 ) );
NAND2_X1 _u10_u7_U955  ( .A1(_u10_u7_n1967 ), .A2(_u10_u7_n3119 ), .ZN(_u10_u7_n3099 ) );
NAND2_X1 _u10_u7_U954  ( .A1(_u10_u7_n3118 ), .A2(_u10_u7_n3001 ), .ZN(_u10_u7_n3117 ) );
NAND2_X1 _u10_u7_U953  ( .A1(_u10_u7_n2446 ), .A2(_u10_u7_n3117 ), .ZN(_u10_u7_n3116 ) );
NAND2_X1 _u10_u7_U952  ( .A1(_u10_u7_n2445 ), .A2(_u10_u7_n3116 ), .ZN(_u10_u7_n3100 ) );
OR2_X1 _u10_u7_U951  ( .A1(_u10_u7_n3115 ), .A2(_u10_u7_n2687 ), .ZN(_u10_u7_n3114 ) );
AND3_X1 _u10_u7_U950  ( .A1(_u10_u7_n2061 ), .A2(_u10_u7_n2166 ), .A3(_u10_u7_n3114 ), .ZN(_u10_u7_n3045 ) );
NOR2_X1 _u10_u7_U949  ( .A1(1'b0), .A2(_u10_u7_n3045 ), .ZN(_u10_u7_n3113 ));
NOR2_X1 _u10_u7_U948  ( .A1(_u10_u7_n3113 ), .A2(1'b0), .ZN(_u10_u7_n3112 ));
NOR2_X1 _u10_u7_U947  ( .A1(_u10_u7_n3112 ), .A2(_u10_u7_n2356 ), .ZN(_u10_u7_n3102 ) );
NAND2_X1 _u10_u7_U946  ( .A1(_u10_u7_n2571 ), .A2(_u10_u7_n2165 ), .ZN(_u10_u7_n3078 ) );
NAND2_X1 _u10_u7_U945  ( .A1(_u10_u7_n2365 ), .A2(_u10_u7_n3078 ), .ZN(_u10_u7_n2241 ) );
NOR2_X1 _u10_u7_U944  ( .A1(_u10_u7_n2377 ), .A2(_u10_u7_n2241 ), .ZN(_u10_u7_n3111 ) );
NOR2_X1 _u10_u7_U943  ( .A1(_u10_u7_n3111 ), .A2(_u10_u7_n1869 ), .ZN(_u10_u7_n3103 ) );
NOR2_X1 _u10_u7_U942  ( .A1(_u10_u7_n2999 ), .A2(_u10_u7_n2977 ), .ZN(_u10_u7_n3061 ) );
NOR2_X1 _u10_u7_U941  ( .A1(_u10_u7_n3061 ), .A2(_u10_u7_n2367 ), .ZN(_u10_u7_n3106 ) );
NAND2_X1 _u10_u7_U940  ( .A1(_u10_u7_n2977 ), .A2(_u10_u7_n3000 ), .ZN(_u10_u7_n3110 ) );
NAND2_X1 _u10_u7_U939  ( .A1(_u10_u7_n3109 ), .A2(_u10_u7_n3110 ), .ZN(_u10_u7_n1924 ) );
AND2_X1 _u10_u7_U938  ( .A1(_u10_u7_n1924 ), .A2(_u10_u7_n3108 ), .ZN(_u10_u7_n3107 ) );
NOR2_X1 _u10_u7_U937  ( .A1(_u10_u7_n3106 ), .A2(_u10_u7_n3107 ), .ZN(_u10_u7_n3105 ) );
NOR2_X1 _u10_u7_U936  ( .A1(_u10_u7_n3105 ), .A2(_u10_u7_n2008 ), .ZN(_u10_u7_n3104 ) );
NOR3_X1 _u10_u7_U935  ( .A1(_u10_u7_n3102 ), .A2(_u10_u7_n3103 ), .A3(_u10_u7_n3104 ), .ZN(_u10_u7_n3101 ) );
NAND4_X1 _u10_u7_U934  ( .A1(_u10_u7_n3098 ), .A2(_u10_u7_n3099 ), .A3(_u10_u7_n3100 ), .A4(_u10_u7_n3101 ), .ZN(_u10_u7_n3071 ) );
NOR2_X1 _u10_u7_U933  ( .A1(_u10_u7_n1926 ), .A2(_u10_u7_n2980 ), .ZN(_u10_u7_n2218 ) );
INV_X1 _u10_u7_U932  ( .A(_u10_u7_n2721 ), .ZN(_u10_u7_n2910 ) );
NAND2_X1 _u10_u7_U931  ( .A1(_u10_u7_n2910 ), .A2(_u10_u7_n1869 ), .ZN(_u10_u7_n2779 ) );
NAND2_X1 _u10_u7_U930  ( .A1(_u10_u7_n2218 ), .A2(_u10_u7_n2779 ), .ZN(_u10_u7_n3081 ) );
NAND2_X1 _u10_u7_U929  ( .A1(_u10_u7_n1922 ), .A2(_u10_u7_n1864 ), .ZN(_u10_u7_n2179 ) );
NOR3_X1 _u10_u7_U928  ( .A1(_u10_u7_n1961 ), .A2(_u10_u7_n1918 ), .A3(_u10_u7_n2179 ), .ZN(_u10_u7_n2693 ) );
NAND2_X1 _u10_u7_U927  ( .A1(_u10_u7_n3097 ), .A2(_u10_u7_n1924 ), .ZN(_u10_u7_n3096 ) );
NAND2_X1 _u10_u7_U926  ( .A1(_u10_u7_n1984 ), .A2(_u10_u7_n3096 ), .ZN(_u10_u7_n2506 ) );
INV_X1 _u10_u7_U925  ( .A(_u10_u7_n2506 ), .ZN(_u10_u7_n2366 ) );
NAND2_X1 _u10_u7_U924  ( .A1(_u10_u7_n2366 ), .A2(_u10_u7_n2375 ), .ZN(_u10_u7_n2236 ) );
NAND2_X1 _u10_u7_U923  ( .A1(_u10_u7_n2693 ), .A2(_u10_u7_n2236 ), .ZN(_u10_u7_n3082 ) );
NAND2_X1 _u10_u7_U922  ( .A1(1'b0), .A2(_u10_u7_n2126 ), .ZN(_u10_u7_n3095 ));
NAND2_X1 _u10_u7_U921  ( .A1(_u10_u7_n1956 ), .A2(_u10_u7_n3095 ), .ZN(_u10_u7_n2907 ) );
OR2_X1 _u10_u7_U920  ( .A1(_u10_u7_n2902 ), .A2(_u10_u7_n2907 ), .ZN(_u10_u7_n3085 ) );
NAND2_X1 _u10_u7_U919  ( .A1(_u10_u7_n2256 ), .A2(_u10_u7_n2113 ), .ZN(_u10_u7_n3094 ) );
NAND2_X1 _u10_u7_U918  ( .A1(_u10_u7_n2688 ), .A2(_u10_u7_n3094 ), .ZN(_u10_u7_n3092 ) );
NAND2_X1 _u10_u7_U917  ( .A1(_u10_u7_n3093 ), .A2(_u10_u7_n3092 ), .ZN(_u10_u7_n3086 ) );
INV_X1 _u10_u7_U916  ( .A(_u10_u7_n2159 ), .ZN(_u10_u7_n1894 ) );
NAND2_X1 _u10_u7_U915  ( .A1(_u10_u7_n3067 ), .A2(_u10_u7_n1894 ), .ZN(_u10_u7_n3091 ) );
INV_X1 _u10_u7_U914  ( .A(_u10_u7_n3092 ), .ZN(_u10_u7_n2234 ) );
NAND3_X1 _u10_u7_U913  ( .A1(_u10_u7_n3091 ), .A2(_u10_u7_n2126 ), .A3(_u10_u7_n2234 ), .ZN(_u10_u7_n3090 ) );
NAND2_X1 _u10_u7_U912  ( .A1(1'b0), .A2(_u10_u7_n3090 ), .ZN(_u10_u7_n3087 ));
NAND3_X1 _u10_u7_U911  ( .A1(_u10_u7_n2329 ), .A2(_u10_u7_n3089 ), .A3(_u10_u7_n2549 ), .ZN(_u10_u7_n3088 ) );
NAND4_X1 _u10_u7_U910  ( .A1(_u10_u7_n3085 ), .A2(_u10_u7_n3086 ), .A3(_u10_u7_n3087 ), .A4(_u10_u7_n3088 ), .ZN(_u10_u7_n3084 ) );
NAND2_X1 _u10_u7_U909  ( .A1(_u10_u7_n3084 ), .A2(_u10_u7_n2803 ), .ZN(_u10_u7_n3083 ) );
NAND3_X1 _u10_u7_U908  ( .A1(_u10_u7_n3081 ), .A2(_u10_u7_n3082 ), .A3(_u10_u7_n3083 ), .ZN(_u10_u7_n3072 ) );
INV_X1 _u10_u7_U907  ( .A(_u10_u7_n2689 ), .ZN(_u10_u7_n1955 ) );
NOR3_X1 _u10_u7_U906  ( .A1(_u10_u7_n1955 ), .A2(_u10_u7_n2813 ), .A3(_u10_u7_n2488 ), .ZN(_u10_u7_n3080 ) );
NOR2_X1 _u10_u7_U905  ( .A1(_u10_u7_n3080 ), .A2(_u10_u7_n2485 ), .ZN(_u10_u7_n3073 ) );
NAND3_X1 _u10_u7_U904  ( .A1(_u10_u7_n2621 ), .A2(_u10_u7_n2202 ), .A3(_u10_u7_n3079 ), .ZN(_u10_u7_n2110 ) );
NOR2_X1 _u10_u7_U903  ( .A1(_u10_u7_n2110 ), .A2(_u10_u7_n2218 ), .ZN(_u10_u7_n2775 ) );
INV_X1 _u10_u7_U902  ( .A(_u10_u7_n2775 ), .ZN(_u10_u7_n3024 ) );
INV_X1 _u10_u7_U901  ( .A(_u10_u7_n3078 ), .ZN(_u10_u7_n2133 ) );
INV_X1 _u10_u7_U900  ( .A(_u10_u7_n2007 ), .ZN(_u10_u7_n2358 ) );
NAND2_X1 _u10_u7_U899  ( .A1(_u10_u7_n2358 ), .A2(_u10_u7_n2886 ), .ZN(_u10_u7_n2240 ) );
INV_X1 _u10_u7_U898  ( .A(_u10_u7_n2240 ), .ZN(_u10_u7_n2083 ) );
NOR3_X1 _u10_u7_U897  ( .A1(_u10_u7_n2952 ), .A2(_u10_u7_n2004 ), .A3(_u10_u7_n1891 ), .ZN(_u10_u7_n3077 ) );
NAND3_X1 _u10_u7_U896  ( .A1(_u10_u7_n2083 ), .A2(_u10_u7_n2938 ), .A3(_u10_u7_n3077 ), .ZN(_u10_u7_n1886 ) );
NOR3_X1 _u10_u7_U895  ( .A1(_u10_u7_n3024 ), .A2(_u10_u7_n2133 ), .A3(_u10_u7_n1886 ), .ZN(_u10_u7_n3075 ) );
NOR2_X1 _u10_u7_U894  ( .A1(_u10_u7_n3075 ), .A2(_u10_u7_n3076 ), .ZN(_u10_u7_n3074 ) );
NOR4_X1 _u10_u7_U893  ( .A1(_u10_u7_n3071 ), .A2(_u10_u7_n3072 ), .A3(_u10_u7_n3073 ), .A4(_u10_u7_n3074 ), .ZN(_u10_u7_n3017 ) );
INV_X1 _u10_u7_U892  ( .A(_u10_u7_n3065 ), .ZN(_u10_u7_n3043 ) );
NAND2_X1 _u10_u7_U891  ( .A1(_u10_u7_n3043 ), .A2(_u10_u7_n2106 ), .ZN(_u10_u7_n3070 ) );
NAND2_X1 _u10_u7_U890  ( .A1(_u10_u7_n3070 ), .A2(_u10_u7_n2038 ), .ZN(_u10_u7_n3068 ) );
NAND2_X1 _u10_u7_U889  ( .A1(_u10_u7_n2344 ), .A2(_u10_u7_n2584 ), .ZN(_u10_u7_n3069 ) );
NAND3_X1 _u10_u7_U888  ( .A1(_u10_u7_n3068 ), .A2(_u10_u7_n1930 ), .A3(_u10_u7_n3069 ), .ZN(_u10_u7_n3047 ) );
NAND2_X1 _u10_u7_U887  ( .A1(_u10_u7_n2835 ), .A2(_u10_u7_n2466 ), .ZN(_u10_u7_n2130 ) );
INV_X1 _u10_u7_U886  ( .A(_u10_u7_n2130 ), .ZN(_u10_u7_n2168 ) );
NAND3_X1 _u10_u7_U885  ( .A1(_u10_u7_n3067 ), .A2(_u10_u7_n2329 ), .A3(_u10_u7_n2168 ), .ZN(_u10_u7_n2665 ) );
NAND3_X1 _u10_u7_U884  ( .A1(_u10_u7_n3065 ), .A2(_u10_u7_n3066 ), .A3(_u10_u7_n2342 ), .ZN(_u10_u7_n3064 ) );
NAND3_X1 _u10_u7_U883  ( .A1(_u10_u7_n3064 ), .A2(_u10_u7_n2175 ), .A3(_u10_u7_n2987 ), .ZN(_u10_u7_n3048 ) );
NOR3_X1 _u10_u7_U882  ( .A1(_u10_u7_n1849 ), .A2(1'b0), .A3(_u10_u7_n3063 ),.ZN(_u10_u7_n3050 ) );
NOR3_X1 _u10_u7_U881  ( .A1(_u10_u7_n2406 ), .A2(1'b0), .A3(_u10_u7_n3062 ),.ZN(_u10_u7_n3060 ) );
NOR3_X1 _u10_u7_U880  ( .A1(_u10_u7_n3060 ), .A2(1'b0), .A3(_u10_u7_n3061 ),.ZN(_u10_u7_n3051 ) );
NAND2_X1 _u10_u7_U879  ( .A1(_u10_u7_n3059 ), .A2(_u10_u7_n2049 ), .ZN(_u10_u7_n3056 ) );
NAND3_X1 _u10_u7_U878  ( .A1(_u10_u7_n3056 ), .A2(_u10_u7_n3057 ), .A3(_u10_u7_n3058 ), .ZN(_u10_u7_n3054 ) );
NOR4_X1 _u10_u7_U877  ( .A1(_u10_u7_n3054 ), .A2(_u10_u7_n3055 ), .A3(_u10_u7_n2055 ), .A4(_u10_u7_n2056 ), .ZN(_u10_u7_n3053 ) );
NOR3_X1 _u10_u7_U876  ( .A1(_u10_u7_n2346 ), .A2(1'b0), .A3(_u10_u7_n3053 ),.ZN(_u10_u7_n3052 ) );
NOR3_X1 _u10_u7_U875  ( .A1(_u10_u7_n3050 ), .A2(_u10_u7_n3051 ), .A3(_u10_u7_n3052 ), .ZN(_u10_u7_n3049 ) );
NAND4_X1 _u10_u7_U874  ( .A1(_u10_u7_n3047 ), .A2(_u10_u7_n2665 ), .A3(_u10_u7_n3048 ), .A4(_u10_u7_n3049 ), .ZN(_u10_u7_n3019 ) );
NAND2_X1 _u10_u7_U873  ( .A1(_u10_u7_n2056 ), .A2(_u10_u7_n2019 ), .ZN(_u10_u7_n3046 ) );
NAND2_X1 _u10_u7_U872  ( .A1(_u10_u7_n3045 ), .A2(_u10_u7_n3046 ), .ZN(_u10_u7_n3044 ) );
NAND2_X1 _u10_u7_U871  ( .A1(_u10_u7_n3044 ), .A2(_u10_u7_n2165 ), .ZN(_u10_u7_n3028 ) );
OR2_X1 _u10_u7_U870  ( .A1(_u10_u7_n2179 ), .A2(_u10_u7_n1961 ), .ZN(_u10_u7_n3037 ) );
NAND2_X1 _u10_u7_U869  ( .A1(_u10_u7_n3043 ), .A2(_u10_u7_n2336 ), .ZN(_u10_u7_n3042 ) );
NAND2_X1 _u10_u7_U868  ( .A1(_u10_u7_n3042 ), .A2(_u10_u7_n3006 ), .ZN(_u10_u7_n3041 ) );
NAND2_X1 _u10_u7_U867  ( .A1(_u10_u7_n3040 ), .A2(_u10_u7_n3041 ), .ZN(_u10_u7_n3026 ) );
NAND4_X1 _u10_u7_U866  ( .A1(_u10_u7_n3026 ), .A2(_u10_u7_n2520 ), .A3(_u10_u7_n1962 ), .A4(_u10_u7_n1864 ), .ZN(_u10_u7_n3039 ) );
NAND2_X1 _u10_u7_U865  ( .A1(_u10_u7_n3039 ), .A2(_u10_u7_n1922 ), .ZN(_u10_u7_n3038 ) );
NAND2_X1 _u10_u7_U864  ( .A1(_u10_u7_n3037 ), .A2(_u10_u7_n3038 ), .ZN(_u10_u7_n3035 ) );
NAND2_X1 _u10_u7_U863  ( .A1(_u10_u7_n2985 ), .A2(_u10_u7_n3036 ), .ZN(_u10_u7_n2432 ) );
NAND2_X1 _u10_u7_U862  ( .A1(_u10_u7_n3035 ), .A2(_u10_u7_n2432 ), .ZN(_u10_u7_n3029 ) );
INV_X1 _u10_u7_U861  ( .A(_u10_u7_n3034 ), .ZN(_u10_u7_n2777 ) );
INV_X1 _u10_u7_U860  ( .A(_u10_u7_n2772 ), .ZN(_u10_u7_n3032 ) );
NAND2_X1 _u10_u7_U859  ( .A1(_u10_u7_n1982 ), .A2(_u10_u7_n2978 ), .ZN(_u10_u7_n3033 ) );
NAND2_X1 _u10_u7_U858  ( .A1(_u10_u7_n3032 ), .A2(_u10_u7_n3033 ), .ZN(_u10_u7_n3031 ) );
NAND2_X1 _u10_u7_U857  ( .A1(_u10_u7_n2777 ), .A2(_u10_u7_n3031 ), .ZN(_u10_u7_n3030 ) );
NAND3_X1 _u10_u7_U856  ( .A1(_u10_u7_n3028 ), .A2(_u10_u7_n3029 ), .A3(_u10_u7_n3030 ), .ZN(_u10_u7_n3020 ) );
NOR3_X1 _u10_u7_U855  ( .A1(_u10_u7_n2179 ), .A2(1'b0), .A3(_u10_u7_n2375 ),.ZN(_u10_u7_n3027 ) );
NOR2_X1 _u10_u7_U854  ( .A1(_u10_u7_n3027 ), .A2(_u10_u7_n2177 ), .ZN(_u10_u7_n3025 ) );
NOR2_X1 _u10_u7_U853  ( .A1(_u10_u7_n3025 ), .A2(_u10_u7_n3026 ), .ZN(_u10_u7_n3021 ) );
NOR2_X1 _u10_u7_U852  ( .A1(_u10_u7_n2256 ), .A2(_u10_u7_n3024 ), .ZN(_u10_u7_n3023 ) );
NOR2_X1 _u10_u7_U851  ( .A1(_u10_u7_n3023 ), .A2(_u10_u7_n1868 ), .ZN(_u10_u7_n3022 ) );
NOR4_X1 _u10_u7_U850  ( .A1(_u10_u7_n3019 ), .A2(_u10_u7_n3020 ), .A3(_u10_u7_n3021 ), .A4(_u10_u7_n3022 ), .ZN(_u10_u7_n3018 ) );
NAND4_X1 _u10_u7_U849  ( .A1(_u10_u7_n3015 ), .A2(_u10_u7_n3016 ), .A3(_u10_u7_n3017 ), .A4(_u10_u7_n3018 ), .ZN(_u10_u7_n2958 ) );
NOR2_X1 _u10_u7_U848  ( .A1(1'b0), .A2(_u10_u7_n2573 ), .ZN(_u10_u7_n3011 ));
NOR2_X1 _u10_u7_U847  ( .A1(1'b0), .A2(_u10_u7_n2359 ), .ZN(_u10_u7_n3012 ));
NOR2_X1 _u10_u7_U846  ( .A1(1'b0), .A2(_u10_u7_n1859 ), .ZN(_u10_u7_n3013 ));
NOR2_X1 _u10_u7_U845  ( .A1(1'b0), .A2(_u10_u7_n1836 ), .ZN(_u10_u7_n3014 ));
NOR4_X1 _u10_u7_U844  ( .A1(_u10_u7_n3011 ), .A2(_u10_u7_n3012 ), .A3(_u10_u7_n3013 ), .A4(_u10_u7_n3014 ), .ZN(_u10_u7_n2959 ) );
NOR2_X1 _u10_u7_U843  ( .A1(1'b0), .A2(_u10_u7_n2025 ), .ZN(_u10_u7_n3007 ));
NOR2_X1 _u10_u7_U842  ( .A1(1'b0), .A2(_u10_u7_n2085 ), .ZN(_u10_u7_n3008 ));
NOR2_X1 _u10_u7_U841  ( .A1(1'b0), .A2(_u10_u7_n2607 ), .ZN(_u10_u7_n3009 ));
NOR2_X1 _u10_u7_U840  ( .A1(1'b0), .A2(_u10_u7_n2071 ), .ZN(_u10_u7_n3010 ));
NOR4_X1 _u10_u7_U839  ( .A1(_u10_u7_n3007 ), .A2(_u10_u7_n3008 ), .A3(_u10_u7_n3009 ), .A4(_u10_u7_n3010 ), .ZN(_u10_u7_n2960 ) );
NAND2_X1 _u10_u7_U838  ( .A1(_u10_u7_n1894 ), .A2(_u10_u7_n2466 ), .ZN(_u10_u7_n3002 ) );
NAND2_X1 _u10_u7_U837  ( .A1(_u10_u7_n2830 ), .A2(_u10_u7_n2600 ), .ZN(_u10_u7_n3003 ) );
NAND2_X1 _u10_u7_U836  ( .A1(_u10_u7_n1960 ), .A2(_u10_u7_n2431 ), .ZN(_u10_u7_n3004 ) );
NAND2_X1 _u10_u7_U835  ( .A1(_u10_u7_n2002 ), .A2(_u10_u7_n3006 ), .ZN(_u10_u7_n3005 ) );
NAND4_X1 _u10_u7_U834  ( .A1(_u10_u7_n3002 ), .A2(_u10_u7_n3003 ), .A3(_u10_u7_n3004 ), .A4(_u10_u7_n3005 ), .ZN(_u10_u7_n2992 ) );
NAND2_X1 _u10_u7_U833  ( .A1(_u10_u7_n2461 ), .A2(_u10_u7_n3001 ), .ZN(_u10_u7_n2997 ) );
NAND2_X1 _u10_u7_U832  ( .A1(_u10_u7_n2999 ), .A2(_u10_u7_n3000 ), .ZN(_u10_u7_n2998 ) );
NAND2_X1 _u10_u7_U831  ( .A1(_u10_u7_n2997 ), .A2(_u10_u7_n2998 ), .ZN(_u10_u7_n2993 ) );
NOR2_X1 _u10_u7_U830  ( .A1(_u10_SYNOPSYS_UNCONNECTED_29 ), .A2(_u10_u7_n2996 ), .ZN(_u10_u7_n2995 ) );
NOR2_X1 _u10_u7_U829  ( .A1(_u10_u7_n2995 ), .A2(_u10_u7_n2126 ), .ZN(_u10_u7_n2994 ) );
NOR4_X1 _u10_u7_U828  ( .A1(_u10_u7_n2992 ), .A2(_u10_u7_n2993 ), .A3(next_ch), .A4(_u10_u7_n2994 ), .ZN(_u10_u7_n2961 ) );
NAND2_X1 _u10_u7_U827  ( .A1(_u10_u7_n2445 ), .A2(_u10_u7_n2803 ), .ZN(_u10_u7_n2988 ) );
OR2_X1 _u10_u7_U826  ( .A1(_u10_u7_n2584 ), .A2(1'b0), .ZN(_u10_u7_n2989 ));
NAND2_X1 _u10_u7_U825  ( .A1(_u10_u7_n2709 ), .A2(_u10_u7_n2080 ), .ZN(_u10_u7_n2990 ) );
NAND2_X1 _u10_u7_U824  ( .A1(_u10_u7_n2183 ), .A2(_u10_u7_n2166 ), .ZN(_u10_u7_n2991 ) );
NAND4_X1 _u10_u7_U823  ( .A1(_u10_u7_n2988 ), .A2(_u10_u7_n2989 ), .A3(_u10_u7_n2990 ), .A4(_u10_u7_n2991 ), .ZN(_u10_u7_n2963 ) );
NAND2_X1 _u10_u7_U822  ( .A1(_u10_u7_n2987 ), .A2(_u10_u7_n1930 ), .ZN(_u10_u7_n2981 ) );
NAND2_X1 _u10_u7_U821  ( .A1(_u10_u7_n2986 ), .A2(_u10_u7_n2038 ), .ZN(_u10_u7_n2982 ) );
OR2_X1 _u10_u7_U820  ( .A1(_u10_u7_n2985 ), .A2(1'b0), .ZN(_u10_u7_n2983 ));
NAND2_X1 _u10_u7_U819  ( .A1(_u10_u7_n2169 ), .A2(_u10_u7_n2113 ), .ZN(_u10_u7_n2984 ) );
NAND4_X1 _u10_u7_U818  ( .A1(_u10_u7_n2981 ), .A2(_u10_u7_n2982 ), .A3(_u10_u7_n2983 ), .A4(_u10_u7_n2984 ), .ZN(_u10_u7_n2964 ) );
NAND2_X1 _u10_u7_U817  ( .A1(_u10_u7_n2509 ), .A2(_u10_u7_n1864 ), .ZN(_u10_u7_n2973 ) );
INV_X1 _u10_u7_U816  ( .A(_u10_u7_n2980 ), .ZN(_u10_u7_n1861 ) );
NAND2_X1 _u10_u7_U815  ( .A1(_u10_u7_n1861 ), .A2(_u10_u7_n1922 ), .ZN(_u10_u7_n2974 ) );
NAND2_X1 _u10_u7_U814  ( .A1(_u10_u7_n2979 ), .A2(_u10_u7_n2405 ), .ZN(_u10_u7_n2975 ) );
NAND2_X1 _u10_u7_U813  ( .A1(_u10_u7_n2977 ), .A2(_u10_u7_n2978 ), .ZN(_u10_u7_n2976 ) );
NAND4_X1 _u10_u7_U812  ( .A1(_u10_u7_n2973 ), .A2(_u10_u7_n2974 ), .A3(_u10_u7_n2975 ), .A4(_u10_u7_n2976 ), .ZN(_u10_u7_n2965 ) );
NAND2_X1 _u10_u7_U811  ( .A1(_u10_u7_n2507 ), .A2(_u10_u7_n2972 ), .ZN(_u10_u7_n2967 ) );
NAND2_X1 _u10_u7_U810  ( .A1(_u10_u7_n2043 ), .A2(_u10_u7_n1965 ), .ZN(_u10_u7_n2968 ) );
NAND2_X1 _u10_u7_U809  ( .A1(_u10_u7_n2063 ), .A2(_u10_u7_n1853 ), .ZN(_u10_u7_n2969 ) );
NAND2_X1 _u10_u7_U808  ( .A1(_u10_u7_n2971 ), .A2(_u10_u7_n2175 ), .ZN(_u10_u7_n2970 ) );
NAND4_X1 _u10_u7_U807  ( .A1(_u10_u7_n2967 ), .A2(_u10_u7_n2968 ), .A3(_u10_u7_n2969 ), .A4(_u10_u7_n2970 ), .ZN(_u10_u7_n2966 ) );
NOR4_X1 _u10_u7_U806  ( .A1(_u10_u7_n2963 ), .A2(_u10_u7_n2964 ), .A3(_u10_u7_n2965 ), .A4(_u10_u7_n2966 ), .ZN(_u10_u7_n2962 ) );
AND4_X1 _u10_u7_U805  ( .A1(_u10_u7_n2959 ), .A2(_u10_u7_n2960 ), .A3(_u10_u7_n2961 ), .A4(_u10_u7_n2962 ), .ZN(_u10_u7_n1819 ) );
MUX2_X1 _u10_u7_U804  ( .A(_u10_u7_n2958 ), .B(_u10_SYNOPSYS_UNCONNECTED_33 ), .S(_u10_u7_n1819 ), .Z(_u10_u7_n1808 ) );
NOR2_X1 _u10_u7_U803  ( .A1(_u10_u7_n2531 ), .A2(_u10_u7_n2607 ), .ZN(_u10_u7_n1911 ) );
NAND2_X1 _u10_u7_U802  ( .A1(_u10_u7_n1911 ), .A2(_u10_u7_n2957 ), .ZN(_u10_u7_n2954 ) );
NAND2_X1 _u10_u7_U801  ( .A1(_u10_u7_n1853 ), .A2(_u10_u7_n1965 ), .ZN(_u10_u7_n2956 ) );
NAND2_X1 _u10_u7_U800  ( .A1(_u10_u7_n1966 ), .A2(_u10_u7_n2956 ), .ZN(_u10_u7_n2955 ) );
NAND2_X1 _u10_u7_U799  ( .A1(_u10_u7_n2954 ), .A2(_u10_u7_n2955 ), .ZN(_u10_u7_n2670 ) );
NOR3_X1 _u10_u7_U798  ( .A1(_u10_u7_n1852 ), .A2(1'b0), .A3(_u10_u7_n1853 ),.ZN(_u10_u7_n2708 ) );
NAND2_X1 _u10_u7_U797  ( .A1(_u10_u7_n2708 ), .A2(_u10_u7_n2080 ), .ZN(_u10_u7_n2355 ) );
NOR2_X1 _u10_u7_U796  ( .A1(_u10_u7_n2355 ), .A2(1'b0), .ZN(_u10_u7_n2599 ));
NAND2_X1 _u10_u7_U795  ( .A1(_u10_u7_n2953 ), .A2(_u10_u7_n2599 ), .ZN(_u10_u7_n2423 ) );
OR2_X1 _u10_u7_U794  ( .A1(_u10_u7_n2423 ), .A2(_u10_u7_n2359 ), .ZN(_u10_u7_n2949 ) );
NAND3_X1 _u10_u7_U793  ( .A1(_u10_u7_n2105 ), .A2(_u10_u7_n1936 ), .A3(_u10_u7_n2952 ), .ZN(_u10_u7_n2950 ) );
NAND3_X1 _u10_u7_U792  ( .A1(_u10_u7_n2549 ), .A2(_u10_u7_n1936 ), .A3(1'b0),.ZN(_u10_u7_n2096 ) );
INV_X1 _u10_u7_U791  ( .A(_u10_u7_n2096 ), .ZN(_u10_u7_n2301 ) );
NAND2_X1 _u10_u7_U790  ( .A1(_u10_u7_n2301 ), .A2(_u10_u7_n2446 ), .ZN(_u10_u7_n2368 ) );
INV_X1 _u10_u7_U789  ( .A(_u10_u7_n2368 ), .ZN(_u10_u7_n2326 ) );
NAND2_X1 _u10_u7_U788  ( .A1(_u10_u7_n2326 ), .A2(_u10_u7_n2941 ), .ZN(_u10_u7_n2800 ) );
INV_X1 _u10_u7_U787  ( .A(_u10_u7_n2800 ), .ZN(_u10_u7_n2081 ) );
NAND2_X1 _u10_u7_U786  ( .A1(_u10_u7_n2081 ), .A2(_u10_u7_n2049 ), .ZN(_u10_u7_n2855 ) );
INV_X1 _u10_u7_U785  ( .A(_u10_u7_n2855 ), .ZN(_u10_u7_n2347 ) );
NAND2_X1 _u10_u7_U784  ( .A1(_u10_u7_n2347 ), .A2(_u10_u7_n2063 ), .ZN(_u10_u7_n2951 ) );
NAND3_X1 _u10_u7_U783  ( .A1(_u10_u7_n2949 ), .A2(_u10_u7_n2950 ), .A3(_u10_u7_n2951 ), .ZN(_u10_u7_n1997 ) );
INV_X1 _u10_u7_U782  ( .A(_u10_u7_n1997 ), .ZN(_u10_u7_n2917 ) );
AND2_X1 _u10_u7_U781  ( .A1(_u10_u7_n2709 ), .A2(_u10_u7_n2708 ), .ZN(_u10_u7_n2942 ) );
INV_X1 _u10_u7_U780  ( .A(_u10_u7_n2907 ), .ZN(_u10_u7_n2737 ) );
NAND2_X1 _u10_u7_U779  ( .A1(_u10_u7_n2737 ), .A2(_u10_u7_n2803 ), .ZN(_u10_u7_n1888 ) );
NOR2_X1 _u10_u7_U778  ( .A1(_u10_u7_n2001 ), .A2(_u10_u7_n1888 ), .ZN(_u10_u7_n2943 ) );
NAND4_X1 _u10_u7_U777  ( .A1(1'b0), .A2(_u10_u7_n2078 ), .A3(_u10_u7_n2059 ),.A4(_u10_u7_n2031 ), .ZN(_u10_u7_n2578 ) );
NOR3_X1 _u10_u7_U776  ( .A1(_u10_u7_n2719 ), .A2(_u10_u7_n2130 ), .A3(_u10_u7_n2305 ), .ZN(_u10_u7_n2386 ) );
NAND2_X1 _u10_u7_U775  ( .A1(_u10_u7_n2386 ), .A2(_u10_u7_n2669 ), .ZN(_u10_u7_n2948 ) );
NAND3_X1 _u10_u7_U774  ( .A1(_u10_u7_n2578 ), .A2(_u10_u7_n2947 ), .A3(_u10_u7_n2948 ), .ZN(_u10_u7_n2750 ) );
NOR2_X1 _u10_u7_U773  ( .A1(_u10_u7_n2274 ), .A2(_u10_u7_n2852 ), .ZN(_u10_u7_n2946 ) );
NOR3_X1 _u10_u7_U772  ( .A1(_u10_u7_n2750 ), .A2(1'b0), .A3(_u10_u7_n2946 ),.ZN(_u10_u7_n2945 ) );
NOR2_X1 _u10_u7_U771  ( .A1(_u10_u7_n2945 ), .A2(_u10_u7_n2359 ), .ZN(_u10_u7_n2944 ) );
NOR3_X1 _u10_u7_U770  ( .A1(_u10_u7_n2942 ), .A2(_u10_u7_n2943 ), .A3(_u10_u7_n2944 ), .ZN(_u10_u7_n2919 ) );
NOR2_X1 _u10_u7_U769  ( .A1(_u10_u7_n2423 ), .A2(1'b0), .ZN(_u10_u7_n1979 ));
NAND3_X1 _u10_u7_U768  ( .A1(_u10_u7_n2549 ), .A2(_u10_u7_n1936 ), .A3(_u10_u7_n1979 ), .ZN(_u10_u7_n2328 ) );
INV_X1 _u10_u7_U767  ( .A(_u10_u7_n2328 ), .ZN(_u10_u7_n2554 ) );
NAND3_X1 _u10_u7_U766  ( .A1(_u10_u7_n2941 ), .A2(_u10_u7_n2446 ), .A3(_u10_u7_n2554 ), .ZN(_u10_u7_n2115 ) );
NOR2_X1 _u10_u7_U765  ( .A1(_u10_u7_n2578 ), .A2(_u10_u7_n2030 ), .ZN(_u10_u7_n2553 ) );
INV_X1 _u10_u7_U764  ( .A(_u10_u7_n2553 ), .ZN(_u10_u7_n2269 ) );
NOR2_X1 _u10_u7_U763  ( .A1(_u10_u7_n2269 ), .A2(_u10_u7_n2790 ), .ZN(_u10_u7_n2657 ) );
INV_X1 _u10_u7_U762  ( .A(_u10_u7_n2657 ), .ZN(_u10_u7_n2210 ) );
NOR2_X1 _u10_u7_U761  ( .A1(_u10_u7_n2210 ), .A2(_u10_u7_n2911 ), .ZN(_u10_u7_n2213 ) );
INV_X1 _u10_u7_U760  ( .A(_u10_u7_n2213 ), .ZN(_u10_u7_n2456 ) );
NAND2_X1 _u10_u7_U759  ( .A1(_u10_u7_n2115 ), .A2(_u10_u7_n2456 ), .ZN(_u10_u7_n2634 ) );
INV_X1 _u10_u7_U758  ( .A(_u10_u7_n2634 ), .ZN(_u10_u7_n2220 ) );
NOR2_X1 _u10_u7_U757  ( .A1(_u10_u7_n2081 ), .A2(_u10_u7_n2386 ), .ZN(_u10_u7_n2131 ) );
NAND2_X1 _u10_u7_U756  ( .A1(_u10_u7_n2940 ), .A2(_u10_u7_n2131 ), .ZN(_u10_u7_n2138 ) );
INV_X1 _u10_u7_U755  ( .A(_u10_u7_n2138 ), .ZN(_u10_u7_n2927 ) );
NAND2_X1 _u10_u7_U754  ( .A1(_u10_u7_n2220 ), .A2(_u10_u7_n2927 ), .ZN(_u10_u7_n2939 ) );
NAND2_X1 _u10_u7_U753  ( .A1(_u10_u7_n1885 ), .A2(_u10_u7_n2939 ), .ZN(_u10_u7_n2931 ) );
NAND3_X1 _u10_u7_U752  ( .A1(_u10_u7_n1859 ), .A2(_u10_u7_n2365 ), .A3(_u10_u7_n2938 ), .ZN(_u10_u7_n2935 ) );
NAND3_X1 _u10_u7_U751  ( .A1(_u10_u7_n2927 ), .A2(_u10_u7_n2937 ), .A3(_u10_u7_n2220 ), .ZN(_u10_u7_n2936 ) );
NAND2_X1 _u10_u7_U750  ( .A1(_u10_u7_n2935 ), .A2(_u10_u7_n2936 ), .ZN(_u10_u7_n2932 ) );
INV_X1 _u10_u7_U749  ( .A(_u10_u7_n1937 ), .ZN(_u10_u7_n2350 ) );
NAND2_X1 _u10_u7_U748  ( .A1(_u10_u7_n1913 ), .A2(_u10_u7_n2350 ), .ZN(_u10_u7_n2934 ) );
NAND2_X1 _u10_u7_U747  ( .A1(_u10_u7_n2386 ), .A2(_u10_u7_n2934 ), .ZN(_u10_u7_n2933 ) );
NAND3_X1 _u10_u7_U746  ( .A1(_u10_u7_n2931 ), .A2(_u10_u7_n2932 ), .A3(_u10_u7_n2933 ), .ZN(_u10_u7_n2921 ) );
OR2_X1 _u10_u7_U745  ( .A1(_u10_u7_n2213 ), .A2(_u10_u7_n2386 ), .ZN(_u10_u7_n2930 ) );
NAND2_X1 _u10_u7_U744  ( .A1(_u10_u7_n2049 ), .A2(_u10_u7_n2930 ), .ZN(_u10_u7_n2228 ) );
AND2_X1 _u10_u7_U743  ( .A1(_u10_u7_n2228 ), .A2(_u10_u7_n2699 ), .ZN(_u10_u7_n2929 ) );
NOR2_X1 _u10_u7_U742  ( .A1(_u10_u7_n2929 ), .A2(_u10_u7_n2495 ), .ZN(_u10_u7_n2922 ) );
NOR2_X1 _u10_u7_U741  ( .A1(_u10_u7_n2633 ), .A2(_u10_u7_n2877 ), .ZN(_u10_u7_n2928 ) );
NOR2_X1 _u10_u7_U740  ( .A1(_u10_u7_n2928 ), .A2(_u10_u7_n2886 ), .ZN(_u10_u7_n2923 ) );
NOR2_X1 _u10_u7_U739  ( .A1(_u10_u7_n2927 ), .A2(_u10_u7_n2531 ), .ZN(_u10_u7_n2926 ) );
NOR2_X1 _u10_u7_U738  ( .A1(_u10_u7_n2926 ), .A2(_u10_u7_n2687 ), .ZN(_u10_u7_n2925 ) );
NOR2_X1 _u10_u7_U737  ( .A1(_u10_u7_n2925 ), .A2(_u10_u7_n1849 ), .ZN(_u10_u7_n2924 ) );
NOR4_X1 _u10_u7_U736  ( .A1(_u10_u7_n2921 ), .A2(_u10_u7_n2922 ), .A3(_u10_u7_n2923 ), .A4(_u10_u7_n2924 ), .ZN(_u10_u7_n2920 ) );
NAND4_X1 _u10_u7_U735  ( .A1(_u10_u7_n2917 ), .A2(_u10_u7_n2918 ), .A3(_u10_u7_n2919 ), .A4(_u10_u7_n2920 ), .ZN(_u10_u7_n2312 ) );
NOR2_X1 _u10_u7_U734  ( .A1(_u10_u7_n2600 ), .A2(_u10_u7_n2686 ), .ZN(_u10_u7_n2401 ) );
NAND2_X1 _u10_u7_U733  ( .A1(_u10_u7_n2401 ), .A2(_u10_u7_n2549 ), .ZN(_u10_u7_n2547 ) );
INV_X1 _u10_u7_U732  ( .A(_u10_u7_n2547 ), .ZN(_u10_u7_n2794 ) );
NAND3_X1 _u10_u7_U731  ( .A1(_u10_u7_n2364 ), .A2(_u10_u7_n2667 ), .A3(_u10_u7_n2794 ), .ZN(_u10_u7_n2535 ) );
INV_X1 _u10_u7_U730  ( .A(_u10_u7_n2535 ), .ZN(_u10_u7_n2586 ) );
NAND2_X1 _u10_u7_U729  ( .A1(_u10_u7_n2586 ), .A2(_u10_u7_n2571 ), .ZN(_u10_u7_n2916 ) );
NAND2_X1 _u10_u7_U728  ( .A1(_u10_u7_n2837 ), .A2(_u10_u7_n2916 ), .ZN(_u10_u7_n2436 ) );
NAND2_X1 _u10_u7_U727  ( .A1(_u10_u7_n2915 ), .A2(_u10_u7_n2571 ), .ZN(_u10_u7_n2914 ) );
NAND2_X1 _u10_u7_U726  ( .A1(_u10_u7_n2166 ), .A2(_u10_u7_n2914 ), .ZN(_u10_u7_n2017 ) );
NOR2_X1 _u10_u7_U725  ( .A1(_u10_u7_n2485 ), .A2(_u10_u7_n1841 ), .ZN(_u10_u7_n2913 ) );
OR4_X1 _u10_u7_U724  ( .A1(_u10_u7_n2436 ), .A2(_u10_u7_n2017 ), .A3(_u10_u7_n2913 ), .A4(_u10_u7_n2442 ), .ZN(_u10_u7_n2912 ) );
NAND2_X1 _u10_u7_U723  ( .A1(_u10_u7_n2709 ), .A2(_u10_u7_n2912 ), .ZN(_u10_u7_n2888 ) );
NAND3_X1 _u10_u7_U722  ( .A1(_u10_u7_n2078 ), .A2(_u10_u7_n2031 ), .A3(1'b0),.ZN(_u10_u7_n2580 ) );
INV_X1 _u10_u7_U721  ( .A(_u10_u7_n2580 ), .ZN(_u10_u7_n2680 ) );
AND2_X1 _u10_u7_U720  ( .A1(_u10_u7_n2680 ), .A2(_u10_u7_n2668 ), .ZN(_u10_u7_n1950 ) );
NAND2_X1 _u10_u7_U719  ( .A1(_u10_u7_n1950 ), .A2(_u10_u7_n2089 ), .ZN(_u10_u7_n2095 ) );
INV_X1 _u10_u7_U718  ( .A(_u10_u7_n2095 ), .ZN(_u10_u7_n2542 ) );
NAND2_X1 _u10_u7_U717  ( .A1(_u10_u7_n2542 ), .A2(_u10_u7_n2446 ), .ZN(_u10_u7_n1887 ) );
NOR2_X1 _u10_u7_U716  ( .A1(_u10_u7_n1887 ), .A2(_u10_u7_n2911 ), .ZN(_u10_u7_n2114 ) );
INV_X1 _u10_u7_U715  ( .A(_u10_u7_n2114 ), .ZN(_u10_u7_n1940 ) );
NAND3_X1 _u10_u7_U714  ( .A1(_u10_u7_n2535 ), .A2(_u10_u7_n1940 ), .A3(_u10_u7_n2910 ), .ZN(_u10_u7_n2524 ) );
NAND2_X1 _u10_u7_U713  ( .A1(_u10_u7_n2524 ), .A2(_u10_u7_n2488 ), .ZN(_u10_u7_n2889 ) );
NAND2_X1 _u10_u7_U712  ( .A1(_u10_u7_n2220 ), .A2(_u10_u7_n1940 ), .ZN(_u10_u7_n2763 ) );
NOR2_X1 _u10_u7_U711  ( .A1(_u10_u7_n2763 ), .A2(_u10_u7_n2586 ), .ZN(_u10_u7_n2808 ) );
NOR2_X1 _u10_u7_U710  ( .A1(_u10_u7_n2808 ), .A2(_u10_u7_n2350 ), .ZN(_u10_u7_n2908 ) );
NOR2_X1 _u10_u7_U709  ( .A1(_u10_u7_n2544 ), .A2(_u10_u7_n1950 ), .ZN(_u10_u7_n2899 ) );
NOR2_X1 _u10_u7_U708  ( .A1(_u10_u7_n2899 ), .A2(_u10_u7_n2159 ), .ZN(_u10_u7_n2909 ) );
NOR2_X1 _u10_u7_U707  ( .A1(_u10_u7_n2908 ), .A2(_u10_u7_n2909 ), .ZN(_u10_u7_n2890 ) );
NOR3_X1 _u10_u7_U706  ( .A1(_u10_u7_n2547 ), .A2(_u10_u7_n1846 ), .A3(_u10_u7_n2907 ), .ZN(_u10_u7_n2892 ) );
NOR3_X1 _u10_u7_U705  ( .A1(_u10_u7_n2240 ), .A2(_u10_u7_n2377 ), .A3(_u10_u7_n1911 ), .ZN(_u10_u7_n2906 ) );
NOR2_X1 _u10_u7_U704  ( .A1(_u10_u7_n2906 ), .A2(_u10_u7_n2535 ), .ZN(_u10_u7_n2893 ) );
NAND2_X1 _u10_u7_U703  ( .A1(_u10_u7_n2554 ), .A2(_u10_u7_n2446 ), .ZN(_u10_u7_n2903 ) );
AND3_X1 _u10_u7_U702  ( .A1(_u10_u7_n2210 ), .A2(_u10_u7_n2905 ), .A3(_u10_u7_n1887 ), .ZN(_u10_u7_n2904 ) );
NAND4_X1 _u10_u7_U701  ( .A1(_u10_u7_n2902 ), .A2(_u10_u7_n2498 ), .A3(_u10_u7_n2903 ), .A4(_u10_u7_n2904 ), .ZN(_u10_u7_n2788 ) );
INV_X1 _u10_u7_U700  ( .A(_u10_u7_n2788 ), .ZN(_u10_u7_n2901 ) );
NOR2_X1 _u10_u7_U699  ( .A1(_u10_u7_n2901 ), .A2(_u10_u7_n1888 ), .ZN(_u10_u7_n2894 ) );
NOR2_X1 _u10_u7_U698  ( .A1(_u10_u7_n2401 ), .A2(_u10_u7_n2553 ), .ZN(_u10_u7_n2900 ) );
NOR2_X1 _u10_u7_U697  ( .A1(_u10_u7_n2900 ), .A2(_u10_u7_n1954 ), .ZN(_u10_u7_n2897 ) );
NOR2_X1 _u10_u7_U696  ( .A1(1'b0), .A2(_u10_u7_n2899 ), .ZN(_u10_u7_n2898 ));
NOR2_X1 _u10_u7_U695  ( .A1(_u10_u7_n2897 ), .A2(_u10_u7_n2898 ), .ZN(_u10_u7_n2896 ) );
NOR2_X1 _u10_u7_U694  ( .A1(_u10_u7_n2896 ), .A2(_u10_u7_n1843 ), .ZN(_u10_u7_n2895 ) );
NOR4_X1 _u10_u7_U693  ( .A1(_u10_u7_n2892 ), .A2(_u10_u7_n2893 ), .A3(_u10_u7_n2894 ), .A4(_u10_u7_n2895 ), .ZN(_u10_u7_n2891 ) );
NAND4_X1 _u10_u7_U692  ( .A1(_u10_u7_n2888 ), .A2(_u10_u7_n2889 ), .A3(_u10_u7_n2890 ), .A4(_u10_u7_n2891 ), .ZN(_u10_u7_n2610 ) );
NOR4_X1 _u10_u7_U691  ( .A1(_u10_u7_n2670 ), .A2(_u10_u7_n2312 ), .A3(_u10_u7_n2610 ), .A4(_u10_u7_n2887 ), .ZN(_u10_u7_n2724 ) );
NOR2_X1 _u10_u7_U690  ( .A1(_u10_u7_n2883 ), .A2(_u10_u7_n2535 ), .ZN(_u10_u7_n2861 ) );
NOR2_X1 _u10_u7_U689  ( .A1(_u10_u7_n1855 ), .A2(_u10_u7_n1869 ), .ZN(_u10_u7_n2862 ) );
NOR2_X1 _u10_u7_U688  ( .A1(_u10_u7_n2886 ), .A2(_u10_u7_n2695 ), .ZN(_u10_u7_n2863 ) );
NAND2_X1 _u10_u7_U687  ( .A1(_u10_u7_n2813 ), .A2(_u10_u7_n2885 ), .ZN(_u10_u7_n2864 ) );
NAND2_X1 _u10_u7_U686  ( .A1(_u10_u7_n2114 ), .A2(_u10_u7_n2884 ), .ZN(_u10_u7_n2865 ) );
NAND2_X1 _u10_u7_U685  ( .A1(1'b0), .A2(_u10_u7_n2667 ), .ZN(_u10_u7_n2112 ));
NOR3_X1 _u10_u7_U684  ( .A1(_u10_u7_n2883 ), .A2(_u10_u7_n2112 ), .A3(_u10_u7_n2719 ), .ZN(_u10_u7_n2878 ) );
INV_X1 _u10_u7_U683  ( .A(_u10_u7_n2112 ), .ZN(_u10_u7_n1856 ) );
NAND2_X1 _u10_u7_U682  ( .A1(_u10_u7_n2364 ), .A2(_u10_u7_n1856 ), .ZN(_u10_u7_n2882 ) );
NAND2_X1 _u10_u7_U681  ( .A1(_u10_u7_n2882 ), .A2(_u10_u7_n1869 ), .ZN(_u10_u7_n2050 ) );
INV_X1 _u10_u7_U680  ( .A(_u10_u7_n2050 ), .ZN(_u10_u7_n1939 ) );
NOR2_X1 _u10_u7_U679  ( .A1(_u10_u7_n1939 ), .A2(_u10_u7_n1841 ), .ZN(_u10_u7_n2881 ) );
NOR2_X1 _u10_u7_U678  ( .A1(_u10_u7_n2881 ), .A2(_u10_u7_n2840 ), .ZN(_u10_u7_n2880 ) );
NOR2_X1 _u10_u7_U677  ( .A1(_u10_u7_n2880 ), .A2(_u10_u7_n1836 ), .ZN(_u10_u7_n2879 ) );
NOR2_X1 _u10_u7_U676  ( .A1(_u10_u7_n2878 ), .A2(_u10_u7_n2879 ), .ZN(_u10_u7_n2866 ) );
NOR2_X1 _u10_u7_U675  ( .A1(_u10_u7_n2081 ), .A2(_u10_u7_n2877 ), .ZN(_u10_u7_n1840 ) );
NAND2_X1 _u10_u7_U674  ( .A1(_u10_u7_n1840 ), .A2(_u10_u7_n2115 ), .ZN(_u10_u7_n1873 ) );
NAND2_X1 _u10_u7_U673  ( .A1(_u10_u7_n2695 ), .A2(_u10_u7_n1940 ), .ZN(_u10_u7_n1874 ) );
NOR3_X1 _u10_u7_U672  ( .A1(_u10_u7_n2050 ), .A2(_u10_u7_n1873 ), .A3(_u10_u7_n1874 ), .ZN(_u10_u7_n2876 ) );
NOR2_X1 _u10_u7_U671  ( .A1(_u10_u7_n2876 ), .A2(_u10_u7_n1913 ), .ZN(_u10_u7_n2868 ) );
NAND2_X1 _u10_u7_U670  ( .A1(_u10_u7_n2875 ), .A2(_u10_u7_n2466 ), .ZN(_u10_u7_n2872 ) );
INV_X1 _u10_u7_U669  ( .A(_u10_u7_n1979 ), .ZN(_u10_u7_n2746 ) );
NAND2_X1 _u10_u7_U668  ( .A1(_u10_u7_n2874 ), .A2(_u10_u7_n2746 ), .ZN(_u10_u7_n1935 ) );
NAND3_X1 _u10_u7_U667  ( .A1(_u10_u7_n1935 ), .A2(_u10_u7_n1936 ), .A3(_u10_u7_n2467 ), .ZN(_u10_u7_n2873 ) );
NAND2_X1 _u10_u7_U666  ( .A1(_u10_u7_n2872 ), .A2(_u10_u7_n2873 ), .ZN(_u10_u7_n2264 ) );
AND2_X1 _u10_u7_U665  ( .A1(_u10_u7_n2264 ), .A2(_u10_u7_n2461 ), .ZN(_u10_u7_n2869 ) );
AND2_X1 _u10_u7_U664  ( .A1(_u10_u7_n1966 ), .A2(_u10_u7_n2761 ), .ZN(_u10_u7_n2870 ) );
NOR2_X1 _u10_u7_U663  ( .A1(_u10_u7_n2159 ), .A2(_u10_u7_n2163 ), .ZN(_u10_u7_n2871 ) );
NOR4_X1 _u10_u7_U662  ( .A1(_u10_u7_n2868 ), .A2(_u10_u7_n2869 ), .A3(_u10_u7_n2870 ), .A4(_u10_u7_n2871 ), .ZN(_u10_u7_n2867 ) );
NAND4_X1 _u10_u7_U661  ( .A1(_u10_u7_n2864 ), .A2(_u10_u7_n2865 ), .A3(_u10_u7_n2866 ), .A4(_u10_u7_n2867 ), .ZN(_u10_u7_n1992 ) );
NOR4_X1 _u10_u7_U660  ( .A1(_u10_u7_n2861 ), .A2(_u10_u7_n2862 ), .A3(_u10_u7_n2863 ), .A4(_u10_u7_n1992 ), .ZN(_u10_u7_n2725 ) );
NAND2_X1 _u10_u7_U659  ( .A1(_u10_u7_n2364 ), .A2(_u10_u7_n1846 ), .ZN(_u10_u7_n2744 ) );
NAND4_X1 _u10_u7_U658  ( .A1(_u10_u7_n2765 ), .A2(_u10_u7_n1939 ), .A3(_u10_u7_n2744 ), .A4(_u10_u7_n2535 ), .ZN(_u10_u7_n2860 ) );
NAND2_X1 _u10_u7_U657  ( .A1(_u10_u7_n2049 ), .A2(_u10_u7_n2860 ), .ZN(_u10_u7_n2856 ) );
NOR4_X1 _u10_u7_U656  ( .A1(1'b0), .A2(_u10_u7_n2858 ), .A3(_u10_u7_n2859 ),.A4(_u10_u7_n2051 ), .ZN(_u10_u7_n2857 ) );
NAND4_X1 _u10_u7_U655  ( .A1(_u10_u7_n2228 ), .A2(_u10_u7_n2855 ), .A3(_u10_u7_n2856 ), .A4(_u10_u7_n2857 ), .ZN(_u10_u7_n2854 ) );
NAND2_X1 _u10_u7_U654  ( .A1(_u10_u7_n2043 ), .A2(_u10_u7_n2854 ), .ZN(_u10_u7_n2821 ) );
INV_X1 _u10_u7_U653  ( .A(_u10_u7_n2071 ), .ZN(_u10_u7_n2279 ) );
INV_X1 _u10_u7_U652  ( .A(_u10_u7_n2599 ), .ZN(_u10_u7_n2357 ) );
OR2_X1 _u10_u7_U651  ( .A1(_u10_u7_n2744 ), .A2(_u10_u7_n2853 ), .ZN(_u10_u7_n2844 ) );
NAND2_X1 _u10_u7_U650  ( .A1(_u10_u7_n2131 ), .A2(_u10_u7_n2852 ), .ZN(_u10_u7_n2851 ) );
NAND2_X1 _u10_u7_U649  ( .A1(_u10_u7_n2082 ), .A2(_u10_u7_n2851 ), .ZN(_u10_u7_n2848 ) );
NAND2_X1 _u10_u7_U648  ( .A1(_u10_u7_n2850 ), .A2(_u10_u7_n2600 ), .ZN(_u10_u7_n2849 ) );
NAND3_X1 _u10_u7_U647  ( .A1(_u10_u7_n2848 ), .A2(_u10_u7_n2077 ), .A3(_u10_u7_n2849 ), .ZN(_u10_u7_n2287 ) );
NAND2_X1 _u10_u7_U646  ( .A1(_u10_u7_n2082 ), .A2(_u10_u7_n2050 ), .ZN(_u10_u7_n2847 ) );
NAND2_X1 _u10_u7_U645  ( .A1(_u10_u7_n2846 ), .A2(_u10_u7_n2847 ), .ZN(_u10_u7_n2074 ) );
NOR3_X1 _u10_u7_U644  ( .A1(_u10_u7_n2287 ), .A2(_u10_u7_n2596 ), .A3(_u10_u7_n2074 ), .ZN(_u10_u7_n2845 ) );
NAND4_X1 _u10_u7_U643  ( .A1(_u10_u7_n2357 ), .A2(_u10_u7_n2837 ), .A3(_u10_u7_n2844 ), .A4(_u10_u7_n2845 ), .ZN(_u10_u7_n2843 ) );
NAND2_X1 _u10_u7_U642  ( .A1(_u10_u7_n2279 ), .A2(_u10_u7_n2843 ), .ZN(_u10_u7_n2822 ) );
NOR3_X1 _u10_u7_U641  ( .A1(_u10_u7_n1925 ), .A2(_u10_u7_n2842 ), .A3(_u10_u7_n2686 ), .ZN(_u10_u7_n2841 ) );
NOR3_X1 _u10_u7_U640  ( .A1(_u10_u7_n2840 ), .A2(_u10_u7_n2599 ), .A3(_u10_u7_n2841 ), .ZN(_u10_u7_n2839 ) );
AND4_X1 _u10_u7_U639  ( .A1(_u10_u7_n2836 ), .A2(_u10_u7_n2837 ), .A3(_u10_u7_n2838 ), .A4(_u10_u7_n2839 ), .ZN(_u10_u7_n2454 ) );
NOR2_X1 _u10_u7_U638  ( .A1(_u10_u7_n2719 ), .A2(_u10_u7_n2835 ), .ZN(_u10_u7_n2773 ) );
NOR2_X1 _u10_u7_U637  ( .A1(_u10_u7_n2138 ), .A2(_u10_u7_n2773 ), .ZN(_u10_u7_n2814 ) );
NAND2_X1 _u10_u7_U636  ( .A1(_u10_u7_n2814 ), .A2(_u10_u7_n1869 ), .ZN(_u10_u7_n2834 ) );
NAND2_X1 _u10_u7_U635  ( .A1(_u10_u7_n2833 ), .A2(_u10_u7_n2834 ), .ZN(_u10_u7_n2832 ) );
NAND2_X1 _u10_u7_U634  ( .A1(_u10_u7_n2454 ), .A2(_u10_u7_n2832 ), .ZN(_u10_u7_n2831 ) );
NAND2_X1 _u10_u7_U633  ( .A1(_u10_u7_n2830 ), .A2(_u10_u7_n2831 ), .ZN(_u10_u7_n2823 ) );
INV_X1 _u10_u7_U632  ( .A(_u10_u7_n2025 ), .ZN(_u10_u7_n2470 ) );
NAND2_X1 _u10_u7_U631  ( .A1(_u10_u7_n1979 ), .A2(_u10_u7_n1936 ), .ZN(_u10_u7_n2829 ) );
AND2_X1 _u10_u7_U630  ( .A1(_u10_u7_n2828 ), .A2(_u10_u7_n2829 ), .ZN(_u10_u7_n2469 ) );
NAND2_X1 _u10_u7_U629  ( .A1(_u10_u7_n2469 ), .A2(_u10_u7_n2269 ), .ZN(_u10_u7_n2161 ) );
INV_X1 _u10_u7_U628  ( .A(_u10_u7_n2161 ), .ZN(_u10_u7_n2276 ) );
NOR2_X1 _u10_u7_U627  ( .A1(_u10_u7_n2274 ), .A2(_u10_u7_n2719 ), .ZN(_u10_u7_n2827 ) );
NOR3_X1 _u10_u7_U626  ( .A1(_u10_u7_n2827 ), .A2(_u10_u7_n2742 ), .A3(_u10_u7_n2680 ), .ZN(_u10_u7_n2826 ) );
NAND3_X1 _u10_u7_U625  ( .A1(_u10_u7_n2276 ), .A2(_u10_u7_n2108 ), .A3(_u10_u7_n2826 ), .ZN(_u10_u7_n2825 ) );
NAND2_X1 _u10_u7_U624  ( .A1(_u10_u7_n2470 ), .A2(_u10_u7_n2825 ), .ZN(_u10_u7_n2824 ) );
NAND4_X1 _u10_u7_U623  ( .A1(_u10_u7_n2821 ), .A2(_u10_u7_n2822 ), .A3(_u10_u7_n2823 ), .A4(_u10_u7_n2824 ), .ZN(_u10_u7_n2804 ) );
NAND2_X1 _u10_u7_U622  ( .A1(_u10_u7_n2131 ), .A2(_u10_u7_n2744 ), .ZN(_u10_u7_n2820 ) );
NAND2_X1 _u10_u7_U621  ( .A1(_u10_u7_n2571 ), .A2(_u10_u7_n2820 ), .ZN(_u10_u7_n2817 ) );
NOR2_X1 _u10_u7_U620  ( .A1(_u10_u7_n2819 ), .A2(_u10_u7_n2436 ), .ZN(_u10_u7_n2818 ) );
NAND4_X1 _u10_u7_U619  ( .A1(_u10_u7_n2437 ), .A2(_u10_u7_n2355 ), .A3(_u10_u7_n2817 ), .A4(_u10_u7_n2818 ), .ZN(_u10_u7_n2816 ) );
NAND2_X1 _u10_u7_U618  ( .A1(_u10_u7_n2815 ), .A2(_u10_u7_n2816 ), .ZN(_u10_u7_n2809 ) );
INV_X1 _u10_u7_U617  ( .A(_u10_u7_n2814 ), .ZN(_u10_u7_n2812 ) );
OR2_X1 _u10_u7_U616  ( .A1(_u10_u7_n1911 ), .A2(_u10_u7_n2813 ), .ZN(_u10_u7_n1884 ) );
NAND2_X1 _u10_u7_U615  ( .A1(_u10_u7_n2812 ), .A2(_u10_u7_n1884 ), .ZN(_u10_u7_n2810 ) );
NOR2_X1 _u10_u7_U614  ( .A1(_u10_u7_n1894 ), .A2(_u10_u7_n2461 ), .ZN(_u10_u7_n1948 ) );
OR2_X1 _u10_u7_U613  ( .A1(_u10_u7_n1847 ), .A2(_u10_u7_n1948 ), .ZN(_u10_u7_n2811 ) );
NAND3_X1 _u10_u7_U612  ( .A1(_u10_u7_n2809 ), .A2(_u10_u7_n2810 ), .A3(_u10_u7_n2811 ), .ZN(_u10_u7_n2805 ) );
NOR2_X1 _u10_u7_U611  ( .A1(_u10_u7_n2808 ), .A2(_u10_u7_n2775 ), .ZN(_u10_u7_n2806 ) );
AND2_X1 _u10_u7_U610  ( .A1(_u10_u7_n2721 ), .A2(_u10_u7_n1911 ), .ZN(_u10_u7_n2807 ) );
NOR4_X1 _u10_u7_U609  ( .A1(_u10_u7_n2804 ), .A2(_u10_u7_n2805 ), .A3(_u10_u7_n2806 ), .A4(_u10_u7_n2807 ), .ZN(_u10_u7_n2726 ) );
NAND2_X1 _u10_u7_U608  ( .A1(_u10_u7_n2803 ), .A2(_u10_u7_n2112 ), .ZN(_u10_u7_n2802 ) );
NAND2_X1 _u10_u7_U607  ( .A1(_u10_u7_n2364 ), .A2(_u10_u7_n2802 ), .ZN(_u10_u7_n2801 ) );
NAND2_X1 _u10_u7_U606  ( .A1(_u10_u7_n2800 ), .A2(_u10_u7_n2801 ), .ZN(_u10_u7_n2799 ) );
NAND2_X1 _u10_u7_U605  ( .A1(_u10_u7_n1937 ), .A2(_u10_u7_n2799 ), .ZN(_u10_u7_n2780 ) );
NAND2_X1 _u10_u7_U604  ( .A1(_u10_u7_n2775 ), .A2(_u10_u7_n2798 ), .ZN(_u10_u7_n2796 ) );
INV_X1 _u10_u7_U603  ( .A(_u10_u7_n2131 ), .ZN(_u10_u7_n2797 ) );
NAND2_X1 _u10_u7_U602  ( .A1(_u10_u7_n2796 ), .A2(_u10_u7_n2797 ), .ZN(_u10_u7_n2781 ) );
OR4_X1 _u10_u7_U601  ( .A1(_u10_u7_n2795 ), .A2(_u10_u7_n2303 ), .A3(_u10_u7_n2553 ), .A4(_u10_u7_n2554 ), .ZN(_u10_u7_n2792 ) );
NAND3_X1 _u10_u7_U600  ( .A1(_u10_u7_n1847 ), .A2(_u10_u7_n2097 ), .A3(_u10_u7_n2096 ), .ZN(_u10_u7_n2793 ) );
NOR4_X1 _u10_u7_U599  ( .A1(_u10_u7_n2792 ), .A2(_u10_u7_n2793 ), .A3(_u10_u7_n2542 ), .A4(_u10_u7_n2794 ), .ZN(_u10_u7_n2791 ) );
NOR2_X1 _u10_u7_U598  ( .A1(_u10_u7_n2791 ), .A2(_u10_u7_n2085 ), .ZN(_u10_u7_n2783 ) );
NAND2_X1 _u10_u7_U597  ( .A1(_u10_u7_n2114 ), .A2(_u10_u7_n2049 ), .ZN(_u10_u7_n2700 ) );
INV_X1 _u10_u7_U596  ( .A(_u10_u7_n2700 ), .ZN(_u10_u7_n2784 ) );
NAND4_X1 _u10_u7_U595  ( .A1(_u10_u7_n2001 ), .A2(_u10_u7_n2547 ), .A3(_u10_u7_n2368 ), .A4(_u10_u7_n1847 ), .ZN(_u10_u7_n2787 ) );
NOR4_X1 _u10_u7_U594  ( .A1(_u10_u7_n2787 ), .A2(_u10_u7_n2788 ), .A3(_u10_u7_n2789 ), .A4(_u10_u7_n2790 ), .ZN(_u10_u7_n2786 ) );
NOR2_X1 _u10_u7_U593  ( .A1(_u10_u7_n2786 ), .A2(_u10_u7_n2000 ), .ZN(_u10_u7_n2785 ) );
NOR3_X1 _u10_u7_U592  ( .A1(_u10_u7_n2783 ), .A2(_u10_u7_n2784 ), .A3(_u10_u7_n2785 ), .ZN(_u10_u7_n2782 ) );
NAND3_X1 _u10_u7_U591  ( .A1(_u10_u7_n2780 ), .A2(_u10_u7_n2781 ), .A3(_u10_u7_n2782 ), .ZN(_u10_u7_n2728 ) );
OR3_X1 _u10_u7_U590  ( .A1(_u10_u7_n2138 ), .A2(_u10_u7_n2633 ), .A3(_u10_u7_n2779 ), .ZN(_u10_u7_n2778 ) );
NAND2_X1 _u10_u7_U589  ( .A1(_u10_u7_n2777 ), .A2(_u10_u7_n2778 ), .ZN(_u10_u7_n2767 ) );
NAND3_X1 _u10_u7_U588  ( .A1(_u10_u7_n2775 ), .A2(_u10_u7_n2083 ), .A3(_u10_u7_n2776 ), .ZN(_u10_u7_n2774 ) );
NAND2_X1 _u10_u7_U587  ( .A1(_u10_u7_n2773 ), .A2(_u10_u7_n2774 ), .ZN(_u10_u7_n2768 ) );
NAND2_X1 _u10_u7_U586  ( .A1(_u10_u7_n2218 ), .A2(_u10_u7_n2772 ), .ZN(_u10_u7_n2769 ) );
NAND2_X1 _u10_u7_U585  ( .A1(_u10_u7_n2302 ), .A2(_u10_u7_n2467 ), .ZN(_u10_u7_n2771 ) );
NAND2_X1 _u10_u7_U584  ( .A1(_u10_u7_n2461 ), .A2(_u10_u7_n2771 ), .ZN(_u10_u7_n2770 ) );
NAND4_X1 _u10_u7_U583  ( .A1(_u10_u7_n2767 ), .A2(_u10_u7_n2768 ), .A3(_u10_u7_n2769 ), .A4(_u10_u7_n2770 ), .ZN(_u10_u7_n2729 ) );
NAND3_X1 _u10_u7_U582  ( .A1(_u10_u7_n2668 ), .A2(_u10_u7_n2600 ), .A3(_u10_u7_n2276 ), .ZN(_u10_u7_n2766 ) );
NAND2_X1 _u10_u7_U581  ( .A1(_u10_u7_n1894 ), .A2(_u10_u7_n2766 ), .ZN(_u10_u7_n2753 ) );
NAND3_X1 _u10_u7_U580  ( .A1(_u10_u7_n2456 ), .A2(_u10_u7_n2744 ), .A3(_u10_u7_n2765 ), .ZN(_u10_u7_n2764 ) );
NAND2_X1 _u10_u7_U579  ( .A1(_u10_u7_n2377 ), .A2(_u10_u7_n2764 ), .ZN(_u10_u7_n2754 ) );
NAND2_X1 _u10_u7_U578  ( .A1(_u10_u7_n2763 ), .A2(_u10_u7_n2007 ), .ZN(_u10_u7_n2755 ) );
NOR2_X1 _u10_u7_U577  ( .A1(_u10_u7_n2531 ), .A2(_u10_u7_n2744 ), .ZN(_u10_u7_n2760 ) );
INV_X1 _u10_u7_U576  ( .A(_u10_u7_n2762 ), .ZN(_u10_u7_n2189 ) );
NOR3_X1 _u10_u7_U575  ( .A1(_u10_u7_n2760 ), .A2(_u10_u7_n2761 ), .A3(_u10_u7_n2189 ), .ZN(_u10_u7_n2759 ) );
NOR2_X1 _u10_u7_U574  ( .A1(_u10_u7_n2759 ), .A2(_u10_u7_n1849 ), .ZN(_u10_u7_n2757 ) );
NOR2_X1 _u10_u7_U573  ( .A1(_u10_u7_n1817 ), .A2(_u10_u7_n2665 ), .ZN(_u10_u7_n2758 ) );
NOR2_X1 _u10_u7_U572  ( .A1(_u10_u7_n2757 ), .A2(_u10_u7_n2758 ), .ZN(_u10_u7_n2756 ) );
NAND4_X1 _u10_u7_U571  ( .A1(_u10_u7_n2753 ), .A2(_u10_u7_n2754 ), .A3(_u10_u7_n2755 ), .A4(_u10_u7_n2756 ), .ZN(_u10_u7_n2730 ) );
INV_X1 _u10_u7_U570  ( .A(_u10_u7_n2359 ), .ZN(_u10_u7_n1899 ) );
NAND4_X1 _u10_u7_U569  ( .A1(_u10_u7_n2078 ), .A2(_u10_u7_n2580 ), .A3(_u10_u7_n2748 ), .A4(_u10_u7_n2752 ), .ZN(_u10_u7_n2751 ) );
NAND2_X1 _u10_u7_U568  ( .A1(_u10_u7_n1899 ), .A2(_u10_u7_n2751 ), .ZN(_u10_u7_n2732 ) );
INV_X1 _u10_u7_U567  ( .A(_u10_u7_n2750 ), .ZN(_u10_u7_n2379 ) );
NAND3_X1 _u10_u7_U566  ( .A1(_u10_u7_n1856 ), .A2(_u10_u7_n2669 ), .A3(_u10_u7_n2364 ), .ZN(_u10_u7_n2749 ) );
AND2_X1 _u10_u7_U565  ( .A1(_u10_u7_n2748 ), .A2(_u10_u7_n2749 ), .ZN(_u10_u7_n2034 ) );
NAND2_X1 _u10_u7_U564  ( .A1(_u10_u7_n2105 ), .A2(_u10_u7_n2669 ), .ZN(_u10_u7_n2745 ) );
AND3_X1 _u10_u7_U563  ( .A1(_u10_u7_n2745 ), .A2(_u10_u7_n2746 ), .A3(_u10_u7_n2747 ), .ZN(_u10_u7_n2380 ) );
NOR2_X1 _u10_u7_U562  ( .A1(_u10_u7_n2274 ), .A2(_u10_u7_n2744 ), .ZN(_u10_u7_n2743 ) );
NOR4_X1 _u10_u7_U561  ( .A1(_u10_u7_n2742 ), .A2(_u10_u7_n2680 ), .A3(_u10_u7_n2743 ), .A4(_u10_u7_n2428 ), .ZN(_u10_u7_n2741 ) );
NAND4_X1 _u10_u7_U560  ( .A1(_u10_u7_n2379 ), .A2(_u10_u7_n2034 ), .A3(_u10_u7_n2380 ), .A4(_u10_u7_n2741 ), .ZN(_u10_u7_n2740 ) );
NAND2_X1 _u10_u7_U559  ( .A1(_u10_u7_n1967 ), .A2(_u10_u7_n2740 ), .ZN(_u10_u7_n2733 ) );
NAND3_X1 _u10_u7_U558  ( .A1(_u10_u7_n2739 ), .A2(_u10_u7_n2368 ), .A3(_u10_u7_n2255 ), .ZN(_u10_u7_n2738 ) );
NAND2_X1 _u10_u7_U557  ( .A1(_u10_u7_n2737 ), .A2(_u10_u7_n2738 ), .ZN(_u10_u7_n2734 ) );
NAND2_X1 _u10_u7_U556  ( .A1(_u10_u7_n2736 ), .A2(_u10_u7_n2524 ), .ZN(_u10_u7_n2735 ) );
NAND4_X1 _u10_u7_U555  ( .A1(_u10_u7_n2732 ), .A2(_u10_u7_n2733 ), .A3(_u10_u7_n2734 ), .A4(_u10_u7_n2735 ), .ZN(_u10_u7_n2731 ) );
NOR4_X1 _u10_u7_U554  ( .A1(_u10_u7_n2728 ), .A2(_u10_u7_n2729 ), .A3(_u10_u7_n2730 ), .A4(_u10_u7_n2731 ), .ZN(_u10_u7_n2727 ) );
NAND4_X1 _u10_u7_U553  ( .A1(_u10_u7_n2724 ), .A2(_u10_u7_n2725 ), .A3(_u10_u7_n2726 ), .A4(_u10_u7_n2727 ), .ZN(_u10_u7_n2723 ) );
MUX2_X1 _u10_u7_U552  ( .A(_u10_u7_n2723 ), .B(_u10_SYNOPSYS_UNCONNECTED_29 ), .S(_u10_u7_n1819 ), .Z(_u10_u7_n1809 ) );
NAND2_X1 _u10_u7_U551  ( .A1(_u10_u7_n2002 ), .A2(_u10_u7_n2722 ), .ZN(_u10_u7_n2713 ) );
NAND2_X1 _u10_u7_U550  ( .A1(_u10_u7_n2720 ), .A2(_u10_u7_n2721 ), .ZN(_u10_u7_n2714 ) );
NAND2_X1 _u10_u7_U549  ( .A1(_u10_u7_n2256 ), .A2(_u10_u7_n2719 ), .ZN(_u10_u7_n2715 ) );
NOR2_X1 _u10_u7_U548  ( .A1(_u10_u7_n2106 ), .A2(_u10_u7_n2037 ), .ZN(_u10_u7_n2717 ) );
AND2_X1 _u10_u7_U547  ( .A1(_u10_u7_n1966 ), .A2(_u10_u7_n2054 ), .ZN(_u10_u7_n2718 ) );
NOR2_X1 _u10_u7_U546  ( .A1(_u10_u7_n2717 ), .A2(_u10_u7_n2718 ), .ZN(_u10_u7_n2716 ) );
NAND4_X1 _u10_u7_U545  ( .A1(_u10_u7_n2713 ), .A2(_u10_u7_n2714 ), .A3(_u10_u7_n2715 ), .A4(_u10_u7_n2716 ), .ZN(_u10_u7_n2608 ) );
NAND2_X1 _u10_u7_U544  ( .A1(1'b0), .A2(_u10_u7_n2669 ), .ZN(_u10_u7_n2385 ));
INV_X1 _u10_u7_U543  ( .A(_u10_u7_n2385 ), .ZN(_u10_u7_n1977 ) );
NAND2_X1 _u10_u7_U542  ( .A1(_u10_u7_n1977 ), .A2(_u10_u7_n2668 ), .ZN(_u10_u7_n2712 ) );
NAND2_X1 _u10_u7_U541  ( .A1(_u10_u7_n2712 ), .A2(_u10_u7_n2092 ), .ZN(_u10_u7_n1844 ) );
NAND2_X1 _u10_u7_U540  ( .A1(_u10_u7_n1894 ), .A2(_u10_u7_n1844 ), .ZN(_u10_u7_n2705 ) );
NAND2_X1 _u10_u7_U539  ( .A1(_u10_u7_n1894 ), .A2(_u10_u7_n2305 ), .ZN(_u10_u7_n2711 ) );
NAND2_X1 _u10_u7_U538  ( .A1(_u10_u7_n2711 ), .A2(_u10_u7_n2025 ), .ZN(_u10_u7_n1932 ) );
NAND2_X1 _u10_u7_U537  ( .A1(_u10_u7_n2710 ), .A2(_u10_u7_n1932 ), .ZN(_u10_u7_n2706 ) );
NAND2_X1 _u10_u7_U536  ( .A1(_u10_u7_n2708 ), .A2(_u10_u7_n2709 ), .ZN(_u10_u7_n2707 ) );
NAND3_X1 _u10_u7_U535  ( .A1(_u10_u7_n2705 ), .A2(_u10_u7_n2706 ), .A3(_u10_u7_n2707 ), .ZN(_u10_u7_n2701 ) );
NOR2_X1 _u10_u7_U534  ( .A1(_u10_u7_n1843 ), .A2(_u10_u7_n2545 ), .ZN(_u10_u7_n2702 ) );
NOR2_X1 _u10_u7_U533  ( .A1(_u10_u7_n2346 ), .A2(_u10_u7_n2700 ), .ZN(_u10_u7_n2703 ) );
NOR2_X1 _u10_u7_U532  ( .A1(_u10_u7_n2000 ), .A2(_u10_u7_n1887 ), .ZN(_u10_u7_n2704 ) );
NOR4_X1 _u10_u7_U531  ( .A1(_u10_u7_n2701 ), .A2(_u10_u7_n2702 ), .A3(_u10_u7_n2703 ), .A4(_u10_u7_n2704 ), .ZN(_u10_u7_n2671 ) );
NAND2_X1 _u10_u7_U530  ( .A1(_u10_u7_n2699 ), .A2(_u10_u7_n2700 ), .ZN(_u10_u7_n2698 ) );
NAND2_X1 _u10_u7_U529  ( .A1(_u10_u7_n2063 ), .A2(_u10_u7_n2698 ), .ZN(_u10_u7_n2682 ) );
NAND2_X1 _u10_u7_U528  ( .A1(_u10_u7_n2697 ), .A2(_u10_u7_n2103 ), .ZN(_u10_u7_n2696 ) );
NAND2_X1 _u10_u7_U527  ( .A1(_u10_u7_n2695 ), .A2(_u10_u7_n2696 ), .ZN(_u10_u7_n2694 ) );
NAND2_X1 _u10_u7_U526  ( .A1(_u10_u7_n1937 ), .A2(_u10_u7_n2694 ), .ZN(_u10_u7_n2683 ) );
INV_X1 _u10_u7_U525  ( .A(_u10_u7_n2693 ), .ZN(_u10_u7_n2691 ) );
NAND3_X1 _u10_u7_U524  ( .A1(_u10_u7_n2103 ), .A2(_u10_u7_n2502 ), .A3(1'b0),.ZN(_u10_u7_n2692 ) );
NAND2_X1 _u10_u7_U523  ( .A1(_u10_u7_n2691 ), .A2(_u10_u7_n2692 ), .ZN(_u10_u7_n2690 ) );
NAND2_X1 _u10_u7_U522  ( .A1(_u10_u7_n2236 ), .A2(_u10_u7_n2690 ), .ZN(_u10_u7_n2684 ) );
NAND3_X1 _u10_u7_U521  ( .A1(_u10_u7_n2688 ), .A2(_u10_u7_n1913 ), .A3(_u10_u7_n2689 ), .ZN(_u10_u7_n2335 ) );
NAND3_X1 _u10_u7_U520  ( .A1(_u10_u7_n2536 ), .A2(_u10_u7_n2103 ), .A3(1'b0),.ZN(_u10_u7_n2052 ) );
NOR2_X1 _u10_u7_U519  ( .A1(_u10_u7_n2052 ), .A2(_u10_u7_n2687 ), .ZN(_u10_u7_n1851 ) );
NAND2_X1 _u10_u7_U518  ( .A1(_u10_u7_n1851 ), .A2(_u10_u7_n2078 ), .ZN(_u10_u7_n2582 ) );
NOR2_X1 _u10_u7_U517  ( .A1(_u10_u7_n2686 ), .A2(_u10_u7_n2582 ), .ZN(_u10_u7_n2094 ) );
NAND3_X1 _u10_u7_U516  ( .A1(_u10_u7_n2251 ), .A2(_u10_u7_n2335 ), .A3(_u10_u7_n2094 ), .ZN(_u10_u7_n2685 ) );
NAND4_X1 _u10_u7_U515  ( .A1(_u10_u7_n2682 ), .A2(_u10_u7_n2683 ), .A3(_u10_u7_n2684 ), .A4(_u10_u7_n2685 ), .ZN(_u10_u7_n2673 ) );
INV_X1 _u10_u7_U514  ( .A(_u10_u7_n2291 ), .ZN(_u10_u7_n2057 ) );
AND2_X1 _u10_u7_U513  ( .A1(_u10_u7_n1851 ), .A2(_u10_u7_n2057 ), .ZN(_u10_u7_n2674 ) );
INV_X1 _u10_u7_U512  ( .A(_u10_u7_n1874 ), .ZN(_u10_u7_n2681 ) );
NOR2_X1 _u10_u7_U511  ( .A1(_u10_u7_n2007 ), .A2(_u10_u7_n1911 ), .ZN(_u10_u7_n2486 ) );
NOR2_X1 _u10_u7_U510  ( .A1(_u10_u7_n2681 ), .A2(_u10_u7_n2486 ), .ZN(_u10_u7_n2675 ) );
NOR2_X1 _u10_u7_U509  ( .A1(_u10_u7_n1977 ), .A2(_u10_u7_n2680 ), .ZN(_u10_u7_n2679 ) );
NOR2_X1 _u10_u7_U508  ( .A1(_u10_u7_n2679 ), .A2(_u10_u7_n2030 ), .ZN(_u10_u7_n2678 ) );
NOR2_X1 _u10_u7_U507  ( .A1(_u10_u7_n2678 ), .A2(_u10_u7_n2094 ), .ZN(_u10_u7_n2677 ) );
NOR2_X1 _u10_u7_U506  ( .A1(_u10_u7_n2677 ), .A2(_u10_u7_n2025 ), .ZN(_u10_u7_n2676 ) );
NOR4_X1 _u10_u7_U505  ( .A1(_u10_u7_n2673 ), .A2(_u10_u7_n2674 ), .A3(_u10_u7_n2675 ), .A4(_u10_u7_n2676 ), .ZN(_u10_u7_n2672 ) );
AND2_X1 _u10_u7_U504  ( .A1(_u10_u7_n2671 ), .A2(_u10_u7_n2672 ), .ZN(_u10_u7_n1990 ) );
INV_X1 _u10_u7_U503  ( .A(_u10_u7_n2670 ), .ZN(_u10_u7_n2660 ) );
NAND4_X1 _u10_u7_U502  ( .A1(_u10_u7_n2251 ), .A2(_u10_u7_n2669 ), .A3(_u10_u7_n2162 ), .A4(_u10_u7_n2169 ), .ZN(_u10_u7_n2664 ) );
AND3_X1 _u10_u7_U501  ( .A1(_u10_u7_n1977 ), .A2(_u10_u7_n2668 ), .A3(_u10_u7_n2089 ), .ZN(_u10_u7_n2555 ) );
NAND2_X1 _u10_u7_U500  ( .A1(_u10_u7_n2555 ), .A2(_u10_u7_n2667 ), .ZN(_u10_u7_n2666 ) );
NAND3_X1 _u10_u7_U499  ( .A1(_u10_u7_n2664 ), .A2(_u10_u7_n2665 ), .A3(_u10_u7_n2666 ), .ZN(_u10_u7_n1988 ) );
INV_X1 _u10_u7_U498  ( .A(_u10_u7_n1988 ), .ZN(_u10_u7_n2661 ) );
NAND2_X1 _u10_u7_U497  ( .A1(1'b0), .A2(_u10_u7_n2043 ), .ZN(_u10_u7_n2662 ));
NAND2_X1 _u10_u7_U496  ( .A1(_u10_u7_n2169 ), .A2(1'b0), .ZN(_u10_u7_n2663 ));
NAND4_X1 _u10_u7_U495  ( .A1(_u10_u7_n2660 ), .A2(_u10_u7_n2661 ), .A3(_u10_u7_n2662 ), .A4(_u10_u7_n2663 ), .ZN(_u10_u7_n2650 ) );
NAND2_X1 _u10_u7_U494  ( .A1(_u10_u7_n2659 ), .A2(1'b0), .ZN(_u10_u7_n2193 ));
INV_X1 _u10_u7_U493  ( .A(_u10_u7_n2193 ), .ZN(_u10_u7_n2143 ) );
NAND2_X1 _u10_u7_U492  ( .A1(_u10_u7_n2143 ), .A2(_u10_u7_n2036 ), .ZN(_u10_u7_n2286 ) );
INV_X1 _u10_u7_U491  ( .A(_u10_u7_n2286 ), .ZN(_u10_u7_n2577 ) );
NAND2_X1 _u10_u7_U490  ( .A1(_u10_u7_n2577 ), .A2(_u10_u7_n2278 ), .ZN(_u10_u7_n2474 ) );
INV_X1 _u10_u7_U489  ( .A(_u10_u7_n2474 ), .ZN(_u10_u7_n2306 ) );
NAND2_X1 _u10_u7_U488  ( .A1(_u10_u7_n2306 ), .A2(_u10_u7_n2251 ), .ZN(_u10_u7_n2654 ) );
NAND2_X1 _u10_u7_U487  ( .A1(_u10_u7_n2649 ), .A2(_u10_u7_n2658 ), .ZN(_u10_u7_n2655 ) );
NAND2_X1 _u10_u7_U486  ( .A1(_u10_u7_n2657 ), .A2(_u10_u7_n2445 ), .ZN(_u10_u7_n2656 ) );
NAND3_X1 _u10_u7_U485  ( .A1(_u10_u7_n2654 ), .A2(_u10_u7_n2655 ), .A3(_u10_u7_n2656 ), .ZN(_u10_u7_n2651 ) );
NOR2_X1 _u10_u7_U484  ( .A1(_u10_u7_n2366 ), .A2(_u10_u7_n2376 ), .ZN(_u10_u7_n2652 ) );
AND2_X1 _u10_u7_U483  ( .A1(_u10_u7_n1966 ), .A2(_u10_u7_n2528 ), .ZN(_u10_u7_n2653 ) );
NOR4_X1 _u10_u7_U482  ( .A1(_u10_u7_n2650 ), .A2(_u10_u7_n2651 ), .A3(_u10_u7_n2652 ), .A4(_u10_u7_n2653 ), .ZN(_u10_u7_n2613 ) );
NAND2_X1 _u10_u7_U481  ( .A1(_u10_u7_n1891 ), .A2(1'b0), .ZN(_u10_u7_n2636 ));
NAND2_X1 _u10_u7_U480  ( .A1(_u10_u7_n1868 ), .A2(_u10_u7_n2113 ), .ZN(_u10_u7_n2101 ) );
NOR4_X1 _u10_u7_U479  ( .A1(_u10_u7_n2649 ), .A2(_u10_u7_n2216 ), .A3(_u10_u7_n2101 ), .A4(_u10_u7_n2634 ), .ZN(_u10_u7_n2648 ) );
NOR2_X1 _u10_u7_U478  ( .A1(_u10_u7_n2648 ), .A2(_u10_u7_n2254 ), .ZN(_u10_u7_n2638 ) );
NOR2_X1 _u10_u7_U477  ( .A1(_u10_u7_n2106 ), .A2(_u10_u7_n2643 ), .ZN(_u10_u7_n2645 ) );
NAND2_X1 _u10_u7_U476  ( .A1(1'b0), .A2(_u10_u7_n2049 ), .ZN(_u10_u7_n2647 ));
NAND2_X1 _u10_u7_U475  ( .A1(_u10_u7_n2646 ), .A2(_u10_u7_n2647 ), .ZN(_u10_u7_n2348 ) );
NOR2_X1 _u10_u7_U474  ( .A1(_u10_u7_n2645 ), .A2(_u10_u7_n2348 ), .ZN(_u10_u7_n2644 ) );
NOR2_X1 _u10_u7_U473  ( .A1(_u10_u7_n2644 ), .A2(_u10_u7_n2495 ), .ZN(_u10_u7_n2639 ) );
NOR2_X1 _u10_u7_U472  ( .A1(_u10_u7_n2643 ), .A2(_u10_u7_n2203 ), .ZN(_u10_u7_n2642 ) );
NOR3_X1 _u10_u7_U471  ( .A1(_u10_u7_n2101 ), .A2(1'b0), .A3(_u10_u7_n2642 ),.ZN(_u10_u7_n2641 ) );
NOR2_X1 _u10_u7_U470  ( .A1(_u10_u7_n2641 ), .A2(_u10_u7_n2253 ), .ZN(_u10_u7_n2640 ) );
NOR3_X1 _u10_u7_U469  ( .A1(_u10_u7_n2638 ), .A2(_u10_u7_n2639 ), .A3(_u10_u7_n2640 ), .ZN(_u10_u7_n2637 ) );
NAND3_X1 _u10_u7_U468  ( .A1(_u10_u7_n2635 ), .A2(_u10_u7_n2636 ), .A3(_u10_u7_n2637 ), .ZN(_u10_u7_n2615 ) );
NOR3_X1 _u10_u7_U467  ( .A1(_u10_u7_n2174 ), .A2(_u10_u7_n2175 ), .A3(_u10_u7_n2179 ), .ZN(_u10_u7_n2631 ) );
NAND3_X1 _u10_u7_U466  ( .A1(_u10_u7_n2223 ), .A2(_u10_u7_n2236 ), .A3(_u10_u7_n2631 ), .ZN(_u10_u7_n2622 ) );
OR2_X1 _u10_u7_U465  ( .A1(_u10_u7_n1960 ), .A2(_u10_u7_n1959 ), .ZN(_u10_u7_n2625 ) );
NOR3_X1 _u10_u7_U464  ( .A1(_u10_u7_n2101 ), .A2(_u10_u7_n2633 ), .A3(_u10_u7_n2634 ), .ZN(_u10_u7_n2523 ) );
OR2_X1 _u10_u7_U463  ( .A1(_u10_u7_n2632 ), .A2(_u10_u7_n2523 ), .ZN(_u10_u7_n2627 ) );
INV_X1 _u10_u7_U462  ( .A(_u10_u7_n2631 ), .ZN(_u10_u7_n2628 ) );
NAND2_X1 _u10_u7_U461  ( .A1(_u10_u7_n2630 ), .A2(_u10_u7_n1922 ), .ZN(_u10_u7_n2629 ) );
NAND3_X1 _u10_u7_U460  ( .A1(_u10_u7_n2627 ), .A2(_u10_u7_n2628 ), .A3(_u10_u7_n2629 ), .ZN(_u10_u7_n2626 ) );
NAND2_X1 _u10_u7_U459  ( .A1(_u10_u7_n2625 ), .A2(_u10_u7_n2626 ), .ZN(_u10_u7_n2624 ) );
NAND3_X1 _u10_u7_U458  ( .A1(_u10_u7_n2622 ), .A2(_u10_u7_n2623 ), .A3(_u10_u7_n2624 ), .ZN(_u10_u7_n2616 ) );
AND2_X1 _u10_u7_U457  ( .A1(_u10_u7_n2621 ), .A2(_u10_u7_n2358 ), .ZN(_u10_u7_n2620 ) );
NOR2_X1 _u10_u7_U456  ( .A1(_u10_u7_n2523 ), .A2(_u10_u7_n2620 ), .ZN(_u10_u7_n2617 ) );
INV_X1 _u10_u7_U455  ( .A(_u10_u7_n2101 ), .ZN(_u10_u7_n2221 ) );
NOR2_X1 _u10_u7_U454  ( .A1(_u10_u7_n1911 ), .A2(_u10_u7_n2488 ), .ZN(_u10_u7_n2619 ) );
NOR2_X1 _u10_u7_U453  ( .A1(_u10_u7_n2221 ), .A2(_u10_u7_n2619 ), .ZN(_u10_u7_n2618 ) );
NOR4_X1 _u10_u7_U452  ( .A1(_u10_u7_n2615 ), .A2(_u10_u7_n2616 ), .A3(_u10_u7_n2617 ), .A4(_u10_u7_n2618 ), .ZN(_u10_u7_n2614 ) );
AND2_X1 _u10_u7_U451  ( .A1(_u10_u7_n2613 ), .A2(_u10_u7_n2614 ), .ZN(_u10_u7_n2314 ) );
NAND3_X1 _u10_u7_U450  ( .A1(_u10_u7_n2612 ), .A2(_u10_u7_n1990 ), .A3(_u10_u7_n2314 ), .ZN(_u10_u7_n2609 ) );
NOR4_X1 _u10_u7_U449  ( .A1(_u10_u7_n2608 ), .A2(_u10_u7_n2609 ), .A3(_u10_u7_n2610 ), .A4(_u10_u7_n2611 ), .ZN(_u10_u7_n2388 ) );
NAND2_X1 _u10_u7_U448  ( .A1(_u10_u7_n2346 ), .A2(_u10_u7_n2607 ), .ZN(_u10_u7_n2191 ) );
NAND2_X1 _u10_u7_U447  ( .A1(_u10_u7_n2143 ), .A2(_u10_u7_n2191 ), .ZN(_u10_u7_n2556 ) );
INV_X1 _u10_u7_U446  ( .A(_u10_u7_n2348 ), .ZN(_u10_u7_n2603 ) );
NAND3_X1 _u10_u7_U445  ( .A1(_u10_u7_n2535 ), .A2(_u10_u7_n2485 ), .A3(_u10_u7_n2456 ), .ZN(_u10_u7_n2606 ) );
NAND2_X1 _u10_u7_U444  ( .A1(_u10_u7_n2049 ), .A2(_u10_u7_n2606 ), .ZN(_u10_u7_n2604 ) );
NAND3_X1 _u10_u7_U443  ( .A1(_u10_u7_n2603 ), .A2(_u10_u7_n2604 ), .A3(_u10_u7_n2605 ), .ZN(_u10_u7_n2602 ) );
NAND2_X1 _u10_u7_U442  ( .A1(_u10_u7_n2043 ), .A2(_u10_u7_n2602 ), .ZN(_u10_u7_n2557 ) );
INV_X1 _u10_u7_U441  ( .A(_u10_u7_n2601 ), .ZN(_u10_u7_n2590 ) );
NAND2_X1 _u10_u7_U440  ( .A1(_u10_u7_n2599 ), .A2(_u10_u7_n2600 ), .ZN(_u10_u7_n2597 ) );
NAND2_X1 _u10_u7_U439  ( .A1(_u10_u7_n2082 ), .A2(_u10_u7_n2101 ), .ZN(_u10_u7_n2598 ) );
AND2_X1 _u10_u7_U438  ( .A1(_u10_u7_n2597 ), .A2(_u10_u7_n2598 ), .ZN(_u10_u7_n2281 ) );
NAND3_X1 _u10_u7_U437  ( .A1(_u10_u7_n1969 ), .A2(_u10_u7_n2582 ), .A3(_u10_u7_n2281 ), .ZN(_u10_u7_n2073 ) );
INV_X1 _u10_u7_U436  ( .A(_u10_u7_n2073 ), .ZN(_u10_u7_n2591 ) );
NOR2_X1 _u10_u7_U435  ( .A1(_u10_u7_n1816 ), .A2(_u10_u7_n2077 ), .ZN(_u10_u7_n2595 ) );
NOR2_X1 _u10_u7_U434  ( .A1(_u10_u7_n2595 ), .A2(_u10_u7_n2596 ), .ZN(_u10_u7_n2592 ) );
NAND3_X1 _u10_u7_U433  ( .A1(_u10_u7_n2107 ), .A2(_u10_u7_n2536 ), .A3(1'b0),.ZN(_u10_u7_n2438 ) );
INV_X1 _u10_u7_U432  ( .A(_u10_u7_n2438 ), .ZN(_u10_u7_n2427 ) );
NOR4_X1 _u10_u7_U431  ( .A1(1'b0), .A2(_u10_u7_n2594 ), .A3(_u10_u7_n2577 ),.A4(_u10_u7_n2427 ), .ZN(_u10_u7_n2593 ) );
NAND4_X1 _u10_u7_U430  ( .A1(_u10_u7_n2590 ), .A2(_u10_u7_n2591 ), .A3(_u10_u7_n2592 ), .A4(_u10_u7_n2593 ), .ZN(_u10_u7_n2589 ) );
NAND2_X1 _u10_u7_U429  ( .A1(_u10_u7_n2279 ), .A2(_u10_u7_n2589 ), .ZN(_u10_u7_n2558 ) );
NAND3_X1 _u10_u7_U428  ( .A1(_u10_u7_n2587 ), .A2(_u10_u7_n2115 ), .A3(_u10_u7_n2588 ), .ZN(_u10_u7_n2585 ) );
NOR4_X1 _u10_u7_U427  ( .A1(_u10_u7_n2585 ), .A2(_u10_u7_n2586 ), .A3(1'b0),.A4(_u10_u7_n2114 ), .ZN(_u10_u7_n2583 ) );
NOR2_X1 _u10_u7_U426  ( .A1(_u10_u7_n2583 ), .A2(_u10_u7_n2584 ), .ZN(_u10_u7_n2560 ) );
OR2_X1 _u10_u7_U425  ( .A1(_u10_u7_n2582 ), .A2(1'b0), .ZN(_u10_u7_n2581 ));
NAND2_X1 _u10_u7_U424  ( .A1(_u10_u7_n2580 ), .A2(_u10_u7_n2581 ), .ZN(_u10_u7_n1974 ) );
INV_X1 _u10_u7_U423  ( .A(_u10_u7_n1974 ), .ZN(_u10_u7_n1901 ) );
AND4_X1 _u10_u7_U422  ( .A1(_u10_u7_n1901 ), .A2(_u10_u7_n2385 ), .A3(_u10_u7_n2578 ), .A4(_u10_u7_n2579 ), .ZN(_u10_u7_n2424 ) );
NOR2_X1 _u10_u7_U421  ( .A1(1'b0), .A2(_u10_u7_n2424 ), .ZN(_u10_u7_n2574 ));
NOR3_X1 _u10_u7_U420  ( .A1(_u10_u7_n2427 ), .A2(1'b0), .A3(_u10_u7_n2577 ),.ZN(_u10_u7_n2576 ) );
NOR2_X1 _u10_u7_U419  ( .A1(_u10_u7_n2576 ), .A2(_u10_u7_n1976 ), .ZN(_u10_u7_n2575 ) );
NOR3_X1 _u10_u7_U418  ( .A1(_u10_u7_n2574 ), .A2(_u10_u7_n1979 ), .A3(_u10_u7_n2575 ), .ZN(_u10_u7_n2572 ) );
NOR2_X1 _u10_u7_U417  ( .A1(_u10_u7_n2572 ), .A2(_u10_u7_n2573 ), .ZN(_u10_u7_n2561 ) );
INV_X1 _u10_u7_U416  ( .A(_u10_u7_n2061 ), .ZN(_u10_u7_n2453 ) );
NOR2_X1 _u10_u7_U415  ( .A1(_u10_u7_n2453 ), .A2(_u10_u7_n1851 ), .ZN(_u10_u7_n2018 ) );
NAND2_X1 _u10_u7_U414  ( .A1(1'b0), .A2(_u10_u7_n2571 ), .ZN(_u10_u7_n2570 ));
NAND2_X1 _u10_u7_U413  ( .A1(_u10_u7_n2018 ), .A2(_u10_u7_n2570 ), .ZN(_u10_u7_n1837 ) );
INV_X1 _u10_u7_U412  ( .A(_u10_u7_n1837 ), .ZN(_u10_u7_n2568 ) );
NAND2_X1 _u10_u7_U411  ( .A1(1'b0), .A2(_u10_u7_n2536 ), .ZN(_u10_u7_n2569 ));
NAND2_X1 _u10_u7_U410  ( .A1(_u10_u7_n2568 ), .A2(_u10_u7_n2569 ), .ZN(_u10_u7_n2564 ) );
NOR2_X1 _u10_u7_U409  ( .A1(_u10_u7_n1841 ), .A2(_u10_u7_n1868 ), .ZN(_u10_u7_n2565 ) );
INV_X1 _u10_u7_U408  ( .A(_u10_u7_n2567 ), .ZN(_u10_u7_n2566 ) );
NOR4_X1 _u10_u7_U407  ( .A1(_u10_u7_n2564 ), .A2(_u10_u7_n2565 ), .A3(_u10_u7_n2143 ), .A4(_u10_u7_n2566 ), .ZN(_u10_u7_n2563 ) );
NOR2_X1 _u10_u7_U406  ( .A1(_u10_u7_n2563 ), .A2(_u10_u7_n2014 ), .ZN(_u10_u7_n2562 ) );
NOR3_X1 _u10_u7_U405  ( .A1(_u10_u7_n2560 ), .A2(_u10_u7_n2561 ), .A3(_u10_u7_n2562 ), .ZN(_u10_u7_n2559 ) );
NAND4_X1 _u10_u7_U404  ( .A1(_u10_u7_n2556 ), .A2(_u10_u7_n2557 ), .A3(_u10_u7_n2558 ), .A4(_u10_u7_n2559 ), .ZN(_u10_u7_n2511 ) );
INV_X1 _u10_u7_U403  ( .A(_u10_u7_n2085 ), .ZN(_u10_u7_n2293 ) );
NOR2_X1 _u10_u7_U402  ( .A1(_u10_u7_n2554 ), .A2(_u10_u7_n2555 ), .ZN(_u10_u7_n2444 ) );
NAND2_X1 _u10_u7_U401  ( .A1(_u10_u7_n2553 ), .A2(_u10_u7_n2549 ), .ZN(_u10_u7_n2552 ) );
AND2_X1 _u10_u7_U400  ( .A1(_u10_u7_n2444 ), .A2(_u10_u7_n2552 ), .ZN(_u10_u7_n2295 ) );
NAND2_X1 _u10_u7_U399  ( .A1(_u10_u7_n2551 ), .A2(_u10_u7_n2549 ), .ZN(_u10_u7_n2538 ) );
AND2_X1 _u10_u7_U398  ( .A1(_u10_u7_n2427 ), .A2(_u10_u7_n2108 ), .ZN(_u10_u7_n2460 ) );
NOR4_X1 _u10_u7_U397  ( .A1(_u10_u7_n2460 ), .A2(_u10_u7_n2306 ), .A3(_u10_u7_n2094 ), .A4(_u10_u7_n2550 ), .ZN(_u10_u7_n2409 ) );
INV_X1 _u10_u7_U396  ( .A(_u10_u7_n2409 ), .ZN(_u10_u7_n2407 ) );
NAND2_X1 _u10_u7_U395  ( .A1(_u10_u7_n2549 ), .A2(_u10_u7_n2407 ), .ZN(_u10_u7_n2546 ) );
NAND3_X1 _u10_u7_U394  ( .A1(_u10_u7_n2546 ), .A2(_u10_u7_n2547 ), .A3(_u10_u7_n2548 ), .ZN(_u10_u7_n2501 ) );
INV_X1 _u10_u7_U393  ( .A(_u10_u7_n2501 ), .ZN(_u10_u7_n2539 ) );
NOR2_X1 _u10_u7_U392  ( .A1(1'b0), .A2(_u10_u7_n2545 ), .ZN(_u10_u7_n2541 ));
AND2_X1 _u10_u7_U391  ( .A1(_u10_u7_n2544 ), .A2(_u10_u7_n2089 ), .ZN(_u10_u7_n2543 ) );
NOR3_X1 _u10_u7_U390  ( .A1(_u10_u7_n2541 ), .A2(_u10_u7_n2542 ), .A3(_u10_u7_n2543 ), .ZN(_u10_u7_n2540 ) );
NAND4_X1 _u10_u7_U389  ( .A1(_u10_u7_n2295 ), .A2(_u10_u7_n2538 ), .A3(_u10_u7_n2539 ), .A4(_u10_u7_n2540 ), .ZN(_u10_u7_n2537 ) );
NAND2_X1 _u10_u7_U388  ( .A1(_u10_u7_n2293 ), .A2(_u10_u7_n2537 ), .ZN(_u10_u7_n2515 ) );
NAND2_X1 _u10_u7_U387  ( .A1(_u10_u7_n2536 ), .A2(_u10_u7_n2508 ), .ZN(_u10_u7_n2526 ) );
NAND2_X1 _u10_u7_U386  ( .A1(_u10_u7_n2535 ), .A2(_u10_u7_n1940 ), .ZN(_u10_u7_n2532 ) );
NOR4_X1 _u10_u7_U385  ( .A1(_u10_u7_n2532 ), .A2(_u10_u7_n2533 ), .A3(1'b0),.A4(_u10_u7_n2534 ), .ZN(_u10_u7_n2530 ) );
NOR2_X1 _u10_u7_U384  ( .A1(_u10_u7_n2530 ), .A2(_u10_u7_n2531 ), .ZN(_u10_u7_n2529 ) );
NOR4_X1 _u10_u7_U383  ( .A1(_u10_u7_n2528 ), .A2(_u10_u7_n2143 ), .A3(_u10_u7_n2189 ), .A4(_u10_u7_n2529 ), .ZN(_u10_u7_n2527 ) );
NAND4_X1 _u10_u7_U382  ( .A1(_u10_u7_n2019 ), .A2(_u10_u7_n2526 ), .A3(_u10_u7_n2018 ), .A4(_u10_u7_n2527 ), .ZN(_u10_u7_n2525 ) );
NAND2_X1 _u10_u7_U381  ( .A1(_u10_u7_n2183 ), .A2(_u10_u7_n2525 ), .ZN(_u10_u7_n2516 ) );
INV_X1 _u10_u7_U380  ( .A(_u10_u7_n2524 ), .ZN(_u10_u7_n2396 ) );
NAND2_X1 _u10_u7_U379  ( .A1(_u10_u7_n2396 ), .A2(_u10_u7_n2523 ), .ZN(_u10_u7_n2522 ) );
NAND2_X1 _u10_u7_U378  ( .A1(_u10_u7_n1866 ), .A2(_u10_u7_n2522 ), .ZN(_u10_u7_n2519 ) );
AND2_X1 _u10_u7_U377  ( .A1(_u10_u7_n2493 ), .A2(_u10_u7_n1961 ), .ZN(_u10_u7_n2429 ) );
NAND2_X1 _u10_u7_U376  ( .A1(_u10_u7_n2429 ), .A2(_u10_u7_n2175 ), .ZN(_u10_u7_n2510 ) );
NAND2_X1 _u10_u7_U375  ( .A1(_u10_u7_n2510 ), .A2(_u10_u7_n1864 ), .ZN(_u10_u7_n2521 ) );
NAND3_X1 _u10_u7_U374  ( .A1(_u10_u7_n2519 ), .A2(_u10_u7_n2520 ), .A3(_u10_u7_n2521 ), .ZN(_u10_u7_n2518 ) );
NAND2_X1 _u10_u7_U373  ( .A1(_u10_u7_n1861 ), .A2(_u10_u7_n2518 ), .ZN(_u10_u7_n2517 ) );
NAND3_X1 _u10_u7_U372  ( .A1(_u10_u7_n2515 ), .A2(_u10_u7_n2516 ), .A3(_u10_u7_n2517 ), .ZN(_u10_u7_n2512 ) );
NOR2_X1 _u10_u7_U371  ( .A1(_u10_u7_n1913 ), .A2(_u10_u7_n1940 ), .ZN(_u10_u7_n2513 ) );
NOR2_X1 _u10_u7_U370  ( .A1(_u10_u7_n2113 ), .A2(_u10_u7_n2350 ), .ZN(_u10_u7_n2514 ) );
NOR4_X1 _u10_u7_U369  ( .A1(_u10_u7_n2511 ), .A2(_u10_u7_n2512 ), .A3(_u10_u7_n2513 ), .A4(_u10_u7_n2514 ), .ZN(_u10_u7_n2389 ) );
NAND2_X1 _u10_u7_U368  ( .A1(_u10_u7_n2509 ), .A2(_u10_u7_n2510 ), .ZN(_u10_u7_n2477 ) );
NAND2_X1 _u10_u7_U367  ( .A1(_u10_u7_n2507 ), .A2(_u10_u7_n2508 ), .ZN(_u10_u7_n2504 ) );
NAND2_X1 _u10_u7_U366  ( .A1(1'b0), .A2(_u10_u7_n2506 ), .ZN(_u10_u7_n2505 ));
NAND2_X1 _u10_u7_U365  ( .A1(_u10_u7_n2504 ), .A2(_u10_u7_n2505 ), .ZN(_u10_u7_n2503 ) );
NAND2_X1 _u10_u7_U364  ( .A1(_u10_u7_n2502 ), .A2(_u10_u7_n2503 ), .ZN(_u10_u7_n2478 ) );
NAND2_X1 _u10_u7_U363  ( .A1(_u10_u7_n2501 ), .A2(_u10_u7_n2446 ), .ZN(_u10_u7_n2497 ) );
INV_X1 _u10_u7_U362  ( .A(_u10_u7_n2500 ), .ZN(_u10_u7_n2499 ) );
NAND3_X1 _u10_u7_U361  ( .A1(_u10_u7_n2497 ), .A2(_u10_u7_n2498 ), .A3(_u10_u7_n2499 ), .ZN(_u10_u7_n2496 ) );
NAND2_X1 _u10_u7_U360  ( .A1(_u10_u7_n2445 ), .A2(_u10_u7_n2496 ), .ZN(_u10_u7_n2479 ) );
NOR2_X1 _u10_u7_U359  ( .A1(_u10_u7_n2429 ), .A2(_u10_u7_n2495 ), .ZN(_u10_u7_n2491 ) );
INV_X1 _u10_u7_U358  ( .A(_u10_u7_n2191 ), .ZN(_u10_u7_n2494 ) );
NOR2_X1 _u10_u7_U357  ( .A1(_u10_u7_n2493 ), .A2(_u10_u7_n2494 ), .ZN(_u10_u7_n2492 ) );
NOR2_X1 _u10_u7_U356  ( .A1(_u10_u7_n2491 ), .A2(_u10_u7_n2492 ), .ZN(_u10_u7_n2489 ) );
NOR2_X1 _u10_u7_U355  ( .A1(_u10_u7_n2489 ), .A2(_u10_u7_n2490 ), .ZN(_u10_u7_n2481 ) );
NAND2_X1 _u10_u7_U354  ( .A1(_u10_u7_n2253 ), .A2(_u10_u7_n1859 ), .ZN(_u10_u7_n2398 ) );
NOR2_X1 _u10_u7_U353  ( .A1(_u10_u7_n2488 ), .A2(_u10_u7_n2398 ), .ZN(_u10_u7_n2487 ) );
NOR2_X1 _u10_u7_U352  ( .A1(_u10_u7_n2220 ), .A2(_u10_u7_n2487 ), .ZN(_u10_u7_n2482 ) );
AND2_X1 _u10_u7_U351  ( .A1(_u10_u7_n2350 ), .A2(_u10_u7_n2486 ), .ZN(_u10_u7_n2484 ) );
NOR2_X1 _u10_u7_U350  ( .A1(_u10_u7_n2484 ), .A2(_u10_u7_n2485 ), .ZN(_u10_u7_n2483 ) );
NOR3_X1 _u10_u7_U349  ( .A1(_u10_u7_n2481 ), .A2(_u10_u7_n2482 ), .A3(_u10_u7_n2483 ), .ZN(_u10_u7_n2480 ) );
NAND4_X1 _u10_u7_U348  ( .A1(_u10_u7_n2477 ), .A2(_u10_u7_n2478 ), .A3(_u10_u7_n2479 ), .A4(_u10_u7_n2480 ), .ZN(_u10_u7_n2447 ) );
NAND2_X1 _u10_u7_U347  ( .A1(_u10_u7_n2476 ), .A2(_u10_u7_n1936 ), .ZN(_u10_u7_n2472 ) );
NAND2_X1 _u10_u7_U346  ( .A1(_u10_u7_n2427 ), .A2(_u10_u7_n2278 ), .ZN(_u10_u7_n2473 ) );
NAND4_X1 _u10_u7_U345  ( .A1(_u10_u7_n2472 ), .A2(_u10_u7_n2473 ), .A3(_u10_u7_n2474 ), .A4(_u10_u7_n2475 ), .ZN(_u10_u7_n2471 ) );
NAND2_X1 _u10_u7_U344  ( .A1(_u10_u7_n2470 ), .A2(_u10_u7_n2471 ), .ZN(_u10_u7_n2457 ) );
NAND2_X1 _u10_u7_U343  ( .A1(_u10_u7_n2409 ), .A2(_u10_u7_n2469 ), .ZN(_u10_u7_n2468 ) );
NAND2_X1 _u10_u7_U342  ( .A1(_u10_u7_n2467 ), .A2(_u10_u7_n2468 ), .ZN(_u10_u7_n2463 ) );
NAND2_X1 _u10_u7_U341  ( .A1(_u10_u7_n1844 ), .A2(_u10_u7_n2466 ), .ZN(_u10_u7_n2465 ) );
NAND3_X1 _u10_u7_U340  ( .A1(_u10_u7_n2463 ), .A2(_u10_u7_n2464 ), .A3(_u10_u7_n2465 ), .ZN(_u10_u7_n2462 ) );
NAND2_X1 _u10_u7_U339  ( .A1(_u10_u7_n2461 ), .A2(_u10_u7_n2462 ), .ZN(_u10_u7_n2458 ) );
NAND2_X1 _u10_u7_U338  ( .A1(_u10_u7_n2460 ), .A2(_u10_u7_n2251 ), .ZN(_u10_u7_n2459 ) );
NAND3_X1 _u10_u7_U337  ( .A1(_u10_u7_n2457 ), .A2(_u10_u7_n2458 ), .A3(_u10_u7_n2459 ), .ZN(_u10_u7_n2448 ) );
NOR2_X1 _u10_u7_U336  ( .A1(_u10_u7_n2455 ), .A2(_u10_u7_n2456 ), .ZN(_u10_u7_n2449 ) );
NAND2_X1 _u10_u7_U335  ( .A1(_u10_u7_n2454 ), .A2(_u10_u7_n2438 ), .ZN(_u10_u7_n2452 ) );
NOR4_X1 _u10_u7_U334  ( .A1(_u10_u7_n2452 ), .A2(_u10_u7_n2453 ), .A3(_u10_u7_n2443 ), .A4(_u10_u7_n2143 ), .ZN(_u10_u7_n2451 ) );
NOR2_X1 _u10_u7_U333  ( .A1(_u10_u7_n2451 ), .A2(_u10_u7_n2356 ), .ZN(_u10_u7_n2450 ) );
NOR4_X1 _u10_u7_U332  ( .A1(_u10_u7_n2447 ), .A2(_u10_u7_n2448 ), .A3(_u10_u7_n2449 ), .A4(_u10_u7_n2450 ), .ZN(_u10_u7_n2390 ) );
NAND2_X1 _u10_u7_U331  ( .A1(_u10_u7_n2445 ), .A2(_u10_u7_n2446 ), .ZN(_u10_u7_n2155 ) );
INV_X1 _u10_u7_U330  ( .A(_u10_u7_n2155 ), .ZN(_u10_u7_n1892 ) );
INV_X1 _u10_u7_U329  ( .A(_u10_u7_n2444 ), .ZN(_u10_u7_n2088 ) );
NAND2_X1 _u10_u7_U328  ( .A1(_u10_u7_n1892 ), .A2(_u10_u7_n2088 ), .ZN(_u10_u7_n2337 ) );
NOR3_X1 _u10_u7_U327  ( .A1(_u10_u7_n2441 ), .A2(_u10_u7_n2442 ), .A3(_u10_u7_n2443 ), .ZN(_u10_u7_n2440 ) );
NAND4_X1 _u10_u7_U326  ( .A1(_u10_u7_n2193 ), .A2(_u10_u7_n2355 ), .A3(_u10_u7_n2439 ), .A4(_u10_u7_n2440 ), .ZN(_u10_u7_n2434 ) );
NAND3_X1 _u10_u7_U325  ( .A1(_u10_u7_n2437 ), .A2(_u10_u7_n2438 ), .A3(_u10_u7_n2059 ), .ZN(_u10_u7_n2435 ) );
NOR4_X1 _u10_u7_U324  ( .A1(_u10_u7_n2434 ), .A2(_u10_u7_n2435 ), .A3(_u10_u7_n1837 ), .A4(_u10_u7_n2436 ), .ZN(_u10_u7_n2433 ) );
NOR2_X1 _u10_u7_U323  ( .A1(_u10_u7_n2433 ), .A2(_u10_u7_n1836 ), .ZN(_u10_u7_n2415 ) );
INV_X1 _u10_u7_U322  ( .A(_u10_u7_n2432 ), .ZN(_u10_u7_n2178 ) );
NOR2_X1 _u10_u7_U321  ( .A1(_u10_u7_n1960 ), .A2(_u10_u7_n2431 ), .ZN(_u10_u7_n2430 ) );
NOR4_X1 _u10_u7_U320  ( .A1(_u10_u7_n2178 ), .A2(_u10_u7_n2429 ), .A3(_u10_u7_n2430 ), .A4(_u10_u7_n2179 ), .ZN(_u10_u7_n2416 ) );
NOR2_X1 _u10_u7_U319  ( .A1(_u10_u7_n2427 ), .A2(_u10_u7_n2428 ), .ZN(_u10_u7_n2426 ) );
NAND4_X1 _u10_u7_U318  ( .A1(_u10_u7_n2286 ), .A2(_u10_u7_n1969 ), .A3(_u10_u7_n2282 ), .A4(_u10_u7_n2426 ), .ZN(_u10_u7_n2425 ) );
NAND2_X1 _u10_u7_U317  ( .A1(_u10_u7_n2031 ), .A2(_u10_u7_n2425 ), .ZN(_u10_u7_n2422 ) );
NAND3_X1 _u10_u7_U316  ( .A1(_u10_u7_n2422 ), .A2(_u10_u7_n2423 ), .A3(_u10_u7_n2424 ), .ZN(_u10_u7_n2419 ) );
NOR4_X1 _u10_u7_U315  ( .A1(_u10_u7_n2419 ), .A2(_u10_u7_n1978 ), .A3(_u10_u7_n2420 ), .A4(_u10_u7_n2421 ), .ZN(_u10_u7_n2418 ) );
NOR2_X1 _u10_u7_U314  ( .A1(_u10_u7_n2418 ), .A2(_u10_u7_n2359 ), .ZN(_u10_u7_n2417 ) );
NOR3_X1 _u10_u7_U313  ( .A1(_u10_u7_n2415 ), .A2(_u10_u7_n2416 ), .A3(_u10_u7_n2417 ), .ZN(_u10_u7_n2414 ) );
NAND4_X1 _u10_u7_U312  ( .A1(_u10_u7_n2337 ), .A2(_u10_u7_n2412 ), .A3(_u10_u7_n2413 ), .A4(_u10_u7_n2414 ), .ZN(_u10_u7_n2392 ) );
NAND2_X1 _u10_u7_U311  ( .A1(_u10_u7_n2411 ), .A2(_u10_u7_n1936 ), .ZN(_u10_u7_n2410 ) );
NAND2_X1 _u10_u7_U310  ( .A1(_u10_u7_n2409 ), .A2(_u10_u7_n2410 ), .ZN(_u10_u7_n2408 ) );
NAND3_X1 _u10_u7_U309  ( .A1(_u10_u7_n2408 ), .A2(_u10_u7_n2305 ), .A3(_u10_u7_n1894 ), .ZN(_u10_u7_n2402 ) );
NAND3_X1 _u10_u7_U308  ( .A1(_u10_u7_n2329 ), .A2(_u10_u7_n2407 ), .A3(_u10_u7_n2255 ), .ZN(_u10_u7_n2403 ) );
NAND3_X1 _u10_u7_U307  ( .A1(_u10_u7_n1924 ), .A2(_u10_u7_n2405 ), .A3(_u10_u7_n2406 ), .ZN(_u10_u7_n2404 ) );
NAND3_X1 _u10_u7_U306  ( .A1(_u10_u7_n2402 ), .A2(_u10_u7_n2403 ), .A3(_u10_u7_n2404 ), .ZN(_u10_u7_n2393 ) );
INV_X1 _u10_u7_U305  ( .A(_u10_u7_n1932 ), .ZN(_u10_u7_n2399 ) );
NOR2_X1 _u10_u7_U304  ( .A1(_u10_u7_n2401 ), .A2(_u10_u7_n2161 ), .ZN(_u10_u7_n2400 ) );
NOR2_X1 _u10_u7_U303  ( .A1(_u10_u7_n2399 ), .A2(_u10_u7_n2400 ), .ZN(_u10_u7_n2394 ) );
NOR2_X1 _u10_u7_U302  ( .A1(_u10_u7_n2110 ), .A2(_u10_u7_n2398 ), .ZN(_u10_u7_n2397 ) );
NOR2_X1 _u10_u7_U301  ( .A1(_u10_u7_n2396 ), .A2(_u10_u7_n2397 ), .ZN(_u10_u7_n2395 ) );
NOR4_X1 _u10_u7_U300  ( .A1(_u10_u7_n2392 ), .A2(_u10_u7_n2393 ), .A3(_u10_u7_n2394 ), .A4(_u10_u7_n2395 ), .ZN(_u10_u7_n2391 ) );
NAND4_X1 _u10_u7_U299  ( .A1(_u10_u7_n2388 ), .A2(_u10_u7_n2389 ), .A3(_u10_u7_n2390 ), .A4(_u10_u7_n2391 ), .ZN(_u10_u7_n2387 ) );
MUX2_X1 _u10_u7_U298  ( .A(_u10_u7_n2387 ), .B(_u10_SYNOPSYS_UNCONNECTED_30 ), .S(_u10_u7_n1819 ), .Z(_u10_u7_n1810 ) );
NAND2_X1 _u10_u7_U297  ( .A1(_u10_u7_n2386 ), .A2(_u10_u7_n2007 ), .ZN(_u10_u7_n2369 ) );
AND2_X1 _u10_u7_U296  ( .A1(1'b0), .A2(_u10_u7_n2195 ), .ZN(_u10_u7_n2308 ));
NAND2_X1 _u10_u7_U295  ( .A1(_u10_u7_n2308 ), .A2(_u10_u7_n2036 ), .ZN(_u10_u7_n2384 ) );
AND2_X1 _u10_u7_U294  ( .A1(_u10_u7_n2384 ), .A2(_u10_u7_n2385 ), .ZN(_u10_u7_n2275 ) );
AND4_X1 _u10_u7_U293  ( .A1(_u10_u7_n2275 ), .A2(_u10_u7_n2286 ), .A3(_u10_u7_n2383 ), .A4(_u10_u7_n2285 ), .ZN(_u10_u7_n2225 ) );
NAND3_X1 _u10_u7_U292  ( .A1(_u10_u7_n2195 ), .A2(_u10_u7_n2223 ), .A3(1'b0),.ZN(_u10_u7_n2021 ) );
INV_X1 _u10_u7_U291  ( .A(_u10_u7_n2021 ), .ZN(_u10_u7_n2167 ) );
NAND2_X1 _u10_u7_U290  ( .A1(_u10_u7_n2036 ), .A2(_u10_u7_n2167 ), .ZN(_u10_u7_n1970 ) );
AND3_X1 _u10_u7_U289  ( .A1(_u10_u7_n1970 ), .A2(_u10_u7_n2164 ), .A3(_u10_u7_n2382 ), .ZN(_u10_u7_n2381 ) );
NAND4_X1 _u10_u7_U288  ( .A1(_u10_u7_n2225 ), .A2(_u10_u7_n2379 ), .A3(_u10_u7_n2380 ), .A4(_u10_u7_n2381 ), .ZN(_u10_u7_n2378 ) );
NAND2_X1 _u10_u7_U287  ( .A1(_u10_u7_n1967 ), .A2(_u10_u7_n2378 ), .ZN(_u10_u7_n2370 ) );
NAND2_X1 _u10_u7_U286  ( .A1(_u10_u7_n2081 ), .A2(_u10_u7_n2377 ), .ZN(_u10_u7_n2371 ) );
NOR2_X1 _u10_u7_U285  ( .A1(_u10_u7_n2375 ), .A2(_u10_u7_n2376 ), .ZN(_u10_u7_n2373 ) );
NOR2_X1 _u10_u7_U284  ( .A1(_u10_u7_n2373 ), .A2(_u10_u7_n2374 ), .ZN(_u10_u7_n2372 ) );
NAND4_X1 _u10_u7_U283  ( .A1(_u10_u7_n2369 ), .A2(_u10_u7_n2370 ), .A3(_u10_u7_n2371 ), .A4(_u10_u7_n2372 ), .ZN(_u10_u7_n2309 ) );
NOR2_X1 _u10_u7_U282  ( .A1(_u10_u7_n2000 ), .A2(_u10_u7_n2368 ), .ZN(_u10_u7_n2360 ) );
NOR2_X1 _u10_u7_U281  ( .A1(_u10_u7_n2366 ), .A2(_u10_u7_n2367 ), .ZN(_u10_u7_n2361 ) );
NOR2_X1 _u10_u7_U280  ( .A1(_u10_u7_n1868 ), .A2(_u10_u7_n2365 ), .ZN(_u10_u7_n2362 ) );
NOR2_X1 _u10_u7_U279  ( .A1(_u10_u7_n2364 ), .A2(_u10_u7_n1859 ), .ZN(_u10_u7_n2363 ) );
NOR4_X1 _u10_u7_U278  ( .A1(_u10_u7_n2360 ), .A2(_u10_u7_n2361 ), .A3(_u10_u7_n2362 ), .A4(_u10_u7_n2363 ), .ZN(_u10_u7_n2316 ) );
NOR2_X1 _u10_u7_U277  ( .A1(_u10_u7_n2359 ), .A2(_u10_u7_n1970 ), .ZN(_u10_u7_n2351 ) );
NOR2_X1 _u10_u7_U276  ( .A1(_u10_u7_n2358 ), .A2(_u10_u7_n1840 ), .ZN(_u10_u7_n2352 ) );
NOR2_X1 _u10_u7_U275  ( .A1(_u10_u7_n2356 ), .A2(_u10_u7_n2357 ), .ZN(_u10_u7_n2353 ) );
NOR2_X1 _u10_u7_U274  ( .A1(_u10_u7_n1836 ), .A2(_u10_u7_n2355 ), .ZN(_u10_u7_n2354 ) );
NOR4_X1 _u10_u7_U273  ( .A1(_u10_u7_n2351 ), .A2(_u10_u7_n2352 ), .A3(_u10_u7_n2353 ), .A4(_u10_u7_n2354 ), .ZN(_u10_u7_n2317 ) );
NOR2_X1 _u10_u7_U272  ( .A1(_u10_u7_n1873 ), .A2(_u10_u7_n2101 ), .ZN(_u10_u7_n2349 ) );
NOR2_X1 _u10_u7_U271  ( .A1(_u10_u7_n2349 ), .A2(_u10_u7_n2350 ), .ZN(_u10_u7_n2338 ) );
NOR2_X1 _u10_u7_U270  ( .A1(_u10_u7_n2347 ), .A2(_u10_u7_n2348 ), .ZN(_u10_u7_n2345 ) );
NOR2_X1 _u10_u7_U269  ( .A1(_u10_u7_n2345 ), .A2(_u10_u7_n2346 ), .ZN(_u10_u7_n2339 ) );
NOR2_X1 _u10_u7_U268  ( .A1(_u10_u7_n2344 ), .A2(_u10_u7_n2142 ), .ZN(_u10_u7_n2340 ) );
NOR2_X1 _u10_u7_U267  ( .A1(_u10_u7_n2342 ), .A2(_u10_u7_n2343 ), .ZN(_u10_u7_n2341 ) );
NOR4_X1 _u10_u7_U266  ( .A1(_u10_u7_n2338 ), .A2(_u10_u7_n2339 ), .A3(_u10_u7_n2340 ), .A4(_u10_u7_n2341 ), .ZN(_u10_u7_n2318 ) );
INV_X1 _u10_u7_U265  ( .A(_u10_u7_n2337 ), .ZN(_u10_u7_n2320 ) );
NOR2_X1 _u10_u7_U264  ( .A1(_u10_u7_n1970 ), .A2(1'b0), .ZN(_u10_u7_n2027 ));
INV_X1 _u10_u7_U263  ( .A(_u10_u7_n2027 ), .ZN(_u10_u7_n2331 ) );
NOR2_X1 _u10_u7_U262  ( .A1(_u10_u7_n2174 ), .A2(_u10_u7_n2216 ), .ZN(_u10_u7_n2333 ) );
AND2_X1 _u10_u7_U261  ( .A1(_u10_u7_n1928 ), .A2(_u10_u7_n2336 ), .ZN(_u10_u7_n2334 ) );
NOR4_X1 _u10_u7_U260  ( .A1(_u10_u7_n1937 ), .A2(_u10_u7_n2333 ), .A3(_u10_u7_n2334 ), .A4(_u10_u7_n2335 ), .ZN(_u10_u7_n2332 ) );
NOR3_X1 _u10_u7_U259  ( .A1(_u10_u7_n2331 ), .A2(_u10_u7_n2332 ), .A3(_u10_u7_n1915 ), .ZN(_u10_u7_n2321 ) );
NOR3_X1 _u10_u7_U258  ( .A1(_u10_u7_n2291 ), .A2(_u10_u7_n2330 ), .A3(_u10_u7_n2021 ), .ZN(_u10_u7_n2322 ) );
NOR2_X1 _u10_u7_U257  ( .A1(_u10_u7_n2329 ), .A2(_u10_u7_n2169 ), .ZN(_u10_u7_n2324 ) );
NOR2_X1 _u10_u7_U256  ( .A1(1'b0), .A2(_u10_u7_n2328 ), .ZN(_u10_u7_n2327 ));
NOR2_X1 _u10_u7_U255  ( .A1(_u10_u7_n2326 ), .A2(_u10_u7_n2327 ), .ZN(_u10_u7_n2325 ) );
NOR3_X1 _u10_u7_U254  ( .A1(_u10_u7_n2324 ), .A2(1'b0), .A3(_u10_u7_n2325 ),.ZN(_u10_u7_n2323 ) );
NOR4_X1 _u10_u7_U253  ( .A1(_u10_u7_n2320 ), .A2(_u10_u7_n2321 ), .A3(_u10_u7_n2322 ), .A4(_u10_u7_n2323 ), .ZN(_u10_u7_n2319 ) );
AND4_X1 _u10_u7_U252  ( .A1(_u10_u7_n2316 ), .A2(_u10_u7_n2317 ), .A3(_u10_u7_n2318 ), .A4(_u10_u7_n2319 ), .ZN(_u10_u7_n1991 ) );
INV_X1 _u10_u7_U251  ( .A(_u10_u7_n2315 ), .ZN(_u10_u7_n2313 ) );
NAND3_X1 _u10_u7_U250  ( .A1(_u10_u7_n1991 ), .A2(_u10_u7_n2313 ), .A3(_u10_u7_n2314 ), .ZN(_u10_u7_n2310 ) );
NOR4_X1 _u10_u7_U249  ( .A1(_u10_u7_n2309 ), .A2(_u10_u7_n2310 ), .A3(_u10_u7_n2311 ), .A4(_u10_u7_n2312 ), .ZN(_u10_u7_n2117 ) );
NAND3_X1 _u10_u7_U248  ( .A1(_u10_u7_n2108 ), .A2(_u10_u7_n2107 ), .A3(_u10_u7_n2308 ), .ZN(_u10_u7_n2217 ) );
NOR3_X1 _u10_u7_U247  ( .A1(_u10_u7_n2306 ), .A2(_u10_u7_n2307 ), .A3(_u10_u7_n2027 ), .ZN(_u10_u7_n2277 ) );
NAND3_X1 _u10_u7_U246  ( .A1(_u10_u7_n2217 ), .A2(_u10_u7_n2305 ), .A3(_u10_u7_n2277 ), .ZN(_u10_u7_n2157 ) );
NAND2_X1 _u10_u7_U245  ( .A1(_u10_u7_n2089 ), .A2(_u10_u7_n2157 ), .ZN(_u10_u7_n2296 ) );
INV_X1 _u10_u7_U244  ( .A(_u10_u7_n2304 ), .ZN(_u10_u7_n2297 ) );
NOR2_X1 _u10_u7_U243  ( .A1(_u10_u7_n2302 ), .A2(_u10_u7_n2303 ), .ZN(_u10_u7_n2299 ) );
NOR3_X1 _u10_u7_U242  ( .A1(_u10_u7_n2299 ), .A2(_u10_u7_n2300 ), .A3(_u10_u7_n2301 ), .ZN(_u10_u7_n2298 ) );
NAND4_X1 _u10_u7_U241  ( .A1(_u10_u7_n2295 ), .A2(_u10_u7_n2296 ), .A3(_u10_u7_n2297 ), .A4(_u10_u7_n2298 ), .ZN(_u10_u7_n2294 ) );
NAND2_X1 _u10_u7_U240  ( .A1(_u10_u7_n2293 ), .A2(_u10_u7_n2294 ), .ZN(_u10_u7_n2257 ) );
NAND2_X1 _u10_u7_U239  ( .A1(_u10_u7_n2165 ), .A2(_u10_u7_n2166 ), .ZN(_u10_u7_n2288 ) );
NAND2_X1 _u10_u7_U238  ( .A1(_u10_u7_n2078 ), .A2(_u10_u7_n2279 ), .ZN(_u10_u7_n2292 ) );
NAND2_X1 _u10_u7_U237  ( .A1(_u10_u7_n2291 ), .A2(_u10_u7_n2292 ), .ZN(_u10_u7_n2290 ) );
NAND2_X1 _u10_u7_U236  ( .A1(_u10_u7_n2059 ), .A2(_u10_u7_n2290 ), .ZN(_u10_u7_n2289 ) );
NAND2_X1 _u10_u7_U235  ( .A1(_u10_u7_n2288 ), .A2(_u10_u7_n2289 ), .ZN(_u10_u7_n2201 ) );
NAND2_X1 _u10_u7_U234  ( .A1(1'b0), .A2(_u10_u7_n2201 ), .ZN(_u10_u7_n2258 ));
INV_X1 _u10_u7_U233  ( .A(_u10_u7_n2287 ), .ZN(_u10_u7_n2283 ) );
AND4_X1 _u10_u7_U232  ( .A1(_u10_u7_n2285 ), .A2(_u10_u7_n2226 ), .A3(_u10_u7_n1970 ), .A4(_u10_u7_n2286 ), .ZN(_u10_u7_n2284 ) );
NAND4_X1 _u10_u7_U231  ( .A1(_u10_u7_n2281 ), .A2(_u10_u7_n2282 ), .A3(_u10_u7_n2283 ), .A4(_u10_u7_n2284 ), .ZN(_u10_u7_n2280 ) );
NAND2_X1 _u10_u7_U230  ( .A1(_u10_u7_n2279 ), .A2(_u10_u7_n2280 ), .ZN(_u10_u7_n2259 ) );
NAND4_X1 _u10_u7_U229  ( .A1(_u10_u7_n2275 ), .A2(_u10_u7_n2276 ), .A3(_u10_u7_n2277 ), .A4(_u10_u7_n2278 ), .ZN(_u10_u7_n2271 ) );
NAND2_X1 _u10_u7_U228  ( .A1(_u10_u7_n1933 ), .A2(_u10_u7_n2164 ), .ZN(_u10_u7_n2272 ) );
NOR2_X1 _u10_u7_U227  ( .A1(_u10_u7_n2274 ), .A2(_u10_u7_n2130 ), .ZN(_u10_u7_n2273 ) );
NOR4_X1 _u10_u7_U226  ( .A1(_u10_u7_n2271 ), .A2(_u10_u7_n2272 ), .A3(_u10_u7_n1978 ), .A4(_u10_u7_n2273 ), .ZN(_u10_u7_n2270 ) );
NOR2_X1 _u10_u7_U225  ( .A1(_u10_u7_n2270 ), .A2(_u10_u7_n2025 ), .ZN(_u10_u7_n2261 ) );
NAND3_X1 _u10_u7_U224  ( .A1(_u10_u7_n1933 ), .A2(_u10_u7_n1936 ), .A3(_u10_u7_n2269 ), .ZN(_u10_u7_n2268 ) );
NOR3_X1 _u10_u7_U223  ( .A1(_u10_u7_n2268 ), .A2(_u10_u7_n1844 ), .A3(_u10_u7_n2157 ), .ZN(_u10_u7_n2267 ) );
NOR2_X1 _u10_u7_U222  ( .A1(1'b0), .A2(_u10_u7_n2267 ), .ZN(_u10_u7_n2265 ));
NOR3_X1 _u10_u7_U221  ( .A1(_u10_u7_n2264 ), .A2(_u10_u7_n2265 ), .A3(_u10_u7_n2266 ), .ZN(_u10_u7_n2263 ) );
NOR2_X1 _u10_u7_U220  ( .A1(_u10_u7_n2263 ), .A2(_u10_u7_n1843 ), .ZN(_u10_u7_n2262 ) );
NOR2_X1 _u10_u7_U219  ( .A1(_u10_u7_n2261 ), .A2(_u10_u7_n2262 ), .ZN(_u10_u7_n2260 ) );
NAND4_X1 _u10_u7_U218  ( .A1(_u10_u7_n2257 ), .A2(_u10_u7_n2258 ), .A3(_u10_u7_n2259 ), .A4(_u10_u7_n2260 ), .ZN(_u10_u7_n2230 ) );
INV_X1 _u10_u7_U217  ( .A(_u10_u7_n2217 ), .ZN(_u10_u7_n2242 ) );
NAND2_X1 _u10_u7_U216  ( .A1(_u10_u7_n2168 ), .A2(_u10_u7_n2169 ), .ZN(_u10_u7_n2244 ) );
NAND2_X1 _u10_u7_U215  ( .A1(_u10_u7_n2255 ), .A2(_u10_u7_n2256 ), .ZN(_u10_u7_n2245 ) );
NAND2_X1 _u10_u7_U214  ( .A1(_u10_u7_n2253 ), .A2(_u10_u7_n2254 ), .ZN(_u10_u7_n2252 ) );
NAND2_X1 _u10_u7_U213  ( .A1(_u10_u7_n2251 ), .A2(_u10_u7_n2252 ), .ZN(_u10_u7_n2246 ) );
NAND2_X1 _u10_u7_U212  ( .A1(_u10_u7_n2152 ), .A2(_u10_u7_n1928 ), .ZN(_u10_u7_n2250 ) );
NAND2_X1 _u10_u7_U211  ( .A1(_u10_u7_n2249 ), .A2(_u10_u7_n2250 ), .ZN(_u10_u7_n2248 ) );
NAND2_X1 _u10_u7_U210  ( .A1(_u10_u7_n2105 ), .A2(_u10_u7_n2248 ), .ZN(_u10_u7_n2247 ) );
NAND4_X1 _u10_u7_U209  ( .A1(_u10_u7_n2244 ), .A2(_u10_u7_n2245 ), .A3(_u10_u7_n2246 ), .A4(_u10_u7_n2247 ), .ZN(_u10_u7_n2243 ) );
NAND2_X1 _u10_u7_U208  ( .A1(_u10_u7_n2242 ), .A2(_u10_u7_n2243 ), .ZN(_u10_u7_n2237 ) );
NAND2_X1 _u10_u7_U207  ( .A1(1'b0), .A2(_u10_u7_n2241 ), .ZN(_u10_u7_n2238 ));
NAND2_X1 _u10_u7_U206  ( .A1(_u10_u7_n2214 ), .A2(_u10_u7_n2240 ), .ZN(_u10_u7_n2239 ) );
NAND3_X1 _u10_u7_U205  ( .A1(_u10_u7_n2237 ), .A2(_u10_u7_n2238 ), .A3(_u10_u7_n2239 ), .ZN(_u10_u7_n2231 ) );
AND2_X1 _u10_u7_U204  ( .A1(_u10_u7_n2200 ), .A2(_u10_u7_n2236 ), .ZN(_u10_u7_n2232 ) );
NOR2_X1 _u10_u7_U203  ( .A1(_u10_u7_n2234 ), .A2(_u10_u7_n2235 ), .ZN(_u10_u7_n2233 ) );
NOR4_X1 _u10_u7_U202  ( .A1(_u10_u7_n2230 ), .A2(_u10_u7_n2231 ), .A3(_u10_u7_n2232 ), .A4(_u10_u7_n2233 ), .ZN(_u10_u7_n2118 ) );
NAND2_X1 _u10_u7_U201  ( .A1(_u10_u7_n2214 ), .A2(_u10_u7_n2049 ), .ZN(_u10_u7_n2229 ) );
NAND2_X1 _u10_u7_U200  ( .A1(_u10_u7_n2228 ), .A2(_u10_u7_n2229 ), .ZN(_u10_u7_n2227 ) );
NAND2_X1 _u10_u7_U199  ( .A1(_u10_u7_n2043 ), .A2(_u10_u7_n2227 ), .ZN(_u10_u7_n2204 ) );
NAND2_X1 _u10_u7_U198  ( .A1(_u10_u7_n2225 ), .A2(_u10_u7_n2226 ), .ZN(_u10_u7_n2224 ) );
NAND2_X1 _u10_u7_U197  ( .A1(_u10_u7_n1899 ), .A2(_u10_u7_n2224 ), .ZN(_u10_u7_n2205 ) );
NAND2_X1 _u10_u7_U196  ( .A1(_u10_u7_n2222 ), .A2(_u10_u7_n2223 ), .ZN(_u10_u7_n1870 ) );
NAND4_X1 _u10_u7_U195  ( .A1(_u10_u7_n2220 ), .A2(_u10_u7_n2131 ), .A3(_u10_u7_n2221 ), .A4(_u10_u7_n1870 ), .ZN(_u10_u7_n2219 ) );
NAND2_X1 _u10_u7_U194  ( .A1(_u10_u7_n2218 ), .A2(_u10_u7_n2219 ), .ZN(_u10_u7_n2206 ) );
NOR2_X1 _u10_u7_U193  ( .A1(_u10_u7_n1925 ), .A2(_u10_u7_n2217 ), .ZN(_u10_u7_n2215 ) );
NOR4_X1 _u10_u7_U192  ( .A1(_u10_u7_n2213 ), .A2(_u10_u7_n2214 ), .A3(_u10_u7_n2215 ), .A4(_u10_u7_n2216 ), .ZN(_u10_u7_n2211 ) );
NOR2_X1 _u10_u7_U191  ( .A1(_u10_u7_n2211 ), .A2(_u10_u7_n2212 ), .ZN(_u10_u7_n2208 ) );
NOR2_X1 _u10_u7_U190  ( .A1(_u10_u7_n1888 ), .A2(_u10_u7_n2210 ), .ZN(_u10_u7_n2209 ) );
NOR2_X1 _u10_u7_U189  ( .A1(_u10_u7_n2208 ), .A2(_u10_u7_n2209 ), .ZN(_u10_u7_n2207 ) );
NAND4_X1 _u10_u7_U188  ( .A1(_u10_u7_n2204 ), .A2(_u10_u7_n2205 ), .A3(_u10_u7_n2206 ), .A4(_u10_u7_n2207 ), .ZN(_u10_u7_n2170 ) );
OR2_X1 _u10_u7_U187  ( .A1(_u10_u7_n2202 ), .A2(_u10_u7_n2203 ), .ZN(_u10_u7_n2197 ) );
NAND2_X1 _u10_u7_U186  ( .A1(1'b0), .A2(_u10_u7_n2201 ), .ZN(_u10_u7_n2198 ));
NAND2_X1 _u10_u7_U185  ( .A1(_u10_u7_n2063 ), .A2(_u10_u7_n2200 ), .ZN(_u10_u7_n2199 ) );
NAND3_X1 _u10_u7_U184  ( .A1(_u10_u7_n2197 ), .A2(_u10_u7_n2198 ), .A3(_u10_u7_n2199 ), .ZN(_u10_u7_n2196 ) );
NAND2_X1 _u10_u7_U183  ( .A1(_u10_u7_n2195 ), .A2(_u10_u7_n2196 ), .ZN(_u10_u7_n2180 ) );
NAND2_X1 _u10_u7_U182  ( .A1(_u10_u7_n2195 ), .A2(_u10_u7_n1918 ), .ZN(_u10_u7_n2192 ) );
NAND4_X1 _u10_u7_U181  ( .A1(_u10_u7_n2192 ), .A2(_u10_u7_n2021 ), .A3(_u10_u7_n2193 ), .A4(_u10_u7_n2194 ), .ZN(_u10_u7_n2188 ) );
NAND2_X1 _u10_u7_U180  ( .A1(_u10_u7_n2188 ), .A2(_u10_u7_n2191 ), .ZN(_u10_u7_n2181 ) );
NAND2_X1 _u10_u7_U179  ( .A1(1'b0), .A2(_u10_u7_n2190 ), .ZN(_u10_u7_n2185 ));
NAND2_X1 _u10_u7_U178  ( .A1(_u10_u7_n2189 ), .A2(_u10_SYNOPSYS_UNCONNECTED_31 ), .ZN(_u10_u7_n2186 ) );
INV_X1 _u10_u7_U177  ( .A(_u10_u7_n2188 ), .ZN(_u10_u7_n2187 ) );
NAND3_X1 _u10_u7_U176  ( .A1(_u10_u7_n2185 ), .A2(_u10_u7_n2186 ), .A3(_u10_u7_n2187 ), .ZN(_u10_u7_n2184 ) );
NAND2_X1 _u10_u7_U175  ( .A1(_u10_u7_n2183 ), .A2(_u10_u7_n2184 ), .ZN(_u10_u7_n2182 ) );
NAND3_X1 _u10_u7_U174  ( .A1(_u10_u7_n2180 ), .A2(_u10_u7_n2181 ), .A3(_u10_u7_n2182 ), .ZN(_u10_u7_n2171 ) );
INV_X1 _u10_u7_U173  ( .A(_u10_u7_n2179 ), .ZN(_u10_u7_n1963 ) );
NOR2_X1 _u10_u7_U172  ( .A1(_u10_u7_n1963 ), .A2(_u10_u7_n2178 ), .ZN(_u10_u7_n2172 ) );
INV_X1 _u10_u7_U171  ( .A(_u10_u7_n2177 ), .ZN(_u10_u7_n2176 ) );
NOR3_X1 _u10_u7_U170  ( .A1(_u10_u7_n2174 ), .A2(_u10_u7_n2175 ), .A3(_u10_u7_n2176 ), .ZN(_u10_u7_n2173 ) );
NOR4_X1 _u10_u7_U169  ( .A1(_u10_u7_n2170 ), .A2(_u10_u7_n2171 ), .A3(_u10_u7_n2172 ), .A4(_u10_u7_n2173 ), .ZN(_u10_u7_n2119 ) );
NAND3_X1 _u10_u7_U168  ( .A1(_u10_u7_n2168 ), .A2(_u10_u7_n2169 ), .A3(1'b0),.ZN(_u10_u7_n2148 ) );
NAND3_X1 _u10_u7_U167  ( .A1(_u10_u7_n2165 ), .A2(_u10_u7_n2166 ), .A3(_u10_u7_n2167 ), .ZN(_u10_u7_n2149 ) );
NAND4_X1 _u10_u7_U166  ( .A1(_u10_u7_n2162 ), .A2(_u10_u7_n1933 ), .A3(_u10_u7_n2163 ), .A4(_u10_u7_n2164 ), .ZN(_u10_u7_n2160 ) );
NOR4_X1 _u10_u7_U165  ( .A1(_u10_u7_n2160 ), .A2(_u10_u7_n2157 ), .A3(_u10_u7_n1844 ), .A4(_u10_u7_n2161 ), .ZN(_u10_u7_n2158 ) );
NOR2_X1 _u10_u7_U164  ( .A1(_u10_u7_n2158 ), .A2(_u10_u7_n2159 ), .ZN(_u10_u7_n2153 ) );
INV_X1 _u10_u7_U163  ( .A(_u10_u7_n2157 ), .ZN(_u10_u7_n2129 ) );
NOR3_X1 _u10_u7_U162  ( .A1(_u10_u7_n2155 ), .A2(_u10_u7_n2129 ), .A3(_u10_u7_n2156 ), .ZN(_u10_u7_n2154 ) );
NOR2_X1 _u10_u7_U161  ( .A1(_u10_u7_n2153 ), .A2(_u10_u7_n2154 ), .ZN(_u10_u7_n2150 ) );
NAND3_X1 _u10_u7_U160  ( .A1(1'b0), .A2(_u10_u7_n1928 ), .A3(_u10_u7_n2152 ),.ZN(_u10_u7_n2151 ) );
NAND4_X1 _u10_u7_U159  ( .A1(_u10_u7_n2148 ), .A2(_u10_u7_n2149 ), .A3(_u10_u7_n2150 ), .A4(_u10_u7_n2151 ), .ZN(_u10_u7_n2121 ) );
NAND2_X1 _u10_u7_U158  ( .A1(_u10_u7_n2107 ), .A2(_u10_u7_n2147 ), .ZN(_u10_u7_n2146 ) );
NAND2_X1 _u10_u7_U157  ( .A1(_u10_u7_n2145 ), .A2(_u10_u7_n2146 ), .ZN(_u10_u7_n2144 ) );
NAND2_X1 _u10_u7_U156  ( .A1(_u10_u7_n2143 ), .A2(_u10_u7_n2144 ), .ZN(_u10_u7_n2134 ) );
NAND2_X1 _u10_u7_U155  ( .A1(_u10_u7_n2141 ), .A2(_u10_u7_n2142 ), .ZN(_u10_u7_n2140 ) );
NAND2_X1 _u10_u7_U154  ( .A1(_u10_u7_n2139 ), .A2(_u10_u7_n2140 ), .ZN(_u10_u7_n2135 ) );
OR2_X1 _u10_u7_U153  ( .A1(_u10_u7_n2110 ), .A2(_u10_u7_n1911 ), .ZN(_u10_u7_n2137 ) );
NAND2_X1 _u10_u7_U152  ( .A1(_u10_u7_n2137 ), .A2(_u10_u7_n2138 ), .ZN(_u10_u7_n2136 ) );
NAND3_X1 _u10_u7_U151  ( .A1(_u10_u7_n2134 ), .A2(_u10_u7_n2135 ), .A3(_u10_u7_n2136 ), .ZN(_u10_u7_n2122 ) );
NOR2_X1 _u10_u7_U150  ( .A1(_u10_u7_n2133 ), .A2(_u10_u7_n1891 ), .ZN(_u10_u7_n2132 ) );
NOR2_X1 _u10_u7_U149  ( .A1(_u10_u7_n2131 ), .A2(_u10_u7_n2132 ), .ZN(_u10_u7_n2123 ) );
NOR2_X1 _u10_u7_U148  ( .A1(_u10_u7_n2129 ), .A2(_u10_u7_n2130 ), .ZN(_u10_u7_n2127 ) );
NOR2_X1 _u10_u7_U147  ( .A1(_u10_u7_n2127 ), .A2(_u10_u7_n2128 ), .ZN(_u10_u7_n2125 ) );
NOR2_X1 _u10_u7_U146  ( .A1(_u10_u7_n2125 ), .A2(_u10_u7_n2126 ), .ZN(_u10_u7_n2124 ) );
NOR4_X1 _u10_u7_U145  ( .A1(_u10_u7_n2121 ), .A2(_u10_u7_n2122 ), .A3(_u10_u7_n2123 ), .A4(_u10_u7_n2124 ), .ZN(_u10_u7_n2120 ) );
NAND4_X1 _u10_u7_U144  ( .A1(_u10_u7_n2117 ), .A2(_u10_u7_n2118 ), .A3(_u10_u7_n2119 ), .A4(_u10_u7_n2120 ), .ZN(_u10_u7_n2116 ) );
MUX2_X1 _u10_u7_U143  ( .A(_u10_u7_n2116 ), .B(_u10_SYNOPSYS_UNCONNECTED_31 ), .S(_u10_u7_n1819 ), .Z(_u10_u7_n1811 ) );
INV_X1 _u10_u7_U142  ( .A(_u10_u7_n2115 ), .ZN(_u10_u7_n2006 ) );
NOR3_X1 _u10_u7_U141  ( .A1(_u10_u7_n2006 ), .A2(_u10_u7_n2114 ), .A3(_u10_u7_n2081 ), .ZN(_u10_u7_n1854 ) );
NAND2_X1 _u10_u7_U140  ( .A1(_u10_u7_n2112 ), .A2(_u10_u7_n2113 ), .ZN(_u10_u7_n1872 ) );
INV_X1 _u10_u7_U139  ( .A(_u10_u7_n1872 ), .ZN(_u10_u7_n1882 ) );
NAND4_X1 _u10_u7_U138  ( .A1(_u10_u7_n1854 ), .A2(_u10_u7_n1882 ), .A3(_u10_u7_n2111 ), .A4(_u10_u7_n1868 ), .ZN(_u10_u7_n2109 ) );
NAND2_X1 _u10_u7_U137  ( .A1(_u10_u7_n2109 ), .A2(_u10_u7_n2110 ), .ZN(_u10_u7_n2098 ) );
NAND2_X1 _u10_u7_U136  ( .A1(1'b0), .A2(_u10_u7_n1983 ), .ZN(_u10_u7_n2023 ));
INV_X1 _u10_u7_U135  ( .A(_u10_u7_n2023 ), .ZN(_u10_u7_n2035 ) );
NAND3_X1 _u10_u7_U134  ( .A1(_u10_u7_n2035 ), .A2(_u10_u7_n2107 ), .A3(_u10_u7_n2108 ), .ZN(_u10_u7_n1916 ) );
INV_X1 _u10_u7_U133  ( .A(_u10_u7_n1916 ), .ZN(_u10_u7_n2093 ) );
NAND3_X1 _u10_u7_U132  ( .A1(_u10_u7_n2105 ), .A2(_u10_u7_n2106 ), .A3(_u10_u7_n2093 ), .ZN(_u10_u7_n2039 ) );
NAND2_X1 _u10_u7_U131  ( .A1(_u10_u7_n2039 ), .A2(_u10_u7_n1930 ), .ZN(_u10_u7_n2104 ) );
NAND2_X1 _u10_u7_U130  ( .A1(_u10_u7_n2103 ), .A2(_u10_u7_n2104 ), .ZN(_u10_u7_n1863 ) );
OR2_X1 _u10_u7_U129  ( .A1(_u10_u7_n1863 ), .A2(_u10_u7_n2102 ), .ZN(_u10_u7_n2099 ) );
NAND2_X1 _u10_u7_U128  ( .A1(_u10_u7_n1890 ), .A2(_u10_u7_n2101 ), .ZN(_u10_u7_n2100 ) );
NAND3_X1 _u10_u7_U127  ( .A1(_u10_u7_n2098 ), .A2(_u10_u7_n2099 ), .A3(_u10_u7_n2100 ), .ZN(_u10_u7_n2066 ) );
NAND4_X1 _u10_u7_U126  ( .A1(_u10_u7_n2095 ), .A2(_u10_u7_n2096 ), .A3(_u10_u7_n1896 ), .A4(_u10_u7_n2097 ), .ZN(_u10_u7_n2086 ) );
NOR4_X1 _u10_u7_U125  ( .A1(_u10_u7_n2093 ), .A2(_u10_u7_n2027 ), .A3(_u10_u7_n2094 ), .A4(_u10_u7_n2026 ), .ZN(_u10_u7_n1952 ) );
NOR2_X1 _u10_u7_U124  ( .A1(1'b0), .A2(_u10_u7_n1952 ), .ZN(_u10_u7_n1951 ));
INV_X1 _u10_u7_U123  ( .A(_u10_u7_n1951 ), .ZN(_u10_u7_n2090 ) );
NAND4_X1 _u10_u7_U122  ( .A1(_u10_u7_n2089 ), .A2(_u10_u7_n2090 ), .A3(_u10_u7_n2091 ), .A4(_u10_u7_n2092 ), .ZN(_u10_u7_n1893 ) );
NOR4_X1 _u10_u7_U121  ( .A1(_u10_u7_n2086 ), .A2(_u10_u7_n1893 ), .A3(_u10_u7_n2087 ), .A4(_u10_u7_n2088 ), .ZN(_u10_u7_n2084 ) );
NOR2_X1 _u10_u7_U120  ( .A1(_u10_u7_n2084 ), .A2(_u10_u7_n2085 ), .ZN(_u10_u7_n2067 ) );
NOR2_X1 _u10_u7_U119  ( .A1(_u10_u7_n2083 ), .A2(_u10_u7_n1869 ), .ZN(_u10_u7_n2068 ) );
NAND2_X1 _u10_u7_U118  ( .A1(_u10_u7_n2081 ), .A2(_u10_u7_n2082 ), .ZN(_u10_u7_n2075 ) );
NAND2_X1 _u10_u7_U117  ( .A1(_u10_u7_n2035 ), .A2(_u10_u7_n2019 ), .ZN(_u10_u7_n2060 ) );
NAND2_X1 _u10_u7_U116  ( .A1(_u10_u7_n2080 ), .A2(_u10_u7_n2060 ), .ZN(_u10_u7_n2079 ) );
NAND2_X1 _u10_u7_U115  ( .A1(_u10_u7_n2078 ), .A2(_u10_u7_n2079 ), .ZN(_u10_u7_n2076 ) );
NAND4_X1 _u10_u7_U114  ( .A1(_u10_u7_n2075 ), .A2(_u10_u7_n2076 ), .A3(_u10_u7_n1970 ), .A4(_u10_u7_n2077 ), .ZN(_u10_u7_n2072 ) );
NOR4_X1 _u10_u7_U113  ( .A1(_u10_u7_n2072 ), .A2(_u10_u7_n2073 ), .A3(_u10_u7_n1975 ), .A4(_u10_u7_n2074 ), .ZN(_u10_u7_n2070 ) );
NOR2_X1 _u10_u7_U112  ( .A1(_u10_u7_n2070 ), .A2(_u10_u7_n2071 ), .ZN(_u10_u7_n2069 ) );
NOR4_X1 _u10_u7_U111  ( .A1(_u10_u7_n2066 ), .A2(_u10_u7_n2067 ), .A3(_u10_u7_n2068 ), .A4(_u10_u7_n2069 ), .ZN(_u10_u7_n1820 ) );
NAND2_X1 _u10_u7_U110  ( .A1(1'b0), .A2(_u10_u7_n1983 ), .ZN(_u10_u7_n2065 ));
NAND4_X1 _u10_u7_U109  ( .A1(_u10_u7_n2065 ), .A2(_u10_u7_n2023 ), .A3(_u10_u7_n2021 ), .A4(_u10_u7_n2052 ), .ZN(_u10_u7_n2064 ) );
NAND2_X1 _u10_u7_U108  ( .A1(_u10_u7_n2063 ), .A2(_u10_u7_n2064 ), .ZN(_u10_u7_n2040 ) );
NAND4_X1 _u10_u7_U107  ( .A1(_u10_u7_n2059 ), .A2(_u10_u7_n2060 ), .A3(_u10_u7_n2061 ), .A4(_u10_u7_n2062 ), .ZN(_u10_u7_n2058 ) );
NAND2_X1 _u10_u7_U106  ( .A1(_u10_u7_n2057 ), .A2(_u10_u7_n2058 ), .ZN(_u10_u7_n2041 ) );
NOR4_X1 _u10_u7_U105  ( .A1(1'b0), .A2(_u10_u7_n2054 ), .A3(_u10_u7_n2055 ),.A4(_u10_u7_n2056 ), .ZN(_u10_u7_n2053 ) );
NAND4_X1 _u10_u7_U104  ( .A1(_u10_u7_n2021 ), .A2(_u10_u7_n2052 ), .A3(_u10_u7_n2023 ), .A4(_u10_u7_n2053 ), .ZN(_u10_u7_n1964 ) );
INV_X1 _u10_u7_U103  ( .A(_u10_u7_n1964 ), .ZN(_u10_u7_n2045 ) );
NAND2_X1 _u10_u7_U102  ( .A1(_u10_u7_n2051 ), .A2(_u10_SYNOPSYS_UNCONNECTED_32 ), .ZN(_u10_u7_n2046 ) );
NAND2_X1 _u10_u7_U101  ( .A1(_u10_u7_n2049 ), .A2(_u10_u7_n2050 ), .ZN(_u10_u7_n2047 ) );
NAND4_X1 _u10_u7_U100  ( .A1(_u10_u7_n2045 ), .A2(_u10_u7_n2046 ), .A3(_u10_u7_n2047 ), .A4(_u10_u7_n2048 ), .ZN(_u10_u7_n2044 ) );
NAND2_X1 _u10_u7_U99  ( .A1(_u10_u7_n2043 ), .A2(_u10_u7_n2044 ), .ZN(_u10_u7_n2042 ) );
NAND3_X1 _u10_u7_U98  ( .A1(_u10_u7_n2040 ), .A2(_u10_u7_n2041 ), .A3(_u10_u7_n2042 ), .ZN(_u10_u7_n2009 ) );
AND2_X1 _u10_u7_U97  ( .A1(_u10_u7_n2038 ), .A2(_u10_u7_n2039 ), .ZN(_u10_u7_n1929 ) );
NOR2_X1 _u10_u7_U96  ( .A1(_u10_u7_n1929 ), .A2(_u10_u7_n2037 ), .ZN(_u10_u7_n2010 ) );
NAND2_X1 _u10_u7_U95  ( .A1(_u10_u7_n2035 ), .A2(_u10_u7_n2036 ), .ZN(_u10_u7_n1902 ) );
NAND3_X1 _u10_u7_U94  ( .A1(_u10_u7_n1902 ), .A2(_u10_u7_n2033 ), .A3(_u10_u7_n2034 ), .ZN(_u10_u7_n1973 ) );
NOR2_X1 _u10_u7_U93  ( .A1(_u10_u7_n1978 ), .A2(_u10_u7_n1973 ), .ZN(_u10_u7_n2032 ) );
NOR2_X1 _u10_u7_U92  ( .A1(1'b0), .A2(_u10_u7_n2032 ), .ZN(_u10_u7_n2028 ));
NOR2_X1 _u10_u7_U91  ( .A1(_u10_u7_n2030 ), .A2(_u10_u7_n2031 ), .ZN(_u10_u7_n2029 ) );
NOR4_X1 _u10_u7_U90  ( .A1(_u10_u7_n2026 ), .A2(_u10_u7_n2027 ), .A3(_u10_u7_n2028 ), .A4(_u10_u7_n2029 ), .ZN(_u10_u7_n2024 ) );
NOR2_X1 _u10_u7_U89  ( .A1(_u10_u7_n2024 ), .A2(_u10_u7_n2025 ), .ZN(_u10_u7_n2011 ) );
NAND3_X1 _u10_u7_U88  ( .A1(_u10_u7_n2021 ), .A2(_u10_u7_n2022 ), .A3(_u10_u7_n2023 ), .ZN(_u10_u7_n2020 ) );
AND2_X1 _u10_u7_U87  ( .A1(_u10_u7_n2019 ), .A2(_u10_u7_n2020 ), .ZN(_u10_u7_n1838 ) );
INV_X1 _u10_u7_U86  ( .A(_u10_u7_n2018 ), .ZN(_u10_u7_n2016 ) );
NOR4_X1 _u10_u7_U85  ( .A1(_u10_u7_n2015 ), .A2(_u10_u7_n1838 ), .A3(_u10_u7_n2016 ), .A4(_u10_u7_n2017 ), .ZN(_u10_u7_n2013 ) );
NOR2_X1 _u10_u7_U84  ( .A1(_u10_u7_n2013 ), .A2(_u10_u7_n2014 ), .ZN(_u10_u7_n2012 ) );
NOR4_X1 _u10_u7_U83  ( .A1(_u10_u7_n2009 ), .A2(_u10_u7_n2010 ), .A3(_u10_u7_n2011 ), .A4(_u10_u7_n2012 ), .ZN(_u10_u7_n1821 ) );
NAND2_X1 _u10_u7_U82  ( .A1(_u10_u7_n1924 ), .A2(_u10_u7_n2008 ), .ZN(_u10_u7_n1993 ) );
NAND2_X1 _u10_u7_U81  ( .A1(_u10_u7_n2006 ), .A2(_u10_u7_n2007 ), .ZN(_u10_u7_n1994 ) );
NAND2_X1 _u10_u7_U80  ( .A1(_u10_u7_n2004 ), .A2(_u10_u7_n2005 ), .ZN(_u10_u7_n1995 ) );
AND2_X1 _u10_u7_U79  ( .A1(_u10_u7_n2002 ), .A2(_u10_u7_n2003 ), .ZN(_u10_u7_n1998 ) );
NOR2_X1 _u10_u7_U78  ( .A1(_u10_u7_n2000 ), .A2(_u10_u7_n2001 ), .ZN(_u10_u7_n1999 ) );
NOR3_X1 _u10_u7_U77  ( .A1(_u10_u7_n1997 ), .A2(_u10_u7_n1998 ), .A3(_u10_u7_n1999 ), .ZN(_u10_u7_n1996 ) );
NAND4_X1 _u10_u7_U76  ( .A1(_u10_u7_n1993 ), .A2(_u10_u7_n1994 ), .A3(_u10_u7_n1995 ), .A4(_u10_u7_n1996 ), .ZN(_u10_u7_n1985 ) );
INV_X1 _u10_u7_U75  ( .A(_u10_u7_n1992 ), .ZN(_u10_u7_n1989 ) );
NAND3_X1 _u10_u7_U74  ( .A1(_u10_u7_n1989 ), .A2(_u10_u7_n1990 ), .A3(_u10_u7_n1991 ), .ZN(_u10_u7_n1986 ) );
NOR4_X1 _u10_u7_U73  ( .A1(_u10_u7_n1985 ), .A2(_u10_u7_n1986 ), .A3(_u10_u7_n1987 ), .A4(_u10_u7_n1988 ), .ZN(_u10_u7_n1822 ) );
INV_X1 _u10_u7_U72  ( .A(_u10_u7_n1984 ), .ZN(_u10_u7_n1980 ) );
NAND4_X1 _u10_u7_U71  ( .A1(_u10_u7_n1980 ), .A2(_u10_u7_n1981 ), .A3(_u10_u7_n1982 ), .A4(_u10_u7_n1983 ), .ZN(_u10_u7_n1941 ) );
NOR3_X1 _u10_u7_U70  ( .A1(_u10_u7_n1977 ), .A2(_u10_u7_n1978 ), .A3(_u10_u7_n1979 ), .ZN(_u10_u7_n1971 ) );
NOR4_X1 _u10_u7_U69  ( .A1(_u10_u7_n1973 ), .A2(_u10_u7_n1974 ), .A3(_u10_u7_n1975 ), .A4(_u10_u7_n1976 ), .ZN(_u10_u7_n1972 ) );
NAND4_X1 _u10_u7_U68  ( .A1(_u10_u7_n1969 ), .A2(_u10_u7_n1970 ), .A3(_u10_u7_n1971 ), .A4(_u10_u7_n1972 ), .ZN(_u10_u7_n1968 ) );
NAND2_X1 _u10_u7_U67  ( .A1(_u10_u7_n1967 ), .A2(_u10_u7_n1968 ), .ZN(_u10_u7_n1942 ) );
NAND3_X1 _u10_u7_U66  ( .A1(_u10_u7_n1964 ), .A2(_u10_u7_n1965 ), .A3(_u10_u7_n1966 ), .ZN(_u10_u7_n1943 ) );
AND4_X1 _u10_u7_U65  ( .A1(_u10_u7_n1961 ), .A2(_u10_u7_n1863 ), .A3(_u10_u7_n1962 ), .A4(_u10_u7_n1963 ), .ZN(_u10_u7_n1957 ) );
NOR2_X1 _u10_u7_U64  ( .A1(_u10_u7_n1959 ), .A2(_u10_u7_n1960 ), .ZN(_u10_u7_n1958 ) );
NOR2_X1 _u10_u7_U63  ( .A1(_u10_u7_n1957 ), .A2(_u10_u7_n1958 ), .ZN(_u10_u7_n1945 ) );
NOR2_X1 _u10_u7_U62  ( .A1(_u10_u7_n1955 ), .A2(_u10_u7_n1956 ), .ZN(_u10_u7_n1953 ) );
NOR4_X1 _u10_u7_U61  ( .A1(_u10_u7_n1952 ), .A2(_u10_u7_n1953 ), .A3(_u10_u7_n1846 ), .A4(_u10_u7_n1954 ), .ZN(_u10_u7_n1946 ) );
NOR2_X1 _u10_u7_U60  ( .A1(_u10_u7_n1950 ), .A2(_u10_u7_n1951 ), .ZN(_u10_u7_n1949 ) );
NOR2_X1 _u10_u7_U59  ( .A1(_u10_u7_n1948 ), .A2(_u10_u7_n1949 ), .ZN(_u10_u7_n1947 ) );
NOR3_X1 _u10_u7_U58  ( .A1(_u10_u7_n1945 ), .A2(_u10_u7_n1946 ), .A3(_u10_u7_n1947 ), .ZN(_u10_u7_n1944 ) );
NAND4_X1 _u10_u7_U57  ( .A1(_u10_u7_n1941 ), .A2(_u10_u7_n1942 ), .A3(_u10_u7_n1943 ), .A4(_u10_u7_n1944 ), .ZN(_u10_u7_n1824 ) );
NAND2_X1 _u10_u7_U56  ( .A1(_u10_u7_n1939 ), .A2(_u10_u7_n1940 ), .ZN(_u10_u7_n1938 ) );
NAND2_X1 _u10_u7_U55  ( .A1(_u10_u7_n1937 ), .A2(_u10_u7_n1938 ), .ZN(_u10_u7_n1903 ) );
NAND2_X1 _u10_u7_U54  ( .A1(_u10_u7_n1935 ), .A2(_u10_u7_n1936 ), .ZN(_u10_u7_n1934 ) );
NAND2_X1 _u10_u7_U53  ( .A1(_u10_u7_n1933 ), .A2(_u10_u7_n1934 ), .ZN(_u10_u7_n1931 ) );
NAND2_X1 _u10_u7_U52  ( .A1(_u10_u7_n1931 ), .A2(_u10_u7_n1932 ), .ZN(_u10_u7_n1904 ) );
NAND2_X1 _u10_u7_U51  ( .A1(_u10_u7_n1929 ), .A2(_u10_u7_n1930 ), .ZN(_u10_u7_n1927 ) );
NAND2_X1 _u10_u7_U50  ( .A1(_u10_u7_n1927 ), .A2(_u10_u7_n1928 ), .ZN(_u10_u7_n1905 ) );
NOR3_X1 _u10_u7_U49  ( .A1(_u10_u7_n1916 ), .A2(_u10_u7_n1925 ), .A3(_u10_u7_n1926 ), .ZN(_u10_u7_n1919 ) );
NOR2_X1 _u10_u7_U48  ( .A1(_u10_u7_n1923 ), .A2(_u10_u7_n1924 ), .ZN(_u10_u7_n1921 ) );
NOR2_X1 _u10_u7_U47  ( .A1(_u10_u7_n1921 ), .A2(_u10_u7_n1922 ), .ZN(_u10_u7_n1920 ) );
NOR2_X1 _u10_u7_U46  ( .A1(_u10_u7_n1919 ), .A2(_u10_u7_n1920 ), .ZN(_u10_u7_n1917 ) );
NOR2_X1 _u10_u7_U45  ( .A1(_u10_u7_n1917 ), .A2(_u10_u7_n1918 ), .ZN(_u10_u7_n1907 ) );
NOR2_X1 _u10_u7_U44  ( .A1(_u10_u7_n1915 ), .A2(_u10_u7_n1916 ), .ZN(_u10_u7_n1914 ) );
NOR2_X1 _u10_u7_U43  ( .A1(_u10_u7_n1914 ), .A2(1'b0), .ZN(_u10_u7_n1912 ));
NOR2_X1 _u10_u7_U42  ( .A1(_u10_u7_n1912 ), .A2(_u10_u7_n1913 ), .ZN(_u10_u7_n1908 ) );
NOR2_X1 _u10_u7_U41  ( .A1(_u10_u7_n1891 ), .A2(_u10_u7_n1911 ), .ZN(_u10_u7_n1910 ) );
NOR2_X1 _u10_u7_U40  ( .A1(_u10_u7_n1910 ), .A2(_u10_u7_n1868 ), .ZN(_u10_u7_n1909 ) );
NOR3_X1 _u10_u7_U39  ( .A1(_u10_u7_n1907 ), .A2(_u10_u7_n1908 ), .A3(_u10_u7_n1909 ), .ZN(_u10_u7_n1906 ) );
NAND4_X1 _u10_u7_U38  ( .A1(_u10_u7_n1903 ), .A2(_u10_u7_n1904 ), .A3(_u10_u7_n1905 ), .A4(_u10_u7_n1906 ), .ZN(_u10_u7_n1825 ) );
NAND2_X1 _u10_u7_U37  ( .A1(_u10_u7_n1901 ), .A2(_u10_u7_n1902 ), .ZN(_u10_u7_n1900 ) );
NAND2_X1 _u10_u7_U36  ( .A1(_u10_u7_n1899 ), .A2(_u10_u7_n1900 ), .ZN(_u10_u7_n1875 ) );
OR2_X1 _u10_u7_U35  ( .A1(_u10_u7_n1847 ), .A2(_u10_u7_n1898 ), .ZN(_u10_u7_n1897 ) );
NAND2_X1 _u10_u7_U34  ( .A1(_u10_u7_n1896 ), .A2(_u10_u7_n1897 ), .ZN(_u10_u7_n1895 ) );
NAND2_X1 _u10_u7_U33  ( .A1(_u10_u7_n1894 ), .A2(_u10_u7_n1895 ), .ZN(_u10_u7_n1876 ) );
NAND2_X1 _u10_u7_U32  ( .A1(_u10_u7_n1892 ), .A2(_u10_u7_n1893 ), .ZN(_u10_u7_n1877 ) );
NOR3_X1 _u10_u7_U31  ( .A1(_u10_u7_n1884 ), .A2(_u10_u7_n1890 ), .A3(_u10_u7_n1891 ), .ZN(_u10_u7_n1889 ) );
NOR2_X1 _u10_u7_U30  ( .A1(_u10_u7_n1840 ), .A2(_u10_u7_n1889 ), .ZN(_u10_u7_n1879 ) );
NOR2_X1 _u10_u7_U29  ( .A1(_u10_u7_n1887 ), .A2(_u10_u7_n1888 ), .ZN(_u10_u7_n1880 ) );
NOR3_X1 _u10_u7_U28  ( .A1(_u10_u7_n1884 ), .A2(_u10_u7_n1885 ), .A3(_u10_u7_n1886 ), .ZN(_u10_u7_n1883 ) );
NOR2_X1 _u10_u7_U27  ( .A1(_u10_u7_n1882 ), .A2(_u10_u7_n1883 ), .ZN(_u10_u7_n1881 ) );
NOR3_X1 _u10_u7_U26  ( .A1(_u10_u7_n1879 ), .A2(_u10_u7_n1880 ), .A3(_u10_u7_n1881 ), .ZN(_u10_u7_n1878 ) );
NAND4_X1 _u10_u7_U25  ( .A1(_u10_u7_n1875 ), .A2(_u10_u7_n1876 ), .A3(_u10_u7_n1877 ), .A4(_u10_u7_n1878 ), .ZN(_u10_u7_n1826 ) );
NOR3_X1 _u10_u7_U24  ( .A1(_u10_u7_n1872 ), .A2(_u10_u7_n1873 ), .A3(_u10_u7_n1874 ), .ZN(_u10_u7_n1871 ) );
NAND4_X1 _u10_u7_U23  ( .A1(_u10_u7_n1868 ), .A2(_u10_u7_n1869 ), .A3(_u10_u7_n1870 ), .A4(_u10_u7_n1871 ), .ZN(_u10_u7_n1867 ) );
NAND2_X1 _u10_u7_U22  ( .A1(_u10_u7_n1866 ), .A2(_u10_u7_n1867 ), .ZN(_u10_u7_n1865 ) );
NAND3_X1 _u10_u7_U21  ( .A1(_u10_u7_n1863 ), .A2(_u10_u7_n1864 ), .A3(_u10_u7_n1865 ), .ZN(_u10_u7_n1862 ) );
NAND2_X1 _u10_u7_U20  ( .A1(_u10_u7_n1861 ), .A2(_u10_u7_n1862 ), .ZN(_u10_u7_n1828 ) );
NAND3_X1 _u10_u7_U19  ( .A1(_u10_u7_n1858 ), .A2(_u10_u7_n1859 ), .A3(_u10_u7_n1860 ), .ZN(_u10_u7_n1857 ) );
NAND2_X1 _u10_u7_U18  ( .A1(_u10_u7_n1856 ), .A2(_u10_u7_n1857 ), .ZN(_u10_u7_n1829 ) );
OR2_X1 _u10_u7_U17  ( .A1(_u10_u7_n1854 ), .A2(_u10_u7_n1855 ), .ZN(_u10_u7_n1830 ) );
NOR2_X1 _u10_u7_U16  ( .A1(_u10_u7_n1852 ), .A2(_u10_u7_n1853 ), .ZN(_u10_u7_n1850 ) );
NOR3_X1 _u10_u7_U15  ( .A1(_u10_u7_n1850 ), .A2(_u10_u7_n1851 ), .A3(_u10_u7_n1838 ), .ZN(_u10_u7_n1848 ) );
NOR2_X1 _u10_u7_U14  ( .A1(_u10_u7_n1848 ), .A2(_u10_u7_n1849 ), .ZN(_u10_u7_n1832 ) );
NOR2_X1 _u10_u7_U13  ( .A1(_u10_u7_n1846 ), .A2(_u10_u7_n1847 ), .ZN(_u10_u7_n1845 ) );
NOR3_X1 _u10_u7_U12  ( .A1(_u10_u7_n1844 ), .A2(1'b0), .A3(_u10_u7_n1845 ),.ZN(_u10_u7_n1842 ) );
NOR2_X1 _u10_u7_U11  ( .A1(_u10_u7_n1842 ), .A2(_u10_u7_n1843 ), .ZN(_u10_u7_n1833 ) );
NOR2_X1 _u10_u7_U10  ( .A1(_u10_u7_n1840 ), .A2(_u10_u7_n1841 ), .ZN(_u10_u7_n1839 ) );
NOR3_X1 _u10_u7_U9  ( .A1(_u10_u7_n1837 ), .A2(_u10_u7_n1838 ), .A3(_u10_u7_n1839 ), .ZN(_u10_u7_n1835 ) );
NOR2_X1 _u10_u7_U8  ( .A1(_u10_u7_n1835 ), .A2(_u10_u7_n1836 ), .ZN(_u10_u7_n1834 ) );
NOR3_X1 _u10_u7_U7  ( .A1(_u10_u7_n1832 ), .A2(_u10_u7_n1833 ), .A3(_u10_u7_n1834 ), .ZN(_u10_u7_n1831 ) );
NAND4_X1 _u10_u7_U6  ( .A1(_u10_u7_n1828 ), .A2(_u10_u7_n1829 ), .A3(_u10_u7_n1830 ), .A4(_u10_u7_n1831 ), .ZN(_u10_u7_n1827 ) );
NOR4_X1 _u10_u7_U5  ( .A1(_u10_u7_n1824 ), .A2(_u10_u7_n1825 ), .A3(_u10_u7_n1826 ), .A4(_u10_u7_n1827 ), .ZN(_u10_u7_n1823 ) );
NAND4_X1 _u10_u7_U4  ( .A1(_u10_u7_n1820 ), .A2(_u10_u7_n1821 ), .A3(_u10_u7_n1822 ), .A4(_u10_u7_n1823 ), .ZN(_u10_u7_n1818 ) );
MUX2_X1 _u10_u7_U3  ( .A(_u10_u7_n1818 ), .B(_u10_SYNOPSYS_UNCONNECTED_32 ),.S(_u10_u7_n1819 ), .Z(_u10_u7_n1812 ) );
DFFR_X1 _u10_u7_state_reg_1_  ( .D(_u10_u7_n1812 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_32 ), .QN(_u10_u7_n1814 ));
DFFR_X1 _u10_u7_state_reg_2_  ( .D(_u10_u7_n1811 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_31 ), .QN(_u10_u7_n1815 ));
DFFR_X1 _u10_u7_state_reg_3_  ( .D(_u10_u7_n1810 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_30 ), .QN(_u10_u7_n1816 ));
DFFR_X1 _u10_u7_state_reg_4_  ( .D(_u10_u7_n1809 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_29 ), .QN(_u10_u7_n1817 ));
DFFR_X1 _u10_u7_state_reg_0_  ( .D(_u10_u7_n1808 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_33 ), .QN(_u10_u7_n1813 ));
NOR2_X1 _u10_u8_U1606  ( .A1(_u10_SYNOPSYS_UNCONNECTED_36 ), .A2(_u10_u8_n1814 ), .ZN(_u10_u8_n3174 ) );
NOR3_X1 _u10_u8_U1605  ( .A1(_u10_SYNOPSYS_UNCONNECTED_35 ), .A2(_u10_u8_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_38 ), .ZN(_u10_u8_n3328 ) );
NAND2_X1 _u10_u8_U1604  ( .A1(_u10_u8_n3174 ), .A2(_u10_u8_n3328 ), .ZN(_u10_u8_n1843 ) );
INV_X1 _u10_u8_U1603  ( .A(_u10_u8_n1843 ), .ZN(_u10_u8_n2461 ) );
INV_X1 _u10_u8_U1602  ( .A(1'b0), .ZN(_u10_u8_n2466 ) );
INV_X1 _u10_u8_U1601  ( .A(1'b0), .ZN(_u10_u8_n2305 ) );
NAND2_X1 _u10_u8_U1600  ( .A1(_u10_u8_n2466 ), .A2(_u10_u8_n2305 ), .ZN(_u10_u8_n1954 ) );
INV_X1 _u10_u8_U1599  ( .A(_u10_u8_n1954 ), .ZN(_u10_u8_n2467 ) );
INV_X1 _u10_u8_U1598  ( .A(1'b0), .ZN(_u10_u8_n1936 ) );
NOR2_X1 _u10_u8_U1597  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u8_n2223 ) );
INV_X1 _u10_u8_U1596  ( .A(1'b0), .ZN(_u10_u8_n1922 ) );
NAND2_X1 _u10_u8_U1595  ( .A1(_u10_u8_n2223 ), .A2(_u10_u8_n1922 ), .ZN(_u10_u8_n2200 ) );
NOR2_X1 _u10_u8_U1594  ( .A1(_u10_u8_n2200 ), .A2(1'b0), .ZN(_u10_u8_n2502 ));
INV_X1 _u10_u8_U1593  ( .A(1'b0), .ZN(_u10_u8_n2978 ) );
INV_X1 _u10_u8_U1592  ( .A(1'b0), .ZN(_u10_u8_n3000 ) );
NAND2_X1 _u10_u8_U1591  ( .A1(_u10_u8_n2978 ), .A2(_u10_u8_n3000 ), .ZN(_u10_u8_n3356 ) );
INV_X1 _u10_u8_U1590  ( .A(1'b0), .ZN(_u10_u8_n2405 ) );
INV_X1 _u10_u8_U1589  ( .A(1'b0), .ZN(_u10_u8_n2972 ) );
NAND2_X1 _u10_u8_U1588  ( .A1(_u10_u8_n2405 ), .A2(_u10_u8_n2972 ), .ZN(_u10_u8_n2008 ) );
NOR2_X1 _u10_u8_U1587  ( .A1(_u10_u8_n3356 ), .A2(_u10_u8_n2008 ), .ZN(_u10_u8_n2195 ) );
NAND2_X1 _u10_u8_U1586  ( .A1(_u10_u8_n2502 ), .A2(_u10_u8_n2195 ), .ZN(_u10_u8_n2490 ) );
INV_X1 _u10_u8_U1585  ( .A(1'b0), .ZN(_u10_u8_n3040 ) );
INV_X1 _u10_u8_U1584  ( .A(1'b0), .ZN(_u10_u8_n3006 ) );
NAND2_X1 _u10_u8_U1583  ( .A1(_u10_u8_n3040 ), .A2(_u10_u8_n3006 ), .ZN(_u10_u8_n2508 ) );
NOR2_X1 _u10_u8_U1582  ( .A1(_u10_u8_n2508 ), .A2(1'b0), .ZN(_u10_u8_n2493 ));
INV_X1 _u10_u8_U1581  ( .A(1'b0), .ZN(_u10_u8_n2038 ) );
NAND2_X1 _u10_u8_U1580  ( .A1(_u10_u8_n2493 ), .A2(_u10_u8_n2038 ), .ZN(_u10_u8_n2174 ) );
NOR2_X1 _u10_u8_U1579  ( .A1(_u10_u8_n2490 ), .A2(_u10_u8_n2174 ), .ZN(_u10_u8_n2659 ) );
INV_X1 _u10_u8_U1578  ( .A(1'b0), .ZN(_u10_u8_n2175 ) );
NAND3_X1 _u10_u8_U1577  ( .A1(_u10_u8_n2659 ), .A2(_u10_u8_n2175 ), .A3(1'b0), .ZN(_u10_u8_n3189 ) );
NOR2_X1 _u10_u8_U1576  ( .A1(_u10_u8_n3189 ), .A2(1'b0), .ZN(_u10_u8_n2528 ));
INV_X1 _u10_u8_U1575  ( .A(1'b0), .ZN(_u10_u8_n2837 ) );
NAND2_X1 _u10_u8_U1574  ( .A1(_u10_u8_n2528 ), .A2(_u10_u8_n2837 ), .ZN(_u10_u8_n2567 ) );
INV_X1 _u10_u8_U1573  ( .A(1'b0), .ZN(_u10_u8_n2080 ) );
INV_X1 _u10_u8_U1572  ( .A(1'b0), .ZN(_u10_u8_n2166 ) );
NAND2_X1 _u10_u8_U1571  ( .A1(_u10_u8_n2080 ), .A2(_u10_u8_n2166 ), .ZN(_u10_u8_n2840 ) );
NOR2_X1 _u10_u8_U1570  ( .A1(_u10_u8_n2567 ), .A2(_u10_u8_n2840 ), .ZN(_u10_u8_n2443 ) );
INV_X1 _u10_u8_U1569  ( .A(1'b0), .ZN(_u10_u8_n2600 ) );
INV_X1 _u10_u8_U1568  ( .A(1'b0), .ZN(_u10_u8_n2836 ) );
NAND2_X1 _u10_u8_U1567  ( .A1(_u10_u8_n2600 ), .A2(_u10_u8_n2836 ), .ZN(_u10_u8_n2428 ) );
INV_X1 _u10_u8_U1566  ( .A(_u10_u8_n2428 ), .ZN(_u10_u8_n2078 ) );
NAND2_X1 _u10_u8_U1565  ( .A1(_u10_u8_n2443 ), .A2(_u10_u8_n2078 ), .ZN(_u10_u8_n2282 ) );
INV_X1 _u10_u8_U1564  ( .A(1'b0), .ZN(_u10_u8_n2874 ) );
INV_X1 _u10_u8_U1563  ( .A(1'b0), .ZN(_u10_u8_n2031 ) );
NAND2_X1 _u10_u8_U1562  ( .A1(_u10_u8_n2874 ), .A2(_u10_u8_n2031 ), .ZN(_u10_u8_n1976 ) );
NOR2_X1 _u10_u8_U1561  ( .A1(_u10_u8_n2282 ), .A2(_u10_u8_n1976 ), .ZN(_u10_u8_n2411 ) );
NAND3_X1 _u10_u8_U1560  ( .A1(_u10_u8_n2467 ), .A2(_u10_u8_n1936 ), .A3(_u10_u8_n2411 ), .ZN(_u10_u8_n2464 ) );
NAND3_X1 _u10_u8_U1559  ( .A1(_u10_u8_n2166 ), .A2(_u10_u8_n2837 ), .A3(1'b0), .ZN(_u10_u8_n3276 ) );
INV_X1 _u10_u8_U1558  ( .A(_u10_u8_n3276 ), .ZN(_u10_u8_n2442 ) );
NAND3_X1 _u10_u8_U1557  ( .A1(_u10_u8_n2836 ), .A2(_u10_u8_n2080 ), .A3(_u10_u8_n2442 ), .ZN(_u10_u8_n2838 ) );
INV_X1 _u10_u8_U1556  ( .A(_u10_u8_n2838 ), .ZN(_u10_u8_n2850 ) );
NOR2_X1 _u10_u8_U1555  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u8_n2953 ) );
NAND2_X1 _u10_u8_U1554  ( .A1(_u10_u8_n2850 ), .A2(_u10_u8_n2953 ), .ZN(_u10_u8_n2947 ) );
INV_X1 _u10_u8_U1553  ( .A(_u10_u8_n2947 ), .ZN(_u10_u8_n2420 ) );
NAND2_X1 _u10_u8_U1552  ( .A1(_u10_u8_n1936 ), .A2(_u10_u8_n2874 ), .ZN(_u10_u8_n2030 ) );
INV_X1 _u10_u8_U1551  ( .A(_u10_u8_n2030 ), .ZN(_u10_u8_n2162 ) );
NAND2_X1 _u10_u8_U1550  ( .A1(_u10_u8_n2420 ), .A2(_u10_u8_n2162 ), .ZN(_u10_u8_n2828 ) );
INV_X1 _u10_u8_U1549  ( .A(_u10_u8_n2828 ), .ZN(_u10_u8_n2551 ) );
NAND2_X1 _u10_u8_U1548  ( .A1(_u10_u8_n2551 ), .A2(_u10_u8_n2467 ), .ZN(_u10_u8_n3416 ) );
NAND2_X1 _u10_u8_U1547  ( .A1(_u10_u8_n2464 ), .A2(_u10_u8_n3416 ), .ZN(_u10_u8_n2266 ) );
INV_X1 _u10_u8_U1546  ( .A(_u10_u8_n2266 ), .ZN(_u10_u8_n3410 ) );
NAND2_X1 _u10_u8_U1545  ( .A1(1'b0), .A2(_u10_u8_n2305 ), .ZN(_u10_u8_n3411 ) );
INV_X1 _u10_u8_U1544  ( .A(_u10_u8_n3356 ), .ZN(_u10_u8_n1983 ) );
NAND3_X1 _u10_u8_U1543  ( .A1(_u10_u8_n1983 ), .A2(_u10_u8_n2405 ), .A3(1'b0), .ZN(_u10_u8_n2022 ) );
INV_X1 _u10_u8_U1542  ( .A(_u10_u8_n2022 ), .ZN(_u10_u8_n2056 ) );
INV_X1 _u10_u8_U1541  ( .A(_u10_u8_n2840 ), .ZN(_u10_u8_n2059 ) );
INV_X1 _u10_u8_U1540  ( .A(1'b0), .ZN(_u10_u8_n1965 ) );
NAND2_X1 _u10_u8_U1539  ( .A1(_u10_u8_n2837 ), .A2(_u10_u8_n1965 ), .ZN(_u10_u8_n1852 ) );
INV_X1 _u10_u8_U1538  ( .A(_u10_u8_n1852 ), .ZN(_u10_u8_n3190 ) );
INV_X1 _u10_u8_U1537  ( .A(1'b0), .ZN(_u10_u8_n1853 ) );
NAND2_X1 _u10_u8_U1536  ( .A1(_u10_u8_n3190 ), .A2(_u10_u8_n1853 ), .ZN(_u10_u8_n2687 ) );
INV_X1 _u10_u8_U1535  ( .A(_u10_u8_n2687 ), .ZN(_u10_u8_n2019 ) );
NAND2_X1 _u10_u8_U1534  ( .A1(_u10_u8_n2059 ), .A2(_u10_u8_n2019 ), .ZN(_u10_u8_n2330 ) );
NOR2_X1 _u10_u8_U1533  ( .A1(_u10_u8_n2428 ), .A2(_u10_u8_n2330 ), .ZN(_u10_u8_n2036 ) );
NAND2_X1 _u10_u8_U1532  ( .A1(_u10_u8_n2056 ), .A2(_u10_u8_n2036 ), .ZN(_u10_u8_n3379 ) );
NOR2_X1 _u10_u8_U1531  ( .A1(_u10_u8_n3379 ), .A2(_u10_u8_n2030 ), .ZN(_u10_u8_n2026 ) );
INV_X1 _u10_u8_U1530  ( .A(1'b0), .ZN(_u10_u8_n2431 ) );
NOR2_X1 _u10_u8_U1529  ( .A1(_u10_u8_n2431 ), .A2(1'b0), .ZN(_u10_u8_n3062 ));
NAND2_X1 _u10_u8_U1528  ( .A1(_u10_u8_n3062 ), .A2(_u10_u8_n2195 ), .ZN(_u10_u8_n3407 ) );
NOR3_X1 _u10_u8_U1527  ( .A1(_u10_u8_n2687 ), .A2(1'b0), .A3(_u10_u8_n3407 ),.ZN(_u10_u8_n3275 ) );
NAND3_X1 _u10_u8_U1526  ( .A1(_u10_u8_n2836 ), .A2(_u10_u8_n2080 ), .A3(_u10_u8_n3275 ), .ZN(_u10_u8_n3297 ) );
INV_X1 _u10_u8_U1525  ( .A(_u10_u8_n3297 ), .ZN(_u10_u8_n3172 ) );
NAND2_X1 _u10_u8_U1524  ( .A1(_u10_u8_n3172 ), .A2(_u10_u8_n2600 ), .ZN(_u10_u8_n2226 ) );
NOR2_X1 _u10_u8_U1523  ( .A1(_u10_u8_n2226 ), .A2(1'b0), .ZN(_u10_u8_n2307 ));
INV_X1 _u10_u8_U1522  ( .A(_u10_u8_n2490 ), .ZN(_u10_u8_n2536 ) );
NAND3_X1 _u10_u8_U1521  ( .A1(_u10_u8_n2536 ), .A2(_u10_u8_n3040 ), .A3(1'b0), .ZN(_u10_u8_n3226 ) );
NOR2_X1 _u10_u8_U1520  ( .A1(_u10_u8_n3226 ), .A2(_u10_u8_n2330 ), .ZN(_u10_u8_n2441 ) );
NAND2_X1 _u10_u8_U1519  ( .A1(_u10_u8_n2441 ), .A2(_u10_u8_n2953 ), .ZN(_u10_u8_n2579 ) );
NOR2_X1 _u10_u8_U1518  ( .A1(_u10_u8_n2579 ), .A2(_u10_u8_n2030 ), .ZN(_u10_u8_n2550 ) );
NOR3_X1 _u10_u8_U1517  ( .A1(_u10_u8_n2026 ), .A2(_u10_u8_n2307 ), .A3(_u10_u8_n2550 ), .ZN(_u10_u8_n3394 ) );
NAND2_X1 _u10_u8_U1516  ( .A1(1'b0), .A2(_u10_u8_n2978 ), .ZN(_u10_u8_n3115 ) );
NOR2_X1 _u10_u8_U1515  ( .A1(_u10_u8_n3115 ), .A2(_u10_u8_n2330 ), .ZN(_u10_u8_n3126 ) );
NAND2_X1 _u10_u8_U1514  ( .A1(_u10_u8_n2162 ), .A2(_u10_u8_n2031 ), .ZN(_u10_u8_n2686 ) );
NOR2_X1 _u10_u8_U1513  ( .A1(_u10_u8_n2686 ), .A2(_u10_u8_n2428 ), .ZN(_u10_u8_n2108 ) );
NAND2_X1 _u10_u8_U1512  ( .A1(_u10_u8_n3126 ), .A2(_u10_u8_n2108 ), .ZN(_u10_u8_n3415 ) );
NAND2_X1 _u10_u8_U1511  ( .A1(_u10_u8_n3394 ), .A2(_u10_u8_n3415 ), .ZN(_u10_u8_n3089 ) );
NAND2_X1 _u10_u8_U1510  ( .A1(_u10_u8_n3089 ), .A2(_u10_u8_n2305 ), .ZN(_u10_u8_n3414 ) );
NAND2_X1 _u10_u8_U1509  ( .A1(_u10_u8_n2466 ), .A2(_u10_u8_n3414 ), .ZN(_u10_u8_n3118 ) );
NAND2_X1 _u10_u8_U1508  ( .A1(_u10_u8_n2078 ), .A2(_u10_u8_n2080 ), .ZN(_u10_u8_n2596 ) );
NAND2_X1 _u10_u8_U1507  ( .A1(1'b0), .A2(_u10_u8_n2493 ), .ZN(_u10_u8_n1961 ) );
NOR3_X1 _u10_u8_U1506  ( .A1(_u10_u8_n2490 ), .A2(1'b0), .A3(_u10_u8_n1961 ),.ZN(_u10_u8_n2054 ) );
NAND2_X1 _u10_u8_U1505  ( .A1(_u10_u8_n2054 ), .A2(_u10_u8_n3190 ), .ZN(_u10_u8_n2061 ) );
OR2_X1 _u10_u8_U1504  ( .A1(_u10_u8_n2596 ), .A2(_u10_u8_n2061 ), .ZN(_u10_u8_n1969 ) );
NOR3_X1 _u10_u8_U1503  ( .A1(_u10_u8_n1976 ), .A2(1'b0), .A3(_u10_u8_n1969 ),.ZN(_u10_u8_n2710 ) );
NAND2_X1 _u10_u8_U1502  ( .A1(_u10_u8_n2710 ), .A2(_u10_u8_n2467 ), .ZN(_u10_u8_n2545 ) );
INV_X1 _u10_u8_U1501  ( .A(_u10_u8_n2545 ), .ZN(_u10_u8_n2087 ) );
NOR2_X1 _u10_u8_U1500  ( .A1(_u10_u8_n3118 ), .A2(_u10_u8_n2087 ), .ZN(_u10_u8_n3145 ) );
NOR2_X1 _u10_u8_U1499  ( .A1(_u10_u8_n2030 ), .A2(1'b0), .ZN(_u10_u8_n2668 ));
NAND2_X1 _u10_u8_U1498  ( .A1(1'b0), .A2(_u10_u8_n2668 ), .ZN(_u10_u8_n2163 ) );
INV_X1 _u10_u8_U1497  ( .A(_u10_u8_n2163 ), .ZN(_u10_u8_n2875 ) );
INV_X1 _u10_u8_U1496  ( .A(_u10_u8_n1976 ), .ZN(_u10_u8_n2747 ) );
NAND3_X1 _u10_u8_U1495  ( .A1(_u10_u8_n2747 ), .A2(_u10_u8_n2600 ), .A3(1'b0), .ZN(_u10_u8_n3393 ) );
NOR3_X1 _u10_u8_U1494  ( .A1(1'b0), .A2(1'b0), .A3(_u10_u8_n3393 ), .ZN(_u10_u8_n3180 ) );
INV_X1 _u10_u8_U1493  ( .A(1'b0), .ZN(_u10_u8_n2113 ) );
INV_X1 _u10_u8_U1492  ( .A(1'b0), .ZN(_u10_u8_n3066 ) );
NAND2_X1 _u10_u8_U1491  ( .A1(_u10_u8_n2175 ), .A2(_u10_u8_n3066 ), .ZN(_u10_u8_n2216 ) );
INV_X1 _u10_u8_U1490  ( .A(_u10_u8_n2659 ), .ZN(_u10_u8_n2643 ) );
NOR2_X1 _u10_u8_U1489  ( .A1(_u10_u8_n2216 ), .A2(_u10_u8_n2643 ), .ZN(_u10_u8_n2049 ) );
AND2_X1 _u10_u8_U1488  ( .A1(_u10_u8_n2049 ), .A2(_u10_u8_n1853 ), .ZN(_u10_u8_n3223 ) );
NAND2_X1 _u10_u8_U1487  ( .A1(_u10_u8_n3223 ), .A2(_u10_u8_n1965 ), .ZN(_u10_u8_n2531 ) );
NOR2_X1 _u10_u8_U1486  ( .A1(_u10_u8_n2531 ), .A2(1'b0), .ZN(_u10_u8_n2884 ));
NAND2_X1 _u10_u8_U1485  ( .A1(_u10_u8_n2884 ), .A2(_u10_u8_n2166 ), .ZN(_u10_u8_n1841 ) );
NOR2_X1 _u10_u8_U1484  ( .A1(_u10_u8_n1841 ), .A2(1'b0), .ZN(_u10_u8_n3129 ));
NAND2_X1 _u10_u8_U1483  ( .A1(_u10_u8_n3129 ), .A2(_u10_u8_n2836 ), .ZN(_u10_u8_n2842 ) );
INV_X1 _u10_u8_U1482  ( .A(_u10_u8_n2842 ), .ZN(_u10_u8_n2833 ) );
NAND2_X1 _u10_u8_U1481  ( .A1(_u10_u8_n2833 ), .A2(_u10_u8_n2600 ), .ZN(_u10_u8_n2853 ) );
INV_X1 _u10_u8_U1480  ( .A(_u10_u8_n2853 ), .ZN(_u10_u8_n2082 ) );
NAND2_X1 _u10_u8_U1479  ( .A1(_u10_u8_n2082 ), .A2(_u10_u8_n2031 ), .ZN(_u10_u8_n2274 ) );
INV_X1 _u10_u8_U1478  ( .A(_u10_u8_n2274 ), .ZN(_u10_u8_n2669 ) );
NAND3_X1 _u10_u8_U1477  ( .A1(_u10_u8_n2668 ), .A2(_u10_u8_n2113 ), .A3(_u10_u8_n2669 ), .ZN(_u10_u8_n1858 ) );
INV_X1 _u10_u8_U1476  ( .A(_u10_u8_n1858 ), .ZN(_u10_u8_n3067 ) );
NAND2_X1 _u10_u8_U1475  ( .A1(_u10_u8_n3067 ), .A2(1'b0), .ZN(_u10_u8_n2092 ) );
INV_X1 _u10_u8_U1474  ( .A(_u10_u8_n2092 ), .ZN(_u10_u8_n3294 ) );
INV_X1 _u10_u8_U1473  ( .A(1'b0), .ZN(_u10_u8_n2446 ) );
INV_X1 _u10_u8_U1472  ( .A(1'b0), .ZN(_u10_u8_n2996 ) );
NAND2_X1 _u10_u8_U1471  ( .A1(_u10_u8_n3067 ), .A2(_u10_u8_n2996 ), .ZN(_u10_u8_n1847 ) );
NOR3_X1 _u10_u8_U1470  ( .A1(_u10_u8_n2446 ), .A2(1'b0), .A3(_u10_u8_n1847 ),.ZN(_u10_u8_n3413 ) );
NOR4_X1 _u10_u8_U1469  ( .A1(_u10_u8_n2875 ), .A2(_u10_u8_n3180 ), .A3(_u10_u8_n3294 ), .A4(_u10_u8_n3413 ), .ZN(_u10_u8_n3412 ) );
NAND4_X1 _u10_u8_U1468  ( .A1(_u10_u8_n3410 ), .A2(_u10_u8_n3411 ), .A3(_u10_u8_n3145 ), .A4(_u10_u8_n3412 ), .ZN(_u10_u8_n3409 ) );
NAND2_X1 _u10_u8_U1467  ( .A1(_u10_u8_n2461 ), .A2(_u10_u8_n3409 ), .ZN(_u10_u8_n3380 ) );
NOR2_X1 _u10_u8_U1466  ( .A1(_u10_u8_n1817 ), .A2(_u10_u8_n1816 ), .ZN(_u10_u8_n3368 ) );
AND2_X1 _u10_u8_U1465  ( .A1(_u10_u8_n3368 ), .A2(_u10_u8_n1813 ), .ZN(_u10_u8_n3320 ) );
NOR2_X1 _u10_u8_U1464  ( .A1(_u10_SYNOPSYS_UNCONNECTED_37 ), .A2(_u10_u8_n1815 ), .ZN(_u10_u8_n3236 ) );
NAND2_X1 _u10_u8_U1463  ( .A1(_u10_u8_n3320 ), .A2(_u10_u8_n3236 ), .ZN(_u10_u8_n2607 ) );
INV_X1 _u10_u8_U1462  ( .A(_u10_u8_n2607 ), .ZN(_u10_u8_n1966 ) );
INV_X1 _u10_u8_U1461  ( .A(_u10_u8_n2200 ), .ZN(_u10_u8_n3216 ) );
NAND2_X1 _u10_u8_U1460  ( .A1(1'b0), .A2(_u10_u8_n3216 ), .ZN(_u10_u8_n2367 ) );
INV_X1 _u10_u8_U1459  ( .A(_u10_u8_n2367 ), .ZN(_u10_u8_n3183 ) );
NAND2_X1 _u10_u8_U1458  ( .A1(_u10_u8_n3183 ), .A2(_u10_u8_n2195 ), .ZN(_u10_u8_n2194 ) );
INV_X1 _u10_u8_U1457  ( .A(_u10_u8_n2194 ), .ZN(_u10_u8_n2055 ) );
NAND2_X1 _u10_u8_U1456  ( .A1(_u10_u8_n2055 ), .A2(_u10_u8_n1853 ), .ZN(_u10_u8_n3401 ) );
INV_X1 _u10_u8_U1455  ( .A(_u10_u8_n2531 ), .ZN(_u10_u8_n2190 ) );
INV_X1 _u10_u8_U1454  ( .A(1'b0), .ZN(_u10_u8_n3001 ) );
NAND2_X1 _u10_u8_U1453  ( .A1(_u10_u8_n3001 ), .A2(_u10_u8_n2466 ), .ZN(_u10_u8_n2156 ) );
NOR2_X1 _u10_u8_U1452  ( .A1(_u10_u8_n2166 ), .A2(_u10_u8_n2596 ), .ZN(_u10_u8_n2594 ) );
NAND2_X1 _u10_u8_U1451  ( .A1(_u10_u8_n2594 ), .A2(_u10_u8_n2031 ), .ZN(_u10_u8_n2752 ) );
INV_X1 _u10_u8_U1450  ( .A(_u10_u8_n2752 ), .ZN(_u10_u8_n2421 ) );
NAND2_X1 _u10_u8_U1449  ( .A1(_u10_u8_n2421 ), .A2(_u10_u8_n2874 ), .ZN(_u10_u8_n2033 ) );
INV_X1 _u10_u8_U1448  ( .A(_u10_u8_n2033 ), .ZN(_u10_u8_n2742 ) );
NAND3_X1 _u10_u8_U1447  ( .A1(_u10_u8_n2305 ), .A2(_u10_u8_n1936 ), .A3(_u10_u8_n2742 ), .ZN(_u10_u8_n1896 ) );
OR3_X1 _u10_u8_U1446  ( .A1(_u10_u8_n2156 ), .A2(1'b0), .A3(_u10_u8_n1896 ),.ZN(_u10_u8_n2905 ) );
NAND2_X1 _u10_u8_U1445  ( .A1(_u10_u8_n2113 ), .A2(_u10_u8_n2996 ), .ZN(_u10_u8_n2719 ) );
NOR2_X1 _u10_u8_U1444  ( .A1(_u10_u8_n2719 ), .A2(1'b0), .ZN(_u10_u8_n2941 ));
INV_X1 _u10_u8_U1443  ( .A(_u10_u8_n2941 ), .ZN(_u10_u8_n2911 ) );
NOR2_X1 _u10_u8_U1442  ( .A1(_u10_u8_n2905 ), .A2(_u10_u8_n2911 ), .ZN(_u10_u8_n3222 ) );
INV_X1 _u10_u8_U1441  ( .A(_u10_u8_n3222 ), .ZN(_u10_u8_n2695 ) );
INV_X1 _u10_u8_U1440  ( .A(_u10_u8_n2156 ), .ZN(_u10_u8_n2089 ) );
NAND3_X1 _u10_u8_U1439  ( .A1(_u10_u8_n2089 ), .A2(_u10_u8_n2446 ), .A3(_u10_u8_n3180 ), .ZN(_u10_u8_n2902 ) );
NOR2_X1 _u10_u8_U1438  ( .A1(_u10_u8_n2902 ), .A2(_u10_u8_n2911 ), .ZN(_u10_u8_n2533 ) );
INV_X1 _u10_u8_U1437  ( .A(_u10_u8_n2533 ), .ZN(_u10_u8_n2485 ) );
NAND2_X1 _u10_u8_U1436  ( .A1(_u10_u8_n2695 ), .A2(_u10_u8_n2485 ), .ZN(_u10_u8_n2721 ) );
NAND2_X1 _u10_u8_U1435  ( .A1(1'b0), .A2(_u10_u8_n2113 ), .ZN(_u10_u8_n1868 ) );
INV_X1 _u10_u8_U1434  ( .A(_u10_u8_n1868 ), .ZN(_u10_u8_n2534 ) );
NOR2_X1 _u10_u8_U1433  ( .A1(_u10_u8_n2721 ), .A2(_u10_u8_n2534 ), .ZN(_u10_u8_n3231 ) );
NAND2_X1 _u10_u8_U1432  ( .A1(_u10_u8_n2467 ), .A2(_u10_u8_n3001 ), .ZN(_u10_u8_n2303 ) );
INV_X1 _u10_u8_U1431  ( .A(_u10_u8_n2303 ), .ZN(_u10_u8_n2549 ) );
INV_X1 _u10_u8_U1430  ( .A(1'b0), .ZN(_u10_u8_n2803 ) );
NAND2_X1 _u10_u8_U1429  ( .A1(_u10_u8_n2803 ), .A2(_u10_u8_n2446 ), .ZN(_u10_u8_n1846 ) );
INV_X1 _u10_u8_U1428  ( .A(_u10_u8_n1846 ), .ZN(_u10_u8_n2667 ) );
NAND3_X1 _u10_u8_U1427  ( .A1(_u10_u8_n2549 ), .A2(_u10_u8_n2667 ), .A3(1'b0), .ZN(_u10_u8_n2739 ) );
INV_X1 _u10_u8_U1426  ( .A(_u10_u8_n2739 ), .ZN(_u10_u8_n3272 ) );
INV_X1 _u10_u8_U1425  ( .A(_u10_u8_n2719 ), .ZN(_u10_u8_n2364 ) );
NAND2_X1 _u10_u8_U1424  ( .A1(_u10_u8_n3272 ), .A2(_u10_u8_n2364 ), .ZN(_u10_u8_n2852 ) );
INV_X1 _u10_u8_U1423  ( .A(_u10_u8_n2852 ), .ZN(_u10_u8_n2214 ) );
NAND2_X1 _u10_u8_U1422  ( .A1(_u10_u8_n2875 ), .A2(_u10_u8_n2089 ), .ZN(_u10_u8_n2097 ) );
INV_X1 _u10_u8_U1421  ( .A(_u10_u8_n2097 ), .ZN(_u10_u8_n2300 ) );
NAND2_X1 _u10_u8_U1420  ( .A1(_u10_u8_n2300 ), .A2(_u10_u8_n2446 ), .ZN(_u10_u8_n2001 ) );
NOR2_X1 _u10_u8_U1419  ( .A1(_u10_u8_n2001 ), .A2(_u10_u8_n2911 ), .ZN(_u10_u8_n2877 ) );
NOR2_X1 _u10_u8_U1418  ( .A1(_u10_u8_n2214 ), .A2(_u10_u8_n2877 ), .ZN(_u10_u8_n2940 ) );
NAND2_X1 _u10_u8_U1417  ( .A1(_u10_u8_n3231 ), .A2(_u10_u8_n2940 ), .ZN(_u10_u8_n3408 ) );
NAND2_X1 _u10_u8_U1416  ( .A1(_u10_u8_n2190 ), .A2(_u10_u8_n3408 ), .ZN(_u10_u8_n3402 ) );
NOR2_X1 _u10_u8_U1415  ( .A1(_u10_u8_n2446 ), .A2(_u10_u8_n2911 ), .ZN(_u10_u8_n3059 ) );
NAND2_X1 _u10_u8_U1414  ( .A1(_u10_u8_n3059 ), .A2(_u10_u8_n2190 ), .ZN(_u10_u8_n3404 ) );
AND3_X1 _u10_u8_U1413  ( .A1(_u10_u8_n3407 ), .A2(_u10_u8_n3226 ), .A3(_u10_u8_n3115 ), .ZN(_u10_u8_n3058 ) );
NAND2_X1 _u10_u8_U1412  ( .A1(_u10_u8_n3058 ), .A2(_u10_u8_n2022 ), .ZN(_u10_u8_n3406 ) );
NAND2_X1 _u10_u8_U1411  ( .A1(_u10_u8_n1853 ), .A2(_u10_u8_n3406 ), .ZN(_u10_u8_n3405 ) );
AND3_X1 _u10_u8_U1410  ( .A1(_u10_u8_n3404 ), .A2(_u10_u8_n1965 ), .A3(_u10_u8_n3405 ), .ZN(_u10_u8_n3063 ) );
NAND2_X1 _u10_u8_U1409  ( .A1(_u10_u8_n2667 ), .A2(_u10_u8_n3001 ), .ZN(_u10_u8_n1898 ) );
INV_X1 _u10_u8_U1408  ( .A(_u10_u8_n1898 ), .ZN(_u10_u8_n2835 ) );
NAND3_X1 _u10_u8_U1407  ( .A1(_u10_u8_n2364 ), .A2(_u10_u8_n2835 ), .A3(1'b0), .ZN(_u10_u8_n1869 ) );
NOR2_X1 _u10_u8_U1406  ( .A1(_u10_u8_n1869 ), .A2(_u10_u8_n2531 ), .ZN(_u10_u8_n2761 ) );
NOR3_X1 _u10_u8_U1405  ( .A1(_u10_u8_n2761 ), .A2(_u10_u8_n2528 ), .A3(_u10_u8_n2054 ), .ZN(_u10_u8_n3403 ) );
NAND4_X1 _u10_u8_U1404  ( .A1(_u10_u8_n3401 ), .A2(_u10_u8_n3402 ), .A3(_u10_u8_n3063 ), .A4(_u10_u8_n3403 ), .ZN(_u10_u8_n3400 ) );
NAND2_X1 _u10_u8_U1403  ( .A1(_u10_u8_n1966 ), .A2(_u10_u8_n3400 ), .ZN(_u10_u8_n3381 ) );
AND2_X1 _u10_u8_U1402  ( .A1(_u10_u8_n3368 ), .A2(_u10_SYNOPSYS_UNCONNECTED_38 ), .ZN(_u10_u8_n3319 ) );
NAND2_X1 _u10_u8_U1401  ( .A1(_u10_u8_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_37 ), .ZN(_u10_u8_n1849 ) );
INV_X1 _u10_u8_U1400  ( .A(_u10_u8_n1849 ), .ZN(_u10_u8_n2183 ) );
NAND2_X1 _u10_u8_U1399  ( .A1(_u10_u8_n2884 ), .A2(_u10_u8_n2183 ), .ZN(_u10_u8_n2883 ) );
INV_X1 _u10_u8_U1398  ( .A(_u10_u8_n2883 ), .ZN(_u10_u8_n1890 ) );
INV_X1 _u10_u8_U1397  ( .A(_u10_u8_n2940 ), .ZN(_u10_u8_n3278 ) );
NAND2_X1 _u10_u8_U1396  ( .A1(_u10_u8_n1890 ), .A2(_u10_u8_n3278 ), .ZN(_u10_u8_n3382 ) );
NAND2_X1 _u10_u8_U1395  ( .A1(_u10_u8_n3059 ), .A2(_u10_u8_n2669 ), .ZN(_u10_u8_n3399 ) );
NAND2_X1 _u10_u8_U1394  ( .A1(_u10_u8_n2031 ), .A2(_u10_u8_n3399 ), .ZN(_u10_u8_n3398 ) );
NAND2_X1 _u10_u8_U1393  ( .A1(_u10_u8_n2162 ), .A2(_u10_u8_n3398 ), .ZN(_u10_u8_n3395 ) );
NAND3_X1 _u10_u8_U1392  ( .A1(_u10_u8_n2747 ), .A2(_u10_u8_n2078 ), .A3(_u10_u8_n3126 ), .ZN(_u10_u8_n3396 ) );
NAND2_X1 _u10_u8_U1391  ( .A1(_u10_u8_n2055 ), .A2(_u10_u8_n2036 ), .ZN(_u10_u8_n2285 ) );
NOR2_X1 _u10_u8_U1390  ( .A1(_u10_u8_n2285 ), .A2(_u10_u8_n2030 ), .ZN(_u10_u8_n3349 ) );
INV_X1 _u10_u8_U1389  ( .A(_u10_u8_n3349 ), .ZN(_u10_u8_n1933 ) );
INV_X1 _u10_u8_U1388  ( .A(_u10_u8_n2710 ), .ZN(_u10_u8_n3397 ) );
NAND4_X1 _u10_u8_U1387  ( .A1(_u10_u8_n3395 ), .A2(_u10_u8_n3396 ), .A3(_u10_u8_n1933 ), .A4(_u10_u8_n3397 ), .ZN(_u10_u8_n3389 ) );
NAND2_X1 _u10_u8_U1386  ( .A1(_u10_u8_n1936 ), .A2(_u10_u8_n2828 ), .ZN(_u10_u8_n3141 ) );
INV_X1 _u10_u8_U1385  ( .A(_u10_u8_n3141 ), .ZN(_u10_u8_n2302 ) );
NAND2_X1 _u10_u8_U1384  ( .A1(_u10_u8_n3394 ), .A2(_u10_u8_n2302 ), .ZN(_u10_u8_n3390 ) );
NOR2_X1 _u10_u8_U1383  ( .A1(_u10_u8_n1869 ), .A2(_u10_u8_n2274 ), .ZN(_u10_u8_n3378 ) );
INV_X1 _u10_u8_U1382  ( .A(_u10_u8_n3378 ), .ZN(_u10_u8_n2748 ) );
NOR2_X1 _u10_u8_U1381  ( .A1(1'b0), .A2(_u10_u8_n2748 ), .ZN(_u10_u8_n3391 ));
NAND2_X1 _u10_u8_U1380  ( .A1(_u10_u8_n2534 ), .A2(_u10_u8_n2669 ), .ZN(_u10_u8_n2383 ) );
INV_X1 _u10_u8_U1379  ( .A(_u10_u8_n2383 ), .ZN(_u10_u8_n1978 ) );
NAND2_X1 _u10_u8_U1378  ( .A1(_u10_u8_n1978 ), .A2(_u10_u8_n2874 ), .ZN(_u10_u8_n3392 ) );
INV_X1 _u10_u8_U1377  ( .A(_u10_u8_n2411 ), .ZN(_u10_u8_n2164 ) );
NAND4_X1 _u10_u8_U1376  ( .A1(_u10_u8_n3392 ), .A2(_u10_u8_n3393 ), .A3(_u10_u8_n2033 ), .A4(_u10_u8_n2164 ), .ZN(_u10_u8_n2476 ) );
NOR4_X1 _u10_u8_U1375  ( .A1(_u10_u8_n3389 ), .A2(_u10_u8_n3390 ), .A3(_u10_u8_n3391 ), .A4(_u10_u8_n2476 ), .ZN(_u10_u8_n3388 ) );
NAND2_X1 _u10_u8_U1374  ( .A1(_u10_u8_n3236 ), .A2(_u10_u8_n3328 ), .ZN(_u10_u8_n2025 ) );
NOR2_X1 _u10_u8_U1373  ( .A1(_u10_u8_n3388 ), .A2(_u10_u8_n2025 ), .ZN(_u10_u8_n3384 ) );
NOR2_X1 _u10_u8_U1372  ( .A1(1'b0), .A2(1'b0), .ZN(_u10_u8_n2152 ) );
NAND2_X1 _u10_u8_U1371  ( .A1(_u10_u8_n2152 ), .A2(_u10_u8_n2175 ), .ZN(_u10_u8_n2722 ) );
INV_X1 _u10_u8_U1370  ( .A(_u10_u8_n2722 ), .ZN(_u10_u8_n2588 ) );
NAND2_X1 _u10_u8_U1369  ( .A1(_u10_u8_n2549 ), .A2(_u10_u8_n3349 ), .ZN(_u10_u8_n2091 ) );
NOR2_X1 _u10_u8_U1368  ( .A1(_u10_u8_n2091 ), .A2(_u10_u8_n1846 ), .ZN(_u10_u8_n2128 ) );
NAND3_X1 _u10_u8_U1367  ( .A1(_u10_u8_n3066 ), .A2(_u10_u8_n2113 ), .A3(_u10_u8_n2128 ), .ZN(_u10_u8_n2342 ) );
INV_X1 _u10_u8_U1366  ( .A(_u10_u8_n2342 ), .ZN(_u10_u8_n3316 ) );
NAND2_X1 _u10_u8_U1365  ( .A1(_u10_u8_n2588 ), .A2(_u10_u8_n3316 ), .ZN(_u10_u8_n2142 ) );
NOR2_X1 _u10_u8_U1364  ( .A1(_u10_u8_n1954 ), .A2(_u10_u8_n1898 ), .ZN(_u10_u8_n2255 ) );
NAND2_X1 _u10_u8_U1363  ( .A1(_u10_u8_n2255 ), .A2(_u10_u8_n2996 ), .ZN(_u10_u8_n1915 ) );
INV_X1 _u10_u8_U1362  ( .A(_u10_u8_n1915 ), .ZN(_u10_u8_n2251 ) );
NAND2_X1 _u10_u8_U1361  ( .A1(_u10_u8_n2251 ), .A2(_u10_u8_n2113 ), .ZN(_u10_u8_n1925 ) );
INV_X1 _u10_u8_U1360  ( .A(_u10_u8_n2026 ), .ZN(_u10_u8_n3340 ) );
NOR3_X1 _u10_u8_U1359  ( .A1(_u10_u8_n1925 ), .A2(_u10_u8_n2216 ), .A3(_u10_u8_n3340 ), .ZN(_u10_u8_n2003 ) );
INV_X1 _u10_u8_U1358  ( .A(1'b0), .ZN(_u10_u8_n1930 ) );
NAND2_X1 _u10_u8_U1357  ( .A1(_u10_u8_n2003 ), .A2(_u10_u8_n1930 ), .ZN(_u10_u8_n3387 ) );
AND2_X1 _u10_u8_U1356  ( .A1(_u10_u8_n2142 ), .A2(_u10_u8_n3387 ), .ZN(_u10_u8_n3366 ) );
NOR3_X1 _u10_u8_U1355  ( .A1(_u10_u8_n1813 ), .A2(_u10_u8_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_34 ), .ZN(_u10_u8_n3360 ) );
NOR2_X1 _u10_u8_U1354  ( .A1(_u10_SYNOPSYS_UNCONNECTED_36 ), .A2(_u10_SYNOPSYS_UNCONNECTED_37 ), .ZN(_u10_u8_n3136 ) );
NAND2_X1 _u10_u8_U1353  ( .A1(_u10_u8_n3360 ), .A2(_u10_u8_n3136 ), .ZN(_u10_u8_n2344 ) );
NOR2_X1 _u10_u8_U1352  ( .A1(_u10_u8_n3366 ), .A2(_u10_u8_n2344 ), .ZN(_u10_u8_n3385 ) );
NOR3_X1 _u10_u8_U1351  ( .A1(_u10_SYNOPSYS_UNCONNECTED_34 ), .A2(_u10_u8_n1816 ), .A3(_u10_SYNOPSYS_UNCONNECTED_38 ), .ZN(_u10_u8_n3342 ) );
NAND2_X1 _u10_u8_U1350  ( .A1(_u10_u8_n3342 ), .A2(_u10_u8_n3136 ), .ZN(_u10_u8_n2584 ) );
NOR2_X1 _u10_u8_U1349  ( .A1(_u10_u8_n2584 ), .A2(1'b0), .ZN(_u10_u8_n2139 ));
INV_X1 _u10_u8_U1348  ( .A(_u10_u8_n2216 ), .ZN(_u10_u8_n2106 ) );
AND2_X1 _u10_u8_U1347  ( .A1(_u10_u8_n2152 ), .A2(_u10_u8_n2106 ), .ZN(_u10_u8_n2336 ) );
NAND2_X1 _u10_u8_U1346  ( .A1(_u10_u8_n2139 ), .A2(_u10_u8_n2336 ), .ZN(_u10_u8_n2365 ) );
INV_X1 _u10_u8_U1345  ( .A(_u10_u8_n2365 ), .ZN(_u10_u8_n2004 ) );
AND2_X1 _u10_u8_U1344  ( .A1(_u10_u8_n2877 ), .A2(_u10_u8_n2004 ), .ZN(_u10_u8_n3386 ) );
NOR3_X1 _u10_u8_U1343  ( .A1(_u10_u8_n3384 ), .A2(_u10_u8_n3385 ), .A3(_u10_u8_n3386 ), .ZN(_u10_u8_n3383 ) );
NAND4_X1 _u10_u8_U1342  ( .A1(_u10_u8_n3380 ), .A2(_u10_u8_n3381 ), .A3(_u10_u8_n3382 ), .A4(_u10_u8_n3383 ), .ZN(_u10_u8_n3191 ) );
NAND2_X1 _u10_u8_U1341  ( .A1(_u10_u8_n2285 ), .A2(_u10_u8_n3379 ), .ZN(_u10_u8_n1975 ) );
NOR3_X1 _u10_u8_U1340  ( .A1(_u10_u8_n3378 ), .A2(1'b0), .A3(_u10_u8_n1975 ),.ZN(_u10_u8_n3122 ) );
AND4_X1 _u10_u8_U1339  ( .A1(_u10_u8_n2752 ), .A2(_u10_u8_n2383 ), .A3(_u10_u8_n1969 ), .A4(_u10_u8_n3122 ), .ZN(_u10_u8_n3377 ) );
NOR2_X1 _u10_u8_U1338  ( .A1(_u10_u8_n1814 ), .A2(_u10_u8_n1815 ), .ZN(_u10_u8_n3147 ) );
NAND2_X1 _u10_u8_U1337  ( .A1(_u10_u8_n3328 ), .A2(_u10_u8_n3147 ), .ZN(_u10_u8_n2359 ) );
NOR2_X1 _u10_u8_U1336  ( .A1(_u10_u8_n3377 ), .A2(_u10_u8_n2359 ), .ZN(_u10_u8_n3362 ) );
INV_X1 _u10_u8_U1335  ( .A(_u10_u8_n2008 ), .ZN(_u10_u8_n3097 ) );
NOR3_X1 _u10_u8_U1334  ( .A1(_u10_SYNOPSYS_UNCONNECTED_34 ), .A2(_u10_u8_n1813 ), .A3(_u10_SYNOPSYS_UNCONNECTED_35 ), .ZN(_u10_u8_n3269 ) );
NAND2_X1 _u10_u8_U1333  ( .A1(_u10_u8_n3269 ), .A2(_u10_u8_n3136 ), .ZN(_u10_u8_n3109 ) );
INV_X1 _u10_u8_U1332  ( .A(_u10_u8_n3109 ), .ZN(_u10_u8_n2999 ) );
INV_X1 _u10_u8_U1331  ( .A(_u10_u8_n2508 ), .ZN(_u10_u8_n2103 ) );
NAND2_X1 _u10_u8_U1330  ( .A1(_u10_u8_n2336 ), .A2(_u10_u8_n2103 ), .ZN(_u10_u8_n2249 ) );
NOR2_X1 _u10_u8_U1329  ( .A1(_u10_u8_n2249 ), .A2(1'b0), .ZN(_u10_u8_n1866 ));
NAND2_X1 _u10_u8_U1328  ( .A1(_u10_u8_n1866 ), .A2(_u10_u8_n1922 ), .ZN(_u10_u8_n2632 ) );
INV_X1 _u10_u8_U1327  ( .A(_u10_u8_n2223 ), .ZN(_u10_u8_n1918 ) );
NOR2_X1 _u10_u8_U1326  ( .A1(_u10_u8_n2632 ), .A2(_u10_u8_n1918 ), .ZN(_u10_u8_n1981 ) );
NAND3_X1 _u10_u8_U1325  ( .A1(_u10_u8_n3097 ), .A2(_u10_u8_n2999 ), .A3(_u10_u8_n1981 ), .ZN(_u10_u8_n3034 ) );
NOR3_X1 _u10_u8_U1324  ( .A1(_u10_SYNOPSYS_UNCONNECTED_35 ), .A2(_u10_SYNOPSYS_UNCONNECTED_34 ), .A3(_u10_SYNOPSYS_UNCONNECTED_38 ),.ZN(_u10_u8_n3302 ) );
NAND2_X1 _u10_u8_U1323  ( .A1(_u10_u8_n3302 ), .A2(_u10_u8_n3174 ), .ZN(_u10_u8_n3162 ) );
INV_X1 _u10_u8_U1322  ( .A(_u10_u8_n3162 ), .ZN(_u10_u8_n2979 ) );
NAND2_X1 _u10_u8_U1321  ( .A1(_u10_u8_n2979 ), .A2(_u10_u8_n2972 ), .ZN(_u10_u8_n1984 ) );
AND2_X1 _u10_u8_U1320  ( .A1(_u10_u8_n3302 ), .A2(_u10_u8_n3136 ), .ZN(_u10_u8_n2977 ) );
NAND3_X1 _u10_u8_U1319  ( .A1(_u10_u8_n2977 ), .A2(_u10_u8_n3000 ), .A3(_u10_u8_n3097 ), .ZN(_u10_u8_n3376 ) );
NAND2_X1 _u10_u8_U1318  ( .A1(_u10_u8_n1984 ), .A2(_u10_u8_n3376 ), .ZN(_u10_u8_n3375 ) );
NAND2_X1 _u10_u8_U1317  ( .A1(_u10_u8_n1981 ), .A2(_u10_u8_n3375 ), .ZN(_u10_u8_n2798 ) );
NAND2_X1 _u10_u8_U1316  ( .A1(_u10_u8_n3034 ), .A2(_u10_u8_n2798 ), .ZN(_u10_u8_n2007 ) );
NAND2_X1 _u10_u8_U1315  ( .A1(_u10_u8_n3269 ), .A2(_u10_u8_n3147 ), .ZN(_u10_u8_n2102 ) );
NOR2_X1 _u10_u8_U1314  ( .A1(_u10_u8_n2249 ), .A2(_u10_u8_n2102 ), .ZN(_u10_u8_n3323 ) );
INV_X1 _u10_u8_U1313  ( .A(_u10_u8_n3323 ), .ZN(_u10_u8_n3374 ) );
INV_X1 _u10_u8_U1312  ( .A(_u10_u8_n2344 ), .ZN(_u10_u8_n2002 ) );
NAND2_X1 _u10_u8_U1311  ( .A1(_u10_u8_n2336 ), .A2(_u10_u8_n2002 ), .ZN(_u10_u8_n3225 ) );
NAND2_X1 _u10_u8_U1310  ( .A1(_u10_u8_n3374 ), .A2(_u10_u8_n3225 ), .ZN(_u10_u8_n2488 ) );
NAND2_X1 _u10_u8_U1309  ( .A1(_u10_u8_n3342 ), .A2(_u10_u8_n3236 ), .ZN(_u10_u8_n2253 ) );
NOR2_X1 _u10_u8_U1308  ( .A1(_u10_u8_n2253 ), .A2(1'b0), .ZN(_u10_u8_n1885 ));
NAND2_X1 _u10_u8_U1307  ( .A1(_u10_u8_n3360 ), .A2(_u10_u8_n3174 ), .ZN(_u10_u8_n2254 ) );
INV_X1 _u10_u8_U1306  ( .A(_u10_u8_n2254 ), .ZN(_u10_u8_n2986 ) );
NAND2_X1 _u10_u8_U1305  ( .A1(_u10_u8_n2106 ), .A2(_u10_u8_n2986 ), .ZN(_u10_u8_n1913 ) );
INV_X1 _u10_u8_U1304  ( .A(_u10_u8_n1913 ), .ZN(_u10_u8_n2377 ) );
OR4_X1 _u10_u8_U1303  ( .A1(_u10_u8_n2007 ), .A2(_u10_u8_n2488 ), .A3(_u10_u8_n1885 ), .A4(_u10_u8_n2377 ), .ZN(_u10_u8_n3373 ) );
NAND2_X1 _u10_u8_U1302  ( .A1(_u10_u8_n2534 ), .A2(_u10_u8_n3373 ), .ZN(_u10_u8_n3370 ) );
NAND2_X1 _u10_u8_U1301  ( .A1(_u10_u8_n3342 ), .A2(_u10_u8_n3174 ), .ZN(_u10_u8_n2037 ) );
NAND2_X1 _u10_u8_U1300  ( .A1(_u10_u8_n2037 ), .A2(_u10_u8_n2254 ), .ZN(_u10_u8_n3372 ) );
NAND2_X1 _u10_u8_U1299  ( .A1(_u10_u8_n2003 ), .A2(_u10_u8_n3372 ), .ZN(_u10_u8_n3371 ) );
NAND2_X1 _u10_u8_U1298  ( .A1(_u10_u8_n3370 ), .A2(_u10_u8_n3371 ), .ZN(_u10_u8_n3363 ) );
NOR2_X1 _u10_u8_U1297  ( .A1(_u10_u8_n2490 ), .A2(_u10_u8_n1961 ), .ZN(_u10_u8_n3369 ) );
NAND2_X1 _u10_u8_U1296  ( .A1(_u10_u8_n2534 ), .A2(_u10_u8_n2049 ), .ZN(_u10_u8_n2646 ) );
INV_X1 _u10_u8_U1295  ( .A(_u10_u8_n2646 ), .ZN(_u10_u8_n3055 ) );
NOR2_X1 _u10_u8_U1294  ( .A1(_u10_u8_n3369 ), .A2(_u10_u8_n3055 ), .ZN(_u10_u8_n3367 ) );
NAND2_X1 _u10_u8_U1293  ( .A1(_u10_u8_n3368 ), .A2(_u10_u8_n3147 ), .ZN(_u10_u8_n2495 ) );
NOR2_X1 _u10_u8_U1292  ( .A1(_u10_u8_n3367 ), .A2(_u10_u8_n2495 ), .ZN(_u10_u8_n3364 ) );
INV_X1 _u10_u8_U1291  ( .A(_u10_u8_n2139 ), .ZN(_u10_u8_n3254 ) );
NOR2_X1 _u10_u8_U1290  ( .A1(_u10_u8_n3366 ), .A2(_u10_u8_n3254 ), .ZN(_u10_u8_n3365 ) );
NOR4_X1 _u10_u8_U1289  ( .A1(_u10_u8_n3362 ), .A2(_u10_u8_n3363 ), .A3(_u10_u8_n3364 ), .A4(_u10_u8_n3365 ), .ZN(_u10_u8_n3305 ) );
NAND2_X1 _u10_u8_U1288  ( .A1(_u10_u8_n3302 ), .A2(_u10_u8_n3147 ), .ZN(_u10_u8_n2980 ) );
NAND2_X1 _u10_u8_U1287  ( .A1(_u10_u8_n2102 ), .A2(_u10_u8_n2980 ), .ZN(_u10_u8_n2177 ) );
NAND2_X1 _u10_u8_U1286  ( .A1(_u10_u8_n2003 ), .A2(_u10_u8_n2493 ), .ZN(_u10_u8_n1962 ) );
NAND2_X1 _u10_u8_U1285  ( .A1(_u10_u8_n1961 ), .A2(_u10_u8_n1962 ), .ZN(_u10_u8_n3361 ) );
NAND2_X1 _u10_u8_U1284  ( .A1(_u10_u8_n2177 ), .A2(_u10_u8_n3361 ), .ZN(_u10_u8_n3357 ) );
NAND2_X1 _u10_u8_U1283  ( .A1(_u10_u8_n3236 ), .A2(_u10_u8_n3360 ), .ZN(_u10_u8_n1859 ) );
INV_X1 _u10_u8_U1282  ( .A(_u10_u8_n1859 ), .ZN(_u10_u8_n2256 ) );
NAND3_X1 _u10_u8_U1281  ( .A1(_u10_u8_n2256 ), .A2(_u10_u8_n2113 ), .A3(_u10_u8_n2128 ), .ZN(_u10_u8_n3358 ) );
NOR2_X1 _u10_u8_U1280  ( .A1(_u10_u8_n2877 ), .A2(_u10_u8_n3222 ), .ZN(_u10_u8_n3347 ) );
NAND2_X1 _u10_u8_U1279  ( .A1(_u10_u8_n3347 ), .A2(_u10_u8_n1869 ), .ZN(_u10_u8_n2005 ) );
NAND2_X1 _u10_u8_U1278  ( .A1(_u10_u8_n2488 ), .A2(_u10_u8_n2005 ), .ZN(_u10_u8_n3359 ) );
NAND3_X1 _u10_u8_U1277  ( .A1(_u10_u8_n3357 ), .A2(_u10_u8_n3358 ), .A3(_u10_u8_n3359 ), .ZN(_u10_u8_n3352 ) );
NAND2_X1 _u10_u8_U1276  ( .A1(_u10_u8_n3320 ), .A2(_u10_u8_n3136 ), .ZN(_u10_u8_n2356 ) );
INV_X1 _u10_u8_U1275  ( .A(_u10_u8_n2356 ), .ZN(_u10_u8_n2830 ) );
NAND2_X1 _u10_u8_U1274  ( .A1(_u10_u8_n2830 ), .A2(_u10_u8_n2836 ), .ZN(_u10_u8_n2291 ) );
NOR3_X1 _u10_u8_U1273  ( .A1(_u10_u8_n2291 ), .A2(_u10_u8_n2330 ), .A3(_u10_u8_n2022 ), .ZN(_u10_u8_n3353 ) );
INV_X1 _u10_u8_U1272  ( .A(_u10_u8_n1925 ), .ZN(_u10_u8_n2105 ) );
AND2_X1 _u10_u8_U1271  ( .A1(_u10_u8_n2108 ), .A2(_u10_u8_n2105 ), .ZN(_u10_u8_n2915 ) );
INV_X1 _u10_u8_U1270  ( .A(_u10_u8_n2330 ), .ZN(_u10_u8_n2107 ) );
NAND2_X1 _u10_u8_U1269  ( .A1(_u10_u8_n2915 ), .A2(_u10_u8_n2107 ), .ZN(_u10_u8_n2203 ) );
INV_X1 _u10_u8_U1268  ( .A(_u10_u8_n2203 ), .ZN(_u10_u8_n1982 ) );
NAND2_X1 _u10_u8_U1267  ( .A1(_u10_u8_n1982 ), .A2(_u10_u8_n2536 ), .ZN(_u10_u8_n2587 ) );
INV_X1 _u10_u8_U1266  ( .A(_u10_u8_n2587 ), .ZN(_u10_u8_n2697 ) );
NAND3_X1 _u10_u8_U1265  ( .A1(_u10_u8_n2697 ), .A2(_u10_u8_n2493 ), .A3(_u10_u8_n2377 ), .ZN(_u10_u8_n2412 ) );
INV_X1 _u10_u8_U1264  ( .A(_u10_u8_n2412 ), .ZN(_u10_u8_n3354 ) );
NAND2_X1 _u10_u8_U1263  ( .A1(_u10_u8_n3174 ), .A2(_u10_u8_n3269 ), .ZN(_u10_u8_n2375 ) );
INV_X1 _u10_u8_U1262  ( .A(_u10_u8_n2375 ), .ZN(_u10_u8_n2507 ) );
NAND2_X1 _u10_u8_U1261  ( .A1(_u10_u8_n1981 ), .A2(_u10_u8_n2507 ), .ZN(_u10_u8_n2621 ) );
NOR4_X1 _u10_u8_U1260  ( .A1(1'b0), .A2(_u10_u8_n3356 ), .A3(_u10_u8_n2203 ),.A4(_u10_u8_n2621 ), .ZN(_u10_u8_n3355 ) );
NOR4_X1 _u10_u8_U1259  ( .A1(_u10_u8_n3352 ), .A2(_u10_u8_n3353 ), .A3(_u10_u8_n3354 ), .A4(_u10_u8_n3355 ), .ZN(_u10_u8_n3306 ) );
NOR2_X1 _u10_u8_U1258  ( .A1(_u10_u8_n2842 ), .A2(_u10_u8_n2356 ), .ZN(_u10_u8_n1891 ) );
INV_X1 _u10_u8_U1257  ( .A(_u10_u8_n1869 ), .ZN(_u10_u8_n2885 ) );
NAND2_X1 _u10_u8_U1256  ( .A1(_u10_u8_n1891 ), .A2(_u10_u8_n2885 ), .ZN(_u10_u8_n3330 ) );
NAND2_X1 _u10_u8_U1255  ( .A1(_u10_u8_n2761 ), .A2(_u10_u8_n2837 ), .ZN(_u10_u8_n3351 ) );
NAND3_X1 _u10_u8_U1254  ( .A1(_u10_u8_n2884 ), .A2(_u10_u8_n2080 ), .A3(_u10_u8_n2915 ), .ZN(_u10_u8_n2762 ) );
NAND2_X1 _u10_u8_U1253  ( .A1(_u10_u8_n2055 ), .A2(_u10_u8_n2019 ), .ZN(_u10_u8_n3259 ) );
NAND4_X1 _u10_u8_U1252  ( .A1(_u10_u8_n3351 ), .A2(_u10_u8_n2762 ), .A3(_u10_u8_n2061 ), .A4(_u10_u8_n3259 ), .ZN(_u10_u8_n3350 ) );
NAND2_X1 _u10_u8_U1251  ( .A1(_u10_u8_n2183 ), .A2(_u10_u8_n3350 ), .ZN(_u10_u8_n3331 ) );
NAND2_X1 _u10_u8_U1250  ( .A1(_u10_u8_n3349 ), .A2(_u10_u8_n2305 ), .ZN(_u10_u8_n3348 ) );
NAND2_X1 _u10_u8_U1249  ( .A1(_u10_u8_n1896 ), .A2(_u10_u8_n3348 ), .ZN(_u10_u8_n3176 ) );
NAND2_X1 _u10_u8_U1248  ( .A1(_u10_u8_n2461 ), .A2(_u10_u8_n3176 ), .ZN(_u10_u8_n3332 ) );
INV_X1 _u10_u8_U1247  ( .A(_u10_u8_n2495 ), .ZN(_u10_u8_n2063 ) );
NAND2_X1 _u10_u8_U1246  ( .A1(_u10_u8_n2049 ), .A2(_u10_u8_n2063 ), .ZN(_u10_u8_n2886 ) );
NOR2_X1 _u10_u8_U1245  ( .A1(_u10_u8_n3347 ), .A2(_u10_u8_n2886 ), .ZN(_u10_u8_n3334 ) );
NAND2_X1 _u10_u8_U1244  ( .A1(1'b0), .A2(_u10_u8_n2835 ), .ZN(_u10_u8_n3344 ) );
NAND2_X1 _u10_u8_U1243  ( .A1(_u10_u8_n2001 ), .A2(_u10_u8_n2905 ), .ZN(_u10_u8_n3346 ) );
NAND2_X1 _u10_u8_U1242  ( .A1(_u10_u8_n3346 ), .A2(_u10_u8_n2803 ), .ZN(_u10_u8_n3345 ) );
NAND2_X1 _u10_u8_U1241  ( .A1(_u10_u8_n2087 ), .A2(_u10_u8_n2835 ), .ZN(_u10_u8_n2413 ) );
INV_X1 _u10_u8_U1240  ( .A(_u10_u8_n2128 ), .ZN(_u10_u8_n2235 ) );
NAND4_X1 _u10_u8_U1239  ( .A1(_u10_u8_n3344 ), .A2(_u10_u8_n3345 ), .A3(_u10_u8_n2413 ), .A4(_u10_u8_n2235 ), .ZN(_u10_u8_n3329 ) );
NOR2_X1 _u10_u8_U1238  ( .A1(_u10_u8_n1915 ), .A2(_u10_u8_n3340 ), .ZN(_u10_u8_n3343 ) );
NOR3_X1 _u10_u8_U1237  ( .A1(_u10_u8_n3329 ), .A2(1'b0), .A3(_u10_u8_n3343 ),.ZN(_u10_u8_n3341 ) );
NAND2_X1 _u10_u8_U1236  ( .A1(_u10_u8_n3342 ), .A2(_u10_u8_n3147 ), .ZN(_u10_u8_n2688 ) );
NOR2_X1 _u10_u8_U1235  ( .A1(_u10_u8_n3341 ), .A2(_u10_u8_n2688 ), .ZN(_u10_u8_n3335 ) );
NOR2_X1 _u10_u8_U1234  ( .A1(_u10_u8_n2256 ), .A2(_u10_u8_n1885 ), .ZN(_u10_u8_n2689 ) );
NOR2_X1 _u10_u8_U1233  ( .A1(1'b0), .A2(_u10_u8_n2413 ), .ZN(_u10_u8_n3338 ));
NOR2_X1 _u10_u8_U1232  ( .A1(_u10_u8_n1925 ), .A2(_u10_u8_n3340 ), .ZN(_u10_u8_n3339 ) );
NOR3_X1 _u10_u8_U1231  ( .A1(_u10_u8_n2005 ), .A2(_u10_u8_n3338 ), .A3(_u10_u8_n3339 ), .ZN(_u10_u8_n3337 ) );
NOR2_X1 _u10_u8_U1230  ( .A1(_u10_u8_n2689 ), .A2(_u10_u8_n3337 ), .ZN(_u10_u8_n3336 ) );
NOR3_X1 _u10_u8_U1229  ( .A1(_u10_u8_n3334 ), .A2(_u10_u8_n3335 ), .A3(_u10_u8_n3336 ), .ZN(_u10_u8_n3333 ) );
NAND4_X1 _u10_u8_U1228  ( .A1(_u10_u8_n3330 ), .A2(_u10_u8_n3331 ), .A3(_u10_u8_n3332 ), .A4(_u10_u8_n3333 ), .ZN(_u10_u8_n3308 ) );
NAND3_X1 _u10_u8_U1227  ( .A1(_u10_SYNOPSYS_UNCONNECTED_38 ), .A2(_u10_SYNOPSYS_UNCONNECTED_35 ), .A3(_u10_u8_n3147 ), .ZN(_u10_u8_n2126 ) );
INV_X1 _u10_u8_U1226  ( .A(_u10_u8_n2126 ), .ZN(_u10_u8_n2329 ) );
NAND2_X1 _u10_u8_U1225  ( .A1(_u10_u8_n2329 ), .A2(_u10_u8_n3329 ), .ZN(_u10_u8_n3324 ) );
NAND2_X1 _u10_u8_U1224  ( .A1(_u10_u8_n3328 ), .A2(_u10_u8_n3136 ), .ZN(_u10_u8_n2000 ) );
INV_X1 _u10_u8_U1223  ( .A(_u10_u8_n2000 ), .ZN(_u10_u8_n2445 ) );
NAND3_X1 _u10_u8_U1222  ( .A1(_u10_u8_n2446 ), .A2(_u10_u8_n3001 ), .A3(_u10_u8_n2087 ), .ZN(_u10_u8_n3327 ) );
NAND2_X1 _u10_u8_U1221  ( .A1(_u10_u8_n3327 ), .A2(_u10_u8_n2905 ), .ZN(_u10_u8_n2500 ) );
NAND2_X1 _u10_u8_U1220  ( .A1(_u10_u8_n2445 ), .A2(_u10_u8_n2500 ), .ZN(_u10_u8_n3325 ) );
NAND2_X1 _u10_u8_U1219  ( .A1(1'b0), .A2(_u10_u8_n2979 ), .ZN(_u10_u8_n3326 ) );
NAND3_X1 _u10_u8_U1218  ( .A1(_u10_u8_n3324 ), .A2(_u10_u8_n3325 ), .A3(_u10_u8_n3326 ), .ZN(_u10_u8_n3309 ) );
AND2_X1 _u10_u8_U1217  ( .A1(_u10_u8_n2877 ), .A2(_u10_u8_n3223 ), .ZN(_u10_u8_n2858 ) );
NAND2_X1 _u10_u8_U1216  ( .A1(_u10_u8_n3319 ), .A2(_u10_SYNOPSYS_UNCONNECTED_36 ), .ZN(_u10_u8_n2346 ) );
INV_X1 _u10_u8_U1215  ( .A(_u10_u8_n2346 ), .ZN(_u10_u8_n2043 ) );
NAND2_X1 _u10_u8_U1214  ( .A1(_u10_u8_n2858 ), .A2(_u10_u8_n2043 ), .ZN(_u10_u8_n3321 ) );
NAND2_X1 _u10_u8_U1213  ( .A1(_u10_u8_n1982 ), .A2(_u10_u8_n2195 ), .ZN(_u10_u8_n3268 ) );
INV_X1 _u10_u8_U1212  ( .A(_u10_u8_n3268 ), .ZN(_u10_u8_n2222 ) );
NAND3_X1 _u10_u8_U1211  ( .A1(_u10_u8_n3323 ), .A2(_u10_u8_n3216 ), .A3(_u10_u8_n2222 ), .ZN(_u10_u8_n3322 ) );
NAND2_X1 _u10_u8_U1210  ( .A1(_u10_u8_n3321 ), .A2(_u10_u8_n3322 ), .ZN(_u10_u8_n2374 ) );
NAND2_X1 _u10_u8_U1209  ( .A1(_u10_u8_n3320 ), .A2(_u10_u8_n3174 ), .ZN(_u10_u8_n2014 ) );
NOR2_X1 _u10_u8_U1208  ( .A1(_u10_u8_n1841 ), .A2(_u10_u8_n2014 ), .ZN(_u10_u8_n2813 ) );
NAND2_X1 _u10_u8_U1207  ( .A1(_u10_u8_n2813 ), .A2(_u10_u8_n2534 ), .ZN(_u10_u8_n3310 ) );
NAND2_X1 _u10_u8_U1206  ( .A1(_u10_u8_n3319 ), .A2(_u10_u8_n3136 ), .ZN(_u10_u8_n1836 ) );
INV_X1 _u10_u8_U1205  ( .A(_u10_u8_n1836 ), .ZN(_u10_u8_n2815 ) );
NAND2_X1 _u10_u8_U1204  ( .A1(_u10_u8_n2534 ), .A2(_u10_u8_n3129 ), .ZN(_u10_u8_n2439 ) );
NAND2_X1 _u10_u8_U1203  ( .A1(_u10_u8_n2055 ), .A2(_u10_u8_n2107 ), .ZN(_u10_u8_n2062 ) );
NAND2_X1 _u10_u8_U1202  ( .A1(_u10_u8_n2439 ), .A2(_u10_u8_n2062 ), .ZN(_u10_u8_n3318 ) );
NAND2_X1 _u10_u8_U1201  ( .A1(_u10_u8_n2815 ), .A2(_u10_u8_n3318 ), .ZN(_u10_u8_n3311 ) );
NAND2_X1 _u10_u8_U1200  ( .A1(_u10_u8_n2986 ), .A2(_u10_u8_n2175 ), .ZN(_u10_u8_n3317 ) );
NAND2_X1 _u10_u8_U1199  ( .A1(_u10_u8_n2253 ), .A2(_u10_u8_n3317 ), .ZN(_u10_u8_n3157 ) );
NAND2_X1 _u10_u8_U1198  ( .A1(_u10_u8_n3316 ), .A2(_u10_u8_n3157 ), .ZN(_u10_u8_n3312 ) );
NOR2_X1 _u10_u8_U1197  ( .A1(_u10_u8_n2495 ), .A2(_u10_u8_n2194 ), .ZN(_u10_u8_n3314 ) );
NOR2_X1 _u10_u8_U1196  ( .A1(_u10_u8_n2375 ), .A2(_u10_u8_n2367 ), .ZN(_u10_u8_n3315 ) );
NOR2_X1 _u10_u8_U1195  ( .A1(_u10_u8_n3314 ), .A2(_u10_u8_n3315 ), .ZN(_u10_u8_n3313 ) );
NAND4_X1 _u10_u8_U1194  ( .A1(_u10_u8_n3310 ), .A2(_u10_u8_n3311 ), .A3(_u10_u8_n3312 ), .A4(_u10_u8_n3313 ), .ZN(_u10_u8_n2315 ) );
NOR4_X1 _u10_u8_U1193  ( .A1(_u10_u8_n3308 ), .A2(_u10_u8_n3309 ), .A3(_u10_u8_n2374 ), .A4(_u10_u8_n2315 ), .ZN(_u10_u8_n3307 ) );
NAND3_X1 _u10_u8_U1192  ( .A1(_u10_u8_n3305 ), .A2(_u10_u8_n3306 ), .A3(_u10_u8_n3307 ), .ZN(_u10_u8_n1987 ) );
AND2_X1 _u10_u8_U1191  ( .A1(1'b0), .A2(_u10_u8_n2977 ), .ZN(_u10_u8_n3240 ));
NAND2_X1 _u10_u8_U1190  ( .A1(_u10_u8_n1891 ), .A2(_u10_u8_n2534 ), .ZN(_u10_u8_n3303 ) );
NAND4_X1 _u10_u8_U1189  ( .A1(_u10_u8_n1982 ), .A2(_u10_u8_n2659 ), .A3(_u10_u8_n2256 ), .A4(_u10_u8_n2175 ), .ZN(_u10_u8_n3304 ) );
AND2_X1 _u10_u8_U1188  ( .A1(_u10_u8_n3303 ), .A2(_u10_u8_n3304 ), .ZN(_u10_u8_n2612 ) );
NAND2_X1 _u10_u8_U1187  ( .A1(_u10_u8_n3302 ), .A2(_u10_u8_n3236 ), .ZN(_u10_u8_n2985 ) );
OR2_X1 _u10_u8_U1186  ( .A1(_u10_u8_n2431 ), .A2(_u10_u8_n2985 ), .ZN(_u10_u8_n3299 ) );
OR2_X1 _u10_u8_U1185  ( .A1(_u10_u8_n2282 ), .A2(_u10_u8_n2359 ), .ZN(_u10_u8_n3300 ) );
NAND2_X1 _u10_u8_U1184  ( .A1(_u10_u8_n1890 ), .A2(_u10_u8_n2534 ), .ZN(_u10_u8_n3301 ) );
NAND4_X1 _u10_u8_U1183  ( .A1(_u10_u8_n2612 ), .A2(_u10_u8_n3299 ), .A3(_u10_u8_n3300 ), .A4(_u10_u8_n3301 ), .ZN(_u10_u8_n3279 ) );
INV_X1 _u10_u8_U1182  ( .A(_u10_u8_n2464 ), .ZN(_u10_u8_n3295 ) );
NAND2_X1 _u10_u8_U1181  ( .A1(_u10_u8_n3295 ), .A2(_u10_u8_n2835 ), .ZN(_u10_u8_n2623 ) );
INV_X1 _u10_u8_U1180  ( .A(_u10_u8_n2623 ), .ZN(_u10_u8_n3185 ) );
INV_X1 _u10_u8_U1179  ( .A(_u10_u8_n2688 ), .ZN(_u10_u8_n2169 ) );
NAND2_X1 _u10_u8_U1178  ( .A1(_u10_u8_n3185 ), .A2(_u10_u8_n2169 ), .ZN(_u10_u8_n3286 ) );
NAND2_X1 _u10_u8_U1177  ( .A1(_u10_u8_n2833 ), .A2(_u10_u8_n3278 ), .ZN(_u10_u8_n3298 ) );
NAND3_X1 _u10_u8_U1176  ( .A1(_u10_u8_n3297 ), .A2(_u10_u8_n2838 ), .A3(_u10_u8_n3298 ), .ZN(_u10_u8_n3296 ) );
NAND2_X1 _u10_u8_U1175  ( .A1(_u10_u8_n2830 ), .A2(_u10_u8_n3296 ), .ZN(_u10_u8_n3287 ) );
NAND2_X1 _u10_u8_U1174  ( .A1(_u10_u8_n3295 ), .A2(_u10_u8_n3001 ), .ZN(_u10_u8_n3292 ) );
NAND2_X1 _u10_u8_U1173  ( .A1(_u10_u8_n3294 ), .A2(_u10_u8_n2089 ), .ZN(_u10_u8_n3293 ) );
AND2_X1 _u10_u8_U1172  ( .A1(_u10_u8_n3292 ), .A2(_u10_u8_n3293 ), .ZN(_u10_u8_n2548 ) );
NAND2_X1 _u10_u8_U1171  ( .A1(_u10_u8_n2548 ), .A2(_u10_u8_n2091 ), .ZN(_u10_u8_n2304 ) );
NAND2_X1 _u10_u8_U1170  ( .A1(_u10_u8_n2304 ), .A2(_u10_u8_n2446 ), .ZN(_u10_u8_n3290 ) );
NAND2_X1 _u10_u8_U1169  ( .A1(_u10_u8_n2549 ), .A2(_u10_u8_n2446 ), .ZN(_u10_u8_n2790 ) );
NOR2_X1 _u10_u8_U1168  ( .A1(_u10_u8_n1936 ), .A2(_u10_u8_n2790 ), .ZN(_u10_u8_n2789 ) );
INV_X1 _u10_u8_U1167  ( .A(_u10_u8_n2789 ), .ZN(_u10_u8_n3291 ) );
OR2_X1 _u10_u8_U1166  ( .A1(_u10_u8_n2828 ), .A2(_u10_u8_n2790 ), .ZN(_u10_u8_n2498 ) );
NAND4_X1 _u10_u8_U1165  ( .A1(_u10_u8_n3290 ), .A2(_u10_u8_n3291 ), .A3(_u10_u8_n2498 ), .A4(_u10_u8_n2001 ), .ZN(_u10_u8_n3289 ) );
NAND2_X1 _u10_u8_U1164  ( .A1(_u10_u8_n2445 ), .A2(_u10_u8_n3289 ), .ZN(_u10_u8_n3288 ) );
NAND3_X1 _u10_u8_U1163  ( .A1(_u10_u8_n3286 ), .A2(_u10_u8_n3287 ), .A3(_u10_u8_n3288 ), .ZN(_u10_u8_n3280 ) );
NOR2_X1 _u10_u8_U1162  ( .A1(_u10_u8_n2940 ), .A2(_u10_u8_n1913 ), .ZN(_u10_u8_n3281 ) );
INV_X1 _u10_u8_U1161  ( .A(1'b0), .ZN(_u10_u8_n1864 ) );
NAND2_X1 _u10_u8_U1160  ( .A1(1'b0), .A2(_u10_u8_n2588 ), .ZN(_u10_u8_n2141 ) );
INV_X1 _u10_u8_U1159  ( .A(_u10_u8_n2141 ), .ZN(_u10_u8_n3159 ) );
NAND3_X1 _u10_u8_U1158  ( .A1(_u10_u8_n2103 ), .A2(_u10_u8_n1864 ), .A3(_u10_u8_n3159 ), .ZN(_u10_u8_n2520 ) );
INV_X1 _u10_u8_U1157  ( .A(_u10_u8_n2520 ), .ZN(_u10_u8_n2630 ) );
INV_X1 _u10_u8_U1156  ( .A(_u10_u8_n2307 ), .ZN(_u10_u8_n2382 ) );
NOR4_X1 _u10_u8_U1155  ( .A1(_u10_u8_n2382 ), .A2(_u10_u8_n2722 ), .A3(_u10_u8_n1925 ), .A4(_u10_u8_n2508 ), .ZN(_u10_u8_n3260 ) );
NOR2_X1 _u10_u8_U1154  ( .A1(_u10_u8_n2498 ), .A2(_u10_u8_n2911 ), .ZN(_u10_u8_n2633 ) );
NOR2_X1 _u10_u8_U1153  ( .A1(_u10_u8_n2633 ), .A2(_u10_u8_n3278 ), .ZN(_u10_u8_n3285 ) );
INV_X1 _u10_u8_U1152  ( .A(_u10_u8_n1866 ), .ZN(_u10_u8_n1926 ) );
NOR2_X1 _u10_u8_U1151  ( .A1(_u10_u8_n3285 ), .A2(_u10_u8_n1926 ), .ZN(_u10_u8_n3284 ) );
NOR4_X1 _u10_u8_U1150  ( .A1(1'b0), .A2(_u10_u8_n2630 ), .A3(_u10_u8_n3260 ),.A4(_u10_u8_n3284 ), .ZN(_u10_u8_n3283 ) );
NOR2_X1 _u10_u8_U1149  ( .A1(_u10_u8_n3283 ), .A2(_u10_u8_n2980 ), .ZN(_u10_u8_n3282 ) );
NOR4_X1 _u10_u8_U1148  ( .A1(_u10_u8_n3279 ), .A2(_u10_u8_n3280 ), .A3(_u10_u8_n3281 ), .A4(_u10_u8_n3282 ), .ZN(_u10_u8_n3241 ) );
NAND2_X1 _u10_u8_U1147  ( .A1(_u10_u8_n1836 ), .A2(_u10_u8_n2291 ), .ZN(_u10_u8_n2147 ) );
NAND2_X1 _u10_u8_U1146  ( .A1(_u10_u8_n2443 ), .A2(_u10_u8_n2147 ), .ZN(_u10_u8_n3261 ) );
INV_X1 _u10_u8_U1145  ( .A(_u10_u8_n1841 ), .ZN(_u10_u8_n2571 ) );
NAND2_X1 _u10_u8_U1144  ( .A1(_u10_u8_n2571 ), .A2(_u10_u8_n3278 ), .ZN(_u10_u8_n3277 ) );
NAND2_X1 _u10_u8_U1143  ( .A1(_u10_u8_n3276 ), .A2(_u10_u8_n3277 ), .ZN(_u10_u8_n2819 ) );
OR2_X1 _u10_u8_U1142  ( .A1(_u10_u8_n2819 ), .A2(_u10_u8_n3275 ), .ZN(_u10_u8_n3273 ) );
NAND2_X1 _u10_u8_U1141  ( .A1(_u10_u8_n2815 ), .A2(_u10_u8_n2080 ), .ZN(_u10_u8_n3274 ) );
NAND2_X1 _u10_u8_U1140  ( .A1(_u10_u8_n2014 ), .A2(_u10_u8_n3274 ), .ZN(_u10_u8_n2165 ) );
NAND2_X1 _u10_u8_U1139  ( .A1(_u10_u8_n3273 ), .A2(_u10_u8_n2165 ), .ZN(_u10_u8_n3262 ) );
NAND2_X1 _u10_u8_U1138  ( .A1(_u10_u8_n2688 ), .A2(_u10_u8_n2126 ), .ZN(_u10_u8_n1956 ) );
INV_X1 _u10_u8_U1137  ( .A(_u10_u8_n1956 ), .ZN(_u10_u8_n1860 ) );
NOR2_X1 _u10_u8_U1136  ( .A1(1'b0), .A2(_u10_u8_n2498 ), .ZN(_u10_u8_n3271 ));
NOR2_X1 _u10_u8_U1135  ( .A1(_u10_u8_n3271 ), .A2(_u10_u8_n3272 ), .ZN(_u10_u8_n3270 ) );
NOR2_X1 _u10_u8_U1134  ( .A1(_u10_u8_n1860 ), .A2(_u10_u8_n3270 ), .ZN(_u10_u8_n3264 ) );
INV_X1 _u10_u8_U1133  ( .A(_u10_u8_n2632 ), .ZN(_u10_u8_n3202 ) );
NAND2_X1 _u10_u8_U1132  ( .A1(_u10_u8_n3236 ), .A2(_u10_u8_n3269 ), .ZN(_u10_u8_n3036 ) );
INV_X1 _u10_u8_U1131  ( .A(_u10_u8_n3036 ), .ZN(_u10_u8_n1960 ) );
NAND2_X1 _u10_u8_U1130  ( .A1(_u10_u8_n3202 ), .A2(_u10_u8_n1960 ), .ZN(_u10_u8_n3079 ) );
NOR3_X1 _u10_u8_U1129  ( .A1(_u10_u8_n3079 ), .A2(1'b0), .A3(_u10_u8_n3268 ),.ZN(_u10_u8_n3265 ) );
INV_X1 _u10_u8_U1128  ( .A(_u10_u8_n2014 ), .ZN(_u10_u8_n2709 ) );
NAND2_X1 _u10_u8_U1127  ( .A1(_u10_u8_n2709 ), .A2(_u10_u8_n2166 ), .ZN(_u10_u8_n2145 ) );
INV_X1 _u10_u8_U1126  ( .A(_u10_u8_n2145 ), .ZN(_u10_u8_n3258 ) );
NOR2_X1 _u10_u8_U1125  ( .A1(_u10_u8_n3258 ), .A2(_u10_u8_n2183 ), .ZN(_u10_u8_n3267 ) );
NOR2_X1 _u10_u8_U1124  ( .A1(_u10_u8_n3267 ), .A2(_u10_u8_n2567 ), .ZN(_u10_u8_n3266 ) );
NOR3_X1 _u10_u8_U1123  ( .A1(_u10_u8_n3264 ), .A2(_u10_u8_n3265 ), .A3(_u10_u8_n3266 ), .ZN(_u10_u8_n3263 ) );
NAND3_X1 _u10_u8_U1122  ( .A1(_u10_u8_n3261 ), .A2(_u10_u8_n3262 ), .A3(_u10_u8_n3263 ), .ZN(_u10_u8_n3243 ) );
INV_X1 _u10_u8_U1121  ( .A(_u10_u8_n2102 ), .ZN(_u10_u8_n2509 ) );
NAND2_X1 _u10_u8_U1120  ( .A1(_u10_u8_n3260 ), .A2(_u10_u8_n2509 ), .ZN(_u10_u8_n3247 ) );
INV_X1 _u10_u8_U1119  ( .A(_u10_u8_n3259 ), .ZN(_u10_u8_n2015 ) );
NAND2_X1 _u10_u8_U1118  ( .A1(_u10_u8_n2015 ), .A2(_u10_u8_n3258 ), .ZN(_u10_u8_n3248 ) );
NAND2_X1 _u10_u8_U1117  ( .A1(_u10_u8_n2251 ), .A2(_u10_u8_n2169 ), .ZN(_u10_u8_n3255 ) );
OR2_X1 _u10_u8_U1116  ( .A1(_u10_u8_n3157 ), .A2(_u10_u8_n2256 ), .ZN(_u10_u8_n3257 ) );
NAND2_X1 _u10_u8_U1115  ( .A1(_u10_u8_n2105 ), .A2(_u10_u8_n3257 ), .ZN(_u10_u8_n3256 ) );
AND2_X1 _u10_u8_U1114  ( .A1(_u10_u8_n3255 ), .A2(_u10_u8_n3256 ), .ZN(_u10_u8_n3212 ) );
INV_X1 _u10_u8_U1113  ( .A(_u10_u8_n2037 ), .ZN(_u10_u8_n2987 ) );
NAND2_X1 _u10_u8_U1112  ( .A1(_u10_u8_n2987 ), .A2(_u10_u8_n2038 ), .ZN(_u10_u8_n2212 ) );
NOR2_X1 _u10_u8_U1111  ( .A1(_u10_u8_n2212 ), .A2(1'b0), .ZN(_u10_u8_n2658 ));
INV_X1 _u10_u8_U1110  ( .A(_u10_u8_n2658 ), .ZN(_u10_u8_n2343 ) );
NAND2_X1 _u10_u8_U1109  ( .A1(_u10_u8_n2344 ), .A2(_u10_u8_n3254 ), .ZN(_u10_u8_n1928 ) );
NAND2_X1 _u10_u8_U1108  ( .A1(_u10_u8_n2588 ), .A2(_u10_u8_n1928 ), .ZN(_u10_u8_n3253 ) );
NAND2_X1 _u10_u8_U1107  ( .A1(_u10_u8_n2343 ), .A2(_u10_u8_n3253 ), .ZN(_u10_u8_n3252 ) );
NAND2_X1 _u10_u8_U1106  ( .A1(_u10_u8_n2105 ), .A2(_u10_u8_n3252 ), .ZN(_u10_u8_n3251 ) );
NAND2_X1 _u10_u8_U1105  ( .A1(_u10_u8_n3212 ), .A2(_u10_u8_n3251 ), .ZN(_u10_u8_n3250 ) );
NAND2_X1 _u10_u8_U1104  ( .A1(_u10_u8_n2307 ), .A2(_u10_u8_n3250 ), .ZN(_u10_u8_n3249 ) );
NAND3_X1 _u10_u8_U1103  ( .A1(_u10_u8_n3247 ), .A2(_u10_u8_n3248 ), .A3(_u10_u8_n3249 ), .ZN(_u10_u8_n3244 ) );
AND2_X1 _u10_u8_U1102  ( .A1(_u10_u8_n2915 ), .A2(_u10_u8_n2059 ), .ZN(_u10_u8_n2957 ) );
AND3_X1 _u10_u8_U1101  ( .A1(_u10_u8_n3223 ), .A2(_u10_u8_n2837 ), .A3(_u10_u8_n2957 ), .ZN(_u10_u8_n2051 ) );
NOR2_X1 _u10_u8_U1100  ( .A1(_u10_u8_n2528 ), .A2(_u10_u8_n2051 ), .ZN(_u10_u8_n2605 ) );
NOR2_X1 _u10_u8_U1099  ( .A1(_u10_u8_n2605 ), .A2(_u10_u8_n2346 ), .ZN(_u10_u8_n3245 ) );
NOR2_X1 _u10_u8_U1098  ( .A1(_u10_u8_n2291 ), .A2(_u10_u8_n2062 ), .ZN(_u10_u8_n3246 ) );
NOR4_X1 _u10_u8_U1097  ( .A1(_u10_u8_n3243 ), .A2(_u10_u8_n3244 ), .A3(_u10_u8_n3245 ), .A4(_u10_u8_n3246 ), .ZN(_u10_u8_n3242 ) );
NAND2_X1 _u10_u8_U1096  ( .A1(_u10_u8_n3241 ), .A2(_u10_u8_n3242 ), .ZN(_u10_u8_n2311 ) );
OR3_X1 _u10_u8_U1095  ( .A1(_u10_u8_n1987 ), .A2(_u10_u8_n3240 ), .A3(_u10_u8_n2311 ), .ZN(_u10_u8_n3192 ) );
INV_X1 _u10_u8_U1094  ( .A(_u10_u8_n2886 ), .ZN(_u10_u8_n2720 ) );
NOR2_X1 _u10_u8_U1093  ( .A1(_u10_u8_n2004 ), .A2(_u10_u8_n2720 ), .ZN(_u10_u8_n2455 ) );
INV_X1 _u10_u8_U1092  ( .A(_u10_u8_n2488 ), .ZN(_u10_u8_n2938 ) );
AND3_X1 _u10_u8_U1091  ( .A1(_u10_u8_n2455 ), .A2(_u10_u8_n1859 ), .A3(_u10_u8_n2938 ), .ZN(_u10_u8_n3239 ) );
INV_X1 _u10_u8_U1090  ( .A(_u10_u8_n2633 ), .ZN(_u10_u8_n2937 ) );
NOR2_X1 _u10_u8_U1089  ( .A1(_u10_u8_n3239 ), .A2(_u10_u8_n2937 ), .ZN(_u10_u8_n3227 ) );
NOR2_X1 _u10_u8_U1088  ( .A1(_u10_u8_n1976 ), .A2(_u10_u8_n1969 ), .ZN(_u10_u8_n3237 ) );
NOR2_X1 _u10_u8_U1087  ( .A1(1'b0), .A2(_u10_u8_n2947 ), .ZN(_u10_u8_n3238 ));
NOR3_X1 _u10_u8_U1086  ( .A1(_u10_u8_n2476 ), .A2(_u10_u8_n3237 ), .A3(_u10_u8_n3238 ), .ZN(_u10_u8_n3235 ) );
NOR3_X1 _u10_u8_U1085  ( .A1(_u10_u8_n1813 ), .A2(_u10_u8_n1817 ), .A3(_u10_SYNOPSYS_UNCONNECTED_35 ), .ZN(_u10_u8_n3135 ) );
NAND2_X1 _u10_u8_U1084  ( .A1(_u10_u8_n3135 ), .A2(_u10_u8_n3236 ), .ZN(_u10_u8_n2573 ) );
NOR2_X1 _u10_u8_U1083  ( .A1(_u10_u8_n3235 ), .A2(_u10_u8_n2573 ), .ZN(_u10_u8_n3228 ) );
NOR2_X1 _u10_u8_U1082  ( .A1(_u10_u8_n2216 ), .A2(_u10_u8_n1868 ), .ZN(_u10_u8_n3233 ) );
INV_X1 _u10_u8_U1081  ( .A(_u10_u8_n2550 ), .ZN(_u10_u8_n2475 ) );
NOR3_X1 _u10_u8_U1080  ( .A1(_u10_u8_n2475 ), .A2(1'b0), .A3(_u10_u8_n1925 ),.ZN(_u10_u8_n3234 ) );
NOR3_X1 _u10_u8_U1079  ( .A1(_u10_u8_n3233 ), .A2(1'b0), .A3(_u10_u8_n3234 ),.ZN(_u10_u8_n3232 ) );
NOR2_X1 _u10_u8_U1078  ( .A1(_u10_u8_n3232 ), .A2(_u10_u8_n2037 ), .ZN(_u10_u8_n3229 ) );
NOR2_X1 _u10_u8_U1077  ( .A1(_u10_u8_n3231 ), .A2(_u10_u8_n2365 ), .ZN(_u10_u8_n3230 ) );
NOR4_X1 _u10_u8_U1076  ( .A1(_u10_u8_n3227 ), .A2(_u10_u8_n3228 ), .A3(_u10_u8_n3229 ), .A4(_u10_u8_n3230 ), .ZN(_u10_u8_n3205 ) );
NOR3_X1 _u10_u8_U1075  ( .A1(_u10_u8_n3226 ), .A2(_u10_u8_n2687 ), .A3(_u10_u8_n2145 ), .ZN(_u10_u8_n3217 ) );
NOR3_X1 _u10_u8_U1074  ( .A1(_u10_u8_n3225 ), .A2(1'b0), .A3(_u10_u8_n2587 ),.ZN(_u10_u8_n3218 ) );
NOR2_X1 _u10_u8_U1073  ( .A1(_u10_u8_n3159 ), .A2(1'b0), .ZN(_u10_u8_n3224 ));
NOR2_X1 _u10_u8_U1072  ( .A1(_u10_u8_n3224 ), .A2(_u10_u8_n2584 ), .ZN(_u10_u8_n3219 ) );
NAND2_X1 _u10_u8_U1071  ( .A1(_u10_u8_n3222 ), .A2(_u10_u8_n3223 ), .ZN(_u10_u8_n2048 ) );
INV_X1 _u10_u8_U1070  ( .A(_u10_u8_n2048 ), .ZN(_u10_u8_n2859 ) );
NOR2_X1 _u10_u8_U1069  ( .A1(_u10_u8_n2859 ), .A2(_u10_u8_n2054 ), .ZN(_u10_u8_n3221 ) );
NOR2_X1 _u10_u8_U1068  ( .A1(_u10_u8_n3221 ), .A2(_u10_u8_n2346 ), .ZN(_u10_u8_n3220 ) );
NOR4_X1 _u10_u8_U1067  ( .A1(_u10_u8_n3217 ), .A2(_u10_u8_n3218 ), .A3(_u10_u8_n3219 ), .A4(_u10_u8_n3220 ), .ZN(_u10_u8_n3206 ) );
NAND2_X1 _u10_u8_U1066  ( .A1(_u10_u8_n2377 ), .A2(_u10_u8_n2721 ), .ZN(_u10_u8_n3213 ) );
AND4_X1 _u10_u8_U1065  ( .A1(1'b0), .A2(_u10_u8_n2502 ), .A3(_u10_u8_n2972 ),.A4(_u10_u8_n3040 ), .ZN(_u10_u8_n2406 ) );
NAND2_X1 _u10_u8_U1064  ( .A1(_u10_u8_n2406 ), .A2(_u10_u8_n2979 ), .ZN(_u10_u8_n3214 ) );
NAND2_X1 _u10_u8_U1063  ( .A1(_u10_u8_n2630 ), .A2(_u10_u8_n3216 ), .ZN(_u10_u8_n2376 ) );
INV_X1 _u10_u8_U1062  ( .A(_u10_u8_n2376 ), .ZN(_u10_u8_n3108 ) );
NAND2_X1 _u10_u8_U1061  ( .A1(_u10_u8_n3108 ), .A2(_u10_u8_n2507 ), .ZN(_u10_u8_n3215 ) );
NOR2_X1 _u10_u8_U1060  ( .A1(_u10_u8_n2937 ), .A2(1'b0), .ZN(_u10_u8_n2649 ));
INV_X1 _u10_u8_U1059  ( .A(_u10_u8_n2253 ), .ZN(_u10_u8_n2971 ) );
NAND2_X1 _u10_u8_U1058  ( .A1(_u10_u8_n2649 ), .A2(_u10_u8_n2971 ), .ZN(_u10_u8_n2918 ) );
NAND4_X1 _u10_u8_U1057  ( .A1(_u10_u8_n3213 ), .A2(_u10_u8_n3214 ), .A3(_u10_u8_n3215 ), .A4(_u10_u8_n2918 ), .ZN(_u10_u8_n3208 ) );
NOR2_X1 _u10_u8_U1056  ( .A1(_u10_u8_n2000 ), .A2(_u10_u8_n2902 ), .ZN(_u10_u8_n3209 ) );
NOR2_X1 _u10_u8_U1055  ( .A1(_u10_u8_n3212 ), .A2(_u10_u8_n2475 ), .ZN(_u10_u8_n3210 ) );
INV_X1 _u10_u8_U1054  ( .A(_u10_u8_n2441 ), .ZN(_u10_u8_n3128 ) );
NOR2_X1 _u10_u8_U1053  ( .A1(_u10_u8_n2356 ), .A2(_u10_u8_n3128 ), .ZN(_u10_u8_n3211 ) );
NOR4_X1 _u10_u8_U1052  ( .A1(_u10_u8_n3208 ), .A2(_u10_u8_n3209 ), .A3(_u10_u8_n3210 ), .A4(_u10_u8_n3211 ), .ZN(_u10_u8_n3207 ) );
NAND3_X1 _u10_u8_U1051  ( .A1(_u10_u8_n3205 ), .A2(_u10_u8_n3206 ), .A3(_u10_u8_n3207 ), .ZN(_u10_u8_n2611 ) );
NOR2_X1 _u10_u8_U1050  ( .A1(_u10_u8_n2212 ), .A2(_u10_u8_n2216 ), .ZN(_u10_u8_n1937 ) );
NOR2_X1 _u10_u8_U1049  ( .A1(_u10_u8_n2533 ), .A2(_u10_u8_n2214 ), .ZN(_u10_u8_n2765 ) );
INV_X1 _u10_u8_U1048  ( .A(_u10_u8_n2005 ), .ZN(_u10_u8_n2111 ) );
AND2_X1 _u10_u8_U1047  ( .A1(_u10_u8_n2765 ), .A2(_u10_u8_n2111 ), .ZN(_u10_u8_n3201 ) );
INV_X1 _u10_u8_U1046  ( .A(_u10_u8_n3059 ), .ZN(_u10_u8_n3076 ) );
NAND2_X1 _u10_u8_U1045  ( .A1(_u10_u8_n3201 ), .A2(_u10_u8_n3076 ), .ZN(_u10_u8_n3204 ) );
NAND2_X1 _u10_u8_U1044  ( .A1(_u10_u8_n1937 ), .A2(_u10_u8_n3204 ), .ZN(_u10_u8_n3193 ) );
NAND2_X1 _u10_u8_U1043  ( .A1(_u10_u8_n2254 ), .A2(_u10_u8_n2212 ), .ZN(_u10_u8_n3203 ) );
NAND3_X1 _u10_u8_U1042  ( .A1(_u10_u8_n3203 ), .A2(_u10_u8_n2175 ), .A3(_u10_u8_n2649 ), .ZN(_u10_u8_n3194 ) );
NOR2_X1 _u10_u8_U1041  ( .A1(_u10_u8_n2985 ), .A2(1'b0), .ZN(_u10_u8_n1959 ));
NAND2_X1 _u10_u8_U1040  ( .A1(_u10_u8_n1959 ), .A2(_u10_u8_n3202 ), .ZN(_u10_u8_n2202 ) );
NAND4_X1 _u10_u8_U1039  ( .A1(_u10_u8_n3079 ), .A2(_u10_u8_n2621 ), .A3(_u10_u8_n2202 ), .A4(_u10_u8_n2798 ), .ZN(_u10_u8_n3200 ) );
NAND2_X1 _u10_u8_U1038  ( .A1(_u10_u8_n3201 ), .A2(_u10_u8_n2937 ), .ZN(_u10_u8_n2772 ) );
NAND2_X1 _u10_u8_U1037  ( .A1(_u10_u8_n3200 ), .A2(_u10_u8_n2772 ), .ZN(_u10_u8_n3195 ) );
NAND2_X1 _u10_u8_U1036  ( .A1(_u10_u8_n2765 ), .A2(_u10_u8_n1869 ), .ZN(_u10_u8_n3199 ) );
NAND2_X1 _u10_u8_U1035  ( .A1(_u10_u8_n2049 ), .A2(_u10_u8_n3199 ), .ZN(_u10_u8_n3057 ) );
NOR2_X1 _u10_u8_U1034  ( .A1(_u10_u8_n2495 ), .A2(_u10_u8_n3057 ), .ZN(_u10_u8_n3197 ) );
NOR2_X1 _u10_u8_U1033  ( .A1(_u10_u8_n2883 ), .A2(_u10_u8_n2485 ), .ZN(_u10_u8_n3198 ) );
NOR2_X1 _u10_u8_U1032  ( .A1(_u10_u8_n3197 ), .A2(_u10_u8_n3198 ), .ZN(_u10_u8_n3196 ) );
NAND4_X1 _u10_u8_U1031  ( .A1(_u10_u8_n3193 ), .A2(_u10_u8_n3194 ), .A3(_u10_u8_n3195 ), .A4(_u10_u8_n3196 ), .ZN(_u10_u8_n2887 ) );
NOR4_X1 _u10_u8_U1030  ( .A1(_u10_u8_n3191 ), .A2(_u10_u8_n3192 ), .A3(_u10_u8_n2611 ), .A4(_u10_u8_n2887 ), .ZN(_u10_u8_n3015 ) );
NAND3_X1 _u10_u8_U1029  ( .A1(_u10_u8_n3190 ), .A2(_u10_u8_n2049 ), .A3(_u10_u8_n2957 ), .ZN(_u10_u8_n2699 ) );
OR2_X1 _u10_u8_U1028  ( .A1(_u10_u8_n2699 ), .A2(_u10_u8_n1813 ), .ZN(_u10_u8_n3187 ) );
NAND3_X1 _u10_u8_U1027  ( .A1(_u10_u8_n2978 ), .A2(_u10_u8_n2405 ), .A3(1'b0), .ZN(_u10_u8_n3188 ) );
NAND4_X1 _u10_u8_U1026  ( .A1(_u10_u8_n3058 ), .A2(_u10_u8_n3187 ), .A3(_u10_u8_n3188 ), .A4(_u10_u8_n3189 ), .ZN(_u10_u8_n3186 ) );
NAND2_X1 _u10_u8_U1025  ( .A1(_u10_u8_n2063 ), .A2(_u10_u8_n3186 ), .ZN(_u10_u8_n3163 ) );
NAND2_X1 _u10_u8_U1024  ( .A1(_u10_u8_n3185 ), .A2(_u10_u8_n2329 ), .ZN(_u10_u8_n3164 ) );
NAND2_X1 _u10_u8_U1023  ( .A1(_u10_u8_n2689 ), .A2(_u10_u8_n2365 ), .ZN(_u10_u8_n2736 ) );
NOR2_X1 _u10_u8_U1022  ( .A1(_u10_u8_n2736 ), .A2(_u10_u8_n2488 ), .ZN(_u10_u8_n1855 ) );
INV_X1 _u10_u8_U1021  ( .A(_u10_u8_n1855 ), .ZN(_u10_u8_n3184 ) );
NOR2_X1 _u10_u8_U1020  ( .A1(_u10_u8_n2274 ), .A2(_u10_u8_n2359 ), .ZN(_u10_u8_n2952 ) );
NOR2_X1 _u10_u8_U1019  ( .A1(_u10_u8_n3184 ), .A2(_u10_u8_n2952 ), .ZN(_u10_u8_n2776 ) );
OR2_X1 _u10_u8_U1018  ( .A1(_u10_u8_n2852 ), .A2(_u10_u8_n2776 ), .ZN(_u10_u8_n3165 ) );
NAND2_X1 _u10_u8_U1017  ( .A1(_u10_u8_n3126 ), .A2(_u10_u8_n2915 ), .ZN(_u10_u8_n3065 ) );
NOR3_X1 _u10_u8_U1016  ( .A1(_u10_u8_n3065 ), .A2(1'b0), .A3(_u10_u8_n2632 ),.ZN(_u10_u8_n3182 ) );
NOR3_X1 _u10_u8_U1015  ( .A1(_u10_u8_n3182 ), .A2(_u10_u8_n3183 ), .A3(_u10_u8_n3108 ), .ZN(_u10_u8_n3181 ) );
NOR2_X1 _u10_u8_U1014  ( .A1(_u10_u8_n3181 ), .A2(_u10_u8_n3162 ), .ZN(_u10_u8_n3167 ) );
INV_X1 _u10_u8_U1013  ( .A(_u10_u8_n3180 ), .ZN(_u10_u8_n3140 ) );
NAND3_X1 _u10_u8_U1012  ( .A1(_u10_u8_n3140 ), .A2(_u10_u8_n2163 ), .A3(_u10_u8_n2092 ), .ZN(_u10_u8_n3175 ) );
NOR4_X1 _u10_u8_U1011  ( .A1(_u10_u8_n2411 ), .A2(_u10_u8_n2710 ), .A3(_u10_u8_n3141 ), .A4(_u10_u8_n3089 ), .ZN(_u10_u8_n3179 ) );
NOR2_X1 _u10_u8_U1010  ( .A1(1'b0), .A2(_u10_u8_n3179 ), .ZN(_u10_u8_n3177 ));
NOR2_X1 _u10_u8_U1009  ( .A1(_u10_u8_n1898 ), .A2(_u10_u8_n1847 ), .ZN(_u10_u8_n3178 ) );
NOR4_X1 _u10_u8_U1008  ( .A1(_u10_u8_n3175 ), .A2(_u10_u8_n3176 ), .A3(_u10_u8_n3177 ), .A4(_u10_u8_n3178 ), .ZN(_u10_u8_n3173 ) );
NAND2_X1 _u10_u8_U1007  ( .A1(_u10_u8_n3135 ), .A2(_u10_u8_n3174 ), .ZN(_u10_u8_n2159 ) );
NOR2_X1 _u10_u8_U1006  ( .A1(_u10_u8_n3173 ), .A2(_u10_u8_n2159 ), .ZN(_u10_u8_n3168 ) );
OR3_X1 _u10_u8_U1005  ( .A1(_u10_u8_n3172 ), .A2(1'b0), .A3(_u10_u8_n3126 ),.ZN(_u10_u8_n3171 ) );
NAND2_X1 _u10_u8_U1004  ( .A1(_u10_u8_n2600 ), .A2(_u10_u8_n3171 ), .ZN(_u10_u8_n3153 ) );
AND3_X1 _u10_u8_U1003  ( .A1(_u10_u8_n3153 ), .A2(_u10_u8_n2947 ), .A3(_u10_u8_n2579 ), .ZN(_u10_u8_n3170 ) );
NOR2_X1 _u10_u8_U1002  ( .A1(_u10_u8_n3170 ), .A2(_u10_u8_n2359 ), .ZN(_u10_u8_n3169 ) );
NOR3_X1 _u10_u8_U1001  ( .A1(_u10_u8_n3167 ), .A2(_u10_u8_n3168 ), .A3(_u10_u8_n3169 ), .ZN(_u10_u8_n3166 ) );
NAND4_X1 _u10_u8_U1000  ( .A1(_u10_u8_n3163 ), .A2(_u10_u8_n3164 ), .A3(_u10_u8_n3165 ), .A4(_u10_u8_n3166 ), .ZN(_u10_u8_n3130 ) );
NAND2_X1 _u10_u8_U999  ( .A1(_u10_u8_n2375 ), .A2(_u10_u8_n3162 ), .ZN(_u10_u8_n1923 ) );
NAND2_X1 _u10_u8_U998  ( .A1(_u10_u8_n3062 ), .A2(_u10_u8_n1923 ), .ZN(_u10_u8_n3154 ) );
NAND2_X1 _u10_u8_U997  ( .A1(_u10_u8_n2103 ), .A2(_u10_u8_n2509 ), .ZN(_u10_u8_n3161 ) );
NAND2_X1 _u10_u8_U996  ( .A1(_u10_u8_n2344 ), .A2(_u10_u8_n3161 ), .ZN(_u10_u8_n3160 ) );
NAND2_X1 _u10_u8_U995  ( .A1(_u10_u8_n3159 ), .A2(_u10_u8_n3160 ), .ZN(_u10_u8_n2635 ) );
AND3_X1 _u10_u8_U994  ( .A1(_u10_u8_n2549 ), .A2(_u10_u8_n2108 ), .A3(_u10_u8_n3126 ), .ZN(_u10_u8_n3093 ) );
NAND2_X1 _u10_u8_U993  ( .A1(_u10_u8_n3093 ), .A2(_u10_u8_n2941 ), .ZN(_u10_u8_n3158 ) );
NAND3_X1 _u10_u8_U992  ( .A1(_u10_u8_n3076 ), .A2(_u10_u8_n3066 ), .A3(_u10_u8_n3158 ), .ZN(_u10_u8_n3156 ) );
NAND2_X1 _u10_u8_U991  ( .A1(_u10_u8_n3156 ), .A2(_u10_u8_n3157 ), .ZN(_u10_u8_n3155 ) );
NAND3_X1 _u10_u8_U990  ( .A1(_u10_u8_n3154 ), .A2(_u10_u8_n2635 ), .A3(_u10_u8_n3155 ), .ZN(_u10_u8_n3131 ) );
INV_X1 _u10_u8_U989  ( .A(_u10_u8_n2594 ), .ZN(_u10_u8_n2846 ) );
NAND3_X1 _u10_u8_U988  ( .A1(_u10_u8_n2162 ), .A2(_u10_u8_n2082 ), .A3(_u10_u8_n2105 ), .ZN(_u10_u8_n2077 ) );
NAND4_X1 _u10_u8_U987  ( .A1(_u10_u8_n3153 ), .A2(_u10_u8_n1969 ), .A3(_u10_u8_n2846 ), .A4(_u10_u8_n2077 ), .ZN(_u10_u8_n3148 ) );
NAND2_X1 _u10_u8_U986  ( .A1(_u10_u8_n2838 ), .A2(_u10_u8_n3128 ), .ZN(_u10_u8_n3152 ) );
NAND2_X1 _u10_u8_U985  ( .A1(_u10_u8_n3152 ), .A2(_u10_u8_n2600 ), .ZN(_u10_u8_n3151 ) );
NAND2_X1 _u10_u8_U984  ( .A1(_u10_u8_n2282 ), .A2(_u10_u8_n3151 ), .ZN(_u10_u8_n2601 ) );
NOR4_X1 _u10_u8_U983  ( .A1(_u10_u8_n2885 ), .A2(_u10_u8_n2534 ), .A3(_u10_u8_n2214 ), .A4(_u10_u8_n3059 ), .ZN(_u10_u8_n3150 ) );
NOR2_X1 _u10_u8_U982  ( .A1(_u10_u8_n3150 ), .A2(_u10_u8_n2853 ), .ZN(_u10_u8_n3149 ) );
NOR4_X1 _u10_u8_U981  ( .A1(_u10_u8_n3148 ), .A2(_u10_u8_n2601 ), .A3(_u10_u8_n3149 ), .A4(_u10_u8_n1975 ), .ZN(_u10_u8_n3146 ) );
NAND3_X1 _u10_u8_U980  ( .A1(_u10_SYNOPSYS_UNCONNECTED_38 ), .A2(_u10_SYNOPSYS_UNCONNECTED_34 ), .A3(_u10_u8_n3147 ), .ZN(_u10_u8_n2071 ) );
NOR2_X1 _u10_u8_U979  ( .A1(_u10_u8_n3146 ), .A2(_u10_u8_n2071 ), .ZN(_u10_u8_n3132 ) );
NOR2_X1 _u10_u8_U978  ( .A1(1'b0), .A2(_u10_u8_n1847 ), .ZN(_u10_u8_n3143 ));
INV_X1 _u10_u8_U977  ( .A(_u10_u8_n3145 ), .ZN(_u10_u8_n3144 ) );
NOR2_X1 _u10_u8_U976  ( .A1(_u10_u8_n3143 ), .A2(_u10_u8_n3144 ), .ZN(_u10_u8_n3142 ) );
NOR2_X1 _u10_u8_U975  ( .A1(1'b0), .A2(_u10_u8_n3142 ), .ZN(_u10_u8_n3137 ));
NAND2_X1 _u10_u8_U974  ( .A1(_u10_u8_n2549 ), .A2(_u10_u8_n3141 ), .ZN(_u10_u8_n3138 ) );
NAND2_X1 _u10_u8_U973  ( .A1(_u10_u8_n1896 ), .A2(_u10_u8_n3140 ), .ZN(_u10_u8_n2544 ) );
NAND2_X1 _u10_u8_U972  ( .A1(_u10_u8_n2089 ), .A2(_u10_u8_n2544 ), .ZN(_u10_u8_n3139 ) );
NAND2_X1 _u10_u8_U971  ( .A1(_u10_u8_n3138 ), .A2(_u10_u8_n3139 ), .ZN(_u10_u8_n2795 ) );
NOR4_X1 _u10_u8_U970  ( .A1(_u10_u8_n2300 ), .A2(_u10_u8_n3137 ), .A3(_u10_u8_n2304 ), .A4(_u10_u8_n2795 ), .ZN(_u10_u8_n3134 ) );
NAND2_X1 _u10_u8_U969  ( .A1(_u10_u8_n3135 ), .A2(_u10_u8_n3136 ), .ZN(_u10_u8_n2085 ) );
NOR2_X1 _u10_u8_U968  ( .A1(_u10_u8_n3134 ), .A2(_u10_u8_n2085 ), .ZN(_u10_u8_n3133 ) );
NOR4_X1 _u10_u8_U967  ( .A1(_u10_u8_n3130 ), .A2(_u10_u8_n3131 ), .A3(_u10_u8_n3132 ), .A4(_u10_u8_n3133 ), .ZN(_u10_u8_n3016 ) );
INV_X1 _u10_u8_U966  ( .A(_u10_u8_n2686 ), .ZN(_u10_u8_n2278 ) );
NAND4_X1 _u10_u8_U965  ( .A1(_u10_u8_n2105 ), .A2(_u10_u8_n2278 ), .A3(_u10_u8_n3129 ), .A4(_u10_u8_n2600 ), .ZN(_u10_u8_n2437 ) );
NAND2_X1 _u10_u8_U964  ( .A1(_u10_u8_n3128 ), .A2(_u10_u8_n2437 ), .ZN(_u10_u8_n3127 ) );
NAND2_X1 _u10_u8_U963  ( .A1(_u10_u8_n2815 ), .A2(_u10_u8_n3127 ), .ZN(_u10_u8_n3098 ) );
INV_X1 _u10_u8_U962  ( .A(_u10_u8_n2573 ), .ZN(_u10_u8_n1967 ) );
NAND2_X1 _u10_u8_U961  ( .A1(_u10_u8_n3126 ), .A2(_u10_u8_n2078 ), .ZN(_u10_u8_n3123 ) );
NAND2_X1 _u10_u8_U960  ( .A1(_u10_u8_n3076 ), .A2(_u10_u8_n1925 ), .ZN(_u10_u8_n3125 ) );
NAND2_X1 _u10_u8_U959  ( .A1(_u10_u8_n2669 ), .A2(_u10_u8_n3125 ), .ZN(_u10_u8_n3124 ) );
NAND4_X1 _u10_u8_U958  ( .A1(_u10_u8_n3122 ), .A2(_u10_u8_n3123 ), .A3(_u10_u8_n3124 ), .A4(_u10_u8_n2579 ), .ZN(_u10_u8_n3121 ) );
NAND2_X1 _u10_u8_U957  ( .A1(_u10_u8_n3121 ), .A2(_u10_u8_n2874 ), .ZN(_u10_u8_n3120 ) );
NAND2_X1 _u10_u8_U956  ( .A1(_u10_u8_n2382 ), .A2(_u10_u8_n3120 ), .ZN(_u10_u8_n3119 ) );
NAND2_X1 _u10_u8_U955  ( .A1(_u10_u8_n1967 ), .A2(_u10_u8_n3119 ), .ZN(_u10_u8_n3099 ) );
NAND2_X1 _u10_u8_U954  ( .A1(_u10_u8_n3118 ), .A2(_u10_u8_n3001 ), .ZN(_u10_u8_n3117 ) );
NAND2_X1 _u10_u8_U953  ( .A1(_u10_u8_n2446 ), .A2(_u10_u8_n3117 ), .ZN(_u10_u8_n3116 ) );
NAND2_X1 _u10_u8_U952  ( .A1(_u10_u8_n2445 ), .A2(_u10_u8_n3116 ), .ZN(_u10_u8_n3100 ) );
OR2_X1 _u10_u8_U951  ( .A1(_u10_u8_n3115 ), .A2(_u10_u8_n2687 ), .ZN(_u10_u8_n3114 ) );
AND3_X1 _u10_u8_U950  ( .A1(_u10_u8_n2061 ), .A2(_u10_u8_n2166 ), .A3(_u10_u8_n3114 ), .ZN(_u10_u8_n3045 ) );
NOR2_X1 _u10_u8_U949  ( .A1(1'b0), .A2(_u10_u8_n3045 ), .ZN(_u10_u8_n3113 ));
NOR2_X1 _u10_u8_U948  ( .A1(_u10_u8_n3113 ), .A2(1'b0), .ZN(_u10_u8_n3112 ));
NOR2_X1 _u10_u8_U947  ( .A1(_u10_u8_n3112 ), .A2(_u10_u8_n2356 ), .ZN(_u10_u8_n3102 ) );
NAND2_X1 _u10_u8_U946  ( .A1(_u10_u8_n2571 ), .A2(_u10_u8_n2165 ), .ZN(_u10_u8_n3078 ) );
NAND2_X1 _u10_u8_U945  ( .A1(_u10_u8_n2365 ), .A2(_u10_u8_n3078 ), .ZN(_u10_u8_n2241 ) );
NOR2_X1 _u10_u8_U944  ( .A1(_u10_u8_n2377 ), .A2(_u10_u8_n2241 ), .ZN(_u10_u8_n3111 ) );
NOR2_X1 _u10_u8_U943  ( .A1(_u10_u8_n3111 ), .A2(_u10_u8_n1869 ), .ZN(_u10_u8_n3103 ) );
NOR2_X1 _u10_u8_U942  ( .A1(_u10_u8_n2999 ), .A2(_u10_u8_n2977 ), .ZN(_u10_u8_n3061 ) );
NOR2_X1 _u10_u8_U941  ( .A1(_u10_u8_n3061 ), .A2(_u10_u8_n2367 ), .ZN(_u10_u8_n3106 ) );
NAND2_X1 _u10_u8_U940  ( .A1(_u10_u8_n2977 ), .A2(_u10_u8_n3000 ), .ZN(_u10_u8_n3110 ) );
NAND2_X1 _u10_u8_U939  ( .A1(_u10_u8_n3109 ), .A2(_u10_u8_n3110 ), .ZN(_u10_u8_n1924 ) );
AND2_X1 _u10_u8_U938  ( .A1(_u10_u8_n1924 ), .A2(_u10_u8_n3108 ), .ZN(_u10_u8_n3107 ) );
NOR2_X1 _u10_u8_U937  ( .A1(_u10_u8_n3106 ), .A2(_u10_u8_n3107 ), .ZN(_u10_u8_n3105 ) );
NOR2_X1 _u10_u8_U936  ( .A1(_u10_u8_n3105 ), .A2(_u10_u8_n2008 ), .ZN(_u10_u8_n3104 ) );
NOR3_X1 _u10_u8_U935  ( .A1(_u10_u8_n3102 ), .A2(_u10_u8_n3103 ), .A3(_u10_u8_n3104 ), .ZN(_u10_u8_n3101 ) );
NAND4_X1 _u10_u8_U934  ( .A1(_u10_u8_n3098 ), .A2(_u10_u8_n3099 ), .A3(_u10_u8_n3100 ), .A4(_u10_u8_n3101 ), .ZN(_u10_u8_n3071 ) );
NOR2_X1 _u10_u8_U933  ( .A1(_u10_u8_n1926 ), .A2(_u10_u8_n2980 ), .ZN(_u10_u8_n2218 ) );
INV_X1 _u10_u8_U932  ( .A(_u10_u8_n2721 ), .ZN(_u10_u8_n2910 ) );
NAND2_X1 _u10_u8_U931  ( .A1(_u10_u8_n2910 ), .A2(_u10_u8_n1869 ), .ZN(_u10_u8_n2779 ) );
NAND2_X1 _u10_u8_U930  ( .A1(_u10_u8_n2218 ), .A2(_u10_u8_n2779 ), .ZN(_u10_u8_n3081 ) );
NAND2_X1 _u10_u8_U929  ( .A1(_u10_u8_n1922 ), .A2(_u10_u8_n1864 ), .ZN(_u10_u8_n2179 ) );
NOR3_X1 _u10_u8_U928  ( .A1(_u10_u8_n1961 ), .A2(_u10_u8_n1918 ), .A3(_u10_u8_n2179 ), .ZN(_u10_u8_n2693 ) );
NAND2_X1 _u10_u8_U927  ( .A1(_u10_u8_n3097 ), .A2(_u10_u8_n1924 ), .ZN(_u10_u8_n3096 ) );
NAND2_X1 _u10_u8_U926  ( .A1(_u10_u8_n1984 ), .A2(_u10_u8_n3096 ), .ZN(_u10_u8_n2506 ) );
INV_X1 _u10_u8_U925  ( .A(_u10_u8_n2506 ), .ZN(_u10_u8_n2366 ) );
NAND2_X1 _u10_u8_U924  ( .A1(_u10_u8_n2366 ), .A2(_u10_u8_n2375 ), .ZN(_u10_u8_n2236 ) );
NAND2_X1 _u10_u8_U923  ( .A1(_u10_u8_n2693 ), .A2(_u10_u8_n2236 ), .ZN(_u10_u8_n3082 ) );
NAND2_X1 _u10_u8_U922  ( .A1(1'b0), .A2(_u10_u8_n2126 ), .ZN(_u10_u8_n3095 ));
NAND2_X1 _u10_u8_U921  ( .A1(_u10_u8_n1956 ), .A2(_u10_u8_n3095 ), .ZN(_u10_u8_n2907 ) );
OR2_X1 _u10_u8_U920  ( .A1(_u10_u8_n2902 ), .A2(_u10_u8_n2907 ), .ZN(_u10_u8_n3085 ) );
NAND2_X1 _u10_u8_U919  ( .A1(_u10_u8_n2256 ), .A2(_u10_u8_n2113 ), .ZN(_u10_u8_n3094 ) );
NAND2_X1 _u10_u8_U918  ( .A1(_u10_u8_n2688 ), .A2(_u10_u8_n3094 ), .ZN(_u10_u8_n3092 ) );
NAND2_X1 _u10_u8_U917  ( .A1(_u10_u8_n3093 ), .A2(_u10_u8_n3092 ), .ZN(_u10_u8_n3086 ) );
INV_X1 _u10_u8_U916  ( .A(_u10_u8_n2159 ), .ZN(_u10_u8_n1894 ) );
NAND2_X1 _u10_u8_U915  ( .A1(_u10_u8_n3067 ), .A2(_u10_u8_n1894 ), .ZN(_u10_u8_n3091 ) );
INV_X1 _u10_u8_U914  ( .A(_u10_u8_n3092 ), .ZN(_u10_u8_n2234 ) );
NAND3_X1 _u10_u8_U913  ( .A1(_u10_u8_n3091 ), .A2(_u10_u8_n2126 ), .A3(_u10_u8_n2234 ), .ZN(_u10_u8_n3090 ) );
NAND2_X1 _u10_u8_U912  ( .A1(1'b0), .A2(_u10_u8_n3090 ), .ZN(_u10_u8_n3087 ));
NAND3_X1 _u10_u8_U911  ( .A1(_u10_u8_n2329 ), .A2(_u10_u8_n3089 ), .A3(_u10_u8_n2549 ), .ZN(_u10_u8_n3088 ) );
NAND4_X1 _u10_u8_U910  ( .A1(_u10_u8_n3085 ), .A2(_u10_u8_n3086 ), .A3(_u10_u8_n3087 ), .A4(_u10_u8_n3088 ), .ZN(_u10_u8_n3084 ) );
NAND2_X1 _u10_u8_U909  ( .A1(_u10_u8_n3084 ), .A2(_u10_u8_n2803 ), .ZN(_u10_u8_n3083 ) );
NAND3_X1 _u10_u8_U908  ( .A1(_u10_u8_n3081 ), .A2(_u10_u8_n3082 ), .A3(_u10_u8_n3083 ), .ZN(_u10_u8_n3072 ) );
INV_X1 _u10_u8_U907  ( .A(_u10_u8_n2689 ), .ZN(_u10_u8_n1955 ) );
NOR3_X1 _u10_u8_U906  ( .A1(_u10_u8_n1955 ), .A2(_u10_u8_n2813 ), .A3(_u10_u8_n2488 ), .ZN(_u10_u8_n3080 ) );
NOR2_X1 _u10_u8_U905  ( .A1(_u10_u8_n3080 ), .A2(_u10_u8_n2485 ), .ZN(_u10_u8_n3073 ) );
NAND3_X1 _u10_u8_U904  ( .A1(_u10_u8_n2621 ), .A2(_u10_u8_n2202 ), .A3(_u10_u8_n3079 ), .ZN(_u10_u8_n2110 ) );
NOR2_X1 _u10_u8_U903  ( .A1(_u10_u8_n2110 ), .A2(_u10_u8_n2218 ), .ZN(_u10_u8_n2775 ) );
INV_X1 _u10_u8_U902  ( .A(_u10_u8_n2775 ), .ZN(_u10_u8_n3024 ) );
INV_X1 _u10_u8_U901  ( .A(_u10_u8_n3078 ), .ZN(_u10_u8_n2133 ) );
INV_X1 _u10_u8_U900  ( .A(_u10_u8_n2007 ), .ZN(_u10_u8_n2358 ) );
NAND2_X1 _u10_u8_U899  ( .A1(_u10_u8_n2358 ), .A2(_u10_u8_n2886 ), .ZN(_u10_u8_n2240 ) );
INV_X1 _u10_u8_U898  ( .A(_u10_u8_n2240 ), .ZN(_u10_u8_n2083 ) );
NOR3_X1 _u10_u8_U897  ( .A1(_u10_u8_n2952 ), .A2(_u10_u8_n2004 ), .A3(_u10_u8_n1891 ), .ZN(_u10_u8_n3077 ) );
NAND3_X1 _u10_u8_U896  ( .A1(_u10_u8_n2083 ), .A2(_u10_u8_n2938 ), .A3(_u10_u8_n3077 ), .ZN(_u10_u8_n1886 ) );
NOR3_X1 _u10_u8_U895  ( .A1(_u10_u8_n3024 ), .A2(_u10_u8_n2133 ), .A3(_u10_u8_n1886 ), .ZN(_u10_u8_n3075 ) );
NOR2_X1 _u10_u8_U894  ( .A1(_u10_u8_n3075 ), .A2(_u10_u8_n3076 ), .ZN(_u10_u8_n3074 ) );
NOR4_X1 _u10_u8_U893  ( .A1(_u10_u8_n3071 ), .A2(_u10_u8_n3072 ), .A3(_u10_u8_n3073 ), .A4(_u10_u8_n3074 ), .ZN(_u10_u8_n3017 ) );
INV_X1 _u10_u8_U892  ( .A(_u10_u8_n3065 ), .ZN(_u10_u8_n3043 ) );
NAND2_X1 _u10_u8_U891  ( .A1(_u10_u8_n3043 ), .A2(_u10_u8_n2106 ), .ZN(_u10_u8_n3070 ) );
NAND2_X1 _u10_u8_U890  ( .A1(_u10_u8_n3070 ), .A2(_u10_u8_n2038 ), .ZN(_u10_u8_n3068 ) );
NAND2_X1 _u10_u8_U889  ( .A1(_u10_u8_n2344 ), .A2(_u10_u8_n2584 ), .ZN(_u10_u8_n3069 ) );
NAND3_X1 _u10_u8_U888  ( .A1(_u10_u8_n3068 ), .A2(_u10_u8_n1930 ), .A3(_u10_u8_n3069 ), .ZN(_u10_u8_n3047 ) );
NAND2_X1 _u10_u8_U887  ( .A1(_u10_u8_n2835 ), .A2(_u10_u8_n2466 ), .ZN(_u10_u8_n2130 ) );
INV_X1 _u10_u8_U886  ( .A(_u10_u8_n2130 ), .ZN(_u10_u8_n2168 ) );
NAND3_X1 _u10_u8_U885  ( .A1(_u10_u8_n3067 ), .A2(_u10_u8_n2329 ), .A3(_u10_u8_n2168 ), .ZN(_u10_u8_n2665 ) );
NAND3_X1 _u10_u8_U884  ( .A1(_u10_u8_n3065 ), .A2(_u10_u8_n3066 ), .A3(_u10_u8_n2342 ), .ZN(_u10_u8_n3064 ) );
NAND3_X1 _u10_u8_U883  ( .A1(_u10_u8_n3064 ), .A2(_u10_u8_n2175 ), .A3(_u10_u8_n2987 ), .ZN(_u10_u8_n3048 ) );
NOR3_X1 _u10_u8_U882  ( .A1(_u10_u8_n1849 ), .A2(1'b0), .A3(_u10_u8_n3063 ),.ZN(_u10_u8_n3050 ) );
NOR3_X1 _u10_u8_U881  ( .A1(_u10_u8_n2406 ), .A2(1'b0), .A3(_u10_u8_n3062 ),.ZN(_u10_u8_n3060 ) );
NOR3_X1 _u10_u8_U880  ( .A1(_u10_u8_n3060 ), .A2(1'b0), .A3(_u10_u8_n3061 ),.ZN(_u10_u8_n3051 ) );
NAND2_X1 _u10_u8_U879  ( .A1(_u10_u8_n3059 ), .A2(_u10_u8_n2049 ), .ZN(_u10_u8_n3056 ) );
NAND3_X1 _u10_u8_U878  ( .A1(_u10_u8_n3056 ), .A2(_u10_u8_n3057 ), .A3(_u10_u8_n3058 ), .ZN(_u10_u8_n3054 ) );
NOR4_X1 _u10_u8_U877  ( .A1(_u10_u8_n3054 ), .A2(_u10_u8_n3055 ), .A3(_u10_u8_n2055 ), .A4(_u10_u8_n2056 ), .ZN(_u10_u8_n3053 ) );
NOR3_X1 _u10_u8_U876  ( .A1(_u10_u8_n2346 ), .A2(1'b0), .A3(_u10_u8_n3053 ),.ZN(_u10_u8_n3052 ) );
NOR3_X1 _u10_u8_U875  ( .A1(_u10_u8_n3050 ), .A2(_u10_u8_n3051 ), .A3(_u10_u8_n3052 ), .ZN(_u10_u8_n3049 ) );
NAND4_X1 _u10_u8_U874  ( .A1(_u10_u8_n3047 ), .A2(_u10_u8_n2665 ), .A3(_u10_u8_n3048 ), .A4(_u10_u8_n3049 ), .ZN(_u10_u8_n3019 ) );
NAND2_X1 _u10_u8_U873  ( .A1(_u10_u8_n2056 ), .A2(_u10_u8_n2019 ), .ZN(_u10_u8_n3046 ) );
NAND2_X1 _u10_u8_U872  ( .A1(_u10_u8_n3045 ), .A2(_u10_u8_n3046 ), .ZN(_u10_u8_n3044 ) );
NAND2_X1 _u10_u8_U871  ( .A1(_u10_u8_n3044 ), .A2(_u10_u8_n2165 ), .ZN(_u10_u8_n3028 ) );
OR2_X1 _u10_u8_U870  ( .A1(_u10_u8_n2179 ), .A2(_u10_u8_n1961 ), .ZN(_u10_u8_n3037 ) );
NAND2_X1 _u10_u8_U869  ( .A1(_u10_u8_n3043 ), .A2(_u10_u8_n2336 ), .ZN(_u10_u8_n3042 ) );
NAND2_X1 _u10_u8_U868  ( .A1(_u10_u8_n3042 ), .A2(_u10_u8_n3006 ), .ZN(_u10_u8_n3041 ) );
NAND2_X1 _u10_u8_U867  ( .A1(_u10_u8_n3040 ), .A2(_u10_u8_n3041 ), .ZN(_u10_u8_n3026 ) );
NAND4_X1 _u10_u8_U866  ( .A1(_u10_u8_n3026 ), .A2(_u10_u8_n2520 ), .A3(_u10_u8_n1962 ), .A4(_u10_u8_n1864 ), .ZN(_u10_u8_n3039 ) );
NAND2_X1 _u10_u8_U865  ( .A1(_u10_u8_n3039 ), .A2(_u10_u8_n1922 ), .ZN(_u10_u8_n3038 ) );
NAND2_X1 _u10_u8_U864  ( .A1(_u10_u8_n3037 ), .A2(_u10_u8_n3038 ), .ZN(_u10_u8_n3035 ) );
NAND2_X1 _u10_u8_U863  ( .A1(_u10_u8_n2985 ), .A2(_u10_u8_n3036 ), .ZN(_u10_u8_n2432 ) );
NAND2_X1 _u10_u8_U862  ( .A1(_u10_u8_n3035 ), .A2(_u10_u8_n2432 ), .ZN(_u10_u8_n3029 ) );
INV_X1 _u10_u8_U861  ( .A(_u10_u8_n3034 ), .ZN(_u10_u8_n2777 ) );
INV_X1 _u10_u8_U860  ( .A(_u10_u8_n2772 ), .ZN(_u10_u8_n3032 ) );
NAND2_X1 _u10_u8_U859  ( .A1(_u10_u8_n1982 ), .A2(_u10_u8_n2978 ), .ZN(_u10_u8_n3033 ) );
NAND2_X1 _u10_u8_U858  ( .A1(_u10_u8_n3032 ), .A2(_u10_u8_n3033 ), .ZN(_u10_u8_n3031 ) );
NAND2_X1 _u10_u8_U857  ( .A1(_u10_u8_n2777 ), .A2(_u10_u8_n3031 ), .ZN(_u10_u8_n3030 ) );
NAND3_X1 _u10_u8_U856  ( .A1(_u10_u8_n3028 ), .A2(_u10_u8_n3029 ), .A3(_u10_u8_n3030 ), .ZN(_u10_u8_n3020 ) );
NOR3_X1 _u10_u8_U855  ( .A1(_u10_u8_n2179 ), .A2(1'b0), .A3(_u10_u8_n2375 ),.ZN(_u10_u8_n3027 ) );
NOR2_X1 _u10_u8_U854  ( .A1(_u10_u8_n3027 ), .A2(_u10_u8_n2177 ), .ZN(_u10_u8_n3025 ) );
NOR2_X1 _u10_u8_U853  ( .A1(_u10_u8_n3025 ), .A2(_u10_u8_n3026 ), .ZN(_u10_u8_n3021 ) );
NOR2_X1 _u10_u8_U852  ( .A1(_u10_u8_n2256 ), .A2(_u10_u8_n3024 ), .ZN(_u10_u8_n3023 ) );
NOR2_X1 _u10_u8_U851  ( .A1(_u10_u8_n3023 ), .A2(_u10_u8_n1868 ), .ZN(_u10_u8_n3022 ) );
NOR4_X1 _u10_u8_U850  ( .A1(_u10_u8_n3019 ), .A2(_u10_u8_n3020 ), .A3(_u10_u8_n3021 ), .A4(_u10_u8_n3022 ), .ZN(_u10_u8_n3018 ) );
NAND4_X1 _u10_u8_U849  ( .A1(_u10_u8_n3015 ), .A2(_u10_u8_n3016 ), .A3(_u10_u8_n3017 ), .A4(_u10_u8_n3018 ), .ZN(_u10_u8_n2958 ) );
NOR2_X1 _u10_u8_U848  ( .A1(1'b0), .A2(_u10_u8_n2573 ), .ZN(_u10_u8_n3011 ));
NOR2_X1 _u10_u8_U847  ( .A1(1'b0), .A2(_u10_u8_n2359 ), .ZN(_u10_u8_n3012 ));
NOR2_X1 _u10_u8_U846  ( .A1(1'b0), .A2(_u10_u8_n1859 ), .ZN(_u10_u8_n3013 ));
NOR2_X1 _u10_u8_U845  ( .A1(1'b0), .A2(_u10_u8_n1836 ), .ZN(_u10_u8_n3014 ));
NOR4_X1 _u10_u8_U844  ( .A1(_u10_u8_n3011 ), .A2(_u10_u8_n3012 ), .A3(_u10_u8_n3013 ), .A4(_u10_u8_n3014 ), .ZN(_u10_u8_n2959 ) );
NOR2_X1 _u10_u8_U843  ( .A1(1'b0), .A2(_u10_u8_n2025 ), .ZN(_u10_u8_n3007 ));
NOR2_X1 _u10_u8_U842  ( .A1(1'b0), .A2(_u10_u8_n2085 ), .ZN(_u10_u8_n3008 ));
NOR2_X1 _u10_u8_U841  ( .A1(1'b0), .A2(_u10_u8_n2607 ), .ZN(_u10_u8_n3009 ));
NOR2_X1 _u10_u8_U840  ( .A1(1'b0), .A2(_u10_u8_n2071 ), .ZN(_u10_u8_n3010 ));
NOR4_X1 _u10_u8_U839  ( .A1(_u10_u8_n3007 ), .A2(_u10_u8_n3008 ), .A3(_u10_u8_n3009 ), .A4(_u10_u8_n3010 ), .ZN(_u10_u8_n2960 ) );
NAND2_X1 _u10_u8_U838  ( .A1(_u10_u8_n1894 ), .A2(_u10_u8_n2466 ), .ZN(_u10_u8_n3002 ) );
NAND2_X1 _u10_u8_U837  ( .A1(_u10_u8_n2830 ), .A2(_u10_u8_n2600 ), .ZN(_u10_u8_n3003 ) );
NAND2_X1 _u10_u8_U836  ( .A1(_u10_u8_n1960 ), .A2(_u10_u8_n2431 ), .ZN(_u10_u8_n3004 ) );
NAND2_X1 _u10_u8_U835  ( .A1(_u10_u8_n2002 ), .A2(_u10_u8_n3006 ), .ZN(_u10_u8_n3005 ) );
NAND4_X1 _u10_u8_U834  ( .A1(_u10_u8_n3002 ), .A2(_u10_u8_n3003 ), .A3(_u10_u8_n3004 ), .A4(_u10_u8_n3005 ), .ZN(_u10_u8_n2992 ) );
NAND2_X1 _u10_u8_U833  ( .A1(_u10_u8_n2461 ), .A2(_u10_u8_n3001 ), .ZN(_u10_u8_n2997 ) );
NAND2_X1 _u10_u8_U832  ( .A1(_u10_u8_n2999 ), .A2(_u10_u8_n3000 ), .ZN(_u10_u8_n2998 ) );
NAND2_X1 _u10_u8_U831  ( .A1(_u10_u8_n2997 ), .A2(_u10_u8_n2998 ), .ZN(_u10_u8_n2993 ) );
NOR2_X1 _u10_u8_U830  ( .A1(_u10_SYNOPSYS_UNCONNECTED_34 ), .A2(_u10_u8_n2996 ), .ZN(_u10_u8_n2995 ) );
NOR2_X1 _u10_u8_U829  ( .A1(_u10_u8_n2995 ), .A2(_u10_u8_n2126 ), .ZN(_u10_u8_n2994 ) );
NOR4_X1 _u10_u8_U828  ( .A1(_u10_u8_n2992 ), .A2(_u10_u8_n2993 ), .A3(next_ch), .A4(_u10_u8_n2994 ), .ZN(_u10_u8_n2961 ) );
NAND2_X1 _u10_u8_U827  ( .A1(_u10_u8_n2445 ), .A2(_u10_u8_n2803 ), .ZN(_u10_u8_n2988 ) );
OR2_X1 _u10_u8_U826  ( .A1(_u10_u8_n2584 ), .A2(1'b0), .ZN(_u10_u8_n2989 ));
NAND2_X1 _u10_u8_U825  ( .A1(_u10_u8_n2709 ), .A2(_u10_u8_n2080 ), .ZN(_u10_u8_n2990 ) );
NAND2_X1 _u10_u8_U824  ( .A1(_u10_u8_n2183 ), .A2(_u10_u8_n2166 ), .ZN(_u10_u8_n2991 ) );
NAND4_X1 _u10_u8_U823  ( .A1(_u10_u8_n2988 ), .A2(_u10_u8_n2989 ), .A3(_u10_u8_n2990 ), .A4(_u10_u8_n2991 ), .ZN(_u10_u8_n2963 ) );
NAND2_X1 _u10_u8_U822  ( .A1(_u10_u8_n2987 ), .A2(_u10_u8_n1930 ), .ZN(_u10_u8_n2981 ) );
NAND2_X1 _u10_u8_U821  ( .A1(_u10_u8_n2986 ), .A2(_u10_u8_n2038 ), .ZN(_u10_u8_n2982 ) );
OR2_X1 _u10_u8_U820  ( .A1(_u10_u8_n2985 ), .A2(1'b0), .ZN(_u10_u8_n2983 ));
NAND2_X1 _u10_u8_U819  ( .A1(_u10_u8_n2169 ), .A2(_u10_u8_n2113 ), .ZN(_u10_u8_n2984 ) );
NAND4_X1 _u10_u8_U818  ( .A1(_u10_u8_n2981 ), .A2(_u10_u8_n2982 ), .A3(_u10_u8_n2983 ), .A4(_u10_u8_n2984 ), .ZN(_u10_u8_n2964 ) );
NAND2_X1 _u10_u8_U817  ( .A1(_u10_u8_n2509 ), .A2(_u10_u8_n1864 ), .ZN(_u10_u8_n2973 ) );
INV_X1 _u10_u8_U816  ( .A(_u10_u8_n2980 ), .ZN(_u10_u8_n1861 ) );
NAND2_X1 _u10_u8_U815  ( .A1(_u10_u8_n1861 ), .A2(_u10_u8_n1922 ), .ZN(_u10_u8_n2974 ) );
NAND2_X1 _u10_u8_U814  ( .A1(_u10_u8_n2979 ), .A2(_u10_u8_n2405 ), .ZN(_u10_u8_n2975 ) );
NAND2_X1 _u10_u8_U813  ( .A1(_u10_u8_n2977 ), .A2(_u10_u8_n2978 ), .ZN(_u10_u8_n2976 ) );
NAND4_X1 _u10_u8_U812  ( .A1(_u10_u8_n2973 ), .A2(_u10_u8_n2974 ), .A3(_u10_u8_n2975 ), .A4(_u10_u8_n2976 ), .ZN(_u10_u8_n2965 ) );
NAND2_X1 _u10_u8_U811  ( .A1(_u10_u8_n2507 ), .A2(_u10_u8_n2972 ), .ZN(_u10_u8_n2967 ) );
NAND2_X1 _u10_u8_U810  ( .A1(_u10_u8_n2043 ), .A2(_u10_u8_n1965 ), .ZN(_u10_u8_n2968 ) );
NAND2_X1 _u10_u8_U809  ( .A1(_u10_u8_n2063 ), .A2(_u10_u8_n1853 ), .ZN(_u10_u8_n2969 ) );
NAND2_X1 _u10_u8_U808  ( .A1(_u10_u8_n2971 ), .A2(_u10_u8_n2175 ), .ZN(_u10_u8_n2970 ) );
NAND4_X1 _u10_u8_U807  ( .A1(_u10_u8_n2967 ), .A2(_u10_u8_n2968 ), .A3(_u10_u8_n2969 ), .A4(_u10_u8_n2970 ), .ZN(_u10_u8_n2966 ) );
NOR4_X1 _u10_u8_U806  ( .A1(_u10_u8_n2963 ), .A2(_u10_u8_n2964 ), .A3(_u10_u8_n2965 ), .A4(_u10_u8_n2966 ), .ZN(_u10_u8_n2962 ) );
AND4_X1 _u10_u8_U805  ( .A1(_u10_u8_n2959 ), .A2(_u10_u8_n2960 ), .A3(_u10_u8_n2961 ), .A4(_u10_u8_n2962 ), .ZN(_u10_u8_n1819 ) );
MUX2_X1 _u10_u8_U804  ( .A(_u10_u8_n2958 ), .B(_u10_SYNOPSYS_UNCONNECTED_38 ), .S(_u10_u8_n1819 ), .Z(_u10_u8_n1808 ) );
NOR2_X1 _u10_u8_U803  ( .A1(_u10_u8_n2531 ), .A2(_u10_u8_n2607 ), .ZN(_u10_u8_n1911 ) );
NAND2_X1 _u10_u8_U802  ( .A1(_u10_u8_n1911 ), .A2(_u10_u8_n2957 ), .ZN(_u10_u8_n2954 ) );
NAND2_X1 _u10_u8_U801  ( .A1(_u10_u8_n1853 ), .A2(_u10_u8_n1965 ), .ZN(_u10_u8_n2956 ) );
NAND2_X1 _u10_u8_U800  ( .A1(_u10_u8_n1966 ), .A2(_u10_u8_n2956 ), .ZN(_u10_u8_n2955 ) );
NAND2_X1 _u10_u8_U799  ( .A1(_u10_u8_n2954 ), .A2(_u10_u8_n2955 ), .ZN(_u10_u8_n2670 ) );
NOR3_X1 _u10_u8_U798  ( .A1(_u10_u8_n1852 ), .A2(1'b0), .A3(_u10_u8_n1853 ),.ZN(_u10_u8_n2708 ) );
NAND2_X1 _u10_u8_U797  ( .A1(_u10_u8_n2708 ), .A2(_u10_u8_n2080 ), .ZN(_u10_u8_n2355 ) );
NOR2_X1 _u10_u8_U796  ( .A1(_u10_u8_n2355 ), .A2(1'b0), .ZN(_u10_u8_n2599 ));
NAND2_X1 _u10_u8_U795  ( .A1(_u10_u8_n2953 ), .A2(_u10_u8_n2599 ), .ZN(_u10_u8_n2423 ) );
OR2_X1 _u10_u8_U794  ( .A1(_u10_u8_n2423 ), .A2(_u10_u8_n2359 ), .ZN(_u10_u8_n2949 ) );
NAND3_X1 _u10_u8_U793  ( .A1(_u10_u8_n2105 ), .A2(_u10_u8_n1936 ), .A3(_u10_u8_n2952 ), .ZN(_u10_u8_n2950 ) );
NAND3_X1 _u10_u8_U792  ( .A1(_u10_u8_n2549 ), .A2(_u10_u8_n1936 ), .A3(1'b0),.ZN(_u10_u8_n2096 ) );
INV_X1 _u10_u8_U791  ( .A(_u10_u8_n2096 ), .ZN(_u10_u8_n2301 ) );
NAND2_X1 _u10_u8_U790  ( .A1(_u10_u8_n2301 ), .A2(_u10_u8_n2446 ), .ZN(_u10_u8_n2368 ) );
INV_X1 _u10_u8_U789  ( .A(_u10_u8_n2368 ), .ZN(_u10_u8_n2326 ) );
NAND2_X1 _u10_u8_U788  ( .A1(_u10_u8_n2326 ), .A2(_u10_u8_n2941 ), .ZN(_u10_u8_n2800 ) );
INV_X1 _u10_u8_U787  ( .A(_u10_u8_n2800 ), .ZN(_u10_u8_n2081 ) );
NAND2_X1 _u10_u8_U786  ( .A1(_u10_u8_n2081 ), .A2(_u10_u8_n2049 ), .ZN(_u10_u8_n2855 ) );
INV_X1 _u10_u8_U785  ( .A(_u10_u8_n2855 ), .ZN(_u10_u8_n2347 ) );
NAND2_X1 _u10_u8_U784  ( .A1(_u10_u8_n2347 ), .A2(_u10_u8_n2063 ), .ZN(_u10_u8_n2951 ) );
NAND3_X1 _u10_u8_U783  ( .A1(_u10_u8_n2949 ), .A2(_u10_u8_n2950 ), .A3(_u10_u8_n2951 ), .ZN(_u10_u8_n1997 ) );
INV_X1 _u10_u8_U782  ( .A(_u10_u8_n1997 ), .ZN(_u10_u8_n2917 ) );
AND2_X1 _u10_u8_U781  ( .A1(_u10_u8_n2709 ), .A2(_u10_u8_n2708 ), .ZN(_u10_u8_n2942 ) );
INV_X1 _u10_u8_U780  ( .A(_u10_u8_n2907 ), .ZN(_u10_u8_n2737 ) );
NAND2_X1 _u10_u8_U779  ( .A1(_u10_u8_n2737 ), .A2(_u10_u8_n2803 ), .ZN(_u10_u8_n1888 ) );
NOR2_X1 _u10_u8_U778  ( .A1(_u10_u8_n2001 ), .A2(_u10_u8_n1888 ), .ZN(_u10_u8_n2943 ) );
NAND4_X1 _u10_u8_U777  ( .A1(1'b0), .A2(_u10_u8_n2078 ), .A3(_u10_u8_n2059 ),.A4(_u10_u8_n2031 ), .ZN(_u10_u8_n2578 ) );
NOR3_X1 _u10_u8_U776  ( .A1(_u10_u8_n2719 ), .A2(_u10_u8_n2130 ), .A3(_u10_u8_n2305 ), .ZN(_u10_u8_n2386 ) );
NAND2_X1 _u10_u8_U775  ( .A1(_u10_u8_n2386 ), .A2(_u10_u8_n2669 ), .ZN(_u10_u8_n2948 ) );
NAND3_X1 _u10_u8_U774  ( .A1(_u10_u8_n2578 ), .A2(_u10_u8_n2947 ), .A3(_u10_u8_n2948 ), .ZN(_u10_u8_n2750 ) );
NOR2_X1 _u10_u8_U773  ( .A1(_u10_u8_n2274 ), .A2(_u10_u8_n2852 ), .ZN(_u10_u8_n2946 ) );
NOR3_X1 _u10_u8_U772  ( .A1(_u10_u8_n2750 ), .A2(1'b0), .A3(_u10_u8_n2946 ),.ZN(_u10_u8_n2945 ) );
NOR2_X1 _u10_u8_U771  ( .A1(_u10_u8_n2945 ), .A2(_u10_u8_n2359 ), .ZN(_u10_u8_n2944 ) );
NOR3_X1 _u10_u8_U770  ( .A1(_u10_u8_n2942 ), .A2(_u10_u8_n2943 ), .A3(_u10_u8_n2944 ), .ZN(_u10_u8_n2919 ) );
NOR2_X1 _u10_u8_U769  ( .A1(_u10_u8_n2423 ), .A2(1'b0), .ZN(_u10_u8_n1979 ));
NAND3_X1 _u10_u8_U768  ( .A1(_u10_u8_n2549 ), .A2(_u10_u8_n1936 ), .A3(_u10_u8_n1979 ), .ZN(_u10_u8_n2328 ) );
INV_X1 _u10_u8_U767  ( .A(_u10_u8_n2328 ), .ZN(_u10_u8_n2554 ) );
NAND3_X1 _u10_u8_U766  ( .A1(_u10_u8_n2941 ), .A2(_u10_u8_n2446 ), .A3(_u10_u8_n2554 ), .ZN(_u10_u8_n2115 ) );
NOR2_X1 _u10_u8_U765  ( .A1(_u10_u8_n2578 ), .A2(_u10_u8_n2030 ), .ZN(_u10_u8_n2553 ) );
INV_X1 _u10_u8_U764  ( .A(_u10_u8_n2553 ), .ZN(_u10_u8_n2269 ) );
NOR2_X1 _u10_u8_U763  ( .A1(_u10_u8_n2269 ), .A2(_u10_u8_n2790 ), .ZN(_u10_u8_n2657 ) );
INV_X1 _u10_u8_U762  ( .A(_u10_u8_n2657 ), .ZN(_u10_u8_n2210 ) );
NOR2_X1 _u10_u8_U761  ( .A1(_u10_u8_n2210 ), .A2(_u10_u8_n2911 ), .ZN(_u10_u8_n2213 ) );
INV_X1 _u10_u8_U760  ( .A(_u10_u8_n2213 ), .ZN(_u10_u8_n2456 ) );
NAND2_X1 _u10_u8_U759  ( .A1(_u10_u8_n2115 ), .A2(_u10_u8_n2456 ), .ZN(_u10_u8_n2634 ) );
INV_X1 _u10_u8_U758  ( .A(_u10_u8_n2634 ), .ZN(_u10_u8_n2220 ) );
NOR2_X1 _u10_u8_U757  ( .A1(_u10_u8_n2081 ), .A2(_u10_u8_n2386 ), .ZN(_u10_u8_n2131 ) );
NAND2_X1 _u10_u8_U756  ( .A1(_u10_u8_n2940 ), .A2(_u10_u8_n2131 ), .ZN(_u10_u8_n2138 ) );
INV_X1 _u10_u8_U755  ( .A(_u10_u8_n2138 ), .ZN(_u10_u8_n2927 ) );
NAND2_X1 _u10_u8_U754  ( .A1(_u10_u8_n2220 ), .A2(_u10_u8_n2927 ), .ZN(_u10_u8_n2939 ) );
NAND2_X1 _u10_u8_U753  ( .A1(_u10_u8_n1885 ), .A2(_u10_u8_n2939 ), .ZN(_u10_u8_n2931 ) );
NAND3_X1 _u10_u8_U752  ( .A1(_u10_u8_n1859 ), .A2(_u10_u8_n2365 ), .A3(_u10_u8_n2938 ), .ZN(_u10_u8_n2935 ) );
NAND3_X1 _u10_u8_U751  ( .A1(_u10_u8_n2927 ), .A2(_u10_u8_n2937 ), .A3(_u10_u8_n2220 ), .ZN(_u10_u8_n2936 ) );
NAND2_X1 _u10_u8_U750  ( .A1(_u10_u8_n2935 ), .A2(_u10_u8_n2936 ), .ZN(_u10_u8_n2932 ) );
INV_X1 _u10_u8_U749  ( .A(_u10_u8_n1937 ), .ZN(_u10_u8_n2350 ) );
NAND2_X1 _u10_u8_U748  ( .A1(_u10_u8_n1913 ), .A2(_u10_u8_n2350 ), .ZN(_u10_u8_n2934 ) );
NAND2_X1 _u10_u8_U747  ( .A1(_u10_u8_n2386 ), .A2(_u10_u8_n2934 ), .ZN(_u10_u8_n2933 ) );
NAND3_X1 _u10_u8_U746  ( .A1(_u10_u8_n2931 ), .A2(_u10_u8_n2932 ), .A3(_u10_u8_n2933 ), .ZN(_u10_u8_n2921 ) );
OR2_X1 _u10_u8_U745  ( .A1(_u10_u8_n2213 ), .A2(_u10_u8_n2386 ), .ZN(_u10_u8_n2930 ) );
NAND2_X1 _u10_u8_U744  ( .A1(_u10_u8_n2049 ), .A2(_u10_u8_n2930 ), .ZN(_u10_u8_n2228 ) );
AND2_X1 _u10_u8_U743  ( .A1(_u10_u8_n2228 ), .A2(_u10_u8_n2699 ), .ZN(_u10_u8_n2929 ) );
NOR2_X1 _u10_u8_U742  ( .A1(_u10_u8_n2929 ), .A2(_u10_u8_n2495 ), .ZN(_u10_u8_n2922 ) );
NOR2_X1 _u10_u8_U741  ( .A1(_u10_u8_n2633 ), .A2(_u10_u8_n2877 ), .ZN(_u10_u8_n2928 ) );
NOR2_X1 _u10_u8_U740  ( .A1(_u10_u8_n2928 ), .A2(_u10_u8_n2886 ), .ZN(_u10_u8_n2923 ) );
NOR2_X1 _u10_u8_U739  ( .A1(_u10_u8_n2927 ), .A2(_u10_u8_n2531 ), .ZN(_u10_u8_n2926 ) );
NOR2_X1 _u10_u8_U738  ( .A1(_u10_u8_n2926 ), .A2(_u10_u8_n2687 ), .ZN(_u10_u8_n2925 ) );
NOR2_X1 _u10_u8_U737  ( .A1(_u10_u8_n2925 ), .A2(_u10_u8_n1849 ), .ZN(_u10_u8_n2924 ) );
NOR4_X1 _u10_u8_U736  ( .A1(_u10_u8_n2921 ), .A2(_u10_u8_n2922 ), .A3(_u10_u8_n2923 ), .A4(_u10_u8_n2924 ), .ZN(_u10_u8_n2920 ) );
NAND4_X1 _u10_u8_U735  ( .A1(_u10_u8_n2917 ), .A2(_u10_u8_n2918 ), .A3(_u10_u8_n2919 ), .A4(_u10_u8_n2920 ), .ZN(_u10_u8_n2312 ) );
NOR2_X1 _u10_u8_U734  ( .A1(_u10_u8_n2600 ), .A2(_u10_u8_n2686 ), .ZN(_u10_u8_n2401 ) );
NAND2_X1 _u10_u8_U733  ( .A1(_u10_u8_n2401 ), .A2(_u10_u8_n2549 ), .ZN(_u10_u8_n2547 ) );
INV_X1 _u10_u8_U732  ( .A(_u10_u8_n2547 ), .ZN(_u10_u8_n2794 ) );
NAND3_X1 _u10_u8_U731  ( .A1(_u10_u8_n2364 ), .A2(_u10_u8_n2667 ), .A3(_u10_u8_n2794 ), .ZN(_u10_u8_n2535 ) );
INV_X1 _u10_u8_U730  ( .A(_u10_u8_n2535 ), .ZN(_u10_u8_n2586 ) );
NAND2_X1 _u10_u8_U729  ( .A1(_u10_u8_n2586 ), .A2(_u10_u8_n2571 ), .ZN(_u10_u8_n2916 ) );
NAND2_X1 _u10_u8_U728  ( .A1(_u10_u8_n2837 ), .A2(_u10_u8_n2916 ), .ZN(_u10_u8_n2436 ) );
NAND2_X1 _u10_u8_U727  ( .A1(_u10_u8_n2915 ), .A2(_u10_u8_n2571 ), .ZN(_u10_u8_n2914 ) );
NAND2_X1 _u10_u8_U726  ( .A1(_u10_u8_n2166 ), .A2(_u10_u8_n2914 ), .ZN(_u10_u8_n2017 ) );
NOR2_X1 _u10_u8_U725  ( .A1(_u10_u8_n2485 ), .A2(_u10_u8_n1841 ), .ZN(_u10_u8_n2913 ) );
OR4_X1 _u10_u8_U724  ( .A1(_u10_u8_n2436 ), .A2(_u10_u8_n2017 ), .A3(_u10_u8_n2913 ), .A4(_u10_u8_n2442 ), .ZN(_u10_u8_n2912 ) );
NAND2_X1 _u10_u8_U723  ( .A1(_u10_u8_n2709 ), .A2(_u10_u8_n2912 ), .ZN(_u10_u8_n2888 ) );
NAND3_X1 _u10_u8_U722  ( .A1(_u10_u8_n2078 ), .A2(_u10_u8_n2031 ), .A3(1'b0),.ZN(_u10_u8_n2580 ) );
INV_X1 _u10_u8_U721  ( .A(_u10_u8_n2580 ), .ZN(_u10_u8_n2680 ) );
AND2_X1 _u10_u8_U720  ( .A1(_u10_u8_n2680 ), .A2(_u10_u8_n2668 ), .ZN(_u10_u8_n1950 ) );
NAND2_X1 _u10_u8_U719  ( .A1(_u10_u8_n1950 ), .A2(_u10_u8_n2089 ), .ZN(_u10_u8_n2095 ) );
INV_X1 _u10_u8_U718  ( .A(_u10_u8_n2095 ), .ZN(_u10_u8_n2542 ) );
NAND2_X1 _u10_u8_U717  ( .A1(_u10_u8_n2542 ), .A2(_u10_u8_n2446 ), .ZN(_u10_u8_n1887 ) );
NOR2_X1 _u10_u8_U716  ( .A1(_u10_u8_n1887 ), .A2(_u10_u8_n2911 ), .ZN(_u10_u8_n2114 ) );
INV_X1 _u10_u8_U715  ( .A(_u10_u8_n2114 ), .ZN(_u10_u8_n1940 ) );
NAND3_X1 _u10_u8_U714  ( .A1(_u10_u8_n2535 ), .A2(_u10_u8_n1940 ), .A3(_u10_u8_n2910 ), .ZN(_u10_u8_n2524 ) );
NAND2_X1 _u10_u8_U713  ( .A1(_u10_u8_n2524 ), .A2(_u10_u8_n2488 ), .ZN(_u10_u8_n2889 ) );
NAND2_X1 _u10_u8_U712  ( .A1(_u10_u8_n2220 ), .A2(_u10_u8_n1940 ), .ZN(_u10_u8_n2763 ) );
NOR2_X1 _u10_u8_U711  ( .A1(_u10_u8_n2763 ), .A2(_u10_u8_n2586 ), .ZN(_u10_u8_n2808 ) );
NOR2_X1 _u10_u8_U710  ( .A1(_u10_u8_n2808 ), .A2(_u10_u8_n2350 ), .ZN(_u10_u8_n2908 ) );
NOR2_X1 _u10_u8_U709  ( .A1(_u10_u8_n2544 ), .A2(_u10_u8_n1950 ), .ZN(_u10_u8_n2899 ) );
NOR2_X1 _u10_u8_U708  ( .A1(_u10_u8_n2899 ), .A2(_u10_u8_n2159 ), .ZN(_u10_u8_n2909 ) );
NOR2_X1 _u10_u8_U707  ( .A1(_u10_u8_n2908 ), .A2(_u10_u8_n2909 ), .ZN(_u10_u8_n2890 ) );
NOR3_X1 _u10_u8_U706  ( .A1(_u10_u8_n2547 ), .A2(_u10_u8_n1846 ), .A3(_u10_u8_n2907 ), .ZN(_u10_u8_n2892 ) );
NOR3_X1 _u10_u8_U705  ( .A1(_u10_u8_n2240 ), .A2(_u10_u8_n2377 ), .A3(_u10_u8_n1911 ), .ZN(_u10_u8_n2906 ) );
NOR2_X1 _u10_u8_U704  ( .A1(_u10_u8_n2906 ), .A2(_u10_u8_n2535 ), .ZN(_u10_u8_n2893 ) );
NAND2_X1 _u10_u8_U703  ( .A1(_u10_u8_n2554 ), .A2(_u10_u8_n2446 ), .ZN(_u10_u8_n2903 ) );
AND3_X1 _u10_u8_U702  ( .A1(_u10_u8_n2210 ), .A2(_u10_u8_n2905 ), .A3(_u10_u8_n1887 ), .ZN(_u10_u8_n2904 ) );
NAND4_X1 _u10_u8_U701  ( .A1(_u10_u8_n2902 ), .A2(_u10_u8_n2498 ), .A3(_u10_u8_n2903 ), .A4(_u10_u8_n2904 ), .ZN(_u10_u8_n2788 ) );
INV_X1 _u10_u8_U700  ( .A(_u10_u8_n2788 ), .ZN(_u10_u8_n2901 ) );
NOR2_X1 _u10_u8_U699  ( .A1(_u10_u8_n2901 ), .A2(_u10_u8_n1888 ), .ZN(_u10_u8_n2894 ) );
NOR2_X1 _u10_u8_U698  ( .A1(_u10_u8_n2401 ), .A2(_u10_u8_n2553 ), .ZN(_u10_u8_n2900 ) );
NOR2_X1 _u10_u8_U697  ( .A1(_u10_u8_n2900 ), .A2(_u10_u8_n1954 ), .ZN(_u10_u8_n2897 ) );
NOR2_X1 _u10_u8_U696  ( .A1(1'b0), .A2(_u10_u8_n2899 ), .ZN(_u10_u8_n2898 ));
NOR2_X1 _u10_u8_U695  ( .A1(_u10_u8_n2897 ), .A2(_u10_u8_n2898 ), .ZN(_u10_u8_n2896 ) );
NOR2_X1 _u10_u8_U694  ( .A1(_u10_u8_n2896 ), .A2(_u10_u8_n1843 ), .ZN(_u10_u8_n2895 ) );
NOR4_X1 _u10_u8_U693  ( .A1(_u10_u8_n2892 ), .A2(_u10_u8_n2893 ), .A3(_u10_u8_n2894 ), .A4(_u10_u8_n2895 ), .ZN(_u10_u8_n2891 ) );
NAND4_X1 _u10_u8_U692  ( .A1(_u10_u8_n2888 ), .A2(_u10_u8_n2889 ), .A3(_u10_u8_n2890 ), .A4(_u10_u8_n2891 ), .ZN(_u10_u8_n2610 ) );
NOR4_X1 _u10_u8_U691  ( .A1(_u10_u8_n2670 ), .A2(_u10_u8_n2312 ), .A3(_u10_u8_n2610 ), .A4(_u10_u8_n2887 ), .ZN(_u10_u8_n2724 ) );
NOR2_X1 _u10_u8_U690  ( .A1(_u10_u8_n2883 ), .A2(_u10_u8_n2535 ), .ZN(_u10_u8_n2861 ) );
NOR2_X1 _u10_u8_U689  ( .A1(_u10_u8_n1855 ), .A2(_u10_u8_n1869 ), .ZN(_u10_u8_n2862 ) );
NOR2_X1 _u10_u8_U688  ( .A1(_u10_u8_n2886 ), .A2(_u10_u8_n2695 ), .ZN(_u10_u8_n2863 ) );
NAND2_X1 _u10_u8_U687  ( .A1(_u10_u8_n2813 ), .A2(_u10_u8_n2885 ), .ZN(_u10_u8_n2864 ) );
NAND2_X1 _u10_u8_U686  ( .A1(_u10_u8_n2114 ), .A2(_u10_u8_n2884 ), .ZN(_u10_u8_n2865 ) );
NAND2_X1 _u10_u8_U685  ( .A1(1'b0), .A2(_u10_u8_n2667 ), .ZN(_u10_u8_n2112 ));
NOR3_X1 _u10_u8_U684  ( .A1(_u10_u8_n2883 ), .A2(_u10_u8_n2112 ), .A3(_u10_u8_n2719 ), .ZN(_u10_u8_n2878 ) );
INV_X1 _u10_u8_U683  ( .A(_u10_u8_n2112 ), .ZN(_u10_u8_n1856 ) );
NAND2_X1 _u10_u8_U682  ( .A1(_u10_u8_n2364 ), .A2(_u10_u8_n1856 ), .ZN(_u10_u8_n2882 ) );
NAND2_X1 _u10_u8_U681  ( .A1(_u10_u8_n2882 ), .A2(_u10_u8_n1869 ), .ZN(_u10_u8_n2050 ) );
INV_X1 _u10_u8_U680  ( .A(_u10_u8_n2050 ), .ZN(_u10_u8_n1939 ) );
NOR2_X1 _u10_u8_U679  ( .A1(_u10_u8_n1939 ), .A2(_u10_u8_n1841 ), .ZN(_u10_u8_n2881 ) );
NOR2_X1 _u10_u8_U678  ( .A1(_u10_u8_n2881 ), .A2(_u10_u8_n2840 ), .ZN(_u10_u8_n2880 ) );
NOR2_X1 _u10_u8_U677  ( .A1(_u10_u8_n2880 ), .A2(_u10_u8_n1836 ), .ZN(_u10_u8_n2879 ) );
NOR2_X1 _u10_u8_U676  ( .A1(_u10_u8_n2878 ), .A2(_u10_u8_n2879 ), .ZN(_u10_u8_n2866 ) );
NOR2_X1 _u10_u8_U675  ( .A1(_u10_u8_n2081 ), .A2(_u10_u8_n2877 ), .ZN(_u10_u8_n1840 ) );
NAND2_X1 _u10_u8_U674  ( .A1(_u10_u8_n1840 ), .A2(_u10_u8_n2115 ), .ZN(_u10_u8_n1873 ) );
NAND2_X1 _u10_u8_U673  ( .A1(_u10_u8_n2695 ), .A2(_u10_u8_n1940 ), .ZN(_u10_u8_n1874 ) );
NOR3_X1 _u10_u8_U672  ( .A1(_u10_u8_n2050 ), .A2(_u10_u8_n1873 ), .A3(_u10_u8_n1874 ), .ZN(_u10_u8_n2876 ) );
NOR2_X1 _u10_u8_U671  ( .A1(_u10_u8_n2876 ), .A2(_u10_u8_n1913 ), .ZN(_u10_u8_n2868 ) );
NAND2_X1 _u10_u8_U670  ( .A1(_u10_u8_n2875 ), .A2(_u10_u8_n2466 ), .ZN(_u10_u8_n2872 ) );
INV_X1 _u10_u8_U669  ( .A(_u10_u8_n1979 ), .ZN(_u10_u8_n2746 ) );
NAND2_X1 _u10_u8_U668  ( .A1(_u10_u8_n2874 ), .A2(_u10_u8_n2746 ), .ZN(_u10_u8_n1935 ) );
NAND3_X1 _u10_u8_U667  ( .A1(_u10_u8_n1935 ), .A2(_u10_u8_n1936 ), .A3(_u10_u8_n2467 ), .ZN(_u10_u8_n2873 ) );
NAND2_X1 _u10_u8_U666  ( .A1(_u10_u8_n2872 ), .A2(_u10_u8_n2873 ), .ZN(_u10_u8_n2264 ) );
AND2_X1 _u10_u8_U665  ( .A1(_u10_u8_n2264 ), .A2(_u10_u8_n2461 ), .ZN(_u10_u8_n2869 ) );
AND2_X1 _u10_u8_U664  ( .A1(_u10_u8_n1966 ), .A2(_u10_u8_n2761 ), .ZN(_u10_u8_n2870 ) );
NOR2_X1 _u10_u8_U663  ( .A1(_u10_u8_n2159 ), .A2(_u10_u8_n2163 ), .ZN(_u10_u8_n2871 ) );
NOR4_X1 _u10_u8_U662  ( .A1(_u10_u8_n2868 ), .A2(_u10_u8_n2869 ), .A3(_u10_u8_n2870 ), .A4(_u10_u8_n2871 ), .ZN(_u10_u8_n2867 ) );
NAND4_X1 _u10_u8_U661  ( .A1(_u10_u8_n2864 ), .A2(_u10_u8_n2865 ), .A3(_u10_u8_n2866 ), .A4(_u10_u8_n2867 ), .ZN(_u10_u8_n1992 ) );
NOR4_X1 _u10_u8_U660  ( .A1(_u10_u8_n2861 ), .A2(_u10_u8_n2862 ), .A3(_u10_u8_n2863 ), .A4(_u10_u8_n1992 ), .ZN(_u10_u8_n2725 ) );
NAND2_X1 _u10_u8_U659  ( .A1(_u10_u8_n2364 ), .A2(_u10_u8_n1846 ), .ZN(_u10_u8_n2744 ) );
NAND4_X1 _u10_u8_U658  ( .A1(_u10_u8_n2765 ), .A2(_u10_u8_n1939 ), .A3(_u10_u8_n2744 ), .A4(_u10_u8_n2535 ), .ZN(_u10_u8_n2860 ) );
NAND2_X1 _u10_u8_U657  ( .A1(_u10_u8_n2049 ), .A2(_u10_u8_n2860 ), .ZN(_u10_u8_n2856 ) );
NOR4_X1 _u10_u8_U656  ( .A1(1'b0), .A2(_u10_u8_n2858 ), .A3(_u10_u8_n2859 ),.A4(_u10_u8_n2051 ), .ZN(_u10_u8_n2857 ) );
NAND4_X1 _u10_u8_U655  ( .A1(_u10_u8_n2228 ), .A2(_u10_u8_n2855 ), .A3(_u10_u8_n2856 ), .A4(_u10_u8_n2857 ), .ZN(_u10_u8_n2854 ) );
NAND2_X1 _u10_u8_U654  ( .A1(_u10_u8_n2043 ), .A2(_u10_u8_n2854 ), .ZN(_u10_u8_n2821 ) );
INV_X1 _u10_u8_U653  ( .A(_u10_u8_n2071 ), .ZN(_u10_u8_n2279 ) );
INV_X1 _u10_u8_U652  ( .A(_u10_u8_n2599 ), .ZN(_u10_u8_n2357 ) );
OR2_X1 _u10_u8_U651  ( .A1(_u10_u8_n2744 ), .A2(_u10_u8_n2853 ), .ZN(_u10_u8_n2844 ) );
NAND2_X1 _u10_u8_U650  ( .A1(_u10_u8_n2131 ), .A2(_u10_u8_n2852 ), .ZN(_u10_u8_n2851 ) );
NAND2_X1 _u10_u8_U649  ( .A1(_u10_u8_n2082 ), .A2(_u10_u8_n2851 ), .ZN(_u10_u8_n2848 ) );
NAND2_X1 _u10_u8_U648  ( .A1(_u10_u8_n2850 ), .A2(_u10_u8_n2600 ), .ZN(_u10_u8_n2849 ) );
NAND3_X1 _u10_u8_U647  ( .A1(_u10_u8_n2848 ), .A2(_u10_u8_n2077 ), .A3(_u10_u8_n2849 ), .ZN(_u10_u8_n2287 ) );
NAND2_X1 _u10_u8_U646  ( .A1(_u10_u8_n2082 ), .A2(_u10_u8_n2050 ), .ZN(_u10_u8_n2847 ) );
NAND2_X1 _u10_u8_U645  ( .A1(_u10_u8_n2846 ), .A2(_u10_u8_n2847 ), .ZN(_u10_u8_n2074 ) );
NOR3_X1 _u10_u8_U644  ( .A1(_u10_u8_n2287 ), .A2(_u10_u8_n2596 ), .A3(_u10_u8_n2074 ), .ZN(_u10_u8_n2845 ) );
NAND4_X1 _u10_u8_U643  ( .A1(_u10_u8_n2357 ), .A2(_u10_u8_n2837 ), .A3(_u10_u8_n2844 ), .A4(_u10_u8_n2845 ), .ZN(_u10_u8_n2843 ) );
NAND2_X1 _u10_u8_U642  ( .A1(_u10_u8_n2279 ), .A2(_u10_u8_n2843 ), .ZN(_u10_u8_n2822 ) );
NOR3_X1 _u10_u8_U641  ( .A1(_u10_u8_n1925 ), .A2(_u10_u8_n2842 ), .A3(_u10_u8_n2686 ), .ZN(_u10_u8_n2841 ) );
NOR3_X1 _u10_u8_U640  ( .A1(_u10_u8_n2840 ), .A2(_u10_u8_n2599 ), .A3(_u10_u8_n2841 ), .ZN(_u10_u8_n2839 ) );
AND4_X1 _u10_u8_U639  ( .A1(_u10_u8_n2836 ), .A2(_u10_u8_n2837 ), .A3(_u10_u8_n2838 ), .A4(_u10_u8_n2839 ), .ZN(_u10_u8_n2454 ) );
NOR2_X1 _u10_u8_U638  ( .A1(_u10_u8_n2719 ), .A2(_u10_u8_n2835 ), .ZN(_u10_u8_n2773 ) );
NOR2_X1 _u10_u8_U637  ( .A1(_u10_u8_n2138 ), .A2(_u10_u8_n2773 ), .ZN(_u10_u8_n2814 ) );
NAND2_X1 _u10_u8_U636  ( .A1(_u10_u8_n2814 ), .A2(_u10_u8_n1869 ), .ZN(_u10_u8_n2834 ) );
NAND2_X1 _u10_u8_U635  ( .A1(_u10_u8_n2833 ), .A2(_u10_u8_n2834 ), .ZN(_u10_u8_n2832 ) );
NAND2_X1 _u10_u8_U634  ( .A1(_u10_u8_n2454 ), .A2(_u10_u8_n2832 ), .ZN(_u10_u8_n2831 ) );
NAND2_X1 _u10_u8_U633  ( .A1(_u10_u8_n2830 ), .A2(_u10_u8_n2831 ), .ZN(_u10_u8_n2823 ) );
INV_X1 _u10_u8_U632  ( .A(_u10_u8_n2025 ), .ZN(_u10_u8_n2470 ) );
NAND2_X1 _u10_u8_U631  ( .A1(_u10_u8_n1979 ), .A2(_u10_u8_n1936 ), .ZN(_u10_u8_n2829 ) );
AND2_X1 _u10_u8_U630  ( .A1(_u10_u8_n2828 ), .A2(_u10_u8_n2829 ), .ZN(_u10_u8_n2469 ) );
NAND2_X1 _u10_u8_U629  ( .A1(_u10_u8_n2469 ), .A2(_u10_u8_n2269 ), .ZN(_u10_u8_n2161 ) );
INV_X1 _u10_u8_U628  ( .A(_u10_u8_n2161 ), .ZN(_u10_u8_n2276 ) );
NOR2_X1 _u10_u8_U627  ( .A1(_u10_u8_n2274 ), .A2(_u10_u8_n2719 ), .ZN(_u10_u8_n2827 ) );
NOR3_X1 _u10_u8_U626  ( .A1(_u10_u8_n2827 ), .A2(_u10_u8_n2742 ), .A3(_u10_u8_n2680 ), .ZN(_u10_u8_n2826 ) );
NAND3_X1 _u10_u8_U625  ( .A1(_u10_u8_n2276 ), .A2(_u10_u8_n2108 ), .A3(_u10_u8_n2826 ), .ZN(_u10_u8_n2825 ) );
NAND2_X1 _u10_u8_U624  ( .A1(_u10_u8_n2470 ), .A2(_u10_u8_n2825 ), .ZN(_u10_u8_n2824 ) );
NAND4_X1 _u10_u8_U623  ( .A1(_u10_u8_n2821 ), .A2(_u10_u8_n2822 ), .A3(_u10_u8_n2823 ), .A4(_u10_u8_n2824 ), .ZN(_u10_u8_n2804 ) );
NAND2_X1 _u10_u8_U622  ( .A1(_u10_u8_n2131 ), .A2(_u10_u8_n2744 ), .ZN(_u10_u8_n2820 ) );
NAND2_X1 _u10_u8_U621  ( .A1(_u10_u8_n2571 ), .A2(_u10_u8_n2820 ), .ZN(_u10_u8_n2817 ) );
NOR2_X1 _u10_u8_U620  ( .A1(_u10_u8_n2819 ), .A2(_u10_u8_n2436 ), .ZN(_u10_u8_n2818 ) );
NAND4_X1 _u10_u8_U619  ( .A1(_u10_u8_n2437 ), .A2(_u10_u8_n2355 ), .A3(_u10_u8_n2817 ), .A4(_u10_u8_n2818 ), .ZN(_u10_u8_n2816 ) );
NAND2_X1 _u10_u8_U618  ( .A1(_u10_u8_n2815 ), .A2(_u10_u8_n2816 ), .ZN(_u10_u8_n2809 ) );
INV_X1 _u10_u8_U617  ( .A(_u10_u8_n2814 ), .ZN(_u10_u8_n2812 ) );
OR2_X1 _u10_u8_U616  ( .A1(_u10_u8_n1911 ), .A2(_u10_u8_n2813 ), .ZN(_u10_u8_n1884 ) );
NAND2_X1 _u10_u8_U615  ( .A1(_u10_u8_n2812 ), .A2(_u10_u8_n1884 ), .ZN(_u10_u8_n2810 ) );
NOR2_X1 _u10_u8_U614  ( .A1(_u10_u8_n1894 ), .A2(_u10_u8_n2461 ), .ZN(_u10_u8_n1948 ) );
OR2_X1 _u10_u8_U613  ( .A1(_u10_u8_n1847 ), .A2(_u10_u8_n1948 ), .ZN(_u10_u8_n2811 ) );
NAND3_X1 _u10_u8_U612  ( .A1(_u10_u8_n2809 ), .A2(_u10_u8_n2810 ), .A3(_u10_u8_n2811 ), .ZN(_u10_u8_n2805 ) );
NOR2_X1 _u10_u8_U611  ( .A1(_u10_u8_n2808 ), .A2(_u10_u8_n2775 ), .ZN(_u10_u8_n2806 ) );
AND2_X1 _u10_u8_U610  ( .A1(_u10_u8_n2721 ), .A2(_u10_u8_n1911 ), .ZN(_u10_u8_n2807 ) );
NOR4_X1 _u10_u8_U609  ( .A1(_u10_u8_n2804 ), .A2(_u10_u8_n2805 ), .A3(_u10_u8_n2806 ), .A4(_u10_u8_n2807 ), .ZN(_u10_u8_n2726 ) );
NAND2_X1 _u10_u8_U608  ( .A1(_u10_u8_n2803 ), .A2(_u10_u8_n2112 ), .ZN(_u10_u8_n2802 ) );
NAND2_X1 _u10_u8_U607  ( .A1(_u10_u8_n2364 ), .A2(_u10_u8_n2802 ), .ZN(_u10_u8_n2801 ) );
NAND2_X1 _u10_u8_U606  ( .A1(_u10_u8_n2800 ), .A2(_u10_u8_n2801 ), .ZN(_u10_u8_n2799 ) );
NAND2_X1 _u10_u8_U605  ( .A1(_u10_u8_n1937 ), .A2(_u10_u8_n2799 ), .ZN(_u10_u8_n2780 ) );
NAND2_X1 _u10_u8_U604  ( .A1(_u10_u8_n2775 ), .A2(_u10_u8_n2798 ), .ZN(_u10_u8_n2796 ) );
INV_X1 _u10_u8_U603  ( .A(_u10_u8_n2131 ), .ZN(_u10_u8_n2797 ) );
NAND2_X1 _u10_u8_U602  ( .A1(_u10_u8_n2796 ), .A2(_u10_u8_n2797 ), .ZN(_u10_u8_n2781 ) );
OR4_X1 _u10_u8_U601  ( .A1(_u10_u8_n2795 ), .A2(_u10_u8_n2303 ), .A3(_u10_u8_n2553 ), .A4(_u10_u8_n2554 ), .ZN(_u10_u8_n2792 ) );
NAND3_X1 _u10_u8_U600  ( .A1(_u10_u8_n1847 ), .A2(_u10_u8_n2097 ), .A3(_u10_u8_n2096 ), .ZN(_u10_u8_n2793 ) );
NOR4_X1 _u10_u8_U599  ( .A1(_u10_u8_n2792 ), .A2(_u10_u8_n2793 ), .A3(_u10_u8_n2542 ), .A4(_u10_u8_n2794 ), .ZN(_u10_u8_n2791 ) );
NOR2_X1 _u10_u8_U598  ( .A1(_u10_u8_n2791 ), .A2(_u10_u8_n2085 ), .ZN(_u10_u8_n2783 ) );
NAND2_X1 _u10_u8_U597  ( .A1(_u10_u8_n2114 ), .A2(_u10_u8_n2049 ), .ZN(_u10_u8_n2700 ) );
INV_X1 _u10_u8_U596  ( .A(_u10_u8_n2700 ), .ZN(_u10_u8_n2784 ) );
NAND4_X1 _u10_u8_U595  ( .A1(_u10_u8_n2001 ), .A2(_u10_u8_n2547 ), .A3(_u10_u8_n2368 ), .A4(_u10_u8_n1847 ), .ZN(_u10_u8_n2787 ) );
NOR4_X1 _u10_u8_U594  ( .A1(_u10_u8_n2787 ), .A2(_u10_u8_n2788 ), .A3(_u10_u8_n2789 ), .A4(_u10_u8_n2790 ), .ZN(_u10_u8_n2786 ) );
NOR2_X1 _u10_u8_U593  ( .A1(_u10_u8_n2786 ), .A2(_u10_u8_n2000 ), .ZN(_u10_u8_n2785 ) );
NOR3_X1 _u10_u8_U592  ( .A1(_u10_u8_n2783 ), .A2(_u10_u8_n2784 ), .A3(_u10_u8_n2785 ), .ZN(_u10_u8_n2782 ) );
NAND3_X1 _u10_u8_U591  ( .A1(_u10_u8_n2780 ), .A2(_u10_u8_n2781 ), .A3(_u10_u8_n2782 ), .ZN(_u10_u8_n2728 ) );
OR3_X1 _u10_u8_U590  ( .A1(_u10_u8_n2138 ), .A2(_u10_u8_n2633 ), .A3(_u10_u8_n2779 ), .ZN(_u10_u8_n2778 ) );
NAND2_X1 _u10_u8_U589  ( .A1(_u10_u8_n2777 ), .A2(_u10_u8_n2778 ), .ZN(_u10_u8_n2767 ) );
NAND3_X1 _u10_u8_U588  ( .A1(_u10_u8_n2775 ), .A2(_u10_u8_n2083 ), .A3(_u10_u8_n2776 ), .ZN(_u10_u8_n2774 ) );
NAND2_X1 _u10_u8_U587  ( .A1(_u10_u8_n2773 ), .A2(_u10_u8_n2774 ), .ZN(_u10_u8_n2768 ) );
NAND2_X1 _u10_u8_U586  ( .A1(_u10_u8_n2218 ), .A2(_u10_u8_n2772 ), .ZN(_u10_u8_n2769 ) );
NAND2_X1 _u10_u8_U585  ( .A1(_u10_u8_n2302 ), .A2(_u10_u8_n2467 ), .ZN(_u10_u8_n2771 ) );
NAND2_X1 _u10_u8_U584  ( .A1(_u10_u8_n2461 ), .A2(_u10_u8_n2771 ), .ZN(_u10_u8_n2770 ) );
NAND4_X1 _u10_u8_U583  ( .A1(_u10_u8_n2767 ), .A2(_u10_u8_n2768 ), .A3(_u10_u8_n2769 ), .A4(_u10_u8_n2770 ), .ZN(_u10_u8_n2729 ) );
NAND3_X1 _u10_u8_U582  ( .A1(_u10_u8_n2668 ), .A2(_u10_u8_n2600 ), .A3(_u10_u8_n2276 ), .ZN(_u10_u8_n2766 ) );
NAND2_X1 _u10_u8_U581  ( .A1(_u10_u8_n1894 ), .A2(_u10_u8_n2766 ), .ZN(_u10_u8_n2753 ) );
NAND3_X1 _u10_u8_U580  ( .A1(_u10_u8_n2456 ), .A2(_u10_u8_n2744 ), .A3(_u10_u8_n2765 ), .ZN(_u10_u8_n2764 ) );
NAND2_X1 _u10_u8_U579  ( .A1(_u10_u8_n2377 ), .A2(_u10_u8_n2764 ), .ZN(_u10_u8_n2754 ) );
NAND2_X1 _u10_u8_U578  ( .A1(_u10_u8_n2763 ), .A2(_u10_u8_n2007 ), .ZN(_u10_u8_n2755 ) );
NOR2_X1 _u10_u8_U577  ( .A1(_u10_u8_n2531 ), .A2(_u10_u8_n2744 ), .ZN(_u10_u8_n2760 ) );
INV_X1 _u10_u8_U576  ( .A(_u10_u8_n2762 ), .ZN(_u10_u8_n2189 ) );
NOR3_X1 _u10_u8_U575  ( .A1(_u10_u8_n2760 ), .A2(_u10_u8_n2761 ), .A3(_u10_u8_n2189 ), .ZN(_u10_u8_n2759 ) );
NOR2_X1 _u10_u8_U574  ( .A1(_u10_u8_n2759 ), .A2(_u10_u8_n1849 ), .ZN(_u10_u8_n2757 ) );
NOR2_X1 _u10_u8_U573  ( .A1(_u10_u8_n1817 ), .A2(_u10_u8_n2665 ), .ZN(_u10_u8_n2758 ) );
NOR2_X1 _u10_u8_U572  ( .A1(_u10_u8_n2757 ), .A2(_u10_u8_n2758 ), .ZN(_u10_u8_n2756 ) );
NAND4_X1 _u10_u8_U571  ( .A1(_u10_u8_n2753 ), .A2(_u10_u8_n2754 ), .A3(_u10_u8_n2755 ), .A4(_u10_u8_n2756 ), .ZN(_u10_u8_n2730 ) );
INV_X1 _u10_u8_U570  ( .A(_u10_u8_n2359 ), .ZN(_u10_u8_n1899 ) );
NAND4_X1 _u10_u8_U569  ( .A1(_u10_u8_n2078 ), .A2(_u10_u8_n2580 ), .A3(_u10_u8_n2748 ), .A4(_u10_u8_n2752 ), .ZN(_u10_u8_n2751 ) );
NAND2_X1 _u10_u8_U568  ( .A1(_u10_u8_n1899 ), .A2(_u10_u8_n2751 ), .ZN(_u10_u8_n2732 ) );
INV_X1 _u10_u8_U567  ( .A(_u10_u8_n2750 ), .ZN(_u10_u8_n2379 ) );
NAND3_X1 _u10_u8_U566  ( .A1(_u10_u8_n1856 ), .A2(_u10_u8_n2669 ), .A3(_u10_u8_n2364 ), .ZN(_u10_u8_n2749 ) );
AND2_X1 _u10_u8_U565  ( .A1(_u10_u8_n2748 ), .A2(_u10_u8_n2749 ), .ZN(_u10_u8_n2034 ) );
NAND2_X1 _u10_u8_U564  ( .A1(_u10_u8_n2105 ), .A2(_u10_u8_n2669 ), .ZN(_u10_u8_n2745 ) );
AND3_X1 _u10_u8_U563  ( .A1(_u10_u8_n2745 ), .A2(_u10_u8_n2746 ), .A3(_u10_u8_n2747 ), .ZN(_u10_u8_n2380 ) );
NOR2_X1 _u10_u8_U562  ( .A1(_u10_u8_n2274 ), .A2(_u10_u8_n2744 ), .ZN(_u10_u8_n2743 ) );
NOR4_X1 _u10_u8_U561  ( .A1(_u10_u8_n2742 ), .A2(_u10_u8_n2680 ), .A3(_u10_u8_n2743 ), .A4(_u10_u8_n2428 ), .ZN(_u10_u8_n2741 ) );
NAND4_X1 _u10_u8_U560  ( .A1(_u10_u8_n2379 ), .A2(_u10_u8_n2034 ), .A3(_u10_u8_n2380 ), .A4(_u10_u8_n2741 ), .ZN(_u10_u8_n2740 ) );
NAND2_X1 _u10_u8_U559  ( .A1(_u10_u8_n1967 ), .A2(_u10_u8_n2740 ), .ZN(_u10_u8_n2733 ) );
NAND3_X1 _u10_u8_U558  ( .A1(_u10_u8_n2739 ), .A2(_u10_u8_n2368 ), .A3(_u10_u8_n2255 ), .ZN(_u10_u8_n2738 ) );
NAND2_X1 _u10_u8_U557  ( .A1(_u10_u8_n2737 ), .A2(_u10_u8_n2738 ), .ZN(_u10_u8_n2734 ) );
NAND2_X1 _u10_u8_U556  ( .A1(_u10_u8_n2736 ), .A2(_u10_u8_n2524 ), .ZN(_u10_u8_n2735 ) );
NAND4_X1 _u10_u8_U555  ( .A1(_u10_u8_n2732 ), .A2(_u10_u8_n2733 ), .A3(_u10_u8_n2734 ), .A4(_u10_u8_n2735 ), .ZN(_u10_u8_n2731 ) );
NOR4_X1 _u10_u8_U554  ( .A1(_u10_u8_n2728 ), .A2(_u10_u8_n2729 ), .A3(_u10_u8_n2730 ), .A4(_u10_u8_n2731 ), .ZN(_u10_u8_n2727 ) );
NAND4_X1 _u10_u8_U553  ( .A1(_u10_u8_n2724 ), .A2(_u10_u8_n2725 ), .A3(_u10_u8_n2726 ), .A4(_u10_u8_n2727 ), .ZN(_u10_u8_n2723 ) );
MUX2_X1 _u10_u8_U552  ( .A(_u10_u8_n2723 ), .B(_u10_SYNOPSYS_UNCONNECTED_34 ), .S(_u10_u8_n1819 ), .Z(_u10_u8_n1809 ) );
NAND2_X1 _u10_u8_U551  ( .A1(_u10_u8_n2002 ), .A2(_u10_u8_n2722 ), .ZN(_u10_u8_n2713 ) );
NAND2_X1 _u10_u8_U550  ( .A1(_u10_u8_n2720 ), .A2(_u10_u8_n2721 ), .ZN(_u10_u8_n2714 ) );
NAND2_X1 _u10_u8_U549  ( .A1(_u10_u8_n2256 ), .A2(_u10_u8_n2719 ), .ZN(_u10_u8_n2715 ) );
NOR2_X1 _u10_u8_U548  ( .A1(_u10_u8_n2106 ), .A2(_u10_u8_n2037 ), .ZN(_u10_u8_n2717 ) );
AND2_X1 _u10_u8_U547  ( .A1(_u10_u8_n1966 ), .A2(_u10_u8_n2054 ), .ZN(_u10_u8_n2718 ) );
NOR2_X1 _u10_u8_U546  ( .A1(_u10_u8_n2717 ), .A2(_u10_u8_n2718 ), .ZN(_u10_u8_n2716 ) );
NAND4_X1 _u10_u8_U545  ( .A1(_u10_u8_n2713 ), .A2(_u10_u8_n2714 ), .A3(_u10_u8_n2715 ), .A4(_u10_u8_n2716 ), .ZN(_u10_u8_n2608 ) );
NAND2_X1 _u10_u8_U544  ( .A1(1'b0), .A2(_u10_u8_n2669 ), .ZN(_u10_u8_n2385 ));
INV_X1 _u10_u8_U543  ( .A(_u10_u8_n2385 ), .ZN(_u10_u8_n1977 ) );
NAND2_X1 _u10_u8_U542  ( .A1(_u10_u8_n1977 ), .A2(_u10_u8_n2668 ), .ZN(_u10_u8_n2712 ) );
NAND2_X1 _u10_u8_U541  ( .A1(_u10_u8_n2712 ), .A2(_u10_u8_n2092 ), .ZN(_u10_u8_n1844 ) );
NAND2_X1 _u10_u8_U540  ( .A1(_u10_u8_n1894 ), .A2(_u10_u8_n1844 ), .ZN(_u10_u8_n2705 ) );
NAND2_X1 _u10_u8_U539  ( .A1(_u10_u8_n1894 ), .A2(_u10_u8_n2305 ), .ZN(_u10_u8_n2711 ) );
NAND2_X1 _u10_u8_U538  ( .A1(_u10_u8_n2711 ), .A2(_u10_u8_n2025 ), .ZN(_u10_u8_n1932 ) );
NAND2_X1 _u10_u8_U537  ( .A1(_u10_u8_n2710 ), .A2(_u10_u8_n1932 ), .ZN(_u10_u8_n2706 ) );
NAND2_X1 _u10_u8_U536  ( .A1(_u10_u8_n2708 ), .A2(_u10_u8_n2709 ), .ZN(_u10_u8_n2707 ) );
NAND3_X1 _u10_u8_U535  ( .A1(_u10_u8_n2705 ), .A2(_u10_u8_n2706 ), .A3(_u10_u8_n2707 ), .ZN(_u10_u8_n2701 ) );
NOR2_X1 _u10_u8_U534  ( .A1(_u10_u8_n1843 ), .A2(_u10_u8_n2545 ), .ZN(_u10_u8_n2702 ) );
NOR2_X1 _u10_u8_U533  ( .A1(_u10_u8_n2346 ), .A2(_u10_u8_n2700 ), .ZN(_u10_u8_n2703 ) );
NOR2_X1 _u10_u8_U532  ( .A1(_u10_u8_n2000 ), .A2(_u10_u8_n1887 ), .ZN(_u10_u8_n2704 ) );
NOR4_X1 _u10_u8_U531  ( .A1(_u10_u8_n2701 ), .A2(_u10_u8_n2702 ), .A3(_u10_u8_n2703 ), .A4(_u10_u8_n2704 ), .ZN(_u10_u8_n2671 ) );
NAND2_X1 _u10_u8_U530  ( .A1(_u10_u8_n2699 ), .A2(_u10_u8_n2700 ), .ZN(_u10_u8_n2698 ) );
NAND2_X1 _u10_u8_U529  ( .A1(_u10_u8_n2063 ), .A2(_u10_u8_n2698 ), .ZN(_u10_u8_n2682 ) );
NAND2_X1 _u10_u8_U528  ( .A1(_u10_u8_n2697 ), .A2(_u10_u8_n2103 ), .ZN(_u10_u8_n2696 ) );
NAND2_X1 _u10_u8_U527  ( .A1(_u10_u8_n2695 ), .A2(_u10_u8_n2696 ), .ZN(_u10_u8_n2694 ) );
NAND2_X1 _u10_u8_U526  ( .A1(_u10_u8_n1937 ), .A2(_u10_u8_n2694 ), .ZN(_u10_u8_n2683 ) );
INV_X1 _u10_u8_U525  ( .A(_u10_u8_n2693 ), .ZN(_u10_u8_n2691 ) );
NAND3_X1 _u10_u8_U524  ( .A1(_u10_u8_n2103 ), .A2(_u10_u8_n2502 ), .A3(1'b0),.ZN(_u10_u8_n2692 ) );
NAND2_X1 _u10_u8_U523  ( .A1(_u10_u8_n2691 ), .A2(_u10_u8_n2692 ), .ZN(_u10_u8_n2690 ) );
NAND2_X1 _u10_u8_U522  ( .A1(_u10_u8_n2236 ), .A2(_u10_u8_n2690 ), .ZN(_u10_u8_n2684 ) );
NAND3_X1 _u10_u8_U521  ( .A1(_u10_u8_n2688 ), .A2(_u10_u8_n1913 ), .A3(_u10_u8_n2689 ), .ZN(_u10_u8_n2335 ) );
NAND3_X1 _u10_u8_U520  ( .A1(_u10_u8_n2536 ), .A2(_u10_u8_n2103 ), .A3(1'b0),.ZN(_u10_u8_n2052 ) );
NOR2_X1 _u10_u8_U519  ( .A1(_u10_u8_n2052 ), .A2(_u10_u8_n2687 ), .ZN(_u10_u8_n1851 ) );
NAND2_X1 _u10_u8_U518  ( .A1(_u10_u8_n1851 ), .A2(_u10_u8_n2078 ), .ZN(_u10_u8_n2582 ) );
NOR2_X1 _u10_u8_U517  ( .A1(_u10_u8_n2686 ), .A2(_u10_u8_n2582 ), .ZN(_u10_u8_n2094 ) );
NAND3_X1 _u10_u8_U516  ( .A1(_u10_u8_n2251 ), .A2(_u10_u8_n2335 ), .A3(_u10_u8_n2094 ), .ZN(_u10_u8_n2685 ) );
NAND4_X1 _u10_u8_U515  ( .A1(_u10_u8_n2682 ), .A2(_u10_u8_n2683 ), .A3(_u10_u8_n2684 ), .A4(_u10_u8_n2685 ), .ZN(_u10_u8_n2673 ) );
INV_X1 _u10_u8_U514  ( .A(_u10_u8_n2291 ), .ZN(_u10_u8_n2057 ) );
AND2_X1 _u10_u8_U513  ( .A1(_u10_u8_n1851 ), .A2(_u10_u8_n2057 ), .ZN(_u10_u8_n2674 ) );
INV_X1 _u10_u8_U512  ( .A(_u10_u8_n1874 ), .ZN(_u10_u8_n2681 ) );
NOR2_X1 _u10_u8_U511  ( .A1(_u10_u8_n2007 ), .A2(_u10_u8_n1911 ), .ZN(_u10_u8_n2486 ) );
NOR2_X1 _u10_u8_U510  ( .A1(_u10_u8_n2681 ), .A2(_u10_u8_n2486 ), .ZN(_u10_u8_n2675 ) );
NOR2_X1 _u10_u8_U509  ( .A1(_u10_u8_n1977 ), .A2(_u10_u8_n2680 ), .ZN(_u10_u8_n2679 ) );
NOR2_X1 _u10_u8_U508  ( .A1(_u10_u8_n2679 ), .A2(_u10_u8_n2030 ), .ZN(_u10_u8_n2678 ) );
NOR2_X1 _u10_u8_U507  ( .A1(_u10_u8_n2678 ), .A2(_u10_u8_n2094 ), .ZN(_u10_u8_n2677 ) );
NOR2_X1 _u10_u8_U506  ( .A1(_u10_u8_n2677 ), .A2(_u10_u8_n2025 ), .ZN(_u10_u8_n2676 ) );
NOR4_X1 _u10_u8_U505  ( .A1(_u10_u8_n2673 ), .A2(_u10_u8_n2674 ), .A3(_u10_u8_n2675 ), .A4(_u10_u8_n2676 ), .ZN(_u10_u8_n2672 ) );
AND2_X1 _u10_u8_U504  ( .A1(_u10_u8_n2671 ), .A2(_u10_u8_n2672 ), .ZN(_u10_u8_n1990 ) );
INV_X1 _u10_u8_U503  ( .A(_u10_u8_n2670 ), .ZN(_u10_u8_n2660 ) );
NAND4_X1 _u10_u8_U502  ( .A1(_u10_u8_n2251 ), .A2(_u10_u8_n2669 ), .A3(_u10_u8_n2162 ), .A4(_u10_u8_n2169 ), .ZN(_u10_u8_n2664 ) );
AND3_X1 _u10_u8_U501  ( .A1(_u10_u8_n1977 ), .A2(_u10_u8_n2668 ), .A3(_u10_u8_n2089 ), .ZN(_u10_u8_n2555 ) );
NAND2_X1 _u10_u8_U500  ( .A1(_u10_u8_n2555 ), .A2(_u10_u8_n2667 ), .ZN(_u10_u8_n2666 ) );
NAND3_X1 _u10_u8_U499  ( .A1(_u10_u8_n2664 ), .A2(_u10_u8_n2665 ), .A3(_u10_u8_n2666 ), .ZN(_u10_u8_n1988 ) );
INV_X1 _u10_u8_U498  ( .A(_u10_u8_n1988 ), .ZN(_u10_u8_n2661 ) );
NAND2_X1 _u10_u8_U497  ( .A1(1'b0), .A2(_u10_u8_n2043 ), .ZN(_u10_u8_n2662 ));
NAND2_X1 _u10_u8_U496  ( .A1(_u10_u8_n2169 ), .A2(1'b0), .ZN(_u10_u8_n2663 ));
NAND4_X1 _u10_u8_U495  ( .A1(_u10_u8_n2660 ), .A2(_u10_u8_n2661 ), .A3(_u10_u8_n2662 ), .A4(_u10_u8_n2663 ), .ZN(_u10_u8_n2650 ) );
NAND2_X1 _u10_u8_U494  ( .A1(_u10_u8_n2659 ), .A2(1'b0), .ZN(_u10_u8_n2193 ));
INV_X1 _u10_u8_U493  ( .A(_u10_u8_n2193 ), .ZN(_u10_u8_n2143 ) );
NAND2_X1 _u10_u8_U492  ( .A1(_u10_u8_n2143 ), .A2(_u10_u8_n2036 ), .ZN(_u10_u8_n2286 ) );
INV_X1 _u10_u8_U491  ( .A(_u10_u8_n2286 ), .ZN(_u10_u8_n2577 ) );
NAND2_X1 _u10_u8_U490  ( .A1(_u10_u8_n2577 ), .A2(_u10_u8_n2278 ), .ZN(_u10_u8_n2474 ) );
INV_X1 _u10_u8_U489  ( .A(_u10_u8_n2474 ), .ZN(_u10_u8_n2306 ) );
NAND2_X1 _u10_u8_U488  ( .A1(_u10_u8_n2306 ), .A2(_u10_u8_n2251 ), .ZN(_u10_u8_n2654 ) );
NAND2_X1 _u10_u8_U487  ( .A1(_u10_u8_n2649 ), .A2(_u10_u8_n2658 ), .ZN(_u10_u8_n2655 ) );
NAND2_X1 _u10_u8_U486  ( .A1(_u10_u8_n2657 ), .A2(_u10_u8_n2445 ), .ZN(_u10_u8_n2656 ) );
NAND3_X1 _u10_u8_U485  ( .A1(_u10_u8_n2654 ), .A2(_u10_u8_n2655 ), .A3(_u10_u8_n2656 ), .ZN(_u10_u8_n2651 ) );
NOR2_X1 _u10_u8_U484  ( .A1(_u10_u8_n2366 ), .A2(_u10_u8_n2376 ), .ZN(_u10_u8_n2652 ) );
AND2_X1 _u10_u8_U483  ( .A1(_u10_u8_n1966 ), .A2(_u10_u8_n2528 ), .ZN(_u10_u8_n2653 ) );
NOR4_X1 _u10_u8_U482  ( .A1(_u10_u8_n2650 ), .A2(_u10_u8_n2651 ), .A3(_u10_u8_n2652 ), .A4(_u10_u8_n2653 ), .ZN(_u10_u8_n2613 ) );
NAND2_X1 _u10_u8_U481  ( .A1(_u10_u8_n1891 ), .A2(1'b0), .ZN(_u10_u8_n2636 ));
NAND2_X1 _u10_u8_U480  ( .A1(_u10_u8_n1868 ), .A2(_u10_u8_n2113 ), .ZN(_u10_u8_n2101 ) );
NOR4_X1 _u10_u8_U479  ( .A1(_u10_u8_n2649 ), .A2(_u10_u8_n2216 ), .A3(_u10_u8_n2101 ), .A4(_u10_u8_n2634 ), .ZN(_u10_u8_n2648 ) );
NOR2_X1 _u10_u8_U478  ( .A1(_u10_u8_n2648 ), .A2(_u10_u8_n2254 ), .ZN(_u10_u8_n2638 ) );
NOR2_X1 _u10_u8_U477  ( .A1(_u10_u8_n2106 ), .A2(_u10_u8_n2643 ), .ZN(_u10_u8_n2645 ) );
NAND2_X1 _u10_u8_U476  ( .A1(1'b0), .A2(_u10_u8_n2049 ), .ZN(_u10_u8_n2647 ));
NAND2_X1 _u10_u8_U475  ( .A1(_u10_u8_n2646 ), .A2(_u10_u8_n2647 ), .ZN(_u10_u8_n2348 ) );
NOR2_X1 _u10_u8_U474  ( .A1(_u10_u8_n2645 ), .A2(_u10_u8_n2348 ), .ZN(_u10_u8_n2644 ) );
NOR2_X1 _u10_u8_U473  ( .A1(_u10_u8_n2644 ), .A2(_u10_u8_n2495 ), .ZN(_u10_u8_n2639 ) );
NOR2_X1 _u10_u8_U472  ( .A1(_u10_u8_n2643 ), .A2(_u10_u8_n2203 ), .ZN(_u10_u8_n2642 ) );
NOR3_X1 _u10_u8_U471  ( .A1(_u10_u8_n2101 ), .A2(1'b0), .A3(_u10_u8_n2642 ),.ZN(_u10_u8_n2641 ) );
NOR2_X1 _u10_u8_U470  ( .A1(_u10_u8_n2641 ), .A2(_u10_u8_n2253 ), .ZN(_u10_u8_n2640 ) );
NOR3_X1 _u10_u8_U469  ( .A1(_u10_u8_n2638 ), .A2(_u10_u8_n2639 ), .A3(_u10_u8_n2640 ), .ZN(_u10_u8_n2637 ) );
NAND3_X1 _u10_u8_U468  ( .A1(_u10_u8_n2635 ), .A2(_u10_u8_n2636 ), .A3(_u10_u8_n2637 ), .ZN(_u10_u8_n2615 ) );
NOR3_X1 _u10_u8_U467  ( .A1(_u10_u8_n2174 ), .A2(_u10_u8_n2175 ), .A3(_u10_u8_n2179 ), .ZN(_u10_u8_n2631 ) );
NAND3_X1 _u10_u8_U466  ( .A1(_u10_u8_n2223 ), .A2(_u10_u8_n2236 ), .A3(_u10_u8_n2631 ), .ZN(_u10_u8_n2622 ) );
OR2_X1 _u10_u8_U465  ( .A1(_u10_u8_n1960 ), .A2(_u10_u8_n1959 ), .ZN(_u10_u8_n2625 ) );
NOR3_X1 _u10_u8_U464  ( .A1(_u10_u8_n2101 ), .A2(_u10_u8_n2633 ), .A3(_u10_u8_n2634 ), .ZN(_u10_u8_n2523 ) );
OR2_X1 _u10_u8_U463  ( .A1(_u10_u8_n2632 ), .A2(_u10_u8_n2523 ), .ZN(_u10_u8_n2627 ) );
INV_X1 _u10_u8_U462  ( .A(_u10_u8_n2631 ), .ZN(_u10_u8_n2628 ) );
NAND2_X1 _u10_u8_U461  ( .A1(_u10_u8_n2630 ), .A2(_u10_u8_n1922 ), .ZN(_u10_u8_n2629 ) );
NAND3_X1 _u10_u8_U460  ( .A1(_u10_u8_n2627 ), .A2(_u10_u8_n2628 ), .A3(_u10_u8_n2629 ), .ZN(_u10_u8_n2626 ) );
NAND2_X1 _u10_u8_U459  ( .A1(_u10_u8_n2625 ), .A2(_u10_u8_n2626 ), .ZN(_u10_u8_n2624 ) );
NAND3_X1 _u10_u8_U458  ( .A1(_u10_u8_n2622 ), .A2(_u10_u8_n2623 ), .A3(_u10_u8_n2624 ), .ZN(_u10_u8_n2616 ) );
AND2_X1 _u10_u8_U457  ( .A1(_u10_u8_n2621 ), .A2(_u10_u8_n2358 ), .ZN(_u10_u8_n2620 ) );
NOR2_X1 _u10_u8_U456  ( .A1(_u10_u8_n2523 ), .A2(_u10_u8_n2620 ), .ZN(_u10_u8_n2617 ) );
INV_X1 _u10_u8_U455  ( .A(_u10_u8_n2101 ), .ZN(_u10_u8_n2221 ) );
NOR2_X1 _u10_u8_U454  ( .A1(_u10_u8_n1911 ), .A2(_u10_u8_n2488 ), .ZN(_u10_u8_n2619 ) );
NOR2_X1 _u10_u8_U453  ( .A1(_u10_u8_n2221 ), .A2(_u10_u8_n2619 ), .ZN(_u10_u8_n2618 ) );
NOR4_X1 _u10_u8_U452  ( .A1(_u10_u8_n2615 ), .A2(_u10_u8_n2616 ), .A3(_u10_u8_n2617 ), .A4(_u10_u8_n2618 ), .ZN(_u10_u8_n2614 ) );
AND2_X1 _u10_u8_U451  ( .A1(_u10_u8_n2613 ), .A2(_u10_u8_n2614 ), .ZN(_u10_u8_n2314 ) );
NAND3_X1 _u10_u8_U450  ( .A1(_u10_u8_n2612 ), .A2(_u10_u8_n1990 ), .A3(_u10_u8_n2314 ), .ZN(_u10_u8_n2609 ) );
NOR4_X1 _u10_u8_U449  ( .A1(_u10_u8_n2608 ), .A2(_u10_u8_n2609 ), .A3(_u10_u8_n2610 ), .A4(_u10_u8_n2611 ), .ZN(_u10_u8_n2388 ) );
NAND2_X1 _u10_u8_U448  ( .A1(_u10_u8_n2346 ), .A2(_u10_u8_n2607 ), .ZN(_u10_u8_n2191 ) );
NAND2_X1 _u10_u8_U447  ( .A1(_u10_u8_n2143 ), .A2(_u10_u8_n2191 ), .ZN(_u10_u8_n2556 ) );
INV_X1 _u10_u8_U446  ( .A(_u10_u8_n2348 ), .ZN(_u10_u8_n2603 ) );
NAND3_X1 _u10_u8_U445  ( .A1(_u10_u8_n2535 ), .A2(_u10_u8_n2485 ), .A3(_u10_u8_n2456 ), .ZN(_u10_u8_n2606 ) );
NAND2_X1 _u10_u8_U444  ( .A1(_u10_u8_n2049 ), .A2(_u10_u8_n2606 ), .ZN(_u10_u8_n2604 ) );
NAND3_X1 _u10_u8_U443  ( .A1(_u10_u8_n2603 ), .A2(_u10_u8_n2604 ), .A3(_u10_u8_n2605 ), .ZN(_u10_u8_n2602 ) );
NAND2_X1 _u10_u8_U442  ( .A1(_u10_u8_n2043 ), .A2(_u10_u8_n2602 ), .ZN(_u10_u8_n2557 ) );
INV_X1 _u10_u8_U441  ( .A(_u10_u8_n2601 ), .ZN(_u10_u8_n2590 ) );
NAND2_X1 _u10_u8_U440  ( .A1(_u10_u8_n2599 ), .A2(_u10_u8_n2600 ), .ZN(_u10_u8_n2597 ) );
NAND2_X1 _u10_u8_U439  ( .A1(_u10_u8_n2082 ), .A2(_u10_u8_n2101 ), .ZN(_u10_u8_n2598 ) );
AND2_X1 _u10_u8_U438  ( .A1(_u10_u8_n2597 ), .A2(_u10_u8_n2598 ), .ZN(_u10_u8_n2281 ) );
NAND3_X1 _u10_u8_U437  ( .A1(_u10_u8_n1969 ), .A2(_u10_u8_n2582 ), .A3(_u10_u8_n2281 ), .ZN(_u10_u8_n2073 ) );
INV_X1 _u10_u8_U436  ( .A(_u10_u8_n2073 ), .ZN(_u10_u8_n2591 ) );
NOR2_X1 _u10_u8_U435  ( .A1(_u10_u8_n1816 ), .A2(_u10_u8_n2077 ), .ZN(_u10_u8_n2595 ) );
NOR2_X1 _u10_u8_U434  ( .A1(_u10_u8_n2595 ), .A2(_u10_u8_n2596 ), .ZN(_u10_u8_n2592 ) );
NAND3_X1 _u10_u8_U433  ( .A1(_u10_u8_n2107 ), .A2(_u10_u8_n2536 ), .A3(1'b0),.ZN(_u10_u8_n2438 ) );
INV_X1 _u10_u8_U432  ( .A(_u10_u8_n2438 ), .ZN(_u10_u8_n2427 ) );
NOR4_X1 _u10_u8_U431  ( .A1(1'b0), .A2(_u10_u8_n2594 ), .A3(_u10_u8_n2577 ),.A4(_u10_u8_n2427 ), .ZN(_u10_u8_n2593 ) );
NAND4_X1 _u10_u8_U430  ( .A1(_u10_u8_n2590 ), .A2(_u10_u8_n2591 ), .A3(_u10_u8_n2592 ), .A4(_u10_u8_n2593 ), .ZN(_u10_u8_n2589 ) );
NAND2_X1 _u10_u8_U429  ( .A1(_u10_u8_n2279 ), .A2(_u10_u8_n2589 ), .ZN(_u10_u8_n2558 ) );
NAND3_X1 _u10_u8_U428  ( .A1(_u10_u8_n2587 ), .A2(_u10_u8_n2115 ), .A3(_u10_u8_n2588 ), .ZN(_u10_u8_n2585 ) );
NOR4_X1 _u10_u8_U427  ( .A1(_u10_u8_n2585 ), .A2(_u10_u8_n2586 ), .A3(1'b0),.A4(_u10_u8_n2114 ), .ZN(_u10_u8_n2583 ) );
NOR2_X1 _u10_u8_U426  ( .A1(_u10_u8_n2583 ), .A2(_u10_u8_n2584 ), .ZN(_u10_u8_n2560 ) );
OR2_X1 _u10_u8_U425  ( .A1(_u10_u8_n2582 ), .A2(1'b0), .ZN(_u10_u8_n2581 ));
NAND2_X1 _u10_u8_U424  ( .A1(_u10_u8_n2580 ), .A2(_u10_u8_n2581 ), .ZN(_u10_u8_n1974 ) );
INV_X1 _u10_u8_U423  ( .A(_u10_u8_n1974 ), .ZN(_u10_u8_n1901 ) );
AND4_X1 _u10_u8_U422  ( .A1(_u10_u8_n1901 ), .A2(_u10_u8_n2385 ), .A3(_u10_u8_n2578 ), .A4(_u10_u8_n2579 ), .ZN(_u10_u8_n2424 ) );
NOR2_X1 _u10_u8_U421  ( .A1(1'b0), .A2(_u10_u8_n2424 ), .ZN(_u10_u8_n2574 ));
NOR3_X1 _u10_u8_U420  ( .A1(_u10_u8_n2427 ), .A2(1'b0), .A3(_u10_u8_n2577 ),.ZN(_u10_u8_n2576 ) );
NOR2_X1 _u10_u8_U419  ( .A1(_u10_u8_n2576 ), .A2(_u10_u8_n1976 ), .ZN(_u10_u8_n2575 ) );
NOR3_X1 _u10_u8_U418  ( .A1(_u10_u8_n2574 ), .A2(_u10_u8_n1979 ), .A3(_u10_u8_n2575 ), .ZN(_u10_u8_n2572 ) );
NOR2_X1 _u10_u8_U417  ( .A1(_u10_u8_n2572 ), .A2(_u10_u8_n2573 ), .ZN(_u10_u8_n2561 ) );
INV_X1 _u10_u8_U416  ( .A(_u10_u8_n2061 ), .ZN(_u10_u8_n2453 ) );
NOR2_X1 _u10_u8_U415  ( .A1(_u10_u8_n2453 ), .A2(_u10_u8_n1851 ), .ZN(_u10_u8_n2018 ) );
NAND2_X1 _u10_u8_U414  ( .A1(1'b0), .A2(_u10_u8_n2571 ), .ZN(_u10_u8_n2570 ));
NAND2_X1 _u10_u8_U413  ( .A1(_u10_u8_n2018 ), .A2(_u10_u8_n2570 ), .ZN(_u10_u8_n1837 ) );
INV_X1 _u10_u8_U412  ( .A(_u10_u8_n1837 ), .ZN(_u10_u8_n2568 ) );
NAND2_X1 _u10_u8_U411  ( .A1(1'b0), .A2(_u10_u8_n2536 ), .ZN(_u10_u8_n2569 ));
NAND2_X1 _u10_u8_U410  ( .A1(_u10_u8_n2568 ), .A2(_u10_u8_n2569 ), .ZN(_u10_u8_n2564 ) );
NOR2_X1 _u10_u8_U409  ( .A1(_u10_u8_n1841 ), .A2(_u10_u8_n1868 ), .ZN(_u10_u8_n2565 ) );
INV_X1 _u10_u8_U408  ( .A(_u10_u8_n2567 ), .ZN(_u10_u8_n2566 ) );
NOR4_X1 _u10_u8_U407  ( .A1(_u10_u8_n2564 ), .A2(_u10_u8_n2565 ), .A3(_u10_u8_n2143 ), .A4(_u10_u8_n2566 ), .ZN(_u10_u8_n2563 ) );
NOR2_X1 _u10_u8_U406  ( .A1(_u10_u8_n2563 ), .A2(_u10_u8_n2014 ), .ZN(_u10_u8_n2562 ) );
NOR3_X1 _u10_u8_U405  ( .A1(_u10_u8_n2560 ), .A2(_u10_u8_n2561 ), .A3(_u10_u8_n2562 ), .ZN(_u10_u8_n2559 ) );
NAND4_X1 _u10_u8_U404  ( .A1(_u10_u8_n2556 ), .A2(_u10_u8_n2557 ), .A3(_u10_u8_n2558 ), .A4(_u10_u8_n2559 ), .ZN(_u10_u8_n2511 ) );
INV_X1 _u10_u8_U403  ( .A(_u10_u8_n2085 ), .ZN(_u10_u8_n2293 ) );
NOR2_X1 _u10_u8_U402  ( .A1(_u10_u8_n2554 ), .A2(_u10_u8_n2555 ), .ZN(_u10_u8_n2444 ) );
NAND2_X1 _u10_u8_U401  ( .A1(_u10_u8_n2553 ), .A2(_u10_u8_n2549 ), .ZN(_u10_u8_n2552 ) );
AND2_X1 _u10_u8_U400  ( .A1(_u10_u8_n2444 ), .A2(_u10_u8_n2552 ), .ZN(_u10_u8_n2295 ) );
NAND2_X1 _u10_u8_U399  ( .A1(_u10_u8_n2551 ), .A2(_u10_u8_n2549 ), .ZN(_u10_u8_n2538 ) );
AND2_X1 _u10_u8_U398  ( .A1(_u10_u8_n2427 ), .A2(_u10_u8_n2108 ), .ZN(_u10_u8_n2460 ) );
NOR4_X1 _u10_u8_U397  ( .A1(_u10_u8_n2460 ), .A2(_u10_u8_n2306 ), .A3(_u10_u8_n2094 ), .A4(_u10_u8_n2550 ), .ZN(_u10_u8_n2409 ) );
INV_X1 _u10_u8_U396  ( .A(_u10_u8_n2409 ), .ZN(_u10_u8_n2407 ) );
NAND2_X1 _u10_u8_U395  ( .A1(_u10_u8_n2549 ), .A2(_u10_u8_n2407 ), .ZN(_u10_u8_n2546 ) );
NAND3_X1 _u10_u8_U394  ( .A1(_u10_u8_n2546 ), .A2(_u10_u8_n2547 ), .A3(_u10_u8_n2548 ), .ZN(_u10_u8_n2501 ) );
INV_X1 _u10_u8_U393  ( .A(_u10_u8_n2501 ), .ZN(_u10_u8_n2539 ) );
NOR2_X1 _u10_u8_U392  ( .A1(1'b0), .A2(_u10_u8_n2545 ), .ZN(_u10_u8_n2541 ));
AND2_X1 _u10_u8_U391  ( .A1(_u10_u8_n2544 ), .A2(_u10_u8_n2089 ), .ZN(_u10_u8_n2543 ) );
NOR3_X1 _u10_u8_U390  ( .A1(_u10_u8_n2541 ), .A2(_u10_u8_n2542 ), .A3(_u10_u8_n2543 ), .ZN(_u10_u8_n2540 ) );
NAND4_X1 _u10_u8_U389  ( .A1(_u10_u8_n2295 ), .A2(_u10_u8_n2538 ), .A3(_u10_u8_n2539 ), .A4(_u10_u8_n2540 ), .ZN(_u10_u8_n2537 ) );
NAND2_X1 _u10_u8_U388  ( .A1(_u10_u8_n2293 ), .A2(_u10_u8_n2537 ), .ZN(_u10_u8_n2515 ) );
NAND2_X1 _u10_u8_U387  ( .A1(_u10_u8_n2536 ), .A2(_u10_u8_n2508 ), .ZN(_u10_u8_n2526 ) );
NAND2_X1 _u10_u8_U386  ( .A1(_u10_u8_n2535 ), .A2(_u10_u8_n1940 ), .ZN(_u10_u8_n2532 ) );
NOR4_X1 _u10_u8_U385  ( .A1(_u10_u8_n2532 ), .A2(_u10_u8_n2533 ), .A3(1'b0),.A4(_u10_u8_n2534 ), .ZN(_u10_u8_n2530 ) );
NOR2_X1 _u10_u8_U384  ( .A1(_u10_u8_n2530 ), .A2(_u10_u8_n2531 ), .ZN(_u10_u8_n2529 ) );
NOR4_X1 _u10_u8_U383  ( .A1(_u10_u8_n2528 ), .A2(_u10_u8_n2143 ), .A3(_u10_u8_n2189 ), .A4(_u10_u8_n2529 ), .ZN(_u10_u8_n2527 ) );
NAND4_X1 _u10_u8_U382  ( .A1(_u10_u8_n2019 ), .A2(_u10_u8_n2526 ), .A3(_u10_u8_n2018 ), .A4(_u10_u8_n2527 ), .ZN(_u10_u8_n2525 ) );
NAND2_X1 _u10_u8_U381  ( .A1(_u10_u8_n2183 ), .A2(_u10_u8_n2525 ), .ZN(_u10_u8_n2516 ) );
INV_X1 _u10_u8_U380  ( .A(_u10_u8_n2524 ), .ZN(_u10_u8_n2396 ) );
NAND2_X1 _u10_u8_U379  ( .A1(_u10_u8_n2396 ), .A2(_u10_u8_n2523 ), .ZN(_u10_u8_n2522 ) );
NAND2_X1 _u10_u8_U378  ( .A1(_u10_u8_n1866 ), .A2(_u10_u8_n2522 ), .ZN(_u10_u8_n2519 ) );
AND2_X1 _u10_u8_U377  ( .A1(_u10_u8_n2493 ), .A2(_u10_u8_n1961 ), .ZN(_u10_u8_n2429 ) );
NAND2_X1 _u10_u8_U376  ( .A1(_u10_u8_n2429 ), .A2(_u10_u8_n2175 ), .ZN(_u10_u8_n2510 ) );
NAND2_X1 _u10_u8_U375  ( .A1(_u10_u8_n2510 ), .A2(_u10_u8_n1864 ), .ZN(_u10_u8_n2521 ) );
NAND3_X1 _u10_u8_U374  ( .A1(_u10_u8_n2519 ), .A2(_u10_u8_n2520 ), .A3(_u10_u8_n2521 ), .ZN(_u10_u8_n2518 ) );
NAND2_X1 _u10_u8_U373  ( .A1(_u10_u8_n1861 ), .A2(_u10_u8_n2518 ), .ZN(_u10_u8_n2517 ) );
NAND3_X1 _u10_u8_U372  ( .A1(_u10_u8_n2515 ), .A2(_u10_u8_n2516 ), .A3(_u10_u8_n2517 ), .ZN(_u10_u8_n2512 ) );
NOR2_X1 _u10_u8_U371  ( .A1(_u10_u8_n1913 ), .A2(_u10_u8_n1940 ), .ZN(_u10_u8_n2513 ) );
NOR2_X1 _u10_u8_U370  ( .A1(_u10_u8_n2113 ), .A2(_u10_u8_n2350 ), .ZN(_u10_u8_n2514 ) );
NOR4_X1 _u10_u8_U369  ( .A1(_u10_u8_n2511 ), .A2(_u10_u8_n2512 ), .A3(_u10_u8_n2513 ), .A4(_u10_u8_n2514 ), .ZN(_u10_u8_n2389 ) );
NAND2_X1 _u10_u8_U368  ( .A1(_u10_u8_n2509 ), .A2(_u10_u8_n2510 ), .ZN(_u10_u8_n2477 ) );
NAND2_X1 _u10_u8_U367  ( .A1(_u10_u8_n2507 ), .A2(_u10_u8_n2508 ), .ZN(_u10_u8_n2504 ) );
NAND2_X1 _u10_u8_U366  ( .A1(1'b0), .A2(_u10_u8_n2506 ), .ZN(_u10_u8_n2505 ));
NAND2_X1 _u10_u8_U365  ( .A1(_u10_u8_n2504 ), .A2(_u10_u8_n2505 ), .ZN(_u10_u8_n2503 ) );
NAND2_X1 _u10_u8_U364  ( .A1(_u10_u8_n2502 ), .A2(_u10_u8_n2503 ), .ZN(_u10_u8_n2478 ) );
NAND2_X1 _u10_u8_U363  ( .A1(_u10_u8_n2501 ), .A2(_u10_u8_n2446 ), .ZN(_u10_u8_n2497 ) );
INV_X1 _u10_u8_U362  ( .A(_u10_u8_n2500 ), .ZN(_u10_u8_n2499 ) );
NAND3_X1 _u10_u8_U361  ( .A1(_u10_u8_n2497 ), .A2(_u10_u8_n2498 ), .A3(_u10_u8_n2499 ), .ZN(_u10_u8_n2496 ) );
NAND2_X1 _u10_u8_U360  ( .A1(_u10_u8_n2445 ), .A2(_u10_u8_n2496 ), .ZN(_u10_u8_n2479 ) );
NOR2_X1 _u10_u8_U359  ( .A1(_u10_u8_n2429 ), .A2(_u10_u8_n2495 ), .ZN(_u10_u8_n2491 ) );
INV_X1 _u10_u8_U358  ( .A(_u10_u8_n2191 ), .ZN(_u10_u8_n2494 ) );
NOR2_X1 _u10_u8_U357  ( .A1(_u10_u8_n2493 ), .A2(_u10_u8_n2494 ), .ZN(_u10_u8_n2492 ) );
NOR2_X1 _u10_u8_U356  ( .A1(_u10_u8_n2491 ), .A2(_u10_u8_n2492 ), .ZN(_u10_u8_n2489 ) );
NOR2_X1 _u10_u8_U355  ( .A1(_u10_u8_n2489 ), .A2(_u10_u8_n2490 ), .ZN(_u10_u8_n2481 ) );
NAND2_X1 _u10_u8_U354  ( .A1(_u10_u8_n2253 ), .A2(_u10_u8_n1859 ), .ZN(_u10_u8_n2398 ) );
NOR2_X1 _u10_u8_U353  ( .A1(_u10_u8_n2488 ), .A2(_u10_u8_n2398 ), .ZN(_u10_u8_n2487 ) );
NOR2_X1 _u10_u8_U352  ( .A1(_u10_u8_n2220 ), .A2(_u10_u8_n2487 ), .ZN(_u10_u8_n2482 ) );
AND2_X1 _u10_u8_U351  ( .A1(_u10_u8_n2350 ), .A2(_u10_u8_n2486 ), .ZN(_u10_u8_n2484 ) );
NOR2_X1 _u10_u8_U350  ( .A1(_u10_u8_n2484 ), .A2(_u10_u8_n2485 ), .ZN(_u10_u8_n2483 ) );
NOR3_X1 _u10_u8_U349  ( .A1(_u10_u8_n2481 ), .A2(_u10_u8_n2482 ), .A3(_u10_u8_n2483 ), .ZN(_u10_u8_n2480 ) );
NAND4_X1 _u10_u8_U348  ( .A1(_u10_u8_n2477 ), .A2(_u10_u8_n2478 ), .A3(_u10_u8_n2479 ), .A4(_u10_u8_n2480 ), .ZN(_u10_u8_n2447 ) );
NAND2_X1 _u10_u8_U347  ( .A1(_u10_u8_n2476 ), .A2(_u10_u8_n1936 ), .ZN(_u10_u8_n2472 ) );
NAND2_X1 _u10_u8_U346  ( .A1(_u10_u8_n2427 ), .A2(_u10_u8_n2278 ), .ZN(_u10_u8_n2473 ) );
NAND4_X1 _u10_u8_U345  ( .A1(_u10_u8_n2472 ), .A2(_u10_u8_n2473 ), .A3(_u10_u8_n2474 ), .A4(_u10_u8_n2475 ), .ZN(_u10_u8_n2471 ) );
NAND2_X1 _u10_u8_U344  ( .A1(_u10_u8_n2470 ), .A2(_u10_u8_n2471 ), .ZN(_u10_u8_n2457 ) );
NAND2_X1 _u10_u8_U343  ( .A1(_u10_u8_n2409 ), .A2(_u10_u8_n2469 ), .ZN(_u10_u8_n2468 ) );
NAND2_X1 _u10_u8_U342  ( .A1(_u10_u8_n2467 ), .A2(_u10_u8_n2468 ), .ZN(_u10_u8_n2463 ) );
NAND2_X1 _u10_u8_U341  ( .A1(_u10_u8_n1844 ), .A2(_u10_u8_n2466 ), .ZN(_u10_u8_n2465 ) );
NAND3_X1 _u10_u8_U340  ( .A1(_u10_u8_n2463 ), .A2(_u10_u8_n2464 ), .A3(_u10_u8_n2465 ), .ZN(_u10_u8_n2462 ) );
NAND2_X1 _u10_u8_U339  ( .A1(_u10_u8_n2461 ), .A2(_u10_u8_n2462 ), .ZN(_u10_u8_n2458 ) );
NAND2_X1 _u10_u8_U338  ( .A1(_u10_u8_n2460 ), .A2(_u10_u8_n2251 ), .ZN(_u10_u8_n2459 ) );
NAND3_X1 _u10_u8_U337  ( .A1(_u10_u8_n2457 ), .A2(_u10_u8_n2458 ), .A3(_u10_u8_n2459 ), .ZN(_u10_u8_n2448 ) );
NOR2_X1 _u10_u8_U336  ( .A1(_u10_u8_n2455 ), .A2(_u10_u8_n2456 ), .ZN(_u10_u8_n2449 ) );
NAND2_X1 _u10_u8_U335  ( .A1(_u10_u8_n2454 ), .A2(_u10_u8_n2438 ), .ZN(_u10_u8_n2452 ) );
NOR4_X1 _u10_u8_U334  ( .A1(_u10_u8_n2452 ), .A2(_u10_u8_n2453 ), .A3(_u10_u8_n2443 ), .A4(_u10_u8_n2143 ), .ZN(_u10_u8_n2451 ) );
NOR2_X1 _u10_u8_U333  ( .A1(_u10_u8_n2451 ), .A2(_u10_u8_n2356 ), .ZN(_u10_u8_n2450 ) );
NOR4_X1 _u10_u8_U332  ( .A1(_u10_u8_n2447 ), .A2(_u10_u8_n2448 ), .A3(_u10_u8_n2449 ), .A4(_u10_u8_n2450 ), .ZN(_u10_u8_n2390 ) );
NAND2_X1 _u10_u8_U331  ( .A1(_u10_u8_n2445 ), .A2(_u10_u8_n2446 ), .ZN(_u10_u8_n2155 ) );
INV_X1 _u10_u8_U330  ( .A(_u10_u8_n2155 ), .ZN(_u10_u8_n1892 ) );
INV_X1 _u10_u8_U329  ( .A(_u10_u8_n2444 ), .ZN(_u10_u8_n2088 ) );
NAND2_X1 _u10_u8_U328  ( .A1(_u10_u8_n1892 ), .A2(_u10_u8_n2088 ), .ZN(_u10_u8_n2337 ) );
NOR3_X1 _u10_u8_U327  ( .A1(_u10_u8_n2441 ), .A2(_u10_u8_n2442 ), .A3(_u10_u8_n2443 ), .ZN(_u10_u8_n2440 ) );
NAND4_X1 _u10_u8_U326  ( .A1(_u10_u8_n2193 ), .A2(_u10_u8_n2355 ), .A3(_u10_u8_n2439 ), .A4(_u10_u8_n2440 ), .ZN(_u10_u8_n2434 ) );
NAND3_X1 _u10_u8_U325  ( .A1(_u10_u8_n2437 ), .A2(_u10_u8_n2438 ), .A3(_u10_u8_n2059 ), .ZN(_u10_u8_n2435 ) );
NOR4_X1 _u10_u8_U324  ( .A1(_u10_u8_n2434 ), .A2(_u10_u8_n2435 ), .A3(_u10_u8_n1837 ), .A4(_u10_u8_n2436 ), .ZN(_u10_u8_n2433 ) );
NOR2_X1 _u10_u8_U323  ( .A1(_u10_u8_n2433 ), .A2(_u10_u8_n1836 ), .ZN(_u10_u8_n2415 ) );
INV_X1 _u10_u8_U322  ( .A(_u10_u8_n2432 ), .ZN(_u10_u8_n2178 ) );
NOR2_X1 _u10_u8_U321  ( .A1(_u10_u8_n1960 ), .A2(_u10_u8_n2431 ), .ZN(_u10_u8_n2430 ) );
NOR4_X1 _u10_u8_U320  ( .A1(_u10_u8_n2178 ), .A2(_u10_u8_n2429 ), .A3(_u10_u8_n2430 ), .A4(_u10_u8_n2179 ), .ZN(_u10_u8_n2416 ) );
NOR2_X1 _u10_u8_U319  ( .A1(_u10_u8_n2427 ), .A2(_u10_u8_n2428 ), .ZN(_u10_u8_n2426 ) );
NAND4_X1 _u10_u8_U318  ( .A1(_u10_u8_n2286 ), .A2(_u10_u8_n1969 ), .A3(_u10_u8_n2282 ), .A4(_u10_u8_n2426 ), .ZN(_u10_u8_n2425 ) );
NAND2_X1 _u10_u8_U317  ( .A1(_u10_u8_n2031 ), .A2(_u10_u8_n2425 ), .ZN(_u10_u8_n2422 ) );
NAND3_X1 _u10_u8_U316  ( .A1(_u10_u8_n2422 ), .A2(_u10_u8_n2423 ), .A3(_u10_u8_n2424 ), .ZN(_u10_u8_n2419 ) );
NOR4_X1 _u10_u8_U315  ( .A1(_u10_u8_n2419 ), .A2(_u10_u8_n1978 ), .A3(_u10_u8_n2420 ), .A4(_u10_u8_n2421 ), .ZN(_u10_u8_n2418 ) );
NOR2_X1 _u10_u8_U314  ( .A1(_u10_u8_n2418 ), .A2(_u10_u8_n2359 ), .ZN(_u10_u8_n2417 ) );
NOR3_X1 _u10_u8_U313  ( .A1(_u10_u8_n2415 ), .A2(_u10_u8_n2416 ), .A3(_u10_u8_n2417 ), .ZN(_u10_u8_n2414 ) );
NAND4_X1 _u10_u8_U312  ( .A1(_u10_u8_n2337 ), .A2(_u10_u8_n2412 ), .A3(_u10_u8_n2413 ), .A4(_u10_u8_n2414 ), .ZN(_u10_u8_n2392 ) );
NAND2_X1 _u10_u8_U311  ( .A1(_u10_u8_n2411 ), .A2(_u10_u8_n1936 ), .ZN(_u10_u8_n2410 ) );
NAND2_X1 _u10_u8_U310  ( .A1(_u10_u8_n2409 ), .A2(_u10_u8_n2410 ), .ZN(_u10_u8_n2408 ) );
NAND3_X1 _u10_u8_U309  ( .A1(_u10_u8_n2408 ), .A2(_u10_u8_n2305 ), .A3(_u10_u8_n1894 ), .ZN(_u10_u8_n2402 ) );
NAND3_X1 _u10_u8_U308  ( .A1(_u10_u8_n2329 ), .A2(_u10_u8_n2407 ), .A3(_u10_u8_n2255 ), .ZN(_u10_u8_n2403 ) );
NAND3_X1 _u10_u8_U307  ( .A1(_u10_u8_n1924 ), .A2(_u10_u8_n2405 ), .A3(_u10_u8_n2406 ), .ZN(_u10_u8_n2404 ) );
NAND3_X1 _u10_u8_U306  ( .A1(_u10_u8_n2402 ), .A2(_u10_u8_n2403 ), .A3(_u10_u8_n2404 ), .ZN(_u10_u8_n2393 ) );
INV_X1 _u10_u8_U305  ( .A(_u10_u8_n1932 ), .ZN(_u10_u8_n2399 ) );
NOR2_X1 _u10_u8_U304  ( .A1(_u10_u8_n2401 ), .A2(_u10_u8_n2161 ), .ZN(_u10_u8_n2400 ) );
NOR2_X1 _u10_u8_U303  ( .A1(_u10_u8_n2399 ), .A2(_u10_u8_n2400 ), .ZN(_u10_u8_n2394 ) );
NOR2_X1 _u10_u8_U302  ( .A1(_u10_u8_n2110 ), .A2(_u10_u8_n2398 ), .ZN(_u10_u8_n2397 ) );
NOR2_X1 _u10_u8_U301  ( .A1(_u10_u8_n2396 ), .A2(_u10_u8_n2397 ), .ZN(_u10_u8_n2395 ) );
NOR4_X1 _u10_u8_U300  ( .A1(_u10_u8_n2392 ), .A2(_u10_u8_n2393 ), .A3(_u10_u8_n2394 ), .A4(_u10_u8_n2395 ), .ZN(_u10_u8_n2391 ) );
NAND4_X1 _u10_u8_U299  ( .A1(_u10_u8_n2388 ), .A2(_u10_u8_n2389 ), .A3(_u10_u8_n2390 ), .A4(_u10_u8_n2391 ), .ZN(_u10_u8_n2387 ) );
MUX2_X1 _u10_u8_U298  ( .A(_u10_u8_n2387 ), .B(_u10_SYNOPSYS_UNCONNECTED_35 ), .S(_u10_u8_n1819 ), .Z(_u10_u8_n1810 ) );
NAND2_X1 _u10_u8_U297  ( .A1(_u10_u8_n2386 ), .A2(_u10_u8_n2007 ), .ZN(_u10_u8_n2369 ) );
AND2_X1 _u10_u8_U296  ( .A1(1'b0), .A2(_u10_u8_n2195 ), .ZN(_u10_u8_n2308 ));
NAND2_X1 _u10_u8_U295  ( .A1(_u10_u8_n2308 ), .A2(_u10_u8_n2036 ), .ZN(_u10_u8_n2384 ) );
AND2_X1 _u10_u8_U294  ( .A1(_u10_u8_n2384 ), .A2(_u10_u8_n2385 ), .ZN(_u10_u8_n2275 ) );
AND4_X1 _u10_u8_U293  ( .A1(_u10_u8_n2275 ), .A2(_u10_u8_n2286 ), .A3(_u10_u8_n2383 ), .A4(_u10_u8_n2285 ), .ZN(_u10_u8_n2225 ) );
NAND3_X1 _u10_u8_U292  ( .A1(_u10_u8_n2195 ), .A2(_u10_u8_n2223 ), .A3(1'b0),.ZN(_u10_u8_n2021 ) );
INV_X1 _u10_u8_U291  ( .A(_u10_u8_n2021 ), .ZN(_u10_u8_n2167 ) );
NAND2_X1 _u10_u8_U290  ( .A1(_u10_u8_n2036 ), .A2(_u10_u8_n2167 ), .ZN(_u10_u8_n1970 ) );
AND3_X1 _u10_u8_U289  ( .A1(_u10_u8_n1970 ), .A2(_u10_u8_n2164 ), .A3(_u10_u8_n2382 ), .ZN(_u10_u8_n2381 ) );
NAND4_X1 _u10_u8_U288  ( .A1(_u10_u8_n2225 ), .A2(_u10_u8_n2379 ), .A3(_u10_u8_n2380 ), .A4(_u10_u8_n2381 ), .ZN(_u10_u8_n2378 ) );
NAND2_X1 _u10_u8_U287  ( .A1(_u10_u8_n1967 ), .A2(_u10_u8_n2378 ), .ZN(_u10_u8_n2370 ) );
NAND2_X1 _u10_u8_U286  ( .A1(_u10_u8_n2081 ), .A2(_u10_u8_n2377 ), .ZN(_u10_u8_n2371 ) );
NOR2_X1 _u10_u8_U285  ( .A1(_u10_u8_n2375 ), .A2(_u10_u8_n2376 ), .ZN(_u10_u8_n2373 ) );
NOR2_X1 _u10_u8_U284  ( .A1(_u10_u8_n2373 ), .A2(_u10_u8_n2374 ), .ZN(_u10_u8_n2372 ) );
NAND4_X1 _u10_u8_U283  ( .A1(_u10_u8_n2369 ), .A2(_u10_u8_n2370 ), .A3(_u10_u8_n2371 ), .A4(_u10_u8_n2372 ), .ZN(_u10_u8_n2309 ) );
NOR2_X1 _u10_u8_U282  ( .A1(_u10_u8_n2000 ), .A2(_u10_u8_n2368 ), .ZN(_u10_u8_n2360 ) );
NOR2_X1 _u10_u8_U281  ( .A1(_u10_u8_n2366 ), .A2(_u10_u8_n2367 ), .ZN(_u10_u8_n2361 ) );
NOR2_X1 _u10_u8_U280  ( .A1(_u10_u8_n1868 ), .A2(_u10_u8_n2365 ), .ZN(_u10_u8_n2362 ) );
NOR2_X1 _u10_u8_U279  ( .A1(_u10_u8_n2364 ), .A2(_u10_u8_n1859 ), .ZN(_u10_u8_n2363 ) );
NOR4_X1 _u10_u8_U278  ( .A1(_u10_u8_n2360 ), .A2(_u10_u8_n2361 ), .A3(_u10_u8_n2362 ), .A4(_u10_u8_n2363 ), .ZN(_u10_u8_n2316 ) );
NOR2_X1 _u10_u8_U277  ( .A1(_u10_u8_n2359 ), .A2(_u10_u8_n1970 ), .ZN(_u10_u8_n2351 ) );
NOR2_X1 _u10_u8_U276  ( .A1(_u10_u8_n2358 ), .A2(_u10_u8_n1840 ), .ZN(_u10_u8_n2352 ) );
NOR2_X1 _u10_u8_U275  ( .A1(_u10_u8_n2356 ), .A2(_u10_u8_n2357 ), .ZN(_u10_u8_n2353 ) );
NOR2_X1 _u10_u8_U274  ( .A1(_u10_u8_n1836 ), .A2(_u10_u8_n2355 ), .ZN(_u10_u8_n2354 ) );
NOR4_X1 _u10_u8_U273  ( .A1(_u10_u8_n2351 ), .A2(_u10_u8_n2352 ), .A3(_u10_u8_n2353 ), .A4(_u10_u8_n2354 ), .ZN(_u10_u8_n2317 ) );
NOR2_X1 _u10_u8_U272  ( .A1(_u10_u8_n1873 ), .A2(_u10_u8_n2101 ), .ZN(_u10_u8_n2349 ) );
NOR2_X1 _u10_u8_U271  ( .A1(_u10_u8_n2349 ), .A2(_u10_u8_n2350 ), .ZN(_u10_u8_n2338 ) );
NOR2_X1 _u10_u8_U270  ( .A1(_u10_u8_n2347 ), .A2(_u10_u8_n2348 ), .ZN(_u10_u8_n2345 ) );
NOR2_X1 _u10_u8_U269  ( .A1(_u10_u8_n2345 ), .A2(_u10_u8_n2346 ), .ZN(_u10_u8_n2339 ) );
NOR2_X1 _u10_u8_U268  ( .A1(_u10_u8_n2344 ), .A2(_u10_u8_n2142 ), .ZN(_u10_u8_n2340 ) );
NOR2_X1 _u10_u8_U267  ( .A1(_u10_u8_n2342 ), .A2(_u10_u8_n2343 ), .ZN(_u10_u8_n2341 ) );
NOR4_X1 _u10_u8_U266  ( .A1(_u10_u8_n2338 ), .A2(_u10_u8_n2339 ), .A3(_u10_u8_n2340 ), .A4(_u10_u8_n2341 ), .ZN(_u10_u8_n2318 ) );
INV_X1 _u10_u8_U265  ( .A(_u10_u8_n2337 ), .ZN(_u10_u8_n2320 ) );
NOR2_X1 _u10_u8_U264  ( .A1(_u10_u8_n1970 ), .A2(1'b0), .ZN(_u10_u8_n2027 ));
INV_X1 _u10_u8_U263  ( .A(_u10_u8_n2027 ), .ZN(_u10_u8_n2331 ) );
NOR2_X1 _u10_u8_U262  ( .A1(_u10_u8_n2174 ), .A2(_u10_u8_n2216 ), .ZN(_u10_u8_n2333 ) );
AND2_X1 _u10_u8_U261  ( .A1(_u10_u8_n1928 ), .A2(_u10_u8_n2336 ), .ZN(_u10_u8_n2334 ) );
NOR4_X1 _u10_u8_U260  ( .A1(_u10_u8_n1937 ), .A2(_u10_u8_n2333 ), .A3(_u10_u8_n2334 ), .A4(_u10_u8_n2335 ), .ZN(_u10_u8_n2332 ) );
NOR3_X1 _u10_u8_U259  ( .A1(_u10_u8_n2331 ), .A2(_u10_u8_n2332 ), .A3(_u10_u8_n1915 ), .ZN(_u10_u8_n2321 ) );
NOR3_X1 _u10_u8_U258  ( .A1(_u10_u8_n2291 ), .A2(_u10_u8_n2330 ), .A3(_u10_u8_n2021 ), .ZN(_u10_u8_n2322 ) );
NOR2_X1 _u10_u8_U257  ( .A1(_u10_u8_n2329 ), .A2(_u10_u8_n2169 ), .ZN(_u10_u8_n2324 ) );
NOR2_X1 _u10_u8_U256  ( .A1(1'b0), .A2(_u10_u8_n2328 ), .ZN(_u10_u8_n2327 ));
NOR2_X1 _u10_u8_U255  ( .A1(_u10_u8_n2326 ), .A2(_u10_u8_n2327 ), .ZN(_u10_u8_n2325 ) );
NOR3_X1 _u10_u8_U254  ( .A1(_u10_u8_n2324 ), .A2(1'b0), .A3(_u10_u8_n2325 ),.ZN(_u10_u8_n2323 ) );
NOR4_X1 _u10_u8_U253  ( .A1(_u10_u8_n2320 ), .A2(_u10_u8_n2321 ), .A3(_u10_u8_n2322 ), .A4(_u10_u8_n2323 ), .ZN(_u10_u8_n2319 ) );
AND4_X1 _u10_u8_U252  ( .A1(_u10_u8_n2316 ), .A2(_u10_u8_n2317 ), .A3(_u10_u8_n2318 ), .A4(_u10_u8_n2319 ), .ZN(_u10_u8_n1991 ) );
INV_X1 _u10_u8_U251  ( .A(_u10_u8_n2315 ), .ZN(_u10_u8_n2313 ) );
NAND3_X1 _u10_u8_U250  ( .A1(_u10_u8_n1991 ), .A2(_u10_u8_n2313 ), .A3(_u10_u8_n2314 ), .ZN(_u10_u8_n2310 ) );
NOR4_X1 _u10_u8_U249  ( .A1(_u10_u8_n2309 ), .A2(_u10_u8_n2310 ), .A3(_u10_u8_n2311 ), .A4(_u10_u8_n2312 ), .ZN(_u10_u8_n2117 ) );
NAND3_X1 _u10_u8_U248  ( .A1(_u10_u8_n2108 ), .A2(_u10_u8_n2107 ), .A3(_u10_u8_n2308 ), .ZN(_u10_u8_n2217 ) );
NOR3_X1 _u10_u8_U247  ( .A1(_u10_u8_n2306 ), .A2(_u10_u8_n2307 ), .A3(_u10_u8_n2027 ), .ZN(_u10_u8_n2277 ) );
NAND3_X1 _u10_u8_U246  ( .A1(_u10_u8_n2217 ), .A2(_u10_u8_n2305 ), .A3(_u10_u8_n2277 ), .ZN(_u10_u8_n2157 ) );
NAND2_X1 _u10_u8_U245  ( .A1(_u10_u8_n2089 ), .A2(_u10_u8_n2157 ), .ZN(_u10_u8_n2296 ) );
INV_X1 _u10_u8_U244  ( .A(_u10_u8_n2304 ), .ZN(_u10_u8_n2297 ) );
NOR2_X1 _u10_u8_U243  ( .A1(_u10_u8_n2302 ), .A2(_u10_u8_n2303 ), .ZN(_u10_u8_n2299 ) );
NOR3_X1 _u10_u8_U242  ( .A1(_u10_u8_n2299 ), .A2(_u10_u8_n2300 ), .A3(_u10_u8_n2301 ), .ZN(_u10_u8_n2298 ) );
NAND4_X1 _u10_u8_U241  ( .A1(_u10_u8_n2295 ), .A2(_u10_u8_n2296 ), .A3(_u10_u8_n2297 ), .A4(_u10_u8_n2298 ), .ZN(_u10_u8_n2294 ) );
NAND2_X1 _u10_u8_U240  ( .A1(_u10_u8_n2293 ), .A2(_u10_u8_n2294 ), .ZN(_u10_u8_n2257 ) );
NAND2_X1 _u10_u8_U239  ( .A1(_u10_u8_n2165 ), .A2(_u10_u8_n2166 ), .ZN(_u10_u8_n2288 ) );
NAND2_X1 _u10_u8_U238  ( .A1(_u10_u8_n2078 ), .A2(_u10_u8_n2279 ), .ZN(_u10_u8_n2292 ) );
NAND2_X1 _u10_u8_U237  ( .A1(_u10_u8_n2291 ), .A2(_u10_u8_n2292 ), .ZN(_u10_u8_n2290 ) );
NAND2_X1 _u10_u8_U236  ( .A1(_u10_u8_n2059 ), .A2(_u10_u8_n2290 ), .ZN(_u10_u8_n2289 ) );
NAND2_X1 _u10_u8_U235  ( .A1(_u10_u8_n2288 ), .A2(_u10_u8_n2289 ), .ZN(_u10_u8_n2201 ) );
NAND2_X1 _u10_u8_U234  ( .A1(1'b0), .A2(_u10_u8_n2201 ), .ZN(_u10_u8_n2258 ));
INV_X1 _u10_u8_U233  ( .A(_u10_u8_n2287 ), .ZN(_u10_u8_n2283 ) );
AND4_X1 _u10_u8_U232  ( .A1(_u10_u8_n2285 ), .A2(_u10_u8_n2226 ), .A3(_u10_u8_n1970 ), .A4(_u10_u8_n2286 ), .ZN(_u10_u8_n2284 ) );
NAND4_X1 _u10_u8_U231  ( .A1(_u10_u8_n2281 ), .A2(_u10_u8_n2282 ), .A3(_u10_u8_n2283 ), .A4(_u10_u8_n2284 ), .ZN(_u10_u8_n2280 ) );
NAND2_X1 _u10_u8_U230  ( .A1(_u10_u8_n2279 ), .A2(_u10_u8_n2280 ), .ZN(_u10_u8_n2259 ) );
NAND4_X1 _u10_u8_U229  ( .A1(_u10_u8_n2275 ), .A2(_u10_u8_n2276 ), .A3(_u10_u8_n2277 ), .A4(_u10_u8_n2278 ), .ZN(_u10_u8_n2271 ) );
NAND2_X1 _u10_u8_U228  ( .A1(_u10_u8_n1933 ), .A2(_u10_u8_n2164 ), .ZN(_u10_u8_n2272 ) );
NOR2_X1 _u10_u8_U227  ( .A1(_u10_u8_n2274 ), .A2(_u10_u8_n2130 ), .ZN(_u10_u8_n2273 ) );
NOR4_X1 _u10_u8_U226  ( .A1(_u10_u8_n2271 ), .A2(_u10_u8_n2272 ), .A3(_u10_u8_n1978 ), .A4(_u10_u8_n2273 ), .ZN(_u10_u8_n2270 ) );
NOR2_X1 _u10_u8_U225  ( .A1(_u10_u8_n2270 ), .A2(_u10_u8_n2025 ), .ZN(_u10_u8_n2261 ) );
NAND3_X1 _u10_u8_U224  ( .A1(_u10_u8_n1933 ), .A2(_u10_u8_n1936 ), .A3(_u10_u8_n2269 ), .ZN(_u10_u8_n2268 ) );
NOR3_X1 _u10_u8_U223  ( .A1(_u10_u8_n2268 ), .A2(_u10_u8_n1844 ), .A3(_u10_u8_n2157 ), .ZN(_u10_u8_n2267 ) );
NOR2_X1 _u10_u8_U222  ( .A1(1'b0), .A2(_u10_u8_n2267 ), .ZN(_u10_u8_n2265 ));
NOR3_X1 _u10_u8_U221  ( .A1(_u10_u8_n2264 ), .A2(_u10_u8_n2265 ), .A3(_u10_u8_n2266 ), .ZN(_u10_u8_n2263 ) );
NOR2_X1 _u10_u8_U220  ( .A1(_u10_u8_n2263 ), .A2(_u10_u8_n1843 ), .ZN(_u10_u8_n2262 ) );
NOR2_X1 _u10_u8_U219  ( .A1(_u10_u8_n2261 ), .A2(_u10_u8_n2262 ), .ZN(_u10_u8_n2260 ) );
NAND4_X1 _u10_u8_U218  ( .A1(_u10_u8_n2257 ), .A2(_u10_u8_n2258 ), .A3(_u10_u8_n2259 ), .A4(_u10_u8_n2260 ), .ZN(_u10_u8_n2230 ) );
INV_X1 _u10_u8_U217  ( .A(_u10_u8_n2217 ), .ZN(_u10_u8_n2242 ) );
NAND2_X1 _u10_u8_U216  ( .A1(_u10_u8_n2168 ), .A2(_u10_u8_n2169 ), .ZN(_u10_u8_n2244 ) );
NAND2_X1 _u10_u8_U215  ( .A1(_u10_u8_n2255 ), .A2(_u10_u8_n2256 ), .ZN(_u10_u8_n2245 ) );
NAND2_X1 _u10_u8_U214  ( .A1(_u10_u8_n2253 ), .A2(_u10_u8_n2254 ), .ZN(_u10_u8_n2252 ) );
NAND2_X1 _u10_u8_U213  ( .A1(_u10_u8_n2251 ), .A2(_u10_u8_n2252 ), .ZN(_u10_u8_n2246 ) );
NAND2_X1 _u10_u8_U212  ( .A1(_u10_u8_n2152 ), .A2(_u10_u8_n1928 ), .ZN(_u10_u8_n2250 ) );
NAND2_X1 _u10_u8_U211  ( .A1(_u10_u8_n2249 ), .A2(_u10_u8_n2250 ), .ZN(_u10_u8_n2248 ) );
NAND2_X1 _u10_u8_U210  ( .A1(_u10_u8_n2105 ), .A2(_u10_u8_n2248 ), .ZN(_u10_u8_n2247 ) );
NAND4_X1 _u10_u8_U209  ( .A1(_u10_u8_n2244 ), .A2(_u10_u8_n2245 ), .A3(_u10_u8_n2246 ), .A4(_u10_u8_n2247 ), .ZN(_u10_u8_n2243 ) );
NAND2_X1 _u10_u8_U208  ( .A1(_u10_u8_n2242 ), .A2(_u10_u8_n2243 ), .ZN(_u10_u8_n2237 ) );
NAND2_X1 _u10_u8_U207  ( .A1(1'b0), .A2(_u10_u8_n2241 ), .ZN(_u10_u8_n2238 ));
NAND2_X1 _u10_u8_U206  ( .A1(_u10_u8_n2214 ), .A2(_u10_u8_n2240 ), .ZN(_u10_u8_n2239 ) );
NAND3_X1 _u10_u8_U205  ( .A1(_u10_u8_n2237 ), .A2(_u10_u8_n2238 ), .A3(_u10_u8_n2239 ), .ZN(_u10_u8_n2231 ) );
AND2_X1 _u10_u8_U204  ( .A1(_u10_u8_n2200 ), .A2(_u10_u8_n2236 ), .ZN(_u10_u8_n2232 ) );
NOR2_X1 _u10_u8_U203  ( .A1(_u10_u8_n2234 ), .A2(_u10_u8_n2235 ), .ZN(_u10_u8_n2233 ) );
NOR4_X1 _u10_u8_U202  ( .A1(_u10_u8_n2230 ), .A2(_u10_u8_n2231 ), .A3(_u10_u8_n2232 ), .A4(_u10_u8_n2233 ), .ZN(_u10_u8_n2118 ) );
NAND2_X1 _u10_u8_U201  ( .A1(_u10_u8_n2214 ), .A2(_u10_u8_n2049 ), .ZN(_u10_u8_n2229 ) );
NAND2_X1 _u10_u8_U200  ( .A1(_u10_u8_n2228 ), .A2(_u10_u8_n2229 ), .ZN(_u10_u8_n2227 ) );
NAND2_X1 _u10_u8_U199  ( .A1(_u10_u8_n2043 ), .A2(_u10_u8_n2227 ), .ZN(_u10_u8_n2204 ) );
NAND2_X1 _u10_u8_U198  ( .A1(_u10_u8_n2225 ), .A2(_u10_u8_n2226 ), .ZN(_u10_u8_n2224 ) );
NAND2_X1 _u10_u8_U197  ( .A1(_u10_u8_n1899 ), .A2(_u10_u8_n2224 ), .ZN(_u10_u8_n2205 ) );
NAND2_X1 _u10_u8_U196  ( .A1(_u10_u8_n2222 ), .A2(_u10_u8_n2223 ), .ZN(_u10_u8_n1870 ) );
NAND4_X1 _u10_u8_U195  ( .A1(_u10_u8_n2220 ), .A2(_u10_u8_n2131 ), .A3(_u10_u8_n2221 ), .A4(_u10_u8_n1870 ), .ZN(_u10_u8_n2219 ) );
NAND2_X1 _u10_u8_U194  ( .A1(_u10_u8_n2218 ), .A2(_u10_u8_n2219 ), .ZN(_u10_u8_n2206 ) );
NOR2_X1 _u10_u8_U193  ( .A1(_u10_u8_n1925 ), .A2(_u10_u8_n2217 ), .ZN(_u10_u8_n2215 ) );
NOR4_X1 _u10_u8_U192  ( .A1(_u10_u8_n2213 ), .A2(_u10_u8_n2214 ), .A3(_u10_u8_n2215 ), .A4(_u10_u8_n2216 ), .ZN(_u10_u8_n2211 ) );
NOR2_X1 _u10_u8_U191  ( .A1(_u10_u8_n2211 ), .A2(_u10_u8_n2212 ), .ZN(_u10_u8_n2208 ) );
NOR2_X1 _u10_u8_U190  ( .A1(_u10_u8_n1888 ), .A2(_u10_u8_n2210 ), .ZN(_u10_u8_n2209 ) );
NOR2_X1 _u10_u8_U189  ( .A1(_u10_u8_n2208 ), .A2(_u10_u8_n2209 ), .ZN(_u10_u8_n2207 ) );
NAND4_X1 _u10_u8_U188  ( .A1(_u10_u8_n2204 ), .A2(_u10_u8_n2205 ), .A3(_u10_u8_n2206 ), .A4(_u10_u8_n2207 ), .ZN(_u10_u8_n2170 ) );
OR2_X1 _u10_u8_U187  ( .A1(_u10_u8_n2202 ), .A2(_u10_u8_n2203 ), .ZN(_u10_u8_n2197 ) );
NAND2_X1 _u10_u8_U186  ( .A1(1'b0), .A2(_u10_u8_n2201 ), .ZN(_u10_u8_n2198 ));
NAND2_X1 _u10_u8_U185  ( .A1(_u10_u8_n2063 ), .A2(_u10_u8_n2200 ), .ZN(_u10_u8_n2199 ) );
NAND3_X1 _u10_u8_U184  ( .A1(_u10_u8_n2197 ), .A2(_u10_u8_n2198 ), .A3(_u10_u8_n2199 ), .ZN(_u10_u8_n2196 ) );
NAND2_X1 _u10_u8_U183  ( .A1(_u10_u8_n2195 ), .A2(_u10_u8_n2196 ), .ZN(_u10_u8_n2180 ) );
NAND2_X1 _u10_u8_U182  ( .A1(_u10_u8_n2195 ), .A2(_u10_u8_n1918 ), .ZN(_u10_u8_n2192 ) );
NAND4_X1 _u10_u8_U181  ( .A1(_u10_u8_n2192 ), .A2(_u10_u8_n2021 ), .A3(_u10_u8_n2193 ), .A4(_u10_u8_n2194 ), .ZN(_u10_u8_n2188 ) );
NAND2_X1 _u10_u8_U180  ( .A1(_u10_u8_n2188 ), .A2(_u10_u8_n2191 ), .ZN(_u10_u8_n2181 ) );
NAND2_X1 _u10_u8_U179  ( .A1(1'b0), .A2(_u10_u8_n2190 ), .ZN(_u10_u8_n2185 ));
NAND2_X1 _u10_u8_U178  ( .A1(_u10_u8_n2189 ), .A2(_u10_SYNOPSYS_UNCONNECTED_36 ), .ZN(_u10_u8_n2186 ) );
INV_X1 _u10_u8_U177  ( .A(_u10_u8_n2188 ), .ZN(_u10_u8_n2187 ) );
NAND3_X1 _u10_u8_U176  ( .A1(_u10_u8_n2185 ), .A2(_u10_u8_n2186 ), .A3(_u10_u8_n2187 ), .ZN(_u10_u8_n2184 ) );
NAND2_X1 _u10_u8_U175  ( .A1(_u10_u8_n2183 ), .A2(_u10_u8_n2184 ), .ZN(_u10_u8_n2182 ) );
NAND3_X1 _u10_u8_U174  ( .A1(_u10_u8_n2180 ), .A2(_u10_u8_n2181 ), .A3(_u10_u8_n2182 ), .ZN(_u10_u8_n2171 ) );
INV_X1 _u10_u8_U173  ( .A(_u10_u8_n2179 ), .ZN(_u10_u8_n1963 ) );
NOR2_X1 _u10_u8_U172  ( .A1(_u10_u8_n1963 ), .A2(_u10_u8_n2178 ), .ZN(_u10_u8_n2172 ) );
INV_X1 _u10_u8_U171  ( .A(_u10_u8_n2177 ), .ZN(_u10_u8_n2176 ) );
NOR3_X1 _u10_u8_U170  ( .A1(_u10_u8_n2174 ), .A2(_u10_u8_n2175 ), .A3(_u10_u8_n2176 ), .ZN(_u10_u8_n2173 ) );
NOR4_X1 _u10_u8_U169  ( .A1(_u10_u8_n2170 ), .A2(_u10_u8_n2171 ), .A3(_u10_u8_n2172 ), .A4(_u10_u8_n2173 ), .ZN(_u10_u8_n2119 ) );
NAND3_X1 _u10_u8_U168  ( .A1(_u10_u8_n2168 ), .A2(_u10_u8_n2169 ), .A3(1'b0),.ZN(_u10_u8_n2148 ) );
NAND3_X1 _u10_u8_U167  ( .A1(_u10_u8_n2165 ), .A2(_u10_u8_n2166 ), .A3(_u10_u8_n2167 ), .ZN(_u10_u8_n2149 ) );
NAND4_X1 _u10_u8_U166  ( .A1(_u10_u8_n2162 ), .A2(_u10_u8_n1933 ), .A3(_u10_u8_n2163 ), .A4(_u10_u8_n2164 ), .ZN(_u10_u8_n2160 ) );
NOR4_X1 _u10_u8_U165  ( .A1(_u10_u8_n2160 ), .A2(_u10_u8_n2157 ), .A3(_u10_u8_n1844 ), .A4(_u10_u8_n2161 ), .ZN(_u10_u8_n2158 ) );
NOR2_X1 _u10_u8_U164  ( .A1(_u10_u8_n2158 ), .A2(_u10_u8_n2159 ), .ZN(_u10_u8_n2153 ) );
INV_X1 _u10_u8_U163  ( .A(_u10_u8_n2157 ), .ZN(_u10_u8_n2129 ) );
NOR3_X1 _u10_u8_U162  ( .A1(_u10_u8_n2155 ), .A2(_u10_u8_n2129 ), .A3(_u10_u8_n2156 ), .ZN(_u10_u8_n2154 ) );
NOR2_X1 _u10_u8_U161  ( .A1(_u10_u8_n2153 ), .A2(_u10_u8_n2154 ), .ZN(_u10_u8_n2150 ) );
NAND3_X1 _u10_u8_U160  ( .A1(1'b0), .A2(_u10_u8_n1928 ), .A3(_u10_u8_n2152 ),.ZN(_u10_u8_n2151 ) );
NAND4_X1 _u10_u8_U159  ( .A1(_u10_u8_n2148 ), .A2(_u10_u8_n2149 ), .A3(_u10_u8_n2150 ), .A4(_u10_u8_n2151 ), .ZN(_u10_u8_n2121 ) );
NAND2_X1 _u10_u8_U158  ( .A1(_u10_u8_n2107 ), .A2(_u10_u8_n2147 ), .ZN(_u10_u8_n2146 ) );
NAND2_X1 _u10_u8_U157  ( .A1(_u10_u8_n2145 ), .A2(_u10_u8_n2146 ), .ZN(_u10_u8_n2144 ) );
NAND2_X1 _u10_u8_U156  ( .A1(_u10_u8_n2143 ), .A2(_u10_u8_n2144 ), .ZN(_u10_u8_n2134 ) );
NAND2_X1 _u10_u8_U155  ( .A1(_u10_u8_n2141 ), .A2(_u10_u8_n2142 ), .ZN(_u10_u8_n2140 ) );
NAND2_X1 _u10_u8_U154  ( .A1(_u10_u8_n2139 ), .A2(_u10_u8_n2140 ), .ZN(_u10_u8_n2135 ) );
OR2_X1 _u10_u8_U153  ( .A1(_u10_u8_n2110 ), .A2(_u10_u8_n1911 ), .ZN(_u10_u8_n2137 ) );
NAND2_X1 _u10_u8_U152  ( .A1(_u10_u8_n2137 ), .A2(_u10_u8_n2138 ), .ZN(_u10_u8_n2136 ) );
NAND3_X1 _u10_u8_U151  ( .A1(_u10_u8_n2134 ), .A2(_u10_u8_n2135 ), .A3(_u10_u8_n2136 ), .ZN(_u10_u8_n2122 ) );
NOR2_X1 _u10_u8_U150  ( .A1(_u10_u8_n2133 ), .A2(_u10_u8_n1891 ), .ZN(_u10_u8_n2132 ) );
NOR2_X1 _u10_u8_U149  ( .A1(_u10_u8_n2131 ), .A2(_u10_u8_n2132 ), .ZN(_u10_u8_n2123 ) );
NOR2_X1 _u10_u8_U148  ( .A1(_u10_u8_n2129 ), .A2(_u10_u8_n2130 ), .ZN(_u10_u8_n2127 ) );
NOR2_X1 _u10_u8_U147  ( .A1(_u10_u8_n2127 ), .A2(_u10_u8_n2128 ), .ZN(_u10_u8_n2125 ) );
NOR2_X1 _u10_u8_U146  ( .A1(_u10_u8_n2125 ), .A2(_u10_u8_n2126 ), .ZN(_u10_u8_n2124 ) );
NOR4_X1 _u10_u8_U145  ( .A1(_u10_u8_n2121 ), .A2(_u10_u8_n2122 ), .A3(_u10_u8_n2123 ), .A4(_u10_u8_n2124 ), .ZN(_u10_u8_n2120 ) );
NAND4_X1 _u10_u8_U144  ( .A1(_u10_u8_n2117 ), .A2(_u10_u8_n2118 ), .A3(_u10_u8_n2119 ), .A4(_u10_u8_n2120 ), .ZN(_u10_u8_n2116 ) );
MUX2_X1 _u10_u8_U143  ( .A(_u10_u8_n2116 ), .B(_u10_SYNOPSYS_UNCONNECTED_36 ), .S(_u10_u8_n1819 ), .Z(_u10_u8_n1811 ) );
INV_X1 _u10_u8_U142  ( .A(_u10_u8_n2115 ), .ZN(_u10_u8_n2006 ) );
NOR3_X1 _u10_u8_U141  ( .A1(_u10_u8_n2006 ), .A2(_u10_u8_n2114 ), .A3(_u10_u8_n2081 ), .ZN(_u10_u8_n1854 ) );
NAND2_X1 _u10_u8_U140  ( .A1(_u10_u8_n2112 ), .A2(_u10_u8_n2113 ), .ZN(_u10_u8_n1872 ) );
INV_X1 _u10_u8_U139  ( .A(_u10_u8_n1872 ), .ZN(_u10_u8_n1882 ) );
NAND4_X1 _u10_u8_U138  ( .A1(_u10_u8_n1854 ), .A2(_u10_u8_n1882 ), .A3(_u10_u8_n2111 ), .A4(_u10_u8_n1868 ), .ZN(_u10_u8_n2109 ) );
NAND2_X1 _u10_u8_U137  ( .A1(_u10_u8_n2109 ), .A2(_u10_u8_n2110 ), .ZN(_u10_u8_n2098 ) );
NAND2_X1 _u10_u8_U136  ( .A1(1'b0), .A2(_u10_u8_n1983 ), .ZN(_u10_u8_n2023 ));
INV_X1 _u10_u8_U135  ( .A(_u10_u8_n2023 ), .ZN(_u10_u8_n2035 ) );
NAND3_X1 _u10_u8_U134  ( .A1(_u10_u8_n2035 ), .A2(_u10_u8_n2107 ), .A3(_u10_u8_n2108 ), .ZN(_u10_u8_n1916 ) );
INV_X1 _u10_u8_U133  ( .A(_u10_u8_n1916 ), .ZN(_u10_u8_n2093 ) );
NAND3_X1 _u10_u8_U132  ( .A1(_u10_u8_n2105 ), .A2(_u10_u8_n2106 ), .A3(_u10_u8_n2093 ), .ZN(_u10_u8_n2039 ) );
NAND2_X1 _u10_u8_U131  ( .A1(_u10_u8_n2039 ), .A2(_u10_u8_n1930 ), .ZN(_u10_u8_n2104 ) );
NAND2_X1 _u10_u8_U130  ( .A1(_u10_u8_n2103 ), .A2(_u10_u8_n2104 ), .ZN(_u10_u8_n1863 ) );
OR2_X1 _u10_u8_U129  ( .A1(_u10_u8_n1863 ), .A2(_u10_u8_n2102 ), .ZN(_u10_u8_n2099 ) );
NAND2_X1 _u10_u8_U128  ( .A1(_u10_u8_n1890 ), .A2(_u10_u8_n2101 ), .ZN(_u10_u8_n2100 ) );
NAND3_X1 _u10_u8_U127  ( .A1(_u10_u8_n2098 ), .A2(_u10_u8_n2099 ), .A3(_u10_u8_n2100 ), .ZN(_u10_u8_n2066 ) );
NAND4_X1 _u10_u8_U126  ( .A1(_u10_u8_n2095 ), .A2(_u10_u8_n2096 ), .A3(_u10_u8_n1896 ), .A4(_u10_u8_n2097 ), .ZN(_u10_u8_n2086 ) );
NOR4_X1 _u10_u8_U125  ( .A1(_u10_u8_n2093 ), .A2(_u10_u8_n2027 ), .A3(_u10_u8_n2094 ), .A4(_u10_u8_n2026 ), .ZN(_u10_u8_n1952 ) );
NOR2_X1 _u10_u8_U124  ( .A1(1'b0), .A2(_u10_u8_n1952 ), .ZN(_u10_u8_n1951 ));
INV_X1 _u10_u8_U123  ( .A(_u10_u8_n1951 ), .ZN(_u10_u8_n2090 ) );
NAND4_X1 _u10_u8_U122  ( .A1(_u10_u8_n2089 ), .A2(_u10_u8_n2090 ), .A3(_u10_u8_n2091 ), .A4(_u10_u8_n2092 ), .ZN(_u10_u8_n1893 ) );
NOR4_X1 _u10_u8_U121  ( .A1(_u10_u8_n2086 ), .A2(_u10_u8_n1893 ), .A3(_u10_u8_n2087 ), .A4(_u10_u8_n2088 ), .ZN(_u10_u8_n2084 ) );
NOR2_X1 _u10_u8_U120  ( .A1(_u10_u8_n2084 ), .A2(_u10_u8_n2085 ), .ZN(_u10_u8_n2067 ) );
NOR2_X1 _u10_u8_U119  ( .A1(_u10_u8_n2083 ), .A2(_u10_u8_n1869 ), .ZN(_u10_u8_n2068 ) );
NAND2_X1 _u10_u8_U118  ( .A1(_u10_u8_n2081 ), .A2(_u10_u8_n2082 ), .ZN(_u10_u8_n2075 ) );
NAND2_X1 _u10_u8_U117  ( .A1(_u10_u8_n2035 ), .A2(_u10_u8_n2019 ), .ZN(_u10_u8_n2060 ) );
NAND2_X1 _u10_u8_U116  ( .A1(_u10_u8_n2080 ), .A2(_u10_u8_n2060 ), .ZN(_u10_u8_n2079 ) );
NAND2_X1 _u10_u8_U115  ( .A1(_u10_u8_n2078 ), .A2(_u10_u8_n2079 ), .ZN(_u10_u8_n2076 ) );
NAND4_X1 _u10_u8_U114  ( .A1(_u10_u8_n2075 ), .A2(_u10_u8_n2076 ), .A3(_u10_u8_n1970 ), .A4(_u10_u8_n2077 ), .ZN(_u10_u8_n2072 ) );
NOR4_X1 _u10_u8_U113  ( .A1(_u10_u8_n2072 ), .A2(_u10_u8_n2073 ), .A3(_u10_u8_n1975 ), .A4(_u10_u8_n2074 ), .ZN(_u10_u8_n2070 ) );
NOR2_X1 _u10_u8_U112  ( .A1(_u10_u8_n2070 ), .A2(_u10_u8_n2071 ), .ZN(_u10_u8_n2069 ) );
NOR4_X1 _u10_u8_U111  ( .A1(_u10_u8_n2066 ), .A2(_u10_u8_n2067 ), .A3(_u10_u8_n2068 ), .A4(_u10_u8_n2069 ), .ZN(_u10_u8_n1820 ) );
NAND2_X1 _u10_u8_U110  ( .A1(1'b0), .A2(_u10_u8_n1983 ), .ZN(_u10_u8_n2065 ));
NAND4_X1 _u10_u8_U109  ( .A1(_u10_u8_n2065 ), .A2(_u10_u8_n2023 ), .A3(_u10_u8_n2021 ), .A4(_u10_u8_n2052 ), .ZN(_u10_u8_n2064 ) );
NAND2_X1 _u10_u8_U108  ( .A1(_u10_u8_n2063 ), .A2(_u10_u8_n2064 ), .ZN(_u10_u8_n2040 ) );
NAND4_X1 _u10_u8_U107  ( .A1(_u10_u8_n2059 ), .A2(_u10_u8_n2060 ), .A3(_u10_u8_n2061 ), .A4(_u10_u8_n2062 ), .ZN(_u10_u8_n2058 ) );
NAND2_X1 _u10_u8_U106  ( .A1(_u10_u8_n2057 ), .A2(_u10_u8_n2058 ), .ZN(_u10_u8_n2041 ) );
NOR4_X1 _u10_u8_U105  ( .A1(1'b0), .A2(_u10_u8_n2054 ), .A3(_u10_u8_n2055 ),.A4(_u10_u8_n2056 ), .ZN(_u10_u8_n2053 ) );
NAND4_X1 _u10_u8_U104  ( .A1(_u10_u8_n2021 ), .A2(_u10_u8_n2052 ), .A3(_u10_u8_n2023 ), .A4(_u10_u8_n2053 ), .ZN(_u10_u8_n1964 ) );
INV_X1 _u10_u8_U103  ( .A(_u10_u8_n1964 ), .ZN(_u10_u8_n2045 ) );
NAND2_X1 _u10_u8_U102  ( .A1(_u10_u8_n2051 ), .A2(_u10_SYNOPSYS_UNCONNECTED_37 ), .ZN(_u10_u8_n2046 ) );
NAND2_X1 _u10_u8_U101  ( .A1(_u10_u8_n2049 ), .A2(_u10_u8_n2050 ), .ZN(_u10_u8_n2047 ) );
NAND4_X1 _u10_u8_U100  ( .A1(_u10_u8_n2045 ), .A2(_u10_u8_n2046 ), .A3(_u10_u8_n2047 ), .A4(_u10_u8_n2048 ), .ZN(_u10_u8_n2044 ) );
NAND2_X1 _u10_u8_U99  ( .A1(_u10_u8_n2043 ), .A2(_u10_u8_n2044 ), .ZN(_u10_u8_n2042 ) );
NAND3_X1 _u10_u8_U98  ( .A1(_u10_u8_n2040 ), .A2(_u10_u8_n2041 ), .A3(_u10_u8_n2042 ), .ZN(_u10_u8_n2009 ) );
AND2_X1 _u10_u8_U97  ( .A1(_u10_u8_n2038 ), .A2(_u10_u8_n2039 ), .ZN(_u10_u8_n1929 ) );
NOR2_X1 _u10_u8_U96  ( .A1(_u10_u8_n1929 ), .A2(_u10_u8_n2037 ), .ZN(_u10_u8_n2010 ) );
NAND2_X1 _u10_u8_U95  ( .A1(_u10_u8_n2035 ), .A2(_u10_u8_n2036 ), .ZN(_u10_u8_n1902 ) );
NAND3_X1 _u10_u8_U94  ( .A1(_u10_u8_n1902 ), .A2(_u10_u8_n2033 ), .A3(_u10_u8_n2034 ), .ZN(_u10_u8_n1973 ) );
NOR2_X1 _u10_u8_U93  ( .A1(_u10_u8_n1978 ), .A2(_u10_u8_n1973 ), .ZN(_u10_u8_n2032 ) );
NOR2_X1 _u10_u8_U92  ( .A1(1'b0), .A2(_u10_u8_n2032 ), .ZN(_u10_u8_n2028 ));
NOR2_X1 _u10_u8_U91  ( .A1(_u10_u8_n2030 ), .A2(_u10_u8_n2031 ), .ZN(_u10_u8_n2029 ) );
NOR4_X1 _u10_u8_U90  ( .A1(_u10_u8_n2026 ), .A2(_u10_u8_n2027 ), .A3(_u10_u8_n2028 ), .A4(_u10_u8_n2029 ), .ZN(_u10_u8_n2024 ) );
NOR2_X1 _u10_u8_U89  ( .A1(_u10_u8_n2024 ), .A2(_u10_u8_n2025 ), .ZN(_u10_u8_n2011 ) );
NAND3_X1 _u10_u8_U88  ( .A1(_u10_u8_n2021 ), .A2(_u10_u8_n2022 ), .A3(_u10_u8_n2023 ), .ZN(_u10_u8_n2020 ) );
AND2_X1 _u10_u8_U87  ( .A1(_u10_u8_n2019 ), .A2(_u10_u8_n2020 ), .ZN(_u10_u8_n1838 ) );
INV_X1 _u10_u8_U86  ( .A(_u10_u8_n2018 ), .ZN(_u10_u8_n2016 ) );
NOR4_X1 _u10_u8_U85  ( .A1(_u10_u8_n2015 ), .A2(_u10_u8_n1838 ), .A3(_u10_u8_n2016 ), .A4(_u10_u8_n2017 ), .ZN(_u10_u8_n2013 ) );
NOR2_X1 _u10_u8_U84  ( .A1(_u10_u8_n2013 ), .A2(_u10_u8_n2014 ), .ZN(_u10_u8_n2012 ) );
NOR4_X1 _u10_u8_U83  ( .A1(_u10_u8_n2009 ), .A2(_u10_u8_n2010 ), .A3(_u10_u8_n2011 ), .A4(_u10_u8_n2012 ), .ZN(_u10_u8_n1821 ) );
NAND2_X1 _u10_u8_U82  ( .A1(_u10_u8_n1924 ), .A2(_u10_u8_n2008 ), .ZN(_u10_u8_n1993 ) );
NAND2_X1 _u10_u8_U81  ( .A1(_u10_u8_n2006 ), .A2(_u10_u8_n2007 ), .ZN(_u10_u8_n1994 ) );
NAND2_X1 _u10_u8_U80  ( .A1(_u10_u8_n2004 ), .A2(_u10_u8_n2005 ), .ZN(_u10_u8_n1995 ) );
AND2_X1 _u10_u8_U79  ( .A1(_u10_u8_n2002 ), .A2(_u10_u8_n2003 ), .ZN(_u10_u8_n1998 ) );
NOR2_X1 _u10_u8_U78  ( .A1(_u10_u8_n2000 ), .A2(_u10_u8_n2001 ), .ZN(_u10_u8_n1999 ) );
NOR3_X1 _u10_u8_U77  ( .A1(_u10_u8_n1997 ), .A2(_u10_u8_n1998 ), .A3(_u10_u8_n1999 ), .ZN(_u10_u8_n1996 ) );
NAND4_X1 _u10_u8_U76  ( .A1(_u10_u8_n1993 ), .A2(_u10_u8_n1994 ), .A3(_u10_u8_n1995 ), .A4(_u10_u8_n1996 ), .ZN(_u10_u8_n1985 ) );
INV_X1 _u10_u8_U75  ( .A(_u10_u8_n1992 ), .ZN(_u10_u8_n1989 ) );
NAND3_X1 _u10_u8_U74  ( .A1(_u10_u8_n1989 ), .A2(_u10_u8_n1990 ), .A3(_u10_u8_n1991 ), .ZN(_u10_u8_n1986 ) );
NOR4_X1 _u10_u8_U73  ( .A1(_u10_u8_n1985 ), .A2(_u10_u8_n1986 ), .A3(_u10_u8_n1987 ), .A4(_u10_u8_n1988 ), .ZN(_u10_u8_n1822 ) );
INV_X1 _u10_u8_U72  ( .A(_u10_u8_n1984 ), .ZN(_u10_u8_n1980 ) );
NAND4_X1 _u10_u8_U71  ( .A1(_u10_u8_n1980 ), .A2(_u10_u8_n1981 ), .A3(_u10_u8_n1982 ), .A4(_u10_u8_n1983 ), .ZN(_u10_u8_n1941 ) );
NOR3_X1 _u10_u8_U70  ( .A1(_u10_u8_n1977 ), .A2(_u10_u8_n1978 ), .A3(_u10_u8_n1979 ), .ZN(_u10_u8_n1971 ) );
NOR4_X1 _u10_u8_U69  ( .A1(_u10_u8_n1973 ), .A2(_u10_u8_n1974 ), .A3(_u10_u8_n1975 ), .A4(_u10_u8_n1976 ), .ZN(_u10_u8_n1972 ) );
NAND4_X1 _u10_u8_U68  ( .A1(_u10_u8_n1969 ), .A2(_u10_u8_n1970 ), .A3(_u10_u8_n1971 ), .A4(_u10_u8_n1972 ), .ZN(_u10_u8_n1968 ) );
NAND2_X1 _u10_u8_U67  ( .A1(_u10_u8_n1967 ), .A2(_u10_u8_n1968 ), .ZN(_u10_u8_n1942 ) );
NAND3_X1 _u10_u8_U66  ( .A1(_u10_u8_n1964 ), .A2(_u10_u8_n1965 ), .A3(_u10_u8_n1966 ), .ZN(_u10_u8_n1943 ) );
AND4_X1 _u10_u8_U65  ( .A1(_u10_u8_n1961 ), .A2(_u10_u8_n1863 ), .A3(_u10_u8_n1962 ), .A4(_u10_u8_n1963 ), .ZN(_u10_u8_n1957 ) );
NOR2_X1 _u10_u8_U64  ( .A1(_u10_u8_n1959 ), .A2(_u10_u8_n1960 ), .ZN(_u10_u8_n1958 ) );
NOR2_X1 _u10_u8_U63  ( .A1(_u10_u8_n1957 ), .A2(_u10_u8_n1958 ), .ZN(_u10_u8_n1945 ) );
NOR2_X1 _u10_u8_U62  ( .A1(_u10_u8_n1955 ), .A2(_u10_u8_n1956 ), .ZN(_u10_u8_n1953 ) );
NOR4_X1 _u10_u8_U61  ( .A1(_u10_u8_n1952 ), .A2(_u10_u8_n1953 ), .A3(_u10_u8_n1846 ), .A4(_u10_u8_n1954 ), .ZN(_u10_u8_n1946 ) );
NOR2_X1 _u10_u8_U60  ( .A1(_u10_u8_n1950 ), .A2(_u10_u8_n1951 ), .ZN(_u10_u8_n1949 ) );
NOR2_X1 _u10_u8_U59  ( .A1(_u10_u8_n1948 ), .A2(_u10_u8_n1949 ), .ZN(_u10_u8_n1947 ) );
NOR3_X1 _u10_u8_U58  ( .A1(_u10_u8_n1945 ), .A2(_u10_u8_n1946 ), .A3(_u10_u8_n1947 ), .ZN(_u10_u8_n1944 ) );
NAND4_X1 _u10_u8_U57  ( .A1(_u10_u8_n1941 ), .A2(_u10_u8_n1942 ), .A3(_u10_u8_n1943 ), .A4(_u10_u8_n1944 ), .ZN(_u10_u8_n1824 ) );
NAND2_X1 _u10_u8_U56  ( .A1(_u10_u8_n1939 ), .A2(_u10_u8_n1940 ), .ZN(_u10_u8_n1938 ) );
NAND2_X1 _u10_u8_U55  ( .A1(_u10_u8_n1937 ), .A2(_u10_u8_n1938 ), .ZN(_u10_u8_n1903 ) );
NAND2_X1 _u10_u8_U54  ( .A1(_u10_u8_n1935 ), .A2(_u10_u8_n1936 ), .ZN(_u10_u8_n1934 ) );
NAND2_X1 _u10_u8_U53  ( .A1(_u10_u8_n1933 ), .A2(_u10_u8_n1934 ), .ZN(_u10_u8_n1931 ) );
NAND2_X1 _u10_u8_U52  ( .A1(_u10_u8_n1931 ), .A2(_u10_u8_n1932 ), .ZN(_u10_u8_n1904 ) );
NAND2_X1 _u10_u8_U51  ( .A1(_u10_u8_n1929 ), .A2(_u10_u8_n1930 ), .ZN(_u10_u8_n1927 ) );
NAND2_X1 _u10_u8_U50  ( .A1(_u10_u8_n1927 ), .A2(_u10_u8_n1928 ), .ZN(_u10_u8_n1905 ) );
NOR3_X1 _u10_u8_U49  ( .A1(_u10_u8_n1916 ), .A2(_u10_u8_n1925 ), .A3(_u10_u8_n1926 ), .ZN(_u10_u8_n1919 ) );
NOR2_X1 _u10_u8_U48  ( .A1(_u10_u8_n1923 ), .A2(_u10_u8_n1924 ), .ZN(_u10_u8_n1921 ) );
NOR2_X1 _u10_u8_U47  ( .A1(_u10_u8_n1921 ), .A2(_u10_u8_n1922 ), .ZN(_u10_u8_n1920 ) );
NOR2_X1 _u10_u8_U46  ( .A1(_u10_u8_n1919 ), .A2(_u10_u8_n1920 ), .ZN(_u10_u8_n1917 ) );
NOR2_X1 _u10_u8_U45  ( .A1(_u10_u8_n1917 ), .A2(_u10_u8_n1918 ), .ZN(_u10_u8_n1907 ) );
NOR2_X1 _u10_u8_U44  ( .A1(_u10_u8_n1915 ), .A2(_u10_u8_n1916 ), .ZN(_u10_u8_n1914 ) );
NOR2_X1 _u10_u8_U43  ( .A1(_u10_u8_n1914 ), .A2(1'b0), .ZN(_u10_u8_n1912 ));
NOR2_X1 _u10_u8_U42  ( .A1(_u10_u8_n1912 ), .A2(_u10_u8_n1913 ), .ZN(_u10_u8_n1908 ) );
NOR2_X1 _u10_u8_U41  ( .A1(_u10_u8_n1891 ), .A2(_u10_u8_n1911 ), .ZN(_u10_u8_n1910 ) );
NOR2_X1 _u10_u8_U40  ( .A1(_u10_u8_n1910 ), .A2(_u10_u8_n1868 ), .ZN(_u10_u8_n1909 ) );
NOR3_X1 _u10_u8_U39  ( .A1(_u10_u8_n1907 ), .A2(_u10_u8_n1908 ), .A3(_u10_u8_n1909 ), .ZN(_u10_u8_n1906 ) );
NAND4_X1 _u10_u8_U38  ( .A1(_u10_u8_n1903 ), .A2(_u10_u8_n1904 ), .A3(_u10_u8_n1905 ), .A4(_u10_u8_n1906 ), .ZN(_u10_u8_n1825 ) );
NAND2_X1 _u10_u8_U37  ( .A1(_u10_u8_n1901 ), .A2(_u10_u8_n1902 ), .ZN(_u10_u8_n1900 ) );
NAND2_X1 _u10_u8_U36  ( .A1(_u10_u8_n1899 ), .A2(_u10_u8_n1900 ), .ZN(_u10_u8_n1875 ) );
OR2_X1 _u10_u8_U35  ( .A1(_u10_u8_n1847 ), .A2(_u10_u8_n1898 ), .ZN(_u10_u8_n1897 ) );
NAND2_X1 _u10_u8_U34  ( .A1(_u10_u8_n1896 ), .A2(_u10_u8_n1897 ), .ZN(_u10_u8_n1895 ) );
NAND2_X1 _u10_u8_U33  ( .A1(_u10_u8_n1894 ), .A2(_u10_u8_n1895 ), .ZN(_u10_u8_n1876 ) );
NAND2_X1 _u10_u8_U32  ( .A1(_u10_u8_n1892 ), .A2(_u10_u8_n1893 ), .ZN(_u10_u8_n1877 ) );
NOR3_X1 _u10_u8_U31  ( .A1(_u10_u8_n1884 ), .A2(_u10_u8_n1890 ), .A3(_u10_u8_n1891 ), .ZN(_u10_u8_n1889 ) );
NOR2_X1 _u10_u8_U30  ( .A1(_u10_u8_n1840 ), .A2(_u10_u8_n1889 ), .ZN(_u10_u8_n1879 ) );
NOR2_X1 _u10_u8_U29  ( .A1(_u10_u8_n1887 ), .A2(_u10_u8_n1888 ), .ZN(_u10_u8_n1880 ) );
NOR3_X1 _u10_u8_U28  ( .A1(_u10_u8_n1884 ), .A2(_u10_u8_n1885 ), .A3(_u10_u8_n1886 ), .ZN(_u10_u8_n1883 ) );
NOR2_X1 _u10_u8_U27  ( .A1(_u10_u8_n1882 ), .A2(_u10_u8_n1883 ), .ZN(_u10_u8_n1881 ) );
NOR3_X1 _u10_u8_U26  ( .A1(_u10_u8_n1879 ), .A2(_u10_u8_n1880 ), .A3(_u10_u8_n1881 ), .ZN(_u10_u8_n1878 ) );
NAND4_X1 _u10_u8_U25  ( .A1(_u10_u8_n1875 ), .A2(_u10_u8_n1876 ), .A3(_u10_u8_n1877 ), .A4(_u10_u8_n1878 ), .ZN(_u10_u8_n1826 ) );
NOR3_X1 _u10_u8_U24  ( .A1(_u10_u8_n1872 ), .A2(_u10_u8_n1873 ), .A3(_u10_u8_n1874 ), .ZN(_u10_u8_n1871 ) );
NAND4_X1 _u10_u8_U23  ( .A1(_u10_u8_n1868 ), .A2(_u10_u8_n1869 ), .A3(_u10_u8_n1870 ), .A4(_u10_u8_n1871 ), .ZN(_u10_u8_n1867 ) );
NAND2_X1 _u10_u8_U22  ( .A1(_u10_u8_n1866 ), .A2(_u10_u8_n1867 ), .ZN(_u10_u8_n1865 ) );
NAND3_X1 _u10_u8_U21  ( .A1(_u10_u8_n1863 ), .A2(_u10_u8_n1864 ), .A3(_u10_u8_n1865 ), .ZN(_u10_u8_n1862 ) );
NAND2_X1 _u10_u8_U20  ( .A1(_u10_u8_n1861 ), .A2(_u10_u8_n1862 ), .ZN(_u10_u8_n1828 ) );
NAND3_X1 _u10_u8_U19  ( .A1(_u10_u8_n1858 ), .A2(_u10_u8_n1859 ), .A3(_u10_u8_n1860 ), .ZN(_u10_u8_n1857 ) );
NAND2_X1 _u10_u8_U18  ( .A1(_u10_u8_n1856 ), .A2(_u10_u8_n1857 ), .ZN(_u10_u8_n1829 ) );
OR2_X1 _u10_u8_U17  ( .A1(_u10_u8_n1854 ), .A2(_u10_u8_n1855 ), .ZN(_u10_u8_n1830 ) );
NOR2_X1 _u10_u8_U16  ( .A1(_u10_u8_n1852 ), .A2(_u10_u8_n1853 ), .ZN(_u10_u8_n1850 ) );
NOR3_X1 _u10_u8_U15  ( .A1(_u10_u8_n1850 ), .A2(_u10_u8_n1851 ), .A3(_u10_u8_n1838 ), .ZN(_u10_u8_n1848 ) );
NOR2_X1 _u10_u8_U14  ( .A1(_u10_u8_n1848 ), .A2(_u10_u8_n1849 ), .ZN(_u10_u8_n1832 ) );
NOR2_X1 _u10_u8_U13  ( .A1(_u10_u8_n1846 ), .A2(_u10_u8_n1847 ), .ZN(_u10_u8_n1845 ) );
NOR3_X1 _u10_u8_U12  ( .A1(_u10_u8_n1844 ), .A2(1'b0), .A3(_u10_u8_n1845 ),.ZN(_u10_u8_n1842 ) );
NOR2_X1 _u10_u8_U11  ( .A1(_u10_u8_n1842 ), .A2(_u10_u8_n1843 ), .ZN(_u10_u8_n1833 ) );
NOR2_X1 _u10_u8_U10  ( .A1(_u10_u8_n1840 ), .A2(_u10_u8_n1841 ), .ZN(_u10_u8_n1839 ) );
NOR3_X1 _u10_u8_U9  ( .A1(_u10_u8_n1837 ), .A2(_u10_u8_n1838 ), .A3(_u10_u8_n1839 ), .ZN(_u10_u8_n1835 ) );
NOR2_X1 _u10_u8_U8  ( .A1(_u10_u8_n1835 ), .A2(_u10_u8_n1836 ), .ZN(_u10_u8_n1834 ) );
NOR3_X1 _u10_u8_U7  ( .A1(_u10_u8_n1832 ), .A2(_u10_u8_n1833 ), .A3(_u10_u8_n1834 ), .ZN(_u10_u8_n1831 ) );
NAND4_X1 _u10_u8_U6  ( .A1(_u10_u8_n1828 ), .A2(_u10_u8_n1829 ), .A3(_u10_u8_n1830 ), .A4(_u10_u8_n1831 ), .ZN(_u10_u8_n1827 ) );
NOR4_X1 _u10_u8_U5  ( .A1(_u10_u8_n1824 ), .A2(_u10_u8_n1825 ), .A3(_u10_u8_n1826 ), .A4(_u10_u8_n1827 ), .ZN(_u10_u8_n1823 ) );
NAND4_X1 _u10_u8_U4  ( .A1(_u10_u8_n1820 ), .A2(_u10_u8_n1821 ), .A3(_u10_u8_n1822 ), .A4(_u10_u8_n1823 ), .ZN(_u10_u8_n1818 ) );
MUX2_X1 _u10_u8_U3  ( .A(_u10_u8_n1818 ), .B(_u10_SYNOPSYS_UNCONNECTED_37 ),.S(_u10_u8_n1819 ), .Z(_u10_u8_n1812 ) );
DFFR_X1 _u10_u8_state_reg_1_  ( .D(_u10_u8_n1812 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_37 ), .QN(_u10_u8_n1814 ));
DFFR_X1 _u10_u8_state_reg_2_  ( .D(_u10_u8_n1811 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_36 ), .QN(_u10_u8_n1815 ));
DFFR_X1 _u10_u8_state_reg_3_  ( .D(_u10_u8_n1810 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_35 ), .QN(_u10_u8_n1816 ));
DFFR_X1 _u10_u8_state_reg_4_  ( .D(_u10_u8_n1809 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_34 ), .QN(_u10_u8_n1817 ));
DFFR_X1 _u10_u8_state_reg_0_  ( .D(_u10_u8_n1808 ), .CK(clk_i), .RN(_u10_n12357 ), .Q(_u10_SYNOPSYS_UNCONNECTED_38 ), .QN(_u10_u8_n1813 ));
INV_X1 _u2_U1058  ( .A(csr[2]), .ZN(_u2_n1284 ) );
MUX2_X1 _u2_U1057  ( .A(mast1_drdy), .B(mast0_drdy), .S(_u2_n1284 ), .Z(_u2_n1267 ) );
NOR3_X1 _u2_U1056  ( .A1(_u2_n1267 ), .A2(dma_err), .A3(_u2_n722 ), .ZN(_u2_n1234 ) );
INV_X1 _u2_U1055  ( .A(_u2_n1234 ), .ZN(_u2_n1556 ) );
NOR3_X1 _u2_U1054  ( .A1(_u2_tsz_cnt[0] ), .A2(_u2_tsz_cnt[11] ), .A3(_u2_tsz_cnt[10] ), .ZN(_u2_n1560 ) );
NOR3_X1 _u2_U1053  ( .A1(_u2_tsz_cnt[1] ), .A2(_u2_tsz_cnt[3] ), .A3(_u2_tsz_cnt[2] ), .ZN(_u2_n1561 ) );
NOR3_X1 _u2_U1052  ( .A1(_u2_tsz_cnt[4] ), .A2(_u2_tsz_cnt[6] ), .A3(_u2_tsz_cnt[5] ), .ZN(_u2_n1562 ) );
NOR4_X1 _u2_U1051  ( .A1(txsz[15]), .A2(_u2_tsz_cnt[9] ), .A3(_u2_tsz_cnt[8] ), .A4(_u2_tsz_cnt[7] ), .ZN(_u2_n1563 ) );
NAND4_X1 _u2_U1050  ( .A1(_u2_n1560 ), .A2(_u2_n1561 ), .A3(_u2_n1562 ),.A4(_u2_n1563 ), .ZN(_u2_n765 ) );
NOR3_X1 _u2_U1049  ( .A1(_u2_chunk_cnt[6] ), .A2(_u2_chunk_cnt[8] ), .A3(_u2_chunk_cnt[7] ), .ZN(_u2_n1558 ) );
NOR4_X1 _u2_U1048  ( .A1(_u2_chunk_cnt[0] ), .A2(_u2_chunk_cnt[2] ), .A3(_u2_chunk_cnt[3] ), .A4(_u2_chunk_cnt[4] ), .ZN(_u2_n1559 ) );
AND4_X1 _u2_U1047  ( .A1(_u2_n1053 ), .A2(_u2_n1052 ), .A3(_u2_n1558 ), .A4(_u2_n1559 ), .ZN(_u2_n1044 ) );
NAND2_X1 _u2_U1046  ( .A1(_u2_n1044 ), .A2(_u2_n931 ), .ZN(_u2_n1557 ) );
NAND2_X1 _u2_U1045  ( .A1(_u2_n765 ), .A2(_u2_n1557 ), .ZN(_u2_n1165 ) );
INV_X1 _u2_U1044  ( .A(_u2_n1165 ), .ZN(_u2_n1274 ) );
MUX2_X1 _u2_U1043  ( .A(mast0_drdy), .B(mast1_drdy), .S(csr[1]), .Z(_u2_n1246 ) );
NAND4_X1 _u2_U1042  ( .A1(_u2_state_2_ ), .A2(_u2_n1006 ), .A3(_u2_n1274 ),.A4(_u2_n1246 ), .ZN(_u2_n1153 ) );
NOR2_X1 _u2_U1041  ( .A1(_u2_read_r ), .A2(_u2_n1418 ), .ZN(_u2_N232 ) );
OR3_X1 _u2_U1040  ( .A1(mast1_err), .A2(mast0_err), .A3(dma_abort), .ZN(_u2_N236 ) );
NAND3_X1 _u2_U1039  ( .A1(csr[8]), .A2(csr[7]), .A3(ndr), .ZN(_u2_n1148 ) );
NOR2_X1 _u2_U1038  ( .A1(_u2_n1148 ), .A2(_u2_n719 ), .ZN(_u2_n1151 ) );
NOR2_X1 _u2_U1037  ( .A1(_u2_n1151 ), .A2(_u2_state_9_ ), .ZN(_u2_n1551 ) );
NOR4_X1 _u2_U1036  ( .A1(_u2_state_4_ ), .A2(_u2_state_5_ ), .A3(_u2_state_6_ ), .A4(_u2_state_7_ ), .ZN(_u2_n1369 ) );
NAND2_X1 _u2_U1035  ( .A1(_u2_n1551 ), .A2(_u2_n728 ), .ZN(_u2_n1552 ) );
INV_X1 _u2_U1034  ( .A(_u2_n1151 ), .ZN(_u2_n1554 ) );
NOR3_X1 _u2_U1033  ( .A1(_u2_state_4_ ), .A2(_u2_state_6_ ), .A3(_u2_state_5_ ), .ZN(_u2_n1555 ) );
NAND3_X1 _u2_U1032  ( .A1(mast0_drdy), .A2(_u2_n1554 ), .A3(_u2_n1555 ),.ZN(_u2_n1553 ) );
NAND2_X1 _u2_U1031  ( .A1(_u2_n1552 ), .A2(_u2_n1553 ), .ZN(_u2_n1278 ) );
INV_X1 _u2_U1030  ( .A(_u2_n1278 ), .ZN(_u2_n1280 ) );
NAND2_X1 _u2_U1029  ( .A1(_u2_n1280 ), .A2(_u2_n1288 ), .ZN(_u2_n1275 ) );
AND2_X1 _u2_U1028  ( .A1(pointer_s[0]), .A2(_u2_n1429 ), .ZN(_u2_N277 ) );
AND2_X1 _u2_U1027  ( .A1(pointer_s[1]), .A2(_u2_n1429 ), .ZN(_u2_N278 ) );
NAND2_X1 _u2_U1026  ( .A1(pointer_s[2]), .A2(_u2_n1429 ), .ZN(_u2_n1544 ) );
NAND2_X1 _u2_U1025  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[0] ), .ZN(_u2_n1545 ) );
NAND2_X1 _u2_U1024  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[0] ), .ZN(_u2_n1546 ) );
NOR2_X1 _u2_U1023  ( .A1(_u2_state_4_ ), .A2(_u2_state_6_ ), .ZN(_u2_n1550 ));
MUX2_X1 _u2_U1022  ( .A(_u2_n723 ), .B(_u2_n1550 ), .S(mast0_drdy), .Z(_u2_n1549 ) );
NAND2_X1 _u2_U1021  ( .A1(_u2_n1549 ), .A2(_u2_n718 ), .ZN(_u2_n1548 ) );
NAND2_X1 _u2_U1020  ( .A1(_u2_n1426 ), .A2(_u2_n1548 ), .ZN(_u2_n1547 ) );
NAND4_X1 _u2_U1019  ( .A1(_u2_n1544 ), .A2(_u2_n1545 ), .A3(_u2_n1546 ),.A4(_u2_n1547 ), .ZN(_u2_N279 ) );
NAND2_X1 _u2_U1018  ( .A1(pointer_s[3]), .A2(_u2_n1429 ), .ZN(_u2_n1538 ) );
NAND2_X1 _u2_U1017  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[1] ), .ZN(_u2_n1539 ) );
NAND2_X1 _u2_U1016  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[1] ), .ZN(_u2_n1540 ) );
NAND2_X1 _u2_U1015  ( .A1(_u2_state_5_ ), .A2(mast0_drdy), .ZN(_u2_n1543 ));
NAND3_X1 _u2_U1014  ( .A1(_u2_n724 ), .A2(_u2_n718 ), .A3(_u2_n1543 ), .ZN(_u2_n1542 ) );
NAND2_X1 _u2_U1013  ( .A1(_u2_n1426 ), .A2(_u2_n1542 ), .ZN(_u2_n1541 ) );
NAND4_X1 _u2_U1012  ( .A1(_u2_n1538 ), .A2(_u2_n1539 ), .A3(_u2_n1540 ),.A4(_u2_n1541 ), .ZN(_u2_N280 ) );
NAND2_X1 _u2_U1011  ( .A1(pointer_s[4]), .A2(_u2_n1429 ), .ZN(_u2_n1534 ) );
NAND2_X1 _u2_U1010  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[2] ), .ZN(_u2_n1535 ) );
NAND2_X1 _u2_U1009  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[2] ), .ZN(_u2_n1536 ) );
NAND2_X1 _u2_U1008  ( .A1(pointer[4]), .A2(_u2_n1426 ), .ZN(_u2_n1537 ) );
NAND4_X1 _u2_U1007  ( .A1(_u2_n1534 ), .A2(_u2_n1535 ), .A3(_u2_n1536 ),.A4(_u2_n1537 ), .ZN(_u2_N281 ) );
NAND2_X1 _u2_U1006  ( .A1(pointer_s[5]), .A2(_u2_n1429 ), .ZN(_u2_n1530 ) );
NAND2_X1 _u2_U1005  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[3] ), .ZN(_u2_n1531 ) );
NAND2_X1 _u2_U1004  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[3] ), .ZN(_u2_n1532 ) );
NAND2_X1 _u2_U1003  ( .A1(pointer[5]), .A2(_u2_n1426 ), .ZN(_u2_n1533 ) );
NAND4_X1 _u2_U1002  ( .A1(_u2_n1530 ), .A2(_u2_n1531 ), .A3(_u2_n1532 ),.A4(_u2_n1533 ), .ZN(_u2_N282 ) );
NAND2_X1 _u2_U1001  ( .A1(pointer_s[6]), .A2(_u2_n1429 ), .ZN(_u2_n1526 ) );
NAND2_X1 _u2_U1000  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[4] ), .ZN(_u2_n1527 ) );
NAND2_X1 _u2_U999  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[4] ), .ZN(_u2_n1528 ));
NAND2_X1 _u2_U998  ( .A1(pointer[6]), .A2(_u2_n1426 ), .ZN(_u2_n1529 ) );
NAND4_X1 _u2_U997  ( .A1(_u2_n1526 ), .A2(_u2_n1527 ), .A3(_u2_n1528 ), .A4(_u2_n1529 ), .ZN(_u2_N283 ) );
NAND2_X1 _u2_U996  ( .A1(pointer_s[7]), .A2(_u2_n1429 ), .ZN(_u2_n1522 ) );
NAND2_X1 _u2_U995  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[5] ), .ZN(_u2_n1523 ));
NAND2_X1 _u2_U994  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[5] ), .ZN(_u2_n1524 ));
NAND2_X1 _u2_U993  ( .A1(pointer[7]), .A2(_u2_n1426 ), .ZN(_u2_n1525 ) );
NAND4_X1 _u2_U992  ( .A1(_u2_n1522 ), .A2(_u2_n1523 ), .A3(_u2_n1524 ), .A4(_u2_n1525 ), .ZN(_u2_N284 ) );
NAND2_X1 _u2_U991  ( .A1(pointer_s[8]), .A2(_u2_n1429 ), .ZN(_u2_n1518 ) );
NAND2_X1 _u2_U990  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[6] ), .ZN(_u2_n1519 ));
NAND2_X1 _u2_U989  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[6] ), .ZN(_u2_n1520 ));
NAND2_X1 _u2_U988  ( .A1(pointer[8]), .A2(_u2_n1426 ), .ZN(_u2_n1521 ) );
NAND4_X1 _u2_U987  ( .A1(_u2_n1518 ), .A2(_u2_n1519 ), .A3(_u2_n1520 ), .A4(_u2_n1521 ), .ZN(_u2_N285 ) );
NAND2_X1 _u2_U986  ( .A1(pointer_s[9]), .A2(_u2_n1429 ), .ZN(_u2_n1514 ) );
NAND2_X1 _u2_U985  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[7] ), .ZN(_u2_n1515 ));
NAND2_X1 _u2_U984  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[7] ), .ZN(_u2_n1516 ));
NAND2_X1 _u2_U983  ( .A1(pointer[9]), .A2(_u2_n1426 ), .ZN(_u2_n1517 ) );
NAND4_X1 _u2_U982  ( .A1(_u2_n1514 ), .A2(_u2_n1515 ), .A3(_u2_n1516 ), .A4(_u2_n1517 ), .ZN(_u2_N286 ) );
NAND2_X1 _u2_U981  ( .A1(pointer_s[10]), .A2(_u2_n1429 ), .ZN(_u2_n1510 ) );
NAND2_X1 _u2_U980  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[8] ), .ZN(_u2_n1511 ));
NAND2_X1 _u2_U979  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[8] ), .ZN(_u2_n1512 ));
NAND2_X1 _u2_U978  ( .A1(pointer[10]), .A2(_u2_n1426 ), .ZN(_u2_n1513 ) );
NAND4_X1 _u2_U977  ( .A1(_u2_n1510 ), .A2(_u2_n1511 ), .A3(_u2_n1512 ), .A4(_u2_n1513 ), .ZN(_u2_N287 ) );
NAND2_X1 _u2_U976  ( .A1(pointer_s[11]), .A2(_u2_n1429 ), .ZN(_u2_n1506 ) );
NAND2_X1 _u2_U975  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[9] ), .ZN(_u2_n1507 ));
NAND2_X1 _u2_U974  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[9] ), .ZN(_u2_n1508 ));
NAND2_X1 _u2_U973  ( .A1(pointer[11]), .A2(_u2_n1426 ), .ZN(_u2_n1509 ) );
NAND4_X1 _u2_U972  ( .A1(_u2_n1506 ), .A2(_u2_n1507 ), .A3(_u2_n1508 ), .A4(_u2_n1509 ), .ZN(_u2_N288 ) );
NAND2_X1 _u2_U971  ( .A1(pointer_s[12]), .A2(_u2_n1429 ), .ZN(_u2_n1502 ) );
NAND2_X1 _u2_U970  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[10] ), .ZN(_u2_n1503 ) );
NAND2_X1 _u2_U969  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[10] ), .ZN(_u2_n1504 ) );
NAND2_X1 _u2_U968  ( .A1(pointer[12]), .A2(_u2_n1426 ), .ZN(_u2_n1505 ) );
NAND4_X1 _u2_U967  ( .A1(_u2_n1502 ), .A2(_u2_n1503 ), .A3(_u2_n1504 ), .A4(_u2_n1505 ), .ZN(_u2_N289 ) );
NAND2_X1 _u2_U966  ( .A1(pointer_s[13]), .A2(_u2_n1429 ), .ZN(_u2_n1498 ) );
NAND2_X1 _u2_U965  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[11] ), .ZN(_u2_n1499 ) );
NAND2_X1 _u2_U964  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[11] ), .ZN(_u2_n1500 ) );
NAND2_X1 _u2_U963  ( .A1(pointer[13]), .A2(_u2_n1426 ), .ZN(_u2_n1501 ) );
NAND4_X1 _u2_U962  ( .A1(_u2_n1498 ), .A2(_u2_n1499 ), .A3(_u2_n1500 ), .A4(_u2_n1501 ), .ZN(_u2_N290 ) );
NAND2_X1 _u2_U961  ( .A1(pointer_s[14]), .A2(_u2_n1429 ), .ZN(_u2_n1494 ) );
NAND2_X1 _u2_U960  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[12] ), .ZN(_u2_n1495 ) );
NAND2_X1 _u2_U959  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[12] ), .ZN(_u2_n1496 ) );
NAND2_X1 _u2_U958  ( .A1(pointer[14]), .A2(_u2_n1426 ), .ZN(_u2_n1497 ) );
NAND4_X1 _u2_U957  ( .A1(_u2_n1494 ), .A2(_u2_n1495 ), .A3(_u2_n1496 ), .A4(_u2_n1497 ), .ZN(_u2_N291 ) );
NAND2_X1 _u2_U956  ( .A1(pointer_s[15]), .A2(_u2_n1429 ), .ZN(_u2_n1490 ) );
NAND2_X1 _u2_U955  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[13] ), .ZN(_u2_n1491 ) );
NAND2_X1 _u2_U954  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[13] ), .ZN(_u2_n1492 ) );
NAND2_X1 _u2_U953  ( .A1(pointer[15]), .A2(_u2_n1426 ), .ZN(_u2_n1493 ) );
NAND4_X1 _u2_U952  ( .A1(_u2_n1490 ), .A2(_u2_n1491 ), .A3(_u2_n1492 ), .A4(_u2_n1493 ), .ZN(_u2_N292 ) );
NAND2_X1 _u2_U951  ( .A1(pointer_s[16]), .A2(_u2_n1429 ), .ZN(_u2_n1486 ) );
NAND2_X1 _u2_U950  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[14] ), .ZN(_u2_n1487 ) );
NAND2_X1 _u2_U949  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[14] ), .ZN(_u2_n1488 ) );
NAND2_X1 _u2_U948  ( .A1(pointer[16]), .A2(_u2_n1426 ), .ZN(_u2_n1489 ) );
NAND4_X1 _u2_U947  ( .A1(_u2_n1486 ), .A2(_u2_n1487 ), .A3(_u2_n1488 ), .A4(_u2_n1489 ), .ZN(_u2_N293 ) );
NAND2_X1 _u2_U946  ( .A1(pointer_s[17]), .A2(_u2_n1429 ), .ZN(_u2_n1482 ) );
NAND2_X1 _u2_U945  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[15] ), .ZN(_u2_n1483 ) );
NAND2_X1 _u2_U944  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[15] ), .ZN(_u2_n1484 ) );
NAND2_X1 _u2_U943  ( .A1(pointer[17]), .A2(_u2_n1426 ), .ZN(_u2_n1485 ) );
NAND4_X1 _u2_U942  ( .A1(_u2_n1482 ), .A2(_u2_n1483 ), .A3(_u2_n1484 ), .A4(_u2_n1485 ), .ZN(_u2_N294 ) );
NAND2_X1 _u2_U941  ( .A1(pointer_s[18]), .A2(_u2_n1429 ), .ZN(_u2_n1478 ) );
NAND2_X1 _u2_U940  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[16] ), .ZN(_u2_n1479 ) );
NAND2_X1 _u2_U939  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[16] ), .ZN(_u2_n1480 ) );
NAND2_X1 _u2_U938  ( .A1(pointer[18]), .A2(_u2_n1426 ), .ZN(_u2_n1481 ) );
NAND4_X1 _u2_U937  ( .A1(_u2_n1478 ), .A2(_u2_n1479 ), .A3(_u2_n1480 ), .A4(_u2_n1481 ), .ZN(_u2_N295 ) );
NAND2_X1 _u2_U936  ( .A1(pointer_s[19]), .A2(_u2_n1429 ), .ZN(_u2_n1474 ) );
NAND2_X1 _u2_U935  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[17] ), .ZN(_u2_n1475 ) );
NAND2_X1 _u2_U934  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[17] ), .ZN(_u2_n1476 ) );
NAND2_X1 _u2_U933  ( .A1(pointer[19]), .A2(_u2_n1426 ), .ZN(_u2_n1477 ) );
NAND4_X1 _u2_U932  ( .A1(_u2_n1474 ), .A2(_u2_n1475 ), .A3(_u2_n1476 ), .A4(_u2_n1477 ), .ZN(_u2_N296 ) );
NAND2_X1 _u2_U931  ( .A1(pointer_s[20]), .A2(_u2_n1429 ), .ZN(_u2_n1470 ) );
NAND2_X1 _u2_U930  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[18] ), .ZN(_u2_n1471 ) );
NAND2_X1 _u2_U929  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[18] ), .ZN(_u2_n1472 ) );
NAND2_X1 _u2_U928  ( .A1(pointer[20]), .A2(_u2_n1426 ), .ZN(_u2_n1473 ) );
NAND4_X1 _u2_U927  ( .A1(_u2_n1470 ), .A2(_u2_n1471 ), .A3(_u2_n1472 ), .A4(_u2_n1473 ), .ZN(_u2_N297 ) );
NAND2_X1 _u2_U926  ( .A1(pointer_s[21]), .A2(_u2_n1429 ), .ZN(_u2_n1466 ) );
NAND2_X1 _u2_U925  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[19] ), .ZN(_u2_n1467 ) );
NAND2_X1 _u2_U924  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[19] ), .ZN(_u2_n1468 ) );
NAND2_X1 _u2_U923  ( .A1(pointer[21]), .A2(_u2_n1426 ), .ZN(_u2_n1469 ) );
NAND4_X1 _u2_U922  ( .A1(_u2_n1466 ), .A2(_u2_n1467 ), .A3(_u2_n1468 ), .A4(_u2_n1469 ), .ZN(_u2_N298 ) );
NAND2_X1 _u2_U921  ( .A1(pointer_s[22]), .A2(_u2_n1429 ), .ZN(_u2_n1462 ) );
NAND2_X1 _u2_U920  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[20] ), .ZN(_u2_n1463 ) );
NAND2_X1 _u2_U919  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[20] ), .ZN(_u2_n1464 ) );
NAND2_X1 _u2_U918  ( .A1(pointer[22]), .A2(_u2_n1426 ), .ZN(_u2_n1465 ) );
NAND4_X1 _u2_U917  ( .A1(_u2_n1462 ), .A2(_u2_n1463 ), .A3(_u2_n1464 ), .A4(_u2_n1465 ), .ZN(_u2_N299 ) );
NAND2_X1 _u2_U916  ( .A1(pointer_s[23]), .A2(_u2_n1429 ), .ZN(_u2_n1458 ) );
NAND2_X1 _u2_U915  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[21] ), .ZN(_u2_n1459 ) );
NAND2_X1 _u2_U914  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[21] ), .ZN(_u2_n1460 ) );
NAND2_X1 _u2_U913  ( .A1(pointer[23]), .A2(_u2_n1426 ), .ZN(_u2_n1461 ) );
NAND4_X1 _u2_U912  ( .A1(_u2_n1458 ), .A2(_u2_n1459 ), .A3(_u2_n1460 ), .A4(_u2_n1461 ), .ZN(_u2_N300 ) );
NAND2_X1 _u2_U911  ( .A1(pointer_s[24]), .A2(_u2_n1429 ), .ZN(_u2_n1454 ) );
NAND2_X1 _u2_U910  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[22] ), .ZN(_u2_n1455 ) );
NAND2_X1 _u2_U909  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[22] ), .ZN(_u2_n1456 ) );
NAND2_X1 _u2_U908  ( .A1(pointer[24]), .A2(_u2_n1426 ), .ZN(_u2_n1457 ) );
NAND4_X1 _u2_U907  ( .A1(_u2_n1454 ), .A2(_u2_n1455 ), .A3(_u2_n1456 ), .A4(_u2_n1457 ), .ZN(_u2_N301 ) );
NAND2_X1 _u2_U906  ( .A1(pointer_s[25]), .A2(_u2_n1429 ), .ZN(_u2_n1450 ) );
NAND2_X1 _u2_U905  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[23] ), .ZN(_u2_n1451 ) );
NAND2_X1 _u2_U904  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[23] ), .ZN(_u2_n1452 ) );
NAND2_X1 _u2_U903  ( .A1(pointer[25]), .A2(_u2_n1426 ), .ZN(_u2_n1453 ) );
NAND4_X1 _u2_U902  ( .A1(_u2_n1450 ), .A2(_u2_n1451 ), .A3(_u2_n1452 ), .A4(_u2_n1453 ), .ZN(_u2_N302 ) );
NAND2_X1 _u2_U901  ( .A1(pointer_s[26]), .A2(_u2_n1429 ), .ZN(_u2_n1446 ) );
NAND2_X1 _u2_U900  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[24] ), .ZN(_u2_n1447 ) );
NAND2_X1 _u2_U899  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[24] ), .ZN(_u2_n1448 ) );
NAND2_X1 _u2_U898  ( .A1(pointer[26]), .A2(_u2_n1426 ), .ZN(_u2_n1449 ) );
NAND4_X1 _u2_U897  ( .A1(_u2_n1446 ), .A2(_u2_n1447 ), .A3(_u2_n1448 ), .A4(_u2_n1449 ), .ZN(_u2_N303 ) );
NAND2_X1 _u2_U896  ( .A1(pointer_s[27]), .A2(_u2_n1429 ), .ZN(_u2_n1442 ) );
NAND2_X1 _u2_U895  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[25] ), .ZN(_u2_n1443 ) );
NAND2_X1 _u2_U894  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[25] ), .ZN(_u2_n1444 ) );
NAND2_X1 _u2_U893  ( .A1(pointer[27]), .A2(_u2_n1426 ), .ZN(_u2_n1445 ) );
NAND4_X1 _u2_U892  ( .A1(_u2_n1442 ), .A2(_u2_n1443 ), .A3(_u2_n1444 ), .A4(_u2_n1445 ), .ZN(_u2_N304 ) );
NAND2_X1 _u2_U891  ( .A1(pointer_s[28]), .A2(_u2_n1429 ), .ZN(_u2_n1438 ) );
NAND2_X1 _u2_U890  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[26] ), .ZN(_u2_n1439 ) );
NAND2_X1 _u2_U889  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[26] ), .ZN(_u2_n1440 ) );
NAND2_X1 _u2_U888  ( .A1(pointer[28]), .A2(_u2_n1426 ), .ZN(_u2_n1441 ) );
NAND4_X1 _u2_U887  ( .A1(_u2_n1438 ), .A2(_u2_n1439 ), .A3(_u2_n1440 ), .A4(_u2_n1441 ), .ZN(_u2_N305 ) );
NAND2_X1 _u2_U886  ( .A1(pointer_s[29]), .A2(_u2_n1429 ), .ZN(_u2_n1434 ) );
NAND2_X1 _u2_U885  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[27] ), .ZN(_u2_n1435 ) );
NAND2_X1 _u2_U884  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[27] ), .ZN(_u2_n1436 ) );
NAND2_X1 _u2_U883  ( .A1(pointer[29]), .A2(_u2_n1426 ), .ZN(_u2_n1437 ) );
NAND4_X1 _u2_U882  ( .A1(_u2_n1434 ), .A2(_u2_n1435 ), .A3(_u2_n1436 ), .A4(_u2_n1437 ), .ZN(_u2_N306 ) );
NAND2_X1 _u2_U881  ( .A1(pointer_s[30]), .A2(_u2_n1429 ), .ZN(_u2_n1430 ) );
NAND2_X1 _u2_U880  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[28] ), .ZN(_u2_n1431 ) );
NAND2_X1 _u2_U879  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[28] ), .ZN(_u2_n1432 ) );
NAND2_X1 _u2_U878  ( .A1(pointer[30]), .A2(_u2_n1426 ), .ZN(_u2_n1433 ) );
NAND4_X1 _u2_U877  ( .A1(_u2_n1430 ), .A2(_u2_n1431 ), .A3(_u2_n1432 ), .A4(_u2_n1433 ), .ZN(_u2_N307 ) );
NAND2_X1 _u2_U876  ( .A1(pointer_s[31]), .A2(_u2_n1429 ), .ZN(_u2_n1422 ) );
NAND2_X1 _u2_U875  ( .A1(_u2_n1428 ), .A2(_u2_adr0_cnt[29] ), .ZN(_u2_n1423 ) );
NAND2_X1 _u2_U874  ( .A1(_u2_n1427 ), .A2(_u2_adr1_cnt[29] ), .ZN(_u2_n1424 ) );
NAND2_X1 _u2_U873  ( .A1(pointer[31]), .A2(_u2_n1426 ), .ZN(_u2_n1425 ) );
NAND4_X1 _u2_U872  ( .A1(_u2_n1422 ), .A2(_u2_n1423 ), .A3(_u2_n1424 ), .A4(_u2_n1425 ), .ZN(_u2_N308 ) );
MUX2_X1 _u2_U871  ( .A(_u2_adr0_cnt[0] ), .B(_u2_adr1_cnt[0] ), .S(_u2_n1418 ), .Z(_u2_N312 ) );
MUX2_X1 _u2_U870  ( .A(_u2_adr0_cnt[1] ), .B(_u2_adr1_cnt[1] ), .S(_u2_n1418 ), .Z(_u2_N313 ) );
MUX2_X1 _u2_U869  ( .A(_u2_adr0_cnt[2] ), .B(_u2_adr1_cnt[2] ), .S(_u2_n1418 ), .Z(_u2_N314 ) );
MUX2_X1 _u2_U868  ( .A(_u2_adr0_cnt[3] ), .B(_u2_adr1_cnt[3] ), .S(_u2_n1418 ), .Z(_u2_N315 ) );
MUX2_X1 _u2_U867  ( .A(_u2_adr0_cnt[4] ), .B(_u2_adr1_cnt[4] ), .S(_u2_n1418 ), .Z(_u2_N316 ) );
MUX2_X1 _u2_U866  ( .A(_u2_adr0_cnt[5] ), .B(_u2_adr1_cnt[5] ), .S(_u2_n1418 ), .Z(_u2_N317 ) );
MUX2_X1 _u2_U865  ( .A(_u2_adr0_cnt[6] ), .B(_u2_adr1_cnt[6] ), .S(_u2_n1418 ), .Z(_u2_N318 ) );
MUX2_X1 _u2_U864  ( .A(_u2_adr0_cnt[7] ), .B(_u2_adr1_cnt[7] ), .S(_u2_n1418 ), .Z(_u2_N319 ) );
MUX2_X1 _u2_U863  ( .A(_u2_adr0_cnt[8] ), .B(_u2_adr1_cnt[8] ), .S(_u2_n1418 ), .Z(_u2_N320 ) );
MUX2_X1 _u2_U862  ( .A(_u2_adr0_cnt[9] ), .B(_u2_adr1_cnt[9] ), .S(_u2_n1418 ), .Z(_u2_N321 ) );
MUX2_X1 _u2_U861  ( .A(_u2_adr0_cnt[10] ), .B(_u2_adr1_cnt[10] ), .S(_u2_n1418 ), .Z(_u2_N322 ) );
MUX2_X1 _u2_U860  ( .A(_u2_adr0_cnt[11] ), .B(_u2_adr1_cnt[11] ), .S(_u2_n1418 ), .Z(_u2_N323 ) );
MUX2_X1 _u2_U859  ( .A(_u2_adr0_cnt[12] ), .B(_u2_adr1_cnt[12] ), .S(_u2_n1418 ), .Z(_u2_N324 ) );
MUX2_X1 _u2_U858  ( .A(_u2_adr0_cnt[13] ), .B(_u2_adr1_cnt[13] ), .S(_u2_n1418 ), .Z(_u2_N325 ) );
MUX2_X1 _u2_U857  ( .A(_u2_adr0_cnt[14] ), .B(_u2_adr1_cnt[14] ), .S(_u2_n1418 ), .Z(_u2_N326 ) );
MUX2_X1 _u2_U856  ( .A(_u2_adr0_cnt[15] ), .B(_u2_adr1_cnt[15] ), .S(_u2_n1418 ), .Z(_u2_N327 ) );
MUX2_X1 _u2_U855  ( .A(_u2_adr0_cnt[16] ), .B(_u2_adr1_cnt[16] ), .S(_u2_n1418 ), .Z(_u2_N328 ) );
MUX2_X1 _u2_U854  ( .A(_u2_adr0_cnt[17] ), .B(_u2_adr1_cnt[17] ), .S(_u2_n1418 ), .Z(_u2_N329 ) );
MUX2_X1 _u2_U853  ( .A(_u2_adr0_cnt[18] ), .B(_u2_adr1_cnt[18] ), .S(_u2_n1418 ), .Z(_u2_N330 ) );
MUX2_X1 _u2_U852  ( .A(_u2_adr0_cnt[19] ), .B(_u2_adr1_cnt[19] ), .S(_u2_n1418 ), .Z(_u2_N331 ) );
MUX2_X1 _u2_U851  ( .A(_u2_adr0_cnt[20] ), .B(_u2_adr1_cnt[20] ), .S(_u2_n1418 ), .Z(_u2_N332 ) );
MUX2_X1 _u2_U850  ( .A(_u2_adr0_cnt[21] ), .B(_u2_adr1_cnt[21] ), .S(_u2_n1418 ), .Z(_u2_N333 ) );
MUX2_X1 _u2_U849  ( .A(_u2_adr0_cnt[22] ), .B(_u2_adr1_cnt[22] ), .S(_u2_n1418 ), .Z(_u2_N334 ) );
MUX2_X1 _u2_U848  ( .A(_u2_adr0_cnt[23] ), .B(_u2_adr1_cnt[23] ), .S(_u2_n1418 ), .Z(_u2_N335 ) );
MUX2_X1 _u2_U847  ( .A(_u2_adr0_cnt[24] ), .B(_u2_adr1_cnt[24] ), .S(_u2_n1418 ), .Z(_u2_N336 ) );
MUX2_X1 _u2_U846  ( .A(_u2_adr0_cnt[25] ), .B(_u2_adr1_cnt[25] ), .S(_u2_n1418 ), .Z(_u2_N337 ) );
MUX2_X1 _u2_U845  ( .A(_u2_adr0_cnt[26] ), .B(_u2_adr1_cnt[26] ), .S(_u2_n1418 ), .Z(_u2_N338 ) );
MUX2_X1 _u2_U844  ( .A(_u2_adr0_cnt[27] ), .B(_u2_adr1_cnt[27] ), .S(_u2_n1418 ), .Z(_u2_N339 ) );
MUX2_X1 _u2_U843  ( .A(_u2_adr0_cnt[28] ), .B(_u2_adr1_cnt[28] ), .S(_u2_n1418 ), .Z(_u2_N340 ) );
MUX2_X1 _u2_U842  ( .A(_u2_adr0_cnt[29] ), .B(_u2_adr1_cnt[29] ), .S(_u2_n1418 ), .Z(_u2_N341 ) );
NAND2_X1 _u2_U841  ( .A1(_u2_state_1_ ), .A2(_u2_n1267 ), .ZN(_u2_n1420 ) );
INV_X1 _u2_U840  ( .A(_u2_n1246 ), .ZN(_u2_n1421 ) );
NAND2_X1 _u2_U839  ( .A1(_u2_n1421 ), .A2(_u2_state_2_ ), .ZN(_u2_n1239 ) );
NAND2_X1 _u2_U838  ( .A1(_u2_n1420 ), .A2(_u2_n1239 ), .ZN(_u2_n1419 ) );
NAND2_X1 _u2_U837  ( .A1(_u2_n1006 ), .A2(_u2_n1419 ), .ZN(_u2_n1270 ) );
NAND2_X1 _u2_U836  ( .A1(_u2_n1270 ), .A2(_u2_n1418 ), .ZN(_u2_N342 ) );
NAND2_X1 _u2_U835  ( .A1(_u2_n727 ), .A2(_u2_n720 ), .ZN(de_fetch_descr) );
INV_X1 _u2_U834  ( .A(de_fetch_descr), .ZN(_u2_n1415 ) );
NOR2_X1 _u2_U833  ( .A1(_u2_state_9_ ), .A2(paused), .ZN(_u2_n1146 ) );
INV_X1 _u2_U832  ( .A(_u2_n1146 ), .ZN(_u2_n1417 ) );
OR2_X1 _u2_U831  ( .A1(_u2_state_2_ ), .A2(_u2_state_1_ ), .ZN(_u2_n1164 ));
NOR2_X1 _u2_U830  ( .A1(_u2_n1417 ), .A2(_u2_n1164 ), .ZN(_u2_n1416 ) );
NOR2_X1 _u2_U829  ( .A1(_u2_n1274 ), .A2(_u2_n719 ), .ZN(de_ack) );
NAND2_X1 _u2_U828  ( .A1(mast0_dout[0]), .A2(_u2_n726 ), .ZN(_u2_n1390 ) );
INV_X1 _u2_U827  ( .A(_u2_n1390 ), .ZN(de_adr0[0]) );
NAND2_X1 _u2_U826  ( .A1(mast0_dout[10]), .A2(_u2_n726 ), .ZN(_u2_n1388 ) );
NAND2_X1 _u2_U825  ( .A1(_u2_n728 ), .A2(_u2_adr0_cnt[8] ), .ZN(_u2_n1414 ));
NAND2_X1 _u2_U824  ( .A1(_u2_n1388 ), .A2(_u2_n1414 ), .ZN(de_adr0[10]) );
NAND2_X1 _u2_U823  ( .A1(mast0_dout[11]), .A2(_u2_n726 ), .ZN(_u2_n1386 ) );
NAND2_X1 _u2_U822  ( .A1(_u2_n729 ), .A2(_u2_adr0_cnt[9] ), .ZN(_u2_n1413 ));
NAND2_X1 _u2_U821  ( .A1(_u2_n1386 ), .A2(_u2_n1413 ), .ZN(de_adr0[11]) );
MUX2_X1 _u2_U820  ( .A(mast0_dout[12]), .B(_u2_adr0_cnt[10] ), .S(_u2_n727 ),.Z(de_adr0[12]) );
MUX2_X1 _u2_U819  ( .A(mast0_dout[13]), .B(_u2_adr0_cnt[11] ), .S(_u2_n728 ),.Z(de_adr0[13]) );
MUX2_X1 _u2_U818  ( .A(mast0_dout[14]), .B(_u2_adr0_cnt[12] ), .S(_u2_n729 ),.Z(de_adr0[14]) );
MUX2_X1 _u2_U817  ( .A(mast0_dout[15]), .B(_u2_adr0_cnt[13] ), .S(_u2_n1369 ), .Z(de_adr0[15]) );
MUX2_X1 _u2_U816  ( .A(mast0_dout[16]), .B(_u2_adr0_cnt[14] ), .S(_u2_n727 ),.Z(de_adr0[16]) );
MUX2_X1 _u2_U815  ( .A(mast0_dout[17]), .B(_u2_adr0_cnt[15] ), .S(_u2_n728 ),.Z(de_adr0[17]) );
MUX2_X1 _u2_U814  ( .A(mast0_dout[18]), .B(_u2_adr0_cnt[16] ), .S(_u2_n729 ),.Z(de_adr0[18]) );
MUX2_X1 _u2_U813  ( .A(mast0_dout[19]), .B(_u2_adr0_cnt[17] ), .S(_u2_n1369 ), .Z(de_adr0[19]) );
NAND2_X1 _u2_U812  ( .A1(mast0_dout[1]), .A2(_u2_n726 ), .ZN(_u2_n1384 ) );
INV_X1 _u2_U811  ( .A(_u2_n1384 ), .ZN(de_adr0[1]) );
MUX2_X1 _u2_U810  ( .A(mast0_dout[20]), .B(_u2_adr0_cnt[18] ), .S(_u2_n727 ),.Z(de_adr0[20]) );
MUX2_X1 _u2_U809  ( .A(mast0_dout[21]), .B(_u2_adr0_cnt[19] ), .S(_u2_n728 ),.Z(de_adr0[21]) );
MUX2_X1 _u2_U808  ( .A(mast0_dout[22]), .B(_u2_adr0_cnt[20] ), .S(_u2_n729 ),.Z(de_adr0[22]) );
MUX2_X1 _u2_U807  ( .A(mast0_dout[23]), .B(_u2_adr0_cnt[21] ), .S(_u2_n1369 ), .Z(de_adr0[23]) );
MUX2_X1 _u2_U806  ( .A(mast0_dout[24]), .B(_u2_adr0_cnt[22] ), .S(_u2_n727 ),.Z(de_adr0[24]) );
MUX2_X1 _u2_U805  ( .A(mast0_dout[25]), .B(_u2_adr0_cnt[23] ), .S(_u2_n728 ),.Z(de_adr0[25]) );
MUX2_X1 _u2_U804  ( .A(mast0_dout[26]), .B(_u2_adr0_cnt[24] ), .S(_u2_n729 ),.Z(de_adr0[26]) );
MUX2_X1 _u2_U803  ( .A(mast0_dout[27]), .B(_u2_adr0_cnt[25] ), .S(_u2_n1369 ), .Z(de_adr0[27]) );
MUX2_X1 _u2_U802  ( .A(mast0_dout[28]), .B(_u2_adr0_cnt[26] ), .S(_u2_n727 ),.Z(de_adr0[28]) );
MUX2_X1 _u2_U801  ( .A(mast0_dout[29]), .B(_u2_adr0_cnt[27] ), .S(_u2_n728 ),.Z(de_adr0[29]) );
NAND2_X1 _u2_U800  ( .A1(mast0_dout[2]), .A2(_u2_n726 ), .ZN(_u2_n1382 ) );
NAND2_X1 _u2_U799  ( .A1(_u2_n1369 ), .A2(_u2_adr0_cnt[0] ), .ZN(_u2_n1412 ));
NAND2_X1 _u2_U798  ( .A1(_u2_n1382 ), .A2(_u2_n1412 ), .ZN(de_adr0[2]) );
MUX2_X1 _u2_U797  ( .A(mast0_dout[30]), .B(_u2_adr0_cnt[28] ), .S(_u2_n729 ),.Z(de_adr0[30]) );
MUX2_X1 _u2_U796  ( .A(mast0_dout[31]), .B(_u2_adr0_cnt[29] ), .S(_u2_n1369 ), .Z(de_adr0[31]) );
NAND2_X1 _u2_U795  ( .A1(mast0_dout[3]), .A2(_u2_n726 ), .ZN(_u2_n1380 ) );
NAND2_X1 _u2_U794  ( .A1(_u2_n727 ), .A2(_u2_adr0_cnt[1] ), .ZN(_u2_n1411 ));
NAND2_X1 _u2_U793  ( .A1(_u2_n1380 ), .A2(_u2_n1411 ), .ZN(de_adr0[3]) );
NAND2_X1 _u2_U792  ( .A1(mast0_dout[4]), .A2(_u2_n726 ), .ZN(_u2_n1378 ) );
NAND2_X1 _u2_U791  ( .A1(_u2_n728 ), .A2(_u2_adr0_cnt[2] ), .ZN(_u2_n1410 ));
NAND2_X1 _u2_U790  ( .A1(_u2_n1378 ), .A2(_u2_n1410 ), .ZN(de_adr0[4]) );
NAND2_X1 _u2_U789  ( .A1(mast0_dout[5]), .A2(_u2_n726 ), .ZN(_u2_n1376 ) );
NAND2_X1 _u2_U788  ( .A1(_u2_n729 ), .A2(_u2_adr0_cnt[3] ), .ZN(_u2_n1409 ));
NAND2_X1 _u2_U787  ( .A1(_u2_n1376 ), .A2(_u2_n1409 ), .ZN(de_adr0[5]) );
NAND2_X1 _u2_U786  ( .A1(mast0_dout[6]), .A2(_u2_n726 ), .ZN(_u2_n1374 ) );
NAND2_X1 _u2_U785  ( .A1(_u2_n1369 ), .A2(_u2_adr0_cnt[4] ), .ZN(_u2_n1408 ));
NAND2_X1 _u2_U784  ( .A1(_u2_n1374 ), .A2(_u2_n1408 ), .ZN(de_adr0[6]) );
NAND2_X1 _u2_U783  ( .A1(mast0_dout[7]), .A2(_u2_n726 ), .ZN(_u2_n1372 ) );
NAND2_X1 _u2_U782  ( .A1(_u2_n727 ), .A2(_u2_adr0_cnt[5] ), .ZN(_u2_n1407 ));
NAND2_X1 _u2_U781  ( .A1(_u2_n1372 ), .A2(_u2_n1407 ), .ZN(de_adr0[7]) );
NAND2_X1 _u2_U780  ( .A1(mast0_dout[8]), .A2(_u2_n726 ), .ZN(_u2_n1370 ) );
NAND2_X1 _u2_U779  ( .A1(_u2_n728 ), .A2(_u2_adr0_cnt[6] ), .ZN(_u2_n1406 ));
NAND2_X1 _u2_U778  ( .A1(_u2_n1370 ), .A2(_u2_n1406 ), .ZN(de_adr0[8]) );
NAND2_X1 _u2_U777  ( .A1(mast0_dout[9]), .A2(_u2_n726 ), .ZN(_u2_n1367 ) );
NAND2_X1 _u2_U776  ( .A1(_u2_n729 ), .A2(_u2_adr0_cnt[7] ), .ZN(_u2_n1405 ));
NAND2_X1 _u2_U775  ( .A1(_u2_n1367 ), .A2(_u2_n1405 ), .ZN(de_adr0[9]) );
NAND2_X1 _u2_U774  ( .A1(_u2_n1564 ), .A2(_u2_state_6_ ), .ZN(_u2_n1404 ) );
NAND2_X1 _u2_U773  ( .A1(_u2_n719 ), .A2(_u2_n1404 ), .ZN(de_adr0_we) );
NAND2_X1 _u2_U772  ( .A1(_u2_n1369 ), .A2(_u2_adr1_cnt[8] ), .ZN(_u2_n1403 ));
NAND2_X1 _u2_U771  ( .A1(_u2_n1388 ), .A2(_u2_n1403 ), .ZN(de_adr1[10]) );
NAND2_X1 _u2_U770  ( .A1(_u2_n727 ), .A2(_u2_adr1_cnt[9] ), .ZN(_u2_n1402 ));
NAND2_X1 _u2_U769  ( .A1(_u2_n1386 ), .A2(_u2_n1402 ), .ZN(de_adr1[11]) );
MUX2_X1 _u2_U768  ( .A(mast0_dout[12]), .B(_u2_adr1_cnt[10] ), .S(_u2_n727 ),.Z(de_adr1[12]) );
MUX2_X1 _u2_U767  ( .A(mast0_dout[13]), .B(_u2_adr1_cnt[11] ), .S(_u2_n728 ),.Z(de_adr1[13]) );
MUX2_X1 _u2_U766  ( .A(mast0_dout[14]), .B(_u2_adr1_cnt[12] ), .S(_u2_n729 ),.Z(de_adr1[14]) );
MUX2_X1 _u2_U765  ( .A(mast0_dout[15]), .B(_u2_adr1_cnt[13] ), .S(_u2_n1369 ), .Z(de_adr1[15]) );
MUX2_X1 _u2_U764  ( .A(mast0_dout[16]), .B(_u2_adr1_cnt[14] ), .S(_u2_n727 ),.Z(de_adr1[16]) );
MUX2_X1 _u2_U763  ( .A(mast0_dout[17]), .B(_u2_adr1_cnt[15] ), .S(_u2_n728 ),.Z(de_adr1[17]) );
MUX2_X1 _u2_U762  ( .A(mast0_dout[18]), .B(_u2_adr1_cnt[16] ), .S(_u2_n729 ),.Z(de_adr1[18]) );
MUX2_X1 _u2_U761  ( .A(mast0_dout[19]), .B(_u2_adr1_cnt[17] ), .S(_u2_n1369 ), .Z(de_adr1[19]) );
MUX2_X1 _u2_U760  ( .A(mast0_dout[20]), .B(_u2_adr1_cnt[18] ), .S(_u2_n727 ),.Z(de_adr1[20]) );
MUX2_X1 _u2_U759  ( .A(mast0_dout[21]), .B(_u2_adr1_cnt[19] ), .S(_u2_n728 ),.Z(de_adr1[21]) );
MUX2_X1 _u2_U758  ( .A(mast0_dout[22]), .B(_u2_adr1_cnt[20] ), .S(_u2_n729 ),.Z(de_adr1[22]) );
MUX2_X1 _u2_U757  ( .A(mast0_dout[23]), .B(_u2_adr1_cnt[21] ), .S(_u2_n1369 ), .Z(de_adr1[23]) );
MUX2_X1 _u2_U756  ( .A(mast0_dout[24]), .B(_u2_adr1_cnt[22] ), .S(_u2_n727 ),.Z(de_adr1[24]) );
MUX2_X1 _u2_U755  ( .A(mast0_dout[25]), .B(_u2_adr1_cnt[23] ), .S(_u2_n728 ),.Z(de_adr1[25]) );
MUX2_X1 _u2_U754  ( .A(mast0_dout[26]), .B(_u2_adr1_cnt[24] ), .S(_u2_n729 ),.Z(de_adr1[26]) );
MUX2_X1 _u2_U753  ( .A(mast0_dout[27]), .B(_u2_adr1_cnt[25] ), .S(_u2_n1369 ), .Z(de_adr1[27]) );
MUX2_X1 _u2_U752  ( .A(mast0_dout[28]), .B(_u2_adr1_cnt[26] ), .S(_u2_n727 ),.Z(de_adr1[28]) );
MUX2_X1 _u2_U751  ( .A(mast0_dout[29]), .B(_u2_adr1_cnt[27] ), .S(_u2_n728 ),.Z(de_adr1[29]) );
NAND2_X1 _u2_U750  ( .A1(_u2_n728 ), .A2(_u2_adr1_cnt[0] ), .ZN(_u2_n1401 ));
NAND2_X1 _u2_U749  ( .A1(_u2_n1382 ), .A2(_u2_n1401 ), .ZN(de_adr1[2]) );
MUX2_X1 _u2_U748  ( .A(mast0_dout[30]), .B(_u2_adr1_cnt[28] ), .S(_u2_n729 ),.Z(de_adr1[30]) );
MUX2_X1 _u2_U747  ( .A(mast0_dout[31]), .B(_u2_adr1_cnt[29] ), .S(_u2_n1369 ), .Z(de_adr1[31]) );
NAND2_X1 _u2_U746  ( .A1(_u2_n729 ), .A2(_u2_adr1_cnt[1] ), .ZN(_u2_n1400 ));
NAND2_X1 _u2_U745  ( .A1(_u2_n1380 ), .A2(_u2_n1400 ), .ZN(de_adr1[3]) );
NAND2_X1 _u2_U744  ( .A1(_u2_n1369 ), .A2(_u2_adr1_cnt[2] ), .ZN(_u2_n1399 ));
NAND2_X1 _u2_U743  ( .A1(_u2_n1378 ), .A2(_u2_n1399 ), .ZN(de_adr1[4]) );
NAND2_X1 _u2_U742  ( .A1(_u2_n727 ), .A2(_u2_adr1_cnt[3] ), .ZN(_u2_n1398 ));
NAND2_X1 _u2_U741  ( .A1(_u2_n1376 ), .A2(_u2_n1398 ), .ZN(de_adr1[5]) );
NAND2_X1 _u2_U740  ( .A1(_u2_n728 ), .A2(_u2_adr1_cnt[4] ), .ZN(_u2_n1397 ));
NAND2_X1 _u2_U739  ( .A1(_u2_n1374 ), .A2(_u2_n1397 ), .ZN(de_adr1[6]) );
NAND2_X1 _u2_U738  ( .A1(_u2_n729 ), .A2(_u2_adr1_cnt[5] ), .ZN(_u2_n1396 ));
NAND2_X1 _u2_U737  ( .A1(_u2_n1372 ), .A2(_u2_n1396 ), .ZN(de_adr1[7]) );
NAND2_X1 _u2_U736  ( .A1(_u2_n1369 ), .A2(_u2_adr1_cnt[6] ), .ZN(_u2_n1395 ));
NAND2_X1 _u2_U735  ( .A1(_u2_n1370 ), .A2(_u2_n1395 ), .ZN(de_adr1[8]) );
NAND2_X1 _u2_U734  ( .A1(_u2_n727 ), .A2(_u2_adr1_cnt[7] ), .ZN(_u2_n1394 ));
NAND2_X1 _u2_U733  ( .A1(_u2_n1367 ), .A2(_u2_n1394 ), .ZN(de_adr1[9]) );
NAND2_X1 _u2_U732  ( .A1(_u2_n1564 ), .A2(_u2_state_7_ ), .ZN(_u2_n1393 ) );
NAND2_X1 _u2_U731  ( .A1(_u2_n719 ), .A2(_u2_n1393 ), .ZN(de_adr1_we) );
AND2_X1 _u2_U730  ( .A1(_u2_n1564 ), .A2(_u2_state_5_ ), .ZN(_u2_n1392 ) );
NOR2_X1 _u2_U729  ( .A1(_u2_state_4_ ), .A2(_u2_n1392 ), .ZN(_u2_n1366 ) );
INV_X1 _u2_U728  ( .A(_u2_n1366 ), .ZN(de_csr_we) );
NAND2_X1 _u2_U727  ( .A1(_u2_tsz_cnt[0] ), .A2(_u2_n729 ), .ZN(_u2_n1391 ));
NAND2_X1 _u2_U726  ( .A1(_u2_n1390 ), .A2(_u2_n1391 ), .ZN(de_txsz[0]) );
NAND2_X1 _u2_U725  ( .A1(_u2_tsz_cnt[10] ), .A2(_u2_n727 ), .ZN(_u2_n1389 ));
NAND2_X1 _u2_U724  ( .A1(_u2_n1388 ), .A2(_u2_n1389 ), .ZN(de_txsz[10]) );
NAND2_X1 _u2_U723  ( .A1(_u2_tsz_cnt[11] ), .A2(_u2_n728 ), .ZN(_u2_n1387 ));
NAND2_X1 _u2_U722  ( .A1(_u2_n1386 ), .A2(_u2_n1387 ), .ZN(de_txsz[11]) );
NAND2_X1 _u2_U721  ( .A1(_u2_tsz_cnt[1] ), .A2(_u2_n729 ), .ZN(_u2_n1385 ));
NAND2_X1 _u2_U720  ( .A1(_u2_n1384 ), .A2(_u2_n1385 ), .ZN(de_txsz[1]) );
NAND2_X1 _u2_U719  ( .A1(_u2_tsz_cnt[2] ), .A2(_u2_n729 ), .ZN(_u2_n1383 ));
NAND2_X1 _u2_U718  ( .A1(_u2_n1382 ), .A2(_u2_n1383 ), .ZN(de_txsz[2]) );
NAND2_X1 _u2_U717  ( .A1(_u2_tsz_cnt[3] ), .A2(_u2_n727 ), .ZN(_u2_n1381 ));
NAND2_X1 _u2_U716  ( .A1(_u2_n1380 ), .A2(_u2_n1381 ), .ZN(de_txsz[3]) );
NAND2_X1 _u2_U715  ( .A1(_u2_tsz_cnt[4] ), .A2(_u2_n728 ), .ZN(_u2_n1379 ));
NAND2_X1 _u2_U714  ( .A1(_u2_n1378 ), .A2(_u2_n1379 ), .ZN(de_txsz[4]) );
NAND2_X1 _u2_U713  ( .A1(_u2_tsz_cnt[5] ), .A2(_u2_n729 ), .ZN(_u2_n1377 ));
NAND2_X1 _u2_U712  ( .A1(_u2_n1376 ), .A2(_u2_n1377 ), .ZN(de_txsz[5]) );
NAND2_X1 _u2_U711  ( .A1(_u2_tsz_cnt[6] ), .A2(_u2_n728 ), .ZN(_u2_n1375 ));
NAND2_X1 _u2_U710  ( .A1(_u2_n1374 ), .A2(_u2_n1375 ), .ZN(de_txsz[6]) );
NAND2_X1 _u2_U709  ( .A1(_u2_tsz_cnt[7] ), .A2(_u2_n727 ), .ZN(_u2_n1373 ));
NAND2_X1 _u2_U708  ( .A1(_u2_n1372 ), .A2(_u2_n1373 ), .ZN(de_txsz[7]) );
NAND2_X1 _u2_U707  ( .A1(_u2_tsz_cnt[8] ), .A2(_u2_n728 ), .ZN(_u2_n1371 ));
NAND2_X1 _u2_U706  ( .A1(_u2_n1370 ), .A2(_u2_n1371 ), .ZN(de_txsz[8]) );
NAND2_X1 _u2_U705  ( .A1(_u2_tsz_cnt[9] ), .A2(_u2_n729 ), .ZN(_u2_n1368 ));
NAND2_X1 _u2_U704  ( .A1(_u2_n1367 ), .A2(_u2_n1368 ), .ZN(de_txsz[9]) );
NAND2_X1 _u2_U703  ( .A1(_u2_n1366 ), .A2(_u2_n719 ), .ZN(de_txsz_we) );
AND2_X1 _u2_U702  ( .A1(_u2_n1044 ), .A2(ndr), .ZN(_u2_n1365 ) );
NOR2_X1 _u2_U701  ( .A1(_u2_n1365 ), .A2(_u2_tsz_cnt_is_0_r ), .ZN(_u2_n1364 ) );
NOR2_X1 _u2_U700  ( .A1(_u2_n1364 ), .A2(_u2_n719 ), .ZN(dma_done_all) );
NAND2_X1 _u2_U699  ( .A1(_u2_n1290 ), .A2(mast1_dout[0]), .ZN(_u2_n1361 ) );
NAND2_X1 _u2_U698  ( .A1(_u2_n1289 ), .A2(mast0_dout[0]), .ZN(_u2_n1362 ) );
NAND2_X1 _u2_U697  ( .A1(_u2_tsz_cnt[0] ), .A2(_u2_n1288 ), .ZN(_u2_n1363 ));
NAND3_X1 _u2_U696  ( .A1(_u2_n1361 ), .A2(_u2_n1362 ), .A3(_u2_n1363 ), .ZN(mast0_din[0]) );
NAND2_X1 _u2_U695  ( .A1(_u2_n1290 ), .A2(mast1_dout[10]), .ZN(_u2_n1358 ));
NAND2_X1 _u2_U694  ( .A1(_u2_n1289 ), .A2(mast0_dout[10]), .ZN(_u2_n1359 ));
NAND2_X1 _u2_U693  ( .A1(_u2_tsz_cnt[10] ), .A2(_u2_n1288 ), .ZN(_u2_n1360 ));
NAND3_X1 _u2_U692  ( .A1(_u2_n1358 ), .A2(_u2_n1359 ), .A3(_u2_n1360 ), .ZN(mast0_din[10]) );
NAND2_X1 _u2_U691  ( .A1(_u2_n1290 ), .A2(mast1_dout[11]), .ZN(_u2_n1355 ));
NAND2_X1 _u2_U690  ( .A1(_u2_n1289 ), .A2(mast0_dout[11]), .ZN(_u2_n1356 ));
NAND2_X1 _u2_U689  ( .A1(_u2_tsz_cnt[11] ), .A2(_u2_n1288 ), .ZN(_u2_n1357 ));
NAND3_X1 _u2_U688  ( .A1(_u2_n1355 ), .A2(_u2_n1356 ), .A3(_u2_n1357 ), .ZN(mast0_din[11]) );
NAND2_X1 _u2_U687  ( .A1(_u2_n1290 ), .A2(mast1_dout[12]), .ZN(_u2_n1353 ));
NAND2_X1 _u2_U686  ( .A1(_u2_n1289 ), .A2(mast0_dout[12]), .ZN(_u2_n1354 ));
NAND2_X1 _u2_U685  ( .A1(_u2_n1353 ), .A2(_u2_n1354 ), .ZN(mast0_din[12]) );
NAND2_X1 _u2_U684  ( .A1(_u2_n1290 ), .A2(mast1_dout[13]), .ZN(_u2_n1351 ));
NAND2_X1 _u2_U683  ( .A1(_u2_n1289 ), .A2(mast0_dout[13]), .ZN(_u2_n1352 ));
NAND2_X1 _u2_U682  ( .A1(_u2_n1351 ), .A2(_u2_n1352 ), .ZN(mast0_din[13]) );
NAND2_X1 _u2_U681  ( .A1(_u2_n1290 ), .A2(mast1_dout[14]), .ZN(_u2_n1349 ));
NAND2_X1 _u2_U680  ( .A1(_u2_n1289 ), .A2(mast0_dout[14]), .ZN(_u2_n1350 ));
NAND2_X1 _u2_U679  ( .A1(_u2_n1349 ), .A2(_u2_n1350 ), .ZN(mast0_din[14]) );
NAND2_X1 _u2_U678  ( .A1(_u2_n1290 ), .A2(mast1_dout[15]), .ZN(_u2_n1347 ));
NAND2_X1 _u2_U677  ( .A1(_u2_n1289 ), .A2(mast0_dout[15]), .ZN(_u2_n1348 ));
NAND2_X1 _u2_U676  ( .A1(_u2_n1347 ), .A2(_u2_n1348 ), .ZN(mast0_din[15]) );
NAND2_X1 _u2_U675  ( .A1(_u2_n1290 ), .A2(mast1_dout[16]), .ZN(_u2_n1345 ));
NAND2_X1 _u2_U674  ( .A1(_u2_n1289 ), .A2(mast0_dout[16]), .ZN(_u2_n1346 ));
NAND2_X1 _u2_U673  ( .A1(_u2_n1345 ), .A2(_u2_n1346 ), .ZN(mast0_din[16]) );
NAND2_X1 _u2_U672  ( .A1(_u2_n1290 ), .A2(mast1_dout[17]), .ZN(_u2_n1343 ));
NAND2_X1 _u2_U671  ( .A1(_u2_n1289 ), .A2(mast0_dout[17]), .ZN(_u2_n1344 ));
NAND2_X1 _u2_U670  ( .A1(_u2_n1343 ), .A2(_u2_n1344 ), .ZN(mast0_din[17]) );
NAND2_X1 _u2_U669  ( .A1(_u2_n1290 ), .A2(mast1_dout[18]), .ZN(_u2_n1341 ));
NAND2_X1 _u2_U668  ( .A1(_u2_n1289 ), .A2(mast0_dout[18]), .ZN(_u2_n1342 ));
NAND2_X1 _u2_U667  ( .A1(_u2_n1341 ), .A2(_u2_n1342 ), .ZN(mast0_din[18]) );
NAND2_X1 _u2_U666  ( .A1(_u2_n1290 ), .A2(mast1_dout[19]), .ZN(_u2_n1339 ));
NAND2_X1 _u2_U665  ( .A1(_u2_n1289 ), .A2(mast0_dout[19]), .ZN(_u2_n1340 ));
NAND2_X1 _u2_U664  ( .A1(_u2_n1339 ), .A2(_u2_n1340 ), .ZN(mast0_din[19]) );
NAND2_X1 _u2_U663  ( .A1(_u2_n1290 ), .A2(mast1_dout[1]), .ZN(_u2_n1336 ) );
NAND2_X1 _u2_U662  ( .A1(_u2_n1289 ), .A2(mast0_dout[1]), .ZN(_u2_n1337 ) );
NAND2_X1 _u2_U661  ( .A1(_u2_tsz_cnt[1] ), .A2(_u2_n1288 ), .ZN(_u2_n1338 ));
NAND3_X1 _u2_U660  ( .A1(_u2_n1336 ), .A2(_u2_n1337 ), .A3(_u2_n1338 ), .ZN(mast0_din[1]) );
NAND2_X1 _u2_U659  ( .A1(_u2_n1290 ), .A2(mast1_dout[20]), .ZN(_u2_n1334 ));
NAND2_X1 _u2_U658  ( .A1(_u2_n1289 ), .A2(mast0_dout[20]), .ZN(_u2_n1335 ));
NAND2_X1 _u2_U657  ( .A1(_u2_n1334 ), .A2(_u2_n1335 ), .ZN(mast0_din[20]) );
NAND2_X1 _u2_U656  ( .A1(_u2_n1290 ), .A2(mast1_dout[21]), .ZN(_u2_n1332 ));
NAND2_X1 _u2_U655  ( .A1(_u2_n1289 ), .A2(mast0_dout[21]), .ZN(_u2_n1333 ));
NAND2_X1 _u2_U654  ( .A1(_u2_n1332 ), .A2(_u2_n1333 ), .ZN(mast0_din[21]) );
NAND2_X1 _u2_U653  ( .A1(_u2_n1290 ), .A2(mast1_dout[22]), .ZN(_u2_n1330 ));
NAND2_X1 _u2_U652  ( .A1(_u2_n1289 ), .A2(mast0_dout[22]), .ZN(_u2_n1331 ));
NAND2_X1 _u2_U651  ( .A1(_u2_n1330 ), .A2(_u2_n1331 ), .ZN(mast0_din[22]) );
NAND2_X1 _u2_U650  ( .A1(_u2_n1290 ), .A2(mast1_dout[23]), .ZN(_u2_n1328 ));
NAND2_X1 _u2_U649  ( .A1(_u2_n1289 ), .A2(mast0_dout[23]), .ZN(_u2_n1329 ));
NAND2_X1 _u2_U648  ( .A1(_u2_n1328 ), .A2(_u2_n1329 ), .ZN(mast0_din[23]) );
NAND2_X1 _u2_U647  ( .A1(_u2_n1290 ), .A2(mast1_dout[24]), .ZN(_u2_n1326 ));
NAND2_X1 _u2_U646  ( .A1(_u2_n1289 ), .A2(mast0_dout[24]), .ZN(_u2_n1327 ));
NAND2_X1 _u2_U645  ( .A1(_u2_n1326 ), .A2(_u2_n1327 ), .ZN(mast0_din[24]) );
NAND2_X1 _u2_U644  ( .A1(_u2_n1290 ), .A2(mast1_dout[25]), .ZN(_u2_n1324 ));
NAND2_X1 _u2_U643  ( .A1(_u2_n1289 ), .A2(mast0_dout[25]), .ZN(_u2_n1325 ));
NAND2_X1 _u2_U642  ( .A1(_u2_n1324 ), .A2(_u2_n1325 ), .ZN(mast0_din[25]) );
NAND2_X1 _u2_U641  ( .A1(_u2_n1290 ), .A2(mast1_dout[26]), .ZN(_u2_n1322 ));
NAND2_X1 _u2_U640  ( .A1(_u2_n1289 ), .A2(mast0_dout[26]), .ZN(_u2_n1323 ));
NAND2_X1 _u2_U639  ( .A1(_u2_n1322 ), .A2(_u2_n1323 ), .ZN(mast0_din[26]) );
NAND2_X1 _u2_U638  ( .A1(_u2_n1290 ), .A2(mast1_dout[27]), .ZN(_u2_n1320 ));
NAND2_X1 _u2_U637  ( .A1(_u2_n1289 ), .A2(mast0_dout[27]), .ZN(_u2_n1321 ));
NAND2_X1 _u2_U636  ( .A1(_u2_n1320 ), .A2(_u2_n1321 ), .ZN(mast0_din[27]) );
NAND2_X1 _u2_U635  ( .A1(_u2_n1290 ), .A2(mast1_dout[28]), .ZN(_u2_n1318 ));
NAND2_X1 _u2_U634  ( .A1(_u2_n1289 ), .A2(mast0_dout[28]), .ZN(_u2_n1319 ));
NAND2_X1 _u2_U633  ( .A1(_u2_n1318 ), .A2(_u2_n1319 ), .ZN(mast0_din[28]) );
NAND2_X1 _u2_U632  ( .A1(_u2_n1290 ), .A2(mast1_dout[29]), .ZN(_u2_n1316 ));
NAND2_X1 _u2_U631  ( .A1(_u2_n1289 ), .A2(mast0_dout[29]), .ZN(_u2_n1317 ));
NAND2_X1 _u2_U630  ( .A1(_u2_n1316 ), .A2(_u2_n1317 ), .ZN(mast0_din[29]) );
NAND2_X1 _u2_U629  ( .A1(_u2_n1290 ), .A2(mast1_dout[2]), .ZN(_u2_n1313 ) );
NAND2_X1 _u2_U628  ( .A1(_u2_n1289 ), .A2(mast0_dout[2]), .ZN(_u2_n1314 ) );
NAND2_X1 _u2_U627  ( .A1(_u2_tsz_cnt[2] ), .A2(_u2_n1288 ), .ZN(_u2_n1315 ));
NAND3_X1 _u2_U626  ( .A1(_u2_n1313 ), .A2(_u2_n1314 ), .A3(_u2_n1315 ), .ZN(mast0_din[2]) );
NAND2_X1 _u2_U625  ( .A1(_u2_n1290 ), .A2(mast1_dout[30]), .ZN(_u2_n1311 ));
NAND2_X1 _u2_U624  ( .A1(_u2_n1289 ), .A2(mast0_dout[30]), .ZN(_u2_n1312 ));
NAND2_X1 _u2_U623  ( .A1(_u2_n1311 ), .A2(_u2_n1312 ), .ZN(mast0_din[30]) );
NAND2_X1 _u2_U622  ( .A1(_u2_n1290 ), .A2(mast1_dout[31]), .ZN(_u2_n1309 ));
NAND2_X1 _u2_U621  ( .A1(_u2_n1289 ), .A2(mast0_dout[31]), .ZN(_u2_n1310 ));
NAND2_X1 _u2_U620  ( .A1(_u2_n1309 ), .A2(_u2_n1310 ), .ZN(mast0_din[31]) );
NAND2_X1 _u2_U619  ( .A1(_u2_n1290 ), .A2(mast1_dout[3]), .ZN(_u2_n1306 ) );
NAND2_X1 _u2_U618  ( .A1(_u2_n1289 ), .A2(mast0_dout[3]), .ZN(_u2_n1307 ) );
NAND2_X1 _u2_U617  ( .A1(_u2_tsz_cnt[3] ), .A2(_u2_n1288 ), .ZN(_u2_n1308 ));
NAND3_X1 _u2_U616  ( .A1(_u2_n1306 ), .A2(_u2_n1307 ), .A3(_u2_n1308 ), .ZN(mast0_din[3]) );
NAND2_X1 _u2_U615  ( .A1(_u2_n1290 ), .A2(mast1_dout[4]), .ZN(_u2_n1303 ) );
NAND2_X1 _u2_U614  ( .A1(_u2_n1289 ), .A2(mast0_dout[4]), .ZN(_u2_n1304 ) );
NAND2_X1 _u2_U613  ( .A1(_u2_tsz_cnt[4] ), .A2(_u2_n1288 ), .ZN(_u2_n1305 ));
NAND3_X1 _u2_U612  ( .A1(_u2_n1303 ), .A2(_u2_n1304 ), .A3(_u2_n1305 ), .ZN(mast0_din[4]) );
NAND2_X1 _u2_U611  ( .A1(_u2_n1290 ), .A2(mast1_dout[5]), .ZN(_u2_n1300 ) );
NAND2_X1 _u2_U610  ( .A1(_u2_n1289 ), .A2(mast0_dout[5]), .ZN(_u2_n1301 ) );
NAND2_X1 _u2_U609  ( .A1(_u2_tsz_cnt[5] ), .A2(_u2_n1288 ), .ZN(_u2_n1302 ));
NAND3_X1 _u2_U608  ( .A1(_u2_n1300 ), .A2(_u2_n1301 ), .A3(_u2_n1302 ), .ZN(mast0_din[5]) );
NAND2_X1 _u2_U607  ( .A1(_u2_n1290 ), .A2(mast1_dout[6]), .ZN(_u2_n1297 ) );
NAND2_X1 _u2_U606  ( .A1(_u2_n1289 ), .A2(mast0_dout[6]), .ZN(_u2_n1298 ) );
NAND2_X1 _u2_U605  ( .A1(_u2_tsz_cnt[6] ), .A2(_u2_n1288 ), .ZN(_u2_n1299 ));
NAND3_X1 _u2_U604  ( .A1(_u2_n1297 ), .A2(_u2_n1298 ), .A3(_u2_n1299 ), .ZN(mast0_din[6]) );
NAND2_X1 _u2_U603  ( .A1(_u2_n1290 ), .A2(mast1_dout[7]), .ZN(_u2_n1294 ) );
NAND2_X1 _u2_U602  ( .A1(_u2_n1289 ), .A2(mast0_dout[7]), .ZN(_u2_n1295 ) );
NAND2_X1 _u2_U601  ( .A1(_u2_tsz_cnt[7] ), .A2(_u2_n1288 ), .ZN(_u2_n1296 ));
NAND3_X1 _u2_U600  ( .A1(_u2_n1294 ), .A2(_u2_n1295 ), .A3(_u2_n1296 ), .ZN(mast0_din[7]) );
NAND2_X1 _u2_U599  ( .A1(_u2_n1290 ), .A2(mast1_dout[8]), .ZN(_u2_n1291 ) );
NAND2_X1 _u2_U598  ( .A1(_u2_n1289 ), .A2(mast0_dout[8]), .ZN(_u2_n1292 ) );
NAND2_X1 _u2_U597  ( .A1(_u2_tsz_cnt[8] ), .A2(_u2_n1288 ), .ZN(_u2_n1293 ));
NAND3_X1 _u2_U596  ( .A1(_u2_n1291 ), .A2(_u2_n1292 ), .A3(_u2_n1293 ), .ZN(mast0_din[8]) );
NAND2_X1 _u2_U595  ( .A1(_u2_n1290 ), .A2(mast1_dout[9]), .ZN(_u2_n1285 ) );
NAND2_X1 _u2_U594  ( .A1(_u2_n1289 ), .A2(mast0_dout[9]), .ZN(_u2_n1286 ) );
NAND2_X1 _u2_U593  ( .A1(_u2_tsz_cnt[9] ), .A2(_u2_n1288 ), .ZN(_u2_n1287 ));
NAND3_X1 _u2_U592  ( .A1(_u2_n1285 ), .A2(_u2_n1286 ), .A3(_u2_n1287 ), .ZN(mast0_din[9]) );
INV_X1 _u2_U591  ( .A(csr[1]), .ZN(_u2_n1271 ) );
NAND3_X1 _u2_U590  ( .A1(_u2_N342 ), .A2(_u2_n1271 ), .A3(_u2_write_hold_r ),.ZN(_u2_n1282 ) );
INV_X1 _u2_U589  ( .A(_u2_n1270 ), .ZN(_u2_n1566 ) );
NAND3_X1 _u2_U588  ( .A1(_u2_n1274 ), .A2(_u2_n1284 ), .A3(_u2_n1566 ), .ZN(_u2_n1283 ) );
NAND2_X1 _u2_U587  ( .A1(_u2_n1284 ), .A2(_u2_read ), .ZN(_u2_n1281 ) );
NAND4_X1 _u2_U586  ( .A1(_u2_n1282 ), .A2(_u2_n1283 ), .A3(_u2_n1281 ), .A4(_u2_n1278 ), .ZN(mast0_go) );
INV_X1 _u2_U585  ( .A(_u2_n1281 ), .ZN(_u2_n1279 ) );
NOR2_X1 _u2_U584  ( .A1(_u2_n1270 ), .A2(csr[1]), .ZN(_u2_n1277 ) );
NOR3_X1 _u2_U583  ( .A1(_u2_n1279 ), .A2(_u2_n1280 ), .A3(_u2_n1277 ), .ZN(mast0_wait) );
NAND2_X1 _u2_U582  ( .A1(_u2_n1277 ), .A2(_u2_n1278 ), .ZN(_u2_n1276 ) );
NAND2_X1 _u2_U581  ( .A1(_u2_n1275 ), .A2(_u2_n1276 ), .ZN(mast0_we) );
MUX2_X1 _u2_U580  ( .A(mast0_dout[0]), .B(mast1_dout[0]), .S(csr[2]), .Z(mast1_din[0]) );
MUX2_X1 _u2_U579  ( .A(mast0_dout[10]), .B(mast1_dout[10]), .S(csr[2]), .Z(mast1_din[10]) );
MUX2_X1 _u2_U578  ( .A(mast0_dout[11]), .B(mast1_dout[11]), .S(csr[2]), .Z(mast1_din[11]) );
MUX2_X1 _u2_U577  ( .A(mast0_dout[12]), .B(mast1_dout[12]), .S(csr[2]), .Z(mast1_din[12]) );
MUX2_X1 _u2_U576  ( .A(mast0_dout[13]), .B(mast1_dout[13]), .S(csr[2]), .Z(mast1_din[13]) );
MUX2_X1 _u2_U575  ( .A(mast0_dout[14]), .B(mast1_dout[14]), .S(csr[2]), .Z(mast1_din[14]) );
MUX2_X1 _u2_U574  ( .A(mast0_dout[15]), .B(mast1_dout[15]), .S(csr[2]), .Z(mast1_din[15]) );
MUX2_X1 _u2_U573  ( .A(mast0_dout[16]), .B(mast1_dout[16]), .S(csr[2]), .Z(mast1_din[16]) );
MUX2_X1 _u2_U572  ( .A(mast0_dout[17]), .B(mast1_dout[17]), .S(csr[2]), .Z(mast1_din[17]) );
MUX2_X1 _u2_U571  ( .A(mast0_dout[18]), .B(mast1_dout[18]), .S(csr[2]), .Z(mast1_din[18]) );
MUX2_X1 _u2_U570  ( .A(mast0_dout[19]), .B(mast1_dout[19]), .S(csr[2]), .Z(mast1_din[19]) );
MUX2_X1 _u2_U569  ( .A(mast0_dout[1]), .B(mast1_dout[1]), .S(csr[2]), .Z(mast1_din[1]) );
MUX2_X1 _u2_U568  ( .A(mast0_dout[20]), .B(mast1_dout[20]), .S(csr[2]), .Z(mast1_din[20]) );
MUX2_X1 _u2_U567  ( .A(mast0_dout[21]), .B(mast1_dout[21]), .S(csr[2]), .Z(mast1_din[21]) );
MUX2_X1 _u2_U566  ( .A(mast0_dout[22]), .B(mast1_dout[22]), .S(csr[2]), .Z(mast1_din[22]) );
MUX2_X1 _u2_U565  ( .A(mast0_dout[23]), .B(mast1_dout[23]), .S(csr[2]), .Z(mast1_din[23]) );
MUX2_X1 _u2_U564  ( .A(mast0_dout[24]), .B(mast1_dout[24]), .S(csr[2]), .Z(mast1_din[24]) );
MUX2_X1 _u2_U563  ( .A(mast0_dout[25]), .B(mast1_dout[25]), .S(csr[2]), .Z(mast1_din[25]) );
MUX2_X1 _u2_U562  ( .A(mast0_dout[26]), .B(mast1_dout[26]), .S(csr[2]), .Z(mast1_din[26]) );
MUX2_X1 _u2_U561  ( .A(mast0_dout[27]), .B(mast1_dout[27]), .S(csr[2]), .Z(mast1_din[27]) );
MUX2_X1 _u2_U560  ( .A(mast0_dout[28]), .B(mast1_dout[28]), .S(csr[2]), .Z(mast1_din[28]) );
MUX2_X1 _u2_U559  ( .A(mast0_dout[29]), .B(mast1_dout[29]), .S(csr[2]), .Z(mast1_din[29]) );
MUX2_X1 _u2_U558  ( .A(mast0_dout[2]), .B(mast1_dout[2]), .S(csr[2]), .Z(mast1_din[2]) );
MUX2_X1 _u2_U557  ( .A(mast0_dout[30]), .B(mast1_dout[30]), .S(csr[2]), .Z(mast1_din[30]) );
MUX2_X1 _u2_U556  ( .A(mast0_dout[31]), .B(mast1_dout[31]), .S(csr[2]), .Z(mast1_din[31]) );
MUX2_X1 _u2_U555  ( .A(mast0_dout[3]), .B(mast1_dout[3]), .S(csr[2]), .Z(mast1_din[3]) );
MUX2_X1 _u2_U554  ( .A(mast0_dout[4]), .B(mast1_dout[4]), .S(csr[2]), .Z(mast1_din[4]) );
MUX2_X1 _u2_U553  ( .A(mast0_dout[5]), .B(mast1_dout[5]), .S(csr[2]), .Z(mast1_din[5]) );
MUX2_X1 _u2_U552  ( .A(mast0_dout[6]), .B(mast1_dout[6]), .S(csr[2]), .Z(mast1_din[6]) );
MUX2_X1 _u2_U551  ( .A(mast0_dout[7]), .B(mast1_dout[7]), .S(csr[2]), .Z(mast1_din[7]) );
MUX2_X1 _u2_U550  ( .A(mast0_dout[8]), .B(mast1_dout[8]), .S(csr[2]), .Z(mast1_din[8]) );
MUX2_X1 _u2_U549  ( .A(mast0_dout[9]), .B(mast1_dout[9]), .S(csr[2]), .Z(mast1_din[9]) );
NAND3_X1 _u2_U548  ( .A1(csr[2]), .A2(_u2_n1274 ), .A3(_u2_n1566 ), .ZN(_u2_n1272 ) );
NAND2_X1 _u2_U547  ( .A1(csr[2]), .A2(_u2_read ), .ZN(_u2_n1269 ) );
NAND3_X1 _u2_U546  ( .A1(csr[1]), .A2(_u2_N342 ), .A3(_u2_write_hold_r ),.ZN(_u2_n1273 ) );
NAND3_X1 _u2_U545  ( .A1(_u2_n1272 ), .A2(_u2_n1269 ), .A3(_u2_n1273 ), .ZN(mast1_go) );
NOR2_X1 _u2_U544  ( .A1(_u2_n1270 ), .A2(_u2_n1271 ), .ZN(mast1_we) );
INV_X1 _u2_U543  ( .A(_u2_n1269 ), .ZN(_u2_n1268 ) );
NOR2_X1 _u2_U542  ( .A1(mast1_we), .A2(_u2_n1268 ), .ZN(mast1_wait) );
INV_X1 _u2_U541  ( .A(de_start), .ZN(_u2_n1230 ) );
NAND2_X1 _u2_U540  ( .A1(_u2_n720 ), .A2(_u2_n1230 ), .ZN(_u2_n892 ) );
INV_X1 _u2_U539  ( .A(_u2_n892 ), .ZN(_u2_n1245 ) );
NOR2_X1 _u2_U538  ( .A1(_u2_n892 ), .A2(_u2_n770 ), .ZN(_u2_n893 ) );
OR2_X1 _u2_U537  ( .A1(_u2_n769 ), .A2(am0[28]), .ZN(_u2_n1266 ) );
NAND2_X1 _u2_U536  ( .A1(_u2_n772 ), .A2(_u2_n1266 ), .ZN(_u2_n1265 ) );
NAND2_X1 _u2_U535  ( .A1(_u2_adr0_cnt[26] ), .A2(_u2_n1265 ), .ZN(_u2_n1262 ) );
NAND3_X1 _u2_U534  ( .A1(_u2_adr0_cnt_next1[26]), .A2(_u2_n770 ), .A3(am0[28]), .ZN(_u2_n1263 ) );
NAND2_X1 _u2_U533  ( .A1(adr0[28]), .A2(_u2_n769 ), .ZN(_u2_n1264 ) );
NAND3_X1 _u2_U532  ( .A1(_u2_n1262 ), .A2(_u2_n1263 ), .A3(_u2_n1264 ), .ZN(_u2_n1000 ) );
OR2_X1 _u2_U531  ( .A1(_u2_n769 ), .A2(am0[29]), .ZN(_u2_n1261 ) );
NAND2_X1 _u2_U530  ( .A1(_u2_n772 ), .A2(_u2_n1261 ), .ZN(_u2_n1260 ) );
NAND2_X1 _u2_U529  ( .A1(_u2_adr0_cnt[27] ), .A2(_u2_n1260 ), .ZN(_u2_n1257 ) );
NAND3_X1 _u2_U528  ( .A1(_u2_adr0_cnt_next1[27]), .A2(_u2_n770 ), .A3(am0[29]), .ZN(_u2_n1258 ) );
NAND2_X1 _u2_U527  ( .A1(adr0[29]), .A2(_u2_n769 ), .ZN(_u2_n1259 ) );
NAND3_X1 _u2_U526  ( .A1(_u2_n1257 ), .A2(_u2_n1258 ), .A3(_u2_n1259 ), .ZN(_u2_n1001 ) );
OR2_X1 _u2_U525  ( .A1(_u2_n769 ), .A2(am0[30]), .ZN(_u2_n1256 ) );
NAND2_X1 _u2_U524  ( .A1(_u2_n772 ), .A2(_u2_n1256 ), .ZN(_u2_n1255 ) );
NAND2_X1 _u2_U523  ( .A1(_u2_adr0_cnt[28] ), .A2(_u2_n1255 ), .ZN(_u2_n1252 ) );
NAND3_X1 _u2_U522  ( .A1(_u2_adr0_cnt_next1[28]), .A2(_u2_n770 ), .A3(am0[30]), .ZN(_u2_n1253 ) );
NAND2_X1 _u2_U521  ( .A1(adr0[30]), .A2(_u2_n769 ), .ZN(_u2_n1254 ) );
NAND3_X1 _u2_U520  ( .A1(_u2_n1252 ), .A2(_u2_n1253 ), .A3(_u2_n1254 ), .ZN(_u2_n1002 ) );
OR2_X1 _u2_U519  ( .A1(_u2_n769 ), .A2(am0[31]), .ZN(_u2_n1251 ) );
NAND2_X1 _u2_U518  ( .A1(_u2_n772 ), .A2(_u2_n1251 ), .ZN(_u2_n1250 ) );
NAND2_X1 _u2_U517  ( .A1(_u2_adr0_cnt[29] ), .A2(_u2_n1250 ), .ZN(_u2_n1247 ) );
NAND3_X1 _u2_U516  ( .A1(_u2_adr0_cnt_next1[29]), .A2(_u2_n770 ), .A3(am0[31]), .ZN(_u2_n1248 ) );
NAND2_X1 _u2_U515  ( .A1(adr0[31]), .A2(_u2_n769 ), .ZN(_u2_n1249 ) );
NAND3_X1 _u2_U514  ( .A1(_u2_n1247 ), .A2(_u2_n1248 ), .A3(_u2_n1249 ), .ZN(_u2_n1003 ) );
NOR2_X1 _u2_U513  ( .A1(_u2_n892 ), .A2(_u2_n901 ), .ZN(_u2_n1138 ) );
OR2_X1 _u2_U512  ( .A1(_u2_n900 ), .A2(am1[31]), .ZN(_u2_n1244 ) );
NAND2_X1 _u2_U511  ( .A1(_u2_n903 ), .A2(_u2_n1244 ), .ZN(_u2_n1243 ) );
NAND2_X1 _u2_U510  ( .A1(_u2_adr1_cnt[29] ), .A2(_u2_n1243 ), .ZN(_u2_n1240 ) );
NAND3_X1 _u2_U509  ( .A1(_u2_adr1_cnt_next1[29]), .A2(_u2_n901 ), .A3(am1[31]), .ZN(_u2_n1241 ) );
NAND2_X1 _u2_U508  ( .A1(adr1[31]), .A2(_u2_n900 ), .ZN(_u2_n1242 ) );
NAND3_X1 _u2_U507  ( .A1(_u2_n1240 ), .A2(_u2_n1241 ), .A3(_u2_n1242 ), .ZN(_u2_n1004 ) );
NOR2_X1 _u2_U506  ( .A1(dma_err), .A2(_u2_n722 ), .ZN(_u2_n1231 ) );
NOR2_X1 _u2_U505  ( .A1(dma_err), .A2(_u2_n1239 ), .ZN(_u2_n1232 ) );
NOR2_X1 _u2_U504  ( .A1(csr[12]), .A2(_u2_n1230 ), .ZN(_u2_n1238 ) );
NOR2_X1 _u2_U503  ( .A1(_u2_n1238 ), .A2(_u2_n721 ), .ZN(_u2_n1237 ) );
MUX2_X1 _u2_U502  ( .A(_u2_n1237 ), .B(paused), .S(pause_req), .Z(_u2_n1233 ) );
NOR2_X1 _u2_U501  ( .A1(_u2_state_9_ ), .A2(_u2_n726 ), .ZN(_u2_n1236 ) );
NOR2_X1 _u2_U500  ( .A1(mast0_drdy), .A2(_u2_n1236 ), .ZN(_u2_n1235 ) );
NOR4_X1 _u2_U499  ( .A1(_u2_n1232 ), .A2(_u2_n1233 ), .A3(_u2_n1234 ), .A4(_u2_n1235 ), .ZN(_u2_n1145 ) );
MUX2_X1 _u2_U498  ( .A(_u2_state_2_ ), .B(_u2_n1231 ), .S(_u2_n1145 ), .Z(_u2_n1011 ) );
AND3_X1 _u2_U497  ( .A1(_u2_chunk_dec ), .A2(_u2_n934 ), .A3(_u2_n1230 ),.ZN(_u2_n1205 ) );
NAND2_X1 _u2_U496  ( .A1(_u2_N188 ), .A2(_u2_n1205 ), .ZN(_u2_n1227 ) );
NOR2_X1 _u2_U495  ( .A1(_u2_n1205 ), .A2(de_start), .ZN(_u2_n1204 ) );
NAND2_X1 _u2_U494  ( .A1(_u2_n1204 ), .A2(_u2_chunk_cnt[8] ), .ZN(_u2_n1228 ) );
NAND2_X1 _u2_U493  ( .A1(txsz[24]), .A2(de_start), .ZN(_u2_n1229 ) );
NAND3_X1 _u2_U492  ( .A1(_u2_n1227 ), .A2(_u2_n1228 ), .A3(_u2_n1229 ), .ZN(_u2_n1012 ) );
NAND2_X1 _u2_U491  ( .A1(_u2_N187 ), .A2(_u2_n1205 ), .ZN(_u2_n1224 ) );
NAND2_X1 _u2_U490  ( .A1(_u2_n1204 ), .A2(_u2_chunk_cnt[7] ), .ZN(_u2_n1225 ) );
NAND2_X1 _u2_U489  ( .A1(txsz[23]), .A2(de_start), .ZN(_u2_n1226 ) );
NAND3_X1 _u2_U488  ( .A1(_u2_n1224 ), .A2(_u2_n1225 ), .A3(_u2_n1226 ), .ZN(_u2_n1013 ) );
NAND2_X1 _u2_U487  ( .A1(_u2_N186 ), .A2(_u2_n1205 ), .ZN(_u2_n1221 ) );
NAND2_X1 _u2_U486  ( .A1(_u2_n1204 ), .A2(_u2_chunk_cnt[6] ), .ZN(_u2_n1222 ) );
NAND2_X1 _u2_U485  ( .A1(txsz[22]), .A2(de_start), .ZN(_u2_n1223 ) );
NAND3_X1 _u2_U484  ( .A1(_u2_n1221 ), .A2(_u2_n1222 ), .A3(_u2_n1223 ), .ZN(_u2_n1014 ) );
NAND2_X1 _u2_U483  ( .A1(_u2_N185 ), .A2(_u2_n1205 ), .ZN(_u2_n1218 ) );
NAND2_X1 _u2_U482  ( .A1(_u2_n1204 ), .A2(_u2_chunk_cnt[5] ), .ZN(_u2_n1219 ) );
NAND2_X1 _u2_U481  ( .A1(txsz[21]), .A2(de_start), .ZN(_u2_n1220 ) );
NAND3_X1 _u2_U480  ( .A1(_u2_n1218 ), .A2(_u2_n1219 ), .A3(_u2_n1220 ), .ZN(_u2_n1015 ) );
NAND2_X1 _u2_U479  ( .A1(_u2_N184 ), .A2(_u2_n1205 ), .ZN(_u2_n1215 ) );
NAND2_X1 _u2_U478  ( .A1(_u2_n1204 ), .A2(_u2_chunk_cnt[4] ), .ZN(_u2_n1216 ) );
NAND2_X1 _u2_U477  ( .A1(txsz[20]), .A2(de_start), .ZN(_u2_n1217 ) );
NAND3_X1 _u2_U476  ( .A1(_u2_n1215 ), .A2(_u2_n1216 ), .A3(_u2_n1217 ), .ZN(_u2_n1016 ) );
NAND2_X1 _u2_U475  ( .A1(_u2_N183 ), .A2(_u2_n1205 ), .ZN(_u2_n1212 ) );
NAND2_X1 _u2_U474  ( .A1(_u2_n1204 ), .A2(_u2_chunk_cnt[3] ), .ZN(_u2_n1213 ) );
NAND2_X1 _u2_U473  ( .A1(txsz[19]), .A2(de_start), .ZN(_u2_n1214 ) );
NAND3_X1 _u2_U472  ( .A1(_u2_n1212 ), .A2(_u2_n1213 ), .A3(_u2_n1214 ), .ZN(_u2_n1017 ) );
NAND2_X1 _u2_U471  ( .A1(_u2_N182 ), .A2(_u2_n1205 ), .ZN(_u2_n1209 ) );
NAND2_X1 _u2_U470  ( .A1(_u2_n1204 ), .A2(_u2_chunk_cnt[2] ), .ZN(_u2_n1210 ) );
NAND2_X1 _u2_U469  ( .A1(txsz[18]), .A2(de_start), .ZN(_u2_n1211 ) );
NAND3_X1 _u2_U468  ( .A1(_u2_n1209 ), .A2(_u2_n1210 ), .A3(_u2_n1211 ), .ZN(_u2_n1018 ) );
NAND2_X1 _u2_U467  ( .A1(_u2_N181 ), .A2(_u2_n1205 ), .ZN(_u2_n1206 ) );
NAND2_X1 _u2_U466  ( .A1(_u2_n1204 ), .A2(_u2_chunk_cnt[1] ), .ZN(_u2_n1207 ) );
NAND2_X1 _u2_U465  ( .A1(txsz[17]), .A2(de_start), .ZN(_u2_n1208 ) );
NAND3_X1 _u2_U464  ( .A1(_u2_n1206 ), .A2(_u2_n1207 ), .A3(_u2_n1208 ), .ZN(_u2_n1019 ) );
NAND2_X1 _u2_U463  ( .A1(_u2_N180 ), .A2(_u2_n1205 ), .ZN(_u2_n1201 ) );
NAND2_X1 _u2_U462  ( .A1(_u2_n1204 ), .A2(_u2_chunk_cnt[0] ), .ZN(_u2_n1202 ) );
NAND2_X1 _u2_U461  ( .A1(txsz[16]), .A2(de_start), .ZN(_u2_n1203 ) );
NAND3_X1 _u2_U460  ( .A1(_u2_n1201 ), .A2(_u2_n1202 ), .A3(_u2_n1203 ), .ZN(_u2_n1020 ) );
NOR3_X1 _u2_U459  ( .A1(_u2_n725 ), .A2(_u2_tsz_cnt_is_0_r ), .A3(_u2_n892 ),.ZN(_u2_n1160 ) );
NAND2_X1 _u2_U458  ( .A1(_u2_N204 ), .A2(_u2_n1160 ), .ZN(_u2_n1198 ) );
NOR2_X1 _u2_U457  ( .A1(_u2_n892 ), .A2(_u2_n1160 ), .ZN(_u2_n1159 ) );
NAND2_X1 _u2_U456  ( .A1(_u2_tsz_cnt[0] ), .A2(_u2_n1159 ), .ZN(_u2_n1199 ));
NAND2_X1 _u2_U455  ( .A1(txsz[0]), .A2(_u2_n892 ), .ZN(_u2_n1200 ) );
NAND3_X1 _u2_U454  ( .A1(_u2_n1198 ), .A2(_u2_n1199 ), .A3(_u2_n1200 ), .ZN(_u2_n1021 ) );
NAND2_X1 _u2_U453  ( .A1(_u2_N205 ), .A2(_u2_n1160 ), .ZN(_u2_n1195 ) );
NAND2_X1 _u2_U452  ( .A1(_u2_tsz_cnt[1] ), .A2(_u2_n1159 ), .ZN(_u2_n1196 ));
NAND2_X1 _u2_U451  ( .A1(txsz[1]), .A2(_u2_n892 ), .ZN(_u2_n1197 ) );
NAND3_X1 _u2_U450  ( .A1(_u2_n1195 ), .A2(_u2_n1196 ), .A3(_u2_n1197 ), .ZN(_u2_n1022 ) );
NAND2_X1 _u2_U449  ( .A1(_u2_N206 ), .A2(_u2_n1160 ), .ZN(_u2_n1192 ) );
NAND2_X1 _u2_U448  ( .A1(_u2_tsz_cnt[2] ), .A2(_u2_n1159 ), .ZN(_u2_n1193 ));
NAND2_X1 _u2_U447  ( .A1(txsz[2]), .A2(_u2_n892 ), .ZN(_u2_n1194 ) );
NAND3_X1 _u2_U446  ( .A1(_u2_n1192 ), .A2(_u2_n1193 ), .A3(_u2_n1194 ), .ZN(_u2_n1023 ) );
NAND2_X1 _u2_U445  ( .A1(_u2_N207 ), .A2(_u2_n1160 ), .ZN(_u2_n1189 ) );
NAND2_X1 _u2_U444  ( .A1(_u2_tsz_cnt[3] ), .A2(_u2_n1159 ), .ZN(_u2_n1190 ));
NAND2_X1 _u2_U443  ( .A1(txsz[3]), .A2(_u2_n892 ), .ZN(_u2_n1191 ) );
NAND3_X1 _u2_U442  ( .A1(_u2_n1189 ), .A2(_u2_n1190 ), .A3(_u2_n1191 ), .ZN(_u2_n1024 ) );
NAND2_X1 _u2_U441  ( .A1(_u2_N208 ), .A2(_u2_n1160 ), .ZN(_u2_n1186 ) );
NAND2_X1 _u2_U440  ( .A1(_u2_tsz_cnt[4] ), .A2(_u2_n1159 ), .ZN(_u2_n1187 ));
NAND2_X1 _u2_U439  ( .A1(txsz[4]), .A2(_u2_n892 ), .ZN(_u2_n1188 ) );
NAND3_X1 _u2_U438  ( .A1(_u2_n1186 ), .A2(_u2_n1187 ), .A3(_u2_n1188 ), .ZN(_u2_n1025 ) );
NAND2_X1 _u2_U437  ( .A1(_u2_N209 ), .A2(_u2_n1160 ), .ZN(_u2_n1183 ) );
NAND2_X1 _u2_U436  ( .A1(_u2_tsz_cnt[5] ), .A2(_u2_n1159 ), .ZN(_u2_n1184 ));
NAND2_X1 _u2_U435  ( .A1(txsz[5]), .A2(_u2_n892 ), .ZN(_u2_n1185 ) );
NAND3_X1 _u2_U434  ( .A1(_u2_n1183 ), .A2(_u2_n1184 ), .A3(_u2_n1185 ), .ZN(_u2_n1026 ) );
NAND2_X1 _u2_U433  ( .A1(_u2_N210 ), .A2(_u2_n1160 ), .ZN(_u2_n1180 ) );
NAND2_X1 _u2_U432  ( .A1(_u2_tsz_cnt[6] ), .A2(_u2_n1159 ), .ZN(_u2_n1181 ));
NAND2_X1 _u2_U431  ( .A1(txsz[6]), .A2(_u2_n892 ), .ZN(_u2_n1182 ) );
NAND3_X1 _u2_U430  ( .A1(_u2_n1180 ), .A2(_u2_n1181 ), .A3(_u2_n1182 ), .ZN(_u2_n1027 ) );
NAND2_X1 _u2_U429  ( .A1(_u2_N211 ), .A2(_u2_n1160 ), .ZN(_u2_n1177 ) );
NAND2_X1 _u2_U428  ( .A1(_u2_tsz_cnt[7] ), .A2(_u2_n1159 ), .ZN(_u2_n1178 ));
NAND2_X1 _u2_U427  ( .A1(txsz[7]), .A2(_u2_n892 ), .ZN(_u2_n1179 ) );
NAND3_X1 _u2_U426  ( .A1(_u2_n1177 ), .A2(_u2_n1178 ), .A3(_u2_n1179 ), .ZN(_u2_n1028 ) );
NAND2_X1 _u2_U425  ( .A1(_u2_N212 ), .A2(_u2_n1160 ), .ZN(_u2_n1174 ) );
NAND2_X1 _u2_U424  ( .A1(_u2_tsz_cnt[8] ), .A2(_u2_n1159 ), .ZN(_u2_n1175 ));
NAND2_X1 _u2_U423  ( .A1(txsz[8]), .A2(_u2_n892 ), .ZN(_u2_n1176 ) );
NAND3_X1 _u2_U422  ( .A1(_u2_n1174 ), .A2(_u2_n1175 ), .A3(_u2_n1176 ), .ZN(_u2_n1029 ) );
NAND2_X1 _u2_U421  ( .A1(_u2_N213 ), .A2(_u2_n1160 ), .ZN(_u2_n1171 ) );
NAND2_X1 _u2_U420  ( .A1(_u2_tsz_cnt[9] ), .A2(_u2_n1159 ), .ZN(_u2_n1172 ));
NAND2_X1 _u2_U419  ( .A1(txsz[9]), .A2(_u2_n892 ), .ZN(_u2_n1173 ) );
NAND3_X1 _u2_U418  ( .A1(_u2_n1171 ), .A2(_u2_n1172 ), .A3(_u2_n1173 ), .ZN(_u2_n1030 ) );
NAND2_X1 _u2_U417  ( .A1(_u2_N214 ), .A2(_u2_n1160 ), .ZN(_u2_n1168 ) );
NAND2_X1 _u2_U416  ( .A1(_u2_tsz_cnt[10] ), .A2(_u2_n1159 ), .ZN(_u2_n1169 ));
NAND2_X1 _u2_U415  ( .A1(txsz[10]), .A2(_u2_n892 ), .ZN(_u2_n1170 ) );
NAND3_X1 _u2_U414  ( .A1(_u2_n1168 ), .A2(_u2_n1169 ), .A3(_u2_n1170 ), .ZN(_u2_n1031 ) );
MUX2_X1 _u2_U413  ( .A(ptr_set), .B(_u2_state_7_ ), .S(_u2_n1145 ), .Z(_u2_n1032 ) );
MUX2_X1 _u2_U412  ( .A(_u2_state_7_ ), .B(_u2_state_6_ ), .S(_u2_n1145 ),.Z(_u2_n1033 ) );
MUX2_X1 _u2_U411  ( .A(_u2_state_6_ ), .B(_u2_state_5_ ), .S(_u2_n1145 ),.Z(_u2_n1034 ) );
MUX2_X1 _u2_U410  ( .A(_u2_state_5_ ), .B(_u2_state_4_ ), .S(_u2_n1145 ),.Z(_u2_n1035 ) );
INV_X1 _u2_U409  ( .A(pointer[0]), .ZN(_u2_n1167 ) );
NAND2_X1 _u2_U408  ( .A1(_u2_n1167 ), .A2(csr[7]), .ZN(_u2_n1155 ) );
NOR3_X1 _u2_U407  ( .A1(_u2_n1155 ), .A2(pause_req), .A3(_u2_n721 ), .ZN(_u2_n1166 ) );
MUX2_X1 _u2_U406  ( .A(_u2_state_4_ ), .B(_u2_n1166 ), .S(_u2_n1145 ), .Z(_u2_n1036 ) );
NAND2_X1 _u2_U405  ( .A1(_u2_state_2_ ), .A2(_u2_n1165 ), .ZN(_u2_n1162 ) );
NAND2_X1 _u2_U404  ( .A1(_u2_n1164 ), .A2(dma_err), .ZN(_u2_n1163 ) );
NAND2_X1 _u2_U403  ( .A1(_u2_n1162 ), .A2(_u2_n1163 ), .ZN(_u2_n1161 ) );
MUX2_X1 _u2_U402  ( .A(_u2_state_3_ ), .B(_u2_n1161 ), .S(_u2_n1145 ), .Z(_u2_n1037 ) );
NAND2_X1 _u2_U401  ( .A1(_u2_N215 ), .A2(_u2_n1160 ), .ZN(_u2_n1156 ) );
NAND2_X1 _u2_U400  ( .A1(_u2_tsz_cnt[11] ), .A2(_u2_n1159 ), .ZN(_u2_n1157 ));
NAND2_X1 _u2_U399  ( .A1(txsz[11]), .A2(_u2_n892 ), .ZN(_u2_n1158 ) );
NAND3_X1 _u2_U398  ( .A1(_u2_n1156 ), .A2(_u2_n1157 ), .A3(_u2_n1158 ), .ZN(_u2_n1038 ) );
INV_X1 _u2_U397  ( .A(pause_req), .ZN(_u2_n1150 ) );
NAND3_X1 _u2_U396  ( .A1(_u2_n1155 ), .A2(_u2_n1150 ), .A3(_u2_state_0_ ),.ZN(_u2_n1154 ) );
NAND3_X1 _u2_U395  ( .A1(_u2_n1153 ), .A2(_u2_n720 ), .A3(_u2_n1154 ), .ZN(_u2_n1152 ) );
MUX2_X1 _u2_U394  ( .A(_u2_state_1_ ), .B(_u2_n1152 ), .S(_u2_n1145 ), .Z(_u2_n1039 ) );
MUX2_X1 _u2_U393  ( .A(_u2_state_9_ ), .B(_u2_n1151 ), .S(_u2_n1145 ), .Z(_u2_n1040 ) );
NOR2_X1 _u2_U392  ( .A1(_u2_n1150 ), .A2(_u2_n721 ), .ZN(_u2_n1149 ) );
MUX2_X1 _u2_U391  ( .A(paused), .B(_u2_n1149 ), .S(_u2_n1145 ), .Z(_u2_n1041 ) );
NAND2_X1 _u2_U390  ( .A1(_u2_state_3_ ), .A2(_u2_n1148 ), .ZN(_u2_n1147 ) );
NAND2_X1 _u2_U389  ( .A1(_u2_n1146 ), .A2(_u2_n1147 ), .ZN(_u2_n1144 ) );
MUX2_X1 _u2_U388  ( .A(_u2_state_0_ ), .B(_u2_n1144 ), .S(_u2_n1145 ), .Z(_u2_n1042 ) );
OR4_X1 _u2_U387  ( .A1(txsz[16]), .A2(txsz[17]), .A3(txsz[18]), .A4(txsz[19]), .ZN(_u2_n1142 ) );
OR3_X1 _u2_U386  ( .A1(txsz[23]), .A2(txsz[24]), .A3(txsz[22]), .ZN(_u2_n1143 ) );
NOR4_X1 _u2_U385  ( .A1(_u2_n1142 ), .A2(_u2_n1143 ), .A3(txsz[21]), .A4(txsz[20]), .ZN(_u2_n1045 ) );
NAND2_X1 _u2_U384  ( .A1(_u2_adr1_cnt_next1[0]), .A2(_u2_n901 ), .ZN(_u2_n1139 ) );
NAND2_X1 _u2_U383  ( .A1(_u2_adr1_cnt[0] ), .A2(_u2_n1138 ), .ZN(_u2_n1140 ));
NAND2_X1 _u2_U382  ( .A1(adr1[2]), .A2(_u2_n892 ), .ZN(_u2_n1141 ) );
NAND3_X1 _u2_U381  ( .A1(_u2_n1139 ), .A2(_u2_n1140 ), .A3(_u2_n1141 ), .ZN(_u2_n945 ) );
NAND2_X1 _u2_U380  ( .A1(_u2_adr1_cnt_next1[1]), .A2(_u2_n901 ), .ZN(_u2_n1135 ) );
NAND2_X1 _u2_U379  ( .A1(_u2_adr1_cnt[1] ), .A2(_u2_n1138 ), .ZN(_u2_n1136 ));
NAND2_X1 _u2_U378  ( .A1(adr1[3]), .A2(_u2_n892 ), .ZN(_u2_n1137 ) );
NAND3_X1 _u2_U377  ( .A1(_u2_n1135 ), .A2(_u2_n1136 ), .A3(_u2_n1137 ), .ZN(_u2_n946 ) );
OR2_X1 _u2_U376  ( .A1(_u2_n900 ), .A2(am1[4]), .ZN(_u2_n1134 ) );
NAND2_X1 _u2_U375  ( .A1(_u2_n903 ), .A2(_u2_n1134 ), .ZN(_u2_n1133 ) );
NAND2_X1 _u2_U374  ( .A1(_u2_adr1_cnt[2] ), .A2(_u2_n1133 ), .ZN(_u2_n1130 ));
NAND3_X1 _u2_U373  ( .A1(_u2_adr1_cnt_next1[2]), .A2(_u2_n901 ), .A3(am1[4]), .ZN(_u2_n1131 ) );
NAND2_X1 _u2_U372  ( .A1(adr1[4]), .A2(_u2_n900 ), .ZN(_u2_n1132 ) );
NAND3_X1 _u2_U371  ( .A1(_u2_n1130 ), .A2(_u2_n1131 ), .A3(_u2_n1132 ), .ZN(_u2_n947 ) );
OR2_X1 _u2_U370  ( .A1(_u2_n900 ), .A2(am1[5]), .ZN(_u2_n1129 ) );
NAND2_X1 _u2_U369  ( .A1(_u2_n903 ), .A2(_u2_n1129 ), .ZN(_u2_n1128 ) );
NAND2_X1 _u2_U368  ( .A1(_u2_adr1_cnt[3] ), .A2(_u2_n1128 ), .ZN(_u2_n1125 ));
NAND3_X1 _u2_U367  ( .A1(_u2_adr1_cnt_next1[3]), .A2(_u2_n901 ), .A3(am1[5]), .ZN(_u2_n1126 ) );
NAND2_X1 _u2_U366  ( .A1(adr1[5]), .A2(_u2_n900 ), .ZN(_u2_n1127 ) );
NAND3_X1 _u2_U365  ( .A1(_u2_n1125 ), .A2(_u2_n1126 ), .A3(_u2_n1127 ), .ZN(_u2_n948 ) );
OR2_X1 _u2_U364  ( .A1(_u2_n900 ), .A2(am1[6]), .ZN(_u2_n1124 ) );
NAND2_X1 _u2_U363  ( .A1(_u2_n903 ), .A2(_u2_n1124 ), .ZN(_u2_n1123 ) );
NAND2_X1 _u2_U362  ( .A1(_u2_adr1_cnt[4] ), .A2(_u2_n1123 ), .ZN(_u2_n1120 ));
NAND3_X1 _u2_U361  ( .A1(_u2_adr1_cnt_next1[4]), .A2(_u2_n901 ), .A3(am1[6]), .ZN(_u2_n1121 ) );
NAND2_X1 _u2_U360  ( .A1(adr1[6]), .A2(_u2_n900 ), .ZN(_u2_n1122 ) );
NAND3_X1 _u2_U359  ( .A1(_u2_n1120 ), .A2(_u2_n1121 ), .A3(_u2_n1122 ), .ZN(_u2_n949 ) );
OR2_X1 _u2_U358  ( .A1(_u2_n900 ), .A2(am1[7]), .ZN(_u2_n1119 ) );
NAND2_X1 _u2_U357  ( .A1(_u2_n903 ), .A2(_u2_n1119 ), .ZN(_u2_n1118 ) );
NAND2_X1 _u2_U356  ( .A1(_u2_adr1_cnt[5] ), .A2(_u2_n1118 ), .ZN(_u2_n1115 ));
NAND3_X1 _u2_U355  ( .A1(_u2_adr1_cnt_next1[5]), .A2(_u2_n901 ), .A3(am1[7]), .ZN(_u2_n1116 ) );
NAND2_X1 _u2_U354  ( .A1(adr1[7]), .A2(_u2_n900 ), .ZN(_u2_n1117 ) );
NAND3_X1 _u2_U353  ( .A1(_u2_n1115 ), .A2(_u2_n1116 ), .A3(_u2_n1117 ), .ZN(_u2_n950 ) );
OR2_X1 _u2_U352  ( .A1(_u2_n900 ), .A2(am1[8]), .ZN(_u2_n1114 ) );
NAND2_X1 _u2_U351  ( .A1(_u2_n903 ), .A2(_u2_n1114 ), .ZN(_u2_n1113 ) );
NAND2_X1 _u2_U350  ( .A1(_u2_adr1_cnt[6] ), .A2(_u2_n1113 ), .ZN(_u2_n1110 ));
NAND3_X1 _u2_U349  ( .A1(_u2_adr1_cnt_next1[6]), .A2(_u2_n901 ), .A3(am1[8]), .ZN(_u2_n1111 ) );
NAND2_X1 _u2_U348  ( .A1(adr1[8]), .A2(_u2_n900 ), .ZN(_u2_n1112 ) );
NAND3_X1 _u2_U347  ( .A1(_u2_n1110 ), .A2(_u2_n1111 ), .A3(_u2_n1112 ), .ZN(_u2_n951 ) );
OR2_X1 _u2_U346  ( .A1(_u2_n900 ), .A2(am1[9]), .ZN(_u2_n1109 ) );
NAND2_X1 _u2_U345  ( .A1(_u2_n903 ), .A2(_u2_n1109 ), .ZN(_u2_n1108 ) );
NAND2_X1 _u2_U344  ( .A1(_u2_adr1_cnt[7] ), .A2(_u2_n1108 ), .ZN(_u2_n1105 ));
NAND3_X1 _u2_U343  ( .A1(_u2_adr1_cnt_next1[7]), .A2(_u2_n901 ), .A3(am1[9]), .ZN(_u2_n1106 ) );
NAND2_X1 _u2_U342  ( .A1(adr1[9]), .A2(_u2_n900 ), .ZN(_u2_n1107 ) );
NAND3_X1 _u2_U341  ( .A1(_u2_n1105 ), .A2(_u2_n1106 ), .A3(_u2_n1107 ), .ZN(_u2_n952 ) );
OR2_X1 _u2_U340  ( .A1(_u2_n900 ), .A2(am1[10]), .ZN(_u2_n1104 ) );
NAND2_X1 _u2_U339  ( .A1(_u2_n903 ), .A2(_u2_n1104 ), .ZN(_u2_n1103 ) );
NAND2_X1 _u2_U338  ( .A1(_u2_adr1_cnt[8] ), .A2(_u2_n1103 ), .ZN(_u2_n1100 ));
NAND3_X1 _u2_U337  ( .A1(_u2_adr1_cnt_next1[8]), .A2(_u2_n901 ), .A3(am1[10]), .ZN(_u2_n1101 ) );
NAND2_X1 _u2_U336  ( .A1(adr1[10]), .A2(_u2_n900 ), .ZN(_u2_n1102 ) );
NAND3_X1 _u2_U335  ( .A1(_u2_n1100 ), .A2(_u2_n1101 ), .A3(_u2_n1102 ), .ZN(_u2_n953 ) );
OR2_X1 _u2_U334  ( .A1(_u2_n900 ), .A2(am1[11]), .ZN(_u2_n1099 ) );
NAND2_X1 _u2_U333  ( .A1(_u2_n903 ), .A2(_u2_n1099 ), .ZN(_u2_n1098 ) );
NAND2_X1 _u2_U332  ( .A1(_u2_adr1_cnt[9] ), .A2(_u2_n1098 ), .ZN(_u2_n1095 ));
NAND3_X1 _u2_U331  ( .A1(_u2_adr1_cnt_next1[9]), .A2(_u2_n901 ), .A3(am1[11]), .ZN(_u2_n1096 ) );
NAND2_X1 _u2_U330  ( .A1(adr1[11]), .A2(_u2_n900 ), .ZN(_u2_n1097 ) );
NAND3_X1 _u2_U329  ( .A1(_u2_n1095 ), .A2(_u2_n1096 ), .A3(_u2_n1097 ), .ZN(_u2_n954 ) );
OR2_X1 _u2_U328  ( .A1(_u2_n900 ), .A2(am1[12]), .ZN(_u2_n1094 ) );
NAND2_X1 _u2_U327  ( .A1(_u2_n903 ), .A2(_u2_n1094 ), .ZN(_u2_n1093 ) );
NAND2_X1 _u2_U326  ( .A1(_u2_adr1_cnt[10] ), .A2(_u2_n1093 ), .ZN(_u2_n1090 ) );
NAND3_X1 _u2_U325  ( .A1(_u2_adr1_cnt_next1[10]), .A2(_u2_n901 ), .A3(am1[12]), .ZN(_u2_n1091 ) );
NAND2_X1 _u2_U324  ( .A1(adr1[12]), .A2(_u2_n900 ), .ZN(_u2_n1092 ) );
NAND3_X1 _u2_U323  ( .A1(_u2_n1090 ), .A2(_u2_n1091 ), .A3(_u2_n1092 ), .ZN(_u2_n955 ) );
OR2_X1 _u2_U322  ( .A1(_u2_n900 ), .A2(am1[13]), .ZN(_u2_n1089 ) );
NAND2_X1 _u2_U321  ( .A1(_u2_n903 ), .A2(_u2_n1089 ), .ZN(_u2_n1088 ) );
NAND2_X1 _u2_U320  ( .A1(_u2_adr1_cnt[11] ), .A2(_u2_n1088 ), .ZN(_u2_n1085 ) );
NAND3_X1 _u2_U319  ( .A1(_u2_adr1_cnt_next1[11]), .A2(_u2_n901 ), .A3(am1[13]), .ZN(_u2_n1086 ) );
NAND2_X1 _u2_U318  ( .A1(adr1[13]), .A2(_u2_n900 ), .ZN(_u2_n1087 ) );
NAND3_X1 _u2_U317  ( .A1(_u2_n1085 ), .A2(_u2_n1086 ), .A3(_u2_n1087 ), .ZN(_u2_n956 ) );
OR2_X1 _u2_U316  ( .A1(_u2_n900 ), .A2(am1[14]), .ZN(_u2_n1084 ) );
NAND2_X1 _u2_U315  ( .A1(_u2_n903 ), .A2(_u2_n1084 ), .ZN(_u2_n1083 ) );
NAND2_X1 _u2_U314  ( .A1(_u2_adr1_cnt[12] ), .A2(_u2_n1083 ), .ZN(_u2_n1080 ) );
NAND3_X1 _u2_U313  ( .A1(_u2_adr1_cnt_next1[12]), .A2(_u2_n901 ), .A3(am1[14]), .ZN(_u2_n1081 ) );
NAND2_X1 _u2_U312  ( .A1(adr1[14]), .A2(_u2_n900 ), .ZN(_u2_n1082 ) );
NAND3_X1 _u2_U311  ( .A1(_u2_n1080 ), .A2(_u2_n1081 ), .A3(_u2_n1082 ), .ZN(_u2_n957 ) );
OR2_X1 _u2_U310  ( .A1(_u2_n900 ), .A2(am1[15]), .ZN(_u2_n1079 ) );
NAND2_X1 _u2_U309  ( .A1(_u2_n903 ), .A2(_u2_n1079 ), .ZN(_u2_n1078 ) );
NAND2_X1 _u2_U308  ( .A1(_u2_adr1_cnt[13] ), .A2(_u2_n1078 ), .ZN(_u2_n1075 ) );
NAND3_X1 _u2_U307  ( .A1(_u2_adr1_cnt_next1[13]), .A2(_u2_n901 ), .A3(am1[15]), .ZN(_u2_n1076 ) );
NAND2_X1 _u2_U306  ( .A1(adr1[15]), .A2(_u2_n900 ), .ZN(_u2_n1077 ) );
NAND3_X1 _u2_U305  ( .A1(_u2_n1075 ), .A2(_u2_n1076 ), .A3(_u2_n1077 ), .ZN(_u2_n958 ) );
OR2_X1 _u2_U304  ( .A1(_u2_n900 ), .A2(am1[16]), .ZN(_u2_n1074 ) );
NAND2_X1 _u2_U303  ( .A1(_u2_n903 ), .A2(_u2_n1074 ), .ZN(_u2_n1073 ) );
NAND2_X1 _u2_U302  ( .A1(_u2_adr1_cnt[14] ), .A2(_u2_n1073 ), .ZN(_u2_n1070 ) );
NAND3_X1 _u2_U301  ( .A1(_u2_adr1_cnt_next1[14]), .A2(_u2_n901 ), .A3(am1[16]), .ZN(_u2_n1071 ) );
NAND2_X1 _u2_U300  ( .A1(adr1[16]), .A2(_u2_n900 ), .ZN(_u2_n1072 ) );
NAND3_X1 _u2_U299  ( .A1(_u2_n1070 ), .A2(_u2_n1071 ), .A3(_u2_n1072 ), .ZN(_u2_n959 ) );
OR2_X1 _u2_U298  ( .A1(_u2_n900 ), .A2(am1[17]), .ZN(_u2_n1069 ) );
NAND2_X1 _u2_U297  ( .A1(_u2_n903 ), .A2(_u2_n1069 ), .ZN(_u2_n1068 ) );
NAND2_X1 _u2_U296  ( .A1(_u2_adr1_cnt[15] ), .A2(_u2_n1068 ), .ZN(_u2_n1065 ) );
NAND3_X1 _u2_U295  ( .A1(_u2_adr1_cnt_next1[15]), .A2(_u2_n901 ), .A3(am1[17]), .ZN(_u2_n1066 ) );
NAND2_X1 _u2_U294  ( .A1(adr1[17]), .A2(_u2_n900 ), .ZN(_u2_n1067 ) );
NAND3_X1 _u2_U293  ( .A1(_u2_n1065 ), .A2(_u2_n1066 ), .A3(_u2_n1067 ), .ZN(_u2_n960 ) );
OR2_X1 _u2_U292  ( .A1(_u2_n900 ), .A2(am1[18]), .ZN(_u2_n1064 ) );
NAND2_X1 _u2_U291  ( .A1(_u2_n903 ), .A2(_u2_n1064 ), .ZN(_u2_n1063 ) );
NAND2_X1 _u2_U290  ( .A1(_u2_adr1_cnt[16] ), .A2(_u2_n1063 ), .ZN(_u2_n1060 ) );
NAND3_X1 _u2_U289  ( .A1(_u2_adr1_cnt_next1[16]), .A2(_u2_n901 ), .A3(am1[18]), .ZN(_u2_n1061 ) );
NAND2_X1 _u2_U288  ( .A1(adr1[18]), .A2(_u2_n900 ), .ZN(_u2_n1062 ) );
NAND3_X1 _u2_U287  ( .A1(_u2_n1060 ), .A2(_u2_n1061 ), .A3(_u2_n1062 ), .ZN(_u2_n961 ) );
OR2_X1 _u2_U286  ( .A1(_u2_n900 ), .A2(am1[19]), .ZN(_u2_n1059 ) );
NAND2_X1 _u2_U285  ( .A1(_u2_n903 ), .A2(_u2_n1059 ), .ZN(_u2_n1058 ) );
NAND2_X1 _u2_U284  ( .A1(_u2_adr1_cnt[17] ), .A2(_u2_n1058 ), .ZN(_u2_n1055 ) );
NAND3_X1 _u2_U283  ( .A1(_u2_adr1_cnt_next1[17]), .A2(_u2_n901 ), .A3(am1[19]), .ZN(_u2_n1056 ) );
NAND2_X1 _u2_U282  ( .A1(adr1[19]), .A2(_u2_n900 ), .ZN(_u2_n1057 ) );
NAND3_X1 _u2_U281  ( .A1(_u2_n1055 ), .A2(_u2_n1056 ), .A3(_u2_n1057 ), .ZN(_u2_n962 ) );
OR2_X1 _u2_U280  ( .A1(_u2_n900 ), .A2(am1[20]), .ZN(_u2_n1054 ) );
NAND2_X1 _u2_U279  ( .A1(_u2_n903 ), .A2(_u2_n1054 ), .ZN(_u2_n1051 ) );
NAND2_X1 _u2_U278  ( .A1(_u2_adr1_cnt[18] ), .A2(_u2_n1051 ), .ZN(_u2_n1048 ) );
NAND3_X1 _u2_U277  ( .A1(_u2_adr1_cnt_next1[18]), .A2(_u2_n901 ), .A3(am1[20]), .ZN(_u2_n1049 ) );
NAND2_X1 _u2_U276  ( .A1(adr1[20]), .A2(_u2_n900 ), .ZN(_u2_n1050 ) );
NAND3_X1 _u2_U275  ( .A1(_u2_n1048 ), .A2(_u2_n1049 ), .A3(_u2_n1050 ), .ZN(_u2_n963 ) );
OR2_X1 _u2_U274  ( .A1(_u2_n900 ), .A2(am1[21]), .ZN(_u2_n1047 ) );
NAND2_X1 _u2_U273  ( .A1(_u2_n903 ), .A2(_u2_n1047 ), .ZN(_u2_n1046 ) );
NAND2_X1 _u2_U272  ( .A1(_u2_adr1_cnt[19] ), .A2(_u2_n1046 ), .ZN(_u2_n1009 ) );
NAND3_X1 _u2_U271  ( .A1(_u2_adr1_cnt_next1[19]), .A2(_u2_n901 ), .A3(am1[21]), .ZN(_u2_n1010 ) );
NAND2_X1 _u2_U270  ( .A1(adr1[21]), .A2(_u2_n900 ), .ZN(_u2_n1043 ) );
NAND3_X1 _u2_U269  ( .A1(_u2_n1009 ), .A2(_u2_n1010 ), .A3(_u2_n1043 ), .ZN(_u2_n964 ) );
OR2_X1 _u2_U268  ( .A1(_u2_n900 ), .A2(am1[22]), .ZN(_u2_n1008 ) );
NAND2_X1 _u2_U267  ( .A1(_u2_n903 ), .A2(_u2_n1008 ), .ZN(_u2_n1007 ) );
NAND2_X1 _u2_U266  ( .A1(_u2_adr1_cnt[20] ), .A2(_u2_n1007 ), .ZN(_u2_n942 ));
NAND3_X1 _u2_U265  ( .A1(_u2_adr1_cnt_next1[20]), .A2(_u2_n901 ), .A3(am1[22]), .ZN(_u2_n943 ) );
NAND2_X1 _u2_U264  ( .A1(adr1[22]), .A2(_u2_n900 ), .ZN(_u2_n1005 ) );
NAND3_X1 _u2_U263  ( .A1(_u2_n942 ), .A2(_u2_n943 ), .A3(_u2_n1005 ), .ZN(_u2_n965 ) );
OR2_X1 _u2_U262  ( .A1(_u2_n900 ), .A2(am1[23]), .ZN(_u2_n941 ) );
NAND2_X1 _u2_U261  ( .A1(_u2_n903 ), .A2(_u2_n941 ), .ZN(_u2_n940 ) );
NAND2_X1 _u2_U260  ( .A1(_u2_adr1_cnt[21] ), .A2(_u2_n940 ), .ZN(_u2_n937 ));
NAND3_X1 _u2_U259  ( .A1(_u2_adr1_cnt_next1[21]), .A2(_u2_n901 ), .A3(am1[23]), .ZN(_u2_n938 ) );
NAND2_X1 _u2_U258  ( .A1(adr1[23]), .A2(_u2_n900 ), .ZN(_u2_n939 ) );
NAND3_X1 _u2_U257  ( .A1(_u2_n937 ), .A2(_u2_n938 ), .A3(_u2_n939 ), .ZN(_u2_n966 ) );
OR2_X1 _u2_U256  ( .A1(_u2_n900 ), .A2(am1[24]), .ZN(_u2_n936 ) );
NAND2_X1 _u2_U255  ( .A1(_u2_n903 ), .A2(_u2_n936 ), .ZN(_u2_n935 ) );
NAND2_X1 _u2_U254  ( .A1(_u2_adr1_cnt[22] ), .A2(_u2_n935 ), .ZN(_u2_n930 ));
NAND3_X1 _u2_U253  ( .A1(_u2_adr1_cnt_next1[22]), .A2(_u2_n901 ), .A3(am1[24]), .ZN(_u2_n932 ) );
NAND2_X1 _u2_U252  ( .A1(adr1[24]), .A2(_u2_n900 ), .ZN(_u2_n933 ) );
NAND3_X1 _u2_U251  ( .A1(_u2_n930 ), .A2(_u2_n932 ), .A3(_u2_n933 ), .ZN(_u2_n967 ) );
OR2_X1 _u2_U250  ( .A1(_u2_n900 ), .A2(am1[25]), .ZN(_u2_n929 ) );
NAND2_X1 _u2_U249  ( .A1(_u2_n903 ), .A2(_u2_n929 ), .ZN(_u2_n928 ) );
NAND2_X1 _u2_U248  ( .A1(_u2_adr1_cnt[23] ), .A2(_u2_n928 ), .ZN(_u2_n925 ));
NAND3_X1 _u2_U247  ( .A1(_u2_adr1_cnt_next1[23]), .A2(_u2_n901 ), .A3(am1[25]), .ZN(_u2_n926 ) );
NAND2_X1 _u2_U246  ( .A1(adr1[25]), .A2(_u2_n900 ), .ZN(_u2_n927 ) );
NAND3_X1 _u2_U245  ( .A1(_u2_n925 ), .A2(_u2_n926 ), .A3(_u2_n927 ), .ZN(_u2_n968 ) );
OR2_X1 _u2_U244  ( .A1(_u2_n900 ), .A2(am1[26]), .ZN(_u2_n924 ) );
NAND2_X1 _u2_U243  ( .A1(_u2_n903 ), .A2(_u2_n924 ), .ZN(_u2_n923 ) );
NAND2_X1 _u2_U242  ( .A1(_u2_adr1_cnt[24] ), .A2(_u2_n923 ), .ZN(_u2_n920 ));
NAND3_X1 _u2_U241  ( .A1(_u2_adr1_cnt_next1[24]), .A2(_u2_n901 ), .A3(am1[26]), .ZN(_u2_n921 ) );
NAND2_X1 _u2_U240  ( .A1(adr1[26]), .A2(_u2_n900 ), .ZN(_u2_n922 ) );
NAND3_X1 _u2_U239  ( .A1(_u2_n920 ), .A2(_u2_n921 ), .A3(_u2_n922 ), .ZN(_u2_n969 ) );
OR2_X1 _u2_U238  ( .A1(_u2_n900 ), .A2(am1[27]), .ZN(_u2_n919 ) );
NAND2_X1 _u2_U237  ( .A1(_u2_n903 ), .A2(_u2_n919 ), .ZN(_u2_n918 ) );
NAND2_X1 _u2_U236  ( .A1(_u2_adr1_cnt[25] ), .A2(_u2_n918 ), .ZN(_u2_n915 ));
NAND3_X1 _u2_U235  ( .A1(_u2_adr1_cnt_next1[25]), .A2(_u2_n901 ), .A3(am1[27]), .ZN(_u2_n916 ) );
NAND2_X1 _u2_U234  ( .A1(adr1[27]), .A2(_u2_n900 ), .ZN(_u2_n917 ) );
NAND3_X1 _u2_U233  ( .A1(_u2_n915 ), .A2(_u2_n916 ), .A3(_u2_n917 ), .ZN(_u2_n970 ) );
OR2_X1 _u2_U232  ( .A1(_u2_n900 ), .A2(am1[28]), .ZN(_u2_n914 ) );
NAND2_X1 _u2_U231  ( .A1(_u2_n903 ), .A2(_u2_n914 ), .ZN(_u2_n913 ) );
NAND2_X1 _u2_U230  ( .A1(_u2_adr1_cnt[26] ), .A2(_u2_n913 ), .ZN(_u2_n910 ));
NAND3_X1 _u2_U229  ( .A1(_u2_adr1_cnt_next1[26]), .A2(_u2_n901 ), .A3(am1[28]), .ZN(_u2_n911 ) );
NAND2_X1 _u2_U228  ( .A1(adr1[28]), .A2(_u2_n900 ), .ZN(_u2_n912 ) );
NAND3_X1 _u2_U227  ( .A1(_u2_n910 ), .A2(_u2_n911 ), .A3(_u2_n912 ), .ZN(_u2_n971 ) );
OR2_X1 _u2_U226  ( .A1(_u2_n900 ), .A2(am1[29]), .ZN(_u2_n909 ) );
NAND2_X1 _u2_U225  ( .A1(_u2_n903 ), .A2(_u2_n909 ), .ZN(_u2_n908 ) );
NAND2_X1 _u2_U224  ( .A1(_u2_adr1_cnt[27] ), .A2(_u2_n908 ), .ZN(_u2_n905 ));
NAND3_X1 _u2_U223  ( .A1(_u2_adr1_cnt_next1[27]), .A2(_u2_n901 ), .A3(am1[29]), .ZN(_u2_n906 ) );
NAND2_X1 _u2_U222  ( .A1(adr1[29]), .A2(_u2_n900 ), .ZN(_u2_n907 ) );
NAND3_X1 _u2_U221  ( .A1(_u2_n905 ), .A2(_u2_n906 ), .A3(_u2_n907 ), .ZN(_u2_n972 ) );
OR2_X1 _u2_U220  ( .A1(_u2_n900 ), .A2(am1[30]), .ZN(_u2_n904 ) );
NAND2_X1 _u2_U219  ( .A1(_u2_n903 ), .A2(_u2_n904 ), .ZN(_u2_n902 ) );
NAND2_X1 _u2_U218  ( .A1(_u2_adr1_cnt[28] ), .A2(_u2_n902 ), .ZN(_u2_n897 ));
NAND3_X1 _u2_U217  ( .A1(_u2_adr1_cnt_next1[28]), .A2(_u2_n901 ), .A3(am1[30]), .ZN(_u2_n898 ) );
NAND2_X1 _u2_U216  ( .A1(adr1[30]), .A2(_u2_n900 ), .ZN(_u2_n899 ) );
NAND3_X1 _u2_U215  ( .A1(_u2_n897 ), .A2(_u2_n898 ), .A3(_u2_n899 ), .ZN(_u2_n973 ) );
NAND2_X1 _u2_U214  ( .A1(_u2_adr0_cnt_next1[0]), .A2(_u2_n770 ), .ZN(_u2_n894 ) );
NAND2_X1 _u2_U213  ( .A1(_u2_adr0_cnt[0] ), .A2(_u2_n893 ), .ZN(_u2_n895 ));
NAND2_X1 _u2_U212  ( .A1(adr0[2]), .A2(_u2_n892 ), .ZN(_u2_n896 ) );
NAND3_X1 _u2_U211  ( .A1(_u2_n894 ), .A2(_u2_n895 ), .A3(_u2_n896 ), .ZN(_u2_n974 ) );
NAND2_X1 _u2_U210  ( .A1(_u2_adr0_cnt_next1[1]), .A2(_u2_n770 ), .ZN(_u2_n889 ) );
NAND2_X1 _u2_U209  ( .A1(_u2_adr0_cnt[1] ), .A2(_u2_n893 ), .ZN(_u2_n890 ));
NAND2_X1 _u2_U208  ( .A1(adr0[3]), .A2(_u2_n892 ), .ZN(_u2_n891 ) );
NAND3_X1 _u2_U207  ( .A1(_u2_n889 ), .A2(_u2_n890 ), .A3(_u2_n891 ), .ZN(_u2_n975 ) );
OR2_X1 _u2_U206  ( .A1(_u2_n769 ), .A2(am0[4]), .ZN(_u2_n888 ) );
NAND2_X1 _u2_U205  ( .A1(_u2_n772 ), .A2(_u2_n888 ), .ZN(_u2_n887 ) );
NAND2_X1 _u2_U204  ( .A1(_u2_adr0_cnt[2] ), .A2(_u2_n887 ), .ZN(_u2_n884 ));
NAND3_X1 _u2_U203  ( .A1(_u2_adr0_cnt_next1[2]), .A2(_u2_n770 ), .A3(am0[4]), .ZN(_u2_n885 ) );
NAND2_X1 _u2_U202  ( .A1(adr0[4]), .A2(_u2_n769 ), .ZN(_u2_n886 ) );
NAND3_X1 _u2_U201  ( .A1(_u2_n884 ), .A2(_u2_n885 ), .A3(_u2_n886 ), .ZN(_u2_n976 ) );
OR2_X1 _u2_U200  ( .A1(_u2_n769 ), .A2(am0[5]), .ZN(_u2_n883 ) );
NAND2_X1 _u2_U199  ( .A1(_u2_n772 ), .A2(_u2_n883 ), .ZN(_u2_n882 ) );
NAND2_X1 _u2_U198  ( .A1(_u2_adr0_cnt[3] ), .A2(_u2_n882 ), .ZN(_u2_n879 ));
NAND3_X1 _u2_U197  ( .A1(_u2_adr0_cnt_next1[3]), .A2(_u2_n770 ), .A3(am0[5]), .ZN(_u2_n880 ) );
NAND2_X1 _u2_U196  ( .A1(adr0[5]), .A2(_u2_n769 ), .ZN(_u2_n881 ) );
NAND3_X1 _u2_U195  ( .A1(_u2_n879 ), .A2(_u2_n880 ), .A3(_u2_n881 ), .ZN(_u2_n977 ) );
OR2_X1 _u2_U194  ( .A1(_u2_n769 ), .A2(am0[6]), .ZN(_u2_n878 ) );
NAND2_X1 _u2_U193  ( .A1(_u2_n772 ), .A2(_u2_n878 ), .ZN(_u2_n877 ) );
NAND2_X1 _u2_U192  ( .A1(_u2_adr0_cnt[4] ), .A2(_u2_n877 ), .ZN(_u2_n874 ));
NAND3_X1 _u2_U191  ( .A1(_u2_adr0_cnt_next1[4]), .A2(_u2_n770 ), .A3(am0[6]), .ZN(_u2_n875 ) );
NAND2_X1 _u2_U190  ( .A1(adr0[6]), .A2(_u2_n769 ), .ZN(_u2_n876 ) );
NAND3_X1 _u2_U189  ( .A1(_u2_n874 ), .A2(_u2_n875 ), .A3(_u2_n876 ), .ZN(_u2_n978 ) );
OR2_X1 _u2_U188  ( .A1(_u2_n769 ), .A2(am0[7]), .ZN(_u2_n873 ) );
NAND2_X1 _u2_U187  ( .A1(_u2_n772 ), .A2(_u2_n873 ), .ZN(_u2_n872 ) );
NAND2_X1 _u2_U186  ( .A1(_u2_adr0_cnt[5] ), .A2(_u2_n872 ), .ZN(_u2_n869 ));
NAND3_X1 _u2_U185  ( .A1(_u2_adr0_cnt_next1[5]), .A2(_u2_n770 ), .A3(am0[7]), .ZN(_u2_n870 ) );
NAND2_X1 _u2_U184  ( .A1(adr0[7]), .A2(_u2_n769 ), .ZN(_u2_n871 ) );
NAND3_X1 _u2_U183  ( .A1(_u2_n869 ), .A2(_u2_n870 ), .A3(_u2_n871 ), .ZN(_u2_n979 ) );
OR2_X1 _u2_U182  ( .A1(_u2_n769 ), .A2(am0[8]), .ZN(_u2_n868 ) );
NAND2_X1 _u2_U181  ( .A1(_u2_n772 ), .A2(_u2_n868 ), .ZN(_u2_n867 ) );
NAND2_X1 _u2_U180  ( .A1(_u2_adr0_cnt[6] ), .A2(_u2_n867 ), .ZN(_u2_n864 ));
NAND3_X1 _u2_U179  ( .A1(_u2_adr0_cnt_next1[6]), .A2(_u2_n770 ), .A3(am0[8]), .ZN(_u2_n865 ) );
NAND2_X1 _u2_U178  ( .A1(adr0[8]), .A2(_u2_n769 ), .ZN(_u2_n866 ) );
NAND3_X1 _u2_U177  ( .A1(_u2_n864 ), .A2(_u2_n865 ), .A3(_u2_n866 ), .ZN(_u2_n980 ) );
OR2_X1 _u2_U176  ( .A1(_u2_n769 ), .A2(am0[9]), .ZN(_u2_n863 ) );
NAND2_X1 _u2_U175  ( .A1(_u2_n772 ), .A2(_u2_n863 ), .ZN(_u2_n862 ) );
NAND2_X1 _u2_U174  ( .A1(_u2_adr0_cnt[7] ), .A2(_u2_n862 ), .ZN(_u2_n859 ));
NAND3_X1 _u2_U173  ( .A1(_u2_adr0_cnt_next1[7]), .A2(_u2_n770 ), .A3(am0[9]), .ZN(_u2_n860 ) );
NAND2_X1 _u2_U172  ( .A1(adr0[9]), .A2(_u2_n769 ), .ZN(_u2_n861 ) );
NAND3_X1 _u2_U171  ( .A1(_u2_n859 ), .A2(_u2_n860 ), .A3(_u2_n861 ), .ZN(_u2_n981 ) );
OR2_X1 _u2_U170  ( .A1(_u2_n769 ), .A2(am0[10]), .ZN(_u2_n858 ) );
NAND2_X1 _u2_U169  ( .A1(_u2_n772 ), .A2(_u2_n858 ), .ZN(_u2_n857 ) );
NAND2_X1 _u2_U168  ( .A1(_u2_adr0_cnt[8] ), .A2(_u2_n857 ), .ZN(_u2_n854 ));
NAND3_X1 _u2_U167  ( .A1(_u2_adr0_cnt_next1[8]), .A2(_u2_n770 ), .A3(am0[10]), .ZN(_u2_n855 ) );
NAND2_X1 _u2_U166  ( .A1(adr0[10]), .A2(_u2_n769 ), .ZN(_u2_n856 ) );
NAND3_X1 _u2_U165  ( .A1(_u2_n854 ), .A2(_u2_n855 ), .A3(_u2_n856 ), .ZN(_u2_n982 ) );
OR2_X1 _u2_U164  ( .A1(_u2_n769 ), .A2(am0[11]), .ZN(_u2_n853 ) );
NAND2_X1 _u2_U163  ( .A1(_u2_n772 ), .A2(_u2_n853 ), .ZN(_u2_n852 ) );
NAND2_X1 _u2_U162  ( .A1(_u2_adr0_cnt[9] ), .A2(_u2_n852 ), .ZN(_u2_n849 ));
NAND3_X1 _u2_U161  ( .A1(_u2_adr0_cnt_next1[9]), .A2(_u2_n770 ), .A3(am0[11]), .ZN(_u2_n850 ) );
NAND2_X1 _u2_U160  ( .A1(adr0[11]), .A2(_u2_n769 ), .ZN(_u2_n851 ) );
NAND3_X1 _u2_U159  ( .A1(_u2_n849 ), .A2(_u2_n850 ), .A3(_u2_n851 ), .ZN(_u2_n983 ) );
OR2_X1 _u2_U158  ( .A1(_u2_n769 ), .A2(am0[12]), .ZN(_u2_n848 ) );
NAND2_X1 _u2_U157  ( .A1(_u2_n772 ), .A2(_u2_n848 ), .ZN(_u2_n847 ) );
NAND2_X1 _u2_U156  ( .A1(_u2_adr0_cnt[10] ), .A2(_u2_n847 ), .ZN(_u2_n844 ));
NAND3_X1 _u2_U155  ( .A1(_u2_adr0_cnt_next1[10]), .A2(_u2_n770 ), .A3(am0[12]), .ZN(_u2_n845 ) );
NAND2_X1 _u2_U154  ( .A1(adr0[12]), .A2(_u2_n769 ), .ZN(_u2_n846 ) );
NAND3_X1 _u2_U153  ( .A1(_u2_n844 ), .A2(_u2_n845 ), .A3(_u2_n846 ), .ZN(_u2_n984 ) );
OR2_X1 _u2_U152  ( .A1(_u2_n769 ), .A2(am0[13]), .ZN(_u2_n843 ) );
NAND2_X1 _u2_U151  ( .A1(_u2_n772 ), .A2(_u2_n843 ), .ZN(_u2_n842 ) );
NAND2_X1 _u2_U150  ( .A1(_u2_adr0_cnt[11] ), .A2(_u2_n842 ), .ZN(_u2_n839 ));
NAND3_X1 _u2_U149  ( .A1(_u2_adr0_cnt_next1[11]), .A2(_u2_n770 ), .A3(am0[13]), .ZN(_u2_n840 ) );
NAND2_X1 _u2_U148  ( .A1(adr0[13]), .A2(_u2_n769 ), .ZN(_u2_n841 ) );
NAND3_X1 _u2_U147  ( .A1(_u2_n839 ), .A2(_u2_n840 ), .A3(_u2_n841 ), .ZN(_u2_n985 ) );
OR2_X1 _u2_U146  ( .A1(_u2_n769 ), .A2(am0[14]), .ZN(_u2_n838 ) );
NAND2_X1 _u2_U145  ( .A1(_u2_n772 ), .A2(_u2_n838 ), .ZN(_u2_n837 ) );
NAND2_X1 _u2_U144  ( .A1(_u2_adr0_cnt[12] ), .A2(_u2_n837 ), .ZN(_u2_n834 ));
NAND3_X1 _u2_U143  ( .A1(_u2_adr0_cnt_next1[12]), .A2(_u2_n770 ), .A3(am0[14]), .ZN(_u2_n835 ) );
NAND2_X1 _u2_U142  ( .A1(adr0[14]), .A2(_u2_n769 ), .ZN(_u2_n836 ) );
NAND3_X1 _u2_U141  ( .A1(_u2_n834 ), .A2(_u2_n835 ), .A3(_u2_n836 ), .ZN(_u2_n986 ) );
OR2_X1 _u2_U140  ( .A1(_u2_n769 ), .A2(am0[15]), .ZN(_u2_n833 ) );
NAND2_X1 _u2_U139  ( .A1(_u2_n772 ), .A2(_u2_n833 ), .ZN(_u2_n832 ) );
NAND2_X1 _u2_U138  ( .A1(_u2_adr0_cnt[13] ), .A2(_u2_n832 ), .ZN(_u2_n829 ));
NAND3_X1 _u2_U137  ( .A1(_u2_adr0_cnt_next1[13]), .A2(_u2_n770 ), .A3(am0[15]), .ZN(_u2_n830 ) );
NAND2_X1 _u2_U136  ( .A1(adr0[15]), .A2(_u2_n769 ), .ZN(_u2_n831 ) );
NAND3_X1 _u2_U135  ( .A1(_u2_n829 ), .A2(_u2_n830 ), .A3(_u2_n831 ), .ZN(_u2_n987 ) );
OR2_X1 _u2_U134  ( .A1(_u2_n769 ), .A2(am0[16]), .ZN(_u2_n828 ) );
NAND2_X1 _u2_U133  ( .A1(_u2_n772 ), .A2(_u2_n828 ), .ZN(_u2_n827 ) );
NAND2_X1 _u2_U132  ( .A1(_u2_adr0_cnt[14] ), .A2(_u2_n827 ), .ZN(_u2_n824 ));
NAND3_X1 _u2_U131  ( .A1(_u2_adr0_cnt_next1[14]), .A2(_u2_n770 ), .A3(am0[16]), .ZN(_u2_n825 ) );
NAND2_X1 _u2_U130  ( .A1(adr0[16]), .A2(_u2_n769 ), .ZN(_u2_n826 ) );
NAND3_X1 _u2_U129  ( .A1(_u2_n824 ), .A2(_u2_n825 ), .A3(_u2_n826 ), .ZN(_u2_n988 ) );
OR2_X1 _u2_U128  ( .A1(_u2_n769 ), .A2(am0[17]), .ZN(_u2_n823 ) );
NAND2_X1 _u2_U127  ( .A1(_u2_n772 ), .A2(_u2_n823 ), .ZN(_u2_n822 ) );
NAND2_X1 _u2_U126  ( .A1(_u2_adr0_cnt[15] ), .A2(_u2_n822 ), .ZN(_u2_n819 ));
NAND3_X1 _u2_U125  ( .A1(_u2_adr0_cnt_next1[15]), .A2(_u2_n770 ), .A3(am0[17]), .ZN(_u2_n820 ) );
NAND2_X1 _u2_U124  ( .A1(adr0[17]), .A2(_u2_n769 ), .ZN(_u2_n821 ) );
NAND3_X1 _u2_U123  ( .A1(_u2_n819 ), .A2(_u2_n820 ), .A3(_u2_n821 ), .ZN(_u2_n989 ) );
OR2_X1 _u2_U122  ( .A1(_u2_n769 ), .A2(am0[18]), .ZN(_u2_n818 ) );
NAND2_X1 _u2_U121  ( .A1(_u2_n772 ), .A2(_u2_n818 ), .ZN(_u2_n817 ) );
NAND2_X1 _u2_U120  ( .A1(_u2_adr0_cnt[16] ), .A2(_u2_n817 ), .ZN(_u2_n814 ));
NAND3_X1 _u2_U119  ( .A1(_u2_adr0_cnt_next1[16]), .A2(_u2_n770 ), .A3(am0[18]), .ZN(_u2_n815 ) );
NAND2_X1 _u2_U118  ( .A1(adr0[18]), .A2(_u2_n769 ), .ZN(_u2_n816 ) );
NAND3_X1 _u2_U117  ( .A1(_u2_n814 ), .A2(_u2_n815 ), .A3(_u2_n816 ), .ZN(_u2_n990 ) );
OR2_X1 _u2_U116  ( .A1(_u2_n769 ), .A2(am0[19]), .ZN(_u2_n813 ) );
NAND2_X1 _u2_U115  ( .A1(_u2_n772 ), .A2(_u2_n813 ), .ZN(_u2_n812 ) );
NAND2_X1 _u2_U114  ( .A1(_u2_adr0_cnt[17] ), .A2(_u2_n812 ), .ZN(_u2_n809 ));
NAND3_X1 _u2_U113  ( .A1(_u2_adr0_cnt_next1[17]), .A2(_u2_n770 ), .A3(am0[19]), .ZN(_u2_n810 ) );
NAND2_X1 _u2_U112  ( .A1(adr0[19]), .A2(_u2_n769 ), .ZN(_u2_n811 ) );
NAND3_X1 _u2_U111  ( .A1(_u2_n809 ), .A2(_u2_n810 ), .A3(_u2_n811 ), .ZN(_u2_n991 ) );
OR2_X1 _u2_U110  ( .A1(_u2_n769 ), .A2(am0[20]), .ZN(_u2_n808 ) );
NAND2_X1 _u2_U109  ( .A1(_u2_n772 ), .A2(_u2_n808 ), .ZN(_u2_n807 ) );
NAND2_X1 _u2_U108  ( .A1(_u2_adr0_cnt[18] ), .A2(_u2_n807 ), .ZN(_u2_n804 ));
NAND3_X1 _u2_U107  ( .A1(_u2_adr0_cnt_next1[18]), .A2(_u2_n770 ), .A3(am0[20]), .ZN(_u2_n805 ) );
NAND2_X1 _u2_U106  ( .A1(adr0[20]), .A2(_u2_n769 ), .ZN(_u2_n806 ) );
NAND3_X1 _u2_U105  ( .A1(_u2_n804 ), .A2(_u2_n805 ), .A3(_u2_n806 ), .ZN(_u2_n992 ) );
OR2_X1 _u2_U104  ( .A1(_u2_n769 ), .A2(am0[21]), .ZN(_u2_n803 ) );
NAND2_X1 _u2_U103  ( .A1(_u2_n772 ), .A2(_u2_n803 ), .ZN(_u2_n802 ) );
NAND2_X1 _u2_U102  ( .A1(_u2_adr0_cnt[19] ), .A2(_u2_n802 ), .ZN(_u2_n799 ));
NAND3_X1 _u2_U101  ( .A1(_u2_adr0_cnt_next1[19]), .A2(_u2_n770 ), .A3(am0[21]), .ZN(_u2_n800 ) );
NAND2_X1 _u2_U100  ( .A1(adr0[21]), .A2(_u2_n769 ), .ZN(_u2_n801 ) );
NAND3_X1 _u2_U99  ( .A1(_u2_n799 ), .A2(_u2_n800 ), .A3(_u2_n801 ), .ZN(_u2_n993 ) );
OR2_X1 _u2_U98  ( .A1(_u2_n769 ), .A2(am0[22]), .ZN(_u2_n798 ) );
NAND2_X1 _u2_U97  ( .A1(_u2_n772 ), .A2(_u2_n798 ), .ZN(_u2_n797 ) );
NAND2_X1 _u2_U96  ( .A1(_u2_adr0_cnt[20] ), .A2(_u2_n797 ), .ZN(_u2_n794 ));
NAND3_X1 _u2_U95  ( .A1(_u2_adr0_cnt_next1[20]), .A2(_u2_n770 ), .A3(am0[22]), .ZN(_u2_n795 ) );
NAND2_X1 _u2_U94  ( .A1(adr0[22]), .A2(_u2_n769 ), .ZN(_u2_n796 ) );
NAND3_X1 _u2_U93  ( .A1(_u2_n794 ), .A2(_u2_n795 ), .A3(_u2_n796 ), .ZN(_u2_n994 ) );
OR2_X1 _u2_U92  ( .A1(_u2_n769 ), .A2(am0[23]), .ZN(_u2_n793 ) );
NAND2_X1 _u2_U91  ( .A1(_u2_n772 ), .A2(_u2_n793 ), .ZN(_u2_n792 ) );
NAND2_X1 _u2_U90  ( .A1(_u2_adr0_cnt[21] ), .A2(_u2_n792 ), .ZN(_u2_n789 ));
NAND3_X1 _u2_U89  ( .A1(_u2_adr0_cnt_next1[21]), .A2(_u2_n770 ), .A3(am0[23]), .ZN(_u2_n790 ) );
NAND2_X1 _u2_U88  ( .A1(adr0[23]), .A2(_u2_n769 ), .ZN(_u2_n791 ) );
NAND3_X1 _u2_U87  ( .A1(_u2_n789 ), .A2(_u2_n790 ), .A3(_u2_n791 ), .ZN(_u2_n995 ) );
OR2_X1 _u2_U86  ( .A1(_u2_n769 ), .A2(am0[24]), .ZN(_u2_n788 ) );
NAND2_X1 _u2_U85  ( .A1(_u2_n772 ), .A2(_u2_n788 ), .ZN(_u2_n787 ) );
NAND2_X1 _u2_U84  ( .A1(_u2_adr0_cnt[22] ), .A2(_u2_n787 ), .ZN(_u2_n784 ));
NAND3_X1 _u2_U83  ( .A1(_u2_adr0_cnt_next1[22]), .A2(_u2_n770 ), .A3(am0[24]), .ZN(_u2_n785 ) );
NAND2_X1 _u2_U82  ( .A1(adr0[24]), .A2(_u2_n769 ), .ZN(_u2_n786 ) );
NAND3_X1 _u2_U81  ( .A1(_u2_n784 ), .A2(_u2_n785 ), .A3(_u2_n786 ), .ZN(_u2_n996 ) );
OR2_X1 _u2_U80  ( .A1(_u2_n769 ), .A2(am0[25]), .ZN(_u2_n783 ) );
NAND2_X1 _u2_U79  ( .A1(_u2_n772 ), .A2(_u2_n783 ), .ZN(_u2_n782 ) );
NAND2_X1 _u2_U78  ( .A1(_u2_adr0_cnt[23] ), .A2(_u2_n782 ), .ZN(_u2_n779 ));
NAND3_X1 _u2_U77  ( .A1(_u2_adr0_cnt_next1[23]), .A2(_u2_n770 ), .A3(am0[25]), .ZN(_u2_n780 ) );
NAND2_X1 _u2_U76  ( .A1(adr0[25]), .A2(_u2_n769 ), .ZN(_u2_n781 ) );
NAND3_X1 _u2_U75  ( .A1(_u2_n779 ), .A2(_u2_n780 ), .A3(_u2_n781 ), .ZN(_u2_n997 ) );
OR2_X1 _u2_U74  ( .A1(_u2_n769 ), .A2(am0[26]), .ZN(_u2_n778 ) );
NAND2_X1 _u2_U73  ( .A1(_u2_n772 ), .A2(_u2_n778 ), .ZN(_u2_n777 ) );
NAND2_X1 _u2_U72  ( .A1(_u2_adr0_cnt[24] ), .A2(_u2_n777 ), .ZN(_u2_n774 ));
NAND3_X1 _u2_U71  ( .A1(_u2_adr0_cnt_next1[24]), .A2(_u2_n770 ), .A3(am0[26]), .ZN(_u2_n775 ) );
NAND2_X1 _u2_U70  ( .A1(adr0[26]), .A2(_u2_n769 ), .ZN(_u2_n776 ) );
NAND3_X1 _u2_U69  ( .A1(_u2_n774 ), .A2(_u2_n775 ), .A3(_u2_n776 ), .ZN(_u2_n998 ) );
OR2_X1 _u2_U68  ( .A1(_u2_n769 ), .A2(am0[27]), .ZN(_u2_n773 ) );
NAND2_X1 _u2_U67  ( .A1(_u2_n772 ), .A2(_u2_n773 ), .ZN(_u2_n771 ) );
NAND2_X1 _u2_U66  ( .A1(_u2_adr0_cnt[25] ), .A2(_u2_n771 ), .ZN(_u2_n766 ));
NAND3_X1 _u2_U65  ( .A1(_u2_adr0_cnt_next1[25]), .A2(_u2_n770 ), .A3(am0[27]), .ZN(_u2_n767 ) );
NAND2_X1 _u2_U64  ( .A1(adr0[27]), .A2(_u2_n769 ), .ZN(_u2_n768 ) );
NAND3_X1 _u2_U63  ( .A1(_u2_n766 ), .A2(_u2_n767 ), .A3(_u2_n768 ), .ZN(_u2_n999 ) );
INV_X1 _u2_U62  ( .A(_u2_n765 ), .ZN(_u2_n1565 ) );
CLKBUF_X2 _u2_U61  ( .A(de_ack), .Z(dma_done) );
CLKBUF_X2 _u2_U60  ( .A(mast0_dout[31]), .Z(de_csr[31]) );
CLKBUF_X2 _u2_U59  ( .A(mast0_dout[30]), .Z(de_csr[30]) );
CLKBUF_X2 _u2_U58  ( .A(mast0_dout[29]), .Z(de_csr[29]) );
CLKBUF_X2 _u2_U57  ( .A(mast0_dout[28]), .Z(de_csr[28]) );
CLKBUF_X2 _u2_U56  ( .A(mast0_dout[27]), .Z(de_csr[27]) );
CLKBUF_X2 _u2_U55  ( .A(mast0_dout[26]), .Z(de_csr[26]) );
CLKBUF_X2 _u2_U54  ( .A(mast0_dout[25]), .Z(de_csr[25]) );
CLKBUF_X2 _u2_U53  ( .A(mast0_dout[24]), .Z(de_csr[24]) );
CLKBUF_X2 _u2_U52  ( .A(mast0_dout[23]), .Z(de_csr[23]) );
CLKBUF_X2 _u2_U51  ( .A(mast0_dout[22]), .Z(de_csr[22]) );
CLKBUF_X2 _u2_U50  ( .A(mast0_dout[21]), .Z(de_csr[21]) );
CLKBUF_X2 _u2_U49  ( .A(mast0_dout[20]), .Z(de_csr[20]) );
CLKBUF_X2 _u2_U48  ( .A(mast0_dout[19]), .Z(de_csr[19]) );
CLKBUF_X2 _u2_U47  ( .A(mast0_dout[18]), .Z(de_csr[18]) );
CLKBUF_X2 _u2_U46  ( .A(mast0_dout[17]), .Z(de_csr[17]) );
CLKBUF_X2 _u2_U45  ( .A(mast0_dout[16]), .Z(de_csr[16]) );
CLKBUF_X2 _u2_U44  ( .A(mast0_dout[15]), .Z(de_csr[15]) );
CLKBUF_X2 _u2_U43  ( .A(mast0_dout[14]), .Z(de_csr[14]) );
CLKBUF_X2 _u2_U42  ( .A(mast0_dout[13]), .Z(de_csr[13]) );
CLKBUF_X2 _u2_U41  ( .A(mast0_dout[12]), .Z(de_csr[12]) );
CLKBUF_X2 _u2_U40  ( .A(mast0_dout[11]), .Z(de_csr[11]) );
CLKBUF_X2 _u2_U39  ( .A(mast0_dout[10]), .Z(de_csr[10]) );
CLKBUF_X2 _u2_U38  ( .A(mast0_dout[9]), .Z(de_csr[9]) );
CLKBUF_X2 _u2_U37  ( .A(mast0_dout[8]), .Z(de_csr[8]) );
CLKBUF_X2 _u2_U36  ( .A(mast0_dout[7]), .Z(de_csr[7]) );
CLKBUF_X2 _u2_U35  ( .A(mast0_dout[6]), .Z(de_csr[6]) );
CLKBUF_X2 _u2_U34  ( .A(mast0_dout[5]), .Z(de_csr[5]) );
CLKBUF_X2 _u2_U33  ( .A(mast0_dout[4]), .Z(de_csr[4]) );
CLKBUF_X2 _u2_U32  ( .A(mast0_dout[3]), .Z(de_csr[3]) );
CLKBUF_X2 _u2_U31  ( .A(mast0_dout[2]), .Z(de_csr[2]) );
CLKBUF_X2 _u2_U30  ( .A(mast0_dout[1]), .Z(de_csr[1]) );
CLKBUF_X2 _u2_U29  ( .A(mast0_dout[0]), .Z(de_csr[0]) );
CLKBUF_X2 _u2_U28  ( .A(de_adr0[1]), .Z(de_adr1[1]) );
CLKBUF_X2 _u2_U27  ( .A(de_adr0[0]), .Z(de_adr1[0]) );
NOR2_X4 _u2_U26  ( .A1(_u2_n893 ), .A2(_u2_n770 ), .ZN(_u2_n769 ) );
NOR2_X4 _u2_U25  ( .A1(_u2_n1138 ), .A2(_u2_n901 ), .ZN(_u2_n900 ) );
NAND2_X2 _u2_U24  ( .A1(_u2_n1556 ), .A2(_u2_n1153 ), .ZN(_u2_read ) );
INV_X4 _u2_U23  ( .A(_u2_read ), .ZN(_u2_n1418 ) );
NOR2_X2 _u2_U22  ( .A1(_u2_n1288 ), .A2(_u2_n1284 ), .ZN(_u2_n1290 ) );
NOR2_X2 _u2_U21  ( .A1(_u2_n1280 ), .A2(_u2_read ), .ZN(_u2_n1427 ) );
AND4_X4 _u2_U20  ( .A1(_u2_read_r ), .A2(csr[4]), .A3(_u2_n1245 ), .A4(_u2_n1267 ), .ZN(_u2_n770 ) );
INV_X4 _u2_U19  ( .A(_u2_n1275 ), .ZN(_u2_n1429 ) );
NOR2_X2 _u2_U18  ( .A1(_u2_n1288 ), .A2(csr[2]), .ZN(_u2_n1289 ) );
NOR2_X2 _u2_U17  ( .A1(_u2_n1280 ), .A2(_u2_n1418 ), .ZN(_u2_n1428 ) );
AND4_X4 _u2_U16  ( .A1(csr[3]), .A2(_u2_n1245 ), .A3(_u2_n1246 ), .A4(_u2_n944 ), .ZN(_u2_n901 ) );
INV_X4 _u2_U15  ( .A(_u2_n893 ), .ZN(_u2_n772 ) );
INV_X4 _u2_U14  ( .A(_u2_n1138 ), .ZN(_u2_n903 ) );
INV_X4 _u2_U13  ( .A(_u2_n1551 ), .ZN(_u2_n1288 ) );
NOR2_X2 _u2_U12  ( .A1(_u2_n1278 ), .A2(_u2_n1288 ), .ZN(_u2_n1426 ) );
NAND4_X2 _u2_U11  ( .A1(_u2_n1415 ), .A2(_u2_n719 ), .A3(_u2_state_0_ ),.A4(_u2_n1416 ), .ZN(dma_busy) );
INV_X4 _u2_U10  ( .A(_u2_n726 ), .ZN(_u2_n729 ) );
INV_X4 _u2_U9  ( .A(_u2_n726 ), .ZN(_u2_n728 ) );
INV_X4 _u2_U8  ( .A(_u2_n726 ), .ZN(_u2_n727 ) );
INV_X1 _u2_U7  ( .A(_u2_n1369 ), .ZN(_u2_n726 ) );
INV_X4 _u2_U5  ( .A(1'b1), .ZN(_u2_mast1_adr[1] ) );
INV_X4 _u2_U3  ( .A(1'b1), .ZN(_u2_mast1_adr[0] ) );
DFF_X2 _u2_mast0_adr_reg_0_  ( .D(_u2_N277 ), .CK(clk_i), .Q(mast0_adr[0]),.QN() );
DFF_X2 _u2_mast0_adr_reg_1_  ( .D(_u2_N278 ), .CK(clk_i), .Q(mast0_adr[1]),.QN() );
DFF_X2 _u2_mast0_adr_reg_2_  ( .D(_u2_N279 ), .CK(clk_i), .Q(mast0_adr[2]),.QN() );
DFF_X2 _u2_mast0_adr_reg_3_  ( .D(_u2_N280 ), .CK(clk_i), .Q(mast0_adr[3]),.QN() );
DFF_X2 _u2_mast0_adr_reg_4_  ( .D(_u2_N281 ), .CK(clk_i), .Q(mast0_adr[4]),.QN() );
DFF_X2 _u2_mast0_adr_reg_5_  ( .D(_u2_N282 ), .CK(clk_i), .Q(mast0_adr[5]),.QN() );
DFF_X2 _u2_mast0_adr_reg_6_  ( .D(_u2_N283 ), .CK(clk_i), .Q(mast0_adr[6]),.QN() );
DFF_X2 _u2_mast0_adr_reg_7_  ( .D(_u2_N284 ), .CK(clk_i), .Q(mast0_adr[7]),.QN() );
DFF_X2 _u2_mast0_adr_reg_8_  ( .D(_u2_N285 ), .CK(clk_i), .Q(mast0_adr[8]),.QN() );
DFF_X2 _u2_mast0_adr_reg_9_  ( .D(_u2_N286 ), .CK(clk_i), .Q(mast0_adr[9]),.QN() );
DFF_X2 _u2_mast0_adr_reg_10_  ( .D(_u2_N287 ), .CK(clk_i), .Q(mast0_adr[10]),.QN() );
DFF_X2 _u2_mast0_adr_reg_11_  ( .D(_u2_N288 ), .CK(clk_i), .Q(mast0_adr[11]),.QN() );
DFF_X2 _u2_mast0_adr_reg_12_  ( .D(_u2_N289 ), .CK(clk_i), .Q(mast0_adr[12]),.QN() );
DFF_X2 _u2_mast0_adr_reg_13_  ( .D(_u2_N290 ), .CK(clk_i), .Q(mast0_adr[13]),.QN() );
DFF_X2 _u2_mast0_adr_reg_14_  ( .D(_u2_N291 ), .CK(clk_i), .Q(mast0_adr[14]),.QN() );
DFF_X2 _u2_mast0_adr_reg_15_  ( .D(_u2_N292 ), .CK(clk_i), .Q(mast0_adr[15]),.QN() );
DFF_X2 _u2_mast0_adr_reg_16_  ( .D(_u2_N293 ), .CK(clk_i), .Q(mast0_adr[16]),.QN() );
DFF_X2 _u2_mast0_adr_reg_17_  ( .D(_u2_N294 ), .CK(clk_i), .Q(mast0_adr[17]),.QN() );
DFF_X2 _u2_mast0_adr_reg_18_  ( .D(_u2_N295 ), .CK(clk_i), .Q(mast0_adr[18]),.QN() );
DFF_X2 _u2_mast0_adr_reg_19_  ( .D(_u2_N296 ), .CK(clk_i), .Q(mast0_adr[19]),.QN() );
DFF_X2 _u2_mast0_adr_reg_20_  ( .D(_u2_N297 ), .CK(clk_i), .Q(mast0_adr[20]),.QN() );
DFF_X2 _u2_mast0_adr_reg_21_  ( .D(_u2_N298 ), .CK(clk_i), .Q(mast0_adr[21]),.QN() );
DFF_X2 _u2_mast0_adr_reg_22_  ( .D(_u2_N299 ), .CK(clk_i), .Q(mast0_adr[22]),.QN() );
DFF_X2 _u2_mast0_adr_reg_23_  ( .D(_u2_N300 ), .CK(clk_i), .Q(mast0_adr[23]),.QN() );
DFF_X2 _u2_mast0_adr_reg_24_  ( .D(_u2_N301 ), .CK(clk_i), .Q(mast0_adr[24]),.QN() );
DFF_X2 _u2_mast0_adr_reg_25_  ( .D(_u2_N302 ), .CK(clk_i), .Q(mast0_adr[25]),.QN() );
DFF_X2 _u2_mast0_adr_reg_26_  ( .D(_u2_N303 ), .CK(clk_i), .Q(mast0_adr[26]),.QN() );
DFF_X2 _u2_mast0_adr_reg_27_  ( .D(_u2_N304 ), .CK(clk_i), .Q(mast0_adr[27]),.QN() );
DFF_X2 _u2_mast0_adr_reg_28_  ( .D(_u2_N305 ), .CK(clk_i), .Q(mast0_adr[28]),.QN() );
DFF_X2 _u2_mast0_adr_reg_29_  ( .D(_u2_N306 ), .CK(clk_i), .Q(mast0_adr[29]),.QN() );
DFF_X2 _u2_mast0_adr_reg_30_  ( .D(_u2_N307 ), .CK(clk_i), .Q(mast0_adr[30]),.QN() );
DFF_X2 _u2_mast0_adr_reg_31_  ( .D(_u2_N308 ), .CK(clk_i), .Q(mast0_adr[31]),.QN() );
DFF_X2 _u2_write_hold_r_reg  ( .D(_u2_N342 ), .CK(clk_i), .Q(_u2_write_hold_r ), .QN() );
DFF_X2 _u2_mast1_adr_reg_31_  ( .D(_u2_N341 ), .CK(clk_i), .Q(mast1_adr[31]),.QN() );
DFF_X2 _u2_mast1_adr_reg_2_  ( .D(_u2_N312 ), .CK(clk_i), .Q(mast1_adr[2]),.QN() );
DFF_X2 _u2_mast1_adr_reg_3_  ( .D(_u2_N313 ), .CK(clk_i), .Q(mast1_adr[3]),.QN() );
DFF_X2 _u2_mast1_adr_reg_4_  ( .D(_u2_N314 ), .CK(clk_i), .Q(mast1_adr[4]),.QN() );
DFF_X2 _u2_mast1_adr_reg_5_  ( .D(_u2_N315 ), .CK(clk_i), .Q(mast1_adr[5]),.QN() );
DFF_X2 _u2_mast1_adr_reg_6_  ( .D(_u2_N316 ), .CK(clk_i), .Q(mast1_adr[6]),.QN() );
DFF_X2 _u2_mast1_adr_reg_7_  ( .D(_u2_N317 ), .CK(clk_i), .Q(mast1_adr[7]),.QN() );
DFF_X2 _u2_mast1_adr_reg_8_  ( .D(_u2_N318 ), .CK(clk_i), .Q(mast1_adr[8]),.QN() );
DFF_X2 _u2_mast1_adr_reg_9_  ( .D(_u2_N319 ), .CK(clk_i), .Q(mast1_adr[9]),.QN() );
DFF_X2 _u2_mast1_adr_reg_10_  ( .D(_u2_N320 ), .CK(clk_i), .Q(mast1_adr[10]),.QN() );
DFF_X2 _u2_mast1_adr_reg_11_  ( .D(_u2_N321 ), .CK(clk_i), .Q(mast1_adr[11]),.QN() );
DFF_X2 _u2_mast1_adr_reg_12_  ( .D(_u2_N322 ), .CK(clk_i), .Q(mast1_adr[12]),.QN() );
DFF_X2 _u2_mast1_adr_reg_13_  ( .D(_u2_N323 ), .CK(clk_i), .Q(mast1_adr[13]),.QN() );
DFF_X2 _u2_mast1_adr_reg_14_  ( .D(_u2_N324 ), .CK(clk_i), .Q(mast1_adr[14]),.QN() );
DFF_X2 _u2_mast1_adr_reg_15_  ( .D(_u2_N325 ), .CK(clk_i), .Q(mast1_adr[15]),.QN() );
DFF_X2 _u2_mast1_adr_reg_16_  ( .D(_u2_N326 ), .CK(clk_i), .Q(mast1_adr[16]),.QN() );
DFF_X2 _u2_mast1_adr_reg_17_  ( .D(_u2_N327 ), .CK(clk_i), .Q(mast1_adr[17]),.QN() );
DFF_X2 _u2_mast1_adr_reg_18_  ( .D(_u2_N328 ), .CK(clk_i), .Q(mast1_adr[18]),.QN() );
DFF_X2 _u2_mast1_adr_reg_19_  ( .D(_u2_N329 ), .CK(clk_i), .Q(mast1_adr[19]),.QN() );
DFF_X2 _u2_mast1_adr_reg_20_  ( .D(_u2_N330 ), .CK(clk_i), .Q(mast1_adr[20]),.QN() );
DFF_X2 _u2_mast1_adr_reg_21_  ( .D(_u2_N331 ), .CK(clk_i), .Q(mast1_adr[21]),.QN() );
DFF_X2 _u2_mast1_adr_reg_22_  ( .D(_u2_N332 ), .CK(clk_i), .Q(mast1_adr[22]),.QN() );
DFF_X2 _u2_mast1_adr_reg_23_  ( .D(_u2_N333 ), .CK(clk_i), .Q(mast1_adr[23]),.QN() );
DFF_X2 _u2_mast1_adr_reg_24_  ( .D(_u2_N334 ), .CK(clk_i), .Q(mast1_adr[24]),.QN() );
DFF_X2 _u2_mast1_adr_reg_25_  ( .D(_u2_N335 ), .CK(clk_i), .Q(mast1_adr[25]),.QN() );
DFF_X2 _u2_mast1_adr_reg_26_  ( .D(_u2_N336 ), .CK(clk_i), .Q(mast1_adr[26]),.QN() );
DFF_X2 _u2_mast1_adr_reg_27_  ( .D(_u2_N337 ), .CK(clk_i), .Q(mast1_adr[27]),.QN() );
DFF_X2 _u2_mast1_adr_reg_28_  ( .D(_u2_N338 ), .CK(clk_i), .Q(mast1_adr[28]),.QN() );
DFF_X2 _u2_mast1_adr_reg_29_  ( .D(_u2_N339 ), .CK(clk_i), .Q(mast1_adr[29]),.QN() );
DFF_X2 _u2_mast1_adr_reg_30_  ( .D(_u2_N340 ), .CK(clk_i), .Q(mast1_adr[30]),.QN() );
DFF_X2 _u2_next_ch_reg  ( .D(de_ack), .CK(clk_i), .Q(next_ch), .QN() );
DFF_X2 _u2_chunk_cnt_is_0_r_reg  ( .D(_u2_n1044 ), .CK(clk_i), .Q(), .QN(_u2_n934 ) );
DFF_X2 _u2_chunk_cnt_reg_8_  ( .D(_u2_n1012 ), .CK(clk_i), .Q(_u2_chunk_cnt[8] ), .QN() );
DFF_X2 _u2_chunk_cnt_reg_7_  ( .D(_u2_n1013 ), .CK(clk_i), .Q(_u2_chunk_cnt[7] ), .QN() );
DFF_X2 _u2_chunk_cnt_reg_6_  ( .D(_u2_n1014 ), .CK(clk_i), .Q(_u2_chunk_cnt[6] ), .QN() );
DFF_X2 _u2_chunk_cnt_reg_5_  ( .D(_u2_n1015 ), .CK(clk_i), .Q(_u2_chunk_cnt[5] ), .QN(_u2_n1052 ) );
DFF_X2 _u2_chunk_cnt_reg_4_  ( .D(_u2_n1016 ), .CK(clk_i), .Q(_u2_chunk_cnt[4] ), .QN() );
DFF_X2 _u2_chunk_cnt_reg_3_  ( .D(_u2_n1017 ), .CK(clk_i), .Q(_u2_chunk_cnt[3] ), .QN() );
DFF_X2 _u2_chunk_cnt_reg_2_  ( .D(_u2_n1018 ), .CK(clk_i), .Q(_u2_chunk_cnt[2] ), .QN() );
DFF_X2 _u2_chunk_cnt_reg_1_  ( .D(_u2_n1019 ), .CK(clk_i), .Q(_u2_chunk_cnt[1] ), .QN(_u2_n1053 ) );
DFF_X2 _u2_chunk_cnt_reg_0_  ( .D(_u2_n1020 ), .CK(clk_i), .Q(_u2_chunk_cnt[0] ), .QN() );
DFF_X2 _u2_chunk_dec_reg  ( .D(_u2_N232 ), .CK(clk_i), .Q(_u2_chunk_dec ),.QN() );
DFF_X2 _u2_tsz_cnt_is_0_r_reg  ( .D(_u2_n1565 ), .CK(clk_i), .Q(_u2_tsz_cnt_is_0_r ), .QN() );
DFF_X2 _u2_tsz_cnt_reg_10_  ( .D(_u2_n1031 ), .CK(clk_i), .Q(_u2_tsz_cnt[10] ), .QN() );
DFF_X2 _u2_tsz_cnt_reg_9_  ( .D(_u2_n1030 ), .CK(clk_i), .Q(_u2_tsz_cnt[9] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_8_  ( .D(_u2_n1029 ), .CK(clk_i), .Q(_u2_tsz_cnt[8] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_7_  ( .D(_u2_n1028 ), .CK(clk_i), .Q(_u2_tsz_cnt[7] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_6_  ( .D(_u2_n1027 ), .CK(clk_i), .Q(_u2_tsz_cnt[6] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_5_  ( .D(_u2_n1026 ), .CK(clk_i), .Q(_u2_tsz_cnt[5] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_4_  ( .D(_u2_n1025 ), .CK(clk_i), .Q(_u2_tsz_cnt[4] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_3_  ( .D(_u2_n1024 ), .CK(clk_i), .Q(_u2_tsz_cnt[3] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_2_  ( .D(_u2_n1023 ), .CK(clk_i), .Q(_u2_tsz_cnt[2] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_1_  ( .D(_u2_n1022 ), .CK(clk_i), .Q(_u2_tsz_cnt[1] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_0_  ( .D(_u2_n1021 ), .CK(clk_i), .Q(_u2_tsz_cnt[0] ),.QN() );
DFF_X2 _u2_tsz_cnt_reg_11_  ( .D(_u2_n1038 ), .CK(clk_i), .Q(_u2_tsz_cnt[11] ), .QN() );
DFF_X2 _u2_tsz_dec_reg  ( .D(_u2_N232 ), .CK(clk_i), .Q(), .QN(_u2_n725 ) );
DFF_X2 _u2_adr1_cnt_reg_0_  ( .D(_u2_n945 ), .CK(clk_i), .Q(_u2_adr1_cnt[0] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_1_  ( .D(_u2_n946 ), .CK(clk_i), .Q(_u2_adr1_cnt[1] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_2_  ( .D(_u2_n947 ), .CK(clk_i), .Q(_u2_adr1_cnt[2] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_3_  ( .D(_u2_n948 ), .CK(clk_i), .Q(_u2_adr1_cnt[3] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_4_  ( .D(_u2_n949 ), .CK(clk_i), .Q(_u2_adr1_cnt[4] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_5_  ( .D(_u2_n950 ), .CK(clk_i), .Q(_u2_adr1_cnt[5] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_6_  ( .D(_u2_n951 ), .CK(clk_i), .Q(_u2_adr1_cnt[6] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_7_  ( .D(_u2_n952 ), .CK(clk_i), .Q(_u2_adr1_cnt[7] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_8_  ( .D(_u2_n953 ), .CK(clk_i), .Q(_u2_adr1_cnt[8] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_9_  ( .D(_u2_n954 ), .CK(clk_i), .Q(_u2_adr1_cnt[9] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_10_  ( .D(_u2_n955 ), .CK(clk_i), .Q(_u2_adr1_cnt[10] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_11_  ( .D(_u2_n956 ), .CK(clk_i), .Q(_u2_adr1_cnt[11] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_12_  ( .D(_u2_n957 ), .CK(clk_i), .Q(_u2_adr1_cnt[12] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_13_  ( .D(_u2_n958 ), .CK(clk_i), .Q(_u2_adr1_cnt[13] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_14_  ( .D(_u2_n959 ), .CK(clk_i), .Q(_u2_adr1_cnt[14] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_15_  ( .D(_u2_n960 ), .CK(clk_i), .Q(_u2_adr1_cnt[15] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_16_  ( .D(_u2_n961 ), .CK(clk_i), .Q(_u2_adr1_cnt[16] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_17_  ( .D(_u2_n962 ), .CK(clk_i), .Q(_u2_adr1_cnt[17] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_18_  ( .D(_u2_n963 ), .CK(clk_i), .Q(_u2_adr1_cnt[18] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_19_  ( .D(_u2_n964 ), .CK(clk_i), .Q(_u2_adr1_cnt[19] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_20_  ( .D(_u2_n965 ), .CK(clk_i), .Q(_u2_adr1_cnt[20] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_21_  ( .D(_u2_n966 ), .CK(clk_i), .Q(_u2_adr1_cnt[21] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_22_  ( .D(_u2_n967 ), .CK(clk_i), .Q(_u2_adr1_cnt[22] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_23_  ( .D(_u2_n968 ), .CK(clk_i), .Q(_u2_adr1_cnt[23] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_24_  ( .D(_u2_n969 ), .CK(clk_i), .Q(_u2_adr1_cnt[24] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_25_  ( .D(_u2_n970 ), .CK(clk_i), .Q(_u2_adr1_cnt[25] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_26_  ( .D(_u2_n971 ), .CK(clk_i), .Q(_u2_adr1_cnt[26] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_27_  ( .D(_u2_n972 ), .CK(clk_i), .Q(_u2_adr1_cnt[27] ), .QN() );
DFF_X2 _u2_adr1_cnt_reg_28_  ( .D(_u2_n973 ), .CK(clk_i), .Q(_u2_adr1_cnt[28] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_0_  ( .D(_u2_n974 ), .CK(clk_i), .Q(_u2_adr0_cnt[0] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_1_  ( .D(_u2_n975 ), .CK(clk_i), .Q(_u2_adr0_cnt[1] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_2_  ( .D(_u2_n976 ), .CK(clk_i), .Q(_u2_adr0_cnt[2] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_3_  ( .D(_u2_n977 ), .CK(clk_i), .Q(_u2_adr0_cnt[3] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_4_  ( .D(_u2_n978 ), .CK(clk_i), .Q(_u2_adr0_cnt[4] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_5_  ( .D(_u2_n979 ), .CK(clk_i), .Q(_u2_adr0_cnt[5] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_6_  ( .D(_u2_n980 ), .CK(clk_i), .Q(_u2_adr0_cnt[6] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_7_  ( .D(_u2_n981 ), .CK(clk_i), .Q(_u2_adr0_cnt[7] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_8_  ( .D(_u2_n982 ), .CK(clk_i), .Q(_u2_adr0_cnt[8] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_9_  ( .D(_u2_n983 ), .CK(clk_i), .Q(_u2_adr0_cnt[9] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_10_  ( .D(_u2_n984 ), .CK(clk_i), .Q(_u2_adr0_cnt[10] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_11_  ( .D(_u2_n985 ), .CK(clk_i), .Q(_u2_adr0_cnt[11] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_12_  ( .D(_u2_n986 ), .CK(clk_i), .Q(_u2_adr0_cnt[12] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_13_  ( .D(_u2_n987 ), .CK(clk_i), .Q(_u2_adr0_cnt[13] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_14_  ( .D(_u2_n988 ), .CK(clk_i), .Q(_u2_adr0_cnt[14] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_15_  ( .D(_u2_n989 ), .CK(clk_i), .Q(_u2_adr0_cnt[15] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_16_  ( .D(_u2_n990 ), .CK(clk_i), .Q(_u2_adr0_cnt[16] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_17_  ( .D(_u2_n991 ), .CK(clk_i), .Q(_u2_adr0_cnt[17] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_18_  ( .D(_u2_n992 ), .CK(clk_i), .Q(_u2_adr0_cnt[18] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_19_  ( .D(_u2_n993 ), .CK(clk_i), .Q(_u2_adr0_cnt[19] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_20_  ( .D(_u2_n994 ), .CK(clk_i), .Q(_u2_adr0_cnt[20] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_21_  ( .D(_u2_n995 ), .CK(clk_i), .Q(_u2_adr0_cnt[21] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_22_  ( .D(_u2_n996 ), .CK(clk_i), .Q(_u2_adr0_cnt[22] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_23_  ( .D(_u2_n997 ), .CK(clk_i), .Q(_u2_adr0_cnt[23] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_24_  ( .D(_u2_n998 ), .CK(clk_i), .Q(_u2_adr0_cnt[24] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_25_  ( .D(_u2_n999 ), .CK(clk_i), .Q(_u2_adr0_cnt[25] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_26_  ( .D(_u2_n1000 ), .CK(clk_i), .Q(_u2_adr0_cnt[26] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_27_  ( .D(_u2_n1001 ), .CK(clk_i), .Q(_u2_adr0_cnt[27] ), .QN() );
DFF_X2 _u2_adr0_cnt_reg_28_  ( .D(_u2_n1002 ), .CK(clk_i), .Q(_u2_adr0_cnt[28] ), .QN() );
DFF_X2 _u2_mast0_drdy_r_reg  ( .D(mast0_drdy), .CK(clk_i), .Q(_u2_n1564 ),.QN() );
DFF_X2 _u2_dma_abort_r_reg  ( .D(_u2_N236 ), .CK(clk_i), .Q(dma_err), .QN(_u2_n1006 ) );
DFF_X2 _u2_chunk_0_reg  ( .D(_u2_n1045 ), .CK(clk_i), .Q(), .QN(_u2_n931 ));
DFF_X2 _u2_adr0_cnt_reg_29_  ( .D(_u2_n1003 ), .CK(clk_i), .Q(_u2_adr0_cnt[29] ), .QN() );
DFF_X2 _u2_read_r_reg  ( .D(_u2_read ), .CK(clk_i), .Q(_u2_read_r ), .QN());
DFF_X2 _u2_adr1_cnt_reg_29_  ( .D(_u2_n1004 ), .CK(clk_i), .Q(_u2_adr1_cnt[29] ), .QN() );
DFF_X2 _u2_write_r_reg  ( .D(_u2_n1566 ), .CK(clk_i), .Q(_u2_n944 ), .QN());
DFFR_X1 _u2_state_reg_9_  ( .D(_u2_n1040 ), .CK(clk_i), .RN(n5), .Q(_u2_state_9_ ), .QN() );
DFFR_X1 _u2_state_reg_3_  ( .D(_u2_n1037 ), .CK(clk_i), .RN(n5), .Q(_u2_state_3_ ), .QN(_u2_n719 ) );
DFFR_X1 _u2_state_reg_8_  ( .D(_u2_n1032 ), .CK(clk_i), .RN(n5), .Q(ptr_set),.QN(_u2_n720 ) );
DFFR_X1 _u2_state_reg_7_  ( .D(_u2_n1033 ), .CK(clk_i), .RN(n5), .Q(_u2_state_7_ ), .QN(_u2_n718 ) );
DFFR_X1 _u2_state_reg_6_  ( .D(_u2_n1034 ), .CK(clk_i), .RN(n5), .Q(_u2_state_6_ ), .QN(_u2_n724 ) );
DFFR_X1 _u2_state_reg_5_  ( .D(_u2_n1035 ), .CK(clk_i), .RN(n5), .Q(_u2_state_5_ ), .QN(_u2_n723 ) );
DFFR_X1 _u2_state_reg_4_  ( .D(_u2_n1036 ), .CK(clk_i), .RN(n5), .Q(_u2_state_4_ ), .QN() );
DFFR_X1 _u2_state_reg_2_  ( .D(_u2_n1011 ), .CK(clk_i), .RN(n5), .Q(_u2_state_2_ ), .QN() );
DFFR_X1 _u2_state_reg_1_  ( .D(_u2_n1039 ), .CK(clk_i), .RN(n5), .Q(_u2_state_1_ ), .QN(_u2_n722 ) );
DFFR_X1 _u2_state_reg_10_  ( .D(_u2_n1041 ), .CK(clk_i), .RN(n5), .Q(paused),.QN() );
DFFS_X1 _u2_state_reg_0_  ( .D(_u2_n1042 ), .CK(clk_i), .SN(n5), .Q(_u2_state_0_ ), .QN(_u2_n721 ) );
NOR2_X2 _u2_sub_360_S2_U20  ( .A1(_u2_tsz_cnt[10] ), .A2(_u2_sub_360_S2_n21 ), .ZN(_u2_sub_360_S2_n39 ) );
INV_X4 _u2_sub_360_S2_U31  ( .A(_u2_tsz_cnt[0] ), .ZN(_u2_N204 ) );
OR2_X2 _u2_sub_360_S2_U30  ( .A1(_u2_tsz_cnt[1] ), .A2(_u2_tsz_cnt[0] ),.ZN(_u2_sub_360_S2_n37 ) );
OR2_X2 _u2_sub_360_S2_U29  ( .A1(_u2_sub_360_S2_n37 ), .A2(_u2_tsz_cnt[2] ),.ZN(_u2_sub_360_S2_n35 ) );
OR2_X2 _u2_sub_360_S2_U28  ( .A1(_u2_sub_360_S2_n35 ), .A2(_u2_tsz_cnt[3] ),.ZN(_u2_sub_360_S2_n33 ) );
OR2_X2 _u2_sub_360_S2_U27  ( .A1(_u2_sub_360_S2_n33 ), .A2(_u2_tsz_cnt[4] ),.ZN(_u2_sub_360_S2_n31 ) );
OR2_X2 _u2_sub_360_S2_U26  ( .A1(_u2_sub_360_S2_n31 ), .A2(_u2_tsz_cnt[5] ),.ZN(_u2_sub_360_S2_n29 ) );
OR2_X2 _u2_sub_360_S2_U25  ( .A1(_u2_sub_360_S2_n29 ), .A2(_u2_tsz_cnt[6] ),.ZN(_u2_sub_360_S2_n27 ) );
OR2_X2 _u2_sub_360_S2_U24  ( .A1(_u2_sub_360_S2_n27 ), .A2(_u2_tsz_cnt[7] ),.ZN(_u2_sub_360_S2_n25 ) );
OR2_X2 _u2_sub_360_S2_U23  ( .A1(_u2_sub_360_S2_n25 ), .A2(_u2_tsz_cnt[8] ),.ZN(_u2_sub_360_S2_n23 ) );
OR2_X2 _u2_sub_360_S2_U22  ( .A1(_u2_sub_360_S2_n23 ), .A2(_u2_tsz_cnt[9] ),.ZN(_u2_sub_360_S2_n21 ) );
XNOR2_X2 _u2_sub_360_S2_U21  ( .A(_u2_tsz_cnt[10] ), .B(_u2_sub_360_S2_n21 ),.ZN(_u2_N214 ) );
XOR2_X2 _u2_sub_360_S2_U19  ( .A(_u2_tsz_cnt[11] ), .B(_u2_sub_360_S2_n39 ),.Z(_u2_N215 ) );
NAND2_X2 _u2_sub_360_S2_U18  ( .A1(_u2_tsz_cnt[1] ), .A2(_u2_tsz_cnt[0] ),.ZN(_u2_sub_360_S2_n38 ) );
NAND2_X2 _u2_sub_360_S2_U17  ( .A1(_u2_sub_360_S2_n37 ), .A2(_u2_sub_360_S2_n38 ), .ZN(_u2_N205 ) );
NAND2_X2 _u2_sub_360_S2_U16  ( .A1(_u2_tsz_cnt[2] ), .A2(_u2_sub_360_S2_n37 ), .ZN(_u2_sub_360_S2_n36 ) );
NAND2_X2 _u2_sub_360_S2_U15  ( .A1(_u2_sub_360_S2_n35 ), .A2(_u2_sub_360_S2_n36 ), .ZN(_u2_N206 ) );
NAND2_X2 _u2_sub_360_S2_U14  ( .A1(_u2_tsz_cnt[3] ), .A2(_u2_sub_360_S2_n35 ), .ZN(_u2_sub_360_S2_n34 ) );
NAND2_X2 _u2_sub_360_S2_U13  ( .A1(_u2_sub_360_S2_n33 ), .A2(_u2_sub_360_S2_n34 ), .ZN(_u2_N207 ) );
NAND2_X2 _u2_sub_360_S2_U12  ( .A1(_u2_tsz_cnt[4] ), .A2(_u2_sub_360_S2_n33 ), .ZN(_u2_sub_360_S2_n32 ) );
NAND2_X2 _u2_sub_360_S2_U11  ( .A1(_u2_sub_360_S2_n31 ), .A2(_u2_sub_360_S2_n32 ), .ZN(_u2_N208 ) );
NAND2_X2 _u2_sub_360_S2_U10  ( .A1(_u2_tsz_cnt[5] ), .A2(_u2_sub_360_S2_n31 ), .ZN(_u2_sub_360_S2_n30 ) );
NAND2_X2 _u2_sub_360_S2_U9  ( .A1(_u2_sub_360_S2_n29 ), .A2(_u2_sub_360_S2_n30 ), .ZN(_u2_N209 ) );
NAND2_X2 _u2_sub_360_S2_U8  ( .A1(_u2_tsz_cnt[6] ), .A2(_u2_sub_360_S2_n29 ),.ZN(_u2_sub_360_S2_n28 ) );
NAND2_X2 _u2_sub_360_S2_U7  ( .A1(_u2_sub_360_S2_n27 ), .A2(_u2_sub_360_S2_n28 ), .ZN(_u2_N210 ) );
NAND2_X2 _u2_sub_360_S2_U6  ( .A1(_u2_tsz_cnt[7] ), .A2(_u2_sub_360_S2_n27 ),.ZN(_u2_sub_360_S2_n26 ) );
NAND2_X2 _u2_sub_360_S2_U5  ( .A1(_u2_sub_360_S2_n25 ), .A2(_u2_sub_360_S2_n26 ), .ZN(_u2_N211 ) );
NAND2_X2 _u2_sub_360_S2_U4  ( .A1(_u2_tsz_cnt[8] ), .A2(_u2_sub_360_S2_n25 ),.ZN(_u2_sub_360_S2_n24 ) );
NAND2_X2 _u2_sub_360_S2_U3  ( .A1(_u2_sub_360_S2_n23 ), .A2(_u2_sub_360_S2_n24 ), .ZN(_u2_N212 ) );
NAND2_X2 _u2_sub_360_S2_U2  ( .A1(_u2_tsz_cnt[9] ), .A2(_u2_sub_360_S2_n23 ),.ZN(_u2_sub_360_S2_n22 ) );
NAND2_X2 _u2_sub_360_S2_U1  ( .A1(_u2_sub_360_S2_n21 ), .A2(_u2_sub_360_S2_n22 ), .ZN(_u2_N213 ) );
NOR2_X2 _u2_sub_349_S2_U2  ( .A1(_u2_chunk_cnt[7] ), .A2(_u2_sub_349_S2_n16 ), .ZN(_u2_sub_349_S2_n15 ) );
INV_X4 _u2_sub_349_S2_U22  ( .A(_u2_chunk_cnt[0] ), .ZN(_u2_N180 ) );
OR2_X2 _u2_sub_349_S2_U21  ( .A1(_u2_chunk_cnt[1] ), .A2(_u2_chunk_cnt[0] ),.ZN(_u2_sub_349_S2_n26 ) );
NAND2_X2 _u2_sub_349_S2_U20  ( .A1(_u2_chunk_cnt[1] ), .A2(_u2_chunk_cnt[0] ), .ZN(_u2_sub_349_S2_n27 ) );
NAND2_X2 _u2_sub_349_S2_U19  ( .A1(_u2_sub_349_S2_n26 ), .A2(_u2_sub_349_S2_n27 ), .ZN(_u2_N181 ) );
OR2_X2 _u2_sub_349_S2_U18  ( .A1(_u2_sub_349_S2_n26 ), .A2(_u2_chunk_cnt[2] ), .ZN(_u2_sub_349_S2_n24 ) );
NAND2_X2 _u2_sub_349_S2_U17  ( .A1(_u2_chunk_cnt[2] ), .A2(_u2_sub_349_S2_n26 ), .ZN(_u2_sub_349_S2_n25 ) );
NAND2_X2 _u2_sub_349_S2_U16  ( .A1(_u2_sub_349_S2_n24 ), .A2(_u2_sub_349_S2_n25 ), .ZN(_u2_N182 ) );
OR2_X2 _u2_sub_349_S2_U15  ( .A1(_u2_sub_349_S2_n24 ), .A2(_u2_chunk_cnt[3] ), .ZN(_u2_sub_349_S2_n22 ) );
NAND2_X2 _u2_sub_349_S2_U14  ( .A1(_u2_chunk_cnt[3] ), .A2(_u2_sub_349_S2_n24 ), .ZN(_u2_sub_349_S2_n23 ) );
NAND2_X2 _u2_sub_349_S2_U13  ( .A1(_u2_sub_349_S2_n22 ), .A2(_u2_sub_349_S2_n23 ), .ZN(_u2_N183 ) );
OR2_X2 _u2_sub_349_S2_U12  ( .A1(_u2_sub_349_S2_n22 ), .A2(_u2_chunk_cnt[4] ), .ZN(_u2_sub_349_S2_n20 ) );
NAND2_X2 _u2_sub_349_S2_U11  ( .A1(_u2_chunk_cnt[4] ), .A2(_u2_sub_349_S2_n22 ), .ZN(_u2_sub_349_S2_n21 ) );
NAND2_X2 _u2_sub_349_S2_U10  ( .A1(_u2_sub_349_S2_n20 ), .A2(_u2_sub_349_S2_n21 ), .ZN(_u2_N184 ) );
OR2_X2 _u2_sub_349_S2_U9  ( .A1(_u2_sub_349_S2_n20 ), .A2(_u2_chunk_cnt[5] ),.ZN(_u2_sub_349_S2_n18 ) );
NAND2_X2 _u2_sub_349_S2_U8  ( .A1(_u2_chunk_cnt[5] ), .A2(_u2_sub_349_S2_n20 ), .ZN(_u2_sub_349_S2_n19 ) );
NAND2_X2 _u2_sub_349_S2_U7  ( .A1(_u2_sub_349_S2_n18 ), .A2(_u2_sub_349_S2_n19 ), .ZN(_u2_N185 ) );
OR2_X2 _u2_sub_349_S2_U6  ( .A1(_u2_sub_349_S2_n18 ), .A2(_u2_chunk_cnt[6] ),.ZN(_u2_sub_349_S2_n16 ) );
NAND2_X2 _u2_sub_349_S2_U5  ( .A1(_u2_chunk_cnt[6] ), .A2(_u2_sub_349_S2_n18 ), .ZN(_u2_sub_349_S2_n17 ) );
NAND2_X2 _u2_sub_349_S2_U4  ( .A1(_u2_sub_349_S2_n16 ), .A2(_u2_sub_349_S2_n17 ), .ZN(_u2_N186 ) );
XNOR2_X2 _u2_sub_349_S2_U3  ( .A(_u2_chunk_cnt[7] ), .B(_u2_sub_349_S2_n16 ),.ZN(_u2_N187 ) );
XOR2_X2 _u2_sub_349_S2_U1  ( .A(_u2_chunk_cnt[8] ), .B(_u2_sub_349_S2_n15 ),.Z(_u2_N188 ) );
INV_X1 _u3_u0_U146  ( .A(mast0_go), .ZN(_u3_u0_n42 ) );
NOR2_X1 _u3_u0_U145  ( .A1(mast0_wait), .A2(_u3_u0_n42 ), .ZN(_u3_u0_N3 ) );
MUX2_X1 _u3_u0_U144  ( .A(mast0_dout[0]), .B(wb0s_data_i[0]), .S(wb0_ack_i),.Z(_u3_u0_n202 ) );
MUX2_X1 _u3_u0_U143  ( .A(mast0_dout[1]), .B(wb0s_data_i[1]), .S(wb0_ack_i),.Z(_u3_u0_n203 ) );
MUX2_X1 _u3_u0_U142  ( .A(mast0_dout[2]), .B(wb0s_data_i[2]), .S(wb0_ack_i),.Z(_u3_u0_n204 ) );
MUX2_X1 _u3_u0_U141  ( .A(mast0_dout[3]), .B(wb0s_data_i[3]), .S(wb0_ack_i),.Z(_u3_u0_n205 ) );
MUX2_X1 _u3_u0_U140  ( .A(mast0_dout[4]), .B(wb0s_data_i[4]), .S(wb0_ack_i),.Z(_u3_u0_n206 ) );
MUX2_X1 _u3_u0_U139  ( .A(mast0_dout[5]), .B(wb0s_data_i[5]), .S(wb0_ack_i),.Z(_u3_u0_n207 ) );
MUX2_X1 _u3_u0_U138  ( .A(mast0_dout[6]), .B(wb0s_data_i[6]), .S(wb0_ack_i),.Z(_u3_u0_n208 ) );
MUX2_X1 _u3_u0_U137  ( .A(mast0_dout[7]), .B(wb0s_data_i[7]), .S(wb0_ack_i),.Z(_u3_u0_n209 ) );
MUX2_X1 _u3_u0_U136  ( .A(mast0_dout[8]), .B(wb0s_data_i[8]), .S(wb0_ack_i),.Z(_u3_u0_n210 ) );
MUX2_X1 _u3_u0_U135  ( .A(mast0_dout[9]), .B(wb0s_data_i[9]), .S(wb0_ack_i),.Z(_u3_u0_n211 ) );
MUX2_X1 _u3_u0_U134  ( .A(mast0_dout[10]), .B(wb0s_data_i[10]), .S(wb0_ack_i), .Z(_u3_u0_n212 ) );
MUX2_X1 _u3_u0_U133  ( .A(mast0_dout[11]), .B(wb0s_data_i[11]), .S(wb0_ack_i), .Z(_u3_u0_n213 ) );
MUX2_X1 _u3_u0_U132  ( .A(mast0_dout[12]), .B(wb0s_data_i[12]), .S(wb0_ack_i), .Z(_u3_u0_n214 ) );
MUX2_X1 _u3_u0_U131  ( .A(mast0_dout[13]), .B(wb0s_data_i[13]), .S(wb0_ack_i), .Z(_u3_u0_n215 ) );
MUX2_X1 _u3_u0_U130  ( .A(mast0_dout[14]), .B(wb0s_data_i[14]), .S(wb0_ack_i), .Z(_u3_u0_n216 ) );
MUX2_X1 _u3_u0_U129  ( .A(mast0_dout[15]), .B(wb0s_data_i[15]), .S(wb0_ack_i), .Z(_u3_u0_n217 ) );
MUX2_X1 _u3_u0_U128  ( .A(mast0_dout[16]), .B(wb0s_data_i[16]), .S(wb0_ack_i), .Z(_u3_u0_n218 ) );
MUX2_X1 _u3_u0_U127  ( .A(mast0_dout[17]), .B(wb0s_data_i[17]), .S(wb0_ack_i), .Z(_u3_u0_n219 ) );
MUX2_X1 _u3_u0_U126  ( .A(mast0_dout[18]), .B(wb0s_data_i[18]), .S(wb0_ack_i), .Z(_u3_u0_n220 ) );
MUX2_X1 _u3_u0_U125  ( .A(mast0_dout[19]), .B(wb0s_data_i[19]), .S(wb0_ack_i), .Z(_u3_u0_n221 ) );
MUX2_X1 _u3_u0_U124  ( .A(mast0_dout[20]), .B(wb0s_data_i[20]), .S(wb0_ack_i), .Z(_u3_u0_n222 ) );
MUX2_X1 _u3_u0_U123  ( .A(mast0_dout[21]), .B(wb0s_data_i[21]), .S(wb0_ack_i), .Z(_u3_u0_n223 ) );
MUX2_X1 _u3_u0_U122  ( .A(mast0_dout[22]), .B(wb0s_data_i[22]), .S(wb0_ack_i), .Z(_u3_u0_n224 ) );
MUX2_X1 _u3_u0_U121  ( .A(mast0_dout[23]), .B(wb0s_data_i[23]), .S(wb0_ack_i), .Z(_u3_u0_n225 ) );
MUX2_X1 _u3_u0_U120  ( .A(mast0_dout[24]), .B(wb0s_data_i[24]), .S(wb0_ack_i), .Z(_u3_u0_n226 ) );
MUX2_X1 _u3_u0_U119  ( .A(mast0_dout[25]), .B(wb0s_data_i[25]), .S(wb0_ack_i), .Z(_u3_u0_n227 ) );
MUX2_X1 _u3_u0_U118  ( .A(mast0_dout[26]), .B(wb0s_data_i[26]), .S(wb0_ack_i), .Z(_u3_u0_n228 ) );
MUX2_X1 _u3_u0_U117  ( .A(mast0_dout[27]), .B(wb0s_data_i[27]), .S(wb0_ack_i), .Z(_u3_u0_n229 ) );
MUX2_X1 _u3_u0_U116  ( .A(mast0_dout[28]), .B(wb0s_data_i[28]), .S(wb0_ack_i), .Z(_u3_u0_n230 ) );
MUX2_X1 _u3_u0_U115  ( .A(mast0_dout[29]), .B(wb0s_data_i[29]), .S(wb0_ack_i), .Z(_u3_u0_n231 ) );
MUX2_X1 _u3_u0_U114  ( .A(mast0_dout[30]), .B(wb0s_data_i[30]), .S(wb0_ack_i), .Z(_u3_u0_n232 ) );
MUX2_X1 _u3_u0_U113  ( .A(mast0_dout[31]), .B(wb0s_data_i[31]), .S(wb0_ack_i), .Z(_u3_u0_n233 ) );
MUX2_X1 _u3_u0_U112  ( .A(mast0_adr[0]), .B(mast0_pt_in[7]), .S(pt0_sel_i),.Z(wb0_addr_o[0]) );
MUX2_X1 _u3_u0_U111  ( .A(mast0_adr[10]), .B(mast0_pt_in[17]), .S(pt0_sel_i),.Z(wb0_addr_o[10]) );
MUX2_X1 _u3_u0_U110  ( .A(mast0_adr[11]), .B(mast0_pt_in[18]), .S(pt0_sel_i),.Z(wb0_addr_o[11]) );
MUX2_X1 _u3_u0_U109  ( .A(mast0_adr[12]), .B(mast0_pt_in[19]), .S(pt0_sel_i),.Z(wb0_addr_o[12]) );
MUX2_X1 _u3_u0_U108  ( .A(mast0_adr[13]), .B(mast0_pt_in[20]), .S(pt0_sel_i),.Z(wb0_addr_o[13]) );
MUX2_X1 _u3_u0_U107  ( .A(mast0_adr[14]), .B(mast0_pt_in[21]), .S(pt0_sel_i),.Z(wb0_addr_o[14]) );
MUX2_X1 _u3_u0_U106  ( .A(mast0_adr[15]), .B(mast0_pt_in[22]), .S(pt0_sel_i),.Z(wb0_addr_o[15]) );
MUX2_X1 _u3_u0_U105  ( .A(mast0_adr[16]), .B(mast0_pt_in[23]), .S(pt0_sel_i),.Z(wb0_addr_o[16]) );
MUX2_X1 _u3_u0_U104  ( .A(mast0_adr[17]), .B(mast0_pt_in[24]), .S(pt0_sel_i),.Z(wb0_addr_o[17]) );
MUX2_X1 _u3_u0_U103  ( .A(mast0_adr[18]), .B(mast0_pt_in[25]), .S(pt0_sel_i),.Z(wb0_addr_o[18]) );
MUX2_X1 _u3_u0_U102  ( .A(mast0_adr[19]), .B(mast0_pt_in[26]), .S(pt0_sel_i),.Z(wb0_addr_o[19]) );
MUX2_X1 _u3_u0_U101  ( .A(mast0_adr[1]), .B(mast0_pt_in[8]), .S(pt0_sel_i),.Z(wb0_addr_o[1]) );
MUX2_X1 _u3_u0_U100  ( .A(mast0_adr[20]), .B(mast0_pt_in[27]), .S(pt0_sel_i),.Z(wb0_addr_o[20]) );
MUX2_X1 _u3_u0_U99  ( .A(mast0_adr[21]), .B(mast0_pt_in[28]), .S(pt0_sel_i),.Z(wb0_addr_o[21]) );
MUX2_X1 _u3_u0_U98  ( .A(mast0_adr[22]), .B(mast0_pt_in[29]), .S(pt0_sel_i),.Z(wb0_addr_o[22]) );
MUX2_X1 _u3_u0_U97  ( .A(mast0_adr[23]), .B(mast0_pt_in[30]), .S(pt0_sel_i),.Z(wb0_addr_o[23]) );
MUX2_X1 _u3_u0_U96  ( .A(mast0_adr[24]), .B(mast0_pt_in[31]), .S(pt0_sel_i),.Z(wb0_addr_o[24]) );
MUX2_X1 _u3_u0_U95  ( .A(mast0_adr[25]), .B(mast0_pt_in[32]), .S(pt0_sel_i),.Z(wb0_addr_o[25]) );
MUX2_X1 _u3_u0_U94  ( .A(mast0_adr[26]), .B(mast0_pt_in[33]), .S(pt0_sel_i),.Z(wb0_addr_o[26]) );
MUX2_X1 _u3_u0_U93  ( .A(mast0_adr[27]), .B(mast0_pt_in[34]), .S(pt0_sel_i),.Z(wb0_addr_o[27]) );
MUX2_X1 _u3_u0_U92  ( .A(mast0_adr[28]), .B(mast0_pt_in[35]), .S(pt0_sel_i),.Z(wb0_addr_o[28]) );
MUX2_X1 _u3_u0_U91  ( .A(mast0_adr[29]), .B(mast0_pt_in[36]), .S(pt0_sel_i),.Z(wb0_addr_o[29]) );
MUX2_X1 _u3_u0_U90  ( .A(mast0_adr[2]), .B(mast0_pt_in[9]), .S(pt0_sel_i),.Z(wb0_addr_o[2]) );
MUX2_X1 _u3_u0_U89  ( .A(mast0_adr[30]), .B(mast0_pt_in[37]), .S(pt0_sel_i),.Z(wb0_addr_o[30]) );
MUX2_X1 _u3_u0_U88  ( .A(mast0_adr[31]), .B(mast0_pt_in[38]), .S(pt0_sel_i),.Z(wb0_addr_o[31]) );
MUX2_X1 _u3_u0_U87  ( .A(mast0_adr[3]), .B(mast0_pt_in[10]), .S(pt0_sel_i),.Z(wb0_addr_o[3]) );
MUX2_X1 _u3_u0_U86  ( .A(mast0_adr[4]), .B(mast0_pt_in[11]), .S(pt0_sel_i),.Z(wb0_addr_o[4]) );
MUX2_X1 _u3_u0_U85  ( .A(mast0_adr[5]), .B(mast0_pt_in[12]), .S(pt0_sel_i),.Z(wb0_addr_o[5]) );
MUX2_X1 _u3_u0_U84  ( .A(mast0_adr[6]), .B(mast0_pt_in[13]), .S(pt0_sel_i),.Z(wb0_addr_o[6]) );
MUX2_X1 _u3_u0_U83  ( .A(mast0_adr[7]), .B(mast0_pt_in[14]), .S(pt0_sel_i),.Z(wb0_addr_o[7]) );
MUX2_X1 _u3_u0_U82  ( .A(mast0_adr[8]), .B(mast0_pt_in[15]), .S(pt0_sel_i),.Z(wb0_addr_o[8]) );
MUX2_X1 _u3_u0_U81  ( .A(mast0_adr[9]), .B(mast0_pt_in[16]), .S(pt0_sel_i),.Z(wb0_addr_o[9]) );
MUX2_X1 _u3_u0_U80  ( .A(_u3_u0_mast_cyc ), .B(mast0_pt_in[1]), .S(pt0_sel_i), .Z(wb0_cyc_o) );
MUX2_X1 _u3_u0_U79  ( .A(mast0_din[0]), .B(mast0_pt_in[39]), .S(pt0_sel_i),.Z(wb0s_data_o[0]) );
MUX2_X1 _u3_u0_U78  ( .A(mast0_din[10]), .B(mast0_pt_in[49]), .S(pt0_sel_i),.Z(wb0s_data_o[10]) );
MUX2_X1 _u3_u0_U77  ( .A(mast0_din[11]), .B(mast0_pt_in[50]), .S(pt0_sel_i),.Z(wb0s_data_o[11]) );
MUX2_X1 _u3_u0_U76  ( .A(mast0_din[12]), .B(mast0_pt_in[51]), .S(pt0_sel_i),.Z(wb0s_data_o[12]) );
MUX2_X1 _u3_u0_U75  ( .A(mast0_din[13]), .B(mast0_pt_in[52]), .S(pt0_sel_i),.Z(wb0s_data_o[13]) );
MUX2_X1 _u3_u0_U74  ( .A(mast0_din[14]), .B(mast0_pt_in[53]), .S(pt0_sel_i),.Z(wb0s_data_o[14]) );
MUX2_X1 _u3_u0_U73  ( .A(mast0_din[15]), .B(mast0_pt_in[54]), .S(pt0_sel_i),.Z(wb0s_data_o[15]) );
MUX2_X1 _u3_u0_U72  ( .A(mast0_din[16]), .B(mast0_pt_in[55]), .S(pt0_sel_i),.Z(wb0s_data_o[16]) );
MUX2_X1 _u3_u0_U71  ( .A(mast0_din[17]), .B(mast0_pt_in[56]), .S(pt0_sel_i),.Z(wb0s_data_o[17]) );
MUX2_X1 _u3_u0_U70  ( .A(mast0_din[18]), .B(mast0_pt_in[57]), .S(pt0_sel_i),.Z(wb0s_data_o[18]) );
MUX2_X1 _u3_u0_U69  ( .A(mast0_din[19]), .B(mast0_pt_in[58]), .S(pt0_sel_i),.Z(wb0s_data_o[19]) );
MUX2_X1 _u3_u0_U68  ( .A(mast0_din[1]), .B(mast0_pt_in[40]), .S(pt0_sel_i),.Z(wb0s_data_o[1]) );
MUX2_X1 _u3_u0_U67  ( .A(mast0_din[20]), .B(mast0_pt_in[59]), .S(pt0_sel_i),.Z(wb0s_data_o[20]) );
MUX2_X1 _u3_u0_U66  ( .A(mast0_din[21]), .B(mast0_pt_in[60]), .S(pt0_sel_i),.Z(wb0s_data_o[21]) );
MUX2_X1 _u3_u0_U65  ( .A(mast0_din[22]), .B(mast0_pt_in[61]), .S(pt0_sel_i),.Z(wb0s_data_o[22]) );
MUX2_X1 _u3_u0_U64  ( .A(mast0_din[23]), .B(mast0_pt_in[62]), .S(pt0_sel_i),.Z(wb0s_data_o[23]) );
MUX2_X1 _u3_u0_U63  ( .A(mast0_din[24]), .B(mast0_pt_in[63]), .S(pt0_sel_i),.Z(wb0s_data_o[24]) );
MUX2_X1 _u3_u0_U62  ( .A(mast0_din[25]), .B(mast0_pt_in[64]), .S(pt0_sel_i),.Z(wb0s_data_o[25]) );
MUX2_X1 _u3_u0_U61  ( .A(mast0_din[26]), .B(mast0_pt_in[65]), .S(pt0_sel_i),.Z(wb0s_data_o[26]) );
MUX2_X1 _u3_u0_U60  ( .A(mast0_din[27]), .B(mast0_pt_in[66]), .S(pt0_sel_i),.Z(wb0s_data_o[27]) );
MUX2_X1 _u3_u0_U59  ( .A(mast0_din[28]), .B(mast0_pt_in[67]), .S(pt0_sel_i),.Z(wb0s_data_o[28]) );
MUX2_X1 _u3_u0_U58  ( .A(mast0_din[29]), .B(mast0_pt_in[68]), .S(pt0_sel_i),.Z(wb0s_data_o[29]) );
MUX2_X1 _u3_u0_U57  ( .A(mast0_din[2]), .B(mast0_pt_in[41]), .S(pt0_sel_i),.Z(wb0s_data_o[2]) );
MUX2_X1 _u3_u0_U56  ( .A(mast0_din[30]), .B(mast0_pt_in[69]), .S(pt0_sel_i),.Z(wb0s_data_o[30]) );
MUX2_X1 _u3_u0_U55  ( .A(mast0_din[31]), .B(mast0_pt_in[70]), .S(pt0_sel_i),.Z(wb0s_data_o[31]) );
MUX2_X1 _u3_u0_U54  ( .A(mast0_din[3]), .B(mast0_pt_in[42]), .S(pt0_sel_i),.Z(wb0s_data_o[3]) );
MUX2_X1 _u3_u0_U53  ( .A(mast0_din[4]), .B(mast0_pt_in[43]), .S(pt0_sel_i),.Z(wb0s_data_o[4]) );
MUX2_X1 _u3_u0_U52  ( .A(mast0_din[5]), .B(mast0_pt_in[44]), .S(pt0_sel_i),.Z(wb0s_data_o[5]) );
MUX2_X1 _u3_u0_U51  ( .A(mast0_din[6]), .B(mast0_pt_in[45]), .S(pt0_sel_i),.Z(wb0s_data_o[6]) );
MUX2_X1 _u3_u0_U50  ( .A(mast0_din[7]), .B(mast0_pt_in[46]), .S(pt0_sel_i),.Z(wb0s_data_o[7]) );
MUX2_X1 _u3_u0_U49  ( .A(mast0_din[8]), .B(mast0_pt_in[47]), .S(pt0_sel_i),.Z(wb0s_data_o[8]) );
MUX2_X1 _u3_u0_U48  ( .A(mast0_din[9]), .B(mast0_pt_in[48]), .S(pt0_sel_i),.Z(wb0s_data_o[9]) );
INV_X1 _u3_u0_U47  ( .A(pt0_sel_i), .ZN(_u3_u0_n41 ) );
OR2_X1 _u3_u0_U46  ( .A1(mast0_pt_in[3]), .A2(_u3_u0_n41 ), .ZN(wb0_sel_o[0]) );
OR2_X1 _u3_u0_U45  ( .A1(mast0_pt_in[4]), .A2(_u3_u0_n41 ), .ZN(wb0_sel_o[1]) );
OR2_X1 _u3_u0_U44  ( .A1(mast0_pt_in[5]), .A2(_u3_u0_n41 ), .ZN(wb0_sel_o[2]) );
OR2_X1 _u3_u0_U43  ( .A1(mast0_pt_in[6]), .A2(_u3_u0_n41 ), .ZN(wb0_sel_o[3]) );
MUX2_X1 _u3_u0_U42  ( .A(_u3_u0_mast_stb ), .B(mast0_pt_in[0]), .S(pt0_sel_i), .Z(wb0_stb_o) );
MUX2_X1 _u3_u0_U41  ( .A(_u3_u0_mast_we_r ), .B(mast0_pt_in[2]), .S(pt0_sel_i), .Z(wb0_we_o) );
CLKBUF_X2 _u3_u0_U40  ( .A(wb0s_data_i[31]), .Z(slv1_pt_in[34]) );
CLKBUF_X2 _u3_u0_U39  ( .A(wb0s_data_i[30]), .Z(slv1_pt_in[33]) );
CLKBUF_X2 _u3_u0_U38  ( .A(wb0s_data_i[29]), .Z(slv1_pt_in[32]) );
CLKBUF_X2 _u3_u0_U37  ( .A(wb0s_data_i[28]), .Z(slv1_pt_in[31]) );
CLKBUF_X2 _u3_u0_U36  ( .A(wb0s_data_i[27]), .Z(slv1_pt_in[30]) );
CLKBUF_X2 _u3_u0_U35  ( .A(wb0s_data_i[26]), .Z(slv1_pt_in[29]) );
CLKBUF_X2 _u3_u0_U34  ( .A(wb0s_data_i[25]), .Z(slv1_pt_in[28]) );
CLKBUF_X2 _u3_u0_U33  ( .A(wb0s_data_i[24]), .Z(slv1_pt_in[27]) );
CLKBUF_X2 _u3_u0_U32  ( .A(wb0s_data_i[23]), .Z(slv1_pt_in[26]) );
CLKBUF_X2 _u3_u0_U31  ( .A(wb0s_data_i[22]), .Z(slv1_pt_in[25]) );
CLKBUF_X2 _u3_u0_U30  ( .A(wb0s_data_i[21]), .Z(slv1_pt_in[24]) );
CLKBUF_X2 _u3_u0_U29  ( .A(wb0s_data_i[20]), .Z(slv1_pt_in[23]) );
CLKBUF_X2 _u3_u0_U28  ( .A(wb0s_data_i[19]), .Z(slv1_pt_in[22]) );
CLKBUF_X2 _u3_u0_U27  ( .A(wb0s_data_i[18]), .Z(slv1_pt_in[21]) );
CLKBUF_X2 _u3_u0_U26  ( .A(wb0s_data_i[17]), .Z(slv1_pt_in[20]) );
CLKBUF_X2 _u3_u0_U25  ( .A(wb0s_data_i[16]), .Z(slv1_pt_in[19]) );
CLKBUF_X2 _u3_u0_U24  ( .A(wb0s_data_i[15]), .Z(slv1_pt_in[18]) );
CLKBUF_X2 _u3_u0_U23  ( .A(wb0s_data_i[14]), .Z(slv1_pt_in[17]) );
CLKBUF_X2 _u3_u0_U22  ( .A(wb0s_data_i[13]), .Z(slv1_pt_in[16]) );
CLKBUF_X2 _u3_u0_U21  ( .A(wb0s_data_i[12]), .Z(slv1_pt_in[15]) );
CLKBUF_X2 _u3_u0_U20  ( .A(wb0s_data_i[11]), .Z(slv1_pt_in[14]) );
CLKBUF_X2 _u3_u0_U19  ( .A(wb0s_data_i[10]), .Z(slv1_pt_in[13]) );
CLKBUF_X2 _u3_u0_U18  ( .A(wb0s_data_i[9]), .Z(slv1_pt_in[12]) );
CLKBUF_X2 _u3_u0_U17  ( .A(wb0s_data_i[8]), .Z(slv1_pt_in[11]) );
CLKBUF_X2 _u3_u0_U16  ( .A(wb0s_data_i[7]), .Z(slv1_pt_in[10]) );
CLKBUF_X2 _u3_u0_U15  ( .A(wb0s_data_i[6]), .Z(slv1_pt_in[9]) );
CLKBUF_X2 _u3_u0_U14  ( .A(wb0s_data_i[5]), .Z(slv1_pt_in[8]) );
CLKBUF_X2 _u3_u0_U13  ( .A(wb0s_data_i[4]), .Z(slv1_pt_in[7]) );
CLKBUF_X2 _u3_u0_U12  ( .A(wb0s_data_i[3]), .Z(slv1_pt_in[6]) );
CLKBUF_X2 _u3_u0_U11  ( .A(wb0s_data_i[2]), .Z(slv1_pt_in[5]) );
CLKBUF_X2 _u3_u0_U10  ( .A(wb0s_data_i[1]), .Z(slv1_pt_in[4]) );
CLKBUF_X2 _u3_u0_U9  ( .A(wb0s_data_i[0]), .Z(slv1_pt_in[3]) );
INV_X4 _u3_u0_U8  ( .A(_u3_u0_n6 ), .ZN(slv1_pt_in[2]) );
INV_X4 _u3_u0_U7  ( .A(_u3_u0_n6 ), .ZN(mast0_drdy) );
INV_X4 _u3_u0_U6  ( .A(wb0_ack_i), .ZN(_u3_u0_n6 ) );
CLKBUF_X2 _u3_u0_U5  ( .A(wb0_err_i), .Z(slv1_pt_in[1]) );
CLKBUF_X2 _u3_u0_U4  ( .A(wb0_err_i), .Z(mast0_err) );
CLKBUF_X2 _u3_u0_U3  ( .A(wb0_rty_i), .Z(slv1_pt_in[0]) );
DFF_X2 _u3_u0_mast_stb_reg  ( .D(_u3_u0_N3 ), .CK(clk_i), .Q(_u3_u0_mast_stb ), .QN() );
DFF_X2 _u3_u0_mast_cyc_reg  ( .D(mast0_go), .CK(clk_i), .Q(_u3_u0_mast_cyc ),.QN() );
DFF_X2 _u3_u0_mast_we_r_reg  ( .D(mast0_we), .CK(clk_i), .Q(_u3_u0_mast_we_r ), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_0_  ( .D(_u3_u0_n202 ), .CK(clk_i), .Q(mast0_dout[0]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_1_  ( .D(_u3_u0_n203 ), .CK(clk_i), .Q(mast0_dout[1]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_2_  ( .D(_u3_u0_n204 ), .CK(clk_i), .Q(mast0_dout[2]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_3_  ( .D(_u3_u0_n205 ), .CK(clk_i), .Q(mast0_dout[3]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_4_  ( .D(_u3_u0_n206 ), .CK(clk_i), .Q(mast0_dout[4]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_5_  ( .D(_u3_u0_n207 ), .CK(clk_i), .Q(mast0_dout[5]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_6_  ( .D(_u3_u0_n208 ), .CK(clk_i), .Q(mast0_dout[6]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_7_  ( .D(_u3_u0_n209 ), .CK(clk_i), .Q(mast0_dout[7]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_8_  ( .D(_u3_u0_n210 ), .CK(clk_i), .Q(mast0_dout[8]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_9_  ( .D(_u3_u0_n211 ), .CK(clk_i), .Q(mast0_dout[9]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_10_  ( .D(_u3_u0_n212 ), .CK(clk_i), .Q(mast0_dout[10]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_11_  ( .D(_u3_u0_n213 ), .CK(clk_i), .Q(mast0_dout[11]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_12_  ( .D(_u3_u0_n214 ), .CK(clk_i), .Q(mast0_dout[12]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_13_  ( .D(_u3_u0_n215 ), .CK(clk_i), .Q(mast0_dout[13]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_14_  ( .D(_u3_u0_n216 ), .CK(clk_i), .Q(mast0_dout[14]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_15_  ( .D(_u3_u0_n217 ), .CK(clk_i), .Q(mast0_dout[15]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_16_  ( .D(_u3_u0_n218 ), .CK(clk_i), .Q(mast0_dout[16]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_17_  ( .D(_u3_u0_n219 ), .CK(clk_i), .Q(mast0_dout[17]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_18_  ( .D(_u3_u0_n220 ), .CK(clk_i), .Q(mast0_dout[18]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_19_  ( .D(_u3_u0_n221 ), .CK(clk_i), .Q(mast0_dout[19]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_20_  ( .D(_u3_u0_n222 ), .CK(clk_i), .Q(mast0_dout[20]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_21_  ( .D(_u3_u0_n223 ), .CK(clk_i), .Q(mast0_dout[21]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_22_  ( .D(_u3_u0_n224 ), .CK(clk_i), .Q(mast0_dout[22]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_23_  ( .D(_u3_u0_n225 ), .CK(clk_i), .Q(mast0_dout[23]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_24_  ( .D(_u3_u0_n226 ), .CK(clk_i), .Q(mast0_dout[24]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_25_  ( .D(_u3_u0_n227 ), .CK(clk_i), .Q(mast0_dout[25]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_26_  ( .D(_u3_u0_n228 ), .CK(clk_i), .Q(mast0_dout[26]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_27_  ( .D(_u3_u0_n229 ), .CK(clk_i), .Q(mast0_dout[27]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_28_  ( .D(_u3_u0_n230 ), .CK(clk_i), .Q(mast0_dout[28]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_29_  ( .D(_u3_u0_n231 ), .CK(clk_i), .Q(mast0_dout[29]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_30_  ( .D(_u3_u0_n232 ), .CK(clk_i), .Q(mast0_dout[30]), .QN() );
DFF_X2 _u3_u0_mast_dout_reg_31_  ( .D(_u3_u0_n233 ), .CK(clk_i), .Q(mast0_dout[31]), .QN() );
NAND3_X1 _u3_u1_U120  ( .A1(wb0_cyc_i), .A2(_u3_u1_n12 ), .A3(wb0_stb_i),.ZN(_u3_u1_n90 ) );
OR4_X1 _u3_u1_U119  ( .A1(wb0_addr_i[29]), .A2(wb0_addr_i[28]), .A3(wb0_addr_i[31]), .A4(wb0_addr_i[30]), .ZN(_u3_u1_n88 ) );
NOR4_X1 _u3_u1_U118  ( .A1(wb0_we_i), .A2(slv0_re), .A3(_u3_u1_n90 ), .A4(_u3_u1_n88 ), .ZN(_u3_u1_N3 ) );
INV_X1 _u3_u1_U117  ( .A(wb0_we_i), .ZN(_u3_u1_n91 ) );
NOR3_X1 _u3_u1_U116  ( .A1(_u3_u1_n91 ), .A2(_u3_u1_n90 ), .A3(_u3_u1_n88 ),.ZN(_u3_u1_N4 ) );
NOR2_X1 _u3_u1_U115  ( .A1(slv0_re), .A2(slv0_we), .ZN(_u3_u1_n89 ) );
NOR2_X1 _u3_u1_U114  ( .A1(_u3_u1_n89 ), .A2(_u3_u1_n90 ), .ZN(_u3_u1_N5 ));
MUX2_X1 _u3_u1_U113  ( .A(_u3_u1_rf_ack ), .B(slv0_pt_in[2]), .S(_u3_u1_n16 ), .Z(wb0_ack_o) );
MUX2_X1 _u3_u1_U112  ( .A(slv0_din[0]), .B(slv0_pt_in[3]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[0]) );
MUX2_X1 _u3_u1_U111  ( .A(slv0_din[10]), .B(slv0_pt_in[13]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[10]) );
MUX2_X1 _u3_u1_U110  ( .A(slv0_din[11]), .B(slv0_pt_in[14]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[11]) );
MUX2_X1 _u3_u1_U109  ( .A(slv0_din[12]), .B(slv0_pt_in[15]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[12]) );
MUX2_X1 _u3_u1_U108  ( .A(slv0_din[13]), .B(slv0_pt_in[16]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[13]) );
MUX2_X1 _u3_u1_U107  ( .A(slv0_din[14]), .B(slv0_pt_in[17]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[14]) );
MUX2_X1 _u3_u1_U106  ( .A(slv0_din[15]), .B(slv0_pt_in[18]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[15]) );
MUX2_X1 _u3_u1_U105  ( .A(slv0_din[16]), .B(slv0_pt_in[19]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[16]) );
MUX2_X1 _u3_u1_U104  ( .A(slv0_din[17]), .B(slv0_pt_in[20]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[17]) );
MUX2_X1 _u3_u1_U103  ( .A(slv0_din[18]), .B(slv0_pt_in[21]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[18]) );
MUX2_X1 _u3_u1_U102  ( .A(slv0_din[19]), .B(slv0_pt_in[22]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[19]) );
MUX2_X1 _u3_u1_U101  ( .A(slv0_din[1]), .B(slv0_pt_in[4]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[1]) );
MUX2_X1 _u3_u1_U100  ( .A(slv0_din[20]), .B(slv0_pt_in[23]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[20]) );
MUX2_X1 _u3_u1_U99  ( .A(slv0_din[21]), .B(slv0_pt_in[24]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[21]) );
MUX2_X1 _u3_u1_U98  ( .A(slv0_din[22]), .B(slv0_pt_in[25]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[22]) );
MUX2_X1 _u3_u1_U97  ( .A(slv0_din[23]), .B(slv0_pt_in[26]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[23]) );
MUX2_X1 _u3_u1_U96  ( .A(slv0_din[24]), .B(slv0_pt_in[27]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[24]) );
MUX2_X1 _u3_u1_U95  ( .A(slv0_din[25]), .B(slv0_pt_in[28]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[25]) );
MUX2_X1 _u3_u1_U94  ( .A(slv0_din[26]), .B(slv0_pt_in[29]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[26]) );
MUX2_X1 _u3_u1_U93  ( .A(slv0_din[27]), .B(slv0_pt_in[30]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[27]) );
MUX2_X1 _u3_u1_U92  ( .A(slv0_din[28]), .B(slv0_pt_in[31]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[28]) );
MUX2_X1 _u3_u1_U91  ( .A(slv0_din[29]), .B(slv0_pt_in[32]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[29]) );
MUX2_X1 _u3_u1_U90  ( .A(slv0_din[2]), .B(slv0_pt_in[5]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[2]) );
MUX2_X1 _u3_u1_U89  ( .A(slv0_din[30]), .B(slv0_pt_in[33]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[30]) );
MUX2_X1 _u3_u1_U88  ( .A(slv0_din[31]), .B(slv0_pt_in[34]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[31]) );
MUX2_X1 _u3_u1_U87  ( .A(slv0_din[3]), .B(slv0_pt_in[6]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[3]) );
MUX2_X1 _u3_u1_U86  ( .A(slv0_din[4]), .B(slv0_pt_in[7]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[4]) );
MUX2_X1 _u3_u1_U85  ( .A(slv0_din[5]), .B(slv0_pt_in[8]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[5]) );
MUX2_X1 _u3_u1_U84  ( .A(slv0_din[6]), .B(slv0_pt_in[9]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[6]) );
MUX2_X1 _u3_u1_U83  ( .A(slv0_din[7]), .B(slv0_pt_in[10]), .S(_u3_u1_n16 ),.Z(wb0m_data_o[7]) );
MUX2_X1 _u3_u1_U82  ( .A(slv0_din[8]), .B(slv0_pt_in[11]), .S(_u3_u1_n14 ),.Z(wb0m_data_o[8]) );
MUX2_X1 _u3_u1_U81  ( .A(slv0_din[9]), .B(slv0_pt_in[12]), .S(_u3_u1_n15 ),.Z(wb0m_data_o[9]) );
AND2_X1 _u3_u1_U80  ( .A1(slv0_pt_in[1]), .A2(_u3_u1_n14 ), .ZN(wb0_err_o));
AND2_X1 _u3_u1_U79  ( .A1(slv0_pt_in[0]), .A2(_u3_u1_n15 ), .ZN(wb0_rty_o));
CLKBUF_X2 _u3_u1_U78  ( .A(wb0_addr_i[31]), .Z(mast1_pt_in[38]) );
CLKBUF_X2 _u3_u1_U77  ( .A(wb0_addr_i[30]), .Z(mast1_pt_in[37]) );
CLKBUF_X2 _u3_u1_U76  ( .A(wb0_addr_i[29]), .Z(mast1_pt_in[36]) );
CLKBUF_X2 _u3_u1_U75  ( .A(wb0_addr_i[28]), .Z(mast1_pt_in[35]) );
CLKBUF_X2 _u3_u1_U74  ( .A(wb0_addr_i[27]), .Z(mast1_pt_in[34]) );
CLKBUF_X2 _u3_u1_U73  ( .A(wb0_addr_i[26]), .Z(mast1_pt_in[33]) );
CLKBUF_X2 _u3_u1_U72  ( .A(wb0_addr_i[25]), .Z(mast1_pt_in[32]) );
CLKBUF_X2 _u3_u1_U71  ( .A(wb0_addr_i[24]), .Z(mast1_pt_in[31]) );
CLKBUF_X2 _u3_u1_U70  ( .A(wb0_addr_i[23]), .Z(mast1_pt_in[30]) );
CLKBUF_X2 _u3_u1_U69  ( .A(wb0_addr_i[22]), .Z(mast1_pt_in[29]) );
CLKBUF_X2 _u3_u1_U68  ( .A(wb0_addr_i[21]), .Z(mast1_pt_in[28]) );
CLKBUF_X2 _u3_u1_U67  ( .A(wb0_addr_i[20]), .Z(mast1_pt_in[27]) );
CLKBUF_X2 _u3_u1_U66  ( .A(wb0_addr_i[19]), .Z(mast1_pt_in[26]) );
CLKBUF_X2 _u3_u1_U65  ( .A(wb0_addr_i[18]), .Z(mast1_pt_in[25]) );
CLKBUF_X2 _u3_u1_U64  ( .A(wb0_addr_i[17]), .Z(mast1_pt_in[24]) );
CLKBUF_X2 _u3_u1_U63  ( .A(wb0_addr_i[16]), .Z(mast1_pt_in[23]) );
CLKBUF_X2 _u3_u1_U62  ( .A(wb0_addr_i[15]), .Z(mast1_pt_in[22]) );
CLKBUF_X2 _u3_u1_U61  ( .A(wb0_addr_i[14]), .Z(mast1_pt_in[21]) );
CLKBUF_X2 _u3_u1_U60  ( .A(wb0_addr_i[13]), .Z(mast1_pt_in[20]) );
CLKBUF_X2 _u3_u1_U59  ( .A(wb0_addr_i[12]), .Z(mast1_pt_in[19]) );
CLKBUF_X2 _u3_u1_U58  ( .A(wb0_addr_i[11]), .Z(mast1_pt_in[18]) );
CLKBUF_X2 _u3_u1_U57  ( .A(wb0_addr_i[10]), .Z(mast1_pt_in[17]) );
CLKBUF_X2 _u3_u1_U56  ( .A(wb0_addr_i[9]), .Z(mast1_pt_in[16]) );
CLKBUF_X2 _u3_u1_U55  ( .A(wb0_addr_i[8]), .Z(mast1_pt_in[15]) );
CLKBUF_X2 _u3_u1_U54  ( .A(wb0_addr_i[7]), .Z(mast1_pt_in[14]) );
CLKBUF_X2 _u3_u1_U53  ( .A(wb0_addr_i[6]), .Z(mast1_pt_in[13]) );
CLKBUF_X2 _u3_u1_U52  ( .A(wb0_addr_i[5]), .Z(mast1_pt_in[12]) );
CLKBUF_X2 _u3_u1_U51  ( .A(wb0_addr_i[4]), .Z(mast1_pt_in[11]) );
CLKBUF_X2 _u3_u1_U50  ( .A(wb0_addr_i[3]), .Z(mast1_pt_in[10]) );
CLKBUF_X2 _u3_u1_U49  ( .A(wb0_addr_i[2]), .Z(mast1_pt_in[9]) );
CLKBUF_X2 _u3_u1_U48  ( .A(wb0_addr_i[1]), .Z(mast1_pt_in[8]) );
CLKBUF_X2 _u3_u1_U47  ( .A(wb0_addr_i[0]), .Z(mast1_pt_in[7]) );
CLKBUF_X2 _u3_u1_U46  ( .A(wb0_sel_i[3]), .Z(mast1_pt_in[6]) );
CLKBUF_X2 _u3_u1_U45  ( .A(wb0_sel_i[2]), .Z(mast1_pt_in[5]) );
CLKBUF_X2 _u3_u1_U44  ( .A(wb0_sel_i[1]), .Z(mast1_pt_in[4]) );
CLKBUF_X2 _u3_u1_U43  ( .A(wb0_sel_i[0]), .Z(mast1_pt_in[3]) );
CLKBUF_X2 _u3_u1_U42  ( .A(wb0_we_i), .Z(mast1_pt_in[2]) );
CLKBUF_X2 _u3_u1_U41  ( .A(wb0_cyc_i), .Z(mast1_pt_in[1]) );
CLKBUF_X2 _u3_u1_U40  ( .A(wb0_stb_i), .Z(mast1_pt_in[0]) );
CLKBUF_X2 _u3_u1_U39  ( .A(wb0m_data_i[31]), .Z(mast1_pt_in[70]) );
CLKBUF_X2 _u3_u1_U38  ( .A(wb0m_data_i[30]), .Z(mast1_pt_in[69]) );
CLKBUF_X2 _u3_u1_U37  ( .A(wb0m_data_i[29]), .Z(mast1_pt_in[68]) );
CLKBUF_X2 _u3_u1_U36  ( .A(wb0m_data_i[28]), .Z(mast1_pt_in[67]) );
CLKBUF_X2 _u3_u1_U35  ( .A(wb0m_data_i[27]), .Z(mast1_pt_in[66]) );
CLKBUF_X2 _u3_u1_U34  ( .A(wb0m_data_i[26]), .Z(mast1_pt_in[65]) );
CLKBUF_X2 _u3_u1_U33  ( .A(wb0m_data_i[25]), .Z(mast1_pt_in[64]) );
CLKBUF_X2 _u3_u1_U32  ( .A(wb0m_data_i[24]), .Z(mast1_pt_in[63]) );
CLKBUF_X2 _u3_u1_U31  ( .A(wb0m_data_i[23]), .Z(mast1_pt_in[62]) );
CLKBUF_X2 _u3_u1_U30  ( .A(wb0m_data_i[22]), .Z(mast1_pt_in[61]) );
CLKBUF_X2 _u3_u1_U29  ( .A(wb0m_data_i[21]), .Z(mast1_pt_in[60]) );
CLKBUF_X2 _u3_u1_U28  ( .A(wb0m_data_i[20]), .Z(mast1_pt_in[59]) );
CLKBUF_X2 _u3_u1_U27  ( .A(wb0m_data_i[19]), .Z(mast1_pt_in[58]) );
CLKBUF_X2 _u3_u1_U26  ( .A(wb0m_data_i[18]), .Z(mast1_pt_in[57]) );
CLKBUF_X2 _u3_u1_U25  ( .A(wb0m_data_i[17]), .Z(mast1_pt_in[56]) );
CLKBUF_X2 _u3_u1_U24  ( .A(wb0m_data_i[16]), .Z(mast1_pt_in[55]) );
CLKBUF_X2 _u3_u1_U23  ( .A(wb0m_data_i[15]), .Z(mast1_pt_in[54]) );
CLKBUF_X2 _u3_u1_U22  ( .A(wb0m_data_i[14]), .Z(mast1_pt_in[53]) );
CLKBUF_X2 _u3_u1_U21  ( .A(wb0m_data_i[13]), .Z(mast1_pt_in[52]) );
CLKBUF_X2 _u3_u1_U20  ( .A(wb0m_data_i[12]), .Z(mast1_pt_in[51]) );
CLKBUF_X2 _u3_u1_U19  ( .A(wb0m_data_i[11]), .Z(mast1_pt_in[50]) );
CLKBUF_X2 _u3_u1_U18  ( .A(wb0m_data_i[10]), .Z(mast1_pt_in[49]) );
CLKBUF_X2 _u3_u1_U17  ( .A(wb0m_data_i[9]), .Z(mast1_pt_in[48]) );
CLKBUF_X2 _u3_u1_U16  ( .A(wb0m_data_i[8]), .Z(mast1_pt_in[47]) );
CLKBUF_X2 _u3_u1_U15  ( .A(wb0m_data_i[7]), .Z(mast1_pt_in[46]) );
CLKBUF_X2 _u3_u1_U14  ( .A(wb0m_data_i[6]), .Z(mast1_pt_in[45]) );
CLKBUF_X2 _u3_u1_U13  ( .A(wb0m_data_i[5]), .Z(mast1_pt_in[44]) );
CLKBUF_X2 _u3_u1_U12  ( .A(wb0m_data_i[4]), .Z(mast1_pt_in[43]) );
CLKBUF_X2 _u3_u1_U11  ( .A(wb0m_data_i[3]), .Z(mast1_pt_in[42]) );
CLKBUF_X2 _u3_u1_U10  ( .A(wb0m_data_i[2]), .Z(mast1_pt_in[41]) );
CLKBUF_X2 _u3_u1_U9  ( .A(wb0m_data_i[1]), .Z(mast1_pt_in[40]) );
CLKBUF_X2 _u3_u1_U8  ( .A(wb0m_data_i[0]), .Z(mast1_pt_in[39]) );
INV_X1 _u3_u1_U7  ( .A(_u3_u1_n11 ), .ZN(_u3_u1_n16 ) );
INV_X1 _u3_u1_U6  ( .A(_u3_u1_n11 ), .ZN(_u3_u1_n15 ) );
INV_X1 _u3_u1_U5  ( .A(_u3_u1_n11 ), .ZN(_u3_u1_n14 ) );
INV_X8 _u3_u1_U4  ( .A(_u3_u1_n11 ), .ZN(pt1_sel_i) );
NAND2_X2 _u3_u1_U3  ( .A1(wb0_cyc_i), .A2(_u3_u1_n88 ), .ZN(_u3_u1_n11 ) );
DFF_X2 _u3_u1_slv_re_reg  ( .D(_u3_u1_N3 ), .CK(clk_i), .Q(slv0_re), .QN());
DFF_X2 _u3_u1_slv_we_reg  ( .D(_u3_u1_N4 ), .CK(clk_i), .Q(slv0_we), .QN());
DFF_X2 _u3_u1_rf_ack_reg  ( .D(_u3_u1_N5 ), .CK(clk_i), .Q(_u3_u1_rf_ack ),.QN(_u3_u1_n12 ) );
DFF_X2 _u3_u1_slv_dout_reg_0_  ( .D(wb0m_data_i[0]), .CK(clk_i), .Q(slv0_dout[0]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_1_  ( .D(wb0m_data_i[1]), .CK(clk_i), .Q(slv0_dout[1]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_2_  ( .D(wb0m_data_i[2]), .CK(clk_i), .Q(slv0_dout[2]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_3_  ( .D(wb0m_data_i[3]), .CK(clk_i), .Q(slv0_dout[3]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_4_  ( .D(wb0m_data_i[4]), .CK(clk_i), .Q(slv0_dout[4]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_5_  ( .D(wb0m_data_i[5]), .CK(clk_i), .Q(slv0_dout[5]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_6_  ( .D(wb0m_data_i[6]), .CK(clk_i), .Q(slv0_dout[6]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_7_  ( .D(wb0m_data_i[7]), .CK(clk_i), .Q(slv0_dout[7]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_8_  ( .D(wb0m_data_i[8]), .CK(clk_i), .Q(slv0_dout[8]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_9_  ( .D(wb0m_data_i[9]), .CK(clk_i), .Q(slv0_dout[9]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_10_  ( .D(wb0m_data_i[10]), .CK(clk_i), .Q(slv0_dout[10]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_11_  ( .D(wb0m_data_i[11]), .CK(clk_i), .Q(slv0_dout[11]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_12_  ( .D(wb0m_data_i[12]), .CK(clk_i), .Q(slv0_dout[12]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_13_  ( .D(wb0m_data_i[13]), .CK(clk_i), .Q(slv0_dout[13]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_14_  ( .D(wb0m_data_i[14]), .CK(clk_i), .Q(slv0_dout[14]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_15_  ( .D(wb0m_data_i[15]), .CK(clk_i), .Q(slv0_dout[15]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_16_  ( .D(wb0m_data_i[16]), .CK(clk_i), .Q(slv0_dout[16]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_17_  ( .D(wb0m_data_i[17]), .CK(clk_i), .Q(slv0_dout[17]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_18_  ( .D(wb0m_data_i[18]), .CK(clk_i), .Q(slv0_dout[18]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_19_  ( .D(wb0m_data_i[19]), .CK(clk_i), .Q(slv0_dout[19]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_20_  ( .D(wb0m_data_i[20]), .CK(clk_i), .Q(slv0_dout[20]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_21_  ( .D(wb0m_data_i[21]), .CK(clk_i), .Q(slv0_dout[21]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_22_  ( .D(wb0m_data_i[22]), .CK(clk_i), .Q(slv0_dout[22]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_23_  ( .D(wb0m_data_i[23]), .CK(clk_i), .Q(slv0_dout[23]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_24_  ( .D(wb0m_data_i[24]), .CK(clk_i), .Q(slv0_dout[24]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_25_  ( .D(wb0m_data_i[25]), .CK(clk_i), .Q(slv0_dout[25]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_26_  ( .D(wb0m_data_i[26]), .CK(clk_i), .Q(slv0_dout[26]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_27_  ( .D(wb0m_data_i[27]), .CK(clk_i), .Q(slv0_dout[27]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_28_  ( .D(wb0m_data_i[28]), .CK(clk_i), .Q(slv0_dout[28]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_29_  ( .D(wb0m_data_i[29]), .CK(clk_i), .Q(slv0_dout[29]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_30_  ( .D(wb0m_data_i[30]), .CK(clk_i), .Q(slv0_dout[30]), .QN() );
DFF_X2 _u3_u1_slv_dout_reg_31_  ( .D(wb0m_data_i[31]), .CK(clk_i), .Q(slv0_dout[31]), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_0_  ( .D(wb0_addr_i[0]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7886), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_1_  ( .D(wb0_addr_i[1]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7885), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_2_  ( .D(wb0_addr_i[2]), .CK(clk_i), .Q(slv0_adr[2]), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_3_  ( .D(wb0_addr_i[3]), .CK(clk_i), .Q(slv0_adr[3]), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_4_  ( .D(wb0_addr_i[4]), .CK(clk_i), .Q(slv0_adr[4]), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_5_  ( .D(wb0_addr_i[5]), .CK(clk_i), .Q(slv0_adr[5]), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_6_  ( .D(wb0_addr_i[6]), .CK(clk_i), .Q(slv0_adr[6]), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_7_  ( .D(wb0_addr_i[7]), .CK(clk_i), .Q(slv0_adr[7]), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_8_  ( .D(wb0_addr_i[8]), .CK(clk_i), .Q(slv0_adr[8]), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_9_  ( .D(wb0_addr_i[9]), .CK(clk_i), .Q(slv0_adr[9]), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_10_  ( .D(wb0_addr_i[10]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7884), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_11_  ( .D(wb0_addr_i[11]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7883), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_12_  ( .D(wb0_addr_i[12]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7882), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_13_  ( .D(wb0_addr_i[13]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7881), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_14_  ( .D(wb0_addr_i[14]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7880), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_15_  ( .D(wb0_addr_i[15]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7879), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_16_  ( .D(wb0_addr_i[16]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7878), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_17_  ( .D(wb0_addr_i[17]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7877), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_18_  ( .D(wb0_addr_i[18]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7876), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_19_  ( .D(wb0_addr_i[19]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7875), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_20_  ( .D(wb0_addr_i[20]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7874), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_21_  ( .D(wb0_addr_i[21]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7873), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_22_  ( .D(wb0_addr_i[22]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7872), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_23_  ( .D(wb0_addr_i[23]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7871), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_24_  ( .D(wb0_addr_i[24]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7870), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_25_  ( .D(wb0_addr_i[25]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7869), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_26_  ( .D(wb0_addr_i[26]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7868), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_27_  ( .D(wb0_addr_i[27]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7867), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_28_  ( .D(wb0_addr_i[28]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7866), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_29_  ( .D(wb0_addr_i[29]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7865), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_30_  ( .D(wb0_addr_i[30]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7864), .QN() );
DFF_X2 _u3_u1_slv_adr_reg_31_  ( .D(wb0_addr_i[31]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7863), .QN() );
INV_X1 _u40_u0_U146  ( .A(mast1_go), .ZN(_u40_u0_n74 ) );
NOR2_X1 _u40_u0_U145  ( .A1(mast1_wait), .A2(_u40_u0_n74 ), .ZN(_u40_u0_N3 ));
MUX2_X1 _u40_u0_U144  ( .A(mast1_dout[24]), .B(wb1s_data_i[24]), .S(wb1_ack_i), .Z(_u40_u0_n10 ) );
MUX2_X1 _u40_u0_U143  ( .A(mast1_dout[23]), .B(wb1s_data_i[23]), .S(wb1_ack_i), .Z(_u40_u0_n11 ) );
MUX2_X1 _u40_u0_U142  ( .A(mast1_dout[22]), .B(wb1s_data_i[22]), .S(wb1_ack_i), .Z(_u40_u0_n12 ) );
MUX2_X1 _u40_u0_U141  ( .A(mast1_dout[21]), .B(wb1s_data_i[21]), .S(wb1_ack_i), .Z(_u40_u0_n13 ) );
MUX2_X1 _u40_u0_U140  ( .A(mast1_dout[20]), .B(wb1s_data_i[20]), .S(wb1_ack_i), .Z(_u40_u0_n14 ) );
MUX2_X1 _u40_u0_U139  ( .A(mast1_dout[19]), .B(wb1s_data_i[19]), .S(wb1_ack_i), .Z(_u40_u0_n15 ) );
MUX2_X1 _u40_u0_U138  ( .A(mast1_dout[18]), .B(wb1s_data_i[18]), .S(wb1_ack_i), .Z(_u40_u0_n16 ) );
MUX2_X1 _u40_u0_U137  ( .A(mast1_dout[17]), .B(wb1s_data_i[17]), .S(wb1_ack_i), .Z(_u40_u0_n17 ) );
MUX2_X1 _u40_u0_U136  ( .A(mast1_dout[16]), .B(wb1s_data_i[16]), .S(wb1_ack_i), .Z(_u40_u0_n18 ) );
MUX2_X1 _u40_u0_U135  ( .A(mast1_dout[15]), .B(wb1s_data_i[15]), .S(wb1_ack_i), .Z(_u40_u0_n19 ) );
MUX2_X1 _u40_u0_U134  ( .A(mast1_dout[14]), .B(wb1s_data_i[14]), .S(wb1_ack_i), .Z(_u40_u0_n20 ) );
MUX2_X1 _u40_u0_U133  ( .A(mast1_dout[13]), .B(wb1s_data_i[13]), .S(wb1_ack_i), .Z(_u40_u0_n21 ) );
MUX2_X1 _u40_u0_U132  ( .A(mast1_dout[12]), .B(wb1s_data_i[12]), .S(wb1_ack_i), .Z(_u40_u0_n22 ) );
MUX2_X1 _u40_u0_U131  ( .A(mast1_dout[11]), .B(wb1s_data_i[11]), .S(wb1_ack_i), .Z(_u40_u0_n23 ) );
MUX2_X1 _u40_u0_U130  ( .A(mast1_dout[10]), .B(wb1s_data_i[10]), .S(wb1_ack_i), .Z(_u40_u0_n24 ) );
MUX2_X1 _u40_u0_U129  ( .A(mast1_dout[9]), .B(wb1s_data_i[9]), .S(wb1_ack_i),.Z(_u40_u0_n25 ) );
MUX2_X1 _u40_u0_U128  ( .A(mast1_dout[8]), .B(wb1s_data_i[8]), .S(wb1_ack_i),.Z(_u40_u0_n26 ) );
MUX2_X1 _u40_u0_U127  ( .A(mast1_dout[7]), .B(wb1s_data_i[7]), .S(wb1_ack_i),.Z(_u40_u0_n27 ) );
MUX2_X1 _u40_u0_U126  ( .A(mast1_dout[6]), .B(wb1s_data_i[6]), .S(wb1_ack_i),.Z(_u40_u0_n28 ) );
MUX2_X1 _u40_u0_U125  ( .A(mast1_dout[5]), .B(wb1s_data_i[5]), .S(wb1_ack_i),.Z(_u40_u0_n29 ) );
MUX2_X1 _u40_u0_U124  ( .A(mast1_dout[31]), .B(wb1s_data_i[31]), .S(wb1_ack_i), .Z(_u40_u0_n300 ) );
MUX2_X1 _u40_u0_U123  ( .A(mast1_dout[4]), .B(wb1s_data_i[4]), .S(wb1_ack_i),.Z(_u40_u0_n301 ) );
MUX2_X1 _u40_u0_U122  ( .A(mast1_dout[3]), .B(wb1s_data_i[3]), .S(wb1_ack_i),.Z(_u40_u0_n31 ) );
MUX2_X1 _u40_u0_U121  ( .A(mast1_dout[2]), .B(wb1s_data_i[2]), .S(wb1_ack_i),.Z(_u40_u0_n32 ) );
MUX2_X1 _u40_u0_U120  ( .A(mast1_dout[1]), .B(wb1s_data_i[1]), .S(wb1_ack_i),.Z(_u40_u0_n33 ) );
MUX2_X1 _u40_u0_U119  ( .A(mast1_dout[0]), .B(wb1s_data_i[0]), .S(wb1_ack_i),.Z(_u40_u0_n34 ) );
MUX2_X1 _u40_u0_U118  ( .A(mast1_dout[30]), .B(wb1s_data_i[30]), .S(wb1_ack_i), .Z(_u40_u0_n4 ) );
MUX2_X1 _u40_u0_U117  ( .A(mast1_dout[29]), .B(wb1s_data_i[29]), .S(wb1_ack_i), .Z(_u40_u0_n5 ) );
MUX2_X1 _u40_u0_U116  ( .A(mast1_dout[28]), .B(wb1s_data_i[28]), .S(wb1_ack_i), .Z(_u40_u0_n6 ) );
MUX2_X1 _u40_u0_U115  ( .A(mast1_dout[27]), .B(wb1s_data_i[27]), .S(wb1_ack_i), .Z(_u40_u0_n7 ) );
MUX2_X1 _u40_u0_U114  ( .A(mast1_dout[26]), .B(wb1s_data_i[26]), .S(wb1_ack_i), .Z(_u40_u0_n8 ) );
MUX2_X1 _u40_u0_U113  ( .A(mast1_dout[25]), .B(wb1s_data_i[25]), .S(wb1_ack_i), .Z(_u40_u0_n9 ) );
MUX2_X1 _u40_u0_U112  ( .A(1'b0), .B(mast1_pt_in[7]), .S(pt1_sel_i), .Z(wb1_addr_o[0]) );
MUX2_X1 _u40_u0_U111  ( .A(mast1_adr[10]), .B(mast1_pt_in[17]), .S(pt1_sel_i), .Z(wb1_addr_o[10]) );
MUX2_X1 _u40_u0_U110  ( .A(mast1_adr[11]), .B(mast1_pt_in[18]), .S(pt1_sel_i), .Z(wb1_addr_o[11]) );
MUX2_X1 _u40_u0_U109  ( .A(mast1_adr[12]), .B(mast1_pt_in[19]), .S(pt1_sel_i), .Z(wb1_addr_o[12]) );
MUX2_X1 _u40_u0_U108  ( .A(mast1_adr[13]), .B(mast1_pt_in[20]), .S(pt1_sel_i), .Z(wb1_addr_o[13]) );
MUX2_X1 _u40_u0_U107  ( .A(mast1_adr[14]), .B(mast1_pt_in[21]), .S(pt1_sel_i), .Z(wb1_addr_o[14]) );
MUX2_X1 _u40_u0_U106  ( .A(mast1_adr[15]), .B(mast1_pt_in[22]), .S(pt1_sel_i), .Z(wb1_addr_o[15]) );
MUX2_X1 _u40_u0_U105  ( .A(mast1_adr[16]), .B(mast1_pt_in[23]), .S(pt1_sel_i), .Z(wb1_addr_o[16]) );
MUX2_X1 _u40_u0_U104  ( .A(mast1_adr[17]), .B(mast1_pt_in[24]), .S(pt1_sel_i), .Z(wb1_addr_o[17]) );
MUX2_X1 _u40_u0_U103  ( .A(mast1_adr[18]), .B(mast1_pt_in[25]), .S(pt1_sel_i), .Z(wb1_addr_o[18]) );
MUX2_X1 _u40_u0_U102  ( .A(mast1_adr[19]), .B(mast1_pt_in[26]), .S(pt1_sel_i), .Z(wb1_addr_o[19]) );
MUX2_X1 _u40_u0_U101  ( .A(1'b0), .B(mast1_pt_in[8]), .S(pt1_sel_i), .Z(wb1_addr_o[1]) );
MUX2_X1 _u40_u0_U100  ( .A(mast1_adr[20]), .B(mast1_pt_in[27]), .S(pt1_sel_i), .Z(wb1_addr_o[20]) );
MUX2_X1 _u40_u0_U99  ( .A(mast1_adr[21]), .B(mast1_pt_in[28]), .S(pt1_sel_i),.Z(wb1_addr_o[21]) );
MUX2_X1 _u40_u0_U98  ( .A(mast1_adr[22]), .B(mast1_pt_in[29]), .S(pt1_sel_i),.Z(wb1_addr_o[22]) );
MUX2_X1 _u40_u0_U97  ( .A(mast1_adr[23]), .B(mast1_pt_in[30]), .S(pt1_sel_i),.Z(wb1_addr_o[23]) );
MUX2_X1 _u40_u0_U96  ( .A(mast1_adr[24]), .B(mast1_pt_in[31]), .S(pt1_sel_i),.Z(wb1_addr_o[24]) );
MUX2_X1 _u40_u0_U95  ( .A(mast1_adr[25]), .B(mast1_pt_in[32]), .S(pt1_sel_i),.Z(wb1_addr_o[25]) );
MUX2_X1 _u40_u0_U94  ( .A(mast1_adr[26]), .B(mast1_pt_in[33]), .S(pt1_sel_i),.Z(wb1_addr_o[26]) );
MUX2_X1 _u40_u0_U93  ( .A(mast1_adr[27]), .B(mast1_pt_in[34]), .S(pt1_sel_i),.Z(wb1_addr_o[27]) );
MUX2_X1 _u40_u0_U92  ( .A(mast1_adr[28]), .B(mast1_pt_in[35]), .S(pt1_sel_i),.Z(wb1_addr_o[28]) );
MUX2_X1 _u40_u0_U91  ( .A(mast1_adr[29]), .B(mast1_pt_in[36]), .S(pt1_sel_i),.Z(wb1_addr_o[29]) );
MUX2_X1 _u40_u0_U90  ( .A(mast1_adr[2]), .B(mast1_pt_in[9]), .S(pt1_sel_i),.Z(wb1_addr_o[2]) );
MUX2_X1 _u40_u0_U89  ( .A(mast1_adr[30]), .B(mast1_pt_in[37]), .S(pt1_sel_i),.Z(wb1_addr_o[30]) );
MUX2_X1 _u40_u0_U88  ( .A(mast1_adr[31]), .B(mast1_pt_in[38]), .S(pt1_sel_i),.Z(wb1_addr_o[31]) );
MUX2_X1 _u40_u0_U87  ( .A(mast1_adr[3]), .B(mast1_pt_in[10]), .S(pt1_sel_i),.Z(wb1_addr_o[3]) );
MUX2_X1 _u40_u0_U86  ( .A(mast1_adr[4]), .B(mast1_pt_in[11]), .S(pt1_sel_i),.Z(wb1_addr_o[4]) );
MUX2_X1 _u40_u0_U85  ( .A(mast1_adr[5]), .B(mast1_pt_in[12]), .S(pt1_sel_i),.Z(wb1_addr_o[5]) );
MUX2_X1 _u40_u0_U84  ( .A(mast1_adr[6]), .B(mast1_pt_in[13]), .S(pt1_sel_i),.Z(wb1_addr_o[6]) );
MUX2_X1 _u40_u0_U83  ( .A(mast1_adr[7]), .B(mast1_pt_in[14]), .S(pt1_sel_i),.Z(wb1_addr_o[7]) );
MUX2_X1 _u40_u0_U82  ( .A(mast1_adr[8]), .B(mast1_pt_in[15]), .S(pt1_sel_i),.Z(wb1_addr_o[8]) );
MUX2_X1 _u40_u0_U81  ( .A(mast1_adr[9]), .B(mast1_pt_in[16]), .S(pt1_sel_i),.Z(wb1_addr_o[9]) );
MUX2_X1 _u40_u0_U80  ( .A(_u40_u0_mast_cyc ), .B(mast1_pt_in[1]), .S(pt1_sel_i), .Z(wb1_cyc_o) );
MUX2_X1 _u40_u0_U79  ( .A(mast1_din[0]), .B(mast1_pt_in[39]), .S(pt1_sel_i),.Z(wb1s_data_o[0]) );
MUX2_X1 _u40_u0_U78  ( .A(mast1_din[10]), .B(mast1_pt_in[49]), .S(pt1_sel_i),.Z(wb1s_data_o[10]) );
MUX2_X1 _u40_u0_U77  ( .A(mast1_din[11]), .B(mast1_pt_in[50]), .S(pt1_sel_i),.Z(wb1s_data_o[11]) );
MUX2_X1 _u40_u0_U76  ( .A(mast1_din[12]), .B(mast1_pt_in[51]), .S(pt1_sel_i),.Z(wb1s_data_o[12]) );
MUX2_X1 _u40_u0_U75  ( .A(mast1_din[13]), .B(mast1_pt_in[52]), .S(pt1_sel_i),.Z(wb1s_data_o[13]) );
MUX2_X1 _u40_u0_U74  ( .A(mast1_din[14]), .B(mast1_pt_in[53]), .S(pt1_sel_i),.Z(wb1s_data_o[14]) );
MUX2_X1 _u40_u0_U73  ( .A(mast1_din[15]), .B(mast1_pt_in[54]), .S(pt1_sel_i),.Z(wb1s_data_o[15]) );
MUX2_X1 _u40_u0_U72  ( .A(mast1_din[16]), .B(mast1_pt_in[55]), .S(pt1_sel_i),.Z(wb1s_data_o[16]) );
MUX2_X1 _u40_u0_U71  ( .A(mast1_din[17]), .B(mast1_pt_in[56]), .S(pt1_sel_i),.Z(wb1s_data_o[17]) );
MUX2_X1 _u40_u0_U70  ( .A(mast1_din[18]), .B(mast1_pt_in[57]), .S(pt1_sel_i),.Z(wb1s_data_o[18]) );
MUX2_X1 _u40_u0_U69  ( .A(mast1_din[19]), .B(mast1_pt_in[58]), .S(pt1_sel_i),.Z(wb1s_data_o[19]) );
MUX2_X1 _u40_u0_U68  ( .A(mast1_din[1]), .B(mast1_pt_in[40]), .S(pt1_sel_i),.Z(wb1s_data_o[1]) );
MUX2_X1 _u40_u0_U67  ( .A(mast1_din[20]), .B(mast1_pt_in[59]), .S(pt1_sel_i),.Z(wb1s_data_o[20]) );
MUX2_X1 _u40_u0_U66  ( .A(mast1_din[21]), .B(mast1_pt_in[60]), .S(pt1_sel_i),.Z(wb1s_data_o[21]) );
MUX2_X1 _u40_u0_U65  ( .A(mast1_din[22]), .B(mast1_pt_in[61]), .S(pt1_sel_i),.Z(wb1s_data_o[22]) );
MUX2_X1 _u40_u0_U64  ( .A(mast1_din[23]), .B(mast1_pt_in[62]), .S(pt1_sel_i),.Z(wb1s_data_o[23]) );
MUX2_X1 _u40_u0_U63  ( .A(mast1_din[24]), .B(mast1_pt_in[63]), .S(pt1_sel_i),.Z(wb1s_data_o[24]) );
MUX2_X1 _u40_u0_U62  ( .A(mast1_din[25]), .B(mast1_pt_in[64]), .S(pt1_sel_i),.Z(wb1s_data_o[25]) );
MUX2_X1 _u40_u0_U61  ( .A(mast1_din[26]), .B(mast1_pt_in[65]), .S(pt1_sel_i),.Z(wb1s_data_o[26]) );
MUX2_X1 _u40_u0_U60  ( .A(mast1_din[27]), .B(mast1_pt_in[66]), .S(pt1_sel_i),.Z(wb1s_data_o[27]) );
MUX2_X1 _u40_u0_U59  ( .A(mast1_din[28]), .B(mast1_pt_in[67]), .S(pt1_sel_i),.Z(wb1s_data_o[28]) );
MUX2_X1 _u40_u0_U58  ( .A(mast1_din[29]), .B(mast1_pt_in[68]), .S(pt1_sel_i),.Z(wb1s_data_o[29]) );
MUX2_X1 _u40_u0_U57  ( .A(mast1_din[2]), .B(mast1_pt_in[41]), .S(pt1_sel_i),.Z(wb1s_data_o[2]) );
MUX2_X1 _u40_u0_U56  ( .A(mast1_din[30]), .B(mast1_pt_in[69]), .S(pt1_sel_i),.Z(wb1s_data_o[30]) );
MUX2_X1 _u40_u0_U55  ( .A(mast1_din[31]), .B(mast1_pt_in[70]), .S(pt1_sel_i),.Z(wb1s_data_o[31]) );
MUX2_X1 _u40_u0_U54  ( .A(mast1_din[3]), .B(mast1_pt_in[42]), .S(pt1_sel_i),.Z(wb1s_data_o[3]) );
MUX2_X1 _u40_u0_U53  ( .A(mast1_din[4]), .B(mast1_pt_in[43]), .S(pt1_sel_i),.Z(wb1s_data_o[4]) );
MUX2_X1 _u40_u0_U52  ( .A(mast1_din[5]), .B(mast1_pt_in[44]), .S(pt1_sel_i),.Z(wb1s_data_o[5]) );
MUX2_X1 _u40_u0_U51  ( .A(mast1_din[6]), .B(mast1_pt_in[45]), .S(pt1_sel_i),.Z(wb1s_data_o[6]) );
MUX2_X1 _u40_u0_U50  ( .A(mast1_din[7]), .B(mast1_pt_in[46]), .S(pt1_sel_i),.Z(wb1s_data_o[7]) );
MUX2_X1 _u40_u0_U49  ( .A(mast1_din[8]), .B(mast1_pt_in[47]), .S(pt1_sel_i),.Z(wb1s_data_o[8]) );
MUX2_X1 _u40_u0_U48  ( .A(mast1_din[9]), .B(mast1_pt_in[48]), .S(pt1_sel_i),.Z(wb1s_data_o[9]) );
INV_X1 _u40_u0_U47  ( .A(pt1_sel_i), .ZN(_u40_u0_n73 ) );
OR2_X1 _u40_u0_U46  ( .A1(mast1_pt_in[3]), .A2(_u40_u0_n73 ), .ZN(wb1_sel_o[0]) );
OR2_X1 _u40_u0_U45  ( .A1(mast1_pt_in[4]), .A2(_u40_u0_n73 ), .ZN(wb1_sel_o[1]) );
OR2_X1 _u40_u0_U44  ( .A1(mast1_pt_in[5]), .A2(_u40_u0_n73 ), .ZN(wb1_sel_o[2]) );
OR2_X1 _u40_u0_U43  ( .A1(mast1_pt_in[6]), .A2(_u40_u0_n73 ), .ZN(wb1_sel_o[3]) );
MUX2_X1 _u40_u0_U42  ( .A(_u40_u0_mast_stb ), .B(mast1_pt_in[0]), .S(pt1_sel_i), .Z(wb1_stb_o) );
MUX2_X1 _u40_u0_U41  ( .A(_u40_u0_mast_we_r ), .B(mast1_pt_in[2]), .S(pt1_sel_i), .Z(wb1_we_o) );
CLKBUF_X2 _u40_u0_U40  ( .A(wb1s_data_i[31]), .Z(slv0_pt_in[34]) );
CLKBUF_X2 _u40_u0_U39  ( .A(wb1s_data_i[30]), .Z(slv0_pt_in[33]) );
CLKBUF_X2 _u40_u0_U38  ( .A(wb1s_data_i[29]), .Z(slv0_pt_in[32]) );
CLKBUF_X2 _u40_u0_U37  ( .A(wb1s_data_i[28]), .Z(slv0_pt_in[31]) );
CLKBUF_X2 _u40_u0_U36  ( .A(wb1s_data_i[27]), .Z(slv0_pt_in[30]) );
CLKBUF_X2 _u40_u0_U35  ( .A(wb1s_data_i[26]), .Z(slv0_pt_in[29]) );
CLKBUF_X2 _u40_u0_U34  ( .A(wb1s_data_i[25]), .Z(slv0_pt_in[28]) );
CLKBUF_X2 _u40_u0_U33  ( .A(wb1s_data_i[24]), .Z(slv0_pt_in[27]) );
CLKBUF_X2 _u40_u0_U32  ( .A(wb1s_data_i[23]), .Z(slv0_pt_in[26]) );
CLKBUF_X2 _u40_u0_U31  ( .A(wb1s_data_i[22]), .Z(slv0_pt_in[25]) );
CLKBUF_X2 _u40_u0_U30  ( .A(wb1s_data_i[21]), .Z(slv0_pt_in[24]) );
CLKBUF_X2 _u40_u0_U29  ( .A(wb1s_data_i[20]), .Z(slv0_pt_in[23]) );
CLKBUF_X2 _u40_u0_U28  ( .A(wb1s_data_i[19]), .Z(slv0_pt_in[22]) );
CLKBUF_X2 _u40_u0_U27  ( .A(wb1s_data_i[18]), .Z(slv0_pt_in[21]) );
CLKBUF_X2 _u40_u0_U26  ( .A(wb1s_data_i[17]), .Z(slv0_pt_in[20]) );
CLKBUF_X2 _u40_u0_U25  ( .A(wb1s_data_i[16]), .Z(slv0_pt_in[19]) );
CLKBUF_X2 _u40_u0_U24  ( .A(wb1s_data_i[15]), .Z(slv0_pt_in[18]) );
CLKBUF_X2 _u40_u0_U23  ( .A(wb1s_data_i[14]), .Z(slv0_pt_in[17]) );
CLKBUF_X2 _u40_u0_U22  ( .A(wb1s_data_i[13]), .Z(slv0_pt_in[16]) );
CLKBUF_X2 _u40_u0_U21  ( .A(wb1s_data_i[12]), .Z(slv0_pt_in[15]) );
CLKBUF_X2 _u40_u0_U20  ( .A(wb1s_data_i[11]), .Z(slv0_pt_in[14]) );
CLKBUF_X2 _u40_u0_U19  ( .A(wb1s_data_i[10]), .Z(slv0_pt_in[13]) );
CLKBUF_X2 _u40_u0_U18  ( .A(wb1s_data_i[9]), .Z(slv0_pt_in[12]) );
CLKBUF_X2 _u40_u0_U17  ( .A(wb1s_data_i[8]), .Z(slv0_pt_in[11]) );
CLKBUF_X2 _u40_u0_U16  ( .A(wb1s_data_i[7]), .Z(slv0_pt_in[10]) );
CLKBUF_X2 _u40_u0_U15  ( .A(wb1s_data_i[6]), .Z(slv0_pt_in[9]) );
CLKBUF_X2 _u40_u0_U14  ( .A(wb1s_data_i[5]), .Z(slv0_pt_in[8]) );
CLKBUF_X2 _u40_u0_U13  ( .A(wb1s_data_i[4]), .Z(slv0_pt_in[7]) );
CLKBUF_X2 _u40_u0_U12  ( .A(wb1s_data_i[3]), .Z(slv0_pt_in[6]) );
CLKBUF_X2 _u40_u0_U11  ( .A(wb1s_data_i[2]), .Z(slv0_pt_in[5]) );
CLKBUF_X2 _u40_u0_U10  ( .A(wb1s_data_i[1]), .Z(slv0_pt_in[4]) );
CLKBUF_X2 _u40_u0_U9  ( .A(wb1s_data_i[0]), .Z(slv0_pt_in[3]) );
INV_X4 _u40_u0_U8  ( .A(_u40_u0_n38 ), .ZN(slv0_pt_in[2]) );
INV_X4 _u40_u0_U7  ( .A(_u40_u0_n38 ), .ZN(mast1_drdy) );
INV_X4 _u40_u0_U6  ( .A(wb1_ack_i), .ZN(_u40_u0_n38 ) );
CLKBUF_X2 _u40_u0_U5  ( .A(wb1_err_i), .Z(slv0_pt_in[1]) );
CLKBUF_X2 _u40_u0_U4  ( .A(wb1_err_i), .Z(mast1_err) );
CLKBUF_X2 _u40_u0_U3  ( .A(wb1_rty_i), .Z(slv0_pt_in[0]) );
DFF_X2 _u40_u0_mast_stb_reg  ( .D(_u40_u0_N3 ), .CK(clk_i), .Q(_u40_u0_mast_stb ), .QN() );
DFF_X2 _u40_u0_mast_cyc_reg  ( .D(mast1_go), .CK(clk_i), .Q(_u40_u0_mast_cyc ), .QN() );
DFF_X2 _u40_u0_mast_we_r_reg  ( .D(mast1_we), .CK(clk_i), .Q(_u40_u0_mast_we_r ), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_0_  ( .D(_u40_u0_n34 ), .CK(clk_i), .Q(mast1_dout[0]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_1_  ( .D(_u40_u0_n33 ), .CK(clk_i), .Q(mast1_dout[1]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_2_  ( .D(_u40_u0_n32 ), .CK(clk_i), .Q(mast1_dout[2]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_3_  ( .D(_u40_u0_n31 ), .CK(clk_i), .Q(mast1_dout[3]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_4_  ( .D(_u40_u0_n301 ), .CK(clk_i), .Q(mast1_dout[4]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_5_  ( .D(_u40_u0_n29 ), .CK(clk_i), .Q(mast1_dout[5]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_6_  ( .D(_u40_u0_n28 ), .CK(clk_i), .Q(mast1_dout[6]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_7_  ( .D(_u40_u0_n27 ), .CK(clk_i), .Q(mast1_dout[7]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_8_  ( .D(_u40_u0_n26 ), .CK(clk_i), .Q(mast1_dout[8]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_9_  ( .D(_u40_u0_n25 ), .CK(clk_i), .Q(mast1_dout[9]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_10_  ( .D(_u40_u0_n24 ), .CK(clk_i), .Q(mast1_dout[10]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_11_  ( .D(_u40_u0_n23 ), .CK(clk_i), .Q(mast1_dout[11]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_12_  ( .D(_u40_u0_n22 ), .CK(clk_i), .Q(mast1_dout[12]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_13_  ( .D(_u40_u0_n21 ), .CK(clk_i), .Q(mast1_dout[13]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_14_  ( .D(_u40_u0_n20 ), .CK(clk_i), .Q(mast1_dout[14]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_15_  ( .D(_u40_u0_n19 ), .CK(clk_i), .Q(mast1_dout[15]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_16_  ( .D(_u40_u0_n18 ), .CK(clk_i), .Q(mast1_dout[16]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_17_  ( .D(_u40_u0_n17 ), .CK(clk_i), .Q(mast1_dout[17]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_18_  ( .D(_u40_u0_n16 ), .CK(clk_i), .Q(mast1_dout[18]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_19_  ( .D(_u40_u0_n15 ), .CK(clk_i), .Q(mast1_dout[19]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_20_  ( .D(_u40_u0_n14 ), .CK(clk_i), .Q(mast1_dout[20]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_21_  ( .D(_u40_u0_n13 ), .CK(clk_i), .Q(mast1_dout[21]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_22_  ( .D(_u40_u0_n12 ), .CK(clk_i), .Q(mast1_dout[22]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_23_  ( .D(_u40_u0_n11 ), .CK(clk_i), .Q(mast1_dout[23]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_24_  ( .D(_u40_u0_n10 ), .CK(clk_i), .Q(mast1_dout[24]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_25_  ( .D(_u40_u0_n9 ), .CK(clk_i), .Q(mast1_dout[25]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_26_  ( .D(_u40_u0_n8 ), .CK(clk_i), .Q(mast1_dout[26]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_27_  ( .D(_u40_u0_n7 ), .CK(clk_i), .Q(mast1_dout[27]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_28_  ( .D(_u40_u0_n6 ), .CK(clk_i), .Q(mast1_dout[28]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_29_  ( .D(_u40_u0_n5 ), .CK(clk_i), .Q(mast1_dout[29]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_30_  ( .D(_u40_u0_n4 ), .CK(clk_i), .Q(mast1_dout[30]), .QN() );
DFF_X2 _u40_u0_mast_dout_reg_31_  ( .D(_u40_u0_n300 ), .CK(clk_i), .Q(mast1_dout[31]), .QN() );
NAND3_X1 _u40_u1_U120  ( .A1(wb1_cyc_i), .A2(_u40_u1_n12 ), .A3(wb1_stb_i),.ZN(_u40_u1_n90 ) );
OR4_X1 _u40_u1_U119  ( .A1(wb1_addr_i[29]), .A2(wb1_addr_i[28]), .A3(wb1_addr_i[31]), .A4(wb1_addr_i[30]), .ZN(_u40_u1_n88 ) );
NOR4_X1 _u40_u1_U118  ( .A1(wb1_we_i), .A2(_u40_slv_re ), .A3(_u40_u1_n90 ),.A4(_u40_u1_n88 ), .ZN(_u40_u1_N3 ) );
INV_X1 _u40_u1_U117  ( .A(wb1_we_i), .ZN(_u40_u1_n91 ) );
NOR3_X1 _u40_u1_U116  ( .A1(_u40_u1_n91 ), .A2(_u40_u1_n90 ), .A3(_u40_u1_n88 ), .ZN(_u40_u1_N4 ) );
NOR2_X1 _u40_u1_U115  ( .A1(_u40_slv_re ), .A2(_u40_slv_we ), .ZN(_u40_u1_n89 ) );
NOR2_X1 _u40_u1_U114  ( .A1(_u40_u1_n89 ), .A2(_u40_u1_n90 ), .ZN(_u40_u1_N5 ) );
MUX2_X1 _u40_u1_U113  ( .A(_u40_u1_rf_ack ), .B(slv1_pt_in[2]), .S(_u40_u1_n16 ), .Z(wb1_ack_o) );
MUX2_X1 _u40_u1_U112  ( .A(1'b0), .B(slv1_pt_in[3]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[0]) );
MUX2_X1 _u40_u1_U111  ( .A(1'b0), .B(slv1_pt_in[13]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[10]) );
MUX2_X1 _u40_u1_U110  ( .A(1'b0), .B(slv1_pt_in[14]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[11]) );
MUX2_X1 _u40_u1_U109  ( .A(1'b0), .B(slv1_pt_in[15]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[12]) );
MUX2_X1 _u40_u1_U108  ( .A(1'b0), .B(slv1_pt_in[16]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[13]) );
MUX2_X1 _u40_u1_U107  ( .A(1'b0), .B(slv1_pt_in[17]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[14]) );
MUX2_X1 _u40_u1_U106  ( .A(1'b0), .B(slv1_pt_in[18]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[15]) );
MUX2_X1 _u40_u1_U105  ( .A(1'b0), .B(slv1_pt_in[19]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[16]) );
MUX2_X1 _u40_u1_U104  ( .A(1'b0), .B(slv1_pt_in[20]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[17]) );
MUX2_X1 _u40_u1_U103  ( .A(1'b0), .B(slv1_pt_in[21]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[18]) );
MUX2_X1 _u40_u1_U102  ( .A(1'b0), .B(slv1_pt_in[22]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[19]) );
MUX2_X1 _u40_u1_U101  ( .A(1'b0), .B(slv1_pt_in[4]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[1]) );
MUX2_X1 _u40_u1_U100  ( .A(1'b0), .B(slv1_pt_in[23]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[20]) );
MUX2_X1 _u40_u1_U99  ( .A(1'b0), .B(slv1_pt_in[24]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[21]) );
MUX2_X1 _u40_u1_U98  ( .A(1'b0), .B(slv1_pt_in[25]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[22]) );
MUX2_X1 _u40_u1_U97  ( .A(1'b0), .B(slv1_pt_in[26]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[23]) );
MUX2_X1 _u40_u1_U96  ( .A(1'b0), .B(slv1_pt_in[27]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[24]) );
MUX2_X1 _u40_u1_U95  ( .A(1'b0), .B(slv1_pt_in[28]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[25]) );
MUX2_X1 _u40_u1_U94  ( .A(1'b0), .B(slv1_pt_in[29]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[26]) );
MUX2_X1 _u40_u1_U93  ( .A(1'b0), .B(slv1_pt_in[30]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[27]) );
MUX2_X1 _u40_u1_U92  ( .A(1'b0), .B(slv1_pt_in[31]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[28]) );
MUX2_X1 _u40_u1_U91  ( .A(1'b0), .B(slv1_pt_in[32]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[29]) );
MUX2_X1 _u40_u1_U90  ( .A(1'b0), .B(slv1_pt_in[5]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[2]) );
MUX2_X1 _u40_u1_U89  ( .A(1'b0), .B(slv1_pt_in[33]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[30]) );
MUX2_X1 _u40_u1_U88  ( .A(1'b0), .B(slv1_pt_in[34]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[31]) );
MUX2_X1 _u40_u1_U87  ( .A(1'b0), .B(slv1_pt_in[6]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[3]) );
MUX2_X1 _u40_u1_U86  ( .A(1'b0), .B(slv1_pt_in[7]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[4]) );
MUX2_X1 _u40_u1_U85  ( .A(1'b0), .B(slv1_pt_in[8]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[5]) );
MUX2_X1 _u40_u1_U84  ( .A(1'b0), .B(slv1_pt_in[9]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[6]) );
MUX2_X1 _u40_u1_U83  ( .A(1'b0), .B(slv1_pt_in[10]), .S(_u40_u1_n16 ), .Z(wb1m_data_o[7]) );
MUX2_X1 _u40_u1_U82  ( .A(1'b0), .B(slv1_pt_in[11]), .S(_u40_u1_n14 ), .Z(wb1m_data_o[8]) );
MUX2_X1 _u40_u1_U81  ( .A(1'b0), .B(slv1_pt_in[12]), .S(_u40_u1_n15 ), .Z(wb1m_data_o[9]) );
AND2_X1 _u40_u1_U80  ( .A1(slv1_pt_in[1]), .A2(_u40_u1_n14 ), .ZN(wb1_err_o));
AND2_X1 _u40_u1_U79  ( .A1(slv1_pt_in[0]), .A2(_u40_u1_n15 ), .ZN(wb1_rty_o));
CLKBUF_X2 _u40_u1_U78  ( .A(wb1_addr_i[31]), .Z(mast0_pt_in[38]) );
CLKBUF_X2 _u40_u1_U77  ( .A(wb1_addr_i[30]), .Z(mast0_pt_in[37]) );
CLKBUF_X2 _u40_u1_U76  ( .A(wb1_addr_i[29]), .Z(mast0_pt_in[36]) );
CLKBUF_X2 _u40_u1_U75  ( .A(wb1_addr_i[28]), .Z(mast0_pt_in[35]) );
CLKBUF_X2 _u40_u1_U74  ( .A(wb1_addr_i[27]), .Z(mast0_pt_in[34]) );
CLKBUF_X2 _u40_u1_U73  ( .A(wb1_addr_i[26]), .Z(mast0_pt_in[33]) );
CLKBUF_X2 _u40_u1_U72  ( .A(wb1_addr_i[25]), .Z(mast0_pt_in[32]) );
CLKBUF_X2 _u40_u1_U71  ( .A(wb1_addr_i[24]), .Z(mast0_pt_in[31]) );
CLKBUF_X2 _u40_u1_U70  ( .A(wb1_addr_i[23]), .Z(mast0_pt_in[30]) );
CLKBUF_X2 _u40_u1_U69  ( .A(wb1_addr_i[22]), .Z(mast0_pt_in[29]) );
CLKBUF_X2 _u40_u1_U68  ( .A(wb1_addr_i[21]), .Z(mast0_pt_in[28]) );
CLKBUF_X2 _u40_u1_U67  ( .A(wb1_addr_i[20]), .Z(mast0_pt_in[27]) );
CLKBUF_X2 _u40_u1_U66  ( .A(wb1_addr_i[19]), .Z(mast0_pt_in[26]) );
CLKBUF_X2 _u40_u1_U65  ( .A(wb1_addr_i[18]), .Z(mast0_pt_in[25]) );
CLKBUF_X2 _u40_u1_U64  ( .A(wb1_addr_i[17]), .Z(mast0_pt_in[24]) );
CLKBUF_X2 _u40_u1_U63  ( .A(wb1_addr_i[16]), .Z(mast0_pt_in[23]) );
CLKBUF_X2 _u40_u1_U62  ( .A(wb1_addr_i[15]), .Z(mast0_pt_in[22]) );
CLKBUF_X2 _u40_u1_U61  ( .A(wb1_addr_i[14]), .Z(mast0_pt_in[21]) );
CLKBUF_X2 _u40_u1_U60  ( .A(wb1_addr_i[13]), .Z(mast0_pt_in[20]) );
CLKBUF_X2 _u40_u1_U59  ( .A(wb1_addr_i[12]), .Z(mast0_pt_in[19]) );
CLKBUF_X2 _u40_u1_U58  ( .A(wb1_addr_i[11]), .Z(mast0_pt_in[18]) );
CLKBUF_X2 _u40_u1_U57  ( .A(wb1_addr_i[10]), .Z(mast0_pt_in[17]) );
CLKBUF_X2 _u40_u1_U56  ( .A(wb1_addr_i[9]), .Z(mast0_pt_in[16]) );
CLKBUF_X2 _u40_u1_U55  ( .A(wb1_addr_i[8]), .Z(mast0_pt_in[15]) );
CLKBUF_X2 _u40_u1_U54  ( .A(wb1_addr_i[7]), .Z(mast0_pt_in[14]) );
CLKBUF_X2 _u40_u1_U53  ( .A(wb1_addr_i[6]), .Z(mast0_pt_in[13]) );
CLKBUF_X2 _u40_u1_U52  ( .A(wb1_addr_i[5]), .Z(mast0_pt_in[12]) );
CLKBUF_X2 _u40_u1_U51  ( .A(wb1_addr_i[4]), .Z(mast0_pt_in[11]) );
CLKBUF_X2 _u40_u1_U50  ( .A(wb1_addr_i[3]), .Z(mast0_pt_in[10]) );
CLKBUF_X2 _u40_u1_U49  ( .A(wb1_addr_i[2]), .Z(mast0_pt_in[9]) );
CLKBUF_X2 _u40_u1_U48  ( .A(wb1_addr_i[1]), .Z(mast0_pt_in[8]) );
CLKBUF_X2 _u40_u1_U47  ( .A(wb1_addr_i[0]), .Z(mast0_pt_in[7]) );
CLKBUF_X2 _u40_u1_U46  ( .A(wb1_sel_i[3]), .Z(mast0_pt_in[6]) );
CLKBUF_X2 _u40_u1_U45  ( .A(wb1_sel_i[2]), .Z(mast0_pt_in[5]) );
CLKBUF_X2 _u40_u1_U44  ( .A(wb1_sel_i[1]), .Z(mast0_pt_in[4]) );
CLKBUF_X2 _u40_u1_U43  ( .A(wb1_sel_i[0]), .Z(mast0_pt_in[3]) );
CLKBUF_X2 _u40_u1_U42  ( .A(wb1_we_i), .Z(mast0_pt_in[2]) );
CLKBUF_X2 _u40_u1_U41  ( .A(wb1_cyc_i), .Z(mast0_pt_in[1]) );
CLKBUF_X2 _u40_u1_U40  ( .A(wb1_stb_i), .Z(mast0_pt_in[0]) );
CLKBUF_X2 _u40_u1_U39  ( .A(wb1m_data_i[31]), .Z(mast0_pt_in[70]) );
CLKBUF_X2 _u40_u1_U38  ( .A(wb1m_data_i[30]), .Z(mast0_pt_in[69]) );
CLKBUF_X2 _u40_u1_U37  ( .A(wb1m_data_i[29]), .Z(mast0_pt_in[68]) );
CLKBUF_X2 _u40_u1_U36  ( .A(wb1m_data_i[28]), .Z(mast0_pt_in[67]) );
CLKBUF_X2 _u40_u1_U35  ( .A(wb1m_data_i[27]), .Z(mast0_pt_in[66]) );
CLKBUF_X2 _u40_u1_U34  ( .A(wb1m_data_i[26]), .Z(mast0_pt_in[65]) );
CLKBUF_X2 _u40_u1_U33  ( .A(wb1m_data_i[25]), .Z(mast0_pt_in[64]) );
CLKBUF_X2 _u40_u1_U32  ( .A(wb1m_data_i[24]), .Z(mast0_pt_in[63]) );
CLKBUF_X2 _u40_u1_U31  ( .A(wb1m_data_i[23]), .Z(mast0_pt_in[62]) );
CLKBUF_X2 _u40_u1_U30  ( .A(wb1m_data_i[22]), .Z(mast0_pt_in[61]) );
CLKBUF_X2 _u40_u1_U29  ( .A(wb1m_data_i[21]), .Z(mast0_pt_in[60]) );
CLKBUF_X2 _u40_u1_U28  ( .A(wb1m_data_i[20]), .Z(mast0_pt_in[59]) );
CLKBUF_X2 _u40_u1_U27  ( .A(wb1m_data_i[19]), .Z(mast0_pt_in[58]) );
CLKBUF_X2 _u40_u1_U26  ( .A(wb1m_data_i[18]), .Z(mast0_pt_in[57]) );
CLKBUF_X2 _u40_u1_U25  ( .A(wb1m_data_i[17]), .Z(mast0_pt_in[56]) );
CLKBUF_X2 _u40_u1_U24  ( .A(wb1m_data_i[16]), .Z(mast0_pt_in[55]) );
CLKBUF_X2 _u40_u1_U23  ( .A(wb1m_data_i[15]), .Z(mast0_pt_in[54]) );
CLKBUF_X2 _u40_u1_U22  ( .A(wb1m_data_i[14]), .Z(mast0_pt_in[53]) );
CLKBUF_X2 _u40_u1_U21  ( .A(wb1m_data_i[13]), .Z(mast0_pt_in[52]) );
CLKBUF_X2 _u40_u1_U20  ( .A(wb1m_data_i[12]), .Z(mast0_pt_in[51]) );
CLKBUF_X2 _u40_u1_U19  ( .A(wb1m_data_i[11]), .Z(mast0_pt_in[50]) );
CLKBUF_X2 _u40_u1_U18  ( .A(wb1m_data_i[10]), .Z(mast0_pt_in[49]) );
CLKBUF_X2 _u40_u1_U17  ( .A(wb1m_data_i[9]), .Z(mast0_pt_in[48]) );
CLKBUF_X2 _u40_u1_U16  ( .A(wb1m_data_i[8]), .Z(mast0_pt_in[47]) );
CLKBUF_X2 _u40_u1_U15  ( .A(wb1m_data_i[7]), .Z(mast0_pt_in[46]) );
CLKBUF_X2 _u40_u1_U14  ( .A(wb1m_data_i[6]), .Z(mast0_pt_in[45]) );
CLKBUF_X2 _u40_u1_U13  ( .A(wb1m_data_i[5]), .Z(mast0_pt_in[44]) );
CLKBUF_X2 _u40_u1_U12  ( .A(wb1m_data_i[4]), .Z(mast0_pt_in[43]) );
CLKBUF_X2 _u40_u1_U11  ( .A(wb1m_data_i[3]), .Z(mast0_pt_in[42]) );
CLKBUF_X2 _u40_u1_U10  ( .A(wb1m_data_i[2]), .Z(mast0_pt_in[41]) );
CLKBUF_X2 _u40_u1_U9  ( .A(wb1m_data_i[1]), .Z(mast0_pt_in[40]) );
CLKBUF_X2 _u40_u1_U8  ( .A(wb1m_data_i[0]), .Z(mast0_pt_in[39]) );
INV_X1 _u40_u1_U7  ( .A(_u40_u1_n11 ), .ZN(_u40_u1_n16 ) );
INV_X1 _u40_u1_U6  ( .A(_u40_u1_n11 ), .ZN(_u40_u1_n15 ) );
INV_X1 _u40_u1_U5  ( .A(_u40_u1_n11 ), .ZN(_u40_u1_n14 ) );
INV_X8 _u40_u1_U4  ( .A(_u40_u1_n11 ), .ZN(pt0_sel_i) );
NAND2_X2 _u40_u1_U3  ( .A1(wb1_cyc_i), .A2(_u40_u1_n88 ), .ZN(_u40_u1_n11 ));
DFF_X2 _u40_u1_slv_re_reg  ( .D(_u40_u1_N3 ), .CK(clk_i), .Q(_u40_slv_re ),.QN() );
DFF_X2 _u40_u1_slv_we_reg  ( .D(_u40_u1_N4 ), .CK(clk_i), .Q(_u40_slv_we ),.QN() );
DFF_X2 _u40_u1_rf_ack_reg  ( .D(_u40_u1_N5 ), .CK(clk_i), .Q(_u40_u1_rf_ack ), .QN(_u40_u1_n12 ) );
DFF_X2 _u40_u1_slv_dout_reg_0_  ( .D(wb1m_data_i[0]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7950), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_1_  ( .D(wb1m_data_i[1]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7949), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_2_  ( .D(wb1m_data_i[2]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7948), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_3_  ( .D(wb1m_data_i[3]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7947), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_4_  ( .D(wb1m_data_i[4]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7946), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_5_  ( .D(wb1m_data_i[5]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7945), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_6_  ( .D(wb1m_data_i[6]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7944), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_7_  ( .D(wb1m_data_i[7]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7943), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_8_  ( .D(wb1m_data_i[8]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7942), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_9_  ( .D(wb1m_data_i[9]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7941), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_10_  ( .D(wb1m_data_i[10]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7940), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_11_  ( .D(wb1m_data_i[11]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7939), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_12_  ( .D(wb1m_data_i[12]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7938), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_13_  ( .D(wb1m_data_i[13]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7937), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_14_  ( .D(wb1m_data_i[14]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7936), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_15_  ( .D(wb1m_data_i[15]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7935), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_16_  ( .D(wb1m_data_i[16]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7934), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_17_  ( .D(wb1m_data_i[17]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7933), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_18_  ( .D(wb1m_data_i[18]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7932), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_19_  ( .D(wb1m_data_i[19]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7931), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_20_  ( .D(wb1m_data_i[20]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7930), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_21_  ( .D(wb1m_data_i[21]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7929), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_22_  ( .D(wb1m_data_i[22]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7928), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_23_  ( .D(wb1m_data_i[23]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7927), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_24_  ( .D(wb1m_data_i[24]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7926), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_25_  ( .D(wb1m_data_i[25]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7925), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_26_  ( .D(wb1m_data_i[26]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7924), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_27_  ( .D(wb1m_data_i[27]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7923), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_28_  ( .D(wb1m_data_i[28]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7922), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_29_  ( .D(wb1m_data_i[29]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7921), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_30_  ( .D(wb1m_data_i[30]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7920), .QN() );
DFF_X2 _u40_u1_slv_dout_reg_31_  ( .D(wb1m_data_i[31]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7919), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_0_  ( .D(wb1_addr_i[0]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7918), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_1_  ( .D(wb1_addr_i[1]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7917), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_2_  ( .D(wb1_addr_i[2]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7916), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_3_  ( .D(wb1_addr_i[3]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7915), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_4_  ( .D(wb1_addr_i[4]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7914), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_5_  ( .D(wb1_addr_i[5]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7913), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_6_  ( .D(wb1_addr_i[6]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7912), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_7_  ( .D(wb1_addr_i[7]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7911), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_8_  ( .D(wb1_addr_i[8]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7910), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_9_  ( .D(wb1_addr_i[9]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7909), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_10_  ( .D(wb1_addr_i[10]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7908), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_11_  ( .D(wb1_addr_i[11]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7907), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_12_  ( .D(wb1_addr_i[12]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7906), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_13_  ( .D(wb1_addr_i[13]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7905), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_14_  ( .D(wb1_addr_i[14]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7904), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_15_  ( .D(wb1_addr_i[15]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7903), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_16_  ( .D(wb1_addr_i[16]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7902), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_17_  ( .D(wb1_addr_i[17]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7901), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_18_  ( .D(wb1_addr_i[18]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7900), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_19_  ( .D(wb1_addr_i[19]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7899), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_20_  ( .D(wb1_addr_i[20]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7898), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_21_  ( .D(wb1_addr_i[21]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7897), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_22_  ( .D(wb1_addr_i[22]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7896), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_23_  ( .D(wb1_addr_i[23]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7895), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_24_  ( .D(wb1_addr_i[24]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7894), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_25_  ( .D(wb1_addr_i[25]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7893), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_26_  ( .D(wb1_addr_i[26]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7892), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_27_  ( .D(wb1_addr_i[27]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7891), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_28_  ( .D(wb1_addr_i[28]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7890), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_29_  ( .D(wb1_addr_i[29]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7889), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_30_  ( .D(wb1_addr_i[30]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7888), .QN() );
DFF_X2 _u40_u1_slv_adr_reg_31_  ( .D(wb1_addr_i[31]), .CK(clk_i), .Q(SYNOPSYS_UNCONNECTED_7887), .QN() );
endmodule
