module s9234_1(blif_clk_net, blif_reset_net, g89, g94, g98, g102,g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561,g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38,g46, g36, g47, g40, g37, g41, g22, g44, g23, g2584, g3222, g3600,g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282,g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374,g6728, g1290, g4121, g4108, g4106, g4103, g1293, g4099, g4102,g4109, g4100, g4112, g4105, g4101, g4110, g4104, g4107, g4098);
input blif_clk_net, blif_reset_net, g89, g94, g98, g102, g107, g301,g306, g310, g314, g319, g557, g558, g559, g560, g561, g562,g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38,g46, g36, g47, g40, g37, g41, g22, g44, g23;
output g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468,g5469, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368,g6370, g6372, g6374, g6728, g1290, g4121, g4108, g4106, g4103,g1293, g4099, g4102, g4109, g4100, g4112, g4105, g4101, g4110,g4104, g4107, g4098;
wire blif_clk_net, blif_reset_net, g89, g94, g98, g102, g107, g301,g306, g310, g314, g319, g557, g558, g559, g560, g561, g562,g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38,g46, g36, g47, g40, g37, g41, g22, g44, g23;
wire g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468,g5469, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368,g6370, g6372, g6374, g6728, g1290, g4121, g4108, g4106, g4103,g1293, g4099, g4102, g4109, g4100, g4112, g4105, g4101, g4110,g4104, g4107, g4098;
wire g18, g24, g48, g204, g206, g207, g209, g210;
wire g211, g212, g218, g224, g230, g236, g242, g248;
wire g254, g260, g266, g269, g276, g277, g278, g279;
wire g280, g281, g282, g283, g293, g297, g402, g406;
wire g410, g414, g418, g422, g426, g430, g434, g437;
wire g441, g445, g449, g453, g457, g461, g465, g471;
wire g478, g486, g489, g492, g496, g500, g504, g508;
wire g512, g516, g520, g524, g528, g532, g536, g541;
wire g545, g548, g551, g554, g571, g574, g578, g586;
wire g590, g594, g598, g602, g606, g610, g613, g616;
wire g619, g622, g625, g628, g631, g634, g638, g642;
wire g646, g650, g654, g658, g662, g663, g664, g665;
wire g667, g669, g672, g675, g676, g677, g678, g679;
wire g680, g681, g682, g683, g684, g685, g687, g688;
wire g689, g690, g691, g692, g693, g694, g695, g696;
wire g697, g698, g_739, g_895, g_1196, g_1210, g_1775, g_1998;
wire g_2315, g_3105, g_4303, g_4304, g_4325, g_4785, g_4890, g_5464;
wire g_5709, g_6081, n_0, n_1, n_2, n_4, n_5, n_6;
wire n_7, n_8, n_10, n_11, n_13, n_15, n_16, n_18;
wire n_20, n_21, n_26, n_27, n_30, n_31, n_32, n_38;
wire n_39, n_40, n_41, n_46, n_49, n_50, n_57, n_58;
wire n_60, n_62, n_64, n_66, n_67, n_69, n_70, n_73;
wire n_74, n_75, n_76, n_77, n_82, n_86, n_90, n_93;
wire n_94, n_95, n_96, n_98, n_101, n_103, n_104, n_105;
wire n_106, n_107, n_108, n_109, n_115, n_116, n_117, n_119;
wire n_120, n_122, n_126, n_127, n_128, n_129, n_130, n_131;
wire n_133, n_136, n_137, n_139, n_141, n_143, n_144, n_145;
wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
wire n_162, n_163, n_164, n_167, n_168, n_169, n_170, n_172;
wire n_175, n_179, n_180, n_181, n_182, n_183, n_184, n_186;
wire n_187, n_188, n_189, n_190, n_191, n_192, n_194, n_195;
wire n_196, n_197, n_198, n_199, n_200, n_210, n_211, n_213;
wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_224;
wire n_225, n_226, n_227, n_228, n_231, n_232, n_233, n_234;
wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
wire n_243, n_244, n_245, n_246, n_247, n_248, n_250, n_251;
wire n_252, n_253, n_255, n_256, n_266, n_267, n_269, n_270;
wire n_271, n_272, n_273, n_275, n_278, n_279, n_280, n_281;
wire n_282, n_283, n_285, n_286, n_287, n_288, n_291, n_292;
wire n_293, n_295, n_298, n_300, n_301, n_302, n_303, n_304;
wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
wire n_320, n_321, n_322, n_328, n_329, n_330, n_331, n_332;
wire n_334, n_337, n_341, n_342, n_343, n_344, n_345, n_347;
wire n_348, n_351, n_352, n_353, n_354, n_355, n_356, n_358;
wire n_359, n_360, n_364, n_365, n_366, n_367, n_368, n_369;
wire n_370, n_371, n_372, n_374, n_376, n_377, n_378, n_380;
wire n_381, n_383, n_384, n_385, n_388, n_389, n_390, n_391;
wire n_392, n_393, n_397, n_398, n_399, n_404, n_405, n_406;
wire n_407, n_409, n_410, n_411, n_412, n_413, n_415, n_417;
wire n_418, n_420, n_422, n_423, n_424, n_425, n_426, n_427;
wire n_428, n_429, n_430, n_431, n_432, n_433, n_435, n_436;
wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
wire n_455, n_456, n_457, n_460, n_461, n_463, n_464, n_465;
wire n_466, n_467, n_468, n_469, n_472, n_473, n_474, n_475;
wire n_476, n_478, n_479, n_481, n_482, n_485, n_486, n_488;
wire n_489, n_490, n_491, n_494, n_495, n_496, n_497, n_498;
wire n_499, n_501, n_502, n_503, n_504, n_505, n_506, n_507;
wire n_508, n_509, n_510, n_511, n_512, n_513, n_515, n_516;
wire n_517, n_518, n_519, n_521, n_522, n_523, n_525, n_527;
wire n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535;
wire n_536, n_538, n_540, n_541, n_542, n_543, n_544, n_545;
wire n_546, n_547, n_548, n_550, n_551, n_553, n_557, n_559;
wire n_560, n_561, n_562, n_563, n_564, n_567, n_568, n_569;
wire n_571, n_572, n_573, n_575, n_576, n_577, n_578, n_579;
wire n_580, n_581, n_583, n_586, n_587, n_588, n_589, n_590;
wire n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
wire n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606;
wire n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614;
wire n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622;
wire n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630;
wire n_631, n_632, n_635, n_636, n_637, n_638, n_639, n_640;
wire n_642, n_644, n_645, n_646, n_647, n_648, n_649, n_651;
wire n_652, n_654, n_655, n_656, n_657, n_658, n_659, n_660;
wire n_661, n_663, n_665, n_666, n_667, n_668, n_669, n_672;
wire n_673, n_674, n_675, n_677, n_678, n_679, n_680, n_681;
wire n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_692;
wire n_693, n_694, n_696, n_698, n_701, n_703, n_704, n_710;
wire n_711, n_712, n_713, n_714, n_717, n_719, n_720, n_721;
wire n_724, n_725, n_729, n_730, n_731, n_732, n_733, n_734;
wire n_735, n_738, n_740, n_741, n_742, n_746, n_749, n_750;
wire n_752, n_753, n_754, n_755, n_756, n_759, n_760, n_762;
wire n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770;
wire n_771, n_772, n_773, n_774, n_776, n_779, n_784, n_786;
wire n_787, n_788, n_790, n_792, n_793, n_795, n_797, n_798;
wire n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809;
wire n_812, n_815, n_817, n_820, n_821, n_823, n_826, n_827;
wire n_829, n_830, n_831, n_832, n_833, n_836, n_839, n_840;
wire n_842, n_843, n_844, n_846, n_847, n_850, n_851, n_853;
wire n_854, n_855, n_856, n_857, n_858, n_861, n_862, n_863;
wire n_864, n_865, n_867, n_868, n_871, n_872, n_874, n_876;
wire n_877, n_878, n_879, n_881, n_882, n_883, n_884, n_885;
wire n_887, n_888, n_890, n_892, n_895, n_897, n_898, n_899;
wire n_900, n_902, n_903, n_905, n_906, n_907, n_908, n_909;
wire n_910, n_912, n_914, n_916, n_918, n_920, n_922, n_923;
wire n_924, n_926, n_928, n_929, n_930, n_932, n_934, n_939;
wire n_940, n_942, n_943, n_944, n_945, n_946, n_949, n_950;
wire n_951, n_955, n_959, n_960, n_961, n_962, n_985, n_986;
wire n_987, n_988, n_989, n_1003, n_1004, n_1006, n_1007, n_1008;
wire n_1009, n_1012, n_1013, n_1014, n_1018, n_1019, n_1020, n_1030;
wire n_1031, n_1032, n_1036, n_1038, n_1039, n_1041, n_1042, n_1050;
wire n_1051, n_1052, n_1053, n_1054, n_1056, n_1062, n_1064, n_1071;
wire n_1072, n_1073, n_1075, n_1076, n_1081, n_1082, n_1086, n_1087;
wire n_1089, n_1091, n_1092, n_1093, n_1094, n_1095, n_1097, n_1098;
wire n_1099, n_1100, n_1102, n_1104, n_1105, n_1106, n_1109, n_1111;
wire n_1112, n_1113, n_1115, n_1117, n_1118, n_1119, n_1120, n_1121;
wire n_1122, n_1123, n_1124, n_1125, n_1127, n_1128, n_1129, n_1130;
wire n_1132, n_1134, n_1135, n_1137, n_1138, n_1139, n_1140, n_1141;
wire n_1142, n_1143, n_1144, n_1146, n_1147, n_1148, n_1149, n_1150;
wire n_1158, n_1160, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167;
wire n_1168, n_1169, n_1170, n_1171, n_1174, n_1175, n_1176, n_1178;
wire n_1179, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187;
wire n_1188, n_1189, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196;
wire n_1197, n_1198, n_1199, n_1202, n_1203, n_1204, n_1212, n_1215;
wire n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1224;
wire n_1225, n_1226, n_1227, n_1228, n_1230, n_1232, n_1233, n_1235;
wire n_1236, n_1237, n_1238, n_1239, n_1241, n_1242, n_1243, n_1244;
wire n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252;
wire n_1253, n_1254, n_1255, n_1256, n_1257;
assign g4098 = g23;
assign g4107 = g44;
assign g4104 = g22;
assign g4110 = g41;
assign g4101 = g37;
assign g4105 = g40;
assign g4112 = g47;
assign g4100 = g36;
assign g4109 = g46;
assign g4102 = g38;
assign g4099 = g32;
assign g4103 = g39;
assign g4106 = g42;
assign g4108 = g45;
assign g6728 = 1'b0;
assign g5692 = 1'b0;
assign g5469 = g4321;
assign g5468 = g4307;
assign g5137 = g3600;
assign g4422 = g564;
assign g3222 = g705;
DFFSRX1 g48_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_934), .Q (g48), .QN ());
MX2X1 g10574(.A (g6284), .B (n_932), .S0 (n_1164), .Y (n_934));
OR2X1 g10577(.A (n_1164), .B (n_932), .Y (g6284));
XOR2X1 g10580(.A (n_929), .B (n_923), .Y (n_932));
DFFSRX1 g28_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_928), .Q (g_4785), .QN ());
XOR2X1 g10583(.A (n_908), .B (n_924), .Y (n_929));
DFFSRX1 g24_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_926), .Q (g24), .QN ());
MX2X1 g10587(.A (g6366), .B (g_1210), .S0 (n_1164), .Y (n_928));
MX2X1 g10595(.A (g6362), .B (g_3105), .S0 (n_1164), .Y (n_926));
XOR2X1 g10598(.A (g_3105), .B (g_1210), .Y (n_924));
OR2X1 g10599(.A (n_1164), .B (g_1210), .Y (g6366));
DFFSRX1 g10_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_920), .Q (g_739), .QN ());
DFFSRX1 g6_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_922), .Q (g_5709), .QN ());
DFFSRX1 g1_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_918), .Q (g_5464), .QN ());
XOR2X1 g10589(.A (n_910), .B (n_907), .Y (n_923));
DFFSRX1 g2_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_914), .Q (g_1196), .QN ());
DFFSRX1 g14_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_916), .Q (g_6081), .QN ());
DFFSRX1 g18_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_912), .Q (g18), .QN ());
MX2X1 g10596(.A (g6370), .B (g_1775), .S0 (n_1164), .Y (n_922));
MX2X1 g10597(.A (g6372), .B (g_895), .S0 (n_1164), .Y (n_920));
MX2X1 g10603(.A (g6364), .B (n_906), .S0 (n_1164), .Y (n_918));
OR2X1 g10606(.A (n_1164), .B (g_3105), .Y (g6362));
DFFSRX1 g33_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_909), .Q (g_1210), .QN ());
MX2X1 g10600(.A (g6374), .B (g_4304), .S0 (n_1164), .Y (n_916));
MX2X1 g10601(.A (g6368), .B (g_1998), .S0 (n_1164), .Y (n_914));
MX2X1 g10602(.A (g6360), .B (g_4303), .S0 (n_1164), .Y (n_912));
XOR2X1 g10604(.A (g_1775), .B (g_895), .Y (n_910));
DFFSRX1 g29_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_905), .Q (g_3105), .QN ());
OR4X1 g10616(.A (n_862), .B (n_1130), .C (n_1129), .D (n_879), .Y(n_909));
OR2X1 g10607(.A (n_1164), .B (g_1775), .Y (g6370));
OR2X1 g10608(.A (n_1164), .B (g_895), .Y (g6372));
XOR2X1 g10610(.A (g_4304), .B (g_4303), .Y (n_908));
XOR2X1 g10611(.A (g_1998), .B (g_2315), .Y (n_907));
OR2X1 g10619(.A (n_1164), .B (n_906), .Y (g6364));
OR2X1 g10621(.A (n_1164), .B (g_4304), .Y (g6374));
OR4X1 g10627(.A (n_864), .B (n_1132), .C (n_1251), .D (n_1250), .Y(n_905));
OR2X1 g10618(.A (n_1164), .B (g_4303), .Y (g6360));
OR2X1 g10620(.A (n_1164), .B (g_1998), .Y (g6368));
INVX1 g10625(.A (g_2315), .Y (n_906));
NAND3X1 g10634(.A (n_943), .B (n_944), .C (n_892), .Y (n_1129));
DFFSRX1 g11_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_903), .Q (g_1775), .QN ());
DFFSRX1 g15_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_902), .Q (g_895), .QN ());
DFFSRX1 g7_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_899), .Q (g_1998), .QN ());
DFFSRX1 g25_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_900), .Q (g_4303), .QN ());
DFFSRX1 g19_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_897), .Q (g_4304), .QN ());
DFFSRX1 g3_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_898), .Q (), .QN (g_2315));
OR4X1 g10629(.A (n_857), .B (n_559), .C (n_590), .D (n_1147), .Y(n_903));
OR4X1 g10630(.A (n_861), .B (n_823), .C (n_589), .D (n_890), .Y(n_902));
OR4X1 g10633(.A (n_865), .B (n_844), .C (n_573), .D (n_881), .Y(n_900));
OR4X1 g10635(.A (n_661), .B (n_649), .C (n_847), .D (n_883), .Y(n_899));
OR4X1 g10636(.A (n_660), .B (n_668), .C (n_846), .D (n_884), .Y(n_898));
OR4X1 g10637(.A (n_868), .B (n_1255), .C (n_1254), .D (n_878), .Y(n_897));
NAND2X1 g10650(.A (n_830), .B (n_895), .Y (n_943));
DFFSRX1 g211_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_895), .Q (g211), .QN ());
DFFSRX1 g548_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_887), .Q (), .QN (g548));
DFFSRX1 g210_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_1054), .Q (g210), .QN ());
DFFSRX1 g668_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_877), .Q (g4321), .QN ());
NAND2X2 g10673(.A (n_959), .B (n_960), .Y (n_895));
NAND2X1 g10651(.A (n_888), .B (n_872), .Y (n_892));
NAND3X1 g10654(.A (n_645), .B (n_632), .C (n_1256), .Y (n_890));
DFFSRX1 g283_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_888), .Q (g283), .QN ());
DFFSRX1 g545_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_876), .Q (), .QN (g545));
MX2X1 g10674(.A (n_885), .B (n_571), .S0 (n_874), .Y (n_887));
NAND2X2 g10687(.A (n_885), .B (g_4325), .Y (n_959));
NAND2X1 g10662(.A (n_882), .B (n_856), .Y (n_884));
NAND2X1 g10664(.A (n_882), .B (n_843), .Y (n_883));
DFFSRX1 g554_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_867), .Q (), .QN (g554));
NAND2X1 g10667(.A (n_644), .B (n_1256), .Y (n_881));
NAND2X1 g10668(.A (n_656), .B (n_1257), .Y (n_1251));
NAND2X1 g10669(.A (n_663), .B (n_1257), .Y (n_879));
NAND2X1 g10670(.A (n_665), .B (n_1257), .Y (n_878));
NAND2X1 g10683(.A (n_885), .B (n_1056), .Y (n_877));
MX2X1 g10698(.A (n_1056), .B (n_561), .S0 (n_874), .Y (n_876));
DFFSRX1 g485_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_858), .Q (g4307), .QN ());
DFFSRX1 g282_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_871), .Q (g282), .QN ());
NAND2X2 g10672(.A (n_1233), .B (n_949), .Y (n_888));
NAND2X2 g10703(.A (n_850), .B (n_851), .Y (n_885));
OAI21X1 g10663(.A0 (n_805), .A1 (n_226), .B0 (n_855), .Y (n_868));
DFFSRX1 g551_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_853), .Q (), .QN (g551));
MX2X1 g10675(.A (n_1232), .B (n_563), .S0 (n_874), .Y (n_867));
NAND3X1 g10685(.A (n_1150), .B (n_692), .C (n_498), .Y (n_882));
OAI21X1 g10689(.A0 (n_863), .A1 (n_581), .B0 (n_542), .Y (n_865));
OAI21X1 g10690(.A0 (n_863), .A1 (n_141), .B0 (n_545), .Y (n_864));
OAI21X1 g10691(.A0 (n_863), .A1 (n_271), .B0 (n_544), .Y (n_862));
NAND2X2 g10695(.A (n_1241), .B (n_955), .Y (n_871));
NAND3X1 g10678(.A (n_821), .B (n_842), .C (n_531), .Y (n_861));
NAND2X1 g10686(.A (n_1232), .B (n_1239), .Y (n_858));
NAND3X1 g10688(.A (n_945), .B (n_833), .C (n_946), .Y (n_857));
AOI21X1 g10692(.A0 (n_854), .A1 (n_767), .B0 (n_809), .Y (n_856));
AOI22X1 g10693(.A0 (n_854), .A1 (n_312), .B0 (n_628), .B1 (g560), .Y(n_855));
MX2X1 g10697(.A (n_1239), .B (n_567), .S0 (n_874), .Y (n_853));
INVX1 g10737(.A (n_1227), .Y (n_850));
NAND2X1 g10729(.A (n_831), .B (n_629), .Y (n_847));
NAND2X1 g10733(.A (n_829), .B (n_631), .Y (n_846));
DFFSRX1 g536_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_836), .Q (), .QN (g536));
NAND3X1 g10679(.A (n_950), .B (n_802), .C (n_951), .Y (n_844));
AOI21X1 g10707(.A0 (n_826), .A1 (n_765), .B0 (n_820), .Y (n_843));
INVX2 g10723(.A (n_854), .Y (n_863));
NAND2X1 g10732(.A (n_840), .B (n_1092), .Y (n_842));
NAND2X1 g10735(.A (n_840), .B (n_832), .Y (n_946));
AOI21X1 g10750(.A0 (n_657), .A1 (n_1220), .B0 (n_1228), .Y (n_839));
OAI21X1 g10704(.A0 (n_760), .A1 (n_368), .B0 (n_815), .Y (n_836));
INVX2 g10724(.A (n_827), .Y (n_854));
NAND2X1 g10736(.A (n_812), .B (n_832), .Y (n_833));
AOI21X1 g10759(.A0 (n_830), .A1 (n_683), .B0 (n_806), .Y (n_831));
AOI21X1 g10761(.A0 (n_830), .A1 (n_693), .B0 (n_779), .Y (n_829));
AOI21X1 g10765(.A0 (n_872), .A1 (n_666), .B0 (n_808), .Y (n_945));
DFFSRX1 g541_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_1094), .Q (), .QN (g541));
DFFSRX1 g496_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_817), .Q (), .QN (g496));
NOR2X1 g10725(.A (n_754), .B (n_826), .Y (n_827));
NAND2X1 g10727(.A (n_684), .B (n_1008), .Y (n_950));
DFFSRX1 g594_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_803), .Q (), .QN (g594));
OAI22X1 g10739(.A0 (n_1007), .A1 (n_679), .B0 (n_1248), .B1 (n_1091),.Y (n_823));
DFFSRX1 g532_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_788), .Q (g532), .QN ());
INVX1 g10753(.A (n_1138), .Y (n_840));
AOI21X1 g10760(.A0 (n_872), .A1 (n_659), .B0 (n_784), .Y (n_821));
NAND2X1 g10763(.A (n_755), .B (n_787), .Y (n_820));
OAI22X1 g10764(.A0 (n_730), .A1 (n_680), .B0 (n_1007), .B1 (n_703),.Y (n_1254));
DFFSRX1 g582_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_786), .Q (n_432), .QN ());
DFFSRX1 g578_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_798), .Q (g578), .QN ());
DFFSRX1 g586_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_804), .Q (), .QN (g586));
DFFSRX1 g465_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_797), .Q (), .QN (g465));
DFFSRX1 g520_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_795), .Q (g520), .QN ());
DFFSRX1 g524_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_793), .Q (g524), .QN ());
DFFSRX1 g528_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_790), .Q (g528), .QN ());
DFFSRX1 g492_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_807), .Q (), .QN (g492));
NAND3X1 g10827(.A (n_1222), .B (n_746), .C (g496), .Y (n_817));
AOI22X1 g10740(.A0 (n_759), .A1 (n_874), .B0 (n_1086), .B1 (n_832),.Y (n_815));
INVX1 g10751(.A (n_1071), .Y (n_812));
DFFSRX1 g574_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_770), .Q (), .QN (g574));
DFFSRX1 g590_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_756), .Q (), .QN (g590));
DFFSRX1 g500_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_768), .Q (g500), .QN ());
DFFSRX1 g504_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_766), .Q (g504), .QN ());
DFFSRX1 g512_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_763), .Q (g512), .QN ());
DFFSRX1 g508_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_764), .Q (g508), .QN ());
NOR2X1 g10783(.A (n_655), .B (n_752), .Y (n_809));
NOR2X1 g10795(.A (n_776), .B (n_651), .Y (n_808));
DFFSRX1 g516_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_762), .Q (g516), .QN ());
NAND2X1 g10826(.A (n_749), .B (n_1109), .Y (n_807));
NOR2X1 g10829(.A (n_805), .B (n_214), .Y (n_806));
INVX1 g10563(.A (n_774), .Y (n_804));
INVX1 g10565(.A (n_771), .Y (n_803));
NAND2X1 g10726(.A (n_658), .B (n_872), .Y (n_802));
NAND2X1 g10756(.A (n_1073), .B (n_1248), .Y (n_826));
INVX1 g10568(.A (n_769), .Y (n_798));
MX2X1 g10767(.A (n_383), .B (n_765), .S0 (n_1087), .Y (n_797));
OAI21X1 g10773(.A0 (n_792), .A1 (n_581), .B0 (n_742), .Y (n_795));
OAI21X1 g10774(.A0 (n_792), .A1 (n_141), .B0 (n_741), .Y (n_793));
OAI21X1 g10775(.A0 (n_792), .A1 (n_271), .B0 (n_740), .Y (n_790));
MX2X1 g10776(.A (g532), .B (n_767), .S0 (n_1087), .Y (n_788));
NAND2X1 g10788(.A (n_872), .B (n_682), .Y (n_787));
INVX1 g10561(.A (n_773), .Y (n_786));
OR2X1 g10806(.A (n_805), .B (n_581), .Y (n_951));
NOR2X1 g10809(.A (n_805), .B (n_1091), .Y (n_784));
OR2X1 g10811(.A (n_805), .B (n_271), .Y (n_944));
NOR2X1 g10812(.A (n_805), .B (n_172), .Y (n_779));
INVX2 g10817(.A (n_1007), .Y (n_830));
INVX1 g10821(.A (n_1006), .Y (n_776));
NAND2X1 g10564(.A (n_642), .B (n_772), .Y (n_774));
NAND2X1 g10562(.A (n_588), .B (n_772), .Y (n_773));
NAND2X1 g10566(.A (n_720), .B (n_772), .Y (n_771));
NAND2X1 g10567(.A (n_686), .B (n_772), .Y (n_770));
NAND2X1 g10569(.A (n_512), .B (n_772), .Y (n_769));
MX2X1 g10768(.A (n_767), .B (g500), .S0 (n_792), .Y (n_768));
MX2X1 g10769(.A (n_765), .B (g504), .S0 (n_792), .Y (n_766));
MX2X1 g10770(.A (n_832), .B (g508), .S0 (n_792), .Y (n_764));
MX2X1 g10771(.A (n_1092), .B (g512), .S0 (n_792), .Y (n_763));
MX2X1 g10772(.A (n_312), .B (g516), .S0 (n_792), .Y (n_762));
DFFSRX1 g269_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_735), .Q (g269), .QN ());
DFFSRX1 g297_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_732), .Q (), .QN (g297));
DFFSRX1 g197_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_731), .Q (g_4325), .QN ());
DFFSRX1 g293_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_734), .Q (), .QN (g293));
INVX1 g10792(.A (n_759), .Y (n_760));
NAND2X1 g10560(.A (n_714), .B (n_772), .Y (n_756));
NAND2X1 g10807(.A (n_754), .B (n_765), .Y (n_755));
NOR2X1 g10808(.A (n_550), .B (n_1111), .Y (n_753));
INVX1 g10813(.A (n_872), .Y (n_752));
INVX2 g10844(.A (n_750), .Y (n_805));
NOR2X1 g10852(.A (n_725), .B (n_507), .Y (n_749));
INVX1 g10862(.A (n_1199), .Y (n_746));
NAND2X1 g10789(.A (n_792), .B (g520), .Y (n_742));
NAND2X1 g10790(.A (n_792), .B (g524), .Y (n_741));
NAND2X1 g10791(.A (n_792), .B (g528), .Y (n_740));
NOR2X1 g10793(.A (n_1086), .B (g536), .Y (n_759));
INVX2 g10815(.A (n_730), .Y (n_872));
INVX1 g10845(.A (n_738), .Y (n_750));
INVX1 g10850(.A (n_1072), .Y (n_754));
INVX1 g10570(.A (n_721), .Y (n_772));
MX2X1 g10800(.A (n_1230), .B (n_765), .S0 (n_733), .Y (n_735));
MX2X1 g10801(.A (n_516), .B (n_832), .S0 (n_733), .Y (n_734));
MX2X1 g10802(.A (n_518), .B (n_1092), .S0 (n_733), .Y (n_732));
MX2X1 g10803(.A (n_675), .B (n_767), .S0 (n_733), .Y (n_731));
NAND2X1 g10816(.A (n_989), .B (n_311), .Y (n_730));
NAND2X2 g10828(.A (n_729), .B (g677), .Y (n_792));
INVX1 g10841(.A (n_989), .Y (n_939));
NAND2X1 g10846(.A (n_322), .B (n_712), .Y (n_738));
INVX1 g10869(.A (n_724), .Y (n_725));
OAI21X1 g10571(.A0 (n_719), .A1 (g594), .B0 (g639), .Y (n_721));
XOR2X1 g10572(.A (g594), .B (n_719), .Y (n_720));
INVX1 g10848(.A (n_1243), .Y (n_717));
NAND2X1 g10870(.A (n_1106), .B (n_696), .Y (n_724));
XOR2X1 g10575(.A (n_150), .B (n_688), .Y (n_714));
NAND3X1 g10933(.A (n_694), .B (n_425), .C (n_359), .Y (n_851));
DFFSRX1 g208_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_704), .Q (n_371), .QN ());
DFFSRX1 g669_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_701), .Q (), .QN (g669));
NOR2X1 g10837(.A (n_448), .B (n_713), .Y (n_733));
NOR2X1 g10838(.A (n_407), .B (n_713), .Y (n_729));
INVX1 g10872(.A (n_711), .Y (n_712));
INVX1 g10873(.A (n_711), .Y (n_710));
OR2X1 g10865(.A (n_1160), .B (n_248), .Y (g6282));
INVX1 g10831(.A (n_703), .Y (n_704));
INVX2 g10874(.A (n_1249), .Y (n_711));
OR2X1 g10904(.A (n_677), .B (n_630), .Y (n_701));
NAND2X1 g10576(.A (n_687), .B (n_150), .Y (n_719));
NAND2X1 g10926(.A (n_1171), .B (n_696), .Y (n_698));
DFFSRX1 g280_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_681), .Q (g280), .QN ());
INVX1 g10994(.A (n_1195), .Y (n_694));
DFFSRX1 g204_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_693), .Q (g204), .QN ());
DFFSRX1 g672_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_672), .Q (), .QN (g672));
AOI21X1 g10832(.A0 (n_640), .A1 (n_66), .B0 (n_270), .Y (n_703));
OR2X1 g10866(.A (n_285), .B (n_1160), .Y (n_713));
AND2X1 g10871(.A (n_637), .B (n_648), .Y (n_692));
INVX1 g10578(.A (n_687), .Y (n_688));
XOR2X1 g10579(.A (n_168), .B (n_674), .Y (n_686));
INVX1 g10984(.A (n_1171), .Y (n_685));
DFFSRX1 g209_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_684), .Q (g209), .QN ());
DFFSRX1 g207_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_678), .Q (g207), .QN ());
DFFSRX1 g205_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_683), .Q (g_4890), .QN ());
DFFSRX1 g206_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_652), .Q (g206), .QN ());
DFFSRX1 g277_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_682), .Q (g277), .QN ());
DFFSRX1 g430_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_611), .Q (), .QN (g430));
INVX1 g10833(.A (n_680), .Y (n_681));
DFFSRX1 g445_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_604), .Q (), .QN (g445));
INVX1 g10914(.A (n_678), .Y (n_679));
DFFSRX1 g422_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_615), .Q (), .QN (g422));
NOR2X1 g10928(.A (n_667), .B (g22), .Y (n_677));
DFFSRX1 g457_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_598), .Q (), .QN (g457));
OAI21X1 g10940(.A0 (n_172), .A1 (n_675), .B0 (n_592), .Y (n_693));
DFFSRX1 g449_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_602), .Q (), .QN (g449));
NOR2X1 g10581(.A (n_674), .B (g574), .Y (n_687));
NAND2X1 g10975(.A (n_498), .B (n_587), .Y (n_673));
OR2X1 g10980(.A (n_593), .B (n_626), .Y (n_672));
INVX1 g11012(.A (n_646), .Y (n_668));
DFFSRX1 g406_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_624), .Q (), .QN (g406));
DFFSRX1 g276_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_654), .Q (g276), .QN ());
DFFSRX1 g402_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_625), .Q (), .QN (g402));
DFFSRX1 g410_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_621), .Q (), .QN (g410));
DFFSRX1 g414_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_619), .Q (), .QN (g414));
DFFSRX1 g418_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_617), .Q (), .QN (g418));
DFFSRX1 g426_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_613), .Q (), .QN (g426));
DFFSRX1 g434_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_609), .Q (), .QN (g434));
DFFSRX1 g441_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_606), .Q (), .QN (g441));
DFFSRX1 g437_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_608), .Q (), .QN (g437));
DFFSRX1 g453_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_600), .Q (), .QN (g453));
DFFSRX1 g461_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_596), .Q (), .QN (g461));
DFFSRX1 g676_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_667), .Q (g676), .QN ());
DFFSRX1 g278_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_666), .Q (g278), .QN ());
OR2X1 g11023(.A (n_13), .B (n_481), .Y (n_665));
AOI21X1 g10834(.A0 (n_551), .A1 (n_1230), .B0 (n_269), .Y (n_680));
OR2X1 g11026(.A (n_20), .B (n_481), .Y (n_663));
NAND4X1 g10905(.A (n_572), .B (n_508), .C (n_503), .D (n_504), .Y(n_661));
NAND4X1 g10907(.A (n_562), .B (n_506), .C (n_501), .D (n_502), .Y(n_660));
DFFSRX1 g279_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_659), .Q (g279), .QN ());
OAI22X1 g10915(.A0 (n_538), .A1 (n_499), .B0 (n_1091), .B1 (n_66), .Y(n_678));
DFFSRX1 g281_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_658), .Q (g281), .QN ());
AND2X1 g10930(.A (n_578), .B (g210), .Y (n_657));
OR2X1 g11025(.A (n_1), .B (n_481), .Y (n_656));
INVX1 g10937(.A (n_654), .Y (n_655));
OAI21X1 g10939(.A0 (n_214), .A1 (g269), .B0 (n_580), .Y (n_682));
OAI21X1 g10941(.A0 (n_675), .A1 (n_256), .B0 (n_576), .Y (n_683));
INVX1 g10943(.A (n_651), .Y (n_652));
OAI21X1 g10758(.A0 (n_581), .A1 (g_4325), .B0 (n_553), .Y (n_684));
INVX1 g11018(.A (n_639), .Y (n_649));
NOR2X1 g10989(.A (n_647), .B (n_586), .Y (n_648));
AOI22X1 g11013(.A0 (g500), .A1 (n_557), .B0 (g532), .B1 (n_638), .Y(n_646));
DFFSRX1 g571_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_583), .Q (), .QN (g571));
OR2X1 g11027(.A (n_7), .B (n_481), .Y (n_645));
OR2X1 g11029(.A (n_8), .B (n_481), .Y (n_644));
XOR2X1 g10588(.A (n_27), .B (n_1039), .Y (n_642));
NAND2X1 g10594(.A (n_1039), .B (n_27), .Y (n_674));
NAND2X1 g10878(.A (n_412), .B (n_591), .Y (n_640));
AOI22X1 g11019(.A0 (n_638), .A1 (n_383), .B0 (n_557), .B1 (g504), .Y(n_639));
NOR2X1 g10906(.A (n_636), .B (n_635), .Y (n_637));
OAI21X1 g10938(.A0 (n_347), .A1 (n_1230), .B0 (n_541), .Y (n_654));
OAI21X1 g10942(.A0 (n_579), .A1 (n_365), .B0 (n_275), .Y (n_666));
AOI21X1 g10944(.A0 (n_575), .A1 (n_295), .B0 (n_225), .Y (n_651));
AND2X1 g10946(.A (n_543), .B (n_519), .Y (n_632));
AOI22X1 g10948(.A0 (n_628), .A1 (g564), .B0 (n_627), .B1 (n_630), .Y(n_631));
AOI22X1 g10949(.A0 (n_628), .A1 (g563), .B0 (n_627), .B1 (n_626), .Y(n_629));
MX2X1 g10951(.A (n_623), .B (n_384), .S0 (n_622), .Y (n_625));
MX2X1 g10952(.A (n_620), .B (n_623), .S0 (n_622), .Y (n_624));
MX2X1 g10953(.A (n_618), .B (n_620), .S0 (n_622), .Y (n_621));
MX2X1 g10954(.A (n_616), .B (n_618), .S0 (n_622), .Y (n_619));
MX2X1 g10955(.A (n_614), .B (n_616), .S0 (n_622), .Y (n_617));
MX2X1 g10956(.A (n_612), .B (n_614), .S0 (n_622), .Y (n_615));
MX2X1 g10957(.A (n_610), .B (n_612), .S0 (n_622), .Y (n_613));
MX2X1 g10958(.A (n_594), .B (n_610), .S0 (n_622), .Y (n_611));
MX2X1 g10959(.A (n_528), .B (n_607), .S0 (n_622), .Y (n_609));
MX2X1 g10960(.A (n_607), .B (n_605), .S0 (n_622), .Y (n_608));
MX2X1 g10961(.A (n_605), .B (n_603), .S0 (n_622), .Y (n_606));
XOR2X1 g11020(.A (g48), .B (n_494), .Y (n_667));
MX2X1 g10962(.A (n_603), .B (n_601), .S0 (n_622), .Y (n_604));
MX2X1 g10963(.A (n_601), .B (n_599), .S0 (n_622), .Y (n_602));
MX2X1 g10964(.A (n_599), .B (n_597), .S0 (n_622), .Y (n_600));
MX2X1 g10965(.A (n_597), .B (n_595), .S0 (n_622), .Y (n_598));
MX2X1 g10966(.A (n_595), .B (n_594), .S0 (n_622), .Y (n_596));
NOR2X1 g11024(.A (n_119), .B (n_521), .Y (n_593));
NAND3X1 g10990(.A (n_591), .B (n_217), .C (g_4325), .Y (n_592));
INVX1 g11004(.A (n_569), .Y (n_590));
INVX1 g11010(.A (n_564), .Y (n_589));
DFFSRX1 g631_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_547), .Q (g631), .QN ());
DFFSRX1 g43_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_523), .Q (g3600), .QN ());
XOR2X1 g10609(.A (n_432), .B (n_515), .Y (n_588));
INVX1 g11041(.A (n_586), .Y (n_587));
NAND2X2 g11055(.A (n_522), .B (n_497), .Y (n_669));
NAND2X1 g10628(.A (n_511), .B (n_513), .Y (n_583));
OAI22X1 g10913(.A0 (n_491), .A1 (n_466), .B0 (n_1091), .B1 (n_1230),.Y (n_659));
OAI21X1 g10757(.A0 (n_581), .A1 (g269), .B0 (n_496), .Y (n_658));
OR2X1 g10979(.A (n_579), .B (n_190), .Y (n_580));
INVX1 g10981(.A (n_577), .Y (n_578));
NAND3X1 g10991(.A (n_575), .B (n_143), .C (n_1097), .Y (n_576));
INVX1 g10997(.A (n_535), .Y (n_1255));
INVX1 g10999(.A (n_534), .Y (n_573));
AOI22X1 g11001(.A0 (n_568), .A1 (n_571), .B0 (n_560), .B1 (n_1230),.Y (n_572));
AOI22X1 g11005(.A0 (n_568), .A1 (n_567), .B0 (n_465), .B1 (n_638), .Y(n_569));
INVX1 g11006(.A (n_530), .Y (n_1132));
INVX1 g11008(.A (n_529), .Y (n_1130));
AOI22X1 g11011(.A0 (n_568), .A1 (n_563), .B0 (n_536), .B1 (n_638), .Y(n_564));
AOI22X1 g11014(.A0 (n_568), .A1 (n_561), .B0 (n_560), .B1 (n_675), .Y(n_562));
INVX1 g11016(.A (n_527), .Y (n_559));
DFFSRX1 g654_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_509), .Q (), .QN (g654));
OR2X1 g11042(.A (n_638), .B (n_557), .Y (n_586));
NAND3X1 g10799(.A (n_457), .B (n_525), .C (n_66), .Y (n_553));
NAND2X1 g10879(.A (n_430), .B (n_540), .Y (n_551));
NAND2X1 g10925(.A (n_548), .B (g282), .Y (n_550));
NAND3X1 g10931(.A (n_452), .B (n_475), .C (n_485), .Y (n_636));
AND2X1 g10641(.A (n_489), .B (g639), .Y (n_547));
NAND2X1 g10968(.A (n_628), .B (g562), .Y (n_546));
NAND2X1 g10969(.A (n_628), .B (g558), .Y (n_545));
NAND2X1 g10970(.A (n_628), .B (g557), .Y (n_544));
NAND2X1 g10971(.A (n_628), .B (g561), .Y (n_543));
NAND2X1 g10972(.A (n_628), .B (g559), .Y (n_542));
NAND3X1 g10978(.A (n_540), .B (n_232), .C (n_1230), .Y (n_541));
NAND2X1 g10982(.A (n_488), .B (n_468), .Y (n_577));
AND2X1 g10988(.A (n_343), .B (n_525), .Y (n_538));
AOI22X1 g10998(.A0 (n_614), .A1 (n_533), .B0 (n_603), .B1 (n_532), .Y(n_535));
AOI22X1 g11000(.A0 (n_612), .A1 (n_533), .B0 (n_605), .B1 (n_532), .Y(n_534));
AOI22X1 g11003(.A0 (n_616), .A1 (n_533), .B0 (n_601), .B1 (n_532), .Y(n_531));
AOI22X1 g11007(.A0 (n_610), .A1 (n_533), .B0 (n_607), .B1 (n_532), .Y(n_530));
AOI22X1 g11009(.A0 (n_528), .A1 (n_532), .B0 (n_594), .B1 (n_533), .Y(n_529));
AOI22X1 g11017(.A0 (n_618), .A1 (n_533), .B0 (n_599), .B1 (n_532), .Y(n_527));
AND2X1 g11038(.A (n_1062), .B (n_525), .Y (n_591));
AOI21X1 g11051(.A0 (n_151), .A1 (n_460), .B0 (n_292), .Y (n_523));
NAND2X1 g11079(.A (n_478), .B (n_255), .Y (n_522));
INVX1 g11091(.A (n_1135), .Y (n_521));
NAND2X1 g11106(.A (n_560), .B (n_518), .Y (n_519));
NAND2X1 g11110(.A (n_560), .B (n_516), .Y (n_517));
INVX1 g10631(.A (n_1042), .Y (n_515));
DFFSRX1 g628_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_463), .Q (g628), .QN ());
NAND4X1 g10638(.A (n_510), .B (n_473), .C (g638), .D (n_31), .Y(n_513));
XOR2X1 g10639(.A (g578), .B (n_1041), .Y (n_512));
NAND3X1 g10644(.A (n_510), .B (n_39), .C (g638), .Y (n_511));
AND2X1 g10649(.A (n_474), .B (g638), .Y (n_509));
DFFSRX1 g650_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_472), .Q (g650), .QN ());
AOI22X1 g11002(.A0 (n_635), .A1 (g489), .B0 (n_647), .B1 (n_507), .Y(n_508));
AOI22X1 g11015(.A0 (n_635), .A1 (g486), .B0 (n_647), .B1 (n_40), .Y(n_506));
AND2X1 g11028(.A (g541), .B (n_505), .Y (n_622));
NAND2X1 g11030(.A (n_467), .B (n_495), .Y (n_579));
NAND2X1 g11031(.A (n_533), .B (n_620), .Y (n_504));
NAND2X1 g11032(.A (n_532), .B (n_597), .Y (n_503));
NAND2X1 g11035(.A (n_595), .B (n_532), .Y (n_502));
NAND2X1 g11036(.A (n_623), .B (n_533), .Y (n_501));
NOR2X1 g11044(.A (n_499), .B (n_482), .Y (n_575));
INVX1 g11049(.A (n_498), .Y (n_627));
INVX1 g11070(.A (n_481), .Y (n_557));
NAND3X1 g11078(.A (g471), .B (n_1219), .C (n_476), .Y (n_497));
NAND3X1 g10798(.A (n_461), .B (n_495), .C (g269), .Y (n_496));
XOR2X1 g11090(.A (n_334), .B (n_1188), .Y (n_494));
AOI21X1 g10983(.A0 (n_355), .A1 (n_469), .B0 (n_455), .Y (n_548));
AND2X1 g10987(.A (n_369), .B (n_495), .Y (n_491));
DFFSRX1 g625_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_456), .Q (g625), .QN ());
AND2X1 g11037(.A (n_490), .B (n_495), .Y (n_540));
XOR2X1 g10671(.A (g631), .B (n_446), .Y (n_489));
NAND2X1 g11040(.A (n_360), .B (n_486), .Y (n_488));
INVX1 g11045(.A (n_485), .Y (n_628));
NAND2X1 g11050(.A (n_454), .B (n_183), .Y (n_498));
INVX1 g11060(.A (n_482), .Y (n_525));
NAND2X2 g11071(.A (n_451), .B (g677), .Y (n_481));
NAND2X1 g11119(.A (n_1179), .B (n_1194), .Y (n_479));
NAND2X1 g11120(.A (n_1219), .B (n_476), .Y (n_478));
INVX1 g11129(.A (n_475), .Y (n_560));
XOR2X1 g10694(.A (n_31), .B (n_473), .Y (n_474));
DFFSRX1 g646_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_442), .Q (g646), .QN ());
AND2X1 g10700(.A (n_443), .B (g638), .Y (n_472));
AOI22X1 g11199(.A0 (g486), .A1 (n_40), .B0 (g489), .B1 (n_507), .Y(g4809));
NAND3X1 g10652(.A (n_39), .B (n_473), .C (n_31), .Y (n_510));
NAND4X1 g11047(.A (n_440), .B (g680), .C (g678), .D (g679), .Y(n_485));
NAND2X1 g11061(.A (n_1196), .B (n_468), .Y (n_482));
INVX1 g11064(.A (n_466), .Y (n_467));
NOR2X1 g11073(.A (n_450), .B (g677), .Y (n_638));
NOR2X1 g11074(.A (n_874), .B (n_465), .Y (n_505));
NOR2X1 g11075(.A (n_464), .B (g677), .Y (n_532));
NOR2X1 g11076(.A (n_464), .B (n_175), .Y (n_533));
AND2X1 g10680(.A (n_444), .B (g639), .Y (n_463));
NAND2X1 g10805(.A (n_447), .B (n_490), .Y (n_461));
MX2X1 g11118(.A (n_433), .B (n_405), .S0 (n_27), .Y (n_460));
NAND2X1 g11130(.A (n_449), .B (n_441), .Y (n_475));
NAND2X1 g10825(.A (n_431), .B (n_1062), .Y (n_457));
AND2X1 g10748(.A (n_435), .B (g639), .Y (n_456));
NOR2X1 g11058(.A (n_696), .B (n_455), .Y (n_495));
NAND2X1 g11063(.A (n_1062), .B (g_4325), .Y (n_499));
NAND2X1 g11065(.A (n_490), .B (g269), .Y (n_466));
NOR2X1 g11077(.A (n_453), .B (g680), .Y (n_454));
NOR2X1 g11081(.A (n_281), .B (n_453), .Y (n_647));
NOR2X1 g11083(.A (n_282), .B (n_453), .Y (n_635));
INVX1 g11084(.A (n_452), .Y (n_568));
NAND2X1 g11089(.A (n_422), .B (n_409), .Y (n_486));
INVX1 g11099(.A (n_450), .Y (n_451));
DFFSRX1 g606_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_413), .Q (g606), .QN ());
NAND3X1 g11137(.A (n_940), .B (n_381), .C (g206), .Y (n_476));
INVX1 g11165(.A (n_448), .Y (n_449));
XOR2X1 g10857(.A (g281), .B (n_429), .Y (n_447));
INVX1 g10708(.A (n_445), .Y (n_446));
DFFSRX1 g622_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_417), .Q (g622), .QN ());
XOR2X1 g10741(.A (g628), .B (n_428), .Y (n_444));
XOR2X1 g10766(.A (g650), .B (n_427), .Y (n_443));
AND2X1 g10782(.A (n_415), .B (g638), .Y (n_442));
NAND4X1 g11085(.A (n_439), .B (n_392), .C (n_139), .D (g682), .Y(n_452));
NAND2X1 g11088(.A (n_391), .B (n_410), .Y (n_469));
NAND2X1 g11100(.A (n_436), .B (n_441), .Y (n_450));
NAND2X1 g11103(.A (n_424), .B (n_389), .Y (n_468));
NAND3X1 g11113(.A (n_420), .B (n_242), .C (n_245), .Y (n_874));
INVX1 g11115(.A (n_453), .Y (n_440));
NAND2X1 g11117(.A (n_418), .B (n_439), .Y (n_464));
XOR2X1 g10830(.A (g625), .B (n_378), .Y (n_435));
NAND3X1 g11166(.A (n_392), .B (g683), .C (g684), .Y (n_448));
AOI22X1 g11169(.A0 (n_376), .A1 (n_432), .B0 (n_352), .B1 (n_404), .Y(n_433));
XOR2X1 g10858(.A (g209), .B (n_411), .Y (n_431));
DFFSRX1 g489_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_214), .Q (), .QN (g489));
OAI21X1 g10936(.A0 (n_342), .A1 (g280), .B0 (n_429), .Y (n_430));
NAND2X1 g10749(.A (n_428), .B (g628), .Y (n_445));
DFFSRX1 g619_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_397), .Q (g619), .QN ());
AND2X1 g10781(.A (n_427), .B (g650), .Y (n_473));
MX2X1 g11086(.A (n_425), .B (n_696), .S0 (n_383), .Y (n_426));
NOR2X1 g11105(.A (n_286), .B (n_423), .Y (n_455));
NAND2X1 g11108(.A (n_287), .B (n_423), .Y (n_490));
NAND2X1 g11114(.A (n_337), .B (n_255), .Y (n_422));
NAND3X1 g11116(.A (n_283), .B (n_441), .C (g688), .Y (n_453));
AND2X1 g11135(.A (n_441), .B (n_406), .Y (n_439));
NOR2X1 g11138(.A (n_364), .B (n_385), .Y (n_420));
INVX1 g11146(.A (n_407), .Y (n_436));
NOR2X1 g11159(.A (n_393), .B (g682), .Y (n_418));
AND2X1 g10836(.A (n_374), .B (g639), .Y (n_417));
XOR2X1 g10856(.A (g646), .B (n_398), .Y (n_415));
AND2X1 g10868(.A (n_372), .B (g638), .Y (n_413));
OAI21X1 g10935(.A0 (n_301), .A1 (n_371), .B0 (n_411), .Y (n_412));
DFFSRX1 g642_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_370), .Q (g642), .QN ());
NAND2X1 g11102(.A (n_388), .B (g478), .Y (n_410));
NAND2X1 g11112(.A (n_389), .B (g471), .Y (n_409));
NAND4X1 g11147(.A (n_380), .B (n_406), .C (g681), .D (g682), .Y(n_407));
NOR2X1 g10839(.A (n_377), .B (n_2), .Y (n_428));
AOI22X1 g11170(.A0 (n_316), .A1 (n_432), .B0 (n_317), .B1 (n_404), .Y(n_405));
NAND2X1 g11185(.A (n_353), .B (g_4890), .Y (n_940));
INVX1 g11203(.A (n_399), .Y (n_1253));
AND2X1 g10867(.A (n_398), .B (g646), .Y (n_427));
DFFSRX1 g486_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_347), .Q (), .QN (g486));
AND2X1 g10922(.A (n_344), .B (g639), .Y (n_397));
NAND2X1 g10974(.A (n_342), .B (g280), .Y (n_429));
INVX1 g11195(.A (n_393), .Y (n_392));
NAND2X1 g11104(.A (n_367), .B (n_390), .Y (n_391));
INVX1 g11131(.A (n_388), .Y (n_423));
INVX1 g11141(.A (n_1196), .Y (n_425));
NAND2X1 g11157(.A (n_1036), .B (n_330), .Y (n_441));
NAND4X1 g11171(.A (n_278), .B (n_243), .C (n_246), .D (n_194), .Y(n_385));
MX2X1 g11172(.A (n_255), .B (n_390), .S0 (n_383), .Y (n_384));
NAND2X1 g11192(.A (n_318), .B (n_1212), .Y (n_381));
INVX1 g11197(.A (n_380), .Y (n_393));
NAND2X1 g11204(.A (n_328), .B (n_288), .Y (n_399));
INVX1 g10880(.A (n_377), .Y (n_378));
OAI21X1 g11238(.A0 (g578), .A1 (n_581), .B0 (n_313), .Y (n_376));
XOR2X1 g10918(.A (g622), .B (n_348), .Y (n_374));
XOR2X1 g10947(.A (g606), .B (n_345), .Y (n_372));
NAND2X1 g10973(.A (n_301), .B (n_371), .Y (n_411));
AND2X1 g10977(.A (n_303), .B (g638), .Y (n_370));
DFFSRX1 g634_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_298), .Q (g634), .QN ());
OAI21X1 g11082(.A0 (n_302), .A1 (g279), .B0 (n_341), .Y (n_369));
DFFSRX1 g616_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_304), .Q (g616), .QN ());
AOI22X1 g11122(.A0 (n_1099), .A1 (g465), .B0 (n_358), .B1 (n_383), .Y(n_368));
INVX1 g11127(.A (n_337), .Y (n_389));
INVX1 g11132(.A (n_367), .Y (n_388));
OR2X1 g11139(.A (n_128), .B (n_1165), .Y (n_366));
OAI21X1 g11163(.A0 (n_164), .A1 (g278), .B0 (n_291), .Y (n_365));
NAND3X1 g11168(.A (n_279), .B (n_241), .C (n_244), .Y (n_364));
AND2X1 g11191(.A (n_240), .B (n_359), .Y (n_360));
NAND2X1 g11133(.A (n_358), .B (n_1018), .Y (n_367));
NOR2X1 g11198(.A (n_1245), .B (g685), .Y (n_380));
INVX1 g11201(.A (n_356), .Y (n_1252));
AND2X1 g11217(.A (n_1018), .B (n_354), .Y (n_355));
NAND2X1 g11232(.A (n_267), .B (n_239), .Y (n_353));
OAI21X1 g11234(.A0 (g578), .A1 (n_271), .B0 (n_231), .Y (n_352));
NAND2X1 g11237(.A (n_238), .B (n_266), .Y (n_351));
NAND2X1 g11280(.A (g697), .B (n_1242), .Y (n_949));
NAND2X1 g11314(.A (g697), .B (n_220), .Y (n_960));
NAND2X1 g10924(.A (n_348), .B (g622), .Y (n_377));
INVX1 g11412(.A (n_767), .Y (n_347));
AND2X1 g10976(.A (n_345), .B (g606), .Y (n_398));
XOR2X1 g11052(.A (g619), .B (n_199), .Y (n_344));
OAI21X1 g11080(.A0 (n_293), .A1 (g207), .B0 (n_300), .Y (n_343));
INVX1 g11093(.A (n_341), .Y (n_342));
NAND2X1 g11128(.A (n_1099), .B (n_240), .Y (n_337));
XOR2X1 g11150(.A (n_62), .B (n_195), .Y (n_334));
AND2X1 g11187(.A (n_331), .B (n_359), .Y (n_332));
AND2X1 g11189(.A (n_21), .B (g471), .Y (n_424));
NAND4X1 g11200(.A (g266), .B (n_329), .C (g41), .D (n_159), .Y(n_330));
MX2X1 g11202(.A (n_182), .B (n_181), .S0 (n_148), .Y (n_356));
NAND2X1 g11210(.A (n_179), .B (n_210), .Y (n_328));
AND2X1 g11224(.A (n_320), .B (g687), .Y (n_322));
AND2X1 g11226(.A (n_320), .B (n_104), .Y (n_321));
NAND2X1 g11233(.A (n_218), .B (n_219), .Y (n_318));
MX2X1 g11235(.A (n_1092), .B (n_832), .S0 (g578), .Y (n_317));
MX2X1 g11236(.A (n_765), .B (n_767), .S0 (g578), .Y (n_316));
INVX1 g11270(.A (n_273), .Y (n_315));
INVX1 g11276(.A (n_272), .Y (n_314));
NAND2X1 g11288(.A (g578), .B (n_312), .Y (n_313));
INVX1 g11318(.A (n_985), .Y (n_311));
INVX1 g11161(.A (n_1165), .Y (n_696));
DFFSRX1 g613_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_251), .Q (g613), .QN ());
AND2X1 g11057(.A (n_252), .B (g639), .Y (n_304));
XOR2X1 g11087(.A (g642), .B (n_253), .Y (n_303));
DFFSRX1 g598_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_200), .Q (g598), .QN ());
NAND2X1 g11095(.A (n_302), .B (g279), .Y (n_341));
INVX1 g11096(.A (n_300), .Y (n_301));
DFFSRX1 g610_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_247), .Q (g610), .QN ());
AND2X1 g11109(.A (n_250), .B (g638), .Y (n_298));
NAND2X1 g11155(.A (n_162), .B (n_1204), .Y (n_358));
NOR2X1 g11316(.A (g683), .B (n_1247), .Y (n_406));
AOI21X1 g11164(.A0 (n_1097), .A1 (n_1218), .B0 (n_293), .Y (n_295));
NOR2X1 g11167(.A (n_192), .B (n_169), .Y (n_292));
INVX1 g11175(.A (n_302), .Y (n_291));
NAND2X1 g11211(.A (n_180), .B (n_1140), .Y (n_288));
INVX1 g11213(.A (n_286), .Y (n_287));
NAND2X1 g11216(.A (n_329), .B (n_1183), .Y (n_285));
NAND2X1 g11223(.A (n_280), .B (g678), .Y (n_282));
NAND2X1 g11225(.A (n_280), .B (n_147), .Y (n_281));
AOI21X1 g11242(.A0 (g260), .A1 (g532), .B0 (n_187), .Y (n_279));
AOI21X1 g11245(.A0 (g254), .A1 (g528), .B0 (n_189), .Y (n_278));
NAND2X1 g11267(.A (n_832), .B (n_1242), .Y (n_275));
NOR2X1 g11271(.A (n_271), .B (n_215), .Y (n_273));
NOR2X1 g11277(.A (n_271), .B (n_235), .Y (n_272));
NOR2X1 g11286(.A (n_226), .B (g_4325), .Y (n_270));
NOR2X1 g11302(.A (n_226), .B (n_1230), .Y (n_269));
INVX1 g11310(.A (n_216), .Y (n_267));
INVX1 g11312(.A (n_213), .Y (n_266));
NAND2X1 g11320(.A (n_211), .B (n_146), .Y (n_942));
INVX1 g11208(.A (g471), .Y (n_255));
NOR2X1 g11062(.A (n_198), .B (n_6), .Y (n_348));
NAND2X1 g11098(.A (n_293), .B (g207), .Y (n_300));
AND2X1 g11101(.A (n_253), .B (g642), .Y (n_345));
XOR2X1 g11148(.A (g616), .B (n_197), .Y (n_252));
NAND2X1 g11156(.A (n_167), .B (g639), .Y (n_251));
XOR2X1 g11173(.A (g634), .B (n_196), .Y (n_250));
AND2X1 g11176(.A (n_164), .B (g278), .Y (n_302));
NAND2X1 g11214(.A (n_116), .B (g478), .Y (n_286));
NAND2X1 g11219(.A (n_154), .B (n_137), .Y (n_247));
AOI21X1 g11228(.A0 (g520), .A1 (n_106), .B0 (n_170), .Y (n_246));
AOI21X1 g11240(.A0 (g224), .A1 (g508), .B0 (n_152), .Y (n_245));
AOI21X1 g11241(.A0 (g218), .A1 (g504), .B0 (n_156), .Y (n_244));
AOI21X1 g11243(.A0 (g248), .A1 (g524), .B0 (n_157), .Y (n_243));
AOI21X1 g11244(.A0 (g230), .A1 (g512), .B0 (n_158), .Y (n_242));
AOI21X1 g11246(.A0 (g500), .A1 (g212), .B0 (n_155), .Y (n_241));
INVX1 g11249(.A (n_240), .Y (n_331));
OR2X1 g11269(.A (n_172), .B (n_217), .Y (n_239));
OR2X1 g11273(.A (n_226), .B (n_217), .Y (n_238));
NAND2X1 g11275(.A (n_232), .B (n_214), .Y (n_237));
NAND2X1 g11281(.A (n_172), .B (n_235), .Y (n_236));
INVX1 g11292(.A (n_188), .Y (n_234));
OR2X1 g11295(.A (n_224), .B (n_232), .Y (n_233));
NAND2X1 g11296(.A (g578), .B (g696), .Y (n_231));
NAND2X1 g11297(.A (g696), .B (n_1242), .Y (n_955));
NAND2X1 g11299(.A (n_581), .B (n_232), .Y (n_228));
NAND2X1 g11301(.A (n_226), .B (n_235), .Y (n_227));
NOR2X1 g11303(.A (n_224), .B (g_4325), .Y (n_225));
INVX1 g11306(.A (n_186), .Y (n_219));
OR2X1 g11309(.A (n_224), .B (n_217), .Y (n_218));
NOR2X1 g11311(.A (n_215), .B (n_214), .Y (n_216));
NOR2X1 g11313(.A (n_581), .B (n_215), .Y (n_213));
NOR2X1 g11317(.A (n_211), .B (g698), .Y (n_320));
INVX1 g11327(.A (n_1139), .Y (n_210));
INVX1 g11347(.A (n_226), .Y (n_312));
INVX1 g11426(.A (n_765), .Y (n_256));
DFFSRX1 g471_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g664), .Q (), .QN (g471));
NAND2X1 g11215(.A (g638), .B (g567), .Y (g4121));
AND2X1 g11193(.A (n_103), .B (g638), .Y (n_200));
INVX1 g11121(.A (n_198), .Y (n_199));
NAND2X1 g11154(.A (n_197), .B (g616), .Y (n_198));
NOR2X1 g11177(.A (n_1097), .B (n_1218), .Y (n_293));
AND2X1 g11178(.A (n_196), .B (g634), .Y (n_253));
XOR2X1 g11205(.A (n_95), .B (n_94), .Y (n_195));
AOI22X1 g11227(.A0 (n_8), .A1 (g242), .B0 (g236), .B1 (g516), .Y(n_194));
INVX1 g11428(.A (n_214), .Y (n_765));
INVX1 g11258(.A (g478), .Y (n_390));
NAND3X1 g11268(.A (g578), .B (n_432), .C (n_27), .Y (n_192));
OR2X1 g11272(.A (n_141), .B (n_217), .Y (n_191));
OAI21X1 g11274(.A0 (n_235), .A1 (n_82), .B0 (n_1203), .Y (n_190));
NOR2X1 g11278(.A (n_11), .B (n_136), .Y (n_329));
NOR2X1 g11291(.A (g254), .B (g528), .Y (n_189));
NOR2X1 g11293(.A (n_1091), .B (n_235), .Y (n_188));
NOR2X1 g11294(.A (g260), .B (g532), .Y (n_187));
NOR2X1 g11307(.A (n_1091), .B (n_215), .Y (n_186));
OR2X1 g11308(.A (n_141), .B (n_232), .Y (n_184));
NOR2X1 g11315(.A (n_211), .B (n_146), .Y (n_283));
NOR2X1 g11321(.A (g679), .B (g678), .Y (n_183));
NOR2X1 g11322(.A (n_105), .B (g679), .Y (n_280));
NAND2X2 g11326(.A (n_107), .B (n_1102), .Y (n_240));
INVX1 g11331(.A (n_181), .Y (n_182));
INVX1 g11333(.A (n_179), .Y (n_180));
INVX2 g11366(.A (g697), .Y (n_271));
INVX1 g11352(.A (n_224), .Y (n_832));
INVX1 g11417(.A (n_172), .Y (n_767));
NOR2X1 g11305(.A (g236), .B (g516), .Y (n_170));
NAND2X1 g11190(.A (n_149), .B (n_168), .Y (n_169));
XOR2X1 g11229(.A (g613), .B (n_133), .Y (n_167));
INVX1 g11384(.A (g677), .Y (n_175));
DFFSRX1 g602_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_153), .Q (g602), .QN ());
INVX1 g11251(.A (n_1203), .Y (n_164));
DFFSRX1 g638_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g667), .Q (g638), .QN ());
AND2X1 g11265(.A (g280), .B (n_161), .Y (n_163));
AND2X1 g11282(.A (n_126), .B (n_161), .Y (n_162));
AND2X1 g11283(.A (n_159), .B (g662), .Y (n_160));
NOR2X1 g11284(.A (g230), .B (g512), .Y (n_158));
OR2X1 g11285(.A (g22), .B (g675), .Y (n_248));
NOR2X1 g11287(.A (g248), .B (g524), .Y (n_157));
NOR2X1 g11289(.A (g218), .B (g504), .Y (n_156));
NOR2X1 g11290(.A (g500), .B (g212), .Y (n_155));
INVX2 g11435(.A (g695), .Y (n_581));
NAND2X1 g11298(.A (n_153), .B (g610), .Y (n_154));
NOR2X1 g11300(.A (g224), .B (g508), .Y (n_152));
AOI21X1 g11324(.A0 (n_150), .A1 (g594), .B0 (n_149), .Y (n_151));
AOI21X1 g11325(.A0 (n_74), .A1 (n_73), .B0 (n_75), .Y (n_148));
NAND2X1 g11332(.A (n_961), .B (n_962), .Y (n_181));
NAND2X1 g11334(.A (n_67), .B (n_90), .Y (n_179));
INVX1 g11349(.A (g694), .Y (n_226));
INVX1 g11353(.A (g692), .Y (n_224));
INVX1 g11355(.A (g678), .Y (n_147));
DFFSRX1 g697_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_144), .Q (g697), .QN ());
DFFSRX1 g684_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_144), .Q (g684), .QN ());
INVX1 g11429(.A (g691), .Y (n_214));
DFFSRX1 g266_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_70), .Q (g266), .QN ());
NAND2X1 g11471(.A (n_1212), .B (n_217), .Y (n_143));
DFFSRX1 g664_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g663), .Q (g664), .QN ());
DFFSRX1 g478_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g665), .Q (), .QN (g478));
INVX1 g11418(.A (g690), .Y (n_172));
DFFSRX1 g658_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_98), .Q (g658), .QN ());
INVX1 g11398(.A (g681), .Y (n_139));
DFFSRX1 g260_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_39), .Q (), .QN (g260));
NAND3X1 g11279(.A (g639), .B (g602), .C (n_0), .Y (n_137));
INVX1 g11340(.A (g1293), .Y (n_136));
DFFSRX1 g254_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_31), .Q (), .QN (g254));
NOR2X1 g11266(.A (n_133), .B (n_46), .Y (n_197));
INVX1 g11392(.A (g689), .Y (n_211));
DFFSRX1 g679_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_117), .Q (g679), .QN ());
DFFSRX1 g681_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_115), .Q (), .QN (g681));
INVX1 g11403(.A (g688), .Y (n_145));
DFFSRX1 g695_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_120), .Q (g695), .QN ());
NAND2X1 g11444(.A (g280), .B (n_86), .Y (n_131));
OR2X1 g11446(.A (n_129), .B (g210), .Y (n_130));
NAND2X1 g11447(.A (g283), .B (n_96), .Y (n_128));
NAND2X1 g11454(.A (n_126), .B (g281), .Y (n_127));
NAND2X2 g11445(.A (n_101), .B (n_15), .Y (n_122));
INVX1 g11550(.A (n_1051), .Y (n_675));
INVX1 g11360(.A (g698), .Y (n_146));
DFFSRX1 g678_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_109), .Q (g678), .QN ());
DFFSRX1 g682_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_120), .Q (), .QN (g682));
DFFSRX1 g690_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_108), .Q (g690), .QN ());
OR2X1 g11461(.A (g41), .B (g22), .Y (n_119));
DFFSRX1 g692_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_117), .Q (g692), .QN ());
NOR2X1 g11470(.A (g283), .B (g282), .Y (n_116));
DFFSRX1 g694_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_115), .Q (g694), .QN ());
DFFSRX1 g691_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_109), .Q (g691), .QN ());
DFFSRX1 g677_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_108), .Q (g677), .QN ());
INVX1 g11410(.A (g696), .Y (n_141));
NAND2X1 g11443(.A (n_371), .B (n_60), .Y (n_107));
INVX1 g11394(.A (g242), .Y (n_106));
INVX1 g11386(.A (g680), .Y (n_105));
INVX1 g11390(.A (g687), .Y (n_104));
INVX1 g11547(.A (n_66), .Y (n_220));
XOR2X1 g11253(.A (g598), .B (g567), .Y (n_103));
OR2X1 g11253_or(.A (g598), .B (g567), .Y (n_196));
NAND2X1 g11458(.A (n_18), .B (g_5709), .Y (n_961));
CLKBUFX1 g11570(.A (n_101), .Y (n_144));
AND2X1 g11442(.A (n_159), .B (g45), .Y (n_98));
DFFSRX1 g663_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g42), .Q (g663), .QN ());
XOR2X1 g11329(.A (g36), .B (g32), .Y (n_95));
XOR2X1 g11330(.A (g38), .B (g37), .Y (n_94));
DFFSRX1 g698_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g40), .Q (g698), .QN ());
DFFSRX1 g662_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_69), .Q (g662), .QN ());
DFFSRX1 g693_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_93), .Q (g693), .QN ());
DFFSRX1 g680_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_93), .Q (), .QN (g680));
DFFSRX1 g683_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_76), .Q (), .QN (g683));
DFFSRX1 g218_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g598), .Q (), .QN (g218));
DFFSRX1 g675_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g702), .Q (), .QN (g675));
NAND2X1 g11450(.A (n_30), .B (g_6081), .Y (n_90));
NOR2X1 g11448(.A (n_49), .B (g602), .Y (n_153));
DFFSRX1 g248_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g650), .Q (), .QN (g248));
NOR2X1 g11460(.A (g283), .B (n_96), .Y (n_354));
NOR2X1 g11465(.A (n_1181), .B (n_86), .Y (n_161));
INVX1 g11481(.A (n_1191), .Y (n_82));
DFFSRX1 g230_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g642), .Q (), .QN (g230));
DFFSRX1 g666_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g46), .Q (g1290), .QN ());
NOR2X1 g11449(.A (n_10), .B (g102), .Y (g2584));
INVX2 g11615(.A (n_77), .Y (n_217));
DFFSRX1 g696_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_76), .Q (g696), .QN ());
DFFSRX1 g685_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g32), .Q (), .QN (g685));
NOR2X1 g11463(.A (n_74), .B (n_73), .Y (n_75));
DFFSRX1 g699_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(n_4), .Q (g1293), .QN ());
AND2X1 g11452(.A (n_69), .B (g45), .Y (n_70));
DFFSRX1 g667_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g45), .Q (g667), .QN ());
NAND2X1 g11453(.A (g18), .B (n_57), .Y (n_67));
DFFSRX1 g689_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g39), .Q (g689), .QN ());
DFFSRX1 g688_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g38), .Q (g688), .QN ());
DFFSRX1 g236_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g606), .Q (), .QN (g236));
DFFSRX1 g212_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g567), .Q (), .QN (g212));
DFFSRX1 g242_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g646), .Q (g242), .QN ());
DFFSRX1 g687_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g37), .Q (g687), .QN ());
DFFSRX1 g665_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g42), .Q (g665), .QN ());
NAND2X1 g11457(.A (n_41), .B (g24), .Y (n_64));
AND2X1 g11441(.A (n_129), .B (g210), .Y (n_359));
XOR2X1 g11335(.A (g39), .B (g40), .Y (n_62));
DFFSRX1 g224_reg(.RN (n_930), .SN (1'b1), .CK (blif_clk_net), .D(g634), .Q (), .QN (g224));
NOR2X1 g11451(.A (n_150), .B (g594), .Y (n_149));
NAND2X1 g11459(.A (n_32), .B (g_739), .Y (n_962));
INVX1 g11501(.A (n_57), .Y (n_115));
INVX1 g11496(.A (n_74), .Y (n_108));
INVX1 g11514(.A (n_73), .Y (n_109));
INVX2 g11488(.A (n_232), .Y (n_235));
INVX2 g11571(.A (n_41), .Y (n_101));
INVX2 g11616(.A (n_38), .Y (n_77));
INVX1 g11617(.A (n_38), .Y (n_215));
INVX1 g11593(.A (n_32), .Y (n_117));
NAND2X1 g11467(.A (g602), .B (g610), .Y (n_133));
INVX1 g11519(.A (n_30), .Y (n_120));
INVX1 g11549(.A (n_1051), .Y (n_66));
NOR2X1 g11464(.A (g211), .B (g210), .Y (n_21));
INVX1 g11581(.A (g430), .Y (n_594));
INVX1 g11631(.A (n_371), .Y (n_26));
INVX1 g11580(.A (g283), .Y (n_58));
INVX1 g11475(.A (g551), .Y (n_567));
INVX2 g11572(.A (g_4785), .Y (n_41));
INVX1 g11508(.A (g528), .Y (n_20));
INVX1 g11521(.A (g449), .Y (n_601));
INVX1 g11583(.A (g541), .Y (n_536));
INVX1 g11591(.A (g281), .Y (n_86));
INVX1 g11561(.A (g434), .Y (n_528));
INVX1 g11528(.A (g536), .Y (n_465));
INVX1 g11585(.A (blif_reset_net), .Y (n_930));
INVX1 g11562(.A (g426), .Y (n_610));
INVX1 g11608(.A (g_739), .Y (n_18));
INVX1 g11536(.A (g654), .Y (n_31));
INVX1 g11566(.A (g422), .Y (n_612));
INVX1 g11582(.A (g554), .Y (n_563));
INVX1 g11589(.A (g571), .Y (n_39));
INVX1 g11609(.A (g590), .Y (n_150));
INVX1 g11477(.A (g639), .Y (n_49));
INVX1 g11473(.A (g508), .Y (n_16));
INVX1 g11594(.A (g_5709), .Y (n_32));
INVX1 g11524(.A (g24), .Y (n_15));
INVX1 g11576(.A (g437), .Y (n_607));
INVX2 g11618(.A (g204), .Y (n_38));
INVX1 g11596(.A (g414), .Y (n_616));
INVX1 g11502(.A (g_6081), .Y (n_57));
INVX1 g11574(.A (g209), .Y (n_60));
INVX1 g11529(.A (g293), .Y (n_516));
INVX1 g11592(.A (g266), .Y (n_69));
INVX1 g11601(.A (g282), .Y (n_96));
INVX1 g11480(.A (g496), .Y (n_40));
INVX1 g11564(.A (g418), .Y (n_614));
INVX1 g11558(.A (g658), .Y (n_159));
INVX1 g11500(.A (g280), .Y (n_126));
INVX1 g11497(.A (g_5464), .Y (n_74));
INVX1 g11587(.A (g445), .Y (n_603));
INVX1 g11624(.A (g516), .Y (n_13));
INVX1 g11492(.A (g672), .Y (n_626));
INVX1 g11522(.A (g702), .Y (n_11));
INVX1 g11575(.A (g545), .Y (n_561));
INVX1 g11598(.A (g89), .Y (n_10));
INVX1 g11560(.A (g410), .Y (n_618));
INVX1 g11586(.A (g457), .Y (n_597));
INVX1 g11504(.A (g586), .Y (n_27));
INVX1 g11517(.A (g520), .Y (n_8));
INVX1 g11602(.A (g492), .Y (n_507));
INVX1 g11518(.A (g402), .Y (n_623));
INVX1 g11474(.A (g669), .Y (n_630));
INVX1 g11577(.A (g512), .Y (n_7));
INVX1 g11567(.A (g619), .Y (n_6));
INVX1 g11546(.A (g631), .Y (n_5));
INVX1 g11559(.A (g47), .Y (n_4));
INVX1 g11557(.A (g210), .Y (n_50));
INVX1 g11606(.A (g461), .Y (n_595));
INVX1 g11515(.A (g_1196), .Y (n_73));
INVX1 g11520(.A (g18), .Y (n_30));
INVX1 g11563(.A (g625), .Y (n_2));
INVX1 g11595(.A (g453), .Y (n_599));
INVX1 g11526(.A (g613), .Y (n_46));
INVX1 g11623(.A (g406), .Y (n_620));
INVX1 g11632(.A (g524), .Y (n_1));
CLKBUFX1 g11523(.A (g24), .Y (n_76));
CLKBUFX1 g11607(.A (g_739), .Y (n_93));
INVX1 g11597(.A (g441), .Y (n_605));
INVX1 g11584(.A (g297), .Y (n_518));
INVX1 g11611(.A (g211), .Y (n_129));
INVX1 g11621(.A (g465), .Y (n_383));
INVX1 g11565(.A (g610), .Y (n_0));
INVX1 g11534(.A (g574), .Y (n_168));
INVX1 g11568(.A (g548), .Y (n_571));
INVX1 g11787(.A (n_987), .Y (n_988));
AND2X1 g11788(.A (n_985), .B (n_986), .Y (n_987));
NAND2X1 g53(.A (n_145), .B (g687), .Y (n_985));
NAND2X1 g52(.A (n_145), .B (n_104), .Y (n_986));
NOR2X1 g49(.A (n_942), .B (n_711), .Y (n_989));
NAND2X1 g27(.A (n_1004), .B (n_1009), .Y (n_1250));
AOI21X1 g29(.A0 (n_871), .A1 (n_872), .B0 (n_1003), .Y (n_1004));
NOR2X1 g30(.A (n_141), .B (n_805), .Y (n_1003));
NAND2X1 g28(.A (n_1054), .B (n_1008), .Y (n_1009));
INVX2 g31(.A (n_1007), .Y (n_1008));
INVX2 g11794(.A (n_1006), .Y (n_1007));
NOR2X1 g33(.A (n_986), .B (n_939), .Y (n_1006));
INVX1 g11797(.A (n_1013), .Y (n_1014));
NAND3X1 g11798(.A (n_127), .B (n_131), .C (n_1012), .Y (n_1013));
NOR2X1 g11799(.A (n_96), .B (n_58), .Y (n_1012));
INVX1 g11801(.A (n_1018), .Y (n_1019));
NAND2X1 g11802(.A (n_127), .B (n_131), .Y (n_1018));
AND2X1 g11805(.A (g209), .B (n_371), .Y (n_1020));
INVX1 g19(.A (n_1031), .Y (n_1032));
NAND3X1 g20(.A (n_160), .B (n_1030), .C (g676), .Y (n_1031));
AND2X1 g11812(.A (n_329), .B (g41), .Y (n_1030));
NAND2X1 g21(.A (n_1030), .B (n_160), .Y (n_1036));
NOR2X1 g16(.A (n_445), .B (n_1038), .Y (n_1039));
NAND3X1 g17(.A (g631), .B (n_432), .C (g578), .Y (n_1038));
NAND2X1 g11816(.A (n_1041), .B (g578), .Y (n_1042));
NOR2X1 g11817(.A (n_445), .B (n_5), .Y (n_1041));
INVX1 g11818(.A (n_432), .Y (n_404));
INVX2 g11823(.A (n_1053), .Y (n_1054));
NOR2X1 g11824(.A (n_1050), .B (n_1052), .Y (n_1053));
AND2X1 g11825(.A (n_220), .B (g696), .Y (n_1050));
AOI21X1 g11826(.A0 (n_839), .A1 (n_851), .B0 (n_1051), .Y (n_1052));
INVX1 g11827(.A (g_4325), .Y (n_1051));
NAND2X1 g11829(.A (n_851), .B (n_839), .Y (n_1056));
NAND2X1 g11836(.A (n_424), .B (n_337), .Y (n_1062));
OR2X1 g11837(.A (n_130), .B (n_1196), .Y (n_1064));
INVX2 g13(.A (g276), .Y (n_232));
AND2X1 g11841(.A (n_738), .B (n_1134), .Y (n_1071));
NAND2X2 g11843(.A (n_710), .B (n_321), .Y (n_1072));
NAND3X1 g11844(.A (n_717), .B (n_1246), .C (g684), .Y (n_1073));
NAND2X1 g11845(.A (n_988), .B (n_989), .Y (n_1075));
NOR2X1 g11846(.A (n_532), .B (n_533), .Y (n_1076));
NAND2X2 g11851(.A (n_1252), .B (n_1253), .Y (n_1081));
NAND2X1 g11852(.A (n_399), .B (n_356), .Y (n_1082));
OAI21X1 g11853(.A0 (n_1087), .A1 (n_1089), .B0 (n_1093), .Y (n_1094));
CLKBUFX3 g26(.A (n_1086), .Y (n_1087));
AND2X1 g11854(.A (n_175), .B (n_729), .Y (n_1086));
AOI21X1 g11855(.A0 (n_426), .A1 (n_505), .B0 (n_536), .Y (n_1089));
NAND2X1 g11856(.A (n_1092), .B (n_1087), .Y (n_1093));
INVX1 g11857(.A (n_1091), .Y (n_1092));
INVX1 g11859(.A (g693), .Y (n_1091));
OR2X1 g11860(.A (n_1097), .B (n_1098), .Y (n_1099));
NAND2X2 g11861(.A (n_1095), .B (g_4890), .Y (n_1097));
INVX1 g11862(.A (n_38), .Y (n_1095));
NAND4X1 g11864(.A (n_26), .B (g209), .C (g207), .D (g206), .Y(n_1098));
INVX1 g11866(.A (g207), .Y (n_1100));
NAND2X1 g11867(.A (n_26), .B (g209), .Y (n_1102));
NAND2X2 g11869(.A (n_1104), .B (n_1105), .Y (n_1106));
NAND2X1 g11870(.A (n_1167), .B (n_1014), .Y (n_1104));
NAND3X1 g11871(.A (n_469), .B (n_1018), .C (n_1012), .Y (n_1105));
INVX1 g11874(.A (n_1111), .Y (n_1112));
NAND2X2 g11875(.A (n_1109), .B (n_1170), .Y (n_1111));
NAND2X2 g11876(.A (n_1106), .B (n_1165), .Y (n_1109));
NAND4X1 g34(.A (n_1128), .B (n_724), .C (n_548), .D (n_698), .Y(n_1115));
AND2X1 g11878(.A (n_1113), .B (g283), .Y (n_1128));
AND2X1 g11879(.A (n_490), .B (n_366), .Y (n_1113));
NAND3X1 g11880(.A (n_698), .B (n_724), .C (n_1113), .Y (n_1117));
INVX1 g11882(.A (n_1121), .Y (n_1122));
NAND3X1 g11883(.A (n_1118), .B (n_1119), .C (n_1120), .Y (n_1121));
AND2X1 g11884(.A (n_1020), .B (g206), .Y (n_1118));
NOR2X1 g11885(.A (n_1100), .B (n_1097), .Y (n_1119));
NOR2X1 g11886(.A (n_129), .B (n_50), .Y (n_1120));
NAND2X1 g37_dup(.A (n_1123), .B (n_1124), .Y (n_1125));
NAND2X1 g11887(.A (n_486), .B (n_240), .Y (n_1123));
NAND2X2 g11888(.A (n_669), .B (n_331), .Y (n_1124));
NAND2X1 g11889(.A (n_1124), .B (n_1123), .Y (n_1127));
NAND3X1 g10786_dup(.A (n_1244), .B (n_1246), .C (n_1247), .Y(n_1134));
MX2X1 g11891(.A (n_1187), .B (g48), .S0 (n_1188), .Y (n_1135));
AND2X1 g11892(.A (n_1072), .B (n_1073), .Y (n_1137));
AND2X1 g11842_dup(.A (n_1072), .B (n_1073), .Y (n_1138));
NAND2X1 g11893(.A (n_122), .B (n_64), .Y (n_1139));
NAND2X1 g11328_dup(.A (n_122), .B (n_64), .Y (n_1140));
NAND4X1 g11894(.A (n_1256), .B (n_1146), .C (n_546), .D (n_517), .Y(n_1147));
AND2X1 g11896(.A (n_1076), .B (n_1143), .Y (n_1144));
NOR2X1 g11897(.A (n_673), .B (n_1142), .Y (n_1143));
OR2X1 g11898(.A (n_647), .B (n_1141), .Y (n_1142));
OR2X1 g11899(.A (n_635), .B (n_636), .Y (n_1141));
OR2X1 g51(.A (n_16), .B (n_481), .Y (n_1146));
NOR2X1 g50(.A (n_1148), .B (n_1149), .Y (n_1150));
NAND2X1 g11900(.A (n_1075), .B (n_1076), .Y (n_1148));
NAND2X1 g54(.A (n_1137), .B (n_1071), .Y (n_1149));
NAND2X2 g11907(.A (n_1162), .B (n_1163), .Y (n_1164));
INVX1 g11908(.A (n_1160), .Y (n_1162));
NAND2X1 g11910(.A (n_1158), .B (g676), .Y (n_1160));
NAND2X1 g11911(.A (n_1135), .B (n_1183), .Y (n_1158));
NOR2X1 g11914(.A (n_1183), .B (n_248), .Y (n_1163));
NAND2X1 g11915(.A (n_1165), .B (n_1169), .Y (n_1170));
NAND2X1 g11916(.A (n_1204), .B (n_163), .Y (n_1165));
NOR2X1 g25_dup(.A (n_1166), .B (n_1168), .Y (n_1169));
NAND2X1 g11917(.A (n_1019), .B (n_354), .Y (n_1166));
INVX1 g11918(.A (n_1167), .Y (n_1168));
MX2X1 g11919(.A (g478), .B (n_390), .S0 (n_479), .Y (n_1167));
NOR2X1 g11920(.A (n_1166), .B (n_1168), .Y (n_1171));
NAND2X1 g11921(.A (n_1175), .B (n_1178), .Y (n_1179));
AND2X1 g11922(.A (n_1181), .B (n_1174), .Y (n_1175));
NAND3X1 g11924(.A (n_228), .B (n_227), .C (g277), .Y (n_1174));
NAND2X1 g11926(.A (n_1176), .B (n_1191), .Y (n_1178));
NAND2X1 g11927(.A (n_184), .B (n_314), .Y (n_1176));
INVX1 g11930(.A (g278), .Y (n_1181));
OR2X1 g11931(.A (n_1182), .B (n_1185), .Y (n_1186));
AOI21X1 g11932(.A0 (n_1081), .A1 (n_1082), .B0 (g48), .Y (n_1182));
NAND2X1 g11933(.A (n_1183), .B (n_1184), .Y (n_1185));
INVX1 g11934(.A (g41), .Y (n_1183));
NAND3X1 g11935(.A (n_1081), .B (n_1082), .C (g48), .Y (n_1184));
INVX1 g11936(.A (g48), .Y (n_1187));
NAND2X1 g11937(.A (n_1082), .B (n_1081), .Y (n_1188));
NAND3X1 g11938(.A (n_1192), .B (n_1193), .C (g278), .Y (n_1194));
NAND2X1 g11939(.A (n_1189), .B (n_1191), .Y (n_1192));
NAND2X1 g11940(.A (n_233), .B (n_234), .Y (n_1189));
INVX1 g11941(.A (g277), .Y (n_1191));
NAND3X1 g11943(.A (n_237), .B (n_236), .C (g277), .Y (n_1193));
AND2X1 g11945(.A (n_332), .B (n_669), .Y (n_1195));
NAND2X1 g11946(.A (n_1118), .B (n_1119), .Y (n_1196));
INVX1 g11947(.A (n_1198), .Y (n_1199));
NAND2X1 g11948(.A (n_1127), .B (n_1197), .Y (n_1198));
AND2X1 g11949(.A (n_1196), .B (n_1120), .Y (n_1197));
NOR2X1 g9(.A (n_1202), .B (n_1203), .Y (n_1204));
INVX1 g15(.A (g279), .Y (n_1202));
NAND2X1 g11951(.A (g277), .B (g276), .Y (n_1203));
NAND3X1 g11958(.A (n_1215), .B (n_1217), .C (n_1218), .Y (n_1219));
NAND2X1 g11959(.A (n_351), .B (g_4890), .Y (n_1215));
INVX1 g11962(.A (g_4890), .Y (n_1212));
NAND2X1 g11963(.A (n_1216), .B (n_1212), .Y (n_1217));
NAND2X1 g11964(.A (n_191), .B (n_315), .Y (n_1216));
INVX1 g11965(.A (g206), .Y (n_1218));
NAND2X1 g35(.A (n_1220), .B (n_1226), .Y (n_1227));
AOI21X1 g11966(.A0 (n_1195), .A1 (n_1196), .B0 (n_1199), .Y (n_1220));
NAND3X1 g11967(.A (n_1221), .B (n_1222), .C (n_1225), .Y (n_1226));
NAND2X1 g11968(.A (n_1195), .B (n_425), .Y (n_1221));
NAND2X1 g11969(.A (n_1125), .B (n_1122), .Y (n_1222));
NOR2X1 g11970(.A (n_577), .B (n_1224), .Y (n_1225));
NAND3X1 g11971(.A (n_1064), .B (n_1062), .C (g211), .Y (n_1224));
NAND4X1 g11973(.A (n_1221), .B (n_1222), .C (n_1064), .D (n_1062), .Y(n_1228));
NAND2X2 g11974(.A (n_1230), .B (n_1232), .Y (n_1233));
INVX1 g11975(.A (n_1242), .Y (n_1230));
NAND3X1 g11977(.A (n_1115), .B (n_1112), .C (n_1235), .Y (n_1232));
NAND2X2 g11980(.A (n_1239), .B (g269), .Y (n_1241));
NAND2X2 g11981(.A (n_1237), .B (n_1238), .Y (n_1239));
NOR2X1 g11982(.A (n_1236), .B (n_753), .Y (n_1237));
INVX1 g11983(.A (n_1235), .Y (n_1236));
NAND3X1 g11984(.A (n_685), .B (n_696), .C (n_354), .Y (n_1235));
INVX1 g11985(.A (n_1117), .Y (n_1238));
INVX1 g11987(.A (g269), .Y (n_1242));
NAND3X1 g11988(.A (n_1244), .B (n_1246), .C (n_1247), .Y (n_1248));
INVX1 g11989(.A (n_1243), .Y (n_1244));
NAND3X1 g11990(.A (g685), .B (n_1032), .C (n_1186), .Y (n_1243));
INVX1 g11991(.A (n_1245), .Y (n_1246));
NAND2X1 g11992(.A (n_283), .B (n_145), .Y (n_1245));
INVX1 g11993(.A (g684), .Y (n_1247));
AND2X1 g11994(.A (n_1186), .B (n_1032), .Y (n_1249));
NAND4X1 g11995(.A (n_1144), .B (n_1071), .C (n_1137), .D (n_1075), .Y(n_1256));
NAND4X1 g11895_dup(.A (n_1144), .B (n_1071), .C (n_1137), .D(n_1075), .Y (n_1257));
endmodule
