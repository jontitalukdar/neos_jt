module s35932(blif_clk_net, blif_reset_net, DATA_0_31, DATA_0_30, DATA_0_29, DATA_0_28, DATA_0_27, DATA_0_26, DATA_0_25, DATA_0_24, DATA_0_23, DATA_0_22, DATA_0_21, DATA_0_20, DATA_0_19, DATA_0_18, DATA_0_17, DATA_0_16, DATA_0_15, DATA_0_14, DATA_0_13, DATA_0_12, DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8, DATA_0_7, DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2, DATA_0_1, DATA_0_0, RESET, TM1, TM0, DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27, DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22, DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17, DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12, DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7, DATA_9_6, DATA_9_5, DATA_9_4, DATA_9_3, DATA_9_2, DATA_9_1, DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2, CRC_OUT_9_3, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30, CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2, CRC_OUT_7_3, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2, CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2, CRC_OUT_2_3, CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_2, CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31, d_out_1, q_in_1, d_out_2, q_in_2, d_out_3, q_in_3, d_out_4, q_in_4, d_out_5, q_in_5, d_out_6, q_in_6, d_out_7, q_in_7, d_out_8, q_in_8, d_out_9, q_in_9, d_out_10, q_in_10, d_out_11, q_in_11, d_out_12, q_in_12, d_out_13, q_in_13, d_out_14, q_in_14, d_out_15, q_in_15, d_out_16, q_in_16, d_out_17, q_in_17, d_out_18, q_in_18, d_out_19, q_in_19, d_out_20, q_in_20, d_out_21, q_in_21, d_out_22, q_in_22, d_out_23, q_in_23, d_out_24, qn_in_24, d_out_25, qn_in_25, d_out_26, q_in_26, d_out_27, q_in_27, d_out_28, q_in_28, d_out_29, qn_in_29, d_out_30, qn_in_30, d_out_31, q_in_31, d_out_32, q_in_32, d_out_33, q_in_33, d_out_34, q_in_34, d_out_35, qn_in_35, d_out_36, qn_in_36, d_out_37, q_in_37, d_out_38, q_in_38, d_out_39, q_in_39, d_out_40, q_in_40, d_out_41, qn_in_41, d_out_42, qn_in_42, d_out_43, q_in_43, d_out_44, q_in_44, d_out_45, q_in_45, d_out_46, q_in_46, d_out_47, qn_in_47, d_out_48, qn_in_48, d_out_49, q_in_49, d_out_50, q_in_50, d_out_51, q_in_51, d_out_52, qn_in_52, d_out_53, qn_in_53, d_out_54, q_in_54, d_out_55, q_in_55, d_out_56, q_in_56, d_out_57, q_in_57, d_out_58, qn_in_58, d_out_59, qn_in_59, d_out_60, q_in_60, d_out_61, q_in_61, d_out_62, q_in_62, d_out_63, q_in_63, d_out_64, qn_in_64, d_out_65, qn_in_65, d_out_66, q_in_66, d_out_67, q_in_67, d_out_68, q_in_68, d_out_69, q_in_69, d_out_70, q_in_70, d_out_71, q_in_71, d_out_72, q_in_72, d_out_73, qn_in_73, d_out_74, qn_in_74, d_out_75, q_in_75, d_out_76, q_in_76, d_out_77, q_in_77, d_out_78, q_in_78, d_out_79, q_in_79, d_out_80, q_in_80, d_out_81, q_in_81, d_out_82, q_in_82, d_out_83, qn_in_83, d_out_84, qn_in_84, d_out_85, q_in_85, d_out_86, q_in_86, d_out_87, q_in_87, d_out_88, q_in_88, d_out_89, q_in_89, d_out_90, qn_in_90, d_out_91, q_in_91, d_out_92, q_in_92, d_out_93, q_in_93, d_out_94, q_in_94, d_out_95, q_in_95, d_out_96, q_in_96, d_out_97, qn_in_97, d_out_98, qn_in_98, d_out_99, q_in_99, d_out_100, q_in_100, d_out_101, q_in_101, d_out_102, q_in_102, d_out_103, q_in_103, d_out_104, qn_in_104, d_out_105, qn_in_105, d_out_106, q_in_106, d_out_107, q_in_107, d_out_108, q_in_108, d_out_109, q_in_109, d_out_110, q_in_110, d_out_111, qn_in_111, d_out_112, qn_in_112, d_out_113, q_in_113, d_out_114, q_in_114, d_out_115, q_in_115, d_out_116, q_in_116, d_out_117, q_in_117, d_out_118, q_in_118, d_out_119, q_in_119, d_out_120, q_in_120, d_out_121, qn_in_121, d_out_122, qn_in_122, d_out_123, qn_in_123, d_out_124, q_in_124, d_out_125, q_in_125, d_out_126, q_in_126, d_out_127, q_in_127, d_out_128, qn_in_128, d_out_129, qn_in_129, d_out_130, q_in_130, d_out_131, q_in_131, d_out_132, q_in_132, d_out_133, q_in_133, d_out_134, q_in_134, d_out_135, q_in_135, d_out_136, q_in_136, d_out_137, qn_in_137, d_out_138, qn_in_138, d_out_139, qn_in_139, d_out_140, qn_in_140, d_out_141, q_in_141, d_out_142, q_in_142, d_out_143, q_in_143, d_out_144, q_in_144, d_out_145, q_in_145, d_out_146, qn_in_146, d_out_147, qn_in_147, d_out_148, qn_in_148, d_out_149, q_in_149, d_out_150, q_in_150, d_out_151, q_in_151, d_out_152, q_in_152, d_out_153, q_in_153, d_out_154, q_in_154, d_out_155, qn_in_155, d_out_156, qn_in_156, d_out_157, qn_in_157, d_out_158, qn_in_158, d_out_159, qn_in_159, d_out_160, q_in_160, d_out_161, q_in_161, d_out_162, q_in_162, d_out_163, q_in_163, d_out_164, qn_in_164, d_out_165, qn_in_165, d_out_166, qn_in_166, d_out_167, q_in_167, d_out_168, q_in_168, d_out_169, q_in_169, d_out_170, q_in_170, d_out_171, q_in_171, d_out_172, qn_in_172, d_out_173, qn_in_173, d_out_174, qn_in_174, d_out_175, qn_in_175, d_out_176, qn_in_176, d_out_177, q_in_177, d_out_178, q_in_178, d_out_179, q_in_179, d_out_180, q_in_180, d_out_181, qn_in_181, d_out_182, qn_in_182, d_out_183, qn_in_183, d_out_184, q_in_184, d_out_185, q_in_185, d_out_186, q_in_186, d_out_187, q_in_187, d_out_188, q_in_188, d_out_189, q_in_189, d_out_190, q_in_190, d_out_191, qn_in_191, d_out_192, qn_in_192, d_out_193, qn_in_193, d_out_194, qn_in_194, d_out_195, q_in_195, d_out_196, q_in_196, d_out_197, q_in_197, d_out_198, qn_in_198, d_out_199, qn_in_199, d_out_200, q_in_200, d_out_201, qn_in_201, d_out_202, qn_in_202, d_out_203, q_in_203, d_out_204, q_in_204, d_out_205, q_in_205, d_out_206, q_in_206, d_out_207, q_in_207, d_out_208, q_in_208, d_out_209, q_in_209, d_out_210, q_in_210, d_out_211, qn_in_211, d_out_212, qn_in_212, d_out_213, qn_in_213, d_out_214, qn_in_214, d_out_215, qn_in_215, d_out_216, q_in_216, d_out_217, q_in_217, d_out_218, q_in_218, d_out_219, qn_in_219, d_out_220, qn_in_220, d_out_221, qn_in_221, d_out_222, qn_in_222, d_out_223, q_in_223, d_out_224, q_in_224, d_out_225, q_in_225, d_out_226, q_in_226, d_out_227, qn_in_227, d_out_228, q_in_228, d_out_229, q_in_229, d_out_230, q_in_230, d_out_231, q_in_231, d_out_232, q_in_232, d_out_233, qn_in_233, d_out_234, qn_in_234, d_out_235, qn_in_235, d_out_236, q_in_236, d_out_237, qn_in_237, d_out_238, qn_in_238, d_out_239, q_in_239, d_out_240, q_in_240, d_out_241, q_in_241, d_out_242, qn_in_242, d_out_243, qn_in_243, d_out_244, qn_in_244, d_out_245, qn_in_245, d_out_246, q_in_246, d_out_247, q_in_247, d_out_248, q_in_248, d_out_249, q_in_249, d_out_250, qn_in_250, d_out_251, qn_in_251, d_out_252, q_in_252, d_out_253, q_in_253, d_out_254, q_in_254, d_out_255, q_in_255, d_out_256, q_in_256, d_out_257, qn_in_257, d_out_258, q_in_258, d_out_259, qn_in_259, d_out_260, qn_in_260, d_out_261, qn_in_261, d_out_262, qn_in_262, d_out_263, q_in_263, d_out_264, q_in_264, d_out_265, q_in_265, d_out_266, qn_in_266, d_out_267, qn_in_267, d_out_268, qn_in_268, d_out_269, q_in_269, d_out_270, qn_in_270, d_out_271, q_in_271, d_out_272, q_in_272, d_out_273, q_in_273, d_out_274, q_in_274, d_out_275, q_in_275, d_out_276, qn_in_276, d_out_277, qn_in_277, d_out_278, qn_in_278, d_out_279, q_in_279, d_out_280, q_in_280, d_out_281, q_in_281, d_out_282, q_in_282, d_out_283, q_in_283, d_out_284, qn_in_284, d_out_285, qn_in_285, d_out_286, qn_in_286, d_out_287, qn_in_287, d_out_288, qn_in_288, d_out_289, qn_in_289, d_out_290, q_in_290, d_out_291, q_in_291, d_out_292, q_in_292, d_out_293, q_in_293, d_out_294, qn_in_294, d_out_295, qn_in_295, d_out_296, qn_in_296, d_out_297, q_in_297, d_out_298, q_in_298, d_out_299, q_in_299, d_out_300, q_in_300, d_out_301, q_in_301, d_out_302, q_in_302, d_out_303, q_in_303, d_out_304, qn_in_304, d_out_305, qn_in_305, d_out_306, qn_in_306, d_out_307, qn_in_307, d_out_308, q_in_308, d_out_309, q_in_309, d_out_310, q_in_310, d_out_311, q_in_311, d_out_312, q_in_312, d_out_313, qn_in_313, d_out_314, qn_in_314, d_out_315, qn_in_315, d_out_316, qn_in_316, d_out_317, qn_in_317, d_out_318, q_in_318, d_out_319, q_in_319, d_out_320, qn_in_320, d_out_321, q_in_321, d_out_322, qn_in_322, d_out_323, qn_in_323, d_out_324, qn_in_324, d_out_325, q_in_325, d_out_326, q_in_326, d_out_327, q_in_327, d_out_328, q_in_328, d_out_329, q_in_329, d_out_330, q_in_330, d_out_331, q_in_331, d_out_332, qn_in_332, d_out_333, qn_in_333, d_out_334, qn_in_334, d_out_335, qn_in_335, d_out_336, qn_in_336, d_out_337, q_in_337, d_out_338, q_in_338, d_out_339, q_in_339, d_out_340, q_in_340, d_out_341, q_in_341, d_out_342, q_in_342, d_out_343, qn_in_343, d_out_344, qn_in_344, d_out_345, qn_in_345, d_out_346, qn_in_346, d_out_347, qn_in_347, d_out_348, qn_in_348, d_out_349, q_in_349, d_out_350, q_in_350, d_out_351, q_in_351, d_out_352, qn_in_352, d_out_353, qn_in_353, d_out_354, qn_in_354, d_out_355, q_in_355, d_out_356, q_in_356, d_out_357, q_in_357, d_out_358, q_in_358, d_out_359, q_in_359, d_out_360, q_in_360, d_out_361, q_in_361, d_out_362, qn_in_362, d_out_363, qn_in_363, d_out_364, qn_in_364, d_out_365, qn_in_365, d_out_366, qn_in_366, d_out_367, qn_in_367, d_out_368, q_in_368, d_out_369, q_in_369, d_out_370, q_in_370, d_out_371, q_in_371, d_out_372, q_in_372, d_out_373, qn_in_373, d_out_374, qn_in_374, d_out_375, q_in_375, d_out_376, qn_in_376, d_out_377, qn_in_377, d_out_378, qn_in_378, d_out_379, q_in_379, d_out_380, q_in_380, d_out_381, q_in_381, d_out_382, qn_in_382, d_out_383, qn_in_383, d_out_384, qn_in_384, d_out_385, q_in_385, d_out_386, q_in_386, d_out_387, q_in_387, d_out_388, q_in_388, d_out_389, q_in_389, d_out_390, q_in_390, d_out_391, qn_in_391, d_out_392, qn_in_392, d_out_393, qn_in_393, d_out_394, qn_in_394, d_out_395, qn_in_395, d_out_396, qn_in_396, d_out_397, q_in_397, d_out_398, q_in_398, d_out_399, q_in_399, d_out_400, q_in_400, d_out_401, q_in_401, d_out_402, q_in_402, d_out_403, qn_in_403, d_out_404, qn_in_404, d_out_405, qn_in_405, d_out_406, qn_in_406, d_out_407, qn_in_407, d_out_408, q_in_408, d_out_409, q_in_409, d_out_410, q_in_410, d_out_411, qn_in_411, d_out_412, qn_in_412, d_out_413, qn_in_413, d_out_414, q_in_414, d_out_415, q_in_415, d_out_416, q_in_416, d_out_417, q_in_417, d_out_418, q_in_418, d_out_419, q_in_419, d_out_420, q_in_420, d_out_421, q_in_421, d_out_422, q_in_422, d_out_423, q_in_423, d_out_424, q_in_424, d_out_425, q_in_425, d_out_426, qn_in_426, d_out_427, qn_in_427, d_out_428, qn_in_428, d_out_429, qn_in_429, d_out_430, qn_in_430, d_out_431, qn_in_431, d_out_432, q_in_432, d_out_433, q_in_433, d_out_434, q_in_434, d_out_435, q_in_435, d_out_436, qn_in_436, d_out_437, qn_in_437, d_out_438, qn_in_438, d_out_439, qn_in_439, d_out_440, q_in_440, d_out_441, q_in_441, d_out_442, q_in_442, d_out_443, qn_in_443, d_out_444, qn_in_444, d_out_445, qn_in_445, d_out_446, qn_in_446, d_out_447, q_in_447, d_out_448, q_in_448, d_out_449, q_in_449, d_out_450, q_in_450, d_out_451, q_in_451, d_out_452, q_in_452, d_out_453, q_in_453, d_out_454, qn_in_454, d_out_455, qn_in_455, d_out_456, qn_in_456, d_out_457, qn_in_457, d_out_458, qn_in_458, d_out_459, qn_in_459, d_out_460, q_in_460, d_out_461, q_in_461, d_out_462, q_in_462, d_out_463, q_in_463, d_out_464, q_in_464, d_out_465, q_in_465, d_out_466, q_in_466, d_out_467, q_in_467, d_out_468, q_in_468, d_out_469, qn_in_469, d_out_470, qn_in_470, d_out_471, qn_in_471, d_out_472, q_in_472, d_out_473, q_in_473, d_out_474, q_in_474, d_out_475, q_in_475, d_out_476, q_in_476, d_out_477, q_in_477, d_out_478, q_in_478, d_out_479, q_in_479, d_out_480, q_in_480, d_out_481, q_in_481, d_out_482, q_in_482, d_out_483, q_in_483, d_out_484, q_in_484, d_out_485, q_in_485, d_out_486, q_in_486, d_out_487, q_in_487, d_out_488, q_in_488, d_out_489, q_in_489, d_out_490, q_in_490, d_out_491, q_in_491, d_out_492, q_in_492, d_out_493, q_in_493, d_out_494, q_in_494, d_out_495, q_in_495, d_out_496, q_in_496, d_out_497, q_in_497, d_out_498, q_in_498, d_out_499, q_in_499, d_out_500, q_in_500, d_out_501, q_in_501, d_out_502, q_in_502, d_out_503, q_in_503, d_out_504, qn_in_504, d_out_505, q_in_505, d_out_506, q_in_506, d_out_507, qn_in_507, d_out_508, q_in_508, d_out_509, qn_in_509, d_out_510, qn_in_510, d_out_511, qn_in_511, d_out_512, q_in_512, d_out_513, q_in_513, d_out_514, q_in_514, d_out_515, q_in_515, d_out_516, q_in_516, d_out_517, q_in_517, d_out_518, qn_in_518, d_out_519, qn_in_519, d_out_520, qn_in_520, d_out_521, qn_in_521, d_out_522, qn_in_522, d_out_523, qn_in_523, d_out_524, qn_in_524, d_out_525, qn_in_525, d_out_526, qn_in_526, d_out_527, qn_in_527, d_out_528, qn_in_528, d_out_529, qn_in_529, d_out_530, qn_in_530, d_out_531, qn_in_531, d_out_532, qn_in_532, d_out_533, qn_in_533, d_out_534, qn_in_534, d_out_535, qn_in_535, d_out_536, qn_in_536, d_out_537, qn_in_537, d_out_538, qn_in_538, d_out_539, qn_in_539, d_out_540, q_in_540, d_out_541, qn_in_541, d_out_542, qn_in_542, d_out_543, qn_in_543, d_out_544, qn_in_544, d_out_545, qn_in_545, d_out_546, qn_in_546, d_out_547, q_in_547, d_out_548, q_in_548, d_out_549, q_in_549, d_out_550, qn_in_550, d_out_551, qn_in_551, d_out_552, qn_in_552, d_out_553, qn_in_553, d_out_554, qn_in_554, d_out_555, qn_in_555, d_out_556, qn_in_556, d_out_557, qn_in_557, d_out_558, q_in_558, d_out_559, qn_in_559, d_out_560, q_in_560, d_out_561, q_in_561, d_out_562, q_in_562, d_out_563, qn_in_563, d_out_564, q_in_564, d_out_565, q_in_565, d_out_566, q_in_566, d_out_567, q_in_567, d_out_568, q_in_568, d_out_569, q_in_569, d_out_570, q_in_570, d_out_571, q_in_571, d_out_572, q_in_572, d_out_573, q_in_573, d_out_574, q_in_574, d_out_575, q_in_575, d_out_576, q_in_576, d_out_577, q_in_577, d_out_578, q_in_578, d_out_579, q_in_579, d_out_580, q_in_580, d_out_581, q_in_581, d_out_582, q_in_582, d_out_583, q_in_583, d_out_584, q_in_584, d_out_585, qn_in_585, d_out_586, qn_in_586, d_out_587, qn_in_587, d_out_588, q_in_588, d_out_589, q_in_589, d_out_590, q_in_590, d_out_591, q_in_591, d_out_592, q_in_592, d_out_593, q_in_593, d_out_594, q_in_594, d_out_595, q_in_595, d_out_596, q_in_596, d_out_597, q_in_597, d_out_598, q_in_598, d_out_599, q_in_599, d_out_600, q_in_600, d_out_601, q_in_601, d_out_602, q_in_602, d_out_603, q_in_603, d_out_604, q_in_604, d_out_605, q_in_605, d_out_606, q_in_606, d_out_607, q_in_607, d_out_608, q_in_608, d_out_609, q_in_609, d_out_610, q_in_610, d_out_611, q_in_611, d_out_612, q_in_612, d_out_613, q_in_613, d_out_614, q_in_614, d_out_615, q_in_615, d_out_616, q_in_616, d_out_617, q_in_617, d_out_618, q_in_618, d_out_619, q_in_619, d_out_620, q_in_620, d_out_621, q_in_621, d_out_622, q_in_622, d_out_623, q_in_623, d_out_624, q_in_624, d_out_625, q_in_625, d_out_626, q_in_626, d_out_627, q_in_627, d_out_628, q_in_628, d_out_629, q_in_629, d_out_630, q_in_630, d_out_631, q_in_631, d_out_632, q_in_632, d_out_633, q_in_633, d_out_634, q_in_634, d_out_635, q_in_635, d_out_636, q_in_636, d_out_637, q_in_637, d_out_638, q_in_638, d_out_639, q_in_639, d_out_640, q_in_640, d_out_641, q_in_641, d_out_642, q_in_642, d_out_643, q_in_643, d_out_644, q_in_644, d_out_645, q_in_645, d_out_646, qn_in_646, d_out_647, q_in_647, d_out_648, q_in_648, d_out_649, q_in_649, d_out_650, q_in_650, d_out_651, q_in_651, d_out_652, q_in_652, d_out_653, q_in_653, d_out_654, q_in_654, d_out_655, q_in_655, d_out_656, q_in_656, d_out_657, q_in_657, d_out_658, q_in_658, d_out_659, q_in_659, d_out_660, q_in_660, d_out_661, q_in_661, d_out_662, q_in_662, d_out_663, q_in_663, d_out_664, q_in_664, d_out_665, q_in_665, d_out_666, q_in_666, d_out_667, q_in_667, d_out_668, q_in_668, d_out_669, q_in_669, d_out_670, q_in_670, d_out_671, q_in_671, d_out_672, q_in_672, d_out_673, q_in_673, d_out_674, q_in_674, d_out_675, q_in_675, d_out_676, q_in_676, d_out_677, q_in_677, d_out_678, q_in_678, d_out_679, q_in_679, d_out_680, q_in_680, d_out_681, q_in_681, d_out_682, q_in_682, d_out_683, q_in_683, d_out_684, q_in_684, d_out_685, q_in_685, d_out_686, q_in_686, d_out_687, q_in_687, d_out_688, q_in_688, d_out_689, q_in_689, d_out_690, q_in_690, d_out_691, q_in_691, d_out_692, q_in_692, d_out_693, q_in_693, d_out_694, q_in_694, d_out_695, q_in_695, d_out_696, q_in_696, d_out_697, q_in_697, d_out_698, q_in_698, d_out_699, q_in_699, d_out_700, q_in_700, d_out_701, q_in_701, d_out_702, q_in_702, d_out_703, q_in_703, d_out_704, q_in_704, d_out_705, q_in_705, d_out_706, q_in_706, d_out_707, q_in_707, d_out_708, q_in_708, d_out_709, q_in_709, d_out_710, q_in_710, d_out_711, q_in_711, d_out_712, q_in_712, d_out_713, q_in_713, d_out_714, q_in_714, d_out_715, q_in_715, d_out_716, q_in_716, d_out_717, q_in_717, d_out_718, q_in_718, d_out_719, q_in_719, d_out_720, q_in_720, d_out_721, q_in_721, d_out_722, q_in_722, d_out_723, q_in_723, d_out_724, q_in_724, d_out_725, q_in_725, d_out_726, q_in_726, d_out_727, q_in_727, d_out_728, q_in_728, d_out_729, q_in_729, d_out_730, q_in_730, d_out_731, q_in_731, d_out_732, q_in_732, d_out_733, q_in_733, d_out_734, qn_in_734, d_out_735, q_in_735, d_out_736, q_in_736, d_out_737, qn_in_737, d_out_738, q_in_738, d_out_739, q_in_739, d_out_740, q_in_740, d_out_741, q_in_741, d_out_742, q_in_742, d_out_743, q_in_743, d_out_744, q_in_744, d_out_745, q_in_745, d_out_746, q_in_746, d_out_747, qn_in_747, d_out_748, q_in_748, d_out_749, q_in_749, d_out_750, q_in_750, d_out_751, q_in_751, d_out_752, q_in_752, d_out_753, q_in_753, d_out_754, q_in_754, d_out_755, q_in_755, d_out_756, q_in_756, d_out_757, q_in_757, d_out_758, q_in_758, d_out_759, q_in_759, d_out_760, q_in_760, d_out_761, q_in_761, d_out_762, q_in_762, d_out_763, q_in_763, d_out_764, q_in_764, d_out_765, q_in_765, d_out_766, q_in_766, d_out_767, q_in_767, d_out_768, q_in_768, d_out_769, q_in_769, d_out_770, q_in_770, d_out_771, q_in_771, d_out_772, q_in_772, d_out_773, q_in_773, d_out_774, q_in_774, d_out_775, q_in_775, d_out_776, q_in_776, d_out_777, q_in_777, d_out_778, q_in_778, d_out_779, q_in_779, d_out_780, q_in_780, d_out_781, q_in_781, d_out_782, q_in_782, d_out_783, q_in_783, d_out_784, q_in_784, d_out_785, q_in_785, d_out_786, q_in_786, d_out_787, q_in_787, d_out_788, q_in_788, d_out_789, q_in_789, d_out_790, q_in_790, d_out_791, q_in_791, d_out_792, q_in_792, d_out_793, q_in_793, d_out_794, q_in_794, d_out_795, q_in_795, d_out_796, q_in_796, d_out_797, q_in_797, d_out_798, q_in_798, d_out_799, q_in_799, d_out_800, q_in_800, d_out_801, q_in_801, d_out_802, q_in_802, d_out_803, q_in_803, d_out_804, q_in_804, d_out_805, q_in_805, d_out_806, q_in_806, d_out_807, q_in_807, d_out_808, q_in_808, d_out_809, q_in_809, d_out_810, q_in_810, d_out_811, q_in_811, d_out_812, q_in_812, d_out_813, q_in_813, d_out_814, q_in_814, d_out_815, q_in_815, d_out_816, q_in_816, d_out_817, q_in_817, d_out_818, q_in_818, d_out_819, q_in_819, d_out_820, q_in_820, d_out_821, q_in_821, d_out_822, q_in_822, d_out_823, q_in_823, d_out_824, q_in_824, d_out_825, q_in_825, d_out_826, q_in_826, d_out_827, q_in_827, d_out_828, q_in_828, d_out_829, q_in_829, d_out_830, q_in_830, d_out_831, q_in_831, d_out_832, q_in_832, d_out_833, q_in_833, d_out_834, q_in_834, d_out_835, q_in_835, d_out_836, q_in_836, d_out_837, q_in_837, d_out_838, q_in_838, d_out_839, q_in_839, d_out_840, q_in_840, d_out_841, q_in_841, d_out_842, q_in_842, d_out_843, q_in_843, d_out_844, q_in_844, d_out_845, q_in_845, d_out_846, q_in_846, d_out_847, q_in_847, d_out_848, q_in_848, d_out_849, q_in_849, d_out_850, q_in_850, d_out_851, q_in_851, d_out_852, q_in_852, d_out_853, q_in_853, d_out_854, q_in_854, d_out_855, q_in_855, d_out_856, q_in_856, d_out_857, q_in_857, d_out_858, q_in_858, d_out_859, q_in_859, d_out_860, q_in_860, d_out_861, q_in_861, d_out_862, q_in_862, d_out_863, q_in_863, d_out_864, q_in_864, d_out_865, q_in_865, d_out_866, q_in_866, d_out_867, q_in_867, d_out_868, q_in_868, d_out_869, q_in_869, d_out_870, q_in_870, d_out_871, q_in_871, d_out_872, q_in_872, d_out_873, q_in_873, d_out_874, q_in_874, d_out_875, q_in_875, d_out_876, q_in_876, d_out_877, q_in_877, d_out_878, q_in_878, d_out_879, q_in_879, d_out_880, q_in_880, d_out_881, q_in_881, d_out_882, q_in_882, d_out_883, q_in_883, d_out_884, q_in_884, d_out_885, q_in_885, d_out_886, q_in_886, d_out_887, q_in_887, d_out_888, q_in_888, d_out_889, q_in_889, d_out_890, q_in_890, d_out_891, q_in_891, d_out_892, q_in_892, d_out_893, q_in_893, d_out_894, q_in_894, d_out_895, q_in_895, d_out_896, q_in_896, d_out_897, q_in_897, d_out_898, q_in_898, d_out_899, q_in_899, d_out_900, q_in_900, d_out_901, q_in_901, d_out_902, q_in_902, d_out_903, q_in_903, d_out_904, q_in_904, d_out_905, q_in_905, d_out_906, q_in_906, d_out_907, q_in_907, d_out_908, q_in_908, d_out_909, q_in_909, d_out_910, q_in_910, d_out_911, q_in_911, d_out_912, q_in_912, d_out_913, q_in_913, d_out_914, q_in_914, d_out_915, q_in_915, d_out_916, q_in_916, d_out_917, q_in_917, d_out_918, q_in_918, d_out_919, q_in_919, d_out_920, q_in_920, d_out_921, q_in_921, d_out_922, q_in_922, d_out_923, q_in_923, d_out_924, q_in_924, d_out_925, q_in_925, d_out_926, q_in_926, d_out_927, q_in_927, d_out_928, q_in_928, d_out_929, q_in_929, d_out_930, q_in_930, d_out_931, q_in_931, d_out_932, q_in_932, d_out_933, q_in_933, d_out_934, q_in_934, d_out_935, q_in_935, d_out_936, q_in_936, d_out_937, q_in_937, d_out_938, q_in_938, d_out_939, q_in_939, d_out_940, q_in_940, d_out_941, q_in_941, d_out_942, q_in_942, d_out_943, q_in_943, d_out_944, q_in_944, d_out_945, q_in_945, d_out_946, q_in_946, d_out_947, q_in_947, d_out_948, q_in_948, d_out_949, q_in_949, d_out_950, q_in_950, d_out_951, q_in_951, d_out_952, q_in_952, d_out_953, q_in_953, d_out_954, q_in_954, d_out_955, q_in_955, d_out_956, q_in_956, d_out_957, qn_in_957, d_out_958, q_in_958, d_out_959, q_in_959, d_out_960, q_in_960, d_out_961, q_in_961, d_out_962, q_in_962, d_out_963, q_in_963, d_out_964, q_in_964, d_out_965, q_in_965, d_out_966, q_in_966, d_out_967, q_in_967, d_out_968, q_in_968, d_out_969, q_in_969, d_out_970, q_in_970, d_out_971, q_in_971, d_out_972, q_in_972, d_out_973, q_in_973, d_out_974, q_in_974, d_out_975, q_in_975, d_out_976, q_in_976, d_out_977, q_in_977, d_out_978, q_in_978, d_out_979, q_in_979, d_out_980, q_in_980, d_out_981, q_in_981, d_out_982, q_in_982, d_out_983, q_in_983, d_out_984, q_in_984, d_out_985, q_in_985, d_out_986, q_in_986, d_out_987, q_in_987, d_out_988, q_in_988, d_out_989, q_in_989, d_out_990, q_in_990, d_out_991, q_in_991, d_out_992, q_in_992, d_out_993, q_in_993, d_out_994, q_in_994, d_out_995, q_in_995, d_out_996, q_in_996, d_out_997, q_in_997, d_out_998, q_in_998, d_out_999, q_in_999, d_out_1000, q_in_1000, d_out_1001, q_in_1001, d_out_1002, q_in_1002, d_out_1003, q_in_1003, d_out_1004, q_in_1004, d_out_1005, q_in_1005, d_out_1006, q_in_1006, d_out_1007, q_in_1007, d_out_1008, q_in_1008, d_out_1009, q_in_1009, d_out_1010, q_in_1010, d_out_1011, q_in_1011, d_out_1012, q_in_1012, d_out_1013, q_in_1013, d_out_1014, q_in_1014, d_out_1015, q_in_1015, d_out_1016, q_in_1016, d_out_1017, q_in_1017, d_out_1018, q_in_1018, d_out_1019, q_in_1019, d_out_1020, q_in_1020, d_out_1021, q_in_1021, d_out_1022, q_in_1022, d_out_1023, q_in_1023, d_out_1024, q_in_1024, d_out_1025, q_in_1025, d_out_1026, q_in_1026, d_out_1027, q_in_1027, d_out_1028, q_in_1028, d_out_1029, q_in_1029, d_out_1030, q_in_1030, d_out_1031, q_in_1031, d_out_1032, q_in_1032, d_out_1033, q_in_1033, d_out_1034, q_in_1034, d_out_1035, q_in_1035, d_out_1036, q_in_1036, d_out_1037, q_in_1037, d_out_1038, q_in_1038, d_out_1039, q_in_1039, d_out_1040, q_in_1040, d_out_1041, q_in_1041, d_out_1042, q_in_1042, d_out_1043, q_in_1043, d_out_1044, q_in_1044, d_out_1045, q_in_1045, d_out_1046, q_in_1046, d_out_1047, q_in_1047, d_out_1048, q_in_1048, d_out_1049, q_in_1049, d_out_1050, q_in_1050, d_out_1051, q_in_1051, d_out_1052, q_in_1052, d_out_1053, q_in_1053, d_out_1054, q_in_1054, d_out_1055, q_in_1055, d_out_1056, q_in_1056, d_out_1057, q_in_1057, d_out_1058, q_in_1058, d_out_1059, q_in_1059, d_out_1060, q_in_1060, d_out_1061, q_in_1061, d_out_1062, q_in_1062, d_out_1063, q_in_1063, d_out_1064, q_in_1064, d_out_1065, q_in_1065, d_out_1066, q_in_1066, d_out_1067, q_in_1067, d_out_1068, q_in_1068, d_out_1069, q_in_1069, d_out_1070, q_in_1070, d_out_1071, q_in_1071, d_out_1072, q_in_1072, d_out_1073, q_in_1073, d_out_1074, q_in_1074, d_out_1075, q_in_1075, d_out_1076, q_in_1076, d_out_1077, q_in_1077, d_out_1078, q_in_1078, d_out_1079, q_in_1079, d_out_1080, q_in_1080, d_out_1081, q_in_1081, d_out_1082, q_in_1082, d_out_1083, q_in_1083, d_out_1084, q_in_1084, d_out_1085, q_in_1085, d_out_1086, q_in_1086, d_out_1087, q_in_1087, d_out_1088, q_in_1088, d_out_1089, q_in_1089, d_out_1090, q_in_1090, d_out_1091, q_in_1091, d_out_1092, q_in_1092, d_out_1093, q_in_1093, d_out_1094, q_in_1094, d_out_1095, q_in_1095, d_out_1096, q_in_1096, d_out_1097, q_in_1097, d_out_1098, q_in_1098, d_out_1099, q_in_1099, d_out_1100, q_in_1100, d_out_1101, q_in_1101, d_out_1102, q_in_1102, d_out_1103, q_in_1103, d_out_1104, q_in_1104, d_out_1105, q_in_1105, d_out_1106, q_in_1106, d_out_1107, q_in_1107, d_out_1108, q_in_1108, d_out_1109, q_in_1109, d_out_1110, q_in_1110, d_out_1111, q_in_1111, d_out_1112, q_in_1112, d_out_1113, q_in_1113, d_out_1114, q_in_1114, d_out_1115, q_in_1115, d_out_1116, q_in_1116, d_out_1117, q_in_1117, d_out_1118, q_in_1118, d_out_1119, q_in_1119, d_out_1120, q_in_1120, d_out_1121, q_in_1121, d_out_1122, q_in_1122, d_out_1123, q_in_1123, d_out_1124, q_in_1124, d_out_1125, q_in_1125, d_out_1126, q_in_1126, d_out_1127, q_in_1127, d_out_1128, q_in_1128, d_out_1129, q_in_1129, d_out_1130, q_in_1130, d_out_1131, q_in_1131, d_out_1132, q_in_1132, d_out_1133, q_in_1133, d_out_1134, q_in_1134, d_out_1135, q_in_1135, d_out_1136, q_in_1136, d_out_1137, q_in_1137, d_out_1138, q_in_1138, d_out_1139, q_in_1139, d_out_1140, q_in_1140, d_out_1141, q_in_1141, d_out_1142, q_in_1142, d_out_1143, q_in_1143, d_out_1144, q_in_1144, d_out_1145, q_in_1145, d_out_1146, q_in_1146, d_out_1147, q_in_1147, d_out_1148, q_in_1148, d_out_1149, q_in_1149, d_out_1150, q_in_1150, d_out_1151, q_in_1151, d_out_1152, q_in_1152, d_out_1153, q_in_1153, d_out_1154, q_in_1154, d_out_1155, q_in_1155, d_out_1156, q_in_1156, d_out_1157, q_in_1157, d_out_1158, q_in_1158, d_out_1159, q_in_1159, d_out_1160, q_in_1160, d_out_1161, q_in_1161, d_out_1162, q_in_1162, d_out_1163, q_in_1163, d_out_1164, q_in_1164, d_out_1165, q_in_1165, d_out_1166, q_in_1166, d_out_1167, q_in_1167, d_out_1168, q_in_1168, d_out_1169, q_in_1169, d_out_1170, q_in_1170, d_out_1171, q_in_1171, d_out_1172, q_in_1172, d_out_1173, q_in_1173, d_out_1174, q_in_1174, d_out_1175, q_in_1175, d_out_1176, q_in_1176, d_out_1177, q_in_1177, d_out_1178, q_in_1178, d_out_1179, q_in_1179, d_out_1180, q_in_1180, d_out_1181, q_in_1181, d_out_1182, q_in_1182, d_out_1183, q_in_1183, d_out_1184, q_in_1184, d_out_1185, q_in_1185, d_out_1186, q_in_1186, d_out_1187, q_in_1187, d_out_1188, q_in_1188, d_out_1189, q_in_1189, d_out_1190, q_in_1190, d_out_1191, q_in_1191, d_out_1192, q_in_1192, d_out_1193, q_in_1193, d_out_1194, q_in_1194, d_out_1195, q_in_1195, d_out_1196, q_in_1196, d_out_1197, q_in_1197, d_out_1198, q_in_1198, d_out_1199, q_in_1199, d_out_1200, q_in_1200, d_out_1201, q_in_1201, d_out_1202, q_in_1202, d_out_1203, q_in_1203, d_out_1204, q_in_1204, d_out_1205, q_in_1205, d_out_1206, q_in_1206, d_out_1207, q_in_1207, d_out_1208, q_in_1208, d_out_1209, q_in_1209, d_out_1210, q_in_1210, d_out_1211, q_in_1211, d_out_1212, q_in_1212, d_out_1213, q_in_1213, d_out_1214, q_in_1214, d_out_1215, q_in_1215, d_out_1216, q_in_1216, d_out_1217, q_in_1217, d_out_1218, q_in_1218, d_out_1219, q_in_1219, d_out_1220, q_in_1220, d_out_1221, q_in_1221, d_out_1222, q_in_1222, d_out_1223, q_in_1223, d_out_1224, q_in_1224, d_out_1225, q_in_1225, d_out_1226, q_in_1226, d_out_1227, q_in_1227, d_out_1228, q_in_1228, d_out_1229, q_in_1229, d_out_1230, q_in_1230, d_out_1231, q_in_1231, d_out_1232, q_in_1232, d_out_1233, q_in_1233, d_out_1234, q_in_1234, d_out_1235, q_in_1235, d_out_1236, q_in_1236, d_out_1237, q_in_1237, d_out_1238, q_in_1238, d_out_1239, q_in_1239, d_out_1240, q_in_1240, d_out_1241, q_in_1241, d_out_1242, q_in_1242, d_out_1243, q_in_1243, d_out_1244, q_in_1244, d_out_1245, q_in_1245, d_out_1246, q_in_1246, d_out_1247, q_in_1247, d_out_1248, q_in_1248, d_out_1249, q_in_1249, d_out_1250, q_in_1250, d_out_1251, q_in_1251, d_out_1252, q_in_1252, d_out_1253, q_in_1253, d_out_1254, q_in_1254, d_out_1255, q_in_1255, d_out_1256, q_in_1256, d_out_1257, q_in_1257, d_out_1258, q_in_1258, d_out_1259, q_in_1259, d_out_1260, q_in_1260, d_out_1261, q_in_1261, d_out_1262, q_in_1262, d_out_1263, q_in_1263, d_out_1264, q_in_1264, d_out_1265, q_in_1265, d_out_1266, q_in_1266, d_out_1267, q_in_1267, d_out_1268, q_in_1268, d_out_1269, q_in_1269, d_out_1270, q_in_1270, d_out_1271, q_in_1271, d_out_1272, q_in_1272, d_out_1273, q_in_1273, d_out_1274, q_in_1274, d_out_1275, q_in_1275, d_out_1276, q_in_1276, d_out_1277, q_in_1277, d_out_1278, q_in_1278, d_out_1279, q_in_1279, d_out_1280, q_in_1280, d_out_1281, q_in_1281, d_out_1282, q_in_1282, d_out_1283, q_in_1283, d_out_1284, q_in_1284, d_out_1285, q_in_1285, d_out_1286, q_in_1286, d_out_1287, q_in_1287, d_out_1288, q_in_1288, d_out_1289, q_in_1289, d_out_1290, q_in_1290, d_out_1291, q_in_1291, d_out_1292, q_in_1292, d_out_1293, q_in_1293, d_out_1294, q_in_1294, d_out_1295, q_in_1295, d_out_1296, q_in_1296, d_out_1297, q_in_1297, d_out_1298, q_in_1298, d_out_1299, q_in_1299, d_out_1300, q_in_1300, d_out_1301, q_in_1301, d_out_1302, q_in_1302, d_out_1303, q_in_1303, d_out_1304, q_in_1304, d_out_1305, q_in_1305, d_out_1306, q_in_1306, d_out_1307, q_in_1307, d_out_1308, q_in_1308, d_out_1309, q_in_1309, d_out_1310, q_in_1310, d_out_1311, q_in_1311, d_out_1312, q_in_1312, d_out_1313, q_in_1313, d_out_1314, q_in_1314, d_out_1315, q_in_1315, d_out_1316, q_in_1316, d_out_1317, q_in_1317, d_out_1318, q_in_1318, d_out_1319, q_in_1319, d_out_1320, q_in_1320, d_out_1321, q_in_1321, d_out_1322, q_in_1322, d_out_1323, q_in_1323, d_out_1324, q_in_1324, d_out_1325, q_in_1325, d_out_1326, q_in_1326, d_out_1327, q_in_1327, d_out_1328, q_in_1328, d_out_1329, q_in_1329, d_out_1330, q_in_1330, d_out_1331, q_in_1331, d_out_1332, q_in_1332, d_out_1333, q_in_1333, d_out_1334, q_in_1334, d_out_1335, q_in_1335, d_out_1336, q_in_1336, d_out_1337, q_in_1337, d_out_1338, q_in_1338, d_out_1339, q_in_1339, d_out_1340, q_in_1340, d_out_1341, q_in_1341, d_out_1342, q_in_1342, d_out_1343, q_in_1343, d_out_1344, q_in_1344, d_out_1345, q_in_1345, d_out_1346, q_in_1346, d_out_1347, q_in_1347, d_out_1348, q_in_1348, d_out_1349, q_in_1349, d_out_1350, q_in_1350, d_out_1351, q_in_1351, d_out_1352, q_in_1352, d_out_1353, q_in_1353, d_out_1354, q_in_1354, d_out_1355, q_in_1355, d_out_1356, q_in_1356, d_out_1357, q_in_1357, d_out_1358, q_in_1358, d_out_1359, q_in_1359, d_out_1360, q_in_1360, d_out_1361, q_in_1361, d_out_1362, q_in_1362, d_out_1363, q_in_1363, d_out_1364, q_in_1364, d_out_1365, q_in_1365, d_out_1366, q_in_1366, d_out_1367, q_in_1367, d_out_1368, q_in_1368, d_out_1369, q_in_1369, d_out_1370, q_in_1370, d_out_1371, q_in_1371, d_out_1372, q_in_1372, d_out_1373, q_in_1373, d_out_1374, q_in_1374, d_out_1375, q_in_1375, d_out_1376, q_in_1376, d_out_1377, q_in_1377, d_out_1378, q_in_1378, d_out_1379, q_in_1379, d_out_1380, q_in_1380, d_out_1381, q_in_1381, d_out_1382, q_in_1382, d_out_1383, q_in_1383, d_out_1384, q_in_1384, d_out_1385, q_in_1385, d_out_1386, q_in_1386, d_out_1387, q_in_1387, d_out_1388, q_in_1388, d_out_1389, q_in_1389, d_out_1390, q_in_1390, d_out_1391, q_in_1391, d_out_1392, q_in_1392, d_out_1393, q_in_1393, d_out_1394, q_in_1394, d_out_1395, q_in_1395, d_out_1396, q_in_1396, d_out_1397, q_in_1397, d_out_1398, q_in_1398, d_out_1399, q_in_1399, d_out_1400, q_in_1400, d_out_1401, q_in_1401, d_out_1402, q_in_1402, d_out_1403, q_in_1403, d_out_1404, q_in_1404, d_out_1405, q_in_1405, d_out_1406, q_in_1406, d_out_1407, q_in_1407, d_out_1408, q_in_1408, d_out_1409, q_in_1409, d_out_1410, q_in_1410, d_out_1411, q_in_1411, d_out_1412, q_in_1412, d_out_1413, q_in_1413, d_out_1414, q_in_1414, d_out_1415, q_in_1415, d_out_1416, q_in_1416, d_out_1417, q_in_1417, d_out_1418, q_in_1418, d_out_1419, q_in_1419, d_out_1420, q_in_1420, d_out_1421, q_in_1421, d_out_1422, q_in_1422, d_out_1423, q_in_1423, d_out_1424, q_in_1424, d_out_1425, q_in_1425, d_out_1426, q_in_1426, d_out_1427, q_in_1427, d_out_1428, q_in_1428, d_out_1429, q_in_1429, d_out_1430, q_in_1430, d_out_1431, q_in_1431, d_out_1432, q_in_1432, d_out_1433, q_in_1433, d_out_1434, q_in_1434, d_out_1435, q_in_1435, d_out_1436, q_in_1436, d_out_1437, q_in_1437, d_out_1438, q_in_1438, d_out_1439, q_in_1439, d_out_1440, q_in_1440, d_out_1441, q_in_1441, d_out_1442, q_in_1442, d_out_1443, q_in_1443, d_out_1444, q_in_1444, d_out_1445, q_in_1445, d_out_1446, q_in_1446, d_out_1447, q_in_1447, d_out_1448, q_in_1448, d_out_1449, q_in_1449, d_out_1450, q_in_1450, d_out_1451, q_in_1451, d_out_1452, q_in_1452, d_out_1453, q_in_1453, d_out_1454, q_in_1454, d_out_1455, q_in_1455, d_out_1456, q_in_1456, d_out_1457, q_in_1457, d_out_1458, q_in_1458, d_out_1459, q_in_1459, d_out_1460, q_in_1460, d_out_1461, q_in_1461, d_out_1462, q_in_1462, d_out_1463, q_in_1463, d_out_1464, q_in_1464, d_out_1465, q_in_1465, d_out_1466, q_in_1466, d_out_1467, q_in_1467, d_out_1468, q_in_1468, d_out_1469, q_in_1469, d_out_1470, q_in_1470, d_out_1471, q_in_1471, d_out_1472, q_in_1472, d_out_1473, q_in_1473, d_out_1474, q_in_1474, d_out_1475, q_in_1475, d_out_1476, q_in_1476, d_out_1477, q_in_1477, d_out_1478, q_in_1478, d_out_1479, q_in_1479, d_out_1480, q_in_1480, d_out_1481, q_in_1481, d_out_1482, q_in_1482, d_out_1483, q_in_1483, d_out_1484, q_in_1484, d_out_1485, q_in_1485, d_out_1486, q_in_1486, d_out_1487, q_in_1487, d_out_1488, q_in_1488, d_out_1489, q_in_1489, d_out_1490, q_in_1490, d_out_1491, q_in_1491, d_out_1492, q_in_1492, d_out_1493, q_in_1493, d_out_1494, q_in_1494, d_out_1495, q_in_1495, d_out_1496, q_in_1496, d_out_1497, q_in_1497, d_out_1498, q_in_1498, d_out_1499, q_in_1499, d_out_1500, q_in_1500, d_out_1501, q_in_1501, d_out_1502, q_in_1502, d_out_1503, q_in_1503, d_out_1504, q_in_1504, d_out_1505, q_in_1505, d_out_1506, q_in_1506, d_out_1507, q_in_1507, d_out_1508, q_in_1508, d_out_1509, q_in_1509, d_out_1510, q_in_1510, d_out_1511, q_in_1511, d_out_1512, q_in_1512, d_out_1513, q_in_1513, d_out_1514, q_in_1514, d_out_1515, q_in_1515, d_out_1516, q_in_1516, d_out_1517, q_in_1517, d_out_1518, q_in_1518, d_out_1519, q_in_1519, d_out_1520, q_in_1520, d_out_1521, q_in_1521, d_out_1522, q_in_1522, d_out_1523, q_in_1523, d_out_1524, q_in_1524, d_out_1525, q_in_1525, d_out_1526, q_in_1526, d_out_1527, q_in_1527, d_out_1528, q_in_1528, d_out_1529, q_in_1529, d_out_1530, q_in_1530, d_out_1531, q_in_1531, d_out_1532, q_in_1532, d_out_1533, q_in_1533, d_out_1534, q_in_1534, d_out_1535, q_in_1535, d_out_1536, q_in_1536, d_out_1537, q_in_1537, d_out_1538, q_in_1538, d_out_1539, q_in_1539, d_out_1540, q_in_1540, d_out_1541, q_in_1541, d_out_1542, q_in_1542, d_out_1543, q_in_1543, d_out_1544, q_in_1544, d_out_1545, q_in_1545, d_out_1546, q_in_1546, d_out_1547, q_in_1547, d_out_1548, q_in_1548, d_out_1549, q_in_1549, d_out_1550, q_in_1550, d_out_1551, q_in_1551, d_out_1552, q_in_1552, d_out_1553, q_in_1553, d_out_1554, q_in_1554, d_out_1555, q_in_1555, d_out_1556, q_in_1556, d_out_1557, q_in_1557, d_out_1558, q_in_1558, d_out_1559, q_in_1559, d_out_1560, q_in_1560, d_out_1561, q_in_1561, d_out_1562, q_in_1562, d_out_1563, q_in_1563, d_out_1564, q_in_1564, d_out_1565, q_in_1565, d_out_1566, q_in_1566, d_out_1567, q_in_1567, d_out_1568, q_in_1568, d_out_1569, q_in_1569, d_out_1570, q_in_1570, d_out_1571, q_in_1571, d_out_1572, q_in_1572, d_out_1573, q_in_1573, d_out_1574, q_in_1574, d_out_1575, q_in_1575, d_out_1576, q_in_1576, d_out_1577, q_in_1577, d_out_1578, q_in_1578, d_out_1579, q_in_1579, d_out_1580, q_in_1580, d_out_1581, qn_in_1581, d_out_1582, qn_in_1582, d_out_1583, q_in_1583, d_out_1584, q_in_1584, d_out_1585, q_in_1585, d_out_1586, q_in_1586, d_out_1587, q_in_1587, d_out_1588, q_in_1588, d_out_1589, q_in_1589, d_out_1590, q_in_1590, d_out_1591, q_in_1591, d_out_1592, q_in_1592, d_out_1593, q_in_1593, d_out_1594, q_in_1594, d_out_1595, q_in_1595, d_out_1596, q_in_1596, d_out_1597, qn_in_1597, d_out_1598, q_in_1598, d_out_1599, q_in_1599, d_out_1600, q_in_1600, d_out_1601, q_in_1601, d_out_1602, q_in_1602, d_out_1603, q_in_1603, d_out_1604, q_in_1604, d_out_1605, q_in_1605, d_out_1606, q_in_1606, d_out_1607, q_in_1607, d_out_1608, q_in_1608, d_out_1609, q_in_1609, d_out_1610, q_in_1610, d_out_1611, q_in_1611, d_out_1612, q_in_1612, d_out_1613, q_in_1613, d_out_1614, q_in_1614, d_out_1615, q_in_1615, d_out_1616, q_in_1616, d_out_1617, q_in_1617, d_out_1618, q_in_1618, d_out_1619, q_in_1619, d_out_1620, q_in_1620, d_out_1621, q_in_1621, d_out_1622, q_in_1622, d_out_1623, q_in_1623, d_out_1624, q_in_1624, d_out_1625, q_in_1625, d_out_1626, q_in_1626, d_out_1627, q_in_1627, d_out_1628, q_in_1628, d_out_1629, q_in_1629, d_out_1630, q_in_1630, d_out_1631, q_in_1631, d_out_1632, q_in_1632, d_out_1633, q_in_1633, d_out_1634, q_in_1634, d_out_1635, q_in_1635, d_out_1636, q_in_1636, d_out_1637, q_in_1637, d_out_1638, q_in_1638, d_out_1639, q_in_1639, d_out_1640, q_in_1640, d_out_1641, q_in_1641, d_out_1642, q_in_1642, d_out_1643, q_in_1643, d_out_1644, q_in_1644, d_out_1645, q_in_1645, d_out_1646, q_in_1646, d_out_1647, q_in_1647, d_out_1648, q_in_1648, d_out_1649, q_in_1649, d_out_1650, q_in_1650, d_out_1651, q_in_1651, d_out_1652, q_in_1652, d_out_1653, q_in_1653, d_out_1654, q_in_1654, d_out_1655, q_in_1655, d_out_1656, q_in_1656, d_out_1657, q_in_1657, d_out_1658, q_in_1658, d_out_1659, q_in_1659, d_out_1660, q_in_1660, d_out_1661, q_in_1661, d_out_1662, q_in_1662, d_out_1663, q_in_1663, d_out_1664, q_in_1664, d_out_1665, q_in_1665, d_out_1666, q_in_1666, d_out_1667, q_in_1667, d_out_1668, q_in_1668, d_out_1669, q_in_1669, d_out_1670, q_in_1670, d_out_1671, q_in_1671, d_out_1672, q_in_1672, d_out_1673, q_in_1673, d_out_1674, q_in_1674, d_out_1675, q_in_1675, d_out_1676, q_in_1676, d_out_1677, q_in_1677, d_out_1678, q_in_1678, d_out_1679, q_in_1679, d_out_1680, q_in_1680, d_out_1681, q_in_1681, d_out_1682, q_in_1682, d_out_1683, q_in_1683, d_out_1684, q_in_1684, d_out_1685, q_in_1685, d_out_1686, q_in_1686, d_out_1687, q_in_1687, d_out_1688, q_in_1688, d_out_1689, q_in_1689, d_out_1690, q_in_1690, d_out_1691, q_in_1691, d_out_1692, q_in_1692, d_out_1693, q_in_1693, d_out_1694, q_in_1694, d_out_1695, q_in_1695, d_out_1696, q_in_1696, d_out_1697, q_in_1697, d_out_1698, q_in_1698, d_out_1699, q_in_1699, d_out_1700, q_in_1700, d_out_1701, q_in_1701, d_out_1702, q_in_1702, d_out_1703, q_in_1703, d_out_1704, q_in_1704, d_out_1705, q_in_1705, d_out_1706, q_in_1706, d_out_1707, q_in_1707, d_out_1708, q_in_1708, d_out_1709, q_in_1709, d_out_1710, q_in_1710, d_out_1711, q_in_1711, d_out_1712, q_in_1712, d_out_1713, q_in_1713, d_out_1714, q_in_1714, d_out_1715, q_in_1715, d_out_1716, q_in_1716, d_out_1717, q_in_1717, d_out_1718, q_in_1718, d_out_1719, q_in_1719, d_out_1720, q_in_1720, d_out_1721, q_in_1721, d_out_1722, q_in_1722, d_out_1723, q_in_1723, d_out_1724, q_in_1724, d_out_1725, q_in_1725, d_out_1726, q_in_1726, d_out_1727, q_in_1727, d_out_1728, q_in_1728);
input q_in_1728;
input q_in_1727;
input q_in_1726;
input q_in_1725;
input q_in_1724;
input q_in_1723;
input q_in_1722;
input q_in_1721;
input q_in_1720;
input q_in_1719;
input q_in_1718;
input q_in_1717;
input q_in_1716;
input q_in_1715;
input q_in_1714;
input q_in_1713;
input q_in_1712;
input q_in_1711;
input q_in_1710;
input q_in_1709;
input q_in_1708;
input q_in_1707;
input q_in_1706;
input q_in_1705;
input q_in_1704;
input q_in_1703;
input q_in_1702;
input q_in_1701;
input q_in_1700;
input q_in_1699;
input q_in_1698;
input q_in_1697;
input q_in_1696;
input q_in_1695;
input q_in_1694;
input q_in_1693;
input q_in_1692;
input q_in_1691;
input q_in_1690;
input q_in_1689;
input q_in_1688;
input q_in_1687;
input q_in_1686;
input q_in_1685;
input q_in_1684;
input q_in_1683;
input q_in_1682;
input q_in_1681;
input q_in_1680;
input q_in_1679;
input q_in_1678;
input q_in_1677;
input q_in_1676;
input q_in_1675;
input q_in_1674;
input q_in_1673;
input q_in_1672;
input q_in_1671;
input q_in_1670;
input q_in_1669;
input q_in_1668;
input q_in_1667;
input q_in_1666;
input q_in_1665;
input q_in_1664;
input q_in_1663;
input q_in_1662;
input q_in_1661;
input q_in_1660;
input q_in_1659;
input q_in_1658;
input q_in_1657;
input q_in_1656;
input q_in_1655;
input q_in_1654;
input q_in_1653;
input q_in_1652;
input q_in_1651;
input q_in_1650;
input q_in_1649;
input q_in_1648;
input q_in_1647;
input q_in_1646;
input q_in_1645;
input q_in_1644;
input q_in_1643;
input q_in_1642;
input q_in_1641;
input q_in_1640;
input q_in_1639;
input q_in_1638;
input q_in_1637;
input q_in_1636;
input q_in_1635;
input q_in_1634;
input q_in_1633;
input q_in_1632;
input q_in_1631;
input q_in_1630;
input q_in_1629;
input q_in_1628;
input q_in_1627;
input q_in_1626;
input q_in_1625;
input q_in_1624;
input q_in_1623;
input q_in_1622;
input q_in_1621;
input q_in_1620;
input q_in_1619;
input q_in_1618;
input q_in_1617;
input q_in_1616;
input q_in_1615;
input q_in_1614;
input q_in_1613;
input q_in_1612;
input q_in_1611;
input q_in_1610;
input q_in_1609;
input q_in_1608;
input q_in_1607;
input q_in_1606;
input q_in_1605;
input q_in_1604;
input q_in_1603;
input q_in_1602;
input q_in_1601;
input q_in_1600;
input q_in_1599;
input q_in_1598;
input qn_in_1597;
input q_in_1596;
input q_in_1595;
input q_in_1594;
input q_in_1593;
input q_in_1592;
input q_in_1591;
input q_in_1590;
input q_in_1589;
input q_in_1588;
input q_in_1587;
input q_in_1586;
input q_in_1585;
input q_in_1584;
input q_in_1583;
input qn_in_1582;
input qn_in_1581;
input q_in_1580;
input q_in_1579;
input q_in_1578;
input q_in_1577;
input q_in_1576;
input q_in_1575;
input q_in_1574;
input q_in_1573;
input q_in_1572;
input q_in_1571;
input q_in_1570;
input q_in_1569;
input q_in_1568;
input q_in_1567;
input q_in_1566;
input q_in_1565;
input q_in_1564;
input q_in_1563;
input q_in_1562;
input q_in_1561;
input q_in_1560;
input q_in_1559;
input q_in_1558;
input q_in_1557;
input q_in_1556;
input q_in_1555;
input q_in_1554;
input q_in_1553;
input q_in_1552;
input q_in_1551;
input q_in_1550;
input q_in_1549;
input q_in_1548;
input q_in_1547;
input q_in_1546;
input q_in_1545;
input q_in_1544;
input q_in_1543;
input q_in_1542;
input q_in_1541;
input q_in_1540;
input q_in_1539;
input q_in_1538;
input q_in_1537;
input q_in_1536;
input q_in_1535;
input q_in_1534;
input q_in_1533;
input q_in_1532;
input q_in_1531;
input q_in_1530;
input q_in_1529;
input q_in_1528;
input q_in_1527;
input q_in_1526;
input q_in_1525;
input q_in_1524;
input q_in_1523;
input q_in_1522;
input q_in_1521;
input q_in_1520;
input q_in_1519;
input q_in_1518;
input q_in_1517;
input q_in_1516;
input q_in_1515;
input q_in_1514;
input q_in_1513;
input q_in_1512;
input q_in_1511;
input q_in_1510;
input q_in_1509;
input q_in_1508;
input q_in_1507;
input q_in_1506;
input q_in_1505;
input q_in_1504;
input q_in_1503;
input q_in_1502;
input q_in_1501;
input q_in_1500;
input q_in_1499;
input q_in_1498;
input q_in_1497;
input q_in_1496;
input q_in_1495;
input q_in_1494;
input q_in_1493;
input q_in_1492;
input q_in_1491;
input q_in_1490;
input q_in_1489;
input q_in_1488;
input q_in_1487;
input q_in_1486;
input q_in_1485;
input q_in_1484;
input q_in_1483;
input q_in_1482;
input q_in_1481;
input q_in_1480;
input q_in_1479;
input q_in_1478;
input q_in_1477;
input q_in_1476;
input q_in_1475;
input q_in_1474;
input q_in_1473;
input q_in_1472;
input q_in_1471;
input q_in_1470;
input q_in_1469;
input q_in_1468;
input q_in_1467;
input q_in_1466;
input q_in_1465;
input q_in_1464;
input q_in_1463;
input q_in_1462;
input q_in_1461;
input q_in_1460;
input q_in_1459;
input q_in_1458;
input q_in_1457;
input q_in_1456;
input q_in_1455;
input q_in_1454;
input q_in_1453;
input q_in_1452;
input q_in_1451;
input q_in_1450;
input q_in_1449;
input q_in_1448;
input q_in_1447;
input q_in_1446;
input q_in_1445;
input q_in_1444;
input q_in_1443;
input q_in_1442;
input q_in_1441;
input q_in_1440;
input q_in_1439;
input q_in_1438;
input q_in_1437;
input q_in_1436;
input q_in_1435;
input q_in_1434;
input q_in_1433;
input q_in_1432;
input q_in_1431;
input q_in_1430;
input q_in_1429;
input q_in_1428;
input q_in_1427;
input q_in_1426;
input q_in_1425;
input q_in_1424;
input q_in_1423;
input q_in_1422;
input q_in_1421;
input q_in_1420;
input q_in_1419;
input q_in_1418;
input q_in_1417;
input q_in_1416;
input q_in_1415;
input q_in_1414;
input q_in_1413;
input q_in_1412;
input q_in_1411;
input q_in_1410;
input q_in_1409;
input q_in_1408;
input q_in_1407;
input q_in_1406;
input q_in_1405;
input q_in_1404;
input q_in_1403;
input q_in_1402;
input q_in_1401;
input q_in_1400;
input q_in_1399;
input q_in_1398;
input q_in_1397;
input q_in_1396;
input q_in_1395;
input q_in_1394;
input q_in_1393;
input q_in_1392;
input q_in_1391;
input q_in_1390;
input q_in_1389;
input q_in_1388;
input q_in_1387;
input q_in_1386;
input q_in_1385;
input q_in_1384;
input q_in_1383;
input q_in_1382;
input q_in_1381;
input q_in_1380;
input q_in_1379;
input q_in_1378;
input q_in_1377;
input q_in_1376;
input q_in_1375;
input q_in_1374;
input q_in_1373;
input q_in_1372;
input q_in_1371;
input q_in_1370;
input q_in_1369;
input q_in_1368;
input q_in_1367;
input q_in_1366;
input q_in_1365;
input q_in_1364;
input q_in_1363;
input q_in_1362;
input q_in_1361;
input q_in_1360;
input q_in_1359;
input q_in_1358;
input q_in_1357;
input q_in_1356;
input q_in_1355;
input q_in_1354;
input q_in_1353;
input q_in_1352;
input q_in_1351;
input q_in_1350;
input q_in_1349;
input q_in_1348;
input q_in_1347;
input q_in_1346;
input q_in_1345;
input q_in_1344;
input q_in_1343;
input q_in_1342;
input q_in_1341;
input q_in_1340;
input q_in_1339;
input q_in_1338;
input q_in_1337;
input q_in_1336;
input q_in_1335;
input q_in_1334;
input q_in_1333;
input q_in_1332;
input q_in_1331;
input q_in_1330;
input q_in_1329;
input q_in_1328;
input q_in_1327;
input q_in_1326;
input q_in_1325;
input q_in_1324;
input q_in_1323;
input q_in_1322;
input q_in_1321;
input q_in_1320;
input q_in_1319;
input q_in_1318;
input q_in_1317;
input q_in_1316;
input q_in_1315;
input q_in_1314;
input q_in_1313;
input q_in_1312;
input q_in_1311;
input q_in_1310;
input q_in_1309;
input q_in_1308;
input q_in_1307;
input q_in_1306;
input q_in_1305;
input q_in_1304;
input q_in_1303;
input q_in_1302;
input q_in_1301;
input q_in_1300;
input q_in_1299;
input q_in_1298;
input q_in_1297;
input q_in_1296;
input q_in_1295;
input q_in_1294;
input q_in_1293;
input q_in_1292;
input q_in_1291;
input q_in_1290;
input q_in_1289;
input q_in_1288;
input q_in_1287;
input q_in_1286;
input q_in_1285;
input q_in_1284;
input q_in_1283;
input q_in_1282;
input q_in_1281;
input q_in_1280;
input q_in_1279;
input q_in_1278;
input q_in_1277;
input q_in_1276;
input q_in_1275;
input q_in_1274;
input q_in_1273;
input q_in_1272;
input q_in_1271;
input q_in_1270;
input q_in_1269;
input q_in_1268;
input q_in_1267;
input q_in_1266;
input q_in_1265;
input q_in_1264;
input q_in_1263;
input q_in_1262;
input q_in_1261;
input q_in_1260;
input q_in_1259;
input q_in_1258;
input q_in_1257;
input q_in_1256;
input q_in_1255;
input q_in_1254;
input q_in_1253;
input q_in_1252;
input q_in_1251;
input q_in_1250;
input q_in_1249;
input q_in_1248;
input q_in_1247;
input q_in_1246;
input q_in_1245;
input q_in_1244;
input q_in_1243;
input q_in_1242;
input q_in_1241;
input q_in_1240;
input q_in_1239;
input q_in_1238;
input q_in_1237;
input q_in_1236;
input q_in_1235;
input q_in_1234;
input q_in_1233;
input q_in_1232;
input q_in_1231;
input q_in_1230;
input q_in_1229;
input q_in_1228;
input q_in_1227;
input q_in_1226;
input q_in_1225;
input q_in_1224;
input q_in_1223;
input q_in_1222;
input q_in_1221;
input q_in_1220;
input q_in_1219;
input q_in_1218;
input q_in_1217;
input q_in_1216;
input q_in_1215;
input q_in_1214;
input q_in_1213;
input q_in_1212;
input q_in_1211;
input q_in_1210;
input q_in_1209;
input q_in_1208;
input q_in_1207;
input q_in_1206;
input q_in_1205;
input q_in_1204;
input q_in_1203;
input q_in_1202;
input q_in_1201;
input q_in_1200;
input q_in_1199;
input q_in_1198;
input q_in_1197;
input q_in_1196;
input q_in_1195;
input q_in_1194;
input q_in_1193;
input q_in_1192;
input q_in_1191;
input q_in_1190;
input q_in_1189;
input q_in_1188;
input q_in_1187;
input q_in_1186;
input q_in_1185;
input q_in_1184;
input q_in_1183;
input q_in_1182;
input q_in_1181;
input q_in_1180;
input q_in_1179;
input q_in_1178;
input q_in_1177;
input q_in_1176;
input q_in_1175;
input q_in_1174;
input q_in_1173;
input q_in_1172;
input q_in_1171;
input q_in_1170;
input q_in_1169;
input q_in_1168;
input q_in_1167;
input q_in_1166;
input q_in_1165;
input q_in_1164;
input q_in_1163;
input q_in_1162;
input q_in_1161;
input q_in_1160;
input q_in_1159;
input q_in_1158;
input q_in_1157;
input q_in_1156;
input q_in_1155;
input q_in_1154;
input q_in_1153;
input q_in_1152;
input q_in_1151;
input q_in_1150;
input q_in_1149;
input q_in_1148;
input q_in_1147;
input q_in_1146;
input q_in_1145;
input q_in_1144;
input q_in_1143;
input q_in_1142;
input q_in_1141;
input q_in_1140;
input q_in_1139;
input q_in_1138;
input q_in_1137;
input q_in_1136;
input q_in_1135;
input q_in_1134;
input q_in_1133;
input q_in_1132;
input q_in_1131;
input q_in_1130;
input q_in_1129;
input q_in_1128;
input q_in_1127;
input q_in_1126;
input q_in_1125;
input q_in_1124;
input q_in_1123;
input q_in_1122;
input q_in_1121;
input q_in_1120;
input q_in_1119;
input q_in_1118;
input q_in_1117;
input q_in_1116;
input q_in_1115;
input q_in_1114;
input q_in_1113;
input q_in_1112;
input q_in_1111;
input q_in_1110;
input q_in_1109;
input q_in_1108;
input q_in_1107;
input q_in_1106;
input q_in_1105;
input q_in_1104;
input q_in_1103;
input q_in_1102;
input q_in_1101;
input q_in_1100;
input q_in_1099;
input q_in_1098;
input q_in_1097;
input q_in_1096;
input q_in_1095;
input q_in_1094;
input q_in_1093;
input q_in_1092;
input q_in_1091;
input q_in_1090;
input q_in_1089;
input q_in_1088;
input q_in_1087;
input q_in_1086;
input q_in_1085;
input q_in_1084;
input q_in_1083;
input q_in_1082;
input q_in_1081;
input q_in_1080;
input q_in_1079;
input q_in_1078;
input q_in_1077;
input q_in_1076;
input q_in_1075;
input q_in_1074;
input q_in_1073;
input q_in_1072;
input q_in_1071;
input q_in_1070;
input q_in_1069;
input q_in_1068;
input q_in_1067;
input q_in_1066;
input q_in_1065;
input q_in_1064;
input q_in_1063;
input q_in_1062;
input q_in_1061;
input q_in_1060;
input q_in_1059;
input q_in_1058;
input q_in_1057;
input q_in_1056;
input q_in_1055;
input q_in_1054;
input q_in_1053;
input q_in_1052;
input q_in_1051;
input q_in_1050;
input q_in_1049;
input q_in_1048;
input q_in_1047;
input q_in_1046;
input q_in_1045;
input q_in_1044;
input q_in_1043;
input q_in_1042;
input q_in_1041;
input q_in_1040;
input q_in_1039;
input q_in_1038;
input q_in_1037;
input q_in_1036;
input q_in_1035;
input q_in_1034;
input q_in_1033;
input q_in_1032;
input q_in_1031;
input q_in_1030;
input q_in_1029;
input q_in_1028;
input q_in_1027;
input q_in_1026;
input q_in_1025;
input q_in_1024;
input q_in_1023;
input q_in_1022;
input q_in_1021;
input q_in_1020;
input q_in_1019;
input q_in_1018;
input q_in_1017;
input q_in_1016;
input q_in_1015;
input q_in_1014;
input q_in_1013;
input q_in_1012;
input q_in_1011;
input q_in_1010;
input q_in_1009;
input q_in_1008;
input q_in_1007;
input q_in_1006;
input q_in_1005;
input q_in_1004;
input q_in_1003;
input q_in_1002;
input q_in_1001;
input q_in_1000;
input q_in_999;
input q_in_998;
input q_in_997;
input q_in_996;
input q_in_995;
input q_in_994;
input q_in_993;
input q_in_992;
input q_in_991;
input q_in_990;
input q_in_989;
input q_in_988;
input q_in_987;
input q_in_986;
input q_in_985;
input q_in_984;
input q_in_983;
input q_in_982;
input q_in_981;
input q_in_980;
input q_in_979;
input q_in_978;
input q_in_977;
input q_in_976;
input q_in_975;
input q_in_974;
input q_in_973;
input q_in_972;
input q_in_971;
input q_in_970;
input q_in_969;
input q_in_968;
input q_in_967;
input q_in_966;
input q_in_965;
input q_in_964;
input q_in_963;
input q_in_962;
input q_in_961;
input q_in_960;
input q_in_959;
input q_in_958;
input qn_in_957;
input q_in_956;
input q_in_955;
input q_in_954;
input q_in_953;
input q_in_952;
input q_in_951;
input q_in_950;
input q_in_949;
input q_in_948;
input q_in_947;
input q_in_946;
input q_in_945;
input q_in_944;
input q_in_943;
input q_in_942;
input q_in_941;
input q_in_940;
input q_in_939;
input q_in_938;
input q_in_937;
input q_in_936;
input q_in_935;
input q_in_934;
input q_in_933;
input q_in_932;
input q_in_931;
input q_in_930;
input q_in_929;
input q_in_928;
input q_in_927;
input q_in_926;
input q_in_925;
input q_in_924;
input q_in_923;
input q_in_922;
input q_in_921;
input q_in_920;
input q_in_919;
input q_in_918;
input q_in_917;
input q_in_916;
input q_in_915;
input q_in_914;
input q_in_913;
input q_in_912;
input q_in_911;
input q_in_910;
input q_in_909;
input q_in_908;
input q_in_907;
input q_in_906;
input q_in_905;
input q_in_904;
input q_in_903;
input q_in_902;
input q_in_901;
input q_in_900;
input q_in_899;
input q_in_898;
input q_in_897;
input q_in_896;
input q_in_895;
input q_in_894;
input q_in_893;
input q_in_892;
input q_in_891;
input q_in_890;
input q_in_889;
input q_in_888;
input q_in_887;
input q_in_886;
input q_in_885;
input q_in_884;
input q_in_883;
input q_in_882;
input q_in_881;
input q_in_880;
input q_in_879;
input q_in_878;
input q_in_877;
input q_in_876;
input q_in_875;
input q_in_874;
input q_in_873;
input q_in_872;
input q_in_871;
input q_in_870;
input q_in_869;
input q_in_868;
input q_in_867;
input q_in_866;
input q_in_865;
input q_in_864;
input q_in_863;
input q_in_862;
input q_in_861;
input q_in_860;
input q_in_859;
input q_in_858;
input q_in_857;
input q_in_856;
input q_in_855;
input q_in_854;
input q_in_853;
input q_in_852;
input q_in_851;
input q_in_850;
input q_in_849;
input q_in_848;
input q_in_847;
input q_in_846;
input q_in_845;
input q_in_844;
input q_in_843;
input q_in_842;
input q_in_841;
input q_in_840;
input q_in_839;
input q_in_838;
input q_in_837;
input q_in_836;
input q_in_835;
input q_in_834;
input q_in_833;
input q_in_832;
input q_in_831;
input q_in_830;
input q_in_829;
input q_in_828;
input q_in_827;
input q_in_826;
input q_in_825;
input q_in_824;
input q_in_823;
input q_in_822;
input q_in_821;
input q_in_820;
input q_in_819;
input q_in_818;
input q_in_817;
input q_in_816;
input q_in_815;
input q_in_814;
input q_in_813;
input q_in_812;
input q_in_811;
input q_in_810;
input q_in_809;
input q_in_808;
input q_in_807;
input q_in_806;
input q_in_805;
input q_in_804;
input q_in_803;
input q_in_802;
input q_in_801;
input q_in_800;
input q_in_799;
input q_in_798;
input q_in_797;
input q_in_796;
input q_in_795;
input q_in_794;
input q_in_793;
input q_in_792;
input q_in_791;
input q_in_790;
input q_in_789;
input q_in_788;
input q_in_787;
input q_in_786;
input q_in_785;
input q_in_784;
input q_in_783;
input q_in_782;
input q_in_781;
input q_in_780;
input q_in_779;
input q_in_778;
input q_in_777;
input q_in_776;
input q_in_775;
input q_in_774;
input q_in_773;
input q_in_772;
input q_in_771;
input q_in_770;
input q_in_769;
input q_in_768;
input q_in_767;
input q_in_766;
input q_in_765;
input q_in_764;
input q_in_763;
input q_in_762;
input q_in_761;
input q_in_760;
input q_in_759;
input q_in_758;
input q_in_757;
input q_in_756;
input q_in_755;
input q_in_754;
input q_in_753;
input q_in_752;
input q_in_751;
input q_in_750;
input q_in_749;
input q_in_748;
input qn_in_747;
input q_in_746;
input q_in_745;
input q_in_744;
input q_in_743;
input q_in_742;
input q_in_741;
input q_in_740;
input q_in_739;
input q_in_738;
input qn_in_737;
input q_in_736;
input q_in_735;
input qn_in_734;
input q_in_733;
input q_in_732;
input q_in_731;
input q_in_730;
input q_in_729;
input q_in_728;
input q_in_727;
input q_in_726;
input q_in_725;
input q_in_724;
input q_in_723;
input q_in_722;
input q_in_721;
input q_in_720;
input q_in_719;
input q_in_718;
input q_in_717;
input q_in_716;
input q_in_715;
input q_in_714;
input q_in_713;
input q_in_712;
input q_in_711;
input q_in_710;
input q_in_709;
input q_in_708;
input q_in_707;
input q_in_706;
input q_in_705;
input q_in_704;
input q_in_703;
input q_in_702;
input q_in_701;
input q_in_700;
input q_in_699;
input q_in_698;
input q_in_697;
input q_in_696;
input q_in_695;
input q_in_694;
input q_in_693;
input q_in_692;
input q_in_691;
input q_in_690;
input q_in_689;
input q_in_688;
input q_in_687;
input q_in_686;
input q_in_685;
input q_in_684;
input q_in_683;
input q_in_682;
input q_in_681;
input q_in_680;
input q_in_679;
input q_in_678;
input q_in_677;
input q_in_676;
input q_in_675;
input q_in_674;
input q_in_673;
input q_in_672;
input q_in_671;
input q_in_670;
input q_in_669;
input q_in_668;
input q_in_667;
input q_in_666;
input q_in_665;
input q_in_664;
input q_in_663;
input q_in_662;
input q_in_661;
input q_in_660;
input q_in_659;
input q_in_658;
input q_in_657;
input q_in_656;
input q_in_655;
input q_in_654;
input q_in_653;
input q_in_652;
input q_in_651;
input q_in_650;
input q_in_649;
input q_in_648;
input q_in_647;
input qn_in_646;
input q_in_645;
input q_in_644;
input q_in_643;
input q_in_642;
input q_in_641;
input q_in_640;
input q_in_639;
input q_in_638;
input q_in_637;
input q_in_636;
input q_in_635;
input q_in_634;
input q_in_633;
input q_in_632;
input q_in_631;
input q_in_630;
input q_in_629;
input q_in_628;
input q_in_627;
input q_in_626;
input q_in_625;
input q_in_624;
input q_in_623;
input q_in_622;
input q_in_621;
input q_in_620;
input q_in_619;
input q_in_618;
input q_in_617;
input q_in_616;
input q_in_615;
input q_in_614;
input q_in_613;
input q_in_612;
input q_in_611;
input q_in_610;
input q_in_609;
input q_in_608;
input q_in_607;
input q_in_606;
input q_in_605;
input q_in_604;
input q_in_603;
input q_in_602;
input q_in_601;
input q_in_600;
input q_in_599;
input q_in_598;
input q_in_597;
input q_in_596;
input q_in_595;
input q_in_594;
input q_in_593;
input q_in_592;
input q_in_591;
input q_in_590;
input q_in_589;
input q_in_588;
input qn_in_587;
input qn_in_586;
input qn_in_585;
input q_in_584;
input q_in_583;
input q_in_582;
input q_in_581;
input q_in_580;
input q_in_579;
input q_in_578;
input q_in_577;
input q_in_576;
input q_in_575;
input q_in_574;
input q_in_573;
input q_in_572;
input q_in_571;
input q_in_570;
input q_in_569;
input q_in_568;
input q_in_567;
input q_in_566;
input q_in_565;
input q_in_564;
input qn_in_563;
input q_in_562;
input q_in_561;
input q_in_560;
input qn_in_559;
input q_in_558;
input qn_in_557;
input qn_in_556;
input qn_in_555;
input qn_in_554;
input qn_in_553;
input qn_in_552;
input qn_in_551;
input qn_in_550;
input q_in_549;
input q_in_548;
input q_in_547;
input qn_in_546;
input qn_in_545;
input qn_in_544;
input qn_in_543;
input qn_in_542;
input qn_in_541;
input q_in_540;
input qn_in_539;
input qn_in_538;
input qn_in_537;
input qn_in_536;
input qn_in_535;
input qn_in_534;
input qn_in_533;
input qn_in_532;
input qn_in_531;
input qn_in_530;
input qn_in_529;
input qn_in_528;
input qn_in_527;
input qn_in_526;
input qn_in_525;
input qn_in_524;
input qn_in_523;
input qn_in_522;
input qn_in_521;
input qn_in_520;
input qn_in_519;
input qn_in_518;
input q_in_517;
input q_in_516;
input q_in_515;
input q_in_514;
input q_in_513;
input q_in_512;
input qn_in_511;
input qn_in_510;
input qn_in_509;
input q_in_508;
input qn_in_507;
input q_in_506;
input q_in_505;
input qn_in_504;
input q_in_503;
input q_in_502;
input q_in_501;
input q_in_500;
input q_in_499;
input q_in_498;
input q_in_497;
input q_in_496;
input q_in_495;
input q_in_494;
input q_in_493;
input q_in_492;
input q_in_491;
input q_in_490;
input q_in_489;
input q_in_488;
input q_in_487;
input q_in_486;
input q_in_485;
input q_in_484;
input q_in_483;
input q_in_482;
input q_in_481;
input q_in_480;
input q_in_479;
input q_in_478;
input q_in_477;
input q_in_476;
input q_in_475;
input q_in_474;
input q_in_473;
input q_in_472;
input qn_in_471;
input qn_in_470;
input qn_in_469;
input q_in_468;
input q_in_467;
input q_in_466;
input q_in_465;
input q_in_464;
input q_in_463;
input q_in_462;
input q_in_461;
input q_in_460;
input qn_in_459;
input qn_in_458;
input qn_in_457;
input qn_in_456;
input qn_in_455;
input qn_in_454;
input q_in_453;
input q_in_452;
input q_in_451;
input q_in_450;
input q_in_449;
input q_in_448;
input q_in_447;
input qn_in_446;
input qn_in_445;
input qn_in_444;
input qn_in_443;
input q_in_442;
input q_in_441;
input q_in_440;
input qn_in_439;
input qn_in_438;
input qn_in_437;
input qn_in_436;
input q_in_435;
input q_in_434;
input q_in_433;
input q_in_432;
input qn_in_431;
input qn_in_430;
input qn_in_429;
input qn_in_428;
input qn_in_427;
input qn_in_426;
input q_in_425;
input q_in_424;
input q_in_423;
input q_in_422;
input q_in_421;
input q_in_420;
input q_in_419;
input q_in_418;
input q_in_417;
input q_in_416;
input q_in_415;
input q_in_414;
input qn_in_413;
input qn_in_412;
input qn_in_411;
input q_in_410;
input q_in_409;
input q_in_408;
input qn_in_407;
input qn_in_406;
input qn_in_405;
input qn_in_404;
input qn_in_403;
input q_in_402;
input q_in_401;
input q_in_400;
input q_in_399;
input q_in_398;
input q_in_397;
input qn_in_396;
input qn_in_395;
input qn_in_394;
input qn_in_393;
input qn_in_392;
input qn_in_391;
input q_in_390;
input q_in_389;
input q_in_388;
input q_in_387;
input q_in_386;
input q_in_385;
input qn_in_384;
input qn_in_383;
input qn_in_382;
input q_in_381;
input q_in_380;
input q_in_379;
input qn_in_378;
input qn_in_377;
input qn_in_376;
input q_in_375;
input qn_in_374;
input qn_in_373;
input q_in_372;
input q_in_371;
input q_in_370;
input q_in_369;
input q_in_368;
input qn_in_367;
input qn_in_366;
input qn_in_365;
input qn_in_364;
input qn_in_363;
input qn_in_362;
input q_in_361;
input q_in_360;
input q_in_359;
input q_in_358;
input q_in_357;
input q_in_356;
input q_in_355;
input qn_in_354;
input qn_in_353;
input qn_in_352;
input q_in_351;
input q_in_350;
input q_in_349;
input qn_in_348;
input qn_in_347;
input qn_in_346;
input qn_in_345;
input qn_in_344;
input qn_in_343;
input q_in_342;
input q_in_341;
input q_in_340;
input q_in_339;
input q_in_338;
input q_in_337;
input qn_in_336;
input qn_in_335;
input qn_in_334;
input qn_in_333;
input qn_in_332;
input q_in_331;
input q_in_330;
input q_in_329;
input q_in_328;
input q_in_327;
input q_in_326;
input q_in_325;
input qn_in_324;
input qn_in_323;
input qn_in_322;
input q_in_321;
input qn_in_320;
input q_in_319;
input q_in_318;
input qn_in_317;
input qn_in_316;
input qn_in_315;
input qn_in_314;
input qn_in_313;
input q_in_312;
input q_in_311;
input q_in_310;
input q_in_309;
input q_in_308;
input qn_in_307;
input qn_in_306;
input qn_in_305;
input qn_in_304;
input q_in_303;
input q_in_302;
input q_in_301;
input q_in_300;
input q_in_299;
input q_in_298;
input q_in_297;
input qn_in_296;
input qn_in_295;
input qn_in_294;
input q_in_293;
input q_in_292;
input q_in_291;
input q_in_290;
input qn_in_289;
input qn_in_288;
input qn_in_287;
input qn_in_286;
input qn_in_285;
input qn_in_284;
input q_in_283;
input q_in_282;
input q_in_281;
input q_in_280;
input q_in_279;
input qn_in_278;
input qn_in_277;
input qn_in_276;
input q_in_275;
input q_in_274;
input q_in_273;
input q_in_272;
input q_in_271;
input qn_in_270;
input q_in_269;
input qn_in_268;
input qn_in_267;
input qn_in_266;
input q_in_265;
input q_in_264;
input q_in_263;
input qn_in_262;
input qn_in_261;
input qn_in_260;
input qn_in_259;
input q_in_258;
input qn_in_257;
input q_in_256;
input q_in_255;
input q_in_254;
input q_in_253;
input q_in_252;
input qn_in_251;
input qn_in_250;
input q_in_249;
input q_in_248;
input q_in_247;
input q_in_246;
input qn_in_245;
input qn_in_244;
input qn_in_243;
input qn_in_242;
input q_in_241;
input q_in_240;
input q_in_239;
input qn_in_238;
input qn_in_237;
input q_in_236;
input qn_in_235;
input qn_in_234;
input qn_in_233;
input q_in_232;
input q_in_231;
input q_in_230;
input q_in_229;
input q_in_228;
input qn_in_227;
input q_in_226;
input q_in_225;
input q_in_224;
input q_in_223;
input qn_in_222;
input qn_in_221;
input qn_in_220;
input qn_in_219;
input q_in_218;
input q_in_217;
input q_in_216;
input qn_in_215;
input qn_in_214;
input qn_in_213;
input qn_in_212;
input qn_in_211;
input q_in_210;
input q_in_209;
input q_in_208;
input q_in_207;
input q_in_206;
input q_in_205;
input q_in_204;
input q_in_203;
input qn_in_202;
input qn_in_201;
input q_in_200;
input qn_in_199;
input qn_in_198;
input q_in_197;
input q_in_196;
input q_in_195;
input qn_in_194;
input qn_in_193;
input qn_in_192;
input qn_in_191;
input q_in_190;
input q_in_189;
input q_in_188;
input q_in_187;
input q_in_186;
input q_in_185;
input q_in_184;
input qn_in_183;
input qn_in_182;
input qn_in_181;
input q_in_180;
input q_in_179;
input q_in_178;
input q_in_177;
input qn_in_176;
input qn_in_175;
input qn_in_174;
input qn_in_173;
input qn_in_172;
input q_in_171;
input q_in_170;
input q_in_169;
input q_in_168;
input q_in_167;
input qn_in_166;
input qn_in_165;
input qn_in_164;
input q_in_163;
input q_in_162;
input q_in_161;
input q_in_160;
input qn_in_159;
input qn_in_158;
input qn_in_157;
input qn_in_156;
input qn_in_155;
input q_in_154;
input q_in_153;
input q_in_152;
input q_in_151;
input q_in_150;
input q_in_149;
input qn_in_148;
input qn_in_147;
input qn_in_146;
input q_in_145;
input q_in_144;
input q_in_143;
input q_in_142;
input q_in_141;
input qn_in_140;
input qn_in_139;
input qn_in_138;
input qn_in_137;
input q_in_136;
input q_in_135;
input q_in_134;
input q_in_133;
input q_in_132;
input q_in_131;
input q_in_130;
input qn_in_129;
input qn_in_128;
input q_in_127;
input q_in_126;
input q_in_125;
input q_in_124;
input qn_in_123;
input qn_in_122;
input qn_in_121;
input q_in_120;
input q_in_119;
input q_in_118;
input q_in_117;
input q_in_116;
input q_in_115;
input q_in_114;
input q_in_113;
input qn_in_112;
input qn_in_111;
input q_in_110;
input q_in_109;
input q_in_108;
input q_in_107;
input q_in_106;
input qn_in_105;
input qn_in_104;
input q_in_103;
input q_in_102;
input q_in_101;
input q_in_100;
input q_in_99;
input qn_in_98;
input qn_in_97;
input q_in_96;
input q_in_95;
input q_in_94;
input q_in_93;
input q_in_92;
input q_in_91;
input qn_in_90;
input q_in_89;
input q_in_88;
input q_in_87;
input q_in_86;
input q_in_85;
input qn_in_84;
input qn_in_83;
input q_in_82;
input q_in_81;
input q_in_80;
input q_in_79;
input q_in_78;
input q_in_77;
input q_in_76;
input q_in_75;
input qn_in_74;
input qn_in_73;
input q_in_72;
input q_in_71;
input q_in_70;
input q_in_69;
input q_in_68;
input q_in_67;
input q_in_66;
input qn_in_65;
input qn_in_64;
input q_in_63;
input q_in_62;
input q_in_61;
input q_in_60;
input qn_in_59;
input qn_in_58;
input q_in_57;
input q_in_56;
input q_in_55;
input q_in_54;
input qn_in_53;
input qn_in_52;
input q_in_51;
input q_in_50;
input q_in_49;
input qn_in_48;
input qn_in_47;
input q_in_46;
input q_in_45;
input q_in_44;
input q_in_43;
input qn_in_42;
input qn_in_41;
input q_in_40;
input q_in_39;
input q_in_38;
input q_in_37;
input qn_in_36;
input qn_in_35;
input q_in_34;
input q_in_33;
input q_in_32;
input q_in_31;
input qn_in_30;
input qn_in_29;
input q_in_28;
input q_in_27;
input q_in_26;
input qn_in_25;
input qn_in_24;
input q_in_23;
input q_in_22;
input q_in_21;
input q_in_20;
input q_in_19;
input q_in_18;
input q_in_17;
input q_in_16;
input q_in_15;
input q_in_14;
input q_in_13;
input q_in_12;
input q_in_11;
input q_in_10;
input q_in_9;
input q_in_8;
input q_in_7;
input q_in_6;
input q_in_5;
input q_in_4;
input q_in_3;
input q_in_2;
input q_in_1;
input blif_clk_net, blif_reset_net, DATA_0_31, DATA_0_30, DATA_0_29, DATA_0_28, DATA_0_27, DATA_0_26, DATA_0_25, DATA_0_24, DATA_0_23, DATA_0_22, DATA_0_21, DATA_0_20, DATA_0_19, DATA_0_18, DATA_0_17, DATA_0_16, DATA_0_15, DATA_0_14, DATA_0_13, DATA_0_12, DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8, DATA_0_7, DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2, DATA_0_1, DATA_0_0, RESET, TM1, TM0;
output d_out_1728;
output d_out_1727;
output d_out_1726;
output d_out_1725;
output d_out_1724;
output d_out_1723;
output d_out_1722;
output d_out_1721;
output d_out_1720;
output d_out_1719;
output d_out_1718;
output d_out_1717;
output d_out_1716;
output d_out_1715;
output d_out_1714;
output d_out_1713;
output d_out_1712;
output d_out_1711;
output d_out_1710;
output d_out_1709;
output d_out_1708;
output d_out_1707;
output d_out_1706;
output d_out_1705;
output d_out_1704;
output d_out_1703;
output d_out_1702;
output d_out_1701;
output d_out_1700;
output d_out_1699;
output d_out_1698;
output d_out_1697;
output d_out_1696;
output d_out_1695;
output d_out_1694;
output d_out_1693;
output d_out_1692;
output d_out_1691;
output d_out_1690;
output d_out_1689;
output d_out_1688;
output d_out_1687;
output d_out_1686;
output d_out_1685;
output d_out_1684;
output d_out_1683;
output d_out_1682;
output d_out_1681;
output d_out_1680;
output d_out_1679;
output d_out_1678;
output d_out_1677;
output d_out_1676;
output d_out_1675;
output d_out_1674;
output d_out_1673;
output d_out_1672;
output d_out_1671;
output d_out_1670;
output d_out_1669;
output d_out_1668;
output d_out_1667;
output d_out_1666;
output d_out_1665;
output d_out_1664;
output d_out_1663;
output d_out_1662;
output d_out_1661;
output d_out_1660;
output d_out_1659;
output d_out_1658;
output d_out_1657;
output d_out_1656;
output d_out_1655;
output d_out_1654;
output d_out_1653;
output d_out_1652;
output d_out_1651;
output d_out_1650;
output d_out_1649;
output d_out_1648;
output d_out_1647;
output d_out_1646;
output d_out_1645;
output d_out_1644;
output d_out_1643;
output d_out_1642;
output d_out_1641;
output d_out_1640;
output d_out_1639;
output d_out_1638;
output d_out_1637;
output d_out_1636;
output d_out_1635;
output d_out_1634;
output d_out_1633;
output d_out_1632;
output d_out_1631;
output d_out_1630;
output d_out_1629;
output d_out_1628;
output d_out_1627;
output d_out_1626;
output d_out_1625;
output d_out_1624;
output d_out_1623;
output d_out_1622;
output d_out_1621;
output d_out_1620;
output d_out_1619;
output d_out_1618;
output d_out_1617;
output d_out_1616;
output d_out_1615;
output d_out_1614;
output d_out_1613;
output d_out_1612;
output d_out_1611;
output d_out_1610;
output d_out_1609;
output d_out_1608;
output d_out_1607;
output d_out_1606;
output d_out_1605;
output d_out_1604;
output d_out_1603;
output d_out_1602;
output d_out_1601;
output d_out_1600;
output d_out_1599;
output d_out_1598;
output d_out_1597;
output d_out_1596;
output d_out_1595;
output d_out_1594;
output d_out_1593;
output d_out_1592;
output d_out_1591;
output d_out_1590;
output d_out_1589;
output d_out_1588;
output d_out_1587;
output d_out_1586;
output d_out_1585;
output d_out_1584;
output d_out_1583;
output d_out_1582;
output d_out_1581;
output d_out_1580;
output d_out_1579;
output d_out_1578;
output d_out_1577;
output d_out_1576;
output d_out_1575;
output d_out_1574;
output d_out_1573;
output d_out_1572;
output d_out_1571;
output d_out_1570;
output d_out_1569;
output d_out_1568;
output d_out_1567;
output d_out_1566;
output d_out_1565;
output d_out_1564;
output d_out_1563;
output d_out_1562;
output d_out_1561;
output d_out_1560;
output d_out_1559;
output d_out_1558;
output d_out_1557;
output d_out_1556;
output d_out_1555;
output d_out_1554;
output d_out_1553;
output d_out_1552;
output d_out_1551;
output d_out_1550;
output d_out_1549;
output d_out_1548;
output d_out_1547;
output d_out_1546;
output d_out_1545;
output d_out_1544;
output d_out_1543;
output d_out_1542;
output d_out_1541;
output d_out_1540;
output d_out_1539;
output d_out_1538;
output d_out_1537;
output d_out_1536;
output d_out_1535;
output d_out_1534;
output d_out_1533;
output d_out_1532;
output d_out_1531;
output d_out_1530;
output d_out_1529;
output d_out_1528;
output d_out_1527;
output d_out_1526;
output d_out_1525;
output d_out_1524;
output d_out_1523;
output d_out_1522;
output d_out_1521;
output d_out_1520;
output d_out_1519;
output d_out_1518;
output d_out_1517;
output d_out_1516;
output d_out_1515;
output d_out_1514;
output d_out_1513;
output d_out_1512;
output d_out_1511;
output d_out_1510;
output d_out_1509;
output d_out_1508;
output d_out_1507;
output d_out_1506;
output d_out_1505;
output d_out_1504;
output d_out_1503;
output d_out_1502;
output d_out_1501;
output d_out_1500;
output d_out_1499;
output d_out_1498;
output d_out_1497;
output d_out_1496;
output d_out_1495;
output d_out_1494;
output d_out_1493;
output d_out_1492;
output d_out_1491;
output d_out_1490;
output d_out_1489;
output d_out_1488;
output d_out_1487;
output d_out_1486;
output d_out_1485;
output d_out_1484;
output d_out_1483;
output d_out_1482;
output d_out_1481;
output d_out_1480;
output d_out_1479;
output d_out_1478;
output d_out_1477;
output d_out_1476;
output d_out_1475;
output d_out_1474;
output d_out_1473;
output d_out_1472;
output d_out_1471;
output d_out_1470;
output d_out_1469;
output d_out_1468;
output d_out_1467;
output d_out_1466;
output d_out_1465;
output d_out_1464;
output d_out_1463;
output d_out_1462;
output d_out_1461;
output d_out_1460;
output d_out_1459;
output d_out_1458;
output d_out_1457;
output d_out_1456;
output d_out_1455;
output d_out_1454;
output d_out_1453;
output d_out_1452;
output d_out_1451;
output d_out_1450;
output d_out_1449;
output d_out_1448;
output d_out_1447;
output d_out_1446;
output d_out_1445;
output d_out_1444;
output d_out_1443;
output d_out_1442;
output d_out_1441;
output d_out_1440;
output d_out_1439;
output d_out_1438;
output d_out_1437;
output d_out_1436;
output d_out_1435;
output d_out_1434;
output d_out_1433;
output d_out_1432;
output d_out_1431;
output d_out_1430;
output d_out_1429;
output d_out_1428;
output d_out_1427;
output d_out_1426;
output d_out_1425;
output d_out_1424;
output d_out_1423;
output d_out_1422;
output d_out_1421;
output d_out_1420;
output d_out_1419;
output d_out_1418;
output d_out_1417;
output d_out_1416;
output d_out_1415;
output d_out_1414;
output d_out_1413;
output d_out_1412;
output d_out_1411;
output d_out_1410;
output d_out_1409;
output d_out_1408;
output d_out_1407;
output d_out_1406;
output d_out_1405;
output d_out_1404;
output d_out_1403;
output d_out_1402;
output d_out_1401;
output d_out_1400;
output d_out_1399;
output d_out_1398;
output d_out_1397;
output d_out_1396;
output d_out_1395;
output d_out_1394;
output d_out_1393;
output d_out_1392;
output d_out_1391;
output d_out_1390;
output d_out_1389;
output d_out_1388;
output d_out_1387;
output d_out_1386;
output d_out_1385;
output d_out_1384;
output d_out_1383;
output d_out_1382;
output d_out_1381;
output d_out_1380;
output d_out_1379;
output d_out_1378;
output d_out_1377;
output d_out_1376;
output d_out_1375;
output d_out_1374;
output d_out_1373;
output d_out_1372;
output d_out_1371;
output d_out_1370;
output d_out_1369;
output d_out_1368;
output d_out_1367;
output d_out_1366;
output d_out_1365;
output d_out_1364;
output d_out_1363;
output d_out_1362;
output d_out_1361;
output d_out_1360;
output d_out_1359;
output d_out_1358;
output d_out_1357;
output d_out_1356;
output d_out_1355;
output d_out_1354;
output d_out_1353;
output d_out_1352;
output d_out_1351;
output d_out_1350;
output d_out_1349;
output d_out_1348;
output d_out_1347;
output d_out_1346;
output d_out_1345;
output d_out_1344;
output d_out_1343;
output d_out_1342;
output d_out_1341;
output d_out_1340;
output d_out_1339;
output d_out_1338;
output d_out_1337;
output d_out_1336;
output d_out_1335;
output d_out_1334;
output d_out_1333;
output d_out_1332;
output d_out_1331;
output d_out_1330;
output d_out_1329;
output d_out_1328;
output d_out_1327;
output d_out_1326;
output d_out_1325;
output d_out_1324;
output d_out_1323;
output d_out_1322;
output d_out_1321;
output d_out_1320;
output d_out_1319;
output d_out_1318;
output d_out_1317;
output d_out_1316;
output d_out_1315;
output d_out_1314;
output d_out_1313;
output d_out_1312;
output d_out_1311;
output d_out_1310;
output d_out_1309;
output d_out_1308;
output d_out_1307;
output d_out_1306;
output d_out_1305;
output d_out_1304;
output d_out_1303;
output d_out_1302;
output d_out_1301;
output d_out_1300;
output d_out_1299;
output d_out_1298;
output d_out_1297;
output d_out_1296;
output d_out_1295;
output d_out_1294;
output d_out_1293;
output d_out_1292;
output d_out_1291;
output d_out_1290;
output d_out_1289;
output d_out_1288;
output d_out_1287;
output d_out_1286;
output d_out_1285;
output d_out_1284;
output d_out_1283;
output d_out_1282;
output d_out_1281;
output d_out_1280;
output d_out_1279;
output d_out_1278;
output d_out_1277;
output d_out_1276;
output d_out_1275;
output d_out_1274;
output d_out_1273;
output d_out_1272;
output d_out_1271;
output d_out_1270;
output d_out_1269;
output d_out_1268;
output d_out_1267;
output d_out_1266;
output d_out_1265;
output d_out_1264;
output d_out_1263;
output d_out_1262;
output d_out_1261;
output d_out_1260;
output d_out_1259;
output d_out_1258;
output d_out_1257;
output d_out_1256;
output d_out_1255;
output d_out_1254;
output d_out_1253;
output d_out_1252;
output d_out_1251;
output d_out_1250;
output d_out_1249;
output d_out_1248;
output d_out_1247;
output d_out_1246;
output d_out_1245;
output d_out_1244;
output d_out_1243;
output d_out_1242;
output d_out_1241;
output d_out_1240;
output d_out_1239;
output d_out_1238;
output d_out_1237;
output d_out_1236;
output d_out_1235;
output d_out_1234;
output d_out_1233;
output d_out_1232;
output d_out_1231;
output d_out_1230;
output d_out_1229;
output d_out_1228;
output d_out_1227;
output d_out_1226;
output d_out_1225;
output d_out_1224;
output d_out_1223;
output d_out_1222;
output d_out_1221;
output d_out_1220;
output d_out_1219;
output d_out_1218;
output d_out_1217;
output d_out_1216;
output d_out_1215;
output d_out_1214;
output d_out_1213;
output d_out_1212;
output d_out_1211;
output d_out_1210;
output d_out_1209;
output d_out_1208;
output d_out_1207;
output d_out_1206;
output d_out_1205;
output d_out_1204;
output d_out_1203;
output d_out_1202;
output d_out_1201;
output d_out_1200;
output d_out_1199;
output d_out_1198;
output d_out_1197;
output d_out_1196;
output d_out_1195;
output d_out_1194;
output d_out_1193;
output d_out_1192;
output d_out_1191;
output d_out_1190;
output d_out_1189;
output d_out_1188;
output d_out_1187;
output d_out_1186;
output d_out_1185;
output d_out_1184;
output d_out_1183;
output d_out_1182;
output d_out_1181;
output d_out_1180;
output d_out_1179;
output d_out_1178;
output d_out_1177;
output d_out_1176;
output d_out_1175;
output d_out_1174;
output d_out_1173;
output d_out_1172;
output d_out_1171;
output d_out_1170;
output d_out_1169;
output d_out_1168;
output d_out_1167;
output d_out_1166;
output d_out_1165;
output d_out_1164;
output d_out_1163;
output d_out_1162;
output d_out_1161;
output d_out_1160;
output d_out_1159;
output d_out_1158;
output d_out_1157;
output d_out_1156;
output d_out_1155;
output d_out_1154;
output d_out_1153;
output d_out_1152;
output d_out_1151;
output d_out_1150;
output d_out_1149;
output d_out_1148;
output d_out_1147;
output d_out_1146;
output d_out_1145;
output d_out_1144;
output d_out_1143;
output d_out_1142;
output d_out_1141;
output d_out_1140;
output d_out_1139;
output d_out_1138;
output d_out_1137;
output d_out_1136;
output d_out_1135;
output d_out_1134;
output d_out_1133;
output d_out_1132;
output d_out_1131;
output d_out_1130;
output d_out_1129;
output d_out_1128;
output d_out_1127;
output d_out_1126;
output d_out_1125;
output d_out_1124;
output d_out_1123;
output d_out_1122;
output d_out_1121;
output d_out_1120;
output d_out_1119;
output d_out_1118;
output d_out_1117;
output d_out_1116;
output d_out_1115;
output d_out_1114;
output d_out_1113;
output d_out_1112;
output d_out_1111;
output d_out_1110;
output d_out_1109;
output d_out_1108;
output d_out_1107;
output d_out_1106;
output d_out_1105;
output d_out_1104;
output d_out_1103;
output d_out_1102;
output d_out_1101;
output d_out_1100;
output d_out_1099;
output d_out_1098;
output d_out_1097;
output d_out_1096;
output d_out_1095;
output d_out_1094;
output d_out_1093;
output d_out_1092;
output d_out_1091;
output d_out_1090;
output d_out_1089;
output d_out_1088;
output d_out_1087;
output d_out_1086;
output d_out_1085;
output d_out_1084;
output d_out_1083;
output d_out_1082;
output d_out_1081;
output d_out_1080;
output d_out_1079;
output d_out_1078;
output d_out_1077;
output d_out_1076;
output d_out_1075;
output d_out_1074;
output d_out_1073;
output d_out_1072;
output d_out_1071;
output d_out_1070;
output d_out_1069;
output d_out_1068;
output d_out_1067;
output d_out_1066;
output d_out_1065;
output d_out_1064;
output d_out_1063;
output d_out_1062;
output d_out_1061;
output d_out_1060;
output d_out_1059;
output d_out_1058;
output d_out_1057;
output d_out_1056;
output d_out_1055;
output d_out_1054;
output d_out_1053;
output d_out_1052;
output d_out_1051;
output d_out_1050;
output d_out_1049;
output d_out_1048;
output d_out_1047;
output d_out_1046;
output d_out_1045;
output d_out_1044;
output d_out_1043;
output d_out_1042;
output d_out_1041;
output d_out_1040;
output d_out_1039;
output d_out_1038;
output d_out_1037;
output d_out_1036;
output d_out_1035;
output d_out_1034;
output d_out_1033;
output d_out_1032;
output d_out_1031;
output d_out_1030;
output d_out_1029;
output d_out_1028;
output d_out_1027;
output d_out_1026;
output d_out_1025;
output d_out_1024;
output d_out_1023;
output d_out_1022;
output d_out_1021;
output d_out_1020;
output d_out_1019;
output d_out_1018;
output d_out_1017;
output d_out_1016;
output d_out_1015;
output d_out_1014;
output d_out_1013;
output d_out_1012;
output d_out_1011;
output d_out_1010;
output d_out_1009;
output d_out_1008;
output d_out_1007;
output d_out_1006;
output d_out_1005;
output d_out_1004;
output d_out_1003;
output d_out_1002;
output d_out_1001;
output d_out_1000;
output d_out_999;
output d_out_998;
output d_out_997;
output d_out_996;
output d_out_995;
output d_out_994;
output d_out_993;
output d_out_992;
output d_out_991;
output d_out_990;
output d_out_989;
output d_out_988;
output d_out_987;
output d_out_986;
output d_out_985;
output d_out_984;
output d_out_983;
output d_out_982;
output d_out_981;
output d_out_980;
output d_out_979;
output d_out_978;
output d_out_977;
output d_out_976;
output d_out_975;
output d_out_974;
output d_out_973;
output d_out_972;
output d_out_971;
output d_out_970;
output d_out_969;
output d_out_968;
output d_out_967;
output d_out_966;
output d_out_965;
output d_out_964;
output d_out_963;
output d_out_962;
output d_out_961;
output d_out_960;
output d_out_959;
output d_out_958;
output d_out_957;
output d_out_956;
output d_out_955;
output d_out_954;
output d_out_953;
output d_out_952;
output d_out_951;
output d_out_950;
output d_out_949;
output d_out_948;
output d_out_947;
output d_out_946;
output d_out_945;
output d_out_944;
output d_out_943;
output d_out_942;
output d_out_941;
output d_out_940;
output d_out_939;
output d_out_938;
output d_out_937;
output d_out_936;
output d_out_935;
output d_out_934;
output d_out_933;
output d_out_932;
output d_out_931;
output d_out_930;
output d_out_929;
output d_out_928;
output d_out_927;
output d_out_926;
output d_out_925;
output d_out_924;
output d_out_923;
output d_out_922;
output d_out_921;
output d_out_920;
output d_out_919;
output d_out_918;
output d_out_917;
output d_out_916;
output d_out_915;
output d_out_914;
output d_out_913;
output d_out_912;
output d_out_911;
output d_out_910;
output d_out_909;
output d_out_908;
output d_out_907;
output d_out_906;
output d_out_905;
output d_out_904;
output d_out_903;
output d_out_902;
output d_out_901;
output d_out_900;
output d_out_899;
output d_out_898;
output d_out_897;
output d_out_896;
output d_out_895;
output d_out_894;
output d_out_893;
output d_out_892;
output d_out_891;
output d_out_890;
output d_out_889;
output d_out_888;
output d_out_887;
output d_out_886;
output d_out_885;
output d_out_884;
output d_out_883;
output d_out_882;
output d_out_881;
output d_out_880;
output d_out_879;
output d_out_878;
output d_out_877;
output d_out_876;
output d_out_875;
output d_out_874;
output d_out_873;
output d_out_872;
output d_out_871;
output d_out_870;
output d_out_869;
output d_out_868;
output d_out_867;
output d_out_866;
output d_out_865;
output d_out_864;
output d_out_863;
output d_out_862;
output d_out_861;
output d_out_860;
output d_out_859;
output d_out_858;
output d_out_857;
output d_out_856;
output d_out_855;
output d_out_854;
output d_out_853;
output d_out_852;
output d_out_851;
output d_out_850;
output d_out_849;
output d_out_848;
output d_out_847;
output d_out_846;
output d_out_845;
output d_out_844;
output d_out_843;
output d_out_842;
output d_out_841;
output d_out_840;
output d_out_839;
output d_out_838;
output d_out_837;
output d_out_836;
output d_out_835;
output d_out_834;
output d_out_833;
output d_out_832;
output d_out_831;
output d_out_830;
output d_out_829;
output d_out_828;
output d_out_827;
output d_out_826;
output d_out_825;
output d_out_824;
output d_out_823;
output d_out_822;
output d_out_821;
output d_out_820;
output d_out_819;
output d_out_818;
output d_out_817;
output d_out_816;
output d_out_815;
output d_out_814;
output d_out_813;
output d_out_812;
output d_out_811;
output d_out_810;
output d_out_809;
output d_out_808;
output d_out_807;
output d_out_806;
output d_out_805;
output d_out_804;
output d_out_803;
output d_out_802;
output d_out_801;
output d_out_800;
output d_out_799;
output d_out_798;
output d_out_797;
output d_out_796;
output d_out_795;
output d_out_794;
output d_out_793;
output d_out_792;
output d_out_791;
output d_out_790;
output d_out_789;
output d_out_788;
output d_out_787;
output d_out_786;
output d_out_785;
output d_out_784;
output d_out_783;
output d_out_782;
output d_out_781;
output d_out_780;
output d_out_779;
output d_out_778;
output d_out_777;
output d_out_776;
output d_out_775;
output d_out_774;
output d_out_773;
output d_out_772;
output d_out_771;
output d_out_770;
output d_out_769;
output d_out_768;
output d_out_767;
output d_out_766;
output d_out_765;
output d_out_764;
output d_out_763;
output d_out_762;
output d_out_761;
output d_out_760;
output d_out_759;
output d_out_758;
output d_out_757;
output d_out_756;
output d_out_755;
output d_out_754;
output d_out_753;
output d_out_752;
output d_out_751;
output d_out_750;
output d_out_749;
output d_out_748;
output d_out_747;
output d_out_746;
output d_out_745;
output d_out_744;
output d_out_743;
output d_out_742;
output d_out_741;
output d_out_740;
output d_out_739;
output d_out_738;
output d_out_737;
output d_out_736;
output d_out_735;
output d_out_734;
output d_out_733;
output d_out_732;
output d_out_731;
output d_out_730;
output d_out_729;
output d_out_728;
output d_out_727;
output d_out_726;
output d_out_725;
output d_out_724;
output d_out_723;
output d_out_722;
output d_out_721;
output d_out_720;
output d_out_719;
output d_out_718;
output d_out_717;
output d_out_716;
output d_out_715;
output d_out_714;
output d_out_713;
output d_out_712;
output d_out_711;
output d_out_710;
output d_out_709;
output d_out_708;
output d_out_707;
output d_out_706;
output d_out_705;
output d_out_704;
output d_out_703;
output d_out_702;
output d_out_701;
output d_out_700;
output d_out_699;
output d_out_698;
output d_out_697;
output d_out_696;
output d_out_695;
output d_out_694;
output d_out_693;
output d_out_692;
output d_out_691;
output d_out_690;
output d_out_689;
output d_out_688;
output d_out_687;
output d_out_686;
output d_out_685;
output d_out_684;
output d_out_683;
output d_out_682;
output d_out_681;
output d_out_680;
output d_out_679;
output d_out_678;
output d_out_677;
output d_out_676;
output d_out_675;
output d_out_674;
output d_out_673;
output d_out_672;
output d_out_671;
output d_out_670;
output d_out_669;
output d_out_668;
output d_out_667;
output d_out_666;
output d_out_665;
output d_out_664;
output d_out_663;
output d_out_662;
output d_out_661;
output d_out_660;
output d_out_659;
output d_out_658;
output d_out_657;
output d_out_656;
output d_out_655;
output d_out_654;
output d_out_653;
output d_out_652;
output d_out_651;
output d_out_650;
output d_out_649;
output d_out_648;
output d_out_647;
output d_out_646;
output d_out_645;
output d_out_644;
output d_out_643;
output d_out_642;
output d_out_641;
output d_out_640;
output d_out_639;
output d_out_638;
output d_out_637;
output d_out_636;
output d_out_635;
output d_out_634;
output d_out_633;
output d_out_632;
output d_out_631;
output d_out_630;
output d_out_629;
output d_out_628;
output d_out_627;
output d_out_626;
output d_out_625;
output d_out_624;
output d_out_623;
output d_out_622;
output d_out_621;
output d_out_620;
output d_out_619;
output d_out_618;
output d_out_617;
output d_out_616;
output d_out_615;
output d_out_614;
output d_out_613;
output d_out_612;
output d_out_611;
output d_out_610;
output d_out_609;
output d_out_608;
output d_out_607;
output d_out_606;
output d_out_605;
output d_out_604;
output d_out_603;
output d_out_602;
output d_out_601;
output d_out_600;
output d_out_599;
output d_out_598;
output d_out_597;
output d_out_596;
output d_out_595;
output d_out_594;
output d_out_593;
output d_out_592;
output d_out_591;
output d_out_590;
output d_out_589;
output d_out_588;
output d_out_587;
output d_out_586;
output d_out_585;
output d_out_584;
output d_out_583;
output d_out_582;
output d_out_581;
output d_out_580;
output d_out_579;
output d_out_578;
output d_out_577;
output d_out_576;
output d_out_575;
output d_out_574;
output d_out_573;
output d_out_572;
output d_out_571;
output d_out_570;
output d_out_569;
output d_out_568;
output d_out_567;
output d_out_566;
output d_out_565;
output d_out_564;
output d_out_563;
output d_out_562;
output d_out_561;
output d_out_560;
output d_out_559;
output d_out_558;
output d_out_557;
output d_out_556;
output d_out_555;
output d_out_554;
output d_out_553;
output d_out_552;
output d_out_551;
output d_out_550;
output d_out_549;
output d_out_548;
output d_out_547;
output d_out_546;
output d_out_545;
output d_out_544;
output d_out_543;
output d_out_542;
output d_out_541;
output d_out_540;
output d_out_539;
output d_out_538;
output d_out_537;
output d_out_536;
output d_out_535;
output d_out_534;
output d_out_533;
output d_out_532;
output d_out_531;
output d_out_530;
output d_out_529;
output d_out_528;
output d_out_527;
output d_out_526;
output d_out_525;
output d_out_524;
output d_out_523;
output d_out_522;
output d_out_521;
output d_out_520;
output d_out_519;
output d_out_518;
output d_out_517;
output d_out_516;
output d_out_515;
output d_out_514;
output d_out_513;
output d_out_512;
output d_out_511;
output d_out_510;
output d_out_509;
output d_out_508;
output d_out_507;
output d_out_506;
output d_out_505;
output d_out_504;
output d_out_503;
output d_out_502;
output d_out_501;
output d_out_500;
output d_out_499;
output d_out_498;
output d_out_497;
output d_out_496;
output d_out_495;
output d_out_494;
output d_out_493;
output d_out_492;
output d_out_491;
output d_out_490;
output d_out_489;
output d_out_488;
output d_out_487;
output d_out_486;
output d_out_485;
output d_out_484;
output d_out_483;
output d_out_482;
output d_out_481;
output d_out_480;
output d_out_479;
output d_out_478;
output d_out_477;
output d_out_476;
output d_out_475;
output d_out_474;
output d_out_473;
output d_out_472;
output d_out_471;
output d_out_470;
output d_out_469;
output d_out_468;
output d_out_467;
output d_out_466;
output d_out_465;
output d_out_464;
output d_out_463;
output d_out_462;
output d_out_461;
output d_out_460;
output d_out_459;
output d_out_458;
output d_out_457;
output d_out_456;
output d_out_455;
output d_out_454;
output d_out_453;
output d_out_452;
output d_out_451;
output d_out_450;
output d_out_449;
output d_out_448;
output d_out_447;
output d_out_446;
output d_out_445;
output d_out_444;
output d_out_443;
output d_out_442;
output d_out_441;
output d_out_440;
output d_out_439;
output d_out_438;
output d_out_437;
output d_out_436;
output d_out_435;
output d_out_434;
output d_out_433;
output d_out_432;
output d_out_431;
output d_out_430;
output d_out_429;
output d_out_428;
output d_out_427;
output d_out_426;
output d_out_425;
output d_out_424;
output d_out_423;
output d_out_422;
output d_out_421;
output d_out_420;
output d_out_419;
output d_out_418;
output d_out_417;
output d_out_416;
output d_out_415;
output d_out_414;
output d_out_413;
output d_out_412;
output d_out_411;
output d_out_410;
output d_out_409;
output d_out_408;
output d_out_407;
output d_out_406;
output d_out_405;
output d_out_404;
output d_out_403;
output d_out_402;
output d_out_401;
output d_out_400;
output d_out_399;
output d_out_398;
output d_out_397;
output d_out_396;
output d_out_395;
output d_out_394;
output d_out_393;
output d_out_392;
output d_out_391;
output d_out_390;
output d_out_389;
output d_out_388;
output d_out_387;
output d_out_386;
output d_out_385;
output d_out_384;
output d_out_383;
output d_out_382;
output d_out_381;
output d_out_380;
output d_out_379;
output d_out_378;
output d_out_377;
output d_out_376;
output d_out_375;
output d_out_374;
output d_out_373;
output d_out_372;
output d_out_371;
output d_out_370;
output d_out_369;
output d_out_368;
output d_out_367;
output d_out_366;
output d_out_365;
output d_out_364;
output d_out_363;
output d_out_362;
output d_out_361;
output d_out_360;
output d_out_359;
output d_out_358;
output d_out_357;
output d_out_356;
output d_out_355;
output d_out_354;
output d_out_353;
output d_out_352;
output d_out_351;
output d_out_350;
output d_out_349;
output d_out_348;
output d_out_347;
output d_out_346;
output d_out_345;
output d_out_344;
output d_out_343;
output d_out_342;
output d_out_341;
output d_out_340;
output d_out_339;
output d_out_338;
output d_out_337;
output d_out_336;
output d_out_335;
output d_out_334;
output d_out_333;
output d_out_332;
output d_out_331;
output d_out_330;
output d_out_329;
output d_out_328;
output d_out_327;
output d_out_326;
output d_out_325;
output d_out_324;
output d_out_323;
output d_out_322;
output d_out_321;
output d_out_320;
output d_out_319;
output d_out_318;
output d_out_317;
output d_out_316;
output d_out_315;
output d_out_314;
output d_out_313;
output d_out_312;
output d_out_311;
output d_out_310;
output d_out_309;
output d_out_308;
output d_out_307;
output d_out_306;
output d_out_305;
output d_out_304;
output d_out_303;
output d_out_302;
output d_out_301;
output d_out_300;
output d_out_299;
output d_out_298;
output d_out_297;
output d_out_296;
output d_out_295;
output d_out_294;
output d_out_293;
output d_out_292;
output d_out_291;
output d_out_290;
output d_out_289;
output d_out_288;
output d_out_287;
output d_out_286;
output d_out_285;
output d_out_284;
output d_out_283;
output d_out_282;
output d_out_281;
output d_out_280;
output d_out_279;
output d_out_278;
output d_out_277;
output d_out_276;
output d_out_275;
output d_out_274;
output d_out_273;
output d_out_272;
output d_out_271;
output d_out_270;
output d_out_269;
output d_out_268;
output d_out_267;
output d_out_266;
output d_out_265;
output d_out_264;
output d_out_263;
output d_out_262;
output d_out_261;
output d_out_260;
output d_out_259;
output d_out_258;
output d_out_257;
output d_out_256;
output d_out_255;
output d_out_254;
output d_out_253;
output d_out_252;
output d_out_251;
output d_out_250;
output d_out_249;
output d_out_248;
output d_out_247;
output d_out_246;
output d_out_245;
output d_out_244;
output d_out_243;
output d_out_242;
output d_out_241;
output d_out_240;
output d_out_239;
output d_out_238;
output d_out_237;
output d_out_236;
output d_out_235;
output d_out_234;
output d_out_233;
output d_out_232;
output d_out_231;
output d_out_230;
output d_out_229;
output d_out_228;
output d_out_227;
output d_out_226;
output d_out_225;
output d_out_224;
output d_out_223;
output d_out_222;
output d_out_221;
output d_out_220;
output d_out_219;
output d_out_218;
output d_out_217;
output d_out_216;
output d_out_215;
output d_out_214;
output d_out_213;
output d_out_212;
output d_out_211;
output d_out_210;
output d_out_209;
output d_out_208;
output d_out_207;
output d_out_206;
output d_out_205;
output d_out_204;
output d_out_203;
output d_out_202;
output d_out_201;
output d_out_200;
output d_out_199;
output d_out_198;
output d_out_197;
output d_out_196;
output d_out_195;
output d_out_194;
output d_out_193;
output d_out_192;
output d_out_191;
output d_out_190;
output d_out_189;
output d_out_188;
output d_out_187;
output d_out_186;
output d_out_185;
output d_out_184;
output d_out_183;
output d_out_182;
output d_out_181;
output d_out_180;
output d_out_179;
output d_out_178;
output d_out_177;
output d_out_176;
output d_out_175;
output d_out_174;
output d_out_173;
output d_out_172;
output d_out_171;
output d_out_170;
output d_out_169;
output d_out_168;
output d_out_167;
output d_out_166;
output d_out_165;
output d_out_164;
output d_out_163;
output d_out_162;
output d_out_161;
output d_out_160;
output d_out_159;
output d_out_158;
output d_out_157;
output d_out_156;
output d_out_155;
output d_out_154;
output d_out_153;
output d_out_152;
output d_out_151;
output d_out_150;
output d_out_149;
output d_out_148;
output d_out_147;
output d_out_146;
output d_out_145;
output d_out_144;
output d_out_143;
output d_out_142;
output d_out_141;
output d_out_140;
output d_out_139;
output d_out_138;
output d_out_137;
output d_out_136;
output d_out_135;
output d_out_134;
output d_out_133;
output d_out_132;
output d_out_131;
output d_out_130;
output d_out_129;
output d_out_128;
output d_out_127;
output d_out_126;
output d_out_125;
output d_out_124;
output d_out_123;
output d_out_122;
output d_out_121;
output d_out_120;
output d_out_119;
output d_out_118;
output d_out_117;
output d_out_116;
output d_out_115;
output d_out_114;
output d_out_113;
output d_out_112;
output d_out_111;
output d_out_110;
output d_out_109;
output d_out_108;
output d_out_107;
output d_out_106;
output d_out_105;
output d_out_104;
output d_out_103;
output d_out_102;
output d_out_101;
output d_out_100;
output d_out_99;
output d_out_98;
output d_out_97;
output d_out_96;
output d_out_95;
output d_out_94;
output d_out_93;
output d_out_92;
output d_out_91;
output d_out_90;
output d_out_89;
output d_out_88;
output d_out_87;
output d_out_86;
output d_out_85;
output d_out_84;
output d_out_83;
output d_out_82;
output d_out_81;
output d_out_80;
output d_out_79;
output d_out_78;
output d_out_77;
output d_out_76;
output d_out_75;
output d_out_74;
output d_out_73;
output d_out_72;
output d_out_71;
output d_out_70;
output d_out_69;
output d_out_68;
output d_out_67;
output d_out_66;
output d_out_65;
output d_out_64;
output d_out_63;
output d_out_62;
output d_out_61;
output d_out_60;
output d_out_59;
output d_out_58;
output d_out_57;
output d_out_56;
output d_out_55;
output d_out_54;
output d_out_53;
output d_out_52;
output d_out_51;
output d_out_50;
output d_out_49;
output d_out_48;
output d_out_47;
output d_out_46;
output d_out_45;
output d_out_44;
output d_out_43;
output d_out_42;
output d_out_41;
output d_out_40;
output d_out_39;
output d_out_38;
output d_out_37;
output d_out_36;
output d_out_35;
output d_out_34;
output d_out_33;
output d_out_32;
output d_out_31;
output d_out_30;
output d_out_29;
output d_out_28;
output d_out_27;
output d_out_26;
output d_out_25;
output d_out_24;
output d_out_23;
output d_out_22;
output d_out_21;
output d_out_20;
output d_out_19;
output d_out_18;
output d_out_17;
output d_out_16;
output d_out_15;
output d_out_14;
output d_out_13;
output d_out_12;
output d_out_11;
output d_out_10;
output d_out_9;
output d_out_8;
output d_out_7;
output d_out_6;
output d_out_5;
output d_out_4;
output d_out_3;
output d_out_2;
output d_out_1;
output DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27, DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22, DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17, DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12, DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7, DATA_9_6, DATA_9_5, DATA_9_4, DATA_9_3, DATA_9_2, DATA_9_1, DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2, CRC_OUT_9_3, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30, CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2, CRC_OUT_7_3, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2, CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2, CRC_OUT_2_3, CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_2, CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31;
wire n_15868;
wire n_15860, n_15861, n_15862, n_15863, n_15864, n_15865, n_15866, n_15867;
wire n_15852, n_15853, n_15854, n_15855, n_15856, n_15857, n_15858, n_15859;
wire n_11621, n_11623, n_11625, n_11626, n_12492, n_12493, n_12494, n_15851;
wire n_11612, n_11613, n_11614, n_11615, n_11616, n_11617, n_11618, n_11619;
wire n_11602, n_11603, n_11604, n_11605, n_11607, n_11608, n_11609, n_11611;
wire n_10746, n_10747, n_11595, n_11596, n_11597, n_11599, n_11600, n_11601;
wire n_10738, n_10739, n_10740, n_10741, n_10742, n_10743, n_10744, n_10745;
wire n_10730, n_10731, n_10732, n_10733, n_10734, n_10735, n_10736, n_10737;
wire n_10722, n_10723, n_10724, n_10725, n_10726, n_10727, n_10728, n_10729;
wire n_10713, n_10714, n_10716, n_10717, n_10718, n_10719, n_10720, n_10721;
wire n_9818, n_9819, n_9820, n_9821, n_9822, n_9823, n_9824, n_10712;
wire n_9797, n_9798, n_9799, n_9800, n_9814, n_9815, n_9816, n_9817;
wire n_9431, n_9432, n_9433, n_9434, n_9435, n_9436, n_9437, n_9438;
wire n_9423, n_9424, n_9425, n_9426, n_9427, n_9428, n_9429, n_9430;
wire n_9414, n_9415, n_9416, n_9418, n_9419, n_9420, n_9421, n_9422;
wire n_9406, n_9407, n_9408, n_9409, n_9410, n_9411, n_9412, n_9413;
wire n_9398, n_9399, n_9400, n_9401, n_9402, n_9403, n_9404, n_9405;
wire n_9390, n_9391, n_9392, n_9393, n_9394, n_9395, n_9396, n_9397;
wire n_8553, n_8554, n_9384, n_9385, n_9386, n_9387, n_9388, n_9389;
wire n_8545, n_8546, n_8547, n_8548, n_8549, n_8550, n_8551, n_8552;
wire n_8355, n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544;
wire n_8347, n_8348, n_8349, n_8350, n_8351, n_8352, n_8353, n_8354;
wire n_8339, n_8340, n_8341, n_8342, n_8343, n_8344, n_8345, n_8346;
wire n_8331, n_8332, n_8333, n_8334, n_8335, n_8336, n_8337, n_8338;
wire n_8323, n_8324, n_8325, n_8326, n_8327, n_8328, n_8329, n_8330;
wire n_8315, n_8316, n_8317, n_8318, n_8319, n_8320, n_8321, n_8322;
wire n_7505, n_7506, n_7507, n_7508, n_7509, n_7510, n_7511, n_8314;
wire n_7482, n_7483, n_7484, n_7485, n_7487, n_7488, n_7490, n_7504;
wire n_7090, n_7092, n_7093, n_7094, n_7281, n_7282, n_7480, n_7481;
wire n_7082, n_7083, n_7084, n_7085, n_7086, n_7087, n_7088, n_7089;
wire n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7080, n_7081;
wire n_7066, n_7067, n_7068, n_7069, n_7070, n_7071, n_7072, n_7073;
wire n_6886, n_7059, n_7060, n_7061, n_7062, n_7063, n_7064, n_7065;
wire n_6696, n_6697, n_6698, n_6699, n_6882, n_6883, n_6884, n_6885;
wire n_6688, n_6689, n_6690, n_6691, n_6692, n_6693, n_6694, n_6695;
wire n_6680, n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687;
wire n_6672, n_6673, n_6674, n_6675, n_6676, n_6677, n_6678, n_6679;
wire n_6664, n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671;
wire n_6644, n_6645, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663;
wire n_6628, n_6629, n_6630, n_6631, n_6632, n_6633, n_6642, n_6643;
wire n_6618, n_6619, n_6620, n_6621, n_6622, n_6623, n_6624, n_6626;
wire n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616, n_6617;
wire n_6585, n_6586, n_6588, n_6589, n_6598, n_6599, n_6600, n_6601;
wire n_6575, n_6576, n_6577, n_6578, n_6580, n_6581, n_6583, n_6584;
wire n_6557, n_6558, n_6560, n_6561, n_6570, n_6571, n_6572, n_6573;
wire n_6548, n_6549, n_6550, n_6551, n_6552, n_6553, n_6555, n_6556;
wire n_6536, n_6537, n_6538, n_6540, n_6541, n_6544, n_6545, n_6546;
wire n_6521, n_6523, n_6524, n_6528, n_6529, n_6530, n_6532, n_6533;
wire n_6510, n_6511, n_6512, n_6513, n_6514, n_6515, n_6519, n_6520;
wire n_6495, n_6497, n_6501, n_6503, n_6504, n_6505, n_6507, n_6508;
wire n_6485, n_6486, n_6487, n_6488, n_6491, n_6492, n_6493, n_6494;
wire n_6472, n_6473, n_6474, n_6475, n_6479, n_6480, n_6482, n_6484;
wire n_6457, n_6458, n_6465, n_6466, n_6467, n_6468, n_6469, n_6471;
wire n_6448, n_6449, n_6450, n_6451, n_6452, n_6454, n_6455, n_6456;
wire n_6432, n_6433, n_6437, n_6438, n_6439, n_6440, n_6446, n_6447;
wire n_6422, n_6423, n_6424, n_6425, n_6428, n_6429, n_6430, n_6431;
wire n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232;
wire n_6217, n_6218, n_6219, n_6220, n_6221, n_6222, n_6223, n_6224;
wire n_6208, n_6209, n_6210, n_6212, n_6213, n_6214, n_6215, n_6216;
wire n_6200, n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207;
wire n_6192, n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199;
wire n_6184, n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191;
wire n_6173, n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183;
wire n_6161, n_6162, n_6163, n_6167, n_6168, n_6169, n_6171, n_6172;
wire n_6152, n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6160;
wire n_6139, n_6141, n_6142, n_6143, n_6146, n_6147, n_6148, n_6150;
wire n_6128, n_6130, n_6131, n_6132, n_6133, n_6136, n_6137, n_6138;
wire n_6117, n_6118, n_6120, n_6121, n_6122, n_6123, n_6126, n_6127;
wire n_6108, n_6109, n_6110, n_6111, n_6112, n_6114, n_6115, n_6116;
wire n_6099, n_6100, n_6102, n_6103, n_6104, n_6105, n_6106, n_6107;
wire n_6088, n_6090, n_6091, n_6092, n_6093, n_6095, n_6096, n_6097;
wire n_6079, n_6080, n_6081, n_6083, n_6084, n_6085, n_6086, n_6087;
wire n_6068, n_6069, n_6070, n_6072, n_6074, n_6075, n_6076, n_6078;
wire n_6058, n_6059, n_6060, n_6061, n_6063, n_6064, n_6066, n_6067;
wire n_6048, n_6050, n_6051, n_6052, n_6053, n_6054, n_6055, n_6057;
wire n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6046, n_6047;
wire n_6027, n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6036;
wire n_6017, n_6019, n_6020, n_6021, n_6022, n_6023, n_6024, n_6025;
wire n_6007, n_6008, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015;
wire n_5996, n_5998, n_5999, n_6000, n_6001, n_6002, n_6003, n_6004;
wire n_5987, n_5988, n_5989, n_5990, n_5991, n_5992, n_5993, n_5995;
wire n_5976, n_5977, n_5978, n_5981, n_5982, n_5983, n_5985, n_5986;
wire n_5966, n_5967, n_5968, n_5969, n_5970, n_5971, n_5973, n_5974;
wire n_5952, n_5954, n_5956, n_5959, n_5961, n_5963, n_5964, n_5965;
wire n_5941, n_5942, n_5944, n_5947, n_5948, n_5949, n_5950, n_5951;
wire n_5931, n_5933, n_5934, n_5936, n_5937, n_5938, n_5939, n_5940;
wire n_5921, n_5922, n_5924, n_5925, n_5926, n_5927, n_5928, n_5929;
wire n_5910, n_5912, n_5914, n_5915, n_5916, n_5917, n_5918, n_5919;
wire n_5894, n_5896, n_5898, n_5899, n_5901, n_5903, n_5905, n_5907;
wire n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892, n_5893;
wire n_5878, n_5879, n_5880, n_5881, n_5882, n_5883, n_5884, n_5885;
wire n_5865, n_5866, n_5867, n_5869, n_5871, n_5872, n_5873, n_5876;
wire n_5853, n_5854, n_5855, n_5856, n_5857, n_5858, n_5860, n_5862;
wire n_5843, n_5844, n_5845, n_5846, n_5847, n_5848, n_5849, n_5851;
wire n_5833, n_5834, n_5835, n_5837, n_5838, n_5840, n_5841, n_5842;
wire n_5822, n_5823, n_5824, n_5825, n_5826, n_5828, n_5830, n_5831;
wire n_5812, n_5813, n_5814, n_5815, n_5816, n_5818, n_5820, n_5821;
wire n_5801, n_5802, n_5803, n_5804, n_5806, n_5807, n_5809, n_5811;
wire n_5789, n_5790, n_5791, n_5792, n_5794, n_5796, n_5798, n_5800;
wire n_5771, n_5773, n_5774, n_5776, n_5777, n_5781, n_5784, n_5788;
wire n_5760, n_5763, n_5765, n_5766, n_5767, n_5768, n_5769, n_5770;
wire n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755, n_5759;
wire n_5737, n_5738, n_5742, n_5743, n_5744, n_5745, n_5747, n_5748;
wire n_5727, n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5735;
wire n_5716, n_5719, n_5720, n_5721, n_5722, n_5723, n_5724, n_5725;
wire n_5706, n_5707, n_5708, n_5709, n_5711, n_5712, n_5713, n_5714;
wire n_5694, n_5695, n_5699, n_5700, n_5701, n_5702, n_5703, n_5705;
wire n_5682, n_5685, n_5686, n_5687, n_5688, n_5689, n_5690, n_5693;
wire n_5667, n_5669, n_5670, n_5671, n_5672, n_5674, n_5676, n_5678;
wire n_5657, n_5658, n_5660, n_5661, n_5662, n_5664, n_5665, n_5666;
wire n_5644, n_5646, n_5648, n_5649, n_5650, n_5651, n_5652, n_5654;
wire n_5631, n_5633, n_5634, n_5637, n_5638, n_5641, n_5642, n_5643;
wire n_5621, n_5622, n_5623, n_5625, n_5627, n_5628, n_5629, n_5630;
wire n_5609, n_5610, n_5612, n_5616, n_5617, n_5618, n_5619, n_5620;
wire n_5599, n_5600, n_5601, n_5603, n_5604, n_5605, n_5606, n_5608;
wire n_5588, n_5591, n_5592, n_5594, n_5595, n_5596, n_5597, n_5598;
wire n_5569, n_5573, n_5576, n_5577, n_5578, n_5579, n_5580, n_5584;
wire n_5560, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568;
wire n_5550, n_5551, n_5553, n_5554, n_5555, n_5556, n_5557, n_5558;
wire n_5540, n_5541, n_5543, n_5545, n_5546, n_5547, n_5548, n_5549;
wire n_5530, n_5532, n_5533, n_5534, n_5535, n_5536, n_5537, n_5539;
wire n_5517, n_5518, n_5519, n_5521, n_5523, n_5525, n_5528, n_5529;
wire n_5503, n_5505, n_5507, n_5509, n_5511, n_5512, n_5513, n_5514;
wire n_5491, n_5492, n_5493, n_5494, n_5496, n_5497, n_5499, n_5500;
wire n_5481, n_5482, n_5483, n_5485, n_5486, n_5488, n_5489, n_5490;
wire n_5472, n_5473, n_5474, n_5475, n_5477, n_5478, n_5479, n_5480;
wire n_5462, n_5463, n_5464, n_5465, n_5467, n_5468, n_5469, n_5471;
wire n_5450, n_5453, n_5454, n_5456, n_5458, n_5459, n_5460, n_5461;
wire n_5437, n_5438, n_5439, n_5440, n_5442, n_5445, n_5446, n_5448;
wire n_5425, n_5426, n_5427, n_5429, n_5430, n_5432, n_5434, n_5436;
wire n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5424;
wire n_5403, n_5404, n_5407, n_5409, n_5410, n_5411, n_5413, n_5414;
wire n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5401;
wire n_5380, n_5382, n_5384, n_5385, n_5386, n_5388, n_5389, n_5390;
wire n_5366, n_5367, n_5368, n_5369, n_5370, n_5371, n_5376, n_5377;
wire n_5354, n_5355, n_5356, n_5358, n_5360, n_5361, n_5362, n_5365;
wire n_5342, n_5343, n_5345, n_5347, n_5348, n_5350, n_5352, n_5353;
wire n_5328, n_5330, n_5331, n_5333, n_5334, n_5335, n_5336, n_5338;
wire n_5316, n_5317, n_5318, n_5319, n_5320, n_5321, n_5323, n_5325;
wire n_5304, n_5305, n_5307, n_5309, n_5310, n_5311, n_5313, n_5314;
wire n_5287, n_5288, n_5289, n_5291, n_5293, n_5294, n_5297, n_5300;
wire n_5274, n_5275, n_5276, n_5278, n_5279, n_5281, n_5282, n_5285;
wire n_5263, n_5264, n_5265, n_5267, n_5269, n_5271, n_5272, n_5273;
wire n_5252, n_5253, n_5254, n_5255, n_5256, n_5257, n_5259, n_5261;
wire n_5241, n_5242, n_5243, n_5245, n_5247, n_5249, n_5250, n_5251;
wire n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240;
wire n_5222, n_5224, n_5225, n_5226, n_5227, n_5228, n_5230, n_5232;
wire n_5208, n_5210, n_5211, n_5212, n_5213, n_5214, n_5217, n_5219;
wire n_5197, n_5198, n_5199, n_5200, n_5201, n_5203, n_5204, n_5207;
wire n_5187, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5196;
wire n_5179, n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186;
wire n_5162, n_5164, n_5165, n_5166, n_5169, n_5171, n_5173, n_5177;
wire n_5153, n_5154, n_5156, n_5157, n_5158, n_5159, n_5160, n_5161;
wire n_5143, n_5144, n_5145, n_5146, n_5148, n_5149, n_5150, n_5152;
wire n_5128, n_5129, n_5132, n_5133, n_5135, n_5136, n_5139, n_5141;
wire n_5117, n_5118, n_5119, n_5121, n_5122, n_5123, n_5126, n_5127;
wire n_5107, n_5109, n_5110, n_5111, n_5112, n_5113, n_5115, n_5116;
wire n_5092, n_5095, n_5097, n_5100, n_5102, n_5104, n_5105, n_5106;
wire n_5083, n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090;
wire n_5074, n_5075, n_5076, n_5078, n_5079, n_5080, n_5081, n_5082;
wire n_5064, n_5065, n_5066, n_5067, n_5069, n_5071, n_5072, n_5073;
wire n_5053, n_5054, n_5055, n_5056, n_5059, n_5060, n_5062, n_5063;
wire n_5041, n_5042, n_5043, n_5045, n_5046, n_5047, n_5050, n_5052;
wire n_5030, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040;
wire n_5016, n_5017, n_5020, n_5022, n_5024, n_5025, n_5027, n_5028;
wire n_5003, n_5004, n_5005, n_5007, n_5009, n_5010, n_5011, n_5012;
wire n_4992, n_4994, n_4995, n_4996, n_4997, n_4998, n_4999, n_5001;
wire n_4978, n_4979, n_4980, n_4984, n_4985, n_4986, n_4988, n_4991;
wire n_4963, n_4964, n_4966, n_4968, n_4970, n_4973, n_4974, n_4976;
wire n_4954, n_4955, n_4956, n_4958, n_4959, n_4960, n_4961, n_4962;
wire n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953;
wire n_4936, n_4938, n_4939, n_4941, n_4942, n_4943, n_4944, n_4945;
wire n_4922, n_4923, n_4924, n_4925, n_4927, n_4930, n_4934, n_4935;
wire n_4912, n_4913, n_4915, n_4916, n_4917, n_4918, n_4920, n_4921;
wire n_4903, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909, n_4911;
wire n_4884, n_4887, n_4888, n_4890, n_4891, n_4893, n_4899, n_4902;
wire n_4875, n_4876, n_4877, n_4879, n_4880, n_4881, n_4882, n_4883;
wire n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4873, n_4874;
wire n_4857, n_4858, n_4859, n_4860, n_4861, n_4863, n_4864, n_4865;
wire n_4842, n_4844, n_4845, n_4848, n_4851, n_4852, n_4853, n_4854;
wire n_4833, n_4834, n_4835, n_4837, n_4838, n_4839, n_4840, n_4841;
wire n_4823, n_4824, n_4825, n_4827, n_4828, n_4829, n_4830, n_4832;
wire n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822;
wire n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814;
wire n_4798, n_4799, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806;
wire n_4790, n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797;
wire n_4779, n_4780, n_4781, n_4783, n_4784, n_4785, n_4786, n_4788;
wire n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4777, n_4778;
wire n_4759, n_4760, n_4761, n_4762, n_4765, n_4766, n_4768, n_4769;
wire n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758;
wire n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750;
wire n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742;
wire n_4725, n_4727, n_4728, n_4729, n_4730, n_4731, n_4733, n_4734;
wire n_4715, n_4716, n_4717, n_4719, n_4720, n_4721, n_4722, n_4723;
wire n_4696, n_4697, n_4698, n_4702, n_4704, n_4706, n_4711, n_4714;
wire n_4686, n_4687, n_4688, n_4689, n_4690, n_4692, n_4693, n_4695;
wire n_4678, n_4679, n_4680, n_4681, n_4682, n_4683, n_4684, n_4685;
wire n_4669, n_4670, n_4671, n_4672, n_4673, n_4674, n_4676, n_4677;
wire n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, n_4665, n_4667;
wire n_4649, n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656;
wire n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648;
wire n_4630, n_4631, n_4633, n_4634, n_4636, n_4638, n_4639, n_4640;
wire n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629;
wire n_4611, n_4613, n_4614, n_4615, n_4616, n_4617, n_4618, n_4620;
wire n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, n_4609, n_4610;
wire n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601, n_4602;
wire n_4587, n_4588, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594;
wire n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584, n_4586;
wire n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4577;
wire n_4560, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568;
wire n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559;
wire n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4551;
wire n_4535, n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542;
wire n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534;
wire n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526;
wire n_4510, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517, n_4518;
wire n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509;
wire n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501;
wire n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493;
wire n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485;
wire n_4468, n_4469, n_4471, n_4472, n_4473, n_4474, n_4476, n_4477;
wire n_4460, n_4461, n_4462, n_4463, n_4464, n_4465, n_4466, n_4467;
wire n_4451, n_4452, n_4454, n_4455, n_4456, n_4457, n_4458, n_4459;
wire n_4441, n_4442, n_4444, n_4446, n_4447, n_4448, n_4449, n_4450;
wire n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440;
wire n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432;
wire n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424;
wire n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415, n_4416;
wire n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4408;
wire n_4389, n_4390, n_4392, n_4394, n_4395, n_4396, n_4398, n_4399;
wire n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388;
wire n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380;
wire n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372;
wire n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364;
wire n_4348, n_4349, n_4350, n_4351, n_4353, n_4354, n_4355, n_4356;
wire n_4339, n_4340, n_4341, n_4342, n_4343, n_4345, n_4346, n_4347;
wire n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338;
wire n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330;
wire n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, n_4322;
wire n_4305, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313;
wire n_4295, n_4297, n_4298, n_4299, n_4301, n_4302, n_4303, n_4304;
wire n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294;
wire n_4277, n_4279, n_4280, n_4281, n_4282, n_4283, n_4285, n_4286;
wire n_4267, n_4269, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276;
wire n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266;
wire n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, n_4258;
wire n_4241, n_4243, n_4244, n_4245, n_4247, n_4248, n_4249, n_4250;
wire n_4232, n_4233, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240;
wire n_4223, n_4224, n_4225, n_4227, n_4228, n_4229, n_4230, n_4231;
wire n_4211, n_4213, n_4215, n_4218, n_4219, n_4220, n_4221, n_4222;
wire n_4201, n_4203, n_4204, n_4205, n_4207, n_4208, n_4209, n_4210;
wire n_4191, n_4192, n_4193, n_4194, n_4195, n_4197, n_4198, n_4199;
wire n_4182, n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4190;
wire n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181;
wire n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173;
wire n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165;
wire n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157;
wire n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149;
wire n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141;
wire n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133;
wire n_4116, n_4117, n_4119, n_4121, n_4122, n_4123, n_4124, n_4125;
wire n_4107, n_4108, n_4109, n_4111, n_4112, n_4113, n_4114, n_4115;
wire n_4096, n_4099, n_4100, n_4101, n_4103, n_4104, n_4105, n_4106;
wire n_4086, n_4087, n_4088, n_4090, n_4092, n_4093, n_4094, n_4095;
wire n_4076, n_4077, n_4078, n_4079, n_4080, n_4082, n_4083, n_4084;
wire n_4064, n_4066, n_4068, n_4069, n_4070, n_4071, n_4072, n_4075;
wire n_4052, n_4053, n_4055, n_4057, n_4058, n_4060, n_4061, n_4062;
wire n_4041, n_4043, n_4044, n_4045, n_4047, n_4049, n_4050, n_4051;
wire n_4029, n_4031, n_4033, n_4035, n_4037, n_4038, n_4039, n_4040;
wire n_4017, n_4018, n_4019, n_4021, n_4023, n_4025, n_4026, n_4027;
wire n_4007, n_4009, n_4011, n_4012, n_4013, n_4014, n_4015, n_4016;
wire n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, n_4005, n_4006;
wire n_3988, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996;
wire n_3977, n_3979, n_3980, n_3981, n_3982, n_3984, n_3985, n_3987;
wire n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976;
wire n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968;
wire n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960;
wire n_3942, n_3943, n_3944, n_3945, n_3947, n_3948, n_3951, n_3952;
wire n_3933, n_3934, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941;
wire n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3930, n_3932;
wire n_3913, n_3914, n_3915, n_3916, n_3917, n_3919, n_3920, n_3921;
wire n_3900, n_3901, n_3903, n_3906, n_3908, n_3910, n_3911, n_3912;
wire n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3898;
wire n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888;
wire n_3872, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880;
wire n_3859, n_3860, n_3863, n_3864, n_3865, n_3868, n_3870, n_3871;
wire n_3846, n_3848, n_3850, n_3853, n_3854, n_3855, n_3856, n_3857;
wire n_3837, n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, n_3845;
wire n_3828, n_3829, n_3830, n_3831, n_3833, n_3834, n_3835, n_3836;
wire n_3817, n_3818, n_3819, n_3821, n_3822, n_3824, n_3826, n_3827;
wire n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3815, n_3816;
wire n_3799, n_3800, n_3801, n_3802, n_3804, n_3805, n_3806, n_3807;
wire n_3786, n_3787, n_3790, n_3792, n_3793, n_3795, n_3796, n_3798;
wire n_3774, n_3775, n_3776, n_3778, n_3781, n_3782, n_3783, n_3785;
wire n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773;
wire n_3755, n_3757, n_3758, n_3759, n_3761, n_3762, n_3764, n_3765;
wire n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753;
wire n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3744;
wire n_3724, n_3726, n_3729, n_3731, n_3732, n_3733, n_3734, n_3735;
wire n_3712, n_3713, n_3714, n_3715, n_3716, n_3718, n_3719, n_3722;
wire n_3701, n_3702, n_3703, n_3707, n_3708, n_3709, n_3710, n_3711;
wire n_3690, n_3691, n_3692, n_3694, n_3695, n_3696, n_3698, n_3699;
wire n_3679, n_3681, n_3682, n_3684, n_3685, n_3686, n_3688, n_3689;
wire n_3658, n_3663, n_3664, n_3666, n_3669, n_3670, n_3676, n_3678;
wire n_3639, n_3642, n_3643, n_3647, n_3648, n_3650, n_3652, n_3653;
wire n_3620, n_3621, n_3622, n_3626, n_3628, n_3632, n_3633, n_3637;
wire n_3601, n_3604, n_3605, n_3606, n_3609, n_3612, n_3614, n_3616;
wire n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600;
wire n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3591, n_3592;
wire n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, n_3583;
wire n_3568, n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575;
wire n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567;
wire n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559;
wire n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551;
wire n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543;
wire n_3527, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535;
wire n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526;
wire n_3510, n_3511, n_3512, n_3513, n_3514, n_3516, n_3517, n_3518;
wire n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509;
wire n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501;
wire n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493;
wire n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485;
wire n_3469, n_3470, n_3471, n_3472, n_3474, n_3475, n_3476, n_3477;
wire n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468;
wire n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460;
wire n_3437, n_3439, n_3443, n_3447, n_3449, n_3450, n_3451, n_3452;
wire n_3421, n_3426, n_3428, n_3431, n_3433, n_3434, n_3435, n_3436;
wire n_3403, n_3404, n_3405, n_3408, n_3409, n_3410, n_3411, n_3414;
wire n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402;
wire n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3393, n_3394;
wire n_3375, n_3376, n_3377, n_3378, n_3379, n_3382, n_3383, n_3384;
wire n_3365, n_3366, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374;
wire n_3353, n_3356, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364;
wire n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3352;
wire n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342;
wire n_3321, n_3322, n_3323, n_3324, n_3327, n_3330, n_3333, n_3334;
wire n_3311, n_3312, n_3313, n_3314, n_3315, n_3318, n_3319, n_3320;
wire n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310;
wire n_3292, n_3293, n_3296, n_3297, n_3299, n_3300, n_3301, n_3302;
wire n_3280, n_3281, n_3282, n_3285, n_3286, n_3287, n_3290, n_3291;
wire n_3264, n_3265, n_3268, n_3269, n_3272, n_3273, n_3276, n_3278;
wire n_3254, n_3255, n_3256, n_3257, n_3260, n_3261, n_3262, n_3263;
wire n_3240, n_3241, n_3242, n_3243, n_3244, n_3249, n_3250, n_3253;
wire n_3231, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239;
wire n_3219, n_3221, n_3222, n_3223, n_3224, n_3225, n_3227, n_3230;
wire n_3210, n_3211, n_3212, n_3213, n_3215, n_3216, n_3217, n_3218;
wire n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3207, n_3208;
wire n_3190, n_3191, n_3192, n_3194, n_3195, n_3197, n_3198, n_3199;
wire n_3179, n_3180, n_3181, n_3183, n_3186, n_3187, n_3188, n_3189;
wire n_3162, n_3163, n_3167, n_3168, n_3169, n_3173, n_3177, n_3178;
wire n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158;
wire n_3138, n_3139, n_3140, n_3141, n_3142, n_3145, n_3147, n_3149;
wire n_3126, n_3127, n_3128, n_3131, n_3134, n_3135, n_3136, n_3137;
wire n_3115, n_3116, n_3117, n_3118, n_3120, n_3121, n_3123, n_3125;
wire n_3105, n_3106, n_3107, n_3108, n_3110, n_3111, n_3113, n_3114;
wire n_3095, n_3096, n_3098, n_3099, n_3101, n_3102, n_3103, n_3104;
wire n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3092, n_3093;
wire n_3072, n_3074, n_3075, n_3076, n_3077, n_3080, n_3081, n_3083;
wire n_3061, n_3062, n_3064, n_3065, n_3066, n_3068, n_3069, n_3071;
wire n_3051, n_3052, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059;
wire n_3040, n_3041, n_3043, n_3044, n_3045, n_3047, n_3048, n_3049;
wire n_3029, n_3030, n_3031, n_3032, n_3034, n_3037, n_3038, n_3039;
wire n_3020, n_3021, n_3022, n_3023, n_3024, n_3026, n_3027, n_3028;
wire n_3007, n_3009, n_3011, n_3012, n_3014, n_3015, n_3017, n_3018;
wire n_2997, n_2998, n_2999, n_3000, n_3001, n_3003, n_3004, n_3005;
wire n_2988, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996;
wire n_2978, n_2979, n_2981, n_2982, n_2984, n_2985, n_2986, n_2987;
wire n_2967, n_2968, n_2969, n_2971, n_2972, n_2974, n_2975, n_2976;
wire n_2955, n_2957, n_2958, n_2960, n_2961, n_2963, n_2965, n_2966;
wire n_2946, n_2947, n_2948, n_2949, n_2950, n_2952, n_2953, n_2954;
wire n_2937, n_2938, n_2939, n_2940, n_2941, n_2943, n_2944, n_2945;
wire n_2928, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936;
wire n_2917, n_2920, n_2921, n_2922, n_2924, n_2925, n_2926, n_2927;
wire n_2906, n_2907, n_2908, n_2909, n_2911, n_2912, n_2914, n_2916;
wire n_2893, n_2894, n_2897, n_2898, n_2900, n_2902, n_2903, n_2905;
wire n_2882, n_2883, n_2884, n_2885, n_2887, n_2888, n_2889, n_2892;
wire n_2870, n_2872, n_2873, n_2875, n_2876, n_2878, n_2879, n_2881;
wire n_2860, n_2861, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868;
wire n_2851, n_2852, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859;
wire n_2840, n_2843, n_2844, n_2846, n_2847, n_2848, n_2849, n_2850;
wire n_2830, n_2831, n_2833, n_2835, n_2836, n_2837, n_2838, n_2839;
wire n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829;
wire n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2820;
wire n_2801, n_2803, n_2805, n_2806, n_2807, n_2809, n_2810, n_2811;
wire n_2792, n_2793, n_2794, n_2795, n_2797, n_2798, n_2799, n_2800;
wire n_2783, n_2784, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791;
wire n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2780, n_2782;
wire n_2763, n_2765, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772;
wire n_2754, n_2755, n_2756, n_2757, n_2759, n_2760, n_2761, n_2762;
wire n_2742, n_2743, n_2744, n_2745, n_2746, n_2749, n_2750, n_2752;
wire n_2732, n_2733, n_2734, n_2736, n_2737, n_2738, n_2739, n_2741;
wire n_2722, n_2724, n_2725, n_2726, n_2728, n_2729, n_2730, n_2731;
wire n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721;
wire n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713;
wire n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705;
wire n_2689, n_2690, n_2691, n_2692, n_2694, n_2695, n_2696, n_2697;
wire n_2678, n_2680, n_2681, n_2682, n_2684, n_2685, n_2686, n_2687;
wire n_2668, n_2669, n_2670, n_2671, n_2673, n_2675, n_2676, n_2677;
wire n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667;
wire n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659;
wire n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651;
wire n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643;
wire n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635;
wire n_2619, n_2620, n_2621, n_2622, n_2624, n_2625, n_2626, n_2627;
wire n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618;
wire n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610;
wire n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602;
wire n_2585, n_2587, n_2588, n_2589, n_2590, n_2591, n_2593, n_2594;
wire n_2575, n_2576, n_2577, n_2579, n_2581, n_2582, n_2583, n_2584;
wire n_2566, n_2567, n_2568, n_2570, n_2571, n_2572, n_2573, n_2574;
wire n_2556, n_2557, n_2558, n_2559, n_2562, n_2563, n_2564, n_2565;
wire n_2546, n_2547, n_2548, n_2551, n_2552, n_2553, n_2554, n_2555;
wire n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545;
wire n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537;
wire n_2521, n_2522, n_2523, n_2524, n_2525, n_2527, n_2528, n_2529;
wire n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520;
wire n_2499, n_2500, n_2503, n_2504, n_2505, n_2508, n_2511, n_2512;
wire n_2487, n_2488, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498;
wire n_2472, n_2473, n_2475, n_2476, n_2477, n_2480, n_2481, n_2484;
wire n_2462, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471;
wire n_2447, n_2448, n_2452, n_2453, n_2454, n_2457, n_2458, n_2459;
wire n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446;
wire n_2424, n_2425, n_2428, n_2431, n_2433, n_2434, n_2437, n_2438;
wire n_2408, n_2409, n_2412, n_2419, n_2420, n_2421, n_2422, n_2423;
wire n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406;
wire n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398;
wire n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390;
wire n_2373, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2382;
wire n_2364, n_2365, n_2366, n_2368, n_2369, n_2370, n_2371, n_2372;
wire n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363;
wire n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2355;
wire n_2338, n_2339, n_2340, n_2341, n_2343, n_2344, n_2345, n_2346;
wire n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337;
wire n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2328, n_2329;
wire n_2311, n_2312, n_2313, n_2315, n_2316, n_2317, n_2318, n_2320;
wire n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310;
wire n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302;
wire n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293;
wire n_2277, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285;
wire n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276;
wire n_2259, n_2260, n_2261, n_2262, n_2264, n_2266, n_2267, n_2268;
wire n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258;
wire n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250;
wire n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242;
wire n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234;
wire n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226;
wire n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218;
wire n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210;
wire n_2194, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202;
wire n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193;
wire n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2185;
wire n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176;
wire n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168;
wire n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160;
wire n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152;
wire n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144;
wire n_2128, n_2129, n_2130, n_2132, n_2133, n_2134, n_2135, n_2136;
wire n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127;
wire n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119;
wire n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111;
wire n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103;
wire n_2087, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095;
wire n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086;
wire n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078;
wire n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070;
wire n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062;
wire n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054;
wire n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046;
wire n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038;
wire n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030;
wire n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022;
wire n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014;
wire n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006;
wire n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998;
wire n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990;
wire n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982;
wire n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974;
wire n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966;
wire n_1950, n_1951, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958;
wire n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949;
wire n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941;
wire n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933;
wire n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925;
wire n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917;
wire n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909;
wire n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901;
wire n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893;
wire n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885;
wire n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877;
wire n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869;
wire n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861;
wire n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853;
wire n_1837, n_1838, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845;
wire n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836;
wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
wire n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820;
wire n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812;
wire n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804;
wire n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796;
wire n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788;
wire n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780;
wire n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772;
wire n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764;
wire n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756;
wire n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748;
wire n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740;
wire n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732;
wire n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724;
wire n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716;
wire n_1698, n_1699, n_1700, n_1701, n_1702, n_1706, n_1707, n_1708;
wire n_1687, n_1688, n_1690, n_1691, n_1693, n_1694, n_1696, n_1697;
wire n_1676, n_1677, n_1678, n_1679, n_1681, n_1682, n_1684, n_1685;
wire n_1666, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1675;
wire n_1656, n_1658, n_1659, n_1660, n_1661, n_1662, n_1664, n_1665;
wire n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1654, n_1655;
wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1644, n_1645, n_1646;
wire n_1628, n_1629, n_1631, n_1632, n_1633, n_1635, n_1636, n_1637;
wire n_1619, n_1620, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627;
wire n_1609, n_1611, n_1612, n_1613, n_1614, n_1615, n_1617, n_1618;
wire n_1600, n_1601, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608;
wire n_1591, n_1592, n_1593, n_1594, n_1595, n_1597, n_1598, n_1599;
wire n_1581, n_1582, n_1583, n_1584, n_1585, n_1587, n_1588, n_1590;
wire n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1579, n_1580;
wire n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1570, n_1571;
wire n_1553, n_1554, n_1555, n_1557, n_1558, n_1559, n_1560, n_1561;
wire n_1544, n_1545, n_1546, n_1547, n_1548, n_1550, n_1551, n_1552;
wire n_1534, n_1535, n_1536, n_1537, n_1539, n_1540, n_1541, n_1542;
wire n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1533;
wire n_1516, n_1517, n_1518, n_1519, n_1521, n_1522, n_1523, n_1524;
wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
wire n_1498, n_1499, n_1500, n_1502, n_1503, n_1504, n_1506, n_1507;
wire n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
wire n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489;
wire n_1472, n_1473, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481;
wire n_1459, n_1460, n_1461, n_1462, n_1464, n_1465, n_1470, n_1471;
wire n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1456, n_1458;
wire n_1440, n_1441, n_1442, n_1443, n_1444, n_1446, n_1447, n_1448;
wire n_1430, n_1431, n_1432, n_1433, n_1435, n_1436, n_1437, n_1438;
wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429;
wire n_1413, n_1414, n_1415, n_1417, n_1418, n_1419, n_1420, n_1421;
wire n_1403, n_1404, n_1405, n_1407, n_1409, n_1410, n_1411, n_1412;
wire n_1391, n_1393, n_1395, n_1396, n_1398, n_1399, n_1400, n_1402;
wire n_1381, n_1382, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
wire n_1372, n_1373, n_1374, n_1375, n_1377, n_1378, n_1379, n_1380;
wire n_1362, n_1364, n_1365, n_1366, n_1367, n_1369, n_1370, n_1371;
wire n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360;
wire n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352;
wire n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1344;
wire n_1327, n_1328, n_1329, n_1330, n_1332, n_1333, n_1334, n_1335;
wire n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326;
wire n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318;
wire n_1294, n_1297, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310;
wire n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291;
wire n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283;
wire n_1262, n_1263, n_1264, n_1265, n_1267, n_1268, n_1272, n_1275;
wire n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261;
wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253;
wire n_1237, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
wire n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236;
wire n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228;
wire n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220;
wire n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212;
wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204;
wire n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196;
wire n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188;
wire n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180;
wire n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172;
wire n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164;
wire n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156;
wire n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148;
wire n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140;
wire n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132;
wire n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124;
wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116;
wire n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108;
wire n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100;
wire n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092;
wire n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084;
wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
wire n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068;
wire n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060;
wire n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052;
wire n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044;
wire n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036;
wire n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028;
wire n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020;
wire n_1003, n_1004, n_1005, n_1006, n_1007, n_1009, n_1011, n_1012;
wire n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002;
wire n_986, n_987, n_988, n_990, n_991, n_992, n_993, n_994;
wire n_977, n_979, n_980, n_981, n_982, n_983, n_984, n_985;
wire n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976;
wire n_959, n_960, n_962, n_963, n_964, n_965, n_966, n_967;
wire n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958;
wire n_942, n_943, n_944, n_945, n_947, n_948, n_949, n_950;
wire n_932, n_933, n_935, n_937, n_938, n_939, n_940, n_941;
wire n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931;
wire n_915, n_916, n_918, n_919, n_920, n_921, n_922, n_923;
wire n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914;
wire n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906;
wire n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898;
wire n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890;
wire n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882;
wire n_858, n_860, n_866, n_867, n_868, n_869, n_873, n_874;
wire n_846, n_847, n_848, n_849, n_850, n_852, n_853, n_857;
wire n_815, n_816, n_817, n_823, n_830, n_831, n_836, n_842;
wire n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814;
wire n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806;
wire n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798;
wire n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790;
wire n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782;
wire n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774;
wire n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766;
wire n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758;
wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
wire n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742;
wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734;
wire n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726;
wire n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718;
wire n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
wire n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702;
wire n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
wire n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685;
wire n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677;
wire n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669;
wire n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661;
wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
wire n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645;
wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
wire n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621;
wire n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613;
wire n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605;
wire n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597;
wire n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589;
wire n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581;
wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
wire n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549;
wire n_532, n_535, n_536, n_537, n_538, n_539, n_540, n_541;
wire n_523, n_524, n_525, n_526, n_527, n_529, n_530, n_531;
wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_514;
wire n_495, n_496, n_497, n_499, n_500, n_501, n_502, n_503;
wire n_482, n_484, n_486, n_488, n_489, n_490, n_491, n_492;
wire n_471, n_472, n_473, n_474, n_476, n_478, n_479, n_480;
wire n_462, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
wire n_451, n_453, n_454, n_456, n_457, n_458, n_460, n_461;
wire n_436, n_438, n_440, n_442, n_443, n_447, n_448, n_450;
wire n_424, n_426, n_427, n_428, n_429, n_431, n_433, n_434;
wire n_415, n_416, n_417, n_418, n_419, n_420, n_422, n_423;
wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
wire n_398, n_399, n_401, n_402, n_403, n_404, n_405, n_406;
wire n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397;
wire n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389;
wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381;
wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
wire n_349, n_350, n_351, n_352, n_353, n_354, n_356, n_357;
wire n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348;
wire n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340;
wire n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332;
wire n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324;
wire n_308, n_310, n_311, n_312, n_313, n_314, n_315, n_316;
wire n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307;
wire n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299;
wire n_283, n_285, n_286, n_287, n_288, n_289, n_290, n_291;
wire n_266, n_268, n_271, n_273, n_276, n_278, n_280, n_282;
wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_264;
wire n_233, n_235, n_236, n_241, n_244, n_247, n_252, n_254;
wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_219;
wire n_198, n_199, n_200, n_201, n_204, n_205, n_206, n_207;
wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_197;
wire n_180, n_181, n_183, n_184, n_185, n_186, n_187, n_188;
wire n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179;
wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
wire n_139, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
wire n_127, n_129, n_130, n_131, n_133, n_135, n_136, n_137;
wire n_112, n_113, n_117, n_118, n_119, n_120, n_124, n_126;
wire n_100, n_101, n_104, n_105, n_106, n_108, n_109, n_111;
wire n_81, n_83, n_85, n_87, n_89, n_95, n_96, n_98;
wire n_65, n_67, n_68, n_69, n_70, n_71, n_73, n_79;
wire n_46, n_48, n_49, n_51, n_52, n_56, n_58, n_63;
wire n_33, n_35, n_36, n_38, n_40, n_41, n_43, n_44;
wire n_18, n_19, n_20, n_21, n_24, n_27, n_28, n_32;
wire n_0, n_2, n_3, n_4, n_5, n_12, n_14, n_16;
wire _2357_, _2358_, _2359_, _2360_, _2361_, _2362_, _2363_, _2364_;
wire _2349_, _2350_, _2351_, _2352_, _2353_, _2354_, _2355_, _2356_;
wire _2341_, _2342_, _2343_, _2344_, _2345_, _2346_, _2347_, _2348_;
wire _2333_, _2334_, _2335_, _2336_, _2337_, _2338_, _2339_, _2340_;
wire _2325_, _2326_, _2327_, _2328_, _2329_, _2330_, _2331_, _2332_;
wire _2317_, _2318_, _2319_, _2320_, _2321_, _2322_, _2323_, _2324_;
wire _2309_, _2310_, _2311_, _2312_, _2313_, _2314_, _2315_, _2316_;
wire _2301_, _2302_, _2303_, _2304_, _2305_, _2306_, _2307_, _2308_;
wire _2293_, _2294_, _2295_, _2296_, _2297_, _2298_, _2299_, _2300_;
wire _2285_, _2286_, _2287_, _2288_, _2289_, _2290_, _2291_, _2292_;
wire _2277_, _2278_, _2279_, _2280_, _2281_, _2282_, _2283_, _2284_;
wire _2269_, _2270_, _2271_, _2272_, _2273_, _2274_, _2275_, _2276_;
wire _2261_, _2262_, _2263_, _2264_, _2265_, _2266_, _2267_, _2268_;
wire _2253_, _2254_, _2255_, _2256_, _2257_, _2258_, _2259_, _2260_;
wire _2245_, _2246_, _2247_, _2248_, _2249_, _2250_, _2251_, _2252_;
wire _2237_, _2238_, _2239_, _2240_, _2241_, _2242_, _2243_, _2244_;
wire _2229_, _2230_, _2231_, _2232_, _2233_, _2234_, _2235_, _2236_;
wire _2221_, _2222_, _2223_, _2224_, _2225_, _2226_, _2227_, _2228_;
wire _2213_, _2214_, _2215_, _2216_, _2217_, _2218_, _2219_, _2220_;
wire _2205_, _2206_, _2207_, _2208_, _2209_, _2210_, _2211_, _2212_;
wire _2197_, _2198_, _2199_, _2200_, _2201_, _2202_, _2203_, _2204_;
wire _2189_, _2190_, _2191_, _2192_, _2193_, _2194_, _2195_, _2196_;
wire _2181_, _2182_, _2183_, _2184_, _2185_, _2186_, _2187_, _2188_;
wire _2173_, _2174_, _2175_, _2176_, _2177_, _2178_, _2179_, _2180_;
wire _2165_, _2166_, _2167_, _2168_, _2169_, _2170_, _2171_, _2172_;
wire _2157_, _2158_, _2159_, _2160_, _2161_, _2162_, _2163_, _2164_;
wire _2149_, _2150_, _2151_, _2152_, _2153_, _2154_, _2155_, _2156_;
wire _2141_, _2142_, _2143_, _2144_, _2145_, _2146_, _2147_, _2148_;
wire _2133_, _2134_, _2135_, _2136_, _2137_, _2138_, _2139_, _2140_;
wire _2125_, _2126_, _2127_, _2128_, _2129_, _2130_, _2131_, _2132_;
wire _2117_, _2118_, _2119_, _2120_, _2121_, _2122_, _2123_, _2124_;
wire _2109_, _2110_, _2111_, _2112_, _2113_, _2114_, _2115_, _2116_;
wire _2101_, _2102_, _2103_, _2104_, _2105_, _2106_, _2107_, _2108_;
wire _2093_, _2094_, _2095_, _2096_, _2097_, _2098_, _2099_, _2100_;
wire _2085_, _2086_, _2087_, _2088_, _2089_, _2090_, _2091_, _2092_;
wire _2077_, _2078_, _2079_, _2080_, _2081_, _2082_, _2083_, _2084_;
wire WX11229, WX11231, WX11233, WX11235, WX11237, WX11239, WX11241, WX11243;
wire WX11213, WX11215, WX11217, WX11219, WX11221, WX11223, WX11225, WX11227;
wire WX11197, WX11199, WX11201, WX11203, WX11205, WX11207, WX11209, WX11211;
wire WX11181, WX11183, WX11185, WX11187, WX11189, WX11191, WX11193, WX11195;
wire WX11165, WX11167, WX11169, WX11171, WX11173, WX11175, WX11177, WX11179;
wire WX11149, WX11151, WX11153, WX11155, WX11157, WX11159, WX11161, WX11163;
wire WX11133, WX11135, WX11137, WX11139, WX11141, WX11143, WX11145, WX11147;
wire WX11117, WX11119, WX11121, WX11123, WX11125, WX11127, WX11129, WX11131;
wire WX11101, WX11103, WX11105, WX11107, WX11109, WX11111, WX11113, WX11115;
wire WX11085, WX11087, WX11089, WX11091, WX11093, WX11095, WX11097, WX11099;
wire WX11069, WX11071, WX11073, WX11075, WX11077, WX11079, WX11081, WX11083;
wire WX11053, WX11055, WX11057, WX11059, WX11061, WX11063, WX11065, WX11067;
wire WX11037, WX11039, WX11041, WX11043, WX11045, WX11047, WX11049, WX11051;
wire WX11021, WX11023, WX11025, WX11027, WX11029, WX11031, WX11033, WX11035;
wire WX11005, WX11007, WX11009, WX11011, WX11013, WX11015, WX11017, WX11019;
wire WX10989, WX10991, WX10993, WX10995, WX10997, WX10999, WX11001, WX11003;
wire WX10877, WX10879, WX10881, WX10883, WX10885, WX10887, WX10889, WX10891;
wire WX10861, WX10863, WX10865, WX10867, WX10869, WX10871, WX10873, WX10875;
wire WX10845, WX10847, WX10849, WX10851, WX10853, WX10855, WX10857, WX10859;
wire WX10829, WX10831, WX10833, WX10835, WX10837, WX10839, WX10841, WX10843;
wire WX9936, WX9938, WX9940, WX9942, WX9944, WX9946, WX9948, WX9950;
wire WX9920, WX9922, WX9924, WX9926, WX9928, WX9930, WX9932, WX9934;
wire WX9904, WX9906, WX9908, WX9910, WX9912, WX9914, WX9916, WX9918;
wire WX9888, WX9890, WX9892, WX9894, WX9896, WX9898, WX9900, WX9902;
wire WX9872, WX9874, WX9876, WX9878, WX9880, WX9882, WX9884, WX9886;
wire WX9856, WX9858, WX9860, WX9862, WX9864, WX9866, WX9868, WX9870;
wire WX9840, WX9842, WX9844, WX9846, WX9848, WX9850, WX9852, WX9854;
wire WX9824, WX9826, WX9828, WX9830, WX9832, WX9834, WX9836, WX9838;
wire WX9808, WX9810, WX9812, WX9814, WX9816, WX9818, WX9820, WX9822;
wire WX9792, WX9794, WX9796, WX9798, WX9800, WX9802, WX9804, WX9806;
wire WX9776, WX9778, WX9780, WX9782, WX9784, WX9786, WX9788, WX9790;
wire WX9760, WX9762, WX9764, WX9766, WX9768, WX9770, WX9772, WX9774;
wire WX9744, WX9746, WX9748, WX9750, WX9752, WX9754, WX9756, WX9758;
wire WX9728, WX9730, WX9732, WX9734, WX9736, WX9738, WX9740, WX9742;
wire WX9712, WX9714, WX9716, WX9718, WX9720, WX9722, WX9724, WX9726;
wire WX9696, WX9698, WX9700, WX9702, WX9704, WX9706, WX9708, WX9710;
wire WX9584, WX9586, WX9588, WX9590, WX9592, WX9594, WX9596, WX9598;
wire WX9568, WX9570, WX9572, WX9574, WX9576, WX9578, WX9580, WX9582;
wire WX9552, WX9554, WX9556, WX9558, WX9560, WX9562, WX9564, WX9566;
wire WX9536, WX9538, WX9540, WX9542, WX9544, WX9546, WX9548, WX9550;
wire WX8643, WX8645, WX8647, WX8649, WX8651, WX8653, WX8655, WX8657;
wire WX8627, WX8629, WX8631, WX8633, WX8635, WX8637, WX8639, WX8641;
wire WX8611, WX8613, WX8615, WX8617, WX8619, WX8621, WX8623, WX8625;
wire WX8595, WX8597, WX8599, WX8601, WX8603, WX8605, WX8607, WX8609;
wire WX8579, WX8581, WX8583, WX8585, WX8587, WX8589, WX8591, WX8593;
wire WX8563, WX8565, WX8567, WX8569, WX8571, WX8573, WX8575, WX8577;
wire WX8547, WX8549, WX8551, WX8553, WX8555, WX8557, WX8559, WX8561;
wire WX8531, WX8533, WX8535, WX8537, WX8539, WX8541, WX8543, WX8545;
wire WX8515, WX8517, WX8519, WX8521, WX8523, WX8525, WX8527, WX8529;
wire WX8499, WX8501, WX8503, WX8505, WX8507, WX8509, WX8511, WX8513;
wire WX8483, WX8485, WX8487, WX8489, WX8491, WX8493, WX8495, WX8497;
wire WX8467, WX8469, WX8471, WX8473, WX8475, WX8477, WX8479, WX8481;
wire WX8451, WX8453, WX8455, WX8457, WX8459, WX8461, WX8463, WX8465;
wire WX8435, WX8437, WX8439, WX8441, WX8443, WX8445, WX8447, WX8449;
wire WX8419, WX8421, WX8423, WX8425, WX8427, WX8429, WX8431, WX8433;
wire WX8403, WX8405, WX8407, WX8409, WX8411, WX8413, WX8415, WX8417;
wire WX8291, WX8293, WX8295, WX8297, WX8299, WX8301, WX8303, WX8305;
wire WX8275, WX8277, WX8279, WX8281, WX8283, WX8285, WX8287, WX8289;
wire WX8259, WX8261, WX8263, WX8265, WX8267, WX8269, WX8271, WX8273;
wire WX8243, WX8245, WX8247, WX8249, WX8251, WX8253, WX8255, WX8257;
wire WX7350, WX7352, WX7354, WX7356, WX7358, WX7360, WX7362, WX7364;
wire WX7334, WX7336, WX7338, WX7340, WX7342, WX7344, WX7346, WX7348;
wire WX7318, WX7320, WX7322, WX7324, WX7326, WX7328, WX7330, WX7332;
wire WX7302, WX7304, WX7306, WX7308, WX7310, WX7312, WX7314, WX7316;
wire WX7286, WX7288, WX7290, WX7292, WX7294, WX7296, WX7298, WX7300;
wire WX7270, WX7272, WX7274, WX7276, WX7278, WX7280, WX7282, WX7284;
wire WX7254, WX7256, WX7258, WX7260, WX7262, WX7264, WX7266, WX7268;
wire WX7238, WX7240, WX7242, WX7244, WX7246, WX7248, WX7250, WX7252;
wire WX7222, WX7224, WX7226, WX7228, WX7230, WX7232, WX7234, WX7236;
wire WX7206, WX7208, WX7210, WX7212, WX7214, WX7216, WX7218, WX7220;
wire WX7190, WX7192, WX7194, WX7196, WX7198, WX7200, WX7202, WX7204;
wire WX7174, WX7176, WX7178, WX7180, WX7182, WX7184, WX7186, WX7188;
wire WX7158, WX7160, WX7162, WX7164, WX7166, WX7168, WX7170, WX7172;
wire WX7142, WX7144, WX7146, WX7148, WX7150, WX7152, WX7154, WX7156;
wire WX7126, WX7128, WX7130, WX7132, WX7134, WX7136, WX7138, WX7140;
wire WX7110, WX7112, WX7114, WX7116, WX7118, WX7120, WX7122, WX7124;
wire WX6998, WX7000, WX7002, WX7004, WX7006, WX7008, WX7010, WX7012;
wire WX6982, WX6984, WX6986, WX6988, WX6990, WX6992, WX6994, WX6996;
wire WX6966, WX6968, WX6970, WX6972, WX6974, WX6976, WX6978, WX6980;
wire WX6950, WX6952, WX6954, WX6956, WX6958, WX6960, WX6962, WX6964;
wire WX6057, WX6059, WX6061, WX6063, WX6065, WX6067, WX6069, WX6071;
wire WX6041, WX6043, WX6045, WX6047, WX6049, WX6051, WX6053, WX6055;
wire WX6025, WX6027, WX6029, WX6031, WX6033, WX6035, WX6037, WX6039;
wire WX6009, WX6011, WX6013, WX6015, WX6017, WX6019, WX6021, WX6023;
wire WX5993, WX5995, WX5997, WX5999, WX6001, WX6003, WX6005, WX6007;
wire WX5977, WX5979, WX5981, WX5983, WX5985, WX5987, WX5989, WX5991;
wire WX5961, WX5963, WX5965, WX5967, WX5969, WX5971, WX5973, WX5975;
wire WX5945, WX5947, WX5949, WX5951, WX5953, WX5955, WX5957, WX5959;
wire WX5929, WX5931, WX5933, WX5935, WX5937, WX5939, WX5941, WX5943;
wire WX5913, WX5915, WX5917, WX5919, WX5921, WX5923, WX5925, WX5927;
wire WX5897, WX5899, WX5901, WX5903, WX5905, WX5907, WX5909, WX5911;
wire WX5881, WX5883, WX5885, WX5887, WX5889, WX5891, WX5893, WX5895;
wire WX5865, WX5867, WX5869, WX5871, WX5873, WX5875, WX5877, WX5879;
wire WX5849, WX5851, WX5853, WX5855, WX5857, WX5859, WX5861, WX5863;
wire WX5833, WX5835, WX5837, WX5839, WX5841, WX5843, WX5845, WX5847;
wire WX5817, WX5819, WX5821, WX5823, WX5825, WX5827, WX5829, WX5831;
wire WX5705, WX5707, WX5709, WX5711, WX5713, WX5715, WX5717, WX5719;
wire WX5689, WX5691, WX5693, WX5695, WX5697, WX5699, WX5701, WX5703;
wire WX5673, WX5675, WX5677, WX5679, WX5681, WX5683, WX5685, WX5687;
wire WX5657, WX5659, WX5661, WX5663, WX5665, WX5667, WX5669, WX5671;
wire WX4764, WX4766, WX4768, WX4770, WX4772, WX4774, WX4776, WX4778;
wire WX4748, WX4750, WX4752, WX4754, WX4756, WX4758, WX4760, WX4762;
wire WX4732, WX4734, WX4736, WX4738, WX4740, WX4742, WX4744, WX4746;
wire WX4716, WX4718, WX4720, WX4722, WX4724, WX4726, WX4728, WX4730;
wire WX4700, WX4702, WX4704, WX4706, WX4708, WX4710, WX4712, WX4714;
wire WX4684, WX4686, WX4688, WX4690, WX4692, WX4694, WX4696, WX4698;
wire WX4668, WX4670, WX4672, WX4674, WX4676, WX4678, WX4680, WX4682;
wire WX4652, WX4654, WX4656, WX4658, WX4660, WX4662, WX4664, WX4666;
wire WX4636, WX4638, WX4640, WX4642, WX4644, WX4646, WX4648, WX4650;
wire WX4620, WX4622, WX4624, WX4626, WX4628, WX4630, WX4632, WX4634;
wire WX4604, WX4606, WX4608, WX4610, WX4612, WX4614, WX4616, WX4618;
wire WX4588, WX4590, WX4592, WX4594, WX4596, WX4598, WX4600, WX4602;
wire WX4572, WX4574, WX4576, WX4578, WX4580, WX4582, WX4584, WX4586;
wire WX4556, WX4558, WX4560, WX4562, WX4564, WX4566, WX4568, WX4570;
wire WX4540, WX4542, WX4544, WX4546, WX4548, WX4550, WX4552, WX4554;
wire WX4524, WX4526, WX4528, WX4530, WX4532, WX4534, WX4536, WX4538;
wire WX4412, WX4414, WX4416, WX4418, WX4420, WX4422, WX4424, WX4426;
wire WX4396, WX4398, WX4400, WX4402, WX4404, WX4406, WX4408, WX4410;
wire WX4380, WX4382, WX4384, WX4386, WX4388, WX4390, WX4392, WX4394;
wire WX4364, WX4366, WX4368, WX4370, WX4372, WX4374, WX4376, WX4378;
wire WX3471, WX3473, WX3475, WX3477, WX3479, WX3481, WX3483, WX3485;
wire WX3455, WX3457, WX3459, WX3461, WX3463, WX3465, WX3467, WX3469;
wire WX3439, WX3441, WX3443, WX3445, WX3447, WX3449, WX3451, WX3453;
wire WX3423, WX3425, WX3427, WX3429, WX3431, WX3433, WX3435, WX3437;
wire WX3407, WX3409, WX3411, WX3413, WX3415, WX3417, WX3419, WX3421;
wire WX3391, WX3393, WX3395, WX3397, WX3399, WX3401, WX3403, WX3405;
wire WX3375, WX3377, WX3379, WX3381, WX3383, WX3385, WX3387, WX3389;
wire WX3359, WX3361, WX3363, WX3365, WX3367, WX3369, WX3371, WX3373;
wire WX3343, WX3345, WX3347, WX3349, WX3351, WX3353, WX3355, WX3357;
wire WX3327, WX3329, WX3331, WX3333, WX3335, WX3337, WX3339, WX3341;
wire WX3311, WX3313, WX3315, WX3317, WX3319, WX3321, WX3323, WX3325;
wire WX3295, WX3297, WX3299, WX3301, WX3303, WX3305, WX3307, WX3309;
wire WX3279, WX3281, WX3283, WX3285, WX3287, WX3289, WX3291, WX3293;
wire WX3263, WX3265, WX3267, WX3269, WX3271, WX3273, WX3275, WX3277;
wire WX3247, WX3249, WX3251, WX3253, WX3255, WX3257, WX3259, WX3261;
wire WX3231, WX3233, WX3235, WX3237, WX3239, WX3241, WX3243, WX3245;
wire WX3119, WX3121, WX3123, WX3125, WX3127, WX3129, WX3131, WX3133;
wire WX3103, WX3105, WX3107, WX3109, WX3111, WX3113, WX3115, WX3117;
wire WX3087, WX3089, WX3091, WX3093, WX3095, WX3097, WX3099, WX3101;
wire WX3071, WX3073, WX3075, WX3077, WX3079, WX3081, WX3083, WX3085;
wire WX2178, WX2180, WX2182, WX2184, WX2186, WX2188, WX2190, WX2192;
wire WX2162, WX2164, WX2166, WX2168, WX2170, WX2172, WX2174, WX2176;
wire WX2146, WX2148, WX2150, WX2152, WX2154, WX2156, WX2158, WX2160;
wire WX2130, WX2132, WX2134, WX2136, WX2138, WX2140, WX2142, WX2144;
wire WX2114, WX2116, WX2118, WX2120, WX2122, WX2124, WX2126, WX2128;
wire WX2098, WX2100, WX2102, WX2104, WX2106, WX2108, WX2110, WX2112;
wire WX2082, WX2084, WX2086, WX2088, WX2090, WX2092, WX2094, WX2096;
wire WX2066, WX2068, WX2070, WX2072, WX2074, WX2076, WX2078, WX2080;
wire WX2050, WX2052, WX2054, WX2056, WX2058, WX2060, WX2062, WX2064;
wire WX2034, WX2036, WX2038, WX2040, WX2042, WX2044, WX2046, WX2048;
wire WX2018, WX2020, WX2022, WX2024, WX2026, WX2028, WX2030, WX2032;
wire WX2002, WX2004, WX2006, WX2008, WX2010, WX2012, WX2014, WX2016;
wire WX1986, WX1988, WX1990, WX1992, WX1994, WX1996, WX1998, WX2000;
wire WX1970, WX1972, WX1974, WX1976, WX1978, WX1980, WX1982, WX1984;
wire WX1954, WX1956, WX1958, WX1960, WX1962, WX1964, WX1966, WX1968;
wire WX1938, WX1940, WX1942, WX1944, WX1946, WX1948, WX1950, WX1952;
wire WX1826, WX1828, WX1830, WX1832, WX1834, WX1836, WX1838, WX1840;
wire WX1810, WX1812, WX1814, WX1816, WX1818, WX1820, WX1822, WX1824;
wire WX1794, WX1796, WX1798, WX1800, WX1802, WX1804, WX1806, WX1808;
wire WX1778, WX1780, WX1782, WX1784, WX1786, WX1788, WX1790, WX1792;
wire WX885, WX887, WX889, WX891, WX893, WX895, WX897, WX899;
wire WX869, WX871, WX873, WX875, WX877, WX879, WX881, WX883;
wire WX853, WX855, WX857, WX859, WX861, WX863, WX865, WX867;
wire WX837, WX839, WX841, WX843, WX845, WX847, WX849, WX851;
wire WX821, WX823, WX825, WX827, WX829, WX831, WX833, WX835;
wire WX805, WX807, WX809, WX811, WX813, WX815, WX817, WX819;
wire WX789, WX791, WX793, WX795, WX797, WX799, WX801, WX803;
wire WX773, WX775, WX777, WX779, WX781, WX783, WX785, WX787;
wire WX757, WX759, WX761, WX763, WX765, WX767, WX769, WX771;
wire WX741, WX743, WX745, WX747, WX749, WX751, WX753, WX755;
wire WX725, WX727, WX729, WX731, WX733, WX735, WX737, WX739;
wire WX709, WX711, WX713, WX715, WX717, WX719, WX721, WX723;
wire WX693, WX695, WX697, WX699, WX701, WX703, WX705, WX707;
wire WX677, WX679, WX681, WX683, WX685, WX687, WX689, WX691;
wire WX661, WX663, WX665, WX667, WX669, WX671, WX673, WX675;
wire WX645, WX647, WX649, WX651, WX653, WX655, WX657, WX659;
wire WX533, WX535, WX537, WX539, WX541, WX543, WX545, WX547;
wire WX517, WX519, WX521, WX523, WX525, WX527, WX529, WX531;
wire WX501, WX503, WX505, WX507, WX509, WX511, WX513, WX515;
wire WX485, WX487, WX489, WX491, WX493, WX495, WX497, WX499;
wire DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27, DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22, DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17, DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12, DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7, DATA_9_6, DATA_9_5, DATA_9_4, DATA_9_3, DATA_9_2, DATA_9_1, DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2, CRC_OUT_9_3, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30, CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2, CRC_OUT_7_3, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2, CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2, CRC_OUT_2_3, CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_2, CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31;
wire blif_clk_net, blif_reset_net, DATA_0_31, DATA_0_30, DATA_0_29, DATA_0_28, DATA_0_27, DATA_0_26, DATA_0_25, DATA_0_24, DATA_0_23, DATA_0_22, DATA_0_21, DATA_0_20, DATA_0_19, DATA_0_18, DATA_0_17, DATA_0_16, DATA_0_15, DATA_0_14, DATA_0_13, DATA_0_12, DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8, DATA_0_7, DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2, DATA_0_1, DATA_0_0, RESET, TM1, TM0;
CLKBUFX1 gbuf_d_1(.A(n_6173), .Y(d_out_1));
CLKBUFX1 gbuf_q_1(.A(q_in_1), .Y(WX651));
NAND2X2 g55802(.A (n_6172), .B (n_4727), .Y (n_6173));
NAND2X1 g55823(.A (n_6615), .B (n_8328), .Y (n_6172));
CLKBUFX1 gbuf_d_2(.A(n_6169), .Y(d_out_2));
CLKBUFX1 gbuf_q_2(.A(q_in_2), .Y(WX653));
OAI21X1 g55843(.A0 (n_6167), .A1 (n_5889), .B0 (n_6156), .Y (n_8328));
NAND2X2 g55841(.A (n_6168), .B (n_4725), .Y (n_6169));
NAND2X1 g55878(.A (n_6555), .B (n_8329), .Y (n_6168));
INVX1 g55905(.A (DATA_9_28), .Y (n_6167));
CLKBUFX1 gbuf_d_3(.A(n_6163), .Y(d_out_3));
CLKBUFX1 gbuf_q_3(.A(q_in_3), .Y(WX655));
OAI21X1 g55906(.A0 (n_6162), .A1 (n_5242), .B0 (n_4070), .Y(DATA_9_28));
OAI21X1 g55903(.A0 (n_6160), .A1 (n_5889), .B0 (n_6146), .Y (n_8329));
NAND2X2 g55901(.A (n_6161), .B (n_4723), .Y (n_6163));
CLKBUFX1 gbuf_d_4(.A(n_6158), .Y(d_out_4));
CLKBUFX1 gbuf_q_4(.A(q_in_4), .Y(WX489));
MX2X1 g55963(.A (n_6157), .B (WX491), .S0 (n_4069), .Y (n_6162));
NAND2X1 g55938(.A (n_6155), .B (n_6583), .Y (n_6161));
INVX1 g55964(.A (DATA_9_27), .Y (n_6160));
NOR2X1 g55992(.A (n_1425), .B (n_6157), .Y (n_6158));
OR2X1 g55996(.A (n_6157), .B (n_5990), .Y (n_6156));
OAI21X1 g55965(.A0 (n_6153), .A1 (n_6091), .B0 (n_4041), .Y(DATA_9_27));
CLKBUFX1 gbuf_d_5(.A(n_6154), .Y(d_out_5));
CLKBUFX1 gbuf_q_5(.A(q_in_5), .Y(WX657));
OAI21X1 g55962(.A0 (n_6150), .A1 (n_5889), .B0 (n_6137), .Y (n_6155));
INVX1 g56007(.A (WX491), .Y (n_6157));
NAND2X2 g55960(.A (n_6152), .B (n_4722), .Y (n_6154));
CLKBUFX1 gbuf_d_6(.A(n_6148), .Y(d_out_6));
CLKBUFX1 gbuf_q_6(.A(q_in_6), .Y(WX491));
MX2X1 g56022(.A (n_6147), .B (WX493), .S0 (n_4040), .Y (n_6153));
NAND2X2 g55997(.A (n_6583), .B (n_6882), .Y (n_6152));
INVX1 g56023(.A (DATA_9_26), .Y (n_6150));
NOR2X1 g56051(.A (n_1425), .B (n_6147), .Y (n_6148));
OR2X1 g56055(.A (n_6147), .B (n_5968), .Y (n_6146));
OAI21X1 g56024(.A0 (n_6142), .A1 (n_5242), .B0 (n_4023), .Y(DATA_9_26));
CLKBUFX1 gbuf_d_7(.A(n_6143), .Y(d_out_7));
CLKBUFX1 gbuf_q_7(.A(q_in_7), .Y(WX659));
INVX1 g56068(.A (WX493), .Y (n_6147));
OAI21X1 g56021(.A0 (n_6141), .A1 (n_5889), .B0 (n_6126), .Y (n_6882));
CLKBUFX1 gbuf_d_8(.A(n_6139), .Y(d_out_8));
CLKBUFX1 gbuf_q_8(.A(q_in_8), .Y(WX493));
NAND2X1 g56019(.A (n_6136), .B (n_4721), .Y (n_6143));
MX2X1 g56081(.A (n_6138), .B (WX495), .S0 (n_7066), .Y (n_6142));
INVX1 g56082(.A (DATA_9_25), .Y (n_6141));
NOR2X1 g56110(.A (n_5181), .B (n_6138), .Y (n_6139));
OR2X1 g56114(.A (n_6138), .B (n_5990), .Y (n_6137));
NAND2X1 g56056(.A (n_6555), .B (n_8330), .Y (n_6136));
OAI21X1 g56083(.A0 (n_6132), .A1 (n_6091), .B0 (n_4072), .Y(DATA_9_25));
CLKBUFX1 gbuf_d_9(.A(n_6133), .Y(d_out_9));
CLKBUFX1 gbuf_q_9(.A(q_in_9), .Y(WX661));
OAI21X1 g56080(.A0 (n_6130), .A1 (n_5889), .B0 (n_6116), .Y (n_8330));
INVX1 g56123(.A (WX495), .Y (n_6138));
NAND2X1 g56078(.A (n_6131), .B (n_4720), .Y (n_6133));
CLKBUFX1 gbuf_d_10(.A(n_6128), .Y(d_out_10));
CLKBUFX1 gbuf_q_10(.A(q_in_10), .Y(WX495));
MX2X1 g56140(.A (n_6127), .B (WX497), .S0 (n_4071), .Y (n_6132));
NAND2X1 g56115(.A (n_6583), .B (n_6883), .Y (n_6131));
INVX1 g56141(.A (DATA_9_24), .Y (n_6130));
NOR2X1 g56169(.A (n_5181), .B (n_6127), .Y (n_6128));
OR2X1 g56173(.A (n_6127), .B (n_5990), .Y (n_6126));
OAI21X1 g56142(.A0 (n_6122), .A1 (n_5242), .B0 (n_4055), .Y(DATA_9_24));
CLKBUFX1 gbuf_d_11(.A(n_6123), .Y(d_out_11));
CLKBUFX1 gbuf_q_11(.A(q_in_11), .Y(WX663));
OAI21X1 g56139(.A0 (n_6120), .A1 (n_5889), .B0 (n_6095), .Y (n_6883));
INVX1 g56184(.A (WX497), .Y (n_6127));
NAND2X1 g56137(.A (n_6121), .B (n_4719), .Y (n_6123));
CLKBUFX1 gbuf_d_12(.A(n_6118), .Y(d_out_12));
CLKBUFX1 gbuf_q_12(.A(q_in_12), .Y(WX497));
CLKBUFX1 gbuf_d_13(.A(n_6115), .Y(d_out_13));
CLKBUFX1 gbuf_q_13(.A(q_in_13), .Y(WX10993));
CLKBUFX1 gbuf_d_14(.A(n_6114), .Y(d_out_14));
CLKBUFX1 gbuf_q_14(.A(q_in_14), .Y(WX1942));
MX2X1 g56199(.A (n_6117), .B (WX499), .S0 (n_10727), .Y (n_6122));
NAND2X1 g56174(.A (n_6110), .B (n_6555), .Y (n_6121));
INVX1 g56200(.A (DATA_9_23), .Y (n_6120));
NOR2X1 g56228(.A (n_5181), .B (n_6117), .Y (n_6118));
OR2X1 g56232(.A (n_6117), .B (n_3828), .Y (n_6116));
OAI21X1 g55842(.A0 (n_3841), .A1 (n_6106), .B0 (n_6111), .Y (n_6115));
OAI21X1 g55836(.A0 (n_4283), .A1 (n_5415), .B0 (n_6112), .Y (n_6114));
OAI21X1 g56201(.A0 (n_6108), .A1 (n_6091), .B0 (n_4043), .Y(DATA_9_23));
CLKBUFX1 gbuf_d_15(.A(n_6109), .Y(d_out_15));
CLKBUFX1 gbuf_q_15(.A(q_in_15), .Y(WX665));
OAI21X1 g55865(.A0 (n_6102), .A1 (n_4195), .B0 (n_5722), .Y (n_6112));
OAI21X1 g55866(.A0 (n_4551), .A1 (n_6177), .B0 (n_5722), .Y (n_6111));
OAI21X1 g56198(.A0 (n_6099), .A1 (n_5889), .B0 (n_6078), .Y (n_6110));
INVX1 g56243(.A (WX499), .Y (n_6117));
CLKBUFX1 gbuf_d_16(.A(n_6105), .Y(d_out_16));
CLKBUFX1 gbuf_q_16(.A(q_in_16), .Y(WX10995));
CLKBUFX1 gbuf_d_17(.A(n_6107), .Y(d_out_17));
CLKBUFX1 gbuf_q_17(.A(q_in_17), .Y(WX1944));
NAND2X1 g56196(.A (n_6100), .B (n_4717), .Y (n_6109));
CLKBUFX1 gbuf_d_18(.A(n_6097), .Y(d_out_18));
CLKBUFX1 gbuf_q_18(.A(q_in_18), .Y(WX499));
CLKBUFX1 gbuf_d_19(.A(n_6104), .Y(d_out_19));
CLKBUFX1 gbuf_q_19(.A(q_in_19), .Y(WX10831));
CLKBUFX1 gbuf_d_20(.A(n_6103), .Y(d_out_20));
CLKBUFX1 gbuf_q_20(.A(q_in_20), .Y(WX1780));
MX2X1 g56258(.A (n_6096), .B (WX501), .S0 (n_7062), .Y (n_6108));
OAI21X1 g55896(.A0 (n_4558), .A1 (n_6106), .B0 (n_6092), .Y (n_6107));
OAI21X1 g55902(.A0 (n_3834), .A1 (n_6050), .B0 (n_6093), .Y (n_6105));
NOR2X1 g55916(.A (WX10833), .B (n_1648), .Y (n_6104));
NOR2X1 g55920(.A (WX1782), .B (n_5181), .Y (n_6103));
NOR2X1 g55923(.A (WX1782), .B (n_5500), .Y (n_6102));
NOR2X1 g55924(.A (WX10833), .B (n_5811), .Y (n_6177));
NAND2X1 g56233(.A (n_6090), .B (n_6583), .Y (n_6100));
INVX1 g56259(.A (DATA_9_22), .Y (n_6099));
NOR2X1 g56287(.A (n_2849), .B (n_6096), .Y (n_6097));
OR2X1 g56291(.A (n_6096), .B (n_5990), .Y (n_6095));
OAI21X1 g55926(.A0 (n_4549), .A1 (n_6184), .B0 (n_5722), .Y (n_6093));
OAI21X1 g55925(.A0 (n_6083), .A1 (n_4193), .B0 (n_4947), .Y (n_6092));
OAI21X1 g56260(.A0 (n_6081), .A1 (n_6091), .B0 (n_4033), .Y(DATA_9_22));
CLKBUFX1 gbuf_d_21(.A(n_6087), .Y(d_out_21));
CLKBUFX1 gbuf_q_21(.A(q_in_21), .Y(WX10997));
CLKBUFX1 gbuf_d_22(.A(n_6088), .Y(d_out_22));
CLKBUFX1 gbuf_q_22(.A(q_in_22), .Y(WX1946));
CLKBUFX1 gbuf_d_23(.A(n_6086), .Y(d_out_23));
CLKBUFX1 gbuf_q_23(.A(q_in_23), .Y(WX667));
CLKBUFX1 gbuf_d_24(.A(n_6085), .Y(d_out_24));
CLKBUFX1 gbuf_qn_24(.A(qn_in_24), .Y(WX10833));
CLKBUFX1 gbuf_d_25(.A(n_6084), .Y(d_out_25));
CLKBUFX1 gbuf_qn_25(.A(qn_in_25), .Y(WX1782));
OAI21X1 g56257(.A0 (n_6072), .A1 (n_5889), .B0 (n_6053), .Y (n_6090));
INVX1 g56303(.A (WX501), .Y (n_6096));
OAI21X1 g55955(.A0 (n_4556), .A1 (n_5600), .B0 (n_6076), .Y (n_6088));
OAI21X1 g55961(.A0 (n_3839), .A1 (n_6106), .B0 (n_6075), .Y (n_6087));
NAND2X1 g56255(.A (n_6074), .B (n_4716), .Y (n_6086));
CLKBUFX1 gbuf_d_26(.A(n_6080), .Y(d_out_26));
CLKBUFX1 gbuf_q_26(.A(q_in_26), .Y(WX501));
NOR2X1 g55975(.A (WX10835), .B (n_2605), .Y (n_6085));
NOR2X1 g55978(.A (WX1784), .B (n_1648), .Y (n_6084));
NOR2X1 g55982(.A (WX1784), .B (n_5479), .Y (n_6083));
NOR2X1 g55984(.A (WX10835), .B (n_5811), .Y (n_6184));
MX2X1 g56317(.A (n_6079), .B (WX503), .S0 (n_7070), .Y (n_6081));
NOR2X1 g56346(.A (n_5181), .B (n_6079), .Y (n_6080));
OR2X1 g56350(.A (n_6079), .B (n_5990), .Y (n_6078));
OAI21X1 g55983(.A0 (n_6064), .A1 (n_4191), .B0 (n_5460), .Y (n_6076));
OAI21X1 g55987(.A0 (n_4547), .A1 (n_6209), .B0 (n_5619), .Y (n_6075));
NAND2X1 g56292(.A (n_6068), .B (n_6615), .Y (n_6074));
CLKBUFX1 gbuf_d_27(.A(n_6069), .Y(d_out_27));
CLKBUFX1 gbuf_q_27(.A(q_in_27), .Y(WX10999));
CLKBUFX1 gbuf_d_28(.A(n_6070), .Y(d_out_28));
CLKBUFX1 gbuf_q_28(.A(q_in_28), .Y(WX1948));
INVX1 g56318(.A (DATA_9_21), .Y (n_6072));
CLKBUFX1 gbuf_d_29(.A(n_6067), .Y(d_out_29));
CLKBUFX1 gbuf_qn_29(.A(qn_in_29), .Y(WX10835));
CLKBUFX1 gbuf_d_30(.A(n_6066), .Y(d_out_30));
CLKBUFX1 gbuf_qn_30(.A(qn_in_30), .Y(WX1784));
CLKBUFX1 gbuf_d_31(.A(n_6063), .Y(d_out_31));
CLKBUFX1 gbuf_q_31(.A(q_in_31), .Y(WX669));
OAI21X1 g56319(.A0 (n_6061), .A1 (n_6091), .B0 (n_4025), .Y(DATA_9_21));
INVX1 g56362(.A (WX503), .Y (n_6079));
OAI21X1 g56014(.A0 (n_4554), .A1 (n_4803), .B0 (n_6060), .Y (n_6070));
OAI21X1 g56020(.A0 (n_3837), .A1 (n_5482), .B0 (n_6059), .Y (n_6069));
OAI21X1 g56316(.A0 (n_6057), .A1 (n_5889), .B0 (n_6033), .Y (n_6068));
CLKBUFX1 gbuf_d_32(.A(n_6055), .Y(d_out_32));
CLKBUFX1 gbuf_q_32(.A(q_in_32), .Y(WX503));
NOR2X1 g56034(.A (WX10837), .B (n_1648), .Y (n_6067));
NOR2X1 g56036(.A (WX1786), .B (n_2605), .Y (n_6066));
NOR2X1 g56041(.A (WX1786), .B (n_5811), .Y (n_6064));
NAND2X1 g56314(.A (n_6058), .B (n_4715), .Y (n_6063));
NOR2X1 g56045(.A (WX10837), .B (n_5811), .Y (n_6209));
MX2X1 g56376(.A (n_6054), .B (WX505), .S0 (n_6553), .Y (n_6061));
CLKBUFX1 gbuf_d_33(.A(n_6051), .Y(d_out_33));
CLKBUFX1 gbuf_q_33(.A(q_in_33), .Y(WX11001));
CLKBUFX1 gbuf_d_34(.A(n_6052), .Y(d_out_34));
CLKBUFX1 gbuf_q_34(.A(q_in_34), .Y(WX1950));
OAI21X1 g56044(.A0 (n_6046), .A1 (n_4188), .B0 (n_4860), .Y (n_6060));
OAI21X1 g56048(.A0 (n_4545), .A1 (n_6210), .B0 (n_5460), .Y (n_6059));
CLKBUFX1 gbuf_d_35(.A(n_6048), .Y(d_out_35));
CLKBUFX1 gbuf_qn_35(.A(qn_in_35), .Y(WX10837));
NAND2X1 g56351(.A (n_6555), .B (n_8331), .Y (n_6058));
CLKBUFX1 gbuf_d_36(.A(n_6047), .Y(d_out_36));
CLKBUFX1 gbuf_qn_36(.A(qn_in_36), .Y(WX1786));
INVX1 g56377(.A (DATA_9_20), .Y (n_6057));
NOR2X1 g56405(.A (n_2849), .B (n_6054), .Y (n_6055));
OR2X1 g56409(.A (n_6054), .B (n_5990), .Y (n_6053));
OAI21X1 g56073(.A0 (n_4522), .A1 (n_5928), .B0 (n_6042), .Y (n_6052));
OAI21X1 g56378(.A0 (n_6040), .A1 (n_5242), .B0 (n_4082), .Y(DATA_9_20));
OAI21X1 g56079(.A0 (n_3822), .A1 (n_6050), .B0 (n_6041), .Y (n_6051));
CLKBUFX1 gbuf_d_37(.A(n_6043), .Y(d_out_37));
CLKBUFX1 gbuf_q_37(.A(q_in_37), .Y(WX671));
OAI21X1 g56375(.A0 (n_6038), .A1 (n_5889), .B0 (n_6013), .Y (n_8331));
NOR2X1 g56093(.A (WX10839), .B (n_2620), .Y (n_6048));
NOR2X1 g56095(.A (WX1788), .B (n_5181), .Y (n_6047));
INVX1 g56423(.A (WX505), .Y (n_6054));
NOR2X1 g56102(.A (WX1788), .B (n_5811), .Y (n_6046));
NOR2X1 g56106(.A (WX10839), .B (n_5811), .Y (n_6210));
NAND2X1 g56373(.A (n_6039), .B (n_4714), .Y (n_6043));
CLKBUFX1 gbuf_d_38(.A(n_6036), .Y(d_out_38));
CLKBUFX1 gbuf_q_38(.A(q_in_38), .Y(WX505));
OAI21X1 g56105(.A0 (n_6027), .A1 (n_4186), .B0 (n_5722), .Y (n_6042));
OAI21X1 g56107(.A0 (n_4543), .A1 (n_6178), .B0 (n_4860), .Y (n_6041));
CLKBUFX1 gbuf_d_39(.A(n_6031), .Y(d_out_39));
CLKBUFX1 gbuf_q_39(.A(q_in_39), .Y(WX11003));
CLKBUFX1 gbuf_d_40(.A(n_6032), .Y(d_out_40));
CLKBUFX1 gbuf_q_40(.A(q_in_40), .Y(WX1952));
MX2X1 g56435(.A (n_6034), .B (WX507), .S0 (n_6645), .Y (n_6040));
CLKBUFX1 gbuf_d_41(.A(n_6030), .Y(d_out_41));
CLKBUFX1 gbuf_qn_41(.A(qn_in_41), .Y(WX10839));
CLKBUFX1 gbuf_d_42(.A(n_6029), .Y(d_out_42));
CLKBUFX1 gbuf_qn_42(.A(qn_in_42), .Y(WX1788));
NAND2X1 g56410(.A (n_6025), .B (n_6583), .Y (n_6039));
INVX1 g56436(.A (DATA_9_19), .Y (n_6038));
NOR2X1 g56464(.A (n_5181), .B (n_6034), .Y (n_6036));
OR2X1 g56468(.A (n_6034), .B (n_5990), .Y (n_6033));
OAI21X1 g56133(.A0 (n_4496), .A1 (n_5918), .B0 (n_6024), .Y (n_6032));
OAI21X1 g56138(.A0 (n_3836), .A1 (n_5879), .B0 (n_6023), .Y (n_6031));
OAI21X1 g56437(.A0 (n_6021), .A1 (n_5843), .B0 (n_4075), .Y(DATA_9_19));
NOR2X1 g56152(.A (WX10841), .B (n_1648), .Y (n_6030));
NOR2X1 g56154(.A (WX1790), .B (n_1648), .Y (n_6029));
NOR2X1 g56163(.A (WX1790), .B (n_5822), .Y (n_6027));
NOR2X1 g56165(.A (WX10841), .B (n_5479), .Y (n_6178));
CLKBUFX1 gbuf_d_43(.A(n_6022), .Y(d_out_43));
CLKBUFX1 gbuf_q_43(.A(q_in_43), .Y(WX673));
OAI21X1 g56434(.A0 (n_6017), .A1 (n_5889), .B0 (n_5991), .Y (n_6025));
INVX1 g56477(.A (WX507), .Y (n_6034));
OAI21X1 g56164(.A0 (n_6010), .A1 (n_4183), .B0 (n_5566), .Y (n_6024));
OAI21X1 g56166(.A0 (n_4541), .A1 (n_6179), .B0 (n_5722), .Y (n_6023));
CLKBUFX1 gbuf_d_44(.A(n_6019), .Y(d_out_44));
CLKBUFX1 gbuf_q_44(.A(q_in_44), .Y(WX11005));
CLKBUFX1 gbuf_d_45(.A(n_6020), .Y(d_out_45));
CLKBUFX1 gbuf_q_45(.A(q_in_45), .Y(WX1954));
NAND2X1 g56432(.A (n_15853), .B (n_15854), .Y (n_6022));
CLKBUFX1 gbuf_d_46(.A(n_6015), .Y(d_out_46));
CLKBUFX1 gbuf_q_46(.A(q_in_46), .Y(WX507));
CLKBUFX1 gbuf_d_47(.A(n_6012), .Y(d_out_47));
CLKBUFX1 gbuf_qn_47(.A(qn_in_47), .Y(WX10841));
CLKBUFX1 gbuf_d_48(.A(n_6011), .Y(d_out_48));
CLKBUFX1 gbuf_qn_48(.A(qn_in_48), .Y(WX1790));
MX2X1 g56494(.A (n_6014), .B (WX509), .S0 (n_10731), .Y (n_6021));
OAI21X1 g56192(.A0 (n_4488), .A1 (n_5834), .B0 (n_6008), .Y (n_6020));
OAI21X1 g56197(.A0 (n_3827), .A1 (n_5841), .B0 (n_6007), .Y (n_6019));
NAND2X1 g56469(.A (n_6615), .B (n_8332), .Y (n_15854));
INVX1 g56495(.A (DATA_9_18), .Y (n_6017));
NOR2X1 g56523(.A (n_1425), .B (n_6014), .Y (n_6015));
OR2X1 g56527(.A (n_6014), .B (n_5968), .Y (n_6013));
NOR2X1 g56211(.A (WX10843), .B (n_5712), .Y (n_6012));
NOR2X1 g56213(.A (WX1792), .B (n_2620), .Y (n_6011));
NOR2X1 g56222(.A (WX1792), .B (n_5427), .Y (n_6010));
NOR2X1 g56224(.A (WX10843), .B (n_5822), .Y (n_6179));
OAI21X1 g56496(.A0 (n_6001), .A1 (n_5965), .B0 (n_4064), .Y(DATA_9_18));
OAI21X1 g56223(.A0 (n_5998), .A1 (n_4181), .B0 (n_4860), .Y (n_6008));
OAI21X1 g56225(.A0 (n_4537), .A1 (n_6439), .B0 (n_6497), .Y (n_6007));
CLKBUFX1 gbuf_d_49(.A(n_6002), .Y(d_out_49));
CLKBUFX1 gbuf_q_49(.A(q_in_49), .Y(WX11007));
CLKBUFX1 gbuf_d_50(.A(n_6003), .Y(d_out_50));
CLKBUFX1 gbuf_q_50(.A(q_in_50), .Y(WX1956));
CLKBUFX1 gbuf_d_51(.A(n_6004), .Y(d_out_51));
CLKBUFX1 gbuf_q_51(.A(q_in_51), .Y(WX675));
OAI21X1 g56493(.A0 (n_5995), .A1 (n_5889), .B0 (n_5969), .Y (n_8332));
INVX1 g56536(.A (WX509), .Y (n_6014));
CLKBUFX1 gbuf_d_52(.A(n_6000), .Y(d_out_52));
CLKBUFX1 gbuf_qn_52(.A(qn_in_52), .Y(WX10843));
CLKBUFX1 gbuf_d_53(.A(n_5999), .Y(d_out_53));
CLKBUFX1 gbuf_qn_53(.A(qn_in_53), .Y(WX1792));
NAND2X2 g56491(.A (n_5996), .B (n_4711), .Y (n_6004));
CLKBUFX1 gbuf_d_54(.A(n_5993), .Y(d_out_54));
CLKBUFX1 gbuf_q_54(.A(q_in_54), .Y(WX509));
OAI21X1 g56251(.A0 (n_4253), .A1 (n_5439), .B0 (n_5989), .Y (n_6003));
OAI21X1 g56256(.A0 (n_3830), .A1 (n_5845), .B0 (n_5988), .Y (n_6002));
MX2X1 g56553(.A (n_5992), .B (WX511), .S0 (n_7074), .Y (n_6001));
NOR2X1 g56270(.A (WX10845), .B (n_1648), .Y (n_6000));
NOR2X1 g56272(.A (WX1794), .B (n_5181), .Y (n_5999));
NOR2X1 g56281(.A (WX1794), .B (n_5662), .Y (n_5998));
NAND2X1 g56528(.A (n_5987), .B (n_6575), .Y (n_5996));
INVX1 g56554(.A (DATA_9_17), .Y (n_5995));
NOR2X1 g56582(.A (n_1425), .B (n_5992), .Y (n_5993));
OR2X1 g56587(.A (n_5992), .B (n_5990), .Y (n_5991));
OAI21X1 g56282(.A0 (n_5981), .A1 (n_4179), .B0 (n_5566), .Y (n_5989));
OAI21X1 g56285(.A0 (n_4625), .A1 (n_6216), .B0 (n_4860), .Y (n_5988));
CLKBUFX1 gbuf_d_55(.A(n_5985), .Y(d_out_55));
CLKBUFX1 gbuf_q_55(.A(q_in_55), .Y(WX11009));
CLKBUFX1 gbuf_d_56(.A(n_5986), .Y(d_out_56));
CLKBUFX1 gbuf_q_56(.A(q_in_56), .Y(WX1958));
OAI21X1 g56555(.A0 (n_5978), .A1 (n_5965), .B0 (n_4057), .Y(DATA_9_17));
CLKBUFX1 gbuf_d_57(.A(n_6524), .Y(d_out_57));
CLKBUFX1 gbuf_q_57(.A(q_in_57), .Y(WX677));
CLKBUFX1 gbuf_d_58(.A(n_5983), .Y(d_out_58));
CLKBUFX1 gbuf_qn_58(.A(qn_in_58), .Y(WX10845));
CLKBUFX1 gbuf_d_59(.A(n_5982), .Y(d_out_59));
CLKBUFX1 gbuf_qn_59(.A(qn_in_59), .Y(WX1794));
OAI21X1 g56552(.A0 (n_5973), .A1 (n_5889), .B0 (n_5940), .Y (n_5987));
INVX1 g56597(.A (WX511), .Y (n_5992));
OAI21X1 g56310(.A0 (n_4251), .A1 (n_5630), .B0 (n_5977), .Y (n_5986));
OAI21X1 g56315(.A0 (n_3833), .A1 (n_5882), .B0 (n_5976), .Y (n_5985));
CLKBUFX1 gbuf_d_60(.A(n_5971), .Y(d_out_60));
CLKBUFX1 gbuf_q_60(.A(q_in_60), .Y(WX511));
CLKBUFX1 gbuf_d_61(.A(n_5974), .Y(d_out_61));
CLKBUFX1 gbuf_q_61(.A(q_in_61), .Y(WX9718));
NOR2X1 g56329(.A (WX10847), .B (n_5712), .Y (n_5983));
NOR2X1 g56331(.A (WX1796), .B (n_1425), .Y (n_5982));
NOR2X1 g56340(.A (WX1796), .B (n_5662), .Y (n_5981));
NOR2X1 g56342(.A (WX10847), .B (n_5811), .Y (n_6216));
MX2X1 g56612(.A (n_5970), .B (WX513), .S0 (n_9800), .Y (n_5978));
CLKBUFX1 gbuf_d_62(.A(n_5966), .Y(d_out_62));
CLKBUFX1 gbuf_q_62(.A(q_in_62), .Y(WX11011));
CLKBUFX1 gbuf_d_63(.A(n_5967), .Y(d_out_63));
CLKBUFX1 gbuf_q_63(.A(q_in_63), .Y(WX1960));
OAI21X1 g56341(.A0 (n_5961), .A1 (n_4176), .B0 (n_7087), .Y (n_5977));
OAI21X1 g56345(.A0 (n_4535), .A1 (n_6217), .B0 (n_5722), .Y (n_5976));
CLKBUFX1 gbuf_d_64(.A(n_5964), .Y(d_out_64));
CLKBUFX1 gbuf_qn_64(.A(qn_in_64), .Y(WX10847));
CLKBUFX1 gbuf_d_65(.A(n_5963), .Y(d_out_65));
CLKBUFX1 gbuf_qn_65(.A(qn_in_65), .Y(WX1796));
OAI21X1 g55798(.A0 (n_4534), .A1 (n_5183), .B0 (n_5959), .Y (n_5974));
INVX1 g56613(.A (DATA_9_16), .Y (n_5973));
NOR2X1 g56641(.A (n_1425), .B (n_5970), .Y (n_5971));
OR2X1 g56647(.A (n_5970), .B (n_5968), .Y (n_5969));
OAI21X1 g56369(.A0 (n_4474), .A1 (n_5418), .B0 (n_5956), .Y (n_5967));
OAI21X1 g56374(.A0 (n_3819), .A1 (n_5892), .B0 (n_5954), .Y (n_5966));
OAI21X1 g56614(.A0 (n_5951), .A1 (n_5965), .B0 (n_4049), .Y(DATA_9_16));
CLKBUFX1 gbuf_d_66(.A(n_6561), .Y(d_out_66));
CLKBUFX1 gbuf_q_66(.A(q_in_66), .Y(WX679));
NOR2X1 g56388(.A (WX10849), .B (n_5712), .Y (n_5964));
NOR2X1 g56390(.A (WX1798), .B (n_1648), .Y (n_5963));
NOR2X1 g56399(.A (WX1798), .B (n_5427), .Y (n_5961));
NOR2X1 g56403(.A (WX10849), .B (n_5479), .Y (n_6217));
OAI21X1 g55820(.A0 (n_4592), .A1 (n_6218), .B0 (n_3183), .Y (n_5959));
INVX1 g56656(.A (WX513), .Y (n_5970));
CLKBUFX1 gbuf_d_67(.A(n_5952), .Y(d_out_67));
CLKBUFX1 gbuf_q_67(.A(q_in_67), .Y(WX8427));
CLKBUFX1 gbuf_d_68(.A(n_5950), .Y(d_out_68));
CLKBUFX1 gbuf_q_68(.A(q_in_68), .Y(WX9720));
OAI21X1 g56400(.A0 (n_5936), .A1 (n_4174), .B0 (n_5722), .Y (n_5956));
OAI21X1 g56404(.A0 (n_4533), .A1 (n_6180), .B0 (n_5722), .Y (n_5954));
CLKBUFX1 gbuf_d_69(.A(n_5942), .Y(d_out_69));
CLKBUFX1 gbuf_q_69(.A(q_in_69), .Y(WX513));
CLKBUFX1 gbuf_d_70(.A(n_5947), .Y(d_out_70));
CLKBUFX1 gbuf_q_70(.A(q_in_70), .Y(WX9556));
CLKBUFX1 gbuf_d_71(.A(n_5948), .Y(d_out_71));
CLKBUFX1 gbuf_q_71(.A(q_in_71), .Y(WX11013));
CLKBUFX1 gbuf_d_72(.A(n_5949), .Y(d_out_72));
CLKBUFX1 gbuf_q_72(.A(q_in_72), .Y(WX1962));
OAI21X1 g55797(.A0 (n_4591), .A1 (n_5886), .B0 (n_5939), .Y (n_5952));
CLKBUFX1 gbuf_d_73(.A(n_5938), .Y(d_out_73));
CLKBUFX1 gbuf_qn_73(.A(qn_in_73), .Y(WX10849));
CLKBUFX1 gbuf_d_74(.A(n_5937), .Y(d_out_74));
CLKBUFX1 gbuf_qn_74(.A(qn_in_74), .Y(WX1798));
MX2X1 g56671(.A (n_5941), .B (WX515), .S0 (n_7078), .Y (n_5951));
OAI21X1 g55837(.A0 (n_4532), .A1 (n_5892), .B0 (n_5934), .Y (n_5950));
OAI21X1 g56428(.A0 (n_4464), .A1 (n_5879), .B0 (n_5933), .Y (n_5949));
OAI21X1 g56433(.A0 (n_3844), .A1 (n_5928), .B0 (n_5931), .Y (n_5948));
AND2X1 g55867(.A (WX9558), .B (n_2383), .Y (n_5947));
AND2X1 g55869(.A (WX9558), .B (n_5828), .Y (n_6218));
INVX1 g56672(.A (DATA_9_15), .Y (n_5944));
NOR2X1 g56700(.A (n_1425), .B (n_5941), .Y (n_5942));
OR2X1 g56706(.A (n_5941), .B (n_4882), .Y (n_5940));
OAI21X1 g55818(.A0 (n_4364), .A1 (n_6658), .B0 (n_5619), .Y (n_5939));
NOR2X1 g56447(.A (WX10851), .B (n_1425), .Y (n_5938));
NOR2X1 g56449(.A (WX1800), .B (n_1648), .Y (n_5937));
NOR2X1 g56458(.A (WX1800), .B (n_5838), .Y (n_5936));
NOR2X1 g56462(.A (WX10851), .B (n_5479), .Y (n_6180));
OAI21X1 g55870(.A0 (n_4590), .A1 (n_6185), .B0 (n_5556), .Y (n_5934));
OAI21X1 g56673(.A0 (n_5917), .A1 (n_5242), .B0 (n_4045), .Y(DATA_9_15));
CLKBUFX1 gbuf_d_75(.A(n_5929), .Y(d_out_75));
CLKBUFX1 gbuf_q_75(.A(q_in_75), .Y(WX7136));
CLKBUFX1 gbuf_d_76(.A(n_5925), .Y(d_out_76));
CLKBUFX1 gbuf_q_76(.A(q_in_76), .Y(WX8429));
CLKBUFX1 gbuf_d_77(.A(n_5926), .Y(d_out_77));
CLKBUFX1 gbuf_q_77(.A(q_in_77), .Y(WX9722));
CLKBUFX1 gbuf_d_78(.A(n_5927), .Y(d_out_78));
CLKBUFX1 gbuf_q_78(.A(q_in_78), .Y(WX681));
OAI21X1 g56459(.A0 (n_5910), .A1 (n_4172), .B0 (n_5722), .Y (n_5933));
OAI21X1 g56463(.A0 (n_4531), .A1 (n_6214), .B0 (n_4860), .Y (n_5931));
CLKBUFX1 gbuf_d_79(.A(n_5924), .Y(d_out_79));
CLKBUFX1 gbuf_q_79(.A(q_in_79), .Y(WX9558));
INVX1 g56715(.A (WX515), .Y (n_5941));
CLKBUFX1 gbuf_d_80(.A(n_5922), .Y(d_out_80));
CLKBUFX1 gbuf_q_80(.A(q_in_80), .Y(WX8265));
CLKBUFX1 gbuf_d_81(.A(n_5919), .Y(d_out_81));
CLKBUFX1 gbuf_q_81(.A(q_in_81), .Y(WX11015));
CLKBUFX1 gbuf_d_82(.A(n_5921), .Y(d_out_82));
CLKBUFX1 gbuf_q_82(.A(q_in_82), .Y(WX1964));
CLKBUFX1 gbuf_d_83(.A(n_5914), .Y(d_out_83));
CLKBUFX1 gbuf_qn_83(.A(qn_in_83), .Y(WX10851));
CLKBUFX1 gbuf_d_84(.A(n_5912), .Y(d_out_84));
CLKBUFX1 gbuf_qn_84(.A(qn_in_84), .Y(WX1800));
OAI21X1 g55801(.A0 (n_4363), .A1 (n_5928), .B0 (n_5907), .Y (n_5929));
NAND2X1 g56668(.A (n_5905), .B (n_4706), .Y (n_5927));
CLKBUFX1 gbuf_d_85(.A(n_5901), .Y(d_out_85));
CLKBUFX1 gbuf_q_85(.A(q_in_85), .Y(WX515));
OAI21X1 g55897(.A0 (n_4530), .A1 (n_5598), .B0 (n_5916), .Y (n_5926));
OAI21X1 g55835(.A0 (n_4589), .A1 (n_5493), .B0 (n_5915), .Y (n_5925));
NOR2X1 g55927(.A (WX9560), .B (n_5712), .Y (n_5924));
NOR2X1 g55929(.A (WX9560), .B (n_5479), .Y (n_6185));
AND2X1 g55858(.A (WX8267), .B (n_2396), .Y (n_5922));
OAI21X1 g56487(.A0 (n_4241), .A1 (n_5830), .B0 (n_5896), .Y (n_5921));
AND2X1 g55861(.A (WX8267), .B (n_5873), .Y (n_6658));
OAI21X1 g56492(.A0 (n_3812), .A1 (n_5918), .B0 (n_5894), .Y (n_5919));
MX2X1 g56730(.A (n_5899), .B (WX517), .S0 (n_4044), .Y (n_5917));
OAI21X1 g55930(.A0 (n_4588), .A1 (n_6187), .B0 (n_5460), .Y (n_5916));
OAI21X1 g55862(.A0 (n_5884), .A1 (n_4362), .B0 (n_5722), .Y (n_5915));
NOR2X1 g56507(.A (WX10853), .B (n_5712), .Y (n_5914));
NOR2X1 g56508(.A (WX1802), .B (n_5712), .Y (n_5912));
NOR2X1 g56517(.A (WX1802), .B (n_5500), .Y (n_5910));
NOR2X1 g56521(.A (WX10853), .B (n_5500), .Y (n_6214));
OAI21X1 g55824(.A0 (n_4413), .A1 (n_6186), .B0 (n_5722), .Y (n_5907));
NAND2X1 g56707(.A (n_5890), .B (n_6575), .Y (n_5905));
INVX1 g56731(.A (DATA_9_14), .Y (n_5903));
NOR2X1 g56758(.A (n_1425), .B (n_5899), .Y (n_5901));
OR2X1 g56764(.A (n_5899), .B (n_5968), .Y (n_5898));
CLKBUFX1 gbuf_d_86(.A(n_5893), .Y(d_out_86));
CLKBUFX1 gbuf_q_86(.A(q_in_86), .Y(WX5845));
CLKBUFX1 gbuf_d_87(.A(n_5887), .Y(d_out_87));
CLKBUFX1 gbuf_q_87(.A(q_in_87), .Y(WX7138));
CLKBUFX1 gbuf_d_88(.A(n_5888), .Y(d_out_88));
CLKBUFX1 gbuf_q_88(.A(q_in_88), .Y(WX8431));
CLKBUFX1 gbuf_d_89(.A(n_5891), .Y(d_out_89));
CLKBUFX1 gbuf_q_89(.A(q_in_89), .Y(WX9724));
CLKBUFX1 gbuf_d_90(.A(n_5878), .Y(d_out_90));
CLKBUFX1 gbuf_qn_90(.A(qn_in_90), .Y(WX9560));
OAI21X1 g56518(.A0 (n_5865), .A1 (n_4170), .B0 (n_4947), .Y (n_5896));
OAI21X1 g56522(.A0 (n_4529), .A1 (n_6215), .B0 (n_7087), .Y (n_5894));
CLKBUFX1 gbuf_d_91(.A(n_5885), .Y(d_out_91));
CLKBUFX1 gbuf_q_91(.A(q_in_91), .Y(WX8267));
OAI21X1 g56732(.A0 (n_5858), .A1 (n_5965), .B0 (n_4039), .Y(DATA_9_14));
CLKBUFX1 gbuf_d_92(.A(n_5883), .Y(d_out_92));
CLKBUFX1 gbuf_q_92(.A(q_in_92), .Y(WX4554));
CLKBUFX1 gbuf_d_93(.A(n_5876), .Y(d_out_93));
CLKBUFX1 gbuf_q_93(.A(q_in_93), .Y(WX6974));
CLKBUFX1 gbuf_d_94(.A(n_5880), .Y(d_out_94));
CLKBUFX1 gbuf_q_94(.A(q_in_94), .Y(WX11017));
CLKBUFX1 gbuf_d_95(.A(n_5881), .Y(d_out_95));
CLKBUFX1 gbuf_q_95(.A(q_in_95), .Y(WX1966));
CLKBUFX1 gbuf_d_96(.A(n_5872), .Y(d_out_96));
CLKBUFX1 gbuf_q_96(.A(q_in_96), .Y(WX683));
OAI21X1 g55800(.A0 (n_4412), .A1 (n_5892), .B0 (n_5869), .Y (n_5893));
OAI21X1 g55956(.A0 (n_4273), .A1 (n_5841), .B0 (n_5862), .Y (n_5891));
CLKBUFX1 gbuf_d_97(.A(n_5867), .Y(d_out_97));
CLKBUFX1 gbuf_qn_97(.A(qn_in_97), .Y(WX10853));
CLKBUFX1 gbuf_d_98(.A(n_5866), .Y(d_out_98));
CLKBUFX1 gbuf_qn_98(.A(qn_in_98), .Y(WX1802));
OAI21X1 g56729(.A0 (n_5853), .A1 (n_5889), .B0 (n_5790), .Y (n_5890));
OAI21X1 g55895(.A0 (n_4303), .A1 (n_5750), .B0 (n_5871), .Y (n_5888));
INVX1 g56775(.A (WX517), .Y (n_5899));
OAI21X1 g55840(.A0 (n_4361), .A1 (n_5886), .B0 (n_5860), .Y (n_5887));
NOR2X1 g55917(.A (WX8269), .B (n_5712), .Y (n_5885));
NOR2X1 g55921(.A (WX8269), .B (n_5838), .Y (n_5884));
OAI21X1 g55799(.A0 (n_4478), .A1 (n_5882), .B0 (n_5857), .Y (n_5883));
OAI21X1 g56547(.A0 (n_4460), .A1 (n_5235), .B0 (n_5856), .Y (n_5881));
OAI21X1 g56551(.A0 (n_3829), .A1 (n_5879), .B0 (n_5855), .Y (n_5880));
NOR2X1 g55985(.A (WX9562), .B (n_1648), .Y (n_5878));
AND2X1 g55879(.A (WX6976), .B (n_2383), .Y (n_5876));
NOR2X1 g55988(.A (WX9562), .B (n_5811), .Y (n_6187));
AND2X1 g55881(.A (WX6976), .B (n_5873), .Y (n_6186));
NAND2X2 g56727(.A (n_5854), .B (n_4704), .Y (n_5872));
CLKBUFX1 gbuf_d_99(.A(n_5851), .Y(d_out_99));
CLKBUFX1 gbuf_q_99(.A(q_in_99), .Y(WX517));
OAI21X1 g55922(.A0 (n_4360), .A1 (n_6189), .B0 (n_5722), .Y (n_5871));
OAI21X1 g55822(.A0 (n_4479), .A1 (n_6188), .B0 (n_5566), .Y (n_5869));
NOR2X1 g56567(.A (WX10855), .B (n_2851), .Y (n_5867));
NOR2X1 g56568(.A (WX1804), .B (n_2851), .Y (n_5866));
NOR2X1 g56577(.A (WX1804), .B (n_5427), .Y (n_5865));
NOR2X1 g56581(.A (WX10855), .B (n_5811), .Y (n_6215));
OAI21X1 g55989(.A0 (n_5823), .A1 (n_4302), .B0 (n_6497), .Y (n_5862));
OAI21X1 g55882(.A0 (n_4411), .A1 (n_6665), .B0 (n_5619), .Y (n_5860));
MX2X1 g56789(.A (n_5849), .B (WX519), .S0 (n_4038), .Y (n_5858));
CLKBUFX1 gbuf_d_100(.A(n_5842), .Y(d_out_100));
CLKBUFX1 gbuf_q_100(.A(q_in_100), .Y(WX5847));
CLKBUFX1 gbuf_d_101(.A(n_5844), .Y(d_out_101));
CLKBUFX1 gbuf_q_101(.A(q_in_101), .Y(WX7140));
CLKBUFX1 gbuf_d_102(.A(n_5847), .Y(d_out_102));
CLKBUFX1 gbuf_q_102(.A(q_in_102), .Y(WX8433));
CLKBUFX1 gbuf_d_103(.A(n_5846), .Y(d_out_103));
CLKBUFX1 gbuf_q_103(.A(q_in_103), .Y(WX9726));
CLKBUFX1 gbuf_d_104(.A(n_5837), .Y(d_out_104));
CLKBUFX1 gbuf_qn_104(.A(qn_in_104), .Y(WX8269));
OAI21X1 g55821(.A0 (n_4623), .A1 (n_6219), .B0 (n_5556), .Y (n_5857));
OAI21X1 g56580(.A0 (n_5813), .A1 (n_4168), .B0 (n_5460), .Y (n_5856));
OAI21X1 g56583(.A0 (n_5812), .A1 (n_4272), .B0 (n_5722), .Y (n_5855));
CLKBUFX1 gbuf_d_105(.A(n_5824), .Y(d_out_105));
CLKBUFX1 gbuf_qn_105(.A(qn_in_105), .Y(WX9562));
CLKBUFX1 gbuf_d_106(.A(n_5840), .Y(d_out_106));
CLKBUFX1 gbuf_q_106(.A(q_in_106), .Y(WX6976));
NAND2X1 g56765(.A (n_6575), .B (n_8333), .Y (n_5854));
INVX1 g56790(.A (DATA_9_13), .Y (n_5853));
CLKBUFX1 gbuf_d_107(.A(n_5826), .Y(d_out_107));
CLKBUFX1 gbuf_q_107(.A(q_in_107), .Y(WX4556));
CLKBUFX1 gbuf_d_108(.A(n_5833), .Y(d_out_108));
CLKBUFX1 gbuf_q_108(.A(q_in_108), .Y(WX5683));
NOR2X1 g56815(.A (n_5181), .B (n_5849), .Y (n_5851));
CLKBUFX1 gbuf_d_109(.A(n_5835), .Y(d_out_109));
CLKBUFX1 gbuf_q_109(.A(q_in_109), .Y(WX1968));
CLKBUFX1 gbuf_d_110(.A(n_5831), .Y(d_out_110));
CLKBUFX1 gbuf_q_110(.A(q_in_110), .Y(WX11019));
OR2X1 g56822(.A (n_5849), .B (n_5990), .Y (n_5848));
OAI21X1 g55954(.A0 (n_4584), .A1 (n_5825), .B0 (n_5818), .Y (n_5847));
CLKBUFX1 gbuf_d_111(.A(n_5816), .Y(d_out_111));
CLKBUFX1 gbuf_qn_111(.A(qn_in_111), .Y(WX10855));
CLKBUFX1 gbuf_d_112(.A(n_5815), .Y(d_out_112));
CLKBUFX1 gbuf_qn_112(.A(qn_in_112), .Y(WX1804));
OAI21X1 g56015(.A0 (n_4526), .A1 (n_5845), .B0 (n_5809), .Y (n_5846));
OAI21X1 g55900(.A0 (n_4357), .A1 (n_5879), .B0 (n_5821), .Y (n_5844));
OAI21X1 g56791(.A0 (n_5803), .A1 (n_5843), .B0 (n_4035), .Y(DATA_9_13));
CLKBUFX1 gbuf_d_113(.A(n_5820), .Y(d_out_113));
CLKBUFX1 gbuf_q_113(.A(q_in_113), .Y(WX4392));
CLKBUFX1 gbuf_d_114(.A(n_6533), .Y(d_out_114));
CLKBUFX1 gbuf_q_114(.A(q_in_114), .Y(WX685));
OAI21X1 g55839(.A0 (n_4410), .A1 (n_5841), .B0 (n_5814), .Y (n_5842));
NOR2X1 g55939(.A (WX6978), .B (n_2620), .Y (n_5840));
NOR2X1 g55941(.A (WX6978), .B (n_5838), .Y (n_6665));
NOR2X1 g55976(.A (WX8271), .B (n_2620), .Y (n_5837));
OAI21X1 g56607(.A0 (n_4452), .A1 (n_5834), .B0 (n_5806), .Y (n_5835));
AND2X1 g55874(.A (WX5685), .B (n_2378), .Y (n_5833));
NOR2X1 g55980(.A (WX8271), .B (n_5838), .Y (n_6189));
OAI21X1 g56610(.A0 (n_3826), .A1 (n_5830), .B0 (n_5804), .Y (n_5831));
AND2X1 g55875(.A (WX5685), .B (n_5828), .Y (n_6188));
OAI21X1 g56788(.A0 (n_5796), .A1 (n_5889), .B0 (n_5743), .Y (n_8333));
OAI21X1 g55838(.A0 (n_4476), .A1 (n_5825), .B0 (n_5807), .Y (n_5826));
INVX1 g56834(.A (WX519), .Y (n_5849));
NOR2X1 g56042(.A (WX9564), .B (n_5712), .Y (n_5824));
NOR2X1 g56046(.A (WX9564), .B (n_5822), .Y (n_5823));
OAI21X1 g55942(.A0 (n_4409), .A1 (n_6671), .B0 (n_5556), .Y (n_5821));
AND2X1 g55868(.A (WX4394), .B (n_2529), .Y (n_5820));
AND2X1 g55871(.A (WX4394), .B (n_5828), .Y (n_6219));
OAI21X1 g55981(.A0 (n_4356), .A1 (n_6220), .B0 (n_5722), .Y (n_5818));
NOR2X1 g56627(.A (WX10857), .B (n_3188), .Y (n_5816));
NOR2X1 g56628(.A (WX1806), .B (n_1648), .Y (n_5815));
OAI21X1 g55876(.A0 (n_4477), .A1 (n_6190), .B0 (n_4860), .Y (n_5814));
NOR2X1 g56639(.A (WX1806), .B (n_5427), .Y (n_5813));
NOR2X1 g56642(.A (WX10857), .B (n_5811), .Y (n_5812));
CLKBUFX1 gbuf_d_115(.A(n_5794), .Y(d_out_115));
CLKBUFX1 gbuf_q_115(.A(q_in_115), .Y(WX3263));
CLKBUFX1 gbuf_d_116(.A(n_5798), .Y(d_out_116));
CLKBUFX1 gbuf_q_116(.A(q_in_116), .Y(WX5849));
CLKBUFX1 gbuf_d_117(.A(n_5801), .Y(d_out_117));
CLKBUFX1 gbuf_q_117(.A(q_in_117), .Y(WX7142));
CLKBUFX1 gbuf_d_118(.A(n_5800), .Y(d_out_118));
CLKBUFX1 gbuf_q_118(.A(q_in_118), .Y(WX8435));
CLKBUFX1 gbuf_d_119(.A(n_5802), .Y(d_out_119));
CLKBUFX1 gbuf_q_119(.A(q_in_119), .Y(WX9728));
CLKBUFX1 gbuf_d_120(.A(n_5792), .Y(d_out_120));
CLKBUFX1 gbuf_q_120(.A(q_in_120), .Y(WX519));
OAI21X1 g56047(.A0 (n_4583), .A1 (n_6659), .B0 (n_5722), .Y (n_5809));
CLKBUFX1 gbuf_d_121(.A(n_5789), .Y(d_out_121));
CLKBUFX1 gbuf_qn_121(.A(qn_in_121), .Y(WX9564));
CLKBUFX1 gbuf_d_122(.A(n_5781), .Y(d_out_122));
CLKBUFX1 gbuf_qn_122(.A(qn_in_122), .Y(WX6978));
OAI21X1 g55872(.A0 (n_5771), .A1 (n_9405), .B0 (n_5556), .Y (n_5807));
OAI21X1 g56640(.A0 (n_5765), .A1 (n_4166), .B0 (n_5460), .Y (n_5806));
OAI21X1 g56644(.A0 (n_4525), .A1 (n_6181), .B0 (n_5722), .Y (n_5804));
CLKBUFX1 gbuf_d_123(.A(n_5776), .Y(d_out_123));
CLKBUFX1 gbuf_qn_123(.A(qn_in_123), .Y(WX8271));
CLKBUFX1 gbuf_d_124(.A(n_5788), .Y(d_out_124));
CLKBUFX1 gbuf_q_124(.A(q_in_124), .Y(WX5685));
CLKBUFX1 gbuf_d_125(.A(n_5777), .Y(d_out_125));
CLKBUFX1 gbuf_q_125(.A(q_in_125), .Y(WX4558));
CLKBUFX1 gbuf_d_126(.A(n_7094), .Y(d_out_126));
CLKBUFX1 gbuf_q_126(.A(q_in_126), .Y(WX11021));
CLKBUFX1 gbuf_d_127(.A(n_5784), .Y(d_out_127));
CLKBUFX1 gbuf_q_127(.A(q_in_127), .Y(WX1970));
MX2X1 g56848(.A (n_5791), .B (WX521), .S0 (n_6573), .Y (n_5803));
OAI21X1 g56074(.A0 (n_4271), .A1 (n_5841), .B0 (n_5769), .Y (n_5802));
OAI21X1 g55959(.A0 (n_4123), .A1 (n_5576), .B0 (n_5766), .Y (n_5801));
CLKBUFX1 gbuf_d_128(.A(n_5768), .Y(d_out_128));
CLKBUFX1 gbuf_qn_128(.A(qn_in_128), .Y(WX10857));
CLKBUFX1 gbuf_d_129(.A(n_5767), .Y(d_out_129));
CLKBUFX1 gbuf_qn_129(.A(qn_in_129), .Y(WX1806));
CLKBUFX1 gbuf_d_130(.A(n_5773), .Y(d_out_130));
CLKBUFX1 gbuf_q_130(.A(q_in_130), .Y(WX4394));
OAI21X1 g56013(.A0 (n_4582), .A1 (n_5439), .B0 (n_5763), .Y (n_5800));
OAI21X1 g55899(.A0 (n_4408), .A1 (n_5549), .B0 (n_5770), .Y (n_5798));
INVX1 g56849(.A (DATA_9_12), .Y (n_5796));
OAI21X1 g55795(.A0 (n_4622), .A1 (n_5183), .B0 (n_5774), .Y (n_5794));
NOR2X1 g56873(.A (n_5181), .B (n_5791), .Y (n_5792));
OR2X1 g56881(.A (n_5791), .B (n_5968), .Y (n_5790));
NOR2X1 g56100(.A (WX9566), .B (n_5181), .Y (n_5789));
NOR2X1 g55934(.A (WX5687), .B (n_5181), .Y (n_5788));
NOR2X1 g55935(.A (WX5687), .B (n_5838), .Y (n_6190));
NOR2X1 g56103(.A (WX9566), .B (n_5500), .Y (n_6659));
OAI21X1 g56666(.A0 (n_4231), .A1 (n_5468), .B0 (n_5759), .Y (n_5784));
NOR2X1 g55998(.A (WX6980), .B (n_2620), .Y (n_5781));
NOR2X1 g56000(.A (WX6980), .B (n_5838), .Y (n_6671));
OAI21X1 g55898(.A0 (n_4249), .A1 (n_5892), .B0 (n_5760), .Y (n_5777));
CLKBUFX1 gbuf_d_131(.A(n_5755), .Y(d_out_131));
CLKBUFX1 gbuf_q_131(.A(q_in_131), .Y(WX687));
NOR2X1 g56035(.A (WX8273), .B (n_1425), .Y (n_5776));
NOR2X1 g56039(.A (WX8273), .B (n_5500), .Y (n_6220));
OAI21X1 g56850(.A0 (n_5748), .A1 (n_5709), .B0 (n_4029), .Y(DATA_9_12));
OAI21X1 g55816(.A0 (n_4230), .A1 (n_8538), .B0 (n_4860), .Y (n_5774));
NOR2X1 g55928(.A (WX4396), .B (n_5712), .Y (n_5773));
NOR2X1 g55931(.A (WX4396), .B (n_5479), .Y (n_5771));
OAI21X1 g55936(.A0 (n_5732), .A1 (n_9421), .B0 (n_4860), .Y (n_5770));
OAI21X1 g56104(.A0 (n_4581), .A1 (n_6685), .B0 (n_5722), .Y (n_5769));
NOR2X1 g56686(.A (WX10859), .B (n_5181), .Y (n_5768));
NOR2X1 g56687(.A (WX1808), .B (n_3188), .Y (n_5767));
OAI21X1 g56001(.A0 (n_5747), .A1 (n_9423), .B0 (n_5706), .Y (n_5766));
NOR2X1 g56698(.A (WX1808), .B (n_4882), .Y (n_5765));
NOR2X1 g56702(.A (WX10859), .B (n_5838), .Y (n_6181));
CLKBUFX1 gbuf_d_132(.A(n_5751), .Y(d_out_132));
CLKBUFX1 gbuf_q_132(.A(q_in_132), .Y(WX3265));
CLKBUFX1 gbuf_d_133(.A(n_5752), .Y(d_out_133));
CLKBUFX1 gbuf_q_133(.A(q_in_133), .Y(WX5851));
CLKBUFX1 gbuf_d_134(.A(n_5749), .Y(d_out_134));
CLKBUFX1 gbuf_q_134(.A(q_in_134), .Y(WX7144));
CLKBUFX1 gbuf_d_135(.A(n_5754), .Y(d_out_135));
CLKBUFX1 gbuf_q_135(.A(q_in_135), .Y(WX8437));
CLKBUFX1 gbuf_d_136(.A(n_5753), .Y(d_out_136));
CLKBUFX1 gbuf_q_136(.A(q_in_136), .Y(WX9730));
OAI21X1 g56040(.A0 (n_4122), .A1 (n_9814), .B0 (n_4947), .Y (n_5763));
INVX1 g56893(.A (WX521), .Y (n_5791));
CLKBUFX1 gbuf_d_137(.A(n_5742), .Y(d_out_137));
CLKBUFX1 gbuf_qn_137(.A(qn_in_137), .Y(WX8273));
OAI21X1 g55932(.A0 (n_15855), .A1 (n_15856), .B0 (n_5722), .Y(n_5760));
CLKBUFX1 gbuf_d_138(.A(n_5733), .Y(d_out_138));
CLKBUFX1 gbuf_qn_138(.A(qn_in_138), .Y(WX5687));
CLKBUFX1 gbuf_d_139(.A(n_5737), .Y(d_out_139));
CLKBUFX1 gbuf_qn_139(.A(qn_in_139), .Y(WX9566));
OAI21X1 g56699(.A0 (n_5711), .A1 (n_4164), .B0 (n_4860), .Y (n_5759));
CLKBUFX1 gbuf_d_140(.A(n_5725), .Y(d_out_140));
CLKBUFX1 gbuf_qn_140(.A(qn_in_140), .Y(WX6980));
CLKBUFX1 gbuf_d_141(.A(n_5735), .Y(d_out_141));
CLKBUFX1 gbuf_q_141(.A(q_in_141), .Y(WX3101));
CLKBUFX1 gbuf_d_142(.A(n_5738), .Y(d_out_142));
CLKBUFX1 gbuf_q_142(.A(q_in_142), .Y(WX4560));
CLKBUFX1 gbuf_d_143(.A(n_5730), .Y(d_out_143));
CLKBUFX1 gbuf_q_143(.A(q_in_143), .Y(WX11023));
CLKBUFX1 gbuf_d_144(.A(n_5731), .Y(d_out_144));
CLKBUFX1 gbuf_q_144(.A(q_in_144), .Y(WX1972));
NAND2X1 g56845(.A (n_5728), .B (n_4702), .Y (n_5755));
CLKBUFX1 gbuf_d_145(.A(n_5745), .Y(d_out_145));
CLKBUFX1 gbuf_q_145(.A(q_in_145), .Y(WX521));
OAI21X1 g56072(.A0 (n_4577), .A1 (n_4868), .B0 (n_5723), .Y (n_5754));
CLKBUFX1 gbuf_d_146(.A(n_5719), .Y(d_out_146));
CLKBUFX1 gbuf_qn_146(.A(qn_in_146), .Y(WX4396));
OAI21X1 g56132(.A0 (n_4524), .A1 (n_5825), .B0 (n_5720), .Y (n_5753));
OAI21X1 g55958(.A0 (n_4406), .A1 (n_5834), .B0 (n_5716), .Y (n_5752));
OAI21X1 g55834(.A0 (n_4322), .A1 (n_5750), .B0 (n_5721), .Y (n_5751));
CLKBUFX1 gbuf_d_147(.A(n_5714), .Y(d_out_147));
CLKBUFX1 gbuf_qn_147(.A(qn_in_147), .Y(WX10859));
CLKBUFX1 gbuf_d_148(.A(n_5713), .Y(d_out_148));
CLKBUFX1 gbuf_qn_148(.A(qn_in_148), .Y(WX1808));
OAI21X1 g56018(.A0 (n_4353), .A1 (n_5393), .B0 (n_5724), .Y (n_5749));
MX2X1 g56907(.A (n_5744), .B (WX523), .S0 (n_10735), .Y (n_5748));
NOR2X1 g56059(.A (WX6982), .B (n_5838), .Y (n_5747));
NOR2X1 g56931(.A (n_1425), .B (n_5744), .Y (n_5745));
OR2X1 g56939(.A (n_5744), .B (n_5990), .Y (n_5743));
NOR2X1 g56094(.A (WX8275), .B (n_3188), .Y (n_5742));
NOR2X1 g56098(.A (WX8275), .B (n_5500), .Y (n_9814));
NOR2X1 g55857(.A (WX3103), .B (n_5479), .Y (n_8538));
OAI21X1 g55957(.A0 (n_4247), .A1 (n_5841), .B0 (n_5708), .Y (n_5738));
NOR2X1 g56159(.A (WX9568), .B (n_3188), .Y (n_5737));
NOR2X1 g56161(.A (WX9568), .B (n_5427), .Y (n_6685));
NOR2X1 g55880(.A (WX3103), .B (n_1648), .Y (n_5735));
NOR2X1 g55993(.A (WX5689), .B (n_5712), .Y (n_5733));
NOR2X1 g55994(.A (WX5689), .B (n_5838), .Y (n_5732));
OAI21X1 g56724(.A0 (n_4450), .A1 (n_5729), .B0 (n_5707), .Y (n_5731));
OAI21X1 g56728(.A0 (n_3824), .A1 (n_5729), .B0 (n_5705), .Y (n_5730));
NAND2X1 g56882(.A (n_6575), .B (n_8334), .Y (n_5728));
INVX1 g56908(.A (DATA_9_11), .Y (n_5727));
NOR2X1 g56057(.A (WX6982), .B (n_1648), .Y (n_5725));
OAI21X1 g56060(.A0 (n_4405), .A1 (n_6686), .B0 (n_4860), .Y (n_5724));
OAI21X1 g56099(.A0 (n_5689), .A1 (n_9407), .B0 (n_5722), .Y (n_5723));
OAI21X1 g55859(.A0 (n_4449), .A1 (n_9815), .B0 (n_5566), .Y (n_5721));
OAI21X1 g56162(.A0 (n_5687), .A1 (n_9409), .B0 (n_4947), .Y (n_5720));
NOR2X1 g55986(.A (WX4398), .B (n_3188), .Y (n_5719));
NOR2X1 g55990(.A (WX4398), .B (n_5662), .Y (n_15856));
OAI21X1 g55995(.A0 (n_4248), .A1 (n_8539), .B0 (n_4860), .Y (n_5716));
NOR2X1 g56745(.A (WX10861), .B (n_1648), .Y (n_5714));
NOR2X1 g56746(.A (WX1810), .B (n_5712), .Y (n_5713));
NOR2X1 g56756(.A (WX1810), .B (n_5838), .Y (n_5711));
CLKBUFX1 gbuf_d_149(.A(n_5700), .Y(d_out_149));
CLKBUFX1 gbuf_q_149(.A(q_in_149), .Y(WX3267));
CLKBUFX1 gbuf_d_150(.A(n_5699), .Y(d_out_150));
CLKBUFX1 gbuf_q_150(.A(q_in_150), .Y(WX5853));
CLKBUFX1 gbuf_d_151(.A(n_5703), .Y(d_out_151));
CLKBUFX1 gbuf_q_151(.A(q_in_151), .Y(WX7146));
CLKBUFX1 gbuf_d_152(.A(n_5702), .Y(d_out_152));
CLKBUFX1 gbuf_q_152(.A(q_in_152), .Y(WX8439));
CLKBUFX1 gbuf_d_153(.A(n_5701), .Y(d_out_153));
CLKBUFX1 gbuf_q_153(.A(q_in_153), .Y(WX9732));
CLKBUFX1 gbuf_d_154(.A(n_6581), .Y(d_out_154));
CLKBUFX1 gbuf_q_154(.A(q_in_154), .Y(WX689));
OAI21X1 g56909(.A0 (n_5695), .A1 (n_5709), .B0 (n_4027), .Y(DATA_9_11));
CLKBUFX1 gbuf_d_155(.A(n_5693), .Y(d_out_155));
CLKBUFX1 gbuf_qn_155(.A(qn_in_155), .Y(WX6982));
INVX1 g56952(.A (WX523), .Y (n_5744));
CLKBUFX1 gbuf_d_156(.A(n_5690), .Y(d_out_156));
CLKBUFX1 gbuf_qn_156(.A(qn_in_156), .Y(WX8275));
CLKBUFX1 gbuf_d_157(.A(n_5688), .Y(d_out_157));
CLKBUFX1 gbuf_qn_157(.A(qn_in_157), .Y(WX9568));
OAI21X1 g55991(.A0 (n_5660), .A1 (n_9411), .B0 (n_4947), .Y (n_5708));
CLKBUFX1 gbuf_d_158(.A(n_5694), .Y(d_out_158));
CLKBUFX1 gbuf_qn_158(.A(qn_in_158), .Y(WX3103));
CLKBUFX1 gbuf_d_159(.A(n_5682), .Y(d_out_159));
CLKBUFX1 gbuf_qn_159(.A(qn_in_159), .Y(WX5689));
OAI21X1 g56757(.A0 (n_5664), .A1 (n_4162), .B0 (n_5706), .Y (n_5707));
OAI21X1 g56761(.A0 (n_4523), .A1 (n_7504), .B0 (n_5619), .Y (n_5705));
CLKBUFX1 gbuf_d_160(.A(n_5686), .Y(d_out_160));
CLKBUFX1 gbuf_q_160(.A(q_in_160), .Y(WX4562));
CLKBUFX1 gbuf_d_161(.A(n_6467), .Y(d_out_161));
CLKBUFX1 gbuf_q_161(.A(q_in_161), .Y(WX11025));
CLKBUFX1 gbuf_d_162(.A(n_5685), .Y(d_out_162));
CLKBUFX1 gbuf_q_162(.A(q_in_162), .Y(WX1974));
OAI21X1 g56906(.A0 (n_5676), .A1 (n_5889), .B0 (n_5608), .Y (n_8334));
CLKBUFX1 gbuf_d_163(.A(n_5674), .Y(d_out_163));
CLKBUFX1 gbuf_q_163(.A(q_in_163), .Y(WX523));
OAI21X1 g56077(.A0 (n_4121), .A1 (n_5235), .B0 (n_5670), .Y (n_5703));
OAI21X1 g56131(.A0 (n_4575), .A1 (n_5830), .B0 (n_5669), .Y (n_5702));
OAI21X1 g56191(.A0 (n_4269), .A1 (n_5834), .B0 (n_5667), .Y (n_5701));
CLKBUFX1 gbuf_d_164(.A(n_5661), .Y(d_out_164));
CLKBUFX1 gbuf_qn_164(.A(qn_in_164), .Y(WX4398));
OAI21X1 g55894(.A0 (n_4620), .A1 (n_5439), .B0 (n_5678), .Y (n_5700));
OAI21X1 g56017(.A0 (n_4404), .A1 (n_6106), .B0 (n_5658), .Y (n_5699));
CLKBUFX1 gbuf_d_165(.A(n_5666), .Y(d_out_165));
CLKBUFX1 gbuf_qn_165(.A(qn_in_165), .Y(WX10861));
CLKBUFX1 gbuf_d_166(.A(n_5665), .Y(d_out_166));
CLKBUFX1 gbuf_qn_166(.A(qn_in_166), .Y(WX1810));
NOR2X1 g55918(.A (WX3105), .B (n_5427), .Y (n_9815));
MX2X1 g56966(.A (n_5672), .B (WX525), .S0 (n_4026), .Y (n_5695));
NOR2X1 g55940(.A (WX3105), .B (n_5712), .Y (n_5694));
NOR2X1 g56116(.A (WX6984), .B (n_2851), .Y (n_5693));
NOR2X1 g56118(.A (WX6984), .B (n_5838), .Y (n_6686));
NOR2X1 g56153(.A (WX8277), .B (n_3690), .Y (n_5690));
NOR2X1 g56157(.A (WX8277), .B (n_5838), .Y (n_5689));
NOR2X1 g56218(.A (WX9570), .B (n_5712), .Y (n_5688));
NOR2X1 g56220(.A (WX9570), .B (n_5811), .Y (n_5687));
OAI21X1 g56016(.A0 (n_4245), .A1 (n_5535), .B0 (n_5654), .Y (n_5686));
OAI21X1 g56783(.A0 (n_4448), .A1 (n_5535), .B0 (n_5657), .Y (n_5685));
NOR2X1 g56052(.A (WX5691), .B (n_1648), .Y (n_5682));
NOR2X1 g56053(.A (WX5691), .B (n_5427), .Y (n_8539));
OAI21X1 g55919(.A0 (n_5638), .A1 (n_4447), .B0 (n_5460), .Y (n_5678));
INVX1 g56967(.A (DATA_9_10), .Y (n_5676));
NOR2X1 g56989(.A (n_5181), .B (n_5672), .Y (n_5674));
OR2X1 g56997(.A (n_5672), .B (n_5990), .Y (n_5671));
OAI21X1 g56119(.A0 (n_4403), .A1 (n_9816), .B0 (n_4947), .Y (n_5670));
OAI21X1 g56158(.A0 (n_15857), .A1 (n_15858), .B0 (n_7087), .Y(n_5669));
OAI21X1 g56221(.A0 (n_4574), .A1 (n_6687), .B0 (n_5460), .Y (n_5667));
NOR2X1 g56804(.A (WX10863), .B (n_1425), .Y (n_5666));
NOR2X1 g56805(.A (WX1812), .B (n_5712), .Y (n_5665));
NOR2X1 g56814(.A (WX1812), .B (n_5811), .Y (n_5664));
CLKBUFX1 gbuf_d_167(.A(n_5651), .Y(d_out_167));
CLKBUFX1 gbuf_q_167(.A(q_in_167), .Y(WX3269));
CLKBUFX1 gbuf_d_168(.A(n_5652), .Y(d_out_168));
CLKBUFX1 gbuf_q_168(.A(q_in_168), .Y(WX5855));
CLKBUFX1 gbuf_d_169(.A(n_5648), .Y(d_out_169));
CLKBUFX1 gbuf_q_169(.A(q_in_169), .Y(WX8441));
CLKBUFX1 gbuf_d_170(.A(n_5650), .Y(d_out_170));
CLKBUFX1 gbuf_q_170(.A(q_in_170), .Y(WX7148));
CLKBUFX1 gbuf_d_171(.A(n_5646), .Y(d_out_171));
CLKBUFX1 gbuf_q_171(.A(q_in_171), .Y(WX9734));
NOR2X1 g56818(.A (WX10863), .B (n_5662), .Y (n_7504));
NOR2X1 g56043(.A (WX4400), .B (n_2620), .Y (n_5661));
NOR2X1 g56049(.A (WX4400), .B (n_5811), .Y (n_5660));
OAI21X1 g56054(.A0 (n_5642), .A1 (n_11608), .B0 (n_3183), .Y(n_5658));
CLKBUFX1 gbuf_d_172(.A(n_5643), .Y(d_out_172));
CLKBUFX1 gbuf_qn_172(.A(qn_in_172), .Y(WX5691));
OAI21X1 g56968(.A0 (n_5628), .A1 (n_6091), .B0 (n_4021), .Y(DATA_9_10));
CLKBUFX1 gbuf_d_173(.A(n_5634), .Y(d_out_173));
CLKBUFX1 gbuf_qn_173(.A(qn_in_173), .Y(WX3105));
CLKBUFX1 gbuf_d_174(.A(n_5641), .Y(d_out_174));
CLKBUFX1 gbuf_qn_174(.A(qn_in_174), .Y(WX6984));
CLKBUFX1 gbuf_d_175(.A(n_5637), .Y(d_out_175));
CLKBUFX1 gbuf_qn_175(.A(qn_in_175), .Y(WX8277));
CLKBUFX1 gbuf_d_176(.A(n_5633), .Y(d_out_176));
CLKBUFX1 gbuf_qn_176(.A(qn_in_176), .Y(WX9570));
CLKBUFX1 gbuf_d_177(.A(n_5644), .Y(d_out_177));
CLKBUFX1 gbuf_q_177(.A(q_in_177), .Y(WX4564));
OAI21X1 g56816(.A0 (n_5616), .A1 (n_4160), .B0 (n_6497), .Y (n_5657));
CLKBUFX1 gbuf_d_178(.A(n_5629), .Y(d_out_178));
CLKBUFX1 gbuf_q_178(.A(q_in_178), .Y(WX11027));
CLKBUFX1 gbuf_d_179(.A(n_5631), .Y(d_out_179));
CLKBUFX1 gbuf_q_179(.A(q_in_179), .Y(WX1976));
CLKBUFX1 gbuf_d_180(.A(n_6541), .Y(d_out_180));
CLKBUFX1 gbuf_q_180(.A(q_in_180), .Y(WX691));
OAI21X1 g56050(.A0 (n_4316), .A1 (n_8547), .B0 (n_6497), .Y (n_5654));
CLKBUFX1 gbuf_d_181(.A(n_5627), .Y(d_out_181));
CLKBUFX1 gbuf_qn_181(.A(qn_in_181), .Y(WX4400));
OAI21X1 g56076(.A0 (n_4402), .A1 (n_5254), .B0 (n_5625), .Y (n_5652));
INVX1 g57013(.A (WX525), .Y (n_5672));
OAI21X1 g55953(.A0 (n_4317), .A1 (n_5649), .B0 (n_5622), .Y (n_5651));
OAI21X1 g56136(.A0 (n_4349), .A1 (n_5649), .B0 (n_5623), .Y (n_5650));
OAI21X1 g56190(.A0 (n_4299), .A1 (n_5841), .B0 (n_5621), .Y (n_5648));
OAI21X1 g56250(.A0 (n_4267), .A1 (n_5439), .B0 (n_5620), .Y (n_5646));
CLKBUFX1 gbuf_d_182(.A(n_5618), .Y(d_out_182));
CLKBUFX1 gbuf_qn_182(.A(qn_in_182), .Y(WX10863));
CLKBUFX1 gbuf_d_183(.A(n_5617), .Y(d_out_183));
CLKBUFX1 gbuf_qn_183(.A(qn_in_183), .Y(WX1812));
OAI21X1 g56075(.A0 (n_4472), .A1 (n_5493), .B0 (n_5606), .Y (n_5644));
CLKBUFX1 gbuf_d_184(.A(n_5610), .Y(d_out_184));
CLKBUFX1 gbuf_q_184(.A(q_in_184), .Y(WX525));
NOR2X1 g56111(.A (WX5693), .B (n_3188), .Y (n_5643));
NOR2X1 g56112(.A (WX5693), .B (n_5662), .Y (n_5642));
NOR2X1 g56175(.A (WX6986), .B (n_1648), .Y (n_5641));
NOR2X1 g56177(.A (WX6986), .B (n_5500), .Y (n_9816));
NOR2X1 g55977(.A (WX3107), .B (n_5811), .Y (n_5638));
NOR2X1 g56212(.A (WX8279), .B (n_1425), .Y (n_5637));
NOR2X1 g56216(.A (WX8279), .B (n_5811), .Y (n_15858));
NOR2X1 g55999(.A (WX3107), .B (n_3690), .Y (n_5634));
NOR2X1 g56277(.A (WX9572), .B (n_5181), .Y (n_5633));
NOR2X1 g56279(.A (WX9572), .B (n_4882), .Y (n_6687));
CLKBUFX1 gbuf_d_185(.A(n_5605), .Y(d_out_185));
CLKBUFX1 gbuf_q_185(.A(q_in_185), .Y(WX3235));
OAI21X1 g56843(.A0 (n_4229), .A1 (n_5630), .B0 (n_5604), .Y (n_5631));
OAI21X1 g56846(.A0 (n_3821), .A1 (n_5630), .B0 (n_5603), .Y (n_5629));
MX2X1 g57025(.A (n_5609), .B (WX527), .S0 (n_10739), .Y (n_5628));
NOR2X1 g56101(.A (WX4402), .B (n_1425), .Y (n_5627));
NOR2X1 g56108(.A (WX4402), .B (n_5052), .Y (n_8547));
OAI21X1 g56113(.A0 (n_4244), .A1 (n_8540), .B0 (n_5722), .Y (n_5625));
OAI21X1 g56178(.A0 (n_4401), .A1 (n_6683), .B0 (n_5619), .Y (n_5623));
OAI21X1 g55979(.A0 (n_4228), .A1 (n_9817), .B0 (n_4947), .Y (n_5622));
OAI21X1 g56217(.A0 (n_4348), .A1 (n_6688), .B0 (n_5566), .Y (n_5621));
OAI21X1 g56280(.A0 (n_4298), .A1 (n_9818), .B0 (n_5619), .Y (n_5620));
CLKBUFX1 gbuf_d_186(.A(n_5597), .Y(d_out_186));
CLKBUFX1 gbuf_q_186(.A(q_in_186), .Y(WX3271));
CLKBUFX1 gbuf_d_187(.A(n_5601), .Y(d_out_187));
CLKBUFX1 gbuf_q_187(.A(q_in_187), .Y(WX5857));
CLKBUFX1 gbuf_d_188(.A(n_5599), .Y(d_out_188));
CLKBUFX1 gbuf_q_188(.A(q_in_188), .Y(WX7150));
CLKBUFX1 gbuf_d_189(.A(n_5596), .Y(d_out_189));
CLKBUFX1 gbuf_q_189(.A(q_in_189), .Y(WX8443));
CLKBUFX1 gbuf_d_190(.A(n_5595), .Y(d_out_190));
CLKBUFX1 gbuf_q_190(.A(q_in_190), .Y(WX9736));
NOR2X1 g56863(.A (WX10865), .B (n_5712), .Y (n_5618));
NOR2X1 g56864(.A (WX1814), .B (n_3188), .Y (n_5617));
NOR2X1 g56874(.A (WX1814), .B (n_5052), .Y (n_5616));
INVX1 g57026(.A (DATA_9_9), .Y (n_5612));
NOR2X1 g57048(.A (n_1425), .B (n_5609), .Y (n_5610));
OR2X1 g57056(.A (n_5609), .B (n_4882), .Y (n_5608));
OAI21X1 g56109(.A0 (n_5568), .A1 (n_4314), .B0 (n_6479), .Y (n_5606));
CLKBUFX1 gbuf_d_191(.A(n_5591), .Y(d_out_191));
CLKBUFX1 gbuf_qn_191(.A(qn_in_191), .Y(WX5693));
CLKBUFX1 gbuf_d_192(.A(n_5588), .Y(d_out_192));
CLKBUFX1 gbuf_qn_192(.A(qn_in_192), .Y(WX6986));
CLKBUFX1 gbuf_d_193(.A(n_5584), .Y(d_out_193));
CLKBUFX1 gbuf_qn_193(.A(qn_in_193), .Y(WX8279));
CLKBUFX1 gbuf_d_194(.A(n_5594), .Y(d_out_194));
CLKBUFX1 gbuf_qn_194(.A(qn_in_194), .Y(WX3107));
CLKBUFX1 gbuf_d_195(.A(n_5592), .Y(d_out_195));
CLKBUFX1 gbuf_q_195(.A(q_in_195), .Y(WX4566));
CLKBUFX1 gbuf_d_196(.A(n_5577), .Y(d_out_196));
CLKBUFX1 gbuf_q_196(.A(q_in_196), .Y(WX11029));
CLKBUFX1 gbuf_d_197(.A(n_5579), .Y(d_out_197));
CLKBUFX1 gbuf_q_197(.A(q_in_197), .Y(WX1978));
CLKBUFX1 gbuf_d_198(.A(n_5578), .Y(d_out_198));
CLKBUFX1 gbuf_qn_198(.A(qn_in_198), .Y(WX9572));
OAI21X1 g56844(.A0 (n_4359), .A1 (n_5630), .B0 (n_5580), .Y (n_5605));
OAI21X1 g56877(.A0 (n_5573), .A1 (n_4158), .B0 (n_5460), .Y (n_5604));
OAI21X1 g56879(.A0 (n_4266), .A1 (n_7506), .B0 (n_4860), .Y (n_5603));
OAI21X1 g57027(.A0 (n_5554), .A1 (n_5843), .B0 (n_4019), .Y(DATA_9_9));
CLKBUFX1 gbuf_d_199(.A(n_5569), .Y(d_out_199));
CLKBUFX1 gbuf_qn_199(.A(qn_in_199), .Y(WX4402));
OAI21X1 g56135(.A0 (n_4400), .A1 (n_5600), .B0 (n_5567), .Y (n_5601));
OAI21X1 g56195(.A0 (n_4119), .A1 (n_5598), .B0 (n_5565), .Y (n_5599));
OAI21X1 g56012(.A0 (n_4315), .A1 (n_5841), .B0 (n_5563), .Y (n_5597));
OAI21X1 g56249(.A0 (n_4573), .A1 (n_5841), .B0 (n_5564), .Y (n_5596));
CLKBUFX1 gbuf_d_200(.A(n_6589), .Y(d_out_200));
CLKBUFX1 gbuf_q_200(.A(q_in_200), .Y(WX693));
OAI21X1 g56309(.A0 (n_4518), .A1 (n_4803), .B0 (n_5562), .Y (n_5595));
CLKBUFX1 gbuf_d_201(.A(n_5560), .Y(d_out_201));
CLKBUFX1 gbuf_qn_201(.A(qn_in_201), .Y(WX10865));
CLKBUFX1 gbuf_d_202(.A(n_5558), .Y(d_out_202));
CLKBUFX1 gbuf_qn_202(.A(qn_in_202), .Y(WX1814));
NOR2X1 g56058(.A (WX3109), .B (n_1648), .Y (n_5594));
INVX1 g57072(.A (WX527), .Y (n_5609));
OAI21X1 g56134(.A0 (n_4243), .A1 (n_5600), .B0 (n_5553), .Y (n_5592));
NOR2X1 g56170(.A (WX5695), .B (n_1648), .Y (n_5591));
NOR2X1 g56171(.A (WX5695), .B (n_5479), .Y (n_8540));
NOR2X1 g56234(.A (WX6988), .B (n_1648), .Y (n_5588));
NOR2X1 g56236(.A (WX6988), .B (n_5500), .Y (n_6683));
NOR2X1 g56271(.A (WX8281), .B (n_5712), .Y (n_5584));
NOR2X1 g56275(.A (WX8281), .B (n_5427), .Y (n_6688));
CLKBUFX1 gbuf_d_203(.A(n_5551), .Y(d_out_203));
CLKBUFX1 gbuf_q_203(.A(q_in_203), .Y(WX4528));
CLKBUFX1 gbuf_d_204(.A(n_5550), .Y(d_out_204));
CLKBUFX1 gbuf_q_204(.A(q_in_204), .Y(WX3237));
NOR2X1 g56037(.A (WX3109), .B (n_5479), .Y (n_9817));
OAI21X1 g56886(.A0 (n_5547), .A1 (n_4282), .B0 (n_4947), .Y (n_5580));
OAI21X1 g56901(.A0 (n_4227), .A1 (n_5535), .B0 (n_5557), .Y (n_5579));
NOR2X1 g56336(.A (WX9574), .B (n_1648), .Y (n_5578));
OAI21X1 g56905(.A0 (n_3817), .A1 (n_5576), .B0 (n_5555), .Y (n_5577));
NOR2X1 g56338(.A (WX9574), .B (n_5427), .Y (n_9818));
NOR2X1 g56935(.A (WX1816), .B (n_5479), .Y (n_5573));
NOR2X1 g56937(.A (WX10867), .B (n_5479), .Y (n_7506));
CLKBUFX1 gbuf_d_205(.A(n_5541), .Y(d_out_205));
CLKBUFX1 gbuf_q_205(.A(q_in_205), .Y(WX527));
NOR2X1 g56160(.A (WX4404), .B (n_1425), .Y (n_5569));
NOR2X1 g56167(.A (WX4404), .B (n_5662), .Y (n_5568));
OAI21X1 g56172(.A0 (n_5518), .A1 (n_9427), .B0 (n_5566), .Y (n_5567));
OAI21X1 g56237(.A0 (n_4399), .A1 (n_9819), .B0 (n_5275), .Y (n_5565));
OAI21X1 g56276(.A0 (n_5513), .A1 (n_11614), .B0 (n_5619), .Y(n_5564));
CLKBUFX1 gbuf_d_206(.A(n_5546), .Y(d_out_206));
CLKBUFX1 gbuf_q_206(.A(q_in_206), .Y(WX3273));
CLKBUFX1 gbuf_d_207(.A(n_5537), .Y(d_out_207));
CLKBUFX1 gbuf_q_207(.A(q_in_207), .Y(WX5859));
CLKBUFX1 gbuf_d_208(.A(n_5536), .Y(d_out_208));
CLKBUFX1 gbuf_q_208(.A(q_in_208), .Y(WX7152));
CLKBUFX1 gbuf_d_209(.A(n_5534), .Y(d_out_209));
CLKBUFX1 gbuf_q_209(.A(q_in_209), .Y(WX8445));
CLKBUFX1 gbuf_d_210(.A(n_5545), .Y(d_out_210));
CLKBUFX1 gbuf_q_210(.A(q_in_210), .Y(WX9738));
CLKBUFX1 gbuf_d_211(.A(n_5548), .Y(d_out_211));
CLKBUFX1 gbuf_qn_211(.A(qn_in_211), .Y(WX3073));
OAI21X1 g56038(.A0 (n_5525), .A1 (n_11612), .B0 (n_5566), .Y(n_5563));
OAI21X1 g56339(.A0 (n_4572), .A1 (n_9820), .B0 (n_4947), .Y (n_5562));
NOR2X1 g56921(.A (WX10867), .B (n_3690), .Y (n_5560));
NOR2X1 g56922(.A (WX1816), .B (n_2605), .Y (n_5558));
OAI21X1 g56936(.A0 (n_5509), .A1 (n_4156), .B0 (n_5556), .Y (n_5557));
OAI21X1 g56938(.A0 (n_4517), .A1 (n_7505), .B0 (n_4860), .Y (n_5555));
CLKBUFX1 gbuf_d_212(.A(n_5528), .Y(d_out_212));
CLKBUFX1 gbuf_qn_212(.A(qn_in_212), .Y(WX9574));
CLKBUFX1 gbuf_d_213(.A(n_5523), .Y(d_out_213));
CLKBUFX1 gbuf_qn_213(.A(qn_in_213), .Y(WX3109));
MX2X1 g57084(.A (n_5540), .B (WX529), .S0 (n_4018), .Y (n_5554));
OAI21X1 g56168(.A0 (n_4310), .A1 (n_8548), .B0 (n_5460), .Y (n_5553));
CLKBUFX1 gbuf_d_214(.A(n_5519), .Y(d_out_214));
CLKBUFX1 gbuf_qn_214(.A(qn_in_214), .Y(WX5695));
CLKBUFX1 gbuf_d_215(.A(n_5517), .Y(d_out_215));
CLKBUFX1 gbuf_qn_215(.A(qn_in_215), .Y(WX6988));
CLKBUFX1 gbuf_d_216(.A(n_5521), .Y(d_out_216));
CLKBUFX1 gbuf_q_216(.A(q_in_216), .Y(WX4568));
CLKBUFX1 gbuf_d_217(.A(n_5529), .Y(d_out_217));
CLKBUFX1 gbuf_q_217(.A(q_in_217), .Y(WX11031));
CLKBUFX1 gbuf_d_218(.A(n_5530), .Y(d_out_218));
CLKBUFX1 gbuf_q_218(.A(q_in_218), .Y(WX1980));
CLKBUFX1 gbuf_d_219(.A(n_5514), .Y(d_out_219));
CLKBUFX1 gbuf_qn_219(.A(qn_in_219), .Y(WX8281));
OAI21X1 g56898(.A0 (n_4520), .A1 (n_5334), .B0 (n_5533), .Y (n_5551));
OAI21X1 g56903(.A0 (n_4355), .A1 (n_5549), .B0 (n_5532), .Y (n_5550));
NOR2X1 g56943(.A (WX3075), .B (n_5181), .Y (n_5548));
NOR2X1 g56944(.A (WX3075), .B (n_5427), .Y (n_5547));
CLKBUFX1 gbuf_d_220(.A(n_5512), .Y(d_out_220));
CLKBUFX1 gbuf_qn_220(.A(qn_in_220), .Y(WX10867));
CLKBUFX1 gbuf_d_221(.A(n_5511), .Y(d_out_221));
CLKBUFX1 gbuf_qn_221(.A(qn_in_221), .Y(WX1816));
OAI21X1 g56071(.A0 (n_4311), .A1 (n_5185), .B0 (n_5505), .Y (n_5546));
OAI21X1 g56368(.A0 (n_4516), .A1 (n_4866), .B0 (n_5507), .Y (n_5545));
INVX1 g57085(.A (DATA_9_8), .Y (n_5543));
NOR2X1 g57107(.A (n_1425), .B (n_5540), .Y (n_5541));
OR2X1 g57115(.A (n_5540), .B (n_3828), .Y (n_5539));
CLKBUFX1 gbuf_d_222(.A(n_5503), .Y(d_out_222));
CLKBUFX1 gbuf_qn_222(.A(qn_in_222), .Y(WX4404));
OAI21X1 g56194(.A0 (n_4220), .A1 (n_5490), .B0 (n_5499), .Y (n_5537));
OAI21X1 g56254(.A0 (n_4345), .A1 (n_5535), .B0 (n_5497), .Y (n_5536));
OAI21X1 g56308(.A0 (n_4293), .A1 (n_5845), .B0 (n_5496), .Y (n_5534));
OAI21X1 g56928(.A0 (n_5480), .A1 (n_4358), .B0 (n_5722), .Y (n_5533));
OAI21X1 g56945(.A0 (n_5477), .A1 (n_4557), .B0 (n_3183), .Y (n_5532));
OAI21X1 g56960(.A0 (n_4425), .A1 (n_5535), .B0 (n_5489), .Y (n_5530));
OAI21X1 g56964(.A0 (n_3816), .A1 (n_5474), .B0 (n_5488), .Y (n_5529));
NOR2X1 g56395(.A (WX9576), .B (n_1648), .Y (n_5528));
NOR2X1 g56398(.A (WX9576), .B (n_5427), .Y (n_9820));
NOR2X1 g56096(.A (WX3111), .B (n_3218), .Y (n_5525));
OAI21X1 g57086(.A0 (n_5473), .A1 (n_5965), .B0 (n_4080), .Y(DATA_9_8));
NOR2X1 g56117(.A (WX3111), .B (n_5712), .Y (n_5523));
OAI21X1 g56193(.A0 (n_4469), .A1 (n_5235), .B0 (n_5485), .Y (n_5521));
NOR2X1 g56229(.A (WX5697), .B (n_1425), .Y (n_5519));
NOR2X1 g56230(.A (WX5697), .B (n_5500), .Y (n_5518));
NOR2X1 g56293(.A (WX6990), .B (n_2620), .Y (n_5517));
CLKBUFX1 gbuf_d_223(.A(n_5492), .Y(d_out_223));
CLKBUFX1 gbuf_q_223(.A(q_in_223), .Y(WX5821));
CLKBUFX1 gbuf_d_224(.A(n_5494), .Y(d_out_224));
CLKBUFX1 gbuf_q_224(.A(q_in_224), .Y(WX4530));
CLKBUFX1 gbuf_d_225(.A(n_5491), .Y(d_out_225));
CLKBUFX1 gbuf_q_225(.A(q_in_225), .Y(WX3239));
CLKBUFX1 gbuf_d_226(.A(n_5486), .Y(d_out_226));
CLKBUFX1 gbuf_q_226(.A(q_in_226), .Y(WX695));
NOR2X1 g56295(.A (WX6990), .B (n_5500), .Y (n_9819));
NOR2X1 g56330(.A (WX8283), .B (n_5712), .Y (n_5514));
NOR2X1 g56334(.A (WX8283), .B (n_5500), .Y (n_5513));
CLKBUFX1 gbuf_d_227(.A(n_5478), .Y(d_out_227));
CLKBUFX1 gbuf_qn_227(.A(qn_in_227), .Y(WX3075));
NOR2X1 g56980(.A (WX10869), .B (n_2849), .Y (n_5512));
NOR2X1 g56981(.A (WX1818), .B (n_2849), .Y (n_5511));
NOR2X1 g56993(.A (WX1818), .B (n_5838), .Y (n_5509));
NOR2X1 g56995(.A (WX10869), .B (n_5662), .Y (n_7505));
OAI21X1 g56397(.A0 (n_4292), .A1 (n_8549), .B0 (n_5722), .Y (n_5507));
OAI21X1 g56097(.A0 (n_4424), .A1 (n_9821), .B0 (n_5722), .Y (n_5505));
INVX1 g57123(.A (WX529), .Y (n_5540));
NOR2X1 g56219(.A (WX4406), .B (n_2851), .Y (n_5503));
NOR2X1 g56226(.A (WX4406), .B (n_5500), .Y (n_8548));
OAI21X1 g56231(.A0 (n_5437), .A1 (n_11616), .B0 (n_4947), .Y(n_5499));
CLKBUFX1 gbuf_d_228(.A(n_5472), .Y(d_out_228));
CLKBUFX1 gbuf_q_228(.A(q_in_228), .Y(WX3275));
CLKBUFX1 gbuf_d_229(.A(n_5471), .Y(d_out_229));
CLKBUFX1 gbuf_q_229(.A(q_in_229), .Y(WX5861));
CLKBUFX1 gbuf_d_230(.A(n_5469), .Y(d_out_230));
CLKBUFX1 gbuf_q_230(.A(q_in_230), .Y(WX7154));
CLKBUFX1 gbuf_d_231(.A(n_5483), .Y(d_out_231));
CLKBUFX1 gbuf_q_231(.A(q_in_231), .Y(WX8447));
CLKBUFX1 gbuf_d_232(.A(n_5475), .Y(d_out_232));
CLKBUFX1 gbuf_q_232(.A(q_in_232), .Y(WX9740));
CLKBUFX1 gbuf_d_233(.A(n_5481), .Y(d_out_233));
CLKBUFX1 gbuf_qn_233(.A(qn_in_233), .Y(WX4366));
OAI21X1 g56296(.A0 (n_5465), .A1 (n_4219), .B0 (n_4947), .Y (n_5497));
OAI21X1 g56335(.A0 (n_5459), .A1 (n_9429), .B0 (n_5460), .Y (n_5496));
CLKBUFX1 gbuf_d_234(.A(n_5462), .Y(d_out_234));
CLKBUFX1 gbuf_qn_234(.A(qn_in_234), .Y(WX8283));
OAI21X1 g56957(.A0 (n_4508), .A1 (n_5493), .B0 (n_5464), .Y (n_5494));
OAI21X1 g56959(.A0 (n_4442), .A1 (n_5415), .B0 (n_5463), .Y (n_5492));
OAI21X1 g56962(.A0 (n_4351), .A1 (n_5490), .B0 (n_5461), .Y (n_5491));
OAI21X1 g56994(.A0 (n_5429), .A1 (n_4154), .B0 (n_5722), .Y (n_5489));
OAI21X1 g56996(.A0 (n_4515), .A1 (n_6678), .B0 (n_4860), .Y (n_5488));
CLKBUFX1 gbuf_d_235(.A(n_5453), .Y(d_out_235));
CLKBUFX1 gbuf_qn_235(.A(qn_in_235), .Y(WX9576));
NAND2X1 g57081(.A (n_5454), .B (n_4698), .Y (n_5486));
CLKBUFX1 gbuf_d_236(.A(n_5448), .Y(d_out_236));
CLKBUFX1 gbuf_q_236(.A(q_in_236), .Y(WX529));
CLKBUFX1 gbuf_d_237(.A(n_5442), .Y(d_out_237));
CLKBUFX1 gbuf_qn_237(.A(qn_in_237), .Y(WX3111));
OAI21X1 g56227(.A0 (n_4308), .A1 (n_8550), .B0 (n_5556), .Y (n_5485));
CLKBUFX1 gbuf_d_238(.A(n_5438), .Y(d_out_238));
CLKBUFX1 gbuf_qn_238(.A(qn_in_238), .Y(WX5697));
CLKBUFX1 gbuf_d_239(.A(n_5440), .Y(d_out_239));
CLKBUFX1 gbuf_q_239(.A(q_in_239), .Y(WX4570));
CLKBUFX1 gbuf_d_240(.A(n_5456), .Y(d_out_240));
CLKBUFX1 gbuf_q_240(.A(q_in_240), .Y(WX11033));
CLKBUFX1 gbuf_d_241(.A(n_5458), .Y(d_out_241));
CLKBUFX1 gbuf_q_241(.A(q_in_241), .Y(WX1982));
CLKBUFX1 gbuf_d_242(.A(n_5467), .Y(d_out_242));
CLKBUFX1 gbuf_qn_242(.A(qn_in_242), .Y(WX6990));
OAI21X1 g56367(.A0 (n_4291), .A1 (n_5482), .B0 (n_5434), .Y (n_5483));
NOR2X1 g56983(.A (WX4368), .B (n_5181), .Y (n_5481));
NOR2X1 g56985(.A (WX4368), .B (n_5479), .Y (n_5480));
NOR2X1 g57002(.A (WX3077), .B (n_5181), .Y (n_5478));
NOR2X1 g57003(.A (WX3077), .B (n_5662), .Y (n_5477));
CLKBUFX1 gbuf_d_243(.A(n_5432), .Y(d_out_243));
CLKBUFX1 gbuf_qn_243(.A(qn_in_243), .Y(WX10869));
CLKBUFX1 gbuf_d_244(.A(n_5430), .Y(d_out_244));
CLKBUFX1 gbuf_qn_244(.A(qn_in_244), .Y(WX1818));
OAI21X1 g56427(.A0 (n_4514), .A1 (n_5474), .B0 (n_5426), .Y (n_5475));
MX2X1 g57143(.A (n_5446), .B (WX531), .S0 (n_4079), .Y (n_5473));
OAI21X1 g56130(.A0 (n_4309), .A1 (n_5105), .B0 (n_5425), .Y (n_5472));
CLKBUFX1 gbuf_d_245(.A(n_5424), .Y(d_out_245));
CLKBUFX1 gbuf_qn_245(.A(qn_in_245), .Y(WX4406));
OAI21X1 g56253(.A0 (n_4218), .A1 (n_4803), .B0 (n_5421), .Y (n_5471));
OAI21X1 g56313(.A0 (n_4117), .A1 (n_5468), .B0 (n_5436), .Y (n_5469));
NOR2X1 g56352(.A (WX6992), .B (n_2851), .Y (n_5467));
NOR2X1 g56354(.A (WX6992), .B (n_5052), .Y (n_5465));
OAI21X1 g56986(.A0 (n_4354), .A1 (n_6191), .B0 (n_5722), .Y (n_5464));
OAI21X1 g56992(.A0 (n_5403), .A1 (n_4519), .B0 (n_3183), .Y (n_5463));
NOR2X1 g56389(.A (WX8285), .B (n_1425), .Y (n_5462));
OAI21X1 g57004(.A0 (n_4555), .A1 (n_6673), .B0 (n_5460), .Y (n_5461));
NOR2X1 g56393(.A (WX8285), .B (n_5500), .Y (n_5459));
OAI21X1 g57019(.A0 (n_4418), .A1 (n_5415), .B0 (n_5414), .Y (n_5458));
OAI21X1 g57023(.A0 (n_3815), .A1 (n_5892), .B0 (n_5413), .Y (n_5456));
NAND2X1 g57117(.A (n_5411), .B (n_6615), .Y (n_5454));
NOR2X1 g56454(.A (WX9578), .B (n_5181), .Y (n_5453));
NOR2X1 g56456(.A (WX9578), .B (n_5427), .Y (n_8549));
INVX1 g57144(.A (DATA_9_7), .Y (n_5450));
NOR2X1 g57167(.A (n_1425), .B (n_5446), .Y (n_5448));
OR2X1 g57175(.A (n_5446), .B (n_4882), .Y (n_5445));
NOR2X1 g56155(.A (WX3113), .B (n_5500), .Y (n_9821));
NOR2X1 g56176(.A (WX3113), .B (n_5712), .Y (n_5442));
OAI21X1 g56252(.A0 (n_4466), .A1 (n_5439), .B0 (n_5410), .Y (n_5440));
NOR2X1 g56288(.A (WX5699), .B (n_1648), .Y (n_5438));
NOR2X1 g56289(.A (WX5699), .B (n_3218), .Y (n_5437));
CLKBUFX1 gbuf_d_246(.A(n_5419), .Y(d_out_246));
CLKBUFX1 gbuf_q_246(.A(q_in_246), .Y(WX5823));
CLKBUFX1 gbuf_d_247(.A(n_5420), .Y(d_out_247));
CLKBUFX1 gbuf_q_247(.A(q_in_247), .Y(WX4532));
CLKBUFX1 gbuf_d_248(.A(n_5417), .Y(d_out_248));
CLKBUFX1 gbuf_q_248(.A(q_in_248), .Y(WX7114));
CLKBUFX1 gbuf_d_249(.A(n_5416), .Y(d_out_249));
CLKBUFX1 gbuf_q_249(.A(q_in_249), .Y(WX3241));
OAI21X1 g56355(.A0 (n_5386), .A1 (n_11618), .B0 (n_5722), .Y(n_5436));
CLKBUFX1 gbuf_d_250(.A(n_5407), .Y(d_out_250));
CLKBUFX1 gbuf_qn_250(.A(qn_in_250), .Y(WX4368));
CLKBUFX1 gbuf_d_251(.A(n_5401), .Y(d_out_251));
CLKBUFX1 gbuf_qn_251(.A(qn_in_251), .Y(WX3077));
OAI21X1 g56394(.A0 (n_4116), .A1 (n_8551), .B0 (n_4860), .Y (n_5434));
NOR2X1 g57040(.A (WX10871), .B (n_3188), .Y (n_5432));
NOR2X1 g57041(.A (WX1820), .B (n_1648), .Y (n_5430));
NOR2X1 g57052(.A (WX1820), .B (n_5838), .Y (n_5429));
NOR2X1 g57054(.A (WX10871), .B (n_5427), .Y (n_6678));
OAI21X1 g56457(.A0 (n_4290), .A1 (n_8552), .B0 (n_5722), .Y (n_5426));
OAI21X1 g57145(.A0 (n_5377), .A1 (n_5965), .B0 (n_4077), .Y(DATA_9_7));
OAI21X1 g56156(.A0 (n_4417), .A1 (n_6689), .B0 (n_5722), .Y (n_5425));
NOR2X1 g56278(.A (WX4408), .B (n_5181), .Y (n_5424));
NOR2X1 g56284(.A (WX4408), .B (n_3218), .Y (n_8550));
OAI21X1 g56290(.A0 (n_4467), .A1 (n_6690), .B0 (n_4947), .Y (n_5421));
CLKBUFX1 gbuf_d_252(.A(n_5395), .Y(d_out_252));
CLKBUFX1 gbuf_q_252(.A(q_in_252), .Y(WX3277));
CLKBUFX1 gbuf_d_253(.A(n_5394), .Y(d_out_253));
CLKBUFX1 gbuf_q_253(.A(q_in_253), .Y(WX5863));
CLKBUFX1 gbuf_d_254(.A(n_5409), .Y(d_out_254));
CLKBUFX1 gbuf_q_254(.A(q_in_254), .Y(WX7156));
CLKBUFX1 gbuf_d_255(.A(n_5398), .Y(d_out_255));
CLKBUFX1 gbuf_q_255(.A(q_in_255), .Y(WX8449));
CLKBUFX1 gbuf_d_256(.A(n_5396), .Y(d_out_256));
CLKBUFX1 gbuf_q_256(.A(q_in_256), .Y(WX9742));
CLKBUFX1 gbuf_d_257(.A(n_5404), .Y(d_out_257));
CLKBUFX1 gbuf_qn_257(.A(qn_in_257), .Y(WX5659));
CLKBUFX1 gbuf_d_258(.A(n_5397), .Y(d_out_258));
CLKBUFX1 gbuf_q_258(.A(q_in_258), .Y(WX697));
CLKBUFX1 gbuf_d_259(.A(n_5388), .Y(d_out_259));
CLKBUFX1 gbuf_qn_259(.A(qn_in_259), .Y(WX6992));
OAI21X1 g57017(.A0 (n_4502), .A1 (n_5841), .B0 (n_5390), .Y (n_5420));
OAI21X1 g57018(.A0 (n_4440), .A1 (n_5418), .B0 (n_5389), .Y (n_5419));
OAI21X1 g57020(.A0 (n_4381), .A1 (n_5439), .B0 (n_5385), .Y (n_5417));
OAI21X1 g57021(.A0 (n_4347), .A1 (n_5415), .B0 (n_5384), .Y (n_5416));
OAI21X1 g57053(.A0 (n_5365), .A1 (n_4152), .B0 (n_5556), .Y (n_5414));
OAI21X1 g57055(.A0 (n_4513), .A1 (n_6679), .B0 (n_4860), .Y (n_5413));
CLKBUFX1 gbuf_d_260(.A(n_5380), .Y(d_out_260));
CLKBUFX1 gbuf_qn_260(.A(qn_in_260), .Y(WX8285));
OAI21X1 g57142(.A0 (n_5360), .A1 (n_5889), .B0 (n_5256), .Y (n_5411));
CLKBUFX1 gbuf_d_261(.A(n_5376), .Y(d_out_261));
CLKBUFX1 gbuf_qn_261(.A(qn_in_261), .Y(WX9578));
INVX1 g57184(.A (WX531), .Y (n_5446));
CLKBUFX1 gbuf_d_262(.A(n_5371), .Y(d_out_262));
CLKBUFX1 gbuf_qn_262(.A(qn_in_262), .Y(WX3113));
CLKBUFX1 gbuf_d_263(.A(n_6486), .Y(d_out_263));
CLKBUFX1 gbuf_q_263(.A(q_in_263), .Y(WX11035));
OAI21X1 g56286(.A0 (n_15851), .A1 (n_15852), .B0 (n_5722), .Y(n_5410));
CLKBUFX1 gbuf_d_264(.A(n_5370), .Y(d_out_264));
CLKBUFX1 gbuf_q_264(.A(q_in_264), .Y(WX4572));
CLKBUFX1 gbuf_d_265(.A(n_5382), .Y(d_out_265));
CLKBUFX1 gbuf_q_265(.A(q_in_265), .Y(WX1984));
CLKBUFX1 gbuf_d_266(.A(n_5392), .Y(d_out_266));
CLKBUFX1 gbuf_qn_266(.A(qn_in_266), .Y(WX5699));
OAI21X1 g56372(.A0 (n_4341), .A1 (n_5105), .B0 (n_5368), .Y (n_5409));
NOR2X1 g57042(.A (WX4370), .B (n_1648), .Y (n_5407));
NOR2X1 g57045(.A (WX4370), .B (n_5662), .Y (n_6191));
NOR2X1 g57049(.A (WX5661), .B (n_1648), .Y (n_5404));
NOR2X1 g57050(.A (WX5661), .B (n_5838), .Y (n_5403));
NOR2X1 g57061(.A (WX3079), .B (n_5181), .Y (n_5401));
NOR2X1 g57062(.A (WX3079), .B (n_5479), .Y (n_6673));
CLKBUFX1 gbuf_d_267(.A(n_5367), .Y(d_out_267));
CLKBUFX1 gbuf_qn_267(.A(qn_in_267), .Y(WX10871));
CLKBUFX1 gbuf_d_268(.A(n_5366), .Y(d_out_268));
CLKBUFX1 gbuf_qn_268(.A(qn_in_268), .Y(WX1820));
OAI21X1 g56426(.A0 (n_4289), .A1 (n_5105), .B0 (n_5362), .Y (n_5398));
NAND2X2 g57140(.A (n_5361), .B (n_4695), .Y (n_5397));
CLKBUFX1 gbuf_d_269(.A(n_5358), .Y(d_out_269));
CLKBUFX1 gbuf_q_269(.A(q_in_269), .Y(WX531));
OAI21X1 g56486(.A0 (n_4512), .A1 (n_5649), .B0 (n_5354), .Y (n_5396));
OAI21X1 g56189(.A0 (n_4307), .A1 (n_5841), .B0 (n_5353), .Y (n_5395));
CLKBUFX1 gbuf_d_270(.A(n_5352), .Y(d_out_270));
CLKBUFX1 gbuf_qn_270(.A(qn_in_270), .Y(WX4408));
OAI21X1 g56312(.A0 (n_4396), .A1 (n_5393), .B0 (n_5369), .Y (n_5394));
NOR2X1 g56347(.A (WX5701), .B (n_1425), .Y (n_5392));
NOR2X1 g56348(.A (WX5701), .B (n_5479), .Y (n_6690));
OAI21X1 g57047(.A0 (n_5331), .A1 (n_4350), .B0 (n_5556), .Y (n_5390));
OAI21X1 g57051(.A0 (n_4507), .A1 (n_6666), .B0 (n_4860), .Y (n_5389));
NOR2X1 g56411(.A (WX6994), .B (n_5181), .Y (n_5388));
NOR2X1 g56413(.A (WX6994), .B (n_5838), .Y (n_5386));
OAI21X1 g57060(.A0 (n_4441), .A1 (n_6192), .B0 (n_5722), .Y (n_5385));
OAI21X1 g57063(.A0 (n_4553), .A1 (n_6193), .B0 (n_4860), .Y (n_5384));
OAI21X1 g57078(.A0 (n_4225), .A1 (n_5918), .B0 (n_5342), .Y (n_5382));
NOR2X1 g56448(.A (WX8287), .B (n_1425), .Y (n_5380));
NOR2X1 g56452(.A (WX8287), .B (n_5838), .Y (n_8551));
MX2X1 g57204(.A (n_5356), .B (WX533), .S0 (n_4076), .Y (n_5377));
NOR2X1 g56513(.A (WX9580), .B (n_1648), .Y (n_5376));
NOR2X1 g56515(.A (WX9580), .B (n_5427), .Y (n_8552));
CLKBUFX1 gbuf_d_271(.A(n_5347), .Y(d_out_271));
CLKBUFX1 gbuf_q_271(.A(q_in_271), .Y(WX5825));
NOR2X1 g56214(.A (WX3115), .B (n_5811), .Y (n_6689));
NOR2X1 g56235(.A (WX3115), .B (n_5181), .Y (n_5371));
CLKBUFX1 gbuf_d_272(.A(n_5350), .Y(d_out_272));
CLKBUFX1 gbuf_q_272(.A(q_in_272), .Y(WX8407));
CLKBUFX1 gbuf_d_273(.A(n_5348), .Y(d_out_273));
CLKBUFX1 gbuf_q_273(.A(q_in_273), .Y(WX4534));
CLKBUFX1 gbuf_d_274(.A(n_5345), .Y(d_out_274));
CLKBUFX1 gbuf_q_274(.A(q_in_274), .Y(WX7116));
CLKBUFX1 gbuf_d_275(.A(n_5343), .Y(d_out_275));
CLKBUFX1 gbuf_q_275(.A(q_in_275), .Y(WX3243));
OAI21X1 g56311(.A0 (n_4462), .A1 (n_5393), .B0 (n_5338), .Y (n_5370));
OAI21X1 g56349(.A0 (n_4465), .A1 (n_6691), .B0 (n_5460), .Y (n_5369));
OAI21X1 g56414(.A0 (n_4395), .A1 (n_6692), .B0 (n_5722), .Y (n_5368));
CLKBUFX1 gbuf_d_276(.A(n_5333), .Y(d_out_276));
CLKBUFX1 gbuf_qn_276(.A(qn_in_276), .Y(WX4370));
CLKBUFX1 gbuf_d_277(.A(n_5330), .Y(d_out_277));
CLKBUFX1 gbuf_qn_277(.A(qn_in_277), .Y(WX5661));
CLKBUFX1 gbuf_d_278(.A(n_5325), .Y(d_out_278));
CLKBUFX1 gbuf_qn_278(.A(qn_in_278), .Y(WX3079));
NOR2X1 g57099(.A (WX10873), .B (n_1648), .Y (n_5367));
NOR2X1 g57100(.A (WX1822), .B (n_1425), .Y (n_5366));
NOR2X1 g57111(.A (WX1822), .B (n_5662), .Y (n_5365));
NOR2X1 g57113(.A (WX10873), .B (n_5662), .Y (n_6679));
OAI21X1 g56453(.A0 (n_4340), .A1 (n_9822), .B0 (n_5566), .Y (n_5362));
NAND2X1 g57177(.A (n_6575), .B (n_8335), .Y (n_5361));
INVX1 g57205(.A (DATA_9_6), .Y (n_5360));
NOR2X1 g57227(.A (n_1425), .B (n_5356), .Y (n_5358));
OR2X1 g57236(.A (n_5356), .B (n_5968), .Y (n_5355));
OAI21X1 g56516(.A0 (n_4288), .A1 (n_9823), .B0 (n_5566), .Y (n_5354));
OAI21X1 g56215(.A0 (n_5294), .A1 (n_4224), .B0 (n_4860), .Y (n_5353));
CLKBUFX1 gbuf_d_279(.A(n_5319), .Y(d_out_279));
CLKBUFX1 gbuf_q_279(.A(q_in_279), .Y(WX3279));
CLKBUFX1 gbuf_d_280(.A(n_5336), .Y(d_out_280));
CLKBUFX1 gbuf_q_280(.A(q_in_280), .Y(WX5865));
CLKBUFX1 gbuf_d_281(.A(n_5335), .Y(d_out_281));
CLKBUFX1 gbuf_q_281(.A(q_in_281), .Y(WX7158));
CLKBUFX1 gbuf_d_282(.A(n_5323), .Y(d_out_282));
CLKBUFX1 gbuf_q_282(.A(q_in_282), .Y(WX8451));
CLKBUFX1 gbuf_d_283(.A(n_5321), .Y(d_out_283));
CLKBUFX1 gbuf_q_283(.A(q_in_283), .Y(WX9744));
CLKBUFX1 gbuf_d_284(.A(n_5328), .Y(d_out_284));
CLKBUFX1 gbuf_qn_284(.A(qn_in_284), .Y(WX6952));
NOR2X1 g56337(.A (WX4410), .B (n_5712), .Y (n_5352));
NOR2X1 g56343(.A (WX4410), .B (n_5662), .Y (n_15852));
CLKBUFX1 gbuf_d_285(.A(n_5316), .Y(d_out_285));
CLKBUFX1 gbuf_qn_285(.A(qn_in_285), .Y(WX5701));
CLKBUFX1 gbuf_d_286(.A(n_5304), .Y(d_out_286));
CLKBUFX1 gbuf_qn_286(.A(qn_in_286), .Y(WX6994));
OAI21X1 g57074(.A0 (n_4616), .A1 (n_5439), .B0 (n_5314), .Y (n_5350));
OAI21X1 g57076(.A0 (n_4500), .A1 (n_5892), .B0 (n_5313), .Y (n_5348));
OAI21X1 g57077(.A0 (n_4437), .A1 (n_5841), .B0 (n_5311), .Y (n_5347));
OAI21X1 g57079(.A0 (n_4379), .A1 (n_5879), .B0 (n_5310), .Y (n_5345));
OAI21X1 g57080(.A0 (n_4343), .A1 (n_5320), .B0 (n_5309), .Y (n_5343));
OAI21X1 g57112(.A0 (n_5285), .A1 (n_4149), .B0 (n_5566), .Y (n_5342));
CLKBUFX1 gbuf_d_287(.A(n_5300), .Y(d_out_287));
CLKBUFX1 gbuf_qn_287(.A(qn_in_287), .Y(WX8287));
OAI21X1 g57206(.A0 (n_5279), .A1 (n_5709), .B0 (n_4068), .Y(DATA_9_6));
CLKBUFX1 gbuf_d_288(.A(n_5297), .Y(d_out_288));
CLKBUFX1 gbuf_qn_288(.A(qn_in_288), .Y(WX9580));
CLKBUFX1 gbuf_d_289(.A(n_5293), .Y(d_out_289));
CLKBUFX1 gbuf_qn_289(.A(qn_in_289), .Y(WX3115));
CLKBUFX1 gbuf_d_290(.A(n_5318), .Y(d_out_290));
CLKBUFX1 gbuf_q_290(.A(q_in_290), .Y(WX4574));
CLKBUFX1 gbuf_d_291(.A(n_5305), .Y(d_out_291));
CLKBUFX1 gbuf_q_291(.A(q_in_291), .Y(WX11037));
CLKBUFX1 gbuf_d_292(.A(n_5307), .Y(d_out_292));
CLKBUFX1 gbuf_q_292(.A(q_in_292), .Y(WX1986));
CLKBUFX1 gbuf_d_293(.A(n_6549), .Y(d_out_293));
CLKBUFX1 gbuf_q_293(.A(q_in_293), .Y(WX699));
OAI21X1 g56344(.A0 (n_4304), .A1 (n_8541), .B0 (n_4947), .Y (n_5338));
CLKBUFX1 gbuf_d_294(.A(n_5291), .Y(d_out_294));
CLKBUFX1 gbuf_qn_294(.A(qn_in_294), .Y(WX4410));
OAI21X1 g56371(.A0 (n_4654), .A1 (n_5317), .B0 (n_5289), .Y (n_5336));
OAI21X1 g56431(.A0 (n_4115), .A1 (n_5334), .B0 (n_5282), .Y (n_5335));
NOR2X1 g57101(.A (WX4372), .B (n_5181), .Y (n_5333));
NOR2X1 g57105(.A (WX4372), .B (n_5479), .Y (n_5331));
NOR2X1 g57108(.A (WX5663), .B (n_1648), .Y (n_5330));
NOR2X1 g57109(.A (WX5663), .B (n_5662), .Y (n_6666));
NOR2X1 g57116(.A (WX6954), .B (n_5712), .Y (n_5328));
NOR2X1 g57118(.A (WX6954), .B (n_5662), .Y (n_6192));
NOR2X1 g57120(.A (WX3081), .B (n_1648), .Y (n_5325));
NOR2X1 g57121(.A (WX3081), .B (n_5811), .Y (n_6193));
CLKBUFX1 gbuf_d_295(.A(n_5288), .Y(d_out_295));
CLKBUFX1 gbuf_qn_295(.A(qn_in_295), .Y(WX10873));
CLKBUFX1 gbuf_d_296(.A(n_5287), .Y(d_out_296));
CLKBUFX1 gbuf_qn_296(.A(qn_in_296), .Y(WX1822));
OAI21X1 g56485(.A0 (n_4287), .A1 (n_5105), .B0 (n_5281), .Y (n_5323));
OAI21X1 g57203(.A0 (n_5261), .A1 (n_5889), .B0 (n_5160), .Y (n_8335));
INVX1 g57247(.A (WX533), .Y (n_5356));
OAI21X1 g56545(.A0 (n_4510), .A1 (n_5320), .B0 (n_5278), .Y (n_5321));
OAI21X1 g56248(.A0 (n_4305), .A1 (n_5535), .B0 (n_5276), .Y (n_5319));
OAI21X1 g56370(.A0 (n_4239), .A1 (n_5317), .B0 (n_5274), .Y (n_5318));
CLKBUFX1 gbuf_d_297(.A(n_5272), .Y(d_out_297));
CLKBUFX1 gbuf_q_297(.A(q_in_297), .Y(WX9700));
NOR2X1 g56406(.A (WX5703), .B (n_2620), .Y (n_5316));
NOR2X1 g56407(.A (WX5703), .B (n_5500), .Y (n_6691));
OAI21X1 g57098(.A0 (n_5252), .A1 (n_4380), .B0 (n_4860), .Y (n_5314));
OAI21X1 g57106(.A0 (n_5250), .A1 (n_4346), .B0 (n_5566), .Y (n_5313));
OAI21X1 g57110(.A0 (n_4501), .A1 (n_6221), .B0 (n_4860), .Y (n_5311));
OAI21X1 g57119(.A0 (n_4438), .A1 (n_6194), .B0 (n_5460), .Y (n_5310));
OAI21X1 g57122(.A0 (n_4521), .A1 (n_6667), .B0 (n_5722), .Y (n_5309));
OAI21X1 g57137(.A0 (n_4223), .A1 (n_5928), .B0 (n_5264), .Y (n_5307));
OAI21X1 g57141(.A0 (n_3813), .A1 (n_5886), .B0 (n_5263), .Y (n_5305));
NOR2X1 g56470(.A (WX6996), .B (n_1648), .Y (n_5304));
NOR2X1 g56472(.A (WX6996), .B (n_5811), .Y (n_6692));
NOR2X1 g56506(.A (WX8289), .B (n_1425), .Y (n_5300));
CLKBUFX1 gbuf_d_298(.A(n_5259), .Y(d_out_298));
CLKBUFX1 gbuf_q_298(.A(q_in_298), .Y(WX533));
NOR2X1 g56511(.A (WX8289), .B (n_5838), .Y (n_9822));
NOR2X1 g56573(.A (WX9582), .B (n_1648), .Y (n_5297));
NOR2X1 g56575(.A (WX9582), .B (n_5822), .Y (n_9823));
NOR2X1 g56273(.A (WX3117), .B (n_5811), .Y (n_5294));
NOR2X1 g56294(.A (WX3117), .B (n_5181), .Y (n_5293));
CLKBUFX1 gbuf_d_299(.A(n_5273), .Y(d_out_299));
CLKBUFX1 gbuf_q_299(.A(q_in_299), .Y(WX8409));
CLKBUFX1 gbuf_d_300(.A(n_5271), .Y(d_out_300));
CLKBUFX1 gbuf_q_300(.A(q_in_300), .Y(WX4536));
CLKBUFX1 gbuf_d_301(.A(n_5269), .Y(d_out_301));
CLKBUFX1 gbuf_q_301(.A(q_in_301), .Y(WX5827));
CLKBUFX1 gbuf_d_302(.A(n_5267), .Y(d_out_302));
CLKBUFX1 gbuf_q_302(.A(q_in_302), .Y(WX7118));
CLKBUFX1 gbuf_d_303(.A(n_5265), .Y(d_out_303));
CLKBUFX1 gbuf_q_303(.A(q_in_303), .Y(WX3245));
NOR2X1 g56396(.A (WX4412), .B (n_3690), .Y (n_5291));
NOR2X1 g56401(.A (WX4412), .B (n_5427), .Y (n_8541));
OAI21X1 g56408(.A0 (n_4461), .A1 (n_6693), .B0 (n_4860), .Y (n_5289));
CLKBUFX1 gbuf_d_304(.A(n_5251), .Y(d_out_304));
CLKBUFX1 gbuf_qn_304(.A(qn_in_304), .Y(WX4372));
CLKBUFX1 gbuf_d_305(.A(n_5249), .Y(d_out_305));
CLKBUFX1 gbuf_qn_305(.A(qn_in_305), .Y(WX5663));
CLKBUFX1 gbuf_d_306(.A(n_5247), .Y(d_out_306));
CLKBUFX1 gbuf_qn_306(.A(qn_in_306), .Y(WX6954));
CLKBUFX1 gbuf_d_307(.A(n_5245), .Y(d_out_307));
CLKBUFX1 gbuf_qn_307(.A(qn_in_307), .Y(WX3081));
NOR2X1 g57159(.A (WX10875), .B (n_2620), .Y (n_5288));
NOR2X1 g57160(.A (WX1824), .B (n_2620), .Y (n_5287));
NOR2X1 g57171(.A (WX1824), .B (n_5838), .Y (n_5285));
OAI21X1 g56473(.A0 (n_4653), .A1 (n_9824), .B0 (n_5722), .Y (n_5282));
OAI21X1 g56512(.A0 (n_4114), .A1 (n_8542), .B0 (n_3183), .Y (n_5281));
MX2X1 g57265(.A (n_5257), .B (WX535), .S0 (n_6601), .Y (n_5279));
OAI21X1 g56576(.A0 (n_4286), .A1 (n_8553), .B0 (n_5460), .Y (n_5278));
OAI21X1 g56274(.A0 (n_5214), .A1 (n_4222), .B0 (n_5275), .Y (n_5276));
CLKBUFX1 gbuf_d_308(.A(n_5238), .Y(d_out_308));
CLKBUFX1 gbuf_q_308(.A(q_in_308), .Y(WX3281));
CLKBUFX1 gbuf_d_309(.A(n_5255), .Y(d_out_309));
CLKBUFX1 gbuf_q_309(.A(q_in_309), .Y(WX5867));
CLKBUFX1 gbuf_d_310(.A(n_5243), .Y(d_out_310));
CLKBUFX1 gbuf_q_310(.A(q_in_310), .Y(WX7160));
CLKBUFX1 gbuf_d_311(.A(n_5241), .Y(d_out_311));
CLKBUFX1 gbuf_q_311(.A(q_in_311), .Y(WX8453));
CLKBUFX1 gbuf_d_312(.A(n_5240), .Y(d_out_312));
CLKBUFX1 gbuf_q_312(.A(q_in_312), .Y(WX9746));
CLKBUFX1 gbuf_d_313(.A(n_5253), .Y(d_out_313));
CLKBUFX1 gbuf_qn_313(.A(qn_in_313), .Y(WX8245));
OAI21X1 g56402(.A0 (n_5212), .A1 (n_9413), .B0 (n_5566), .Y (n_5274));
CLKBUFX1 gbuf_d_314(.A(n_5233), .Y(d_out_314));
CLKBUFX1 gbuf_qn_314(.A(qn_in_314), .Y(WX5703));
OAI21X1 g57133(.A0 (n_4613), .A1 (n_5239), .B0 (n_5234), .Y (n_5273));
OAI21X1 g57134(.A0 (n_4552), .A1 (n_5158), .B0 (n_5232), .Y (n_5272));
OAI21X1 g57135(.A0 (n_4498), .A1 (n_5535), .B0 (n_5230), .Y (n_5271));
OAI21X1 g57136(.A0 (n_4435), .A1 (n_5493), .B0 (n_5228), .Y (n_5269));
OAI21X1 g57138(.A0 (n_4377), .A1 (n_5535), .B0 (n_5227), .Y (n_5267));
OAI21X1 g57139(.A0 (n_4339), .A1 (n_5196), .B0 (n_5226), .Y (n_5265));
OAI21X1 g57172(.A0 (n_5207), .A1 (n_4147), .B0 (n_4947), .Y (n_5264));
OAI21X1 g57174(.A0 (n_4509), .A1 (n_6682), .B0 (n_5460), .Y (n_5263));
CLKBUFX1 gbuf_d_315(.A(n_5222), .Y(d_out_315));
CLKBUFX1 gbuf_qn_315(.A(qn_in_315), .Y(WX6996));
INVX1 g57266(.A (DATA_9_5), .Y (n_5261));
NOR2X1 g57293(.A (n_5181), .B (n_5257), .Y (n_5259));
CLKBUFX1 gbuf_d_316(.A(n_5219), .Y(d_out_316));
CLKBUFX1 gbuf_qn_316(.A(qn_in_316), .Y(WX8289));
OR2X1 g57302(.A (n_5257), .B (n_5968), .Y (n_5256));
CLKBUFX1 gbuf_d_317(.A(n_5217), .Y(d_out_317));
CLKBUFX1 gbuf_qn_317(.A(qn_in_317), .Y(WX9582));
CLKBUFX1 gbuf_d_318(.A(n_5236), .Y(d_out_318));
CLKBUFX1 gbuf_q_318(.A(q_in_318), .Y(WX4576));
CLKBUFX1 gbuf_d_319(.A(n_5225), .Y(d_out_319));
CLKBUFX1 gbuf_q_319(.A(q_in_319), .Y(WX1988));
CLKBUFX1 gbuf_d_320(.A(n_5237), .Y(d_out_320));
CLKBUFX1 gbuf_qn_320(.A(qn_in_320), .Y(WX3117));
CLKBUFX1 gbuf_d_321(.A(n_5224), .Y(d_out_321));
CLKBUFX1 gbuf_q_321(.A(q_in_321), .Y(WX11039));
CLKBUFX1 gbuf_d_322(.A(n_5213), .Y(d_out_322));
CLKBUFX1 gbuf_qn_322(.A(qn_in_322), .Y(WX4412));
OAI21X1 g56430(.A0 (n_4215), .A1 (n_5254), .B0 (n_5211), .Y (n_5255));
NOR2X1 g57156(.A (WX8247), .B (n_5712), .Y (n_5253));
NOR2X1 g57157(.A (WX8247), .B (n_5811), .Y (n_5252));
NOR2X1 g57162(.A (WX4374), .B (n_1425), .Y (n_5251));
NOR2X1 g57165(.A (WX4374), .B (n_5662), .Y (n_5250));
NOR2X1 g57168(.A (WX5665), .B (n_5712), .Y (n_5249));
NOR2X1 g57169(.A (WX5665), .B (n_5838), .Y (n_6221));
NOR2X1 g57176(.A (WX6956), .B (n_5181), .Y (n_5247));
NOR2X1 g57178(.A (WX6956), .B (n_5427), .Y (n_6194));
NOR2X1 g57180(.A (WX3083), .B (n_5181), .Y (n_5245));
NOR2X1 g57181(.A (WX3083), .B (n_5500), .Y (n_6667));
CLKBUFX1 gbuf_d_323(.A(n_5210), .Y(d_out_323));
CLKBUFX1 gbuf_qn_323(.A(qn_in_323), .Y(WX10875));
CLKBUFX1 gbuf_d_324(.A(n_5208), .Y(d_out_324));
CLKBUFX1 gbuf_qn_324(.A(qn_in_324), .Y(WX1824));
OAI21X1 g56490(.A0 (n_4113), .A1 (n_5183), .B0 (n_5203), .Y (n_5243));
OAI21X1 g57267(.A0 (n_5187), .A1 (n_5242), .B0 (n_4066), .Y(DATA_9_5));
OAI21X1 g56544(.A0 (n_4285), .A1 (n_5320), .B0 (n_5201), .Y (n_5241));
OAI21X1 g56605(.A0 (n_4506), .A1 (n_5239), .B0 (n_5200), .Y (n_5240));
CLKBUFX1 gbuf_d_325(.A(n_5204), .Y(d_out_325));
CLKBUFX1 gbuf_q_325(.A(q_in_325), .Y(WX701));
OAI21X1 g56307(.A0 (n_4587), .A1 (n_5085), .B0 (n_5199), .Y (n_5238));
NOR2X1 g56353(.A (WX3119), .B (n_5712), .Y (n_5237));
OAI21X1 g56429(.A0 (n_4237), .A1 (n_5235), .B0 (n_5198), .Y (n_5236));
OAI21X1 g57158(.A0 (n_5180), .A1 (n_4378), .B0 (n_6479), .Y (n_5234));
NOR2X1 g56465(.A (WX5705), .B (n_5181), .Y (n_5233));
OAI21X1 g57164(.A0 (n_4614), .A1 (n_6222), .B0 (n_5722), .Y (n_5232));
NOR2X1 g56466(.A (WX5705), .B (n_5662), .Y (n_6693));
OAI21X1 g57166(.A0 (n_4342), .A1 (n_6223), .B0 (n_5566), .Y (n_5230));
OAI21X1 g57170(.A0 (n_4499), .A1 (n_6224), .B0 (n_4860), .Y (n_5228));
OAI21X1 g57179(.A0 (n_4436), .A1 (n_6674), .B0 (n_6479), .Y (n_5227));
OAI21X1 g57182(.A0 (n_4495), .A1 (n_6225), .B0 (n_4860), .Y (n_5226));
OAI21X1 g57197(.A0 (n_4398), .A1 (n_5493), .B0 (n_5190), .Y (n_5225));
OAI21X1 g57202(.A0 (n_3811), .A1 (n_5535), .B0 (n_5189), .Y (n_5224));
NOR2X1 g56529(.A (WX6998), .B (n_5712), .Y (n_5222));
NOR2X1 g56531(.A (WX6998), .B (n_5811), .Y (n_9824));
INVX1 g57311(.A (WX535), .Y (n_5257));
NOR2X1 g56566(.A (WX8291), .B (n_2620), .Y (n_5219));
NOR2X1 g56571(.A (WX8291), .B (n_4882), .Y (n_8542));
NOR2X1 g56633(.A (WX9584), .B (n_2849), .Y (n_5217));
NOR2X1 g56635(.A (WX9584), .B (n_5427), .Y (n_8553));
CLKBUFX1 gbuf_d_326(.A(n_6505), .Y(d_out_326));
CLKBUFX1 gbuf_q_326(.A(q_in_326), .Y(WX9702));
CLKBUFX1 gbuf_d_327(.A(n_5194), .Y(d_out_327));
CLKBUFX1 gbuf_q_327(.A(q_in_327), .Y(WX4538));
CLKBUFX1 gbuf_d_328(.A(n_5191), .Y(d_out_328));
CLKBUFX1 gbuf_q_328(.A(q_in_328), .Y(WX3247));
CLKBUFX1 gbuf_d_329(.A(n_5193), .Y(d_out_329));
CLKBUFX1 gbuf_q_329(.A(q_in_329), .Y(WX5829));
CLKBUFX1 gbuf_d_330(.A(n_5197), .Y(d_out_330));
CLKBUFX1 gbuf_q_330(.A(q_in_330), .Y(WX8411));
CLKBUFX1 gbuf_d_331(.A(n_5192), .Y(d_out_331));
CLKBUFX1 gbuf_q_331(.A(q_in_331), .Y(WX7120));
NOR2X1 g56332(.A (WX3119), .B (n_5427), .Y (n_5214));
NOR2X1 g56455(.A (WX4414), .B (n_2605), .Y (n_5213));
NOR2X1 g56460(.A (WX4414), .B (n_5662), .Y (n_5212));
OAI21X1 g56467(.A0 (n_4238), .A1 (n_8543), .B0 (n_5722), .Y (n_5211));
CLKBUFX1 gbuf_d_332(.A(n_5182), .Y(d_out_332));
CLKBUFX1 gbuf_qn_332(.A(qn_in_332), .Y(WX8247));
CLKBUFX1 gbuf_d_333(.A(n_5177), .Y(d_out_333));
CLKBUFX1 gbuf_qn_333(.A(qn_in_333), .Y(WX4374));
CLKBUFX1 gbuf_d_334(.A(n_5173), .Y(d_out_334));
CLKBUFX1 gbuf_qn_334(.A(qn_in_334), .Y(WX5665));
CLKBUFX1 gbuf_d_335(.A(n_5171), .Y(d_out_335));
CLKBUFX1 gbuf_qn_335(.A(qn_in_335), .Y(WX6956));
CLKBUFX1 gbuf_d_336(.A(n_5169), .Y(d_out_336));
CLKBUFX1 gbuf_qn_336(.A(qn_in_336), .Y(WX3083));
NOR2X1 g57219(.A (WX10877), .B (n_2620), .Y (n_5210));
NOR2X1 g57220(.A (WX1826), .B (n_2620), .Y (n_5208));
NOR2X1 g57231(.A (WX1826), .B (n_5838), .Y (n_5207));
NOR2X1 g57234(.A (WX10877), .B (n_5662), .Y (n_6682));
NAND2X1 g57262(.A (n_5166), .B (n_4693), .Y (n_5204));
OAI21X1 g56532(.A0 (n_15859), .A1 (n_15860), .B0 (n_5619), .Y(n_5203));
CLKBUFX1 gbuf_d_337(.A(n_5162), .Y(d_out_337));
CLKBUFX1 gbuf_q_337(.A(q_in_337), .Y(WX535));
OAI21X1 g56572(.A0 (n_4112), .A1 (n_8554), .B0 (n_5556), .Y (n_5201));
OAI21X1 g56636(.A0 (n_5135), .A1 (n_11595), .B0 (n_5619), .Y(n_5200));
CLKBUFX1 gbuf_d_338(.A(n_5186), .Y(d_out_338));
CLKBUFX1 gbuf_q_338(.A(q_in_338), .Y(WX3283));
CLKBUFX1 gbuf_d_339(.A(n_5184), .Y(d_out_339));
CLKBUFX1 gbuf_q_339(.A(q_in_339), .Y(WX5869));
CLKBUFX1 gbuf_d_340(.A(n_5165), .Y(d_out_340));
CLKBUFX1 gbuf_q_340(.A(q_in_340), .Y(WX7162));
CLKBUFX1 gbuf_d_341(.A(n_5159), .Y(d_out_341));
CLKBUFX1 gbuf_q_341(.A(q_in_341), .Y(WX8455));
CLKBUFX1 gbuf_d_342(.A(n_5157), .Y(d_out_342));
CLKBUFX1 gbuf_q_342(.A(q_in_342), .Y(WX9748));
CLKBUFX1 gbuf_d_343(.A(n_5179), .Y(d_out_343));
CLKBUFX1 gbuf_qn_343(.A(qn_in_343), .Y(WX9538));
OAI21X1 g56333(.A0 (n_5156), .A1 (n_9415), .B0 (n_5460), .Y (n_5199));
CLKBUFX1 gbuf_d_344(.A(n_5154), .Y(d_out_344));
CLKBUFX1 gbuf_qn_344(.A(qn_in_344), .Y(WX3119));
OAI21X1 g56461(.A0 (n_15861), .A1 (n_15862), .B0 (n_5722), .Y(n_5198));
CLKBUFX1 gbuf_d_345(.A(n_5143), .Y(d_out_345));
CLKBUFX1 gbuf_qn_345(.A(qn_in_345), .Y(WX5705));
OAI21X1 g57193(.A0 (n_4313), .A1 (n_5196), .B0 (n_5152), .Y (n_5197));
OAI21X1 g57195(.A0 (n_4494), .A1 (n_5334), .B0 (n_5150), .Y (n_5194));
OAI21X1 g57196(.A0 (n_4433), .A1 (n_5928), .B0 (n_5149), .Y (n_5193));
OAI21X1 g57198(.A0 (n_4375), .A1 (n_5254), .B0 (n_5148), .Y (n_5192));
OAI21X1 g57199(.A0 (n_4337), .A1 (n_5235), .B0 (n_5146), .Y (n_5191));
OAI21X1 g57232(.A0 (n_5126), .A1 (n_4145), .B0 (n_5722), .Y (n_5190));
OAI21X1 g57235(.A0 (n_4505), .A1 (n_6680), .B0 (n_4860), .Y (n_5189));
CLKBUFX1 gbuf_d_346(.A(n_5141), .Y(d_out_346));
CLKBUFX1 gbuf_qn_346(.A(qn_in_346), .Y(WX6998));
MX2X1 g57334(.A (n_5161), .B (WX537), .S0 (n_10743), .Y (n_5187));
CLKBUFX1 gbuf_d_347(.A(n_5139), .Y(d_out_347));
CLKBUFX1 gbuf_qn_347(.A(qn_in_347), .Y(WX8291));
CLKBUFX1 gbuf_d_348(.A(n_5136), .Y(d_out_348));
CLKBUFX1 gbuf_qn_348(.A(qn_in_348), .Y(WX9584));
CLKBUFX1 gbuf_d_349(.A(n_5153), .Y(d_out_349));
CLKBUFX1 gbuf_q_349(.A(q_in_349), .Y(WX4578));
CLKBUFX1 gbuf_d_350(.A(n_5144), .Y(d_out_350));
CLKBUFX1 gbuf_q_350(.A(q_in_350), .Y(WX11041));
CLKBUFX1 gbuf_d_351(.A(n_5145), .Y(d_out_351));
CLKBUFX1 gbuf_q_351(.A(q_in_351), .Y(WX1990));
OAI21X1 g56366(.A0 (n_4301), .A1 (n_5185), .B0 (n_5133), .Y (n_5186));
CLKBUFX1 gbuf_d_352(.A(n_5132), .Y(d_out_352));
CLKBUFX1 gbuf_qn_352(.A(qn_in_352), .Y(WX4414));
OAI21X1 g56489(.A0 (n_4662), .A1 (n_5183), .B0 (n_5129), .Y (n_5184));
NOR2X1 g57216(.A (WX8249), .B (n_5181), .Y (n_5182));
NOR2X1 g57217(.A (WX8249), .B (n_5500), .Y (n_5180));
NOR2X1 g57221(.A (WX9540), .B (n_2851), .Y (n_5179));
NOR2X1 g57222(.A (WX4376), .B (n_2851), .Y (n_5177));
NOR2X1 g57223(.A (WX9540), .B (n_5500), .Y (n_6222));
NOR2X1 g57225(.A (WX4376), .B (n_5811), .Y (n_6223));
NOR2X1 g57228(.A (WX5667), .B (n_1648), .Y (n_5173));
NOR2X1 g57229(.A (WX5667), .B (n_5811), .Y (n_6224));
NOR2X1 g57237(.A (WX6958), .B (n_5712), .Y (n_5171));
NOR2X1 g57239(.A (WX6958), .B (n_5662), .Y (n_6674));
NOR2X1 g57241(.A (WX3085), .B (n_1648), .Y (n_5169));
NOR2X1 g57242(.A (WX3085), .B (n_5811), .Y (n_6225));
CLKBUFX1 gbuf_d_353(.A(n_5127), .Y(d_out_353));
CLKBUFX1 gbuf_qn_353(.A(qn_in_353), .Y(WX1826));
CLKBUFX1 gbuf_d_354(.A(n_5128), .Y(d_out_354));
CLKBUFX1 gbuf_qn_354(.A(qn_in_354), .Y(WX10877));
NAND2X1 g57303(.A (n_5123), .B (n_6615), .Y (n_5166));
OAI21X1 g56549(.A0 (n_4111), .A1 (n_5928), .B0 (n_5122), .Y (n_5165));
INVX1 g57335(.A (DATA_9_4), .Y (n_5164));
NOR2X1 g57360(.A (n_1425), .B (n_5161), .Y (n_5162));
OR2X1 g57369(.A (n_5161), .B (n_5990), .Y (n_5160));
OAI21X1 g56604(.A0 (n_4281), .A1 (n_5158), .B0 (n_5121), .Y (n_5159));
OAI21X1 g56664(.A0 (n_4265), .A1 (n_5490), .B0 (n_5119), .Y (n_5157));
NOR2X1 g56391(.A (WX3121), .B (n_5427), .Y (n_5156));
NOR2X1 g56412(.A (WX3121), .B (n_3188), .Y (n_5154));
OAI21X1 g56488(.A0 (n_4235), .A1 (n_5825), .B0 (n_5111), .Y (n_5153));
OAI21X1 g57218(.A0 (n_4376), .A1 (n_6227), .B0 (n_4860), .Y (n_5152));
OAI21X1 g57226(.A0 (n_4338), .A1 (n_6195), .B0 (n_5619), .Y (n_5150));
OAI21X1 g57230(.A0 (n_4497), .A1 (n_6226), .B0 (n_5566), .Y (n_5149));
OAI21X1 g57240(.A0 (n_4434), .A1 (n_6228), .B0 (n_4947), .Y (n_5148));
OAI21X1 g57243(.A0 (n_4487), .A1 (n_6675), .B0 (n_3183), .Y (n_5146));
OAI21X1 g57259(.A0 (n_4213), .A1 (n_5254), .B0 (n_5110), .Y (n_5145));
OAI21X1 g57263(.A0 (n_3810), .A1 (n_5320), .B0 (n_5109), .Y (n_5144));
NOR2X1 g56524(.A (WX5707), .B (n_2620), .Y (n_5143));
NOR2X1 g56525(.A (WX5707), .B (n_5838), .Y (n_8543));
OAI21X1 g57336(.A0 (n_5089), .A1 (n_6091), .B0 (n_4062), .Y(DATA_9_4));
NOR2X1 g56589(.A (WX7000), .B (n_5712), .Y (n_5141));
NOR2X1 g56591(.A (WX7000), .B (n_5500), .Y (n_15860));
CLKBUFX1 gbuf_d_355(.A(n_5113), .Y(d_out_355));
CLKBUFX1 gbuf_q_355(.A(q_in_355), .Y(WX5831));
NOR2X1 g56626(.A (WX8293), .B (n_5181), .Y (n_5139));
NOR2X1 g56631(.A (WX8293), .B (n_5479), .Y (n_8554));
NOR2X1 g56692(.A (WX9586), .B (n_1425), .Y (n_5136));
NOR2X1 g56694(.A (WX9586), .B (n_5662), .Y (n_5135));
CLKBUFX1 gbuf_d_356(.A(n_5118), .Y(d_out_356));
CLKBUFX1 gbuf_q_356(.A(q_in_356), .Y(WX3249));
CLKBUFX1 gbuf_d_357(.A(n_5117), .Y(d_out_357));
CLKBUFX1 gbuf_q_357(.A(q_in_357), .Y(WX8413));
CLKBUFX1 gbuf_d_358(.A(n_5116), .Y(d_out_358));
CLKBUFX1 gbuf_q_358(.A(q_in_358), .Y(WX9704));
CLKBUFX1 gbuf_d_359(.A(n_5115), .Y(d_out_359));
CLKBUFX1 gbuf_q_359(.A(q_in_359), .Y(WX4540));
CLKBUFX1 gbuf_d_360(.A(n_5112), .Y(d_out_360));
CLKBUFX1 gbuf_q_360(.A(q_in_360), .Y(WX7122));
CLKBUFX1 gbuf_d_361(.A(n_5107), .Y(d_out_361));
CLKBUFX1 gbuf_q_361(.A(q_in_361), .Y(WX703));
OAI21X1 g56392(.A0 (n_5084), .A1 (n_11626), .B0 (n_5722), .Y(n_5133));
CLKBUFX1 gbuf_d_362(.A(n_5104), .Y(d_out_362));
CLKBUFX1 gbuf_qn_362(.A(qn_in_362), .Y(WX8249));
CLKBUFX1 gbuf_d_363(.A(n_5102), .Y(d_out_363));
CLKBUFX1 gbuf_qn_363(.A(qn_in_363), .Y(WX9540));
CLKBUFX1 gbuf_d_364(.A(n_5100), .Y(d_out_364));
CLKBUFX1 gbuf_qn_364(.A(qn_in_364), .Y(WX4376));
CLKBUFX1 gbuf_d_365(.A(n_5097), .Y(d_out_365));
CLKBUFX1 gbuf_qn_365(.A(qn_in_365), .Y(WX5667));
CLKBUFX1 gbuf_d_366(.A(n_5095), .Y(d_out_366));
CLKBUFX1 gbuf_qn_366(.A(qn_in_366), .Y(WX6958));
CLKBUFX1 gbuf_d_367(.A(n_5092), .Y(d_out_367));
CLKBUFX1 gbuf_qn_367(.A(qn_in_367), .Y(WX3085));
NOR2X1 g56514(.A (WX4416), .B (n_1425), .Y (n_5132));
NOR2X1 g56519(.A (WX4416), .B (n_5500), .Y (n_15862));
OAI21X1 g56526(.A0 (n_4236), .A1 (n_12492), .B0 (n_7087), .Y(n_5129));
NOR2X1 g57285(.A (WX10879), .B (n_1648), .Y (n_5128));
NOR2X1 g57286(.A (WX1828), .B (n_3188), .Y (n_5127));
NOR2X1 g57297(.A (WX1828), .B (n_4882), .Y (n_5126));
NOR2X1 g57299(.A (WX10879), .B (n_5427), .Y (n_6680));
OAI21X1 g57333(.A0 (n_5069), .A1 (n_5889), .B0 (n_4961), .Y (n_5123));
OAI21X1 g56565(.A0 (n_5064), .A1 (n_4661), .B0 (n_5556), .Y (n_5122));
INVX1 g57382(.A (WX537), .Y (n_5161));
OAI21X1 g56632(.A0 (n_5060), .A1 (n_10713), .B0 (n_5556), .Y(n_5121));
OAI21X1 g56695(.A0 (n_4280), .A1 (n_12493), .B0 (n_5619), .Y(n_5119));
CLKBUFX1 gbuf_d_368(.A(n_5106), .Y(d_out_368));
CLKBUFX1 gbuf_q_368(.A(q_in_368), .Y(WX3285));
CLKBUFX1 gbuf_d_369(.A(n_5090), .Y(d_out_369));
CLKBUFX1 gbuf_q_369(.A(q_in_369), .Y(WX5871));
CLKBUFX1 gbuf_d_370(.A(n_5088), .Y(d_out_370));
CLKBUFX1 gbuf_q_370(.A(q_in_370), .Y(WX7164));
CLKBUFX1 gbuf_d_371(.A(n_5087), .Y(d_out_371));
CLKBUFX1 gbuf_q_371(.A(q_in_371), .Y(WX8457));
CLKBUFX1 gbuf_d_372(.A(n_5086), .Y(d_out_372));
CLKBUFX1 gbuf_q_372(.A(q_in_372), .Y(WX9750));
CLKBUFX1 gbuf_d_373(.A(n_5083), .Y(d_out_373));
CLKBUFX1 gbuf_qn_373(.A(qn_in_373), .Y(WX3121));
OAI21X1 g57254(.A0 (n_4647), .A1 (n_5158), .B0 (n_5082), .Y (n_5118));
OAI21X1 g57255(.A0 (n_4611), .A1 (n_5235), .B0 (n_5081), .Y (n_5117));
OAI21X1 g57256(.A0 (n_4548), .A1 (n_5239), .B0 (n_5080), .Y (n_5116));
OAI21X1 g57257(.A0 (n_4492), .A1 (n_5439), .B0 (n_5079), .Y (n_5115));
OAI21X1 g57258(.A0 (n_4431), .A1 (n_5879), .B0 (n_5078), .Y (n_5113));
OAI21X1 g57260(.A0 (n_4132), .A1 (n_5879), .B0 (n_5076), .Y (n_5112));
OAI21X1 g56520(.A0 (n_4578), .A1 (n_6694), .B0 (n_7087), .Y (n_5111));
OAI21X1 g57298(.A0 (n_5053), .A1 (n_4143), .B0 (n_5460), .Y (n_5110));
OAI21X1 g57300(.A0 (n_4264), .A1 (n_7507), .B0 (n_5460), .Y (n_5109));
CLKBUFX1 gbuf_d_374(.A(n_5071), .Y(d_out_374));
CLKBUFX1 gbuf_qn_374(.A(qn_in_374), .Y(WX5707));
NAND2X2 g57326(.A (n_5072), .B (n_4692), .Y (n_5107));
CLKBUFX1 gbuf_d_375(.A(n_5067), .Y(d_out_375));
CLKBUFX1 gbuf_q_375(.A(q_in_375), .Y(WX537));
CLKBUFX1 gbuf_d_376(.A(n_5063), .Y(d_out_376));
CLKBUFX1 gbuf_qn_376(.A(qn_in_376), .Y(WX7000));
CLKBUFX1 gbuf_d_377(.A(n_5062), .Y(d_out_377));
CLKBUFX1 gbuf_qn_377(.A(qn_in_377), .Y(WX8293));
CLKBUFX1 gbuf_d_378(.A(n_5059), .Y(d_out_378));
CLKBUFX1 gbuf_qn_378(.A(qn_in_378), .Y(WX9586));
CLKBUFX1 gbuf_d_379(.A(n_5075), .Y(d_out_379));
CLKBUFX1 gbuf_q_379(.A(q_in_379), .Y(WX4580));
CLKBUFX1 gbuf_d_380(.A(n_5073), .Y(d_out_380));
CLKBUFX1 gbuf_q_380(.A(q_in_380), .Y(WX11043));
CLKBUFX1 gbuf_d_381(.A(n_5074), .Y(d_out_381));
CLKBUFX1 gbuf_q_381(.A(q_in_381), .Y(WX1992));
OAI21X1 g56425(.A0 (n_4580), .A1 (n_5105), .B0 (n_5056), .Y (n_5106));
NOR2X1 g57282(.A (WX8251), .B (n_5712), .Y (n_5104));
NOR2X1 g57283(.A (WX8251), .B (n_5811), .Y (n_6227));
NOR2X1 g57287(.A (WX9542), .B (n_1425), .Y (n_5102));
NOR2X1 g57288(.A (WX4378), .B (n_5181), .Y (n_5100));
NOR2X1 g57291(.A (WX4378), .B (n_4882), .Y (n_6195));
NOR2X1 g57294(.A (WX5669), .B (n_5712), .Y (n_5097));
NOR2X1 g57295(.A (WX5669), .B (n_4882), .Y (n_6226));
NOR2X1 g57301(.A (WX6960), .B (n_5712), .Y (n_5095));
CLKBUFX1 gbuf_d_382(.A(n_5050), .Y(d_out_382));
CLKBUFX1 gbuf_qn_382(.A(qn_in_382), .Y(WX4416));
NOR2X1 g57304(.A (WX6960), .B (n_5822), .Y (n_6228));
NOR2X1 g57305(.A (WX3087), .B (n_1648), .Y (n_5092));
NOR2X1 g57307(.A (WX3087), .B (n_5427), .Y (n_6675));
CLKBUFX1 gbuf_d_383(.A(n_5055), .Y(d_out_383));
CLKBUFX1 gbuf_qn_383(.A(qn_in_383), .Y(WX10879));
CLKBUFX1 gbuf_d_384(.A(n_5054), .Y(d_out_384));
CLKBUFX1 gbuf_qn_384(.A(qn_in_384), .Y(WX1828));
OAI21X1 g56548(.A0 (n_4211), .A1 (n_5649), .B0 (n_5047), .Y (n_5090));
MX2X1 g57400(.A (n_5066), .B (WX539), .S0 (n_4061), .Y (n_5089));
OAI21X1 g56602(.A0 (n_4326), .A1 (n_5841), .B0 (n_5046), .Y (n_5088));
OAI21X1 g56663(.A0 (n_4565), .A1 (n_5576), .B0 (n_5045), .Y (n_5087));
OAI21X1 g56722(.A0 (n_4263), .A1 (n_5085), .B0 (n_5043), .Y (n_5086));
NOR2X1 g56450(.A (WX3123), .B (n_5427), .Y (n_5084));
NOR2X1 g56471(.A (WX3123), .B (n_5712), .Y (n_5083));
OAI21X1 g57281(.A0 (n_5028), .A1 (n_4252), .B0 (n_5566), .Y (n_5082));
OAI21X1 g57284(.A0 (n_4374), .A1 (n_6197), .B0 (n_5460), .Y (n_5081));
OAI21X1 g57290(.A0 (n_5022), .A1 (n_4312), .B0 (n_4947), .Y (n_5080));
OAI21X1 g57292(.A0 (n_4336), .A1 (n_6229), .B0 (n_3183), .Y (n_5079));
OAI21X1 g57296(.A0 (n_4493), .A1 (n_6196), .B0 (n_4860), .Y (n_5078));
OAI21X1 g57306(.A0 (n_4432), .A1 (n_6672), .B0 (n_4947), .Y (n_5076));
OAI21X1 g56546(.A0 (n_4233), .A1 (n_5235), .B0 (n_5034), .Y (n_5075));
OAI21X1 g57324(.A0 (n_4394), .A1 (n_5892), .B0 (n_5036), .Y (n_5074));
OAI21X1 g57330(.A0 (n_3818), .A1 (n_5439), .B0 (n_5035), .Y (n_5073));
NAND2X1 g57371(.A (n_6615), .B (n_8320), .Y (n_5072));
NOR2X1 g56584(.A (WX5709), .B (n_5181), .Y (n_5071));
NOR2X1 g56585(.A (WX5709), .B (n_5052), .Y (n_12492));
INVX1 g57402(.A (DATA_9_3), .Y (n_5069));
NOR2X1 g57450(.A (n_5181), .B (n_5066), .Y (n_5067));
OR2X1 g57457(.A (n_5066), .B (n_3828), .Y (n_5065));
NOR2X1 g56624(.A (WX7002), .B (n_5500), .Y (n_5064));
NOR2X1 g56649(.A (WX7002), .B (n_1425), .Y (n_5063));
NOR2X1 g56685(.A (WX8295), .B (n_5181), .Y (n_5062));
NOR2X1 g56690(.A (WX8295), .B (n_5662), .Y (n_5060));
NOR2X1 g56750(.A (WX9588), .B (n_5712), .Y (n_5059));
NOR2X1 g56752(.A (WX9588), .B (n_5427), .Y (n_12493));
CLKBUFX1 gbuf_d_385(.A(n_5038), .Y(d_out_385));
CLKBUFX1 gbuf_q_385(.A(q_in_385), .Y(WX5833));
CLKBUFX1 gbuf_d_386(.A(n_5042), .Y(d_out_386));
CLKBUFX1 gbuf_q_386(.A(q_in_386), .Y(WX3251));
CLKBUFX1 gbuf_d_387(.A(n_5041), .Y(d_out_387));
CLKBUFX1 gbuf_q_387(.A(q_in_387), .Y(WX8415));
CLKBUFX1 gbuf_d_388(.A(n_5040), .Y(d_out_388));
CLKBUFX1 gbuf_q_388(.A(q_in_388), .Y(WX9706));
CLKBUFX1 gbuf_d_389(.A(n_5039), .Y(d_out_389));
CLKBUFX1 gbuf_q_389(.A(q_in_389), .Y(WX4542));
CLKBUFX1 gbuf_d_390(.A(n_5037), .Y(d_out_390));
CLKBUFX1 gbuf_q_390(.A(q_in_390), .Y(WX7124));
OAI21X1 g56451(.A0 (n_15863), .A1 (n_15864), .B0 (n_5566), .Y(n_5056));
CLKBUFX1 gbuf_d_391(.A(n_5027), .Y(d_out_391));
CLKBUFX1 gbuf_qn_391(.A(qn_in_391), .Y(WX8251));
CLKBUFX1 gbuf_d_392(.A(n_5025), .Y(d_out_392));
CLKBUFX1 gbuf_qn_392(.A(qn_in_392), .Y(WX9542));
CLKBUFX1 gbuf_d_393(.A(n_5024), .Y(d_out_393));
CLKBUFX1 gbuf_qn_393(.A(qn_in_393), .Y(WX4378));
CLKBUFX1 gbuf_d_394(.A(n_5020), .Y(d_out_394));
CLKBUFX1 gbuf_qn_394(.A(qn_in_394), .Y(WX5669));
CLKBUFX1 gbuf_d_395(.A(n_5017), .Y(d_out_395));
CLKBUFX1 gbuf_qn_395(.A(qn_in_395), .Y(WX6960));
CLKBUFX1 gbuf_d_396(.A(n_5016), .Y(d_out_396));
CLKBUFX1 gbuf_qn_396(.A(qn_in_396), .Y(WX3087));
NOR2X1 g57350(.A (WX10881), .B (n_5181), .Y (n_5055));
NOR2X1 g57351(.A (WX1830), .B (n_2620), .Y (n_5054));
NOR2X1 g57364(.A (WX1830), .B (n_5052), .Y (n_5053));
NOR2X1 g57367(.A (WX10881), .B (n_5811), .Y (n_7507));
NOR2X1 g56574(.A (WX4418), .B (n_3188), .Y (n_5050));
NOR2X1 g56578(.A (WX4418), .B (n_5822), .Y (n_6694));
OAI21X1 g56586(.A0 (n_4992), .A1 (n_10717), .B0 (n_6497), .Y(n_5047));
OAI21X1 g57403(.A0 (n_4991), .A1 (n_5965), .B0 (n_4060), .Y(DATA_9_3));
OAI21X1 g56625(.A0 (n_4210), .A1 (n_8544), .B0 (n_4947), .Y (n_5046));
OAI21X1 g56691(.A0 (n_4985), .A1 (n_4325), .B0 (n_5566), .Y (n_5045));
OAI21X1 g56753(.A0 (n_4564), .A1 (n_6695), .B0 (n_5706), .Y (n_5043));
CLKBUFX1 gbuf_d_397(.A(n_5030), .Y(d_out_397));
CLKBUFX1 gbuf_q_397(.A(q_in_397), .Y(WX3287));
CLKBUFX1 gbuf_d_398(.A(n_5012), .Y(d_out_398));
CLKBUFX1 gbuf_q_398(.A(q_in_398), .Y(WX5873));
CLKBUFX1 gbuf_d_399(.A(n_5011), .Y(d_out_399));
CLKBUFX1 gbuf_q_399(.A(q_in_399), .Y(WX7166));
CLKBUFX1 gbuf_d_400(.A(n_5010), .Y(d_out_400));
CLKBUFX1 gbuf_q_400(.A(q_in_400), .Y(WX8459));
CLKBUFX1 gbuf_d_401(.A(n_5009), .Y(d_out_401));
CLKBUFX1 gbuf_q_401(.A(q_in_401), .Y(WX9752));
CLKBUFX1 gbuf_d_402(.A(n_6621), .Y(d_out_402));
CLKBUFX1 gbuf_q_402(.A(q_in_402), .Y(WX705));
CLKBUFX1 gbuf_d_403(.A(n_5007), .Y(d_out_403));
CLKBUFX1 gbuf_qn_403(.A(qn_in_403), .Y(WX3123));
OAI21X1 g57318(.A0 (n_4642), .A1 (n_5879), .B0 (n_5005), .Y (n_5042));
OAI21X1 g57319(.A0 (n_4609), .A1 (n_5474), .B0 (n_5004), .Y (n_5041));
OAI21X1 g57321(.A0 (n_4546), .A1 (n_5841), .B0 (n_5003), .Y (n_5040));
OAI21X1 g57322(.A0 (n_4490), .A1 (n_5105), .B0 (n_5001), .Y (n_5039));
OAI21X1 g57323(.A0 (n_4429), .A1 (n_5493), .B0 (n_4999), .Y (n_5038));
OAI21X1 g57325(.A0 (n_4130), .A1 (n_5183), .B0 (n_4998), .Y (n_5037));
OAI21X1 g57365(.A0 (n_4973), .A1 (n_4141), .B0 (n_5460), .Y (n_5036));
OAI21X1 g57370(.A0 (n_4262), .A1 (n_7508), .B0 (n_4860), .Y (n_5035));
OAI21X1 g56579(.A0 (n_15865), .A1 (n_15866), .B0 (n_5556), .Y(n_5034));
OAI21X1 g57397(.A0 (n_4966), .A1 (n_5889), .B0 (n_4873), .Y (n_8320));
CLKBUFX1 gbuf_d_404(.A(n_4994), .Y(d_out_404));
CLKBUFX1 gbuf_qn_404(.A(qn_in_404), .Y(WX5709));
INVX1 g57468(.A (WX539), .Y (n_5066));
CLKBUFX1 gbuf_d_405(.A(n_4988), .Y(d_out_405));
CLKBUFX1 gbuf_qn_405(.A(qn_in_405), .Y(WX7002));
CLKBUFX1 gbuf_d_406(.A(n_4986), .Y(d_out_406));
CLKBUFX1 gbuf_qn_406(.A(qn_in_406), .Y(WX8295));
CLKBUFX1 gbuf_d_407(.A(n_4984), .Y(d_out_407));
CLKBUFX1 gbuf_qn_407(.A(qn_in_407), .Y(WX9588));
CLKBUFX1 gbuf_d_408(.A(n_4995), .Y(d_out_408));
CLKBUFX1 gbuf_q_408(.A(q_in_408), .Y(WX4582));
CLKBUFX1 gbuf_d_409(.A(n_4996), .Y(d_out_409));
CLKBUFX1 gbuf_q_409(.A(q_in_409), .Y(WX11045));
CLKBUFX1 gbuf_d_410(.A(n_4997), .Y(d_out_410));
CLKBUFX1 gbuf_q_410(.A(q_in_410), .Y(WX1994));
OAI21X1 g56484(.A0 (n_4297), .A1 (n_5928), .B0 (n_4979), .Y (n_5030));
NOR2X1 g57345(.A (WX3089), .B (n_5822), .Y (n_5028));
NOR2X1 g57347(.A (WX8253), .B (n_5712), .Y (n_5027));
NOR2X1 g57348(.A (WX8253), .B (n_5811), .Y (n_6197));
NOR2X1 g57354(.A (WX9544), .B (n_1425), .Y (n_5025));
NOR2X1 g57355(.A (WX4380), .B (n_3188), .Y (n_5024));
NOR2X1 g57356(.A (WX9544), .B (n_5500), .Y (n_5022));
NOR2X1 g57358(.A (WX4380), .B (n_5052), .Y (n_6229));
NOR2X1 g57361(.A (WX5671), .B (n_2620), .Y (n_5020));
NOR2X1 g57362(.A (WX5671), .B (n_5052), .Y (n_6196));
NOR2X1 g57368(.A (WX6962), .B (n_5712), .Y (n_5017));
NOR2X1 g57374(.A (WX3089), .B (n_2849), .Y (n_5016));
NOR2X1 g57375(.A (WX6962), .B (n_5500), .Y (n_6672));
CLKBUFX1 gbuf_d_411(.A(n_4976), .Y(d_out_411));
CLKBUFX1 gbuf_qn_411(.A(qn_in_411), .Y(WX10881));
CLKBUFX1 gbuf_d_412(.A(n_4974), .Y(d_out_412));
CLKBUFX1 gbuf_qn_412(.A(qn_in_412), .Y(WX1830));
CLKBUFX1 gbuf_d_413(.A(n_4970), .Y(d_out_413));
CLKBUFX1 gbuf_qn_413(.A(qn_in_413), .Y(WX4418));
OAI21X1 g56608(.A0 (n_4392), .A1 (n_5886), .B0 (n_4968), .Y (n_5012));
CLKBUFX1 gbuf_d_414(.A(n_4964), .Y(d_out_414));
CLKBUFX1 gbuf_q_414(.A(q_in_414), .Y(WX539));
OAI21X1 g56661(.A0 (n_4324), .A1 (n_5830), .B0 (n_4962), .Y (n_5011));
OAI21X1 g56721(.A0 (n_4563), .A1 (n_5085), .B0 (n_4959), .Y (n_5010));
OAI21X1 g56782(.A0 (n_4504), .A1 (n_4803), .B0 (n_4958), .Y (n_5009));
CLKBUFX1 gbuf_d_415(.A(n_4960), .Y(d_out_415));
CLKBUFX1 gbuf_q_415(.A(q_in_415), .Y(WX649));
CLKBUFX1 gbuf_d_416(.A(n_4956), .Y(d_out_416));
CLKBUFX1 gbuf_q_416(.A(q_in_416), .Y(WX647));
CLKBUFX1 gbuf_d_417(.A(n_4980), .Y(d_out_417));
CLKBUFX1 gbuf_q_417(.A(q_in_417), .Y(WX645));
CLKBUFX1 gbuf_d_418(.A(n_4978), .Y(d_out_418));
CLKBUFX1 gbuf_q_418(.A(q_in_418), .Y(WX707));
NOR2X1 g56509(.A (WX3125), .B (n_5662), .Y (n_15864));
NOR2X1 g56530(.A (WX3125), .B (n_5712), .Y (n_5007));
OAI21X1 g57346(.A0 (n_4939), .A1 (n_4250), .B0 (n_4947), .Y (n_5005));
OAI21X1 g57349(.A0 (n_4936), .A1 (n_4131), .B0 (n_5460), .Y (n_5004));
OAI21X1 g57357(.A0 (n_4610), .A1 (n_6231), .B0 (n_4860), .Y (n_5003));
OAI21X1 g57359(.A0 (n_4646), .A1 (n_6198), .B0 (n_4947), .Y (n_5001));
OAI21X1 g57363(.A0 (n_4491), .A1 (n_6230), .B0 (n_4860), .Y (n_4999));
OAI21X1 g57376(.A0 (n_4924), .A1 (n_4430), .B0 (n_4947), .Y (n_4998));
OAI21X1 g57393(.A0 (n_4205), .A1 (n_5105), .B0 (n_4949), .Y (n_4997));
OAI21X1 g57396(.A0 (n_3809), .A1 (n_5418), .B0 (n_4948), .Y (n_4996));
OAI21X1 g56606(.A0 (n_4458), .A1 (n_5239), .B0 (n_4946), .Y (n_4995));
NOR2X1 g56643(.A (WX5711), .B (n_5181), .Y (n_4994));
NOR2X1 g56645(.A (WX5711), .B (n_5500), .Y (n_4992));
MX2X1 g57508(.A (n_4963), .B (WX541), .S0 (n_6613), .Y (n_4991));
NOR2X1 g56683(.A (WX7004), .B (n_4882), .Y (n_8544));
NOR2X1 g56708(.A (WX7004), .B (n_2620), .Y (n_4988));
CLKBUFX1 gbuf_d_419(.A(n_4950), .Y(d_out_419));
CLKBUFX1 gbuf_q_419(.A(q_in_419), .Y(WX7126));
NOR2X1 g56744(.A (WX8297), .B (n_3690), .Y (n_4986));
NOR2X1 g56748(.A (WX8297), .B (n_5427), .Y (n_4985));
NOR2X1 g56808(.A (WX9590), .B (n_3188), .Y (n_4984));
NOR2X1 g56811(.A (WX9590), .B (n_5662), .Y (n_6695));
CLKBUFX1 gbuf_d_420(.A(n_4954), .Y(d_out_420));
CLKBUFX1 gbuf_q_420(.A(q_in_420), .Y(WX8417));
CLKBUFX1 gbuf_d_421(.A(n_4953), .Y(d_out_421));
CLKBUFX1 gbuf_q_421(.A(q_in_421), .Y(WX9708));
CLKBUFX1 gbuf_d_422(.A(n_4955), .Y(d_out_422));
CLKBUFX1 gbuf_q_422(.A(q_in_422), .Y(WX3253));
CLKBUFX1 gbuf_d_423(.A(n_4951), .Y(d_out_423));
CLKBUFX1 gbuf_q_423(.A(q_in_423), .Y(WX5835));
CLKBUFX1 gbuf_d_424(.A(n_4952), .Y(d_out_424));
CLKBUFX1 gbuf_q_424(.A(q_in_424), .Y(WX4544));
CLKBUFX1 gbuf_d_425(.A(n_4942), .Y(d_out_425));
CLKBUFX1 gbuf_q_425(.A(q_in_425), .Y(WX3289));
NAND2X1 g57200(.A (n_4944), .B (n_4745), .Y (n_4980));
OAI21X1 g56510(.A0 (n_4204), .A1 (n_12494), .B0 (n_5722), .Y(n_4979));
NAND2X2 g57328(.A (n_4941), .B (n_4690), .Y (n_4978));
CLKBUFX1 gbuf_d_426(.A(n_4938), .Y(d_out_426));
CLKBUFX1 gbuf_qn_426(.A(qn_in_426), .Y(WX8253));
CLKBUFX1 gbuf_d_427(.A(n_4935), .Y(d_out_427));
CLKBUFX1 gbuf_qn_427(.A(qn_in_427), .Y(WX9544));
CLKBUFX1 gbuf_d_428(.A(n_4934), .Y(d_out_428));
CLKBUFX1 gbuf_qn_428(.A(qn_in_428), .Y(WX4380));
CLKBUFX1 gbuf_d_429(.A(n_4930), .Y(d_out_429));
CLKBUFX1 gbuf_qn_429(.A(qn_in_429), .Y(WX5671));
CLKBUFX1 gbuf_d_430(.A(n_4927), .Y(d_out_430));
CLKBUFX1 gbuf_qn_430(.A(qn_in_430), .Y(WX6962));
CLKBUFX1 gbuf_d_431(.A(n_4925), .Y(d_out_431));
CLKBUFX1 gbuf_qn_431(.A(qn_in_431), .Y(WX3089));
NOR2X1 g57439(.A (WX10883), .B (n_5712), .Y (n_4976));
NOR2X1 g57440(.A (WX1832), .B (n_5712), .Y (n_4974));
NOR2X1 g57454(.A (WX1832), .B (n_5662), .Y (n_4973));
NOR2X1 g57458(.A (WX10883), .B (n_5479), .Y (n_7508));
NOR2X1 g56634(.A (WX4420), .B (n_5712), .Y (n_4970));
NOR2X1 g56637(.A (WX4420), .B (n_5479), .Y (n_15866));
OAI21X1 g56646(.A0 (n_4905), .A1 (n_4232), .B0 (n_4947), .Y (n_4968));
INVX1 g57510(.A (DATA_9_2), .Y (n_4966));
NOR2X1 g57544(.A (n_2849), .B (n_4963), .Y (n_4964));
OAI21X1 g56684(.A0 (n_4904), .A1 (n_10719), .B0 (n_5566), .Y(n_4962));
OR2X1 g57583(.A (n_4963), .B (n_5968), .Y (n_4961));
NAND2X2 g55783(.A (n_4943), .B (n_4728), .Y (n_4960));
OAI21X1 g56749(.A0 (n_4323), .A1 (n_8545), .B0 (n_5619), .Y (n_4959));
OAI21X1 g56812(.A0 (n_15867), .A1 (n_15868), .B0 (n_4860), .Y(n_4958));
CLKBUFX1 gbuf_d_432(.A(n_4923), .Y(d_out_432));
CLKBUFX1 gbuf_q_432(.A(q_in_432), .Y(WX5875));
CLKBUFX1 gbuf_d_433(.A(n_4922), .Y(d_out_433));
CLKBUFX1 gbuf_q_433(.A(q_in_433), .Y(WX7168));
CLKBUFX1 gbuf_d_434(.A(n_4921), .Y(d_out_434));
CLKBUFX1 gbuf_q_434(.A(q_in_434), .Y(WX8461));
CLKBUFX1 gbuf_d_435(.A(n_4920), .Y(d_out_435));
CLKBUFX1 gbuf_q_435(.A(q_in_435), .Y(WX9754));
NAND2X2 g55780(.A (n_4945), .B (n_4729), .Y (n_4956));
CLKBUFX1 gbuf_d_436(.A(n_4918), .Y(d_out_436));
CLKBUFX1 gbuf_qn_436(.A(qn_in_436), .Y(WX3125));
OAI21X1 g57387(.A0 (n_4636), .A1 (n_5841), .B0 (n_4917), .Y (n_4955));
OAI21X1 g57388(.A0 (n_4606), .A1 (n_5549), .B0 (n_4916), .Y (n_4954));
OAI21X1 g57390(.A0 (n_4544), .A1 (n_5415), .B0 (n_4915), .Y (n_4953));
OAI21X1 g57391(.A0 (n_4486), .A1 (n_5415), .B0 (n_4913), .Y (n_4952));
OAI21X1 g57392(.A0 (n_4427), .A1 (n_5439), .B0 (n_4912), .Y (n_4951));
OAI21X1 g57395(.A0 (n_4128), .A1 (n_5415), .B0 (n_4911), .Y (n_4950));
OAI21X1 g57455(.A0 (n_4887), .A1 (n_4139), .B0 (n_5460), .Y (n_4949));
OAI21X1 g57459(.A0 (n_4503), .A1 (n_6681), .B0 (n_4947), .Y (n_4948));
OAI21X1 g56638(.A0 (n_4883), .A1 (n_4570), .B0 (n_5460), .Y (n_4946));
OAI21X1 g57511(.A0 (n_4876), .A1 (n_5709), .B0 (n_4053), .Y(DATA_9_2));
CLKBUFX1 gbuf_d_437(.A(n_4906), .Y(d_out_437));
CLKBUFX1 gbuf_qn_437(.A(qn_in_437), .Y(WX5711));
CLKBUFX1 gbuf_d_438(.A(n_4903), .Y(d_out_438));
CLKBUFX1 gbuf_qn_438(.A(qn_in_438), .Y(WX7004));
CLKBUFX1 gbuf_d_439(.A(n_4902), .Y(d_out_439));
CLKBUFX1 gbuf_qn_439(.A(qn_in_439), .Y(WX8297));
CLKBUFX1 gbuf_d_440(.A(n_4907), .Y(d_out_440));
CLKBUFX1 gbuf_q_440(.A(q_in_440), .Y(WX4584));
CLKBUFX1 gbuf_d_441(.A(n_4908), .Y(d_out_441));
CLKBUFX1 gbuf_q_441(.A(q_in_441), .Y(WX11047));
CLKBUFX1 gbuf_d_442(.A(n_4909), .Y(d_out_442));
CLKBUFX1 gbuf_q_442(.A(q_in_442), .Y(WX1996));
CLKBUFX1 gbuf_d_443(.A(n_4899), .Y(d_out_443));
CLKBUFX1 gbuf_qn_443(.A(qn_in_443), .Y(WX9590));
NAND2X1 g55782(.A (n_6555), .B (n_8336), .Y (n_4945));
NAND2X1 g57233(.A (n_6583), .B (n_8337), .Y (n_4944));
NAND2X1 g55794(.A (n_4888), .B (n_6555), .Y (n_4943));
OAI21X1 g56543(.A0 (n_4571), .A1 (n_5600), .B0 (n_4893), .Y (n_4942));
NAND2X1 g57373(.A (n_6615), .B (n_8322), .Y (n_4941));
NOR2X1 g57434(.A (WX3091), .B (n_5500), .Y (n_4939));
NOR2X1 g57436(.A (WX8255), .B (n_5712), .Y (n_4938));
NOR2X1 g57437(.A (WX8255), .B (n_5500), .Y (n_4936));
NOR2X1 g57443(.A (WX9546), .B (n_3188), .Y (n_4935));
NOR2X1 g57444(.A (WX4382), .B (n_2851), .Y (n_4934));
NOR2X1 g57445(.A (WX9546), .B (n_4882), .Y (n_6231));
NOR2X1 g57447(.A (WX4382), .B (n_4882), .Y (n_6198));
NOR2X1 g57451(.A (WX5673), .B (n_2851), .Y (n_4930));
NOR2X1 g57452(.A (WX5673), .B (n_5479), .Y (n_6230));
NOR2X1 g57456(.A (WX6964), .B (n_1425), .Y (n_4927));
NOR2X1 g57460(.A (WX3091), .B (n_3188), .Y (n_4925));
NOR2X1 g57461(.A (WX6964), .B (n_5822), .Y (n_4924));
CLKBUFX1 gbuf_d_444(.A(n_4891), .Y(d_out_444));
CLKBUFX1 gbuf_qn_444(.A(qn_in_444), .Y(WX10883));
CLKBUFX1 gbuf_d_445(.A(n_4890), .Y(d_out_445));
CLKBUFX1 gbuf_qn_445(.A(qn_in_445), .Y(WX1832));
CLKBUFX1 gbuf_d_446(.A(n_4884), .Y(d_out_446));
CLKBUFX1 gbuf_qn_446(.A(qn_in_446), .Y(WX4420));
OAI21X1 g56667(.A0 (n_4209), .A1 (n_5468), .B0 (n_4881), .Y (n_4923));
INVX1 g57605(.A (WX541), .Y (n_4963));
OAI21X1 g56720(.A0 (n_4645), .A1 (n_5535), .B0 (n_4880), .Y (n_4922));
OAI21X1 g56780(.A0 (n_4279), .A1 (n_5439), .B0 (n_4879), .Y (n_4921));
OAI21X1 g56841(.A0 (n_4261), .A1 (n_5845), .B0 (n_4877), .Y (n_4920));
NOR2X1 g56569(.A (WX3127), .B (n_5811), .Y (n_12494));
NOR2X1 g56590(.A (WX3127), .B (n_1425), .Y (n_4918));
OAI21X1 g57435(.A0 (n_4473), .A1 (n_6232), .B0 (n_5556), .Y (n_4917));
OAI21X1 g57438(.A0 (n_4853), .A1 (n_4129), .B0 (n_5556), .Y (n_4916));
OAI21X1 g57446(.A0 (n_4607), .A1 (n_6199), .B0 (n_5619), .Y (n_4915));
OAI21X1 g57448(.A0 (n_4641), .A1 (n_6200), .B0 (n_5619), .Y (n_4913));
OAI21X1 g57453(.A0 (n_4489), .A1 (n_6676), .B0 (n_4860), .Y (n_4912));
OAI21X1 g57462(.A0 (n_4842), .A1 (n_4428), .B0 (n_5460), .Y (n_4911));
OAI21X1 g57496(.A0 (n_4203), .A1 (n_6050), .B0 (n_4861), .Y (n_4909));
OAI21X1 g57503(.A0 (n_3808), .A1 (n_5549), .B0 (n_4859), .Y (n_4908));
OAI21X1 g56665(.A0 (n_4456), .A1 (n_5598), .B0 (n_4858), .Y (n_4907));
CLKBUFX1 gbuf_d_447(.A(n_4875), .Y(d_out_447));
CLKBUFX1 gbuf_q_447(.A(q_in_447), .Y(WX541));
NOR2X1 g56701(.A (WX5713), .B (n_1648), .Y (n_4906));
NOR2X1 g56704(.A (WX5713), .B (n_5479), .Y (n_4905));
NOR2X1 g56742(.A (WX7006), .B (n_5662), .Y (n_4904));
NOR2X1 g56766(.A (WX7006), .B (n_5181), .Y (n_4903));
NOR2X1 g56803(.A (WX8299), .B (n_1425), .Y (n_4902));
NOR2X1 g56806(.A (WX8299), .B (n_5479), .Y (n_8545));
CLKBUFX1 gbuf_d_448(.A(n_4871), .Y(d_out_448));
CLKBUFX1 gbuf_q_448(.A(q_in_448), .Y(WX3255));
CLKBUFX1 gbuf_d_449(.A(n_4870), .Y(d_out_449));
CLKBUFX1 gbuf_q_449(.A(q_in_449), .Y(WX8419));
CLKBUFX1 gbuf_d_450(.A(n_4869), .Y(d_out_450));
CLKBUFX1 gbuf_q_450(.A(q_in_450), .Y(WX9710));
CLKBUFX1 gbuf_d_451(.A(n_4867), .Y(d_out_451));
CLKBUFX1 gbuf_q_451(.A(q_in_451), .Y(WX4546));
CLKBUFX1 gbuf_d_452(.A(n_4865), .Y(d_out_452));
CLKBUFX1 gbuf_q_452(.A(q_in_452), .Y(WX5837));
CLKBUFX1 gbuf_d_453(.A(n_4864), .Y(d_out_453));
CLKBUFX1 gbuf_q_453(.A(q_in_453), .Y(WX7128));
NOR2X1 g56867(.A (WX9592), .B (n_2620), .Y (n_4899));
NOR2X1 g56871(.A (WX9592), .B (n_5479), .Y (n_15868));
OAI21X1 g55784(.A0 (n_4790), .A1 (n_5889), .B0 (n_3653), .Y (n_8336));
OAI21X1 g57261(.A0 (n_4827), .A1 (n_5889), .B0 (n_3600), .Y (n_8337));
OAI21X1 g56570(.A0 (n_4819), .A1 (n_11600), .B0 (n_5722), .Y(n_4893));
OAI21X1 g57399(.A0 (n_4801), .A1 (n_5889), .B0 (n_3692), .Y (n_8322));
CLKBUFX1 gbuf_d_454(.A(n_4854), .Y(d_out_454));
CLKBUFX1 gbuf_qn_454(.A(qn_in_454), .Y(WX8255));
CLKBUFX1 gbuf_d_455(.A(n_4852), .Y(d_out_455));
CLKBUFX1 gbuf_qn_455(.A(qn_in_455), .Y(WX9546));
CLKBUFX1 gbuf_d_456(.A(n_4851), .Y(d_out_456));
CLKBUFX1 gbuf_qn_456(.A(qn_in_456), .Y(WX4382));
CLKBUFX1 gbuf_d_457(.A(n_4848), .Y(d_out_457));
CLKBUFX1 gbuf_qn_457(.A(qn_in_457), .Y(WX5673));
CLKBUFX1 gbuf_d_458(.A(n_4845), .Y(d_out_458));
CLKBUFX1 gbuf_qn_458(.A(qn_in_458), .Y(WX6964));
CLKBUFX1 gbuf_d_459(.A(n_4844), .Y(d_out_459));
CLKBUFX1 gbuf_qn_459(.A(qn_in_459), .Y(WX3091));
NOR2X1 g57524(.A (WX10885), .B (n_5712), .Y (n_4891));
NOR2X1 g57526(.A (WX1834), .B (n_3188), .Y (n_4890));
OAI21X1 g55804(.A0 (n_4832), .A1 (n_5889), .B0 (n_3686), .Y (n_4888));
NOR2X1 g57551(.A (WX1834), .B (n_4882), .Y (n_4887));
NOR2X1 g57588(.A (WX10885), .B (n_5838), .Y (n_6681));
NOR2X1 g56693(.A (WX4422), .B (n_3690), .Y (n_4884));
NOR2X1 g56696(.A (WX4422), .B (n_4882), .Y (n_4883));
OAI21X1 g56705(.A0 (n_4786), .A1 (n_4457), .B0 (n_4860), .Y (n_4881));
OAI21X1 g56743(.A0 (n_4208), .A1 (n_9438), .B0 (n_5275), .Y (n_4880));
OAI21X1 g56807(.A0 (n_4775), .A1 (n_4643), .B0 (n_5722), .Y (n_4879));
CLKBUFX1 gbuf_d_460(.A(n_4857), .Y(d_out_460));
CLKBUFX1 gbuf_q_460(.A(q_in_460), .Y(WX3291));
CLKBUFX1 gbuf_d_461(.A(n_4841), .Y(d_out_461));
CLKBUFX1 gbuf_q_461(.A(q_in_461), .Y(WX5877));
CLKBUFX1 gbuf_d_462(.A(n_4840), .Y(d_out_462));
CLKBUFX1 gbuf_q_462(.A(q_in_462), .Y(WX7170));
CLKBUFX1 gbuf_d_463(.A(n_4839), .Y(d_out_463));
CLKBUFX1 gbuf_q_463(.A(q_in_463), .Y(WX8463));
CLKBUFX1 gbuf_d_464(.A(n_4838), .Y(d_out_464));
CLKBUFX1 gbuf_q_464(.A(q_in_464), .Y(WX9756));
OAI21X1 g56872(.A0 (n_4835), .A1 (n_11602), .B0 (n_6497), .Y(n_4877));
MX2X1 g57867(.A (n_4874), .B (WX543), .S0 (n_4052), .Y (n_4876));
NOR2X1 g58169(.A (n_1425), .B (n_4874), .Y (n_4875));
OR2X1 g58174(.A (n_4874), .B (n_5990), .Y (n_4873));
CLKBUFX1 gbuf_d_465(.A(n_4828), .Y(d_out_465));
CLKBUFX1 gbuf_q_465(.A(q_in_465), .Y(WX1938));
CLKBUFX1 gbuf_d_466(.A(n_4816), .Y(d_out_466));
CLKBUFX1 gbuf_q_466(.A(q_in_466), .Y(WX9716));
CLKBUFX1 gbuf_d_467(.A(n_4820), .Y(d_out_467));
CLKBUFX1 gbuf_q_467(.A(q_in_467), .Y(WX8425));
CLKBUFX1 gbuf_d_468(.A(n_4823), .Y(d_out_468));
CLKBUFX1 gbuf_q_468(.A(q_in_468), .Y(WX3261));
CLKBUFX1 gbuf_d_469(.A(n_4802), .Y(d_out_469));
CLKBUFX1 gbuf_qn_469(.A(qn_in_469), .Y(WX3127));
OAI21X1 g57476(.A0 (n_4633), .A1 (n_5317), .B0 (n_4799), .Y (n_4871));
OAI21X1 g57480(.A0 (n_4604), .A1 (n_5317), .B0 (n_4797), .Y (n_4870));
OAI21X1 g57484(.A0 (n_4542), .A1 (n_4868), .B0 (n_4796), .Y (n_4869));
OAI21X1 g57488(.A0 (n_4255), .A1 (n_4866), .B0 (n_4795), .Y (n_4867));
OAI21X1 g57492(.A0 (n_4423), .A1 (n_5185), .B0 (n_4794), .Y (n_4865));
OAI21X1 g57499(.A0 (n_4373), .A1 (n_5482), .B0 (n_4793), .Y (n_4864));
INVX1 g57512(.A (DATA_9_1), .Y (n_4863));
OAI21X1 g57552(.A0 (n_4765), .A1 (n_4137), .B0 (n_4860), .Y (n_4861));
OAI21X1 g57589(.A0 (n_4260), .A1 (n_7509), .B0 (n_5722), .Y (n_4859));
OAI21X1 g56697(.A0 (n_4758), .A1 (n_4568), .B0 (n_4860), .Y (n_4858));
CLKBUFX1 gbuf_d_470(.A(n_4788), .Y(d_out_470));
CLKBUFX1 gbuf_qn_470(.A(qn_in_470), .Y(WX5713));
CLKBUFX1 gbuf_d_471(.A(n_4781), .Y(d_out_471));
CLKBUFX1 gbuf_qn_471(.A(qn_in_471), .Y(WX7006));
CLKBUFX1 gbuf_d_472(.A(n_4798), .Y(d_out_472));
CLKBUFX1 gbuf_q_472(.A(q_in_472), .Y(WX3293));
CLKBUFX1 gbuf_d_473(.A(n_4792), .Y(d_out_473));
CLKBUFX1 gbuf_q_473(.A(q_in_473), .Y(WX4586));
CLKBUFX1 gbuf_d_474(.A(n_4791), .Y(d_out_474));
CLKBUFX1 gbuf_q_474(.A(q_in_474), .Y(WX3231));
CLKBUFX1 gbuf_d_475(.A(n_4785), .Y(d_out_475));
CLKBUFX1 gbuf_q_475(.A(q_in_475), .Y(WX4524));
CLKBUFX1 gbuf_d_476(.A(n_4784), .Y(d_out_476));
CLKBUFX1 gbuf_q_476(.A(q_in_476), .Y(WX5879));
CLKBUFX1 gbuf_d_477(.A(n_4783), .Y(d_out_477));
CLKBUFX1 gbuf_q_477(.A(q_in_477), .Y(WX3233));
CLKBUFX1 gbuf_d_478(.A(n_4780), .Y(d_out_478));
CLKBUFX1 gbuf_q_478(.A(q_in_478), .Y(WX7172));
CLKBUFX1 gbuf_d_479(.A(n_4779), .Y(d_out_479));
CLKBUFX1 gbuf_q_479(.A(q_in_479), .Y(WX4526));
CLKBUFX1 gbuf_d_480(.A(n_4778), .Y(d_out_480));
CLKBUFX1 gbuf_q_480(.A(q_in_480), .Y(WX5817));
CLKBUFX1 gbuf_d_481(.A(n_4774), .Y(d_out_481));
CLKBUFX1 gbuf_q_481(.A(q_in_481), .Y(WX8465));
CLKBUFX1 gbuf_d_482(.A(n_4773), .Y(d_out_482));
CLKBUFX1 gbuf_q_482(.A(q_in_482), .Y(WX5819));
CLKBUFX1 gbuf_d_483(.A(n_4772), .Y(d_out_483));
CLKBUFX1 gbuf_q_483(.A(q_in_483), .Y(WX7110));
CLKBUFX1 gbuf_d_484(.A(n_4834), .Y(d_out_484));
CLKBUFX1 gbuf_q_484(.A(q_in_484), .Y(WX8403));
CLKBUFX1 gbuf_d_485(.A(n_4833), .Y(d_out_485));
CLKBUFX1 gbuf_q_485(.A(q_in_485), .Y(WX7112));
CLKBUFX1 gbuf_d_486(.A(n_4830), .Y(d_out_486));
CLKBUFX1 gbuf_q_486(.A(q_in_486), .Y(WX8405));
CLKBUFX1 gbuf_d_487(.A(n_4829), .Y(d_out_487));
CLKBUFX1 gbuf_q_487(.A(q_in_487), .Y(WX9698));
CLKBUFX1 gbuf_d_488(.A(n_4804), .Y(d_out_488));
CLKBUFX1 gbuf_q_488(.A(q_in_488), .Y(WX11049));
CLKBUFX1 gbuf_d_489(.A(n_4824), .Y(d_out_489));
CLKBUFX1 gbuf_q_489(.A(q_in_489), .Y(WX3259));
CLKBUFX1 gbuf_d_490(.A(n_4825), .Y(d_out_490));
CLKBUFX1 gbuf_q_490(.A(q_in_490), .Y(WX3257));
CLKBUFX1 gbuf_d_491(.A(n_4822), .Y(d_out_491));
CLKBUFX1 gbuf_q_491(.A(q_in_491), .Y(WX8421));
CLKBUFX1 gbuf_d_492(.A(n_4821), .Y(d_out_492));
CLKBUFX1 gbuf_q_492(.A(q_in_492), .Y(WX8423));
CLKBUFX1 gbuf_d_493(.A(n_4817), .Y(d_out_493));
CLKBUFX1 gbuf_q_493(.A(q_in_493), .Y(WX9714));
CLKBUFX1 gbuf_d_494(.A(n_4818), .Y(d_out_494));
CLKBUFX1 gbuf_q_494(.A(q_in_494), .Y(WX9712));
CLKBUFX1 gbuf_d_495(.A(n_4814), .Y(d_out_495));
CLKBUFX1 gbuf_q_495(.A(q_in_495), .Y(WX4550));
CLKBUFX1 gbuf_d_496(.A(n_4815), .Y(d_out_496));
CLKBUFX1 gbuf_q_496(.A(q_in_496), .Y(WX4548));
CLKBUFX1 gbuf_d_497(.A(n_4811), .Y(d_out_497));
CLKBUFX1 gbuf_q_497(.A(q_in_497), .Y(WX5841));
CLKBUFX1 gbuf_d_498(.A(n_4812), .Y(d_out_498));
CLKBUFX1 gbuf_q_498(.A(q_in_498), .Y(WX5839));
CLKBUFX1 gbuf_d_499(.A(n_4809), .Y(d_out_499));
CLKBUFX1 gbuf_q_499(.A(q_in_499), .Y(WX1998));
CLKBUFX1 gbuf_d_500(.A(n_4808), .Y(d_out_500));
CLKBUFX1 gbuf_q_500(.A(q_in_500), .Y(WX2000));
CLKBUFX1 gbuf_d_501(.A(n_4807), .Y(d_out_501));
CLKBUFX1 gbuf_q_501(.A(q_in_501), .Y(WX7130));
CLKBUFX1 gbuf_d_502(.A(n_4806), .Y(d_out_502));
CLKBUFX1 gbuf_q_502(.A(q_in_502), .Y(WX7132));
CLKBUFX1 gbuf_d_503(.A(n_4805), .Y(d_out_503));
CLKBUFX1 gbuf_q_503(.A(q_in_503), .Y(WX7134));
CLKBUFX1 gbuf_d_504(.A(n_4777), .Y(d_out_504));
CLKBUFX1 gbuf_qn_504(.A(qn_in_504), .Y(WX8299));
CLKBUFX1 gbuf_d_505(.A(n_4813), .Y(d_out_505));
CLKBUFX1 gbuf_q_505(.A(q_in_505), .Y(WX4552));
CLKBUFX1 gbuf_d_506(.A(n_4810), .Y(d_out_506));
CLKBUFX1 gbuf_q_506(.A(q_in_506), .Y(WX5843));
CLKBUFX1 gbuf_d_507(.A(n_4837), .Y(d_out_507));
CLKBUFX1 gbuf_qn_507(.A(qn_in_507), .Y(WX9592));
CLKBUFX1 gbuf_d_508(.A(n_4760), .Y(d_out_508));
CLKBUFX1 gbuf_q_508(.A(q_in_508), .Y(WX11051));
OAI21X1 g56603(.A0 (n_4569), .A1 (n_5158), .B0 (n_4761), .Y (n_4857));
OAI21X1 g57513(.A0 (n_4679), .A1 (n_5965), .B0 (n_4051), .Y(DATA_9_1));
NOR2X1 g57516(.A (WX3093), .B (n_5500), .Y (n_6232));
NOR2X1 g57521(.A (WX8257), .B (n_1425), .Y (n_4854));
NOR2X1 g57522(.A (WX8257), .B (n_5500), .Y (n_4853));
NOR2X1 g57529(.A (WX9548), .B (n_1648), .Y (n_4852));
NOR2X1 g57530(.A (WX4384), .B (n_5712), .Y (n_4851));
NOR2X1 g57531(.A (WX9548), .B (n_5500), .Y (n_6199));
NOR2X1 g57536(.A (WX4384), .B (n_5838), .Y (n_6200));
NOR2X1 g57545(.A (WX5675), .B (n_3690), .Y (n_4848));
NOR2X1 g57546(.A (WX5675), .B (n_4882), .Y (n_6676));
NOR2X1 g57580(.A (WX6966), .B (n_3690), .Y (n_4845));
NOR2X1 g57590(.A (WX3093), .B (n_1648), .Y (n_4844));
NOR2X1 g57591(.A (WX6966), .B (n_4670), .Y (n_4842));
CLKBUFX1 gbuf_d_509(.A(n_4768), .Y(d_out_509));
CLKBUFX1 gbuf_qn_509(.A(qn_in_509), .Y(WX1834));
CLKBUFX1 gbuf_d_510(.A(n_4769), .Y(d_out_510));
CLKBUFX1 gbuf_qn_510(.A(qn_in_510), .Y(WX10885));
CLKBUFX1 gbuf_d_511(.A(n_4759), .Y(d_out_511));
CLKBUFX1 gbuf_qn_511(.A(qn_in_511), .Y(WX4422));
OAI21X1 g56725(.A0 (n_4207), .A1 (n_5439), .B0 (n_4756), .Y (n_4841));
OAI21X1 g56779(.A0 (n_4640), .A1 (n_5729), .B0 (n_4755), .Y (n_4840));
CLKBUFX1 gbuf_d_512(.A(n_4762), .Y(d_out_512));
CLKBUFX1 gbuf_q_512(.A(q_in_512), .Y(WX10991));
CLKBUFX1 gbuf_d_513(.A(n_4757), .Y(d_out_513));
CLKBUFX1 gbuf_q_513(.A(q_in_513), .Y(WX1940));
CLKBUFX1 gbuf_d_514(.A(n_4770), .Y(d_out_514));
CLKBUFX1 gbuf_q_514(.A(q_in_514), .Y(WX9758));
OAI21X1 g56839(.A0 (n_4560), .A1 (n_5085), .B0 (n_4754), .Y (n_4839));
CLKBUFX1 gbuf_d_515(.A(n_4766), .Y(d_out_515));
CLKBUFX1 gbuf_q_515(.A(q_in_515), .Y(WX9696));
OAI21X1 g56899(.A0 (n_4259), .A1 (n_5334), .B0 (n_4771), .Y (n_4838));
NOR2X1 g56926(.A (WX9594), .B (n_1425), .Y (n_4837));
NOR2X1 g56929(.A (WX9594), .B (n_5427), .Y (n_4835));
CLKBUFX1 gbuf_d_516(.A(n_4746), .Y(d_out_516));
CLKBUFX1 gbuf_q_516(.A(q_in_516), .Y(WX10989));
OAI21X1 g56956(.A0 (n_4319), .A1 (n_6050), .B0 (n_4750), .Y (n_4834));
OAI21X1 g56961(.A0 (n_4383), .A1 (n_4868), .B0 (n_4749), .Y (n_4833));
INVX1 g55845(.A (DATA_9_29), .Y (n_4832));
OAI21X1 g57015(.A0 (n_4618), .A1 (n_4866), .B0 (n_4748), .Y (n_4830));
INVX1 g58206(.A (WX543), .Y (n_4874));
OAI21X1 g57075(.A0 (n_4275), .A1 (n_5183), .B0 (n_4747), .Y (n_4829));
OAI21X1 g57320(.A0 (n_4596), .A1 (n_5918), .B0 (n_4652), .Y (n_4828));
INVX1 g57331(.A (DATA_9_31), .Y (n_4827));
OAI21X1 g57477(.A0 (n_4631), .A1 (n_5928), .B0 (n_4651), .Y (n_4825));
OAI21X1 g57478(.A0 (n_4629), .A1 (n_5841), .B0 (n_4744), .Y (n_4824));
OAI21X1 g57479(.A0 (n_4624), .A1 (n_5439), .B0 (n_4743), .Y (n_4823));
OAI21X1 g57481(.A0 (n_4601), .A1 (n_4866), .B0 (n_4742), .Y (n_4822));
OAI21X1 g57482(.A0 (n_4598), .A1 (n_5474), .B0 (n_4741), .Y (n_4821));
OAI21X1 g57483(.A0 (n_4594), .A1 (n_5418), .B0 (n_4740), .Y (n_4820));
NOR2X1 g56629(.A (WX3129), .B (n_4882), .Y (n_4819));
OAI21X1 g57485(.A0 (n_4538), .A1 (n_5892), .B0 (n_4739), .Y (n_4818));
OAI21X1 g57486(.A0 (n_4626), .A1 (n_5490), .B0 (n_4738), .Y (n_4817));
OAI21X1 g57487(.A0 (n_4536), .A1 (n_4868), .B0 (n_4737), .Y (n_4816));
OAI21X1 g57489(.A0 (n_4484), .A1 (n_5535), .B0 (n_4736), .Y (n_4815));
OAI21X1 g57490(.A0 (n_4482), .A1 (n_5415), .B0 (n_4735), .Y (n_4814));
OAI21X1 g57491(.A0 (n_4480), .A1 (n_5482), .B0 (n_4734), .Y (n_4813));
OAI21X1 g57493(.A0 (n_4421), .A1 (n_5196), .B0 (n_4650), .Y (n_4812));
OAI21X1 g57494(.A0 (n_4416), .A1 (n_5493), .B0 (n_4733), .Y (n_4811));
OAI21X1 g57495(.A0 (n_4414), .A1 (n_5185), .B0 (n_4731), .Y (n_4810));
OAI21X1 g57497(.A0 (n_4201), .A1 (n_5576), .B0 (n_4730), .Y (n_4809));
OAI21X1 g57498(.A0 (n_4387), .A1 (n_5882), .B0 (n_4649), .Y (n_4808));
OAI21X1 g57500(.A0 (n_4371), .A1 (n_5598), .B0 (n_4689), .Y (n_4807));
OAI21X1 g57501(.A0 (n_4369), .A1 (n_5493), .B0 (n_4687), .Y (n_4806));
OAI21X1 g57502(.A0 (n_4365), .A1 (n_5882), .B0 (n_4686), .Y (n_4805));
OAI21X1 g57504(.A0 (n_3807), .A1 (n_4803), .B0 (n_4688), .Y (n_4804));
NOR2X1 g56650(.A (WX3129), .B (n_1425), .Y (n_4802));
INVX1 g57514(.A (DATA_9_0), .Y (n_4801));
OAI21X1 g57517(.A0 (n_4677), .A1 (n_4463), .B0 (n_5460), .Y (n_4799));
OAI21X1 g56662(.A0 (n_4567), .A1 (n_5235), .B0 (n_4696), .Y (n_4798));
OAI21X1 g57523(.A0 (n_4674), .A1 (n_4127), .B0 (n_5460), .Y (n_4797));
OAI21X1 g57532(.A0 (n_4605), .A1 (n_6660), .B0 (n_5566), .Y (n_4796));
OAI21X1 g57538(.A0 (n_4671), .A1 (n_4634), .B0 (n_5566), .Y (n_4795));
OAI21X1 g57547(.A0 (n_4485), .A1 (n_6201), .B0 (n_4947), .Y (n_4794));
OAI21X1 g57592(.A0 (n_4426), .A1 (n_6668), .B0 (n_4947), .Y (n_4793));
OAI21X1 g56723(.A0 (n_4454), .A1 (n_5729), .B0 (n_4685), .Y (n_4792));
OAI21X1 g56726(.A0 (n_4125), .A1 (n_5439), .B0 (n_4684), .Y (n_4791));
INVX1 g55805(.A (DATA_9_30), .Y (n_4790));
NOR2X1 g56759(.A (WX5715), .B (n_1425), .Y (n_4788));
NOR2X1 g56762(.A (WX5715), .B (n_5427), .Y (n_4786));
OAI21X1 g56781(.A0 (n_4540), .A1 (n_4803), .B0 (n_4419), .Y (n_4785));
OAI21X1 g56784(.A0 (n_4390), .A1 (n_5750), .B0 (n_4683), .Y (n_4784));
OAI21X1 g56785(.A0 (n_4367), .A1 (n_5750), .B0 (n_4388), .Y (n_4783));
NOR2X1 g56801(.A (WX7008), .B (n_5427), .Y (n_9438));
NOR2X1 g56824(.A (WX7008), .B (n_2851), .Y (n_4781));
OAI21X1 g56838(.A0 (n_4638), .A1 (n_5535), .B0 (n_4682), .Y (n_4780));
OAI21X1 g56840(.A0 (n_4528), .A1 (n_5535), .B0 (n_4681), .Y (n_4779));
OAI21X1 g56842(.A0 (n_4446), .A1 (n_4803), .B0 (n_4680), .Y (n_4778));
NOR2X1 g56862(.A (WX8301), .B (n_5712), .Y (n_4777));
NOR2X1 g56865(.A (WX8301), .B (n_5479), .Y (n_4775));
OAI21X1 g56897(.A0 (n_4277), .A1 (n_5393), .B0 (n_4753), .Y (n_4774));
OAI21X1 g56900(.A0 (n_4444), .A1 (n_5535), .B0 (n_4752), .Y (n_4773));
OAI21X1 g56902(.A0 (n_4385), .A1 (n_5468), .B0 (n_4751), .Y (n_4772));
OAI21X1 g56930(.A0 (n_4332), .A1 (n_4559), .B0 (n_4947), .Y (n_4771));
OAI21X1 g56958(.A0 (n_4257), .A1 (n_5196), .B0 (n_4678), .Y (n_4770));
OAI21X1 g55846(.A0 (n_4178), .A1 (n_5843), .B0 (n_4037), .Y(DATA_9_29));
NOR2X1 g58163(.A (WX10887), .B (n_5712), .Y (n_4769));
NOR2X1 g58164(.A (WX1836), .B (n_1648), .Y (n_4768));
OAI21X1 g57016(.A0 (n_4088), .A1 (n_5439), .B0 (n_4660), .Y (n_4766));
NOR2X1 g58172(.A (WX1836), .B (n_4882), .Y (n_4765));
NOR2X1 g58176(.A (WX10887), .B (n_6438), .Y (n_7509));
CLKBUFX1 gbuf_d_517(.A(n_4657), .Y(d_out_517));
CLKBUFX1 gbuf_q_517(.A(q_in_517), .Y(WX543));
OAI21X1 g57332(.A0 (n_4328), .A1 (n_5242), .B0 (n_4086), .Y(DATA_9_31));
OAI21X1 g55803(.A0 (n_3842), .A1 (n_5183), .B0 (n_4658), .Y (n_4762));
OAI21X1 g56630(.A0 (n_4327), .A1 (n_10721), .B0 (n_5556), .Y(n_4761));
OAI21X1 g57505(.A0 (n_3806), .A1 (n_4803), .B0 (n_4648), .Y (n_4760));
OAI21X1 g57515(.A0 (n_4109), .A1 (n_6091), .B0 (n_4047), .Y(DATA_9_0));
CLKBUFX1 gbuf_d_518(.A(n_4676), .Y(d_out_518));
CLKBUFX1 gbuf_qn_518(.A(qn_in_518), .Y(WX8257));
CLKBUFX1 gbuf_d_519(.A(n_4673), .Y(d_out_519));
CLKBUFX1 gbuf_qn_519(.A(qn_in_519), .Y(WX9548));
CLKBUFX1 gbuf_d_520(.A(n_4672), .Y(d_out_520));
CLKBUFX1 gbuf_qn_520(.A(qn_in_520), .Y(WX4384));
CLKBUFX1 gbuf_d_521(.A(n_4669), .Y(d_out_521));
CLKBUFX1 gbuf_qn_521(.A(qn_in_521), .Y(WX5675));
CLKBUFX1 gbuf_d_522(.A(n_4667), .Y(d_out_522));
CLKBUFX1 gbuf_qn_522(.A(qn_in_522), .Y(WX6966));
CLKBUFX1 gbuf_d_523(.A(n_4665), .Y(d_out_523));
CLKBUFX1 gbuf_qn_523(.A(qn_in_523), .Y(WX3093));
OAI21X1 g55806(.A0 (n_4334), .A1 (n_5242), .B0 (n_4031), .Y(DATA_9_30));
NOR2X1 g56751(.A (WX4424), .B (n_5712), .Y (n_4759));
NOR2X1 g56754(.A (WX4424), .B (n_5838), .Y (n_4758));
OAI21X1 g55796(.A0 (n_4295), .A1 (n_5183), .B0 (n_4659), .Y (n_4757));
OAI21X1 g56763(.A0 (n_4455), .A1 (n_6684), .B0 (n_5722), .Y (n_4756));
OAI21X1 g56802(.A0 (n_4126), .A1 (n_11604), .B0 (n_5275), .Y(n_4755));
OAI21X1 g56866(.A0 (n_4335), .A1 (n_4639), .B0 (n_5722), .Y (n_4754));
OAI21X1 g56924(.A0 (n_3845), .A1 (n_9419), .B0 (n_6497), .Y (n_4753));
OAI21X1 g56934(.A0 (n_4527), .A1 (n_6202), .B0 (n_5460), .Y (n_4752));
OAI21X1 g56942(.A0 (n_6886), .A1 (n_6213), .B0 (n_4947), .Y (n_4751));
CLKBUFX1 gbuf_d_524(.A(n_4333), .Y(d_out_524));
CLKBUFX1 gbuf_qn_524(.A(qn_in_524), .Y(WX9594));
OAI21X1 g56979(.A0 (n_4384), .A1 (n_6183), .B0 (n_4947), .Y (n_4750));
OAI21X1 g57001(.A0 (n_3639), .A1 (n_6451), .B0 (n_5566), .Y (n_4749));
OAI21X1 g57039(.A0 (n_4382), .A1 (n_6670), .B0 (n_5460), .Y (n_4748));
OAI21X1 g57104(.A0 (n_4617), .A1 (n_6203), .B0 (n_4860), .Y (n_4747));
OAI21X1 g57329(.A0 (n_3843), .A1 (n_5105), .B0 (n_4331), .Y (n_4746));
OR2X1 g57366(.A (n_4330), .B (n_4697), .Y (n_4745));
OAI21X1 g57519(.A0 (n_3447), .A1 (n_4459), .B0 (n_4947), .Y (n_4744));
CLKBUFX1 gbuf_d_525(.A(n_4320), .Y(d_out_525));
CLKBUFX1 gbuf_qn_525(.A(qn_in_525), .Y(WX3129));
OAI21X1 g57520(.A0 (n_3433), .A1 (n_4451), .B0 (n_5619), .Y (n_4743));
OAI21X1 g57525(.A0 (n_4372), .A1 (n_6662), .B0 (n_5460), .Y (n_4742));
OAI21X1 g57527(.A0 (n_4370), .A1 (n_6663), .B0 (n_5460), .Y (n_4741));
OAI21X1 g57528(.A0 (n_3601), .A1 (n_4368), .B0 (n_5556), .Y (n_4740));
OAI21X1 g57533(.A0 (n_3850), .A1 (n_4602), .B0 (n_4860), .Y (n_4739));
OAI21X1 g57534(.A0 (n_4599), .A1 (n_6204), .B0 (n_3183), .Y (n_4738));
OAI21X1 g57535(.A0 (n_4597), .A1 (n_6661), .B0 (n_4860), .Y (n_4737));
OAI21X1 g57539(.A0 (n_3857), .A1 (n_6632), .B0 (n_5460), .Y (n_4736));
OAI21X1 g57540(.A0 (n_4630), .A1 (n_6205), .B0 (n_5722), .Y (n_4735));
OAI21X1 g57542(.A0 (n_3434), .A1 (n_4627), .B0 (n_5566), .Y (n_4734));
OAI21X1 g57549(.A0 (n_4483), .A1 (n_6206), .B0 (n_6479), .Y (n_4733));
OAI21X1 g57550(.A0 (n_4481), .A1 (n_6208), .B0 (n_4860), .Y (n_4731));
OAI21X1 g57553(.A0 (n_4090), .A1 (n_4135), .B0 (n_5722), .Y (n_4730));
OR2X1 g57554(.A (n_4199), .B (n_4697), .Y (n_4729));
OR2X1 g57555(.A (n_4197), .B (n_4697), .Y (n_4728));
OR2X1 g57556(.A (n_4194), .B (n_4697), .Y (n_4727));
OR2X1 g57557(.A (n_4192), .B (n_4697), .Y (n_4725));
OR2X1 g57558(.A (n_4190), .B (n_4697), .Y (n_4723));
OR2X1 g57559(.A (n_4187), .B (n_4697), .Y (n_4722));
OR2X1 g57560(.A (n_4185), .B (n_4697), .Y (n_4721));
OR2X1 g57561(.A (n_4182), .B (n_4697), .Y (n_4720));
OR2X1 g57563(.A (n_4180), .B (n_4697), .Y (n_4719));
OR2X1 g57564(.A (n_4177), .B (n_4697), .Y (n_4717));
OR2X1 g57565(.A (n_4175), .B (n_4697), .Y (n_4716));
OR2X1 g57566(.A (n_4173), .B (n_4697), .Y (n_4715));
OR2X1 g57567(.A (n_4171), .B (n_4697), .Y (n_4714));
OR2X1 g57568(.A (n_4169), .B (n_4697), .Y (n_15853));
OR2X1 g57569(.A (n_4167), .B (n_4697), .Y (n_4711));
OR2X1 g57572(.A (n_4161), .B (n_4697), .Y (n_4706));
OR2X1 g57573(.A (n_4159), .B (n_4697), .Y (n_4704));
OR2X1 g57575(.A (n_4155), .B (n_4697), .Y (n_4702));
OR2X1 g57579(.A (n_4146), .B (n_4697), .Y (n_4698));
OAI21X1 g56689(.A0 (n_3698), .A1 (n_4386), .B0 (n_5566), .Y (n_4696));
OR2X1 g57581(.A (n_4144), .B (n_4697), .Y (n_4695));
OR2X1 g57584(.A (n_4140), .B (n_4697), .Y (n_4693));
OR2X1 g57585(.A (n_4138), .B (n_4697), .Y (n_4692));
OR2X1 g57587(.A (n_4134), .B (n_4697), .Y (n_4690));
OAI21X1 g57593(.A0 (n_4422), .A1 (n_6207), .B0 (n_5460), .Y (n_4689));
OAI21X1 g57594(.A0 (n_4258), .A1 (n_7510), .B0 (n_5706), .Y (n_4688));
OAI21X1 g57595(.A0 (n_4420), .A1 (n_6677), .B0 (n_4947), .Y (n_4687));
OAI21X1 g57596(.A0 (n_4415), .A1 (n_6664), .B0 (n_5619), .Y (n_4686));
OAI21X1 g56755(.A0 (n_4083), .A1 (n_4566), .B0 (n_5566), .Y (n_4685));
OAI21X1 g56768(.A0 (n_4595), .A1 (n_6182), .B0 (n_4860), .Y (n_4684));
CLKBUFX1 gbuf_d_526(.A(n_4221), .Y(d_out_526));
CLKBUFX1 gbuf_qn_526(.A(qn_in_526), .Y(WX5715));
CLKBUFX1 gbuf_d_527(.A(n_4108), .Y(d_out_527));
CLKBUFX1 gbuf_qn_527(.A(qn_in_527), .Y(WX7008));
OAI21X1 g56821(.A0 (n_3689), .A1 (n_10723), .B0 (n_4860), .Y(n_4683));
OAI21X1 g56861(.A0 (n_3688), .A1 (n_4389), .B0 (n_4860), .Y (n_4682));
OAI21X1 g56870(.A0 (n_4366), .A1 (n_6669), .B0 (n_7087), .Y (n_4681));
OAI21X1 g56876(.A0 (n_4539), .A1 (n_6212), .B0 (n_5722), .Y (n_4680));
MX2X1 g57868(.A (n_4656), .B (WX545), .S0 (n_4050), .Y (n_4679));
CLKBUFX1 gbuf_d_528(.A(n_4107), .Y(d_out_528));
CLKBUFX1 gbuf_qn_528(.A(qn_in_528), .Y(WX8301));
OAI21X1 g56988(.A0 (n_4276), .A1 (n_8546), .B0 (n_4860), .Y (n_4678));
NOR2X1 g58159(.A (WX3095), .B (n_5662), .Y (n_4677));
NOR2X1 g58160(.A (WX8259), .B (n_1648), .Y (n_4676));
NOR2X1 g58161(.A (WX9550), .B (n_6438), .Y (n_6660));
NOR2X1 g58162(.A (WX8259), .B (n_4882), .Y (n_4674));
NOR2X1 g58165(.A (WX9550), .B (n_2851), .Y (n_4673));
NOR2X1 g58166(.A (WX4386), .B (n_2620), .Y (n_4672));
NOR2X1 g58168(.A (WX4386), .B (n_4670), .Y (n_4671));
NOR2X1 g58170(.A (WX5677), .B (n_1648), .Y (n_4669));
NOR2X1 g58171(.A (WX5677), .B (n_4670), .Y (n_6201));
NOR2X1 g58173(.A (WX6968), .B (n_1648), .Y (n_4667));
NOR2X1 g58175(.A (WX3095), .B (n_3690), .Y (n_4665));
NOR2X1 g58177(.A (WX6968), .B (n_6438), .Y (n_6668));
CLKBUFX1 gbuf_d_529(.A(n_4093), .Y(d_out_529));
CLKBUFX1 gbuf_qn_529(.A(qn_in_529), .Y(WX1836));
CLKBUFX1 gbuf_d_530(.A(n_4092), .Y(d_out_530));
CLKBUFX1 gbuf_qn_530(.A(qn_in_530), .Y(WX10887));
AOI21X1 g57785(.A0 (_2210_), .A1 (n_4608), .B0 (n_4661), .Y (n_4662));
OAI21X1 g57044(.A0 (n_3439), .A1 (n_4318), .B0 (n_6479), .Y (n_4660));
OAI21X1 g55817(.A0 (n_3437), .A1 (n_4198), .B0 (n_7087), .Y (n_4659));
OAI21X1 g55819(.A0 (n_3436), .A1 (n_4274), .B0 (n_6479), .Y (n_4658));
NOR2X1 g58609(.A (n_5181), .B (n_4656), .Y (n_4657));
OR2X1 g58614(.A (n_4656), .B (n_5990), .Y (n_4655));
AOI21X1 g57783(.A0 (_2212_), .A1 (n_4468), .B0 (n_4653), .Y (n_4654));
OAI21X1 g57353(.A0 (n_3435), .A1 (n_4329), .B0 (n_4860), .Y (n_4652));
OAI21X1 g57518(.A0 (n_3864), .A1 (n_4240), .B0 (n_4947), .Y (n_4651));
OAI21X1 g57548(.A0 (n_3855), .A1 (n_4254), .B0 (n_5722), .Y (n_4650));
OAI21X1 g57562(.A0 (n_3648), .A1 (n_4133), .B0 (n_4860), .Y (n_4649));
OAI21X1 g57597(.A0 (n_4256), .A1 (n_7511), .B0 (n_4947), .Y (n_4648));
AOI21X1 g57611(.A0 (_2163_), .A1 (n_4644), .B0 (n_4646), .Y (n_4647));
AOI21X1 g57613(.A0 (_2239_), .A1 (n_4644), .B0 (n_4643), .Y (n_4645));
AOI21X1 g57614(.A0 (_2162_), .A1 (n_4644), .B0 (n_4641), .Y (n_4642));
AOI21X1 g57615(.A0 (_2238_), .A1 (n_4562), .B0 (n_4639), .Y (n_4640));
AOI21X1 g57616(.A0 (_2237_), .A1 (n_4628), .B0 (n_9418), .Y (n_4638));
AOI21X1 g57617(.A0 (_2161_), .A1 (n_4562), .B0 (n_4634), .Y (n_4636));
AOI21X1 g57618(.A0 (_2160_), .A1 (n_4644), .B0 (n_6632), .Y (n_4633));
AOI21X1 g57619(.A0 (_2159_), .A1 (n_4644), .B0 (n_4630), .Y (n_4631));
AOI21X1 g57620(.A0 (_2158_), .A1 (n_4628), .B0 (n_4627), .Y (n_4629));
AOI21X1 g57621(.A0 (_2323_), .A1 (n_4628), .B0 (n_4625), .Y (n_4626));
AOI21X1 g57622(.A0 (_2157_), .A1 (n_4628), .B0 (n_4623), .Y (n_4624));
AOI21X1 g57623(.A0 (_2156_), .A1 (n_4562), .B0 (n_9404), .Y (n_4622));
AOI21X1 g57625(.A0 (_2154_), .A1 (n_4615), .B0 (n_9410), .Y (n_4620));
AOI21X1 g57627(.A0 (_2299_), .A1 (n_4603), .B0 (n_4617), .Y (n_4618));
AOI21X1 g57629(.A0 (_2298_), .A1 (n_4615), .B0 (n_4614), .Y (n_4616));
AOI21X1 g57630(.A0 (_2297_), .A1 (n_4615), .B0 (n_6508), .Y (n_4613));
AOI21X1 g57633(.A0 (_2295_), .A1 (n_4615), .B0 (n_4610), .Y (n_4611));
AOI21X1 g57635(.A0 (_2294_), .A1 (n_4608), .B0 (n_4607), .Y (n_4609));
AOI21X1 g57636(.A0 (_2293_), .A1 (n_4600), .B0 (n_4605), .Y (n_4606));
AOI21X1 g57638(.A0 (_2292_), .A1 (n_4603), .B0 (n_4602), .Y (n_4604));
AOI21X1 g57640(.A0 (_2291_), .A1 (n_4600), .B0 (n_4599), .Y (n_4601));
AOI21X1 g57641(.A0 (_2290_), .A1 (n_4593), .B0 (n_4597), .Y (n_4598));
AOI21X1 g57642(.A0 (_2140_), .A1 (n_4586), .B0 (n_4595), .Y (n_4596));
AOI21X1 g57644(.A0 (_2289_), .A1 (n_4593), .B0 (n_4592), .Y (n_4594));
AOI21X1 g57645(.A0 (_2288_), .A1 (n_4593), .B0 (n_4590), .Y (n_4591));
AOI21X1 g57646(.A0 (_2287_), .A1 (n_4615), .B0 (n_4588), .Y (n_4589));
AOI21X1 g57647(.A0 (_2147_), .A1 (n_4586), .B0 (n_9412), .Y (n_4587));
AOI21X1 g57650(.A0 (_2285_), .A1 (n_4600), .B0 (n_4583), .Y (n_4584));
AOI21X1 g57651(.A0 (_2284_), .A1 (n_4579), .B0 (n_4581), .Y (n_4582));
AOI21X1 g57652(.A0 (_2145_), .A1 (n_4579), .B0 (n_4578), .Y (n_4580));
AOI21X1 g57653(.A0 (_2283_), .A1 (n_4579), .B0 (n_9408), .Y (n_4577));
AOI21X1 g57654(.A0 (_2282_), .A1 (n_4615), .B0 (n_4574), .Y (n_4575));
AOI21X1 g57657(.A0 (_2280_), .A1 (n_4600), .B0 (n_4572), .Y (n_4573));
AOI21X1 g57660(.A0 (_2143_), .A1 (n_4579), .B0 (n_4570), .Y (n_4571));
AOI21X1 g57663(.A0 (_2142_), .A1 (n_4579), .B0 (n_4568), .Y (n_4569));
AOI21X1 g57667(.A0 (_2141_), .A1 (n_4603), .B0 (n_4566), .Y (n_4567));
AOI21X1 g57669(.A0 (_2273_), .A1 (n_4562), .B0 (n_4564), .Y (n_4565));
AOI21X1 g57670(.A0 (_2272_), .A1 (n_4562), .B0 (n_9416), .Y (n_4563));
AOI21X1 g57672(.A0 (_2270_), .A1 (n_4586), .B0 (n_4559), .Y (n_4560));
AOI21X1 g57673(.A0 (_2137_), .A1 (n_4579), .B0 (n_4557), .Y (n_4558));
AOI21X1 g57675(.A0 (_2136_), .A1 (n_4579), .B0 (n_4555), .Y (n_4556));
AOI21X1 g57676(.A0 (_2135_), .A1 (n_4579), .B0 (n_4553), .Y (n_4554));
AOI21X1 g57678(.A0 (_2330_), .A1 (n_4562), .B0 (n_4551), .Y (n_4552));
AOI21X1 g57680(.A0 (_2328_), .A1 (n_4593), .B0 (n_4547), .Y (n_4548));
AOI21X1 g57681(.A0 (_2327_), .A1 (n_4593), .B0 (n_4545), .Y (n_4546));
AOI21X1 g57682(.A0 (_2326_), .A1 (n_4593), .B0 (n_4543), .Y (n_4544));
AOI21X1 g57683(.A0 (_2325_), .A1 (n_4593), .B0 (n_4541), .Y (n_4542));
AOI21X1 g57684(.A0 (_2204_), .A1 (n_4586), .B0 (n_4539), .Y (n_4540));
AOI21X1 g57685(.A0 (_2324_), .A1 (n_4562), .B0 (n_4537), .Y (n_4538));
AOI21X1 g57686(.A0 (_2322_), .A1 (n_4562), .B0 (n_4535), .Y (n_4536));
AOI21X1 g57687(.A0 (_2321_), .A1 (n_4608), .B0 (n_4533), .Y (n_4534));
AOI21X1 g57688(.A0 (_2320_), .A1 (n_4608), .B0 (n_4531), .Y (n_4532));
AOI21X1 g57689(.A0 (_2319_), .A1 (n_4600), .B0 (n_4529), .Y (n_4530));
AOI21X1 g57691(.A0 (_2203_), .A1 (n_4608), .B0 (n_4527), .Y (n_4528));
AOI21X1 g57692(.A0 (_2317_), .A1 (n_4608), .B0 (n_4525), .Y (n_4526));
AOI21X1 g57694(.A0 (_2315_), .A1 (n_4562), .B0 (n_4523), .Y (n_4524));
AOI21X1 g57696(.A0 (_2134_), .A1 (n_4608), .B0 (n_4521), .Y (n_4522));
AOI21X1 g57698(.A0 (_2202_), .A1 (n_4600), .B0 (n_4519), .Y (n_4520));
AOI21X1 g57699(.A0 (_2312_), .A1 (n_4600), .B0 (n_4517), .Y (n_4518));
AOI21X1 g57700(.A0 (_2311_), .A1 (n_4600), .B0 (n_4515), .Y (n_4516));
AOI21X1 g57701(.A0 (_2310_), .A1 (n_4562), .B0 (n_4513), .Y (n_4514));
AOI21X1 g57702(.A0 (_2309_), .A1 (n_4562), .B0 (n_6488), .Y (n_4512));
AOI21X1 g57703(.A0 (_2308_), .A1 (n_4608), .B0 (n_4509), .Y (n_4510));
AOI21X1 g57704(.A0 (_2201_), .A1 (n_4608), .B0 (n_4507), .Y (n_4508));
AOI21X1 g57705(.A0 (_2307_), .A1 (n_4608), .B0 (n_4505), .Y (n_4506));
AOI21X1 g57708(.A0 (_2304_), .A1 (n_4628), .B0 (n_4503), .Y (n_4504));
AOI21X1 g57711(.A0 (_2200_), .A1 (n_4644), .B0 (n_4501), .Y (n_4502));
CLKBUFX1 gbuf_d_531(.A(n_4084), .Y(d_out_531));
CLKBUFX1 gbuf_qn_531(.A(qn_in_531), .Y(WX4424));
AOI21X1 g57713(.A0 (_2199_), .A1 (n_4644), .B0 (n_4499), .Y (n_4500));
AOI21X1 g57714(.A0 (_2198_), .A1 (n_4562), .B0 (n_4497), .Y (n_4498));
AOI21X1 g57715(.A0 (_2133_), .A1 (n_4562), .B0 (n_4495), .Y (n_4496));
AOI21X1 g57716(.A0 (_2197_), .A1 (n_4628), .B0 (n_4493), .Y (n_4494));
AOI21X1 g57717(.A0 (_2196_), .A1 (n_4628), .B0 (n_4491), .Y (n_4492));
AOI21X1 g57718(.A0 (_2195_), .A1 (n_4644), .B0 (n_4489), .Y (n_4490));
AOI21X1 g57719(.A0 (_2132_), .A1 (n_4644), .B0 (n_4487), .Y (n_4488));
AOI21X1 g57720(.A0 (_2194_), .A1 (n_4562), .B0 (n_4485), .Y (n_4486));
AOI21X1 g57722(.A0 (_2192_), .A1 (n_4562), .B0 (n_4483), .Y (n_4484));
AOI21X1 g57723(.A0 (_2191_), .A1 (n_4644), .B0 (n_4481), .Y (n_4482));
AOI21X1 g57725(.A0 (_2190_), .A1 (n_4644), .B0 (n_4479), .Y (n_4480));
AOI21X1 g57726(.A0 (_2189_), .A1 (n_4644), .B0 (n_4477), .Y (n_4478));
AOI21X1 g57727(.A0 (_2188_), .A1 (n_4562), .B0 (n_9420), .Y (n_4476));
AOI21X1 g57732(.A0 (_2129_), .A1 (n_4471), .B0 (n_4473), .Y (n_4474));
AOI21X1 g57733(.A0 (_2184_), .A1 (n_4471), .B0 (n_9426), .Y (n_4472));
AOI21X1 g57735(.A0 (_2182_), .A1 (n_4468), .B0 (n_4467), .Y (n_4469));
AOI21X1 g57736(.A0 (_2181_), .A1 (n_4562), .B0 (n_4465), .Y (n_4466));
AOI21X1 g57737(.A0 (_2128_), .A1 (n_4603), .B0 (n_4463), .Y (n_4464));
AOI21X1 g57738(.A0 (_2180_), .A1 (n_4603), .B0 (n_4461), .Y (n_4462));
AOI21X1 g57744(.A0 (_2126_), .A1 (n_4468), .B0 (n_4459), .Y (n_4460));
AOI21X1 g57745(.A0 (_2175_), .A1 (n_4593), .B0 (n_4457), .Y (n_4458));
AOI21X1 g57746(.A0 (_2174_), .A1 (n_4593), .B0 (n_4455), .Y (n_4456));
AOI21X1 g57747(.A0 (_2173_), .A1 (n_4471), .B0 (n_10722), .Y(n_4454));
AOI21X1 g57748(.A0 (_2125_), .A1 (n_4471), .B0 (n_4451), .Y (n_4452));
AOI21X1 g57750(.A0 (_2123_), .A1 (n_4471), .B0 (n_4449), .Y (n_4450));
AOI21X1 g57751(.A0 (_2122_), .A1 (n_4586), .B0 (n_4447), .Y (n_4448));
AOI21X1 g57752(.A0 (_2236_), .A1 (n_4586), .B0 (n_6885), .Y (n_4446));
AOI21X1 g57753(.A0 (_2235_), .A1 (n_4586), .B0 (n_6451), .Y (n_4444));
AOI21X1 g57755(.A0 (_2234_), .A1 (n_4439), .B0 (n_4441), .Y (n_4442));
AOI21X1 g57756(.A0 (_2233_), .A1 (n_4439), .B0 (n_4438), .Y (n_4440));
AOI21X1 g57757(.A0 (_2232_), .A1 (n_4439), .B0 (n_4436), .Y (n_4437));
AOI21X1 g57759(.A0 (_2231_), .A1 (n_4586), .B0 (n_4434), .Y (n_4435));
AOI21X1 g57760(.A0 (_2230_), .A1 (n_4586), .B0 (n_4432), .Y (n_4433));
AOI21X1 g57761(.A0 (_2229_), .A1 (n_4586), .B0 (n_4430), .Y (n_4431));
AOI21X1 g57762(.A0 (_2228_), .A1 (n_4586), .B0 (n_4428), .Y (n_4429));
AOI21X1 g57763(.A0 (_2227_), .A1 (n_4603), .B0 (n_4426), .Y (n_4427));
AOI21X1 g57764(.A0 (_2119_), .A1 (n_4603), .B0 (n_4424), .Y (n_4425));
AOI21X1 g57765(.A0 (_2226_), .A1 (n_4586), .B0 (n_4422), .Y (n_4423));
AOI21X1 g57766(.A0 (_2225_), .A1 (n_4586), .B0 (n_4420), .Y (n_4421));
OAI21X1 g56810(.A0 (n_3642), .A1 (n_4124), .B0 (n_4860), .Y (n_4419));
AOI21X1 g57767(.A0 (_2118_), .A1 (n_4562), .B0 (n_4417), .Y (n_4418));
AOI21X1 g57768(.A0 (_2224_), .A1 (n_4562), .B0 (n_4415), .Y (n_4416));
AOI21X1 g57769(.A0 (_2223_), .A1 (n_4603), .B0 (n_4413), .Y (n_4414));
AOI21X1 g57770(.A0 (_2222_), .A1 (n_4439), .B0 (n_4411), .Y (n_4412));
AOI21X1 g57771(.A0 (_2221_), .A1 (n_4603), .B0 (n_4409), .Y (n_4410));
AOI21X1 g57772(.A0 (_2220_), .A1 (n_4439), .B0 (n_9422), .Y (n_4408));
AOI21X1 g57774(.A0 (_2219_), .A1 (n_4468), .B0 (n_4405), .Y (n_4406));
AOI21X1 g57775(.A0 (_2218_), .A1 (n_4471), .B0 (n_4403), .Y (n_4404));
AOI21X1 g57777(.A0 (_2217_), .A1 (n_4439), .B0 (n_4401), .Y (n_4402));
AOI21X1 g57778(.A0 (_2216_), .A1 (n_4439), .B0 (n_4399), .Y (n_4400));
AOI21X1 g57781(.A0 (_2115_), .A1 (n_4439), .B0 (n_9414), .Y (n_4398));
AOI21X1 g57782(.A0 (_2213_), .A1 (n_4562), .B0 (n_4395), .Y (n_4396));
AOI21X1 g57788(.A0 (_2113_), .A1 (n_4468), .B0 (n_10714), .Y(n_4394));
AOI21X1 g57789(.A0 (_2208_), .A1 (n_4468), .B0 (n_10718), .Y(n_4392));
AOI21X1 g57792(.A0 (_2205_), .A1 (n_4600), .B0 (n_4389), .Y (n_4390));
OAI21X1 g56827(.A0 (n_3443), .A1 (n_4294), .B0 (n_4860), .Y (n_4388));
AOI21X1 g57800(.A0 (_2109_), .A1 (n_4471), .B0 (n_4386), .Y (n_4387));
AOI21X1 g57828(.A0 (_2268_), .A1 (n_4586), .B0 (n_4384), .Y (n_4385));
AOI21X1 g57829(.A0 (_2267_), .A1 (n_4603), .B0 (n_4382), .Y (n_4383));
AOI21X1 g57830(.A0 (_2266_), .A1 (n_4471), .B0 (n_4380), .Y (n_4381));
AOI21X1 g57831(.A0 (_2265_), .A1 (n_4468), .B0 (n_4378), .Y (n_4379));
AOI21X1 g57832(.A0 (_2264_), .A1 (n_4603), .B0 (n_4376), .Y (n_4377));
AOI21X1 g57833(.A0 (_2263_), .A1 (n_4468), .B0 (n_4374), .Y (n_4375));
AOI21X1 g57837(.A0 (_2259_), .A1 (n_4603), .B0 (n_4372), .Y (n_4373));
AOI21X1 g57839(.A0 (_2258_), .A1 (n_4644), .B0 (n_4370), .Y (n_4371));
AOI21X1 g57840(.A0 (_2257_), .A1 (n_4628), .B0 (n_4368), .Y (n_4369));
AOI21X1 g57841(.A0 (_2171_), .A1 (n_4628), .B0 (n_4366), .Y (n_4367));
AOI21X1 g57842(.A0 (_2256_), .A1 (n_4628), .B0 (n_4364), .Y (n_4365));
AOI21X1 g57843(.A0 (_2255_), .A1 (n_4562), .B0 (n_4362), .Y (n_4363));
AOI21X1 g57844(.A0 (_2254_), .A1 (n_4628), .B0 (n_4360), .Y (n_4361));
AOI21X1 g57845(.A0 (_2170_), .A1 (n_4593), .B0 (n_4358), .Y (n_4359));
AOI21X1 g57846(.A0 (_2253_), .A1 (n_4593), .B0 (n_4356), .Y (n_4357));
AOI21X1 g57847(.A0 (_2169_), .A1 (n_4579), .B0 (n_4354), .Y (n_4355));
AOI21X1 g57849(.A0 (_2251_), .A1 (n_4593), .B0 (n_9406), .Y (n_4353));
AOI21X1 g57850(.A0 (_2168_), .A1 (n_4615), .B0 (n_4350), .Y (n_4351));
AOI21X1 g57852(.A0 (_2249_), .A1 (n_4615), .B0 (n_4348), .Y (n_4349));
AOI21X1 g57853(.A0 (_2167_), .A1 (n_4615), .B0 (n_4346), .Y (n_4347));
AOI21X1 g57855(.A0 (_2247_), .A1 (n_4468), .B0 (n_9428), .Y (n_4345));
AOI21X1 g57856(.A0 (_2166_), .A1 (n_4468), .B0 (n_4342), .Y (n_4343));
AOI21X1 g57858(.A0 (_2245_), .A1 (n_4468), .B0 (n_4340), .Y (n_4341));
AOI21X1 g57859(.A0 (_2165_), .A1 (n_4628), .B0 (n_4338), .Y (n_4339));
AOI21X1 g57862(.A0 (_2164_), .A1 (n_4628), .B0 (n_4336), .Y (n_4337));
NOR2X1 g56923(.A (WX8303), .B (n_5479), .Y (n_4335));
MX2X1 g55844(.A (n_2888), .B (WX487), .S0 (n_10747), .Y (n_4334));
NOR2X1 g56984(.A (WX9596), .B (n_1425), .Y (n_4333));
NOR2X1 g56987(.A (WX9596), .B (n_5479), .Y (n_4332));
OAI21X1 g57352(.A0 (n_3431), .A1 (n_4087), .B0 (n_4860), .Y (n_4331));
AOI21X1 g57394(.A0 (_2108_), .A1 (n_4184), .B0 (n_4329), .Y (n_4330));
MX2X1 g57401(.A (n_3599), .B (WX485), .S0 (n_9433), .Y (n_4328));
NOR2X1 g56688(.A (WX3131), .B (n_4670), .Y (n_4327));
AOI21X1 g57610(.A0 (_2241_), .A1 (n_4644), .B0 (n_4325), .Y (n_4326));
AOI21X1 g57612(.A0 (_2240_), .A1 (n_4644), .B0 (n_4323), .Y (n_4324));
AOI21X1 g57624(.A0 (_2155_), .A1 (n_4615), .B0 (n_11605), .Y(n_4322));
NOR2X1 g56709(.A (WX3131), .B (n_3690), .Y (n_4320));
AOI21X1 g57626(.A0 (_2300_), .A1 (n_4562), .B0 (n_4318), .Y (n_4319));
AOI21X1 g57628(.A0 (_2153_), .A1 (n_4615), .B0 (n_4316), .Y (n_4317));
AOI21X1 g57631(.A0 (_2152_), .A1 (n_4603), .B0 (n_4314), .Y (n_4315));
AOI21X1 g57632(.A0 (_2296_), .A1 (n_4615), .B0 (n_4312), .Y (n_4313));
AOI21X1 g57634(.A0 (_2151_), .A1 (n_4615), .B0 (n_4310), .Y (n_4311));
AOI21X1 g57637(.A0 (_2150_), .A1 (n_4600), .B0 (n_4308), .Y (n_4309));
AOI21X1 g57639(.A0 (_2149_), .A1 (n_4600), .B0 (n_11619), .Y(n_4307));
AOI21X1 g57643(.A0 (_2148_), .A1 (n_4593), .B0 (n_4304), .Y (n_4305));
AOI21X1 g57648(.A0 (_2286_), .A1 (n_4615), .B0 (n_4302), .Y (n_4303));
AOI21X1 g57649(.A0 (_2146_), .A1 (n_4600), .B0 (n_11623), .Y(n_4301));
AOI21X1 g57655(.A0 (_2281_), .A1 (n_4615), .B0 (n_4298), .Y (n_4299));
AOI21X1 g57656(.A0 (_2144_), .A1 (n_4600), .B0 (n_11597), .Y(n_4297));
AOI21X1 g57658(.A0 (_2139_), .A1 (n_4579), .B0 (n_4294), .Y (n_4295));
AOI21X1 g57659(.A0 (_2279_), .A1 (n_4579), .B0 (n_4292), .Y (n_4293));
AOI21X1 g57661(.A0 (_2278_), .A1 (n_4579), .B0 (n_4290), .Y (n_4291));
AOI21X1 g57662(.A0 (_2277_), .A1 (n_4579), .B0 (n_4288), .Y (n_4289));
AOI21X1 g57664(.A0 (_2276_), .A1 (n_4579), .B0 (n_4286), .Y (n_4287));
AOI21X1 g57665(.A0 (_2275_), .A1 (n_4579), .B0 (n_11596), .Y(n_4285));
AOI21X1 g57666(.A0 (_2138_), .A1 (n_4603), .B0 (n_4282), .Y (n_4283));
AOI21X1 g57668(.A0 (_2274_), .A1 (n_4603), .B0 (n_4280), .Y (n_4281));
AOI21X1 g57671(.A0 (_2271_), .A1 (n_4586), .B0 (n_11601), .Y(n_4279));
AOI21X1 g57674(.A0 (_2269_), .A1 (n_4579), .B0 (n_4276), .Y (n_4277));
AOI21X1 g57677(.A0 (_2331_), .A1 (n_4562), .B0 (n_4274), .Y (n_4275));
AOI21X1 g57690(.A0 (_2318_), .A1 (n_4600), .B0 (n_4272), .Y (n_4273));
AOI21X1 g57693(.A0 (_2316_), .A1 (n_4562), .B0 (n_7084), .Y (n_4271));
AOI21X1 g57695(.A0 (_2314_), .A1 (n_4608), .B0 (n_6469), .Y (n_4269));
AOI21X1 g57697(.A0 (_2313_), .A1 (n_4600), .B0 (n_4266), .Y (n_4267));
AOI21X1 g57706(.A0 (_2306_), .A1 (n_4608), .B0 (n_4264), .Y (n_4265));
AOI21X1 g57707(.A0 (_2305_), .A1 (n_4628), .B0 (n_4262), .Y (n_4263));
AOI21X1 g57709(.A0 (_2303_), .A1 (n_4562), .B0 (n_4260), .Y (n_4261));
AOI21X1 g57710(.A0 (_2302_), .A1 (n_4562), .B0 (n_4258), .Y (n_4259));
AOI21X1 g57712(.A0 (_2301_), .A1 (n_4593), .B0 (n_4256), .Y (n_4257));
AOI21X1 g57721(.A0 (_2193_), .A1 (n_4562), .B0 (n_4254), .Y (n_4255));
AOI21X1 g57724(.A0 (_2131_), .A1 (n_4644), .B0 (n_4252), .Y (n_4253));
AOI21X1 g57728(.A0 (_2130_), .A1 (n_4562), .B0 (n_4250), .Y (n_4251));
AOI21X1 g57729(.A0 (_2187_), .A1 (n_4468), .B0 (n_4248), .Y (n_4249));
AOI21X1 g57730(.A0 (_2186_), .A1 (n_4608), .B0 (n_11607), .Y(n_4247));
AOI21X1 g57731(.A0 (_2185_), .A1 (n_4608), .B0 (n_4244), .Y (n_4245));
AOI21X1 g57734(.A0 (_2183_), .A1 (n_4468), .B0 (n_11615), .Y(n_4243));
AOI21X1 g57739(.A0 (_2127_), .A1 (n_4471), .B0 (n_4240), .Y (n_4241));
AOI21X1 g57740(.A0 (_2179_), .A1 (n_4471), .B0 (n_4238), .Y (n_4239));
AOI21X1 g57741(.A0 (_2178_), .A1 (n_4439), .B0 (n_4236), .Y (n_4237));
AOI21X1 g57742(.A0 (_2177_), .A1 (n_4439), .B0 (n_10716), .Y(n_4235));
AOI21X1 g57743(.A0 (_2176_), .A1 (n_4593), .B0 (n_4232), .Y (n_4233));
AOI21X1 g57749(.A0 (_2124_), .A1 (n_4471), .B0 (n_4230), .Y (n_4231));
AOI21X1 g57754(.A0 (_2121_), .A1 (n_4439), .B0 (n_4228), .Y (n_4229));
AOI21X1 g57758(.A0 (_2120_), .A1 (n_4439), .B0 (n_11611), .Y(n_4227));
AOI21X1 g57773(.A0 (_2117_), .A1 (n_4439), .B0 (n_4224), .Y (n_4225));
AOI21X1 g57776(.A0 (_2116_), .A1 (n_4439), .B0 (n_4222), .Y (n_4223));
NOR2X1 g56817(.A (WX5717), .B (n_2620), .Y (n_4221));
AOI21X1 g57779(.A0 (_2215_), .A1 (n_4439), .B0 (n_4219), .Y (n_4220));
AOI21X1 g57780(.A0 (_2214_), .A1 (n_4439), .B0 (n_11617), .Y(n_4218));
NOR2X1 g56820(.A (WX5717), .B (n_5052), .Y (n_6684));
AOI21X1 g57784(.A0 (_2211_), .A1 (n_4468), .B0 (n_11621), .Y(n_4215));
AOI21X1 g57786(.A0 (_2114_), .A1 (n_4468), .B0 (n_11625), .Y(n_4213));
AOI21X1 g57787(.A0 (_2209_), .A1 (n_4608), .B0 (n_4210), .Y (n_4211));
AOI21X1 g57790(.A0 (_2207_), .A1 (n_4562), .B0 (n_4208), .Y (n_4209));
AOI21X1 g57791(.A0 (_2206_), .A1 (n_4600), .B0 (n_11603), .Y(n_4207));
AOI21X1 g57793(.A0 (_2112_), .A1 (n_4471), .B0 (n_4204), .Y (n_4205));
AOI21X1 g57794(.A0 (_2111_), .A1 (n_4471), .B0 (n_11599), .Y(n_4203));
AOI21X1 g57795(.A0 (_2110_), .A1 (n_4471), .B0 (n_10720), .Y(n_4201));
AOI21X1 g57796(.A0 (_2107_), .A1 (n_3831), .B0 (n_4198), .Y (n_4199));
AOI21X1 g57797(.A0 (_2106_), .A1 (n_3831), .B0 (n_4195), .Y (n_4197));
AOI21X1 g57798(.A0 (_2105_), .A1 (n_3831), .B0 (n_4193), .Y (n_4194));
AOI21X1 g57799(.A0 (_2104_), .A1 (n_5828), .B0 (n_4191), .Y (n_4192));
AOI21X1 g57801(.A0 (_2103_), .A1 (n_5828), .B0 (n_4188), .Y (n_4190));
AOI21X1 g57802(.A0 (_2102_), .A1 (n_3831), .B0 (n_4186), .Y (n_4187));
AOI21X1 g57803(.A0 (_2101_), .A1 (n_4184), .B0 (n_4183), .Y (n_4185));
AOI21X1 g57804(.A0 (_2100_), .A1 (n_5828), .B0 (n_4181), .Y (n_4182));
AOI21X1 g57805(.A0 (_2099_), .A1 (n_4184), .B0 (n_4179), .Y (n_4180));
MX2X1 g55904(.A (n_3685), .B (WX489), .S0 (n_7082), .Y (n_4178));
AOI21X1 g57806(.A0 (_2098_), .A1 (n_4184), .B0 (n_4176), .Y (n_4177));
AOI21X1 g57807(.A0 (_2097_), .A1 (n_4150), .B0 (n_4174), .Y (n_4175));
AOI21X1 g57808(.A0 (_2096_), .A1 (n_4184), .B0 (n_4172), .Y (n_4173));
AOI21X1 g57809(.A0 (_2095_), .A1 (n_4184), .B0 (n_4170), .Y (n_4171));
AOI21X1 g57810(.A0 (_2094_), .A1 (n_5828), .B0 (n_4168), .Y (n_4169));
AOI21X1 g57811(.A0 (_2093_), .A1 (n_4184), .B0 (n_4166), .Y (n_4167));
AOI21X1 g57812(.A0 (_2092_), .A1 (n_5828), .B0 (n_4164), .Y (n_4165));
AOI21X1 g57813(.A0 (_2091_), .A1 (n_5828), .B0 (n_4162), .Y (n_4163));
AOI21X1 g57814(.A0 (_2090_), .A1 (n_4184), .B0 (n_4160), .Y (n_4161));
AOI21X1 g57815(.A0 (_2089_), .A1 (n_5828), .B0 (n_4158), .Y (n_4159));
AOI21X1 g57816(.A0 (_2088_), .A1 (n_4184), .B0 (n_4156), .Y (n_4157));
AOI21X1 g57817(.A0 (_2087_), .A1 (n_4184), .B0 (n_4154), .Y (n_4155));
AOI21X1 g57818(.A0 (_2086_), .A1 (n_5828), .B0 (n_4152), .Y (n_4153));
AOI21X1 g57819(.A0 (_2085_), .A1 (n_4150), .B0 (n_4149), .Y (n_4151));
AOI21X1 g57820(.A0 (_2084_), .A1 (n_5828), .B0 (n_4147), .Y (n_4148));
AOI21X1 g57821(.A0 (_2083_), .A1 (n_3831), .B0 (n_4145), .Y (n_4146));
AOI21X1 g57822(.A0 (_2082_), .A1 (n_5828), .B0 (n_4143), .Y (n_4144));
AOI21X1 g57823(.A0 (_2081_), .A1 (n_5828), .B0 (n_4141), .Y (n_4142));
AOI21X1 g57824(.A0 (_2080_), .A1 (n_4184), .B0 (n_4139), .Y (n_4140));
AOI21X1 g57825(.A0 (_2079_), .A1 (n_4184), .B0 (n_4137), .Y (n_4138));
AOI21X1 g57826(.A0 (_2078_), .A1 (n_4150), .B0 (n_4135), .Y (n_4136));
AOI21X1 g57827(.A0 (_2077_), .A1 (n_5828), .B0 (n_4133), .Y (n_4134));
AOI21X1 g57834(.A0 (_2262_), .A1 (n_4608), .B0 (n_4131), .Y (n_4132));
AOI21X1 g57835(.A0 (_2261_), .A1 (n_4471), .B0 (n_4129), .Y (n_4130));
AOI21X1 g57836(.A0 (_2260_), .A1 (n_4471), .B0 (n_4127), .Y (n_4128));
NOR2X1 g56860(.A (WX7010), .B (n_5479), .Y (n_4126));
AOI21X1 g57838(.A0 (_2172_), .A1 (n_4562), .B0 (n_4124), .Y (n_4125));
AOI21X1 g57848(.A0 (_2252_), .A1 (n_4593), .B0 (n_4122), .Y (n_4123));
AOI21X1 g57851(.A0 (_2250_), .A1 (n_4603), .B0 (n_11609), .Y(n_4121));
AOI21X1 g57854(.A0 (_2248_), .A1 (n_4615), .B0 (n_11613), .Y(n_4119));
AOI21X1 g57857(.A0 (_2246_), .A1 (n_4468), .B0 (n_4116), .Y (n_4117));
AOI21X1 g57860(.A0 (_2244_), .A1 (n_4628), .B0 (n_4114), .Y (n_4115));
AOI21X1 g57861(.A0 (_2243_), .A1 (n_4628), .B0 (n_4112), .Y (n_4113));
AOI21X1 g57863(.A0 (_2242_), .A1 (n_4562), .B0 (n_10712), .Y(n_4111));
MX2X1 g57869(.A (n_3695), .B (WX547), .S0 (n_9437), .Y (n_4109));
NOR2X1 g56883(.A (WX7010), .B (n_2851), .Y (n_4108));
NOR2X1 g56920(.A (WX8303), .B (n_1648), .Y (n_4107));
AND2X1 g57963(.A (n_3980), .B (n_4106), .Y (n_4566));
AND2X1 g57965(.A (n_3979), .B (n_4106), .Y (n_4564));
AND2X1 g57969(.A (n_3977), .B (n_4105), .Y (n_4559));
AND2X1 g57970(.A (n_3976), .B (n_4105), .Y (n_4557));
AND2X1 g57972(.A (n_3975), .B (n_4101), .Y (n_4551));
AND2X1 g57975(.A (n_3974), .B (n_4103), .Y (n_4549));
AND2X1 g57976(.A (n_3973), .B (n_4104), .Y (n_4555));
AND2X1 g57977(.A (n_3972), .B (n_4105), .Y (n_4553));
AND2X1 g57978(.A (n_3971), .B (n_4106), .Y (n_4539));
AND2X1 g57980(.A (n_3970), .B (n_4104), .Y (n_4547));
AND2X1 g57981(.A (n_3969), .B (n_4105), .Y (n_4527));
AND2X1 g57982(.A (n_3968), .B (n_4106), .Y (n_4521));
AND2X1 g57983(.A (n_3967), .B (n_4103), .Y (n_4519));
AND2X1 g57984(.A (n_3966), .B (n_4096), .Y (n_4507));
AND2X1 g57986(.A (n_3965), .B (n_4104), .Y (n_4501));
AND2X1 g57987(.A (n_3964), .B (n_4104), .Y (n_4545));
AND2X1 g57988(.A (n_3963), .B (n_4104), .Y (n_4499));
AND2X1 g57990(.A (n_3962), .B (n_4106), .Y (n_4497));
AND2X1 g57991(.A (n_3961), .B (n_4100), .Y (n_4495));
AND2X1 g57992(.A (n_3960), .B (n_4103), .Y (n_4493));
AND2X1 g57993(.A (n_3959), .B (n_4096), .Y (n_4491));
AND2X1 g57995(.A (n_3957), .B (n_6452), .Y (n_4543));
AND2X1 g57996(.A (n_3958), .B (n_4101), .Y (n_4489));
AND2X1 g57997(.A (n_3956), .B (n_4101), .Y (n_4487));
AND2X1 g57998(.A (n_3955), .B (n_4100), .Y (n_4485));
AND2X1 g58001(.A (n_3954), .B (n_6633), .Y (n_4483));
AND2X1 g58002(.A (n_3953), .B (n_4099), .Y (n_4541));
AND2X1 g58003(.A (n_3952), .B (n_4099), .Y (n_4481));
AND2X1 g58005(.A (n_3951), .B (n_4096), .Y (n_4479));
AND2X1 g58007(.A (n_4099), .B (n_7281), .Y (n_4477));
AND2X1 g58011(.A (n_3948), .B (n_6452), .Y (n_4537));
AND2X1 g58015(.A (n_3947), .B (n_4101), .Y (n_4473));
AND2X1 g58018(.A (n_3945), .B (n_4099), .Y (n_4625));
AND2X1 g58020(.A (n_3944), .B (n_6452), .Y (n_4467));
AND2X1 g58021(.A (n_3943), .B (n_4099), .Y (n_4465));
AND2X1 g58022(.A (n_3942), .B (n_4106), .Y (n_4463));
AND2X1 g58023(.A (n_3941), .B (n_4104), .Y (n_4461));
AND2X1 g58027(.A (n_3940), .B (n_4106), .Y (n_4535));
AND2X1 g58031(.A (n_3939), .B (n_6633), .Y (n_4459));
AND2X1 g58032(.A (n_3938), .B (n_6452), .Y (n_4457));
AND2X1 g58033(.A (n_3937), .B (n_4099), .Y (n_4533));
AND2X1 g58035(.A (n_3936), .B (n_4096), .Y (n_4455));
AND2X1 g58038(.A (n_3934), .B (n_4106), .Y (n_4451));
AND2X1 g58039(.A (n_3933), .B (n_4095), .Y (n_4531));
AND2X1 g58042(.A (n_3932), .B (n_4099), .Y (n_4529));
AND2X1 g58044(.A (n_4103), .B (n_8340), .Y (n_4449));
AND2X1 g58047(.A (n_3930), .B (n_6452), .Y (n_4447));
AND2X1 g58051(.A (n_3927), .B (n_4100), .Y (n_4441));
AND2X1 g58052(.A (n_3926), .B (n_4100), .Y (n_4438));
AND2X1 g58053(.A (n_3925), .B (n_4096), .Y (n_4525));
AND2X1 g58055(.A (n_3924), .B (n_4100), .Y (n_4436));
AND2X1 g58057(.A (n_3923), .B (n_4096), .Y (n_4434));
AND2X1 g58058(.A (n_3922), .B (n_4100), .Y (n_4432));
AND2X1 g58060(.A (n_3921), .B (n_4100), .Y (n_4430));
AND2X1 g58062(.A (n_3920), .B (n_4096), .Y (n_4428));
AND2X1 g58064(.A (n_3919), .B (n_6452), .Y (n_4426));
AND2X1 g58065(.A (n_6633), .B (n_8346), .Y (n_4424));
AND2X1 g58066(.A (n_3917), .B (n_4105), .Y (n_4422));
AND2X1 g58067(.A (n_3916), .B (n_6633), .Y (n_4420));
AND2X1 g58068(.A (n_3915), .B (n_4105), .Y (n_4523));
AND2X1 g58069(.A (n_3913), .B (n_4095), .Y (n_4417));
AND2X1 g58070(.A (n_3914), .B (n_4099), .Y (n_4415));
AND2X1 g58072(.A (n_3912), .B (n_4095), .Y (n_4413));
AND2X1 g58073(.A (n_3911), .B (n_4104), .Y (n_4411));
AND2X1 g58075(.A (n_3910), .B (n_6633), .Y (n_4409));
AND2X1 g58079(.A (n_3908), .B (n_4104), .Y (n_4405));
AND2X1 g58080(.A (n_4095), .B (n_8341), .Y (n_4403));
AND2X1 g58082(.A (n_3906), .B (n_4095), .Y (n_4401));
AND2X1 g58085(.A (n_4100), .B (n_8344), .Y (n_4399));
AND2X1 g58089(.A (n_3903), .B (n_6452), .Y (n_4395));
AND2X1 g58091(.A (n_3901), .B (n_4100), .Y (n_4517));
AND2X1 g58092(.A (n_6633), .B (n_8349), .Y (n_4653));
AND2X1 g58095(.A (n_3900), .B (n_4101), .Y (n_4661));
AND2X1 g58098(.A (n_3898), .B (n_4017), .Y (n_4515));
AND2X1 g58104(.A (n_4105), .B (n_9403), .Y (n_4389));
AND2X1 g58106(.A (n_3895), .B (n_6633), .Y (n_4513));
AND2X1 g58113(.A (n_3893), .B (n_4104), .Y (n_4509));
AND2X1 g58114(.A (n_3892), .B (n_4104), .Y (n_4386));
AND2X1 g58116(.A (n_3891), .B (n_4101), .Y (n_4505));
AND2X1 g58119(.A (n_3890), .B (n_6633), .Y (n_4384));
AND2X1 g58120(.A (n_3889), .B (n_4103), .Y (n_4382));
AND2X1 g58121(.A (n_3888), .B (n_4094), .Y (n_4380));
AND2X1 g58122(.A (n_3887), .B (n_4094), .Y (n_4503));
AND2X1 g58123(.A (n_3886), .B (n_6452), .Y (n_4378));
AND2X1 g58124(.A (n_3885), .B (n_4096), .Y (n_4376));
AND2X1 g58125(.A (n_3884), .B (n_6633), .Y (n_4374));
AND2X1 g58130(.A (n_3883), .B (n_4096), .Y (n_4372));
AND2X1 g58132(.A (n_3882), .B (n_4095), .Y (n_4370));
AND2X1 g58134(.A (n_3881), .B (n_4096), .Y (n_4368));
AND2X1 g58135(.A (n_3880), .B (n_4096), .Y (n_4366));
AND2X1 g58136(.A (n_3879), .B (n_4095), .Y (n_4364));
AND2X1 g58137(.A (n_3878), .B (n_4095), .Y (n_4362));
AND2X1 g58138(.A (n_3877), .B (n_4095), .Y (n_4360));
AND2X1 g58139(.A (n_3876), .B (n_4096), .Y (n_4358));
AND2X1 g58140(.A (n_3875), .B (n_4096), .Y (n_4356));
AND2X1 g58142(.A (n_3874), .B (n_6452), .Y (n_4354));
AND2X1 g58145(.A (n_3872), .B (n_4094), .Y (n_4350));
AND2X1 g58147(.A (n_3871), .B (n_4094), .Y (n_4348));
AND2X1 g58149(.A (n_3870), .B (n_6452), .Y (n_4346));
AND2X1 g58151(.A (n_3868), .B (n_4096), .Y (n_4342));
AND2X1 g58153(.A (n_4101), .B (n_8347), .Y (n_4340));
AND2X1 g58154(.A (n_4096), .B (n_7282), .Y (n_4338));
AND2X1 g58157(.A (n_3865), .B (n_6633), .Y (n_4336));
CLKBUFX1 gbuf_d_532(.A(n_3863), .Y(d_out_532));
CLKBUFX1 gbuf_qn_532(.A(qn_in_532), .Y(WX8259));
CLKBUFX1 gbuf_d_533(.A(n_3860), .Y(d_out_533));
CLKBUFX1 gbuf_qn_533(.A(qn_in_533), .Y(WX9550));
CLKBUFX1 gbuf_d_534(.A(n_3859), .Y(d_out_534));
CLKBUFX1 gbuf_qn_534(.A(qn_in_534), .Y(WX4386));
CLKBUFX1 gbuf_d_535(.A(n_3856), .Y(d_out_535));
CLKBUFX1 gbuf_qn_535(.A(qn_in_535), .Y(WX5677));
CLKBUFX1 gbuf_d_536(.A(n_3854), .Y(d_out_536));
CLKBUFX1 gbuf_qn_536(.A(qn_in_536), .Y(WX6968));
CLKBUFX1 gbuf_d_537(.A(n_3853), .Y(d_out_537));
CLKBUFX1 gbuf_qn_537(.A(qn_in_537), .Y(WX3095));
NOR2X1 g58604(.A (WX1838), .B (n_2620), .Y (n_4093));
NOR2X1 g58605(.A (WX10889), .B (n_1425), .Y (n_4092));
NOR2X1 g58612(.A (WX1838), .B (n_5479), .Y (n_4090));
NOR2X1 g58618(.A (WX10889), .B (n_5662), .Y (n_7510));
INVX1 g58812(.A (WX545), .Y (n_4656));
AOI21X1 g57389(.A0 (_2332_), .A1 (n_4562), .B0 (n_4087), .Y (n_4088));
NAND2X1 g57449(.A (n_9433), .B (n_4015), .Y (n_4086));
NOR2X1 g56809(.A (WX4426), .B (n_1425), .Y (n_4084));
NOR2X1 g56813(.A (WX4426), .B (n_5479), .Y (n_4083));
NAND2X1 g57874(.A (n_6645), .B (n_4078), .Y (n_4082));
NAND2X1 g57875(.A (n_4079), .B (n_4078), .Y (n_4080));
NAND2X1 g57876(.A (n_4076), .B (n_4078), .Y (n_4077));
NAND2X1 g57877(.A (n_10731), .B (n_4015), .Y (n_4075));
NAND2X1 g57878(.A (n_4071), .B (n_4078), .Y (n_4072));
NAND2X1 g57879(.A (n_4069), .B (n_4078), .Y (n_4070));
NAND2X1 g57880(.A (n_6601), .B (n_4078), .Y (n_4068));
NAND2X1 g57881(.A (n_10743), .B (n_4058), .Y (n_4066));
NAND2X1 g57882(.A (n_7074), .B (n_4078), .Y (n_4064));
NAND2X1 g57883(.A (n_4061), .B (n_4078), .Y (n_4062));
NAND2X1 g57884(.A (n_6613), .B (n_4058), .Y (n_4060));
NAND2X1 g57885(.A (n_9800), .B (n_4058), .Y (n_4057));
NAND2X1 g57886(.A (n_10727), .B (n_4015), .Y (n_4055));
NAND2X1 g57887(.A (n_4052), .B (n_4078), .Y (n_4053));
NAND2X1 g57888(.A (n_4050), .B (n_4078), .Y (n_4051));
NAND2X1 g57889(.A (n_7078), .B (n_4015), .Y (n_4049));
NAND2X1 g57890(.A (n_9437), .B (n_4015), .Y (n_4047));
NAND2X1 g57891(.A (n_4044), .B (n_3173), .Y (n_4045));
NAND2X1 g57892(.A (n_7062), .B (n_4078), .Y (n_4043));
NAND2X1 g57893(.A (n_4040), .B (n_4015), .Y (n_4041));
NAND2X1 g57894(.A (n_4038), .B (n_4078), .Y (n_4039));
NAND2X1 g57895(.A (n_7082), .B (n_4078), .Y (n_4037));
NAND2X1 g57896(.A (n_6573), .B (n_4058), .Y (n_4035));
NAND2X1 g57897(.A (n_7070), .B (n_4078), .Y (n_4033));
NAND2X1 g57898(.A (n_10747), .B (n_4015), .Y (n_4031));
NAND2X1 g57899(.A (n_10735), .B (n_4058), .Y (n_4029));
NAND2X1 g57900(.A (n_4026), .B (n_4058), .Y (n_4027));
NAND2X1 g57901(.A (n_6553), .B (n_4058), .Y (n_4025));
NAND2X1 g57902(.A (n_7066), .B (n_4078), .Y (n_4023));
NAND2X1 g57903(.A (n_10739), .B (n_4078), .Y (n_4021));
NAND2X1 g57904(.A (n_4018), .B (n_4058), .Y (n_4019));
AND2X1 g57906(.A (n_4014), .B (n_4094), .Y (n_4646));
AND2X1 g57908(.A (n_4013), .B (n_4104), .Y (n_4643));
AND2X1 g57909(.A (n_4012), .B (n_4095), .Y (n_4641));
AND2X1 g57910(.A (n_4011), .B (n_4104), .Y (n_4639));
AND2X1 g57912(.A (n_4009), .B (n_4103), .Y (n_4634));
AND2X1 g57914(.A (n_4007), .B (n_4106), .Y (n_4630));
AND2X1 g57915(.A (n_4006), .B (n_4096), .Y (n_4627));
AND2X1 g57916(.A (n_4005), .B (n_4096), .Y (n_4623));
AND2X1 g57921(.A (n_4002), .B (n_6633), .Y (n_4617));
AND2X1 g57923(.A (n_4001), .B (n_4096), .Y (n_4614));
AND2X1 g57927(.A (n_3999), .B (n_4101), .Y (n_4610));
AND2X1 g57929(.A (n_3998), .B (n_4017), .Y (n_4607));
AND2X1 g57930(.A (n_3997), .B (n_4017), .Y (n_4605));
AND2X1 g57932(.A (n_3996), .B (n_4017), .Y (n_4602));
AND2X1 g57934(.A (n_3995), .B (n_4017), .Y (n_4599));
AND2X1 g57935(.A (n_3994), .B (n_4017), .Y (n_4597));
AND2X1 g57936(.A (n_3992), .B (n_4017), .Y (n_4595));
AND2X1 g57938(.A (n_3993), .B (n_4017), .Y (n_4592));
AND2X1 g57939(.A (n_3991), .B (n_4017), .Y (n_4590));
AND2X1 g57940(.A (n_3990), .B (n_4017), .Y (n_4588));
AND2X1 g57944(.A (n_3988), .B (n_4105), .Y (n_4583));
AND2X1 g57945(.A (n_3987), .B (n_4099), .Y (n_4581));
AND2X1 g57946(.A (n_3985), .B (n_4105), .Y (n_4578));
AND2X1 g57949(.A (n_3984), .B (n_4094), .Y (n_4574));
AND2X1 g57952(.A (n_4106), .B (n_8345), .Y (n_4572));
AND2X1 g57955(.A (n_3982), .B (n_4105), .Y (n_4570));
AND2X1 g57959(.A (n_3981), .B (n_6452), .Y (n_4568));
AND2X1 g57964(.A (n_4106), .B (n_9401), .Y (n_4280));
AND2X1 g57966(.A (n_3778), .B (n_4058), .Y (n_4195));
AND2X1 g57971(.A (n_3776), .B (n_4094), .Y (n_4276));
AND2X1 g57973(.A (n_3775), .B (n_4016), .Y (n_4193));
AND2X1 g57974(.A (n_3774), .B (n_4016), .Y (n_4191));
AND2X1 g57979(.A (n_3773), .B (n_4015), .Y (n_4188));
AND2X1 g57985(.A (n_3772), .B (n_4016), .Y (n_4186));
AND2X1 g57989(.A (n_3771), .B (n_4058), .Y (n_4183));
AND2X1 g57994(.A (n_3770), .B (n_4016), .Y (n_4181));
AND2X1 g57999(.A (n_3769), .B (n_6633), .Y (n_4254));
AND2X1 g58000(.A (n_3768), .B (n_4016), .Y (n_4179));
AND2X1 g58004(.A (n_3767), .B (n_4104), .Y (n_4252));
AND2X1 g58006(.A (n_3766), .B (n_4015), .Y (n_4176));
AND2X1 g58009(.A (n_3765), .B (n_4103), .Y (n_4250));
AND2X1 g58010(.A (n_3764), .B (n_6452), .Y (n_4248));
AND2X1 g58013(.A (n_3762), .B (n_4016), .Y (n_4174));
AND2X1 g58014(.A (n_3761), .B (n_4104), .Y (n_4244));
AND2X1 g58019(.A (n_3759), .B (n_4058), .Y (n_4172));
CLKBUFX1 gbuf_d_538(.A(n_3846), .Y(d_out_538));
CLKBUFX1 gbuf_qn_538(.A(qn_in_538), .Y(WX8303));
AND2X1 g58024(.A (n_3757), .B (n_4095), .Y (n_4240));
AND2X1 g58025(.A (n_3758), .B (n_4094), .Y (n_4238));
AND2X1 g58026(.A (n_4103), .B (n_9400), .Y (n_4236));
AND2X1 g58028(.A (n_3755), .B (n_4016), .Y (n_4170));
AND2X1 g58030(.A (n_3753), .B (n_4096), .Y (n_4232));
AND2X1 g58034(.A (n_3752), .B (n_4016), .Y (n_4168));
AND2X1 g58037(.A (n_3751), .B (n_4015), .Y (n_4166));
AND2X1 g58040(.A (n_3750), .B (n_4096), .Y (n_4230));
AND2X1 g58041(.A (n_3749), .B (n_4016), .Y (n_4164));
AND2X1 g58043(.A (n_3748), .B (n_4016), .Y (n_4162));
AND2X1 g58045(.A (n_3747), .B (n_4058), .Y (n_4160));
AND2X1 g58046(.A (n_3746), .B (n_4103), .Y (n_4272));
AND2X1 g58050(.A (n_4100), .B (n_8342), .Y (n_4228));
AND2X1 g58054(.A (n_3744), .B (n_4015), .Y (n_4158));
AND2X1 g58059(.A (n_3742), .B (n_4015), .Y (n_4156));
AND2X1 g58063(.A (n_3740), .B (n_4015), .Y (n_4154));
AND2X1 g58071(.A (n_3739), .B (n_4016), .Y (n_4152));
AND2X1 g58074(.A (n_3738), .B (n_4058), .Y (n_4149));
AND2X1 g58078(.A (n_3736), .B (n_4096), .Y (n_4224));
AND2X1 g58081(.A (n_3735), .B (n_4099), .Y (n_4222));
AND2X1 g58083(.A (n_3733), .B (n_4100), .Y (n_4266));
AND2X1 g58084(.A (n_3734), .B (n_4016), .Y (n_4147));
AND2X1 g58086(.A (n_3732), .B (n_4096), .Y (n_4219));
AND2X1 g58087(.A (n_3731), .B (n_4016), .Y (n_4145));
AND2X1 g58093(.A (n_3729), .B (n_4016), .Y (n_4143));
AND2X1 g58097(.A (n_3726), .B (n_4106), .Y (n_4210));
AND2X1 g58101(.A (n_4099), .B (n_8338), .Y (n_4208));
AND2X1 g58102(.A (n_3724), .B (n_4058), .Y (n_4141));
AND2X1 g58105(.A (n_3722), .B (n_4058), .Y (n_4139));
AND2X1 g58107(.A (n_4103), .B (n_9402), .Y (n_4204));
AND2X1 g58110(.A (n_3719), .B (n_4016), .Y (n_4137));
AND2X1 g58111(.A (n_3718), .B (n_4015), .Y (n_4135));
AND2X1 g58115(.A (n_3716), .B (n_4016), .Y (n_4133));
AND2X1 g58117(.A (n_3715), .B (n_4101), .Y (n_4264));
AND2X1 g58118(.A (n_3714), .B (n_4100), .Y (n_4262));
AND2X1 g58126(.A (n_3713), .B (n_4106), .Y (n_4131));
AND2X1 g58127(.A (n_3712), .B (n_4103), .Y (n_4260));
AND2X1 g58128(.A (n_3711), .B (n_4096), .Y (n_4129));
AND2X1 g58129(.A (n_3710), .B (n_4095), .Y (n_4127));
AND2X1 g58131(.A (n_3709), .B (n_4096), .Y (n_4124));
AND2X1 g58133(.A (n_3708), .B (n_4095), .Y (n_4258));
AND2X1 g58141(.A (n_3707), .B (n_4096), .Y (n_4256));
AND2X1 g58143(.A (n_4101), .B (n_8339), .Y (n_4122));
AND2X1 g58152(.A (n_3703), .B (n_4096), .Y (n_4116));
AND2X1 g58155(.A (n_3702), .B (n_4096), .Y (n_4114));
AND2X1 g58156(.A (n_3701), .B (n_4101), .Y (n_4112));
CLKBUFX1 gbuf_d_539(.A(n_3800), .Y(d_out_539));
CLKBUFX1 gbuf_qn_539(.A(qn_in_539), .Y(WX9596));
CLKBUFX1 gbuf_d_540(.A(n_3696), .Y(d_out_540));
CLKBUFX1 gbuf_q_540(.A(q_in_540), .Y(WX545));
NOR2X1 g57441(.A (n_3699), .B (n_3269), .Y (n_4329));
CLKBUFX1 gbuf_d_541(.A(n_3694), .Y(d_out_541));
CLKBUFX1 gbuf_qn_541(.A(qn_in_541), .Y(WX3131));
CLKBUFX1 gbuf_d_542(.A(n_3691), .Y(d_out_542));
CLKBUFX1 gbuf_qn_542(.A(qn_in_542), .Y(WX5717));
CLKBUFX1 gbuf_d_543(.A(n_3848), .Y(d_out_543));
CLKBUFX1 gbuf_qn_543(.A(qn_in_543), .Y(WX7010));
AND2X1 g57905(.A (n_3805), .B (n_4103), .Y (n_4325));
AND2X1 g57907(.A (n_3804), .B (n_4103), .Y (n_4323));
AND2X1 g57920(.A (n_3802), .B (n_4096), .Y (n_4318));
AND2X1 g57922(.A (n_3801), .B (n_4096), .Y (n_4316));
AND2X1 g57925(.A (n_3799), .B (n_4101), .Y (n_4314));
AND2X1 g57926(.A (n_3798), .B (n_4101), .Y (n_4312));
AND2X1 g57928(.A (n_3796), .B (n_4096), .Y (n_4310));
AND2X1 g57931(.A (n_3795), .B (n_4017), .Y (n_4308));
AND2X1 g57937(.A (n_3793), .B (n_4105), .Y (n_4304));
AND2X1 g57942(.A (n_3792), .B (n_4017), .Y (n_4302));
AND2X1 g57948(.A (n_3790), .B (n_4058), .Y (n_4198));
AND2X1 g57950(.A (n_4099), .B (n_8343), .Y (n_4298));
AND2X1 g57953(.A (n_3787), .B (n_4104), .Y (n_4294));
AND2X1 g57954(.A (n_3786), .B (n_4105), .Y (n_4292));
AND2X1 g57956(.A (n_3785), .B (n_4094), .Y (n_4290));
AND2X1 g57957(.A (n_4094), .B (n_8348), .Y (n_4288));
AND2X1 g57958(.A (n_3783), .B (n_4106), .Y (n_4274));
AND2X1 g57960(.A (n_3782), .B (n_4094), .Y (n_4286));
AND2X1 g57961(.A (n_3781), .B (n_4105), .Y (n_4282));
XOR2X1 g58226(.A (n_812), .B (n_3596), .Y (n_4014));
XOR2X1 g58228(.A (n_811), .B (n_3595), .Y (n_4013));
XOR2X1 g58229(.A (n_810), .B (n_3594), .Y (n_4012));
XOR2X1 g58230(.A (n_507), .B (n_3593), .Y (n_4011));
XOR2X1 g58231(.A (n_809), .B (n_3592), .Y (n_8323));
XOR2X1 g58232(.A (n_770), .B (n_3591), .Y (n_4009));
XOR2X1 g58234(.A (n_508), .B (n_3589), .Y (n_4007));
XOR2X1 g58235(.A (n_807), .B (n_3588), .Y (n_4006));
XOR2X1 g58236(.A (n_803), .B (n_3587), .Y (n_4005));
XOR2X1 g58237(.A (n_806), .B (n_3586), .Y (n_8314));
XOR2X1 g58239(.A (n_515), .B (n_3585), .Y (n_8317));
XOR2X1 g58241(.A (n_801), .B (n_3584), .Y (n_4002));
XOR2X1 g58243(.A (n_799), .B (n_3583), .Y (n_4001));
XOR2X1 g58244(.A (n_798), .B (n_3582), .Y (n_4000));
XOR2X1 g58247(.A (n_794), .B (n_3581), .Y (n_3999));
XOR2X1 g58249(.A (n_791), .B (n_3580), .Y (n_3998));
XOR2X1 g58250(.A (n_619), .B (n_3579), .Y (n_3997));
XOR2X1 g58252(.A (n_790), .B (n_3578), .Y (n_3996));
XOR2X1 g58253(.A (n_623), .B (n_3577), .Y (n_3995));
XOR2X1 g58255(.A (n_643), .B (n_3576), .Y (n_3994));
XOR2X1 g58256(.A (n_670), .B (n_3575), .Y (n_3993));
XOR2X1 g58257(.A (n_787), .B (n_3574), .Y (n_3992));
XOR2X1 g58259(.A (n_789), .B (n_3573), .Y (n_3991));
XOR2X1 g58260(.A (n_786), .B (n_3572), .Y (n_3990));
XOR2X1 g58261(.A (n_785), .B (n_3571), .Y (n_8318));
XOR2X1 g58263(.A (n_757), .B (n_3570), .Y (n_3988));
XOR2X1 g58265(.A (n_783), .B (n_3569), .Y (n_3987));
XOR2X1 g58266(.A (n_793), .B (n_3568), .Y (n_8316));
XOR2X1 g58267(.A (n_781), .B (n_3567), .Y (n_3985));
XOR2X1 g58269(.A (n_780), .B (n_3566), .Y (n_3984));
XOR2X1 g58272(.A (n_778), .B (n_3565), .Y (n_8345));
XOR2X1 g58275(.A (n_637), .B (n_3564), .Y (n_3982));
XOR2X1 g58278(.A (n_688), .B (n_3492), .Y (n_3981));
XOR2X1 g58283(.A (n_802), .B (n_3538), .Y (n_3980));
XOR2X1 g58285(.A (n_755), .B (n_3563), .Y (n_3979));
XOR2X1 g58287(.A (n_768), .B (n_3562), .Y (n_8321));
XOR2X1 g58289(.A (n_765), .B (n_3561), .Y (n_3977));
XOR2X1 g58290(.A (n_503), .B (n_3560), .Y (n_3976));
XOR2X1 g58292(.A (n_530), .B (n_3559), .Y (n_3975));
XOR2X1 g58295(.A (n_723), .B (n_3558), .Y (n_3974));
XOR2X1 g58296(.A (n_762), .B (n_3557), .Y (n_3973));
XOR2X1 g58297(.A (n_758), .B (n_3556), .Y (n_3972));
XOR2X1 g58298(.A (n_756), .B (n_3501), .Y (n_3971));
XOR2X1 g58300(.A (n_750), .B (n_3555), .Y (n_3970));
XOR2X1 g58301(.A (n_752), .B (n_3554), .Y (n_3969));
XOR2X1 g58302(.A (n_748), .B (n_3552), .Y (n_3968));
XOR2X1 g58303(.A (n_749), .B (n_3553), .Y (n_3967));
XOR2X1 g58304(.A (n_746), .B (n_3550), .Y (n_3966));
XOR2X1 g58306(.A (n_671), .B (n_3549), .Y (n_3965));
XOR2X1 g58307(.A (n_650), .B (n_3547), .Y (n_3964));
XOR2X1 g58308(.A (n_782), .B (n_3548), .Y (n_3963));
XOR2X1 g58310(.A (n_702), .B (n_3546), .Y (n_3962));
XOR2X1 g58311(.A (n_742), .B (n_3545), .Y (n_3961));
XOR2X1 g58312(.A (n_743), .B (n_3544), .Y (n_3960));
XOR2X1 g58313(.A (n_715), .B (n_3543), .Y (n_3959));
XOR2X1 g58315(.A (n_531), .B (n_3542), .Y (n_3958));
XOR2X1 g58316(.A (n_700), .B (n_3541), .Y (n_3957));
XOR2X1 g58317(.A (n_706), .B (n_3539), .Y (n_3956));
XOR2X1 g58318(.A (n_741), .B (n_3540), .Y (n_3955));
XOR2X1 g58321(.A (n_535), .B (n_3537), .Y (n_3954));
XOR2X1 g58322(.A (n_766), .B (n_3535), .Y (n_3953));
XOR2X1 g58323(.A (n_731), .B (n_3536), .Y (n_3952));
XOR2X1 g58325(.A (n_737), .B (n_3475), .Y (n_3951));
XOR2X1 g58327(.A (n_647), .B (n_3534), .Y (n_7281));
XOR2X1 g58328(.A (n_759), .B (n_3533), .Y (n_8324));
XOR2X1 g58331(.A (n_730), .B (n_3532), .Y (n_3948));
XOR2X1 g58335(.A (n_727), .B (n_3531), .Y (n_3947));
XOR2X1 g58336(.A (n_720), .B (n_3597), .Y (n_8326));
XOR2X1 g58338(.A (n_722), .B (n_3551), .Y (n_3945));
XOR2X1 g58340(.A (n_526), .B (n_3530), .Y (n_3944));
XOR2X1 g58341(.A (n_725), .B (n_3529), .Y (n_3943));
XOR2X1 g58342(.A (n_602), .B (n_6425), .Y (n_3942));
XOR2X1 g58343(.A (n_740), .B (n_3474), .Y (n_3941));
XOR2X1 g58346(.A (n_504), .B (n_3527), .Y (n_3940));
XOR2X1 g58351(.A (n_788), .B (n_3526), .Y (n_3939));
XOR2X1 g58352(.A (n_721), .B (n_3525), .Y (n_3938));
XOR2X1 g58353(.A (n_519), .B (n_3523), .Y (n_3937));
XOR2X1 g58355(.A (n_760), .B (n_3524), .Y (n_3936));
XOR2X1 g58356(.A (n_625), .B (n_3522), .Y (n_8355));
XOR2X1 g58358(.A (n_734), .B (n_3521), .Y (n_3934));
XOR2X1 g58359(.A (n_719), .B (n_3520), .Y (n_3933));
XOR2X1 g58362(.A (n_714), .B (n_3519), .Y (n_3932));
XOR2X1 g58364(.A (n_713), .B (n_3518), .Y (n_8340));
XOR2X1 g58367(.A (n_709), .B (n_3517), .Y (n_3930));
XOR2X1 g58368(.A (n_711), .B (n_3516), .Y (n_6884));
XOR2X1 g58371(.A (n_708), .B (n_3514), .Y (n_3927));
XOR2X1 g58372(.A (n_705), .B (n_3513), .Y (n_3926));
XOR2X1 g58373(.A (n_701), .B (n_3512), .Y (n_3925));
XOR2X1 g58375(.A (n_703), .B (n_3511), .Y (n_3924));
XOR2X1 g58377(.A (n_763), .B (n_3510), .Y (n_3923));
XOR2X1 g58378(.A (n_698), .B (n_3509), .Y (n_3922));
XOR2X1 g58380(.A (n_696), .B (n_3508), .Y (n_3921));
XOR2X1 g58382(.A (n_695), .B (n_3507), .Y (n_3920));
XOR2X1 g58384(.A (n_690), .B (n_3506), .Y (n_3919));
XOR2X1 g58385(.A (n_689), .B (n_3504), .Y (n_8346));
XOR2X1 g58386(.A (n_491), .B (n_3505), .Y (n_3917));
XOR2X1 g58387(.A (n_492), .B (n_3503), .Y (n_3916));
XOR2X1 g58388(.A (n_685), .B (n_3498), .Y (n_3915));
XOR2X1 g58389(.A (n_686), .B (n_3500), .Y (n_3914));
XOR2X1 g58390(.A (n_495), .B (n_3502), .Y (n_3913));
XOR2X1 g58391(.A (n_684), .B (n_3499), .Y (n_3912));
XOR2X1 g58393(.A (n_681), .B (n_3497), .Y (n_3911));
XOR2X1 g58395(.A (n_496), .B (n_3496), .Y (n_3910));
XOR2X1 g58397(.A (n_678), .B (n_3495), .Y (n_8325));
XOR2X1 g58399(.A (n_675), .B (n_3494), .Y (n_3908));
XOR2X1 g58400(.A (n_497), .B (n_3493), .Y (n_8341));
XOR2X1 g58402(.A (n_672), .B (n_3491), .Y (n_3906));
XOR2X1 g58405(.A (n_669), .B (n_3490), .Y (n_8344));
XOR2X1 g58409(.A (n_662), .B (n_3488), .Y (n_8319));
XOR2X1 g58410(.A (n_728), .B (n_3489), .Y (n_3903));
XOR2X1 g58411(.A (n_661), .B (n_3487), .Y (n_8349));
XOR2X1 g58412(.A (n_659), .B (n_3486), .Y (n_3901));
XOR2X1 g58415(.A (n_657), .B (n_3485), .Y (n_3900));
XOR2X1 g58418(.A (n_654), .B (n_3484), .Y (n_8353));
XOR2X1 g58419(.A (n_651), .B (n_3483), .Y (n_3898));
XOR2X1 g58420(.A (n_653), .B (n_3482), .Y (n_8351));
XOR2X1 g58424(.A (n_645), .B (n_3481), .Y (n_9403));
XOR2X1 g58426(.A (n_641), .B (n_3480), .Y (n_3895));
XOR2X1 g58429(.A (n_500), .B (n_3479), .Y (n_3894));
XOR2X1 g58433(.A (n_501), .B (n_3478), .Y (n_3893));
XOR2X1 g58434(.A (n_638), .B (n_3477), .Y (n_3892));
XOR2X1 g58436(.A (n_636), .B (n_3476), .Y (n_3891));
XOR2X1 g58439(.A (n_630), .B (n_7485), .Y (n_3890));
XOR2X1 g58440(.A (n_735), .B (n_3472), .Y (n_3889));
XOR2X1 g58441(.A (n_629), .B (n_3471), .Y (n_3888));
XOR2X1 g58442(.A (n_626), .B (n_3469), .Y (n_3887));
XOR2X1 g58443(.A (n_764), .B (n_3470), .Y (n_3886));
XOR2X1 g58444(.A (n_627), .B (n_3468), .Y (n_3885));
XOR2X1 g58445(.A (n_808), .B (n_3467), .Y (n_3884));
XOR2X1 g58450(.A (n_617), .B (n_3466), .Y (n_3883));
XOR2X1 g58451(.A (n_616), .B (n_3465), .Y (n_3882));
XOR2X1 g58453(.A (n_506), .B (n_3464), .Y (n_3881));
XOR2X1 g58455(.A (n_509), .B (n_3462), .Y (n_3880));
XOR2X1 g58456(.A (n_614), .B (n_3463), .Y (n_3879));
XOR2X1 g58457(.A (n_612), .B (n_3461), .Y (n_3878));
XOR2X1 g58458(.A (n_510), .B (n_3460), .Y (n_3877));
XOR2X1 g58459(.A (n_610), .B (n_3459), .Y (n_3876));
XOR2X1 g58460(.A (n_609), .B (n_3458), .Y (n_3875));
XOR2X1 g58462(.A (n_607), .B (n_3457), .Y (n_3874));
XOR2X1 g58464(.A (n_514), .B (n_3456), .Y (n_8315));
XOR2X1 g58465(.A (n_604), .B (n_3455), .Y (n_3872));
XOR2X1 g58467(.A (n_516), .B (n_3454), .Y (n_3871));
XOR2X1 g58469(.A (n_634), .B (n_3453), .Y (n_3870));
XOR2X1 g58470(.A (n_603), .B (n_3452), .Y (n_8327));
XOR2X1 g58471(.A (n_601), .B (n_3451), .Y (n_3868));
XOR2X1 g58473(.A (n_600), .B (n_3450), .Y (n_8347));
XOR2X1 g58474(.A (n_683), .B (n_3449), .Y (n_7282));
XOR2X1 g58478(.A (n_815), .B (n_3598), .Y (n_3865));
NAND2X1 g58480(.A (n_3682), .B (n_3633), .Y (n_4079));
NAND2X1 g58481(.A (n_3681), .B (n_3632), .Y (n_4076));
NAND2X2 g58483(.A (n_3678), .B (n_3628), .Y (n_4071));
NAND2X2 g58485(.A (n_3676), .B (n_3621), .Y (n_4069));
NAND2X1 g58488(.A (n_3679), .B (n_3626), .Y (n_4061));
NAND2X2 g58492(.A (n_3670), .B (n_3622), .Y (n_4052));
NAND2X1 g58493(.A (n_3669), .B (n_3620), .Y (n_4050));
NAND2X2 g58496(.A (n_3666), .B (n_3616), .Y (n_4044));
NAND2X2 g58498(.A (n_3664), .B (n_3612), .Y (n_4040));
NAND2X1 g58499(.A (n_3663), .B (n_3614), .Y (n_4038));
NAND2X1 g58505(.A (n_3658), .B (n_3609), .Y (n_4026));
NAND2X1 g58509(.A (n_3684), .B (n_3637), .Y (n_4018));
NOR2X1 g58599(.A (WX3097), .B (n_3218), .Y (n_3864));
NOR2X1 g58601(.A (WX8261), .B (n_5181), .Y (n_3863));
NOR2X1 g58603(.A (WX8261), .B (n_5838), .Y (n_6662));
NOR2X1 g58606(.A (WX9552), .B (n_2851), .Y (n_3860));
NOR2X1 g58607(.A (WX4388), .B (n_1425), .Y (n_3859));
NOR2X1 g58608(.A (WX4388), .B (n_5838), .Y (n_3857));
NOR2X1 g58610(.A (WX5679), .B (n_5712), .Y (n_3856));
NOR2X1 g58611(.A (WX5679), .B (n_5838), .Y (n_3855));
NOR2X1 g58613(.A (WX6970), .B (n_5712), .Y (n_3854));
NOR2X1 g58616(.A (WX3097), .B (n_5712), .Y (n_3853));
NOR2X1 g58617(.A (WX6970), .B (n_5662), .Y (n_6207));
NOR2X1 g58619(.A (WX9552), .B (n_5479), .Y (n_3850));
CLKBUFX1 gbuf_d_544(.A(n_3647), .Y(d_out_544));
CLKBUFX1 gbuf_qn_544(.A(qn_in_544), .Y(WX1838));
CLKBUFX1 gbuf_d_545(.A(n_3650), .Y(d_out_545));
CLKBUFX1 gbuf_qn_545(.A(qn_in_545), .Y(WX10889));
NOR2X1 g57442(.A (n_3652), .B (n_4150), .Y (n_4087));
CLKBUFX1 gbuf_d_546(.A(n_3643), .Y(d_out_546));
CLKBUFX1 gbuf_qn_546(.A(qn_in_546), .Y(WX4426));
NOR2X1 g56941(.A (WX7012), .B (n_1425), .Y (n_3848));
NOR2X1 g56978(.A (WX8305), .B (n_1425), .Y (n_3846));
NOR2X1 g56982(.A (WX8305), .B (n_5479), .Y (n_3845));
AOI22X1 g60674(.A0 (DATA_0_19), .A1 (n_3828), .B0 (_2352_), .B1(n_5873), .Y (n_3844));
AOI22X1 g60675(.A0 (DATA_0_31), .A1 (n_5968), .B0 (_2364_), .B1(n_3831), .Y (n_3843));
AOI22X1 g60676(.A0 (DATA_0_30), .A1 (n_5968), .B0 (_2363_), .B1(n_3840), .Y (n_3842));
AOI22X1 g60677(.A0 (DATA_0_29), .A1 (n_4670), .B0 (_2362_), .B1(n_3840), .Y (n_3841));
AOI22X1 g60678(.A0 (DATA_0_27), .A1 (n_3828), .B0 (_2360_), .B1(n_3840), .Y (n_3839));
AOI22X1 g60679(.A0 (DATA_0_26), .A1 (n_3828), .B0 (_2359_), .B1(n_3835), .Y (n_3837));
AOI22X1 g60680(.A0 (DATA_0_24), .A1 (n_4882), .B0 (_2357_), .B1(n_3835), .Y (n_3836));
AOI22X1 g60681(.A0 (DATA_0_28), .A1 (n_3828), .B0 (_2361_), .B1(n_3831), .Y (n_3834));
AOI22X1 g60682(.A0 (DATA_0_21), .A1 (n_5968), .B0 (_2354_), .B1(n_3831), .Y (n_3833));
AOI22X1 g60683(.A0 (DATA_0_22), .A1 (n_4670), .B0 (_2355_), .B1(n_3831), .Y (n_3830));
AOI22X1 g60684(.A0 (DATA_0_17), .A1 (n_3828), .B0 (_2350_), .B1(n_3835), .Y (n_3829));
AOI22X1 g60685(.A0 (DATA_0_23), .A1 (n_4670), .B0 (_2356_), .B1(n_3835), .Y (n_3827));
AOI22X1 g60686(.A0 (DATA_0_16), .A1 (n_4882), .B0 (_2349_), .B1(n_3835), .Y (n_3826));
AOI22X1 g60688(.A0 (DATA_0_14), .A1 (n_4882), .B0 (_2347_), .B1(n_3835), .Y (n_3824));
AOI22X1 g60690(.A0 (DATA_0_25), .A1 (n_4670), .B0 (_2358_), .B1(n_3835), .Y (n_3822));
AOI22X1 g60691(.A0 (DATA_0_12), .A1 (n_5968), .B0 (_2345_), .B1(n_3840), .Y (n_3821));
AOI22X1 g60692(.A0 (DATA_0_20), .A1 (n_5968), .B0 (_2353_), .B1(n_3840), .Y (n_3819));
AOI22X1 g60693(.A0 (DATA_0_4), .A1 (n_3828), .B0 (_2337_), .B1(n_3840), .Y (n_3818));
AOI22X1 g60694(.A0 (DATA_0_11), .A1 (n_5968), .B0 (_2344_), .B1(n_3840), .Y (n_3817));
AOI22X1 g60695(.A0 (DATA_0_10), .A1 (n_5968), .B0 (_2343_), .B1(n_3840), .Y (n_3816));
AOI22X1 g60696(.A0 (DATA_0_9), .A1 (n_5968), .B0 (_2342_), .B1(n_3840), .Y (n_3815));
AOI22X1 g60698(.A0 (DATA_0_7), .A1 (n_5968), .B0 (_2340_), .B1(n_5873), .Y (n_3813));
AOI22X1 g60699(.A0 (DATA_0_18), .A1 (n_3828), .B0 (_2351_), .B1(n_5873), .Y (n_3812));
AOI22X1 g60700(.A0 (DATA_0_6), .A1 (n_3828), .B0 (_2339_), .B1(n_3840), .Y (n_3811));
AOI22X1 g60701(.A0 (DATA_0_5), .A1 (n_3828), .B0 (_2338_), .B1(n_3840), .Y (n_3810));
AOI22X1 g60702(.A0 (DATA_0_3), .A1 (n_3828), .B0 (_2336_), .B1(n_3835), .Y (n_3809));
AOI22X1 g60703(.A0 (DATA_0_2), .A1 (n_5968), .B0 (_2335_), .B1(n_3835), .Y (n_3808));
AOI22X1 g60704(.A0 (DATA_0_1), .A1 (n_5968), .B0 (_2334_), .B1(n_3840), .Y (n_3807));
AOI22X1 g60705(.A0 (DATA_0_0), .A1 (n_3828), .B0 (_2333_), .B1(n_3835), .Y (n_3806));
XOR2X1 g58225(.A (n_538), .B (n_3409), .Y (n_3805));
XOR2X1 g58227(.A (n_814), .B (n_3408), .Y (n_3804));
XOR2X1 g58238(.A (n_805), .B (n_3403), .Y (n_9389));
XOR2X1 g58240(.A (n_804), .B (n_3402), .Y (n_3802));
XOR2X1 g58242(.A (n_800), .B (n_3401), .Y (n_3801));
NOR2X1 g57043(.A (WX9598), .B (n_5181), .Y (n_3800));
XOR2X1 g58245(.A (n_796), .B (n_3400), .Y (n_3799));
XOR2X1 g58246(.A (n_795), .B (n_3399), .Y (n_3798));
NOR2X1 g57046(.A (WX9598), .B (n_5838), .Y (n_8546));
XOR2X1 g58248(.A (n_792), .B (n_3398), .Y (n_3796));
XOR2X1 g58251(.A (n_736), .B (n_3397), .Y (n_3795));
XOR2X1 g58254(.A (n_521), .B (n_3394), .Y (n_9396));
XOR2X1 g58258(.A (n_522), .B (n_3393), .Y (n_3793));
XOR2X1 g58262(.A (n_784), .B (n_3390), .Y (n_3792));
XOR2X1 g58264(.A (n_773), .B (n_3389), .Y (n_9398));
XOR2X1 g58268(.A (n_813), .B (n_3388), .Y (n_3790));
XOR2X1 g58270(.A (n_744), .B (n_3387), .Y (n_8343));
XOR2X1 g58271(.A (n_779), .B (n_3386), .Y (n_9385));
XOR2X1 g58273(.A (n_525), .B (n_3385), .Y (n_3787));
XOR2X1 g58274(.A (n_631), .B (n_3257), .Y (n_3786));
XOR2X1 g58276(.A (n_777), .B (n_3384), .Y (n_3785));
XOR2X1 g58277(.A (n_674), .B (n_3379), .Y (n_8348));
XOR2X1 g58279(.A (n_772), .B (n_3378), .Y (n_3783));
XOR2X1 g58280(.A (n_527), .B (n_3376), .Y (n_3782));
XOR2X1 g58281(.A (n_775), .B (n_3375), .Y (n_3781));
XOR2X1 g58282(.A (n_776), .B (n_3374), .Y (n_9384));
XOR2X1 g58284(.A (n_774), .B (n_3373), .Y (n_9401));
XOR2X1 g58286(.A (n_767), .B (n_3372), .Y (n_3778));
XOR2X1 g58288(.A (n_529), .B (n_3371), .Y (n_9387));
XOR2X1 g58291(.A (n_599), .B (n_3370), .Y (n_3776));
XOR2X1 g58293(.A (n_691), .B (n_3369), .Y (n_3775));
XOR2X1 g58294(.A (n_754), .B (n_3366), .Y (n_3774));
XOR2X1 g58299(.A (n_753), .B (n_3363), .Y (n_3773));
XOR2X1 g58305(.A (n_745), .B (n_3360), .Y (n_3772));
XOR2X1 g58309(.A (n_532), .B (n_3359), .Y (n_3771));
XOR2X1 g58314(.A (n_628), .B (n_3356), .Y (n_3770));
XOR2X1 g58319(.A (n_739), .B (n_3352), .Y (n_3769));
XOR2X1 g58320(.A (n_667), .B (n_3349), .Y (n_3768));
XOR2X1 g58324(.A (n_738), .B (n_3348), .Y (n_3767));
XOR2X1 g58326(.A (n_632), .B (n_3377), .Y (n_3766));
XOR2X1 g58329(.A (n_733), .B (n_3345), .Y (n_3765));
XOR2X1 g58330(.A (n_633), .B (n_3344), .Y (n_3764));
XOR2X1 g58332(.A (n_732), .B (n_3343), .Y (n_9390));
XOR2X1 g58333(.A (n_747), .B (n_3342), .Y (n_3762));
XOR2X1 g58334(.A (n_729), .B (n_3341), .Y (n_3761));
XOR2X1 g58337(.A (n_518), .B (n_3340), .Y (n_9394));
XOR2X1 g58339(.A (n_726), .B (n_3339), .Y (n_3759));
XOR2X1 g58344(.A (n_536), .B (n_3336), .Y (n_3758));
XOR2X1 g58345(.A (n_724), .B (n_3335), .Y (n_3757));
XOR2X1 g58347(.A (n_505), .B (n_3353), .Y (n_9400));
XOR2X1 g58348(.A (n_537), .B (n_3334), .Y (n_3755));
XOR2X1 g58349(.A (n_797), .B (n_3333), .Y (n_8352));
XOR2X1 g58350(.A (n_751), .B (n_3330), .Y (n_3753));
XOR2X1 g58354(.A (n_622), .B (n_3327), .Y (n_3752));
XOR2X1 g58357(.A (n_761), .B (n_3324), .Y (n_3751));
XOR2X1 g58360(.A (n_611), .B (n_3323), .Y (n_3750));
XOR2X1 g58361(.A (n_718), .B (n_3272), .Y (n_3749));
XOR2X1 g58363(.A (n_717), .B (n_3322), .Y (n_3748));
XOR2X1 g58365(.A (n_712), .B (n_3319), .Y (n_3747));
XOR2X1 g58366(.A (n_710), .B (n_3318), .Y (n_3746));
XOR2X1 g58370(.A (n_707), .B (n_3315), .Y (n_8342));
XOR2X1 g58374(.A (n_704), .B (n_3314), .Y (n_3744));
XOR2X1 g58376(.A (n_699), .B (n_3313), .Y (n_9392));
XOR2X1 g58379(.A (n_697), .B (n_3312), .Y (n_3742));
XOR2X1 g58381(.A (n_693), .B (n_3311), .Y (n_3741));
XOR2X1 g58383(.A (n_692), .B (n_3310), .Y (n_3740));
XOR2X1 g58392(.A (n_682), .B (n_3305), .Y (n_3739));
XOR2X1 g58394(.A (n_680), .B (n_3304), .Y (n_3738));
XOR2X1 g58396(.A (n_677), .B (n_3303), .Y (n_3737));
XOR2X1 g58398(.A (n_676), .B (n_3302), .Y (n_3736));
XOR2X1 g58401(.A (n_673), .B (n_3301), .Y (n_3735));
XOR2X1 g58403(.A (n_668), .B (n_3300), .Y (n_3734));
XOR2X1 g58404(.A (n_665), .B (n_3299), .Y (n_3733));
XOR2X1 g58406(.A (n_666), .B (n_6515), .Y (n_3732));
XOR2X1 g58407(.A (n_664), .B (n_3297), .Y (n_3731));
XOR2X1 g58408(.A (n_663), .B (n_3296), .Y (n_9395));
XOR2X1 g58413(.A (n_658), .B (n_3293), .Y (n_3729));
XOR2X1 g58414(.A (n_660), .B (n_3292), .Y (n_9397));
XOR2X1 g58416(.A (n_655), .B (n_3291), .Y (n_9399));
XOR2X1 g58417(.A (n_499), .B (n_3290), .Y (n_3726));
XOR2X1 g58421(.A (n_652), .B (n_3287), .Y (n_8338));
XOR2X1 g58422(.A (n_648), .B (n_3286), .Y (n_3724));
XOR2X1 g58423(.A (n_649), .B (n_3285), .Y (n_9388));
XOR2X1 g58425(.A (n_644), .B (n_3282), .Y (n_3722));
XOR2X1 g58427(.A (n_642), .B (n_3281), .Y (n_9402));
XOR2X1 g58428(.A (n_687), .B (n_3280), .Y (n_9386));
XOR2X1 g58430(.A (n_656), .B (n_3278), .Y (n_3719));
XOR2X1 g58431(.A (n_640), .B (n_3276), .Y (n_3718));
XOR2X1 g58432(.A (n_639), .B (n_3273), .Y (n_8354));
XOR2X1 g58435(.A (n_502), .B (n_3268), .Y (n_3716));
XOR2X1 g58437(.A (n_635), .B (n_3265), .Y (n_3715));
XOR2X1 g58438(.A (n_716), .B (n_3260), .Y (n_3714));
XOR2X1 g58446(.A (n_831), .B (n_3256), .Y (n_3713));
XOR2X1 g58447(.A (n_618), .B (n_3254), .Y (n_3712));
XOR2X1 g58448(.A (n_621), .B (n_3255), .Y (n_3711));
XOR2X1 g58449(.A (n_620), .B (n_3253), .Y (n_3710));
XOR2X1 g58452(.A (n_615), .B (n_3250), .Y (n_3709));
XOR2X1 g58454(.A (n_613), .B (n_3249), .Y (n_3708));
XOR2X1 g58461(.A (n_606), .B (n_3244), .Y (n_3707));
XOR2X1 g58463(.A (n_608), .B (n_3243), .Y (n_8339));
XOR2X1 g58466(.A (n_605), .B (n_3242), .Y (n_9391));
XOR2X1 g58468(.A (n_624), .B (n_3241), .Y (n_9393));
XOR2X1 g58472(.A (n_646), .B (n_3240), .Y (n_3703));
XOR2X1 g58475(.A (n_679), .B (n_3239), .Y (n_3702));
XOR2X1 g58476(.A (n_598), .B (n_3238), .Y (n_3701));
XOR2X1 g58477(.A (n_816), .B (n_3237), .Y (n_8350));
XOR2X1 g57506(.A (n_850), .B (n_3414), .Y (n_3699));
NOR2X1 g56747(.A (WX3133), .B (n_5662), .Y (n_3698));
NOR2X1 g59506(.A (n_1425), .B (n_3695), .Y (n_3696));
NOR2X1 g56767(.A (WX3133), .B (n_1648), .Y (n_3694));
OR2X1 g59514(.A (n_3695), .B (n_5990), .Y (n_3692));
CLKBUFX1 gbuf_d_547(.A(n_3606), .Y(d_out_547));
CLKBUFX1 gbuf_q_547(.A(q_in_547), .Y(_2081_));
CLKBUFX1 gbuf_d_548(.A(n_3605), .Y(d_out_548));
CLKBUFX1 gbuf_q_548(.A(q_in_548), .Y(_2088_));
CLKBUFX1 gbuf_d_549(.A(n_3604), .Y(d_out_549));
CLKBUFX1 gbuf_q_549(.A(q_in_549), .Y(_2093_));
NOR2X1 g56875(.A (WX5719), .B (n_3690), .Y (n_3691));
NOR2X1 g56880(.A (WX5719), .B (n_5427), .Y (n_3689));
NOR2X1 g56919(.A (WX7012), .B (n_5500), .Y (n_3688));
NOR2X1 g57097(.A (WX8245), .B (n_5662), .Y (n_6670));
OR2X1 g55937(.A (n_3685), .B (n_4882), .Y (n_3686));
NAND2X1 g58510(.A (n_3411), .B (n_2512), .Y (n_3684));
NAND2X1 g58514(.A (n_3405), .B (n_2454), .Y (n_3682));
NAND2X1 g58518(.A (n_3396), .B (n_2499), .Y (n_3681));
NAND2X1 g58520(.A (n_3362), .B (n_2473), .Y (n_3679));
NAND2X2 g58522(.A (n_3383), .B (n_2495), .Y (n_3678));
NAND2X2 g58526(.A (n_3365), .B (n_2447), .Y (n_3676));
NAND2X2 g58539(.A (n_3347), .B (n_2467), .Y (n_3670));
NAND2X1 g58541(.A (n_3338), .B (n_2469), .Y (n_3669));
NAND2X2 g58549(.A (n_3321), .B (n_2459), .Y (n_3666));
NAND2X2 g58552(.A (n_3309), .B (n_2438), .Y (n_3664));
NAND2X1 g58553(.A (n_3307), .B (n_2444), .Y (n_3663));
NAND2X1 g58564(.A (n_3262), .B (n_2423), .Y (n_3658));
CLKBUFX1 gbuf_d_550(.A(n_3236), .Y(d_out_550));
CLKBUFX1 gbuf_qn_550(.A(qn_in_550), .Y(WX8261));
CLKBUFX1 gbuf_d_551(.A(n_3235), .Y(d_out_551));
CLKBUFX1 gbuf_qn_551(.A(qn_in_551), .Y(WX9552));
CLKBUFX1 gbuf_d_552(.A(n_3234), .Y(d_out_552));
CLKBUFX1 gbuf_qn_552(.A(qn_in_552), .Y(WX4388));
CLKBUFX1 gbuf_d_553(.A(n_3233), .Y(d_out_553));
CLKBUFX1 gbuf_qn_553(.A(qn_in_553), .Y(WX5679));
CLKBUFX1 gbuf_d_554(.A(n_3231), .Y(d_out_554));
CLKBUFX1 gbuf_qn_554(.A(qn_in_554), .Y(WX6970));
CLKBUFX1 gbuf_d_555(.A(n_3230), .Y(d_out_555));
CLKBUFX1 gbuf_qn_555(.A(qn_in_555), .Y(WX3097));
OR2X1 g55877(.A (n_2888), .B (n_3828), .Y (n_3653));
XOR2X1 g57507(.A (n_849), .B (n_3178), .Y (n_3652));
NOR2X1 g59503(.A (WX10891), .B (n_1648), .Y (n_3650));
NOR2X1 g59510(.A (WX4390), .B (n_5479), .Y (n_6205));
NOR2X1 g59511(.A (WX1840), .B (n_5479), .Y (n_3648));
NOR2X1 g59515(.A (WX1840), .B (n_1425), .Y (n_3647));
NOR2X1 g59517(.A (WX6972), .B (n_5662), .Y (n_6677));
NOR2X1 g59518(.A (WX10891), .B (n_5662), .Y (n_7511));
NOR2X1 g56868(.A (WX4364), .B (n_2605), .Y (n_3643));
AND2X1 g56869(.A (WX4364), .B (n_5873), .Y (n_3642));
NOR2X1 g56927(.A (WX4366), .B (n_5427), .Y (n_6669));
CLKBUFX1 gbuf_d_556(.A(n_3219), .Y(d_out_556));
CLKBUFX1 gbuf_qn_556(.A(qn_in_556), .Y(WX7012));
INVX1 g60387(.A (WX547), .Y (n_3695));
NOR2X1 g56991(.A (WX5659), .B (n_5838), .Y (n_6202));
CLKBUFX1 gbuf_d_557(.A(n_3217), .Y(d_out_557));
CLKBUFX1 gbuf_qn_557(.A(qn_in_557), .Y(WX8305));
NOR2X1 g57059(.A (WX6952), .B (n_5838), .Y (n_3639));
CLKBUFX1 gbuf_d_558(.A(n_3210), .Y(d_out_558));
CLKBUFX1 gbuf_q_558(.A(q_in_558), .Y(_2152_));
CLKBUFX1 gbuf_d_559(.A(n_3216), .Y(d_out_559));
CLKBUFX1 gbuf_qn_559(.A(qn_in_559), .Y(WX9598));
CLKBUFX1 gbuf_d_560(.A(n_3204), .Y(d_out_560));
CLKBUFX1 gbuf_q_560(.A(q_in_560), .Y(_2189_));
NOR2X1 g57163(.A (WX9538), .B (n_5811), .Y (n_6203));
NAND2X1 g58512(.A (n_3410), .B (n_2511), .Y (n_3637));
NAND2X1 g58517(.A (n_3404), .B (n_2453), .Y (n_3633));
NAND2X1 g58521(.A (n_3395), .B (n_2498), .Y (n_3632));
NAND2X1 g58530(.A (n_3382), .B (n_2494), .Y (n_3628));
NAND2X1 g58532(.A (n_3361), .B (n_2472), .Y (n_3626));
NAND2X1 g58540(.A (n_3346), .B (n_2466), .Y (n_3622));
NAND2X1 g58543(.A (n_3364), .B (n_2446), .Y (n_3621));
NAND2X1 g58544(.A (n_3337), .B (n_2468), .Y (n_3620));
NAND2X1 g58551(.A (n_3320), .B (n_2458), .Y (n_3616));
NAND2X1 g58555(.A (n_3306), .B (n_2443), .Y (n_3614));
NAND2X1 g58561(.A (n_3308), .B (n_2437), .Y (n_3612));
NAND2X1 g58567(.A (n_3261), .B (n_2422), .Y (n_3609));
NOR2X1 g58572(.A (n_3181), .B (n_3690), .Y (n_3606));
NOR2X1 g58573(.A (n_3180), .B (n_5712), .Y (n_3605));
NOR2X1 g58574(.A (n_3179), .B (n_1648), .Y (n_3604));
AND2X1 g61727(.A (WX9556), .B (n_5873), .Y (n_6661));
AND2X1 g62334(.A (WX8265), .B (n_5873), .Y (n_3601));
OR2X1 g62530(.A (n_3599), .B (n_5990), .Y (n_3600));
XOR2X1 g58924(.A (WX4604), .B (n_3157), .Y (n_3598));
XOR2X1 g58927(.A (WX5921), .B (n_2930), .Y (n_3597));
XOR2X1 g58930(.A (WX4606), .B (n_3055), .Y (n_3596));
XOR2X1 g58931(.A (WX8525), .B (n_3155), .Y (n_3595));
XOR2X1 g58932(.A (WX4608), .B (n_3153), .Y (n_3594));
XOR2X1 g58933(.A (WX8527), .B (n_3154), .Y (n_3593));
XOR2X1 g58934(.A (WX8529), .B (n_3152), .Y (n_3592));
XOR2X1 g58935(.A (WX4610), .B (n_3151), .Y (n_3591));
XOR2X1 g58939(.A (WX4614), .B (n_3147), .Y (n_3589));
XOR2X1 g58940(.A (WX4616), .B (n_3145), .Y (n_3588));
XOR2X1 g58941(.A (WX4618), .B (n_3156), .Y (n_3587));
XOR2X1 g58944(.A (WX4620), .B (n_3142), .Y (n_3586));
XOR2X1 g58946(.A (WX4624), .B (n_3139), .Y (n_3585));
XOR2X1 g58948(.A (WX9762), .B (n_3138), .Y (n_3584));
XOR2X1 g58950(.A (WX9764), .B (n_3135), .Y (n_3583));
XOR2X1 g58951(.A (WX9766), .B (n_3134), .Y (n_3582));
XOR2X1 g58954(.A (WX9770), .B (n_3131), .Y (n_3581));
XOR2X1 g58956(.A (WX9772), .B (n_3127), .Y (n_3580));
XOR2X1 g58957(.A (WX9774), .B (n_3096), .Y (n_3579));
XOR2X1 g58959(.A (WX9776), .B (n_3125), .Y (n_3578));
XOR2X1 g58962(.A (WX9778), .B (n_2943), .Y (n_3577));
XOR2X1 g58964(.A (WX9780), .B (n_2972), .Y (n_3576));
XOR2X1 g58965(.A (WX9782), .B (n_3001), .Y (n_3575));
XOR2X1 g58967(.A (WX3295), .B (n_3123), .Y (n_3574));
XOR2X1 g58968(.A (WX9784), .B (n_3017), .Y (n_3573));
XOR2X1 g58969(.A (WX9786), .B (n_3121), .Y (n_3572));
XOR2X1 g58972(.A (WX4638), .B (n_3057), .Y (n_3571));
XOR2X1 g58974(.A (WX9790), .B (n_3118), .Y (n_3570));
XOR2X1 g58976(.A (WX9792), .B (n_3117), .Y (n_3569));
XOR2X1 g58977(.A (WX9794), .B (n_3126), .Y (n_3568));
XOR2X1 g58978(.A (WX4642), .B (n_3116), .Y (n_3567));
XOR2X1 g58980(.A (WX9796), .B (n_2954), .Y (n_3566));
XOR2X1 g58983(.A (WX9800), .B (n_2936), .Y (n_3565));
XOR2X1 g58985(.A (WX4646), .B (n_3113), .Y (n_3564));
XOR2X1 g58998(.A (WX9814), .B (n_3107), .Y (n_3563));
CLKBUFX1 gbuf_d_561(.A(n_3215), .Y(d_out_561));
CLKBUFX1 gbuf_q_561(.A(q_in_561), .Y(_2113_));
XOR2X1 g59000(.A (WX9816), .B (n_3104), .Y (n_3562));
XOR2X1 g59002(.A (WX9820), .B (n_3101), .Y (n_3561));
XOR2X1 g59004(.A (WX3301), .B (n_3099), .Y (n_3560));
XOR2X1 g59005(.A (WX11057), .B (n_3098), .Y (n_3559));
XOR2X1 g59012(.A (WX11059), .B (n_3095), .Y (n_3558));
XOR2X1 g59013(.A (WX3303), .B (n_3093), .Y (n_3557));
XOR2X1 g59014(.A (WX3305), .B (n_3092), .Y (n_3556));
XOR2X1 g59016(.A (WX11061), .B (n_3085), .Y (n_3555));
XOR2X1 g59017(.A (WX5883), .B (n_3087), .Y (n_3554));
XOR2X1 g59018(.A (WX5885), .B (n_2957), .Y (n_3553));
XOR2X1 g59019(.A (WX3307), .B (n_2969), .Y (n_3552));
XOR2X1 g59020(.A (WX11071), .B (n_3111), .Y (n_3551));
XOR2X1 g59023(.A (WX5887), .B (n_3083), .Y (n_3550));
XOR2X1 g59025(.A (WX5889), .B (n_3081), .Y (n_3549));
XOR2X1 g59026(.A (WX5891), .B (n_3022), .Y (n_3548));
XOR2X1 g59027(.A (WX11063), .B (n_2955), .Y (n_3547));
XOR2X1 g59029(.A (WX5893), .B (n_3080), .Y (n_3546));
XOR2X1 g59030(.A (WX3309), .B (n_3043), .Y (n_3545));
XOR2X1 g59033(.A (WX5895), .B (n_3076), .Y (n_3544));
XOR2X1 g59034(.A (WX5897), .B (n_3075), .Y (n_3543));
XOR2X1 g59038(.A (WX5899), .B (n_3029), .Y (n_3542));
XOR2X1 g59039(.A (WX11065), .B (n_2958), .Y (n_3541));
XOR2X1 g59040(.A (WX5901), .B (n_3015), .Y (n_3540));
XOR2X1 g59041(.A (WX3311), .B (n_3074), .Y (n_3539));
XOR2X1 g59046(.A (WX4650), .B (n_3110), .Y (n_3538));
XOR2X1 g59048(.A (WX5905), .B (n_3071), .Y (n_3537));
XOR2X1 g59049(.A (WX5907), .B (n_3069), .Y (n_3536));
XOR2X1 g59050(.A (WX11067), .B (n_3088), .Y (n_3535));
XOR2X1 g59052(.A (WX5911), .B (n_3114), .Y (n_3534));
XOR2X1 g59053(.A (WX5913), .B (n_3128), .Y (n_3533));
XOR2X1 g59058(.A (WX11069), .B (n_3064), .Y (n_3532));
XOR2X1 g59062(.A (WX3317), .B (n_3052), .Y (n_3531));
XOR2X1 g59065(.A (WX5925), .B (n_3062), .Y (n_3530));
XOR2X1 g59066(.A (WX5927), .B (n_3090), .Y (n_3529));
XOR2X1 g59072(.A (WX11073), .B (n_3054), .Y (n_3527));
XOR2X1 g59078(.A (WX3323), .B (n_3051), .Y (n_3526));
XOR2X1 g59079(.A (WX5939), .B (n_3115), .Y (n_3525));
XOR2X1 g59082(.A (WX5941), .B (n_3066), .Y (n_3524));
XOR2X1 g59083(.A (WX11075), .B (n_3049), .Y (n_3523));
XOR2X1 g59087(.A (WX5943), .B (n_3102), .Y (n_3522));
XOR2X1 g59089(.A (WX3325), .B (n_3039), .Y (n_3521));
XOR2X1 g59090(.A (WX11077), .B (n_3065), .Y (n_3520));
XOR2X1 g59092(.A (WX11079), .B (n_3047), .Y (n_3519));
XOR2X1 g59096(.A (WX3329), .B (n_3045), .Y (n_3518));
XOR2X1 g59099(.A (WX3331), .B (n_3037), .Y (n_3517));
XOR2X1 g59100(.A (WX7174), .B (n_3038), .Y (n_3516));
XOR2X1 g59105(.A (WX7178), .B (n_3032), .Y (n_3514));
XOR2X1 g59106(.A (WX7180), .B (n_3030), .Y (n_3513));
XOR2X1 g59108(.A (WX11083), .B (n_3028), .Y (n_3512));
XOR2X1 g59109(.A (WX7182), .B (n_3026), .Y (n_3511));
XOR2X1 g59110(.A (WX7184), .B (n_3024), .Y (n_3510));
XOR2X1 g59112(.A (WX7186), .B (n_3023), .Y (n_3509));
XOR2X1 g59114(.A (WX7188), .B (n_3020), .Y (n_3508));
XOR2X1 g59116(.A (WX7190), .B (n_3018), .Y (n_3507));
XOR2X1 g59118(.A (WX7192), .B (n_3014), .Y (n_3506));
XOR2X1 g59121(.A (WX7194), .B (n_3012), .Y (n_3505));
XOR2X1 g59122(.A (WX3337), .B (n_3011), .Y (n_3504));
XOR2X1 g59125(.A (WX7196), .B (n_3009), .Y (n_3503));
XOR2X1 g59126(.A (WX3339), .B (n_3007), .Y (n_3502));
XOR2X1 g59127(.A (WX5881), .B (n_3077), .Y (n_3501));
XOR2X1 g59128(.A (WX7198), .B (n_3003), .Y (n_3500));
XOR2X1 g59129(.A (WX7200), .B (n_3000), .Y (n_3499));
XOR2X1 g59131(.A (WX11087), .B (n_3005), .Y (n_3498));
XOR2X1 g59132(.A (WX7202), .B (n_2999), .Y (n_3497));
XOR2X1 g59134(.A (WX7204), .B (n_3040), .Y (n_3496));
XOR2X1 g59135(.A (WX7206), .B (n_2997), .Y (n_3495));
XOR2X1 g59138(.A (WX7208), .B (n_2995), .Y (n_3494));
XOR2X1 g59139(.A (WX7210), .B (n_2994), .Y (n_3493));
XOR2X1 g59140(.A (WX4648), .B (n_2998), .Y (n_3492));
XOR2X1 g59142(.A (WX7212), .B (n_2992), .Y (n_3491));
XOR2X1 g59144(.A (WX7214), .B (n_2991), .Y (n_3490));
XOR2X1 g59149(.A (WX7220), .B (n_2990), .Y (n_3489));
XOR2X1 g59150(.A (WX3345), .B (n_2987), .Y (n_3488));
XOR2X1 g59151(.A (WX7222), .B (n_2985), .Y (n_3487));
XOR2X1 g59152(.A (WX11093), .B (n_2984), .Y (n_3486));
XOR2X1 g59157(.A (WX7226), .B (n_2981), .Y (n_3485));
XOR2X1 g59162(.A (WX7230), .B (n_2979), .Y (n_3484));
XOR2X1 g59163(.A (WX11095), .B (n_2975), .Y (n_3483));
XOR2X1 g59164(.A (WX3349), .B (n_2978), .Y (n_3482));
XOR2X1 g59170(.A (WX7236), .B (n_2974), .Y (n_3481));
XOR2X1 g59172(.A (WX11097), .B (n_2971), .Y (n_3480));
XOR2X1 g59176(.A (WX11099), .B (n_3048), .Y (n_3479));
XOR2X1 g59182(.A (WX11101), .B (n_2968), .Y (n_3478));
XOR2X1 g59183(.A (WX3357), .B (n_2967), .Y (n_3477));
XOR2X1 g59185(.A (WX11103), .B (n_2966), .Y (n_3476));
XOR2X1 g59186(.A (WX5909), .B (n_3141), .Y (n_3475));
XOR2X1 g59188(.A (WX5929), .B (n_3059), .Y (n_3474));
XOR2X1 g59193(.A (WX8469), .B (n_2965), .Y (n_3472));
XOR2X1 g59194(.A (WX8471), .B (n_2963), .Y (n_3471));
XOR2X1 g59197(.A (WX8473), .B (n_2961), .Y (n_3470));
XOR2X1 g59198(.A (WX11109), .B (n_3108), .Y (n_3469));
XOR2X1 g59199(.A (WX8475), .B (n_2960), .Y (n_3468));
XOR2X1 g59201(.A (WX8477), .B (n_3136), .Y (n_3467));
XOR2X1 g59206(.A (WX8485), .B (n_2952), .Y (n_3466));
XOR2X1 g59209(.A (WX8487), .B (n_2950), .Y (n_3465));
XOR2X1 g59211(.A (WX8489), .B (n_2949), .Y (n_3464));
XOR2X1 g59215(.A (WX8491), .B (n_3061), .Y (n_3463));
XOR2X1 g59216(.A (WX4590), .B (n_2948), .Y (n_3462));
XOR2X1 g59217(.A (WX8493), .B (n_2947), .Y (n_3461));
XOR2X1 g59220(.A (WX8495), .B (n_2946), .Y (n_3460));
XOR2X1 g59221(.A (WX4592), .B (n_2944), .Y (n_3459));
XOR2X1 g59222(.A (WX8497), .B (n_3068), .Y (n_3458));
XOR2X1 g59224(.A (WX4594), .B (n_2941), .Y (n_3457));
XOR2X1 g59226(.A (WX8501), .B (n_2940), .Y (n_3456));
XOR2X1 g59227(.A (WX4596), .B (n_2939), .Y (n_3455));
XOR2X1 g59229(.A (WX8505), .B (n_2937), .Y (n_3454));
XOR2X1 g59231(.A (WX4598), .B (n_2934), .Y (n_3453));
XOR2X1 g59232(.A (WX8509), .B (n_2933), .Y (n_3452));
XOR2X1 g59234(.A (WX4600), .B (n_2932), .Y (n_3451));
XOR2X1 g59235(.A (WX8513), .B (n_2982), .Y (n_3450));
XOR2X1 g59237(.A (WX4602), .B (n_2931), .Y (n_3449));
CLKBUFX1 gbuf_d_562(.A(n_3200), .Y(d_out_562));
CLKBUFX1 gbuf_q_562(.A(q_in_562), .Y(_2241_));
NOR2X1 g59499(.A (WX3099), .B (n_5500), .Y (n_3447));
NOR2X1 g59502(.A (WX8263), .B (n_5500), .Y (n_6663));
NOR2X1 g59508(.A (WX9554), .B (n_5811), .Y (n_6204));
NOR2X1 g59509(.A (WX5681), .B (n_5811), .Y (n_6206));
CLKBUFX1 gbuf_d_563(.A(n_3167), .Y(d_out_563));
CLKBUFX1 gbuf_qn_563(.A(qn_in_563), .Y(WX3133));
CLKBUFX1 gbuf_d_564(.A(n_3177), .Y(d_out_564));
CLKBUFX1 gbuf_q_564(.A(q_in_564), .Y(WX485));
CLKBUFX1 gbuf_d_565(.A(n_3190), .Y(d_out_565));
CLKBUFX1 gbuf_q_565(.A(q_in_565), .Y(_2317_));
CLKBUFX1 gbuf_d_566(.A(n_3213), .Y(d_out_566));
CLKBUFX1 gbuf_q_566(.A(q_in_566), .Y(_2120_));
CLKBUFX1 gbuf_d_567(.A(n_3212), .Y(d_out_567));
CLKBUFX1 gbuf_q_567(.A(q_in_567), .Y(_2125_));
CLKBUFX1 gbuf_d_568(.A(n_3211), .Y(d_out_568));
CLKBUFX1 gbuf_q_568(.A(q_in_568), .Y(_2145_));
CLKBUFX1 gbuf_d_569(.A(n_3208), .Y(d_out_569));
CLKBUFX1 gbuf_q_569(.A(q_in_569), .Y(_2157_));
CLKBUFX1 gbuf_d_570(.A(n_3207), .Y(d_out_570));
CLKBUFX1 gbuf_q_570(.A(q_in_570), .Y(_2177_));
CLKBUFX1 gbuf_d_571(.A(n_3205), .Y(d_out_571));
CLKBUFX1 gbuf_q_571(.A(q_in_571), .Y(_2184_));
CLKBUFX1 gbuf_d_572(.A(n_3203), .Y(d_out_572));
CLKBUFX1 gbuf_q_572(.A(q_in_572), .Y(_2209_));
CLKBUFX1 gbuf_d_573(.A(n_3202), .Y(d_out_573));
CLKBUFX1 gbuf_q_573(.A(q_in_573), .Y(_2216_));
CLKBUFX1 gbuf_d_574(.A(n_3201), .Y(d_out_574));
CLKBUFX1 gbuf_q_574(.A(q_in_574), .Y(_2221_));
CLKBUFX1 gbuf_d_575(.A(n_3199), .Y(d_out_575));
CLKBUFX1 gbuf_q_575(.A(q_in_575), .Y(_2248_));
CLKBUFX1 gbuf_d_576(.A(n_3197), .Y(d_out_576));
CLKBUFX1 gbuf_q_576(.A(q_in_576), .Y(_2273_));
CLKBUFX1 gbuf_d_577(.A(n_3194), .Y(d_out_577));
CLKBUFX1 gbuf_q_577(.A(q_in_577), .Y(_2285_));
CLKBUFX1 gbuf_d_578(.A(n_3192), .Y(d_out_578));
CLKBUFX1 gbuf_q_578(.A(q_in_578), .Y(_2305_));
CLKBUFX1 gbuf_d_579(.A(n_3191), .Y(d_out_579));
CLKBUFX1 gbuf_q_579(.A(q_in_579), .Y(_2312_));
CLKBUFX1 gbuf_d_580(.A(n_3189), .Y(d_out_580));
CLKBUFX1 gbuf_q_580(.A(q_in_580), .Y(_2337_));
CLKBUFX1 gbuf_d_581(.A(n_3187), .Y(d_out_581));
CLKBUFX1 gbuf_q_581(.A(q_in_581), .Y(_2344_));
CLKBUFX1 gbuf_d_582(.A(n_3186), .Y(d_out_582));
CLKBUFX1 gbuf_q_582(.A(q_in_582), .Y(_2349_));
CLKBUFX1 gbuf_d_583(.A(n_3198), .Y(d_out_583));
CLKBUFX1 gbuf_q_583(.A(q_in_583), .Y(_2253_));
CLKBUFX1 gbuf_d_584(.A(n_3195), .Y(d_out_584));
CLKBUFX1 gbuf_q_584(.A(q_in_584), .Y(_2280_));
NOR2X1 g56885(.A (WX3073), .B (n_5427), .Y (n_3443));
CLKBUFX1 gbuf_d_585(.A(n_3227), .Y(d_out_585));
CLKBUFX1 gbuf_qn_585(.A(qn_in_585), .Y(WX5719));
AND2X1 g56933(.A (WX5657), .B (n_5828), .Y (n_6212));
CLKBUFX1 gbuf_d_586(.A(n_2917), .Y(d_out_586));
CLKBUFX1 gbuf_qn_586(.A(qn_in_586), .Y(WX1840));
CLKBUFX1 gbuf_d_587(.A(n_2928), .Y(d_out_587));
CLKBUFX1 gbuf_qn_587(.A(qn_in_587), .Y(WX10891));
CLKBUFX1 gbuf_d_588(.A(n_2927), .Y(d_out_588));
CLKBUFX1 gbuf_q_588(.A(q_in_588), .Y(WX547));
AND2X1 g57000(.A (WX6950), .B (n_5828), .Y (n_6213));
CLKBUFX1 gbuf_d_589(.A(n_2843), .Y(d_out_589));
CLKBUFX1 gbuf_q_589(.A(q_in_589), .Y(_2087_));
AND2X1 g57038(.A (WX8243), .B (n_5828), .Y (n_6183));
CLKBUFX1 gbuf_d_590(.A(n_2879), .Y(d_out_590));
CLKBUFX1 gbuf_q_590(.A(q_in_590), .Y(_2085_));
AND2X1 g57103(.A (WX9536), .B (n_5828), .Y (n_3439));
CLKBUFX1 gbuf_d_591(.A(n_2881), .Y(d_out_591));
CLKBUFX1 gbuf_q_591(.A(q_in_591), .Y(_2083_));
AND2X1 g61553(.A (WX5683), .B (n_5828), .Y (n_6208));
AND2X1 g55863(.A (WX1780), .B (n_5828), .Y (n_3437));
AND2X1 g55864(.A (WX10831), .B (n_5828), .Y (n_3436));
AND2X1 g61819(.A (WX1778), .B (n_5828), .Y (n_3435));
AND2X1 g61843(.A (WX4392), .B (n_5828), .Y (n_3434));
AND2X1 g62063(.A (WX3101), .B (n_5828), .Y (n_3433));
AND2X1 g62145(.A (WX6974), .B (n_5828), .Y (n_6664));
AND2X1 g62308(.A (WX10829), .B (n_5828), .Y (n_3431));
INVX4 g62383(.A (n_3428), .Y (n_5460));
INVX4 g62393(.A (n_3428), .Y (n_5619));
INVX4 g62398(.A (n_3428), .Y (n_5556));
INVX8 g62403(.A (n_3426), .Y (n_4860));
INVX4 g62439(.A (n_3421), .Y (n_5566));
INVX8 g62441(.A (n_3421), .Y (n_4947));
INVX8 g62445(.A (n_7088), .Y (n_5722));
INVX1 g62449(.A (n_7088), .Y (n_5706));
INVX1 g62452(.A (n_7088), .Y (n_5275));
XOR2X1 g58920(.A (WX2002), .B (n_2811), .Y (n_3414));
INVX1 g58925(.A (n_3410), .Y (n_3411));
XOR2X1 g58928(.A (WX8521), .B (n_2839), .Y (n_3409));
XOR2X1 g58929(.A (WX8523), .B (n_2836), .Y (n_3408));
CLKBUFX1 gbuf_d_592(.A(n_2887), .Y(d_out_592));
CLKBUFX1 gbuf_q_592(.A(q_in_592), .Y(_2077_));
INVX1 g58942(.A (n_3404), .Y (n_3405));
XOR2X1 g58945(.A (WX4622), .B (n_2835), .Y (n_3403));
XOR2X1 g58947(.A (WX9760), .B (n_2831), .Y (n_3402));
XOR2X1 g58949(.A (WX4626), .B (n_2830), .Y (n_3401));
XOR2X1 g58952(.A (WX4628), .B (n_2824), .Y (n_3400));
XOR2X1 g58953(.A (WX9768), .B (n_2823), .Y (n_3399));
XOR2X1 g58955(.A (WX4630), .B (n_2820), .Y (n_3398));
XOR2X1 g58958(.A (WX4632), .B (n_2818), .Y (n_3397));
INVX1 g58960(.A (n_3395), .Y (n_3396));
XOR2X1 g58963(.A (WX4634), .B (n_2816), .Y (n_3394));
XOR2X1 g58966(.A (WX4636), .B (n_2814), .Y (n_3393));
XOR2X1 g58973(.A (WX9788), .B (n_2812), .Y (n_3390));
XOR2X1 g58975(.A (WX4640), .B (n_2810), .Y (n_3389));
XOR2X1 g58979(.A (WX2004), .B (n_2807), .Y (n_3388));
XOR2X1 g58981(.A (WX9798), .B (n_2699), .Y (n_3387));
XOR2X1 g58982(.A (WX4644), .B (n_2711), .Y (n_3386));
XOR2X1 g58984(.A (WX3297), .B (n_2709), .Y (n_3385));
XOR2X1 g58986(.A (WX9804), .B (n_2806), .Y (n_3384));
INVX1 g58987(.A (n_3382), .Y (n_3383));
XOR2X1 g58991(.A (WX9806), .B (n_2805), .Y (n_3379));
XOR2X1 g58992(.A (WX11055), .B (n_2801), .Y (n_3378));
XOR2X1 g58993(.A (WX2022), .B (n_2773), .Y (n_3377));
XOR2X1 g58994(.A (WX9808), .B (n_2749), .Y (n_3376));
XOR2X1 g58995(.A (WX3299), .B (n_2794), .Y (n_3375));
XOR2X1 g58996(.A (WX9810), .B (n_2797), .Y (n_3374));
XOR2X1 g58997(.A (WX9812), .B (n_2793), .Y (n_3373));
XOR2X1 g58999(.A (WX2006), .B (n_2803), .Y (n_3372));
XOR2X1 g59001(.A (WX9818), .B (n_2792), .Y (n_3371));
XOR2X1 g59003(.A (WX9822), .B (n_2694), .Y (n_3370));
XOR2X1 g59006(.A (WX2008), .B (n_2726), .Y (n_3369));
XOR2X1 g59009(.A (WX2010), .B (n_2786), .Y (n_3366));
INVX1 g59010(.A (n_3364), .Y (n_3365));
XOR2X1 g59015(.A (WX2012), .B (n_2791), .Y (n_3363));
INVX1 g59021(.A (n_3361), .Y (n_3362));
XOR2X1 g59024(.A (WX2014), .B (n_2789), .Y (n_3360));
XOR2X1 g59028(.A (WX2016), .B (n_2787), .Y (n_3359));
XOR2X1 g59035(.A (WX2018), .B (n_2714), .Y (n_3356));
XOR2X1 g59042(.A (WX5933), .B (n_2777), .Y (n_3353));
XOR2X1 g59043(.A (WX5903), .B (n_2784), .Y (n_3352));
XOR2X1 g59047(.A (WX2020), .B (n_2700), .Y (n_3349));
XOR2X1 g59051(.A (WX3313), .B (n_2783), .Y (n_3348));
INVX1 g59054(.A (n_3346), .Y (n_3347));
XOR2X1 g59056(.A (WX3315), .B (n_2763), .Y (n_3345));
XOR2X1 g59057(.A (WX5915), .B (n_2769), .Y (n_3344));
XOR2X1 g59059(.A (WX5917), .B (n_2799), .Y (n_3343));
XOR2X1 g59060(.A (WX2024), .B (n_2703), .Y (n_3342));
XOR2X1 g59061(.A (WX5919), .B (n_2822), .Y (n_3341));
XOR2X1 g59063(.A (WX5923), .B (n_2780), .Y (n_3340));
XOR2X1 g59064(.A (WX2026), .B (n_2778), .Y (n_3339));
INVX1 g59067(.A (n_3337), .Y (n_3338));
XOR2X1 g59070(.A (WX5931), .B (n_2771), .Y (n_3336));
XOR2X1 g59071(.A (WX3321), .B (n_2695), .Y (n_3335));
XOR2X1 g59073(.A (WX2028), .B (n_2768), .Y (n_3334));
XOR2X1 g59074(.A (WX5935), .B (n_2790), .Y (n_3333));
XOR2X1 g59077(.A (WX5937), .B (n_2765), .Y (n_3330));
XOR2X1 g59084(.A (WX2030), .B (n_2774), .Y (n_3327));
XOR2X1 g59088(.A (WX2032), .B (n_2827), .Y (n_3324));
XOR2X1 g59091(.A (WX3327), .B (n_2833), .Y (n_3323));
XOR2X1 g59093(.A (WX2036), .B (n_2788), .Y (n_3322));
INVX1 g59094(.A (n_3320), .Y (n_3321));
XOR2X1 g59097(.A (WX2038), .B (n_2767), .Y (n_3319));
XOR2X1 g59098(.A (WX11081), .B (n_2762), .Y (n_3318));
XOR2X1 g59104(.A (WX3333), .B (n_2761), .Y (n_3315));
XOR2X1 g59107(.A (WX2040), .B (n_2759), .Y (n_3314));
XOR2X1 g59111(.A (WX3335), .B (n_2756), .Y (n_3313));
XOR2X1 g59113(.A (WX2042), .B (n_2754), .Y (n_3312));
XOR2X1 g59115(.A (WX11085), .B (n_2752), .Y (n_3311));
XOR2X1 g59117(.A (WX2044), .B (n_2750), .Y (n_3310));
INVX1 g59119(.A (n_3308), .Y (n_3309));
INVX1 g59123(.A (n_3306), .Y (n_3307));
XOR2X1 g59130(.A (WX2046), .B (n_2745), .Y (n_3305));
XOR2X1 g59133(.A (WX2048), .B (n_2743), .Y (n_3304));
XOR2X1 g59136(.A (WX11089), .B (n_2742), .Y (n_3303));
XOR2X1 g59137(.A (WX3341), .B (n_2741), .Y (n_3302));
XOR2X1 g59141(.A (WX3343), .B (n_2738), .Y (n_3301));
XOR2X1 g59143(.A (WX2050), .B (n_2737), .Y (n_3300));
XOR2X1 g59145(.A (WX11091), .B (n_2736), .Y (n_3299));
XOR2X1 g59147(.A (WX2052), .B (n_2733), .Y (n_3297));
XOR2X1 g59148(.A (WX7218), .B (n_2732), .Y (n_3296));
XOR2X1 g59155(.A (WX2054), .B (n_2731), .Y (n_3293));
XOR2X1 g59156(.A (WX7224), .B (n_2730), .Y (n_3292));
XOR2X1 g59158(.A (WX3347), .B (n_2729), .Y (n_3291));
XOR2X1 g59159(.A (WX7228), .B (n_2728), .Y (n_3290));
XOR2X1 g59165(.A (WX7232), .B (n_2725), .Y (n_3287));
XOR2X1 g59166(.A (WX2056), .B (n_2724), .Y (n_3286));
XOR2X1 g59167(.A (WX7234), .B (n_2722), .Y (n_3285));
XOR2X1 g59171(.A (WX2058), .B (n_2721), .Y (n_3282));
XOR2X1 g59173(.A (WX3351), .B (n_2720), .Y (n_3281));
XOR2X1 g59174(.A (WX3353), .B (n_2719), .Y (n_3280));
INVX2 g63085(.A (n_5873), .Y (n_5822));
XOR2X1 g59175(.A (WX2060), .B (n_2718), .Y (n_3278));
INVX2 g63101(.A (n_4150), .Y (n_5052));
INVX4 g63107(.A (n_3221), .Y (n_5968));
XOR2X1 g59177(.A (WX2062), .B (n_2772), .Y (n_3276));
XOR2X1 g59180(.A (WX3355), .B (n_2717), .Y (n_3273));
XOR2X1 g59181(.A (WX2034), .B (n_2782), .Y (n_3272));
INVX8 g63165(.A (n_6440), .Y (n_4882));
INVX4 g63172(.A (n_3269), .Y (n_3828));
XOR2X1 g59184(.A (WX2064), .B (n_2715), .Y (n_3268));
INVX8 g63194(.A (n_3264), .Y (n_5662));
XOR2X1 g59187(.A (WX11105), .B (n_2713), .Y (n_3265));
INVX8 g63212(.A (n_3263), .Y (n_5479));
INVX1 g59189(.A (n_3261), .Y (n_3262));
XOR2X1 g59191(.A (WX11107), .B (n_2710), .Y (n_3260));
XOR2X1 g59200(.A (WX9802), .B (n_2708), .Y (n_3257));
XOR2X1 g59202(.A (WX8479), .B (n_2707), .Y (n_3256));
XOR2X1 g59203(.A (WX8481), .B (n_2706), .Y (n_3255));
XOR2X1 g59204(.A (WX11111), .B (n_2705), .Y (n_3254));
XOR2X1 g59205(.A (WX8483), .B (n_2704), .Y (n_3253));
XOR2X1 g59210(.A (WX4588), .B (n_2702), .Y (n_3250));
XOR2X1 g59212(.A (WX11113), .B (n_2701), .Y (n_3249));
XOR2X1 g59223(.A (WX11115), .B (n_2698), .Y (n_3244));
XOR2X1 g59225(.A (WX8499), .B (n_2697), .Y (n_3243));
XOR2X1 g59228(.A (WX8503), .B (n_2696), .Y (n_3242));
XOR2X1 g59230(.A (WX8507), .B (n_2712), .Y (n_3241));
XOR2X1 g59233(.A (WX8511), .B (n_2734), .Y (n_3240));
XOR2X1 g59236(.A (WX8515), .B (n_2739), .Y (n_3239));
XOR2X1 g59238(.A (WX8517), .B (n_2746), .Y (n_3238));
XOR2X1 g59239(.A (WX8519), .B (n_2760), .Y (n_3237));
NOR2X1 g59501(.A (WX8263), .B (n_5712), .Y (n_3236));
NOR2X1 g59504(.A (WX9554), .B (n_1648), .Y (n_3235));
NOR2X1 g59505(.A (WX4390), .B (n_3188), .Y (n_3234));
NOR2X1 g59507(.A (WX5681), .B (n_5712), .Y (n_3233));
NOR2X1 g59513(.A (WX6972), .B (n_5712), .Y (n_3231));
NOR2X1 g59516(.A (WX3099), .B (n_3188), .Y (n_3230));
CLKBUFX1 gbuf_d_593(.A(n_2872), .Y(d_out_593));
CLKBUFX1 gbuf_q_593(.A(q_in_593), .Y(_2094_));
CLKBUFX1 gbuf_d_594(.A(n_2868), .Y(d_out_594));
CLKBUFX1 gbuf_q_594(.A(q_in_594), .Y(_2099_));
CLKBUFX1 gbuf_d_595(.A(n_2846), .Y(d_out_595));
CLKBUFX1 gbuf_q_595(.A(q_in_595), .Y(_2103_));
CLKBUFX1 gbuf_d_596(.A(n_2898), .Y(d_out_596));
CLKBUFX1 gbuf_q_596(.A(q_in_596), .Y(_2108_));
CLKBUFX1 gbuf_d_597(.A(n_2861), .Y(d_out_597));
CLKBUFX1 gbuf_q_597(.A(q_in_597), .Y(_2118_));
CLKBUFX1 gbuf_d_598(.A(n_2883), .Y(d_out_598));
CLKBUFX1 gbuf_q_598(.A(q_in_598), .Y(_2080_));
CLKBUFX1 gbuf_d_599(.A(n_2885), .Y(d_out_599));
CLKBUFX1 gbuf_q_599(.A(q_in_599), .Y(_2078_));
CLKBUFX1 gbuf_d_600(.A(n_2884), .Y(d_out_600));
CLKBUFX1 gbuf_q_600(.A(q_in_600), .Y(_2079_));
CLKBUFX1 gbuf_d_601(.A(n_2882), .Y(d_out_601));
CLKBUFX1 gbuf_q_601(.A(q_in_601), .Y(_2082_));
CLKBUFX1 gbuf_d_602(.A(n_2850), .Y(d_out_602));
CLKBUFX1 gbuf_q_602(.A(q_in_602), .Y(_2084_));
CLKBUFX1 gbuf_d_603(.A(n_2878), .Y(d_out_603));
CLKBUFX1 gbuf_q_603(.A(q_in_603), .Y(_2086_));
CLKBUFX1 gbuf_d_604(.A(n_2875), .Y(d_out_604));
CLKBUFX1 gbuf_q_604(.A(q_in_604), .Y(_2090_));
CLKBUFX1 gbuf_d_605(.A(n_2852), .Y(d_out_605));
CLKBUFX1 gbuf_q_605(.A(q_in_605), .Y(_2091_));
CLKBUFX1 gbuf_d_606(.A(n_2873), .Y(d_out_606));
CLKBUFX1 gbuf_q_606(.A(q_in_606), .Y(_2092_));
CLKBUFX1 gbuf_d_607(.A(n_2870), .Y(d_out_607));
CLKBUFX1 gbuf_q_607(.A(q_in_607), .Y(_2095_));
CLKBUFX1 gbuf_d_608(.A(n_2844), .Y(d_out_608));
CLKBUFX1 gbuf_q_608(.A(q_in_608), .Y(_2096_));
CLKBUFX1 gbuf_d_609(.A(n_2893), .Y(d_out_609));
CLKBUFX1 gbuf_q_609(.A(q_in_609), .Y(_2098_));
CLKBUFX1 gbuf_d_610(.A(n_2856), .Y(d_out_610));
CLKBUFX1 gbuf_q_610(.A(q_in_610), .Y(_2100_));
CLKBUFX1 gbuf_d_611(.A(n_2867), .Y(d_out_611));
CLKBUFX1 gbuf_q_611(.A(q_in_611), .Y(_2101_));
CLKBUFX1 gbuf_d_612(.A(n_2854), .Y(d_out_612));
CLKBUFX1 gbuf_q_612(.A(q_in_612), .Y(_2102_));
CLKBUFX1 gbuf_d_613(.A(n_2866), .Y(d_out_613));
CLKBUFX1 gbuf_q_613(.A(q_in_613), .Y(_2104_));
CLKBUFX1 gbuf_d_614(.A(n_2865), .Y(d_out_614));
CLKBUFX1 gbuf_q_614(.A(q_in_614), .Y(_2105_));
CLKBUFX1 gbuf_d_615(.A(n_2864), .Y(d_out_615));
CLKBUFX1 gbuf_q_615(.A(q_in_615), .Y(_2106_));
CLKBUFX1 gbuf_d_616(.A(n_2889), .Y(d_out_616));
CLKBUFX1 gbuf_q_616(.A(q_in_616), .Y(_2131_));
AND2X1 g56826(.A (WX3071), .B (n_5828), .Y (n_6182));
CLKBUFX1 gbuf_d_617(.A(n_2860), .Y(d_out_617));
CLKBUFX1 gbuf_q_617(.A(q_in_617), .Y(_2183_));
CLKBUFX1 gbuf_d_618(.A(n_2859), .Y(d_out_618));
CLKBUFX1 gbuf_q_618(.A(q_in_618), .Y(_2185_));
CLKBUFX1 gbuf_d_619(.A(n_2892), .Y(d_out_619));
CLKBUFX1 gbuf_q_619(.A(q_in_619), .Y(_2198_));
CLKBUFX1 gbuf_d_620(.A(n_2858), .Y(d_out_620));
CLKBUFX1 gbuf_q_620(.A(q_in_620), .Y(_2271_));
CLKBUFX1 gbuf_d_621(.A(n_2857), .Y(d_out_621));
CLKBUFX1 gbuf_q_621(.A(q_in_621), .Y(_2272_));
CLKBUFX1 gbuf_d_622(.A(n_2847), .Y(d_out_622));
CLKBUFX1 gbuf_q_622(.A(q_in_622), .Y(_2331_));
CLKBUFX1 gbuf_d_623(.A(n_2848), .Y(d_out_623));
CLKBUFX1 gbuf_q_623(.A(q_in_623), .Y(_2362_));
CLKBUFX1 gbuf_d_624(.A(n_2855), .Y(d_out_624));
CLKBUFX1 gbuf_q_624(.A(q_in_624), .Y(_2097_));
CLKBUFX1 gbuf_d_625(.A(n_2876), .Y(d_out_625));
CLKBUFX1 gbuf_q_625(.A(q_in_625), .Y(_2089_));
CLKBUFX1 gbuf_d_626(.A(n_2863), .Y(d_out_626));
CLKBUFX1 gbuf_q_626(.A(q_in_626), .Y(_2107_));
CLKBUFX1 gbuf_d_627(.A(n_2907), .Y(d_out_627));
CLKBUFX1 gbuf_q_627(.A(q_in_627), .Y(WX721));
CLKBUFX1 gbuf_d_628(.A(n_2914), .Y(d_out_628));
CLKBUFX1 gbuf_q_628(.A(q_in_628), .Y(WX725));
CLKBUFX1 gbuf_d_629(.A(n_2916), .Y(d_out_629));
CLKBUFX1 gbuf_q_629(.A(q_in_629), .Y(WX727));
CLKBUFX1 gbuf_d_630(.A(n_2903), .Y(d_out_630));
CLKBUFX1 gbuf_q_630(.A(q_in_630), .Y(WX745));
CLKBUFX1 gbuf_d_631(.A(n_2911), .Y(d_out_631));
CLKBUFX1 gbuf_q_631(.A(q_in_631), .Y(WX831));
CLKBUFX1 gbuf_d_632(.A(n_2909), .Y(d_out_632));
CLKBUFX1 gbuf_q_632(.A(q_in_632), .Y(WX835));
CLKBUFX1 gbuf_d_633(.A(n_2912), .Y(d_out_633));
CLKBUFX1 gbuf_q_633(.A(q_in_633), .Y(WX899));
CLKBUFX1 gbuf_d_634(.A(n_2908), .Y(d_out_634));
CLKBUFX1 gbuf_q_634(.A(q_in_634), .Y(WX845));
CLKBUFX1 gbuf_d_635(.A(n_2902), .Y(d_out_635));
CLKBUFX1 gbuf_q_635(.A(q_in_635), .Y(WX873));
CLKBUFX1 gbuf_d_636(.A(n_2906), .Y(d_out_636));
CLKBUFX1 gbuf_q_636(.A(q_in_636), .Y(WX895));
CLKBUFX1 gbuf_d_637(.A(n_2900), .Y(d_out_637));
CLKBUFX1 gbuf_q_637(.A(q_in_637), .Y(WX2032));
CLKBUFX1 gbuf_d_638(.A(n_2905), .Y(d_out_638));
CLKBUFX1 gbuf_q_638(.A(q_in_638), .Y(WX715));
CLKBUFX1 gbuf_d_639(.A(n_3163), .Y(d_out_639));
CLKBUFX1 gbuf_q_639(.A(q_in_639), .Y(WX4364));
NOR2X1 g56932(.A (WX5657), .B (n_2605), .Y (n_3227));
CLKBUFX1 gbuf_d_640(.A(n_2583), .Y(d_out_640));
CLKBUFX1 gbuf_q_640(.A(q_in_640), .Y(_2334_));
BUFX3 g63099(.A (n_3221), .Y (n_3840));
BUFX3 g63100(.A (n_3221), .Y (n_3835));
CLKBUFX3 g63103(.A (n_3221), .Y (n_4150));
BUFX3 g63094(.A (n_3221), .Y (n_4600));
BUFX3 g63092(.A (n_3221), .Y (n_4579));
BUFX3 g63093(.A (n_3221), .Y (n_4439));
BUFX3 g63090(.A (n_3221), .Y (n_4608));
NOR2X1 g56999(.A (WX6950), .B (n_2605), .Y (n_3219));
INVX4 g63058(.A (n_3831), .Y (n_3218));
NOR2X1 g57037(.A (WX8243), .B (n_2849), .Y (n_3217));
NOR2X1 g57102(.A (WX9536), .B (n_2605), .Y (n_3216));
CLKBUFX1 gbuf_d_641(.A(n_2567), .Y(d_out_641));
CLKBUFX1 gbuf_q_641(.A(q_in_641), .Y(_2308_));
NOR2X1 g58575(.A (n_2658), .B (n_5712), .Y (n_3215));
NOR2X1 g58576(.A (n_2662), .B (n_5712), .Y (n_3213));
NOR2X1 g58577(.A (n_2656), .B (n_5712), .Y (n_3212));
NOR2X1 g58578(.A (n_2655), .B (n_5181), .Y (n_3211));
NOR2X1 g58579(.A (n_2654), .B (n_1425), .Y (n_3210));
NOR2X1 g58580(.A (n_2653), .B (n_3690), .Y (n_3208));
NOR2X1 g58581(.A (n_2652), .B (n_3690), .Y (n_3207));
NOR2X1 g58582(.A (n_2661), .B (n_2851), .Y (n_3205));
NOR2X1 g58583(.A (n_2651), .B (n_2849), .Y (n_3204));
NOR2X1 g58584(.A (n_2649), .B (n_1425), .Y (n_3203));
NOR2X1 g58585(.A (n_2647), .B (n_5181), .Y (n_3202));
NOR2X1 g58586(.A (n_2646), .B (n_5712), .Y (n_3201));
NOR2X1 g58587(.A (n_2644), .B (n_5712), .Y (n_3200));
NOR2X1 g58588(.A (n_2648), .B (n_1648), .Y (n_3199));
NOR2X1 g58589(.A (n_2643), .B (n_1425), .Y (n_3198));
NOR2X1 g58590(.A (n_2642), .B (n_1648), .Y (n_3197));
NOR2X1 g58591(.A (n_2641), .B (n_1425), .Y (n_3195));
NOR2X1 g58592(.A (n_2657), .B (n_5712), .Y (n_3194));
NOR2X1 g58593(.A (n_2635), .B (n_5712), .Y (n_3192));
NOR2X1 g58594(.A (n_2640), .B (n_3188), .Y (n_3191));
NOR2X1 g58595(.A (n_2634), .B (n_1425), .Y (n_3190));
NOR2X1 g58596(.A (n_2639), .B (n_3188), .Y (n_3189));
NOR2X1 g58597(.A (n_2637), .B (n_1425), .Y (n_3187));
NOR2X1 g58598(.A (n_2636), .B (n_3188), .Y (n_3186));
INVX4 g62395(.A (n_6614), .Y (n_3428));
INVX4 g62406(.A (n_6497), .Y (n_3426));
INVX8 g62432(.A (n_3183), .Y (n_3421));
XOR2X1 g58893(.A (_2080_), .B (n_2544), .Y (n_3181));
XOR2X1 g58898(.A (_2087_), .B (n_2540), .Y (n_3180));
XOR2X1 g58899(.A (_2092_), .B (n_2537), .Y (n_3179));
XOR2X1 g58921(.A (WX11053), .B (n_2496), .Y (n_3178));
MX2X1 g58926(.A (n_18), .B (WX753), .S0 (n_2514), .Y (n_3410));
MX2X1 g58943(.A (n_19), .B (WX755), .S0 (n_2406), .Y (n_3404));
AND2X1 g55873(.A (n_2378), .B (WX487), .Y (n_3177));
MX2X1 g58961(.A (n_67), .B (WX757), .S0 (n_2500), .Y (n_3395));
MX2X1 g58988(.A (n_12), .B (WX721), .S0 (n_2487), .Y (n_3382));
MX2X1 g59011(.A (n_71), .B (WX715), .S0 (n_2471), .Y (n_3364));
MX2X1 g59022(.A (n_112), .B (WX763), .S0 (n_2477), .Y (n_3361));
MX2X1 g59055(.A (n_85), .B (WX767), .S0 (n_2470), .Y (n_3346));
MX2X1 g59068(.A (n_87), .B (WX769), .S0 (n_2480), .Y (n_3337));
MX2X1 g59095(.A (n_20), .B (WX741), .S0 (n_2462), .Y (n_3320));
MX2X1 g59120(.A (n_2), .B (WX717), .S0 (n_2445), .Y (n_3308));
MX2X1 g59124(.A (n_16), .B (WX743), .S0 (n_2448), .Y (n_3306));
INVX8 g63064(.A (n_3173), .Y (n_5889));
INVX2 g63083(.A (n_6626), .Y (n_5873));
BUFX3 g63091(.A (n_3221), .Y (n_4468));
BUFX3 g63095(.A (n_3221), .Y (n_4603));
BUFX3 g63096(.A (n_3221), .Y (n_4586));
BUFX3 g63097(.A (n_3221), .Y (n_4615));
INVX8 g63116(.A (n_3222), .Y (n_5427));
INVX8 g63127(.A (n_3223), .Y (n_5811));
INVX8 g63135(.A (n_3224), .Y (n_5500));
INVX8 g63145(.A (n_3225), .Y (n_5838));
INVX4 g63189(.A (n_3169), .Y (n_4015));
INVX4 g63213(.A (n_3168), .Y (n_3263));
MX2X1 g59190(.A (n_106), .B (WX749), .S0 (n_2424), .Y (n_3261));
CLKBUFX1 gbuf_d_642(.A(n_2585), .Y(d_out_642));
CLKBUFX1 gbuf_q_642(.A(q_in_642), .Y(_2332_));
CLKBUFX1 gbuf_d_643(.A(n_2572), .Y(d_out_643));
CLKBUFX1 gbuf_q_643(.A(q_in_643), .Y(_2363_));
CLKBUFX1 gbuf_d_644(.A(n_2587), .Y(d_out_644));
CLKBUFX1 gbuf_q_644(.A(q_in_644), .Y(_2328_));
CLKBUFX1 gbuf_d_645(.A(n_2631), .Y(d_out_645));
CLKBUFX1 gbuf_q_645(.A(q_in_645), .Y(_2140_));
CLKBUFX1 gbuf_d_646(.A(n_2678), .Y(d_out_646));
CLKBUFX1 gbuf_qn_646(.A(qn_in_646), .Y(WX11181));
CLKBUFX1 gbuf_d_647(.A(n_2571), .Y(d_out_647));
CLKBUFX1 gbuf_q_647(.A(q_in_647), .Y(_2150_));
CLKBUFX1 gbuf_d_648(.A(n_2596), .Y(d_out_648));
CLKBUFX1 gbuf_q_648(.A(q_in_648), .Y(_2293_));
CLKBUFX1 gbuf_d_649(.A(n_2621), .Y(d_out_649));
CLKBUFX1 gbuf_q_649(.A(q_in_649), .Y(_2119_));
CLKBUFX1 gbuf_d_650(.A(n_2619), .Y(d_out_650));
CLKBUFX1 gbuf_q_650(.A(q_in_650), .Y(_2121_));
CLKBUFX1 gbuf_d_651(.A(n_2629), .Y(d_out_651));
CLKBUFX1 gbuf_q_651(.A(q_in_651), .Y(_2139_));
CLKBUFX1 gbuf_d_652(.A(n_2618), .Y(d_out_652));
CLKBUFX1 gbuf_q_652(.A(q_in_652), .Y(_2162_));
CLKBUFX1 gbuf_d_653(.A(n_2617), .Y(d_out_653));
CLKBUFX1 gbuf_q_653(.A(q_in_653), .Y(_2163_));
CLKBUFX1 gbuf_d_654(.A(n_2622), .Y(d_out_654));
CLKBUFX1 gbuf_q_654(.A(q_in_654), .Y(_2171_));
CLKBUFX1 gbuf_d_655(.A(n_2616), .Y(d_out_655));
CLKBUFX1 gbuf_q_655(.A(q_in_655), .Y(_2174_));
CLKBUFX1 gbuf_d_656(.A(n_2615), .Y(d_out_656));
CLKBUFX1 gbuf_q_656(.A(q_in_656), .Y(_2175_));
CLKBUFX1 gbuf_d_657(.A(n_2563), .Y(d_out_657));
CLKBUFX1 gbuf_q_657(.A(q_in_657), .Y(_2181_));
CLKBUFX1 gbuf_d_658(.A(n_2613), .Y(d_out_658));
CLKBUFX1 gbuf_q_658(.A(q_in_658), .Y(_2194_));
CLKBUFX1 gbuf_d_659(.A(n_2612), .Y(d_out_659));
CLKBUFX1 gbuf_q_659(.A(q_in_659), .Y(_2201_));
CLKBUFX1 gbuf_d_660(.A(n_2611), .Y(d_out_660));
CLKBUFX1 gbuf_q_660(.A(q_in_660), .Y(_2202_));
CLKBUFX1 gbuf_d_661(.A(n_2610), .Y(d_out_661));
CLKBUFX1 gbuf_q_661(.A(q_in_661), .Y(_2205_));
CLKBUFX1 gbuf_d_662(.A(n_2609), .Y(d_out_662));
CLKBUFX1 gbuf_q_662(.A(q_in_662), .Y(_2207_));
CLKBUFX1 gbuf_d_663(.A(n_2608), .Y(d_out_663));
CLKBUFX1 gbuf_q_663(.A(q_in_663), .Y(_2218_));
CLKBUFX1 gbuf_d_664(.A(n_2565), .Y(d_out_664));
CLKBUFX1 gbuf_q_664(.A(q_in_664), .Y(_2220_));
CLKBUFX1 gbuf_d_665(.A(n_2607), .Y(d_out_665));
CLKBUFX1 gbuf_q_665(.A(q_in_665), .Y(_2224_));
CLKBUFX1 gbuf_d_666(.A(n_2600), .Y(d_out_666));
CLKBUFX1 gbuf_q_666(.A(q_in_666), .Y(_2232_));
CLKBUFX1 gbuf_d_667(.A(n_2606), .Y(d_out_667));
CLKBUFX1 gbuf_q_667(.A(q_in_667), .Y(_2237_));
CLKBUFX1 gbuf_d_668(.A(n_2604), .Y(d_out_668));
CLKBUFX1 gbuf_q_668(.A(q_in_668), .Y(_2240_));
CLKBUFX1 gbuf_d_669(.A(n_2564), .Y(d_out_669));
CLKBUFX1 gbuf_q_669(.A(q_in_669), .Y(_2244_));
CLKBUFX1 gbuf_d_670(.A(n_2566), .Y(d_out_670));
CLKBUFX1 gbuf_q_670(.A(q_in_670), .Y(_2246_));
CLKBUFX1 gbuf_d_671(.A(n_2625), .Y(d_out_671));
CLKBUFX1 gbuf_q_671(.A(q_in_671), .Y(_2250_));
CLKBUFX1 gbuf_d_672(.A(n_2602), .Y(d_out_672));
CLKBUFX1 gbuf_q_672(.A(q_in_672), .Y(_2258_));
CLKBUFX1 gbuf_d_673(.A(n_2601), .Y(d_out_673));
CLKBUFX1 gbuf_q_673(.A(q_in_673), .Y(_2262_));
CLKBUFX1 gbuf_d_674(.A(n_2626), .Y(d_out_674));
CLKBUFX1 gbuf_q_674(.A(q_in_674), .Y(_2263_));
CLKBUFX1 gbuf_d_675(.A(n_2599), .Y(d_out_675));
CLKBUFX1 gbuf_q_675(.A(q_in_675), .Y(_2268_));
CLKBUFX1 gbuf_d_676(.A(n_2570), .Y(d_out_676));
CLKBUFX1 gbuf_q_676(.A(q_in_676), .Y(_2281_));
CLKBUFX1 gbuf_d_677(.A(n_2598), .Y(d_out_677));
CLKBUFX1 gbuf_q_677(.A(q_in_677), .Y(_2289_));
CLKBUFX1 gbuf_d_678(.A(n_2597), .Y(d_out_678));
CLKBUFX1 gbuf_q_678(.A(q_in_678), .Y(_2292_));
CLKBUFX1 gbuf_d_679(.A(n_2624), .Y(d_out_679));
CLKBUFX1 gbuf_q_679(.A(q_in_679), .Y(_2295_));
CLKBUFX1 gbuf_d_680(.A(n_2628), .Y(d_out_680));
CLKBUFX1 gbuf_q_680(.A(q_in_680), .Y(_2298_));
CLKBUFX1 gbuf_d_681(.A(n_2595), .Y(d_out_681));
CLKBUFX1 gbuf_q_681(.A(q_in_681), .Y(_2301_));
CLKBUFX1 gbuf_d_682(.A(n_2594), .Y(d_out_682));
CLKBUFX1 gbuf_q_682(.A(q_in_682), .Y(_2302_));
CLKBUFX1 gbuf_d_683(.A(n_2593), .Y(d_out_683));
CLKBUFX1 gbuf_q_683(.A(q_in_683), .Y(_2303_));
CLKBUFX1 gbuf_d_684(.A(n_2591), .Y(d_out_684));
CLKBUFX1 gbuf_q_684(.A(q_in_684), .Y(_2306_));
CLKBUFX1 gbuf_d_685(.A(n_2590), .Y(d_out_685));
CLKBUFX1 gbuf_q_685(.A(q_in_685), .Y(_2307_));
CLKBUFX1 gbuf_d_686(.A(n_2627), .Y(d_out_686));
CLKBUFX1 gbuf_q_686(.A(q_in_686), .Y(_2309_));
CLKBUFX1 gbuf_d_687(.A(n_2589), .Y(d_out_687));
CLKBUFX1 gbuf_q_687(.A(q_in_687), .Y(_2319_));
CLKBUFX1 gbuf_d_688(.A(n_2588), .Y(d_out_688));
CLKBUFX1 gbuf_q_688(.A(q_in_688), .Y(_2327_));
CLKBUFX1 gbuf_d_689(.A(n_2584), .Y(d_out_689));
CLKBUFX1 gbuf_q_689(.A(q_in_689), .Y(_2333_));
CLKBUFX1 gbuf_d_690(.A(n_2582), .Y(d_out_690));
CLKBUFX1 gbuf_q_690(.A(q_in_690), .Y(_2335_));
CLKBUFX1 gbuf_d_691(.A(n_2581), .Y(d_out_691));
CLKBUFX1 gbuf_q_691(.A(q_in_691), .Y(_2348_));
CLKBUFX1 gbuf_d_692(.A(n_2579), .Y(d_out_692));
CLKBUFX1 gbuf_q_692(.A(q_in_692), .Y(_2350_));
CLKBUFX1 gbuf_d_693(.A(n_2576), .Y(d_out_693));
CLKBUFX1 gbuf_q_693(.A(q_in_693), .Y(_2352_));
CLKBUFX1 gbuf_d_694(.A(n_2575), .Y(d_out_694));
CLKBUFX1 gbuf_q_694(.A(q_in_694), .Y(_2353_));
CLKBUFX1 gbuf_d_695(.A(n_2574), .Y(d_out_695));
CLKBUFX1 gbuf_q_695(.A(q_in_695), .Y(_2354_));
CLKBUFX1 gbuf_d_696(.A(n_2568), .Y(d_out_696));
CLKBUFX1 gbuf_q_696(.A(q_in_696), .Y(_2264_));
CLKBUFX1 gbuf_d_697(.A(n_2663), .Y(d_out_697));
CLKBUFX1 gbuf_q_697(.A(q_in_697), .Y(WX11115));
CLKBUFX1 gbuf_d_698(.A(n_2689), .Y(d_out_698));
CLKBUFX1 gbuf_q_698(.A(q_in_698), .Y(WX11153));
CLKBUFX1 gbuf_d_699(.A(n_2677), .Y(d_out_699));
CLKBUFX1 gbuf_q_699(.A(q_in_699), .Y(WX7216));
CLKBUFX1 gbuf_d_700(.A(n_2630), .Y(d_out_700));
CLKBUFX1 gbuf_q_700(.A(q_in_700), .Y(WX7272));
CLKBUFX1 gbuf_d_701(.A(n_2682), .Y(d_out_701));
CLKBUFX1 gbuf_q_701(.A(q_in_701), .Y(WX4606));
CLKBUFX1 gbuf_d_702(.A(n_2686), .Y(d_out_702));
CLKBUFX1 gbuf_q_702(.A(q_in_702), .Y(WX11199));
CLKBUFX1 gbuf_d_703(.A(n_2650), .Y(d_out_703));
CLKBUFX1 gbuf_q_703(.A(q_in_703), .Y(WX11235));
CLKBUFX1 gbuf_d_704(.A(n_2690), .Y(d_out_704));
CLKBUFX1 gbuf_q_704(.A(q_in_704), .Y(WX11239));
CLKBUFX1 gbuf_d_705(.A(n_2665), .Y(d_out_705));
CLKBUFX1 gbuf_q_705(.A(q_in_705), .Y(WX4674));
CLKBUFX1 gbuf_d_706(.A(n_2666), .Y(d_out_706));
CLKBUFX1 gbuf_q_706(.A(q_in_706), .Y(WX3369));
CLKBUFX1 gbuf_d_707(.A(n_2645), .Y(d_out_707));
CLKBUFX1 gbuf_q_707(.A(q_in_707), .Y(WX3401));
CLKBUFX1 gbuf_d_708(.A(n_2667), .Y(d_out_708));
CLKBUFX1 gbuf_q_708(.A(q_in_708), .Y(WX3433));
CLKBUFX1 gbuf_d_709(.A(n_2668), .Y(d_out_709));
CLKBUFX1 gbuf_q_709(.A(q_in_709), .Y(WX3439));
CLKBUFX1 gbuf_d_710(.A(n_2680), .Y(d_out_710));
CLKBUFX1 gbuf_q_710(.A(q_in_710), .Y(WX11169));
CLKBUFX1 gbuf_d_711(.A(n_2660), .Y(d_out_711));
CLKBUFX1 gbuf_q_711(.A(q_in_711), .Y(WX8649));
CLKBUFX1 gbuf_d_712(.A(n_2659), .Y(d_out_712));
CLKBUFX1 gbuf_q_712(.A(q_in_712), .Y(WX8651));
CLKBUFX1 gbuf_d_713(.A(n_2562), .Y(d_out_713));
CLKBUFX1 gbuf_q_713(.A(q_in_713), .Y(WX9804));
CLKBUFX1 gbuf_d_714(.A(n_2671), .Y(d_out_714));
CLKBUFX1 gbuf_q_714(.A(q_in_714), .Y(WX9828));
CLKBUFX1 gbuf_d_715(.A(n_2687), .Y(d_out_715));
CLKBUFX1 gbuf_q_715(.A(q_in_715), .Y(WX9834));
CLKBUFX1 gbuf_d_716(.A(n_2681), .Y(d_out_716));
CLKBUFX1 gbuf_q_716(.A(q_in_716), .Y(WX9872));
CLKBUFX1 gbuf_d_717(.A(n_2673), .Y(d_out_717));
CLKBUFX1 gbuf_q_717(.A(q_in_717), .Y(WX9926));
CLKBUFX1 gbuf_d_718(.A(n_2685), .Y(d_out_718));
CLKBUFX1 gbuf_q_718(.A(q_in_718), .Y(WX4620));
CLKBUFX1 gbuf_d_719(.A(n_2614), .Y(d_out_719));
CLKBUFX1 gbuf_q_719(.A(q_in_719), .Y(WX4638));
CLKBUFX1 gbuf_d_720(.A(n_2670), .Y(d_out_720));
CLKBUFX1 gbuf_q_720(.A(q_in_720), .Y(WX4746));
CLKBUFX1 gbuf_d_721(.A(n_2669), .Y(d_out_721));
CLKBUFX1 gbuf_q_721(.A(q_in_721), .Y(WX4754));
CLKBUFX1 gbuf_d_722(.A(n_2638), .Y(d_out_722));
CLKBUFX1 gbuf_q_722(.A(q_in_722), .Y(WX5927));
CLKBUFX1 gbuf_d_723(.A(n_2664), .Y(d_out_723));
CLKBUFX1 gbuf_q_723(.A(q_in_723), .Y(WX6051));
CLKBUFX1 gbuf_d_724(.A(n_2692), .Y(d_out_724));
CLKBUFX1 gbuf_q_724(.A(q_in_724), .Y(WX2050));
CLKBUFX1 gbuf_d_725(.A(n_2676), .Y(d_out_725));
CLKBUFX1 gbuf_q_725(.A(q_in_725), .Y(WX2064));
CLKBUFX1 gbuf_d_726(.A(n_2633), .Y(d_out_726));
CLKBUFX1 gbuf_q_726(.A(q_in_726), .Y(WX2098));
CLKBUFX1 gbuf_d_727(.A(n_2632), .Y(d_out_727));
CLKBUFX1 gbuf_q_727(.A(q_in_727), .Y(WX2146));
CLKBUFX1 gbuf_d_728(.A(n_2684), .Y(d_out_728));
CLKBUFX1 gbuf_q_728(.A(q_in_728), .Y(WX11207));
INVX4 g63208(.A (n_3168), .Y (n_3264));
CLKBUFX1 gbuf_d_729(.A(n_2603), .Y(d_out_729));
CLKBUFX1 gbuf_q_729(.A(q_in_729), .Y(_2242_));
NOR2X1 g56825(.A (WX3071), .B (n_2849), .Y (n_3167));
CLKBUFX1 gbuf_d_730(.A(n_2573), .Y(d_out_730));
CLKBUFX1 gbuf_q_730(.A(q_in_730), .Y(_2355_));
CLKBUFX1 gbuf_d_731(.A(n_2577), .Y(d_out_731));
CLKBUFX1 gbuf_q_731(.A(q_in_731), .Y(_2351_));
INVX2 g63177(.A (n_4184), .Y (n_5990));
INVX2 g63174(.A (n_4670), .Y (n_3269));
INVX2 g63162(.A (n_6438), .Y (n_6440));
CLKBUFX1 gbuf_d_732(.A(n_1678), .Y(d_out_732));
CLKBUFX1 gbuf_q_732(.A(q_in_732), .Y(WX9816));
NOR2X1 g56925(.A (WX4366), .B (n_2849), .Y (n_3163));
CLKBUFX1 gbuf_d_733(.A(n_2307), .Y(d_out_733));
CLKBUFX1 gbuf_q_733(.A(q_in_733), .Y(WX9924));
CLKBUFX1 gbuf_d_734(.A(n_1487), .Y(d_out_734));
CLKBUFX1 gbuf_qn_734(.A(qn_in_734), .Y(WX8263));
CLKBUFX1 gbuf_d_735(.A(n_1956), .Y(d_out_735));
CLKBUFX1 gbuf_q_735(.A(q_in_735), .Y(WX7206));
CLKBUFX1 gbuf_d_736(.A(n_1830), .Y(d_out_736));
CLKBUFX1 gbuf_q_736(.A(q_in_736), .Y(WX11237));
CLKBUFX1 gbuf_d_737(.A(n_1720), .Y(d_out_737));
CLKBUFX1 gbuf_qn_737(.A(qn_in_737), .Y(WX6972));
BUFX3 g63138(.A (n_3162), .Y (n_3224));
CLKBUFX1 gbuf_d_738(.A(n_2196), .Y(d_out_738));
CLKBUFX1 gbuf_q_738(.A(q_in_738), .Y(WX7202));
CLKBUFX1 gbuf_d_739(.A(n_2405), .Y(d_out_739));
CLKBUFX1 gbuf_q_739(.A(q_in_739), .Y(WX1778));
CLKBUFX1 gbuf_d_740(.A(n_1524), .Y(d_out_740));
CLKBUFX1 gbuf_q_740(.A(q_in_740), .Y(_2346_));
CLKBUFX1 gbuf_d_741(.A(n_1928), .Y(d_out_741));
CLKBUFX1 gbuf_q_741(.A(q_in_741), .Y(WX4758));
CLKBUFX1 gbuf_d_742(.A(n_1565), .Y(d_out_742));
CLKBUFX1 gbuf_q_742(.A(q_in_742), .Y(_2270_));
CLKBUFX1 gbuf_d_743(.A(n_1688), .Y(d_out_743));
CLKBUFX1 gbuf_q_743(.A(q_in_743), .Y(_2296_));
CLKBUFX1 gbuf_d_744(.A(n_1694), .Y(d_out_744));
CLKBUFX1 gbuf_q_744(.A(q_in_744), .Y(_2347_));
BUFX3 g63129(.A (n_3162), .Y (n_3223));
CLKBUFX1 gbuf_d_745(.A(n_1605), .Y(d_out_745));
CLKBUFX1 gbuf_q_745(.A(q_in_745), .Y(_2196_));
CLKBUFX1 gbuf_d_746(.A(n_1905), .Y(d_out_746));
CLKBUFX1 gbuf_q_746(.A(q_in_746), .Y(WX6025));
CLKBUFX1 gbuf_d_747(.A(n_1900), .Y(d_out_747));
CLKBUFX1 gbuf_qn_747(.A(qn_in_747), .Y(WX3099));
CLKBUFX1 gbuf_d_748(.A(n_1582), .Y(d_out_748));
CLKBUFX1 gbuf_q_748(.A(q_in_748), .Y(_2235_));
CLKBUFX1 gbuf_d_749(.A(n_2094), .Y(d_out_749));
CLKBUFX1 gbuf_q_749(.A(q_in_749), .Y(WX8631));
BUFX3 g63120(.A (n_3162), .Y (n_3222));
INVX4 g63109(.A (n_6626), .Y (n_3221));
CLKBUFX1 gbuf_d_750(.A(n_2055), .Y(d_out_750));
CLKBUFX1 gbuf_q_750(.A(q_in_750), .Y(WX2166));
CLKBUFX1 gbuf_d_751(.A(n_1633), .Y(d_out_751));
CLKBUFX1 gbuf_q_751(.A(q_in_751), .Y(_2161_));
CLKBUFX1 gbuf_d_752(.A(n_1658), .Y(d_out_752));
CLKBUFX1 gbuf_q_752(.A(q_in_752), .Y(_2127_));
CLKBUFX1 gbuf_d_753(.A(n_2085), .Y(d_out_753));
CLKBUFX1 gbuf_q_753(.A(q_in_753), .Y(WX11079));
CLKBUFX1 gbuf_d_754(.A(n_2525), .Y(d_out_754));
CLKBUFX1 gbuf_q_754(.A(q_in_754), .Y(WX5893));
CLKBUFX1 gbuf_d_755(.A(n_1891), .Y(d_out_755));
CLKBUFX1 gbuf_q_755(.A(q_in_755), .Y(WX8543));
CLKBUFX1 gbuf_d_756(.A(n_1615), .Y(d_out_756));
CLKBUFX1 gbuf_q_756(.A(q_in_756), .Y(_2182_));
CLKBUFX1 gbuf_d_757(.A(n_1636), .Y(d_out_757));
CLKBUFX1 gbuf_q_757(.A(q_in_757), .Y(_2158_));
CLKBUFX1 gbuf_d_758(.A(n_1922), .Y(d_out_758));
CLKBUFX1 gbuf_q_758(.A(q_in_758), .Y(WX2174));
CLKBUFX1 gbuf_d_759(.A(n_2002), .Y(d_out_759));
CLKBUFX1 gbuf_q_759(.A(q_in_759), .Y(WX2156));
CLKBUFX1 gbuf_d_760(.A(n_1660), .Y(d_out_760));
CLKBUFX1 gbuf_q_760(.A(q_in_760), .Y(_2124_));
CLKBUFX1 gbuf_d_761(.A(n_1503), .Y(d_out_761));
CLKBUFX1 gbuf_q_761(.A(q_in_761), .Y(_2160_));
BUFX3 g63074(.A (n_4562), .Y (n_4628));
BUFX3 g63088(.A (n_6626), .Y (n_4105));
CLKBUFX1 gbuf_d_762(.A(n_2013), .Y(d_out_762));
CLKBUFX1 gbuf_q_762(.A(q_in_762), .Y(WX11063));
CLKBUFX1 gbuf_d_763(.A(n_1604), .Y(d_out_763));
CLKBUFX1 gbuf_q_763(.A(q_in_763), .Y(_2197_));
CLKBUFX1 gbuf_d_764(.A(n_2247), .Y(d_out_764));
CLKBUFX1 gbuf_q_764(.A(q_in_764), .Y(WX2192));
CLKBUFX1 gbuf_d_765(.A(n_2194), .Y(d_out_765));
CLKBUFX1 gbuf_q_765(.A(q_in_765), .Y(WX2182));
BUFX3 g63076(.A (n_4562), .Y (n_4471));
CLKBUFX1 gbuf_d_766(.A(n_1581), .Y(d_out_766));
CLKBUFX1 gbuf_q_766(.A(q_in_766), .Y(_2236_));
CLKBUFX1 gbuf_d_767(.A(n_1951), .Y(d_out_767));
CLKBUFX1 gbuf_q_767(.A(q_in_767), .Y(WX11129));
INVX2 g63065(.A (n_3158), .Y (n_3173));
CLKBUFX1 gbuf_d_768(.A(n_2067), .Y(d_out_768));
CLKBUFX1 gbuf_q_768(.A(q_in_768), .Y(WX4734));
CLKBUFX1 gbuf_d_769(.A(n_1737), .Y(d_out_769));
CLKBUFX1 gbuf_q_769(.A(q_in_769), .Y(WX11071));
CLKBUFX1 gbuf_d_770(.A(n_2172), .Y(d_out_770));
CLKBUFX1 gbuf_q_770(.A(q_in_770), .Y(WX2124));
CLKBUFX1 gbuf_d_771(.A(n_1597), .Y(d_out_771));
CLKBUFX1 gbuf_q_771(.A(q_in_771), .Y(_2212_));
CLKBUFX1 gbuf_d_772(.A(n_2193), .Y(d_out_772));
CLKBUFX1 gbuf_q_772(.A(q_in_772), .Y(WX4690));
CLKBUFX1 gbuf_d_773(.A(n_1723), .Y(d_out_773));
CLKBUFX1 gbuf_q_773(.A(q_in_773), .Y(WX4596));
CLKBUFX1 gbuf_d_774(.A(n_2143), .Y(d_out_774));
CLKBUFX1 gbuf_q_774(.A(q_in_774), .Y(WX4716));
CLKBUFX3 g63060(.A (n_3158), .Y (n_3831));
MX2X1 g60707(.A (n_3027), .B (n_6422), .S0 (WX4540), .Y (n_3157));
MX2X1 g60711(.A (n_3140), .B (n_2938), .S0 (WX4554), .Y (n_3156));
CLKBUFX1 gbuf_d_775(.A(n_2035), .Y(d_out_775));
CLKBUFX1 gbuf_q_775(.A(q_in_775), .Y(WX4612));
MX2X1 g60716(.A (n_3058), .B (n_2775), .S0 (WX8461), .Y (n_3155));
MX2X1 g60718(.A (n_3106), .B (n_2837), .S0 (WX8463), .Y (n_3154));
MX2X1 g60719(.A (n_3137), .B (n_3086), .S0 (WX4544), .Y (n_3153));
MX2X1 g60722(.A (n_2776), .B (n_2996), .S0 (WX8465), .Y (n_3152));
MX2X1 g60726(.A (n_3137), .B (n_2938), .S0 (WX4546), .Y (n_3151));
CLKBUFX1 gbuf_d_776(.A(n_1500), .Y(d_out_776));
CLKBUFX1 gbuf_q_776(.A(q_in_776), .Y(_2278_));
MX2X1 g60729(.A (n_3137), .B (n_3072), .S0 (WX4548), .Y (n_3149));
MX2X1 g60733(.A (n_3021), .B (n_3086), .S0 (WX4550), .Y (n_3147));
MX2X1 g60735(.A (n_3021), .B (n_3041), .S0 (WX4552), .Y (n_3145));
MX2X1 g60739(.A (n_2798), .B (n_3004), .S0 (WX4556), .Y (n_3142));
CLKBUFX1 gbuf_d_777(.A(n_2159), .Y(d_out_777));
CLKBUFX1 gbuf_q_777(.A(q_in_777), .Y(WX4652));
MX2X1 g60745(.A (n_3140), .B (n_3086), .S0 (WX5845), .Y (n_3141));
MX2X1 g60746(.A (n_2986), .B (n_3056), .S0 (WX4560), .Y (n_3139));
MX2X1 g60751(.A (n_3137), .B (n_3086), .S0 (WX9698), .Y (n_3138));
CLKBUFX1 gbuf_d_778(.A(n_1870), .Y(d_out_778));
CLKBUFX1 gbuf_q_778(.A(q_in_778), .Y(WX4654));
MX2X1 g60755(.A (n_3137), .B (n_7488), .S0 (WX8413), .Y (n_3136));
MX2X1 g60758(.A (n_3031), .B (n_2938), .S0 (WX9700), .Y (n_3135));
MX2X1 g60761(.A (n_3031), .B (n_3041), .S0 (WX9702), .Y (n_3134));
MX2X1 g60769(.A (n_3027), .B (n_6422), .S0 (WX9706), .Y (n_3131));
MX2X1 g60774(.A (n_2815), .B (n_2976), .S0 (WX5849), .Y (n_3128));
MX2X1 g60776(.A (n_3137), .B (n_2945), .S0 (WX9708), .Y (n_3127));
MX2X1 g60780(.A (n_2838), .B (n_3044), .S0 (WX9730), .Y (n_3126));
CLKBUFX1 gbuf_d_779(.A(n_1672), .Y(d_out_779));
CLKBUFX1 gbuf_q_779(.A(q_in_779), .Y(WX7244));
CLKBUFX1 gbuf_d_780(.A(n_2138), .Y(d_out_780));
CLKBUFX1 gbuf_q_780(.A(q_in_780), .Y(WX9786));
MX2X1 g60782(.A (n_3137), .B (n_6422), .S0 (WX9712), .Y (n_3125));
MX2X1 g60788(.A (n_3120), .B (n_7488), .S0 (WX3231), .Y (n_3123));
MX2X1 g60793(.A (n_3120), .B (n_3086), .S0 (WX9722), .Y (n_3121));
MX2X1 g60801(.A (n_3140), .B (n_3072), .S0 (WX9726), .Y (n_3118));
CLKBUFX1 gbuf_d_781(.A(n_1557), .Y(d_out_781));
CLKBUFX1 gbuf_q_781(.A(q_in_781), .Y(_2287_));
MX2X1 g60805(.A (n_3058), .B (n_3105), .S0 (WX9728), .Y (n_3117));
MX2X1 g60810(.A (n_3106), .B (n_3103), .S0 (WX4578), .Y (n_3116));
CLKBUFX1 gbuf_d_782(.A(n_2305), .Y(d_out_782));
CLKBUFX1 gbuf_q_782(.A(q_in_782), .Y(WX7290));
MX2X1 g60811(.A (n_3106), .B (n_2775), .S0 (WX5875), .Y (n_3115));
MX2X1 g60816(.A (n_3031), .B (n_2945), .S0 (WX5847), .Y (n_3114));
MX2X1 g60821(.A (n_3058), .B (n_2837), .S0 (WX4582), .Y (n_3113));
CLKBUFX1 gbuf_d_783(.A(n_2320), .Y(d_out_783));
CLKBUFX1 gbuf_q_783(.A(q_in_783), .Y(WX7294));
MX2X1 g60828(.A (n_3031), .B (n_3041), .S0 (WX11007), .Y (n_3111));
CLKBUFX1 gbuf_d_784(.A(n_1709), .Y(d_out_784));
CLKBUFX1 gbuf_q_784(.A(q_in_784), .Y(WX7330));
CLKBUFX1 gbuf_d_785(.A(n_2233), .Y(d_out_785));
CLKBUFX1 gbuf_q_785(.A(q_in_785), .Y(WX4702));
MX2X1 g60838(.A (n_3106), .B (n_2837), .S0 (WX4586), .Y (n_3110));
MX2X1 g60843(.A (n_3106), .B (n_3089), .S0 (WX11045), .Y (n_3108));
MX2X1 g60846(.A (n_3106), .B (n_3105), .S0 (WX9750), .Y (n_3107));
MX2X1 g60848(.A (n_2935), .B (n_3103), .S0 (WX9752), .Y (n_3104));
MX2X1 g60856(.A (n_2798), .B (n_3105), .S0 (WX5879), .Y (n_3102));
MX2X1 g60857(.A (n_3106), .B (n_3089), .S0 (WX9756), .Y (n_3101));
CLKBUFX1 gbuf_d_786(.A(n_2181), .Y(d_out_786));
CLKBUFX1 gbuf_q_786(.A(q_in_786), .Y(WX7196));
MX2X1 g60860(.A (n_3027), .B (n_3041), .S0 (WX3237), .Y (n_3099));
MX2X1 g60861(.A (n_3027), .B (n_2945), .S0 (WX10993), .Y (n_3098));
MX2X1 g60866(.A (n_3027), .B (n_3072), .S0 (WX9710), .Y (n_3096));
MX2X1 g60867(.A (n_3027), .B (n_2945), .S0 (WX10995), .Y (n_3095));
MX2X1 g60868(.A (n_3027), .B (n_3072), .S0 (WX3239), .Y (n_3093));
MX2X1 g60874(.A (n_3027), .B (n_2945), .S0 (WX3241), .Y (n_3092));
MX2X1 g60875(.A (n_3058), .B (n_3089), .S0 (WX5863), .Y (n_3090));
MX2X1 g60877(.A (n_3021), .B (n_2945), .S0 (WX11003), .Y (n_3088));
MX2X1 g60884(.A (n_3021), .B (n_3086), .S0 (WX5819), .Y (n_3087));
MX2X1 g60885(.A (n_3120), .B (n_3072), .S0 (WX10997), .Y (n_3085));
CLKBUFX1 gbuf_d_787(.A(n_2300), .Y(d_out_787));
CLKBUFX1 gbuf_q_787(.A(q_in_787), .Y(WX7286));
CLKBUFX1 gbuf_d_788(.A(n_1931), .Y(d_out_788));
CLKBUFX1 gbuf_q_788(.A(q_in_788), .Y(WX4636));
MX2X1 g60897(.A (n_3120), .B (n_3072), .S0 (WX5823), .Y (n_3083));
CLKBUFX1 gbuf_d_789(.A(n_2240), .Y(d_out_789));
CLKBUFX1 gbuf_q_789(.A(q_in_789), .Y(WX11163));
MX2X1 g60900(.A (n_3027), .B (n_3041), .S0 (WX5825), .Y (n_3081));
MX2X1 g60910(.A (n_3027), .B (n_3072), .S0 (WX5829), .Y (n_3080));
MX2X1 g60911(.A (n_3137), .B (n_3041), .S0 (WX5817), .Y (n_3077));
MX2X1 g60912(.A (n_3137), .B (n_3086), .S0 (WX5831), .Y (n_3076));
MX2X1 g60916(.A (n_3137), .B (n_3072), .S0 (WX5833), .Y (n_3075));
CLKBUFX1 gbuf_d_790(.A(n_1515), .Y(d_out_790));
CLKBUFX1 gbuf_q_790(.A(q_in_790), .Y(_2267_));
MX2X1 g60918(.A (n_3137), .B (n_3072), .S0 (WX3247), .Y (n_3074));
MX2X1 g60922(.A (n_3027), .B (n_2945), .S0 (WX5841), .Y (n_3071));
CLKBUFX1 gbuf_d_791(.A(n_2015), .Y(d_out_791));
CLKBUFX1 gbuf_q_791(.A(q_in_791), .Y(WX8601));
MX2X1 g60924(.A (n_3137), .B (n_2945), .S0 (WX5843), .Y (n_3069));
MX2X1 g60925(.A (n_3137), .B (n_3072), .S0 (WX8433), .Y (n_3068));
CLKBUFX1 gbuf_d_792(.A(n_2201), .Y(d_out_792));
CLKBUFX1 gbuf_q_792(.A(q_in_792), .Y(WX3365));
MX2X1 g60929(.A (n_3106), .B (n_2988), .S0 (WX5877), .Y (n_3066));
MX2X1 g60932(.A (n_3021), .B (n_3072), .S0 (WX11013), .Y (n_3065));
MX2X1 g60936(.A (n_3021), .B (n_3072), .S0 (WX11005), .Y (n_3064));
CLKBUFX1 gbuf_d_793(.A(n_1801), .Y(d_out_793));
CLKBUFX1 gbuf_q_793(.A(q_in_793), .Y(WX2092));
MX2X1 g60946(.A (n_3106), .B (n_3089), .S0 (WX5861), .Y (n_3062));
MX2X1 g60948(.A (n_3021), .B (n_3072), .S0 (WX8427), .Y (n_3061));
MX2X1 g60952(.A (n_3058), .B (n_2953), .S0 (WX5865), .Y (n_3059));
MX2X1 g60953(.A (n_2829), .B (n_3056), .S0 (WX4574), .Y (n_3057));
MX2X1 g60954(.A (n_3021), .B (n_2945), .S0 (WX4542), .Y (n_3055));
MX2X1 g60958(.A (n_3021), .B (n_3041), .S0 (WX11009), .Y (n_3054));
MX2X1 g60960(.A (n_3137), .B (n_3041), .S0 (WX3253), .Y (n_3052));
CLKBUFX1 gbuf_d_794(.A(n_1885), .Y(d_out_794));
CLKBUFX1 gbuf_q_794(.A(q_in_794), .Y(WX2086));
MX2X1 g60962(.A (n_3137), .B (n_2938), .S0 (WX3259), .Y (n_3051));
MX2X1 g60967(.A (n_3120), .B (n_2945), .S0 (WX11011), .Y (n_3049));
CLKBUFX1 gbuf_d_795(.A(n_2080), .Y(d_out_795));
CLKBUFX1 gbuf_q_795(.A(q_in_795), .Y(WX2150));
CLKBUFX1 gbuf_d_796(.A(n_1988), .Y(d_out_796));
CLKBUFX1 gbuf_q_796(.A(q_in_796), .Y(WX11125));
MX2X1 g60980(.A (n_2986), .B (n_3056), .S0 (WX11035), .Y (n_3048));
MX2X1 g60983(.A (n_3120), .B (n_3072), .S0 (WX11015), .Y (n_3047));
MX2X1 g60989(.A (n_2829), .B (n_3044), .S0 (WX3265), .Y (n_3045));
CLKBUFX1 gbuf_d_797(.A(n_2205), .Y(d_out_797));
CLKBUFX1 gbuf_q_797(.A(q_in_797), .Y(WX3385));
CLKBUFX1 gbuf_d_798(.A(n_2197), .Y(d_out_798));
CLKBUFX1 gbuf_q_798(.A(q_in_798), .Y(WX7336));
CLKBUFX1 gbuf_d_799(.A(n_1948), .Y(d_out_799));
CLKBUFX1 gbuf_q_799(.A(q_in_799), .Y(WX2138));
MX2X1 g60992(.A (n_6423), .B (n_3041), .S0 (WX3245), .Y (n_3043));
MX2X1 g60993(.A (n_3137), .B (n_3072), .S0 (WX7140), .Y (n_3040));
MX2X1 g60994(.A (n_3137), .B (n_3041), .S0 (WX3261), .Y (n_3039));
CLKBUFX1 gbuf_d_800(.A(n_1999), .Y(d_out_800));
CLKBUFX1 gbuf_q_800(.A(q_in_800), .Y(WX7332));
MX2X1 g61003(.A (n_7483), .B (n_3072), .S0 (WX7110), .Y (n_3038));
MX2X1 g61004(.A (n_3058), .B (n_2828), .S0 (WX3267), .Y (n_3037));
MX2X1 g61009(.A (n_3031), .B (n_3072), .S0 (WX7112), .Y (n_3034));
MX2X1 g61014(.A (n_3031), .B (n_3086), .S0 (WX7114), .Y (n_3032));
MX2X1 g61018(.A (n_3031), .B (n_2945), .S0 (WX7116), .Y (n_3030));
MX2X1 g61023(.A (n_3027), .B (n_3072), .S0 (WX5835), .Y (n_3029));
MX2X1 g61024(.A (n_3027), .B (n_3086), .S0 (WX11019), .Y (n_3028));
MX2X1 g61026(.A (n_7483), .B (n_3072), .S0 (WX7118), .Y (n_3026));
MX2X1 g61031(.A (n_7483), .B (n_3041), .S0 (WX7120), .Y (n_3024));
MX2X1 g61037(.A (n_3021), .B (n_3072), .S0 (WX7122), .Y (n_3023));
MX2X1 g61039(.A (n_3021), .B (n_3072), .S0 (WX5827), .Y (n_3022));
MX2X1 g61041(.A (n_3021), .B (n_3041), .S0 (WX7124), .Y (n_3020));
MX2X1 g61045(.A (n_3021), .B (n_3041), .S0 (WX7126), .Y (n_3018));
MX2X1 g61046(.A (n_3021), .B (n_7488), .S0 (WX9720), .Y (n_3017));
MX2X1 g61049(.A (n_3021), .B (n_3086), .S0 (WX5837), .Y (n_3015));
MX2X1 g61053(.A (n_3021), .B (n_3072), .S0 (WX7128), .Y (n_3014));
CLKBUFX1 gbuf_d_801(.A(n_2299), .Y(d_out_801));
CLKBUFX1 gbuf_q_801(.A(q_in_801), .Y(WX9920));
CLKBUFX1 gbuf_d_802(.A(n_1509), .Y(d_out_802));
CLKBUFX1 gbuf_q_802(.A(q_in_802), .Y(_2304_));
CLKBUFX1 gbuf_d_803(.A(n_1913), .Y(d_out_803));
CLKBUFX1 gbuf_q_803(.A(q_in_803), .Y(WX8605));
MX2X1 g61059(.A (n_3027), .B (n_3086), .S0 (WX7130), .Y (n_3012));
MX2X1 g61060(.A (n_2986), .B (n_3044), .S0 (WX3273), .Y (n_3011));
MX2X1 g61067(.A (n_3027), .B (n_3072), .S0 (WX7132), .Y (n_3009));
CLKBUFX1 gbuf_d_804(.A(n_1510), .Y(d_out_804));
CLKBUFX1 gbuf_q_804(.A(q_in_804), .Y(_2117_));
MX2X1 g61070(.A (n_3058), .B (n_2993), .S0 (WX3275), .Y (n_3007));
MX2X1 g61071(.A (n_2776), .B (n_3004), .S0 (WX11023), .Y (n_3005));
MX2X1 g61072(.A (n_3021), .B (n_3072), .S0 (WX7134), .Y (n_3003));
MX2X1 g61076(.A (n_3021), .B (n_3041), .S0 (WX9718), .Y (n_3001));
MX2X1 g61077(.A (n_3021), .B (n_3086), .S0 (WX7136), .Y (n_3000));
MX2X1 g61082(.A (n_3021), .B (n_3072), .S0 (WX7138), .Y (n_2999));
MX2X1 g61087(.A (n_3106), .B (n_2817), .S0 (WX4584), .Y (n_2998));
MX2X1 g61094(.A (n_3058), .B (n_2996), .S0 (WX7142), .Y (n_2997));
MX2X1 g61099(.A (n_3106), .B (n_3105), .S0 (WX7144), .Y (n_2995));
MX2X1 g61104(.A (n_2813), .B (n_2993), .S0 (WX7146), .Y (n_2994));
MX2X1 g61108(.A (n_3106), .B (n_2770), .S0 (WX7148), .Y (n_2992));
CLKBUFX1 gbuf_d_805(.A(n_1807), .Y(d_out_805));
CLKBUFX1 gbuf_q_805(.A(q_in_805), .Y(WX7242));
CLKBUFX1 gbuf_d_806(.A(n_1529), .Y(d_out_806));
CLKBUFX1 gbuf_q_806(.A(q_in_806), .Y(_2341_));
MX2X1 g61112(.A (n_2986), .B (n_2996), .S0 (WX7150), .Y (n_2991));
MX2X1 g61126(.A (n_3058), .B (n_2988), .S0 (WX7156), .Y (n_2990));
CLKBUFX1 gbuf_d_807(.A(n_1691), .Y(d_out_807));
CLKBUFX1 gbuf_q_807(.A(q_in_807), .Y(_2153_));
MX2X1 g61127(.A (n_2986), .B (n_3103), .S0 (WX3281), .Y (n_2987));
MX2X1 g61129(.A (n_6513), .B (n_3004), .S0 (WX7158), .Y (n_2985));
MX2X1 g61131(.A (n_2798), .B (n_3103), .S0 (WX11029), .Y (n_2984));
MX2X1 g61132(.A (n_2986), .B (n_2993), .S0 (WX8449), .Y (n_2982));
CLKBUFX1 gbuf_d_808(.A(n_1611), .Y(d_out_808));
CLKBUFX1 gbuf_q_808(.A(q_in_808), .Y(_2190_));
CLKBUFX1 gbuf_d_809(.A(n_1986), .Y(d_out_809));
CLKBUFX1 gbuf_q_809(.A(q_in_809), .Y(WX8633));
MX2X1 g61139(.A (n_3106), .B (n_2755), .S0 (WX7162), .Y (n_2981));
MX2X1 g61147(.A (n_3106), .B (n_3056), .S0 (WX7166), .Y (n_2979));
MX2X1 g61149(.A (n_2829), .B (n_2976), .S0 (WX3285), .Y (n_2978));
MX2X1 g61150(.A (n_3058), .B (n_2755), .S0 (WX11031), .Y (n_2975));
CLKBUFX1 gbuf_d_810(.A(n_2392), .Y(d_out_810));
CLKBUFX1 gbuf_q_810(.A(q_in_810), .Y(WX9916));
CLKBUFX1 gbuf_d_811(.A(n_1964), .Y(d_out_811));
CLKBUFX1 gbuf_q_811(.A(q_in_811), .Y(WX8493));
MX2X1 g61166(.A (n_3058), .B (n_2795), .S0 (WX7172), .Y (n_2974));
MX2X1 g61169(.A (n_3021), .B (n_3072), .S0 (WX9716), .Y (n_2972));
MX2X1 g61171(.A (n_3058), .B (n_2755), .S0 (WX11033), .Y (n_2971));
CLKBUFX1 gbuf_d_812(.A(n_2179), .Y(d_out_812));
CLKBUFX1 gbuf_q_812(.A(q_in_812), .Y(WX3345));
MX2X1 g61187(.A (n_3137), .B (n_3072), .S0 (WX3243), .Y (n_2969));
MX2X1 g61188(.A (n_3058), .B (n_3044), .S0 (WX11037), .Y (n_2968));
MX2X1 g61189(.A (n_3058), .B (n_2988), .S0 (WX3293), .Y (n_2967));
MX2X1 g61197(.A (n_3058), .B (n_2795), .S0 (WX11039), .Y (n_2966));
CLKBUFX1 gbuf_d_813(.A(n_2253), .Y(d_out_813));
CLKBUFX1 gbuf_q_813(.A(q_in_813), .Y(WX9790));
CLKBUFX1 gbuf_d_814(.A(n_2231), .Y(d_out_814));
CLKBUFX1 gbuf_q_814(.A(q_in_814), .Y(WX9794));
MX2X1 g61212(.A (n_3137), .B (n_3072), .S0 (WX8405), .Y (n_2965));
MX2X1 g61215(.A (n_3137), .B (n_2938), .S0 (WX8407), .Y (n_2963));
CLKBUFX1 gbuf_d_815(.A(n_1965), .Y(d_out_815));
CLKBUFX1 gbuf_q_815(.A(q_in_815), .Y(WX9868));
MX2X1 g61218(.A (n_3021), .B (n_2938), .S0 (WX8409), .Y (n_2961));
CLKBUFX1 gbuf_d_816(.A(n_1584), .Y(d_out_816));
CLKBUFX1 gbuf_q_816(.A(q_in_816), .Y(_2231_));
MX2X1 g61221(.A (n_3021), .B (n_2938), .S0 (WX8411), .Y (n_2960));
CLKBUFX1 gbuf_d_817(.A(n_1551), .Y(d_out_817));
CLKBUFX1 gbuf_q_817(.A(q_in_817), .Y(_2310_));
MX2X1 g61225(.A (n_3137), .B (n_2945), .S0 (WX11001), .Y (n_2958));
MX2X1 g61226(.A (n_3137), .B (n_3041), .S0 (WX5821), .Y (n_2957));
CLKBUFX1 gbuf_d_818(.A(n_2129), .Y(d_out_818));
CLKBUFX1 gbuf_q_818(.A(q_in_818), .Y(WX9824));
MX2X1 g61228(.A (n_3021), .B (n_3072), .S0 (WX10999), .Y (n_2955));
MX2X1 g61238(.A (n_3058), .B (n_2953), .S0 (WX9732), .Y (n_2954));
MX2X1 g61244(.A (n_3137), .B (n_3072), .S0 (WX8421), .Y (n_2952));
CLKBUFX1 gbuf_d_819(.A(n_2124), .Y(d_out_819));
CLKBUFX1 gbuf_q_819(.A(q_in_819), .Y(WX9832));
MX2X1 g61248(.A (n_3137), .B (n_3072), .S0 (WX8423), .Y (n_2950));
CLKBUFX1 gbuf_d_820(.A(n_2379), .Y(d_out_820));
CLKBUFX1 gbuf_q_820(.A(q_in_820), .Y(WX11175));
CLKBUFX1 gbuf_d_821(.A(n_2178), .Y(d_out_821));
CLKBUFX1 gbuf_q_821(.A(q_in_821), .Y(WX3311));
MX2X1 g61252(.A (n_3140), .B (n_2938), .S0 (WX8425), .Y (n_2949));
MX2X1 g61259(.A (n_3137), .B (n_3072), .S0 (WX4526), .Y (n_2948));
CLKBUFX1 gbuf_d_822(.A(n_1895), .Y(d_out_822));
CLKBUFX1 gbuf_q_822(.A(q_in_822), .Y(WX2134));
MX2X1 g61266(.A (n_3137), .B (n_2938), .S0 (WX8429), .Y (n_2947));
MX2X1 g61269(.A (n_3021), .B (n_2945), .S0 (WX8431), .Y (n_2946));
MX2X1 g61272(.A (n_3021), .B (n_3041), .S0 (WX4528), .Y (n_2944));
MX2X1 g61277(.A (n_3021), .B (n_2945), .S0 (WX9714), .Y (n_2943));
MX2X1 g61278(.A (n_3021), .B (n_2945), .S0 (WX4530), .Y (n_2941));
CLKBUFX1 gbuf_d_823(.A(n_1587), .Y(d_out_823));
CLKBUFX1 gbuf_q_823(.A(q_in_823), .Y(_2229_));
MX2X1 g61283(.A (n_2809), .B (n_3004), .S0 (WX8437), .Y (n_2940));
CLKBUFX1 gbuf_d_824(.A(n_1974), .Y(d_out_824));
CLKBUFX1 gbuf_q_824(.A(q_in_824), .Y(WX11121));
MX2X1 g61287(.A (n_3021), .B (n_2938), .S0 (WX4532), .Y (n_2939));
MX2X1 g61291(.A (n_3106), .B (n_2993), .S0 (WX8441), .Y (n_2937));
CLKBUFX1 gbuf_d_825(.A(n_1608), .Y(d_out_825));
CLKBUFX1 gbuf_q_825(.A(q_in_825), .Y(_2192_));
MX2X1 g61293(.A (n_2935), .B (n_2976), .S0 (WX9736), .Y (n_2936));
MX2X1 g61294(.A (n_3021), .B (n_2938), .S0 (WX4534), .Y (n_2934));
MX2X1 g61296(.A (n_3106), .B (n_2976), .S0 (WX8445), .Y (n_2933));
MX2X1 g61299(.A (n_3137), .B (n_2938), .S0 (WX4536), .Y (n_2932));
MX2X1 g61305(.A (n_3031), .B (n_2945), .S0 (WX4538), .Y (n_2931));
MX2X1 g61308(.A (n_6513), .B (n_2996), .S0 (WX5857), .Y (n_2930));
NOR2X1 g61336(.A (WX10829), .B (n_2849), .Y (n_2928));
NOR2X1 g61341(.A (n_2849), .B (WX485), .Y (n_2927));
CLKBUFX1 gbuf_d_826(.A(n_2312), .Y(d_out_826));
CLKBUFX1 gbuf_q_826(.A(q_in_826), .Y(WX9826));
CLKBUFX1 gbuf_d_827(.A(n_1904), .Y(d_out_827));
CLKBUFX1 gbuf_q_827(.A(q_in_827), .Y(WX8575));
CLKBUFX1 gbuf_d_828(.A(n_1750), .Y(d_out_828));
CLKBUFX1 gbuf_q_828(.A(q_in_828), .Y(WX2108));
INVX2 g61376(.A (n_2926), .Y (n_5493));
INVX2 g61377(.A (n_2926), .Y (n_5183));
INVX1 g61378(.A (n_2926), .Y (n_5085));
INVX2 g61379(.A (n_2926), .Y (n_4803));
INVX1 g61380(.A (n_2926), .Y (n_5254));
INVX1 g61385(.A (n_2925), .Y (n_5474));
INVX1 g61386(.A (n_2925), .Y (n_5600));
INVX1 g61387(.A (n_2925), .Y (n_5918));
INVX1 g61388(.A (n_2925), .Y (n_5320));
INVX1 g61389(.A (n_2925), .Y (n_5598));
INVX1 g61390(.A (n_2925), .Y (n_5239));
INVX1 g61391(.A (n_2925), .Y (n_4866));
INVX1 g61392(.A (n_2925), .Y (n_5549));
INVX2 g61395(.A (n_2924), .Y (n_5415));
INVX2 g61396(.A (n_2924), .Y (n_5928));
INVX1 g61397(.A (n_2924), .Y (n_5196));
CLKBUFX1 gbuf_d_829(.A(n_2275), .Y(d_out_829));
CLKBUFX1 gbuf_q_829(.A(q_in_829), .Y(WX3415));
INVX1 g61398(.A (n_2924), .Y (n_5317));
INVX1 g61399(.A (n_2924), .Y (n_4868));
INVX1 g61400(.A (n_2924), .Y (n_5630));
INVX1 g61404(.A (n_6482), .Y (n_5750));
INVX1 g61405(.A (n_6482), .Y (n_5334));
INVX4 g61406(.A (n_6482), .Y (n_5439));
INVX1 g61408(.A (n_6482), .Y (n_5649));
INVX1 g61410(.A (n_6482), .Y (n_5158));
INVX8 g61418(.A (n_2922), .Y (n_4697));
INVX2 g61421(.A (n_2921), .Y (n_5235));
INVX1 g61422(.A (n_2921), .Y (n_5576));
INVX1 g61424(.A (n_2921), .Y (n_5886));
INVX1 g61425(.A (n_2921), .Y (n_5845));
INVX1 g61426(.A (n_2921), .Y (n_5729));
INVX1 g61427(.A (n_2921), .Y (n_5418));
INVX1 g61428(.A (n_2921), .Y (n_5482));
INVX1 g61430(.A (n_7090), .Y (n_5393));
INVX1 g61432(.A (n_7090), .Y (n_5882));
INVX1 g61433(.A (n_7090), .Y (n_5185));
INVX4 g61435(.A (n_7090), .Y (n_5841));
INVX1 g61437(.A (n_7090), .Y (n_6106));
INVX4 g61440(.A (n_6503), .Y (n_5535));
INVX2 g61441(.A (n_6503), .Y (n_5468));
INVX1 g61444(.A (n_6503), .Y (n_5830));
INVX1 g61445(.A (n_6503), .Y (n_6050));
INVX1 g61446(.A (n_6503), .Y (n_5490));
INVX2 g61448(.A (n_2920), .Y (n_5879));
INVX1 g61451(.A (n_2920), .Y (n_5825));
INVX2 g61452(.A (n_2920), .Y (n_5105));
INVX2 g61454(.A (n_2920), .Y (n_5892));
INVX1 g61455(.A (n_2920), .Y (n_5834));
CLKBUFX1 gbuf_d_830(.A(n_1645), .Y(d_out_830));
CLKBUFX1 gbuf_q_830(.A(q_in_830), .Y(_2144_));
NOR2X1 g61468(.A (WX1778), .B (n_2849), .Y (n_2917));
CLKBUFX1 gbuf_d_831(.A(n_1962), .Y(d_out_831));
CLKBUFX1 gbuf_q_831(.A(q_in_831), .Y(WX6065));
CLKBUFX1 gbuf_d_832(.A(n_2323), .Y(d_out_832));
CLKBUFX1 gbuf_q_832(.A(q_in_832), .Y(WX5997));
CLKBUFX1 gbuf_d_833(.A(n_1613), .Y(d_out_833));
CLKBUFX1 gbuf_q_833(.A(q_in_833), .Y(_2187_));
CLKBUFX1 gbuf_d_834(.A(n_1977), .Y(d_out_834));
CLKBUFX1 gbuf_q_834(.A(q_in_834), .Y(WX9944));
CLKBUFX1 gbuf_d_835(.A(n_2353), .Y(d_out_835));
CLKBUFX1 gbuf_q_835(.A(q_in_835), .Y(WX6017));
CLKBUFX1 gbuf_d_836(.A(n_2010), .Y(d_out_836));
CLKBUFX1 gbuf_q_836(.A(q_in_836), .Y(WX3451));
CLKBUFX1 gbuf_d_837(.A(n_2176), .Y(d_out_837));
CLKBUFX1 gbuf_q_837(.A(q_in_837), .Y(WX7190));
CLKBUFX1 gbuf_d_838(.A(n_2110), .Y(d_out_838));
CLKBUFX1 gbuf_q_838(.A(q_in_838), .Y(WX8655));
CLKBUFX1 gbuf_d_839(.A(n_2290), .Y(d_out_839));
CLKBUFX1 gbuf_q_839(.A(q_in_839), .Y(WX7278));
CLKBUFX1 gbuf_d_840(.A(n_1840), .Y(d_out_840));
CLKBUFX1 gbuf_q_840(.A(q_in_840), .Y(WX7232));
CLKBUFX1 gbuf_d_841(.A(n_1671), .Y(d_out_841));
CLKBUFX1 gbuf_q_841(.A(q_in_841), .Y(WX9774));
CLKBUFX1 gbuf_d_842(.A(n_1485), .Y(d_out_842));
CLKBUFX1 gbuf_q_842(.A(q_in_842), .Y(WX8597));
CLKBUFX1 gbuf_d_843(.A(n_2133), .Y(d_out_843));
CLKBUFX1 gbuf_q_843(.A(q_in_843), .Y(WX9860));
CLKBUFX1 gbuf_d_844(.A(n_1791), .Y(d_out_844));
CLKBUFX1 gbuf_q_844(.A(q_in_844), .Y(WX11229));
NOR2X1 g61699(.A (n_2849), .B (n_920), .Y (n_2916));
NOR2X1 g61737(.A (n_2849), .B (n_935), .Y (n_2914));
NOR2X1 g61760(.A (n_2849), .B (n_126), .Y (n_2912));
CLKBUFX1 gbuf_d_845(.A(n_2116), .Y(d_out_845));
CLKBUFX1 gbuf_q_845(.A(q_in_845), .Y(WX8653));
CLKBUFX1 gbuf_d_846(.A(n_1959), .Y(d_out_846));
CLKBUFX1 gbuf_q_846(.A(q_in_846), .Y(WX6053));
NOR2X1 g61771(.A (n_2849), .B (n_85), .Y (n_2911));
CLKBUFX1 gbuf_d_847(.A(n_2363), .Y(d_out_847));
CLKBUFX1 gbuf_q_847(.A(q_in_847), .Y(WX3485));
NOR2X1 g61774(.A (n_2849), .B (n_120), .Y (n_2909));
NOR2X1 g61775(.A (n_2849), .B (n_40), .Y (n_2908));
CLKBUFX1 gbuf_d_848(.A(n_2120), .Y(d_out_848));
CLKBUFX1 gbuf_q_848(.A(q_in_848), .Y(WX9782));
NOR2X1 g61806(.A (n_2849), .B (n_977), .Y (n_2907));
NOR2X1 g61808(.A (n_2849), .B (n_5), .Y (n_2906));
CLKBUFX1 gbuf_d_849(.A(n_2054), .Y(d_out_849));
CLKBUFX1 gbuf_q_849(.A(q_in_849), .Y(WX8619));
CLKBUFX1 gbuf_d_850(.A(n_2057), .Y(d_out_850));
CLKBUFX1 gbuf_q_850(.A(q_in_850), .Y(WX3471));
CLKBUFX1 gbuf_d_851(.A(n_2142), .Y(d_out_851));
CLKBUFX1 gbuf_q_851(.A(q_in_851), .Y(WX6021));
CLKBUFX1 gbuf_d_852(.A(n_2408), .Y(d_out_852));
CLKBUFX1 gbuf_q_852(.A(q_in_852), .Y(WX2100));
CLKBUFX1 gbuf_d_853(.A(n_2258), .Y(d_out_853));
CLKBUFX1 gbuf_q_853(.A(q_in_853), .Y(WX6049));
CLKBUFX1 gbuf_d_854(.A(n_1754), .Y(d_out_854));
CLKBUFX1 gbuf_q_854(.A(q_in_854), .Y(WX2078));
CLKBUFX1 gbuf_d_855(.A(n_2027), .Y(d_out_855));
CLKBUFX1 gbuf_q_855(.A(q_in_855), .Y(WX4666));
CLKBUFX1 gbuf_d_856(.A(n_1620), .Y(d_out_856));
CLKBUFX1 gbuf_q_856(.A(q_in_856), .Y(_2261_));
CLKBUFX1 gbuf_d_857(.A(n_1552), .Y(d_out_857));
CLKBUFX1 gbuf_q_857(.A(q_in_857), .Y(_2300_));
CLKBUFX1 gbuf_d_858(.A(n_1765), .Y(d_out_858));
CLKBUFX1 gbuf_q_858(.A(q_in_858), .Y(WX7236));
CLKBUFX1 gbuf_d_859(.A(n_1590), .Y(d_out_859));
CLKBUFX1 gbuf_q_859(.A(q_in_859), .Y(_2225_));
CLKBUFX1 gbuf_d_860(.A(n_1471), .Y(d_out_860));
CLKBUFX1 gbuf_q_860(.A(q_in_860), .Y(WX5885));
CLKBUFX1 gbuf_d_861(.A(n_2101), .Y(d_out_861));
CLKBUFX1 gbuf_q_861(.A(q_in_861), .Y(WX8623));
NOR2X1 g62112(.A (n_2849), .B (n_927), .Y (n_2905));
NOR2X1 g62114(.A (n_2849), .B (n_924), .Y (n_2903));
CLKBUFX1 gbuf_d_862(.A(n_1738), .Y(d_out_862));
CLKBUFX1 gbuf_q_862(.A(q_in_862), .Y(WX5903));
CLKBUFX1 gbuf_d_863(.A(n_2061), .Y(d_out_863));
CLKBUFX1 gbuf_q_863(.A(q_in_863), .Y(WX4630));
CLKBUFX1 gbuf_d_864(.A(n_2073), .Y(d_out_864));
CLKBUFX1 gbuf_q_864(.A(q_in_864), .Y(WX3399));
CLKBUFX1 gbuf_d_865(.A(n_2394), .Y(d_out_865));
CLKBUFX1 gbuf_q_865(.A(q_in_865), .Y(WX11113));
NOR2X1 g62151(.A (n_2849), .B (n_33), .Y (n_2902));
CLKBUFX1 gbuf_d_866(.A(n_2175), .Y(d_out_866));
CLKBUFX1 gbuf_q_866(.A(q_in_866), .Y(WX6001));
CLKBUFX1 gbuf_d_867(.A(n_1788), .Y(d_out_867));
CLKBUFX1 gbuf_q_867(.A(q_in_867), .Y(WX4592));
CLKBUFX1 gbuf_d_868(.A(n_1787), .Y(d_out_868));
CLKBUFX1 gbuf_q_868(.A(q_in_868), .Y(WX5907));
CLKBUFX1 gbuf_d_869(.A(n_1825), .Y(d_out_869));
CLKBUFX1 gbuf_q_869(.A(q_in_869), .Y(WX5955));
CLKBUFX1 gbuf_d_870(.A(n_1814), .Y(d_out_870));
CLKBUFX1 gbuf_q_870(.A(q_in_870), .Y(WX2082));
CLKBUFX1 gbuf_d_871(.A(n_2117), .Y(d_out_871));
CLKBUFX1 gbuf_q_871(.A(q_in_871), .Y(WX2074));
CLKBUFX1 gbuf_d_872(.A(n_1710), .Y(d_out_872));
CLKBUFX1 gbuf_q_872(.A(q_in_872), .Y(WX8591));
CLKBUFX1 gbuf_d_873(.A(n_1813), .Y(d_out_873));
CLKBUFX1 gbuf_q_873(.A(q_in_873), .Y(WX8567));
CLKBUFX1 gbuf_d_874(.A(n_2160), .Y(d_out_874));
CLKBUFX1 gbuf_q_874(.A(q_in_874), .Y(WX3419));
CLKBUFX1 gbuf_d_875(.A(n_2559), .Y(d_out_875));
CLKBUFX1 gbuf_q_875(.A(q_in_875), .Y(WX7302));
CLKBUFX1 gbuf_d_876(.A(n_1873), .Y(d_out_876));
CLKBUFX1 gbuf_q_876(.A(q_in_876), .Y(WX8565));
CLKBUFX1 gbuf_d_877(.A(n_2068), .Y(d_out_877));
CLKBUFX1 gbuf_q_877(.A(q_in_877), .Y(WX9902));
BUFX3 g62443(.A (n_7086), .Y (n_3183));
CLKBUFX1 gbuf_d_878(.A(n_1883), .Y(d_out_878));
CLKBUFX1 gbuf_q_878(.A(q_in_878), .Y(WX4588));
CLKBUFX1 gbuf_d_879(.A(n_1955), .Y(d_out_879));
CLKBUFX1 gbuf_q_879(.A(q_in_879), .Y(WX9820));
CLKBUFX1 gbuf_d_880(.A(n_2442), .Y(d_out_880));
CLKBUFX1 gbuf_q_880(.A(q_in_880), .Y(WX8539));
CLKBUFX1 gbuf_d_881(.A(n_1483), .Y(d_out_881));
CLKBUFX1 gbuf_q_881(.A(q_in_881), .Y(WX11109));
CLKBUFX1 gbuf_d_882(.A(n_2369), .Y(d_out_882));
CLKBUFX1 gbuf_q_882(.A(q_in_882), .Y(WX8537));
CLKBUFX1 gbuf_d_883(.A(n_1878), .Y(d_out_883));
CLKBUFX1 gbuf_q_883(.A(q_in_883), .Y(WX5979));
CLKBUFX1 gbuf_d_884(.A(n_2167), .Y(d_out_884));
CLKBUFX1 gbuf_q_884(.A(q_in_884), .Y(WX3347));
CLKBUFX1 gbuf_d_885(.A(n_2074), .Y(d_out_885));
CLKBUFX1 gbuf_q_885(.A(q_in_885), .Y(WX4750));
CLKBUFX1 gbuf_d_886(.A(n_1833), .Y(d_out_886));
CLKBUFX1 gbuf_q_886(.A(q_in_886), .Y(WX8467));
CLKBUFX1 gbuf_d_887(.A(n_2136), .Y(d_out_887));
CLKBUFX1 gbuf_q_887(.A(q_in_887), .Y(WX5931));
CLKBUFX1 gbuf_d_888(.A(n_1875), .Y(d_out_888));
CLKBUFX1 gbuf_q_888(.A(q_in_888), .Y(WX8501));
NOR2X1 g62618(.A (n_2825), .B (n_2849), .Y (n_2900));
CLKBUFX1 gbuf_d_889(.A(n_1993), .Y(d_out_889));
CLKBUFX1 gbuf_q_889(.A(q_in_889), .Y(WX3295));
CLKBUFX1 gbuf_d_890(.A(n_1668), .Y(d_out_890));
CLKBUFX1 gbuf_q_890(.A(q_in_890), .Y(_2111_));
CLKBUFX1 gbuf_d_891(.A(n_2228), .Y(d_out_891));
CLKBUFX1 gbuf_q_891(.A(q_in_891), .Y(WX3319));
CLKBUFX1 gbuf_d_892(.A(n_1534), .Y(d_out_892));
CLKBUFX1 gbuf_q_892(.A(q_in_892), .Y(_2336_));
CLKBUFX1 gbuf_d_893(.A(n_1644), .Y(d_out_893));
CLKBUFX1 gbuf_q_893(.A(q_in_893), .Y(_2147_));
CLKBUFX1 gbuf_d_894(.A(n_1665), .Y(d_out_894));
CLKBUFX1 gbuf_q_894(.A(q_in_894), .Y(_2114_));
CLKBUFX1 gbuf_d_895(.A(n_2123), .Y(d_out_895));
CLKBUFX1 gbuf_q_895(.A(q_in_895), .Y(WX4726));
CLKBUFX1 gbuf_d_896(.A(n_2053), .Y(d_out_896));
CLKBUFX1 gbuf_q_896(.A(q_in_896), .Y(WX3359));
CLKBUFX1 gbuf_d_897(.A(n_2147), .Y(d_out_897));
CLKBUFX1 gbuf_q_897(.A(q_in_897), .Y(WX4634));
CLKBUFX1 gbuf_d_898(.A(n_1996), .Y(d_out_898));
CLKBUFX1 gbuf_q_898(.A(q_in_898), .Y(WX4682));
CLKBUFX1 gbuf_d_899(.A(n_1481), .Y(d_out_899));
CLKBUFX1 gbuf_q_899(.A(q_in_899), .Y(WX11105));
CLKBUFX1 gbuf_d_900(.A(n_2113), .Y(d_out_900));
CLKBUFX1 gbuf_q_900(.A(q_in_900), .Y(WX3307));
CLKBUFX1 gbuf_d_901(.A(n_1837), .Y(d_out_901));
CLKBUFX1 gbuf_q_901(.A(q_in_901), .Y(WX3313));
CLKBUFX1 gbuf_d_902(.A(n_2141), .Y(d_out_902));
CLKBUFX1 gbuf_q_902(.A(q_in_902), .Y(WX3351));
CLKBUFX1 gbuf_d_903(.A(n_1531), .Y(d_out_903));
CLKBUFX1 gbuf_q_903(.A(q_in_903), .Y(_2339_));
CLKBUFX1 gbuf_d_904(.A(n_1989), .Y(d_out_904));
CLKBUFX1 gbuf_q_904(.A(q_in_904), .Y(WX3431));
CLKBUFX1 gbuf_d_905(.A(n_1896), .Y(d_out_905));
CLKBUFX1 gbuf_q_905(.A(q_in_905), .Y(WX3379));
CLKBUFX1 gbuf_d_906(.A(n_2095), .Y(d_out_906));
CLKBUFX1 gbuf_q_906(.A(q_in_906), .Y(WX3299));
CLKBUFX1 gbuf_d_907(.A(n_2109), .Y(d_out_907));
CLKBUFX1 gbuf_q_907(.A(q_in_907), .Y(WX3303));
CLKBUFX1 gbuf_d_908(.A(n_1717), .Y(d_out_908));
CLKBUFX1 gbuf_q_908(.A(q_in_908), .Y(WX3355));
CLKBUFX1 gbuf_d_909(.A(n_1650), .Y(d_out_909));
CLKBUFX1 gbuf_q_909(.A(q_in_909), .Y(_2138_));
CLKBUFX1 gbuf_d_910(.A(n_1877), .Y(d_out_910));
CLKBUFX1 gbuf_q_910(.A(q_in_910), .Y(WX8559));
CLKBUFX1 gbuf_d_911(.A(n_2127), .Y(d_out_911));
CLKBUFX1 gbuf_q_911(.A(q_in_911), .Y(WX3459));
CLKBUFX1 gbuf_d_912(.A(n_1958), .Y(d_out_912));
CLKBUFX1 gbuf_q_912(.A(q_in_912), .Y(WX6057));
CLKBUFX1 gbuf_d_913(.A(n_1969), .Y(d_out_913));
CLKBUFX1 gbuf_q_913(.A(q_in_913), .Y(WX8531));
CLKBUFX1 gbuf_d_914(.A(n_1762), .Y(d_out_914));
CLKBUFX1 gbuf_q_914(.A(q_in_914), .Y(WX8579));
CLKBUFX1 gbuf_d_915(.A(n_2111), .Y(d_out_915));
CLKBUFX1 gbuf_q_915(.A(q_in_915), .Y(WX4762));
CLKBUFX1 gbuf_d_916(.A(n_1693), .Y(d_out_916));
CLKBUFX1 gbuf_q_916(.A(q_in_916), .Y(_2219_));
CLKBUFX1 gbuf_d_917(.A(n_1792), .Y(d_out_917));
CLKBUFX1 gbuf_q_917(.A(q_in_917), .Y(WX7248));
CLKBUFX1 gbuf_d_918(.A(n_1991), .Y(d_out_918));
CLKBUFX1 gbuf_q_918(.A(q_in_918), .Y(WX8589));
CLKBUFX1 gbuf_d_919(.A(n_2274), .Y(d_out_919));
CLKBUFX1 gbuf_q_919(.A(q_in_919), .Y(WX4626));
CLKBUFX1 gbuf_d_920(.A(n_1647), .Y(d_out_920));
CLKBUFX1 gbuf_q_920(.A(q_in_920), .Y(_2142_));
CLKBUFX1 gbuf_d_921(.A(n_1491), .Y(d_out_921));
CLKBUFX1 gbuf_q_921(.A(q_in_921), .Y(WX7262));
CLKBUFX1 gbuf_d_922(.A(n_1498), .Y(d_out_922));
CLKBUFX1 gbuf_q_922(.A(q_in_922), .Y(_2252_));
CLKBUFX1 gbuf_d_923(.A(n_2070), .Y(d_out_923));
CLKBUFX1 gbuf_q_923(.A(q_in_923), .Y(WX9852));
CLKBUFX1 gbuf_d_924(.A(n_1517), .Y(d_out_924));
CLKBUFX1 gbuf_q_924(.A(q_in_924), .Y(_2361_));
CLKBUFX1 gbuf_d_925(.A(n_1670), .Y(d_out_925));
CLKBUFX1 gbuf_q_925(.A(q_in_925), .Y(_2109_));
CLKBUFX1 gbuf_d_926(.A(n_2170), .Y(d_out_926));
CLKBUFX1 gbuf_q_926(.A(q_in_926), .Y(WX9806));
CLKBUFX1 gbuf_d_927(.A(n_2356), .Y(d_out_927));
CLKBUFX1 gbuf_q_927(.A(q_in_927), .Y(WX7268));
NOR2X1 g57537(.A (n_1473), .B (n_5181), .Y (n_2898));
CLKBUFX1 gbuf_d_928(.A(n_1593), .Y(d_out_928));
CLKBUFX1 gbuf_q_928(.A(q_in_928), .Y(_2215_));
CLKBUFX1 gbuf_d_929(.A(n_2134), .Y(d_out_929));
CLKBUFX1 gbuf_q_929(.A(q_in_929), .Y(WX7180));
CLKBUFX1 gbuf_d_930(.A(n_1980), .Y(d_out_930));
CLKBUFX1 gbuf_q_930(.A(q_in_930), .Y(WX7364));
BUFX3 g63072(.A (n_4562), .Y (n_4593));
CLKBUFX1 gbuf_d_931(.A(n_2390), .Y(d_out_931));
CLKBUFX1 gbuf_q_931(.A(q_in_931), .Y(WX9940));
BUFX3 g63075(.A (n_4562), .Y (n_4644));
BUFX3 g63080(.A (n_6626), .Y (n_4096));
CLKBUFX1 gbuf_d_932(.A(n_1550), .Y(d_out_932));
CLKBUFX1 gbuf_q_932(.A(q_in_932), .Y(_2313_));
CLKBUFX1 gbuf_d_933(.A(n_2071), .Y(d_out_933));
CLKBUFX1 gbuf_q_933(.A(q_in_933), .Y(WX9894));
BUFX3 g63147(.A (n_3162), .Y (n_3225));
INVX4 g63153(.A (n_2897), .Y (n_5965));
INVX4 g63155(.A (n_2897), .Y (n_6091));
BUFX3 g63159(.A (n_6437), .Y (n_4184));
BUFX3 g63181(.A (n_6437), .Y (n_5828));
BUFX3 g63187(.A (n_6452), .Y (n_4099));
BUFX3 g63215(.A (n_2894), .Y (n_4078));
BUFX3 g63217(.A (n_2894), .Y (n_4016));
CLKBUFX1 gbuf_d_934(.A(n_2243), .Y(d_out_934));
CLKBUFX1 gbuf_q_934(.A(q_in_934), .Y(WX6061));
CLKBUFX1 gbuf_d_935(.A(n_2277), .Y(d_out_935));
CLKBUFX1 gbuf_q_935(.A(q_in_935), .Y(WX9836));
CLKBUFX1 gbuf_d_936(.A(n_1912), .Y(d_out_936));
CLKBUFX1 gbuf_q_936(.A(q_in_936), .Y(WX6033));
CLKBUFX1 gbuf_d_937(.A(n_1920), .Y(d_out_937));
CLKBUFX1 gbuf_q_937(.A(q_in_937), .Y(WX6041));
CLKBUFX1 gbuf_d_938(.A(n_1797), .Y(d_out_938));
CLKBUFX1 gbuf_q_938(.A(q_in_938), .Y(WX6037));
CLKBUFX1 gbuf_d_939(.A(n_1990), .Y(d_out_939));
CLKBUFX1 gbuf_q_939(.A(q_in_939), .Y(WX11223));
CLKBUFX1 gbuf_d_940(.A(n_1724), .Y(d_out_940));
CLKBUFX1 gbuf_q_940(.A(q_in_940), .Y(WX8545));
CLKBUFX1 gbuf_d_941(.A(n_2182), .Y(d_out_941));
CLKBUFX1 gbuf_q_941(.A(q_in_941), .Y(WX7184));
CLKBUFX1 gbuf_d_942(.A(n_1489), .Y(d_out_942));
CLKBUFX1 gbuf_q_942(.A(q_in_942), .Y(WX7326));
CLKBUFX1 gbuf_d_943(.A(n_1617), .Y(d_out_943));
CLKBUFX1 gbuf_q_943(.A(q_in_943), .Y(_2180_));
CLKBUFX1 gbuf_d_944(.A(n_1848), .Y(d_out_944));
CLKBUFX1 gbuf_q_944(.A(q_in_944), .Y(WX9798));
NOR2X1 g59247(.A (n_2535), .B (n_1648), .Y (n_2893));
NOR2X1 g59258(.A (n_1235), .B (n_2605), .Y (n_2892));
CLKBUFX1 gbuf_d_945(.A(n_2276), .Y(d_out_945));
CLKBUFX1 gbuf_q_945(.A(q_in_945), .Y(WX11187));
CLKBUFX1 gbuf_d_946(.A(n_1772), .Y(d_out_946));
CLKBUFX1 gbuf_q_946(.A(q_in_946), .Y(WX8523));
NOR2X1 g59262(.A (n_1026), .B (n_2849), .Y (n_2889));
INVX1 g55889(.A (WX487), .Y (n_2888));
CLKBUFX1 gbuf_d_947(.A(n_2364), .Y(d_out_947));
CLKBUFX1 gbuf_q_947(.A(q_in_947), .Y(WX7224));
CLKBUFX1 gbuf_d_948(.A(n_1504), .Y(d_out_948));
CLKBUFX1 gbuf_q_948(.A(q_in_948), .Y(_2129_));
CLKBUFX1 gbuf_d_949(.A(n_2350), .Y(d_out_949));
CLKBUFX1 gbuf_q_949(.A(q_in_949), .Y(WX7228));
CLKBUFX1 gbuf_d_950(.A(n_1719), .Y(d_out_950));
CLKBUFX1 gbuf_q_950(.A(q_in_950), .Y(WX7270));
NOR2X1 g59268(.A (n_2546), .B (n_1648), .Y (n_2887));
NOR2X1 g59269(.A (n_2523), .B (n_1425), .Y (n_2885));
NOR2X1 g59270(.A (n_2545), .B (n_1425), .Y (n_2884));
NOR2X1 g59271(.A (n_2524), .B (n_5181), .Y (n_2883));
CLKBUFX1 gbuf_d_951(.A(n_2154), .Y(d_out_951));
CLKBUFX1 gbuf_q_951(.A(q_in_951), .Y(WX4700));
NOR2X1 g59272(.A (n_2517), .B (n_1425), .Y (n_2882));
CLKBUFX1 gbuf_d_952(.A(n_1784), .Y(d_out_952));
CLKBUFX1 gbuf_q_952(.A(q_in_952), .Y(WX5899));
NOR2X1 g59273(.A (n_2519), .B (n_1425), .Y (n_2881));
NOR2X1 g59274(.A (n_2542), .B (n_1425), .Y (n_2879));
NOR2X1 g59275(.A (n_2541), .B (n_5181), .Y (n_2878));
NOR2X1 g59276(.A (n_2539), .B (n_2849), .Y (n_2876));
NOR2X1 g59277(.A (n_2516), .B (n_1425), .Y (n_2875));
NOR2X1 g59278(.A (n_2551), .B (n_2849), .Y (n_2873));
NOR2X1 g59279(.A (n_2536), .B (n_1425), .Y (n_2872));
NOR2X1 g59280(.A (n_2518), .B (n_5181), .Y (n_2870));
NOR2X1 g59281(.A (n_2547), .B (n_1425), .Y (n_2868));
NOR2X1 g59282(.A (n_2557), .B (n_1425), .Y (n_2867));
NOR2X1 g59283(.A (n_2532), .B (n_1425), .Y (n_2866));
NOR2X1 g59284(.A (n_2548), .B (n_2849), .Y (n_2865));
CLKBUFX1 gbuf_d_953(.A(n_1721), .Y(d_out_953));
CLKBUFX1 gbuf_q_953(.A(q_in_953), .Y(WX7274));
NOR2X1 g59285(.A (n_2531), .B (n_5712), .Y (n_2864));
NOR2X1 g59286(.A (n_2552), .B (n_5712), .Y (n_2863));
NOR2X1 g59293(.A (n_1029), .B (n_2605), .Y (n_2861));
CLKBUFX1 gbuf_d_954(.A(n_1563), .Y(d_out_954));
CLKBUFX1 gbuf_q_954(.A(q_in_954), .Y(_2277_));
CLKBUFX1 gbuf_d_955(.A(n_2151), .Y(d_out_955));
CLKBUFX1 gbuf_q_955(.A(q_in_955), .Y(WX9936));
CLKBUFX1 gbuf_d_956(.A(n_2248), .Y(d_out_956));
CLKBUFX1 gbuf_q_956(.A(q_in_956), .Y(WX5987));
CLKBUFX1 gbuf_d_957(.A(n_2226), .Y(d_out_957));
CLKBUFX1 gbuf_qn_957(.A(qn_in_957), .Y(WX2130));
NOR2X1 g59338(.A (n_1167), .B (n_2605), .Y (n_2860));
NOR2X1 g59339(.A (n_1234), .B (n_2605), .Y (n_2859));
CLKBUFX1 gbuf_d_958(.A(n_2553), .Y(d_out_958));
CLKBUFX1 gbuf_q_958(.A(q_in_958), .Y(WX11159));
CLKBUFX1 gbuf_d_959(.A(n_1741), .Y(d_out_959));
CLKBUFX1 gbuf_q_959(.A(q_in_959), .Y(WX3375));
CLKBUFX1 gbuf_d_960(.A(n_2322), .Y(d_out_960));
CLKBUFX1 gbuf_q_960(.A(q_in_960), .Y(WX3443));
CLKBUFX1 gbuf_d_961(.A(n_1785), .Y(d_out_961));
CLKBUFX1 gbuf_q_961(.A(q_in_961), .Y(WX7318));
CLKBUFX1 gbuf_d_962(.A(n_1961), .Y(d_out_962));
CLKBUFX1 gbuf_q_962(.A(q_in_962), .Y(WX8585));
CLKBUFX1 gbuf_d_963(.A(n_2107), .Y(d_out_963));
CLKBUFX1 gbuf_q_963(.A(q_in_963), .Y(WX8647));
CLKBUFX1 gbuf_d_964(.A(n_2062), .Y(d_out_964));
CLKBUFX1 gbuf_q_964(.A(q_in_964), .Y(WX9760));
CLKBUFX1 gbuf_d_965(.A(n_2020), .Y(d_out_965));
CLKBUFX1 gbuf_q_965(.A(q_in_965), .Y(WX5963));
CLKBUFX1 gbuf_d_966(.A(n_2046), .Y(d_out_966));
CLKBUFX1 gbuf_q_966(.A(q_in_966), .Y(WX8617));
CLKBUFX1 gbuf_d_967(.A(n_2173), .Y(d_out_967));
CLKBUFX1 gbuf_q_967(.A(q_in_967), .Y(WX3411));
NOR2X1 g59396(.A (n_1121), .B (n_2849), .Y (n_2858));
NOR2X1 g59397(.A (n_1222), .B (n_2849), .Y (n_2857));
CLKBUFX1 gbuf_d_968(.A(n_2344), .Y(d_out_968));
CLKBUFX1 gbuf_q_968(.A(q_in_968), .Y(WX5993));
CLKBUFX1 gbuf_d_969(.A(n_2148), .Y(d_out_969));
CLKBUFX1 gbuf_q_969(.A(q_in_969), .Y(WX8611));
CLKBUFX1 gbuf_d_970(.A(n_2366), .Y(d_out_970));
CLKBUFX1 gbuf_q_970(.A(q_in_970), .Y(WX11157));
CLKBUFX1 gbuf_d_971(.A(n_2528), .Y(d_out_971));
CLKBUFX1 gbuf_q_971(.A(q_in_971), .Y(WX11145));
CLKBUFX1 gbuf_d_972(.A(n_1820), .Y(d_out_972));
CLKBUFX1 gbuf_q_972(.A(q_in_972), .Y(WX9848));
CLKBUFX1 gbuf_d_973(.A(n_2285), .Y(d_out_973));
CLKBUFX1 gbuf_q_973(.A(q_in_973), .Y(WX11171));
CLKBUFX1 gbuf_d_974(.A(n_1898), .Y(d_out_974));
CLKBUFX1 gbuf_q_974(.A(q_in_974), .Y(WX7176));
CLKBUFX1 gbuf_d_975(.A(n_1507), .Y(d_out_975));
CLKBUFX1 gbuf_q_975(.A(q_in_975), .Y(_2257_));
CLKBUFX1 gbuf_d_976(.A(n_1540), .Y(d_out_976));
CLKBUFX1 gbuf_q_976(.A(q_in_976), .Y(_2324_));
CLKBUFX1 gbuf_d_977(.A(n_1535), .Y(d_out_977));
CLKBUFX1 gbuf_q_977(.A(q_in_977), .Y(_2330_));
NOR2X1 g59466(.A (n_2521), .B (n_5712), .Y (n_2856));
NOR2X1 g59467(.A (n_2555), .B (n_5712), .Y (n_2855));
CLKBUFX1 gbuf_d_978(.A(n_2391), .Y(d_out_978));
CLKBUFX1 gbuf_q_978(.A(q_in_978), .Y(WX9766));
NOR2X1 g59470(.A (n_2533), .B (n_5181), .Y (n_2854));
CLKBUFX1 gbuf_d_979(.A(n_1690), .Y(d_out_979));
CLKBUFX1 gbuf_q_979(.A(q_in_979), .Y(_2297_));
CLKBUFX1 gbuf_d_980(.A(n_1889), .Y(d_out_980));
CLKBUFX1 gbuf_q_980(.A(q_in_980), .Y(WX9802));
NOR2X1 g59479(.A (n_2538), .B (n_2851), .Y (n_2852));
NOR2X1 g59480(.A (n_2543), .B (n_2849), .Y (n_2850));
NOR2X1 g59481(.A (n_1043), .B (n_2849), .Y (n_2848));
CLKBUFX1 gbuf_d_981(.A(n_2064), .Y(d_out_981));
CLKBUFX1 gbuf_q_981(.A(q_in_981), .Y(WX7360));
NOR2X1 g59482(.A (n_1042), .B (n_2849), .Y (n_2847));
CLKBUFX1 gbuf_d_982(.A(n_1838), .Y(d_out_982));
CLKBUFX1 gbuf_q_982(.A(q_in_982), .Y(WX5971));
CLKBUFX1 gbuf_d_983(.A(n_1537), .Y(d_out_983));
CLKBUFX1 gbuf_q_983(.A(q_in_983), .Y(_2326_));
NOR2X1 g59488(.A (n_2522), .B (n_5712), .Y (n_2846));
NOR2X1 g59491(.A (n_2520), .B (n_1648), .Y (n_2844));
NOR2X1 g59494(.A (n_2554), .B (n_5712), .Y (n_2843));
CLKBUFX1 gbuf_d_984(.A(n_1555), .Y(d_out_984));
CLKBUFX1 gbuf_q_984(.A(q_in_984), .Y(_2290_));
CLKBUFX1 gbuf_d_985(.A(n_2281), .Y(d_out_985));
CLKBUFX1 gbuf_q_985(.A(q_in_985), .Y(WX3425));
CLKBUFX1 gbuf_d_986(.A(n_1554), .Y(d_out_986));
CLKBUFX1 gbuf_q_986(.A(q_in_986), .Y(_2291_));
CLKBUFX1 gbuf_d_987(.A(n_1729), .Y(d_out_987));
CLKBUFX1 gbuf_q_987(.A(q_in_987), .Y(WX8645));
CLKBUFX1 gbuf_d_988(.A(n_2041), .Y(d_out_988));
CLKBUFX1 gbuf_q_988(.A(q_in_988), .Y(WX8527));
CLKBUFX1 gbuf_d_989(.A(n_1681), .Y(d_out_989));
CLKBUFX1 gbuf_q_989(.A(q_in_989), .Y(_2255_));
CLKBUFX1 gbuf_d_990(.A(n_2308), .Y(d_out_990));
CLKBUFX1 gbuf_q_990(.A(q_in_990), .Y(WX6009));
CLKBUFX1 gbuf_d_991(.A(n_2241), .Y(d_out_991));
CLKBUFX1 gbuf_q_991(.A(q_in_991), .Y(WX3323));
CLKBUFX1 gbuf_d_992(.A(n_1654), .Y(d_out_992));
CLKBUFX1 gbuf_q_992(.A(q_in_992), .Y(_2133_));
CLKBUFX1 gbuf_d_993(.A(n_1508), .Y(d_out_993));
CLKBUFX1 gbuf_q_993(.A(q_in_993), .Y(_2247_));
CLKBUFX1 gbuf_d_994(.A(n_1559), .Y(d_out_994));
CLKBUFX1 gbuf_q_994(.A(q_in_994), .Y(_2283_));
CLKBUFX1 gbuf_d_995(.A(n_1575), .Y(d_out_995));
CLKBUFX1 gbuf_q_995(.A(q_in_995), .Y(_2251_));
CLKBUFX1 gbuf_d_996(.A(n_1514), .Y(d_out_996));
CLKBUFX1 gbuf_q_996(.A(q_in_996), .Y(_2137_));
CLKBUFX1 gbuf_d_997(.A(n_1496), .Y(d_out_997));
CLKBUFX1 gbuf_q_997(.A(q_in_997), .Y(_2199_));
CLKBUFX1 gbuf_d_998(.A(n_2331), .Y(d_out_998));
CLKBUFX1 gbuf_q_998(.A(q_in_998), .Y(WX3341));
CLKBUFX1 gbuf_d_999(.A(n_1545), .Y(d_out_999));
CLKBUFX1 gbuf_q_999(.A(q_in_999), .Y(_2320_));
CLKBUFX1 gbuf_d_1000(.A(n_2303), .Y(d_out_1000));
CLKBUFX1 gbuf_q_1000(.A(q_in_1000), .Y(WX8487));
CLKBUFX1 gbuf_d_1001(.A(n_1984), .Y(d_out_1001));
CLKBUFX1 gbuf_q_1001(.A(q_in_1001), .Y(WX8477));
CLKBUFX1 gbuf_d_1002(.A(n_2166), .Y(d_out_1002));
CLKBUFX1 gbuf_q_1002(.A(q_in_1002), .Y(WX8511));
CLKBUFX1 gbuf_d_1003(.A(n_1493), .Y(d_out_1003));
CLKBUFX1 gbuf_q_1003(.A(q_in_1003), .Y(WX2066));
CLKBUFX1 gbuf_d_1004(.A(n_2264), .Y(d_out_1004));
CLKBUFX1 gbuf_q_1004(.A(q_in_1004), .Y(WX7254));
CLKBUFX1 gbuf_d_1005(.A(n_2270), .Y(d_out_1005));
CLKBUFX1 gbuf_q_1005(.A(q_in_1005), .Y(WX5939));
CLKBUFX1 gbuf_d_1006(.A(n_1725), .Y(d_out_1006));
CLKBUFX1 gbuf_q_1006(.A(q_in_1006), .Y(WX8639));
CLKBUFX1 gbuf_d_1007(.A(n_1847), .Y(d_out_1007));
CLKBUFX1 gbuf_q_1007(.A(q_in_1007), .Y(WX5947));
CLKBUFX1 gbuf_d_1008(.A(n_2207), .Y(d_out_1008));
CLKBUFX1 gbuf_q_1008(.A(q_in_1008), .Y(WX9906));
CLKBUFX1 gbuf_d_1009(.A(n_2221), .Y(d_out_1009));
CLKBUFX1 gbuf_q_1009(.A(q_in_1009), .Y(WX8513));
CLKBUFX1 gbuf_d_1010(.A(n_2309), .Y(d_out_1010));
CLKBUFX1 gbuf_q_1010(.A(q_in_1010), .Y(WX3337));
CLKBUFX1 gbuf_d_1011(.A(n_1972), .Y(d_out_1011));
CLKBUFX1 gbuf_q_1011(.A(q_in_1011), .Y(WX8475));
CLKBUFX1 gbuf_d_1012(.A(n_1580), .Y(d_out_1012));
CLKBUFX1 gbuf_q_1012(.A(q_in_1012), .Y(_2239_));
CLKBUFX1 gbuf_d_1013(.A(n_2132), .Y(d_out_1013));
CLKBUFX1 gbuf_q_1013(.A(q_in_1013), .Y(WX9840));
CLKBUFX1 gbuf_d_1014(.A(n_1924), .Y(d_out_1014));
CLKBUFX1 gbuf_q_1014(.A(q_in_1014), .Y(WX4600));
CLKBUFX1 gbuf_d_1015(.A(n_1925), .Y(d_out_1015));
CLKBUFX1 gbuf_q_1015(.A(q_in_1015), .Y(WX4670));
CLKBUFX1 gbuf_d_1016(.A(n_2399), .Y(d_out_1016));
CLKBUFX1 gbuf_q_1016(.A(q_in_1016), .Y(WX7316));
CLKBUFX1 gbuf_d_1017(.A(n_1992), .Y(d_out_1017));
CLKBUFX1 gbuf_q_1017(.A(q_in_1017), .Y(WX8553));
CLKBUFX1 gbuf_d_1018(.A(n_2393), .Y(d_out_1018));
CLKBUFX1 gbuf_q_1018(.A(q_in_1018), .Y(WX11101));
CLKBUFX1 gbuf_d_1019(.A(n_1732), .Y(d_out_1019));
CLKBUFX1 gbuf_q_1019(.A(q_in_1019), .Y(WX3333));
CLKBUFX1 gbuf_d_1020(.A(n_2452), .Y(d_out_1020));
CLKBUFX1 gbuf_q_1020(.A(q_in_1020), .Y(WX10829));
CLKBUFX1 gbuf_d_1021(.A(n_2036), .Y(d_out_1021));
CLKBUFX1 gbuf_q_1021(.A(q_in_1021), .Y(WX5923));
CLKBUFX1 gbuf_d_1022(.A(n_2096), .Y(d_out_1022));
CLKBUFX1 gbuf_q_1022(.A(q_in_1022), .Y(WX8519));
CLKBUFX1 gbuf_d_1023(.A(n_1856), .Y(d_out_1023));
CLKBUFX1 gbuf_q_1023(.A(q_in_1023), .Y(WX8551));
CLKBUFX1 gbuf_d_1024(.A(n_1519), .Y(d_out_1024));
CLKBUFX1 gbuf_q_1024(.A(q_in_1024), .Y(_2359_));
CLKBUFX1 gbuf_d_1025(.A(n_2237), .Y(d_out_1025));
CLKBUFX1 gbuf_q_1025(.A(q_in_1025), .Y(WX7344));
CLKBUFX1 gbuf_d_1026(.A(n_1901), .Y(d_out_1026));
CLKBUFX1 gbuf_q_1026(.A(q_in_1026), .Y(WX7352));
CLKBUFX1 gbuf_d_1027(.A(n_1696), .Y(d_out_1027));
CLKBUFX1 gbuf_q_1027(.A(q_in_1027), .Y(_2170_));
CLKBUFX1 gbuf_d_1028(.A(n_2337), .Y(d_out_1028));
CLKBUFX1 gbuf_q_1028(.A(q_in_1028), .Y(WX7296));
CLKBUFX1 gbuf_d_1029(.A(n_1624), .Y(d_out_1029));
CLKBUFX1 gbuf_q_1029(.A(q_in_1029), .Y(_2172_));
CLKBUFX1 gbuf_d_1030(.A(n_2206), .Y(d_out_1030));
CLKBUFX1 gbuf_q_1030(.A(q_in_1030), .Y(WX7212));
CLKBUFX1 gbuf_d_1031(.A(n_1676), .Y(d_out_1031));
CLKBUFX1 gbuf_q_1031(.A(q_in_1031), .Y(_2210_));
CLKBUFX1 gbuf_d_1032(.A(n_1594), .Y(d_out_1032));
CLKBUFX1 gbuf_q_1032(.A(q_in_1032), .Y(_2214_));
CLKBUFX1 gbuf_d_1033(.A(n_1818), .Y(d_out_1033));
CLKBUFX1 gbuf_q_1033(.A(q_in_1033), .Y(WX2116));
CLKBUFX1 gbuf_d_1034(.A(n_2011), .Y(d_out_1034));
CLKBUFX1 gbuf_q_1034(.A(q_in_1034), .Y(WX2070));
CLKBUFX1 gbuf_d_1035(.A(n_1935), .Y(d_out_1035));
CLKBUFX1 gbuf_q_1035(.A(q_in_1035), .Y(WX2184));
CLKBUFX1 gbuf_d_1036(.A(n_1522), .Y(d_out_1036));
CLKBUFX1 gbuf_q_1036(.A(q_in_1036), .Y(_2357_));
CLKBUFX1 gbuf_d_1037(.A(n_1623), .Y(d_out_1037));
CLKBUFX1 gbuf_q_1037(.A(q_in_1037), .Y(_2173_));
CLKBUFX1 gbuf_d_1038(.A(n_1673), .Y(d_out_1038));
CLKBUFX1 gbuf_q_1038(.A(q_in_1038), .Y(_2294_));
CLKBUFX1 gbuf_d_1039(.A(n_1706), .Y(d_out_1039));
CLKBUFX1 gbuf_q_1039(.A(q_in_1039), .Y(_2364_));
CLKBUFX1 gbuf_d_1040(.A(n_1622), .Y(d_out_1040));
CLKBUFX1 gbuf_q_1040(.A(q_in_1040), .Y(_2176_));
CLKBUFX1 gbuf_d_1041(.A(n_1579), .Y(d_out_1041));
CLKBUFX1 gbuf_q_1041(.A(q_in_1041), .Y(_2243_));
CLKBUFX1 gbuf_d_1042(.A(n_1495), .Y(d_out_1042));
CLKBUFX1 gbuf_q_1042(.A(q_in_1042), .Y(WX11117));
CLKBUFX1 gbuf_d_1043(.A(n_1669), .Y(d_out_1043));
CLKBUFX1 gbuf_q_1043(.A(q_in_1043), .Y(_2110_));
CLKBUFX1 gbuf_d_1044(.A(n_1666), .Y(d_out_1044));
CLKBUFX1 gbuf_q_1044(.A(q_in_1044), .Y(_2112_));
CLKBUFX1 gbuf_d_1045(.A(n_1512), .Y(d_out_1045));
CLKBUFX1 gbuf_q_1045(.A(q_in_1045), .Y(_2116_));
CLKBUFX1 gbuf_d_1046(.A(n_1664), .Y(d_out_1046));
CLKBUFX1 gbuf_q_1046(.A(q_in_1046), .Y(_2115_));
CLKBUFX1 gbuf_d_1047(.A(n_1662), .Y(d_out_1047));
CLKBUFX1 gbuf_q_1047(.A(q_in_1047), .Y(_2122_));
CLKBUFX1 gbuf_d_1048(.A(n_1661), .Y(d_out_1048));
CLKBUFX1 gbuf_q_1048(.A(q_in_1048), .Y(_2123_));
CLKBUFX1 gbuf_d_1049(.A(n_1659), .Y(d_out_1049));
CLKBUFX1 gbuf_q_1049(.A(q_in_1049), .Y(_2126_));
CLKBUFX1 gbuf_d_1050(.A(n_1656), .Y(d_out_1050));
CLKBUFX1 gbuf_q_1050(.A(q_in_1050), .Y(_2128_));
CLKBUFX1 gbuf_d_1051(.A(n_1516), .Y(d_out_1051));
CLKBUFX1 gbuf_q_1051(.A(q_in_1051), .Y(_2130_));
CLKBUFX1 gbuf_d_1052(.A(n_1655), .Y(d_out_1052));
CLKBUFX1 gbuf_q_1052(.A(q_in_1052), .Y(_2132_));
CLKBUFX1 gbuf_d_1053(.A(n_1652), .Y(d_out_1053));
CLKBUFX1 gbuf_q_1053(.A(q_in_1053), .Y(_2134_));
CLKBUFX1 gbuf_d_1054(.A(n_1651), .Y(d_out_1054));
CLKBUFX1 gbuf_q_1054(.A(q_in_1054), .Y(_2136_));
CLKBUFX1 gbuf_d_1055(.A(n_1682), .Y(d_out_1055));
CLKBUFX1 gbuf_q_1055(.A(q_in_1055), .Y(_2141_));
CLKBUFX1 gbuf_d_1056(.A(n_1646), .Y(d_out_1056));
CLKBUFX1 gbuf_q_1056(.A(q_in_1056), .Y(_2143_));
CLKBUFX1 gbuf_d_1057(.A(n_1697), .Y(d_out_1057));
CLKBUFX1 gbuf_q_1057(.A(q_in_1057), .Y(_2146_));
CLKBUFX1 gbuf_d_1058(.A(n_1642), .Y(d_out_1058));
CLKBUFX1 gbuf_q_1058(.A(q_in_1058), .Y(_2148_));
CLKBUFX1 gbuf_d_1059(.A(n_1641), .Y(d_out_1059));
CLKBUFX1 gbuf_q_1059(.A(q_in_1059), .Y(_2149_));
CLKBUFX1 gbuf_d_1060(.A(n_1640), .Y(d_out_1060));
CLKBUFX1 gbuf_q_1060(.A(q_in_1060), .Y(_2151_));
CLKBUFX1 gbuf_d_1061(.A(n_1639), .Y(d_out_1061));
CLKBUFX1 gbuf_q_1061(.A(q_in_1061), .Y(_2154_));
CLKBUFX1 gbuf_d_1062(.A(n_1638), .Y(d_out_1062));
CLKBUFX1 gbuf_q_1062(.A(q_in_1062), .Y(_2155_));
CLKBUFX1 gbuf_d_1063(.A(n_1637), .Y(d_out_1063));
CLKBUFX1 gbuf_q_1063(.A(q_in_1063), .Y(_2156_));
CLKBUFX1 gbuf_d_1064(.A(n_1635), .Y(d_out_1064));
CLKBUFX1 gbuf_q_1064(.A(q_in_1064), .Y(_2159_));
CLKBUFX1 gbuf_d_1065(.A(n_1631), .Y(d_out_1065));
CLKBUFX1 gbuf_q_1065(.A(q_in_1065), .Y(_2164_));
CLKBUFX1 gbuf_d_1066(.A(n_1629), .Y(d_out_1066));
CLKBUFX1 gbuf_q_1066(.A(q_in_1066), .Y(_2165_));
CLKBUFX1 gbuf_d_1067(.A(n_1627), .Y(d_out_1067));
CLKBUFX1 gbuf_q_1067(.A(q_in_1067), .Y(_2167_));
CLKBUFX1 gbuf_d_1068(.A(n_1625), .Y(d_out_1068));
CLKBUFX1 gbuf_q_1068(.A(q_in_1068), .Y(_2169_));
CLKBUFX1 gbuf_d_1069(.A(n_1619), .Y(d_out_1069));
CLKBUFX1 gbuf_q_1069(.A(q_in_1069), .Y(_2178_));
CLKBUFX1 gbuf_d_1070(.A(n_1618), .Y(d_out_1070));
CLKBUFX1 gbuf_q_1070(.A(q_in_1070), .Y(_2179_));
CLKBUFX1 gbuf_d_1071(.A(n_1614), .Y(d_out_1071));
CLKBUFX1 gbuf_q_1071(.A(q_in_1071), .Y(_2186_));
CLKBUFX1 gbuf_d_1072(.A(n_1612), .Y(d_out_1072));
CLKBUFX1 gbuf_q_1072(.A(q_in_1072), .Y(_2188_));
CLKBUFX1 gbuf_d_1073(.A(n_1609), .Y(d_out_1073));
CLKBUFX1 gbuf_q_1073(.A(q_in_1073), .Y(_2191_));
CLKBUFX1 gbuf_d_1074(.A(n_1607), .Y(d_out_1074));
CLKBUFX1 gbuf_q_1074(.A(q_in_1074), .Y(_2193_));
CLKBUFX1 gbuf_d_1075(.A(n_1606), .Y(d_out_1075));
CLKBUFX1 gbuf_q_1075(.A(q_in_1075), .Y(_2195_));
CLKBUFX1 gbuf_d_1076(.A(n_1603), .Y(d_out_1076));
CLKBUFX1 gbuf_q_1076(.A(q_in_1076), .Y(_2200_));
CLKBUFX1 gbuf_d_1077(.A(n_1601), .Y(d_out_1077));
CLKBUFX1 gbuf_q_1077(.A(q_in_1077), .Y(_2203_));
CLKBUFX1 gbuf_d_1078(.A(n_1558), .Y(d_out_1078));
CLKBUFX1 gbuf_q_1078(.A(q_in_1078), .Y(_2284_));
CLKBUFX1 gbuf_d_1079(.A(n_1599), .Y(d_out_1079));
CLKBUFX1 gbuf_q_1079(.A(q_in_1079), .Y(_2208_));
CLKBUFX1 gbuf_d_1080(.A(n_1598), .Y(d_out_1080));
CLKBUFX1 gbuf_q_1080(.A(q_in_1080), .Y(_2211_));
CLKBUFX1 gbuf_d_1081(.A(n_1595), .Y(d_out_1081));
CLKBUFX1 gbuf_q_1081(.A(q_in_1081), .Y(_2213_));
CLKBUFX1 gbuf_d_1082(.A(n_1592), .Y(d_out_1082));
CLKBUFX1 gbuf_q_1082(.A(q_in_1082), .Y(_2217_));
CLKBUFX1 gbuf_d_1083(.A(n_1591), .Y(d_out_1083));
CLKBUFX1 gbuf_q_1083(.A(q_in_1083), .Y(_2223_));
CLKBUFX1 gbuf_d_1084(.A(n_1687), .Y(d_out_1084));
CLKBUFX1 gbuf_q_1084(.A(q_in_1084), .Y(_2222_));
CLKBUFX1 gbuf_d_1085(.A(n_1588), .Y(d_out_1085));
CLKBUFX1 gbuf_q_1085(.A(q_in_1085), .Y(_2226_));
CLKBUFX1 gbuf_d_1086(.A(n_1568), .Y(d_out_1086));
CLKBUFX1 gbuf_q_1086(.A(q_in_1086), .Y(_2227_));
CLKBUFX1 gbuf_d_1087(.A(n_1577), .Y(d_out_1087));
CLKBUFX1 gbuf_q_1087(.A(q_in_1087), .Y(_2228_));
CLKBUFX1 gbuf_d_1088(.A(n_1585), .Y(d_out_1088));
CLKBUFX1 gbuf_q_1088(.A(q_in_1088), .Y(_2230_));
CLKBUFX1 gbuf_d_1089(.A(n_1583), .Y(d_out_1089));
CLKBUFX1 gbuf_q_1089(.A(q_in_1089), .Y(_2233_));
CLKBUFX1 gbuf_d_1090(.A(n_1506), .Y(d_out_1090));
CLKBUFX1 gbuf_q_1090(.A(q_in_1090), .Y(_2234_));
CLKBUFX1 gbuf_d_1091(.A(n_1946), .Y(d_out_1091));
CLKBUFX1 gbuf_q_1091(.A(q_in_1091), .Y(WX3371));
CLKBUFX1 gbuf_d_1092(.A(n_1684), .Y(d_out_1092));
CLKBUFX1 gbuf_q_1092(.A(q_in_1092), .Y(_2238_));
CLKBUFX1 gbuf_d_1093(.A(n_1649), .Y(d_out_1093));
CLKBUFX1 gbuf_q_1093(.A(q_in_1093), .Y(_2245_));
CLKBUFX1 gbuf_d_1094(.A(n_1677), .Y(d_out_1094));
CLKBUFX1 gbuf_q_1094(.A(q_in_1094), .Y(_2249_));
CLKBUFX1 gbuf_d_1095(.A(n_1574), .Y(d_out_1095));
CLKBUFX1 gbuf_q_1095(.A(q_in_1095), .Y(_2254_));
CLKBUFX1 gbuf_d_1096(.A(n_1573), .Y(d_out_1096));
CLKBUFX1 gbuf_q_1096(.A(q_in_1096), .Y(_2256_));
CLKBUFX1 gbuf_d_1097(.A(n_1572), .Y(d_out_1097));
CLKBUFX1 gbuf_q_1097(.A(q_in_1097), .Y(_2259_));
CLKBUFX1 gbuf_d_1098(.A(n_1571), .Y(d_out_1098));
CLKBUFX1 gbuf_q_1098(.A(q_in_1098), .Y(_2260_));
CLKBUFX1 gbuf_d_1099(.A(n_1567), .Y(d_out_1099));
CLKBUFX1 gbuf_q_1099(.A(q_in_1099), .Y(_2266_));
CLKBUFX1 gbuf_d_1100(.A(n_1675), .Y(d_out_1100));
CLKBUFX1 gbuf_q_1100(.A(q_in_1100), .Y(_2269_));
CLKBUFX1 gbuf_d_1101(.A(n_1576), .Y(d_out_1101));
CLKBUFX1 gbuf_q_1101(.A(q_in_1101), .Y(_2274_));
CLKBUFX1 gbuf_d_1102(.A(n_1564), .Y(d_out_1102));
CLKBUFX1 gbuf_q_1102(.A(q_in_1102), .Y(_2275_));
CLKBUFX1 gbuf_d_1103(.A(n_1561), .Y(d_out_1103));
CLKBUFX1 gbuf_q_1103(.A(q_in_1103), .Y(_2279_));
CLKBUFX1 gbuf_d_1104(.A(n_1560), .Y(d_out_1104));
CLKBUFX1 gbuf_q_1104(.A(q_in_1104), .Y(_2282_));
CLKBUFX1 gbuf_d_1105(.A(n_1685), .Y(d_out_1105));
CLKBUFX1 gbuf_q_1105(.A(q_in_1105), .Y(_2288_));
CLKBUFX1 gbuf_d_1106(.A(n_1511), .Y(d_out_1106));
CLKBUFX1 gbuf_q_1106(.A(q_in_1106), .Y(_2286_));
CLKBUFX1 gbuf_d_1107(.A(n_1553), .Y(d_out_1107));
CLKBUFX1 gbuf_q_1107(.A(q_in_1107), .Y(_2299_));
CLKBUFX1 gbuf_d_1108(.A(n_1679), .Y(d_out_1108));
CLKBUFX1 gbuf_q_1108(.A(q_in_1108), .Y(_2311_));
CLKBUFX1 gbuf_d_1109(.A(n_1502), .Y(d_out_1109));
CLKBUFX1 gbuf_q_1109(.A(q_in_1109), .Y(_2314_));
CLKBUFX1 gbuf_d_1110(.A(n_1547), .Y(d_out_1110));
CLKBUFX1 gbuf_q_1110(.A(q_in_1110), .Y(_2316_));
CLKBUFX1 gbuf_d_1111(.A(n_1544), .Y(d_out_1111));
CLKBUFX1 gbuf_q_1111(.A(q_in_1111), .Y(_2321_));
CLKBUFX1 gbuf_d_1112(.A(n_1542), .Y(d_out_1112));
CLKBUFX1 gbuf_q_1112(.A(q_in_1112), .Y(_2322_));
CLKBUFX1 gbuf_d_1113(.A(n_1541), .Y(d_out_1113));
CLKBUFX1 gbuf_q_1113(.A(q_in_1113), .Y(_2323_));
CLKBUFX1 gbuf_d_1114(.A(n_1539), .Y(d_out_1114));
CLKBUFX1 gbuf_q_1114(.A(q_in_1114), .Y(_2325_));
CLKBUFX1 gbuf_d_1115(.A(n_1536), .Y(d_out_1115));
CLKBUFX1 gbuf_q_1115(.A(q_in_1115), .Y(_2329_));
CLKBUFX1 gbuf_d_1116(.A(n_1533), .Y(d_out_1116));
CLKBUFX1 gbuf_q_1116(.A(q_in_1116), .Y(_2338_));
CLKBUFX1 gbuf_d_1117(.A(n_1530), .Y(d_out_1117));
CLKBUFX1 gbuf_q_1117(.A(q_in_1117), .Y(_2340_));
CLKBUFX1 gbuf_d_1118(.A(n_1528), .Y(d_out_1118));
CLKBUFX1 gbuf_q_1118(.A(q_in_1118), .Y(_2342_));
CLKBUFX1 gbuf_d_1119(.A(n_1527), .Y(d_out_1119));
CLKBUFX1 gbuf_q_1119(.A(q_in_1119), .Y(_2343_));
CLKBUFX1 gbuf_d_1120(.A(n_1525), .Y(d_out_1120));
CLKBUFX1 gbuf_q_1120(.A(q_in_1120), .Y(_2345_));
CLKBUFX1 gbuf_d_1121(.A(n_1523), .Y(d_out_1121));
CLKBUFX1 gbuf_q_1121(.A(q_in_1121), .Y(_2356_));
CLKBUFX1 gbuf_d_1122(.A(n_1521), .Y(d_out_1122));
CLKBUFX1 gbuf_q_1122(.A(q_in_1122), .Y(_2358_));
CLKBUFX1 gbuf_d_1123(.A(n_1518), .Y(d_out_1123));
CLKBUFX1 gbuf_q_1123(.A(q_in_1123), .Y(_2360_));
CLKBUFX1 gbuf_d_1124(.A(n_1499), .Y(d_out_1124));
CLKBUFX1 gbuf_q_1124(.A(q_in_1124), .Y(_2265_));
CLKBUFX1 gbuf_d_1125(.A(n_2168), .Y(d_out_1125));
CLKBUFX1 gbuf_q_1125(.A(q_in_1125), .Y(WX11107));
CLKBUFX1 gbuf_d_1126(.A(n_1906), .Y(d_out_1126));
CLKBUFX1 gbuf_q_1126(.A(q_in_1126), .Y(WX11111));
CLKBUFX1 gbuf_d_1127(.A(n_1970), .Y(d_out_1127));
CLKBUFX1 gbuf_q_1127(.A(q_in_1127), .Y(WX11119));
CLKBUFX1 gbuf_d_1128(.A(n_2404), .Y(d_out_1128));
CLKBUFX1 gbuf_q_1128(.A(q_in_1128), .Y(WX11123));
CLKBUFX1 gbuf_d_1129(.A(n_2043), .Y(d_out_1129));
CLKBUFX1 gbuf_q_1129(.A(q_in_1129), .Y(WX11127));
CLKBUFX1 gbuf_d_1130(.A(n_2164), .Y(d_out_1130));
CLKBUFX1 gbuf_q_1130(.A(q_in_1130), .Y(WX11131));
CLKBUFX1 gbuf_d_1131(.A(n_1482), .Y(d_out_1131));
CLKBUFX1 gbuf_q_1131(.A(q_in_1131), .Y(WX11133));
CLKBUFX1 gbuf_d_1132(.A(n_2130), .Y(d_out_1132));
CLKBUFX1 gbuf_q_1132(.A(q_in_1132), .Y(WX11135));
CLKBUFX1 gbuf_d_1133(.A(n_1742), .Y(d_out_1133));
CLKBUFX1 gbuf_q_1133(.A(q_in_1133), .Y(WX11139));
CLKBUFX1 gbuf_d_1134(.A(n_2376), .Y(d_out_1134));
CLKBUFX1 gbuf_q_1134(.A(q_in_1134), .Y(WX11143));
CLKBUFX1 gbuf_d_1135(.A(n_2375), .Y(d_out_1135));
CLKBUFX1 gbuf_q_1135(.A(q_in_1135), .Y(WX7174));
CLKBUFX1 gbuf_d_1136(.A(n_2387), .Y(d_out_1136));
CLKBUFX1 gbuf_q_1136(.A(q_in_1136), .Y(WX7178));
CLKBUFX1 gbuf_d_1137(.A(n_2372), .Y(d_out_1137));
CLKBUFX1 gbuf_q_1137(.A(q_in_1137), .Y(WX11147));
CLKBUFX1 gbuf_d_1138(.A(n_2297), .Y(d_out_1138));
CLKBUFX1 gbuf_q_1138(.A(q_in_1138), .Y(WX7182));
CLKBUFX1 gbuf_d_1139(.A(n_2203), .Y(d_out_1139));
CLKBUFX1 gbuf_q_1139(.A(q_in_1139), .Y(WX11151));
CLKBUFX1 gbuf_d_1140(.A(n_2155), .Y(d_out_1140));
CLKBUFX1 gbuf_q_1140(.A(q_in_1140), .Y(WX7186));
CLKBUFX1 gbuf_d_1141(.A(n_2202), .Y(d_out_1141));
CLKBUFX1 gbuf_q_1141(.A(q_in_1141), .Y(WX7188));
CLKBUFX1 gbuf_d_1142(.A(n_2174), .Y(d_out_1142));
CLKBUFX1 gbuf_q_1142(.A(q_in_1142), .Y(WX7192));
CLKBUFX1 gbuf_d_1143(.A(n_2169), .Y(d_out_1143));
CLKBUFX1 gbuf_q_1143(.A(q_in_1143), .Y(WX11149));
CLKBUFX1 gbuf_d_1144(.A(n_2171), .Y(d_out_1144));
CLKBUFX1 gbuf_q_1144(.A(q_in_1144), .Y(WX7194));
CLKBUFX1 gbuf_d_1145(.A(n_2212), .Y(d_out_1145));
CLKBUFX1 gbuf_q_1145(.A(q_in_1145), .Y(WX7198));
CLKBUFX1 gbuf_d_1146(.A(n_2000), .Y(d_out_1146));
CLKBUFX1 gbuf_q_1146(.A(q_in_1146), .Y(WX7200));
CLKBUFX1 gbuf_d_1147(.A(n_1699), .Y(d_out_1147));
CLKBUFX1 gbuf_q_1147(.A(q_in_1147), .Y(WX7204));
CLKBUFX1 gbuf_d_1148(.A(n_1894), .Y(d_out_1148));
CLKBUFX1 gbuf_q_1148(.A(q_in_1148), .Y(WX11155));
CLKBUFX1 gbuf_d_1149(.A(n_2208), .Y(d_out_1149));
CLKBUFX1 gbuf_q_1149(.A(q_in_1149), .Y(WX7214));
CLKBUFX1 gbuf_d_1150(.A(n_2214), .Y(d_out_1150));
CLKBUFX1 gbuf_q_1150(.A(q_in_1150), .Y(WX7218));
CLKBUFX1 gbuf_d_1151(.A(n_2215), .Y(d_out_1151));
CLKBUFX1 gbuf_q_1151(.A(q_in_1151), .Y(WX7220));
CLKBUFX1 gbuf_d_1152(.A(n_2220), .Y(d_out_1152));
CLKBUFX1 gbuf_q_1152(.A(q_in_1152), .Y(WX7222));
CLKBUFX1 gbuf_d_1153(.A(n_1865), .Y(d_out_1153));
CLKBUFX1 gbuf_q_1153(.A(q_in_1153), .Y(WX7226));
CLKBUFX1 gbuf_d_1154(.A(n_2266), .Y(d_out_1154));
CLKBUFX1 gbuf_q_1154(.A(q_in_1154), .Y(WX7230));
CLKBUFX1 gbuf_d_1155(.A(n_1828), .Y(d_out_1155));
CLKBUFX1 gbuf_q_1155(.A(q_in_1155), .Y(WX7234));
CLKBUFX1 gbuf_d_1156(.A(n_1824), .Y(d_out_1156));
CLKBUFX1 gbuf_q_1156(.A(q_in_1156), .Y(WX11161));
CLKBUFX1 gbuf_d_1157(.A(n_1730), .Y(d_out_1157));
CLKBUFX1 gbuf_q_1157(.A(q_in_1157), .Y(WX7238));
CLKBUFX1 gbuf_d_1158(.A(n_1815), .Y(d_out_1158));
CLKBUFX1 gbuf_q_1158(.A(q_in_1158), .Y(WX7240));
CLKBUFX1 gbuf_d_1159(.A(n_1773), .Y(d_out_1159));
CLKBUFX1 gbuf_q_1159(.A(q_in_1159), .Y(WX11165));
CLKBUFX1 gbuf_d_1160(.A(n_2360), .Y(d_out_1160));
CLKBUFX1 gbuf_q_1160(.A(q_in_1160), .Y(WX7246));
CLKBUFX1 gbuf_d_1161(.A(n_2250), .Y(d_out_1161));
CLKBUFX1 gbuf_q_1161(.A(q_in_1161), .Y(WX7250));
CLKBUFX1 gbuf_d_1162(.A(n_1713), .Y(d_out_1162));
CLKBUFX1 gbuf_q_1162(.A(q_in_1162), .Y(WX7252));
CLKBUFX1 gbuf_d_1163(.A(n_2359), .Y(d_out_1163));
CLKBUFX1 gbuf_q_1163(.A(q_in_1163), .Y(WX11167));
CLKBUFX1 gbuf_d_1164(.A(n_2257), .Y(d_out_1164));
CLKBUFX1 gbuf_q_1164(.A(q_in_1164), .Y(WX7256));
CLKBUFX1 gbuf_d_1165(.A(n_2357), .Y(d_out_1165));
CLKBUFX1 gbuf_q_1165(.A(q_in_1165), .Y(WX7260));
CLKBUFX1 gbuf_d_1166(.A(n_1731), .Y(d_out_1166));
CLKBUFX1 gbuf_q_1166(.A(q_in_1166), .Y(WX7264));
CLKBUFX1 gbuf_d_1167(.A(n_1632), .Y(d_out_1167));
CLKBUFX1 gbuf_q_1167(.A(q_in_1167), .Y(WX7266));
CLKBUFX1 gbuf_d_1168(.A(n_2304), .Y(d_out_1168));
CLKBUFX1 gbuf_q_1168(.A(q_in_1168), .Y(WX11173));
CLKBUFX1 gbuf_d_1169(.A(n_2008), .Y(d_out_1169));
CLKBUFX1 gbuf_q_1169(.A(q_in_1169), .Y(WX7276));
CLKBUFX1 gbuf_d_1170(.A(n_1886), .Y(d_out_1170));
CLKBUFX1 gbuf_q_1170(.A(q_in_1170), .Y(WX7280));
CLKBUFX1 gbuf_d_1171(.A(n_2296), .Y(d_out_1171));
CLKBUFX1 gbuf_q_1171(.A(q_in_1171), .Y(WX7282));
CLKBUFX1 gbuf_d_1172(.A(n_2384), .Y(d_out_1172));
CLKBUFX1 gbuf_q_1172(.A(q_in_1172), .Y(WX7284));
CLKBUFX1 gbuf_d_1173(.A(n_2295), .Y(d_out_1173));
CLKBUFX1 gbuf_q_1173(.A(q_in_1173), .Y(WX7288));
CLKBUFX1 gbuf_d_1174(.A(n_2306), .Y(d_out_1174));
CLKBUFX1 gbuf_q_1174(.A(q_in_1174), .Y(WX7292));
CLKBUFX1 gbuf_d_1175(.A(n_2395), .Y(d_out_1175));
CLKBUFX1 gbuf_q_1175(.A(q_in_1175), .Y(WX11179));
CLKBUFX1 gbuf_d_1176(.A(n_2347), .Y(d_out_1176));
CLKBUFX1 gbuf_q_1176(.A(q_in_1176), .Y(WX7298));
CLKBUFX1 gbuf_d_1177(.A(n_2348), .Y(d_out_1177));
CLKBUFX1 gbuf_q_1177(.A(q_in_1177), .Y(WX11177));
CLKBUFX1 gbuf_d_1178(.A(n_2373), .Y(d_out_1178));
CLKBUFX1 gbuf_q_1178(.A(q_in_1178), .Y(WX7304));
CLKBUFX1 gbuf_d_1179(.A(n_2343), .Y(d_out_1179));
CLKBUFX1 gbuf_q_1179(.A(q_in_1179), .Y(WX7308));
CLKBUFX1 gbuf_d_1180(.A(n_2211), .Y(d_out_1180));
CLKBUFX1 gbuf_q_1180(.A(q_in_1180), .Y(WX7310));
CLKBUFX1 gbuf_d_1181(.A(n_2341), .Y(d_out_1181));
CLKBUFX1 gbuf_q_1181(.A(q_in_1181), .Y(WX7312));
CLKBUFX1 gbuf_d_1182(.A(n_2012), .Y(d_out_1182));
CLKBUFX1 gbuf_q_1182(.A(q_in_1182), .Y(WX7314));
CLKBUFX1 gbuf_d_1183(.A(n_2389), .Y(d_out_1183));
CLKBUFX1 gbuf_q_1183(.A(q_in_1183), .Y(WX11185));
CLKBUFX1 gbuf_d_1184(.A(n_2260), .Y(d_out_1184));
CLKBUFX1 gbuf_q_1184(.A(q_in_1184), .Y(WX7320));
CLKBUFX1 gbuf_d_1185(.A(n_1976), .Y(d_out_1185));
CLKBUFX1 gbuf_q_1185(.A(q_in_1185), .Y(WX7322));
CLKBUFX1 gbuf_d_1186(.A(n_1954), .Y(d_out_1186));
CLKBUFX1 gbuf_q_1186(.A(q_in_1186), .Y(WX7324));
CLKBUFX1 gbuf_d_1187(.A(n_1967), .Y(d_out_1187));
CLKBUFX1 gbuf_q_1187(.A(q_in_1187), .Y(WX7328));
CLKBUFX1 gbuf_d_1188(.A(n_1985), .Y(d_out_1188));
CLKBUFX1 gbuf_q_1188(.A(q_in_1188), .Y(WX11189));
CLKBUFX1 gbuf_d_1189(.A(n_1960), .Y(d_out_1189));
CLKBUFX1 gbuf_q_1189(.A(q_in_1189), .Y(WX7334));
CLKBUFX1 gbuf_d_1190(.A(n_1921), .Y(d_out_1190));
CLKBUFX1 gbuf_q_1190(.A(q_in_1190), .Y(WX7338));
CLKBUFX1 gbuf_d_1191(.A(n_2332), .Y(d_out_1191));
CLKBUFX1 gbuf_q_1191(.A(q_in_1191), .Y(WX7340));
CLKBUFX1 gbuf_d_1192(.A(n_1804), .Y(d_out_1192));
CLKBUFX1 gbuf_q_1192(.A(q_in_1192), .Y(WX11191));
CLKBUFX1 gbuf_d_1193(.A(n_2244), .Y(d_out_1193));
CLKBUFX1 gbuf_q_1193(.A(q_in_1193), .Y(WX7342));
CLKBUFX1 gbuf_d_1194(.A(n_2022), .Y(d_out_1194));
CLKBUFX1 gbuf_q_1194(.A(q_in_1194), .Y(WX7346));
CLKBUFX1 gbuf_d_1195(.A(n_1494), .Y(d_out_1195));
CLKBUFX1 gbuf_q_1195(.A(q_in_1195), .Y(WX11193));
CLKBUFX1 gbuf_d_1196(.A(n_1472), .Y(d_out_1196));
CLKBUFX1 gbuf_q_1196(.A(q_in_1196), .Y(WX7348));
CLKBUFX1 gbuf_d_1197(.A(n_1774), .Y(d_out_1197));
CLKBUFX1 gbuf_q_1197(.A(q_in_1197), .Y(WX7354));
CLKBUFX1 gbuf_d_1198(.A(n_2349), .Y(d_out_1198));
CLKBUFX1 gbuf_q_1198(.A(q_in_1198), .Y(WX7358));
CLKBUFX1 gbuf_d_1199(.A(n_2288), .Y(d_out_1199));
CLKBUFX1 gbuf_q_1199(.A(q_in_1199), .Y(WX4662));
CLKBUFX1 gbuf_d_1200(.A(n_2328), .Y(d_out_1200));
CLKBUFX1 gbuf_q_1200(.A(q_in_1200), .Y(WX11197));
CLKBUFX1 gbuf_d_1201(.A(n_2326), .Y(d_out_1201));
CLKBUFX1 gbuf_q_1201(.A(q_in_1201), .Y(WX11201));
CLKBUFX1 gbuf_d_1202(.A(n_2145), .Y(d_out_1202));
CLKBUFX1 gbuf_q_1202(.A(q_in_1202), .Y(WX11203));
CLKBUFX1 gbuf_d_1203(.A(n_2190), .Y(d_out_1203));
CLKBUFX1 gbuf_q_1203(.A(q_in_1203), .Y(WX11205));
CLKBUFX1 gbuf_d_1204(.A(n_1745), .Y(d_out_1204));
CLKBUFX1 gbuf_q_1204(.A(q_in_1204), .Y(WX11209));
CLKBUFX1 gbuf_d_1205(.A(n_2156), .Y(d_out_1205));
CLKBUFX1 gbuf_q_1205(.A(q_in_1205), .Y(WX11211));
CLKBUFX1 gbuf_d_1206(.A(n_1761), .Y(d_out_1206));
CLKBUFX1 gbuf_q_1206(.A(q_in_1206), .Y(WX7300));
CLKBUFX1 gbuf_d_1207(.A(n_2140), .Y(d_out_1207));
CLKBUFX1 gbuf_q_1207(.A(q_in_1207), .Y(WX11213));
CLKBUFX1 gbuf_d_1208(.A(n_1822), .Y(d_out_1208));
CLKBUFX1 gbuf_q_1208(.A(q_in_1208), .Y(WX11215));
CLKBUFX1 gbuf_d_1209(.A(n_2361), .Y(d_out_1209));
CLKBUFX1 gbuf_q_1209(.A(q_in_1209), .Y(WX11217));
CLKBUFX1 gbuf_d_1210(.A(n_1490), .Y(d_out_1210));
CLKBUFX1 gbuf_q_1210(.A(q_in_1210), .Y(WX11219));
CLKBUFX1 gbuf_d_1211(.A(n_1978), .Y(d_out_1211));
CLKBUFX1 gbuf_q_1211(.A(q_in_1211), .Y(WX4710));
CLKBUFX1 gbuf_d_1212(.A(n_1861), .Y(d_out_1212));
CLKBUFX1 gbuf_q_1212(.A(q_in_1212), .Y(WX11221));
CLKBUFX1 gbuf_d_1213(.A(n_2324), .Y(d_out_1213));
CLKBUFX1 gbuf_q_1213(.A(q_in_1213), .Y(WX11225));
CLKBUFX1 gbuf_d_1214(.A(n_2280), .Y(d_out_1214));
CLKBUFX1 gbuf_q_1214(.A(q_in_1214), .Y(WX11227));
CLKBUFX1 gbuf_d_1215(.A(n_1470), .Y(d_out_1215));
CLKBUFX1 gbuf_q_1215(.A(q_in_1215), .Y(WX11231));
CLKBUFX1 gbuf_d_1216(.A(n_2513), .Y(d_out_1216));
CLKBUFX1 gbuf_q_1216(.A(q_in_1216), .Y(WX11233));
CLKBUFX1 gbuf_d_1217(.A(n_1944), .Y(d_out_1217));
CLKBUFX1 gbuf_q_1217(.A(q_in_1217), .Y(WX4646));
CLKBUFX1 gbuf_d_1218(.A(n_2329), .Y(d_out_1218));
CLKBUFX1 gbuf_q_1218(.A(q_in_1218), .Y(WX11241));
CLKBUFX1 gbuf_d_1219(.A(n_1746), .Y(d_out_1219));
CLKBUFX1 gbuf_q_1219(.A(q_in_1219), .Y(WX11243));
CLKBUFX1 gbuf_d_1220(.A(n_2351), .Y(d_out_1220));
CLKBUFX1 gbuf_q_1220(.A(q_in_1220), .Y(WX4658));
CLKBUFX1 gbuf_d_1221(.A(n_2267), .Y(d_out_1221));
CLKBUFX1 gbuf_q_1221(.A(q_in_1221), .Y(WX3327));
CLKBUFX1 gbuf_d_1222(.A(n_2398), .Y(d_out_1222));
CLKBUFX1 gbuf_q_1222(.A(q_in_1222), .Y(WX3321));
CLKBUFX1 gbuf_d_1223(.A(n_2128), .Y(d_out_1223));
CLKBUFX1 gbuf_q_1223(.A(q_in_1223), .Y(WX4640));
CLKBUFX1 gbuf_d_1224(.A(n_1936), .Y(d_out_1224));
CLKBUFX1 gbuf_q_1224(.A(q_in_1224), .Y(WX4708));
CLKBUFX1 gbuf_d_1225(.A(n_1914), .Y(d_out_1225));
CLKBUFX1 gbuf_q_1225(.A(q_in_1225), .Y(WX7210));
CLKBUFX1 gbuf_d_1226(.A(n_2098), .Y(d_out_1226));
CLKBUFX1 gbuf_q_1226(.A(q_in_1226), .Y(WX3297));
CLKBUFX1 gbuf_d_1227(.A(n_2318), .Y(d_out_1227));
CLKBUFX1 gbuf_q_1227(.A(q_in_1227), .Y(WX3301));
CLKBUFX1 gbuf_d_1228(.A(n_2112), .Y(d_out_1228));
CLKBUFX1 gbuf_q_1228(.A(q_in_1228), .Y(WX3305));
CLKBUFX1 gbuf_d_1229(.A(n_2118), .Y(d_out_1229));
CLKBUFX1 gbuf_q_1229(.A(q_in_1229), .Y(WX3309));
CLKBUFX1 gbuf_d_1230(.A(n_1714), .Y(d_out_1230));
CLKBUFX1 gbuf_q_1230(.A(q_in_1230), .Y(WX3315));
CLKBUFX1 gbuf_d_1231(.A(n_2066), .Y(d_out_1231));
CLKBUFX1 gbuf_q_1231(.A(q_in_1231), .Y(WX3317));
CLKBUFX1 gbuf_d_1232(.A(n_1793), .Y(d_out_1232));
CLKBUFX1 gbuf_q_1232(.A(q_in_1232), .Y(WX3325));
CLKBUFX1 gbuf_d_1233(.A(n_2191), .Y(d_out_1233));
CLKBUFX1 gbuf_q_1233(.A(q_in_1233), .Y(WX3329));
CLKBUFX1 gbuf_d_1234(.A(n_2183), .Y(d_out_1234));
CLKBUFX1 gbuf_q_1234(.A(q_in_1234), .Y(WX3331));
CLKBUFX1 gbuf_d_1235(.A(n_2403), .Y(d_out_1235));
CLKBUFX1 gbuf_q_1235(.A(q_in_1235), .Y(WX3335));
CLKBUFX1 gbuf_d_1236(.A(n_2433), .Y(d_out_1236));
CLKBUFX1 gbuf_q_1236(.A(q_in_1236), .Y(WX3339));
CLKBUFX1 gbuf_d_1237(.A(n_2355), .Y(d_out_1237));
CLKBUFX1 gbuf_q_1237(.A(q_in_1237), .Y(WX3343));
CLKBUFX1 gbuf_d_1238(.A(n_2352), .Y(d_out_1238));
CLKBUFX1 gbuf_q_1238(.A(q_in_1238), .Y(WX3349));
CLKBUFX1 gbuf_d_1239(.A(n_2234), .Y(d_out_1239));
CLKBUFX1 gbuf_q_1239(.A(q_in_1239), .Y(WX3353));
CLKBUFX1 gbuf_d_1240(.A(n_2086), .Y(d_out_1240));
CLKBUFX1 gbuf_q_1240(.A(q_in_1240), .Y(WX7306));
CLKBUFX1 gbuf_d_1241(.A(n_1783), .Y(d_out_1241));
CLKBUFX1 gbuf_q_1241(.A(q_in_1241), .Y(WX3357));
CLKBUFX1 gbuf_d_1242(.A(n_2048), .Y(d_out_1242));
CLKBUFX1 gbuf_q_1242(.A(q_in_1242), .Y(WX3361));
CLKBUFX1 gbuf_d_1243(.A(n_2038), .Y(d_out_1243));
CLKBUFX1 gbuf_q_1243(.A(q_in_1243), .Y(WX3363));
CLKBUFX1 gbuf_d_1244(.A(n_2026), .Y(d_out_1244));
CLKBUFX1 gbuf_q_1244(.A(q_in_1244), .Y(WX8469));
CLKBUFX1 gbuf_d_1245(.A(n_2149), .Y(d_out_1245));
CLKBUFX1 gbuf_q_1245(.A(q_in_1245), .Y(WX8471));
CLKBUFX1 gbuf_d_1246(.A(n_1997), .Y(d_out_1246));
CLKBUFX1 gbuf_q_1246(.A(q_in_1246), .Y(WX8473));
CLKBUFX1 gbuf_d_1247(.A(n_1957), .Y(d_out_1247));
CLKBUFX1 gbuf_q_1247(.A(q_in_1247), .Y(WX3367));
CLKBUFX1 gbuf_d_1248(.A(n_1734), .Y(d_out_1248));
CLKBUFX1 gbuf_q_1248(.A(q_in_1248), .Y(WX8479));
CLKBUFX1 gbuf_d_1249(.A(n_2282), .Y(d_out_1249));
CLKBUFX1 gbuf_q_1249(.A(q_in_1249), .Y(WX11195));
CLKBUFX1 gbuf_d_1250(.A(n_1790), .Y(d_out_1250));
CLKBUFX1 gbuf_q_1250(.A(q_in_1250), .Y(WX8483));
CLKBUFX1 gbuf_d_1251(.A(n_1735), .Y(d_out_1251));
CLKBUFX1 gbuf_q_1251(.A(q_in_1251), .Y(WX3373));
CLKBUFX1 gbuf_d_1252(.A(n_1829), .Y(d_out_1252));
CLKBUFX1 gbuf_q_1252(.A(q_in_1252), .Y(WX8489));
CLKBUFX1 gbuf_d_1253(.A(n_1930), .Y(d_out_1253));
CLKBUFX1 gbuf_q_1253(.A(q_in_1253), .Y(WX8491));
CLKBUFX1 gbuf_d_1254(.A(n_1876), .Y(d_out_1254));
CLKBUFX1 gbuf_q_1254(.A(q_in_1254), .Y(WX3377));
CLKBUFX1 gbuf_d_1255(.A(n_1903), .Y(d_out_1255));
CLKBUFX1 gbuf_q_1255(.A(q_in_1255), .Y(WX8495));
CLKBUFX1 gbuf_d_1256(.A(n_1907), .Y(d_out_1256));
CLKBUFX1 gbuf_q_1256(.A(q_in_1256), .Y(WX8497));
CLKBUFX1 gbuf_d_1257(.A(n_2016), .Y(d_out_1257));
CLKBUFX1 gbuf_q_1257(.A(q_in_1257), .Y(WX8499));
CLKBUFX1 gbuf_d_1258(.A(n_1755), .Y(d_out_1258));
CLKBUFX1 gbuf_q_1258(.A(q_in_1258), .Y(WX3381));
CLKBUFX1 gbuf_d_1259(.A(n_1890), .Y(d_out_1259));
CLKBUFX1 gbuf_q_1259(.A(q_in_1259), .Y(WX8503));
CLKBUFX1 gbuf_d_1260(.A(n_2249), .Y(d_out_1260));
CLKBUFX1 gbuf_q_1260(.A(q_in_1260), .Y(WX8505));
CLKBUFX1 gbuf_d_1261(.A(n_2289), .Y(d_out_1261));
CLKBUFX1 gbuf_q_1261(.A(q_in_1261), .Y(WX3383));
CLKBUFX1 gbuf_d_1262(.A(n_2255), .Y(d_out_1262));
CLKBUFX1 gbuf_q_1262(.A(q_in_1262), .Y(WX8509));
CLKBUFX1 gbuf_d_1263(.A(n_1816), .Y(d_out_1263));
CLKBUFX1 gbuf_q_1263(.A(q_in_1263), .Y(WX3387));
CLKBUFX1 gbuf_d_1264(.A(n_1764), .Y(d_out_1264));
CLKBUFX1 gbuf_q_1264(.A(q_in_1264), .Y(WX8515));
CLKBUFX1 gbuf_d_1265(.A(n_1767), .Y(d_out_1265));
CLKBUFX1 gbuf_q_1265(.A(q_in_1265), .Y(WX3389));
CLKBUFX1 gbuf_d_1266(.A(n_2163), .Y(d_out_1266));
CLKBUFX1 gbuf_q_1266(.A(q_in_1266), .Y(WX8517));
CLKBUFX1 gbuf_d_1267(.A(n_2302), .Y(d_out_1267));
CLKBUFX1 gbuf_q_1267(.A(q_in_1267), .Y(WX3391));
CLKBUFX1 gbuf_d_1268(.A(n_1849), .Y(d_out_1268));
CLKBUFX1 gbuf_q_1268(.A(q_in_1268), .Y(WX3393));
CLKBUFX1 gbuf_d_1269(.A(n_1513), .Y(d_out_1269));
CLKBUFX1 gbuf_q_1269(.A(q_in_1269), .Y(_2135_));
CLKBUFX1 gbuf_d_1270(.A(n_1850), .Y(d_out_1270));
CLKBUFX1 gbuf_q_1270(.A(q_in_1270), .Y(WX8525));
CLKBUFX1 gbuf_d_1271(.A(n_2039), .Y(d_out_1271));
CLKBUFX1 gbuf_q_1271(.A(q_in_1271), .Y(WX3395));
CLKBUFX1 gbuf_d_1272(.A(n_2004), .Y(d_out_1272));
CLKBUFX1 gbuf_q_1272(.A(q_in_1272), .Y(WX3397));
CLKBUFX1 gbuf_d_1273(.A(n_1775), .Y(d_out_1273));
CLKBUFX1 gbuf_q_1273(.A(q_in_1273), .Y(WX8535));
CLKBUFX1 gbuf_d_1274(.A(n_2530), .Y(d_out_1274));
CLKBUFX1 gbuf_q_1274(.A(q_in_1274), .Y(WX3403));
CLKBUFX1 gbuf_d_1275(.A(n_1880), .Y(d_out_1275));
CLKBUFX1 gbuf_q_1275(.A(q_in_1275), .Y(WX8541));
CLKBUFX1 gbuf_d_1276(.A(n_1817), .Y(d_out_1276));
CLKBUFX1 gbuf_q_1276(.A(q_in_1276), .Y(WX3405));
CLKBUFX1 gbuf_d_1277(.A(n_1947), .Y(d_out_1277));
CLKBUFX1 gbuf_q_1277(.A(q_in_1277), .Y(WX8547));
CLKBUFX1 gbuf_d_1278(.A(n_1899), .Y(d_out_1278));
CLKBUFX1 gbuf_q_1278(.A(q_in_1278), .Y(WX3407));
CLKBUFX1 gbuf_d_1279(.A(n_1726), .Y(d_out_1279));
CLKBUFX1 gbuf_q_1279(.A(q_in_1279), .Y(WX8549));
CLKBUFX1 gbuf_d_1280(.A(n_1853), .Y(d_out_1280));
CLKBUFX1 gbuf_q_1280(.A(q_in_1280), .Y(WX3409));
CLKBUFX1 gbuf_d_1281(.A(n_2370), .Y(d_out_1281));
CLKBUFX1 gbuf_q_1281(.A(q_in_1281), .Y(WX8555));
CLKBUFX1 gbuf_d_1282(.A(n_1860), .Y(d_out_1282));
CLKBUFX1 gbuf_q_1282(.A(q_in_1282), .Y(WX8557));
CLKBUFX1 gbuf_d_1283(.A(n_2362), .Y(d_out_1283));
CLKBUFX1 gbuf_q_1283(.A(q_in_1283), .Y(WX3413));
CLKBUFX1 gbuf_d_1284(.A(n_1863), .Y(d_out_1284));
CLKBUFX1 gbuf_q_1284(.A(q_in_1284), .Y(WX8561));
CLKBUFX1 gbuf_d_1285(.A(n_1867), .Y(d_out_1285));
CLKBUFX1 gbuf_q_1285(.A(q_in_1285), .Y(WX8563));
CLKBUFX1 gbuf_d_1286(.A(n_1933), .Y(d_out_1286));
CLKBUFX1 gbuf_q_1286(.A(q_in_1286), .Y(WX3417));
CLKBUFX1 gbuf_d_1287(.A(n_2558), .Y(d_out_1287));
CLKBUFX1 gbuf_q_1287(.A(q_in_1287), .Y(WX8569));
CLKBUFX1 gbuf_d_1288(.A(n_1918), .Y(d_out_1288));
CLKBUFX1 gbuf_q_1288(.A(q_in_1288), .Y(WX8571));
CLKBUFX1 gbuf_d_1289(.A(n_1908), .Y(d_out_1289));
CLKBUFX1 gbuf_q_1289(.A(q_in_1289), .Y(WX8573));
CLKBUFX1 gbuf_d_1290(.A(n_2180), .Y(d_out_1290));
CLKBUFX1 gbuf_q_1290(.A(q_in_1290), .Y(WX3421));
CLKBUFX1 gbuf_d_1291(.A(n_1909), .Y(d_out_1291));
CLKBUFX1 gbuf_q_1291(.A(q_in_1291), .Y(WX8577));
CLKBUFX1 gbuf_d_1292(.A(n_1492), .Y(d_out_1292));
CLKBUFX1 gbuf_q_1292(.A(q_in_1292), .Y(WX3423));
CLKBUFX1 gbuf_d_1293(.A(n_2279), .Y(d_out_1293));
CLKBUFX1 gbuf_q_1293(.A(q_in_1293), .Y(WX8581));
CLKBUFX1 gbuf_d_1294(.A(n_1998), .Y(d_out_1294));
CLKBUFX1 gbuf_q_1294(.A(q_in_1294), .Y(WX4706));
CLKBUFX1 gbuf_d_1295(.A(n_2242), .Y(d_out_1295));
CLKBUFX1 gbuf_q_1295(.A(q_in_1295), .Y(WX3427));
CLKBUFX1 gbuf_d_1296(.A(n_2283), .Y(d_out_1296));
CLKBUFX1 gbuf_q_1296(.A(q_in_1296), .Y(WX3429));
CLKBUFX1 gbuf_d_1297(.A(n_2224), .Y(d_out_1297));
CLKBUFX1 gbuf_q_1297(.A(q_in_1297), .Y(WX8593));
CLKBUFX1 gbuf_d_1298(.A(n_1973), .Y(d_out_1298));
CLKBUFX1 gbuf_q_1298(.A(q_in_1298), .Y(WX3435));
CLKBUFX1 gbuf_d_1299(.A(n_1911), .Y(d_out_1299));
CLKBUFX1 gbuf_q_1299(.A(q_in_1299), .Y(WX3437));
CLKBUFX1 gbuf_d_1300(.A(n_2031), .Y(d_out_1300));
CLKBUFX1 gbuf_q_1300(.A(q_in_1300), .Y(WX8603));
CLKBUFX1 gbuf_d_1301(.A(n_2177), .Y(d_out_1301));
CLKBUFX1 gbuf_q_1301(.A(q_in_1301), .Y(WX11183));
CLKBUFX1 gbuf_d_1302(.A(n_1893), .Y(d_out_1302));
CLKBUFX1 gbuf_q_1302(.A(q_in_1302), .Y(WX3441));
CLKBUFX1 gbuf_d_1303(.A(n_2037), .Y(d_out_1303));
CLKBUFX1 gbuf_q_1303(.A(q_in_1303), .Y(WX8613));
CLKBUFX1 gbuf_d_1304(.A(n_2256), .Y(d_out_1304));
CLKBUFX1 gbuf_q_1304(.A(q_in_1304), .Y(WX7258));
CLKBUFX1 gbuf_d_1305(.A(n_2152), .Y(d_out_1305));
CLKBUFX1 gbuf_q_1305(.A(q_in_1305), .Y(WX8615));
CLKBUFX1 gbuf_d_1306(.A(n_2262), .Y(d_out_1306));
CLKBUFX1 gbuf_q_1306(.A(q_in_1306), .Y(WX3445));
CLKBUFX1 gbuf_d_1307(.A(n_2102), .Y(d_out_1307));
CLKBUFX1 gbuf_q_1307(.A(q_in_1307), .Y(WX3447));
CLKBUFX1 gbuf_d_1308(.A(n_2139), .Y(d_out_1308));
CLKBUFX1 gbuf_q_1308(.A(q_in_1308), .Y(WX8621));
CLKBUFX1 gbuf_d_1309(.A(n_2083), .Y(d_out_1309));
CLKBUFX1 gbuf_q_1309(.A(q_in_1309), .Y(WX3449));
CLKBUFX1 gbuf_d_1310(.A(n_2077), .Y(d_out_1310));
CLKBUFX1 gbuf_q_1310(.A(q_in_1310), .Y(WX8625));
CLKBUFX1 gbuf_d_1311(.A(n_1736), .Y(d_out_1311));
CLKBUFX1 gbuf_q_1311(.A(q_in_1311), .Y(WX8627));
CLKBUFX1 gbuf_d_1312(.A(n_2104), .Y(d_out_1312));
CLKBUFX1 gbuf_q_1312(.A(q_in_1312), .Y(WX8629));
CLKBUFX1 gbuf_d_1313(.A(n_1698), .Y(d_out_1313));
CLKBUFX1 gbuf_q_1313(.A(q_in_1313), .Y(WX3453));
CLKBUFX1 gbuf_d_1314(.A(n_2090), .Y(d_out_1314));
CLKBUFX1 gbuf_q_1314(.A(q_in_1314), .Y(WX8635));
CLKBUFX1 gbuf_d_1315(.A(n_2093), .Y(d_out_1315));
CLKBUFX1 gbuf_q_1315(.A(q_in_1315), .Y(WX8637));
CLKBUFX1 gbuf_d_1316(.A(n_2097), .Y(d_out_1316));
CLKBUFX1 gbuf_q_1316(.A(q_in_1316), .Y(WX3457));
CLKBUFX1 gbuf_d_1317(.A(n_1708), .Y(d_out_1317));
CLKBUFX1 gbuf_q_1317(.A(q_in_1317), .Y(WX8641));
CLKBUFX1 gbuf_d_1318(.A(n_2103), .Y(d_out_1318));
CLKBUFX1 gbuf_q_1318(.A(q_in_1318), .Y(WX8643));
CLKBUFX1 gbuf_d_1319(.A(n_1981), .Y(d_out_1319));
CLKBUFX1 gbuf_q_1319(.A(q_in_1319), .Y(WX3461));
CLKBUFX1 gbuf_d_1320(.A(n_1776), .Y(d_out_1320));
CLKBUFX1 gbuf_q_1320(.A(q_in_1320), .Y(WX3463));
CLKBUFX1 gbuf_d_1321(.A(n_2045), .Y(d_out_1321));
CLKBUFX1 gbuf_q_1321(.A(q_in_1321), .Y(WX3465));
CLKBUFX1 gbuf_d_1322(.A(n_1975), .Y(d_out_1322));
CLKBUFX1 gbuf_q_1322(.A(q_in_1322), .Y(WX8657));
CLKBUFX1 gbuf_d_1323(.A(n_2397), .Y(d_out_1323));
CLKBUFX1 gbuf_q_1323(.A(q_in_1323), .Y(WX3467));
CLKBUFX1 gbuf_d_1324(.A(n_2119), .Y(d_out_1324));
CLKBUFX1 gbuf_q_1324(.A(q_in_1324), .Y(WX3469));
CLKBUFX1 gbuf_d_1325(.A(n_2200), .Y(d_out_1325));
CLKBUFX1 gbuf_q_1325(.A(q_in_1325), .Y(WX3473));
CLKBUFX1 gbuf_d_1326(.A(n_1864), .Y(d_out_1326));
CLKBUFX1 gbuf_q_1326(.A(q_in_1326), .Y(WX3475));
CLKBUFX1 gbuf_d_1327(.A(n_1718), .Y(d_out_1327));
CLKBUFX1 gbuf_q_1327(.A(q_in_1327), .Y(WX3477));
CLKBUFX1 gbuf_d_1328(.A(n_2229), .Y(d_out_1328));
CLKBUFX1 gbuf_q_1328(.A(q_in_1328), .Y(WX3479));
CLKBUFX1 gbuf_d_1329(.A(n_1919), .Y(d_out_1329));
CLKBUFX1 gbuf_q_1329(.A(q_in_1329), .Y(WX3481));
CLKBUFX1 gbuf_d_1330(.A(n_2034), .Y(d_out_1330));
CLKBUFX1 gbuf_q_1330(.A(q_in_1330), .Y(WX3483));
CLKBUFX1 gbuf_d_1331(.A(n_2059), .Y(d_out_1331));
CLKBUFX1 gbuf_q_1331(.A(q_in_1331), .Y(WX9876));
CLKBUFX1 gbuf_d_1332(.A(n_2137), .Y(d_out_1332));
CLKBUFX1 gbuf_q_1332(.A(q_in_1332), .Y(WX9904));
CLKBUFX1 gbuf_d_1333(.A(n_2042), .Y(d_out_1333));
CLKBUFX1 gbuf_q_1333(.A(q_in_1333), .Y(WX9764));
CLKBUFX1 gbuf_d_1334(.A(n_2084), .Y(d_out_1334));
CLKBUFX1 gbuf_q_1334(.A(q_in_1334), .Y(WX9928));
CLKBUFX1 gbuf_d_1335(.A(n_2284), .Y(d_out_1335));
CLKBUFX1 gbuf_q_1335(.A(q_in_1335), .Y(WX9762));
CLKBUFX1 gbuf_d_1336(.A(n_2252), .Y(d_out_1336));
CLKBUFX1 gbuf_q_1336(.A(q_in_1336), .Y(WX9768));
CLKBUFX1 gbuf_d_1337(.A(n_2114), .Y(d_out_1337));
CLKBUFX1 gbuf_q_1337(.A(q_in_1337), .Y(WX9770));
CLKBUFX1 gbuf_d_1338(.A(n_2556), .Y(d_out_1338));
CLKBUFX1 gbuf_q_1338(.A(q_in_1338), .Y(WX9772));
CLKBUFX1 gbuf_d_1339(.A(n_2345), .Y(d_out_1339));
CLKBUFX1 gbuf_q_1339(.A(q_in_1339), .Y(WX9776));
CLKBUFX1 gbuf_d_1340(.A(n_2475), .Y(d_out_1340));
CLKBUFX1 gbuf_q_1340(.A(q_in_1340), .Y(WX9778));
CLKBUFX1 gbuf_d_1341(.A(n_2316), .Y(d_out_1341));
CLKBUFX1 gbuf_q_1341(.A(q_in_1341), .Y(WX9780));
CLKBUFX1 gbuf_d_1342(.A(n_1917), .Y(d_out_1342));
CLKBUFX1 gbuf_q_1342(.A(q_in_1342), .Y(WX9784));
CLKBUFX1 gbuf_d_1343(.A(n_2158), .Y(d_out_1343));
CLKBUFX1 gbuf_q_1343(.A(q_in_1343), .Y(WX9788));
CLKBUFX1 gbuf_d_1344(.A(n_2121), .Y(d_out_1344));
CLKBUFX1 gbuf_q_1344(.A(q_in_1344), .Y(WX9792));
CLKBUFX1 gbuf_d_1345(.A(n_1805), .Y(d_out_1345));
CLKBUFX1 gbuf_q_1345(.A(q_in_1345), .Y(WX9796));
CLKBUFX1 gbuf_d_1346(.A(n_2209), .Y(d_out_1346));
CLKBUFX1 gbuf_q_1346(.A(q_in_1346), .Y(WX9800));
CLKBUFX1 gbuf_d_1347(.A(n_2313), .Y(d_out_1347));
CLKBUFX1 gbuf_q_1347(.A(q_in_1347), .Y(WX9808));
CLKBUFX1 gbuf_d_1348(.A(n_1766), .Y(d_out_1348));
CLKBUFX1 gbuf_q_1348(.A(q_in_1348), .Y(WX9810));
CLKBUFX1 gbuf_d_1349(.A(n_2321), .Y(d_out_1349));
CLKBUFX1 gbuf_q_1349(.A(q_in_1349), .Y(WX9814));
CLKBUFX1 gbuf_d_1350(.A(n_1982), .Y(d_out_1350));
CLKBUFX1 gbuf_q_1350(.A(q_in_1350), .Y(WX9822));
CLKBUFX1 gbuf_d_1351(.A(n_1897), .Y(d_out_1351));
CLKBUFX1 gbuf_q_1351(.A(q_in_1351), .Y(WX9830));
CLKBUFX1 gbuf_d_1352(.A(n_2261), .Y(d_out_1352));
CLKBUFX1 gbuf_q_1352(.A(q_in_1352), .Y(WX9838));
CLKBUFX1 gbuf_d_1353(.A(n_2199), .Y(d_out_1353));
CLKBUFX1 gbuf_q_1353(.A(q_in_1353), .Y(WX9842));
CLKBUFX1 gbuf_d_1354(.A(n_1727), .Y(d_out_1354));
CLKBUFX1 gbuf_q_1354(.A(q_in_1354), .Y(WX9846));
CLKBUFX1 gbuf_d_1355(.A(n_1480), .Y(d_out_1355));
CLKBUFX1 gbuf_q_1355(.A(q_in_1355), .Y(WX9850));
CLKBUFX1 gbuf_d_1356(.A(n_2125), .Y(d_out_1356));
CLKBUFX1 gbuf_q_1356(.A(q_in_1356), .Y(WX9854));
CLKBUFX1 gbuf_d_1357(.A(n_1868), .Y(d_out_1357));
CLKBUFX1 gbuf_q_1357(.A(q_in_1357), .Y(WX9856));
CLKBUFX1 gbuf_d_1358(.A(n_1488), .Y(d_out_1358));
CLKBUFX1 gbuf_q_1358(.A(q_in_1358), .Y(WX9858));
CLKBUFX1 gbuf_d_1359(.A(n_1712), .Y(d_out_1359));
CLKBUFX1 gbuf_q_1359(.A(q_in_1359), .Y(WX9862));
CLKBUFX1 gbuf_d_1360(.A(n_2238), .Y(d_out_1360));
CLKBUFX1 gbuf_q_1360(.A(q_in_1360), .Y(WX9864));
CLKBUFX1 gbuf_d_1361(.A(n_2386), .Y(d_out_1361));
CLKBUFX1 gbuf_q_1361(.A(q_in_1361), .Y(WX9866));
CLKBUFX1 gbuf_d_1362(.A(n_2504), .Y(d_out_1362));
CLKBUFX1 gbuf_q_1362(.A(q_in_1362), .Y(WX9870));
CLKBUFX1 gbuf_d_1363(.A(n_1733), .Y(d_out_1363));
CLKBUFX1 gbuf_q_1363(.A(q_in_1363), .Y(WX9874));
CLKBUFX1 gbuf_d_1364(.A(n_2213), .Y(d_out_1364));
CLKBUFX1 gbuf_q_1364(.A(q_in_1364), .Y(WX9880));
CLKBUFX1 gbuf_d_1365(.A(n_1740), .Y(d_out_1365));
CLKBUFX1 gbuf_q_1365(.A(q_in_1365), .Y(WX9882));
CLKBUFX1 gbuf_d_1366(.A(n_2287), .Y(d_out_1366));
CLKBUFX1 gbuf_q_1366(.A(q_in_1366), .Y(WX9884));
CLKBUFX1 gbuf_d_1367(.A(n_2385), .Y(d_out_1367));
CLKBUFX1 gbuf_q_1367(.A(q_in_1367), .Y(WX9888));
CLKBUFX1 gbuf_d_1368(.A(n_2003), .Y(d_out_1368));
CLKBUFX1 gbuf_q_1368(.A(q_in_1368), .Y(WX9890));
CLKBUFX1 gbuf_d_1369(.A(n_1859), .Y(d_out_1369));
CLKBUFX1 gbuf_q_1369(.A(q_in_1369), .Y(WX9892));
CLKBUFX1 gbuf_d_1370(.A(n_2222), .Y(d_out_1370));
CLKBUFX1 gbuf_q_1370(.A(q_in_1370), .Y(WX9896));
CLKBUFX1 gbuf_d_1371(.A(n_1887), .Y(d_out_1371));
CLKBUFX1 gbuf_q_1371(.A(q_in_1371), .Y(WX9898));
CLKBUFX1 gbuf_d_1372(.A(n_1971), .Y(d_out_1372));
CLKBUFX1 gbuf_q_1372(.A(q_in_1372), .Y(WX9900));
CLKBUFX1 gbuf_d_1373(.A(n_1768), .Y(d_out_1373));
CLKBUFX1 gbuf_q_1373(.A(q_in_1373), .Y(WX9908));
CLKBUFX1 gbuf_d_1374(.A(n_1782), .Y(d_out_1374));
CLKBUFX1 gbuf_q_1374(.A(q_in_1374), .Y(WX9910));
CLKBUFX1 gbuf_d_1375(.A(n_2377), .Y(d_out_1375));
CLKBUFX1 gbuf_q_1375(.A(q_in_1375), .Y(WX9914));
CLKBUFX1 gbuf_d_1376(.A(n_2014), .Y(d_out_1376));
CLKBUFX1 gbuf_q_1376(.A(q_in_1376), .Y(WX9918));
CLKBUFX1 gbuf_d_1377(.A(n_2135), .Y(d_out_1377));
CLKBUFX1 gbuf_q_1377(.A(q_in_1377), .Y(WX2140));
CLKBUFX1 gbuf_d_1378(.A(n_1945), .Y(d_out_1378));
CLKBUFX1 gbuf_q_1378(.A(q_in_1378), .Y(WX9930));
CLKBUFX1 gbuf_d_1379(.A(n_1846), .Y(d_out_1379));
CLKBUFX1 gbuf_q_1379(.A(q_in_1379), .Y(WX9932));
CLKBUFX1 gbuf_d_1380(.A(n_1968), .Y(d_out_1380));
CLKBUFX1 gbuf_q_1380(.A(q_in_1380), .Y(WX9934));
CLKBUFX1 gbuf_d_1381(.A(n_1484), .Y(d_out_1381));
CLKBUFX1 gbuf_q_1381(.A(q_in_1381), .Y(WX9938));
CLKBUFX1 gbuf_d_1382(.A(n_2380), .Y(d_out_1382));
CLKBUFX1 gbuf_q_1382(.A(q_in_1382), .Y(WX9942));
CLKBUFX1 gbuf_d_1383(.A(n_2340), .Y(d_out_1383));
CLKBUFX1 gbuf_q_1383(.A(q_in_1383), .Y(WX9946));
CLKBUFX1 gbuf_d_1384(.A(n_2021), .Y(d_out_1384));
CLKBUFX1 gbuf_q_1384(.A(q_in_1384), .Y(WX9948));
CLKBUFX1 gbuf_d_1385(.A(n_1810), .Y(d_out_1385));
CLKBUFX1 gbuf_q_1385(.A(q_in_1385), .Y(WX8587));
CLKBUFX1 gbuf_d_1386(.A(n_2033), .Y(d_out_1386));
CLKBUFX1 gbuf_q_1386(.A(q_in_1386), .Y(WX8609));
CLKBUFX1 gbuf_d_1387(.A(n_2019), .Y(d_out_1387));
CLKBUFX1 gbuf_q_1387(.A(q_in_1387), .Y(WX4680));
CLKBUFX1 gbuf_d_1388(.A(n_1949), .Y(d_out_1388));
CLKBUFX1 gbuf_q_1388(.A(q_in_1388), .Y(WX4610));
CLKBUFX1 gbuf_d_1389(.A(n_2009), .Y(d_out_1389));
CLKBUFX1 gbuf_q_1389(.A(q_in_1389), .Y(WX8599));
CLKBUFX1 gbuf_d_1390(.A(n_2056), .Y(d_out_1390));
CLKBUFX1 gbuf_q_1390(.A(q_in_1390), .Y(WX8595));
CLKBUFX1 gbuf_d_1391(.A(n_2236), .Y(d_out_1391));
CLKBUFX1 gbuf_q_1391(.A(q_in_1391), .Y(WX8583));
CLKBUFX1 gbuf_d_1392(.A(n_2126), .Y(d_out_1392));
CLKBUFX1 gbuf_q_1392(.A(q_in_1392), .Y(WX4590));
CLKBUFX1 gbuf_d_1393(.A(n_1826), .Y(d_out_1393));
CLKBUFX1 gbuf_q_1393(.A(q_in_1393), .Y(WX4594));
CLKBUFX1 gbuf_d_1394(.A(n_2162), .Y(d_out_1394));
CLKBUFX1 gbuf_q_1394(.A(q_in_1394), .Y(WX4602));
CLKBUFX1 gbuf_d_1395(.A(n_2273), .Y(d_out_1395));
CLKBUFX1 gbuf_q_1395(.A(q_in_1395), .Y(WX4604));
CLKBUFX1 gbuf_d_1396(.A(n_2293), .Y(d_out_1396));
CLKBUFX1 gbuf_q_1396(.A(q_in_1396), .Y(WX4608));
CLKBUFX1 gbuf_d_1397(.A(n_1841), .Y(d_out_1397));
CLKBUFX1 gbuf_q_1397(.A(q_in_1397), .Y(WX4618));
CLKBUFX1 gbuf_d_1398(.A(n_2338), .Y(d_out_1398));
CLKBUFX1 gbuf_q_1398(.A(q_in_1398), .Y(WX4614));
CLKBUFX1 gbuf_d_1399(.A(n_2310), .Y(d_out_1399));
CLKBUFX1 gbuf_q_1399(.A(q_in_1399), .Y(WX4622));
CLKBUFX1 gbuf_d_1400(.A(n_2292), .Y(d_out_1400));
CLKBUFX1 gbuf_q_1400(.A(q_in_1400), .Y(WX4624));
CLKBUFX1 gbuf_d_1401(.A(n_2165), .Y(d_out_1401));
CLKBUFX1 gbuf_q_1401(.A(q_in_1401), .Y(WX4628));
CLKBUFX1 gbuf_d_1402(.A(n_1716), .Y(d_out_1402));
CLKBUFX1 gbuf_q_1402(.A(q_in_1402), .Y(WX4632));
CLKBUFX1 gbuf_d_1403(.A(n_1806), .Y(d_out_1403));
CLKBUFX1 gbuf_q_1403(.A(q_in_1403), .Y(WX4642));
CLKBUFX1 gbuf_d_1404(.A(n_2122), .Y(d_out_1404));
CLKBUFX1 gbuf_q_1404(.A(q_in_1404), .Y(WX4644));
CLKBUFX1 gbuf_d_1405(.A(n_2185), .Y(d_out_1405));
CLKBUFX1 gbuf_q_1405(.A(q_in_1405), .Y(WX4648));
CLKBUFX1 gbuf_d_1406(.A(n_1566), .Y(d_out_1406));
CLKBUFX1 gbuf_q_1406(.A(q_in_1406), .Y(WX4656));
CLKBUFX1 gbuf_d_1407(.A(n_1942), .Y(d_out_1407));
CLKBUFX1 gbuf_q_1407(.A(q_in_1407), .Y(WX4660));
CLKBUFX1 gbuf_d_1408(.A(n_1966), .Y(d_out_1408));
CLKBUFX1 gbuf_q_1408(.A(q_in_1408), .Y(WX4668));
CLKBUFX1 gbuf_d_1409(.A(n_1879), .Y(d_out_1409));
CLKBUFX1 gbuf_q_1409(.A(q_in_1409), .Y(WX4672));
CLKBUFX1 gbuf_d_1410(.A(n_1995), .Y(d_out_1410));
CLKBUFX1 gbuf_q_1410(.A(q_in_1410), .Y(WX4676));
CLKBUFX1 gbuf_d_1411(.A(n_1770), .Y(d_out_1411));
CLKBUFX1 gbuf_q_1411(.A(q_in_1411), .Y(WX4678));
CLKBUFX1 gbuf_d_1412(.A(n_2058), .Y(d_out_1412));
CLKBUFX1 gbuf_q_1412(.A(q_in_1412), .Y(WX4684));
CLKBUFX1 gbuf_d_1413(.A(n_2032), .Y(d_out_1413));
CLKBUFX1 gbuf_q_1413(.A(q_in_1413), .Y(WX4686));
CLKBUFX1 gbuf_d_1414(.A(n_2001), .Y(d_out_1414));
CLKBUFX1 gbuf_q_1414(.A(q_in_1414), .Y(WX4688));
CLKBUFX1 gbuf_d_1415(.A(n_2153), .Y(d_out_1415));
CLKBUFX1 gbuf_q_1415(.A(q_in_1415), .Y(WX4692));
CLKBUFX1 gbuf_d_1416(.A(n_1836), .Y(d_out_1416));
CLKBUFX1 gbuf_q_1416(.A(q_in_1416), .Y(WX4694));
CLKBUFX1 gbuf_d_1417(.A(n_1799), .Y(d_out_1417));
CLKBUFX1 gbuf_q_1417(.A(q_in_1417), .Y(WX4696));
CLKBUFX1 gbuf_d_1418(.A(n_2024), .Y(d_out_1418));
CLKBUFX1 gbuf_q_1418(.A(q_in_1418), .Y(WX8607));
CLKBUFX1 gbuf_d_1419(.A(n_1943), .Y(d_out_1419));
CLKBUFX1 gbuf_q_1419(.A(q_in_1419), .Y(WX4704));
CLKBUFX1 gbuf_d_1420(.A(n_2025), .Y(d_out_1420));
CLKBUFX1 gbuf_q_1420(.A(q_in_1420), .Y(WX4714));
CLKBUFX1 gbuf_d_1421(.A(n_2005), .Y(d_out_1421));
CLKBUFX1 gbuf_q_1421(.A(q_in_1421), .Y(WX4720));
CLKBUFX1 gbuf_d_1422(.A(n_1778), .Y(d_out_1422));
CLKBUFX1 gbuf_q_1422(.A(q_in_1422), .Y(WX4722));
CLKBUFX1 gbuf_d_1423(.A(n_2063), .Y(d_out_1423));
CLKBUFX1 gbuf_q_1423(.A(q_in_1423), .Y(WX4724));
CLKBUFX1 gbuf_d_1424(.A(n_2065), .Y(d_out_1424));
CLKBUFX1 gbuf_q_1424(.A(q_in_1424), .Y(WX4728));
CLKBUFX1 gbuf_d_1425(.A(n_2072), .Y(d_out_1425));
CLKBUFX1 gbuf_q_1425(.A(q_in_1425), .Y(WX4730));
CLKBUFX1 gbuf_d_1426(.A(n_1771), .Y(d_out_1426));
CLKBUFX1 gbuf_q_1426(.A(q_in_1426), .Y(WX4732));
CLKBUFX1 gbuf_d_1427(.A(n_1769), .Y(d_out_1427));
CLKBUFX1 gbuf_q_1427(.A(q_in_1427), .Y(WX4736));
CLKBUFX1 gbuf_d_1428(.A(n_2069), .Y(d_out_1428));
CLKBUFX1 gbuf_q_1428(.A(q_in_1428), .Y(WX4738));
CLKBUFX1 gbuf_d_1429(.A(n_2217), .Y(d_out_1429));
CLKBUFX1 gbuf_q_1429(.A(q_in_1429), .Y(WX4740));
CLKBUFX1 gbuf_d_1430(.A(n_2079), .Y(d_out_1430));
CLKBUFX1 gbuf_q_1430(.A(q_in_1430), .Y(WX4744));
CLKBUFX1 gbuf_d_1431(.A(n_1929), .Y(d_out_1431));
CLKBUFX1 gbuf_q_1431(.A(q_in_1431), .Y(WX4748));
CLKBUFX1 gbuf_d_1432(.A(n_2115), .Y(d_out_1432));
CLKBUFX1 gbuf_q_1432(.A(q_in_1432), .Y(WX4752));
CLKBUFX1 gbuf_d_1433(.A(n_1759), .Y(d_out_1433));
CLKBUFX1 gbuf_q_1433(.A(q_in_1433), .Y(WX4756));
CLKBUFX1 gbuf_d_1434(.A(n_1869), .Y(d_out_1434));
CLKBUFX1 gbuf_q_1434(.A(q_in_1434), .Y(WX2188));
CLKBUFX1 gbuf_d_1435(.A(n_2078), .Y(d_out_1435));
CLKBUFX1 gbuf_q_1435(.A(q_in_1435), .Y(WX4760));
CLKBUFX1 gbuf_d_1436(.A(n_1760), .Y(d_out_1436));
CLKBUFX1 gbuf_q_1436(.A(q_in_1436), .Y(WX4764));
CLKBUFX1 gbuf_d_1437(.A(n_2108), .Y(d_out_1437));
CLKBUFX1 gbuf_q_1437(.A(q_in_1437), .Y(WX4768));
CLKBUFX1 gbuf_d_1438(.A(n_1821), .Y(d_out_1438));
CLKBUFX1 gbuf_q_1438(.A(q_in_1438), .Y(WX4770));
CLKBUFX1 gbuf_d_1439(.A(n_1751), .Y(d_out_1439));
CLKBUFX1 gbuf_q_1439(.A(q_in_1439), .Y(WX4772));
CLKBUFX1 gbuf_d_1440(.A(n_2105), .Y(d_out_1440));
CLKBUFX1 gbuf_q_1440(.A(q_in_1440), .Y(WX4776));
CLKBUFX1 gbuf_d_1441(.A(n_1844), .Y(d_out_1441));
CLKBUFX1 gbuf_q_1441(.A(q_in_1441), .Y(WX4778));
CLKBUFX1 gbuf_d_1442(.A(n_1941), .Y(d_out_1442));
CLKBUFX1 gbuf_q_1442(.A(q_in_1442), .Y(WX7362));
CLKBUFX1 gbuf_d_1443(.A(n_2204), .Y(d_out_1443));
CLKBUFX1 gbuf_q_1443(.A(q_in_1443), .Y(WX4698));
CLKBUFX1 gbuf_d_1444(.A(n_1927), .Y(d_out_1444));
CLKBUFX1 gbuf_q_1444(.A(q_in_1444), .Y(WX9950));
CLKBUFX1 gbuf_d_1445(.A(n_2006), .Y(d_out_1445));
CLKBUFX1 gbuf_q_1445(.A(q_in_1445), .Y(WX4650));
CLKBUFX1 gbuf_d_1446(.A(n_2028), .Y(d_out_1446));
CLKBUFX1 gbuf_q_1446(.A(q_in_1446), .Y(WX4664));
CLKBUFX1 gbuf_d_1447(.A(n_2230), .Y(d_out_1447));
CLKBUFX1 gbuf_q_1447(.A(q_in_1447), .Y(WX9818));
CLKBUFX1 gbuf_d_1448(.A(n_2382), .Y(d_out_1448));
CLKBUFX1 gbuf_q_1448(.A(q_in_1448), .Y(WX11137));
CLKBUFX1 gbuf_d_1449(.A(n_1802), .Y(d_out_1449));
CLKBUFX1 gbuf_q_1449(.A(q_in_1449), .Y(WX8533));
CLKBUFX1 gbuf_d_1450(.A(n_1477), .Y(d_out_1450));
CLKBUFX1 gbuf_q_1450(.A(q_in_1450), .Y(WX5881));
CLKBUFX1 gbuf_d_1451(.A(n_2291), .Y(d_out_1451));
CLKBUFX1 gbuf_q_1451(.A(q_in_1451), .Y(WX5883));
CLKBUFX1 gbuf_d_1452(.A(n_2515), .Y(d_out_1452));
CLKBUFX1 gbuf_q_1452(.A(q_in_1452), .Y(WX5887));
CLKBUFX1 gbuf_d_1453(.A(n_1777), .Y(d_out_1453));
CLKBUFX1 gbuf_q_1453(.A(q_in_1453), .Y(WX5889));
CLKBUFX1 gbuf_d_1454(.A(n_1786), .Y(d_out_1454));
CLKBUFX1 gbuf_q_1454(.A(q_in_1454), .Y(WX5891));
CLKBUFX1 gbuf_d_1455(.A(n_2235), .Y(d_out_1455));
CLKBUFX1 gbuf_q_1455(.A(q_in_1455), .Y(WX5895));
CLKBUFX1 gbuf_d_1456(.A(n_1795), .Y(d_out_1456));
CLKBUFX1 gbuf_q_1456(.A(q_in_1456), .Y(WX5897));
CLKBUFX1 gbuf_d_1457(.A(n_1827), .Y(d_out_1457));
CLKBUFX1 gbuf_q_1457(.A(q_in_1457), .Y(WX8529));
CLKBUFX1 gbuf_d_1458(.A(n_1476), .Y(d_out_1458));
CLKBUFX1 gbuf_q_1458(.A(q_in_1458), .Y(WX5901));
CLKBUFX1 gbuf_d_1459(.A(n_1798), .Y(d_out_1459));
CLKBUFX1 gbuf_q_1459(.A(q_in_1459), .Y(WX5905));
CLKBUFX1 gbuf_d_1460(.A(n_1728), .Y(d_out_1460));
CLKBUFX1 gbuf_q_1460(.A(q_in_1460), .Y(WX5909));
CLKBUFX1 gbuf_d_1461(.A(n_1803), .Y(d_out_1461));
CLKBUFX1 gbuf_q_1461(.A(q_in_1461), .Y(WX5911));
CLKBUFX1 gbuf_d_1462(.A(n_2047), .Y(d_out_1462));
CLKBUFX1 gbuf_q_1462(.A(q_in_1462), .Y(WX5913));
CLKBUFX1 gbuf_d_1463(.A(n_1882), .Y(d_out_1463));
CLKBUFX1 gbuf_q_1463(.A(q_in_1463), .Y(WX5917));
CLKBUFX1 gbuf_d_1464(.A(n_2017), .Y(d_out_1464));
CLKBUFX1 gbuf_q_1464(.A(q_in_1464), .Y(WX5919));
CLKBUFX1 gbuf_d_1465(.A(n_1789), .Y(d_out_1465));
CLKBUFX1 gbuf_q_1465(.A(q_in_1465), .Y(WX5921));
CLKBUFX1 gbuf_d_1466(.A(n_2150), .Y(d_out_1466));
CLKBUFX1 gbuf_q_1466(.A(q_in_1466), .Y(WX5925));
CLKBUFX1 gbuf_d_1467(.A(n_1809), .Y(d_out_1467));
CLKBUFX1 gbuf_q_1467(.A(q_in_1467), .Y(WX5929));
CLKBUFX1 gbuf_d_1468(.A(n_1747), .Y(d_out_1468));
CLKBUFX1 gbuf_q_1468(.A(q_in_1468), .Y(WX5933));
CLKBUFX1 gbuf_d_1469(.A(n_2315), .Y(d_out_1469));
CLKBUFX1 gbuf_q_1469(.A(q_in_1469), .Y(WX5935));
CLKBUFX1 gbuf_d_1470(.A(n_1702), .Y(d_out_1470));
CLKBUFX1 gbuf_q_1470(.A(q_in_1470), .Y(WX5937));
CLKBUFX1 gbuf_d_1471(.A(n_2330), .Y(d_out_1471));
CLKBUFX1 gbuf_q_1471(.A(q_in_1471), .Y(WX5915));
CLKBUFX1 gbuf_d_1472(.A(n_1963), .Y(d_out_1472));
CLKBUFX1 gbuf_q_1472(.A(q_in_1472), .Y(WX5941));
CLKBUFX1 gbuf_d_1473(.A(n_2271), .Y(d_out_1473));
CLKBUFX1 gbuf_q_1473(.A(q_in_1473), .Y(WX5943));
CLKBUFX1 gbuf_d_1474(.A(n_1937), .Y(d_out_1474));
CLKBUFX1 gbuf_q_1474(.A(q_in_1474), .Y(WX5945));
CLKBUFX1 gbuf_d_1475(.A(n_1808), .Y(d_out_1475));
CLKBUFX1 gbuf_q_1475(.A(q_in_1475), .Y(WX5949));
CLKBUFX1 gbuf_d_1476(.A(n_1834), .Y(d_out_1476));
CLKBUFX1 gbuf_q_1476(.A(q_in_1476), .Y(WX5951));
CLKBUFX1 gbuf_d_1477(.A(n_1881), .Y(d_out_1477));
CLKBUFX1 gbuf_q_1477(.A(q_in_1477), .Y(WX5953));
CLKBUFX1 gbuf_d_1478(.A(n_1781), .Y(d_out_1478));
CLKBUFX1 gbuf_q_1478(.A(q_in_1478), .Y(WX5957));
CLKBUFX1 gbuf_d_1479(.A(n_1835), .Y(d_out_1479));
CLKBUFX1 gbuf_q_1479(.A(q_in_1479), .Y(WX5959));
CLKBUFX1 gbuf_d_1480(.A(n_1831), .Y(d_out_1480));
CLKBUFX1 gbuf_q_1480(.A(q_in_1480), .Y(WX5961));
CLKBUFX1 gbuf_d_1481(.A(n_2420), .Y(d_out_1481));
CLKBUFX1 gbuf_q_1481(.A(q_in_1481), .Y(WX5965));
CLKBUFX1 gbuf_d_1482(.A(n_1953), .Y(d_out_1482));
CLKBUFX1 gbuf_q_1482(.A(q_in_1482), .Y(WX5967));
CLKBUFX1 gbuf_d_1483(.A(n_1854), .Y(d_out_1483));
CLKBUFX1 gbuf_q_1483(.A(q_in_1483), .Y(WX5969));
CLKBUFX1 gbuf_d_1484(.A(n_1763), .Y(d_out_1484));
CLKBUFX1 gbuf_q_1484(.A(q_in_1484), .Y(WX5973));
CLKBUFX1 gbuf_d_1485(.A(n_1858), .Y(d_out_1485));
CLKBUFX1 gbuf_q_1485(.A(q_in_1485), .Y(WX5975));
CLKBUFX1 gbuf_d_1486(.A(n_1855), .Y(d_out_1486));
CLKBUFX1 gbuf_q_1486(.A(q_in_1486), .Y(WX5977));
CLKBUFX1 gbuf_d_1487(.A(n_1862), .Y(d_out_1487));
CLKBUFX1 gbuf_q_1487(.A(q_in_1487), .Y(WX5981));
CLKBUFX1 gbuf_d_1488(.A(n_2365), .Y(d_out_1488));
CLKBUFX1 gbuf_q_1488(.A(q_in_1488), .Y(WX5983));
CLKBUFX1 gbuf_d_1489(.A(n_1701), .Y(d_out_1489));
CLKBUFX1 gbuf_q_1489(.A(q_in_1489), .Y(WX5985));
CLKBUFX1 gbuf_d_1490(.A(n_2358), .Y(d_out_1490));
CLKBUFX1 gbuf_q_1490(.A(q_in_1490), .Y(WX5989));
CLKBUFX1 gbuf_d_1491(.A(n_2018), .Y(d_out_1491));
CLKBUFX1 gbuf_q_1491(.A(q_in_1491), .Y(WX8521));
CLKBUFX1 gbuf_d_1492(.A(n_2335), .Y(d_out_1492));
CLKBUFX1 gbuf_q_1492(.A(q_in_1492), .Y(WX5991));
CLKBUFX1 gbuf_d_1493(.A(n_1871), .Y(d_out_1493));
CLKBUFX1 gbuf_q_1493(.A(q_in_1493), .Y(WX5995));
CLKBUFX1 gbuf_d_1494(.A(n_1874), .Y(d_out_1494));
CLKBUFX1 gbuf_q_1494(.A(q_in_1494), .Y(WX5999));
CLKBUFX1 gbuf_d_1495(.A(n_2317), .Y(d_out_1495));
CLKBUFX1 gbuf_q_1495(.A(q_in_1495), .Y(WX6003));
CLKBUFX1 gbuf_d_1496(.A(n_2534), .Y(d_out_1496));
CLKBUFX1 gbuf_q_1496(.A(q_in_1496), .Y(WX6005));
CLKBUFX1 gbuf_d_1497(.A(n_1892), .Y(d_out_1497));
CLKBUFX1 gbuf_q_1497(.A(q_in_1497), .Y(WX6007));
CLKBUFX1 gbuf_d_1498(.A(n_2189), .Y(d_out_1498));
CLKBUFX1 gbuf_q_1498(.A(q_in_1498), .Y(WX6011));
CLKBUFX1 gbuf_d_1499(.A(n_2192), .Y(d_out_1499));
CLKBUFX1 gbuf_q_1499(.A(q_in_1499), .Y(WX6013));
CLKBUFX1 gbuf_d_1500(.A(n_2050), .Y(d_out_1500));
CLKBUFX1 gbuf_q_1500(.A(q_in_1500), .Y(WX6015));
CLKBUFX1 gbuf_d_1501(.A(n_1811), .Y(d_out_1501));
CLKBUFX1 gbuf_q_1501(.A(q_in_1501), .Y(WX6019));
CLKBUFX1 gbuf_d_1502(.A(n_2161), .Y(d_out_1502));
CLKBUFX1 gbuf_q_1502(.A(q_in_1502), .Y(WX6023));
CLKBUFX1 gbuf_d_1503(.A(n_1910), .Y(d_out_1503));
CLKBUFX1 gbuf_q_1503(.A(q_in_1503), .Y(WX6027));
CLKBUFX1 gbuf_d_1504(.A(n_2157), .Y(d_out_1504));
CLKBUFX1 gbuf_q_1504(.A(q_in_1504), .Y(WX6029));
CLKBUFX1 gbuf_d_1505(.A(n_1915), .Y(d_out_1505));
CLKBUFX1 gbuf_q_1505(.A(q_in_1505), .Y(WX6031));
CLKBUFX1 gbuf_d_1506(.A(n_1916), .Y(d_out_1506));
CLKBUFX1 gbuf_q_1506(.A(q_in_1506), .Y(WX6035));
CLKBUFX1 gbuf_d_1507(.A(n_1923), .Y(d_out_1507));
CLKBUFX1 gbuf_q_1507(.A(q_in_1507), .Y(WX6039));
CLKBUFX1 gbuf_d_1508(.A(n_2286), .Y(d_out_1508));
CLKBUFX1 gbuf_q_1508(.A(q_in_1508), .Y(WX6043));
CLKBUFX1 gbuf_d_1509(.A(n_2007), .Y(d_out_1509));
CLKBUFX1 gbuf_q_1509(.A(q_in_1509), .Y(WX6045));
CLKBUFX1 gbuf_d_1510(.A(n_1932), .Y(d_out_1510));
CLKBUFX1 gbuf_q_1510(.A(q_in_1510), .Y(WX6047));
CLKBUFX1 gbuf_d_1511(.A(n_2269), .Y(d_out_1511));
CLKBUFX1 gbuf_q_1511(.A(q_in_1511), .Y(WX6055));
CLKBUFX1 gbuf_d_1512(.A(n_1794), .Y(d_out_1512));
CLKBUFX1 gbuf_q_1512(.A(q_in_1512), .Y(WX6059));
CLKBUFX1 gbuf_d_1513(.A(n_2254), .Y(d_out_1513));
CLKBUFX1 gbuf_q_1513(.A(q_in_1513), .Y(WX6063));
CLKBUFX1 gbuf_d_1514(.A(n_1979), .Y(d_out_1514));
CLKBUFX1 gbuf_q_1514(.A(q_in_1514), .Y(WX6067));
CLKBUFX1 gbuf_d_1515(.A(n_1812), .Y(d_out_1515));
CLKBUFX1 gbuf_q_1515(.A(q_in_1515), .Y(WX6069));
CLKBUFX1 gbuf_d_1516(.A(n_1752), .Y(d_out_1516));
CLKBUFX1 gbuf_q_1516(.A(q_in_1516), .Y(WX6071));
CLKBUFX1 gbuf_d_1517(.A(n_1934), .Y(d_out_1517));
CLKBUFX1 gbuf_q_1517(.A(q_in_1517), .Y(WX4718));
CLKBUFX1 gbuf_d_1518(.A(n_1758), .Y(d_out_1518));
CLKBUFX1 gbuf_q_1518(.A(q_in_1518), .Y(WX8507));
CLKBUFX1 gbuf_d_1519(.A(n_1852), .Y(d_out_1519));
CLKBUFX1 gbuf_q_1519(.A(q_in_1519), .Y(WX9812));
CLKBUFX1 gbuf_d_1520(.A(n_2476), .Y(d_out_1520));
CLKBUFX1 gbuf_q_1520(.A(q_in_1520), .Y(WX2068));
CLKBUFX1 gbuf_d_1521(.A(n_2087), .Y(d_out_1521));
CLKBUFX1 gbuf_q_1521(.A(q_in_1521), .Y(WX2072));
CLKBUFX1 gbuf_d_1522(.A(n_2081), .Y(d_out_1522));
CLKBUFX1 gbuf_q_1522(.A(q_in_1522), .Y(WX2076));
CLKBUFX1 gbuf_d_1523(.A(n_2044), .Y(d_out_1523));
CLKBUFX1 gbuf_q_1523(.A(q_in_1523), .Y(WX2080));
CLKBUFX1 gbuf_d_1524(.A(n_1753), .Y(d_out_1524));
CLKBUFX1 gbuf_q_1524(.A(q_in_1524), .Y(WX2084));
CLKBUFX1 gbuf_d_1525(.A(n_1832), .Y(d_out_1525));
CLKBUFX1 gbuf_q_1525(.A(q_in_1525), .Y(WX2088));
CLKBUFX1 gbuf_d_1526(.A(n_1926), .Y(d_out_1526));
CLKBUFX1 gbuf_q_1526(.A(q_in_1526), .Y(WX4616));
CLKBUFX1 gbuf_d_1527(.A(n_1739), .Y(d_out_1527));
CLKBUFX1 gbuf_q_1527(.A(q_in_1527), .Y(WX2090));
CLKBUFX1 gbuf_d_1528(.A(n_1757), .Y(d_out_1528));
CLKBUFX1 gbuf_q_1528(.A(q_in_1528), .Y(WX2096));
CLKBUFX1 gbuf_d_1529(.A(n_1743), .Y(d_out_1529));
CLKBUFX1 gbuf_q_1529(.A(q_in_1529), .Y(WX2094));
CLKBUFX1 gbuf_d_1530(.A(n_1939), .Y(d_out_1530));
CLKBUFX1 gbuf_q_1530(.A(q_in_1530), .Y(WX2102));
CLKBUFX1 gbuf_d_1531(.A(n_1857), .Y(d_out_1531));
CLKBUFX1 gbuf_q_1531(.A(q_in_1531), .Y(WX2104));
CLKBUFX1 gbuf_d_1532(.A(n_2301), .Y(d_out_1532));
CLKBUFX1 gbuf_q_1532(.A(q_in_1532), .Y(WX2106));
CLKBUFX1 gbuf_d_1533(.A(n_1749), .Y(d_out_1533));
CLKBUFX1 gbuf_q_1533(.A(q_in_1533), .Y(WX2110));
CLKBUFX1 gbuf_d_1534(.A(n_2029), .Y(d_out_1534));
CLKBUFX1 gbuf_q_1534(.A(q_in_1534), .Y(WX2112));
CLKBUFX1 gbuf_d_1535(.A(n_1779), .Y(d_out_1535));
CLKBUFX1 gbuf_q_1535(.A(q_in_1535), .Y(WX2114));
CLKBUFX1 gbuf_d_1536(.A(n_1497), .Y(d_out_1536));
CLKBUFX1 gbuf_q_1536(.A(q_in_1536), .Y(_2276_));
CLKBUFX1 gbuf_d_1537(.A(n_1748), .Y(d_out_1537));
CLKBUFX1 gbuf_q_1537(.A(q_in_1537), .Y(WX2118));
CLKBUFX1 gbuf_d_1538(.A(n_2268), .Y(d_out_1538));
CLKBUFX1 gbuf_q_1538(.A(q_in_1538), .Y(WX2120));
CLKBUFX1 gbuf_d_1539(.A(n_1851), .Y(d_out_1539));
CLKBUFX1 gbuf_q_1539(.A(q_in_1539), .Y(WX2122));
CLKBUFX1 gbuf_d_1540(.A(n_1983), .Y(d_out_1540));
CLKBUFX1 gbuf_q_1540(.A(q_in_1540), .Y(WX2126));
CLKBUFX1 gbuf_d_1541(.A(n_2336), .Y(d_out_1541));
CLKBUFX1 gbuf_q_1541(.A(q_in_1541), .Y(WX2128));
CLKBUFX1 gbuf_d_1542(.A(n_2368), .Y(d_out_1542));
CLKBUFX1 gbuf_q_1542(.A(q_in_1542), .Y(WX2132));
CLKBUFX1 gbuf_d_1543(.A(n_1479), .Y(d_out_1543));
CLKBUFX1 gbuf_q_1543(.A(q_in_1543), .Y(WX2136));
CLKBUFX1 gbuf_d_1544(.A(n_1940), .Y(d_out_1544));
CLKBUFX1 gbuf_q_1544(.A(q_in_1544), .Y(WX2142));
CLKBUFX1 gbuf_d_1545(.A(n_1744), .Y(d_out_1545));
CLKBUFX1 gbuf_q_1545(.A(q_in_1545), .Y(WX2144));
CLKBUFX1 gbuf_d_1546(.A(n_2259), .Y(d_out_1546));
CLKBUFX1 gbuf_q_1546(.A(q_in_1546), .Y(WX2148));
CLKBUFX1 gbuf_d_1547(.A(n_2239), .Y(d_out_1547));
CLKBUFX1 gbuf_q_1547(.A(q_in_1547), .Y(WX2152));
CLKBUFX1 gbuf_d_1548(.A(n_1843), .Y(d_out_1548));
CLKBUFX1 gbuf_q_1548(.A(q_in_1548), .Y(WX2154));
CLKBUFX1 gbuf_d_1549(.A(n_2030), .Y(d_out_1549));
CLKBUFX1 gbuf_q_1549(.A(q_in_1549), .Y(WX2158));
CLKBUFX1 gbuf_d_1550(.A(n_2040), .Y(d_out_1550));
CLKBUFX1 gbuf_q_1550(.A(q_in_1550), .Y(WX2160));
CLKBUFX1 gbuf_d_1551(.A(n_2049), .Y(d_out_1551));
CLKBUFX1 gbuf_q_1551(.A(q_in_1551), .Y(WX2162));
CLKBUFX1 gbuf_d_1552(.A(n_2052), .Y(d_out_1552));
CLKBUFX1 gbuf_q_1552(.A(q_in_1552), .Y(WX2164));
CLKBUFX1 gbuf_d_1553(.A(n_2100), .Y(d_out_1553));
CLKBUFX1 gbuf_q_1553(.A(q_in_1553), .Y(WX2168));
CLKBUFX1 gbuf_d_1554(.A(n_2075), .Y(d_out_1554));
CLKBUFX1 gbuf_q_1554(.A(q_in_1554), .Y(WX2170));
CLKBUFX1 gbuf_d_1555(.A(n_2089), .Y(d_out_1555));
CLKBUFX1 gbuf_q_1555(.A(q_in_1555), .Y(WX2172));
CLKBUFX1 gbuf_d_1556(.A(n_2232), .Y(d_out_1556));
CLKBUFX1 gbuf_q_1556(.A(q_in_1556), .Y(WX2176));
CLKBUFX1 gbuf_d_1557(.A(n_2186), .Y(d_out_1557));
CLKBUFX1 gbuf_q_1557(.A(q_in_1557), .Y(WX2178));
CLKBUFX1 gbuf_d_1558(.A(n_1823), .Y(d_out_1558));
CLKBUFX1 gbuf_q_1558(.A(q_in_1558), .Y(WX2180));
CLKBUFX1 gbuf_d_1559(.A(n_1486), .Y(d_out_1559));
CLKBUFX1 gbuf_q_1559(.A(q_in_1559), .Y(WX9912));
CLKBUFX1 gbuf_d_1560(.A(n_2225), .Y(d_out_1560));
CLKBUFX1 gbuf_q_1560(.A(q_in_1560), .Y(WX2186));
CLKBUFX1 gbuf_d_1561(.A(n_2245), .Y(d_out_1561));
CLKBUFX1 gbuf_q_1561(.A(q_in_1561), .Y(WX2190));
CLKBUFX1 gbuf_d_1562(.A(n_1722), .Y(d_out_1562));
CLKBUFX1 gbuf_q_1562(.A(q_in_1562), .Y(WX11095));
CLKBUFX1 gbuf_d_1563(.A(n_1845), .Y(d_out_1563));
CLKBUFX1 gbuf_q_1563(.A(q_in_1563), .Y(WX8481));
CLKBUFX1 gbuf_d_1564(.A(n_1866), .Y(d_out_1564));
CLKBUFX1 gbuf_q_1564(.A(q_in_1564), .Y(WX11055));
CLKBUFX1 gbuf_d_1565(.A(n_1707), .Y(d_out_1565));
CLKBUFX1 gbuf_q_1565(.A(q_in_1565), .Y(WX11057));
CLKBUFX1 gbuf_d_1566(.A(n_2023), .Y(d_out_1566));
CLKBUFX1 gbuf_q_1566(.A(q_in_1566), .Y(WX11061));
CLKBUFX1 gbuf_d_1567(.A(n_2091), .Y(d_out_1567));
CLKBUFX1 gbuf_q_1567(.A(q_in_1567), .Y(WX11059));
CLKBUFX1 gbuf_d_1568(.A(n_2060), .Y(d_out_1568));
CLKBUFX1 gbuf_q_1568(.A(q_in_1568), .Y(WX11065));
CLKBUFX1 gbuf_d_1569(.A(n_1938), .Y(d_out_1569));
CLKBUFX1 gbuf_q_1569(.A(q_in_1569), .Y(WX11067));
CLKBUFX1 gbuf_d_1570(.A(n_2441), .Y(d_out_1570));
CLKBUFX1 gbuf_q_1570(.A(q_in_1570), .Y(WX11069));
CLKBUFX1 gbuf_d_1571(.A(n_1872), .Y(d_out_1571));
CLKBUFX1 gbuf_q_1571(.A(q_in_1571), .Y(WX11073));
CLKBUFX1 gbuf_d_1572(.A(n_2219), .Y(d_out_1572));
CLKBUFX1 gbuf_q_1572(.A(q_in_1572), .Y(WX11075));
CLKBUFX1 gbuf_d_1573(.A(n_1819), .Y(d_out_1573));
CLKBUFX1 gbuf_q_1573(.A(q_in_1573), .Y(WX11077));
CLKBUFX1 gbuf_d_1574(.A(n_2051), .Y(d_out_1574));
CLKBUFX1 gbuf_q_1574(.A(q_in_1574), .Y(WX11081));
CLKBUFX1 gbuf_d_1575(.A(n_1800), .Y(d_out_1575));
CLKBUFX1 gbuf_q_1575(.A(q_in_1575), .Y(WX11085));
CLKBUFX1 gbuf_d_1576(.A(n_2187), .Y(d_out_1576));
CLKBUFX1 gbuf_q_1576(.A(q_in_1576), .Y(WX11089));
CLKBUFX1 gbuf_d_1577(.A(n_2106), .Y(d_out_1577));
CLKBUFX1 gbuf_q_1577(.A(q_in_1577), .Y(WX11093));
CLKBUFX1 gbuf_d_1578(.A(n_2401), .Y(d_out_1578));
CLKBUFX1 gbuf_q_1578(.A(q_in_1578), .Y(WX11097));
CLKBUFX1 gbuf_d_1579(.A(n_1715), .Y(d_out_1579));
CLKBUFX1 gbuf_q_1579(.A(q_in_1579), .Y(WX11099));
CLKBUFX1 gbuf_d_1580(.A(n_1711), .Y(d_out_1580));
CLKBUFX1 gbuf_q_1580(.A(q_in_1580), .Y(WX11103));
CLKBUFX1 gbuf_d_1581(.A(n_1526), .Y(d_out_1581));
CLKBUFX1 gbuf_qn_1581(.A(qn_in_1581), .Y(WX9554));
CLKBUFX1 gbuf_d_1582(.A(n_1987), .Y(d_out_1582));
CLKBUFX1 gbuf_qn_1582(.A(qn_in_1582), .Y(WX4390));
CLKBUFX1 gbuf_d_1583(.A(n_2092), .Y(d_out_1583));
CLKBUFX1 gbuf_q_1583(.A(q_in_1583), .Y(WX3455));
CLKBUFX1 gbuf_d_1584(.A(n_1950), .Y(d_out_1584));
CLKBUFX1 gbuf_q_1584(.A(q_in_1584), .Y(WX4598));
CLKBUFX1 gbuf_d_1585(.A(n_1796), .Y(d_out_1585));
CLKBUFX1 gbuf_q_1585(.A(q_in_1585), .Y(WX11083));
CLKBUFX1 gbuf_d_1586(.A(n_1756), .Y(d_out_1586));
CLKBUFX1 gbuf_q_1586(.A(q_in_1586), .Y(WX11087));
CLKBUFX1 gbuf_d_1587(.A(n_1902), .Y(d_out_1587));
CLKBUFX1 gbuf_q_1587(.A(q_in_1587), .Y(WX7350));
CLKBUFX1 gbuf_d_1588(.A(n_2146), .Y(d_out_1588));
CLKBUFX1 gbuf_q_1588(.A(q_in_1588), .Y(WX11091));
CLKBUFX1 gbuf_d_1589(.A(n_1628), .Y(d_out_1589));
CLKBUFX1 gbuf_q_1589(.A(q_in_1589), .Y(_2166_));
CLKBUFX1 gbuf_d_1590(.A(n_1478), .Y(d_out_1590));
CLKBUFX1 gbuf_q_1590(.A(q_in_1590), .Y(WX4712));
CLKBUFX1 gbuf_d_1591(.A(n_1626), .Y(d_out_1591));
CLKBUFX1 gbuf_q_1591(.A(q_in_1591), .Y(_2168_));
CLKBUFX1 gbuf_d_1592(.A(n_1600), .Y(d_out_1592));
CLKBUFX1 gbuf_q_1592(.A(q_in_1592), .Y(_2204_));
CLKBUFX1 gbuf_d_1593(.A(n_1842), .Y(d_out_1593));
CLKBUFX1 gbuf_q_1593(.A(q_in_1593), .Y(WX8485));
BUFX3 g63216(.A (n_2894), .Y (n_4058));
CLKBUFX3 g63214(.A (n_2894), .Y (n_3168));
CLKBUFX1 gbuf_d_1594(.A(n_2334), .Y(d_out_1594));
CLKBUFX1 gbuf_q_1594(.A(q_in_1594), .Y(WX9886));
CLKBUFX1 gbuf_d_1595(.A(n_1548), .Y(d_out_1595));
CLKBUFX1 gbuf_q_1595(.A(q_in_1595), .Y(_2315_));
CLKBUFX1 gbuf_d_1596(.A(n_2099), .Y(d_out_1596));
CLKBUFX1 gbuf_q_1596(.A(q_in_1596), .Y(WX4742));
INVX4 g63152(.A (n_2897), .Y (n_5242));
CLKBUFX1 gbuf_d_1597(.A(n_2144), .Y(d_out_1597));
CLKBUFX1 gbuf_qn_1597(.A(qn_in_1597), .Y(WX5681));
INVX2 g63175(.A (n_6437), .Y (n_4670));
BUFX3 g63192(.A (n_6452), .Y (n_4017));
INVX2 g63190(.A (n_6452), .Y (n_3169));
BUFX3 g63191(.A (n_6452), .Y (n_4095));
CLKBUFX1 gbuf_d_1598(.A(n_2076), .Y(d_out_1598));
CLKBUFX1 gbuf_q_1598(.A(q_in_1598), .Y(WX11141));
BUFX3 g63186(.A (n_6452), .Y (n_4103));
CLKBUFX1 gbuf_d_1599(.A(n_1700), .Y(d_out_1599));
CLKBUFX1 gbuf_q_1599(.A(q_in_1599), .Y(WX9844));
CLKBUFX1 gbuf_d_1600(.A(n_1546), .Y(d_out_1600));
CLKBUFX1 gbuf_q_1600(.A(q_in_1600), .Y(_2318_));
BUFX3 g63185(.A (n_6452), .Y (n_4104));
CLKBUFX1 gbuf_d_1601(.A(n_1570), .Y(d_out_1601));
CLKBUFX1 gbuf_q_1601(.A(q_in_1601), .Y(_2206_));
CLKBUFX1 gbuf_d_1602(.A(n_1994), .Y(d_out_1602));
CLKBUFX1 gbuf_q_1602(.A(q_in_1602), .Y(WX7356));
CLKBUFX1 gbuf_d_1603(.A(n_1888), .Y(d_out_1603));
CLKBUFX1 gbuf_q_1603(.A(q_in_1603), .Y(WX9922));
INVX2 g63154(.A (n_2897), .Y (n_5709));
CLKBUFX1 gbuf_d_1604(.A(n_1780), .Y(d_out_1604));
CLKBUFX1 gbuf_q_1604(.A(q_in_1604), .Y(WX9878));
CLKBUFX1 gbuf_d_1605(.A(n_2082), .Y(d_out_1605));
CLKBUFX1 gbuf_q_1605(.A(q_in_1605), .Y(WX4774));
CLKBUFX1 gbuf_d_1606(.A(n_2210), .Y(d_out_1606));
CLKBUFX1 gbuf_q_1606(.A(q_in_1606), .Y(WX7208));
CLKBUFX1 gbuf_d_1607(.A(n_1884), .Y(d_out_1607));
CLKBUFX1 gbuf_q_1607(.A(q_in_1607), .Y(WX4766));
INVX1 g63156(.A (n_2897), .Y (n_5843));
CLKBUFX1 gbuf_d_1608(.A(n_1287), .Y(d_out_1608));
CLKBUFX1 gbuf_q_1608(.A(q_in_1608), .Y(WX2040));
CLKBUFX1 gbuf_d_1609(.A(n_1464), .Y(d_out_1609));
CLKBUFX1 gbuf_q_1609(.A(q_in_1609), .Y(WX5657));
CLKBUFX1 gbuf_d_1610(.A(n_1280), .Y(d_out_1610));
CLKBUFX1 gbuf_q_1610(.A(q_in_1610), .Y(WX877));
CLKBUFX1 gbuf_d_1611(.A(n_1448), .Y(d_out_1611));
CLKBUFX1 gbuf_q_1611(.A(q_in_1611), .Y(WX887));
CLKBUFX1 gbuf_d_1612(.A(n_1326), .Y(d_out_1612));
CLKBUFX1 gbuf_q_1612(.A(q_in_1612), .Y(WX711));
CLKBUFX1 gbuf_d_1613(.A(n_1366), .Y(d_out_1613));
CLKBUFX1 gbuf_q_1613(.A(q_in_1613), .Y(WX857));
INVX8 g63078(.A (n_2840), .Y (n_4562));
CLKBUFX1 gbuf_d_1614(.A(n_1407), .Y(d_out_1614));
CLKBUFX1 gbuf_q_1614(.A(q_in_1614), .Y(WX799));
CLKBUFX1 gbuf_d_1615(.A(n_1330), .Y(d_out_1615));
CLKBUFX1 gbuf_q_1615(.A(q_in_1615), .Y(WX743));
INVX1 g63071(.A (n_2840), .Y (n_3158));
CLKBUFX1 gbuf_d_1616(.A(n_1459), .Y(d_out_1616));
CLKBUFX1 gbuf_q_1616(.A(q_in_1616), .Y(WX6950));
MX2X1 g60709(.A (n_2838), .B (n_2837), .S0 (WX8457), .Y (n_2839));
MX2X1 g60712(.A (n_2813), .B (n_2953), .S0 (WX8459), .Y (n_2836));
CLKBUFX1 gbuf_d_1617(.A(n_1353), .Y(d_out_1617));
CLKBUFX1 gbuf_q_1617(.A(q_in_1617), .Y(WX875));
MX2X1 g60741(.A (n_2813), .B (n_2817), .S0 (WX4558), .Y (n_2835));
MX2X1 g60744(.A (n_2935), .B (n_2770), .S0 (WX3263), .Y (n_2833));
MX2X1 g60747(.A (n_3140), .B (n_2826), .S0 (WX9696), .Y (n_2831));
CLKBUFX1 gbuf_d_1618(.A(n_1382), .Y(d_out_1618));
CLKBUFX1 gbuf_q_1618(.A(q_in_1618), .Y(WX713));
BUFX3 g63052(.A (n_2840), .Y (n_4100));
MX2X1 g60754(.A (n_2829), .B (n_2828), .S0 (WX4562), .Y (n_2830));
MX2X1 g60757(.A (n_2826), .B (n_860), .S0 (n_2825), .Y (n_2827));
BUFX3 g63050(.A (n_2840), .Y (n_4094));
MX2X1 g60765(.A (n_2838), .B (n_3089), .S0 (WX4564), .Y (n_2824));
MX2X1 g60766(.A (n_3137), .B (n_2800), .S0 (WX9704), .Y (n_2823));
MX2X1 g60770(.A (n_2776), .B (n_2770), .S0 (WX5855), .Y (n_2822));
MX2X1 g60773(.A (n_2809), .B (n_3089), .S0 (WX4566), .Y (n_2820));
MX2X1 g60781(.A (n_2776), .B (n_2817), .S0 (WX4568), .Y (n_2818));
MX2X1 g60784(.A (n_2815), .B (n_2828), .S0 (WX4570), .Y (n_2816));
MX2X1 g60787(.A (n_2813), .B (n_2770), .S0 (WX4572), .Y (n_2814));
MX2X1 g60797(.A (n_3140), .B (n_2826), .S0 (WX9724), .Y (n_2812));
MX2X1 g60800(.A (n_6422), .B (n_3140), .S0 (n_1337), .Y (n_2811));
MX2X1 g60803(.A (n_2809), .B (n_2775), .S0 (WX4576), .Y (n_2810));
MX2X1 g60813(.A (n_2826), .B (n_860), .S0 (n_1335), .Y (n_2807));
MX2X1 g60822(.A (n_2935), .B (n_3089), .S0 (WX9740), .Y (n_2806));
MX2X1 g60827(.A (n_2716), .B (n_2795), .S0 (WX9742), .Y (n_2805));
MX2X1 g60832(.A (n_6422), .B (n_860), .S0 (n_1359), .Y (n_2803));
MX2X1 g60833(.A (n_3120), .B (n_2800), .S0 (WX10991), .Y (n_2801));
MX2X1 g60834(.A (n_2798), .B (n_2795), .S0 (WX5853), .Y (n_2799));
MX2X1 g60835(.A (n_2935), .B (n_2795), .S0 (WX9746), .Y (n_2797));
MX2X1 g60837(.A (n_3120), .B (n_2800), .S0 (WX3235), .Y (n_2794));
MX2X1 g60840(.A (n_2798), .B (n_2770), .S0 (WX9748), .Y (n_2793));
CLKBUFX1 gbuf_d_1619(.A(n_1454), .Y(d_out_1619));
CLKBUFX1 gbuf_q_1619(.A(q_in_1619), .Y(WX8243));
MX2X1 g60853(.A (n_2813), .B (n_2837), .S0 (WX9754), .Y (n_2792));
MX2X1 g60880(.A (n_6422), .B (n_860), .S0 (n_1357), .Y (n_2791));
MX2X1 g60888(.A (n_2815), .B (n_6512), .S0 (WX5871), .Y (n_2790));
MX2X1 g60899(.A (n_2826), .B (n_6432), .S0 (n_1284), .Y (n_2789));
MX2X1 g60905(.A (n_2744), .B (n_2757), .S0 (n_1431), .Y (n_2788));
MX2X1 g60907(.A (n_2826), .B (n_858), .S0 (n_1341), .Y (n_2787));
MX2X1 g60909(.A (n_2826), .B (n_3140), .S0 (n_1412), .Y (n_2786));
CLKBUFX1 gbuf_d_1620(.A(n_1389), .Y(d_out_1620));
CLKBUFX1 gbuf_q_1620(.A(q_in_1620), .Y(WX753));
MX2X1 g60920(.A (n_3027), .B (n_2826), .S0 (WX5839), .Y (n_2784));
MX2X1 g60926(.A (n_3021), .B (n_2826), .S0 (WX3249), .Y (n_2783));
CLKBUFX1 gbuf_d_1621(.A(n_1404), .Y(d_out_1621));
CLKBUFX1 gbuf_q_1621(.A(q_in_1621), .Y(WX733));
MX2X1 g60938(.A (n_2744), .B (n_2757), .S0 (n_1350), .Y (n_2782));
MX2X1 g60944(.A (n_2829), .B (n_2953), .S0 (WX5859), .Y (n_2780));
MX2X1 g60945(.A (n_2826), .B (n_858), .S0 (n_1345), .Y (n_2778));
MX2X1 g60957(.A (n_2776), .B (n_2775), .S0 (WX5869), .Y (n_2777));
CLKBUFX1 gbuf_d_1622(.A(n_1418), .Y(d_out_1622));
CLKBUFX1 gbuf_q_1622(.A(q_in_1622), .Y(WX751));
MX2X1 g60966(.A (n_2826), .B (n_858), .S0 (n_1427), .Y (n_2774));
MX2X1 g60970(.A (n_2826), .B (n_6432), .S0 (n_1419), .Y (n_2773));
MX2X1 g60971(.A (n_2744), .B (n_2757), .S0 (n_1451), .Y (n_2772));
MX2X1 g60975(.A (n_2776), .B (n_2770), .S0 (WX5867), .Y (n_2771));
MX2X1 g60978(.A (n_2776), .B (n_2795), .S0 (WX5851), .Y (n_2769));
MX2X1 g60981(.A (n_2826), .B (n_858), .S0 (n_1323), .Y (n_2768));
MX2X1 g60995(.A (n_2744), .B (n_2757), .S0 (n_1348), .Y (n_2767));
MX2X1 g60996(.A (n_2838), .B (n_2817), .S0 (WX5873), .Y (n_2765));
CLKBUFX1 gbuf_d_1623(.A(n_1319), .Y(d_out_1623));
CLKBUFX1 gbuf_q_1623(.A(q_in_1623), .Y(WX2060));
MX2X1 g61001(.A (n_6423), .B (n_2800), .S0 (WX3251), .Y (n_2763));
MX2X1 g61002(.A (n_6423), .B (n_2800), .S0 (WX11017), .Y (n_2762));
MX2X1 g61013(.A (n_2813), .B (n_2837), .S0 (WX3269), .Y (n_2761));
MX2X1 g61021(.A (n_2716), .B (n_2988), .S0 (WX8455), .Y (n_2760));
MX2X1 g61022(.A (n_2744), .B (n_2757), .S0 (n_1286), .Y (n_2759));
MX2X1 g61032(.A (n_2829), .B (n_2755), .S0 (WX3271), .Y (n_2756));
MX2X1 g61040(.A (n_2744), .B (n_2757), .S0 (n_1374), .Y (n_2754));
MX2X1 g61044(.A (n_2815), .B (n_3089), .S0 (WX11021), .Y (n_2752));
MX2X1 g61048(.A (n_2744), .B (n_2757), .S0 (n_1288), .Y (n_2750));
CLKBUFX1 gbuf_d_1624(.A(n_1340), .Y(d_out_1624));
CLKBUFX1 gbuf_q_1624(.A(q_in_1624), .Y(WX2008));
MX2X1 g61051(.A (n_2809), .B (n_2988), .S0 (WX9744), .Y (n_2749));
MX2X1 g61056(.A (n_2809), .B (n_2817), .S0 (WX8453), .Y (n_2746));
CLKBUFX1 gbuf_d_1625(.A(n_1453), .Y(d_out_1625));
CLKBUFX1 gbuf_q_1625(.A(q_in_1625), .Y(WX9536));
MX2X1 g61080(.A (n_2744), .B (n_2757), .S0 (n_1309), .Y (n_2745));
MX2X1 g61088(.A (n_2744), .B (n_2757), .S0 (n_1282), .Y (n_2743));
MX2X1 g61095(.A (n_2986), .B (n_2953), .S0 (WX11025), .Y (n_2742));
MX2X1 g61097(.A (n_2986), .B (n_6512), .S0 (WX3277), .Y (n_2741));
MX2X1 g61103(.A (n_2776), .B (n_6512), .S0 (WX8451), .Y (n_2739));
MX2X1 g61106(.A (n_6513), .B (n_2770), .S0 (WX3279), .Y (n_2738));
MX2X1 g61113(.A (n_2744), .B (n_2757), .S0 (n_2691), .Y (n_2737));
MX2X1 g61115(.A (n_2813), .B (n_2953), .S0 (WX11027), .Y (n_2736));
MX2X1 g61121(.A (n_2829), .B (n_2953), .S0 (WX8447), .Y (n_2734));
MX2X1 g61122(.A (n_2744), .B (n_2757), .S0 (n_1442), .Y (n_2733));
MX2X1 g61123(.A (n_2798), .B (n_2837), .S0 (WX7154), .Y (n_2732));
MX2X1 g61133(.A (n_2744), .B (n_2757), .S0 (n_1328), .Y (n_2731));
MX2X1 g61134(.A (n_2815), .B (n_2988), .S0 (WX7160), .Y (n_2730));
MX2X1 g61142(.A (n_2935), .B (n_2775), .S0 (WX3283), .Y (n_2729));
MX2X1 g61144(.A (n_2716), .B (n_2817), .S0 (WX7164), .Y (n_2728));
MX2X1 g61146(.A (n_6422), .B (n_860), .S0 (n_1339), .Y (n_2726));
MX2X1 g61154(.A (n_2809), .B (n_2755), .S0 (WX7168), .Y (n_2725));
MX2X1 g61160(.A (n_2744), .B (n_2757), .S0 (n_1437), .Y (n_2724));
MX2X1 g61161(.A (n_2798), .B (n_2775), .S0 (WX7170), .Y (n_2722));
MX2X1 g61170(.A (n_2744), .B (n_2757), .S0 (n_1429), .Y (n_2721));
MX2X1 g61173(.A (n_2815), .B (n_2988), .S0 (WX3287), .Y (n_2720));
CLKBUFX1 gbuf_d_1626(.A(n_1447), .Y(d_out_1626));
CLKBUFX1 gbuf_q_1626(.A(q_in_1626), .Y(WX833));
MX2X1 g61177(.A (n_2716), .B (n_2770), .S0 (WX3289), .Y (n_2719));
MX2X1 g61178(.A (n_2744), .B (n_2757), .S0 (n_1318), .Y (n_2718));
CLKBUFX1 gbuf_d_1627(.A(n_1321), .Y(d_out_1627));
CLKBUFX1 gbuf_q_1627(.A(q_in_1627), .Y(WX2024));
MX2X1 g61184(.A (n_2716), .B (n_2775), .S0 (WX3291), .Y (n_2717));
MX2X1 g61192(.A (n_2744), .B (n_2757), .S0 (n_2675), .Y (n_2715));
CLKBUFX1 gbuf_d_1628(.A(n_1289), .Y(d_out_1628));
CLKBUFX1 gbuf_q_1628(.A(q_in_1628), .Y(WX2044));
MX2X1 g61200(.A (n_2826), .B (n_3140), .S0 (n_1449), .Y (n_2714));
MX2X1 g61201(.A (n_2815), .B (n_2795), .S0 (WX11041), .Y (n_2713));
MX2X1 g61202(.A (n_2798), .B (n_2837), .S0 (WX8443), .Y (n_2712));
MX2X1 g61206(.A (n_2815), .B (n_2817), .S0 (WX4580), .Y (n_2711));
MX2X1 g61208(.A (n_2813), .B (n_2988), .S0 (WX11043), .Y (n_2710));
MX2X1 g61213(.A (n_3137), .B (n_2826), .S0 (WX3233), .Y (n_2709));
MX2X1 g61227(.A (n_2809), .B (n_2828), .S0 (WX9738), .Y (n_2708));
MX2X1 g61230(.A (n_3021), .B (n_2826), .S0 (WX8415), .Y (n_2707));
MX2X1 g61234(.A (n_3137), .B (n_2826), .S0 (WX8417), .Y (n_2706));
MX2X1 g61237(.A (n_2716), .B (n_2795), .S0 (WX11047), .Y (n_2705));
MX2X1 g61239(.A (n_3137), .B (n_2826), .S0 (WX8419), .Y (n_2704));
CLKBUFX1 gbuf_d_1629(.A(n_1388), .Y(d_out_1629));
CLKBUFX1 gbuf_q_1629(.A(q_in_1629), .Y(WX803));
MX2X1 g61246(.A (n_2826), .B (n_3140), .S0 (n_1320), .Y (n_2703));
MX2X1 g61249(.A (n_3140), .B (n_2800), .S0 (WX4524), .Y (n_2702));
MX2X1 g61258(.A (n_2716), .B (n_2775), .S0 (WX11049), .Y (n_2701));
MX2X1 g61265(.A (n_2826), .B (n_6432), .S0 (n_1421), .Y (n_2700));
CLKBUFX1 gbuf_d_1630(.A(n_1452), .Y(d_out_1630));
CLKBUFX1 gbuf_q_1630(.A(q_in_1630), .Y(WX2062));
CLKBUFX1 gbuf_d_1631(.A(n_1365), .Y(d_out_1631));
CLKBUFX1 gbuf_q_1631(.A(q_in_1631), .Y(WX719));
MX2X1 g61274(.A (n_2809), .B (n_2755), .S0 (WX9734), .Y (n_2699));
MX2X1 g61276(.A (n_2829), .B (n_2755), .S0 (WX11051), .Y (n_2698));
MX2X1 g61279(.A (n_2935), .B (n_2817), .S0 (WX8435), .Y (n_2697));
MX2X1 g61288(.A (n_2716), .B (n_2755), .S0 (WX8439), .Y (n_2696));
MX2X1 g61300(.A (n_3137), .B (n_2800), .S0 (WX3257), .Y (n_2695));
MX2X1 g61304(.A (n_2935), .B (n_2953), .S0 (WX9758), .Y (n_2694));
CLKBUFX1 gbuf_d_1632(.A(n_1423), .Y(d_out_1632));
CLKBUFX1 gbuf_q_1632(.A(q_in_1632), .Y(WX723));
CLKBUFX1 gbuf_d_1633(.A(n_1380), .Y(d_out_1633));
CLKBUFX1 gbuf_q_1633(.A(q_in_1633), .Y(WX889));
BUFX3 g61384(.A (n_7089), .Y (n_2926));
BUFX3 g61393(.A (n_7089), .Y (n_2925));
BUFX3 g61402(.A (n_7089), .Y (n_2924));
BUFX3 g61420(.A (n_7089), .Y (n_2922));
BUFX3 g61429(.A (n_7089), .Y (n_2921));
BUFX3 g61456(.A (n_7089), .Y (n_2920));
CLKBUFX1 gbuf_d_1634(.A(n_1324), .Y(d_out_1634));
CLKBUFX1 gbuf_q_1634(.A(q_in_1634), .Y(WX2028));
NOR2X1 g61542(.A (n_2691), .B (n_3188), .Y (n_2692));
CLKBUFX1 gbuf_d_1635(.A(n_1435), .Y(d_out_1635));
CLKBUFX1 gbuf_q_1635(.A(q_in_1635), .Y(WX871));
AND2X1 g61572(.A (WX11175), .B (n_2298), .Y (n_2690));
AND2X1 g61573(.A (WX11089), .B (n_2298), .Y (n_2689));
AND2X1 g61577(.A (WX9770), .B (n_2298), .Y (n_2687));
CLKBUFX1 gbuf_d_1636(.A(n_1399), .Y(d_out_1636));
CLKBUFX1 gbuf_q_1636(.A(q_in_1636), .Y(WX865));
AND2X1 g61638(.A (WX11135), .B (n_2298), .Y (n_2686));
CLKBUFX1 gbuf_d_1637(.A(n_1362), .Y(d_out_1637));
CLKBUFX1 gbuf_q_1637(.A(q_in_1637), .Y(WX897));
AND2X1 g61647(.A (WX4556), .B (n_2298), .Y (n_2685));
AND2X1 g61648(.A (WX11143), .B (n_2298), .Y (n_2684));
CLKBUFX1 gbuf_d_1638(.A(n_1400), .Y(d_out_1638));
CLKBUFX1 gbuf_q_1638(.A(q_in_1638), .Y(WX793));
AND2X1 g61675(.A (WX4542), .B (n_2298), .Y (n_2682));
AND2X1 g61676(.A (WX9808), .B (n_2298), .Y (n_2681));
AND2X1 g61716(.A (WX11105), .B (n_2298), .Y (n_2680));
AND2X1 g58600(.A (WX11117), .B (n_2298), .Y (n_2678));
CLKBUFX1 gbuf_d_1639(.A(n_1398), .Y(d_out_1639));
CLKBUFX1 gbuf_q_1639(.A(q_in_1639), .Y(WX869));
AND2X1 g61801(.A (WX7152), .B (n_2298), .Y (n_2677));
NOR2X1 g61817(.A (n_2675), .B (n_3188), .Y (n_2676));
CLKBUFX1 gbuf_d_1640(.A(n_1338), .Y(d_out_1640));
CLKBUFX1 gbuf_q_1640(.A(q_in_1640), .Y(WX2002));
CLKBUFX1 gbuf_d_1641(.A(n_1422), .Y(d_out_1641));
CLKBUFX1 gbuf_q_1641(.A(q_in_1641), .Y(WX2020));
CLKBUFX1 gbuf_d_1642(.A(n_1279), .Y(d_out_1642));
CLKBUFX1 gbuf_q_1642(.A(q_in_1642), .Y(WX3071));
AND2X1 g61914(.A (WX9862), .B (n_2378), .Y (n_2673));
AND2X1 g61934(.A (WX9764), .B (n_2378), .Y (n_2671));
AND2X1 g61960(.A (WX4682), .B (n_2298), .Y (n_2670));
AND2X1 g61964(.A (WX4690), .B (n_2378), .Y (n_2669));
AND2X1 g62074(.A (WX3375), .B (n_2298), .Y (n_2668));
AND2X1 g62097(.A (WX3369), .B (n_2298), .Y (n_2667));
AND2X1 g62137(.A (WX3305), .B (n_2298), .Y (n_2666));
CLKBUFX1 gbuf_d_1643(.A(n_1329), .Y(d_out_1643));
CLKBUFX1 gbuf_q_1643(.A(q_in_1643), .Y(WX2054));
CLKBUFX1 gbuf_d_1644(.A(n_1438), .Y(d_out_1644));
CLKBUFX1 gbuf_q_1644(.A(q_in_1644), .Y(WX2056));
AND2X1 g62215(.A (WX4610), .B (n_2378), .Y (n_2665));
AND2X1 g62219(.A (WX5987), .B (n_2378), .Y (n_2664));
AND2X1 g62221(.A (WX11051), .B (n_2378), .Y (n_2663));
CLKBUFX1 gbuf_d_1645(.A(n_1327), .Y(d_out_1645));
CLKBUFX1 gbuf_q_1645(.A(q_in_1645), .Y(WX853));
CLKBUFX1 gbuf_d_1646(.A(n_1432), .Y(d_out_1646));
CLKBUFX1 gbuf_q_1646(.A(q_in_1646), .Y(WX2036));
CLKBUFX1 gbuf_d_1647(.A(n_1333), .Y(d_out_1647));
CLKBUFX1 gbuf_q_1647(.A(q_in_1647), .Y(WX849));
XOR2X1 g58894(.A (_2119_), .B (n_1221), .Y (n_2662));
XOR2X1 g58895(.A (_2183_), .B (n_1044), .Y (n_2661));
AND2X1 g62490(.A (WX8585), .B (n_2298), .Y (n_2660));
AND2X1 g62491(.A (WX8587), .B (n_2298), .Y (n_2659));
XOR2X1 g58896(.A (_2112_), .B (n_1254), .Y (n_2658));
XOR2X1 g58897(.A (_2284_), .B (n_1111), .Y (n_2657));
XOR2X1 g58900(.A (_2124_), .B (n_1231), .Y (n_2656));
XOR2X1 g58901(.A (_2144_), .B (n_1047), .Y (n_2655));
XOR2X1 g58902(.A (_2151_), .B (n_1186), .Y (n_2654));
XOR2X1 g58903(.A (_2156_), .B (n_1181), .Y (n_2653));
XOR2X1 g58904(.A (_2176_), .B (n_1210), .Y (n_2652));
XOR2X1 g58905(.A (_2188_), .B (n_1257), .Y (n_2651));
AND2X1 g62520(.A (WX11171), .B (n_2298), .Y (n_2650));
XOR2X1 g58906(.A (_2208_), .B (n_1154), .Y (n_2649));
XOR2X1 g58907(.A (_2247_), .B (n_1237), .Y (n_2648));
XOR2X1 g58908(.A (_2215_), .B (n_1150), .Y (n_2647));
XOR2X1 g58909(.A (_2220_), .B (n_1148), .Y (n_2646));
AND2X1 g62532(.A (WX3337), .B (n_2298), .Y (n_2645));
XOR2X1 g58910(.A (_2240_), .B (n_1135), .Y (n_2644));
XOR2X1 g58911(.A (_2252_), .B (n_1116), .Y (n_2643));
XOR2X1 g58912(.A (_2272_), .B (n_1120), .Y (n_2642));
XOR2X1 g58913(.A (_2279_), .B (n_1114), .Y (n_2641));
XOR2X1 g58914(.A (_2311_), .B (n_1094), .Y (n_2640));
XOR2X1 g58915(.A (_2336_), .B (n_1082), .Y (n_2639));
AND2X1 g62550(.A (WX5863), .B (n_2298), .Y (n_2638));
XOR2X1 g58916(.A (_2343_), .B (n_1079), .Y (n_2637));
XOR2X1 g58917(.A (_2348_), .B (n_1076), .Y (n_2636));
XOR2X1 g58918(.A (_2304_), .B (n_1051), .Y (n_2635));
XOR2X1 g58919(.A (_2316_), .B (n_1091), .Y (n_2634));
CLKBUFX1 gbuf_d_1648(.A(n_1314), .Y(d_out_1648));
CLKBUFX1 gbuf_q_1648(.A(q_in_1648), .Y(WX829));
AND2X1 g62615(.A (WX2034), .B (n_2298), .Y (n_2633));
AND2X1 g62680(.A (WX2082), .B (n_2298), .Y (n_2632));
CLKBUFX1 gbuf_d_1649(.A(n_1458), .Y(d_out_1649));
CLKBUFX1 gbuf_q_1649(.A(q_in_1649), .Y(WX827));
CLKBUFX1 gbuf_d_1650(.A(n_1428), .Y(d_out_1650));
CLKBUFX1 gbuf_q_1650(.A(q_in_1650), .Y(WX2030));
CLKBUFX1 gbuf_d_1651(.A(n_1373), .Y(d_out_1651));
CLKBUFX1 gbuf_q_1651(.A(q_in_1651), .Y(WX747));
CLKBUFX1 gbuf_d_1652(.A(n_1342), .Y(d_out_1652));
CLKBUFX1 gbuf_q_1652(.A(q_in_1652), .Y(WX2016));
CLKBUFX1 gbuf_d_1653(.A(n_1347), .Y(d_out_1653));
CLKBUFX1 gbuf_q_1653(.A(q_in_1653), .Y(WX861));
CLKBUFX1 gbuf_d_1654(.A(n_1415), .Y(d_out_1654));
CLKBUFX1 gbuf_q_1654(.A(q_in_1654), .Y(WX795));
CLKBUFX1 gbuf_d_1655(.A(n_1332), .Y(d_out_1655));
CLKBUFX1 gbuf_q_1655(.A(q_in_1655), .Y(WX735));
CLKBUFX1 gbuf_d_1656(.A(n_1410), .Y(d_out_1656));
CLKBUFX1 gbuf_q_1656(.A(q_in_1656), .Y(WX883));
CLKBUFX1 gbuf_d_1657(.A(n_1378), .Y(d_out_1657));
CLKBUFX1 gbuf_q_1657(.A(q_in_1657), .Y(WX787));
CLKBUFX1 gbuf_d_1658(.A(n_1411), .Y(d_out_1658));
CLKBUFX1 gbuf_q_1658(.A(q_in_1658), .Y(WX825));
CLKBUFX1 g63148(.A (n_6437), .Y (n_3162));
CLKBUFX1 gbuf_d_1659(.A(n_1354), .Y(d_out_1659));
CLKBUFX1 gbuf_q_1659(.A(q_in_1659), .Y(WX839));
CLKBUFX1 gbuf_d_1660(.A(n_1436), .Y(d_out_1660));
CLKBUFX1 gbuf_q_1660(.A(q_in_1660), .Y(WX821));
CLKBUFX1 gbuf_d_1661(.A(n_1409), .Y(d_out_1661));
CLKBUFX1 gbuf_q_1661(.A(q_in_1661), .Y(WX757));
NOR2X1 g57541(.A (n_848), .B (n_3188), .Y (n_2631));
BUFX3 g63051(.A (n_2840), .Y (n_4101));
BUFX3 g63053(.A (n_2840), .Y (n_4106));
CLKBUFX1 gbuf_d_1662(.A(n_1433), .Y(d_out_1662));
CLKBUFX1 gbuf_q_1662(.A(q_in_1662), .Y(WX731));
CLKBUFX1 gbuf_d_1663(.A(n_1444), .Y(d_out_1663));
CLKBUFX1 gbuf_q_1663(.A(q_in_1663), .Y(WX783));
AND2X1 g62721(.A (WX7208), .B (n_2298), .Y (n_2630));
NOR2X1 g59242(.A (n_1195), .B (n_3188), .Y (n_2629));
NOR2X1 g59244(.A (n_1104), .B (n_2620), .Y (n_2628));
CLKBUFX1 gbuf_d_1664(.A(n_1364), .Y(d_out_1664));
CLKBUFX1 gbuf_q_1664(.A(q_in_1664), .Y(WX737));
NOR2X1 g59248(.A (n_1097), .B (n_3188), .Y (n_2627));
NOR2X1 g59249(.A (n_1065), .B (n_3690), .Y (n_2626));
NOR2X1 g59250(.A (n_1131), .B (n_3690), .Y (n_2625));
NOR2X1 g59251(.A (n_1245), .B (n_2851), .Y (n_2624));
NOR2X1 g59257(.A (n_1233), .B (n_3690), .Y (n_2622));
NOR2X1 g59266(.A (n_1205), .B (n_2620), .Y (n_2621));
CLKBUFX1 gbuf_d_1665(.A(n_1456), .Y(d_out_1665));
CLKBUFX1 gbuf_q_1665(.A(q_in_1665), .Y(WX487));
CLKBUFX1 gbuf_d_1666(.A(n_1465), .Y(d_out_1666));
CLKBUFX1 gbuf_q_1666(.A(q_in_1666), .Y(WX855));
CLKBUFX1 gbuf_d_1667(.A(n_1393), .Y(d_out_1667));
CLKBUFX1 gbuf_q_1667(.A(q_in_1667), .Y(WX717));
CLKBUFX1 gbuf_d_1668(.A(n_1424), .Y(d_out_1668));
CLKBUFX1 gbuf_q_1668(.A(q_in_1668), .Y(WX837));
NOR2X1 g59294(.A (n_1023), .B (n_3188), .Y (n_2619));
CLKBUFX1 gbuf_d_1669(.A(n_1377), .Y(d_out_1669));
CLKBUFX1 gbuf_q_1669(.A(q_in_1669), .Y(WX823));
NOR2X1 g59320(.A (n_1176), .B (n_2620), .Y (n_2618));
NOR2X1 g59321(.A (n_1227), .B (n_2620), .Y (n_2617));
NOR2X1 g59330(.A (n_1170), .B (n_2620), .Y (n_2616));
NOR2X1 g59331(.A (n_1066), .B (n_2620), .Y (n_2615));
AND2X1 g62701(.A (WX4574), .B (n_2298), .Y (n_2614));
NOR2X1 g59347(.A (n_1032), .B (n_2620), .Y (n_2613));
NOR2X1 g59352(.A (n_1158), .B (n_2851), .Y (n_2612));
NOR2X1 g59353(.A (n_1119), .B (n_2851), .Y (n_2611));
NOR2X1 g59356(.A (n_1033), .B (n_2605), .Y (n_2610));
NOR2X1 g59357(.A (n_1155), .B (n_2851), .Y (n_2609));
NOR2X1 g59365(.A (n_1019), .B (n_3188), .Y (n_2608));
NOR2X1 g59367(.A (n_1145), .B (n_3188), .Y (n_2607));
NOR2X1 g59376(.A (n_1054), .B (n_2605), .Y (n_2606));
NOR2X1 g59378(.A (n_1136), .B (n_2851), .Y (n_2604));
NOR2X1 g59379(.A (n_1226), .B (n_2851), .Y (n_2603));
NOR2X1 g59386(.A (n_1128), .B (n_2620), .Y (n_2602));
NOR2X1 g59390(.A (n_1055), .B (n_3188), .Y (n_2601));
NOR2X1 g59391(.A (n_1142), .B (n_3188), .Y (n_2600));
NOR2X1 g59394(.A (n_1265), .B (n_2620), .Y (n_2599));
NOR2X1 g59405(.A (n_1108), .B (n_3188), .Y (n_2598));
NOR2X1 g59408(.A (n_1106), .B (n_2851), .Y (n_2597));
NOR2X1 g59409(.A (n_1228), .B (n_2620), .Y (n_2596));
NOR2X1 g59412(.A (n_1102), .B (n_2605), .Y (n_2595));
NOR2X1 g59413(.A (n_1101), .B (n_2851), .Y (n_2594));
NOR2X1 g59414(.A (n_1244), .B (n_3188), .Y (n_2593));
NOR2X1 g59415(.A (n_1182), .B (n_3188), .Y (n_2591));
NOR2X1 g59416(.A (n_1099), .B (n_3188), .Y (n_2590));
NOR2X1 g59422(.A (n_1048), .B (n_3188), .Y (n_2589));
NOR2X1 g59430(.A (n_1086), .B (n_3690), .Y (n_2588));
NOR2X1 g59431(.A (n_1020), .B (n_3690), .Y (n_2587));
NOR2X1 g59434(.A (n_1064), .B (n_3690), .Y (n_2585));
NOR2X1 g59435(.A (n_1084), .B (n_2605), .Y (n_2584));
NOR2X1 g59436(.A (n_1230), .B (n_3690), .Y (n_2583));
NOR2X1 g59437(.A (n_1083), .B (n_3690), .Y (n_2582));
NOR2X1 g59447(.A (n_1264), .B (n_2851), .Y (n_2581));
NOR2X1 g59448(.A (n_1075), .B (n_3690), .Y (n_2579));
NOR2X1 g59449(.A (n_1015), .B (n_3690), .Y (n_2577));
NOR2X1 g59450(.A (n_1074), .B (n_2620), .Y (n_2576));
NOR2X1 g59451(.A (n_1247), .B (n_2851), .Y (n_2575));
NOR2X1 g59452(.A (n_1073), .B (n_2851), .Y (n_2574));
NOR2X1 g59453(.A (n_1072), .B (n_3690), .Y (n_2573));
NOR2X1 g59460(.A (n_1132), .B (n_3690), .Y (n_2572));
NOR2X1 g59464(.A (n_1068), .B (n_2851), .Y (n_2571));
NOR2X1 g59465(.A (n_1113), .B (n_2851), .Y (n_2570));
NOR2X1 g59468(.A (n_1242), .B (n_2851), .Y (n_2568));
NOR2X1 g59469(.A (n_1268), .B (n_2851), .Y (n_2567));
NOR2X1 g59475(.A (n_1035), .B (n_3690), .Y (n_2566));
NOR2X1 g59476(.A (n_1263), .B (n_2851), .Y (n_2565));
NOR2X1 g59477(.A (n_1027), .B (n_2851), .Y (n_2564));
NOR2X1 g59478(.A (n_1168), .B (n_3690), .Y (n_2563));
CLKBUFX1 gbuf_d_1670(.A(n_1355), .Y(d_out_1670));
CLKBUFX1 gbuf_q_1670(.A(q_in_1670), .Y(WX779));
CLKBUFX1 gbuf_d_1671(.A(n_1405), .Y(d_out_1671));
CLKBUFX1 gbuf_q_1671(.A(q_in_1671), .Y(WX819));
CLKBUFX1 gbuf_d_1672(.A(n_1275), .Y(d_out_1672));
CLKBUFX1 gbuf_q_1672(.A(q_in_1672), .Y(WX771));
AND2X1 g62661(.A (WX9740), .B (n_2378), .Y (n_2562));
CLKBUFX1 gbuf_d_1673(.A(n_1344), .Y(d_out_1673));
CLKBUFX1 gbuf_q_1673(.A(q_in_1673), .Y(WX891));
CLKBUFX1 gbuf_d_1674(.A(n_1369), .Y(d_out_1674));
CLKBUFX1 gbuf_q_1674(.A(q_in_1674), .Y(WX879));
CLKBUFX1 gbuf_d_1675(.A(n_1313), .Y(d_out_1675));
CLKBUFX1 gbuf_q_1675(.A(q_in_1675), .Y(WX863));
CLKBUFX1 gbuf_d_1676(.A(n_1290), .Y(d_out_1676));
CLKBUFX1 gbuf_q_1676(.A(q_in_1676), .Y(WX773));
CLKBUFX1 gbuf_d_1677(.A(n_1312), .Y(d_out_1677));
CLKBUFX1 gbuf_q_1677(.A(q_in_1677), .Y(WX805));
CLKBUFX1 gbuf_d_1678(.A(n_1283), .Y(d_out_1678));
CLKBUFX1 gbuf_q_1678(.A(q_in_1678), .Y(WX2048));
CLKBUFX1 gbuf_d_1679(.A(n_1307), .Y(d_out_1679));
CLKBUFX1 gbuf_q_1679(.A(q_in_1679), .Y(WX815));
CLKBUFX1 gbuf_d_1680(.A(n_1311), .Y(d_out_1680));
CLKBUFX1 gbuf_q_1680(.A(q_in_1680), .Y(WX813));
CLKBUFX1 gbuf_d_1681(.A(n_1367), .Y(d_out_1681));
CLKBUFX1 gbuf_q_1681(.A(q_in_1681), .Y(WX741));
CLKBUFX1 gbuf_d_1682(.A(n_1372), .Y(d_out_1682));
CLKBUFX1 gbuf_q_1682(.A(q_in_1682), .Y(WX739));
CLKBUFX1 gbuf_d_1683(.A(n_1403), .Y(d_out_1683));
CLKBUFX1 gbuf_q_1683(.A(q_in_1683), .Y(WX749));
CLKBUFX1 gbuf_d_1684(.A(n_1396), .Y(d_out_1684));
CLKBUFX1 gbuf_q_1684(.A(q_in_1684), .Y(WX755));
CLKBUFX1 gbuf_d_1685(.A(n_1402), .Y(d_out_1685));
CLKBUFX1 gbuf_q_1685(.A(q_in_1685), .Y(WX759));
CLKBUFX1 gbuf_d_1686(.A(n_1291), .Y(d_out_1686));
CLKBUFX1 gbuf_q_1686(.A(q_in_1686), .Y(WX765));
CLKBUFX1 gbuf_d_1687(.A(n_1441), .Y(d_out_1687));
CLKBUFX1 gbuf_q_1687(.A(q_in_1687), .Y(WX769));
CLKBUFX1 gbuf_d_1688(.A(n_1322), .Y(d_out_1688));
CLKBUFX1 gbuf_q_1688(.A(q_in_1688), .Y(WX777));
CLKBUFX1 gbuf_d_1689(.A(n_1306), .Y(d_out_1689));
CLKBUFX1 gbuf_q_1689(.A(q_in_1689), .Y(WX775));
CLKBUFX1 gbuf_d_1690(.A(n_1462), .Y(d_out_1690));
CLKBUFX1 gbuf_q_1690(.A(q_in_1690), .Y(WX781));
CLKBUFX1 gbuf_d_1691(.A(n_1426), .Y(d_out_1691));
CLKBUFX1 gbuf_q_1691(.A(q_in_1691), .Y(WX785));
CLKBUFX1 gbuf_d_1692(.A(n_1334), .Y(d_out_1692));
CLKBUFX1 gbuf_q_1692(.A(q_in_1692), .Y(WX789));
CLKBUFX1 gbuf_d_1693(.A(n_1414), .Y(d_out_1693));
CLKBUFX1 gbuf_q_1693(.A(q_in_1693), .Y(WX791));
CLKBUFX1 gbuf_d_1694(.A(n_1385), .Y(d_out_1694));
CLKBUFX1 gbuf_q_1694(.A(q_in_1694), .Y(WX797));
CLKBUFX1 gbuf_d_1695(.A(n_1325), .Y(d_out_1695));
CLKBUFX1 gbuf_q_1695(.A(q_in_1695), .Y(WX801));
CLKBUFX1 gbuf_d_1696(.A(n_1391), .Y(d_out_1696));
CLKBUFX1 gbuf_q_1696(.A(q_in_1696), .Y(WX807));
CLKBUFX1 gbuf_d_1697(.A(n_1308), .Y(d_out_1697));
CLKBUFX1 gbuf_q_1697(.A(q_in_1697), .Y(WX809));
CLKBUFX1 gbuf_d_1698(.A(n_1356), .Y(d_out_1698));
CLKBUFX1 gbuf_q_1698(.A(q_in_1698), .Y(WX811));
CLKBUFX1 gbuf_d_1699(.A(n_1386), .Y(d_out_1699));
CLKBUFX1 gbuf_q_1699(.A(q_in_1699), .Y(WX817));
CLKBUFX1 gbuf_d_1700(.A(n_1387), .Y(d_out_1700));
CLKBUFX1 gbuf_q_1700(.A(q_in_1700), .Y(WX843));
CLKBUFX1 gbuf_d_1701(.A(n_1316), .Y(d_out_1701));
CLKBUFX1 gbuf_q_1701(.A(q_in_1701), .Y(WX11053));
CLKBUFX1 gbuf_d_1702(.A(n_1417), .Y(d_out_1702));
CLKBUFX1 gbuf_q_1702(.A(q_in_1702), .Y(WX851));
CLKBUFX1 gbuf_d_1703(.A(n_1379), .Y(d_out_1703));
CLKBUFX1 gbuf_q_1703(.A(q_in_1703), .Y(WX859));
CLKBUFX1 gbuf_d_1704(.A(n_1446), .Y(d_out_1704));
CLKBUFX1 gbuf_q_1704(.A(q_in_1704), .Y(WX841));
CLKBUFX1 gbuf_d_1705(.A(n_1371), .Y(d_out_1705));
CLKBUFX1 gbuf_q_1705(.A(q_in_1705), .Y(WX847));
CLKBUFX1 gbuf_d_1706(.A(n_1370), .Y(d_out_1706));
CLKBUFX1 gbuf_q_1706(.A(q_in_1706), .Y(WX881));
CLKBUFX1 gbuf_d_1707(.A(n_1384), .Y(d_out_1707));
CLKBUFX1 gbuf_q_1707(.A(q_in_1707), .Y(WX885));
CLKBUFX1 gbuf_d_1708(.A(n_1381), .Y(d_out_1708));
CLKBUFX1 gbuf_q_1708(.A(q_in_1708), .Y(WX893));
CLKBUFX1 gbuf_d_1709(.A(n_1395), .Y(d_out_1709));
CLKBUFX1 gbuf_q_1709(.A(q_in_1709), .Y(WX867));
CLKBUFX1 gbuf_d_1710(.A(n_1461), .Y(d_out_1710));
CLKBUFX1 gbuf_q_1710(.A(q_in_1710), .Y(WX761));
CLKBUFX1 gbuf_d_1711(.A(n_1440), .Y(d_out_1711));
CLKBUFX1 gbuf_q_1711(.A(q_in_1711), .Y(WX709));
CLKBUFX1 gbuf_d_1712(.A(n_1336), .Y(d_out_1712));
CLKBUFX1 gbuf_q_1712(.A(q_in_1712), .Y(WX2004));
CLKBUFX1 gbuf_d_1713(.A(n_1360), .Y(d_out_1713));
CLKBUFX1 gbuf_q_1713(.A(q_in_1713), .Y(WX2006));
CLKBUFX1 gbuf_d_1714(.A(n_1413), .Y(d_out_1714));
CLKBUFX1 gbuf_q_1714(.A(q_in_1714), .Y(WX2010));
CLKBUFX1 gbuf_d_1715(.A(n_1358), .Y(d_out_1715));
CLKBUFX1 gbuf_q_1715(.A(q_in_1715), .Y(WX2012));
CLKBUFX1 gbuf_d_1716(.A(n_1285), .Y(d_out_1716));
CLKBUFX1 gbuf_q_1716(.A(q_in_1716), .Y(WX2014));
CLKBUFX1 gbuf_d_1717(.A(n_1450), .Y(d_out_1717));
CLKBUFX1 gbuf_q_1717(.A(q_in_1717), .Y(WX2018));
CLKBUFX1 gbuf_d_1718(.A(n_1420), .Y(d_out_1718));
CLKBUFX1 gbuf_q_1718(.A(q_in_1718), .Y(WX2022));
CLKBUFX1 gbuf_d_1719(.A(n_1346), .Y(d_out_1719));
CLKBUFX1 gbuf_q_1719(.A(q_in_1719), .Y(WX2026));
CLKBUFX1 gbuf_d_1720(.A(n_1351), .Y(d_out_1720));
CLKBUFX1 gbuf_q_1720(.A(q_in_1720), .Y(WX2034));
CLKBUFX1 gbuf_d_1721(.A(n_1349), .Y(d_out_1721));
CLKBUFX1 gbuf_q_1721(.A(q_in_1721), .Y(WX2038));
CLKBUFX1 gbuf_d_1722(.A(n_1375), .Y(d_out_1722));
CLKBUFX1 gbuf_q_1722(.A(q_in_1722), .Y(WX2042));
CLKBUFX1 gbuf_d_1723(.A(n_1310), .Y(d_out_1723));
CLKBUFX1 gbuf_q_1723(.A(q_in_1723), .Y(WX2046));
CLKBUFX1 gbuf_d_1724(.A(n_1443), .Y(d_out_1724));
CLKBUFX1 gbuf_q_1724(.A(q_in_1724), .Y(WX2052));
CLKBUFX1 gbuf_d_1725(.A(n_1430), .Y(d_out_1725));
CLKBUFX1 gbuf_q_1725(.A(q_in_1725), .Y(WX2058));
CLKBUFX1 gbuf_d_1726(.A(n_1317), .Y(d_out_1726));
CLKBUFX1 gbuf_q_1726(.A(q_in_1726), .Y(WX763));
CLKBUFX1 gbuf_d_1727(.A(n_1352), .Y(d_out_1727));
CLKBUFX1 gbuf_q_1727(.A(q_in_1727), .Y(WX767));
INVX2 g63218(.A (n_6446), .Y (n_2894));
CLKBUFX1 gbuf_d_1728(.A(n_1277), .Y(d_out_1728));
CLKBUFX1 gbuf_q_1728(.A(q_in_1728), .Y(WX729));
BUFX3 g63157(.A (n_6437), .Y (n_2897));
AND2X1 g61592(.A (WX7238), .B (n_2527), .Y (n_2559));
AND2X1 g62609(.A (WX8505), .B (n_2346), .Y (n_2558));
AOI21X1 g60399(.A0 (_2100_), .A1 (WX851), .B0 (n_897), .Y (n_2557));
AND2X1 g61587(.A (WX9708), .B (n_2400), .Y (n_2556));
AOI21X1 g60402(.A0 (_2096_), .A1 (WX859), .B0 (n_895), .Y (n_2555));
AOI21X1 g60405(.A0 (_2086_), .A1 (WX879), .B0 (n_900), .Y (n_2554));
AND2X1 g61585(.A (WX11095), .B (n_2346), .Y (n_2553));
AOI21X1 g60428(.A0 (_2106_), .A1 (WX839), .B0 (n_883), .Y (n_2552));
AOI21X1 g60431(.A0 (_2091_), .A1 (WX869), .B0 (n_877), .Y (n_2551));
AOI21X1 g60440(.A0 (_2104_), .A1 (WX843), .B0 (n_885), .Y (n_2548));
AOI21X1 g60449(.A0 (_2098_), .A1 (WX855), .B0 (n_875), .Y (n_2547));
AOI21X1 g60451(.A0 (_2108_), .A1 (WX899), .B0 (n_882), .Y (n_2546));
AOI21X1 g60452(.A0 (_2078_), .A1 (WX895), .B0 (n_1272), .Y (n_2545));
AOI21X1 g60453(.A0 (_2108_), .A1 (WX891), .B0 (n_887), .Y (n_2544));
AOI21X1 g60455(.A0 (_2083_), .A1 (WX885), .B0 (n_901), .Y (n_2543));
AOI21X1 g60456(.A0 (_2084_), .A1 (WX883), .B0 (n_852), .Y (n_2542));
AOI21X1 g60457(.A0 (_2085_), .A1 (WX881), .B0 (n_846), .Y (n_2541));
AOI21X1 g60458(.A0 (_2108_), .A1 (WX877), .B0 (n_898), .Y (n_2540));
AOI21X1 g60459(.A0 (_2088_), .A1 (WX875), .B0 (n_892), .Y (n_2539));
AOI21X1 g60460(.A0 (_2090_), .A1 (WX871), .B0 (n_894), .Y (n_2538));
AOI21X1 g60461(.A0 (_2108_), .A1 (WX867), .B0 (n_878), .Y (n_2537));
AOI21X1 g60462(.A0 (_2093_), .A1 (WX865), .B0 (n_890), .Y (n_2536));
AOI21X1 g60463(.A0 (_2097_), .A1 (WX857), .B0 (n_893), .Y (n_2535));
AND2X1 g61580(.A (WX5941), .B (n_2378), .Y (n_2534));
AOI21X1 g60464(.A0 (_2101_), .A1 (WX849), .B0 (n_873), .Y (n_2533));
AOI21X1 g60465(.A0 (_2103_), .A1 (WX845), .B0 (n_886), .Y (n_2532));
AOI21X1 g60466(.A0 (_2105_), .A1 (WX841), .B0 (n_889), .Y (n_2531));
AND2X1 g61570(.A (WX3339), .B (n_2529), .Y (n_2530));
AND2X1 g61566(.A (WX11081), .B (n_2527), .Y (n_2528));
CLKBUFX3 g63079(.A (n_6624), .Y (n_2840));
AND2X1 g62582(.A (WX5829), .B (n_2378), .Y (n_2525));
AOI21X1 g60623(.A0 (_2079_), .A1 (WX893), .B0 (n_881), .Y (n_2524));
AOI21X1 g60635(.A0 (_2077_), .A1 (WX897), .B0 (n_896), .Y (n_2523));
AOI21X1 g60649(.A0 (_2102_), .A1 (WX847), .B0 (n_888), .Y (n_2522));
AOI21X1 g60650(.A0 (_2099_), .A1 (WX853), .B0 (n_879), .Y (n_2521));
AOI21X1 g60657(.A0 (_2095_), .A1 (WX861), .B0 (n_874), .Y (n_2520));
AOI21X1 g60658(.A0 (_2082_), .A1 (WX887), .B0 (n_884), .Y (n_2519));
AOI21X1 g60662(.A0 (_2094_), .A1 (WX863), .B0 (n_876), .Y (n_2518));
AOI21X1 g60672(.A0 (_2081_), .A1 (WX889), .B0 (n_891), .Y (n_2517));
AOI21X1 g60673(.A0 (_2089_), .A1 (WX873), .B0 (n_899), .Y (n_2516));
AND2X1 g62596(.A (WX5823), .B (n_2527), .Y (n_2515));
NAND2X1 g60710(.A (n_1005), .B (n_1003), .Y (n_2514));
AND2X1 g61558(.A (WX11169), .B (n_2227), .Y (n_2513));
INVX1 g60724(.A (n_2511), .Y (n_2512));
NAND2X1 g60731(.A (n_1002), .B (n_999), .Y (n_2508));
NAND2X1 g60743(.A (n_998), .B (n_908), .Y (n_2505));
AND2X1 g61552(.A (WX9806), .B (n_2383), .Y (n_2504));
NAND2X1 g60764(.A (n_988), .B (n_910), .Y (n_2503));
NAND2X1 g60785(.A (n_986), .B (n_984), .Y (n_2500));
INVX1 g60795(.A (n_2498), .Y (n_2499));
NAND2X1 g60802(.A (n_982), .B (n_980), .Y (n_2497));
XOR2X1 g60804(.A (n_1315), .B (n_2800), .Y (n_2496));
INVX1 g60807(.A (n_2494), .Y (n_2495));
NAND2X1 g60818(.A (n_923), .B (n_941), .Y (n_2493));
NAND2X1 g60830(.A (n_976), .B (n_955), .Y (n_2488));
NAND2X1 g60842(.A (n_6696), .B (n_6697), .Y (n_2487));
NAND2X1 g60863(.A (n_969), .B (n_971), .Y (n_2484));
NAND2X1 g60872(.A (n_949), .B (n_904), .Y (n_2481));
NAND2X1 g60889(.A (n_952), .B (n_950), .Y (n_2480));
NAND2X1 g60896(.A (n_974), .B (n_967), .Y (n_2477));
AND2X1 g61532(.A (WX2004), .B (n_2216), .Y (n_2476));
AND2X1 g61531(.A (WX9714), .B (n_2383), .Y (n_2475));
INVX1 g60902(.A (n_2472), .Y (n_2473));
NAND2X1 g60906(.A (n_903), .B (n_928), .Y (n_2471));
NAND2X1 g60933(.A (n_957), .B (n_915), .Y (n_2470));
INVX1 g60950(.A (n_2468), .Y (n_2469));
INVX1 g60964(.A (n_2466), .Y (n_2467));
NAND2X1 g60968(.A (n_945), .B (n_942), .Y (n_2465));
NAND2X1 g60991(.A (n_939), .B (n_937), .Y (n_2462));
INVX1 g61010(.A (n_2458), .Y (n_2459));
NAND2X1 g61020(.A (n_6698), .B (n_6699), .Y (n_2457));
INVX1 g61057(.A (n_2453), .Y (n_2454));
AND2X1 g55856(.A (WX10831), .B (n_2346), .Y (n_2452));
NAND2X1 g61069(.A (n_933), .B (n_931), .Y (n_2448));
INVX1 g61083(.A (n_2446), .Y (n_2447));
NAND2X1 g61086(.A (n_991), .B (n_926), .Y (n_2445));
INVX1 g61091(.A (n_2443), .Y (n_2444));
AND2X1 g62569(.A (WX8475), .B (n_2188), .Y (n_2442));
AND2X1 g62572(.A (WX11005), .B (n_2339), .Y (n_2441));
NAND2X1 g61138(.A (n_925), .B (n_922), .Y (n_2440));
NAND2X1 g61140(.A (n_921), .B (n_919), .Y (n_2439));
INVX1 g61151(.A (n_2437), .Y (n_2438));
NAND2X1 g61167(.A (n_963), .B (n_960), .Y (n_2434));
AND2X1 g62573(.A (WX3275), .B (n_2227), .Y (n_2433));
NAND2X1 g61179(.A (n_930), .B (n_916), .Y (n_2431));
NAND2X1 g61185(.A (n_918), .B (n_965), .Y (n_2428));
NAND2X1 g61196(.A (n_1007), .B (n_947), .Y (n_2425));
NAND2X1 g61209(.A (n_914), .B (n_912), .Y (n_2424));
INVX1 g61219(.A (n_2422), .Y (n_2423));
NAND2X1 g61229(.A (n_954), .B (n_909), .Y (n_2421));
AND2X1 g62571(.A (WX5901), .B (n_2298), .Y (n_2420));
NAND2X1 g61233(.A (n_993), .B (n_911), .Y (n_2419));
NAND2X1 g61271(.A (n_959), .B (n_907), .Y (n_2412));
NAND2X1 g61295(.A (n_906), .B (n_902), .Y (n_2409));
AND2X1 g62567(.A (WX2036), .B (n_2188), .Y (n_2408));
NAND2X1 g61307(.A (n_996), .B (n_994), .Y (n_2406));
AND2X1 g55860(.A (WX1780), .B (n_2402), .Y (n_2405));
AND2X1 g61521(.A (WX11059), .B (n_2346), .Y (n_2404));
AND2X1 g61523(.A (WX3271), .B (n_2402), .Y (n_2403));
AND2X1 g61524(.A (WX11033), .B (n_2400), .Y (n_2401));
AND2X1 g61526(.A (WX7252), .B (n_2227), .Y (n_2399));
AND2X1 g61527(.A (WX3257), .B (n_2378), .Y (n_2398));
AND2X1 g61528(.A (WX3403), .B (n_2396), .Y (n_2397));
AND2X1 g61529(.A (WX11115), .B (n_2400), .Y (n_2395));
AND2X1 g61530(.A (WX11049), .B (n_2227), .Y (n_2394));
AND2X1 g61533(.A (WX11037), .B (n_2402), .Y (n_2393));
AND2X1 g61535(.A (WX9852), .B (n_2402), .Y (n_2392));
AND2X1 g61537(.A (WX9702), .B (n_2371), .Y (n_2391));
AND2X1 g61539(.A (WX9876), .B (n_2388), .Y (n_2390));
AND2X1 g61540(.A (WX11121), .B (n_2388), .Y (n_2389));
AND2X1 g61541(.A (WX7114), .B (n_2346), .Y (n_2387));
AND2X1 g61546(.A (WX9802), .B (n_2346), .Y (n_2386));
AND2X1 g61550(.A (WX9824), .B (n_2383), .Y (n_2385));
AND2X1 g61551(.A (WX7220), .B (n_2383), .Y (n_2384));
AND2X1 g61554(.A (WX11073), .B (n_2383), .Y (n_2382));
AND2X1 g61555(.A (WX9878), .B (n_2383), .Y (n_2380));
AND2X1 g61556(.A (WX11111), .B (n_2378), .Y (n_2379));
AND2X1 g61561(.A (WX9850), .B (n_2227), .Y (n_2377));
AND2X1 g61562(.A (WX11079), .B (n_2227), .Y (n_2376));
AND2X1 g61563(.A (WX7110), .B (n_2227), .Y (n_2375));
AND2X1 g61564(.A (WX7240), .B (n_2527), .Y (n_2373));
AND2X1 g61568(.A (WX11083), .B (n_2371), .Y (n_2372));
AND2X1 g61571(.A (WX8491), .B (n_2371), .Y (n_2370));
AND2X1 g62556(.A (WX8473), .B (n_2216), .Y (n_2369));
AND2X1 g61578(.A (WX2068), .B (n_2378), .Y (n_2368));
AND2X1 g61581(.A (WX11093), .B (n_2378), .Y (n_2366));
AND2X1 g61582(.A (WX5919), .B (n_2188), .Y (n_2365));
AND2X1 g61583(.A (WX7160), .B (n_2346), .Y (n_2364));
AND2X1 g62560(.A (WX3421), .B (n_2402), .Y (n_2363));
AND2X1 g61586(.A (WX3349), .B (n_2378), .Y (n_2362));
AND2X1 g61589(.A (WX11153), .B (n_2383), .Y (n_2361));
AND2X1 g61591(.A (WX7182), .B (n_2383), .Y (n_2360));
AND2X1 g61594(.A (WX11103), .B (n_2400), .Y (n_2359));
AND2X1 g61595(.A (WX5925), .B (n_2527), .Y (n_2358));
AND2X1 g61596(.A (WX7196), .B (n_2402), .Y (n_2357));
AND2X1 g61597(.A (WX7204), .B (n_2402), .Y (n_2356));
AND2X1 g61598(.A (WX3279), .B (n_2378), .Y (n_2355));
AND2X1 g61599(.A (WX5953), .B (n_2378), .Y (n_2353));
AND2X1 g61600(.A (WX3285), .B (n_2378), .Y (n_2352));
AND2X1 g61601(.A (WX4594), .B (n_2227), .Y (n_2351));
AND2X1 g61606(.A (WX7164), .B (n_2400), .Y (n_2350));
AND2X1 g61610(.A (WX7294), .B (n_2227), .Y (n_2349));
AND2X1 g61611(.A (WX11113), .B (n_2378), .Y (n_2348));
AND2X1 g61613(.A (WX7234), .B (n_2346), .Y (n_2347));
AND2X1 g61615(.A (WX9712), .B (n_2378), .Y (n_2345));
AND2X1 g61616(.A (WX5929), .B (n_2346), .Y (n_2344));
AND2X1 g61617(.A (WX7244), .B (n_2346), .Y (n_2343));
AND2X1 g61618(.A (WX7248), .B (n_2223), .Y (n_2341));
AND2X1 g61619(.A (WX9882), .B (n_2339), .Y (n_2340));
AND2X1 g61620(.A (WX4550), .B (n_2378), .Y (n_2338));
AND2X1 g61623(.A (WX7232), .B (n_2378), .Y (n_2337));
AND2X1 g61625(.A (WX2064), .B (n_2378), .Y (n_2336));
AND2X1 g61626(.A (WX5927), .B (n_2333), .Y (n_2335));
AND2X1 g61627(.A (WX9822), .B (n_2333), .Y (n_2334));
AND2X1 g61629(.A (WX7276), .B (n_2325), .Y (n_2332));
AND2X1 g61630(.A (WX3277), .B (n_2272), .Y (n_2331));
AND2X1 g62555(.A (WX5851), .B (n_2378), .Y (n_2330));
AND2X1 g61632(.A (WX11177), .B (n_2527), .Y (n_2329));
AND2X1 g61634(.A (WX11133), .B (n_2378), .Y (n_2328));
AND2X1 g61639(.A (WX11137), .B (n_2325), .Y (n_2326));
AND2X1 g61641(.A (WX11161), .B (n_2378), .Y (n_2324));
AND2X1 g61642(.A (WX5933), .B (n_2388), .Y (n_2323));
AND2X1 g61644(.A (WX3379), .B (n_2378), .Y (n_2322));
AND2X1 g61649(.A (WX9750), .B (n_2311), .Y (n_2321));
AND2X1 g61653(.A (WX7230), .B (n_2383), .Y (n_2320));
AND2X1 g61654(.A (WX3237), .B (n_2188), .Y (n_2318));
AND2X1 g61656(.A (WX5939), .B (n_2188), .Y (n_2317));
AND2X1 g61658(.A (WX9716), .B (n_2188), .Y (n_2316));
AND2X1 g61661(.A (WX5871), .B (n_2188), .Y (n_2315));
AND2X1 g61664(.A (WX9744), .B (n_2188), .Y (n_2313));
AND2X1 g61666(.A (WX9762), .B (n_2311), .Y (n_2312));
AND2X1 g61667(.A (WX4558), .B (n_2311), .Y (n_2310));
AND2X1 g61668(.A (WX3273), .B (n_2188), .Y (n_2309));
AND2X1 g61670(.A (WX5945), .B (n_2311), .Y (n_2308));
AND2X1 g61671(.A (WX9860), .B (n_2311), .Y (n_2307));
AND2X1 g61672(.A (WX7228), .B (n_2383), .Y (n_2306));
AND2X1 g61673(.A (WX7226), .B (n_2383), .Y (n_2305));
AND2X1 g61680(.A (WX11109), .B (n_2311), .Y (n_2304));
AND2X1 g61681(.A (WX8423), .B (n_2311), .Y (n_2303));
AND2X1 g61682(.A (WX3327), .B (n_2311), .Y (n_2302));
AND2X1 g62551(.A (WX2042), .B (n_2388), .Y (n_2301));
AND2X1 g61686(.A (WX7222), .B (n_2383), .Y (n_2300));
AND2X1 g61687(.A (WX9856), .B (n_2298), .Y (n_2299));
AND2X1 g61689(.A (WX7118), .B (n_2383), .Y (n_2297));
AND2X1 g61690(.A (WX7218), .B (n_2346), .Y (n_2296));
AND2X1 g61691(.A (WX7224), .B (n_2346), .Y (n_2295));
AND2X1 g61693(.A (WX4544), .B (n_2188), .Y (n_2293));
AND2X1 g61694(.A (WX4560), .B (n_2378), .Y (n_2292));
AND2X1 g62549(.A (WX5819), .B (n_2346), .Y (n_2291));
AND2X1 g61697(.A (WX7214), .B (n_2378), .Y (n_2290));
AND2X1 g61698(.A (WX3319), .B (n_2246), .Y (n_2289));
AND2X1 g61700(.A (WX4598), .B (n_2188), .Y (n_2288));
AND2X1 g61701(.A (WX9820), .B (n_2188), .Y (n_2287));
AND2X1 g61702(.A (WX5979), .B (n_2346), .Y (n_2286));
AND2X1 g61703(.A (WX11107), .B (n_2346), .Y (n_2285));
AND2X1 g61704(.A (WX9698), .B (n_2346), .Y (n_2284));
AND2X1 g61706(.A (WX3365), .B (n_2311), .Y (n_2283));
AND2X1 g61707(.A (WX11131), .B (n_2325), .Y (n_2282));
AND2X1 g61708(.A (WX3361), .B (n_2298), .Y (n_2281));
AND2X1 g61711(.A (WX11163), .B (n_2227), .Y (n_2280));
AND2X1 g61712(.A (WX8517), .B (n_2227), .Y (n_2279));
AND2X1 g61714(.A (WX9772), .B (n_2346), .Y (n_2277));
AND2X1 g61717(.A (WX11123), .B (n_2346), .Y (n_2276));
AND2X1 g61719(.A (WX3351), .B (n_2227), .Y (n_2275));
AND2X1 g61720(.A (WX4562), .B (n_2227), .Y (n_2274));
AND2X1 g61721(.A (WX4540), .B (n_2272), .Y (n_2273));
AND2X1 g61724(.A (WX5879), .B (n_2333), .Y (n_2271));
AND2X1 g61725(.A (WX5875), .B (n_2333), .Y (n_2270));
AND2X1 g61728(.A (WX5991), .B (n_2227), .Y (n_2269));
AND2X1 g61729(.A (WX2056), .B (n_2227), .Y (n_2268));
AND2X1 g61731(.A (WX3263), .B (n_2227), .Y (n_2267));
AND2X1 g61732(.A (WX7166), .B (n_2378), .Y (n_2266));
AND2X1 g61733(.A (WX7190), .B (n_2346), .Y (n_2264));
AND2X1 g62544(.A (WX3381), .B (n_2378), .Y (n_2262));
AND2X1 g61739(.A (WX9774), .B (n_2346), .Y (n_2261));
AND2X1 g61741(.A (WX7256), .B (n_2272), .Y (n_2260));
AND2X1 g62542(.A (WX2084), .B (n_2346), .Y (n_2259));
AND2X1 g61743(.A (WX5985), .B (n_2272), .Y (n_2258));
AND2X1 g61744(.A (WX7192), .B (n_2246), .Y (n_2257));
AND2X1 g61745(.A (WX7194), .B (n_2346), .Y (n_2256));
AND2X1 g61746(.A (WX8445), .B (n_2346), .Y (n_2255));
AND2X1 g61747(.A (WX5999), .B (n_2333), .Y (n_2254));
AND2X1 g61749(.A (WX9726), .B (n_2251), .Y (n_2253));
AND2X1 g61750(.A (WX9704), .B (n_2251), .Y (n_2252));
AND2X1 g61751(.A (WX7186), .B (n_2272), .Y (n_2250));
AND2X1 g61752(.A (WX8441), .B (n_2272), .Y (n_2249));
AND2X1 g61753(.A (WX5923), .B (n_2333), .Y (n_2248));
AND2X1 g61754(.A (WX2128), .B (n_2246), .Y (n_2247));
AND2X1 g61755(.A (WX2126), .B (n_2246), .Y (n_2245));
AND2X1 g61759(.A (WX7278), .B (n_2333), .Y (n_2244));
AND2X1 g61761(.A (WX5997), .B (n_2396), .Y (n_2243));
AND2X1 g61762(.A (WX3363), .B (n_2396), .Y (n_2242));
AND2X1 g61765(.A (WX3259), .B (n_2346), .Y (n_2241));
AND2X1 g61768(.A (WX11099), .B (n_2383), .Y (n_2240));
AND2X1 g61769(.A (WX2088), .B (n_2383), .Y (n_2239));
AND2X1 g61770(.A (WX9800), .B (n_2188), .Y (n_2238));
AND2X1 g61772(.A (WX7280), .B (n_2383), .Y (n_2237));
AND2X1 g61773(.A (WX8519), .B (n_2188), .Y (n_2236));
AND2X1 g62539(.A (WX5831), .B (n_2188), .Y (n_2235));
AND2X1 g61777(.A (WX3289), .B (n_2188), .Y (n_2234));
AND2X1 g61778(.A (WX4638), .B (n_2378), .Y (n_2233));
AND2X1 g61781(.A (WX2112), .B (n_2346), .Y (n_2232));
AND2X1 g61783(.A (WX9730), .B (n_2346), .Y (n_2231));
AND2X1 g61784(.A (WX9754), .B (n_2188), .Y (n_2230));
AND2X1 g61790(.A (WX3415), .B (n_2378), .Y (n_2229));
AND2X1 g61791(.A (WX3255), .B (n_2227), .Y (n_2228));
AND2X1 g58615(.A (WX2066), .B (n_2346), .Y (n_2226));
AND2X1 g61794(.A (WX2122), .B (n_2227), .Y (n_2225));
AND2X1 g61795(.A (WX8529), .B (n_2223), .Y (n_2224));
AND2X1 g61796(.A (WX9832), .B (n_2378), .Y (n_2222));
AND2X1 g61797(.A (WX8449), .B (n_2223), .Y (n_2221));
AND2X1 g61799(.A (WX7158), .B (n_2218), .Y (n_2220));
AND2X1 g61800(.A (WX11011), .B (n_2218), .Y (n_2219));
AND2X1 g61802(.A (WX4676), .B (n_2216), .Y (n_2217));
AND2X1 g61803(.A (WX7156), .B (n_2216), .Y (n_2215));
AND2X1 g61805(.A (WX7154), .B (n_2223), .Y (n_2214));
AND2X1 g61807(.A (WX9816), .B (n_2383), .Y (n_2213));
AND2X1 g61809(.A (WX7134), .B (n_2223), .Y (n_2212));
AND2X1 g61810(.A (WX7246), .B (n_2246), .Y (n_2211));
AND2X1 g61811(.A (WX7144), .B (n_2371), .Y (n_2210));
AND2X1 g61812(.A (WX9736), .B (n_2246), .Y (n_2209));
AND2X1 g61816(.A (WX7150), .B (n_2371), .Y (n_2208));
AND2X1 g61820(.A (WX9842), .B (n_2371), .Y (n_2207));
AND2X1 g61823(.A (WX7148), .B (n_2371), .Y (n_2206));
AND2X1 g61825(.A (WX3321), .B (n_2383), .Y (n_2205));
AND2X1 g61826(.A (WX4634), .B (n_2396), .Y (n_2204));
AND2X1 g61827(.A (WX11087), .B (n_2198), .Y (n_2203));
AND2X1 g61828(.A (WX7124), .B (n_2227), .Y (n_2202));
AND2X1 g61829(.A (WX3301), .B (n_2218), .Y (n_2201));
AND2X1 g61832(.A (WX3409), .B (n_2371), .Y (n_2200));
AND2X1 g61834(.A (WX9778), .B (n_2198), .Y (n_2199));
AND2X1 g61835(.A (WX7272), .B (n_2218), .Y (n_2197));
AND2X1 g61837(.A (WX7138), .B (n_2216), .Y (n_2196));
AND2X1 g61838(.A (WX2118), .B (n_2218), .Y (n_2194));
AND2X1 g61839(.A (WX4626), .B (n_2529), .Y (n_2193));
AND2X1 g61840(.A (WX5949), .B (n_2383), .Y (n_2192));
AND2X1 g61847(.A (WX3265), .B (n_2529), .Y (n_2191));
AND2X1 g61848(.A (WX11141), .B (n_2383), .Y (n_2190));
AND2X1 g61849(.A (WX5947), .B (n_2188), .Y (n_2189));
AND2X1 g62536(.A (WX11025), .B (n_2227), .Y (n_2187));
AND2X1 g61850(.A (WX2114), .B (n_2188), .Y (n_2186));
AND2X1 g61851(.A (WX4584), .B (n_2227), .Y (n_2185));
AND2X1 g61854(.A (WX3267), .B (n_2227), .Y (n_2183));
AND2X1 g61855(.A (WX7120), .B (n_2383), .Y (n_2182));
AND2X1 g61856(.A (WX7132), .B (n_2227), .Y (n_2181));
AND2X1 g61858(.A (WX3357), .B (n_2227), .Y (n_2180));
AND2X1 g61859(.A (WX3281), .B (n_2227), .Y (n_2179));
AND2X1 g61861(.A (WX3247), .B (n_2188), .Y (n_2178));
AND2X1 g61863(.A (WX11119), .B (n_2198), .Y (n_2177));
AND2X1 g61864(.A (WX7126), .B (n_2198), .Y (n_2176));
AND2X1 g61865(.A (WX5937), .B (n_2216), .Y (n_2175));
AND2X1 g61866(.A (WX7128), .B (n_2227), .Y (n_2174));
AND2X1 g61867(.A (WX3347), .B (n_2339), .Y (n_2173));
AND2X1 g61868(.A (WX2060), .B (n_2251), .Y (n_2172));
AND2X1 g61869(.A (WX7130), .B (n_2251), .Y (n_2171));
AND2X1 g61870(.A (WX9742), .B (n_2396), .Y (n_2170));
AND2X1 g61871(.A (WX11085), .B (n_2383), .Y (n_2169));
AND2X1 g61873(.A (WX11043), .B (n_2251), .Y (n_2168));
AND2X1 g61874(.A (WX3283), .B (n_2378), .Y (n_2167));
AND2X1 g61877(.A (WX8447), .B (n_2198), .Y (n_2166));
AND2X1 g61879(.A (WX4564), .B (n_2227), .Y (n_2165));
AND2X1 g61881(.A (WX11067), .B (n_2198), .Y (n_2164));
AND2X1 g61883(.A (WX8453), .B (n_2216), .Y (n_2163));
AND2X1 g61884(.A (WX4538), .B (n_2216), .Y (n_2162));
AND2X1 g61886(.A (WX5959), .B (n_2529), .Y (n_2161));
AND2X1 g61887(.A (WX3355), .B (n_2298), .Y (n_2160));
AND2X1 g61890(.A (WX4588), .B (n_2227), .Y (n_2159));
AND2X1 g61891(.A (WX9724), .B (n_2227), .Y (n_2158));
AND2X1 g61892(.A (WX5965), .B (n_2223), .Y (n_2157));
AND2X1 g61893(.A (WX11147), .B (n_2383), .Y (n_2156));
AND2X1 g61894(.A (WX7122), .B (n_2216), .Y (n_2155));
AND2X1 g61900(.A (WX4636), .B (n_2216), .Y (n_2154));
AND2X1 g61901(.A (WX4628), .B (n_2333), .Y (n_2153));
AND2X1 g61902(.A (WX8551), .B (n_2298), .Y (n_2152));
AND2X1 g61904(.A (WX9872), .B (n_2223), .Y (n_2151));
AND2X1 g61905(.A (WX5861), .B (n_2227), .Y (n_2150));
AND2X1 g61906(.A (WX8407), .B (n_2246), .Y (n_2149));
AND2X1 g61907(.A (WX8547), .B (n_2198), .Y (n_2148));
AND2X1 g61915(.A (WX4570), .B (n_2227), .Y (n_2147));
AND2X1 g61917(.A (WX11027), .B (n_2383), .Y (n_2146));
AND2X1 g61919(.A (WX11139), .B (n_2251), .Y (n_2145));
AND2X1 g61920(.A (WX5683), .B (n_2198), .Y (n_2144));
AND2X1 g61921(.A (WX4652), .B (n_2246), .Y (n_2143));
AND2X1 g61925(.A (WX5957), .B (n_2251), .Y (n_2142));
AND2X1 g61926(.A (WX3287), .B (n_2346), .Y (n_2141));
AND2X1 g61929(.A (WX11149), .B (n_2383), .Y (n_2140));
AND2X1 g61931(.A (WX8557), .B (n_2227), .Y (n_2139));
AND2X1 g61932(.A (WX9722), .B (n_2218), .Y (n_2138));
AND2X1 g61933(.A (WX9840), .B (n_2396), .Y (n_2137));
AND2X1 g62534(.A (WX5867), .B (n_2383), .Y (n_2136));
AND2X1 g61935(.A (WX2076), .B (n_2371), .Y (n_2135));
AND2X1 g61936(.A (WX7116), .B (n_2378), .Y (n_2134));
AND2X1 g61937(.A (WX9796), .B (n_2298), .Y (n_2133));
AND2X1 g61938(.A (WX9776), .B (n_2246), .Y (n_2132));
AND2X1 g61939(.A (WX11071), .B (n_2383), .Y (n_2130));
AND2X1 g61943(.A (WX9760), .B (n_2216), .Y (n_2129));
AND2X1 g61944(.A (WX4576), .B (n_2346), .Y (n_2128));
AND2X1 g61947(.A (WX3395), .B (n_2346), .Y (n_2127));
AND2X1 g61948(.A (WX4526), .B (n_2216), .Y (n_2126));
AND2X1 g61949(.A (WX9790), .B (n_2383), .Y (n_2125));
AND2X1 g61950(.A (WX9768), .B (n_2216), .Y (n_2124));
AND2X1 g61952(.A (WX4662), .B (n_2216), .Y (n_2123));
AND2X1 g61953(.A (WX4580), .B (n_2216), .Y (n_2122));
AND2X1 g61955(.A (WX9728), .B (n_2188), .Y (n_2121));
AND2X1 g61956(.A (WX9718), .B (n_2383), .Y (n_2120));
AND2X1 g61957(.A (WX3405), .B (n_2346), .Y (n_2119));
AND2X1 g61958(.A (WX3245), .B (n_2227), .Y (n_2118));
AND2X1 g61959(.A (WX2010), .B (n_2333), .Y (n_2117));
AND2X1 g61961(.A (WX8589), .B (n_2325), .Y (n_2116));
AND2X1 g61962(.A (WX4688), .B (n_2246), .Y (n_2115));
AND2X1 g61963(.A (WX9706), .B (n_2527), .Y (n_2114));
AND2X1 g61965(.A (WX3243), .B (n_2298), .Y (n_2113));
AND2X1 g61966(.A (WX3241), .B (n_2383), .Y (n_2112));
AND2X1 g61967(.A (WX4698), .B (n_2346), .Y (n_2111));
AND2X1 g61968(.A (WX8591), .B (n_2339), .Y (n_2110));
AND2X1 g61969(.A (WX3239), .B (n_2402), .Y (n_2109));
AND2X1 g61970(.A (WX4704), .B (n_2223), .Y (n_2108));
AND2X1 g61971(.A (WX8583), .B (n_2383), .Y (n_2107));
AND2X1 g61972(.A (WX11029), .B (n_2396), .Y (n_2106));
AND2X1 g61973(.A (WX4712), .B (n_2246), .Y (n_2105));
AND2X1 g61976(.A (WX8565), .B (n_2383), .Y (n_2104));
AND2X1 g61978(.A (WX8579), .B (n_2339), .Y (n_2103));
AND2X1 g61980(.A (WX3383), .B (n_2378), .Y (n_2102));
AND2X1 g61981(.A (WX8559), .B (n_2396), .Y (n_2101));
AND2X1 g61982(.A (WX2104), .B (n_2311), .Y (n_2100));
AND2X1 g61983(.A (WX4678), .B (n_2346), .Y (n_2099));
AND2X1 g61985(.A (WX3233), .B (n_2339), .Y (n_2098));
AND2X1 g61986(.A (WX3393), .B (n_2378), .Y (n_2097));
AND2X1 g61987(.A (WX8455), .B (n_2188), .Y (n_2096));
AND2X1 g61988(.A (WX3235), .B (n_2378), .Y (n_2095));
AND2X1 g61990(.A (WX8567), .B (n_2227), .Y (n_2094));
AND2X1 g61992(.A (WX8573), .B (n_2227), .Y (n_2093));
AND2X1 g61994(.A (WX3391), .B (n_2227), .Y (n_2092));
AND2X1 g61995(.A (WX10995), .B (n_2227), .Y (n_2091));
AND2X1 g61996(.A (WX8571), .B (n_2227), .Y (n_2090));
AND2X1 g61997(.A (WX2108), .B (n_2227), .Y (n_2089));
AND2X1 g61998(.A (WX2008), .B (n_2396), .Y (n_2087));
AND2X1 g62000(.A (WX7242), .B (n_2227), .Y (n_2086));
AND2X1 g62001(.A (WX11015), .B (n_2346), .Y (n_2085));
AND2X1 g62002(.A (WX9864), .B (n_2346), .Y (n_2084));
AND2X1 g62003(.A (WX3385), .B (n_2339), .Y (n_2083));
AND2X1 g62004(.A (WX4710), .B (n_2339), .Y (n_2082));
AND2X1 g62009(.A (WX2012), .B (n_2378), .Y (n_2081));
AND2X1 g62010(.A (WX2086), .B (n_2346), .Y (n_2080));
AND2X1 g62011(.A (WX4680), .B (n_2251), .Y (n_2079));
AND2X1 g62012(.A (WX4696), .B (n_2383), .Y (n_2078));
AND2X1 g62013(.A (WX8561), .B (n_2400), .Y (n_2077));
AND2X1 g62014(.A (WX11077), .B (n_2227), .Y (n_2076));
AND2X1 g62015(.A (WX2106), .B (n_2227), .Y (n_2075));
AND2X1 g62016(.A (WX4686), .B (n_2396), .Y (n_2074));
AND2X1 g62017(.A (WX3335), .B (n_2388), .Y (n_2073));
AND2X1 g62018(.A (WX4666), .B (n_2383), .Y (n_2072));
AND2X1 g62019(.A (WX9830), .B (n_2272), .Y (n_2071));
AND2X1 g62020(.A (WX9788), .B (n_2529), .Y (n_2070));
AND2X1 g62021(.A (WX4674), .B (n_2388), .Y (n_2069));
AND2X1 g62022(.A (WX9838), .B (n_2396), .Y (n_2068));
AND2X1 g62023(.A (WX4670), .B (n_2227), .Y (n_2067));
AND2X1 g62024(.A (WX3253), .B (n_2529), .Y (n_2066));
AND2X1 g62025(.A (WX4664), .B (n_2227), .Y (n_2065));
AND2X1 g62026(.A (WX7296), .B (n_2216), .Y (n_2064));
AND2X1 g62027(.A (WX4660), .B (n_2383), .Y (n_2063));
AND2X1 g62030(.A (WX9696), .B (n_2529), .Y (n_2062));
AND2X1 g62033(.A (WX4566), .B (n_2529), .Y (n_2061));
AND2X1 g62034(.A (WX11001), .B (n_2227), .Y (n_2060));
AND2X1 g62036(.A (WX9812), .B (n_2227), .Y (n_2059));
AND2X1 g62038(.A (WX4620), .B (n_2383), .Y (n_2058));
AND2X1 g62041(.A (WX3407), .B (n_2227), .Y (n_2057));
AND2X1 g62043(.A (WX8531), .B (n_2383), .Y (n_2056));
AND2X1 g62044(.A (WX2102), .B (n_2383), .Y (n_2055));
AND2X1 g62047(.A (WX8555), .B (n_2346), .Y (n_2054));
AND2X1 g62048(.A (WX3295), .B (n_2346), .Y (n_2053));
AND2X1 g62050(.A (WX2100), .B (n_2227), .Y (n_2052));
AND2X1 g62052(.A (WX11017), .B (n_2346), .Y (n_2051));
AND2X1 g62055(.A (WX5951), .B (n_2378), .Y (n_2050));
AND2X1 g62057(.A (WX2098), .B (n_2396), .Y (n_2049));
AND2X1 g62058(.A (WX3297), .B (n_2188), .Y (n_2048));
AND2X1 g62059(.A (WX5849), .B (n_2198), .Y (n_2047));
AND2X1 g62060(.A (WX8553), .B (n_2529), .Y (n_2046));
AND2X1 g62529(.A (WX3401), .B (n_2298), .Y (n_2045));
AND2X1 g62061(.A (WX2016), .B (n_2529), .Y (n_2044));
AND2X1 g62062(.A (WX11063), .B (n_2188), .Y (n_2043));
AND2X1 g62064(.A (WX9700), .B (n_2216), .Y (n_2042));
AND2X1 g62065(.A (WX8463), .B (n_2227), .Y (n_2041));
AND2X1 g62066(.A (WX2096), .B (n_2325), .Y (n_2040));
AND2X1 g62067(.A (WX3331), .B (n_2188), .Y (n_2039));
AND2X1 g62068(.A (WX3299), .B (n_2371), .Y (n_2038));
AND2X1 g62072(.A (WX8549), .B (n_2378), .Y (n_2037));
AND2X1 g62075(.A (WX5859), .B (n_2400), .Y (n_2036));
AND2X1 g62076(.A (WX4548), .B (n_2346), .Y (n_2035));
AND2X1 g62077(.A (WX3419), .B (n_2378), .Y (n_2034));
AND2X1 g62078(.A (WX8545), .B (n_2383), .Y (n_2033));
AND2X1 g62080(.A (WX4622), .B (n_2272), .Y (n_2032));
AND2X1 g62081(.A (WX8539), .B (n_2378), .Y (n_2031));
AND2X1 g62082(.A (WX2094), .B (n_2402), .Y (n_2030));
AND2X1 g62084(.A (WX2048), .B (n_2396), .Y (n_2029));
AND2X1 g62086(.A (WX4600), .B (n_2346), .Y (n_2028));
AND2X1 g62087(.A (WX4602), .B (n_2251), .Y (n_2027));
AND2X1 g62088(.A (WX8405), .B (n_2400), .Y (n_2026));
AND2X1 g62089(.A (WX4650), .B (n_2218), .Y (n_2025));
AND2X1 g62090(.A (WX8543), .B (n_2223), .Y (n_2024));
AND2X1 g62091(.A (WX10997), .B (n_2383), .Y (n_2023));
AND2X1 g62092(.A (WX7282), .B (n_2216), .Y (n_2022));
AND2X1 g62094(.A (WX9884), .B (n_2346), .Y (n_2021));
AND2X1 g62096(.A (WX5899), .B (n_2223), .Y (n_2020));
AND2X1 g62098(.A (WX4616), .B (n_2346), .Y (n_2019));
AND2X1 g62099(.A (WX8457), .B (n_2402), .Y (n_2018));
AND2X1 g62100(.A (WX5855), .B (n_2339), .Y (n_2017));
AND2X1 g62101(.A (WX8435), .B (n_2388), .Y (n_2016));
AND2X1 g62104(.A (WX8537), .B (n_2402), .Y (n_2015));
AND2X1 g62106(.A (WX9854), .B (n_2188), .Y (n_2014));
AND2X1 g62107(.A (WX10999), .B (n_2388), .Y (n_2013));
AND2X1 g62108(.A (WX7250), .B (n_2383), .Y (n_2012));
AND2X1 g62531(.A (WX2006), .B (n_2188), .Y (n_2011));
AND2X1 g62113(.A (WX3387), .B (n_2527), .Y (n_2010));
AND2X1 g62116(.A (WX8535), .B (n_2272), .Y (n_2009));
AND2X1 g62117(.A (WX7212), .B (n_2402), .Y (n_2008));
AND2X1 g62118(.A (WX5981), .B (n_2378), .Y (n_2007));
AND2X1 g62119(.A (WX4586), .B (n_2272), .Y (n_2006));
AND2X1 g62120(.A (WX4656), .B (n_2383), .Y (n_2005));
AND2X1 g62121(.A (WX3333), .B (n_2188), .Y (n_2004));
AND2X1 g62122(.A (WX9826), .B (n_2383), .Y (n_2003));
AND2X1 g62124(.A (WX2092), .B (n_2311), .Y (n_2002));
AND2X1 g62126(.A (WX4624), .B (n_2388), .Y (n_2001));
AND2X1 g62127(.A (WX7136), .B (n_2388), .Y (n_2000));
AND2X1 g62128(.A (WX7268), .B (n_2346), .Y (n_1999));
AND2X1 g62129(.A (WX4642), .B (n_2527), .Y (n_1998));
AND2X1 g62130(.A (WX8409), .B (n_2346), .Y (n_1997));
AND2X1 g62131(.A (WX4618), .B (n_2246), .Y (n_1996));
AND2X1 g62132(.A (WX4612), .B (n_2298), .Y (n_1995));
AND2X1 g62133(.A (WX7292), .B (n_2378), .Y (n_1994));
AND2X1 g62135(.A (WX3231), .B (n_2378), .Y (n_1993));
AND2X1 g62136(.A (WX8489), .B (n_2346), .Y (n_1992));
AND2X1 g62138(.A (WX8525), .B (n_2325), .Y (n_1991));
AND2X1 g62140(.A (WX11159), .B (n_2346), .Y (n_1990));
AND2X1 g62143(.A (WX3367), .B (n_2383), .Y (n_1989));
AND2X1 g62144(.A (WX11061), .B (n_2227), .Y (n_1988));
AND2X1 g62148(.A (WX4392), .B (n_2227), .Y (n_1987));
AND2X1 g62149(.A (WX8569), .B (n_2188), .Y (n_1986));
AND2X1 g62150(.A (WX11125), .B (n_2246), .Y (n_1985));
AND2X1 g62155(.A (WX8413), .B (n_2246), .Y (n_1984));
AND2X1 g62156(.A (WX2062), .B (n_2272), .Y (n_1983));
AND2X1 g62158(.A (WX9758), .B (n_2251), .Y (n_1982));
AND2X1 g62160(.A (WX3397), .B (n_2346), .Y (n_1981));
AND2X1 g62161(.A (WX7300), .B (n_2346), .Y (n_1980));
AND2X1 g62162(.A (WX6003), .B (n_2333), .Y (n_1979));
AND2X1 g62164(.A (WX4646), .B (n_2333), .Y (n_1978));
AND2X1 g62165(.A (WX9880), .B (n_2346), .Y (n_1977));
AND2X1 g62166(.A (WX7258), .B (n_2325), .Y (n_1976));
AND2X1 g62167(.A (WX8593), .B (n_2227), .Y (n_1975));
AND2X1 g62168(.A (WX11057), .B (n_2227), .Y (n_1974));
AND2X1 g62172(.A (WX3371), .B (n_2346), .Y (n_1973));
AND2X1 g62175(.A (WX8411), .B (n_2227), .Y (n_1972));
AND2X1 g62176(.A (WX9836), .B (n_2227), .Y (n_1971));
AND2X1 g62177(.A (WX11055), .B (n_2378), .Y (n_1970));
AND2X1 g62178(.A (WX8467), .B (n_2227), .Y (n_1969));
AND2X1 g62180(.A (WX9870), .B (n_2378), .Y (n_1968));
AND2X1 g62182(.A (WX7264), .B (n_2227), .Y (n_1967));
AND2X1 g62183(.A (WX4604), .B (n_2223), .Y (n_1966));
AND2X1 g62184(.A (WX9804), .B (n_2218), .Y (n_1965));
AND2X1 g62185(.A (WX8429), .B (n_2527), .Y (n_1964));
AND2X1 g62188(.A (WX5877), .B (n_2188), .Y (n_1963));
AND2X1 g62189(.A (WX6001), .B (n_2378), .Y (n_1962));
AND2X1 g62190(.A (WX8521), .B (n_2378), .Y (n_1961));
AND2X1 g62191(.A (WX7270), .B (n_2216), .Y (n_1960));
AND2X1 g62194(.A (WX5989), .B (n_2218), .Y (n_1959));
AND2X1 g62195(.A (WX5993), .B (n_2383), .Y (n_1958));
AND2X1 g62196(.A (WX3303), .B (n_2198), .Y (n_1957));
AND2X1 g62197(.A (WX7142), .B (n_2216), .Y (n_1956));
AND2X1 g62201(.A (WX9756), .B (n_2383), .Y (n_1955));
AND2X1 g62202(.A (WX7260), .B (n_2216), .Y (n_1954));
AND2X1 g62203(.A (WX5903), .B (n_2383), .Y (n_1953));
AND2X1 g62205(.A (WX11065), .B (n_2223), .Y (n_1951));
AND2X1 g62206(.A (WX4534), .B (n_2223), .Y (n_1950));
AND2X1 g62207(.A (WX4546), .B (n_2383), .Y (n_1949));
AND2X1 g62208(.A (WX2074), .B (n_2346), .Y (n_1948));
AND2X1 g62209(.A (WX8483), .B (n_2383), .Y (n_1947));
AND2X1 g62210(.A (WX3307), .B (n_2227), .Y (n_1946));
AND2X1 g62211(.A (WX9866), .B (n_2378), .Y (n_1945));
AND2X1 g62218(.A (WX4582), .B (n_2216), .Y (n_1944));
AND2X1 g62222(.A (WX4640), .B (n_2383), .Y (n_1943));
AND2X1 g62224(.A (WX4596), .B (n_2383), .Y (n_1942));
AND2X1 g62229(.A (WX7298), .B (n_2227), .Y (n_1941));
AND2X1 g62230(.A (WX2078), .B (n_2227), .Y (n_1940));
AND2X1 g62231(.A (WX2038), .B (n_2227), .Y (n_1939));
AND2X1 g62233(.A (WX11003), .B (n_2378), .Y (n_1938));
AND2X1 g62236(.A (WX5881), .B (n_2346), .Y (n_1937));
AND2X1 g62237(.A (WX4644), .B (n_2383), .Y (n_1936));
AND2X1 g62238(.A (WX2120), .B (n_2378), .Y (n_1935));
AND2X1 g62240(.A (WX4654), .B (n_2371), .Y (n_1934));
AND2X1 g62241(.A (WX3353), .B (n_2383), .Y (n_1933));
AND2X1 g62243(.A (WX5983), .B (n_2383), .Y (n_1932));
AND2X1 g62244(.A (WX4572), .B (n_2383), .Y (n_1931));
AND2X1 g62245(.A (WX8427), .B (n_2346), .Y (n_1930));
AND2X1 g62247(.A (WX4684), .B (n_2339), .Y (n_1929));
AND2X1 g62248(.A (WX4694), .B (n_2346), .Y (n_1928));
AND2X1 g62252(.A (WX9886), .B (n_2227), .Y (n_1927));
AND2X1 g62253(.A (WX4552), .B (n_2227), .Y (n_1926));
AND2X1 g62255(.A (WX4606), .B (n_2378), .Y (n_1925));
AND2X1 g62256(.A (WX4536), .B (n_2227), .Y (n_1924));
AND2X1 g62258(.A (WX5975), .B (n_2188), .Y (n_1923));
AND2X1 g62259(.A (WX2110), .B (n_2402), .Y (n_1922));
AND2X1 g62260(.A (WX7274), .B (n_2346), .Y (n_1921));
AND2X1 g62261(.A (WX5977), .B (n_2272), .Y (n_1920));
AND2X1 g62262(.A (WX3417), .B (n_2378), .Y (n_1919));
AND2X1 g62263(.A (WX8507), .B (n_2371), .Y (n_1918));
AND2X1 g62264(.A (WX9720), .B (n_2383), .Y (n_1917));
AND2X1 g62265(.A (WX5971), .B (n_2346), .Y (n_1916));
AND2X1 g62267(.A (WX5967), .B (n_2227), .Y (n_1915));
AND2X1 g62269(.A (WX7146), .B (n_2383), .Y (n_1914));
AND2X1 g62270(.A (WX8541), .B (n_2198), .Y (n_1913));
AND2X1 g62272(.A (WX5969), .B (n_2346), .Y (n_1912));
AND2X1 g62274(.A (WX3373), .B (n_2371), .Y (n_1911));
AND2X1 g62277(.A (WX5963), .B (n_2333), .Y (n_1910));
AND2X1 g62279(.A (WX8513), .B (n_2346), .Y (n_1909));
AND2X1 g62280(.A (WX8509), .B (n_2383), .Y (n_1908));
AND2X1 g62281(.A (WX8433), .B (n_2383), .Y (n_1907));
AND2X1 g62283(.A (WX11047), .B (n_2346), .Y (n_1906));
AND2X1 g62285(.A (WX5961), .B (n_2198), .Y (n_1905));
AND2X1 g62286(.A (WX8511), .B (n_2298), .Y (n_1904));
AND2X1 g62288(.A (WX8431), .B (n_2198), .Y (n_1903));
AND2X1 g62289(.A (WX7286), .B (n_2216), .Y (n_1902));
AND2X1 g62290(.A (WX7288), .B (n_2216), .Y (n_1901));
AND2X1 g62291(.A (WX3101), .B (n_2216), .Y (n_1900));
AND2X1 g62294(.A (WX3343), .B (n_2227), .Y (n_1899));
AND2X1 g62295(.A (WX7112), .B (n_2371), .Y (n_1898));
AND2X1 g62296(.A (WX9766), .B (n_2227), .Y (n_1897));
AND2X1 g62297(.A (WX3315), .B (n_2383), .Y (n_1896));
AND2X1 g62298(.A (WX2070), .B (n_2198), .Y (n_1895));
AND2X1 g62299(.A (WX11091), .B (n_2339), .Y (n_1894));
AND2X1 g62303(.A (WX3377), .B (n_2218), .Y (n_1893));
AND2X1 g62305(.A (WX5943), .B (n_2227), .Y (n_1892));
AND2X1 g62306(.A (WX8479), .B (n_2227), .Y (n_1891));
AND2X1 g62311(.A (WX8439), .B (n_2346), .Y (n_1890));
AND2X1 g62312(.A (WX9738), .B (n_2251), .Y (n_1889));
AND2X1 g62313(.A (WX9858), .B (n_2383), .Y (n_1888));
AND2X1 g62528(.A (WX9834), .B (n_2527), .Y (n_1887));
AND2X1 g62314(.A (WX7216), .B (n_2325), .Y (n_1886));
AND2X1 g62315(.A (WX2022), .B (n_2246), .Y (n_1885));
AND2X1 g62316(.A (WX4702), .B (n_2527), .Y (n_1884));
AND2X1 g62317(.A (WX4524), .B (n_2527), .Y (n_1883));
AND2X1 g62318(.A (WX5853), .B (n_2529), .Y (n_1882));
AND2X1 g62319(.A (WX5889), .B (n_2227), .Y (n_1881));
AND2X1 g62320(.A (WX8477), .B (n_2378), .Y (n_1880));
AND2X1 g62322(.A (WX4608), .B (n_2227), .Y (n_1879));
AND2X1 g62324(.A (WX5915), .B (n_2216), .Y (n_1878));
AND2X1 g62325(.A (WX8495), .B (n_2371), .Y (n_1877));
AND2X1 g62326(.A (WX3313), .B (n_2198), .Y (n_1876));
AND2X1 g62327(.A (WX8437), .B (n_2216), .Y (n_1875));
AND2X1 g62329(.A (WX5935), .B (n_2246), .Y (n_1874));
AND2X1 g62331(.A (WX8501), .B (n_2246), .Y (n_1873));
AND2X1 g62332(.A (WX11009), .B (n_2218), .Y (n_1872));
AND2X1 g62333(.A (WX5931), .B (n_2218), .Y (n_1871));
AND2X1 g62335(.A (WX4590), .B (n_2246), .Y (n_1870));
AND2X1 g62336(.A (WX2124), .B (n_2378), .Y (n_1869));
AND2X1 g62341(.A (WX9792), .B (n_2216), .Y (n_1868));
AND2X1 g62344(.A (WX8499), .B (n_2378), .Y (n_1867));
AND2X1 g62345(.A (WX10991), .B (n_2383), .Y (n_1866));
AND2X1 g62348(.A (WX7162), .B (n_2227), .Y (n_1865));
AND2X1 g62349(.A (WX3411), .B (n_2188), .Y (n_1864));
AND2X1 g62350(.A (WX8497), .B (n_2246), .Y (n_1863));
AND2X1 g62354(.A (WX5917), .B (n_2246), .Y (n_1862));
AND2X1 g62355(.A (WX11157), .B (n_2383), .Y (n_1861));
AND2X1 g62362(.A (WX8493), .B (n_2227), .Y (n_1860));
AND2X1 g62363(.A (WX9828), .B (n_2227), .Y (n_1859));
AND2X1 g62364(.A (WX5911), .B (n_2378), .Y (n_1858));
AND2X1 g62367(.A (WX2040), .B (n_2346), .Y (n_1857));
AND2X1 g62369(.A (WX8487), .B (n_2251), .Y (n_1856));
AND2X1 g62370(.A (WX5913), .B (n_2333), .Y (n_1855));
AND2X1 g62372(.A (WX5905), .B (n_2325), .Y (n_1854));
AND2X1 g62373(.A (WX3345), .B (n_2188), .Y (n_1853));
AND2X1 g62374(.A (WX9748), .B (n_2346), .Y (n_1852));
AND2X1 g62376(.A (WX2058), .B (n_2227), .Y (n_1851));
AND2X1 g62518(.A (WX8461), .B (n_2378), .Y (n_1850));
AND2X1 g62519(.A (WX3329), .B (n_2400), .Y (n_1849));
AND2X1 g62521(.A (WX9734), .B (n_2383), .Y (n_1848));
AND2X1 g62515(.A (WX5883), .B (n_2396), .Y (n_1847));
AND2X1 g62517(.A (WX9868), .B (n_2400), .Y (n_1846));
AND2X1 g62513(.A (WX8417), .B (n_2333), .Y (n_1845));
AND2X1 g62510(.A (WX4714), .B (n_2346), .Y (n_1844));
AND2X1 g62504(.A (WX2090), .B (n_2346), .Y (n_1843));
AND2X1 g62503(.A (WX8421), .B (n_2346), .Y (n_1842));
AND2X1 g62502(.A (WX4554), .B (n_2346), .Y (n_1841));
AND2X1 g62501(.A (WX7168), .B (n_2378), .Y (n_1840));
AND2X1 g62467(.A (WX5907), .B (n_2378), .Y (n_1838));
AND2X1 g62468(.A (WX3249), .B (n_2227), .Y (n_1837));
AND2X1 g62470(.A (WX4630), .B (n_2378), .Y (n_1836));
AND2X1 g62471(.A (WX5895), .B (n_2246), .Y (n_1835));
AND2X1 g62472(.A (WX5887), .B (n_2346), .Y (n_1834));
AND2X1 g62475(.A (WX8403), .B (n_2298), .Y (n_1833));
AND2X1 g62499(.A (WX2024), .B (n_2388), .Y (n_1832));
AND2X1 g62480(.A (WX5897), .B (n_2325), .Y (n_1831));
AND2X1 g62481(.A (WX11173), .B (n_2246), .Y (n_1830));
AND2X1 g62482(.A (WX8425), .B (n_2383), .Y (n_1829));
AND2X1 g62483(.A (WX7170), .B (n_2378), .Y (n_1828));
AND2X1 g62484(.A (WX8465), .B (n_2298), .Y (n_1827));
AND2X1 g62485(.A (WX4530), .B (n_2311), .Y (n_1826));
AND2X1 g62492(.A (WX5891), .B (n_2339), .Y (n_1825));
AND2X1 g62495(.A (WX11097), .B (n_2325), .Y (n_1824));
AND2X1 g62496(.A (WX2116), .B (n_2402), .Y (n_1823));
AND2X1 g62497(.A (WX11151), .B (n_2339), .Y (n_1822));
AND2X1 g62500(.A (WX4706), .B (n_2402), .Y (n_1821));
AND2X1 g62509(.A (WX9784), .B (n_2188), .Y (n_1820));
AND2X1 g62511(.A (WX11013), .B (n_2346), .Y (n_1819));
AND2X1 g62512(.A (WX2052), .B (n_2378), .Y (n_1818));
AND2X1 g62514(.A (WX3341), .B (n_2227), .Y (n_1817));
AND2X1 g62516(.A (WX3323), .B (n_2298), .Y (n_1816));
AND2X1 g62523(.A (WX7176), .B (n_2227), .Y (n_1815));
AND2X1 g62526(.A (WX2018), .B (n_2378), .Y (n_1814));
AND2X1 g62533(.A (WX8503), .B (n_2346), .Y (n_1813));
AND2X1 g62535(.A (WX6005), .B (n_2188), .Y (n_1812));
AND2X1 g62540(.A (WX5955), .B (n_2346), .Y (n_1811));
AND2X1 g62541(.A (WX8523), .B (n_2383), .Y (n_1810));
AND2X1 g62545(.A (WX5865), .B (n_2378), .Y (n_1809));
AND2X1 g62547(.A (WX5885), .B (n_2188), .Y (n_1808));
AND2X1 g62552(.A (WX7178), .B (n_2388), .Y (n_1807));
AND2X1 g62557(.A (WX4578), .B (n_2223), .Y (n_1806));
AND2X1 g62562(.A (WX9732), .B (n_2218), .Y (n_1805));
AND2X1 g62563(.A (WX11127), .B (n_2246), .Y (n_1804));
AND2X1 g62564(.A (WX5847), .B (n_2227), .Y (n_1803));
AND2X1 g62565(.A (WX8469), .B (n_2223), .Y (n_1802));
AND2X1 g62494(.A (WX2028), .B (n_2388), .Y (n_1801));
AND2X1 g62570(.A (WX11021), .B (n_2378), .Y (n_1800));
AND2X1 g62574(.A (WX4632), .B (n_2378), .Y (n_1799));
AND2X1 g62576(.A (WX5841), .B (n_2188), .Y (n_1798));
AND2X1 g62577(.A (WX5973), .B (n_2346), .Y (n_1797));
AND2X1 g62581(.A (WX11019), .B (n_2227), .Y (n_1796));
AND2X1 g62585(.A (WX5833), .B (n_2251), .Y (n_1795));
AND2X1 g62586(.A (WX5995), .B (n_2383), .Y (n_1794));
AND2X1 g62588(.A (WX3261), .B (n_2378), .Y (n_1793));
AND2X1 g62589(.A (WX7184), .B (n_2227), .Y (n_1792));
AND2X1 g62593(.A (WX11165), .B (n_2298), .Y (n_1791));
AND2X1 g62594(.A (WX8419), .B (n_2298), .Y (n_1790));
AND2X1 g62597(.A (WX5857), .B (n_2383), .Y (n_1789));
AND2X1 g62599(.A (WX4528), .B (n_2218), .Y (n_1788));
AND2X1 g62600(.A (WX5843), .B (n_2388), .Y (n_1787));
AND2X1 g62601(.A (WX5827), .B (n_2400), .Y (n_1786));
AND2X1 g62602(.A (WX7254), .B (n_2188), .Y (n_1785));
AND2X1 g62603(.A (WX5835), .B (n_2272), .Y (n_1784));
AND2X1 g62605(.A (WX3293), .B (n_2400), .Y (n_1783));
AND2X1 g62606(.A (WX9846), .B (n_2333), .Y (n_1782));
AND2X1 g62487(.A (WX5893), .B (n_2325), .Y (n_1781));
AND2X1 g62608(.A (WX9814), .B (n_2216), .Y (n_1780));
AND2X1 g62489(.A (WX2050), .B (n_2388), .Y (n_1779));
AND2X1 g62610(.A (WX4658), .B (n_2402), .Y (n_1778));
AND2X1 g62612(.A (WX5825), .B (n_2388), .Y (n_1777));
AND2X1 g62614(.A (WX3399), .B (n_2246), .Y (n_1776));
AND2X1 g62617(.A (WX8471), .B (n_2378), .Y (n_1775));
AND2X1 g62620(.A (WX7290), .B (n_2227), .Y (n_1774));
AND2X1 g62621(.A (WX11101), .B (n_2227), .Y (n_1773));
AND2X1 g62624(.A (WX8459), .B (n_2378), .Y (n_1772));
AND2X1 g62626(.A (WX4668), .B (n_2383), .Y (n_1771));
AND2X1 g62627(.A (WX4614), .B (n_2246), .Y (n_1770));
AND2X1 g62629(.A (WX4672), .B (n_2216), .Y (n_1769));
AND2X1 g62630(.A (WX9844), .B (n_2227), .Y (n_1768));
AND2X1 g62633(.A (WX3325), .B (n_2227), .Y (n_1767));
AND2X1 g62637(.A (WX9746), .B (n_2346), .Y (n_1766));
AND2X1 g62486(.A (WX7172), .B (n_2246), .Y (n_1765));
AND2X1 g62640(.A (WX8451), .B (n_2529), .Y (n_1764));
AND2X1 g62642(.A (WX5909), .B (n_2246), .Y (n_1763));
AND2X1 g62643(.A (WX8515), .B (n_2378), .Y (n_1762));
AND2X1 g62646(.A (WX7236), .B (n_2251), .Y (n_1761));
AND2X1 g62647(.A (WX4700), .B (n_2188), .Y (n_1760));
AND2X1 g62649(.A (WX4692), .B (n_2378), .Y (n_1759));
AND2X1 g62653(.A (WX8443), .B (n_2298), .Y (n_1758));
AND2X1 g62656(.A (WX2032), .B (n_2227), .Y (n_1757));
AND2X1 g62658(.A (WX11023), .B (n_2378), .Y (n_1756));
AND2X1 g62660(.A (WX3317), .B (n_2346), .Y (n_1755));
AND2X1 g62662(.A (WX2014), .B (n_2227), .Y (n_1754));
AND2X1 g62664(.A (WX2020), .B (n_2378), .Y (n_1753));
AND2X1 g62665(.A (WX6007), .B (n_2218), .Y (n_1752));
AND2X1 g62667(.A (WX4708), .B (n_2378), .Y (n_1751));
AND2X1 g62669(.A (WX2044), .B (n_2383), .Y (n_1750));
AND2X1 g62670(.A (WX2046), .B (n_2346), .Y (n_1749));
AND2X1 g62672(.A (WX2054), .B (n_2246), .Y (n_1748));
AND2X1 g62674(.A (WX5869), .B (n_2272), .Y (n_1747));
AND2X1 g62675(.A (WX11179), .B (n_2346), .Y (n_1746));
AND2X1 g62677(.A (WX11145), .B (n_2272), .Y (n_1745));
AND2X1 g62679(.A (WX2080), .B (n_2246), .Y (n_1744));
AND2X1 g62681(.A (WX2030), .B (n_2346), .Y (n_1743));
AND2X1 g62682(.A (WX11075), .B (n_2325), .Y (n_1742));
AND2X1 g62684(.A (WX3311), .B (n_2188), .Y (n_1741));
AND2X1 g62685(.A (WX9818), .B (n_2311), .Y (n_1740));
AND2X1 g62687(.A (WX2026), .B (n_2188), .Y (n_1739));
AND2X1 g62690(.A (WX5839), .B (n_2378), .Y (n_1738));
AND2X1 g62693(.A (WX11007), .B (n_2339), .Y (n_1737));
AND2X1 g62698(.A (WX8563), .B (n_2383), .Y (n_1736));
AND2X1 g62699(.A (WX3309), .B (n_2339), .Y (n_1735));
AND2X1 g62703(.A (WX8415), .B (n_2339), .Y (n_1734));
AND2X1 g62704(.A (WX9810), .B (n_2378), .Y (n_1733));
AND2X1 g62709(.A (WX3269), .B (n_2188), .Y (n_1732));
AND2X1 g62710(.A (WX7200), .B (n_2346), .Y (n_1731));
AND2X1 g62714(.A (WX7174), .B (n_2400), .Y (n_1730));
AND2X1 g62717(.A (WX8581), .B (n_2400), .Y (n_1729));
AND2X1 g62718(.A (WX5845), .B (n_2227), .Y (n_1728));
AND2X1 g62720(.A (WX9782), .B (n_2188), .Y (n_1727));
AND2X1 g62723(.A (WX8485), .B (n_2216), .Y (n_1726));
AND2X1 g62725(.A (WX8575), .B (n_2383), .Y (n_1725));
AND2X1 g62726(.A (WX8481), .B (n_2188), .Y (n_1724));
AND2X1 g62729(.A (WX4532), .B (n_2378), .Y (n_1723));
AND2X1 g62731(.A (WX11031), .B (n_2188), .Y (n_1722));
AND2X1 g62733(.A (WX7210), .B (n_2227), .Y (n_1721));
AND2X1 g62737(.A (WX6974), .B (n_2529), .Y (n_1720));
AND2X1 g62738(.A (WX7206), .B (n_2311), .Y (n_1719));
AND2X1 g62748(.A (WX3413), .B (n_2529), .Y (n_1718));
AND2X1 g62753(.A (WX3291), .B (n_2383), .Y (n_1717));
AND2X1 g62759(.A (WX4568), .B (n_2383), .Y (n_1716));
AND2X1 g62763(.A (WX11035), .B (n_2216), .Y (n_1715));
AND2X1 g62767(.A (WX3251), .B (n_2227), .Y (n_1714));
AND2X1 g62613(.A (WX7188), .B (n_2378), .Y (n_1713));
AND2X1 g61862(.A (WX9798), .B (n_2188), .Y (n_1712));
AND2X1 g62766(.A (WX11039), .B (n_2396), .Y (n_1711));
AND2X1 g62760(.A (WX8527), .B (n_2218), .Y (n_1710));
AND2X1 g62758(.A (WX7266), .B (n_2227), .Y (n_1709));
AND2X1 g62749(.A (WX8577), .B (n_2529), .Y (n_1708));
AND2X1 g62747(.A (WX10993), .B (n_2227), .Y (n_1707));
NOR2X1 g57543(.A (n_847), .B (n_1648), .Y (n_1706));
AND2X1 g62719(.A (WX5873), .B (n_2400), .Y (n_1702));
AND2X1 g61763(.A (WX5921), .B (n_2188), .Y (n_1701));
AND2X1 g61766(.A (WX9780), .B (n_2188), .Y (n_1700));
AND2X1 g62257(.A (WX7140), .B (n_2251), .Y (n_1699));
AND2X1 g62715(.A (WX3389), .B (n_2246), .Y (n_1698));
NOR2X1 g59240(.A (n_1190), .B (n_5712), .Y (n_1697));
NOR2X1 g59241(.A (n_1172), .B (n_5181), .Y (n_1696));
NOR2X1 g59243(.A (n_1077), .B (n_1425), .Y (n_1694));
NOR2X1 g59245(.A (n_1149), .B (n_1425), .Y (n_1693));
NOR2X1 g59246(.A (n_1185), .B (n_1425), .Y (n_1691));
NOR2X1 g59252(.A (n_1118), .B (n_1425), .Y (n_1690));
NOR2X1 g59253(.A (n_1049), .B (n_1425), .Y (n_1688));
NOR2X1 g59254(.A (n_1147), .B (n_5712), .Y (n_1687));
NOR2X1 g59255(.A (n_1109), .B (n_5712), .Y (n_1685));
NOR2X1 g59256(.A (n_1216), .B (n_1648), .Y (n_1684));
NOR2X1 g59259(.A (n_1194), .B (n_5181), .Y (n_1682));
NOR2X1 g59260(.A (n_1218), .B (n_5181), .Y (n_1681));
NOR2X1 g59261(.A (n_1267), .B (n_5181), .Y (n_1679));
AND2X1 g62711(.A (WX9752), .B (n_2227), .Y (n_1678));
NOR2X1 g59263(.A (n_1239), .B (n_1648), .Y (n_1677));
NOR2X1 g59264(.A (n_1229), .B (n_1425), .Y (n_1676));
NOR2X1 g59265(.A (n_1123), .B (n_5181), .Y (n_1675));
NOR2X1 g59267(.A (n_1217), .B (n_1648), .Y (n_1673));
AND2X1 g61757(.A (WX7180), .B (n_2246), .Y (n_1672));
AND2X1 g62700(.A (WX9710), .B (n_2378), .Y (n_1671));
NOR2X1 g59287(.A (n_1022), .B (n_5181), .Y (n_1670));
NOR2X1 g59288(.A (n_1209), .B (n_5181), .Y (n_1669));
NOR2X1 g59289(.A (n_1059), .B (n_5712), .Y (n_1668));
NOR2X1 g59290(.A (n_1208), .B (n_5712), .Y (n_1666));
NOR2X1 g59291(.A (n_1058), .B (n_5712), .Y (n_1665));
NOR2X1 g59292(.A (n_1207), .B (n_1425), .Y (n_1664));
NOR2X1 g59295(.A (n_1204), .B (n_1648), .Y (n_1662));
NOR2X1 g59296(.A (n_1060), .B (n_1648), .Y (n_1661));
NOR2X1 g59297(.A (n_1203), .B (n_1648), .Y (n_1660));
NOR2X1 g59298(.A (n_1202), .B (n_5712), .Y (n_1659));
NOR2X1 g59299(.A (n_1201), .B (n_5712), .Y (n_1658));
NOR2X1 g59300(.A (n_1045), .B (n_5181), .Y (n_1656));
NOR2X1 g59301(.A (n_1030), .B (n_5181), .Y (n_1655));
NOR2X1 g59302(.A (n_1199), .B (n_1425), .Y (n_1654));
NOR2X1 g59303(.A (n_1014), .B (n_1425), .Y (n_1652));
NOR2X1 g59304(.A (n_1250), .B (n_1648), .Y (n_1651));
NOR2X1 g59305(.A (n_1196), .B (n_1648), .Y (n_1650));
NOR2X1 g59306(.A (n_1062), .B (n_1648), .Y (n_1649));
NOR2X1 g59307(.A (n_1193), .B (n_1648), .Y (n_1647));
NOR2X1 g59308(.A (n_1192), .B (n_5181), .Y (n_1646));
NOR2X1 g59309(.A (n_1191), .B (n_5712), .Y (n_1645));
NOR2X1 g59310(.A (n_1188), .B (n_1648), .Y (n_1644));
NOR2X1 g59311(.A (n_1187), .B (n_1648), .Y (n_1642));
NOR2X1 g59312(.A (n_1251), .B (n_5712), .Y (n_1641));
NOR2X1 g59313(.A (n_1213), .B (n_5712), .Y (n_1640));
NOR2X1 g59314(.A (n_1184), .B (n_1425), .Y (n_1639));
NOR2X1 g59315(.A (n_1183), .B (n_1425), .Y (n_1638));
NOR2X1 g59316(.A (n_1098), .B (n_5181), .Y (n_1637));
NOR2X1 g59317(.A (n_1180), .B (n_5712), .Y (n_1636));
NOR2X1 g59318(.A (n_1179), .B (n_5712), .Y (n_1635));
NOR2X1 g59319(.A (n_1177), .B (n_5712), .Y (n_1633));
AND2X1 g62702(.A (WX7202), .B (n_2378), .Y (n_1632));
NOR2X1 g59322(.A (n_1175), .B (n_1648), .Y (n_1631));
NOR2X1 g59323(.A (n_1256), .B (n_5712), .Y (n_1629));
NOR2X1 g59324(.A (n_1260), .B (n_1648), .Y (n_1628));
NOR2X1 g59325(.A (n_1056), .B (n_1648), .Y (n_1627));
NOR2X1 g59326(.A (n_1057), .B (n_1425), .Y (n_1626));
NOR2X1 g59327(.A (n_1173), .B (n_1425), .Y (n_1625));
NOR2X1 g59328(.A (n_1171), .B (n_5712), .Y (n_1624));
NOR2X1 g59329(.A (n_1017), .B (n_5181), .Y (n_1623));
NOR2X1 g59332(.A (n_1169), .B (n_1648), .Y (n_1622));
NOR2X1 g59333(.A (n_1126), .B (n_1648), .Y (n_1620));
NOR2X1 g59334(.A (n_1253), .B (n_1425), .Y (n_1619));
NOR2X1 g59335(.A (n_1259), .B (n_1425), .Y (n_1618));
NOR2X1 g59336(.A (n_1225), .B (n_1425), .Y (n_1617));
NOR2X1 g59337(.A (n_1105), .B (n_1425), .Y (n_1615));
NOR2X1 g59340(.A (n_1166), .B (n_5712), .Y (n_1614));
NOR2X1 g59341(.A (n_1252), .B (n_5712), .Y (n_1613));
NOR2X1 g59342(.A (n_1164), .B (n_5181), .Y (n_1612));
NOR2X1 g59343(.A (n_1240), .B (n_5181), .Y (n_1611));
NOR2X1 g59344(.A (n_1163), .B (n_5712), .Y (n_1609));
NOR2X1 g59345(.A (n_1162), .B (n_5712), .Y (n_1608));
NOR2X1 g59346(.A (n_1161), .B (n_5181), .Y (n_1607));
NOR2X1 g59348(.A (n_1095), .B (n_5181), .Y (n_1606));
NOR2X1 g59349(.A (n_1262), .B (n_5181), .Y (n_1605));
NOR2X1 g59350(.A (n_1160), .B (n_1425), .Y (n_1604));
NOR2X1 g59351(.A (n_1024), .B (n_1425), .Y (n_1603));
NOR2X1 g59354(.A (n_1157), .B (n_1425), .Y (n_1601));
NOR2X1 g59355(.A (n_1156), .B (n_1425), .Y (n_1600));
NOR2X1 g59358(.A (n_1037), .B (n_1648), .Y (n_1599));
NOR2X1 g59359(.A (n_1258), .B (n_5712), .Y (n_1598));
NOR2X1 g59360(.A (n_1153), .B (n_5712), .Y (n_1597));
NOR2X1 g59361(.A (n_1025), .B (n_5712), .Y (n_1595));
NOR2X1 g59362(.A (n_1151), .B (n_1648), .Y (n_1594));
NOR2X1 g59363(.A (n_1215), .B (n_1648), .Y (n_1593));
NOR2X1 g59364(.A (n_1243), .B (n_5712), .Y (n_1592));
NOR2X1 g59366(.A (n_1146), .B (n_1648), .Y (n_1591));
NOR2X1 g59368(.A (n_1018), .B (n_5181), .Y (n_1590));
NOR2X1 g59369(.A (n_1144), .B (n_5181), .Y (n_1588));
NOR2X1 g59370(.A (n_1214), .B (n_5712), .Y (n_1587));
NOR2X1 g59371(.A (n_1143), .B (n_5712), .Y (n_1585));
NOR2X1 g59372(.A (n_1036), .B (n_5181), .Y (n_1584));
NOR2X1 g59373(.A (n_1034), .B (n_5181), .Y (n_1583));
NOR2X1 g59374(.A (n_1139), .B (n_1648), .Y (n_1582));
NOR2X1 g59375(.A (n_1138), .B (n_1648), .Y (n_1581));
NOR2X1 g59377(.A (n_1137), .B (n_5712), .Y (n_1580));
NOR2X1 g59380(.A (n_1134), .B (n_1648), .Y (n_1579));
NOR2X1 g59381(.A (n_1212), .B (n_1425), .Y (n_1577));
NOR2X1 g59382(.A (n_1117), .B (n_5712), .Y (n_1576));
NOR2X1 g59383(.A (n_1046), .B (n_5181), .Y (n_1575));
NOR2X1 g59384(.A (n_1140), .B (n_1648), .Y (n_1574));
NOR2X1 g59385(.A (n_1255), .B (n_1648), .Y (n_1573));
NOR2X1 g59387(.A (n_1127), .B (n_1425), .Y (n_1572));
NOR2X1 g59388(.A (n_1053), .B (n_5712), .Y (n_1571));
NOR2X1 g59389(.A (n_1261), .B (n_5712), .Y (n_1570));
NOR2X1 g59392(.A (n_1061), .B (n_5712), .Y (n_1568));
NOR2X1 g59393(.A (n_1125), .B (n_5712), .Y (n_1567));
AND2X1 g62226(.A (WX4592), .B (n_2383), .Y (n_1566));
NOR2X1 g59395(.A (n_1122), .B (n_5712), .Y (n_1565));
NOR2X1 g59398(.A (n_1220), .B (n_1425), .Y (n_1564));
NOR2X1 g59399(.A (n_1219), .B (n_1425), .Y (n_1563));
NOR2X1 g59400(.A (n_1152), .B (n_5712), .Y (n_1561));
NOR2X1 g59401(.A (n_1249), .B (n_5712), .Y (n_1560));
NOR2X1 g59402(.A (n_1112), .B (n_1425), .Y (n_1559));
NOR2X1 g59403(.A (n_1211), .B (n_1425), .Y (n_1558));
NOR2X1 g59404(.A (n_1241), .B (n_5712), .Y (n_1557));
NOR2X1 g59406(.A (n_1107), .B (n_5712), .Y (n_1555));
NOR2X1 g59407(.A (n_1040), .B (n_5712), .Y (n_1554));
NOR2X1 g59410(.A (n_1039), .B (n_5181), .Y (n_1553));
NOR2X1 g59411(.A (n_1103), .B (n_5181), .Y (n_1552));
NOR2X1 g59417(.A (n_1096), .B (n_5181), .Y (n_1551));
NOR2X1 g59418(.A (n_1021), .B (n_5712), .Y (n_1550));
NOR2X1 g59419(.A (n_1246), .B (n_5712), .Y (n_1548));
NOR2X1 g59420(.A (n_1092), .B (n_5712), .Y (n_1547));
NOR2X1 g59421(.A (n_1063), .B (n_5181), .Y (n_1546));
NOR2X1 g59423(.A (n_1090), .B (n_1648), .Y (n_1545));
NOR2X1 g59424(.A (n_1089), .B (n_5712), .Y (n_1544));
NOR2X1 g59425(.A (n_1050), .B (n_5712), .Y (n_1542));
NOR2X1 g59426(.A (n_1088), .B (n_5712), .Y (n_1541));
NOR2X1 g59427(.A (n_1165), .B (n_5181), .Y (n_1540));
NOR2X1 g59428(.A (n_1087), .B (n_1425), .Y (n_1539));
NOR2X1 g59429(.A (n_1189), .B (n_1425), .Y (n_1537));
NOR2X1 g59432(.A (n_1085), .B (n_1648), .Y (n_1536));
NOR2X1 g59433(.A (n_1013), .B (n_1425), .Y (n_1535));
NOR2X1 g59438(.A (n_1041), .B (n_5181), .Y (n_1534));
NOR2X1 g59439(.A (n_1081), .B (n_5181), .Y (n_1533));
NOR2X1 g59440(.A (n_1174), .B (n_1648), .Y (n_1531));
NOR2X1 g59441(.A (n_1224), .B (n_5181), .Y (n_1530));
NOR2X1 g59442(.A (n_1052), .B (n_5181), .Y (n_1529));
NOR2X1 g59443(.A (n_1080), .B (n_5181), .Y (n_1528));
NOR2X1 g59444(.A (n_1028), .B (n_5712), .Y (n_1527));
AND2X1 g61735(.A (WX9556), .B (n_2246), .Y (n_1526));
NOR2X1 g59445(.A (n_1078), .B (n_1648), .Y (n_1525));
NOR2X1 g59446(.A (n_1223), .B (n_1648), .Y (n_1524));
NOR2X1 g59454(.A (n_1071), .B (n_1648), .Y (n_1523));
NOR2X1 g59455(.A (n_1236), .B (n_1648), .Y (n_1522));
NOR2X1 g59456(.A (n_1070), .B (n_5181), .Y (n_1521));
NOR2X1 g59457(.A (n_1016), .B (n_5181), .Y (n_1519));
NOR2X1 g59458(.A (n_1069), .B (n_5712), .Y (n_1518));
NOR2X1 g59459(.A (n_1232), .B (n_5712), .Y (n_1517));
NOR2X1 g59461(.A (n_1067), .B (n_1648), .Y (n_1516));
NOR2X1 g59462(.A (n_1124), .B (n_5712), .Y (n_1515));
NOR2X1 g59463(.A (n_1197), .B (n_1648), .Y (n_1514));
NOR2X1 g59471(.A (n_1198), .B (n_5181), .Y (n_1513));
NOR2X1 g59472(.A (n_1031), .B (n_5181), .Y (n_1512));
NOR2X1 g59473(.A (n_1110), .B (n_1425), .Y (n_1511));
NOR2X1 g59474(.A (n_1206), .B (n_1425), .Y (n_1510));
NOR2X1 g59483(.A (n_1100), .B (n_1425), .Y (n_1509));
NOR2X1 g59484(.A (n_1133), .B (n_5712), .Y (n_1508));
NOR2X1 g59485(.A (n_1129), .B (n_5712), .Y (n_1507));
NOR2X1 g59486(.A (n_1141), .B (n_5712), .Y (n_1506));
NOR2X1 g59487(.A (n_1200), .B (n_5712), .Y (n_1504));
NOR2X1 g59489(.A (n_1178), .B (n_5712), .Y (n_1503));
NOR2X1 g59490(.A (n_1093), .B (n_5712), .Y (n_1502));
NOR2X1 g59492(.A (n_1115), .B (n_5712), .Y (n_1500));
NOR2X1 g59493(.A (n_1012), .B (n_5712), .Y (n_1499));
NOR2X1 g59495(.A (n_1130), .B (n_5712), .Y (n_1498));
NOR2X1 g59496(.A (n_1248), .B (n_1648), .Y (n_1497));
NOR2X1 g59497(.A (n_1159), .B (n_5712), .Y (n_1496));
AND2X1 g59498(.A (WX11053), .B (n_2325), .Y (n_1495));
AND2X1 g62676(.A (WX11129), .B (n_2346), .Y (n_1494));
AND2X1 g59512(.A (WX2002), .B (n_2346), .Y (n_1493));
AND2X1 g62671(.A (WX3359), .B (n_2333), .Y (n_1492));
AND2X1 g61705(.A (WX7198), .B (n_2311), .Y (n_1491));
AND2X1 g62663(.A (WX11155), .B (n_2251), .Y (n_1490));
AND2X1 g62181(.A (WX7262), .B (n_2223), .Y (n_1489));
AND2X1 g62548(.A (WX9794), .B (n_2383), .Y (n_1488));
AND2X1 g62659(.A (WX8265), .B (n_2198), .Y (n_1487));
AND2X1 g62657(.A (WX9848), .B (n_2272), .Y (n_1486));
AND2X1 g61684(.A (WX8533), .B (n_2325), .Y (n_1485));
AND2X1 g62638(.A (WX9874), .B (n_2383), .Y (n_1484));
AND2X1 g61663(.A (WX11045), .B (n_2311), .Y (n_1483));
AND2X1 g62636(.A (WX11069), .B (n_2371), .Y (n_1482));
AND2X1 g61655(.A (WX11041), .B (n_2527), .Y (n_1481));
AND2X1 g61650(.A (WX9786), .B (n_2383), .Y (n_1480));
AND2X1 g61640(.A (WX2072), .B (n_2325), .Y (n_1479));
AND2X1 g62632(.A (WX4648), .B (n_2227), .Y (n_1478));
AND2X1 g62625(.A (WX5817), .B (n_2527), .Y (n_1477));
AND2X1 g62622(.A (WX5837), .B (n_2400), .Y (n_1476));
AOI21X1 g57873(.A0 (_2107_), .A1 (WX837), .B0 (n_1038), .Y (n_1473));
AND2X1 g61631(.A (WX7284), .B (n_2527), .Y (n_1472));
AND2X1 g62554(.A (WX5821), .B (n_2227), .Y (n_1471));
AND2X1 g61607(.A (WX11167), .B (n_2227), .Y (n_1470));
INVX4 g63523(.A (n_2227), .Y (n_3690));
NOR2X1 g61584(.A (n_5181), .B (n_35), .Y (n_1465));
NOR2X1 g56990(.A (WX5659), .B (n_1648), .Y (n_1464));
NOR2X1 g62598(.A (n_1425), .B (n_2), .Y (n_1462));
NOR2X1 g62595(.A (n_5181), .B (n_970), .Y (n_1461));
NAND2X1 g60725(.A (n_597), .B (n_596), .Y (n_2511));
NAND2X1 g60796(.A (n_568), .B (n_590), .Y (n_2498));
NAND2X1 g60808(.A (n_582), .B (n_583), .Y (n_2494));
NOR2X1 g57058(.A (WX6952), .B (n_1648), .Y (n_1459));
NOR2X1 g62566(.A (n_5181), .B (n_112), .Y (n_1458));
NOR2X1 g55933(.A (n_1425), .B (n_3685), .Y (n_1456));
NAND2X1 g60903(.A (n_578), .B (n_576), .Y (n_2472));
NAND2X1 g60951(.A (n_548), .B (n_771), .Y (n_2468));
NOR2X1 g57096(.A (WX8245), .B (n_1648), .Y (n_1454));
NAND2X1 g60965(.A (n_570), .B (n_569), .Y (n_2466));
NAND2X1 g61011(.A (n_564), .B (n_563), .Y (n_2458));
NAND2X1 g61058(.A (n_593), .B (n_573), .Y (n_2453));
NAND2X1 g61092(.A (n_559), .B (n_547), .Y (n_2443));
NAND2X1 g61152(.A (n_557), .B (n_555), .Y (n_2437));
NOR2X1 g57161(.A (WX9538), .B (n_1425), .Y (n_1453));
NAND2X1 g61220(.A (n_545), .B (n_544), .Y (n_2422));
NOR2X1 g61559(.A (n_1451), .B (n_1425), .Y (n_1452));
NOR2X1 g61565(.A (n_1449), .B (n_5181), .Y (n_1450));
NOR2X1 g61579(.A (n_5181), .B (n_69), .Y (n_1448));
NOR2X1 g61588(.A (n_5181), .B (n_87), .Y (n_1447));
NOR2X1 g61605(.A (n_1425), .B (n_81), .Y (n_1446));
NOR2X1 g61608(.A (n_1425), .B (n_4), .Y (n_1444));
NOR2X1 g61612(.A (n_1442), .B (n_1425), .Y (n_1443));
NOR2X1 g61624(.A (n_1425), .B (n_951), .Y (n_1441));
NOR2X1 g61633(.A (n_1425), .B (n_1006), .Y (n_1440));
NOR2X1 g61636(.A (n_1437), .B (n_1425), .Y (n_1438));
NOR2X1 g61662(.A (n_5181), .B (n_67), .Y (n_1436));
NOR2X1 g61683(.A (n_1425), .B (n_119), .Y (n_1435));
NOR2X1 g61696(.A (n_5181), .B (n_1001), .Y (n_1433));
NOR2X1 g61736(.A (n_1431), .B (n_5712), .Y (n_1432));
NOR2X1 g61740(.A (n_1429), .B (n_5712), .Y (n_1430));
NOR2X1 g61748(.A (n_1427), .B (n_5181), .Y (n_1428));
NOR2X1 g61758(.A (n_1425), .B (n_12), .Y (n_1426));
NOR2X1 g58602(.A (n_5181), .B (n_0), .Y (n_1424));
NOR2X1 g61764(.A (n_1425), .B (n_940), .Y (n_1423));
NOR2X1 g61767(.A (n_1421), .B (n_1425), .Y (n_1422));
NOR2X1 g61776(.A (n_1419), .B (n_1425), .Y (n_1420));
NOR2X1 g61780(.A (n_1425), .B (n_958), .Y (n_1418));
NOR2X1 g61786(.A (n_1425), .B (n_56), .Y (n_1417));
NOR2X1 g61787(.A (n_1425), .B (n_109), .Y (n_1415));
NOR2X1 g61798(.A (n_5181), .B (n_52), .Y (n_1414));
NOR2X1 g61813(.A (n_1412), .B (n_1648), .Y (n_1413));
NOR2X1 g61818(.A (n_5181), .B (n_32), .Y (n_1411));
NOR2X1 g61822(.A (n_1425), .B (n_96), .Y (n_1410));
NOR2X1 g61844(.A (n_1425), .B (n_985), .Y (n_1409));
NOR2X1 g61853(.A (n_5181), .B (n_14), .Y (n_1407));
NOR2X1 g61875(.A (n_1425), .B (n_19), .Y (n_1405));
NOR2X1 g61878(.A (n_1425), .B (n_981), .Y (n_1404));
NOR2X1 g61880(.A (n_1425), .B (n_913), .Y (n_1403));
NOR2X1 g61895(.A (n_1425), .B (n_975), .Y (n_1402));
NOR2X1 g61924(.A (n_1425), .B (n_101), .Y (n_1400));
NOR2X1 g61927(.A (n_5181), .B (n_28), .Y (n_1399));
NOR2X1 g61928(.A (n_5181), .B (n_118), .Y (n_1398));
NOR2X1 g61930(.A (n_5181), .B (n_995), .Y (n_1396));
NOR2X1 g61945(.A (n_5181), .B (n_117), .Y (n_1395));
NOR2X1 g61951(.A (n_1425), .B (n_990), .Y (n_1393));
NOR2X1 g61974(.A (n_5181), .B (n_16), .Y (n_1391));
NOR2X1 g61984(.A (n_5181), .B (n_1004), .Y (n_1389));
NOR2X1 g61989(.A (n_1425), .B (n_46), .Y (n_1388));
NOR2X1 g62005(.A (n_5181), .B (n_41), .Y (n_1387));
NOR2X1 g62007(.A (n_1425), .B (n_18), .Y (n_1386));
NOR2X1 g62008(.A (n_5181), .B (n_51), .Y (n_1385));
NOR2X1 g62042(.A (n_5181), .B (n_130), .Y (n_1384));
NOR2X1 g62045(.A (n_5181), .B (n_929), .Y (n_1382));
NOR2X1 g62046(.A (n_5181), .B (n_68), .Y (n_1381));
NOR2X1 g62051(.A (n_5181), .B (n_3), .Y (n_1380));
NOR2X1 g62073(.A (n_1425), .B (n_79), .Y (n_1379));
NOR2X1 g62085(.A (n_1425), .B (n_105), .Y (n_1378));
NOR2X1 g62102(.A (n_1425), .B (n_111), .Y (n_1377));
NOR2X1 g62110(.A (n_1374), .B (n_1648), .Y (n_1375));
NOR2X1 g62153(.A (n_1425), .B (n_964), .Y (n_1373));
NOR2X1 g62169(.A (n_1425), .B (n_948), .Y (n_1372));
NOR2X1 g62173(.A (n_1425), .B (n_24), .Y (n_1371));
NOR2X1 g62179(.A (n_1425), .B (n_70), .Y (n_1370));
NOR2X1 g62186(.A (n_1425), .B (n_73), .Y (n_1369));
NOR2X1 g62193(.A (n_1425), .B (n_938), .Y (n_1367));
NOR2X1 g62200(.A (n_5181), .B (n_38), .Y (n_1366));
NOR2X1 g62223(.A (n_1425), .B (n_905), .Y (n_1365));
NOR2X1 g62225(.A (n_5181), .B (n_987), .Y (n_1364));
NOR2X1 g62250(.A (n_1425), .B (n_129), .Y (n_1362));
NOR2X1 g62284(.A (n_1359), .B (n_1425), .Y (n_1360));
NOR2X1 g62307(.A (n_1357), .B (n_5181), .Y (n_1358));
NOR2X1 g62309(.A (n_1425), .B (n_43), .Y (n_1356));
NOR2X1 g62330(.A (n_1425), .B (n_71), .Y (n_1355));
NOR2X1 g62338(.A (n_1425), .B (n_83), .Y (n_1354));
NOR2X1 g62342(.A (n_5181), .B (n_21), .Y (n_1353));
NOR2X1 g62353(.A (n_1425), .B (n_956), .Y (n_1352));
NOR2X1 g62356(.A (n_1350), .B (n_1425), .Y (n_1351));
NOR2X1 g62359(.A (n_1348), .B (n_1425), .Y (n_1349));
NOR2X1 g62365(.A (n_1425), .B (n_89), .Y (n_1347));
NOR2X1 g62366(.A (n_1345), .B (n_5181), .Y (n_1346));
NOR2X1 g62368(.A (n_1425), .B (n_58), .Y (n_1344));
NOR2X1 g62371(.A (n_1341), .B (n_5181), .Y (n_1342));
NOR2X1 g62469(.A (n_1339), .B (n_5181), .Y (n_1340));
NOR2X1 g62473(.A (n_1337), .B (n_1425), .Y (n_1338));
NOR2X1 g62474(.A (n_1335), .B (n_1425), .Y (n_1336));
NOR2X1 g62478(.A (n_5181), .B (n_104), .Y (n_1334));
NOR2X1 g62488(.A (n_1425), .B (n_98), .Y (n_1333));
NOR2X1 g62493(.A (n_5181), .B (n_992), .Y (n_1332));
NOR2X1 g62498(.A (n_1425), .B (n_932), .Y (n_1330));
NOR2X1 g62537(.A (n_1328), .B (n_1425), .Y (n_1329));
NOR2X1 g62543(.A (n_5181), .B (n_27), .Y (n_1327));
NOR2X1 g62584(.A (n_5181), .B (n_997), .Y (n_1326));
NOR2X1 g62604(.A (n_5181), .B (n_48), .Y (n_1325));
NOR2X1 g62607(.A (n_1323), .B (n_1425), .Y (n_1324));
NOR2X1 g62635(.A (n_1425), .B (n_63), .Y (n_1322));
NOR2X1 g62644(.A (n_1320), .B (n_1648), .Y (n_1321));
NOR2X1 g62655(.A (n_1318), .B (n_5181), .Y (n_1319));
NOR2X1 g62678(.A (n_5181), .B (n_973), .Y (n_1317));
NOR2X1 g62741(.A (n_1315), .B (n_5712), .Y (n_1316));
NOR2X1 g62742(.A (n_5181), .B (n_113), .Y (n_1314));
NOR2X1 g62744(.A (n_5181), .B (n_36), .Y (n_1313));
NOR2X1 g62755(.A (n_1425), .B (n_20), .Y (n_1312));
NOR2X1 g62756(.A (n_1425), .B (n_106), .Y (n_1311));
NOR2X1 g62761(.A (n_1309), .B (n_1425), .Y (n_1310));
NOR2X1 g62768(.A (n_1425), .B (n_44), .Y (n_1308));
NOR2X1 g62746(.A (n_1425), .B (n_100), .Y (n_1307));
NOR2X1 g62745(.A (n_5181), .B (n_65), .Y (n_1306));
INVX4 g63039(.A (n_1460), .Y (n_3058));
INVX4 g63043(.A (n_1305), .Y (n_3106));
INVX1 g63227(.A (n_1278), .Y (n_2993));
INVX1 g63230(.A (n_1278), .Y (n_3044));
INVX1 g63231(.A (n_1278), .Y (n_2996));
INVX1 g63233(.A (n_1278), .Y (n_2976));
INVX4 g63503(.A (n_2378), .Y (n_2605));
INVX8 g63530(.A (n_2227), .Y (n_2851));
INVX8 g63543(.A (n_1297), .Y (n_3188));
INVX8 g63554(.A (n_2227), .Y (n_2620));
INVX4 g63584(.A (n_6428), .Y (n_2938));
INVX8 g63599(.A (n_1294), .Y (n_3072));
NOR2X1 g62686(.A (n_5181), .B (n_962), .Y (n_1291));
NOR2X1 g59500(.A (n_1425), .B (n_95), .Y (n_1290));
NOR2X1 g62651(.A (n_1288), .B (n_5712), .Y (n_1289));
NOR2X1 g62650(.A (n_1286), .B (n_1648), .Y (n_1287));
NOR2X1 g62641(.A (n_1284), .B (n_5712), .Y (n_1285));
NOR2X1 g61688(.A (n_1282), .B (n_5712), .Y (n_1283));
INVX4 g63665(.A (n_1281), .Y (n_2945));
INVX4 g63659(.A (n_3120), .Y (n_3086));
NOR2X1 g62553(.A (n_5181), .B (n_49), .Y (n_1280));
NAND2X1 g61084(.A (n_551), .B (n_566), .Y (n_2446));
NOR2X1 g56884(.A (WX3073), .B (n_1648), .Y (n_1279));
INVX1 g63232(.A (n_1278), .Y (n_3004));
INVX1 g63228(.A (n_1278), .Y (n_3056));
INVX1 g63226(.A (n_1278), .Y (n_3105));
INVX1 g63225(.A (n_1278), .Y (n_3103));
NOR2X1 g61621(.A (n_1425), .B (n_953), .Y (n_1277));
INVX4 g63591(.A (n_1276), .Y (n_3041));
NOR2X1 g61609(.A (n_1425), .B (n_944), .Y (n_1275));
NOR2X1 g61593(.A (_2078_), .B (WX895), .Y (n_1272));
AOI21X1 g60389(.A0 (WX9936), .A1 (_2307_), .B0 (n_412), .Y (n_1268));
AOI21X1 g60390(.A0 (WX9930), .A1 (_2310_), .B0 (n_302), .Y (n_1267));
AOI21X1 g60391(.A0 (WX7302), .A1 (_2267_), .B0 (n_419), .Y (n_1265));
AOI21X1 g60392(.A0 (WX11213), .A1 (_2347_), .B0 (n_285), .Y (n_1264));
AOI21X1 g60393(.A0 (WX6041), .A1 (_2219_), .B0 (n_324), .Y (n_1263));
BUFX3 g63475(.A (n_2298), .Y (n_2216));
AOI21X1 g60394(.A0 (WX4732), .A1 (_2195_), .B0 (n_332), .Y (n_1262));
AOI21X1 g60395(.A0 (WX6069), .A1 (_2205_), .B0 (n_328), .Y (n_1261));
AOI21X1 g60396(.A0 (WX3435), .A1 (_2165_), .B0 (n_427), .Y (n_1260));
AOI21X1 g60397(.A0 (WX4766), .A1 (_2178_), .B0 (n_145), .Y (n_1259));
AOI21X1 g60398(.A0 (WX6059), .A1 (_2210_), .B0 (n_200), .Y (n_1258));
AOI21X1 g60400(.A0 (WX4746), .A1 (_2204_), .B0 (n_422), .Y (n_1257));
BUFX3 g63477(.A (n_2298), .Y (n_2188));
AOI21X1 g60401(.A0 (WX3437), .A1 (_2164_), .B0 (n_232), .Y (n_1256));
AOI21X1 g60403(.A0 (WX7326), .A1 (_2255_), .B0 (n_148), .Y (n_1255));
AOI21X1 g60404(.A0 (WX2184), .A1 (_2140_), .B0 (n_469), .Y (n_1254));
AOI21X1 g60406(.A0 (WX4768), .A1 (_2177_), .B0 (n_198), .Y (n_1253));
AOI21X1 g60407(.A0 (WX4750), .A1 (_2186_), .B0 (n_254), .Y (n_1252));
AOI21X1 g60408(.A0 (WX3469), .A1 (_2148_), .B0 (n_377), .Y (n_1251));
AOI21X1 g60409(.A0 (WX2138), .A1 (_2135_), .B0 (n_136), .Y (n_1250));
AOI21X1 g60410(.A0 (WX8631), .A1 (_2281_), .B0 (n_181), .Y (n_1249));
AOI21X1 g60411(.A0 (WX8643), .A1 (_2275_), .B0 (n_415), .Y (n_1248));
AOI21X1 g60412(.A0 (WX11203), .A1 (_2352_), .B0 (n_151), .Y (n_1247));
AOI21X1 g60413(.A0 (WX9922), .A1 (_2314_), .B0 (n_428), .Y (n_1246));
AOI21X1 g60414(.A0 (WX8605), .A1 (_2294_), .B0 (n_317), .Y (n_1245));
AOI21X1 g60415(.A0 (WX9946), .A1 (_2302_), .B0 (n_407), .Y (n_1244));
AOI21X1 g60416(.A0 (WX6047), .A1 (_2216_), .B0 (n_453), .Y (n_1243));
AOI21X1 g60417(.A0 (WX7310), .A1 (_2263_), .B0 (n_433), .Y (n_1242));
AOI21X1 g60418(.A0 (WX8621), .A1 (_2286_), .B0 (n_461), .Y (n_1241));
AOI21X1 g60419(.A0 (WX4744), .A1 (_2189_), .B0 (n_199), .Y (n_1240));
AOI21X1 g60420(.A0 (WX7340), .A1 (_2248_), .B0 (n_157), .Y (n_1239));
INVX4 g63466(.A (n_2298), .Y (n_2849));
AOI21X1 g60421(.A0 (WX7342), .A1 (_2268_), .B0 (n_150), .Y (n_1237));
AOI21X1 g60422(.A0 (WX11195), .A1 (_2356_), .B0 (n_349), .Y (n_1236));
AOI21X1 g60423(.A0 (WX4728), .A1 (_2197_), .B0 (n_479), .Y (n_1235));
AOI21X1 g60424(.A0 (WX4754), .A1 (_2184_), .B0 (n_192), .Y (n_1234));
AOI21X1 g60425(.A0 (WX3425), .A1 (_2170_), .B0 (n_176), .Y (n_1233));
AOI21X1 g60426(.A0 (WX11187), .A1 (_2360_), .B0 (n_405), .Y (n_1232));
AOI21X1 g60427(.A0 (WX2160), .A1 (_2140_), .B0 (n_306), .Y (n_1231));
AOI21X1 g60429(.A0 (WX11241), .A1 (_2333_), .B0 (n_153), .Y (n_1230));
AOI21X1 g60430(.A0 (WX6061), .A1 (_2209_), .B0 (n_178), .Y (n_1229));
AOI21X1 g60432(.A0 (WX8609), .A1 (_2292_), .B0 (n_410), .Y (n_1228));
AOI21X1 g60433(.A0 (WX3441), .A1 (_2162_), .B0 (n_341), .Y (n_1227));
AOI21X1 g60434(.A0 (WX7354), .A1 (_2241_), .B0 (n_316), .Y (n_1226));
AOI21X1 g60435(.A0 (WX4764), .A1 (_2179_), .B0 (n_142), .Y (n_1225));
AOI21X1 g60436(.A0 (WX11229), .A1 (_2339_), .B0 (n_386), .Y (n_1224));
AOI21X1 g60437(.A0 (WX11217), .A1 (_2345_), .B0 (n_194), .Y (n_1223));
AOI21X1 g60438(.A0 (WX8651), .A1 (_2271_), .B0 (n_382), .Y (n_1222));
AOI21X1 g60439(.A0 (WX2170), .A1 (_2140_), .B0 (n_228), .Y (n_1221));
AOI21X1 g60441(.A0 (WX8645), .A1 (_2274_), .B0 (n_440), .Y (n_1220));
AOI21X1 g60442(.A0 (WX8641), .A1 (_2276_), .B0 (n_213), .Y (n_1219));
AOI21X1 g60443(.A0 (WX7328), .A1 (_2254_), .B0 (n_468), .Y (n_1218));
AOI21X1 g60444(.A0 (WX8607), .A1 (_2293_), .B0 (n_362), .Y (n_1217));
AOI21X1 g60445(.A0 (WX7362), .A1 (_2237_), .B0 (n_227), .Y (n_1216));
AOI21X1 g60446(.A0 (WX6051), .A1 (_2214_), .B0 (n_172), .Y (n_1215));
AOI21X1 g60447(.A0 (WX6023), .A1 (_2228_), .B0 (n_295), .Y (n_1214));
AOI21X1 g60448(.A0 (WX3465), .A1 (_2150_), .B0 (n_374), .Y (n_1213));
AOI21X1 g60450(.A0 (WX6025), .A1 (_2227_), .B0 (n_408), .Y (n_1212));
AOI21X1 g60454(.A0 (WX8627), .A1 (_2283_), .B0 (n_318), .Y (n_1211));
AOI21X1 g60467(.A0 (WX4770), .A1 (_2204_), .B0 (n_169), .Y (n_1210));
AOI21X1 g60468(.A0 (WX2190), .A1 (_2109_), .B0 (n_376), .Y (n_1209));
AOI21X1 g60469(.A0 (WX2186), .A1 (_2111_), .B0 (n_291), .Y (n_1208));
AOI21X1 g60470(.A0 (WX2180), .A1 (_2114_), .B0 (n_399), .Y (n_1207));
AOI21X1 g60471(.A0 (WX2176), .A1 (_2116_), .B0 (n_385), .Y (n_1206));
AOI21X1 g60472(.A0 (WX2172), .A1 (_2118_), .B0 (n_185), .Y (n_1205));
AOI21X1 g60473(.A0 (WX2166), .A1 (_2121_), .B0 (n_326), .Y (n_1204));
AOI21X1 g60474(.A0 (WX2162), .A1 (_2123_), .B0 (n_209), .Y (n_1203));
AOI21X1 g60475(.A0 (WX2158), .A1 (_2125_), .B0 (n_235), .Y (n_1202));
AOI21X1 g60476(.A0 (WX2156), .A1 (_2126_), .B0 (n_365), .Y (n_1201));
AOI21X1 g60477(.A0 (WX2152), .A1 (_2128_), .B0 (n_325), .Y (n_1200));
AOI21X1 g60478(.A0 (WX2144), .A1 (_2132_), .B0 (n_205), .Y (n_1199));
AOI21X1 g60479(.A0 (WX2140), .A1 (_2134_), .B0 (n_304), .Y (n_1198));
AOI21X1 g60480(.A0 (WX2136), .A1 (_2136_), .B0 (n_373), .Y (n_1197));
AOI21X1 g60481(.A0 (WX2134), .A1 (_2137_), .B0 (n_247), .Y (n_1196));
AOI21X1 g60482(.A0 (WX2132), .A1 (_2138_), .B0 (n_229), .Y (n_1195));
AOI21X1 g60483(.A0 (WX3485), .A1 (_2172_), .B0 (n_171), .Y (n_1194));
AOI21X1 g60484(.A0 (WX3483), .A1 (_2141_), .B0 (n_402), .Y (n_1193));
AOI21X1 g60485(.A0 (WX3481), .A1 (_2142_), .B0 (n_401), .Y (n_1192));
AOI21X1 g60486(.A0 (WX3479), .A1 (_2143_), .B0 (n_314), .Y (n_1191));
AOI21X1 g60487(.A0 (WX3475), .A1 (_2145_), .B0 (n_464), .Y (n_1190));
AOI21X1 g60488(.A0 (WX9900), .A1 (_2325_), .B0 (n_135), .Y (n_1189));
AOI21X1 g60489(.A0 (WX3473), .A1 (_2146_), .B0 (n_489), .Y (n_1188));
AOI21X1 g60490(.A0 (WX3471), .A1 (_2147_), .B0 (n_313), .Y (n_1187));
AOI21X1 g60491(.A0 (WX3463), .A1 (_2172_), .B0 (n_457), .Y (n_1186));
AOI21X1 g60492(.A0 (WX3461), .A1 (_2152_), .B0 (n_423), .Y (n_1185));
AOI21X1 g60493(.A0 (WX3459), .A1 (_2153_), .B0 (n_488), .Y (n_1184));
AOI21X1 g60494(.A0 (WX3457), .A1 (_2154_), .B0 (n_414), .Y (n_1183));
AOI21X1 g60495(.A0 (WX9940), .A1 (_2305_), .B0 (n_131), .Y (n_1182));
AOI21X1 g60496(.A0 (WX3453), .A1 (_2172_), .B0 (n_356), .Y (n_1181));
AOI21X1 g60497(.A0 (WX3451), .A1 (_2157_), .B0 (n_206), .Y (n_1180));
AOI21X1 g60498(.A0 (WX3449), .A1 (_2158_), .B0 (n_396), .Y (n_1179));
AOI21X1 g60499(.A0 (WX3447), .A1 (_2159_), .B0 (n_170), .Y (n_1178));
AOI21X1 g60500(.A0 (WX3445), .A1 (_2160_), .B0 (n_389), .Y (n_1177));
AOI21X1 g60501(.A0 (WX3443), .A1 (_2161_), .B0 (n_299), .Y (n_1176));
AOI21X1 g60502(.A0 (WX3439), .A1 (_2163_), .B0 (n_395), .Y (n_1175));
AOI21X1 g60503(.A0 (WX11231), .A1 (_2338_), .B0 (n_257), .Y (n_1174));
AOI21X1 g60504(.A0 (WX3429), .A1 (_2168_), .B0 (n_460), .Y (n_1173));
AOI21X1 g60505(.A0 (WX3427), .A1 (_2169_), .B0 (n_387), .Y (n_1172));
AOI21X1 g60506(.A0 (WX3423), .A1 (_2171_), .B0 (n_394), .Y (n_1171));
AOI21X1 g60507(.A0 (WX4776), .A1 (_2173_), .B0 (n_184), .Y (n_1170));
AOI21X1 g60508(.A0 (WX4772), .A1 (_2175_), .B0 (n_391), .Y (n_1169));
AOI21X1 g60509(.A0 (WX4762), .A1 (_2180_), .B0 (n_141), .Y (n_1168));
AOI21X1 g60510(.A0 (WX4758), .A1 (_2182_), .B0 (n_163), .Y (n_1167));
AOI21X1 g60511(.A0 (WX4752), .A1 (_2185_), .B0 (n_322), .Y (n_1166));
AOI21X1 g60512(.A0 (WX9904), .A1 (_2323_), .B0 (n_329), .Y (n_1165));
AOI21X1 g60513(.A0 (WX4748), .A1 (_2187_), .B0 (n_154), .Y (n_1164));
AOI21X1 g60514(.A0 (WX4742), .A1 (_2190_), .B0 (n_189), .Y (n_1163));
AOI21X1 g60515(.A0 (WX4740), .A1 (_2191_), .B0 (n_179), .Y (n_1162));
AOI21X1 g60516(.A0 (WX4738), .A1 (_2192_), .B0 (n_173), .Y (n_1161));
AOI21X1 g60517(.A0 (WX4730), .A1 (_2196_), .B0 (n_353), .Y (n_1160));
AOI21X1 g60518(.A0 (WX4726), .A1 (_2198_), .B0 (n_357), .Y (n_1159));
AOI21X1 g60519(.A0 (WX4722), .A1 (_2200_), .B0 (n_331), .Y (n_1158));
AOI21X1 g60520(.A0 (WX4718), .A1 (_2202_), .B0 (n_162), .Y (n_1157));
AOI21X1 g60521(.A0 (WX4716), .A1 (_2203_), .B0 (n_300), .Y (n_1156));
AOI21X1 g60522(.A0 (WX6067), .A1 (_2206_), .B0 (n_315), .Y (n_1155));
AOI21X1 g60523(.A0 (WX6063), .A1 (_2236_), .B0 (n_212), .Y (n_1154));
AOI21X1 g60524(.A0 (WX6057), .A1 (_2211_), .B0 (n_406), .Y (n_1153));
AOI21X1 g60525(.A0 (WX8637), .A1 (_2278_), .B0 (n_366), .Y (n_1152));
AOI21X1 g60526(.A0 (WX6053), .A1 (_2213_), .B0 (n_397), .Y (n_1151));
AOI21X1 g60527(.A0 (WX6049), .A1 (_2236_), .B0 (n_307), .Y (n_1150));
AOI21X1 g60528(.A0 (WX6043), .A1 (_2218_), .B0 (n_470), .Y (n_1149));
AOI21X1 g60529(.A0 (WX6039), .A1 (_2236_), .B0 (n_347), .Y (n_1148));
AOI21X1 g60530(.A0 (WX6037), .A1 (_2221_), .B0 (n_301), .Y (n_1147));
AOI21X1 g60531(.A0 (WX6035), .A1 (_2222_), .B0 (n_392), .Y (n_1146));
AOI21X1 g60532(.A0 (WX6033), .A1 (_2223_), .B0 (n_164), .Y (n_1145));
AOI21X1 g60533(.A0 (WX6029), .A1 (_2225_), .B0 (n_372), .Y (n_1144));
AOI21X1 g60534(.A0 (WX6021), .A1 (_2229_), .B0 (n_156), .Y (n_1143));
AOI21X1 g60535(.A0 (WX6017), .A1 (_2231_), .B0 (n_418), .Y (n_1142));
AOI21X1 g60536(.A0 (WX6013), .A1 (_2233_), .B0 (n_133), .Y (n_1141));
AOI21X1 g60537(.A0 (WX7330), .A1 (_2253_), .B0 (n_256), .Y (n_1140));
AOI21X1 g60538(.A0 (WX6011), .A1 (_2234_), .B0 (n_339), .Y (n_1139));
AOI21X1 g60539(.A0 (WX6009), .A1 (_2235_), .B0 (n_166), .Y (n_1138));
AOI21X1 g60540(.A0 (WX7360), .A1 (_2238_), .B0 (n_177), .Y (n_1137));
AOI21X1 g60541(.A0 (WX7358), .A1 (_2239_), .B0 (n_211), .Y (n_1136));
AOI21X1 g60542(.A0 (WX7356), .A1 (_2268_), .B0 (n_180), .Y (n_1135));
AOI21X1 g60543(.A0 (WX7352), .A1 (_2242_), .B0 (n_231), .Y (n_1134));
AOI21X1 g60544(.A0 (WX7344), .A1 (_2246_), .B0 (n_350), .Y (n_1133));
AOI21X1 g60545(.A0 (WX11183), .A1 (_2362_), .B0 (n_409), .Y (n_1132));
AOI21X1 g60546(.A0 (WX7338), .A1 (_2249_), .B0 (n_384), .Y (n_1131));
AOI21X1 g60547(.A0 (WX7334), .A1 (_2251_), .B0 (n_167), .Y (n_1130));
AOI21X1 g60548(.A0 (WX7324), .A1 (_2256_), .B0 (n_230), .Y (n_1129));
AOI21X1 g60549(.A0 (WX7322), .A1 (_2257_), .B0 (n_416), .Y (n_1128));
AOI21X1 g60550(.A0 (WX7320), .A1 (_2258_), .B0 (n_233), .Y (n_1127));
AOI21X1 g60551(.A0 (WX7316), .A1 (_2260_), .B0 (n_195), .Y (n_1126));
AOI21X1 g60552(.A0 (WX7306), .A1 (_2265_), .B0 (n_380), .Y (n_1125));
AOI21X1 g60553(.A0 (WX7304), .A1 (_2266_), .B0 (n_334), .Y (n_1124));
AOI21X1 g60554(.A0 (WX8657), .A1 (_2300_), .B0 (n_447), .Y (n_1123));
AOI21X1 g60555(.A0 (WX8655), .A1 (_2269_), .B0 (n_289), .Y (n_1122));
AOI21X1 g60556(.A0 (WX8653), .A1 (_2270_), .B0 (n_146), .Y (n_1121));
AOI21X1 g60557(.A0 (WX8649), .A1 (_2300_), .B0 (n_369), .Y (n_1120));
AOI21X1 g60558(.A0 (WX4720), .A1 (_2201_), .B0 (n_465), .Y (n_1119));
AOI21X1 g60559(.A0 (WX8601), .A1 (_2296_), .B0 (n_147), .Y (n_1118));
AOI21X1 g60560(.A0 (WX8647), .A1 (_2273_), .B0 (n_417), .Y (n_1117));
AOI21X1 g60561(.A0 (WX7332), .A1 (_2268_), .B0 (n_393), .Y (n_1116));
AOI21X1 g60562(.A0 (WX8639), .A1 (_2277_), .B0 (n_288), .Y (n_1115));
AOI21X1 g60563(.A0 (WX8635), .A1 (_2300_), .B0 (n_426), .Y (n_1114));
AOI21X1 g60564(.A0 (WX8633), .A1 (_2280_), .B0 (n_225), .Y (n_1113));
AOI21X1 g60565(.A0 (WX8629), .A1 (_2282_), .B0 (n_187), .Y (n_1112));
AOI21X1 g60566(.A0 (WX8625), .A1 (_2300_), .B0 (n_188), .Y (n_1111));
AOI21X1 g60567(.A0 (WX8623), .A1 (_2285_), .B0 (n_358), .Y (n_1110));
AOI21X1 g60568(.A0 (WX8619), .A1 (_2287_), .B0 (n_197), .Y (n_1109));
AOI21X1 g60569(.A0 (WX8617), .A1 (_2288_), .B0 (n_298), .Y (n_1108));
AOI21X1 g60570(.A0 (WX8615), .A1 (_2289_), .B0 (n_226), .Y (n_1107));
AOI21X1 g60571(.A0 (WX8611), .A1 (_2291_), .B0 (n_403), .Y (n_1106));
AOI21X1 g60572(.A0 (WX4760), .A1 (_2181_), .B0 (n_258), .Y (n_1105));
AOI21X1 g60573(.A0 (WX8599), .A1 (_2297_), .B0 (n_293), .Y (n_1104));
AOI21X1 g60574(.A0 (WX8595), .A1 (_2299_), .B0 (n_330), .Y (n_1103));
AOI21X1 g60575(.A0 (WX9950), .A1 (_2332_), .B0 (n_241), .Y (n_1102));
AOI21X1 g60576(.A0 (WX9948), .A1 (_2301_), .B0 (n_333), .Y (n_1101));
AOI21X1 g60577(.A0 (WX9944), .A1 (_2303_), .B0 (n_207), .Y (n_1100));
AOI21X1 g60578(.A0 (WX9938), .A1 (_2306_), .B0 (n_375), .Y (n_1099));
AOI21X1 g60579(.A0 (WX3455), .A1 (_2155_), .B0 (n_175), .Y (n_1098));
AOI21X1 g60580(.A0 (WX9934), .A1 (_2308_), .B0 (n_337), .Y (n_1097));
AOI21X1 g60581(.A0 (WX9932), .A1 (_2309_), .B0 (n_411), .Y (n_1096));
AOI21X1 g60582(.A0 (WX4734), .A1 (_2194_), .B0 (n_327), .Y (n_1095));
AOI21X1 g60583(.A0 (WX9928), .A1 (_2332_), .B0 (n_305), .Y (n_1094));
AOI21X1 g60584(.A0 (WX9924), .A1 (_2313_), .B0 (n_342), .Y (n_1093));
AOI21X1 g60585(.A0 (WX9920), .A1 (_2315_), .B0 (n_378), .Y (n_1092));
AOI21X1 g60586(.A0 (WX9918), .A1 (_2332_), .B0 (n_282), .Y (n_1091));
AOI21X1 g60587(.A0 (WX9912), .A1 (_2319_), .B0 (n_236), .Y (n_1090));
AOI21X1 g60588(.A0 (WX9910), .A1 (_2320_), .B0 (n_204), .Y (n_1089));
AOI21X1 g60589(.A0 (WX9906), .A1 (_2322_), .B0 (n_361), .Y (n_1088));
AOI21X1 g60590(.A0 (WX9902), .A1 (_2324_), .B0 (n_390), .Y (n_1087));
AOI21X1 g60591(.A0 (WX9898), .A1 (_2326_), .B0 (n_193), .Y (n_1086));
AOI21X1 g60592(.A0 (WX9894), .A1 (_2328_), .B0 (n_379), .Y (n_1085));
AOI21X1 g60593(.A0 (WX11243), .A1 (_2364_), .B0 (n_158), .Y (n_1084));
AOI21X1 g60594(.A0 (WX11239), .A1 (_2334_), .B0 (n_310), .Y (n_1083));
AOI21X1 g60595(.A0 (WX11235), .A1 (_2364_), .B0 (n_294), .Y (n_1082));
AOI21X1 g60596(.A0 (WX11233), .A1 (_2337_), .B0 (n_303), .Y (n_1081));
AOI21X1 g60597(.A0 (WX11225), .A1 (_2341_), .B0 (n_296), .Y (n_1080));
AOI21X1 g60598(.A0 (WX11221), .A1 (_2364_), .B0 (n_208), .Y (n_1079));
AOI21X1 g60599(.A0 (WX11219), .A1 (_2344_), .B0 (n_467), .Y (n_1078));
AOI21X1 g60600(.A0 (WX11215), .A1 (_2346_), .B0 (n_343), .Y (n_1077));
AOI21X1 g60601(.A0 (WX11211), .A1 (_2364_), .B0 (n_371), .Y (n_1076));
AOI21X1 g60602(.A0 (WX11209), .A1 (_2349_), .B0 (n_160), .Y (n_1075));
AOI21X1 g60603(.A0 (WX11205), .A1 (_2351_), .B0 (n_174), .Y (n_1074));
AOI21X1 g60604(.A0 (WX11201), .A1 (_2353_), .B0 (n_260), .Y (n_1073));
AOI21X1 g60605(.A0 (WX11199), .A1 (_2354_), .B0 (n_320), .Y (n_1072));
AOI21X1 g60606(.A0 (WX11197), .A1 (_2355_), .B0 (n_346), .Y (n_1071));
AOI21X1 g60607(.A0 (WX11193), .A1 (_2357_), .B0 (n_442), .Y (n_1070));
AOI21X1 g60608(.A0 (WX11189), .A1 (_2359_), .B0 (n_352), .Y (n_1069));
AOI21X1 g60609(.A0 (WX3467), .A1 (_2149_), .B0 (n_155), .Y (n_1068));
AOI21X1 g60610(.A0 (WX2150), .A1 (_2129_), .B0 (n_360), .Y (n_1067));
AOI21X1 g60611(.A0 (WX4774), .A1 (_2174_), .B0 (n_381), .Y (n_1066));
AOI21X1 g60612(.A0 (WX7312), .A1 (_2262_), .B0 (n_165), .Y (n_1065));
AOI21X1 g60613(.A0 (WX9888), .A1 (_2331_), .B0 (n_413), .Y (n_1064));
AOI21X1 g60614(.A0 (WX9916), .A1 (_2317_), .B0 (n_259), .Y (n_1063));
AOI21X1 g60615(.A0 (WX7348), .A1 (_2244_), .B0 (n_348), .Y (n_1062));
AOI21X1 g60616(.A0 (WX6027), .A1 (_2226_), .B0 (n_335), .Y (n_1061));
AOI21X1 g60617(.A0 (WX2164), .A1 (_2122_), .B0 (n_383), .Y (n_1060));
AOI21X1 g60618(.A0 (WX2188), .A1 (_2110_), .B0 (n_152), .Y (n_1059));
AOI21X1 g60619(.A0 (WX2182), .A1 (_2113_), .B0 (n_149), .Y (n_1058));
AOI21X1 g60620(.A0 (WX3431), .A1 (_2167_), .B0 (n_364), .Y (n_1057));
AOI21X1 g60621(.A0 (WX3433), .A1 (_2166_), .B0 (n_368), .Y (n_1056));
AOI21X1 g60622(.A0 (WX7314), .A1 (_2261_), .B0 (n_159), .Y (n_1055));
AOI21X1 g60624(.A0 (WX7364), .A1 (_2268_), .B0 (n_186), .Y (n_1054));
AOI21X1 g60625(.A0 (WX7318), .A1 (_2259_), .B0 (n_351), .Y (n_1053));
AOI21X1 g60626(.A0 (WX11227), .A1 (_2340_), .B0 (n_363), .Y (n_1052));
AOI21X1 g60627(.A0 (WX9942), .A1 (_2332_), .B0 (n_287), .Y (n_1051));
AOI21X1 g60628(.A0 (WX9908), .A1 (_2321_), .B0 (n_336), .Y (n_1050));
AOI21X1 g60629(.A0 (WX8603), .A1 (_2295_), .B0 (n_292), .Y (n_1049));
AOI21X1 g60630(.A0 (WX9914), .A1 (_2318_), .B0 (n_312), .Y (n_1048));
AOI21X1 g60631(.A0 (WX3477), .A1 (_2172_), .B0 (n_201), .Y (n_1047));
AOI21X1 g60632(.A0 (WX7336), .A1 (_2250_), .B0 (n_191), .Y (n_1046));
AOI21X1 g60633(.A0 (WX2154), .A1 (_2127_), .B0 (n_297), .Y (n_1045));
AOI21X1 g60634(.A0 (WX4756), .A1 (_2204_), .B0 (n_478), .Y (n_1044));
AOI21X1 g60636(.A0 (WX11185), .A1 (_2361_), .B0 (n_168), .Y (n_1043));
AOI21X1 g60637(.A0 (WX9890), .A1 (_2330_), .B0 (n_404), .Y (n_1042));
AOI21X1 g60638(.A0 (WX11237), .A1 (_2335_), .B0 (n_143), .Y (n_1041));
AOI21X1 g60639(.A0 (WX8613), .A1 (_2290_), .B0 (n_319), .Y (n_1040));
AOI21X1 g60640(.A0 (WX8597), .A1 (_2298_), .B0 (n_345), .Y (n_1039));
NOR2X1 g58167(.A (_2107_), .B (WX837), .Y (n_1038));
AOI21X1 g60641(.A0 (WX6065), .A1 (_2207_), .B0 (n_398), .Y (n_1037));
AOI21X1 g60642(.A0 (WX6019), .A1 (_2230_), .B0 (n_137), .Y (n_1036));
AOI21X1 g60643(.A0 (WX7346), .A1 (_2245_), .B0 (n_323), .Y (n_1035));
AOI21X1 g60644(.A0 (WX6015), .A1 (_2232_), .B0 (n_424), .Y (n_1034));
AOI21X1 g60645(.A0 (WX6071), .A1 (_2236_), .B0 (n_344), .Y (n_1033));
AOI21X1 g60646(.A0 (WX4736), .A1 (_2193_), .B0 (n_367), .Y (n_1032));
AOI21X1 g60647(.A0 (WX2178), .A1 (_2115_), .B0 (n_466), .Y (n_1031));
AOI21X1 g60648(.A0 (WX2146), .A1 (_2131_), .B0 (n_255), .Y (n_1030));
AOI21X1 g60651(.A0 (WX2174), .A1 (_2117_), .B0 (n_219), .Y (n_1029));
AOI21X1 g60652(.A0 (WX11223), .A1 (_2342_), .B0 (n_311), .Y (n_1028));
AOI21X1 g60653(.A0 (WX7350), .A1 (_2243_), .B0 (n_290), .Y (n_1027));
AOI21X1 g60654(.A0 (WX2148), .A1 (_2130_), .B0 (n_214), .Y (n_1026));
AOI21X1 g60655(.A0 (WX6055), .A1 (_2212_), .B0 (n_490), .Y (n_1025));
AOI21X1 g60656(.A0 (WX4724), .A1 (_2199_), .B0 (n_190), .Y (n_1024));
AOI21X1 g60659(.A0 (WX2168), .A1 (_2120_), .B0 (n_183), .Y (n_1023));
AOI21X1 g60660(.A0 (WX2192), .A1 (_2140_), .B0 (n_161), .Y (n_1022));
AOI21X1 g60661(.A0 (WX9926), .A1 (_2312_), .B0 (n_370), .Y (n_1021));
AOI21X1 g60663(.A0 (WX9896), .A1 (_2327_), .B0 (n_458), .Y (n_1020));
AOI21X1 g60664(.A0 (WX6045), .A1 (_2217_), .B0 (n_388), .Y (n_1019));
AOI21X1 g60665(.A0 (WX6031), .A1 (_2224_), .B0 (n_321), .Y (n_1018));
AOI21X1 g60666(.A0 (WX4778), .A1 (_2204_), .B0 (n_340), .Y (n_1017));
AOI21X1 g60667(.A0 (WX11191), .A1 (_2358_), .B0 (n_144), .Y (n_1016));
AOI21X1 g60668(.A0 (WX11207), .A1 (_2350_), .B0 (n_210), .Y (n_1015));
AOI21X1 g60669(.A0 (WX2142), .A1 (_2133_), .B0 (n_338), .Y (n_1014));
AOI21X1 g60670(.A0 (WX9892), .A1 (_2329_), .B0 (n_359), .Y (n_1013));
AOI21X1 g60671(.A0 (WX7308), .A1 (_2264_), .B0 (n_286), .Y (n_1012));
CLKBUFX3 g63046(.A (n_1011), .Y (n_1305));
CLKBUFX3 g63041(.A (n_1011), .Y (n_1460));
INVX2 g63023(.A (n_1009), .Y (n_2988));
INVX2 g63024(.A (n_1009), .Y (n_2953));
INVX2 g63018(.A (n_1009), .Y (n_2775));
INVX2 g63012(.A (n_1009), .Y (n_2755));
OR2X1 g61310(.A (n_1006), .B (n_1000), .Y (n_1007));
OR2X1 g61311(.A (n_1004), .B (n_943), .Y (n_1005));
NAND2X1 g61312(.A (n_983), .B (n_1004), .Y (n_1003));
OR2X1 g61315(.A (n_1001), .B (n_1000), .Y (n_1002));
NAND2X1 g61316(.A (n_1001), .B (n_979), .Y (n_999));
OR2X1 g61318(.A (n_997), .B (n_1000), .Y (n_998));
OR2X1 g61320(.A (n_995), .B (n_972), .Y (n_996));
NAND2X1 g61321(.A (n_6511), .B (n_995), .Y (n_994));
OR2X1 g61324(.A (n_992), .B (n_7490), .Y (n_993));
OR2X1 g61325(.A (n_990), .B (n_7490), .Y (n_991));
OR2X1 g61326(.A (n_987), .B (n_7490), .Y (n_988));
OR2X1 g61327(.A (n_985), .B (n_966), .Y (n_986));
NAND2X1 g61328(.A (n_985), .B (n_983), .Y (n_984));
OR2X1 g61331(.A (n_981), .B (n_1000), .Y (n_982));
NAND2X1 g61332(.A (n_981), .B (n_979), .Y (n_980));
OR2X1 g61337(.A (n_977), .B (n_7490), .Y (n_6697));
OR2X1 g61340(.A (n_975), .B (n_943), .Y (n_976));
OR2X1 g61347(.A (n_973), .B (n_972), .Y (n_974));
NAND2X1 g61349(.A (n_970), .B (n_966), .Y (n_971));
OR2X1 g61351(.A (n_970), .B (n_943), .Y (n_969));
NAND2X1 g61352(.A (n_973), .B (n_966), .Y (n_967));
NAND2X1 g61358(.A (n_964), .B (n_966), .Y (n_965));
OR2X1 g61359(.A (n_962), .B (n_966), .Y (n_963));
NAND2X1 g61360(.A (n_962), .B (n_983), .Y (n_960));
OR2X1 g61363(.A (n_958), .B (n_966), .Y (n_959));
OR2X1 g61365(.A (n_956), .B (n_943), .Y (n_957));
NAND2X1 g61370(.A (n_975), .B (n_983), .Y (n_955));
OR2X1 g61371(.A (n_953), .B (n_6432), .Y (n_954));
OR2X1 g61373(.A (n_951), .B (n_943), .Y (n_952));
NAND2X1 g61374(.A (n_951), .B (n_983), .Y (n_950));
OR2X1 g61458(.A (n_948), .B (n_7490), .Y (n_949));
NAND2X1 g61459(.A (n_1006), .B (n_6432), .Y (n_947));
OR2X1 g61460(.A (n_944), .B (n_943), .Y (n_945));
NAND2X1 g61461(.A (n_944), .B (n_966), .Y (n_942));
NAND2X1 g61462(.A (n_940), .B (n_979), .Y (n_941));
OR2X1 g61464(.A (n_938), .B (n_972), .Y (n_939));
NAND2X1 g61465(.A (n_938), .B (n_966), .Y (n_937));
OR2X1 g61469(.A (n_935), .B (n_7490), .Y (n_6699));
NAND2X1 g61470(.A (n_935), .B (n_6433), .Y (n_6698));
OR2X1 g61473(.A (n_932), .B (n_943), .Y (n_933));
NAND2X1 g61474(.A (n_983), .B (n_932), .Y (n_931));
OR2X1 g61477(.A (n_929), .B (n_7490), .Y (n_930));
NAND2X1 g61478(.A (n_927), .B (n_979), .Y (n_928));
NAND2X1 g61479(.A (n_990), .B (n_979), .Y (n_926));
OR2X1 g61480(.A (n_924), .B (n_943), .Y (n_925));
OR2X1 g61481(.A (n_940), .B (n_7490), .Y (n_923));
NAND2X1 g61482(.A (n_924), .B (n_983), .Y (n_922));
OR2X1 g61486(.A (n_920), .B (n_7490), .Y (n_921));
NAND2X1 g61487(.A (n_920), .B (n_6433), .Y (n_919));
OR2X1 g61490(.A (n_964), .B (n_966), .Y (n_918));
NAND2X1 g61492(.A (n_977), .B (n_6433), .Y (n_6696));
NAND2X1 g61499(.A (n_929), .B (n_6433), .Y (n_916));
NAND2X1 g61500(.A (n_956), .B (n_966), .Y (n_915));
OR2X1 g61501(.A (n_913), .B (n_972), .Y (n_914));
NAND2X1 g61503(.A (n_913), .B (n_966), .Y (n_912));
NAND2X1 g61506(.A (n_992), .B (n_6433), .Y (n_911));
NAND2X1 g61508(.A (n_987), .B (n_979), .Y (n_910));
NAND2X1 g61509(.A (n_953), .B (n_6433), .Y (n_909));
NAND2X1 g61511(.A (n_997), .B (n_979), .Y (n_908));
NAND2X1 g61513(.A (n_958), .B (n_966), .Y (n_907));
OR2X1 g61516(.A (n_905), .B (n_7490), .Y (n_906));
NAND2X1 g61517(.A (n_948), .B (n_6433), .Y (n_904));
OR2X1 g61518(.A (n_927), .B (n_7490), .Y (n_903));
NAND2X1 g61519(.A (n_905), .B (n_6433), .Y (n_902));
NOR2X1 g61522(.A (_2083_), .B (WX885), .Y (n_901));
NOR2X1 g61543(.A (_2086_), .B (WX879), .Y (n_900));
NOR2X1 g61547(.A (_2089_), .B (WX873), .Y (n_899));
NOR2X1 g61549(.A (_2108_), .B (WX877), .Y (n_898));
NOR2X1 g61603(.A (_2100_), .B (WX851), .Y (n_897));
INVX2 g63013(.A (n_1009), .Y (n_2770));
NOR2X1 g61831(.A (_2077_), .B (WX897), .Y (n_896));
NOR2X1 g61940(.A (_2096_), .B (WX859), .Y (n_895));
NOR2X1 g61946(.A (_2090_), .B (WX871), .Y (n_894));
NOR2X1 g61979(.A (_2097_), .B (WX857), .Y (n_893));
NOR2X1 g62069(.A (_2088_), .B (WX875), .Y (n_892));
NOR2X1 g62083(.A (_2081_), .B (WX889), .Y (n_891));
NOR2X1 g62103(.A (_2093_), .B (WX865), .Y (n_890));
NOR2X1 g62146(.A (_2105_), .B (WX841), .Y (n_889));
NOR2X1 g62187(.A (_2102_), .B (WX847), .Y (n_888));
NOR2X1 g62214(.A (_2108_), .B (WX891), .Y (n_887));
NOR2X1 g62275(.A (_2103_), .B (WX845), .Y (n_886));
NOR2X1 g62282(.A (_2104_), .B (WX843), .Y (n_885));
NOR2X1 g62301(.A (_2082_), .B (WX887), .Y (n_884));
NOR2X1 g62304(.A (_2106_), .B (WX839), .Y (n_883));
NOR2X1 g62321(.A (_2108_), .B (WX899), .Y (n_882));
NOR2X1 g62337(.A (_2079_), .B (WX893), .Y (n_881));
NOR2X1 g62587(.A (_2099_), .B (WX853), .Y (n_879));
NOR2X1 g62623(.A (_2108_), .B (WX867), .Y (n_878));
NOR2X1 g62689(.A (_2091_), .B (WX869), .Y (n_877));
NOR2X1 g62707(.A (_2094_), .B (WX863), .Y (n_876));
NOR2X1 g62735(.A (_2098_), .B (WX855), .Y (n_875));
NOR2X1 g62751(.A (_2095_), .B (WX861), .Y (n_874));
NOR2X1 g62762(.A (_2101_), .B (WX849), .Y (n_873));
INVX2 g63011(.A (n_1009), .Y (n_2817));
INVX2 g63021(.A (n_1009), .Y (n_3089));
INVX2 g63027(.A (n_1009), .Y (n_2837));
INVX4 g63032(.A (n_880), .Y (n_2744));
INVX2 g63240(.A (n_6512), .Y (n_2986));
INVX1 g63241(.A (n_6512), .Y (n_2838));
INVX4 g63247(.A (n_9424), .Y (n_2795));
INVX4 g63252(.A (n_869), .Y (n_2813));
INVX4 g63253(.A (n_869), .Y (n_2815));
INVX4 g63259(.A (n_868), .Y (n_2716));
INVX4 g63261(.A (n_867), .Y (n_2829));
INVX4 g63263(.A (n_867), .Y (n_2798));
INVX4 g63266(.A (n_866), .Y (n_2935));
INVX4 g63267(.A (n_866), .Y (n_2776));
BUFX3 g63480(.A (n_2298), .Y (n_2246));
BUFX3 g63488(.A (n_2346), .Y (n_2198));
BUFX3 g63489(.A (n_2346), .Y (n_2333));
BUFX3 g63490(.A (n_2346), .Y (n_2223));
BUFX3 g63493(.A (n_2383), .Y (n_2251));
BUFX3 g63494(.A (n_2383), .Y (n_2400));
BUFX3 g63498(.A (n_2383), .Y (n_2218));
BUFX3 g63572(.A (n_2227), .Y (n_2371));
BUFX3 g63574(.A (n_2227), .Y (n_2527));
INVX2 g63592(.A (n_6429), .Y (n_1276));
INVX4 g63612(.A (n_2826), .Y (n_860));
INVX4 g63616(.A (n_2826), .Y (n_858));
INVX2 g63618(.A (n_2826), .Y (n_3031));
INVX8 g63632(.A (n_857), .Y (n_3021));
INVX4 g63646(.A (n_7482), .Y (n_3120));
INVX2 g63652(.A (n_853), .Y (n_3027));
INVX2 g63666(.A (n_7482), .Y (n_1281));
NOR2X1 g61730(.A (_2084_), .B (WX883), .Y (n_852));
INVX4 g63258(.A (n_868), .Y (n_2809));
INVX2 g63248(.A (n_9425), .Y (n_2828));
AOI21X1 g57864(.A0 (WX2066), .A1 (WX2130), .B0 (n_472), .Y (n_850));
AOI21X1 g57865(.A0 (WX11117), .A1 (WX11181), .B0 (n_473), .Y (n_849));
XOR2X1 g57866(.A (n_108), .B (WX2130), .Y (n_848));
XOR2X1 g57870(.A (n_124), .B (WX11181), .Y (n_847));
NOR2X1 g62111(.A (_2085_), .B (WX881), .Y (n_846));
INVX8 g63621(.A (n_857), .Y (n_3137));
INVX4 g63229(.A (n_842), .Y (n_1278));
INVX4 g63222(.A (n_6623), .Y (n_2757));
INVX4 g63598(.A (n_836), .Y (n_1294));
BUFX3 g63571(.A (n_2227), .Y (n_2272));
INVX4 g63581(.A (n_836), .Y (n_3140));
BUFX3 g63573(.A (n_2227), .Y (n_2325));
BUFX3 g63575(.A (n_2227), .Y (n_2529));
BUFX3 g63569(.A (n_2227), .Y (n_2339));
BUFX3 g63570(.A (n_2227), .Y (n_2388));
BUFX3 g63563(.A (n_2227), .Y (n_2396));
BUFX3 g63560(.A (n_2227), .Y (n_2311));
BUFX3 g63561(.A (n_2227), .Y (n_2402));
INVX4 g63516(.A (n_3188), .Y (n_2378));
INVX4 g63501(.A (n_3188), .Y (n_2383));
XOR2X1 g60976(.A (WX8543), .B (WX8607), .Y (n_831));
NAND2X1 g58180(.A (n_0), .B (WX837), .Y (n_830));
INVX8 g63359(.A (n_823), .Y (n_1648));
NAND2X1 g58181(.A (WX773), .B (n_139), .Y (n_817));
INVX2 g63270(.A (n_517), .Y (n_866));
XOR2X1 g60706(.A (WX8583), .B (WX8647), .Y (n_816));
XOR2X1 g60708(.A (WX4668), .B (WX4732), .Y (n_815));
XOR2X1 g60713(.A (WX8587), .B (WX8651), .Y (n_814));
XOR2X1 g60714(.A (WX2068), .B (WX2132), .Y (n_813));
XOR2X1 g60715(.A (WX4670), .B (WX4734), .Y (n_812));
XOR2X1 g60717(.A (WX8589), .B (WX8653), .Y (n_811));
XOR2X1 g60721(.A (WX4672), .B (WX4736), .Y (n_810));
XOR2X1 g60723(.A (WX8593), .B (WX8657), .Y (n_809));
XOR2X1 g60732(.A (WX8541), .B (WX8605), .Y (n_808));
XOR2X1 g60736(.A (WX4680), .B (WX4744), .Y (n_807));
XOR2X1 g60740(.A (WX4684), .B (WX4748), .Y (n_806));
XOR2X1 g60742(.A (WX4686), .B (WX4750), .Y (n_805));
XOR2X1 g60749(.A (WX9824), .B (WX9888), .Y (n_804));
XOR2X1 g60750(.A (WX4682), .B (WX4746), .Y (n_803));
XOR2X1 g60752(.A (WX4714), .B (WX4778), .Y (n_802));
XOR2X1 g60753(.A (WX9826), .B (WX9890), .Y (n_801));
XOR2X1 g60756(.A (WX4690), .B (WX4754), .Y (n_800));
XOR2X1 g60759(.A (WX9828), .B (WX9892), .Y (n_799));
XOR2X1 g60762(.A (WX9830), .B (WX9894), .Y (n_798));
XOR2X1 g60763(.A (WX5999), .B (WX6063), .Y (n_797));
INVX2 g63047(.A (n_520), .Y (n_1011));
XOR2X1 g60767(.A (WX4692), .B (WX4756), .Y (n_796));
XOR2X1 g60768(.A (WX9832), .B (WX9896), .Y (n_795));
XOR2X1 g60771(.A (WX9834), .B (WX9898), .Y (n_794));
XOR2X1 g60772(.A (WX9858), .B (WX9922), .Y (n_793));
XOR2X1 g60775(.A (WX4694), .B (WX4758), .Y (n_792));
XOR2X1 g60777(.A (WX9836), .B (WX9900), .Y (n_791));
XOR2X1 g60783(.A (WX9840), .B (WX9904), .Y (n_790));
XOR2X1 g60790(.A (WX9848), .B (WX9912), .Y (n_789));
XOR2X1 g60791(.A (WX3387), .B (WX3451), .Y (n_788));
XOR2X1 g60792(.A (WX3359), .B (WX3423), .Y (n_787));
XOR2X1 g60794(.A (WX9850), .B (WX9914), .Y (n_786));
XOR2X1 g60798(.A (WX4702), .B (WX4766), .Y (n_785));
XOR2X1 g60799(.A (WX9852), .B (WX9916), .Y (n_784));
XOR2X1 g60806(.A (WX9856), .B (WX9920), .Y (n_783));
XOR2X1 g60809(.A (WX5955), .B (WX6019), .Y (n_782));
XOR2X1 g60812(.A (WX4706), .B (WX4770), .Y (n_781));
XOR2X1 g60814(.A (WX9860), .B (WX9924), .Y (n_780));
XOR2X1 g60815(.A (WX4708), .B (WX4772), .Y (n_779));
XOR2X1 g60817(.A (WX9864), .B (WX9928), .Y (n_778));
XOR2X1 g60824(.A (WX9868), .B (WX9932), .Y (n_777));
XOR2X1 g60836(.A (WX9874), .B (WX9938), .Y (n_776));
XOR2X1 g60839(.A (WX3363), .B (WX3427), .Y (n_775));
XOR2X1 g60841(.A (WX9876), .B (WX9940), .Y (n_774));
XOR2X1 g60844(.A (WX4704), .B (WX4768), .Y (n_773));
XOR2X1 g60845(.A (WX11119), .B (WX11183), .Y (n_772));
NAND2X1 g61520(.A (n_129), .B (WX897), .Y (n_771));
XOR2X1 g60847(.A (WX4674), .B (WX4738), .Y (n_770));
XOR2X1 g60851(.A (WX9880), .B (WX9944), .Y (n_768));
XOR2X1 g60852(.A (WX2070), .B (WX2134), .Y (n_767));
XOR2X1 g60855(.A (WX11131), .B (WX11195), .Y (n_766));
XOR2X1 g60858(.A (WX9884), .B (WX9948), .Y (n_765));
XOR2X1 g60859(.A (WX8537), .B (WX8601), .Y (n_764));
XOR2X1 g61033(.A (WX7248), .B (WX7312), .Y (n_763));
XOR2X1 g60869(.A (WX3367), .B (WX3431), .Y (n_762));
XOR2X1 g60870(.A (WX2096), .B (WX2160), .Y (n_761));
XOR2X1 g60871(.A (WX6005), .B (WX6069), .Y (n_760));
XOR2X1 g60873(.A (WX5977), .B (WX6041), .Y (n_759));
XOR2X1 g60876(.A (WX3369), .B (WX3433), .Y (n_758));
XOR2X1 g60878(.A (WX9854), .B (WX9918), .Y (n_757));
XOR2X1 g60879(.A (WX5945), .B (WX6009), .Y (n_756));
XOR2X1 g60881(.A (WX9878), .B (WX9942), .Y (n_755));
XOR2X1 g60882(.A (WX2074), .B (WX2138), .Y (n_754));
XOR2X1 g60883(.A (WX2076), .B (WX2140), .Y (n_753));
XOR2X1 g60886(.A (WX5947), .B (WX6011), .Y (n_752));
XOR2X1 g60887(.A (WX6001), .B (WX6065), .Y (n_751));
XOR2X1 g60892(.A (WX11125), .B (WX11189), .Y (n_750));
XOR2X1 g60893(.A (WX5949), .B (WX6013), .Y (n_749));
XOR2X1 g60894(.A (WX3371), .B (WX3435), .Y (n_748));
XOR2X1 g60895(.A (WX2088), .B (WX2152), .Y (n_747));
XOR2X1 g60898(.A (WX5951), .B (WX6015), .Y (n_746));
XOR2X1 g60901(.A (WX2078), .B (WX2142), .Y (n_745));
INVX4 g63020(.A (n_769), .Y (n_1009));
XOR2X1 g60913(.A (WX9862), .B (WX9926), .Y (n_744));
XOR2X1 g60914(.A (WX5959), .B (WX6023), .Y (n_743));
XOR2X1 g60915(.A (WX3373), .B (WX3437), .Y (n_742));
XOR2X1 g60917(.A (WX5965), .B (WX6029), .Y (n_741));
XOR2X1 g60919(.A (WX5993), .B (WX6057), .Y (n_740));
XOR2X1 g60921(.A (WX5967), .B (WX6031), .Y (n_739));
XOR2X1 g60927(.A (WX3377), .B (WX3441), .Y (n_738));
XOR2X1 g60928(.A (WX5973), .B (WX6037), .Y (n_737));
XOR2X1 g60930(.A (WX4696), .B (WX4760), .Y (n_736));
XOR2X1 g60931(.A (WX8533), .B (WX8597), .Y (n_735));
XOR2X1 g60934(.A (WX3389), .B (WX3453), .Y (n_734));
XOR2X1 g60935(.A (WX3379), .B (WX3443), .Y (n_733));
XOR2X1 g60937(.A (WX5981), .B (WX6045), .Y (n_732));
XOR2X1 g60939(.A (WX5971), .B (WX6035), .Y (n_731));
XOR2X1 g60940(.A (WX11133), .B (WX11197), .Y (n_730));
XOR2X1 g60941(.A (WX5983), .B (WX6047), .Y (n_729));
XOR2X1 g60942(.A (WX7284), .B (WX7348), .Y (n_728));
XOR2X1 g60943(.A (WX3381), .B (WX3445), .Y (n_727));
XOR2X1 g60947(.A (WX2090), .B (WX2154), .Y (n_726));
XOR2X1 g60949(.A (WX5991), .B (WX6055), .Y (n_725));
XOR2X1 g60956(.A (WX3385), .B (WX3449), .Y (n_724));
XOR2X1 g60961(.A (WX11123), .B (WX11187), .Y (n_723));
XOR2X1 g60963(.A (WX11135), .B (WX11199), .Y (n_722));
XOR2X1 g60969(.A (WX6003), .B (WX6067), .Y (n_721));
XOR2X1 g60977(.A (WX5985), .B (WX6049), .Y (n_720));
XOR2X1 g60979(.A (WX11141), .B (WX11205), .Y (n_719));
XOR2X1 g60982(.A (WX2098), .B (WX2162), .Y (n_718));
XOR2X1 g60984(.A (WX2100), .B (WX2164), .Y (n_717));
XOR2X1 g60985(.A (WX11171), .B (WX11235), .Y (n_716));
XOR2X1 g60986(.A (WX5961), .B (WX6025), .Y (n_715));
XOR2X1 g60987(.A (WX11143), .B (WX11207), .Y (n_714));
XOR2X1 g60990(.A (WX3393), .B (WX3457), .Y (n_713));
XOR2X1 g60997(.A (WX2102), .B (WX2166), .Y (n_712));
XOR2X1 g61005(.A (WX7238), .B (WX7302), .Y (n_711));
XOR2X1 g61006(.A (WX11145), .B (WX11209), .Y (n_710));
XOR2X1 g61007(.A (WX3395), .B (WX3459), .Y (n_709));
XOR2X1 g61015(.A (WX7242), .B (WX7306), .Y (n_708));
XOR2X1 g61016(.A (WX3397), .B (WX3461), .Y (n_707));
XOR2X1 g61017(.A (WX3375), .B (WX3439), .Y (n_706));
XOR2X1 g61019(.A (WX7244), .B (WX7308), .Y (n_705));
XOR2X1 g61025(.A (WX2104), .B (WX2168), .Y (n_704));
XOR2X1 g61027(.A (WX7246), .B (WX7310), .Y (n_703));
XOR2X1 g61028(.A (WX5957), .B (WX6021), .Y (n_702));
XOR2X1 g61029(.A (WX11147), .B (WX11211), .Y (n_701));
XOR2X1 g61030(.A (WX11129), .B (WX11193), .Y (n_700));
XOR2X1 g61036(.A (WX3399), .B (WX3463), .Y (n_699));
XOR2X1 g61038(.A (WX7250), .B (WX7314), .Y (n_698));
XOR2X1 g61042(.A (WX2106), .B (WX2170), .Y (n_697));
XOR2X1 g61043(.A (WX7252), .B (WX7316), .Y (n_696));
XOR2X1 g61047(.A (WX7254), .B (WX7318), .Y (n_695));
XOR2X1 g61050(.A (WX11149), .B (WX11213), .Y (n_693));
XOR2X1 g61052(.A (WX2108), .B (WX2172), .Y (n_692));
XOR2X1 g61054(.A (WX2072), .B (WX2136), .Y (n_691));
XOR2X1 g61055(.A (WX7256), .B (WX7320), .Y (n_690));
XOR2X1 g61064(.A (WX3401), .B (WX3465), .Y (n_689));
XOR2X1 g61065(.A (WX4712), .B (WX4776), .Y (n_688));
XOR2X1 g61066(.A (WX3417), .B (WX3481), .Y (n_687));
XOR2X1 g61074(.A (WX7262), .B (WX7326), .Y (n_686));
XOR2X1 g61075(.A (WX11151), .B (WX11215), .Y (n_685));
XOR2X1 g61078(.A (WX7264), .B (WX7328), .Y (n_684));
XOR2X1 g61079(.A (WX4666), .B (WX4730), .Y (n_683));
XOR2X1 g61081(.A (WX2110), .B (WX2174), .Y (n_682));
XOR2X1 g61085(.A (WX7266), .B (WX7330), .Y (n_681));
XOR2X1 g61090(.A (WX2112), .B (WX2176), .Y (n_680));
XOR2X1 g61093(.A (WX8579), .B (WX8643), .Y (n_679));
XOR2X1 g61096(.A (WX7270), .B (WX7334), .Y (n_678));
XOR2X1 g61098(.A (WX11153), .B (WX11217), .Y (n_677));
XOR2X1 g61100(.A (WX3405), .B (WX3469), .Y (n_676));
XOR2X1 g61101(.A (WX7272), .B (WX7336), .Y (n_675));
XOR2X1 g61102(.A (WX9870), .B (WX9934), .Y (n_674));
XOR2X1 g61107(.A (WX3407), .B (WX3471), .Y (n_673));
XOR2X1 g61109(.A (WX7276), .B (WX7340), .Y (n_672));
XOR2X1 g61110(.A (WX5953), .B (WX6017), .Y (n_671));
XOR2X1 g61111(.A (WX9846), .B (WX9910), .Y (n_670));
XOR2X1 g61114(.A (WX7278), .B (WX7342), .Y (n_669));
XOR2X1 g61116(.A (WX2114), .B (WX2178), .Y (n_668));
XOR2X1 g61118(.A (WX2084), .B (WX2148), .Y (n_667));
XOR2X1 g61119(.A (WX7280), .B (WX7344), .Y (n_666));
XOR2X1 g61120(.A (WX11155), .B (WX11219), .Y (n_665));
XOR2X1 g61124(.A (WX2116), .B (WX2180), .Y (n_664));
XOR2X1 g61125(.A (WX7282), .B (WX7346), .Y (n_663));
XOR2X1 g61128(.A (WX3409), .B (WX3473), .Y (n_662));
XOR2X1 g61130(.A (WX7286), .B (WX7350), .Y (n_661));
XOR2X1 g61135(.A (WX7288), .B (WX7352), .Y (n_660));
XOR2X1 g61136(.A (WX11157), .B (WX11221), .Y (n_659));
XOR2X1 g61137(.A (WX2118), .B (WX2182), .Y (n_658));
XOR2X1 g61141(.A (WX7290), .B (WX7354), .Y (n_657));
XOR2X1 g61000(.A (WX2124), .B (WX2188), .Y (n_656));
XOR2X1 g61143(.A (WX3411), .B (WX3475), .Y (n_655));
XOR2X1 g61148(.A (WX7294), .B (WX7358), .Y (n_654));
XOR2X1 g61153(.A (WX3413), .B (WX3477), .Y (n_653));
XOR2X1 g61155(.A (WX7296), .B (WX7360), .Y (n_652));
XOR2X1 g61158(.A (WX11159), .B (WX11223), .Y (n_651));
XOR2X1 g61159(.A (WX11127), .B (WX11191), .Y (n_650));
XOR2X1 g61162(.A (WX7298), .B (WX7362), .Y (n_649));
XOR2X1 g61163(.A (WX2120), .B (WX2184), .Y (n_648));
XOR2X1 g61164(.A (WX5975), .B (WX6039), .Y (n_647));
XOR2X1 g61165(.A (WX8575), .B (WX8639), .Y (n_646));
XOR2X1 g61168(.A (WX7300), .B (WX7364), .Y (n_645));
XOR2X1 g61172(.A (WX2122), .B (WX2186), .Y (n_644));
XOR2X1 g61174(.A (WX9844), .B (WX9908), .Y (n_643));
XOR2X1 g61175(.A (WX3415), .B (WX3479), .Y (n_642));
XOR2X1 g61176(.A (WX11161), .B (WX11225), .Y (n_641));
XOR2X1 g61181(.A (WX2126), .B (WX2190), .Y (n_640));
XOR2X1 g61186(.A (WX3419), .B (WX3483), .Y (n_639));
XOR2X1 g61191(.A (WX3421), .B (WX3485), .Y (n_638));
XOR2X1 g61198(.A (WX4710), .B (WX4774), .Y (n_637));
XOR2X1 g61199(.A (WX11167), .B (WX11231), .Y (n_636));
XOR2X1 g61203(.A (WX11169), .B (WX11233), .Y (n_635));
XOR2X1 g61204(.A (WX4662), .B (WX4726), .Y (n_634));
XOR2X1 g61205(.A (WX5979), .B (WX6043), .Y (n_633));
XOR2X1 g61207(.A (WX2086), .B (WX2150), .Y (n_632));
XOR2X1 g61210(.A (WX9866), .B (WX9930), .Y (n_631));
XOR2X1 g61211(.A (WX8531), .B (WX8595), .Y (n_630));
XOR2X1 g61216(.A (WX8535), .B (WX8599), .Y (n_629));
XOR2X1 g61217(.A (WX2082), .B (WX2146), .Y (n_628));
XOR2X1 g61222(.A (WX8539), .B (WX8603), .Y (n_627));
XOR2X1 g61223(.A (WX11173), .B (WX11237), .Y (n_626));
XOR2X1 g61224(.A (WX6007), .B (WX6071), .Y (n_625));
XOR2X1 g61231(.A (WX8571), .B (WX8635), .Y (n_624));
XOR2X1 g61232(.A (WX9842), .B (WX9906), .Y (n_623));
XOR2X1 g61235(.A (WX2094), .B (WX2158), .Y (n_622));
XOR2X1 g61236(.A (WX8545), .B (WX8609), .Y (n_621));
XOR2X1 g61241(.A (WX8547), .B (WX8611), .Y (n_620));
XOR2X1 g61242(.A (WX9838), .B (WX9902), .Y (n_619));
XOR2X1 g61243(.A (WX11175), .B (WX11239), .Y (n_618));
XOR2X1 g61245(.A (WX8549), .B (WX8613), .Y (n_617));
XOR2X1 g61250(.A (WX8551), .B (WX8615), .Y (n_616));
XOR2X1 g61251(.A (WX4652), .B (WX4716), .Y (n_615));
XOR2X1 g61260(.A (WX8555), .B (WX8619), .Y (n_614));
XOR2X1 g61264(.A (WX11177), .B (WX11241), .Y (n_613));
XOR2X1 g61267(.A (WX8557), .B (WX8621), .Y (n_612));
XOR2X1 g61268(.A (WX3391), .B (WX3455), .Y (n_611));
XOR2X1 g61273(.A (WX4656), .B (WX4720), .Y (n_610));
XOR2X1 g61275(.A (WX8561), .B (WX8625), .Y (n_609));
XOR2X1 g61280(.A (WX8563), .B (WX8627), .Y (n_608));
XOR2X1 g61281(.A (WX4658), .B (WX4722), .Y (n_607));
XOR2X1 g61282(.A (WX11179), .B (WX11243), .Y (n_606));
XOR2X1 g61289(.A (WX8567), .B (WX8631), .Y (n_605));
XOR2X1 g61290(.A (WX4660), .B (WX4724), .Y (n_604));
XOR2X1 g61297(.A (WX8573), .B (WX8637), .Y (n_603));
XOR2X1 g61298(.A (WX3383), .B (WX3447), .Y (n_602));
XOR2X1 g61301(.A (WX4664), .B (WX4728), .Y (n_601));
XOR2X1 g61302(.A (WX8577), .B (WX8641), .Y (n_600));
XOR2X1 g61303(.A (WX9886), .B (WX9950), .Y (n_599));
XOR2X1 g61309(.A (WX8581), .B (WX8645), .Y (n_598));
NAND2X1 g61313(.A (WX817), .B (n_261), .Y (n_597));
NAND2X1 g61314(.A (n_70), .B (WX881), .Y (n_596));
NAND2X1 g61317(.A (n_69), .B (WX887), .Y (n_595));
NAND2X1 g61319(.A (n_24), .B (WX847), .Y (n_594));
NAND2X1 g61322(.A (WX819), .B (n_484), .Y (n_593));
NAND2X1 g61323(.A (n_79), .B (WX859), .Y (n_592));
NAND2X1 g61329(.A (WX801), .B (n_462), .Y (n_591));
NAND2X1 g61330(.A (n_130), .B (WX885), .Y (n_590));
NAND2X1 g61333(.A (WX795), .B (n_280), .Y (n_589));
NAND2X1 g61334(.A (WX783), .B (n_252), .Y (n_588));
NAND2X1 g61335(.A (WX823), .B (n_266), .Y (n_587));
NAND2X1 g61338(.A (n_117), .B (WX867), .Y (n_586));
NAND2X1 g61339(.A (WX829), .B (n_451), .Y (n_585));
NAND2X1 g61342(.A (WX825), .B (n_268), .Y (n_584));
NAND2X1 g61343(.A (n_98), .B (WX849), .Y (n_583));
NAND2X1 g61344(.A (WX785), .B (n_420), .Y (n_582));
NAND2X1 g61345(.A (WX799), .B (n_438), .Y (n_581));
NAND2X1 g61346(.A (n_3), .B (WX889), .Y (n_580));
NAND2X1 g61348(.A (n_89), .B (WX861), .Y (n_579));
NAND2X1 g61354(.A (WX827), .B (n_448), .Y (n_578));
NAND2X1 g61355(.A (n_81), .B (WX841), .Y (n_577));
NAND2X1 g61356(.A (n_58), .B (WX891), .Y (n_576));
NAND2X1 g61357(.A (WX777), .B (n_273), .Y (n_575));
NAND2X1 g61361(.A (n_68), .B (WX893), .Y (n_574));
NAND2X1 g61362(.A (n_96), .B (WX883), .Y (n_573));
NAND2X1 g61364(.A (WX835), .B (n_480), .Y (n_572));
NAND2X1 g61366(.A (n_28), .B (WX865), .Y (n_571));
NAND2X1 g61367(.A (WX831), .B (n_278), .Y (n_570));
NAND2X1 g61368(.A (n_5), .B (WX895), .Y (n_569));
NAND2X1 g61369(.A (WX821), .B (n_482), .Y (n_568));
NAND2X1 g61372(.A (n_83), .B (WX839), .Y (n_567));
NAND2X1 g61375(.A (n_41), .B (WX843), .Y (n_566));
NAND2X1 g61463(.A (WX787), .B (n_454), .Y (n_565));
NAND2X1 g61466(.A (WX805), .B (n_474), .Y (n_564));
NAND2X1 g61467(.A (n_118), .B (WX869), .Y (n_563));
NAND2X1 g61471(.A (WX789), .B (n_264), .Y (n_562));
NAND2X1 g61472(.A (WX797), .B (n_244), .Y (n_561));
NAND2X1 g61475(.A (n_27), .B (WX853), .Y (n_560));
NAND2X1 g61476(.A (WX807), .B (n_283), .Y (n_559));
NAND2X1 g61483(.A (WX809), .B (n_486), .Y (n_558));
NAND2X1 g61484(.A (WX781), .B (n_308), .Y (n_557));
NAND2X1 g61485(.A (n_33), .B (WX873), .Y (n_556));
NAND2X1 g61488(.A (n_40), .B (WX845), .Y (n_555));
NAND2X1 g61489(.A (WX791), .B (n_434), .Y (n_554));
NAND2X1 g61491(.A (n_35), .B (WX855), .Y (n_553));
NAND2X1 g61493(.A (WX811), .B (n_429), .Y (n_552));
NAND2X1 g61494(.A (WX779), .B (n_436), .Y (n_551));
NAND2X1 g61495(.A (n_126), .B (WX899), .Y (n_550));
NAND2X1 g61496(.A (n_21), .B (WX875), .Y (n_549));
NAND2X1 g61497(.A (WX833), .B (n_443), .Y (n_548));
NAND2X1 g61498(.A (n_119), .B (WX871), .Y (n_547));
NAND2X1 g61502(.A (WX803), .B (n_476), .Y (n_546));
NAND2X1 g61504(.A (WX813), .B (n_271), .Y (n_545));
NAND2X1 g61505(.A (n_49), .B (WX877), .Y (n_544));
NAND2X1 g61507(.A (n_73), .B (WX879), .Y (n_543));
NAND2X1 g61510(.A (n_56), .B (WX851), .Y (n_542));
NAND2X1 g61512(.A (WX793), .B (n_354), .Y (n_541));
NAND2X1 g61514(.A (WX815), .B (n_431), .Y (n_540));
NAND2X1 g61515(.A (n_38), .B (WX857), .Y (n_539));
XOR2X1 g60972(.A (WX8585), .B (WX8649), .Y (n_538));
XOR2X1 g60959(.A (WX2092), .B (WX2156), .Y (n_537));
XOR2X1 g60955(.A (WX5995), .B (WX6059), .Y (n_536));
XOR2X1 g60923(.A (WX5969), .B (WX6033), .Y (n_535));
INVX4 g63483(.A (n_3188), .Y (n_2298));
XOR2X1 g60908(.A (WX2080), .B (WX2144), .Y (n_532));
XOR2X1 g60904(.A (WX5963), .B (WX6027), .Y (n_531));
XOR2X1 g60862(.A (WX11121), .B (WX11185), .Y (n_530));
XOR2X1 g60854(.A (WX9882), .B (WX9946), .Y (n_529));
XOR2X1 g60831(.A (WX9872), .B (WX9936), .Y (n_527));
XOR2X1 g60829(.A (WX5989), .B (WX6053), .Y (n_526));
XOR2X1 g60823(.A (WX3361), .B (WX3425), .Y (n_525));
NAND2X1 g61353(.A (n_36), .B (WX863), .Y (n_524));
NAND2X1 g61350(.A (WX775), .B (n_276), .Y (n_523));
XOR2X1 g60789(.A (WX4700), .B (WX4764), .Y (n_522));
XOR2X1 g60786(.A (WX4698), .B (WX4762), .Y (n_521));
CLKBUFX3 g63036(.A (n_520), .Y (n_880));
XOR2X1 g60760(.A (WX11139), .B (WX11203), .Y (n_519));
XOR2X1 g61306(.A (WX5987), .B (WX6051), .Y (n_518));
INVX2 g63255(.A (n_517), .Y (n_869));
XOR2X1 g61292(.A (WX8569), .B (WX8633), .Y (n_516));
XOR2X1 g60748(.A (WX4688), .B (WX4752), .Y (n_515));
XOR2X1 g61284(.A (WX8565), .B (WX8629), .Y (n_514));
INVX2 g63235(.A (n_943), .Y (n_842));
INVX2 g63260(.A (n_517), .Y (n_868));
INVX2 g63265(.A (n_517), .Y (n_867));
INVX8 g63418(.A (n_471), .Y (n_5712));
INVX4 g63492(.A (n_3188), .Y (n_2346));
XOR2X1 g61270(.A (WX8559), .B (WX8623), .Y (n_510));
XOR2X1 g61263(.A (WX4654), .B (WX4718), .Y (n_509));
XOR2X1 g60734(.A (WX4678), .B (WX4742), .Y (n_508));
XOR2X1 g60720(.A (WX8591), .B (WX8655), .Y (n_507));
XOR2X1 g61253(.A (WX8553), .B (WX8617), .Y (n_506));
INVX8 g63319(.A (n_471), .Y (n_5181));
XOR2X1 g61247(.A (WX5997), .B (WX6061), .Y (n_505));
XOR2X1 g61240(.A (WX11137), .B (WX11201), .Y (n_504));
INVX8 g63447(.A (n_471), .Y (n_1425));
XOR2X1 g61214(.A (WX3365), .B (WX3429), .Y (n_503));
XOR2X1 g61193(.A (WX2128), .B (WX2192), .Y (n_502));
XOR2X1 g61190(.A (WX11165), .B (WX11229), .Y (n_501));
XOR2X1 g61180(.A (WX11163), .B (WX11227), .Y (n_500));
XOR2X1 g61145(.A (WX7292), .B (WX7356), .Y (n_499));
INVX2 g63653(.A (n_7487), .Y (n_853));
XOR2X1 g61105(.A (WX7274), .B (WX7338), .Y (n_497));
INVX1 g63643(.A (n_7487), .Y (n_2800));
XOR2X1 g61089(.A (WX7268), .B (WX7332), .Y (n_496));
XOR2X1 g61073(.A (WX3403), .B (WX3467), .Y (n_495));
INVX4 g63630(.A (n_1000), .Y (n_857));
INVX4 g63604(.A (n_6431), .Y (n_836));
INVX8 g63619(.A (n_6432), .Y (n_2826));
XOR2X1 g61068(.A (WX7260), .B (WX7324), .Y (n_492));
INVX8 g63567(.A (n_3188), .Y (n_2227));
XOR2X1 g61061(.A (WX7258), .B (WX7322), .Y (n_491));
NOR2X1 g62558(.A (WX6055), .B (_2212_), .Y (n_490));
NOR2X1 g62559(.A (WX3473), .B (_2146_), .Y (n_489));
NOR2X1 g62095(.A (WX3459), .B (_2153_), .Y (n_488));
NOR2X1 g61590(.A (WX4728), .B (_2197_), .Y (n_479));
NOR2X1 g61538(.A (WX4756), .B (_2204_), .Y (n_478));
NOR2X1 g58179(.A (WX11117), .B (WX11181), .Y (n_473));
NOR2X1 g58178(.A (WX2066), .B (WX2130), .Y (n_472));
NOR2X1 g62750(.A (WX6043), .B (_2218_), .Y (n_470));
NOR2X1 g61574(.A (WX2184), .B (_2140_), .Y (n_469));
NOR2X1 g61575(.A (WX7328), .B (_2254_), .Y (n_468));
NOR2X1 g61576(.A (WX11219), .B (_2344_), .Y (n_467));
NOR2X1 g62049(.A (WX2178), .B (_2115_), .Y (n_466));
NOR2X1 g61569(.A (WX4720), .B (_2201_), .Y (n_465));
NOR2X1 g61560(.A (WX3475), .B (_2145_), .Y (n_464));
NOR2X1 g62029(.A (WX8621), .B (_2286_), .Y (n_461));
NOR2X1 g62591(.A (WX3429), .B (_2168_), .Y (n_460));
INVX2 g63048(.A (n_456), .Y (n_520));
NOR2X1 g61544(.A (WX9896), .B (_2327_), .Y (n_458));
NOR2X1 g61545(.A (WX3463), .B (_2172_), .Y (n_457));
CLKBUFX3 g63031(.A (n_456), .Y (n_769));
NOR2X1 g62040(.A (WX6047), .B (_2216_), .Y (n_453));
INVX4 g63009(.A (n_450), .Y (n_966));
NOR2X1 g62578(.A (WX8657), .B (_2300_), .Y (n_447));
NOR2X1 g62579(.A (WX11193), .B (_2357_), .Y (n_442));
NOR2X1 g62580(.A (WX8645), .B (_2274_), .Y (n_440));
NOR2X1 g62357(.A (WX7310), .B (_2263_), .Y (n_433));
NOR2X1 g61913(.A (WX9922), .B (_2314_), .Y (n_428));
NOR2X1 g62568(.A (WX3435), .B (_2165_), .Y (n_427));
NOR2X1 g61897(.A (WX8635), .B (_2300_), .Y (n_426));
NOR2X1 g62522(.A (WX6015), .B (_2232_), .Y (n_424));
NOR2X1 g61534(.A (WX3461), .B (_2152_), .Y (n_423));
NOR2X1 g61536(.A (WX4746), .B (_2204_), .Y (n_422));
NOR2X1 g61567(.A (WX7302), .B (_2267_), .Y (n_419));
NOR2X1 g62561(.A (WX6017), .B (_2231_), .Y (n_418));
NOR2X1 g62071(.A (WX8647), .B (_2273_), .Y (n_417));
NOR2X1 g61602(.A (WX7322), .B (_2257_), .Y (n_416));
NOR2X1 g61525(.A (WX8643), .B (_2275_), .Y (n_415));
NOR2X1 g61635(.A (WX3457), .B (_2154_), .Y (n_414));
NOR2X1 g61637(.A (WX9888), .B (_2331_), .Y (n_413));
NOR2X1 g61645(.A (WX9936), .B (_2307_), .Y (n_412));
NOR2X1 g61651(.A (WX9932), .B (_2309_), .Y (n_411));
NOR2X1 g61659(.A (WX8609), .B (_2292_), .Y (n_410));
NOR2X1 g61669(.A (WX11183), .B (_2362_), .Y (n_409));
NOR2X1 g61674(.A (WX6025), .B (_2227_), .Y (n_408));
NOR2X1 g61695(.A (WX9946), .B (_2302_), .Y (n_407));
NOR2X1 g61709(.A (WX6057), .B (_2211_), .Y (n_406));
NOR2X1 g61710(.A (WX11187), .B (_2360_), .Y (n_405));
NOR2X1 g61713(.A (WX9890), .B (_2330_), .Y (n_404));
NOR2X1 g61722(.A (WX8611), .B (_2291_), .Y (n_403));
NOR2X1 g61726(.A (WX3483), .B (_2141_), .Y (n_402));
NOR2X1 g61742(.A (WX3481), .B (_2142_), .Y (n_401));
NOR2X1 g62538(.A (WX2180), .B (_2114_), .Y (n_399));
NOR2X1 g61782(.A (WX6065), .B (_2207_), .Y (n_398));
NOR2X1 g61785(.A (WX6053), .B (_2213_), .Y (n_397));
NOR2X1 g61788(.A (WX3449), .B (_2158_), .Y (n_396));
NOR2X1 g61789(.A (WX3439), .B (_2163_), .Y (n_395));
NOR2X1 g61792(.A (WX3423), .B (_2171_), .Y (n_394));
NOR2X1 g61804(.A (WX7332), .B (_2268_), .Y (n_393));
NOR2X1 g61824(.A (WX6035), .B (_2222_), .Y (n_392));
NOR2X1 g61830(.A (WX4772), .B (_2175_), .Y (n_391));
NOR2X1 g61836(.A (WX9902), .B (_2324_), .Y (n_390));
NOR2X1 g61842(.A (WX3445), .B (_2160_), .Y (n_389));
NOR2X1 g61845(.A (WX6045), .B (_2217_), .Y (n_388));
NOR2X1 g61860(.A (WX3427), .B (_2169_), .Y (n_387));
NOR2X1 g61876(.A (WX11229), .B (_2339_), .Y (n_386));
NOR2X1 g61882(.A (WX2176), .B (_2116_), .Y (n_385));
NOR2X1 g61885(.A (WX7338), .B (_2249_), .Y (n_384));
NOR2X1 g61888(.A (WX2164), .B (_2122_), .Y (n_383));
NOR2X1 g61896(.A (WX8651), .B (_2271_), .Y (n_382));
NOR2X1 g61903(.A (WX4774), .B (_2174_), .Y (n_381));
NOR2X1 g61909(.A (WX7306), .B (_2265_), .Y (n_380));
NOR2X1 g61911(.A (WX9894), .B (_2328_), .Y (n_379));
NOR2X1 g61916(.A (WX9920), .B (_2315_), .Y (n_378));
NOR2X1 g61918(.A (WX3469), .B (_2148_), .Y (n_377));
NOR2X1 g61922(.A (WX2190), .B (_2109_), .Y (n_376));
NOR2X1 g61923(.A (WX9938), .B (_2306_), .Y (n_375));
NOR2X1 g61679(.A (WX3465), .B (_2150_), .Y (n_374));
NOR2X1 g61942(.A (WX2136), .B (_2136_), .Y (n_373));
NOR2X1 g61954(.A (WX6029), .B (_2225_), .Y (n_372));
NOR2X1 g61975(.A (WX11211), .B (_2364_), .Y (n_371));
NOR2X1 g61977(.A (WX9926), .B (_2312_), .Y (n_370));
NOR2X1 g62006(.A (WX8649), .B (_2300_), .Y (n_369));
NOR2X1 g62028(.A (WX3433), .B (_2166_), .Y (n_368));
NOR2X1 g62031(.A (WX4736), .B (_2193_), .Y (n_367));
NOR2X1 g62032(.A (WX8637), .B (_2278_), .Y (n_366));
NOR2X1 g62035(.A (WX2156), .B (_2126_), .Y (n_365));
NOR2X1 g62037(.A (WX3431), .B (_2167_), .Y (n_364));
NOR2X1 g62039(.A (WX11227), .B (_2340_), .Y (n_363));
NOR2X1 g62053(.A (WX8607), .B (_2293_), .Y (n_362));
NOR2X1 g62054(.A (WX9906), .B (_2322_), .Y (n_361));
NOR2X1 g62056(.A (WX2150), .B (_2129_), .Y (n_360));
NOR2X1 g62070(.A (WX9892), .B (_2329_), .Y (n_359));
NOR2X1 g62079(.A (WX8623), .B (_2285_), .Y (n_358));
NOR2X1 g62093(.A (WX4726), .B (_2198_), .Y (n_357));
NOR2X1 g62105(.A (WX3453), .B (_2172_), .Y (n_356));
NOR2X1 g62109(.A (WX4730), .B (_2196_), .Y (n_353));
NOR2X1 g62115(.A (WX11189), .B (_2359_), .Y (n_352));
NOR2X1 g62125(.A (WX7318), .B (_2259_), .Y (n_351));
NOR2X1 g62134(.A (WX7344), .B (_2246_), .Y (n_350));
NOR2X1 g62141(.A (WX11195), .B (_2356_), .Y (n_349));
NOR2X1 g62147(.A (WX7348), .B (_2244_), .Y (n_348));
NOR2X1 g62152(.A (WX6039), .B (_2236_), .Y (n_347));
NOR2X1 g62154(.A (WX11197), .B (_2355_), .Y (n_346));
NOR2X1 g62157(.A (WX8597), .B (_2298_), .Y (n_345));
NOR2X1 g62159(.A (WX6071), .B (_2236_), .Y (n_344));
NOR2X1 g62170(.A (WX11215), .B (_2346_), .Y (n_343));
NOR2X1 g62192(.A (WX9924), .B (_2313_), .Y (n_342));
NOR2X1 g62198(.A (WX3441), .B (_2162_), .Y (n_341));
NOR2X1 g62204(.A (WX4778), .B (_2204_), .Y (n_340));
NOR2X1 g62212(.A (WX6011), .B (_2234_), .Y (n_339));
NOR2X1 g62216(.A (WX2142), .B (_2133_), .Y (n_338));
NOR2X1 g62217(.A (WX9934), .B (_2308_), .Y (n_337));
NOR2X1 g62227(.A (WX9908), .B (_2321_), .Y (n_336));
NOR2X1 g62232(.A (WX6027), .B (_2226_), .Y (n_335));
NOR2X1 g62234(.A (WX7304), .B (_2266_), .Y (n_334));
NOR2X1 g62239(.A (WX9948), .B (_2301_), .Y (n_333));
NOR2X1 g62242(.A (WX4732), .B (_2195_), .Y (n_332));
NOR2X1 g62246(.A (WX4722), .B (_2200_), .Y (n_331));
NOR2X1 g62251(.A (WX8595), .B (_2299_), .Y (n_330));
NOR2X1 g62254(.A (WX9904), .B (_2323_), .Y (n_329));
NOR2X1 g62266(.A (WX6069), .B (_2205_), .Y (n_328));
NOR2X1 g62271(.A (WX4734), .B (_2194_), .Y (n_327));
NOR2X1 g62273(.A (WX2166), .B (_2121_), .Y (n_326));
NOR2X1 g62278(.A (WX2152), .B (_2128_), .Y (n_325));
NOR2X1 g62292(.A (WX6041), .B (_2219_), .Y (n_324));
NOR2X1 g62300(.A (WX7346), .B (_2245_), .Y (n_323));
NOR2X1 g62302(.A (WX4752), .B (_2185_), .Y (n_322));
NOR2X1 g62310(.A (WX6031), .B (_2224_), .Y (n_321));
NOR2X1 g62323(.A (WX11199), .B (_2354_), .Y (n_320));
NOR2X1 g62328(.A (WX8613), .B (_2290_), .Y (n_319));
NOR2X1 g62339(.A (WX8627), .B (_2283_), .Y (n_318));
NOR2X1 g62343(.A (WX8605), .B (_2294_), .Y (n_317));
NOR2X1 g62346(.A (WX7354), .B (_2241_), .Y (n_316));
NOR2X1 g62351(.A (WX6067), .B (_2206_), .Y (n_315));
NOR2X1 g62352(.A (WX3479), .B (_2143_), .Y (n_314));
NOR2X1 g62358(.A (WX3471), .B (_2147_), .Y (n_313));
NOR2X1 g62360(.A (WX9914), .B (_2318_), .Y (n_312));
NOR2X1 g62361(.A (WX11223), .B (_2342_), .Y (n_311));
NOR2X1 g62525(.A (WX11239), .B (_2334_), .Y (n_310));
NOR2X1 g62508(.A (WX6049), .B (_2236_), .Y (n_307));
NOR2X1 g62507(.A (WX2160), .B (_2140_), .Y (n_306));
NOR2X1 g62505(.A (WX9928), .B (_2332_), .Y (n_305));
NOR2X1 g62476(.A (WX2140), .B (_2134_), .Y (n_304));
NOR2X1 g62479(.A (WX11233), .B (_2337_), .Y (n_303));
NOR2X1 g62506(.A (WX9930), .B (_2310_), .Y (n_302));
NOR2X1 g62575(.A (WX6037), .B (_2221_), .Y (n_301));
NOR2X1 g62583(.A (WX4716), .B (_2203_), .Y (n_300));
NOR2X1 g62590(.A (WX3443), .B (_2161_), .Y (n_299));
NOR2X1 g62592(.A (WX8617), .B (_2288_), .Y (n_298));
NOR2X1 g62611(.A (WX2154), .B (_2127_), .Y (n_297));
NOR2X1 g61548(.A (WX11225), .B (_2341_), .Y (n_296));
NOR2X1 g62631(.A (WX6023), .B (_2228_), .Y (n_295));
NOR2X1 g62634(.A (WX11235), .B (_2364_), .Y (n_294));
NOR2X1 g62654(.A (WX8599), .B (_2297_), .Y (n_293));
NOR2X1 g62691(.A (WX8603), .B (_2295_), .Y (n_292));
NOR2X1 g62695(.A (WX2186), .B (_2111_), .Y (n_291));
NOR2X1 g62477(.A (WX7350), .B (_2243_), .Y (n_290));
NOR2X1 g62705(.A (WX8655), .B (_2269_), .Y (n_289));
NOR2X1 g61941(.A (WX8639), .B (_2277_), .Y (n_288));
NOR2X1 g62712(.A (WX9942), .B (_2332_), .Y (n_287));
NOR2X1 g62727(.A (WX7308), .B (_2264_), .Y (n_286));
NOR2X1 g62739(.A (WX11213), .B (_2347_), .Y (n_285));
NOR2X1 g62754(.A (WX9918), .B (_2332_), .Y (n_282));
NOR2X1 g61910(.A (WX11201), .B (_2353_), .Y (n_260));
NOR2X1 g61912(.A (WX9916), .B (_2317_), .Y (n_259));
NOR2X1 g61908(.A (WX4760), .B (_2181_), .Y (n_258));
NOR2X1 g62375(.A (WX11231), .B (_2338_), .Y (n_257));
NOR2X1 g62524(.A (WX7330), .B (_2253_), .Y (n_256));
NOR2X1 g61899(.A (WX2146), .B (_2131_), .Y (n_255));
NOR2X1 g61898(.A (WX4750), .B (_2186_), .Y (n_254));
NOR2X1 g61889(.A (WX2134), .B (_2137_), .Y (n_247));
NOR2X1 g61872(.A (WX9950), .B (_2332_), .Y (n_241));
NOR2X1 g61857(.A (WX9912), .B (_2319_), .Y (n_236));
NOR2X1 g62347(.A (WX2158), .B (_2125_), .Y (n_235));
INVX2 g63272(.A (n_6510), .Y (n_983));
NOR2X1 g62764(.A (WX7320), .B (_2258_), .Y (n_233));
NOR2X1 g62340(.A (WX3437), .B (_2164_), .Y (n_232));
NOR2X1 g62765(.A (WX7352), .B (_2242_), .Y (n_231));
NOR2X1 g61852(.A (WX7324), .B (_2256_), .Y (n_230));
NOR2X1 g62757(.A (WX2132), .B (_2138_), .Y (n_229));
NOR2X1 g61846(.A (WX2170), .B (_2140_), .Y (n_228));
NOR2X1 g61841(.A (WX7362), .B (_2237_), .Y (n_227));
NOR2X1 g62752(.A (WX8615), .B (_2289_), .Y (n_226));
INVX2 g63271(.A (n_6510), .Y (n_517));
NOR2X1 g61833(.A (WX8633), .B (_2280_), .Y (n_225));
NOR2X1 g62527(.A (WX2174), .B (_2117_), .Y (n_219));
NOR2X1 g61821(.A (WX2148), .B (_2130_), .Y (n_214));
NOR2X1 g62743(.A (WX8641), .B (_2276_), .Y (n_213));
NOR2X1 g61815(.A (WX6063), .B (_2236_), .Y (n_212));
NOR2X1 g61814(.A (WX7358), .B (_2239_), .Y (n_211));
NOR2X1 g61991(.A (WX11207), .B (_2350_), .Y (n_210));
NOR2X1 g62293(.A (WX2162), .B (_2123_), .Y (n_209));
NOR2X1 g61793(.A (WX11221), .B (_2364_), .Y (n_208));
NOR2X1 g62740(.A (WX9944), .B (_2303_), .Y (n_207));
NOR2X1 g62287(.A (WX3451), .B (_2157_), .Y (n_206));
NOR2X1 g62734(.A (WX2144), .B (_2132_), .Y (n_205));
NOR2X1 g62736(.A (WX9910), .B (_2320_), .Y (n_204));
INVX2 g63273(.A (n_6510), .Y (n_972));
NOR2X1 g62732(.A (WX3477), .B (_2172_), .Y (n_201));
CLKBUFX1 g63401(.A (n_471), .Y (n_823));
NOR2X1 g62730(.A (WX6059), .B (_2210_), .Y (n_200));
NOR2X1 g62268(.A (WX4744), .B (_2189_), .Y (n_199));
NOR2X1 g62728(.A (WX4768), .B (_2177_), .Y (n_198));
NOR2X1 g62722(.A (WX8619), .B (_2287_), .Y (n_197));
NOR2X1 g62716(.A (WX7316), .B (_2260_), .Y (n_195));
NOR2X1 g62713(.A (WX11217), .B (_2345_), .Y (n_194));
NOR2X1 g61756(.A (WX9898), .B (_2326_), .Y (n_193));
NOR2X1 g62249(.A (WX4754), .B (_2184_), .Y (n_192));
NOR2X1 g62708(.A (WX7336), .B (_2250_), .Y (n_191));
NOR2X1 g62706(.A (WX4724), .B (_2199_), .Y (n_190));
NOR2X1 g61557(.A (WX4742), .B (_2190_), .Y (n_189));
NOR2X1 g61993(.A (WX8625), .B (_2300_), .Y (n_188));
NOR2X1 g62235(.A (WX8629), .B (_2282_), .Y (n_187));
NOR2X1 g62694(.A (WX7364), .B (_2268_), .Y (n_186));
NOR2X1 g62228(.A (WX2172), .B (_2118_), .Y (n_185));
NOR2X1 g62696(.A (WX4776), .B (_2173_), .Y (n_184));
NOR2X1 g62697(.A (WX2168), .B (_2120_), .Y (n_183));
NOR2X1 g61738(.A (WX8631), .B (_2281_), .Y (n_181));
NOR2X1 g62692(.A (WX7356), .B (_2268_), .Y (n_180));
NOR2X1 g62688(.A (WX4740), .B (_2191_), .Y (n_179));
NOR2X1 g62666(.A (WX6061), .B (_2209_), .Y (n_178));
NOR2X1 g62220(.A (WX7360), .B (_2238_), .Y (n_177));
NOR2X1 g61734(.A (WX3425), .B (_2170_), .Y (n_176));
NOR2X1 g62276(.A (WX3455), .B (_2155_), .Y (n_175));
NOR2X1 g62213(.A (WX11205), .B (_2351_), .Y (n_174));
NOR2X1 g62683(.A (WX4738), .B (_2192_), .Y (n_173));
NOR2X1 g61779(.A (WX6051), .B (_2214_), .Y (n_172));
NOR2X1 g61723(.A (WX3485), .B (_2172_), .Y (n_171));
NOR2X1 g62673(.A (WX3447), .B (_2159_), .Y (n_170));
NOR2X1 g61718(.A (WX4770), .B (_2204_), .Y (n_169));
NOR2X1 g62199(.A (WX11185), .B (_2361_), .Y (n_168));
NOR2X1 g61715(.A (WX7334), .B (_2251_), .Y (n_167));
NOR2X1 g62668(.A (WX6009), .B (_2235_), .Y (n_166));
NOR2X1 g61652(.A (WX7312), .B (_2262_), .Y (n_165));
NOR2X1 g61999(.A (WX6033), .B (_2223_), .Y (n_164));
NOR2X1 g62724(.A (WX4758), .B (_2182_), .Y (n_163));
NOR2X1 g62174(.A (WX4718), .B (_2202_), .Y (n_162));
NOR2X1 g62652(.A (WX2192), .B (_2140_), .Y (n_161));
NOR2X1 g62648(.A (WX11209), .B (_2349_), .Y (n_160));
NOR2X1 g62171(.A (WX7314), .B (_2261_), .Y (n_159));
NOR2X1 g62645(.A (WX11243), .B (_2364_), .Y (n_158));
NOR2X1 g62639(.A (WX7340), .B (_2248_), .Y (n_157));
NOR2X1 g62163(.A (WX6021), .B (_2229_), .Y (n_156));
NOR2X1 g61692(.A (WX3467), .B (_2149_), .Y (n_155));
NOR2X1 g62546(.A (WX4748), .B (_2187_), .Y (n_154));
NOR2X1 g61685(.A (WX11241), .B (_2333_), .Y (n_153));
NOR2X1 g61677(.A (WX2188), .B (_2110_), .Y (n_152));
NOR2X1 g61678(.A (WX11203), .B (_2352_), .Y (n_151));
NOR2X1 g61665(.A (WX7342), .B (_2268_), .Y (n_150));
NOR2X1 g61660(.A (WX2182), .B (_2113_), .Y (n_149));
NOR2X1 g62142(.A (WX7326), .B (_2255_), .Y (n_148));
NOR2X1 g61657(.A (WX8601), .B (_2296_), .Y (n_147));
INVX2 g63655(.A (n_7480), .Y (n_979));
NOR2X1 g62139(.A (WX8653), .B (_2270_), .Y (n_146));
INVX4 g63656(.A (n_7480), .Y (n_1000));
NOR2X1 g62619(.A (WX4766), .B (_2178_), .Y (n_145));
NOR2X1 g61646(.A (WX11191), .B (_2358_), .Y (n_144));
NOR2X1 g61643(.A (WX11237), .B (_2335_), .Y (n_143));
NOR2X1 g62628(.A (WX4764), .B (_2179_), .Y (n_142));
NOR2X1 g62123(.A (WX4762), .B (_2180_), .Y (n_141));
INVX4 g63238(.A (n_6622), .Y (n_943));
NOR2X1 g61628(.A (WX6019), .B (_2230_), .Y (n_137));
NOR2X1 g61622(.A (WX2138), .B (_2135_), .Y (n_136));
NOR2X1 g61614(.A (WX9900), .B (_2325_), .Y (n_135));
NOR2X1 g62616(.A (WX6013), .B (_2233_), .Y (n_133));
NOR2X1 g61604(.A (WX9940), .B (_2305_), .Y (n_131));
INVX1 g62887(.A (WX1940), .Y (n_1335));
INVX1 g62969(.A (WX821), .Y (n_130));
INVX1 g62946(.A (WX833), .Y (n_129));
INVX1 g63302(.A (WX845), .Y (n_308));
INVX1 g62856(.A (WX691), .Y (n_995));
INVX1 g62982(.A (WX1980), .Y (n_1288));
INVX1 g62817(.A (WX861), .Y (n_244));
INVX1 g62811(.A (WX863), .Y (n_438));
INVX1 g63579(.A (RESET), .Y (n_127));
INVX1 g62797(.A (WX899), .Y (n_480));
INVX1 g62845(.A (WX835), .Y (n_126));
INVX1 g63294(.A (WX677), .Y (n_938));
INVX1 g62824(.A (_2363_), .Y (n_124));
INVX1 g62967(.A (WX671), .Y (n_992));
INVX1 g62828(.A (WX1960), .Y (n_1320));
INVX1 g63297(.A (WX853), .Y (n_264));
INVX1 g62926(.A (WX659), .Y (n_940));
INVX2 g63049(.A (TM0), .Y (n_456));
INVX1 g62980(.A (WX1992), .Y (n_1437));
INVX1 g63002(.A (WX771), .Y (n_120));
INVX1 g62818(.A (WX699), .Y (n_973));
INVX1 g62771(.A (WX1952), .Y (n_1341));
INVX1 g63305(.A (WX807), .Y (n_119));
INVX1 g62833(.A (WX805), .Y (n_118));
INVX1 g63670(.A (WX803), .Y (n_117));
INVX1 g62908(.A (WX855), .Y (n_434));
INVX1 g62772(.A (WX765), .Y (n_113));
INVX1 g62829(.A (WX763), .Y (n_112));
INVX1 g62837(.A (WX759), .Y (n_111));
INVX1 g62800(.A (WX1950), .Y (n_1284));
INVX1 g62939(.A (WX731), .Y (n_109));
INVX1 g62949(.A (_2139_), .Y (n_108));
INVX1 g62985(.A (WX891), .Y (n_448));
INVX1 g63282(.A (WX1958), .Y (n_1419));
INVX1 g62974(.A (WX749), .Y (n_106));
INVX1 g62914(.A (WX723), .Y (n_105));
INVX1 g62891(.A (WX703), .Y (n_956));
INVX1 g62783(.A (WX725), .Y (n_104));
INVX1 g62781(.A (WX2000), .Y (n_2675));
INVX1 g63280(.A (WX729), .Y (n_101));
INVX1 g62954(.A (WX751), .Y (n_100));
INVX1 g63674(.A (WX1968), .Y (n_2825));
INVX1 g62894(.A (WX785), .Y (n_98));
INVX1 g62794(.A (WX839), .Y (n_276));
INVX1 g62857(.A (WX819), .Y (n_96));
INVX1 g60143(.A (WX709), .Y (n_95));
INVX1 g62938(.A (WX679), .Y (n_932));
INVX1 g62995(.A (WX897), .Y (n_443));
INVX1 g62973(.A (WX867), .Y (n_476));
INVX1 g62924(.A (WX705), .Y (n_951));
INVX1 g62879(.A (WX797), .Y (n_89));
INVX1 g63275(.A (WX1998), .Y (n_1451));
INVX1 g63307(.A (WX1944), .Y (n_1339));
INVX1 g62902(.A (WX665), .Y (n_953));
INVX1 g63308(.A (WX675), .Y (n_948));
INVX1 g62779(.A (WX895), .Y (n_278));
INVX1 g62978(.A (WX769), .Y (n_87));
INVX1 g62996(.A (WX767), .Y (n_85));
INVX1 g63298(.A (WX775), .Y (n_83));
INVX1 g62883(.A (WX673), .Y (n_987));
INVX1 g62898(.A (WX777), .Y (n_81));
INVX1 g62776(.A (WX859), .Y (n_280));
INVX1 g62780(.A (WX651), .Y (n_927));
INVX1 g62862(.A (WX663), .Y (n_920));
INVX1 g62847(.A (WX795), .Y (n_79));
INVX1 g62890(.A (WX847), .Y (n_252));
INVX1 g62945(.A (WX875), .Y (n_429));
INVX1 g62803(.A (WX1974), .Y (n_1348));
INVX1 g62988(.A (WX815), .Y (n_73));
INVX1 g62855(.A (WX647), .Y (n_997));
INVX1 g63293(.A (WX881), .Y (n_261));
INVX1 g62918(.A (WX715), .Y (n_71));
INVX1 g63675(.A (WX817), .Y (n_70));
INVX2 g63010(.A (TM0), .Y (n_450));
INVX1 g63279(.A (WX653), .Y (n_990));
INVX1 g62998(.A (WX1984), .Y (n_1282));
INVX1 g62962(.A (WX869), .Y (n_474));
INVX1 g62966(.A (WX1994), .Y (n_1429));
INVX1 g63303(.A (WX823), .Y (n_69));
INVX1 g62941(.A (WX829), .Y (n_68));
INVX1 g62897(.A (WX1982), .Y (n_1309));
INVX1 g62814(.A (WX701), .Y (n_962));
INVX1 g62788(.A (WX757), .Y (n_67));
INVX1 g62948(.A (WX655), .Y (n_905));
INVX1 g63311(.A (WX683), .Y (n_964));
INVX1 g62957(.A (WX1972), .Y (n_1431));
INVX1 g62968(.A (WX1942), .Y (n_1359));
INVX1 g62922(.A (WX711), .Y (n_65));
INVX1 g62808(.A (WX885), .Y (n_482));
INVX1 g63276(.A (WX713), .Y (n_63));
INVX1 g62896(.A (WX649), .Y (n_929));
INVX1 g62905(.A (WX865), .Y (n_462));
INVX1 g62882(.A (WX1964), .Y (n_1323));
INVX1 g62956(.A (WX1986), .Y (n_2691));
INVX1 g62901(.A (WX645), .Y (n_1006));
INVX1 g62839(.A (WX697), .Y (n_970));
INVX1 g62990(.A (WX667), .Y (n_1001));
BUFX3 g63456(.A (RESET), .Y (n_471));
INVX1 g62886(.A (WX873), .Y (n_486));
INVX1 g62892(.A (WX1954), .Y (n_1449));
INVX1 g62936(.A (WX827), .Y (n_58));
INVX1 g62927(.A (WX1966), .Y (n_1427));
CLKBUFX3 g63578(.A (RESET), .Y (n_1297));
INVX1 g62854(.A (WX689), .Y (n_1004));
INVX1 g63001(.A (WX893), .Y (n_451));
INVX1 g62881(.A (WX1988), .Y (n_1442));
INVX1 g62909(.A (WX787), .Y (n_56));
INVX1 g62866(.A (WX687), .Y (n_958));
INVX1 g62931(.A (WX727), .Y (n_52));
INVX1 g62878(.A (WX695), .Y (n_975));
INVX1 g62769(.A (WX733), .Y (n_51));
INVX1 g62925(.A (WX1956), .Y (n_1421));
INVX1 g62953(.A (WX851), .Y (n_454));
INVX1 g63289(.A (WX813), .Y (n_49));
INVX1 g62831(.A (WX737), .Y (n_48));
INVX1 g62798(.A (WX739), .Y (n_46));
INVX1 g62920(.A (WX745), .Y (n_44));
INVX1 g63006(.A (WX747), .Y (n_43));
INVX1 g62930(.A (WX843), .Y (n_436));
INVX1 g62900(.A (blif_reset_net), .Y (n_6171));
INVX1 g62827(.A (WX841), .Y (n_273));
INVX1 g62782(.A (WX1978), .Y (n_1374));
INVX1 g63679(.A (WX779), .Y (n_41));
INVX1 g62801(.A (WX781), .Y (n_40));
INVX1 g62790(.A (WX793), .Y (n_38));
INVX1 g62819(.A (WX799), .Y (n_36));
INVX1 g62785(.A (WX791), .Y (n_35));
INVX1 g62958(.A (WX809), .Y (n_33));
INVX1 g62981(.A (WX661), .Y (n_935));
INVX1 g62852(.A (WX761), .Y (n_32));
INVX1 g62836(.A (WX485), .Y (n_3599));
INVX1 g62844(.A (WX883), .Y (n_484));
INVX1 g63004(.A (WX801), .Y (n_28));
INVX1 g63309(.A (WX789), .Y (n_27));
INVX1 g62863(.A (WX783), .Y (n_24));
INVX1 g62965(.A (WX849), .Y (n_420));
INVX1 g62851(.A (WX877), .Y (n_271));
INVX1 g62787(.A (WX693), .Y (n_985));
INVX1 g62867(.A (WX811), .Y (n_21));
INVX1 g62986(.A (WX741), .Y (n_20));
INVX1 g62935(.A (WX879), .Y (n_431));
INVX1 g62822(.A (WX755), .Y (n_19));
INVX1 g63286(.A (WX753), .Y (n_18));
INVX1 g62917(.A (WX1962), .Y (n_1345));
INVX1 g62976(.A (WX743), .Y (n_16));
INVX1 g62872(.A (WX707), .Y (n_944));
INVX1 g62870(.A (WX735), .Y (n_14));
INVX1 g62950(.A (WX1990), .Y (n_1328));
INVX1 g63278(.A (WX1970), .Y (n_1350));
INVX1 g62821(.A (WX685), .Y (n_913));
INVX1 g62913(.A (WX857), .Y (n_354));
INVX1 g62812(.A (WX721), .Y (n_12));
INVX1 g62869(.A (WX669), .Y (n_981));
INVX1 g58184(.A (WX837), .Y (n_139));
INVX1 g63678(.A (WX657), .Y (n_977));
INVX1 g62873(.A (WX1946), .Y (n_1412));
INVX1 g63288(.A (WX1996), .Y (n_1318));
INVX1 g62877(.A (WX1976), .Y (n_1286));
INVX1 g63285(.A (WX871), .Y (n_283));
INVX1 g62893(.A (WX1948), .Y (n_1357));
INVX1 g62916(.A (WX681), .Y (n_924));
INVX1 g62840(.A (WX831), .Y (n_5));
INVX1 g62804(.A (WX719), .Y (n_4));
INVX1 g62865(.A (WX10989), .Y (n_1315));
INVX1 g62876(.A (WX887), .Y (n_266));
INVX1 g55946(.A (WX489), .Y (n_3685));
INVX1 g63672(.A (WX825), .Y (n_3));
INVX1 g62991(.A (WX717), .Y (n_2));
INVX1 g62861(.A (WX889), .Y (n_268));
INVX1 g63677(.A (WX1938), .Y (n_1337));
INVX1 g58623(.A (WX773), .Y (n_0));
XOR2X1 g24(.A (WX3319), .B (n_6424), .Y (n_6425));
XOR2X1 g25(.A (WX3255), .B (n_6423), .Y (n_6424));
INVX1 g29(.A (n_6422), .Y (n_6423));
INVX2 g30(.A (n_7487), .Y (n_6422));
CLKBUFX1 g26(.A (n_7487), .Y (n_6428));
INVX1 g27(.A (n_7487), .Y (n_6429));
INVX2 g3(.A (n_6430), .Y (n_6431));
INVX2 g4(.A (TM1), .Y (n_6430));
INVX4 g1(.A (n_6430), .Y (n_6432));
INVX2 g2(.A (n_6430), .Y (n_6433));
NOR2X1 g14(.A (n_6438), .B (WX10845), .Y (n_6439));
INVX1 g65498(.A (n_6437), .Y (n_6438));
INVX4 g65499(.A (n_6624), .Y (n_6437));
NOR3X1 g65504(.A (n_6446), .B (n_6449), .C (n_6450), .Y (n_6451));
INVX2 g46(.A (n_6624), .Y (n_6446));
NOR2X1 g65505(.A (n_6447), .B (n_6448), .Y (n_6449));
XOR2X1 g65506(.A (WX7240), .B (WX7304), .Y (n_6447));
XOR2X1 g65507(.A (WX7176), .B (n_3034), .Y (n_6448));
AND2X1 g65508(.A (n_6448), .B (n_6447), .Y (n_6450));
INVX4 g43(.A (n_6446), .Y (n_6452));
OAI21X1 g40(.A0 (n_6458), .A1 (n_3426), .B0 (n_6466), .Y (n_6467));
INVX1 g42(.A (n_6457), .Y (n_6458));
NAND2X1 g65509(.A (n_6455), .B (n_6456), .Y (n_6457));
NAND2X1 g52(.A (n_3222), .B (n_6454), .Y (n_6455));
INVX1 g57(.A (WX10865), .Y (n_6454));
NAND2X1 g46_dup(.A (n_4100), .B (n_3737), .Y (n_6456));
OR2X1 g41(.A (n_5535), .B (n_6465), .Y (n_6466));
AOI22X1 g44(.A0 (_2346_), .A1 (n_3835), .B0 (n_4670), .B1(DATA_0_13), .Y (n_6465));
INVX1 g45(.A (n_6468), .Y (n_6469));
NAND2X1 g65511(.A (n_4100), .B (n_3737), .Y (n_6468));
OAI21X1 g36(.A0 (n_6475), .A1 (n_6480), .B0 (n_6485), .Y (n_6486));
INVX1 g38(.A (n_6474), .Y (n_6475));
NAND2X1 g39(.A (n_6472), .B (n_6473), .Y (n_6474));
NAND2X1 g65512(.A (n_3225), .B (n_6471), .Y (n_6472));
INVX1 g54(.A (WX10875), .Y (n_6471));
NAND2X1 g42_dup(.A (n_4094), .B (n_3894), .Y (n_6473));
INVX1 g65514(.A (n_6479), .Y (n_6480));
CLKBUFX1 g65515(.A (n_6497), .Y (n_6479));
OR2X1 g37(.A (n_5439), .B (n_6484), .Y (n_6485));
CLKBUFX3 g65520(.A (n_7089), .Y (n_6482));
AOI22X1 g65522(.A0 (_2341_), .A1 (n_5873), .B0 (n_3828), .B1(DATA_0_8), .Y (n_6484));
INVX1 g65523(.A (n_6487), .Y (n_6488));
NAND2X1 g65524(.A (n_4094), .B (n_3894), .Y (n_6487));
OAI21X1 g35(.A0 (n_6495), .A1 (n_6480), .B0 (n_6504), .Y (n_6505));
INVX1 g65526(.A (n_6494), .Y (n_6495));
NAND2X1 g65527(.A (n_6492), .B (n_6493), .Y (n_6494));
NAND2X1 g65528(.A (n_3223), .B (n_6491), .Y (n_6492));
INVX1 g65530(.A (WX9542), .Y (n_6491));
NAND2X1 g41_dup(.A (n_4101), .B (n_4000), .Y (n_6493));
CLKBUFX3 g65534(.A (n_7086), .Y (n_6497));
OAI21X1 g65536(.A0 (n_4549), .A1 (n_6501), .B0 (n_6503), .Y (n_6504));
AND2X1 g65537(.A (n_4586), .B (_2329_), .Y (n_6501));
CLKBUFX3 g51(.A (n_7089), .Y (n_6503));
INVX1 g65540(.A (n_6507), .Y (n_6508));
NAND2X1 g65541(.A (n_4101), .B (n_4000), .Y (n_6507));
XOR2X1 g21(.A (WX7216), .B (n_6514), .Y (n_6515));
XOR2X1 g22(.A (WX7152), .B (n_6513), .Y (n_6514));
INVX2 g65543(.A (n_6512), .Y (n_6513));
INVX4 g65544(.A (n_6511), .Y (n_6512));
INVX2 g65545(.A (n_6510), .Y (n_6511));
INVX2 g65546(.A (TM0), .Y (n_6510));
NAND2X2 g19(.A (n_6520), .B (n_6523), .Y (n_6524));
NAND2X2 g20(.A (n_6555), .B (n_6519), .Y (n_6520));
OAI21X1 g65549(.A0 (n_5944), .A1 (n_5889), .B0 (n_5898), .Y (n_6519));
NAND2X1 g65550(.A (n_6521), .B (n_2922), .Y (n_6523));
INVX1 g65551(.A (n_4165), .Y (n_6521));
NAND2X2 g65554(.A (n_6529), .B (n_6532), .Y (n_6533));
NAND2X2 g65555(.A (n_6575), .B (n_6528), .Y (n_6529));
OAI21X1 g65557(.A0 (n_5727), .A1 (n_5889), .B0 (n_5671), .Y (n_6528));
NAND2X2 g65558(.A (n_6530), .B (n_2922), .Y (n_6532));
INVX1 g65559(.A (n_4157), .Y (n_6530));
NAND2X2 g65561(.A (n_6537), .B (n_6540), .Y (n_6541));
NAND2X2 g65562(.A (n_6575), .B (n_6536), .Y (n_6537));
OAI21X1 g65565(.A0 (n_5543), .A1 (n_5889), .B0 (n_5445), .Y (n_6536));
NAND2X2 g65566(.A (n_6538), .B (n_2922), .Y (n_6540));
INVX1 g65567(.A (n_4151), .Y (n_6538));
NAND2X2 g65569(.A (n_6545), .B (n_6548), .Y (n_6549));
NAND2X2 g65570(.A (n_6583), .B (n_6544), .Y (n_6545));
OAI21X1 g65572(.A0 (n_5164), .A1 (n_5889), .B0 (n_5065), .Y (n_6544));
NAND2X2 g65573(.A (n_6546), .B (n_2922), .Y (n_6548));
INVX1 g65574(.A (n_4142), .Y (n_6546));
MX2X1 g65576(.A (n_6551), .B (n_6550), .S0 (n_6552), .Y (n_6553));
INVX1 g65577(.A (n_6550), .Y (n_6551));
NAND2X1 g65578(.A (n_541), .B (n_539), .Y (n_6550));
MX2X1 g65579(.A (n_101), .B (WX729), .S0 (n_2421), .Y (n_6552));
NAND2X2 g65580(.A (n_6557), .B (n_6560), .Y (n_6561));
NAND2X2 g65581(.A (n_6555), .B (n_6556), .Y (n_6557));
CLKBUFX3 g65582(.A (n_6614), .Y (n_6555));
OAI21X1 g65584(.A0 (n_5903), .A1 (n_5889), .B0 (n_5848), .Y (n_6556));
NAND2X1 g65585(.A (n_6558), .B (n_2922), .Y (n_6560));
INVX1 g65586(.A (n_4163), .Y (n_6558));
MX2X1 g65595(.A (n_6571), .B (n_6570), .S0 (n_6572), .Y (n_6573));
INVX1 g65596(.A (n_6570), .Y (n_6571));
NAND2X1 g65597(.A (n_558), .B (n_556), .Y (n_6570));
MX2X1 g65598(.A (n_44), .B (WX745), .S0 (n_2440), .Y (n_6572));
NAND2X2 g65599(.A (n_6577), .B (n_6580), .Y (n_6581));
NAND2X2 g65600(.A (n_6575), .B (n_6576), .Y (n_6577));
CLKBUFX3 g65601(.A (n_6614), .Y (n_6575));
OAI21X1 g65602(.A0 (n_5612), .A1 (n_5889), .B0 (n_5539), .Y (n_6576));
NAND2X1 g65603(.A (n_6578), .B (n_6619), .Y (n_6580));
INVX1 g65604(.A (n_4153), .Y (n_6578));
NAND2X2 g65606(.A (n_6585), .B (n_6588), .Y (n_6589));
NAND2X2 g65607(.A (n_6583), .B (n_6584), .Y (n_6585));
CLKBUFX3 g65608(.A (n_6614), .Y (n_6583));
OAI21X1 g65610(.A0 (n_5450), .A1 (n_5889), .B0 (n_5355), .Y (n_6584));
NAND2X1 g65611(.A (n_6586), .B (n_6619), .Y (n_6588));
INVX1 g65612(.A (n_4148), .Y (n_6586));
MX2X1 g65621(.A (n_6599), .B (n_6598), .S0 (n_6600), .Y (n_6601));
INVX1 g65622(.A (n_6598), .Y (n_6599));
NAND2X1 g65623(.A (n_587), .B (n_595), .Y (n_6598));
MX2X1 g65624(.A (n_111), .B (WX759), .S0 (n_2488), .Y (n_6600));
MX2X1 g65632(.A (n_6611), .B (n_6610), .S0 (n_6612), .Y (n_6613));
INVX1 g65633(.A (n_6610), .Y (n_6611));
NAND2X1 g65634(.A (n_585), .B (n_574), .Y (n_6610));
MX2X1 g65635(.A (n_113), .B (WX765), .S0 (n_2434), .Y (n_6612));
NAND2X2 g65636(.A (n_6617), .B (n_6620), .Y (n_6621));
NAND2X2 g65637(.A (n_6615), .B (n_6616), .Y (n_6617));
CLKBUFX2 g65638(.A (n_6614), .Y (n_6615));
AND2X1 g23(.A (n_3140), .B (RESET), .Y (n_6614));
OAI21X1 g65639(.A0 (n_4863), .A1 (n_5889), .B0 (n_4655), .Y (n_6616));
NAND2X1 g65640(.A (n_6618), .B (n_6619), .Y (n_6620));
INVX1 g65641(.A (n_4136), .Y (n_6618));
INVX1 g65642(.A (n_4697), .Y (n_6619));
NOR3X1 g65643(.A (n_5873), .B (n_6630), .C (n_6631), .Y (n_6632));
INVX4 g65645(.A (n_6437), .Y (n_6626));
CLKBUFX3 g65647(.A (n_6623), .Y (n_6624));
CLKBUFX3 g65648(.A (n_6622), .Y (n_6623));
INVX2 g65649(.A (TM0), .Y (n_6622));
NOR2X1 g65650(.A (n_6628), .B (n_6629), .Y (n_6630));
XOR2X1 g65651(.A (WX4676), .B (WX4740), .Y (n_6628));
XOR2X1 g65652(.A (WX4612), .B (n_3149), .Y (n_6629));
AND2X1 g65653(.A (n_6629), .B (n_6628), .Y (n_6631));
INVX4 g65654(.A (n_5873), .Y (n_6633));
MX2X1 g65663(.A (n_6643), .B (n_6642), .S0 (n_6644), .Y (n_6645));
INVX1 g65664(.A (n_6642), .Y (n_6643));
NAND2X1 g65665(.A (n_589), .B (n_592), .Y (n_6642));
MX2X1 g65666(.A (n_109), .B (WX731), .S0 (n_2508), .Y (n_6644));
AND2X1 g65763(.A (n_4099), .B (n_6884), .Y (n_6885));
AND2X1 g58048_dup(.A (n_4099), .B (n_6884), .Y (n_6886));
MX2X1 g65840(.A (n_7060), .B (n_7059), .S0 (n_7061), .Y (n_7062));
INVX1 g65841(.A (n_7059), .Y (n_7060));
NAND2X1 g65842(.A (n_562), .B (n_560), .Y (n_7059));
MX2X1 g65843(.A (n_104), .B (WX725), .S0 (n_2457), .Y (n_7061));
MX2X1 g65844(.A (n_7064), .B (n_7063), .S0 (n_7065), .Y (n_7066));
INVX1 g65845(.A (n_7063), .Y (n_7064));
NAND2X1 g65846(.A (n_588), .B (n_594), .Y (n_7063));
MX2X1 g65847(.A (n_4), .B (WX719), .S0 (n_2409), .Y (n_7065));
MX2X1 g65848(.A (n_7068), .B (n_7067), .S0 (n_7069), .Y (n_7070));
INVX1 g65849(.A (n_7067), .Y (n_7068));
NAND2X1 g65850(.A (n_554), .B (n_553), .Y (n_7067));
MX2X1 g65851(.A (n_52), .B (WX727), .S0 (n_2439), .Y (n_7069));
MX2X1 g65852(.A (n_7072), .B (n_7071), .S0 (n_7073), .Y (n_7074));
INVX1 g65853(.A (n_7071), .Y (n_7072));
NAND2X1 g65854(.A (n_581), .B (n_524), .Y (n_7071));
MX2X1 g65855(.A (n_14), .B (WX735), .S0 (n_2419), .Y (n_7073));
MX2X1 g65856(.A (n_7076), .B (n_7075), .S0 (n_7077), .Y (n_7078));
INVX1 g65857(.A (n_7075), .Y (n_7076));
NAND2X1 g65858(.A (n_546), .B (n_586), .Y (n_7075));
MX2X1 g65859(.A (n_46), .B (WX739), .S0 (n_2481), .Y (n_7077));
MX2X1 g65860(.A (n_7080), .B (n_7079), .S0 (n_7081), .Y (n_7082));
INVX1 g65861(.A (n_7079), .Y (n_7080));
NAND2X1 g65862(.A (n_575), .B (n_577), .Y (n_7079));
MX2X1 g65863(.A (n_63), .B (WX713), .S0 (n_2431), .Y (n_7081));
OAI21X1 g65864(.A0 (n_7085), .A1 (n_7088), .B0 (n_7093), .Y (n_7094));
NOR2X1 g65865(.A (n_7083), .B (n_7084), .Y (n_7085));
NOR2X1 g65866(.A (WX10861), .B (n_5427), .Y (n_7083));
AND2X1 g65867(.A (n_3741), .B (n_6633), .Y (n_7084));
INVX8 g65868(.A (n_7087), .Y (n_7088));
CLKBUFX3 g65869(.A (n_7086), .Y (n_7087));
AND2X1 g65870(.A (RESET), .B (n_3140), .Y (n_7086));
OR2X1 g65871(.A (n_5841), .B (n_7092), .Y (n_7093));
CLKBUFX3 g49(.A (n_7089), .Y (n_7090));
NOR2X1 g50(.A (n_3140), .B (n_127), .Y (n_7089));
AOI22X1 g65872(.A0 (_2348_), .A1 (n_3835), .B0 (n_5968), .B1(DATA_0_15), .Y (n_7092));
XOR2X1 g66050(.A (WX8467), .B (n_7484), .Y (n_7485));
XOR2X1 g66051(.A (WX8403), .B (n_7483), .Y (n_7484));
INVX2 g66052(.A (n_7482), .Y (n_7483));
INVX4 g66053(.A (n_7481), .Y (n_7482));
INVX2 g66054(.A (n_7480), .Y (n_7481));
INVX4 g33(.A (TM1), .Y (n_7480));
INVX4 g66056(.A (n_7480), .Y (n_7487));
INVX1 g66057(.A (n_7483), .Y (n_7488));
INVX4 g66059(.A (n_7480), .Y (n_7490));
AND2X1 g66953(.A (n_4017), .B (n_8314), .Y (n_9404));
AND2X1 g57917_dup(.A (n_4017), .B (n_8314), .Y (n_9405));
AND2X1 g66954(.A (n_4101), .B (n_8315), .Y (n_9406));
AND2X1 g58144_dup(.A (n_4101), .B (n_8315), .Y (n_9407));
AND2X1 g66955(.A (n_4099), .B (n_8316), .Y (n_9408));
AND2X1 g57947_dup(.A (n_4099), .B (n_8316), .Y (n_9409));
AND2X1 g66956(.A (n_4096), .B (n_8317), .Y (n_9410));
AND2X1 g57919_dup(.A (n_4096), .B (n_8317), .Y (n_9411));
AND2X1 g66957(.A (n_4017), .B (n_8318), .Y (n_9412));
AND2X1 g57941_dup(.A (n_4017), .B (n_8318), .Y (n_9413));
AND2X1 g66958(.A (n_4100), .B (n_8319), .Y (n_9414));
AND2X1 g58090_dup(.A (n_4100), .B (n_8319), .Y (n_9415));
AND2X1 g66959(.A (n_4106), .B (n_8321), .Y (n_9416));
AND2X1 g57967_dup(.A (n_4106), .B (n_8321), .Y (n_15867));
AND2X1 g66960(.A (n_4105), .B (n_8323), .Y (n_9418));
AND2X1 g57911_dup(.A (n_4105), .B (n_8323), .Y (n_9419));
AND2X1 g66961(.A (n_4103), .B (n_8324), .Y (n_9420));
AND2X1 g58008_dup(.A (n_4103), .B (n_8324), .Y (n_9421));
AND2X1 g66962(.A (n_6633), .B (n_8325), .Y (n_9422));
AND2X1 g58077_dup(.A (n_6633), .B (n_8325), .Y (n_9423));
CLKBUFX2 g66963(.A (n_6511), .Y (n_9424));
CLKBUFX1 g65547_dup(.A (n_6511), .Y (n_9425));
AND2X1 g66964(.A (n_4101), .B (n_8326), .Y (n_9426));
AND2X1 g58016_dup(.A (n_4101), .B (n_8326), .Y (n_9427));
AND2X1 g66965(.A (n_4103), .B (n_8327), .Y (n_9428));
AND2X1 g58150_dup(.A (n_4103), .B (n_8327), .Y (n_9429));
MX2X1 g66966(.A (n_9431), .B (n_9430), .S0 (n_9432), .Y (n_9433));
INVX1 g66967(.A (n_9430), .Y (n_9431));
NAND2X1 g66968(.A (n_817), .B (n_830), .Y (n_9430));
MX2X1 g66969(.A (n_95), .B (WX709), .S0 (n_2425), .Y (n_9432));
MX2X1 g66970(.A (n_9435), .B (n_9434), .S0 (n_9436), .Y (n_9437));
INVX1 g66971(.A (n_9434), .Y (n_9435));
NAND2X1 g66972(.A (n_572), .B (n_550), .Y (n_9434));
MX2X1 g66973(.A (n_120), .B (WX771), .S0 (n_2465), .Y (n_9436));
MX2X1 g67130(.A (n_9798), .B (n_9797), .S0 (n_9799), .Y (n_9800));
INVX1 g67131(.A (n_9797), .Y (n_9798));
NAND2X1 g67132(.A (n_591), .B (n_571), .Y (n_9797));
MX2X1 g67133(.A (n_48), .B (WX737), .S0 (n_2503), .Y (n_9799));
AND2X1 g67587(.A (n_4100), .B (n_8350), .Y (n_10712));
AND2X1 g58158_dup(.A (n_4100), .B (n_8350), .Y (n_10713));
AND2X1 g67588(.A (n_4095), .B (n_8351), .Y (n_10714));
AND2X1 g58100_dup(.A (n_4095), .B (n_8351), .Y (n_15863));
AND2X1 g67589(.A (n_4095), .B (n_8352), .Y (n_10716));
AND2X1 g58029_dup(.A (n_4095), .B (n_8352), .Y (n_10717));
AND2X1 g67590(.A (n_4106), .B (n_8353), .Y (n_10718));
AND2X1 g58099_dup(.A (n_4106), .B (n_8353), .Y (n_10719));
AND2X1 g67591(.A (n_6452), .B (n_8354), .Y (n_10720));
AND2X1 g58112_dup(.A (n_6452), .B (n_8354), .Y (n_10721));
AND2X1 g67592(.A (n_4104), .B (n_8355), .Y (n_10722));
AND2X1 g58036_dup(.A (n_4104), .B (n_8355), .Y (n_10723));
MX2X1 g67593(.A (n_10725), .B (n_10724), .S0 (n_10726), .Y (n_10727));
INVX1 g67594(.A (n_10724), .Y (n_10725));
NAND2X1 g67595(.A (n_565), .B (n_542), .Y (n_10724));
MX2X1 g67596(.A (n_105), .B (WX723), .S0 (n_2493), .Y (n_10726));
MX2X1 g67597(.A (n_10729), .B (n_10728), .S0 (n_10730), .Y (n_10731));
INVX1 g67598(.A (n_10728), .Y (n_10729));
NAND2X1 g67599(.A (n_561), .B (n_579), .Y (n_10728));
MX2X1 g67600(.A (n_51), .B (WX733), .S0 (n_2497), .Y (n_10730));
MX2X1 g67601(.A (n_10733), .B (n_10732), .S0 (n_10734), .Y (n_10735));
INVX1 g67602(.A (n_10732), .Y (n_10733));
NAND2X1 g67603(.A (n_552), .B (n_549), .Y (n_10732));
MX2X1 g67604(.A (n_43), .B (WX747), .S0 (n_2428), .Y (n_10734));
MX2X1 g67605(.A (n_10737), .B (n_10736), .S0 (n_10738), .Y (n_10739));
INVX1 g67606(.A (n_10736), .Y (n_10737));
NAND2X1 g67607(.A (n_540), .B (n_543), .Y (n_10736));
MX2X1 g67608(.A (n_100), .B (WX751), .S0 (n_2412), .Y (n_10738));
MX2X1 g67609(.A (n_10741), .B (n_10740), .S0 (n_10742), .Y (n_10743));
INVX1 g67610(.A (n_10740), .Y (n_10741));
NAND2X1 g67611(.A (n_584), .B (n_580), .Y (n_10740));
MX2X1 g67612(.A (n_32), .B (WX761), .S0 (n_2484), .Y (n_10742));
MX2X1 g67613(.A (n_10745), .B (n_10744), .S0 (n_10746), .Y (n_10747));
INVX1 g67614(.A (n_10744), .Y (n_10745));
NAND2X1 g67615(.A (n_523), .B (n_567), .Y (n_10744));
MX2X1 g67616(.A (n_65), .B (WX711), .S0 (n_2505), .Y (n_10746));
AND2X1 g68036(.A (n_4105), .B (n_9384), .Y (n_11595));
AND2X1 g57962_dup(.A (n_4105), .B (n_9384), .Y (n_11596));
AND2X1 g68037(.A (n_4099), .B (n_9385), .Y (n_11597));
AND2X1 g57951_dup(.A (n_4099), .B (n_9385), .Y (n_15865));
AND2X1 g68038(.A (n_4100), .B (n_9386), .Y (n_11599));
AND2X1 g58108_dup(.A (n_4100), .B (n_9386), .Y (n_11600));
AND2X1 g68039(.A (n_4094), .B (n_9387), .Y (n_11601));
AND2X1 g57968_dup(.A (n_4094), .B (n_9387), .Y (n_11602));
AND2X1 g68040(.A (n_4099), .B (n_9388), .Y (n_11603));
AND2X1 g58103_dup(.A (n_4099), .B (n_9388), .Y (n_11604));
AND2X1 g68041(.A (n_4017), .B (n_9389), .Y (n_11605));
AND2X1 g57918_dup(.A (n_4017), .B (n_9389), .Y (n_15855));
AND2X1 g68042(.A (n_6452), .B (n_9390), .Y (n_11607));
AND2X1 g58012_dup(.A (n_6452), .B (n_9390), .Y (n_11608));
AND2X1 g68043(.A (n_4094), .B (n_9391), .Y (n_11609));
AND2X1 g58146_dup(.A (n_4094), .B (n_9391), .Y (n_15857));
AND2X1 g68044(.A (n_6633), .B (n_9392), .Y (n_11611));
AND2X1 g58056_dup(.A (n_6633), .B (n_9392), .Y (n_11612));
AND2X1 g68045(.A (n_6452), .B (n_9393), .Y (n_11613));
AND2X1 g58148_dup(.A (n_6452), .B (n_9393), .Y (n_11614));
AND2X1 g68046(.A (n_4095), .B (n_9394), .Y (n_11615));
AND2X1 g58017_dup(.A (n_4095), .B (n_9394), .Y (n_11616));
AND2X1 g68047(.A (n_4096), .B (n_9395), .Y (n_11617));
AND2X1 g58088_dup(.A (n_4096), .B (n_9395), .Y (n_11618));
AND2X1 g68048(.A (n_4017), .B (n_9396), .Y (n_11619));
AND2X1 g57933_dup(.A (n_4017), .B (n_9396), .Y (n_15851));
AND2X1 g68049(.A (n_4103), .B (n_9397), .Y (n_11621));
AND2X1 g58094_dup(.A (n_4103), .B (n_9397), .Y (n_15859));
AND2X1 g68050(.A (n_4105), .B (n_9398), .Y (n_11623));
AND2X1 g57943_dup(.A (n_4105), .B (n_9398), .Y (n_15861));
AND2X1 g68051(.A (n_4094), .B (n_9399), .Y (n_11625));
AND2X1 g58096_dup(.A (n_4094), .B (n_9399), .Y (n_11626));
endmodule
