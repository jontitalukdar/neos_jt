
module keccak ( clk, reset, in, in_ready, is_last, byte_num, buffer_full, out, 
        out_ready );
  input [31:0] in;
  input [1:0] byte_num;
  output [511:0] out;
  input clk, reset, in_ready, is_last;
  output buffer_full, out_ready;
  wire   i_22_, state, f_ack, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         padder_out_ready, n4, n50, n900, n1000, n1100, n120, n130, n140, n150,
         n160, n170, n180, n190, n200, n210, n220, n230, n240, n250, n260,
         n270, n28, n29, n30, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n901, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n1001, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n1101, n111, n112, n113, n114, n115, n116,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414,
         SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416,
         SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418,
         SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420,
         SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422,
         SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424,
         SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426,
         SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428,
         SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430,
         SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432,
         SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434,
         SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436,
         SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438,
         SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440,
         SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442,
         SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444,
         SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446,
         SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448,
         SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450,
         SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452,
         SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454,
         SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456,
         SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458,
         SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460,
         SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462,
         SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464,
         SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466,
         SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468,
         SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470,
         SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472,
         SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474,
         SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476,
         SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478,
         SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480,
         SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482,
         SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484,
         SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486,
         SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488,
         SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490,
         SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492,
         SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494,
         SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496,
         SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498,
         SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500,
         SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502,
         SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504,
         SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506,
         SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508,
         SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510,
         SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512,
         SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514,
         SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516,
         SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518,
         SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520,
         SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522,
         SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524,
         SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526,
         SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528,
         SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530,
         SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532,
         SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534,
         SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536,
         SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538,
         SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540,
         SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542,
         SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544,
         SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546,
         SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548,
         SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550,
         SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552,
         SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554,
         SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556,
         SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558,
         SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560,
         SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562,
         SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564,
         SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566,
         SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568,
         SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570,
         SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572,
         SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574,
         SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576,
         SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578,
         SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580,
         SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582,
         SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584,
         SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586,
         SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588,
         SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590,
         SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592,
         SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594,
         SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596,
         SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598,
         SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600,
         SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602,
         SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604,
         SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606,
         SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608,
         SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610,
         SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612,
         SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614,
         SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616,
         SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618,
         SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620,
         SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622,
         SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624,
         SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626,
         SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628,
         SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630,
         SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632,
         SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634,
         SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636,
         SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638,
         SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640,
         SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642,
         SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644,
         SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646,
         SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648,
         SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650,
         SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652,
         SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654,
         SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656,
         SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658,
         SYNOPSYS_UNCONNECTED_659, SYNOPSYS_UNCONNECTED_660,
         SYNOPSYS_UNCONNECTED_661, SYNOPSYS_UNCONNECTED_662,
         SYNOPSYS_UNCONNECTED_663, SYNOPSYS_UNCONNECTED_664,
         SYNOPSYS_UNCONNECTED_665, SYNOPSYS_UNCONNECTED_666,
         SYNOPSYS_UNCONNECTED_667, SYNOPSYS_UNCONNECTED_668,
         SYNOPSYS_UNCONNECTED_669, SYNOPSYS_UNCONNECTED_670,
         SYNOPSYS_UNCONNECTED_671, SYNOPSYS_UNCONNECTED_672,
         SYNOPSYS_UNCONNECTED_673, SYNOPSYS_UNCONNECTED_674,
         SYNOPSYS_UNCONNECTED_675, SYNOPSYS_UNCONNECTED_676,
         SYNOPSYS_UNCONNECTED_677, SYNOPSYS_UNCONNECTED_678,
         SYNOPSYS_UNCONNECTED_679, SYNOPSYS_UNCONNECTED_680,
         SYNOPSYS_UNCONNECTED_681, SYNOPSYS_UNCONNECTED_682,
         SYNOPSYS_UNCONNECTED_683, SYNOPSYS_UNCONNECTED_684,
         SYNOPSYS_UNCONNECTED_685, SYNOPSYS_UNCONNECTED_686,
         SYNOPSYS_UNCONNECTED_687, SYNOPSYS_UNCONNECTED_688,
         SYNOPSYS_UNCONNECTED_689, SYNOPSYS_UNCONNECTED_690,
         SYNOPSYS_UNCONNECTED_691, SYNOPSYS_UNCONNECTED_692,
         SYNOPSYS_UNCONNECTED_693, SYNOPSYS_UNCONNECTED_694,
         SYNOPSYS_UNCONNECTED_695, SYNOPSYS_UNCONNECTED_696,
         SYNOPSYS_UNCONNECTED_697, SYNOPSYS_UNCONNECTED_698,
         SYNOPSYS_UNCONNECTED_699, SYNOPSYS_UNCONNECTED_700,
         SYNOPSYS_UNCONNECTED_701, SYNOPSYS_UNCONNECTED_702,
         SYNOPSYS_UNCONNECTED_703, SYNOPSYS_UNCONNECTED_704,
         SYNOPSYS_UNCONNECTED_705, SYNOPSYS_UNCONNECTED_706,
         SYNOPSYS_UNCONNECTED_707, SYNOPSYS_UNCONNECTED_708,
         SYNOPSYS_UNCONNECTED_709, SYNOPSYS_UNCONNECTED_710,
         SYNOPSYS_UNCONNECTED_711, SYNOPSYS_UNCONNECTED_712,
         SYNOPSYS_UNCONNECTED_713, SYNOPSYS_UNCONNECTED_714,
         SYNOPSYS_UNCONNECTED_715, SYNOPSYS_UNCONNECTED_716,
         SYNOPSYS_UNCONNECTED_717, SYNOPSYS_UNCONNECTED_718,
         SYNOPSYS_UNCONNECTED_719, SYNOPSYS_UNCONNECTED_720,
         SYNOPSYS_UNCONNECTED_721, SYNOPSYS_UNCONNECTED_722,
         SYNOPSYS_UNCONNECTED_723, SYNOPSYS_UNCONNECTED_724,
         SYNOPSYS_UNCONNECTED_725, SYNOPSYS_UNCONNECTED_726,
         SYNOPSYS_UNCONNECTED_727, SYNOPSYS_UNCONNECTED_728,
         SYNOPSYS_UNCONNECTED_729, SYNOPSYS_UNCONNECTED_730,
         SYNOPSYS_UNCONNECTED_731, SYNOPSYS_UNCONNECTED_732,
         SYNOPSYS_UNCONNECTED_733, SYNOPSYS_UNCONNECTED_734,
         SYNOPSYS_UNCONNECTED_735, SYNOPSYS_UNCONNECTED_736,
         SYNOPSYS_UNCONNECTED_737, SYNOPSYS_UNCONNECTED_738,
         SYNOPSYS_UNCONNECTED_739, SYNOPSYS_UNCONNECTED_740,
         SYNOPSYS_UNCONNECTED_741, SYNOPSYS_UNCONNECTED_742,
         SYNOPSYS_UNCONNECTED_743, SYNOPSYS_UNCONNECTED_744,
         SYNOPSYS_UNCONNECTED_745, SYNOPSYS_UNCONNECTED_746,
         SYNOPSYS_UNCONNECTED_747, SYNOPSYS_UNCONNECTED_748,
         SYNOPSYS_UNCONNECTED_749, SYNOPSYS_UNCONNECTED_750,
         SYNOPSYS_UNCONNECTED_751, SYNOPSYS_UNCONNECTED_752,
         SYNOPSYS_UNCONNECTED_753, SYNOPSYS_UNCONNECTED_754,
         SYNOPSYS_UNCONNECTED_755, SYNOPSYS_UNCONNECTED_756,
         SYNOPSYS_UNCONNECTED_757, SYNOPSYS_UNCONNECTED_758,
         SYNOPSYS_UNCONNECTED_759, SYNOPSYS_UNCONNECTED_760,
         SYNOPSYS_UNCONNECTED_761, SYNOPSYS_UNCONNECTED_762,
         SYNOPSYS_UNCONNECTED_763, SYNOPSYS_UNCONNECTED_764,
         SYNOPSYS_UNCONNECTED_765, SYNOPSYS_UNCONNECTED_766,
         SYNOPSYS_UNCONNECTED_767, SYNOPSYS_UNCONNECTED_768,
         SYNOPSYS_UNCONNECTED_769, SYNOPSYS_UNCONNECTED_770,
         SYNOPSYS_UNCONNECTED_771, SYNOPSYS_UNCONNECTED_772,
         SYNOPSYS_UNCONNECTED_773, SYNOPSYS_UNCONNECTED_774,
         SYNOPSYS_UNCONNECTED_775, SYNOPSYS_UNCONNECTED_776,
         SYNOPSYS_UNCONNECTED_777, SYNOPSYS_UNCONNECTED_778,
         SYNOPSYS_UNCONNECTED_779, SYNOPSYS_UNCONNECTED_780,
         SYNOPSYS_UNCONNECTED_781, SYNOPSYS_UNCONNECTED_782,
         SYNOPSYS_UNCONNECTED_783, SYNOPSYS_UNCONNECTED_784,
         SYNOPSYS_UNCONNECTED_785, SYNOPSYS_UNCONNECTED_786,
         SYNOPSYS_UNCONNECTED_787, SYNOPSYS_UNCONNECTED_788,
         SYNOPSYS_UNCONNECTED_789, SYNOPSYS_UNCONNECTED_790,
         SYNOPSYS_UNCONNECTED_791, SYNOPSYS_UNCONNECTED_792,
         SYNOPSYS_UNCONNECTED_793, SYNOPSYS_UNCONNECTED_794,
         SYNOPSYS_UNCONNECTED_795, SYNOPSYS_UNCONNECTED_796,
         SYNOPSYS_UNCONNECTED_797, SYNOPSYS_UNCONNECTED_798,
         SYNOPSYS_UNCONNECTED_799, SYNOPSYS_UNCONNECTED_800,
         SYNOPSYS_UNCONNECTED_801, SYNOPSYS_UNCONNECTED_802,
         SYNOPSYS_UNCONNECTED_803, SYNOPSYS_UNCONNECTED_804,
         SYNOPSYS_UNCONNECTED_805, SYNOPSYS_UNCONNECTED_806,
         SYNOPSYS_UNCONNECTED_807, SYNOPSYS_UNCONNECTED_808,
         SYNOPSYS_UNCONNECTED_809, SYNOPSYS_UNCONNECTED_810,
         SYNOPSYS_UNCONNECTED_811, SYNOPSYS_UNCONNECTED_812,
         SYNOPSYS_UNCONNECTED_813, SYNOPSYS_UNCONNECTED_814,
         SYNOPSYS_UNCONNECTED_815, SYNOPSYS_UNCONNECTED_816,
         SYNOPSYS_UNCONNECTED_817, SYNOPSYS_UNCONNECTED_818,
         SYNOPSYS_UNCONNECTED_819, SYNOPSYS_UNCONNECTED_820,
         SYNOPSYS_UNCONNECTED_821, SYNOPSYS_UNCONNECTED_822,
         SYNOPSYS_UNCONNECTED_823, SYNOPSYS_UNCONNECTED_824,
         SYNOPSYS_UNCONNECTED_825, SYNOPSYS_UNCONNECTED_826,
         SYNOPSYS_UNCONNECTED_827, SYNOPSYS_UNCONNECTED_828,
         SYNOPSYS_UNCONNECTED_829, SYNOPSYS_UNCONNECTED_830,
         SYNOPSYS_UNCONNECTED_831, SYNOPSYS_UNCONNECTED_832,
         SYNOPSYS_UNCONNECTED_833, SYNOPSYS_UNCONNECTED_834,
         SYNOPSYS_UNCONNECTED_835, SYNOPSYS_UNCONNECTED_836,
         SYNOPSYS_UNCONNECTED_837, SYNOPSYS_UNCONNECTED_838,
         SYNOPSYS_UNCONNECTED_839, SYNOPSYS_UNCONNECTED_840,
         SYNOPSYS_UNCONNECTED_841, SYNOPSYS_UNCONNECTED_842,
         SYNOPSYS_UNCONNECTED_843, SYNOPSYS_UNCONNECTED_844,
         SYNOPSYS_UNCONNECTED_845, SYNOPSYS_UNCONNECTED_846,
         SYNOPSYS_UNCONNECTED_847, SYNOPSYS_UNCONNECTED_848,
         SYNOPSYS_UNCONNECTED_849, SYNOPSYS_UNCONNECTED_850,
         SYNOPSYS_UNCONNECTED_851, SYNOPSYS_UNCONNECTED_852,
         SYNOPSYS_UNCONNECTED_853, SYNOPSYS_UNCONNECTED_854,
         SYNOPSYS_UNCONNECTED_855, SYNOPSYS_UNCONNECTED_856,
         SYNOPSYS_UNCONNECTED_857, SYNOPSYS_UNCONNECTED_858,
         SYNOPSYS_UNCONNECTED_859, SYNOPSYS_UNCONNECTED_860,
         SYNOPSYS_UNCONNECTED_861, SYNOPSYS_UNCONNECTED_862,
         SYNOPSYS_UNCONNECTED_863, SYNOPSYS_UNCONNECTED_864,
         SYNOPSYS_UNCONNECTED_865, SYNOPSYS_UNCONNECTED_866,
         SYNOPSYS_UNCONNECTED_867, SYNOPSYS_UNCONNECTED_868,
         SYNOPSYS_UNCONNECTED_869, SYNOPSYS_UNCONNECTED_870,
         SYNOPSYS_UNCONNECTED_871, SYNOPSYS_UNCONNECTED_872,
         SYNOPSYS_UNCONNECTED_873, SYNOPSYS_UNCONNECTED_874,
         SYNOPSYS_UNCONNECTED_875, SYNOPSYS_UNCONNECTED_876,
         SYNOPSYS_UNCONNECTED_877, SYNOPSYS_UNCONNECTED_878,
         SYNOPSYS_UNCONNECTED_879, SYNOPSYS_UNCONNECTED_880,
         SYNOPSYS_UNCONNECTED_881, SYNOPSYS_UNCONNECTED_882,
         SYNOPSYS_UNCONNECTED_883, SYNOPSYS_UNCONNECTED_884,
         SYNOPSYS_UNCONNECTED_885, SYNOPSYS_UNCONNECTED_886,
         SYNOPSYS_UNCONNECTED_887, SYNOPSYS_UNCONNECTED_888,
         SYNOPSYS_UNCONNECTED_889, SYNOPSYS_UNCONNECTED_890,
         SYNOPSYS_UNCONNECTED_891, SYNOPSYS_UNCONNECTED_892,
         SYNOPSYS_UNCONNECTED_893, SYNOPSYS_UNCONNECTED_894,
         SYNOPSYS_UNCONNECTED_895, SYNOPSYS_UNCONNECTED_896,
         SYNOPSYS_UNCONNECTED_897, SYNOPSYS_UNCONNECTED_898,
         SYNOPSYS_UNCONNECTED_899, SYNOPSYS_UNCONNECTED_900,
         SYNOPSYS_UNCONNECTED_901, SYNOPSYS_UNCONNECTED_902,
         SYNOPSYS_UNCONNECTED_903, SYNOPSYS_UNCONNECTED_904,
         SYNOPSYS_UNCONNECTED_905, SYNOPSYS_UNCONNECTED_906,
         SYNOPSYS_UNCONNECTED_907, SYNOPSYS_UNCONNECTED_908,
         SYNOPSYS_UNCONNECTED_909, SYNOPSYS_UNCONNECTED_910,
         SYNOPSYS_UNCONNECTED_911, SYNOPSYS_UNCONNECTED_912,
         SYNOPSYS_UNCONNECTED_913, SYNOPSYS_UNCONNECTED_914,
         SYNOPSYS_UNCONNECTED_915, SYNOPSYS_UNCONNECTED_916,
         SYNOPSYS_UNCONNECTED_917, SYNOPSYS_UNCONNECTED_918,
         SYNOPSYS_UNCONNECTED_919, SYNOPSYS_UNCONNECTED_920,
         SYNOPSYS_UNCONNECTED_921, SYNOPSYS_UNCONNECTED_922,
         SYNOPSYS_UNCONNECTED_923, SYNOPSYS_UNCONNECTED_924,
         SYNOPSYS_UNCONNECTED_925, SYNOPSYS_UNCONNECTED_926,
         SYNOPSYS_UNCONNECTED_927, SYNOPSYS_UNCONNECTED_928,
         SYNOPSYS_UNCONNECTED_929, SYNOPSYS_UNCONNECTED_930,
         SYNOPSYS_UNCONNECTED_931, SYNOPSYS_UNCONNECTED_932,
         SYNOPSYS_UNCONNECTED_933, SYNOPSYS_UNCONNECTED_934,
         SYNOPSYS_UNCONNECTED_935, SYNOPSYS_UNCONNECTED_936,
         SYNOPSYS_UNCONNECTED_937, SYNOPSYS_UNCONNECTED_938,
         SYNOPSYS_UNCONNECTED_939, SYNOPSYS_UNCONNECTED_940,
         SYNOPSYS_UNCONNECTED_941, SYNOPSYS_UNCONNECTED_942,
         SYNOPSYS_UNCONNECTED_943, SYNOPSYS_UNCONNECTED_944,
         SYNOPSYS_UNCONNECTED_945, SYNOPSYS_UNCONNECTED_946,
         SYNOPSYS_UNCONNECTED_947, SYNOPSYS_UNCONNECTED_948,
         SYNOPSYS_UNCONNECTED_949, SYNOPSYS_UNCONNECTED_950,
         SYNOPSYS_UNCONNECTED_951, SYNOPSYS_UNCONNECTED_952,
         SYNOPSYS_UNCONNECTED_953, SYNOPSYS_UNCONNECTED_954,
         SYNOPSYS_UNCONNECTED_955, SYNOPSYS_UNCONNECTED_956,
         SYNOPSYS_UNCONNECTED_957, SYNOPSYS_UNCONNECTED_958,
         SYNOPSYS_UNCONNECTED_959, SYNOPSYS_UNCONNECTED_960,
         SYNOPSYS_UNCONNECTED_961, SYNOPSYS_UNCONNECTED_962,
         SYNOPSYS_UNCONNECTED_963, SYNOPSYS_UNCONNECTED_964,
         SYNOPSYS_UNCONNECTED_965, SYNOPSYS_UNCONNECTED_966,
         SYNOPSYS_UNCONNECTED_967, SYNOPSYS_UNCONNECTED_968,
         SYNOPSYS_UNCONNECTED_969, SYNOPSYS_UNCONNECTED_970,
         SYNOPSYS_UNCONNECTED_971, SYNOPSYS_UNCONNECTED_972,
         SYNOPSYS_UNCONNECTED_973, SYNOPSYS_UNCONNECTED_974,
         SYNOPSYS_UNCONNECTED_975, SYNOPSYS_UNCONNECTED_976,
         SYNOPSYS_UNCONNECTED_977, SYNOPSYS_UNCONNECTED_978,
         SYNOPSYS_UNCONNECTED_979, SYNOPSYS_UNCONNECTED_980,
         SYNOPSYS_UNCONNECTED_981, SYNOPSYS_UNCONNECTED_982,
         SYNOPSYS_UNCONNECTED_983, SYNOPSYS_UNCONNECTED_984,
         SYNOPSYS_UNCONNECTED_985, SYNOPSYS_UNCONNECTED_986,
         SYNOPSYS_UNCONNECTED_987, SYNOPSYS_UNCONNECTED_988,
         SYNOPSYS_UNCONNECTED_989, SYNOPSYS_UNCONNECTED_990,
         SYNOPSYS_UNCONNECTED_991, SYNOPSYS_UNCONNECTED_992,
         SYNOPSYS_UNCONNECTED_993, SYNOPSYS_UNCONNECTED_994,
         SYNOPSYS_UNCONNECTED_995, SYNOPSYS_UNCONNECTED_996,
         SYNOPSYS_UNCONNECTED_997, SYNOPSYS_UNCONNECTED_998,
         SYNOPSYS_UNCONNECTED_999, SYNOPSYS_UNCONNECTED_1000,
         SYNOPSYS_UNCONNECTED_1001, SYNOPSYS_UNCONNECTED_1002,
         SYNOPSYS_UNCONNECTED_1003, SYNOPSYS_UNCONNECTED_1004,
         SYNOPSYS_UNCONNECTED_1005, SYNOPSYS_UNCONNECTED_1006,
         SYNOPSYS_UNCONNECTED_1007, SYNOPSYS_UNCONNECTED_1008,
         SYNOPSYS_UNCONNECTED_1009, SYNOPSYS_UNCONNECTED_1010,
         SYNOPSYS_UNCONNECTED_1011, SYNOPSYS_UNCONNECTED_1012,
         SYNOPSYS_UNCONNECTED_1013, SYNOPSYS_UNCONNECTED_1014,
         SYNOPSYS_UNCONNECTED_1015, SYNOPSYS_UNCONNECTED_1016,
         SYNOPSYS_UNCONNECTED_1017, SYNOPSYS_UNCONNECTED_1018,
         SYNOPSYS_UNCONNECTED_1019, SYNOPSYS_UNCONNECTED_1020,
         SYNOPSYS_UNCONNECTED_1021, SYNOPSYS_UNCONNECTED_1022,
         SYNOPSYS_UNCONNECTED_1023, SYNOPSYS_UNCONNECTED_1024,
         SYNOPSYS_UNCONNECTED_1025, SYNOPSYS_UNCONNECTED_1026,
         SYNOPSYS_UNCONNECTED_1027, SYNOPSYS_UNCONNECTED_1028,
         SYNOPSYS_UNCONNECTED_1029, SYNOPSYS_UNCONNECTED_1030,
         SYNOPSYS_UNCONNECTED_1031, SYNOPSYS_UNCONNECTED_1032,
         SYNOPSYS_UNCONNECTED_1033, SYNOPSYS_UNCONNECTED_1034,
         SYNOPSYS_UNCONNECTED_1035, SYNOPSYS_UNCONNECTED_1036,
         SYNOPSYS_UNCONNECTED_1037, SYNOPSYS_UNCONNECTED_1038,
         SYNOPSYS_UNCONNECTED_1039, SYNOPSYS_UNCONNECTED_1040,
         SYNOPSYS_UNCONNECTED_1041, SYNOPSYS_UNCONNECTED_1042,
         SYNOPSYS_UNCONNECTED_1043, SYNOPSYS_UNCONNECTED_1044,
         SYNOPSYS_UNCONNECTED_1045, SYNOPSYS_UNCONNECTED_1046,
         SYNOPSYS_UNCONNECTED_1047, SYNOPSYS_UNCONNECTED_1048,
         SYNOPSYS_UNCONNECTED_1049, SYNOPSYS_UNCONNECTED_1050,
         SYNOPSYS_UNCONNECTED_1051, SYNOPSYS_UNCONNECTED_1052,
         SYNOPSYS_UNCONNECTED_1053, SYNOPSYS_UNCONNECTED_1054,
         SYNOPSYS_UNCONNECTED_1055, SYNOPSYS_UNCONNECTED_1056,
         SYNOPSYS_UNCONNECTED_1057, SYNOPSYS_UNCONNECTED_1058,
         SYNOPSYS_UNCONNECTED_1059, SYNOPSYS_UNCONNECTED_1060,
         SYNOPSYS_UNCONNECTED_1061, SYNOPSYS_UNCONNECTED_1062,
         SYNOPSYS_UNCONNECTED_1063, SYNOPSYS_UNCONNECTED_1064,
         SYNOPSYS_UNCONNECTED_1065, SYNOPSYS_UNCONNECTED_1066,
         SYNOPSYS_UNCONNECTED_1067, SYNOPSYS_UNCONNECTED_1068,
         SYNOPSYS_UNCONNECTED_1069, SYNOPSYS_UNCONNECTED_1070,
         SYNOPSYS_UNCONNECTED_1071, SYNOPSYS_UNCONNECTED_1072,
         SYNOPSYS_UNCONNECTED_1073, SYNOPSYS_UNCONNECTED_1074,
         SYNOPSYS_UNCONNECTED_1075, SYNOPSYS_UNCONNECTED_1076,
         SYNOPSYS_UNCONNECTED_1077, SYNOPSYS_UNCONNECTED_1078,
         SYNOPSYS_UNCONNECTED_1079, SYNOPSYS_UNCONNECTED_1080,
         SYNOPSYS_UNCONNECTED_1081, SYNOPSYS_UNCONNECTED_1082,
         SYNOPSYS_UNCONNECTED_1083, SYNOPSYS_UNCONNECTED_1084,
         SYNOPSYS_UNCONNECTED_1085, SYNOPSYS_UNCONNECTED_1086,
         SYNOPSYS_UNCONNECTED_1087, SYNOPSYS_UNCONNECTED_1088, _padder__n2571 ,
         _padder__n2570 , _padder__n2569 , _padder__n2568 , _padder__n2567 ,
         _padder__n2566 , _padder__n2565 , _padder__n2564 , _padder__n2563 ,
         _padder__n2562 , _padder__n2561 , _padder__n2560 , _padder__n2559 ,
         _padder__n2558 , _padder__n2557 , _padder__n2556 , _padder__n2555 ,
         _padder__n2554 , _padder__n2553 , _padder__n2552 , _padder__n2551 ,
         _padder__n2550 , _padder__n2549 , _padder__n2548 , _padder__n2547 ,
         _padder__n2546 , _padder__n2545 , _padder__n2544 , _padder__n2543 ,
         _padder__n2542 , _padder__n2541 , _padder__n2540 , _padder__n2539 ,
         _padder__n2538 , _padder__n2537 , _padder__n2536 , _padder__n2535 ,
         _padder__n2534 , _padder__n2533 , _padder__n2532 , _padder__n2531 ,
         _padder__n2530 , _padder__n2529 , _padder__n2528 , _padder__n2527 ,
         _padder__n2526 , _padder__n2525 , _padder__n2524 , _padder__n2523 ,
         _padder__n2522 , _padder__n2521 , _padder__n2520 , _padder__n2519 ,
         _padder__n2518 , _padder__n2517 , _padder__n2516 , _padder__n2515 ,
         _padder__n2514 , _padder__n2513 , _padder__n2512 , _padder__n2511 ,
         _padder__n2510 , _padder__n2509 , _padder__n2508 , _padder__n2507 ,
         _padder__n2506 , _padder__n2505 , _padder__n2504 , _padder__n2503 ,
         _padder__n2502 , _padder__n2501 , _padder__n2500 , _padder__n2499 ,
         _padder__n2498 , _padder__n2497 , _padder__n2496 , _padder__n2495 ,
         _padder__n2494 , _padder__n2493 , _padder__n2492 , _padder__n2491 ,
         _padder__n2490 , _padder__n2489 , _padder__n2488 , _padder__n2487 ,
         _padder__n2486 , _padder__n2485 , _padder__n2484 , _padder__n2483 ,
         _padder__n2482 , _padder__n2480 , _padder__n2479 , _padder__n2478 ,
         _padder__n2477 , _padder__n2476 , _padder__n2475 , _padder__n2474 ,
         _padder__n2473 , _padder__n2472 , _padder__n2471 , _padder__n2470 ,
         _padder__n2469 , _padder__n2468 , _padder__n2467 , _padder__n2466 ,
         _padder__n2465 , _padder__n2464 , _padder__n2463 , _padder__n2462 ,
         _padder__n2461 , _padder__n2460 , _padder__n2459 , _padder__n2458 ,
         _padder__n2457 , _padder__n2456 , _padder__n2455 , _padder__n2454 ,
         _padder__n2453 , _padder__n2452 , _padder__n2451 , _padder__n2450 ,
         _padder__n2449 , _padder__n2448 , _padder__n2447 , _padder__n2446 ,
         _padder__n2445 , _padder__n2444 , _padder__n2443 , _padder__n2442 ,
         _padder__n2441 , _padder__n2440 , _padder__n2439 , _padder__n2438 ,
         _padder__n2437 , _padder__n2436 , _padder__n2435 , _padder__n2434 ,
         _padder__n2433 , _padder__n2432 , _padder__n2431 , _padder__n2430 ,
         _padder__n2429 , _padder__n2428 , _padder__n2427 , _padder__n2426 ,
         _padder__n2425 , _padder__n2424 , _padder__n2423 , _padder__n2422 ,
         _padder__n2421 , _padder__n2420 , _padder__n2419 , _padder__n2418 ,
         _padder__n2417 , _padder__n2416 , _padder__n2415 , _padder__n2414 ,
         _padder__n2413 , _padder__n2412 , _padder__n2411 , _padder__n2410 ,
         _padder__n2409 , _padder__n2408 , _padder__n2407 , _padder__n2406 ,
         _padder__n2405 , _padder__n2404 , _padder__n2403 , _padder__n2402 ,
         _padder__n2401 , _padder__n2400 , _padder__n2399 , _padder__n2398 ,
         _padder__n2397 , _padder__n2396 , _padder__n2395 , _padder__n2394 ,
         _padder__n2393 , _padder__n2392 , _padder__n2391 , _padder__n2390 ,
         _padder__n2389 , _padder__n2388 , _padder__n2387 , _padder__n2386 ,
         _padder__n2385 , _padder__n2384 , _padder__n2383 , _padder__n2382 ,
         _padder__n2381 , _padder__n2380 , _padder__n2379 , _padder__n2378 ,
         _padder__n2377 , _padder__n2376 , _padder__n2375 , _padder__n2374 ,
         _padder__n2373 , _padder__n2372 , _padder__n2371 , _padder__n2370 ,
         _padder__n2369 , _padder__n2368 , _padder__n2367 , _padder__n2366 ,
         _padder__n2365 , _padder__n2364 , _padder__n2363 , _padder__n2362 ,
         _padder__n2361 , _padder__n2360 , _padder__n2359 , _padder__n2358 ,
         _padder__n2357 , _padder__n2356 , _padder__n2355 , _padder__n2354 ,
         _padder__n2353 , _padder__n2352 , _padder__n2351 , _padder__n2350 ,
         _padder__n2349 , _padder__n2348 , _padder__n2347 , _padder__n2346 ,
         _padder__n2345 , _padder__n2344 , _padder__n2343 , _padder__n2342 ,
         _padder__n2341 , _padder__n2340 , _padder__n2339 , _padder__n2338 ,
         _padder__n2337 , _padder__n2336 , _padder__n2335 , _padder__n2334 ,
         _padder__n2333 , _padder__n2332 , _padder__n2331 , _padder__n2330 ,
         _padder__n2329 , _padder__n2328 , _padder__n2327 , _padder__n2326 ,
         _padder__n2325 , _padder__n2324 , _padder__n2323 , _padder__n2322 ,
         _padder__n2321 , _padder__n2320 , _padder__n2319 , _padder__n2318 ,
         _padder__n2317 , _padder__n2316 , _padder__n2315 , _padder__n2314 ,
         _padder__n2313 , _padder__n2312 , _padder__n2311 , _padder__n2310 ,
         _padder__n2309 , _padder__n2308 , _padder__n2307 , _padder__n2306 ,
         _padder__n2305 , _padder__n2304 , _padder__n2303 , _padder__n2302 ,
         _padder__n2301 , _padder__n2300 , _padder__n2299 , _padder__n2298 ,
         _padder__n2297 , _padder__n2296 , _padder__n2295 , _padder__n2294 ,
         _padder__n2293 , _padder__n2292 , _padder__n2291 , _padder__n2290 ,
         _padder__n2289 , _padder__n2288 , _padder__n2287 , _padder__n2286 ,
         _padder__n2285 , _padder__n2284 , _padder__n2283 , _padder__n2282 ,
         _padder__n2281 , _padder__n2280 , _padder__n2279 , _padder__n2278 ,
         _padder__n2277 , _padder__n2276 , _padder__n2275 , _padder__n2274 ,
         _padder__n2273 , _padder__n2272 , _padder__n2271 , _padder__n2270 ,
         _padder__n2269 , _padder__n2268 , _padder__n2267 , _padder__n2266 ,
         _padder__n2265 , _padder__n2264 , _padder__n2263 , _padder__n2262 ,
         _padder__n2261 , _padder__n2260 , _padder__n2259 , _padder__n2258 ,
         _padder__n2257 , _padder__n2256 , _padder__n2255 , _padder__n2254 ,
         _padder__n2253 , _padder__n2252 , _padder__n2251 , _padder__n2250 ,
         _padder__n2249 , _padder__n2248 , _padder__n2247 , _padder__n2246 ,
         _padder__n2245 , _padder__n2244 , _padder__n2243 , _padder__n2242 ,
         _padder__n2241 , _padder__n2240 , _padder__n2239 , _padder__n2238 ,
         _padder__n2237 , _padder__n2236 , _padder__n2235 , _padder__n2234 ,
         _padder__n2233 , _padder__n2232 , _padder__n2231 , _padder__n2230 ,
         _padder__n2229 , _padder__n2228 , _padder__n2227 , _padder__n2226 ,
         _padder__n2225 , _padder__n2224 , _padder__n2223 , _padder__n2222 ,
         _padder__n2221 , _padder__n2220 , _padder__n2219 , _padder__n2218 ,
         _padder__n2217 , _padder__n2216 , _padder__n2215 , _padder__n2214 ,
         _padder__n2213 , _padder__n2212 , _padder__n2211 , _padder__n2210 ,
         _padder__n2209 , _padder__n2208 , _padder__n2207 , _padder__n2206 ,
         _padder__n2205 , _padder__n2204 , _padder__n2203 , _padder__n2202 ,
         _padder__n2201 , _padder__n2200 , _padder__n2199 , _padder__n2198 ,
         _padder__n2197 , _padder__n2196 , _padder__n2195 , _padder__n2194 ,
         _padder__n2193 , _padder__n2192 , _padder__n2191 , _padder__n2190 ,
         _padder__n2189 , _padder__n2188 , _padder__n2187 , _padder__n2186 ,
         _padder__n2185 , _padder__n2184 , _padder__n2183 , _padder__n2182 ,
         _padder__n2181 , _padder__n2180 , _padder__n2179 , _padder__n2178 ,
         _padder__n2177 , _padder__n2176 , _padder__n2175 , _padder__n2174 ,
         _padder__n2173 , _padder__n2172 , _padder__n2171 , _padder__n2170 ,
         _padder__n2169 , _padder__n2168 , _padder__n2167 , _padder__n2166 ,
         _padder__n2165 , _padder__n2164 , _padder__n2163 , _padder__n2162 ,
         _padder__n2161 , _padder__n2160 , _padder__n2159 , _padder__n2158 ,
         _padder__n2157 , _padder__n2156 , _padder__n2155 , _padder__n2154 ,
         _padder__n2153 , _padder__n2152 , _padder__n2151 , _padder__n2150 ,
         _padder__n2149 , _padder__n2148 , _padder__n2147 , _padder__n2146 ,
         _padder__n2145 , _padder__n2144 , _padder__n2143 , _padder__n2142 ,
         _padder__n2141 , _padder__n2140 , _padder__n2139 , _padder__n2138 ,
         _padder__n2137 , _padder__n2136 , _padder__n2135 , _padder__n2134 ,
         _padder__n2133 , _padder__n2132 , _padder__n2131 , _padder__n2130 ,
         _padder__n2129 , _padder__n2128 , _padder__n2127 , _padder__n2126 ,
         _padder__n2125 , _padder__n2124 , _padder__n2123 , _padder__n2122 ,
         _padder__n2121 , _padder__n2120 , _padder__n2119 , _padder__n2118 ,
         _padder__n2117 , _padder__n2116 , _padder__n2115 , _padder__n2114 ,
         _padder__n2113 , _padder__n2112 , _padder__n2111 , _padder__n2110 ,
         _padder__n2109 , _padder__n2108 , _padder__n2107 , _padder__n2106 ,
         _padder__n2105 , _padder__n2104 , _padder__n2103 , _padder__n2102 ,
         _padder__n2101 , _padder__n2100 , _padder__n2099 , _padder__n2098 ,
         _padder__n2097 , _padder__n2096 , _padder__n2095 , _padder__n2094 ,
         _padder__n2093 , _padder__n2092 , _padder__n2091 , _padder__n2090 ,
         _padder__n2089 , _padder__n2088 , _padder__n2087 , _padder__n2086 ,
         _padder__n2085 , _padder__n2084 , _padder__n2083 , _padder__n2082 ,
         _padder__n2081 , _padder__n2080 , _padder__n2079 , _padder__n2078 ,
         _padder__n2077 , _padder__n2076 , _padder__n2075 , _padder__n2074 ,
         _padder__n2073 , _padder__n2072 , _padder__n2071 , _padder__n2070 ,
         _padder__n2069 , _padder__n2068 , _padder__n2067 , _padder__n2066 ,
         _padder__n2065 , _padder__n2064 , _padder__n2063 , _padder__n2062 ,
         _padder__n2061 , _padder__n2060 , _padder__n2059 , _padder__n2058 ,
         _padder__n2057 , _padder__n2056 , _padder__n2055 , _padder__n2054 ,
         _padder__n2053 , _padder__n2052 , _padder__n2051 , _padder__n2050 ,
         _padder__n2049 , _padder__n2048 , _padder__n2047 , _padder__n2046 ,
         _padder__n2045 , _padder__n2044 , _padder__n2043 , _padder__n2042 ,
         _padder__n2041 , _padder__n2040 , _padder__n2039 , _padder__n2038 ,
         _padder__n2037 , _padder__n2036 , _padder__n2035 , _padder__n2034 ,
         _padder__n2033 , _padder__n2032 , _padder__n2031 , _padder__n2030 ,
         _padder__n2029 , _padder__n2028 , _padder__n2027 , _padder__n2026 ,
         _padder__n2025 , _padder__n2024 , _padder__n2023 , _padder__n2022 ,
         _padder__n2021 , _padder__n2020 , _padder__n2019 , _padder__n2018 ,
         _padder__n2017 , _padder__n2016 , _padder__n2015 , _padder__n2014 ,
         _padder__n2013 , _padder__n2012 , _padder__n2011 , _padder__n2010 ,
         _padder__n2009 , _padder__n2008 , _padder__n2007 , _padder__n2006 ,
         _padder__n2005 , _padder__n2004 , _padder__n2003 , _padder__n2002 ,
         _padder__n2001 , _padder__n2000 , _padder__n1999 , _padder__n1998 ,
         _padder__n1997 , _padder__n1996 , _padder__n1995 , _padder__n1994 ,
         _padder__n1993 , _padder__n1992 , _padder__n1991 , _padder__n1990 ,
         _padder__n1989 , _padder__n1988 , _padder__n1987 , _padder__n1986 ,
         _padder__n1985 , _padder__n1984 , _padder__n1983 , _padder__n1982 ,
         _padder__n1981 , _padder__n1980 , _padder__n1979 , _padder__n1978 ,
         _padder__n1977 , _padder__n1976 , _padder__n1975 , _padder__n1974 ,
         _padder__n1973 , _padder__n1972 , _padder__n1971 , _padder__n1970 ,
         _padder__n1969 , _padder__n1968 , _padder__n1967 , _padder__n1966 ,
         _padder__n1965 , _padder__n1964 , _padder__n1963 , _padder__n1962 ,
         _padder__n1960 , _padder__n1959 , _padder__n1958 , _padder__n1957 ,
         _padder__n1956 , _padder__n1955 , _padder__n1954 , _padder__n1953 ,
         _padder__n1952 , _padder__n1951 , _padder__n1950 , _padder__n1949 ,
         _padder__n1948 , _padder__n1947 , _padder__n1946 , _padder__n1945 ,
         _padder__n1944 , _padder__n1943 , _padder__n1942 , _padder__n1941 ,
         _padder__n1940 , _padder__n1939 , _padder__n1938 , _padder__n1937 ,
         _padder__n1936 , _padder__n1935 , _padder__n1934 , _padder__n1933 ,
         _padder__n1932 , _padder__n1931 , _padder__n1930 , _padder__n1929 ,
         _padder__n1928 , _padder__n1927 , _padder__n1926 , _padder__n1925 ,
         _padder__n1924 , _padder__n1923 , _padder__n1922 , _padder__n1921 ,
         _padder__n1920 , _padder__n1919 , _padder__n1918 , _padder__n1917 ,
         _padder__n1916 , _padder__n1915 , _padder__n1914 , _padder__n1913 ,
         _padder__n1912 , _padder__n1911 , _padder__n1910 , _padder__n1909 ,
         _padder__n1908 , _padder__n1907 , _padder__n1906 , _padder__n1905 ,
         _padder__n1904 , _padder__n1903 , _padder__n1902 , _padder__n1901 ,
         _padder__n1900 , _padder__n1899 , _padder__n1898 , _padder__n1897 ,
         _padder__n1896 , _padder__n1895 , _padder__n1894 , _padder__n1893 ,
         _padder__n1892 , _padder__n1891 , _padder__n1890 , _padder__n1889 ,
         _padder__n1888 , _padder__n1887 , _padder__n1886 , _padder__n1885 ,
         _padder__n1884 , _padder__n1883 , _padder__n1882 , _padder__n1881 ,
         _padder__n1880 , _padder__n1879 , _padder__n1878 , _padder__n1877 ,
         _padder__n1876 , _padder__n1875 , _padder__n1874 , _padder__n1873 ,
         _padder__n1872 , _padder__n1871 , _padder__n1870 , _padder__n1869 ,
         _padder__n1868 , _padder__n1867 , _padder__n1866 , _padder__n1865 ,
         _padder__n1864 , _padder__n1863 , _padder__n1862 , _padder__n1861 ,
         _padder__n1860 , _padder__n1859 , _padder__n1858 , _padder__n1857 ,
         _padder__n1856 , _padder__n1855 , _padder__n1854 , _padder__n1853 ,
         _padder__n1852 , _padder__n1851 , _padder__n1850 , _padder__n1849 ,
         _padder__n1848 , _padder__n1847 , _padder__n1846 , _padder__n1845 ,
         _padder__n1844 , _padder__n1843 , _padder__n1842 , _padder__n1841 ,
         _padder__n1840 , _padder__n1839 , _padder__n1838 , _padder__n1837 ,
         _padder__n1240 , _padder__n1239 , _padder__n1238 , _padder__n1237 ,
         _padder__n1236 , _padder__n1235 , _padder__n1234 , _padder__n1233 ,
         _padder__n1232 , _padder__n1231 , _padder__n1230 , _padder__n1229 ,
         _padder__n1228 , _padder__n1227 , _padder__n1226 , _padder__n1225 ,
         _padder__n1224 , _padder__n1223 , _padder__n1222 , _padder__n1221 ,
         _padder__n1220 , _padder__n1219 , _padder__n1218 , _padder__n1217 ,
         _padder__n1216 , _padder__n1215 , _padder__n1214 , _padder__n1213 ,
         _padder__n1212 , _padder__n1211 , _padder__n1210 , _padder__n1209 ,
         _padder__n1208 , _padder__n1207 , _padder__n1206 , _padder__n1205 ,
         _padder__n1204 , _padder__n1203 , _padder__n1202 , _padder__n1201 ,
         _padder__n1200 , _padder__n1199 , _padder__n1198 , _padder__n1197 ,
         _padder__n1196 , _padder__n1195 , _padder__n1194 , _padder__n1193 ,
         _padder__n1192 , _padder__n1191 , _padder__n1190 , _padder__n1189 ,
         _padder__n1188 , _padder__n1187 , _padder__n1186 , _padder__n1185 ,
         _padder__n1184 , _padder__n1183 , _padder__n1182 , _padder__n1181 ,
         _padder__n1180 , _padder__n1179 , _padder__n1178 , _padder__n1177 ,
         _padder__n1176 , _padder__n1175 , _padder__n1174 , _padder__n1173 ,
         _padder__n1172 , _padder__n1171 , _padder__n1170 , _padder__n1169 ,
         _padder__n1168 , _padder__n1167 , _padder__n1166 , _padder__n1165 ,
         _padder__n1164 , _padder__n1163 , _padder__n1162 , _padder__n1161 ,
         _padder__n1160 , _padder__n1159 , _padder__n1158 , _padder__n1157 ,
         _padder__n1156 , _padder__n1155 , _padder__n1154 , _padder__n1153 ,
         _padder__n1152 , _padder__n1151 , _padder__n1150 , _padder__n1149 ,
         _padder__n1148 , _padder__n1147 , _padder__n1146 , _padder__n1145 ,
         _padder__n1144 , _padder__n1143 , _padder__n1142 , _padder__n1141 ,
         _padder__n1140 , _padder__n1139 , _padder__n1138 , _padder__n1137 ,
         _padder__n1136 , _padder__n1135 , _padder__n1134 , _padder__n1133 ,
         _padder__n1132 , _padder__n1131 , _padder__n1130 , _padder__n1129 ,
         _padder__n1128 , _padder__n1127 , _padder__n1126 , _padder__n1125 ,
         _padder__n1124 , _padder__n1123 , _padder__n1122 , _padder__n1121 ,
         _padder__n1120 , _padder__n1119 , _padder__n1118 , _padder__n1117 ,
         _padder__n1116 , _padder__n1115 , _padder__n1114 , _padder__n1113 ,
         _padder__n1112 , _padder__n1111 , _padder__n1110 , _padder__n1109 ,
         _padder__n1108 , _padder__n1107 , _padder__n1106 , _padder__n1105 ,
         _padder__n1104 , _padder__n1103 , _padder__n1102 , _padder__n1101 ,
         _padder__n1100 , _padder__n1099 , _padder__n1098 , _padder__n1097 ,
         _padder__n1096 , _padder__n1095 , _padder__n1094 , _padder__n1093 ,
         _padder__n1092 , _padder__n1091 , _padder__n1090 , _padder__n1089 ,
         _padder__n1088 , _padder__n1087 , _padder__n1086 , _padder__n1085 ,
         _padder__n1084 , _padder__n1083 , _padder__n1082 , _padder__n1081 ,
         _padder__n1080 , _padder__n1079 , _padder__n1078 , _padder__n1077 ,
         _padder__n1076 , _padder__n1075 , _padder__n1074 , _padder__n1073 ,
         _padder__n1072 , _padder__n1071 , _padder__n1070 , _padder__n1069 ,
         _padder__n1068 , _padder__n1067 , _padder__n1066 , _padder__n1065 ,
         _padder__n1064 , _padder__n1063 , _padder__n1062 , _padder__n1061 ,
         _padder__n1060 , _padder__n1059 , _padder__n1058 , _padder__n1057 ,
         _padder__n1056 , _padder__n1055 , _padder__n1054 , _padder__n1053 ,
         _padder__n1052 , _padder__n1051 , _padder__n1050 , _padder__n1049 ,
         _padder__n1048 , _padder__n1047 , _padder__n1046 , _padder__n1045 ,
         _padder__n1044 , _padder__n1043 , _padder__n1042 , _padder__n1041 ,
         _padder__n1040 , _padder__n1039 , _padder__n1038 , _padder__n1037 ,
         _padder__n1036 , _padder__n1035 , _padder__n1034 , _padder__n1033 ,
         _padder__n1032 , _padder__n1031 , _padder__n1030 , _padder__n1029 ,
         _padder__n1028 , _padder__n1027 , _padder__n1026 , _padder__n1025 ,
         _padder__n1024 , _padder__n1023 , _padder__n1022 , _padder__n1021 ,
         _padder__n1020 , _padder__n1019 , _padder__n1018 , _padder__n1017 ,
         _padder__n1016 , _padder__n1015 , _padder__n1014 , _padder__n1013 ,
         _padder__n1012 , _padder__n1011 , _padder__n1010 , _padder__n1009 ,
         _padder__n1008 , _padder__n1007 , _padder__n1006 , _padder__n1005 ,
         _padder__n1004 , _padder__n1003 , _padder__n1002 , _padder__n1001 ,
         _padder__n1000 , _padder__n999 , _padder__n998 , _padder__n997 ,
         _padder__n996 , _padder__n995 , _padder__n994 , _padder__n993 ,
         _padder__n992 , _padder__n991 , _padder__n990 , _padder__n989 ,
         _padder__n988 , _padder__n987 , _padder__n986 , _padder__n985 ,
         _padder__n984 , _padder__n983 , _padder__n982 , _padder__n981 ,
         _padder__n980 , _padder__n979 , _padder__n978 , _padder__n977 ,
         _padder__n976 , _padder__n975 , _padder__n974 , _padder__n973 ,
         _padder__n972 , _padder__n971 , _padder__n970 , _padder__n969 ,
         _padder__n968 , _padder__n967 , _padder__n966 , _padder__n965 ,
         _padder__n964 , _padder__n963 , _padder__n962 , _padder__n961 ,
         _padder__n960 , _padder__n959 , _padder__n958 , _padder__n957 ,
         _padder__n956 , _padder__n955 , _padder__n954 , _padder__n953 ,
         _padder__n952 , _padder__n951 , _padder__n950 , _padder__n949 ,
         _padder__n948 , _padder__n947 , _padder__n946 , _padder__n945 ,
         _padder__n944 , _padder__n943 , _padder__n942 , _padder__n941 ,
         _padder__n940 , _padder__n939 , _padder__n938 , _padder__n937 ,
         _padder__n936 , _padder__n935 , _padder__n934 , _padder__n933 ,
         _padder__n932 , _padder__n931 , _padder__n930 , _padder__n929 ,
         _padder__n928 , _padder__n927 , _padder__n926 , _padder__n925 ,
         _padder__n924 , _padder__n923 , _padder__n922 , _padder__n921 ,
         _padder__n920 , _padder__n919 , _padder__n918 , _padder__n917 ,
         _padder__n916 , _padder__n915 , _padder__n914 , _padder__n913 ,
         _padder__n912 , _padder__n911 , _padder__n910 , _padder__n909 ,
         _padder__n908 , _padder__n907 , _padder__n906 , _padder__n905 ,
         _padder__n904 , _padder__n903 , _padder__n902 , _padder__n901 ,
         _padder__n900 , _padder__n899 , _padder__n898 , _padder__n897 ,
         _padder__n896 , _padder__n895 , _padder__n894 , _padder__n893 ,
         _padder__n892 , _padder__n891 , _padder__n890 , _padder__n889 ,
         _padder__n888 , _padder__n887 , _padder__n886 , _padder__n885 ,
         _padder__n884 , _padder__n883 , _padder__n882 , _padder__n881 ,
         _padder__n880 , _padder__n879 , _padder__n878 , _padder__n877 ,
         _padder__n876 , _padder__n875 , _padder__n874 , _padder__n873 ,
         _padder__n872 , _padder__n871 , _padder__n870 , _padder__n869 ,
         _padder__n868 , _padder__n867 , _padder__n866 , _padder__n865 ,
         _padder__n864 , _padder__n863 , _padder__n862 , _padder__n861 ,
         _padder__n860 , _padder__n859 , _padder__n858 , _padder__n857 ,
         _padder__n856 , _padder__n855 , _padder__n854 , _padder__n853 ,
         _padder__n852 , _padder__n851 , _padder__n850 , _padder__n849 ,
         _padder__n848 , _padder__n847 , _padder__n846 , _padder__n845 ,
         _padder__n844 , _padder__n843 , _padder__n842 , _padder__n841 ,
         _padder__n840 , _padder__n839 , _padder__n838 , _padder__n837 ,
         _padder__n836 , _padder__n835 , _padder__n834 , _padder__n833 ,
         _padder__n832 , _padder__n831 , _padder__n830 , _padder__n829 ,
         _padder__n828 , _padder__n827 , _padder__n826 , _padder__n825 ,
         _padder__n824 , _padder__n823 , _padder__n822 , _padder__n821 ,
         _padder__n820 , _padder__n819 , _padder__n818 , _padder__n817 ,
         _padder__n816 , _padder__n815 , _padder__n814 , _padder__n813 ,
         _padder__n812 , _padder__n811 , _padder__n810 , _padder__n809 ,
         _padder__n808 , _padder__n807 , _padder__n806 , _padder__n805 ,
         _padder__n804 , _padder__n803 , _padder__n802 , _padder__n801 ,
         _padder__n800 , _padder__n799 , _padder__n798 , _padder__n797 ,
         _padder__n796 , _padder__n795 , _padder__n794 , _padder__n793 ,
         _padder__n792 , _padder__n791 , _padder__n790 , _padder__n789 ,
         _padder__n788 , _padder__n787 , _padder__n786 , _padder__n785 ,
         _padder__n784 , _padder__n783 , _padder__n782 , _padder__n781 ,
         _padder__n780 , _padder__n779 , _padder__n778 , _padder__n777 ,
         _padder__n776 , _padder__n775 , _padder__n774 , _padder__n773 ,
         _padder__n772 , _padder__n771 , _padder__n770 , _padder__n769 ,
         _padder__n768 , _padder__n767 , _padder__n766 , _padder__n765 ,
         _padder__n764 , _padder__n763 , _padder__n762 , _padder__n761 ,
         _padder__n760 , _padder__n759 , _padder__n758 , _padder__n757 ,
         _padder__n756 , _padder__n755 , _padder__n754 , _padder__n753 ,
         _padder__n752 , _padder__n751 , _padder__n750 , _padder__n749 ,
         _padder__n748 , _padder__n747 , _padder__n746 , _padder__n745 ,
         _padder__n744 , _padder__n743 , _padder__n742 , _padder__n741 ,
         _padder__n740 , _padder__n739 , _padder__n738 , _padder__n737 ,
         _padder__n736 , _padder__n735 , _padder__n734 , _padder__n733 ,
         _padder__n732 , _padder__n731 , _padder__n730 , _padder__n729 ,
         _padder__n728 , _padder__n727 , _padder__n726 , _padder__n725 ,
         _padder__n724 , _padder__n723 , _padder__n722 , _padder__n721 ,
         _padder__n720 , _padder__n719 , _padder__n718 , _padder__n717 ,
         _padder__n716 , _padder__n715 , _padder__n714 , _padder__n713 ,
         _padder__n712 , _padder__n711 , _padder__n710 , _padder__n709 ,
         _padder__n708 , _padder__n707 , _padder__n706 , _padder__n705 ,
         _padder__n704 , _padder__n703 , _padder__n702 , _padder__n701 ,
         _padder__n700 , _padder__n699 , _padder__n698 , _padder__n697 ,
         _padder__n696 , _padder__n695 , _padder__n694 , _padder__n693 ,
         _padder__n692 , _padder__n691 , _padder__n690 , _padder__n689 ,
         _padder__n688 , _padder__n687 , _padder__n686 , _padder__n685 ,
         _padder__n683 , _padder__n682 , _padder__n681 , _padder__n680 ,
         _padder__n679 , _padder__n678 , _padder__n677 , _padder__n676 ,
         _padder__n675 , _padder__n674 , _padder__n673 , _padder__n672 ,
         _padder__n671 , _padder__n670 , _padder__n669 , _padder__n668 ,
         _padder__n667 , _padder__n666 , _padder__n664 , _padder__n663 ,
         _padder__n662 , _padder__n660 , _padder__n659 , _padder__n658 ,
         _padder__n657 , _padder__n656 , _padder__n655 , _padder__n654 ,
         _padder__n653 , _padder__n652 , _padder__n651 , _padder__n650 ,
         _padder__n649 , _padder__n648 , _padder__n647 , _padder__n646 ,
         _padder__n645 , _padder__n644 , _padder__n643 , _padder__n642 ,
         _padder__n641 , _padder__n640 , _padder__n639 , _padder__n638 ,
         _padder__n637 , _padder__n636 , _padder__n635 , _padder__n634 ,
         _padder__n633 , _padder__n632 , _padder__n631 , _padder__n630 ,
         _padder__n629 , _padder__n628 , _padder__n627 , _padder__n624 ,
         _padder__n623 , _padder__n622 , _padder__n621 , _padder__n619 ,
         _padder__n618 , _padder__n617 , _padder__n616 , _padder__n615 ,
         _padder__n614 , _padder__n613 , _padder__n612 , _padder__n611 ,
         _padder__n610 , _padder__n609 , _padder__n608 , _padder__n607 ,
         _padder__n606 , _padder__n605 , _padder__n604 , _padder__n603 ,
         _padder__n602 , _padder__n598 , _padder__n1961 , _padder__n1836 ,
         _padder__n1835 , _padder__n1834 , _padder__n1833 , _padder__n1832 ,
         _padder__n1831 , _padder__n1830 , _padder__n1829 , _padder__n1828 ,
         _padder__n1827 , _padder__n1826 , _padder__n1825 , _padder__n1824 ,
         _padder__n1823 , _padder__n1822 , _padder__n1821 , _padder__n1820 ,
         _padder__n1819 , _padder__n1818 , _padder__n1817 , _padder__n1816 ,
         _padder__n1815 , _padder__n1814 , _padder__n1813 , _padder__n1812 ,
         _padder__n1811 , _padder__n1810 , _padder__n1808 , _padder__n1807 ,
         _padder__n1806 , _padder__n1805 , _padder__n1804 , _padder__n1803 ,
         _padder__n1802 , _padder__n1801 , _padder__n1800 , _padder__n1799 ,
         _padder__n1798 , _padder__n1797 , _padder__n1796 , _padder__n1795 ,
         _padder__n1794 , _padder__n1793 , _padder__n1792 , _padder__n1791 ,
         _padder__n1790 , _padder__n1789 , _padder__n1788 , _padder__n1787 ,
         _padder__n1786 , _padder__n1785 , _padder__n1784 , _padder__n1783 ,
         _padder__n1782 , _padder__n1781 , _padder__n1780 , _padder__n1779 ,
         _padder__n1778 , _padder__n1777 , _padder__n1776 , _padder__n1775 ,
         _padder__n1774 , _padder__n1773 , _padder__n1772 , _padder__n1771 ,
         _padder__n1770 , _padder__n1769 , _padder__n1768 , _padder__n1767 ,
         _padder__n1766 , _padder__n1765 , _padder__n1764 , _padder__n1763 ,
         _padder__n1762 , _padder__n1761 , _padder__n1760 , _padder__n1759 ,
         _padder__n1758 , _padder__n1757 , _padder__n1756 , _padder__n1755 ,
         _padder__n1754 , _padder__n1753 , _padder__n1752 , _padder__n1751 ,
         _padder__n1750 , _padder__n1749 , _padder__n1748 , _padder__n1747 ,
         _padder__n1746 , _padder__n1745 , _padder__n1744 , _padder__n1743 ,
         _padder__n1742 , _padder__n1741 , _padder__n1740 , _padder__n1739 ,
         _padder__n1738 , _padder__n1737 , _padder__n1736 , _padder__n1735 ,
         _padder__n1734 , _padder__n1733 , _padder__n1732 , _padder__n1731 ,
         _padder__n1730 , _padder__n1729 , _padder__n1728 , _padder__n1727 ,
         _padder__n1726 , _padder__n1725 , _padder__n1724 , _padder__n1723 ,
         _padder__n1722 , _padder__n1721 , _padder__n1720 , _padder__n1719 ,
         _padder__n1718 , _padder__n1717 , _padder__n1716 , _padder__n1715 ,
         _padder__n1714 , _padder__n1713 , _padder__n1712 , _padder__n1711 ,
         _padder__n1710 , _padder__n1709 , _padder__n1708 , _padder__n1707 ,
         _padder__n1706 , _padder__n1705 , _padder__n1704 , _padder__n1703 ,
         _padder__n1702 , _padder__n1701 , _padder__n1700 , _padder__n1699 ,
         _padder__n1698 , _padder__n1697 , _padder__n1696 , _padder__n1695 ,
         _padder__n1694 , _padder__n1693 , _padder__n1692 , _padder__n1691 ,
         _padder__n1690 , _padder__n1689 , _padder__n1688 , _padder__n1687 ,
         _padder__n1686 , _padder__n1685 , _padder__n1684 , _padder__n1683 ,
         _padder__n1682 , _padder__n1681 , _padder__n1680 , _padder__n1679 ,
         _padder__n1678 , _padder__n1677 , _padder__n1676 , _padder__n1675 ,
         _padder__n1674 , _padder__n1673 , _padder__n1672 , _padder__n1671 ,
         _padder__n1670 , _padder__n1669 , _padder__n1668 , _padder__n1667 ,
         _padder__n1666 , _padder__n1665 , _padder__n1664 , _padder__n1663 ,
         _padder__n1662 , _padder__n1661 , _padder__n1660 , _padder__n1659 ,
         _padder__n1658 , _padder__n1657 , _padder__n1656 , _padder__n1655 ,
         _padder__n1654 , _padder__n1653 , _padder__n1652 , _padder__n1651 ,
         _padder__n1650 , _padder__n1649 , _padder__n1648 , _padder__n1647 ,
         _padder__n1646 , _padder__n1645 , _padder__n1644 , _padder__n1643 ,
         _padder__n1642 , _padder__n1641 , _padder__n1640 , _padder__n1639 ,
         _padder__n1638 , _padder__n1637 , _padder__n1636 , _padder__n1635 ,
         _padder__n1634 , _padder__n1633 , _padder__n1632 , _padder__n1631 ,
         _padder__n1630 , _padder__n1629 , _padder__n1628 , _padder__n1627 ,
         _padder__n1626 , _padder__n1625 , _padder__n1624 , _padder__n1623 ,
         _padder__n1622 , _padder__n1621 , _padder__n1620 , _padder__n1619 ,
         _padder__n1618 , _padder__n1617 , _padder__n1616 , _padder__n1615 ,
         _padder__n1614 , _padder__n1613 , _padder__n1612 , _padder__n1611 ,
         _padder__n1610 , _padder__n1609 , _padder__n1608 , _padder__n1607 ,
         _padder__n1606 , _padder__n1605 , _padder__n1604 , _padder__n1603 ,
         _padder__n1602 , _padder__n1601 , _padder__n1600 , _padder__n1599 ,
         _padder__n1598 , _padder__n1597 , _padder__n1596 , _padder__n1595 ,
         _padder__n1594 , _padder__n1593 , _padder__n1592 , _padder__n1591 ,
         _padder__n1590 , _padder__n1589 , _padder__n1588 , _padder__n1587 ,
         _padder__n1586 , _padder__n1585 , _padder__n1584 , _padder__n1583 ,
         _padder__n1582 , _padder__n1581 , _padder__n1580 , _padder__n1579 ,
         _padder__n1578 , _padder__n1577 , _padder__n1576 , _padder__n1575 ,
         _padder__n1574 , _padder__n1573 , _padder__n1572 , _padder__n1571 ,
         _padder__n1570 , _padder__n1569 , _padder__n1568 , _padder__n1567 ,
         _padder__n1566 , _padder__n1565 , _padder__n1564 , _padder__n1563 ,
         _padder__n1562 , _padder__n1561 , _padder__n1560 , _padder__n1559 ,
         _padder__n1558 , _padder__n1557 , _padder__n1556 , _padder__n1555 ,
         _padder__n1554 , _padder__n1553 , _padder__n1552 , _padder__n1551 ,
         _padder__n1550 , _padder__n1549 , _padder__n1548 , _padder__n1547 ,
         _padder__n1546 , _padder__n1545 , _padder__n1544 , _padder__n1543 ,
         _padder__n1542 , _padder__n1541 , _padder__n1540 , _padder__n1539 ,
         _padder__n1538 , _padder__n1537 , _padder__n1536 , _padder__n1535 ,
         _padder__n1534 , _padder__n1533 , _padder__n1532 , _padder__n1531 ,
         _padder__n1530 , _padder__n1529 , _padder__n1528 , _padder__n1527 ,
         _padder__n1526 , _padder__n1525 , _padder__n1524 , _padder__n1523 ,
         _padder__n1522 , _padder__n1521 , _padder__n1520 , _padder__n1519 ,
         _padder__n1518 , _padder__n1517 , _padder__n1516 , _padder__n1515 ,
         _padder__n1514 , _padder__n1513 , _padder__n1512 , _padder__n1511 ,
         _padder__n1510 , _padder__n1509 , _padder__n1508 , _padder__n1507 ,
         _padder__n1506 , _padder__n1505 , _padder__n1504 , _padder__n1503 ,
         _padder__n1502 , _padder__n1501 , _padder__n1500 , _padder__n1499 ,
         _padder__n1498 , _padder__n1497 , _padder__n1496 , _padder__n1495 ,
         _padder__n1494 , _padder__n1493 , _padder__n1492 , _padder__n1491 ,
         _padder__n1490 , _padder__n1489 , _padder__n1488 , _padder__n1487 ,
         _padder__n1486 , _padder__n1485 , _padder__n1484 , _padder__n1483 ,
         _padder__n1482 , _padder__n1481 , _padder__n1480 , _padder__n1479 ,
         _padder__n1478 , _padder__n1477 , _padder__n1476 , _padder__n1475 ,
         _padder__n1474 , _padder__n1473 , _padder__n1472 , _padder__n1471 ,
         _padder__n1470 , _padder__n1469 , _padder__n1468 , _padder__n1467 ,
         _padder__n1466 , _padder__n1465 , _padder__n1464 , _padder__n1463 ,
         _padder__n1462 , _padder__n1461 , _padder__n1460 , _padder__n1459 ,
         _padder__n1458 , _padder__n1457 , _padder__n1456 , _padder__n1455 ,
         _padder__n1454 , _padder__n1453 , _padder__n1452 , _padder__n1451 ,
         _padder__n1450 , _padder__n1449 , _padder__n1448 , _padder__n1447 ,
         _padder__n1446 , _padder__n1445 , _padder__n1444 , _padder__n1443 ,
         _padder__n1442 , _padder__n1441 , _padder__n1440 , _padder__n1439 ,
         _padder__n1438 , _padder__n1437 , _padder__n1436 , _padder__n1435 ,
         _padder__n1434 , _padder__n1433 , _padder__n1432 , _padder__n1431 ,
         _padder__n1430 , _padder__n1429 , _padder__n1428 , _padder__n1427 ,
         _padder__n1426 , _padder__n1425 , _padder__n1424 , _padder__n1423 ,
         _padder__n1422 , _padder__n1421 , _padder__n1420 , _padder__n1419 ,
         _padder__n1418 , _padder__n1417 , _padder__n1416 , _padder__n1415 ,
         _padder__n1414 , _padder__n1413 , _padder__n1412 , _padder__n1411 ,
         _padder__n1410 , _padder__n1409 , _padder__n1408 , _padder__n1407 ,
         _padder__n1406 , _padder__n1405 , _padder__n1404 , _padder__n1403 ,
         _padder__n1402 , _padder__n1401 , _padder__n1400 , _padder__n1399 ,
         _padder__n1398 , _padder__n1397 , _padder__n1396 , _padder__n1395 ,
         _padder__n1394 , _padder__n1393 , _padder__n1392 , _padder__n1391 ,
         _padder__n1390 , _padder__n1389 , _padder__n1388 , _padder__n1387 ,
         _padder__n1386 , _padder__n1385 , _padder__n1384 , _padder__n1383 ,
         _padder__n1382 , _padder__n1381 , _padder__n1380 , _padder__n1379 ,
         _padder__n1378 , _padder__n1377 , _padder__n1376 , _padder__n1375 ,
         _padder__n1374 , _padder__n1373 , _padder__n1372 , _padder__n1371 ,
         _padder__n1370 , _padder__n1369 , _padder__n1368 , _padder__n1367 ,
         _padder__n1366 , _padder__n1365 , _padder__n1364 , _padder__n1363 ,
         _padder__n1362 , _padder__n1361 , _padder__n1360 , _padder__n1359 ,
         _padder__n1358 , _padder__n1357 , _padder__n1356 , _padder__n1355 ,
         _padder__n1354 , _padder__n1353 , _padder__n1352 , _padder__n1351 ,
         _padder__n1350 , _padder__n1349 , _padder__n1348 , _padder__n1347 ,
         _padder__n1346 , _padder__n1345 , _padder__n1344 , _padder__n1343 ,
         _padder__n1342 , _padder__n1341 , _padder__n1340 , _padder__n1339 ,
         _padder__n1338 , _padder__n1337 , _padder__n1336 , _padder__n1335 ,
         _padder__n1334 , _padder__n1333 , _padder__n1332 , _padder__n1331 ,
         _padder__n1330 , _padder__n1329 , _padder__n1328 , _padder__n1327 ,
         _padder__n1326 , _padder__n1325 , _padder__n1324 , _padder__n1323 ,
         _padder__n1322 , _padder__n1321 , _padder__n1320 , _padder__n1319 ,
         _padder__n1318 , _padder__n1317 , _padder__n1316 , _padder__n1315 ,
         _padder__n1314 , _padder__n1313 , _padder__n1312 , _padder__n1311 ,
         _padder__n1310 , _padder__n1309 , _padder__n1308 , _padder__n1307 ,
         _padder__n1306 , _padder__n1305 , _padder__n1304 , _padder__n1303 ,
         _padder__n1302 , _padder__n1301 , _padder__n1300 , _padder__n1299 ,
         _padder__n1298 , _padder__n1297 , _padder__n1296 , _padder__n1295 ,
         _padder__n1294 , _padder__n1293 , _padder__n1292 , _padder__n1291 ,
         _padder__n1290 , _padder__n1289 , _padder__n1288 , _padder__n1287 ,
         _padder__n1286 , _padder__n1285 , _padder__n1284 , _padder__n1283 ,
         _padder__n1282 , _padder__n1281 , _padder__n1280 , _padder__n1279 ,
         _padder__n1278 , _padder__n1277 , _padder__n1276 , _padder__n1275 ,
         _padder__n1274 , _padder__n1273 , _padder__n1272 , _padder__n1271 ,
         _padder__n1270 , _padder__n1269 , _padder__n1268 , _padder__n1267 ,
         _padder__n1266 , _padder__n1265 , _padder__n1264 , _padder__n1263 ,
         _padder__n1262 , _padder__n1261 , _padder__n1260 , _padder__n1259 ,
         _padder__n1258 , _padder__n1257 , _padder__n1256 , _padder__n1255 ,
         _padder__n1254 , _padder__n1253 , _padder__n1252 , _padder__n1251 ,
         _padder__n1250 , _padder__n1249 , _padder__n1248 , _padder__n1247 ,
         _padder__n1246 , _padder__n1245 , _padder__n1244 , _padder__n1243 ,
         _padder__n1242 , _padder__n1241 , _padder__state ,
         _padder__p0_out[7] , _padder__p0_out[6] , _padder__p0_out[5] ,
         _padder__p0_out[4] , _padder__p0_out[3] , _padder__p0_out[2] ,
         _padder__p0_out[1] , _padder__p0_n8 , _padder__p0_n7 ,
         _padder__p0_n6 , _padder__p0_n5 , _padder__p0_n4 , _padder__p0_n3 ,
         _padder__p0_n2 , _padder__p0_n1 , _f_permutation__n7326 ,
         _f_permutation__n7325 , _f_permutation__n7324 ,
         _f_permutation__n7323 , _f_permutation__n7322 ,
         _f_permutation__n7321 , _f_permutation__n7320 ,
         _f_permutation__n7319 , _f_permutation__n7318 ,
         _f_permutation__n7317 , _f_permutation__n7316 ,
         _f_permutation__n7315 , _f_permutation__n7314 ,
         _f_permutation__n7313 , _f_permutation__n7312 ,
         _f_permutation__n7310 , _f_permutation__n7309 ,
         _f_permutation__n7308 , _f_permutation__n7307 ,
         _f_permutation__n7306 , _f_permutation__n7305 ,
         _f_permutation__n7304 , _f_permutation__n7303 ,
         _f_permutation__n7302 , _f_permutation__n7301 ,
         _f_permutation__n7300 , _f_permutation__n7299 ,
         _f_permutation__n7298 , _f_permutation__n7297 ,
         _f_permutation__n7296 , _f_permutation__n7295 ,
         _f_permutation__n7294 , _f_permutation__n7293 ,
         _f_permutation__n7292 , _f_permutation__n7291 ,
         _f_permutation__n7290 , _f_permutation__n7289 ,
         _f_permutation__n7288 , _f_permutation__n7287 ,
         _f_permutation__n7286 , _f_permutation__n7285 ,
         _f_permutation__n7284 , _f_permutation__n7283 ,
         _f_permutation__n7282 , _f_permutation__n7281 ,
         _f_permutation__n7280 , _f_permutation__n7279 ,
         _f_permutation__n7278 , _f_permutation__n7277 ,
         _f_permutation__n7276 , _f_permutation__n7275 ,
         _f_permutation__n7274 , _f_permutation__n7273 ,
         _f_permutation__n7272 , _f_permutation__n7271 ,
         _f_permutation__n7270 , _f_permutation__n7269 ,
         _f_permutation__n7268 , _f_permutation__n7267 ,
         _f_permutation__n7266 , _f_permutation__n7265 ,
         _f_permutation__n7264 , _f_permutation__n7263 ,
         _f_permutation__n7262 , _f_permutation__n7261 ,
         _f_permutation__n7260 , _f_permutation__n7259 ,
         _f_permutation__n7258 , _f_permutation__n7257 ,
         _f_permutation__n7256 , _f_permutation__n7255 ,
         _f_permutation__n7254 , _f_permutation__n7253 ,
         _f_permutation__n7252 , _f_permutation__n7251 ,
         _f_permutation__n7250 , _f_permutation__n7249 ,
         _f_permutation__n7248 , _f_permutation__n7247 ,
         _f_permutation__n7246 , _f_permutation__n7245 ,
         _f_permutation__n7244 , _f_permutation__n7243 ,
         _f_permutation__n7242 , _f_permutation__n7241 ,
         _f_permutation__n7240 , _f_permutation__n7239 ,
         _f_permutation__n7238 , _f_permutation__n7237 ,
         _f_permutation__n7236 , _f_permutation__n7235 ,
         _f_permutation__n7234 , _f_permutation__n7233 ,
         _f_permutation__n7232 , _f_permutation__n7231 ,
         _f_permutation__n7230 , _f_permutation__n7229 ,
         _f_permutation__n7228 , _f_permutation__n7227 ,
         _f_permutation__n7226 , _f_permutation__n7225 ,
         _f_permutation__n7224 , _f_permutation__n7223 ,
         _f_permutation__n7222 , _f_permutation__n7221 ,
         _f_permutation__n7220 , _f_permutation__n7219 ,
         _f_permutation__n7218 , _f_permutation__n7217 ,
         _f_permutation__n7216 , _f_permutation__n7215 ,
         _f_permutation__n7214 , _f_permutation__n7213 ,
         _f_permutation__n7212 , _f_permutation__n7211 ,
         _f_permutation__n7210 , _f_permutation__n7209 ,
         _f_permutation__n7208 , _f_permutation__n7207 ,
         _f_permutation__n7206 , _f_permutation__n7205 ,
         _f_permutation__n7204 , _f_permutation__n7203 ,
         _f_permutation__n7202 , _f_permutation__n7201 ,
         _f_permutation__n7200 , _f_permutation__n7199 ,
         _f_permutation__n7198 , _f_permutation__n7197 ,
         _f_permutation__n7196 , _f_permutation__n7195 ,
         _f_permutation__n7194 , _f_permutation__n7193 ,
         _f_permutation__n7192 , _f_permutation__n7191 ,
         _f_permutation__n7190 , _f_permutation__n7189 ,
         _f_permutation__n7188 , _f_permutation__n7187 ,
         _f_permutation__n7186 , _f_permutation__n7185 ,
         _f_permutation__n7184 , _f_permutation__n7183 ,
         _f_permutation__n7182 , _f_permutation__n7181 ,
         _f_permutation__n7180 , _f_permutation__n7179 ,
         _f_permutation__n7178 , _f_permutation__n7177 ,
         _f_permutation__n7176 , _f_permutation__n7175 ,
         _f_permutation__n7174 , _f_permutation__n7173 ,
         _f_permutation__n7172 , _f_permutation__n7171 ,
         _f_permutation__n7170 , _f_permutation__n7169 ,
         _f_permutation__n7168 , _f_permutation__n7167 ,
         _f_permutation__n7166 , _f_permutation__n7165 ,
         _f_permutation__n7164 , _f_permutation__n7163 ,
         _f_permutation__n7162 , _f_permutation__n7161 ,
         _f_permutation__n7160 , _f_permutation__n7159 ,
         _f_permutation__n7158 , _f_permutation__n7157 ,
         _f_permutation__n7156 , _f_permutation__n7155 ,
         _f_permutation__n7154 , _f_permutation__n7153 ,
         _f_permutation__n7152 , _f_permutation__n7151 ,
         _f_permutation__n7150 , _f_permutation__n7149 ,
         _f_permutation__n7148 , _f_permutation__n7147 ,
         _f_permutation__n7146 , _f_permutation__n7145 ,
         _f_permutation__n7144 , _f_permutation__n7143 ,
         _f_permutation__n7142 , _f_permutation__n7141 ,
         _f_permutation__n7140 , _f_permutation__n7139 ,
         _f_permutation__n7138 , _f_permutation__n7137 ,
         _f_permutation__n7136 , _f_permutation__n7135 ,
         _f_permutation__n7134 , _f_permutation__n7133 ,
         _f_permutation__n7132 , _f_permutation__n7131 ,
         _f_permutation__n7130 , _f_permutation__n7129 ,
         _f_permutation__n7128 , _f_permutation__n7127 ,
         _f_permutation__n7126 , _f_permutation__n7125 ,
         _f_permutation__n7124 , _f_permutation__n7123 ,
         _f_permutation__n7122 , _f_permutation__n7121 ,
         _f_permutation__n7120 , _f_permutation__n7119 ,
         _f_permutation__n7118 , _f_permutation__n7117 ,
         _f_permutation__n7116 , _f_permutation__n7115 ,
         _f_permutation__n7114 , _f_permutation__n7113 ,
         _f_permutation__n7112 , _f_permutation__n7111 ,
         _f_permutation__n7110 , _f_permutation__n7109 ,
         _f_permutation__n7108 , _f_permutation__n7107 ,
         _f_permutation__n7106 , _f_permutation__n7105 ,
         _f_permutation__n7104 , _f_permutation__n7103 ,
         _f_permutation__n7102 , _f_permutation__n7101 ,
         _f_permutation__n7100 , _f_permutation__n7099 ,
         _f_permutation__n7098 , _f_permutation__n7097 ,
         _f_permutation__n7096 , _f_permutation__n7095 ,
         _f_permutation__n7094 , _f_permutation__n7093 ,
         _f_permutation__n7092 , _f_permutation__n7091 ,
         _f_permutation__n7090 , _f_permutation__n7089 ,
         _f_permutation__n7088 , _f_permutation__n7087 ,
         _f_permutation__n7086 , _f_permutation__n7085 ,
         _f_permutation__n7084 , _f_permutation__n7083 ,
         _f_permutation__n7082 , _f_permutation__n7081 ,
         _f_permutation__n7080 , _f_permutation__n7079 ,
         _f_permutation__n7078 , _f_permutation__n7077 ,
         _f_permutation__n7076 , _f_permutation__n7075 ,
         _f_permutation__n7074 , _f_permutation__n7073 ,
         _f_permutation__n7072 , _f_permutation__n7071 ,
         _f_permutation__n7070 , _f_permutation__n7069 ,
         _f_permutation__n7068 , _f_permutation__n7067 ,
         _f_permutation__n7066 , _f_permutation__n7065 ,
         _f_permutation__n7064 , _f_permutation__n7063 ,
         _f_permutation__n7062 , _f_permutation__n7061 ,
         _f_permutation__n7060 , _f_permutation__n7059 ,
         _f_permutation__n7058 , _f_permutation__n7057 ,
         _f_permutation__n7056 , _f_permutation__n7055 ,
         _f_permutation__n7054 , _f_permutation__n7053 ,
         _f_permutation__n7052 , _f_permutation__n7051 ,
         _f_permutation__n7050 , _f_permutation__n7049 ,
         _f_permutation__n7048 , _f_permutation__n7047 ,
         _f_permutation__n7046 , _f_permutation__n7045 ,
         _f_permutation__n7044 , _f_permutation__n7043 ,
         _f_permutation__n7042 , _f_permutation__n7041 ,
         _f_permutation__n7040 , _f_permutation__n7039 ,
         _f_permutation__n7038 , _f_permutation__n7037 ,
         _f_permutation__n7036 , _f_permutation__n7035 ,
         _f_permutation__n7034 , _f_permutation__n7033 ,
         _f_permutation__n7032 , _f_permutation__n7031 ,
         _f_permutation__n7030 , _f_permutation__n7029 ,
         _f_permutation__n7028 , _f_permutation__n7027 ,
         _f_permutation__n7026 , _f_permutation__n7025 ,
         _f_permutation__n7024 , _f_permutation__n7023 ,
         _f_permutation__n7022 , _f_permutation__n7021 ,
         _f_permutation__n7020 , _f_permutation__n7019 ,
         _f_permutation__n7018 , _f_permutation__n7017 ,
         _f_permutation__n7016 , _f_permutation__n7015 ,
         _f_permutation__n7014 , _f_permutation__n7013 ,
         _f_permutation__n7012 , _f_permutation__n7011 ,
         _f_permutation__n7010 , _f_permutation__n7009 ,
         _f_permutation__n7008 , _f_permutation__n7007 ,
         _f_permutation__n7006 , _f_permutation__n7005 ,
         _f_permutation__n7004 , _f_permutation__n7003 ,
         _f_permutation__n7002 , _f_permutation__n7001 ,
         _f_permutation__n7000 , _f_permutation__n6999 ,
         _f_permutation__n6998 , _f_permutation__n6997 ,
         _f_permutation__n6996 , _f_permutation__n6995 ,
         _f_permutation__n6994 , _f_permutation__n6993 ,
         _f_permutation__n6992 , _f_permutation__n6991 ,
         _f_permutation__n6990 , _f_permutation__n6989 ,
         _f_permutation__n6988 , _f_permutation__n6987 ,
         _f_permutation__n6986 , _f_permutation__n6985 ,
         _f_permutation__n6984 , _f_permutation__n6983 ,
         _f_permutation__n6982 , _f_permutation__n6981 ,
         _f_permutation__n6980 , _f_permutation__n6979 ,
         _f_permutation__n6978 , _f_permutation__n6977 ,
         _f_permutation__n6976 , _f_permutation__n6975 ,
         _f_permutation__n6974 , _f_permutation__n6973 ,
         _f_permutation__n6972 , _f_permutation__n6971 ,
         _f_permutation__n6970 , _f_permutation__n6969 ,
         _f_permutation__n6968 , _f_permutation__n6967 ,
         _f_permutation__n6966 , _f_permutation__n6965 ,
         _f_permutation__n6964 , _f_permutation__n6963 ,
         _f_permutation__n6962 , _f_permutation__n6961 ,
         _f_permutation__n6960 , _f_permutation__n6959 ,
         _f_permutation__n6958 , _f_permutation__n6957 ,
         _f_permutation__n6956 , _f_permutation__n6955 ,
         _f_permutation__n6954 , _f_permutation__n6953 ,
         _f_permutation__n6952 , _f_permutation__n6951 ,
         _f_permutation__n6950 , _f_permutation__n6949 ,
         _f_permutation__n6948 , _f_permutation__n6947 ,
         _f_permutation__n6946 , _f_permutation__n6945 ,
         _f_permutation__n6944 , _f_permutation__n6943 ,
         _f_permutation__n6942 , _f_permutation__n6941 ,
         _f_permutation__n6940 , _f_permutation__n6939 ,
         _f_permutation__n6938 , _f_permutation__n6937 ,
         _f_permutation__n6936 , _f_permutation__n6935 ,
         _f_permutation__n6934 , _f_permutation__n6933 ,
         _f_permutation__n6932 , _f_permutation__n6931 ,
         _f_permutation__n6930 , _f_permutation__n6929 ,
         _f_permutation__n6928 , _f_permutation__n6927 ,
         _f_permutation__n6926 , _f_permutation__n6925 ,
         _f_permutation__n6924 , _f_permutation__n6923 ,
         _f_permutation__n6922 , _f_permutation__n6921 ,
         _f_permutation__n6920 , _f_permutation__n6919 ,
         _f_permutation__n6918 , _f_permutation__n6917 ,
         _f_permutation__n6916 , _f_permutation__n6915 ,
         _f_permutation__n6914 , _f_permutation__n6913 ,
         _f_permutation__n6912 , _f_permutation__n6911 ,
         _f_permutation__n6910 , _f_permutation__n6909 ,
         _f_permutation__n6908 , _f_permutation__n6907 ,
         _f_permutation__n6906 , _f_permutation__n6905 ,
         _f_permutation__n6904 , _f_permutation__n6903 ,
         _f_permutation__n6902 , _f_permutation__n6901 ,
         _f_permutation__n6900 , _f_permutation__n6899 ,
         _f_permutation__n6898 , _f_permutation__n6897 ,
         _f_permutation__n6896 , _f_permutation__n6895 ,
         _f_permutation__n6894 , _f_permutation__n6893 ,
         _f_permutation__n6892 , _f_permutation__n6891 ,
         _f_permutation__n6890 , _f_permutation__n6889 ,
         _f_permutation__n6888 , _f_permutation__n6887 ,
         _f_permutation__n6886 , _f_permutation__n6885 ,
         _f_permutation__n6884 , _f_permutation__n6883 ,
         _f_permutation__n6882 , _f_permutation__n6881 ,
         _f_permutation__n6880 , _f_permutation__n6879 ,
         _f_permutation__n6878 , _f_permutation__n6877 ,
         _f_permutation__n6876 , _f_permutation__n6875 ,
         _f_permutation__n6874 , _f_permutation__n6873 ,
         _f_permutation__n6872 , _f_permutation__n6871 ,
         _f_permutation__n6870 , _f_permutation__n6869 ,
         _f_permutation__n6868 , _f_permutation__n6867 ,
         _f_permutation__n6866 , _f_permutation__n6865 ,
         _f_permutation__n6864 , _f_permutation__n6863 ,
         _f_permutation__n6862 , _f_permutation__n6861 ,
         _f_permutation__n6860 , _f_permutation__n6859 ,
         _f_permutation__n6858 , _f_permutation__n6857 ,
         _f_permutation__n6856 , _f_permutation__n6855 ,
         _f_permutation__n6854 , _f_permutation__n6853 ,
         _f_permutation__n6852 , _f_permutation__n6851 ,
         _f_permutation__n6850 , _f_permutation__n6849 ,
         _f_permutation__n6848 , _f_permutation__n6847 ,
         _f_permutation__n6846 , _f_permutation__n6845 ,
         _f_permutation__n6844 , _f_permutation__n6843 ,
         _f_permutation__n6842 , _f_permutation__n6841 ,
         _f_permutation__n6840 , _f_permutation__n6839 ,
         _f_permutation__n6838 , _f_permutation__n6837 ,
         _f_permutation__n6836 , _f_permutation__n6835 ,
         _f_permutation__n6834 , _f_permutation__n6833 ,
         _f_permutation__n6832 , _f_permutation__n6831 ,
         _f_permutation__n6830 , _f_permutation__n6829 ,
         _f_permutation__n6828 , _f_permutation__n6827 ,
         _f_permutation__n6826 , _f_permutation__n6825 ,
         _f_permutation__n6824 , _f_permutation__n6823 ,
         _f_permutation__n6822 , _f_permutation__n6821 ,
         _f_permutation__n6820 , _f_permutation__n6819 ,
         _f_permutation__n6818 , _f_permutation__n6817 ,
         _f_permutation__n6816 , _f_permutation__n6815 ,
         _f_permutation__n6814 , _f_permutation__n6813 ,
         _f_permutation__n6812 , _f_permutation__n6811 ,
         _f_permutation__n6810 , _f_permutation__n6809 ,
         _f_permutation__n6808 , _f_permutation__n6807 ,
         _f_permutation__n6806 , _f_permutation__n6805 ,
         _f_permutation__n6804 , _f_permutation__n6803 ,
         _f_permutation__n6802 , _f_permutation__n6801 ,
         _f_permutation__n6800 , _f_permutation__n6799 ,
         _f_permutation__n6798 , _f_permutation__n6797 ,
         _f_permutation__n6796 , _f_permutation__n6795 ,
         _f_permutation__n6794 , _f_permutation__n6793 ,
         _f_permutation__n6792 , _f_permutation__n6791 ,
         _f_permutation__n6790 , _f_permutation__n6789 ,
         _f_permutation__n6788 , _f_permutation__n6787 ,
         _f_permutation__n6786 , _f_permutation__n6785 ,
         _f_permutation__n6784 , _f_permutation__n6783 ,
         _f_permutation__n6782 , _f_permutation__n6781 ,
         _f_permutation__n6780 , _f_permutation__n6779 ,
         _f_permutation__n6778 , _f_permutation__n6777 ,
         _f_permutation__n6776 , _f_permutation__n6775 ,
         _f_permutation__n6774 , _f_permutation__n6773 ,
         _f_permutation__n6772 , _f_permutation__n6771 ,
         _f_permutation__n6770 , _f_permutation__n6769 ,
         _f_permutation__n6768 , _f_permutation__n6767 ,
         _f_permutation__n6766 , _f_permutation__n6765 ,
         _f_permutation__n6764 , _f_permutation__n6763 ,
         _f_permutation__n6762 , _f_permutation__n6761 ,
         _f_permutation__n6760 , _f_permutation__n6759 ,
         _f_permutation__n6758 , _f_permutation__n6757 ,
         _f_permutation__n6756 , _f_permutation__n6755 ,
         _f_permutation__n6754 , _f_permutation__n6753 ,
         _f_permutation__n6752 , _f_permutation__n6751 ,
         _f_permutation__n6750 , _f_permutation__n6749 ,
         _f_permutation__n6748 , _f_permutation__n6747 ,
         _f_permutation__n6746 , _f_permutation__n6745 ,
         _f_permutation__n6744 , _f_permutation__n6743 ,
         _f_permutation__n6742 , _f_permutation__n6741 ,
         _f_permutation__n6740 , _f_permutation__n6739 ,
         _f_permutation__n6738 , _f_permutation__n6737 ,
         _f_permutation__n6736 , _f_permutation__n6735 ,
         _f_permutation__n6734 , _f_permutation__n6733 ,
         _f_permutation__n6732 , _f_permutation__n6731 ,
         _f_permutation__n6730 , _f_permutation__n6729 ,
         _f_permutation__n6728 , _f_permutation__n6727 ,
         _f_permutation__n6726 , _f_permutation__n6725 ,
         _f_permutation__n6724 , _f_permutation__n6723 ,
         _f_permutation__n6722 , _f_permutation__n6721 ,
         _f_permutation__n6720 , _f_permutation__n6719 ,
         _f_permutation__n6718 , _f_permutation__n6717 ,
         _f_permutation__n6716 , _f_permutation__n6715 ,
         _f_permutation__n6714 , _f_permutation__n6713 ,
         _f_permutation__n6712 , _f_permutation__n6711 ,
         _f_permutation__n6710 , _f_permutation__n6709 ,
         _f_permutation__n6708 , _f_permutation__n6707 ,
         _f_permutation__n6706 , _f_permutation__n6705 ,
         _f_permutation__n6704 , _f_permutation__n6703 ,
         _f_permutation__n6702 , _f_permutation__n6701 ,
         _f_permutation__n6700 , _f_permutation__n6699 ,
         _f_permutation__n6698 , _f_permutation__n6697 ,
         _f_permutation__n6696 , _f_permutation__n6695 ,
         _f_permutation__n6694 , _f_permutation__n6693 ,
         _f_permutation__n6692 , _f_permutation__n6691 ,
         _f_permutation__n6690 , _f_permutation__n6689 ,
         _f_permutation__n6688 , _f_permutation__n6687 ,
         _f_permutation__n6686 , _f_permutation__n6685 ,
         _f_permutation__n6684 , _f_permutation__n6683 ,
         _f_permutation__n6682 , _f_permutation__n6681 ,
         _f_permutation__n6680 , _f_permutation__n6679 ,
         _f_permutation__n6678 , _f_permutation__n6677 ,
         _f_permutation__n6676 , _f_permutation__n6675 ,
         _f_permutation__n6674 , _f_permutation__n6673 ,
         _f_permutation__n6672 , _f_permutation__n6671 ,
         _f_permutation__n6670 , _f_permutation__n6669 ,
         _f_permutation__n6668 , _f_permutation__n6667 ,
         _f_permutation__n6666 , _f_permutation__n6665 ,
         _f_permutation__n6664 , _f_permutation__n6663 ,
         _f_permutation__n6662 , _f_permutation__n6661 ,
         _f_permutation__n6660 , _f_permutation__n6659 ,
         _f_permutation__n6658 , _f_permutation__n6657 ,
         _f_permutation__n6656 , _f_permutation__n6655 ,
         _f_permutation__n6654 , _f_permutation__n6653 ,
         _f_permutation__n6652 , _f_permutation__n6651 ,
         _f_permutation__n6650 , _f_permutation__n6649 ,
         _f_permutation__n6648 , _f_permutation__n6647 ,
         _f_permutation__n6646 , _f_permutation__n6645 ,
         _f_permutation__n6644 , _f_permutation__n6643 ,
         _f_permutation__n6642 , _f_permutation__n6641 ,
         _f_permutation__n6640 , _f_permutation__n6639 ,
         _f_permutation__n6638 , _f_permutation__n6637 ,
         _f_permutation__n6636 , _f_permutation__n6635 ,
         _f_permutation__n6634 , _f_permutation__n6633 ,
         _f_permutation__n6632 , _f_permutation__n6631 ,
         _f_permutation__n6630 , _f_permutation__n6629 ,
         _f_permutation__n6628 , _f_permutation__n6627 ,
         _f_permutation__n6626 , _f_permutation__n6625 ,
         _f_permutation__n6624 , _f_permutation__n6623 ,
         _f_permutation__n6622 , _f_permutation__n6621 ,
         _f_permutation__n6620 , _f_permutation__n6619 ,
         _f_permutation__n6618 , _f_permutation__n6617 ,
         _f_permutation__n6616 , _f_permutation__n6615 ,
         _f_permutation__n6614 , _f_permutation__n6613 ,
         _f_permutation__n6612 , _f_permutation__n6611 ,
         _f_permutation__n6610 , _f_permutation__n6609 ,
         _f_permutation__n6608 , _f_permutation__n6607 ,
         _f_permutation__n6606 , _f_permutation__n6605 ,
         _f_permutation__n6604 , _f_permutation__n6603 ,
         _f_permutation__n6602 , _f_permutation__n6601 ,
         _f_permutation__n6600 , _f_permutation__n6599 ,
         _f_permutation__n6598 , _f_permutation__n6597 ,
         _f_permutation__n6596 , _f_permutation__n6595 ,
         _f_permutation__n6594 , _f_permutation__n6593 ,
         _f_permutation__n6592 , _f_permutation__n6591 ,
         _f_permutation__n6590 , _f_permutation__n6589 ,
         _f_permutation__n6588 , _f_permutation__n6587 ,
         _f_permutation__n6586 , _f_permutation__n6585 ,
         _f_permutation__n6584 , _f_permutation__n6583 ,
         _f_permutation__n6582 , _f_permutation__n6581 ,
         _f_permutation__n6580 , _f_permutation__n6579 ,
         _f_permutation__n6578 , _f_permutation__n6577 ,
         _f_permutation__n6576 , _f_permutation__n6575 ,
         _f_permutation__n6574 , _f_permutation__n6573 ,
         _f_permutation__n6572 , _f_permutation__n6571 ,
         _f_permutation__n6570 , _f_permutation__n6569 ,
         _f_permutation__n6568 , _f_permutation__n6567 ,
         _f_permutation__n6566 , _f_permutation__n6565 ,
         _f_permutation__n6564 , _f_permutation__n6563 ,
         _f_permutation__n6562 , _f_permutation__n6561 ,
         _f_permutation__n6560 , _f_permutation__n6559 ,
         _f_permutation__n6558 , _f_permutation__n6557 ,
         _f_permutation__n6556 , _f_permutation__n6555 ,
         _f_permutation__n6554 , _f_permutation__n6553 ,
         _f_permutation__n6552 , _f_permutation__n6551 ,
         _f_permutation__n6550 , _f_permutation__n6549 ,
         _f_permutation__n6548 , _f_permutation__n6547 ,
         _f_permutation__n6546 , _f_permutation__n6545 ,
         _f_permutation__n6544 , _f_permutation__n6543 ,
         _f_permutation__n6542 , _f_permutation__n6541 ,
         _f_permutation__n6540 , _f_permutation__n6539 ,
         _f_permutation__n6538 , _f_permutation__n6537 ,
         _f_permutation__n6536 , _f_permutation__n6535 ,
         _f_permutation__n6534 , _f_permutation__n6533 ,
         _f_permutation__n6532 , _f_permutation__n6531 ,
         _f_permutation__n6530 , _f_permutation__n6529 ,
         _f_permutation__n6528 , _f_permutation__n6527 ,
         _f_permutation__n6526 , _f_permutation__n6525 ,
         _f_permutation__n6524 , _f_permutation__n6523 ,
         _f_permutation__n6522 , _f_permutation__n6521 ,
         _f_permutation__n6520 , _f_permutation__n6519 ,
         _f_permutation__n6518 , _f_permutation__n6517 ,
         _f_permutation__n6516 , _f_permutation__n6515 ,
         _f_permutation__n6514 , _f_permutation__n6513 ,
         _f_permutation__n6512 , _f_permutation__n6511 ,
         _f_permutation__n6510 , _f_permutation__n6509 ,
         _f_permutation__n6508 , _f_permutation__n6507 ,
         _f_permutation__n6506 , _f_permutation__n6505 ,
         _f_permutation__n6504 , _f_permutation__n6503 ,
         _f_permutation__n6502 , _f_permutation__n6501 ,
         _f_permutation__n6500 , _f_permutation__n6499 ,
         _f_permutation__n6498 , _f_permutation__n6497 ,
         _f_permutation__n6496 , _f_permutation__n6495 ,
         _f_permutation__n6494 , _f_permutation__n6493 ,
         _f_permutation__n6492 , _f_permutation__n6491 ,
         _f_permutation__n6490 , _f_permutation__n6489 ,
         _f_permutation__n6488 , _f_permutation__n6487 ,
         _f_permutation__n6486 , _f_permutation__n6485 ,
         _f_permutation__n6484 , _f_permutation__n6483 ,
         _f_permutation__n6482 , _f_permutation__n6481 ,
         _f_permutation__n6480 , _f_permutation__n6479 ,
         _f_permutation__n6478 , _f_permutation__n6477 ,
         _f_permutation__n6476 , _f_permutation__n6475 ,
         _f_permutation__n6474 , _f_permutation__n6473 ,
         _f_permutation__n6472 , _f_permutation__n6471 ,
         _f_permutation__n6470 , _f_permutation__n6469 ,
         _f_permutation__n6468 , _f_permutation__n6467 ,
         _f_permutation__n6466 , _f_permutation__n6465 ,
         _f_permutation__n6464 , _f_permutation__n6463 ,
         _f_permutation__n6462 , _f_permutation__n6461 ,
         _f_permutation__n6460 , _f_permutation__n6459 ,
         _f_permutation__n6458 , _f_permutation__n6457 ,
         _f_permutation__n6456 , _f_permutation__n6455 ,
         _f_permutation__n6454 , _f_permutation__n6453 ,
         _f_permutation__n6452 , _f_permutation__n6451 ,
         _f_permutation__n6450 , _f_permutation__n6449 ,
         _f_permutation__n6448 , _f_permutation__n6447 ,
         _f_permutation__n6446 , _f_permutation__n6445 ,
         _f_permutation__n6444 , _f_permutation__n6443 ,
         _f_permutation__n6442 , _f_permutation__n6441 ,
         _f_permutation__n6440 , _f_permutation__n6439 ,
         _f_permutation__n6438 , _f_permutation__n6437 ,
         _f_permutation__n6436 , _f_permutation__n6435 ,
         _f_permutation__n6434 , _f_permutation__n6433 ,
         _f_permutation__n6432 , _f_permutation__n6431 ,
         _f_permutation__n6430 , _f_permutation__n6429 ,
         _f_permutation__n6428 , _f_permutation__n6427 ,
         _f_permutation__n6426 , _f_permutation__n6425 ,
         _f_permutation__n6424 , _f_permutation__n6423 ,
         _f_permutation__n6422 , _f_permutation__n6421 ,
         _f_permutation__n6420 , _f_permutation__n6419 ,
         _f_permutation__n6418 , _f_permutation__n6417 ,
         _f_permutation__n6416 , _f_permutation__n6415 ,
         _f_permutation__n6414 , _f_permutation__n6413 ,
         _f_permutation__n6412 , _f_permutation__n6411 ,
         _f_permutation__n6410 , _f_permutation__n6409 ,
         _f_permutation__n6408 , _f_permutation__n6407 ,
         _f_permutation__n6406 , _f_permutation__n6405 ,
         _f_permutation__n6404 , _f_permutation__n6403 ,
         _f_permutation__n6402 , _f_permutation__n6401 ,
         _f_permutation__n6400 , _f_permutation__n6399 ,
         _f_permutation__n6398 , _f_permutation__n6397 ,
         _f_permutation__n6396 , _f_permutation__n6395 ,
         _f_permutation__n6394 , _f_permutation__n6393 ,
         _f_permutation__n6392 , _f_permutation__n6391 ,
         _f_permutation__n6390 , _f_permutation__n6389 ,
         _f_permutation__n6388 , _f_permutation__n6387 ,
         _f_permutation__n6386 , _f_permutation__n6385 ,
         _f_permutation__n6384 , _f_permutation__n6383 ,
         _f_permutation__n6382 , _f_permutation__n6381 ,
         _f_permutation__n6380 , _f_permutation__n6379 ,
         _f_permutation__n6378 , _f_permutation__n6377 ,
         _f_permutation__n6376 , _f_permutation__n6375 ,
         _f_permutation__n6374 , _f_permutation__n6373 ,
         _f_permutation__n6372 , _f_permutation__n6371 ,
         _f_permutation__n6370 , _f_permutation__n6369 ,
         _f_permutation__n6368 , _f_permutation__n6367 ,
         _f_permutation__n6366 , _f_permutation__n6365 ,
         _f_permutation__n6364 , _f_permutation__n6363 ,
         _f_permutation__n6362 , _f_permutation__n6361 ,
         _f_permutation__n6360 , _f_permutation__n6359 ,
         _f_permutation__n6358 , _f_permutation__n6357 ,
         _f_permutation__n6356 , _f_permutation__n6355 ,
         _f_permutation__n6354 , _f_permutation__n6353 ,
         _f_permutation__n6352 , _f_permutation__n6351 ,
         _f_permutation__n6350 , _f_permutation__n6349 ,
         _f_permutation__n6348 , _f_permutation__n6347 ,
         _f_permutation__n6346 , _f_permutation__n6345 ,
         _f_permutation__n6344 , _f_permutation__n6343 ,
         _f_permutation__n6342 , _f_permutation__n6341 ,
         _f_permutation__n6340 , _f_permutation__n6339 ,
         _f_permutation__n6338 , _f_permutation__n6337 ,
         _f_permutation__n6336 , _f_permutation__n6335 ,
         _f_permutation__n6334 , _f_permutation__n6333 ,
         _f_permutation__n6332 , _f_permutation__n6331 ,
         _f_permutation__n6330 , _f_permutation__n6329 ,
         _f_permutation__n6328 , _f_permutation__n6327 ,
         _f_permutation__n6326 , _f_permutation__n6325 ,
         _f_permutation__n6324 , _f_permutation__n6323 ,
         _f_permutation__n6322 , _f_permutation__n6321 ,
         _f_permutation__n6320 , _f_permutation__n6319 ,
         _f_permutation__n6318 , _f_permutation__n6317 ,
         _f_permutation__n6316 , _f_permutation__n6315 ,
         _f_permutation__n6314 , _f_permutation__n6313 ,
         _f_permutation__n6312 , _f_permutation__n6311 ,
         _f_permutation__n6310 , _f_permutation__n6309 ,
         _f_permutation__n6308 , _f_permutation__n6307 ,
         _f_permutation__n6306 , _f_permutation__n6305 ,
         _f_permutation__n6304 , _f_permutation__n6303 ,
         _f_permutation__n6302 , _f_permutation__n6301 ,
         _f_permutation__n6300 , _f_permutation__n6299 ,
         _f_permutation__n6298 , _f_permutation__n6297 ,
         _f_permutation__n6296 , _f_permutation__n6295 ,
         _f_permutation__n6294 , _f_permutation__n6293 ,
         _f_permutation__n6292 , _f_permutation__n6291 ,
         _f_permutation__n6290 , _f_permutation__n6289 ,
         _f_permutation__n6288 , _f_permutation__n6287 ,
         _f_permutation__n6286 , _f_permutation__n6285 ,
         _f_permutation__n6284 , _f_permutation__n6283 ,
         _f_permutation__n6282 , _f_permutation__n6281 ,
         _f_permutation__n6280 , _f_permutation__n6279 ,
         _f_permutation__n6278 , _f_permutation__n6277 ,
         _f_permutation__n6276 , _f_permutation__n6275 ,
         _f_permutation__n6274 , _f_permutation__n6273 ,
         _f_permutation__n6272 , _f_permutation__n6271 ,
         _f_permutation__n6270 , _f_permutation__n6269 ,
         _f_permutation__n6268 , _f_permutation__n6267 ,
         _f_permutation__n6266 , _f_permutation__n6265 ,
         _f_permutation__n6264 , _f_permutation__n6263 ,
         _f_permutation__n6262 , _f_permutation__n6261 ,
         _f_permutation__n6260 , _f_permutation__n6259 ,
         _f_permutation__n6258 , _f_permutation__n6257 ,
         _f_permutation__n6256 , _f_permutation__n6255 ,
         _f_permutation__n6254 , _f_permutation__n6253 ,
         _f_permutation__n6252 , _f_permutation__n6251 ,
         _f_permutation__n6250 , _f_permutation__n6249 ,
         _f_permutation__n6248 , _f_permutation__n6247 ,
         _f_permutation__n6246 , _f_permutation__n6245 ,
         _f_permutation__n6244 , _f_permutation__n6243 ,
         _f_permutation__n6242 , _f_permutation__n6241 ,
         _f_permutation__n6240 , _f_permutation__n6239 ,
         _f_permutation__n6238 , _f_permutation__n6237 ,
         _f_permutation__n6236 , _f_permutation__n6235 ,
         _f_permutation__n6234 , _f_permutation__n6233 ,
         _f_permutation__n6232 , _f_permutation__n6231 ,
         _f_permutation__n6230 , _f_permutation__n6229 ,
         _f_permutation__n6228 , _f_permutation__n6227 ,
         _f_permutation__n6226 , _f_permutation__n6225 ,
         _f_permutation__n6224 , _f_permutation__n6223 ,
         _f_permutation__n6222 , _f_permutation__n6221 ,
         _f_permutation__n6220 , _f_permutation__n6219 ,
         _f_permutation__n6218 , _f_permutation__n6217 ,
         _f_permutation__n6216 , _f_permutation__n6215 ,
         _f_permutation__n6214 , _f_permutation__n6213 ,
         _f_permutation__n6212 , _f_permutation__n6211 ,
         _f_permutation__n6210 , _f_permutation__n6209 ,
         _f_permutation__n6208 , _f_permutation__n6207 ,
         _f_permutation__n6206 , _f_permutation__n6205 ,
         _f_permutation__n6204 , _f_permutation__n6203 ,
         _f_permutation__n6202 , _f_permutation__n6201 ,
         _f_permutation__n6200 , _f_permutation__n6199 ,
         _f_permutation__n6198 , _f_permutation__n6197 ,
         _f_permutation__n6196 , _f_permutation__n6195 ,
         _f_permutation__n6194 , _f_permutation__n6193 ,
         _f_permutation__n6192 , _f_permutation__n6191 ,
         _f_permutation__n6190 , _f_permutation__n6189 ,
         _f_permutation__n6188 , _f_permutation__n6187 ,
         _f_permutation__n6186 , _f_permutation__n6185 ,
         _f_permutation__n6184 , _f_permutation__n6183 ,
         _f_permutation__n6182 , _f_permutation__n6181 ,
         _f_permutation__n6180 , _f_permutation__n6179 ,
         _f_permutation__n6178 , _f_permutation__n6177 ,
         _f_permutation__n6176 , _f_permutation__n6175 ,
         _f_permutation__n6174 , _f_permutation__n6173 ,
         _f_permutation__n6172 , _f_permutation__n6171 ,
         _f_permutation__n6170 , _f_permutation__n6169 ,
         _f_permutation__n6168 , _f_permutation__n6167 ,
         _f_permutation__n6166 , _f_permutation__n6165 ,
         _f_permutation__n6164 , _f_permutation__n6163 ,
         _f_permutation__n6162 , _f_permutation__n6161 ,
         _f_permutation__n6160 , _f_permutation__n6159 ,
         _f_permutation__n6158 , _f_permutation__n6157 ,
         _f_permutation__n6156 , _f_permutation__n6155 ,
         _f_permutation__n6154 , _f_permutation__n6153 ,
         _f_permutation__n6152 , _f_permutation__n6151 ,
         _f_permutation__n6150 , _f_permutation__n6149 ,
         _f_permutation__n6148 , _f_permutation__n6147 ,
         _f_permutation__n6146 , _f_permutation__n6145 ,
         _f_permutation__n6144 , _f_permutation__n6143 ,
         _f_permutation__n6142 , _f_permutation__n6141 ,
         _f_permutation__n6140 , _f_permutation__n6139 ,
         _f_permutation__n6138 , _f_permutation__n6137 ,
         _f_permutation__n6136 , _f_permutation__n6135 ,
         _f_permutation__n6134 , _f_permutation__n6133 ,
         _f_permutation__n6132 , _f_permutation__n6131 ,
         _f_permutation__n6130 , _f_permutation__n6129 ,
         _f_permutation__n6128 , _f_permutation__n6127 ,
         _f_permutation__n6126 , _f_permutation__n6125 ,
         _f_permutation__n6124 , _f_permutation__n6123 ,
         _f_permutation__n6122 , _f_permutation__n6121 ,
         _f_permutation__n6120 , _f_permutation__n6119 ,
         _f_permutation__n6118 , _f_permutation__n6117 ,
         _f_permutation__n6116 , _f_permutation__n6115 ,
         _f_permutation__n6114 , _f_permutation__n6113 ,
         _f_permutation__n6112 , _f_permutation__n6111 ,
         _f_permutation__n6110 , _f_permutation__n6109 ,
         _f_permutation__n6108 , _f_permutation__n6107 ,
         _f_permutation__n6106 , _f_permutation__n6105 ,
         _f_permutation__n6104 , _f_permutation__n6103 ,
         _f_permutation__n6102 , _f_permutation__n6101 ,
         _f_permutation__n6100 , _f_permutation__n6099 ,
         _f_permutation__n6098 , _f_permutation__n6097 ,
         _f_permutation__n6096 , _f_permutation__n6095 ,
         _f_permutation__n6094 , _f_permutation__n6093 ,
         _f_permutation__n6092 , _f_permutation__n6091 ,
         _f_permutation__n6090 , _f_permutation__n6089 ,
         _f_permutation__n6088 , _f_permutation__n6087 ,
         _f_permutation__n6086 , _f_permutation__n6085 ,
         _f_permutation__n6084 , _f_permutation__n6083 ,
         _f_permutation__n6082 , _f_permutation__n6081 ,
         _f_permutation__n6080 , _f_permutation__n6079 ,
         _f_permutation__n6078 , _f_permutation__n6077 ,
         _f_permutation__n6076 , _f_permutation__n6075 ,
         _f_permutation__n6074 , _f_permutation__n6073 ,
         _f_permutation__n6072 , _f_permutation__n6071 ,
         _f_permutation__n6070 , _f_permutation__n6069 ,
         _f_permutation__n6068 , _f_permutation__n6067 ,
         _f_permutation__n6066 , _f_permutation__n6065 ,
         _f_permutation__n6064 , _f_permutation__n6063 ,
         _f_permutation__n6062 , _f_permutation__n6061 ,
         _f_permutation__n6060 , _f_permutation__n6059 ,
         _f_permutation__n6058 , _f_permutation__n6057 ,
         _f_permutation__n6056 , _f_permutation__n6055 ,
         _f_permutation__n6054 , _f_permutation__n6053 ,
         _f_permutation__n6052 , _f_permutation__n6051 ,
         _f_permutation__n6050 , _f_permutation__n6049 ,
         _f_permutation__n6048 , _f_permutation__n6047 ,
         _f_permutation__n6046 , _f_permutation__n6045 ,
         _f_permutation__n6044 , _f_permutation__n6043 ,
         _f_permutation__n6042 , _f_permutation__n6041 ,
         _f_permutation__n6040 , _f_permutation__n6039 ,
         _f_permutation__n6038 , _f_permutation__n6037 ,
         _f_permutation__n6036 , _f_permutation__n6035 ,
         _f_permutation__n6034 , _f_permutation__n6033 ,
         _f_permutation__n6032 , _f_permutation__n6031 ,
         _f_permutation__n6030 , _f_permutation__n6029 ,
         _f_permutation__n6028 , _f_permutation__n6027 ,
         _f_permutation__n6026 , _f_permutation__n6025 ,
         _f_permutation__n6024 , _f_permutation__n6023 ,
         _f_permutation__n6022 , _f_permutation__n6021 ,
         _f_permutation__n6020 , _f_permutation__n6019 ,
         _f_permutation__n6018 , _f_permutation__n6017 ,
         _f_permutation__n6016 , _f_permutation__n6015 ,
         _f_permutation__n6014 , _f_permutation__n6013 ,
         _f_permutation__n6012 , _f_permutation__n6011 ,
         _f_permutation__n6010 , _f_permutation__n6009 ,
         _f_permutation__n6008 , _f_permutation__n6007 ,
         _f_permutation__n6006 , _f_permutation__n6005 ,
         _f_permutation__n6004 , _f_permutation__n6003 ,
         _f_permutation__n6002 , _f_permutation__n6001 ,
         _f_permutation__n6000 , _f_permutation__n5999 ,
         _f_permutation__n5998 , _f_permutation__n5997 ,
         _f_permutation__n5996 , _f_permutation__n5995 ,
         _f_permutation__n5994 , _f_permutation__n5993 ,
         _f_permutation__n5992 , _f_permutation__n5991 ,
         _f_permutation__n5990 , _f_permutation__n5989 ,
         _f_permutation__n5988 , _f_permutation__n5987 ,
         _f_permutation__n5986 , _f_permutation__n5985 ,
         _f_permutation__n5984 , _f_permutation__n5983 ,
         _f_permutation__n5982 , _f_permutation__n5981 ,
         _f_permutation__n5980 , _f_permutation__n5979 ,
         _f_permutation__n5978 , _f_permutation__n5977 ,
         _f_permutation__n5976 , _f_permutation__n5975 ,
         _f_permutation__n5974 , _f_permutation__n5973 ,
         _f_permutation__n5972 , _f_permutation__n5971 ,
         _f_permutation__n5970 , _f_permutation__n5969 ,
         _f_permutation__n5968 , _f_permutation__n5967 ,
         _f_permutation__n5966 , _f_permutation__n5965 ,
         _f_permutation__n5964 , _f_permutation__n5963 ,
         _f_permutation__n5962 , _f_permutation__n5961 ,
         _f_permutation__n5960 , _f_permutation__n5959 ,
         _f_permutation__n5958 , _f_permutation__n5957 ,
         _f_permutation__n5956 , _f_permutation__n5955 ,
         _f_permutation__n5954 , _f_permutation__n5953 ,
         _f_permutation__n5952 , _f_permutation__n5951 ,
         _f_permutation__n5950 , _f_permutation__n5949 ,
         _f_permutation__n5948 , _f_permutation__n5947 ,
         _f_permutation__n5946 , _f_permutation__n5945 ,
         _f_permutation__n5944 , _f_permutation__n5943 ,
         _f_permutation__n5942 , _f_permutation__n5941 ,
         _f_permutation__n5940 , _f_permutation__n5939 ,
         _f_permutation__n5938 , _f_permutation__n5937 ,
         _f_permutation__n5936 , _f_permutation__n5935 ,
         _f_permutation__n5934 , _f_permutation__n5933 ,
         _f_permutation__n5932 , _f_permutation__n5931 ,
         _f_permutation__n5930 , _f_permutation__n5929 ,
         _f_permutation__n5928 , _f_permutation__n5927 ,
         _f_permutation__n5926 , _f_permutation__n5925 ,
         _f_permutation__n5924 , _f_permutation__n5923 ,
         _f_permutation__n5922 , _f_permutation__n5921 ,
         _f_permutation__n5920 , _f_permutation__n5919 ,
         _f_permutation__n5918 , _f_permutation__n5917 ,
         _f_permutation__n5916 , _f_permutation__n5915 ,
         _f_permutation__n5914 , _f_permutation__n5913 ,
         _f_permutation__n5912 , _f_permutation__n5911 ,
         _f_permutation__n5910 , _f_permutation__n5909 ,
         _f_permutation__n5908 , _f_permutation__n5907 ,
         _f_permutation__n5906 , _f_permutation__n5905 ,
         _f_permutation__n5904 , _f_permutation__n5903 ,
         _f_permutation__n5902 , _f_permutation__n5901 ,
         _f_permutation__n5900 , _f_permutation__n5899 ,
         _f_permutation__n5898 , _f_permutation__n5897 ,
         _f_permutation__n5896 , _f_permutation__n5895 ,
         _f_permutation__n5894 , _f_permutation__n5893 ,
         _f_permutation__n5892 , _f_permutation__n5891 ,
         _f_permutation__n5890 , _f_permutation__n5889 ,
         _f_permutation__n5888 , _f_permutation__n5887 ,
         _f_permutation__n5886 , _f_permutation__n5885 ,
         _f_permutation__n5884 , _f_permutation__n5883 ,
         _f_permutation__n5882 , _f_permutation__n5881 ,
         _f_permutation__n5880 , _f_permutation__n5879 ,
         _f_permutation__n5878 , _f_permutation__n5877 ,
         _f_permutation__n5876 , _f_permutation__n5875 ,
         _f_permutation__n5874 , _f_permutation__n5873 ,
         _f_permutation__n5872 , _f_permutation__n5871 ,
         _f_permutation__n5870 , _f_permutation__n5869 ,
         _f_permutation__n5868 , _f_permutation__n5867 ,
         _f_permutation__n5866 , _f_permutation__n5865 ,
         _f_permutation__n5864 , _f_permutation__n5863 ,
         _f_permutation__n5862 , _f_permutation__n5861 ,
         _f_permutation__n5860 , _f_permutation__n5859 ,
         _f_permutation__n5858 , _f_permutation__n5857 ,
         _f_permutation__n5856 , _f_permutation__n5855 ,
         _f_permutation__n5854 , _f_permutation__n5853 ,
         _f_permutation__n5852 , _f_permutation__n5851 ,
         _f_permutation__n5850 , _f_permutation__n5849 ,
         _f_permutation__n5848 , _f_permutation__n5847 ,
         _f_permutation__n5846 , _f_permutation__n5845 ,
         _f_permutation__n5844 , _f_permutation__n5843 ,
         _f_permutation__n5842 , _f_permutation__n5841 ,
         _f_permutation__n5840 , _f_permutation__n5839 ,
         _f_permutation__n5838 , _f_permutation__n5837 ,
         _f_permutation__n5836 , _f_permutation__n5835 ,
         _f_permutation__n5834 , _f_permutation__n5833 ,
         _f_permutation__n5832 , _f_permutation__n5831 ,
         _f_permutation__n5830 , _f_permutation__n5829 ,
         _f_permutation__n5828 , _f_permutation__n5827 ,
         _f_permutation__n5826 , _f_permutation__n5825 ,
         _f_permutation__n5824 , _f_permutation__n5823 ,
         _f_permutation__n5822 , _f_permutation__n5821 ,
         _f_permutation__n5820 , _f_permutation__n5819 ,
         _f_permutation__n5818 , _f_permutation__n5817 ,
         _f_permutation__n5816 , _f_permutation__n5815 ,
         _f_permutation__n5814 , _f_permutation__n5813 ,
         _f_permutation__n5812 , _f_permutation__n5811 ,
         _f_permutation__n5810 , _f_permutation__n5809 ,
         _f_permutation__n5808 , _f_permutation__n5807 ,
         _f_permutation__n5806 , _f_permutation__n5781 ,
         _f_permutation__n5780 , _f_permutation__n5779 ,
         _f_permutation__n5778 , _f_permutation__n5777 ,
         _f_permutation__n5776 , _f_permutation__n5775 ,
         _f_permutation__n5774 , _f_permutation__n5773 ,
         _f_permutation__n5772 , _f_permutation__n5771 ,
         _f_permutation__n5770 , _f_permutation__n5769 ,
         _f_permutation__n5768 , _f_permutation__n5767 ,
         _f_permutation__n5766 , _f_permutation__n5765 ,
         _f_permutation__n5764 , _f_permutation__n5763 ,
         _f_permutation__n5762 , _f_permutation__n5761 ,
         _f_permutation__n5760 , _f_permutation__n5759 ,
         _f_permutation__n5758 , _f_permutation__n5757 ,
         _f_permutation__n5756 , _f_permutation__n5755 ,
         _f_permutation__n5754 , _f_permutation__n5753 ,
         _f_permutation__n5752 , _f_permutation__n5751 ,
         _f_permutation__n5750 , _f_permutation__n5749 ,
         _f_permutation__n5748 , _f_permutation__n5747 ,
         _f_permutation__n5746 , _f_permutation__n5745 ,
         _f_permutation__n5744 , _f_permutation__n5743 ,
         _f_permutation__n5742 , _f_permutation__n5741 ,
         _f_permutation__n5740 , _f_permutation__n5739 ,
         _f_permutation__n5738 , _f_permutation__n5737 ,
         _f_permutation__n5736 , _f_permutation__n5735 ,
         _f_permutation__n5734 , _f_permutation__n5733 ,
         _f_permutation__n5732 , _f_permutation__n5731 ,
         _f_permutation__n5730 , _f_permutation__n5729 ,
         _f_permutation__n5728 , _f_permutation__n5727 ,
         _f_permutation__n5726 , _f_permutation__n5725 ,
         _f_permutation__n5724 , _f_permutation__n5723 ,
         _f_permutation__n5722 , _f_permutation__n5721 ,
         _f_permutation__n5720 , _f_permutation__n5719 ,
         _f_permutation__n5718 , _f_permutation__n5717 ,
         _f_permutation__n5716 , _f_permutation__n5715 ,
         _f_permutation__n5714 , _f_permutation__n5713 ,
         _f_permutation__n5712 , _f_permutation__n5711 ,
         _f_permutation__n5710 , _f_permutation__n5709 ,
         _f_permutation__n5708 , _f_permutation__n5707 ,
         _f_permutation__n5706 , _f_permutation__n5705 ,
         _f_permutation__n5704 , _f_permutation__n5703 ,
         _f_permutation__n5702 , _f_permutation__n5701 ,
         _f_permutation__n5700 , _f_permutation__n5699 ,
         _f_permutation__n5698 , _f_permutation__n5697 ,
         _f_permutation__n5696 , _f_permutation__n5695 ,
         _f_permutation__n5694 , _f_permutation__n5693 ,
         _f_permutation__n5692 , _f_permutation__n5691 ,
         _f_permutation__n5690 , _f_permutation__n5689 ,
         _f_permutation__n5688 , _f_permutation__n5687 ,
         _f_permutation__n5686 , _f_permutation__n5685 ,
         _f_permutation__n5684 , _f_permutation__n5683 ,
         _f_permutation__n5682 , _f_permutation__n5681 ,
         _f_permutation__n5680 , _f_permutation__n5679 ,
         _f_permutation__n5678 , _f_permutation__n5677 ,
         _f_permutation__n5676 , _f_permutation__n5675 ,
         _f_permutation__n5674 , _f_permutation__n5673 ,
         _f_permutation__n5672 , _f_permutation__n5671 ,
         _f_permutation__n5670 , _f_permutation__n5669 ,
         _f_permutation__n5668 , _f_permutation__n5667 ,
         _f_permutation__n5666 , _f_permutation__n5665 ,
         _f_permutation__n5664 , _f_permutation__n5663 ,
         _f_permutation__n5662 , _f_permutation__n5661 ,
         _f_permutation__n5660 , _f_permutation__n5659 ,
         _f_permutation__n5658 , _f_permutation__n5657 ,
         _f_permutation__n5656 , _f_permutation__n5655 ,
         _f_permutation__n5654 , _f_permutation__n5653 ,
         _f_permutation__n5652 , _f_permutation__n5651 ,
         _f_permutation__n5650 , _f_permutation__n5649 ,
         _f_permutation__n5648 , _f_permutation__n5647 ,
         _f_permutation__n5646 , _f_permutation__n5645 ,
         _f_permutation__n5644 , _f_permutation__n5643 ,
         _f_permutation__n5642 , _f_permutation__n5641 ,
         _f_permutation__n5640 , _f_permutation__n5639 ,
         _f_permutation__n5638 , _f_permutation__n5637 ,
         _f_permutation__n5636 , _f_permutation__n5635 ,
         _f_permutation__n5634 , _f_permutation__n5633 ,
         _f_permutation__n5632 , _f_permutation__n5631 ,
         _f_permutation__n5630 , _f_permutation__n5629 ,
         _f_permutation__n5628 , _f_permutation__n5627 ,
         _f_permutation__n5626 , _f_permutation__n5625 ,
         _f_permutation__n5624 , _f_permutation__n5623 ,
         _f_permutation__n5622 , _f_permutation__n5621 ,
         _f_permutation__n5620 , _f_permutation__n5619 ,
         _f_permutation__n5618 , _f_permutation__n5617 ,
         _f_permutation__n5616 , _f_permutation__n5615 ,
         _f_permutation__n5614 , _f_permutation__n5613 ,
         _f_permutation__n5612 , _f_permutation__n5611 ,
         _f_permutation__n5610 , _f_permutation__n5609 ,
         _f_permutation__n5608 , _f_permutation__n5607 ,
         _f_permutation__n5606 , _f_permutation__n5605 ,
         _f_permutation__n5604 , _f_permutation__n5603 ,
         _f_permutation__n5602 , _f_permutation__n5601 ,
         _f_permutation__n5600 , _f_permutation__n5599 ,
         _f_permutation__n5598 , _f_permutation__n5597 ,
         _f_permutation__n5596 , _f_permutation__n5595 ,
         _f_permutation__n5594 , _f_permutation__n5593 ,
         _f_permutation__n5592 , _f_permutation__n5591 ,
         _f_permutation__n5590 , _f_permutation__n5589 ,
         _f_permutation__n5588 , _f_permutation__n5587 ,
         _f_permutation__n5586 , _f_permutation__n5585 ,
         _f_permutation__n5584 , _f_permutation__n5583 ,
         _f_permutation__n5582 , _f_permutation__n5581 ,
         _f_permutation__n5580 , _f_permutation__n5579 ,
         _f_permutation__n5578 , _f_permutation__n5577 ,
         _f_permutation__n5576 , _f_permutation__n5575 ,
         _f_permutation__n5574 , _f_permutation__n5573 ,
         _f_permutation__n5572 , _f_permutation__n5571 ,
         _f_permutation__n5570 , _f_permutation__n5569 ,
         _f_permutation__n5568 , _f_permutation__n5567 ,
         _f_permutation__n5566 , _f_permutation__n5565 ,
         _f_permutation__n5564 , _f_permutation__n5563 ,
         _f_permutation__n5562 , _f_permutation__n5561 ,
         _f_permutation__n5560 , _f_permutation__n5559 ,
         _f_permutation__n5558 , _f_permutation__n5557 ,
         _f_permutation__n5556 , _f_permutation__n5555 ,
         _f_permutation__n5554 , _f_permutation__n5553 ,
         _f_permutation__n5552 , _f_permutation__n5551 ,
         _f_permutation__n5550 , _f_permutation__n5549 ,
         _f_permutation__n5548 , _f_permutation__n5547 ,
         _f_permutation__n5546 , _f_permutation__n5545 ,
         _f_permutation__n5544 , _f_permutation__n5543 ,
         _f_permutation__n5542 , _f_permutation__n5541 ,
         _f_permutation__n5540 , _f_permutation__n5539 ,
         _f_permutation__n5538 , _f_permutation__n5537 ,
         _f_permutation__n5536 , _f_permutation__n5535 ,
         _f_permutation__n5534 , _f_permutation__n5533 ,
         _f_permutation__n5532 , _f_permutation__n5531 ,
         _f_permutation__n5530 , _f_permutation__n5529 ,
         _f_permutation__n5528 , _f_permutation__n5527 ,
         _f_permutation__n5526 , _f_permutation__n5525 ,
         _f_permutation__n5524 , _f_permutation__n5523 ,
         _f_permutation__n5522 , _f_permutation__n5521 ,
         _f_permutation__n5520 , _f_permutation__n5519 ,
         _f_permutation__n5518 , _f_permutation__n5517 ,
         _f_permutation__n5516 , _f_permutation__n5515 ,
         _f_permutation__n5514 , _f_permutation__n5513 ,
         _f_permutation__n5512 , _f_permutation__n5511 ,
         _f_permutation__n5510 , _f_permutation__n5509 ,
         _f_permutation__n5508 , _f_permutation__n5507 ,
         _f_permutation__n5506 , _f_permutation__n5505 ,
         _f_permutation__n5504 , _f_permutation__n5503 ,
         _f_permutation__n5502 , _f_permutation__n5501 ,
         _f_permutation__n5500 , _f_permutation__n5499 ,
         _f_permutation__n5498 , _f_permutation__n5497 ,
         _f_permutation__n5496 , _f_permutation__n5495 ,
         _f_permutation__n5494 , _f_permutation__n5493 ,
         _f_permutation__n5492 , _f_permutation__n5491 ,
         _f_permutation__n5490 , _f_permutation__n5489 ,
         _f_permutation__n5488 , _f_permutation__n5487 ,
         _f_permutation__n5486 , _f_permutation__n5485 ,
         _f_permutation__n5484 , _f_permutation__n5483 ,
         _f_permutation__n5482 , _f_permutation__n5481 ,
         _f_permutation__n5480 , _f_permutation__n5479 ,
         _f_permutation__n5478 , _f_permutation__n5477 ,
         _f_permutation__n5476 , _f_permutation__n5475 ,
         _f_permutation__n5474 , _f_permutation__n5473 ,
         _f_permutation__n5472 , _f_permutation__n5471 ,
         _f_permutation__n5470 , _f_permutation__n5469 ,
         _f_permutation__n5468 , _f_permutation__n5467 ,
         _f_permutation__n5466 , _f_permutation__n5465 ,
         _f_permutation__n5464 , _f_permutation__n5463 ,
         _f_permutation__n5462 , _f_permutation__n5461 ,
         _f_permutation__n5460 , _f_permutation__n5459 ,
         _f_permutation__n5458 , _f_permutation__n5457 ,
         _f_permutation__n5456 , _f_permutation__n5455 ,
         _f_permutation__n5454 , _f_permutation__n5453 ,
         _f_permutation__n5452 , _f_permutation__n5451 ,
         _f_permutation__n5450 , _f_permutation__n5449 ,
         _f_permutation__n5448 , _f_permutation__n5447 ,
         _f_permutation__n5446 , _f_permutation__n5445 ,
         _f_permutation__n5444 , _f_permutation__n5443 ,
         _f_permutation__n5442 , _f_permutation__n5441 ,
         _f_permutation__n5440 , _f_permutation__n5439 ,
         _f_permutation__n5438 , _f_permutation__n5437 ,
         _f_permutation__n5436 , _f_permutation__n5435 ,
         _f_permutation__n5434 , _f_permutation__n5433 ,
         _f_permutation__n5432 , _f_permutation__n5431 ,
         _f_permutation__n5430 , _f_permutation__n5429 ,
         _f_permutation__n5428 , _f_permutation__n5427 ,
         _f_permutation__n5426 , _f_permutation__n5425 ,
         _f_permutation__n5424 , _f_permutation__n5423 ,
         _f_permutation__n5422 , _f_permutation__n5421 ,
         _f_permutation__n5420 , _f_permutation__n5419 ,
         _f_permutation__n5418 , _f_permutation__n5417 ,
         _f_permutation__n5416 , _f_permutation__n5415 ,
         _f_permutation__n5414 , _f_permutation__n5413 ,
         _f_permutation__n5412 , _f_permutation__n5411 ,
         _f_permutation__n5410 , _f_permutation__n5409 ,
         _f_permutation__n5408 , _f_permutation__n5407 ,
         _f_permutation__n5406 , _f_permutation__n5405 ,
         _f_permutation__n5404 , _f_permutation__n5403 ,
         _f_permutation__n5402 , _f_permutation__n5401 ,
         _f_permutation__n5400 , _f_permutation__n5399 ,
         _f_permutation__n5398 , _f_permutation__n5397 ,
         _f_permutation__n5396 , _f_permutation__n5395 ,
         _f_permutation__n5394 , _f_permutation__n5393 ,
         _f_permutation__n5392 , _f_permutation__n5391 ,
         _f_permutation__n5390 , _f_permutation__n5389 ,
         _f_permutation__n3787 , _f_permutation__n3786 ,
         _f_permutation__n3785 , _f_permutation__n3784 ,
         _f_permutation__n3783 , _f_permutation__n3782 ,
         _f_permutation__n3781 , _f_permutation__n3780 ,
         _f_permutation__n3779 , _f_permutation__n3778 ,
         _f_permutation__n3777 , _f_permutation__n3776 ,
         _f_permutation__n3775 , _f_permutation__n3774 ,
         _f_permutation__n3773 , _f_permutation__n3772 ,
         _f_permutation__n3771 , _f_permutation__n3770 ,
         _f_permutation__n3769 , _f_permutation__n3768 ,
         _f_permutation__n3767 , _f_permutation__n3766 ,
         _f_permutation__n3765 , _f_permutation__n3764 ,
         _f_permutation__n3763 , _f_permutation__n3762 ,
         _f_permutation__n3761 , _f_permutation__n3760 ,
         _f_permutation__n3759 , _f_permutation__n3758 ,
         _f_permutation__n3757 , _f_permutation__n3756 ,
         _f_permutation__n3755 , _f_permutation__n3754 ,
         _f_permutation__n3753 , _f_permutation__n3752 ,
         _f_permutation__n3751 , _f_permutation__n3750 ,
         _f_permutation__n3749 , _f_permutation__n3748 ,
         _f_permutation__n3747 , _f_permutation__n3746 ,
         _f_permutation__n3745 , _f_permutation__n3744 ,
         _f_permutation__n3743 , _f_permutation__n3742 ,
         _f_permutation__n3741 , _f_permutation__n3740 ,
         _f_permutation__n3739 , _f_permutation__n3738 ,
         _f_permutation__n3737 , _f_permutation__n3736 ,
         _f_permutation__n3735 , _f_permutation__n3734 ,
         _f_permutation__n3733 , _f_permutation__n3732 ,
         _f_permutation__n3731 , _f_permutation__n3730 ,
         _f_permutation__n3729 , _f_permutation__n3728 ,
         _f_permutation__n3727 , _f_permutation__n3726 ,
         _f_permutation__n3725 , _f_permutation__n3724 ,
         _f_permutation__n3723 , _f_permutation__n3722 ,
         _f_permutation__n3721 , _f_permutation__n3720 ,
         _f_permutation__n3719 , _f_permutation__n3718 ,
         _f_permutation__n3717 , _f_permutation__n3716 ,
         _f_permutation__n3715 , _f_permutation__n3714 ,
         _f_permutation__n3713 , _f_permutation__n3712 ,
         _f_permutation__n3711 , _f_permutation__n3710 ,
         _f_permutation__n3709 , _f_permutation__n3708 ,
         _f_permutation__n3707 , _f_permutation__n3706 ,
         _f_permutation__n3705 , _f_permutation__n3704 ,
         _f_permutation__n3703 , _f_permutation__n3702 ,
         _f_permutation__n3701 , _f_permutation__n3700 ,
         _f_permutation__n3699 , _f_permutation__n3698 ,
         _f_permutation__n3697 , _f_permutation__n3696 ,
         _f_permutation__n3695 , _f_permutation__n3694 ,
         _f_permutation__n3693 , _f_permutation__n3692 ,
         _f_permutation__n3691 , _f_permutation__n3690 ,
         _f_permutation__n3689 , _f_permutation__n3688 ,
         _f_permutation__n3687 , _f_permutation__n3686 ,
         _f_permutation__n3685 , _f_permutation__n3684 ,
         _f_permutation__n3683 , _f_permutation__n3682 ,
         _f_permutation__n3681 , _f_permutation__n3680 ,
         _f_permutation__n3679 , _f_permutation__n3678 ,
         _f_permutation__n3677 , _f_permutation__n3676 ,
         _f_permutation__n3675 , _f_permutation__n3674 ,
         _f_permutation__n3673 , _f_permutation__n3672 ,
         _f_permutation__n3671 , _f_permutation__n3670 ,
         _f_permutation__n3669 , _f_permutation__n3668 ,
         _f_permutation__n3667 , _f_permutation__n3666 ,
         _f_permutation__n3665 , _f_permutation__n3664 ,
         _f_permutation__n3663 , _f_permutation__n3662 ,
         _f_permutation__n3661 , _f_permutation__n3660 ,
         _f_permutation__n3659 , _f_permutation__n3658 ,
         _f_permutation__n3657 , _f_permutation__n3656 ,
         _f_permutation__n3655 , _f_permutation__n3654 ,
         _f_permutation__n3653 , _f_permutation__n3652 ,
         _f_permutation__n3651 , _f_permutation__n3650 ,
         _f_permutation__n3649 , _f_permutation__n3648 ,
         _f_permutation__n3647 , _f_permutation__n3646 ,
         _f_permutation__n3645 , _f_permutation__n3644 ,
         _f_permutation__n3643 , _f_permutation__n3642 ,
         _f_permutation__n3641 , _f_permutation__n3640 ,
         _f_permutation__n3639 , _f_permutation__n3638 ,
         _f_permutation__n3637 , _f_permutation__n3636 ,
         _f_permutation__n3635 , _f_permutation__n3634 ,
         _f_permutation__n3633 , _f_permutation__n3632 ,
         _f_permutation__n3631 , _f_permutation__n3630 ,
         _f_permutation__n3629 , _f_permutation__n3628 ,
         _f_permutation__n3627 , _f_permutation__n3626 ,
         _f_permutation__n3625 , _f_permutation__n3624 ,
         _f_permutation__n3623 , _f_permutation__n3622 ,
         _f_permutation__n3621 , _f_permutation__n3620 ,
         _f_permutation__n3619 , _f_permutation__n3618 ,
         _f_permutation__n3617 , _f_permutation__n3616 ,
         _f_permutation__n3615 , _f_permutation__n3614 ,
         _f_permutation__n3613 , _f_permutation__n3612 ,
         _f_permutation__n3611 , _f_permutation__n3610 ,
         _f_permutation__n3609 , _f_permutation__n3608 ,
         _f_permutation__n3607 , _f_permutation__n3606 ,
         _f_permutation__n3605 , _f_permutation__n3604 ,
         _f_permutation__n3603 , _f_permutation__n3602 ,
         _f_permutation__n3601 , _f_permutation__n3600 ,
         _f_permutation__n3599 , _f_permutation__n3598 ,
         _f_permutation__n3597 , _f_permutation__n3596 ,
         _f_permutation__n3595 , _f_permutation__n3594 ,
         _f_permutation__n3593 , _f_permutation__n3592 ,
         _f_permutation__n3591 , _f_permutation__n3590 ,
         _f_permutation__n3589 , _f_permutation__n3588 ,
         _f_permutation__n3587 , _f_permutation__n3586 ,
         _f_permutation__n3585 , _f_permutation__n3584 ,
         _f_permutation__n3583 , _f_permutation__n3582 ,
         _f_permutation__n3581 , _f_permutation__n3580 ,
         _f_permutation__n3579 , _f_permutation__n3578 ,
         _f_permutation__n3577 , _f_permutation__n3576 ,
         _f_permutation__n3575 , _f_permutation__n3574 ,
         _f_permutation__n3573 , _f_permutation__n3572 ,
         _f_permutation__n3571 , _f_permutation__n3570 ,
         _f_permutation__n3569 , _f_permutation__n3568 ,
         _f_permutation__n3567 , _f_permutation__n3566 ,
         _f_permutation__n3565 , _f_permutation__n3564 ,
         _f_permutation__n3563 , _f_permutation__n3562 ,
         _f_permutation__n3561 , _f_permutation__n3560 ,
         _f_permutation__n3559 , _f_permutation__n3558 ,
         _f_permutation__n3557 , _f_permutation__n3556 ,
         _f_permutation__n3555 , _f_permutation__n3554 ,
         _f_permutation__n3553 , _f_permutation__n3552 ,
         _f_permutation__n3551 , _f_permutation__n3550 ,
         _f_permutation__n3549 , _f_permutation__n3548 ,
         _f_permutation__n3547 , _f_permutation__n3546 ,
         _f_permutation__n3545 , _f_permutation__n3544 ,
         _f_permutation__n3543 , _f_permutation__n3542 ,
         _f_permutation__n3541 , _f_permutation__n3540 ,
         _f_permutation__n3539 , _f_permutation__n3538 ,
         _f_permutation__n3537 , _f_permutation__n3536 ,
         _f_permutation__n3535 , _f_permutation__n3534 ,
         _f_permutation__n3533 , _f_permutation__n3532 ,
         _f_permutation__n3531 , _f_permutation__n3530 ,
         _f_permutation__n3529 , _f_permutation__n3528 ,
         _f_permutation__n3527 , _f_permutation__n3526 ,
         _f_permutation__n3525 , _f_permutation__n3524 ,
         _f_permutation__n3523 , _f_permutation__n3522 ,
         _f_permutation__n3521 , _f_permutation__n3520 ,
         _f_permutation__n3519 , _f_permutation__n3518 ,
         _f_permutation__n3517 , _f_permutation__n3516 ,
         _f_permutation__n3515 , _f_permutation__n3514 ,
         _f_permutation__n3513 , _f_permutation__n3512 ,
         _f_permutation__n3511 , _f_permutation__n3510 ,
         _f_permutation__n3509 , _f_permutation__n3508 ,
         _f_permutation__n3507 , _f_permutation__n3506 ,
         _f_permutation__n3505 , _f_permutation__n3504 ,
         _f_permutation__n3503 , _f_permutation__n3502 ,
         _f_permutation__n3501 , _f_permutation__n3500 ,
         _f_permutation__n3499 , _f_permutation__n3498 ,
         _f_permutation__n3497 , _f_permutation__n3496 ,
         _f_permutation__n3495 , _f_permutation__n3494 ,
         _f_permutation__n3493 , _f_permutation__n3492 ,
         _f_permutation__n3491 , _f_permutation__n3490 ,
         _f_permutation__n3489 , _f_permutation__n3488 ,
         _f_permutation__n3487 , _f_permutation__n3486 ,
         _f_permutation__n3485 , _f_permutation__n3484 ,
         _f_permutation__n3483 , _f_permutation__n3482 ,
         _f_permutation__n3481 , _f_permutation__n3480 ,
         _f_permutation__n3479 , _f_permutation__n3478 ,
         _f_permutation__n3477 , _f_permutation__n3476 ,
         _f_permutation__n3475 , _f_permutation__n3474 ,
         _f_permutation__n3473 , _f_permutation__n3472 ,
         _f_permutation__n3471 , _f_permutation__n3470 ,
         _f_permutation__n3469 , _f_permutation__n3468 ,
         _f_permutation__n3467 , _f_permutation__n3466 ,
         _f_permutation__n3465 , _f_permutation__n3464 ,
         _f_permutation__n3463 , _f_permutation__n3462 ,
         _f_permutation__n3461 , _f_permutation__n3460 ,
         _f_permutation__n3459 , _f_permutation__n3458 ,
         _f_permutation__n3457 , _f_permutation__n3456 ,
         _f_permutation__n3455 , _f_permutation__n3454 ,
         _f_permutation__n3453 , _f_permutation__n3452 ,
         _f_permutation__n3451 , _f_permutation__n3450 ,
         _f_permutation__n3449 , _f_permutation__n3448 ,
         _f_permutation__n3447 , _f_permutation__n3446 ,
         _f_permutation__n3445 , _f_permutation__n3444 ,
         _f_permutation__n3443 , _f_permutation__n3442 ,
         _f_permutation__n3441 , _f_permutation__n3440 ,
         _f_permutation__n3439 , _f_permutation__n3438 ,
         _f_permutation__n3437 , _f_permutation__n3436 ,
         _f_permutation__n3435 , _f_permutation__n3434 ,
         _f_permutation__n3433 , _f_permutation__n3432 ,
         _f_permutation__n3431 , _f_permutation__n3430 ,
         _f_permutation__n3429 , _f_permutation__n3428 ,
         _f_permutation__n3427 , _f_permutation__n3426 ,
         _f_permutation__n3425 , _f_permutation__n3424 ,
         _f_permutation__n3423 , _f_permutation__n3422 ,
         _f_permutation__n3421 , _f_permutation__n3420 ,
         _f_permutation__n3419 , _f_permutation__n3418 ,
         _f_permutation__n3417 , _f_permutation__n3416 ,
         _f_permutation__n3415 , _f_permutation__n3414 ,
         _f_permutation__n3413 , _f_permutation__n3412 ,
         _f_permutation__n3411 , _f_permutation__n3410 ,
         _f_permutation__n3409 , _f_permutation__n3408 ,
         _f_permutation__n3407 , _f_permutation__n3406 ,
         _f_permutation__n3405 , _f_permutation__n3404 ,
         _f_permutation__n3403 , _f_permutation__n3402 ,
         _f_permutation__n3401 , _f_permutation__n3400 ,
         _f_permutation__n3399 , _f_permutation__n3398 ,
         _f_permutation__n3397 , _f_permutation__n3396 ,
         _f_permutation__n3395 , _f_permutation__n3394 ,
         _f_permutation__n3393 , _f_permutation__n3392 ,
         _f_permutation__n3391 , _f_permutation__n3390 ,
         _f_permutation__n3389 , _f_permutation__n3388 ,
         _f_permutation__n3387 , _f_permutation__n3386 ,
         _f_permutation__n3385 , _f_permutation__n3384 ,
         _f_permutation__n3383 , _f_permutation__n3382 ,
         _f_permutation__n3381 , _f_permutation__n3380 ,
         _f_permutation__n3379 , _f_permutation__n3378 ,
         _f_permutation__n3377 , _f_permutation__n3376 ,
         _f_permutation__n3375 , _f_permutation__n3374 ,
         _f_permutation__n3373 , _f_permutation__n3372 ,
         _f_permutation__n3371 , _f_permutation__n3370 ,
         _f_permutation__n3369 , _f_permutation__n3368 ,
         _f_permutation__n3367 , _f_permutation__n3366 ,
         _f_permutation__n3365 , _f_permutation__n3364 ,
         _f_permutation__n3363 , _f_permutation__n3362 ,
         _f_permutation__n3361 , _f_permutation__n3360 ,
         _f_permutation__n3359 , _f_permutation__n3358 ,
         _f_permutation__n3357 , _f_permutation__n3356 ,
         _f_permutation__n3355 , _f_permutation__n3354 ,
         _f_permutation__n3353 , _f_permutation__n3352 ,
         _f_permutation__n3351 , _f_permutation__n3350 ,
         _f_permutation__n3349 , _f_permutation__n3348 ,
         _f_permutation__n3347 , _f_permutation__n3346 ,
         _f_permutation__n3345 , _f_permutation__n3344 ,
         _f_permutation__n3343 , _f_permutation__n3342 ,
         _f_permutation__n3341 , _f_permutation__n3340 ,
         _f_permutation__n3339 , _f_permutation__n3338 ,
         _f_permutation__n3337 , _f_permutation__n3336 ,
         _f_permutation__n3335 , _f_permutation__n3334 ,
         _f_permutation__n3333 , _f_permutation__n3332 ,
         _f_permutation__n3331 , _f_permutation__n3330 ,
         _f_permutation__n3329 , _f_permutation__n3328 ,
         _f_permutation__n3327 , _f_permutation__n3326 ,
         _f_permutation__n3325 , _f_permutation__n3324 ,
         _f_permutation__n3323 , _f_permutation__n3322 ,
         _f_permutation__n3321 , _f_permutation__n3320 ,
         _f_permutation__n3319 , _f_permutation__n3318 ,
         _f_permutation__n3317 , _f_permutation__n3316 ,
         _f_permutation__n3315 , _f_permutation__n3314 ,
         _f_permutation__n3313 , _f_permutation__n3312 ,
         _f_permutation__n3311 , _f_permutation__n3310 ,
         _f_permutation__n3309 , _f_permutation__n3308 ,
         _f_permutation__n3307 , _f_permutation__n3306 ,
         _f_permutation__n3305 , _f_permutation__n3304 ,
         _f_permutation__n3303 , _f_permutation__n3302 ,
         _f_permutation__n3301 , _f_permutation__n3300 ,
         _f_permutation__n3299 , _f_permutation__n3298 ,
         _f_permutation__n3297 , _f_permutation__n3296 ,
         _f_permutation__n3295 , _f_permutation__n3294 ,
         _f_permutation__n3293 , _f_permutation__n3292 ,
         _f_permutation__n3291 , _f_permutation__n3290 ,
         _f_permutation__n3289 , _f_permutation__n3288 ,
         _f_permutation__n3287 , _f_permutation__n3286 ,
         _f_permutation__n3285 , _f_permutation__n3284 ,
         _f_permutation__n3283 , _f_permutation__n3282 ,
         _f_permutation__n3281 , _f_permutation__n3280 ,
         _f_permutation__n3279 , _f_permutation__n3278 ,
         _f_permutation__n3277 , _f_permutation__n3276 ,
         _f_permutation__n3275 , _f_permutation__n3274 ,
         _f_permutation__n3273 , _f_permutation__n3272 ,
         _f_permutation__n3271 , _f_permutation__n3270 ,
         _f_permutation__n3269 , _f_permutation__n3268 ,
         _f_permutation__n3267 , _f_permutation__n3266 ,
         _f_permutation__n3265 , _f_permutation__n3264 ,
         _f_permutation__n3263 , _f_permutation__n3262 ,
         _f_permutation__n3261 , _f_permutation__n3260 ,
         _f_permutation__n3259 , _f_permutation__n3258 ,
         _f_permutation__n3257 , _f_permutation__n3256 ,
         _f_permutation__n3255 , _f_permutation__n3254 ,
         _f_permutation__n3253 , _f_permutation__n3252 ,
         _f_permutation__n3251 , _f_permutation__n3250 ,
         _f_permutation__n3249 , _f_permutation__n3248 ,
         _f_permutation__n3247 , _f_permutation__n3246 ,
         _f_permutation__n3245 , _f_permutation__n3244 ,
         _f_permutation__n3243 , _f_permutation__n3242 ,
         _f_permutation__n3241 , _f_permutation__n3240 ,
         _f_permutation__n3239 , _f_permutation__n3238 ,
         _f_permutation__n3237 , _f_permutation__n3236 ,
         _f_permutation__n3235 , _f_permutation__n3234 ,
         _f_permutation__n3233 , _f_permutation__n3232 ,
         _f_permutation__n3231 , _f_permutation__n3230 ,
         _f_permutation__n3229 , _f_permutation__n3228 ,
         _f_permutation__n3227 , _f_permutation__n3226 ,
         _f_permutation__n3225 , _f_permutation__n3224 ,
         _f_permutation__n3223 , _f_permutation__n3222 ,
         _f_permutation__n3221 , _f_permutation__n3220 ,
         _f_permutation__n3219 , _f_permutation__n3218 ,
         _f_permutation__n3217 , _f_permutation__n3216 ,
         _f_permutation__n3215 , _f_permutation__n3214 ,
         _f_permutation__n3213 , _f_permutation__n3212 ,
         _f_permutation__n3211 , _f_permutation__n3210 ,
         _f_permutation__n3209 , _f_permutation__n3208 ,
         _f_permutation__n3207 , _f_permutation__n3206 ,
         _f_permutation__n3205 , _f_permutation__n3204 ,
         _f_permutation__n3203 , _f_permutation__n3202 ,
         _f_permutation__n3201 , _f_permutation__n3200 ,
         _f_permutation__n3199 , _f_permutation__n3198 ,
         _f_permutation__n3197 , _f_permutation__n3196 ,
         _f_permutation__n3195 , _f_permutation__n3194 ,
         _f_permutation__n3193 , _f_permutation__n3192 ,
         _f_permutation__n3191 , _f_permutation__n3190 ,
         _f_permutation__n3189 , _f_permutation__n3188 ,
         _f_permutation__n3187 , _f_permutation__n3186 ,
         _f_permutation__n3185 , _f_permutation__n3184 ,
         _f_permutation__n3183 , _f_permutation__n3182 ,
         _f_permutation__n3181 , _f_permutation__n3180 ,
         _f_permutation__n3179 , _f_permutation__n3178 ,
         _f_permutation__n3177 , _f_permutation__n3176 ,
         _f_permutation__n3175 , _f_permutation__n3174 ,
         _f_permutation__n3173 , _f_permutation__n3172 ,
         _f_permutation__n3171 , _f_permutation__n3170 ,
         _f_permutation__n3169 , _f_permutation__n3168 ,
         _f_permutation__n3167 , _f_permutation__n3166 ,
         _f_permutation__n3165 , _f_permutation__n3164 ,
         _f_permutation__n3163 , _f_permutation__n3162 ,
         _f_permutation__n3161 , _f_permutation__n3160 ,
         _f_permutation__n3159 , _f_permutation__n3158 ,
         _f_permutation__n3157 , _f_permutation__n3156 ,
         _f_permutation__n3155 , _f_permutation__n3154 ,
         _f_permutation__n3153 , _f_permutation__n3152 ,
         _f_permutation__n3151 , _f_permutation__n3150 ,
         _f_permutation__n3149 , _f_permutation__n3148 ,
         _f_permutation__n3147 , _f_permutation__n3146 ,
         _f_permutation__n3145 , _f_permutation__n3144 ,
         _f_permutation__n3143 , _f_permutation__n3142 ,
         _f_permutation__n3141 , _f_permutation__n3140 ,
         _f_permutation__n3139 , _f_permutation__n3138 ,
         _f_permutation__n3137 , _f_permutation__n3136 ,
         _f_permutation__n3135 , _f_permutation__n3134 ,
         _f_permutation__n3133 , _f_permutation__n3132 ,
         _f_permutation__n3131 , _f_permutation__n3130 ,
         _f_permutation__n3129 , _f_permutation__n3128 ,
         _f_permutation__n3127 , _f_permutation__n3126 ,
         _f_permutation__n3125 , _f_permutation__n3124 ,
         _f_permutation__n3123 , _f_permutation__n3122 ,
         _f_permutation__n3121 , _f_permutation__n3120 ,
         _f_permutation__n3119 , _f_permutation__n3118 ,
         _f_permutation__n3117 , _f_permutation__n3116 ,
         _f_permutation__n3115 , _f_permutation__n3114 ,
         _f_permutation__n3113 , _f_permutation__n3112 ,
         _f_permutation__n3111 , _f_permutation__n3110 ,
         _f_permutation__n3109 , _f_permutation__n3108 ,
         _f_permutation__n3107 , _f_permutation__n3106 ,
         _f_permutation__n3105 , _f_permutation__n3104 ,
         _f_permutation__n3103 , _f_permutation__n3102 ,
         _f_permutation__n3101 , _f_permutation__n3100 ,
         _f_permutation__n3099 , _f_permutation__n3098 ,
         _f_permutation__n3097 , _f_permutation__n3096 ,
         _f_permutation__n3095 , _f_permutation__n3094 ,
         _f_permutation__n3093 , _f_permutation__n3092 ,
         _f_permutation__n3091 , _f_permutation__n3090 ,
         _f_permutation__n3089 , _f_permutation__n3088 ,
         _f_permutation__n3087 , _f_permutation__n3086 ,
         _f_permutation__n3085 , _f_permutation__n3084 ,
         _f_permutation__n3083 , _f_permutation__n3082 ,
         _f_permutation__n3081 , _f_permutation__n3080 ,
         _f_permutation__n3079 , _f_permutation__n3078 ,
         _f_permutation__n3077 , _f_permutation__n3076 ,
         _f_permutation__n3075 , _f_permutation__n3074 ,
         _f_permutation__n3073 , _f_permutation__n3072 ,
         _f_permutation__n3071 , _f_permutation__n3070 ,
         _f_permutation__n3069 , _f_permutation__n3068 ,
         _f_permutation__n3067 , _f_permutation__n3066 ,
         _f_permutation__n3065 , _f_permutation__n3064 ,
         _f_permutation__n3063 , _f_permutation__n3062 ,
         _f_permutation__n3061 , _f_permutation__n3060 ,
         _f_permutation__n3059 , _f_permutation__n3058 ,
         _f_permutation__n3057 , _f_permutation__n3056 ,
         _f_permutation__n3055 , _f_permutation__n3054 ,
         _f_permutation__n3053 , _f_permutation__n3052 ,
         _f_permutation__n3051 , _f_permutation__n3050 ,
         _f_permutation__n3049 , _f_permutation__n3048 ,
         _f_permutation__n3047 , _f_permutation__n3046 ,
         _f_permutation__n3045 , _f_permutation__n3044 ,
         _f_permutation__n3043 , _f_permutation__n3042 ,
         _f_permutation__n3041 , _f_permutation__n3040 ,
         _f_permutation__n3039 , _f_permutation__n3038 ,
         _f_permutation__n3037 , _f_permutation__n3036 ,
         _f_permutation__n3035 , _f_permutation__n3034 ,
         _f_permutation__n3033 , _f_permutation__n3032 ,
         _f_permutation__n3031 , _f_permutation__n3030 ,
         _f_permutation__n3029 , _f_permutation__n3028 ,
         _f_permutation__n3027 , _f_permutation__n3026 ,
         _f_permutation__n3025 , _f_permutation__n3024 ,
         _f_permutation__n3023 , _f_permutation__n3022 ,
         _f_permutation__n3021 , _f_permutation__n3020 ,
         _f_permutation__n3019 , _f_permutation__n3018 ,
         _f_permutation__n3017 , _f_permutation__n3016 ,
         _f_permutation__n3015 , _f_permutation__n3014 ,
         _f_permutation__n3013 , _f_permutation__n3012 ,
         _f_permutation__n3011 , _f_permutation__n3010 ,
         _f_permutation__n3009 , _f_permutation__n3008 ,
         _f_permutation__n3007 , _f_permutation__n3006 ,
         _f_permutation__n3005 , _f_permutation__n3004 ,
         _f_permutation__n3003 , _f_permutation__n3002 ,
         _f_permutation__n3001 , _f_permutation__n3000 ,
         _f_permutation__n2999 , _f_permutation__n2998 ,
         _f_permutation__n2997 , _f_permutation__n2996 ,
         _f_permutation__n2995 , _f_permutation__n2994 ,
         _f_permutation__n2993 , _f_permutation__n2992 ,
         _f_permutation__n2991 , _f_permutation__n2990 ,
         _f_permutation__n2989 , _f_permutation__n2988 ,
         _f_permutation__n2987 , _f_permutation__n2986 ,
         _f_permutation__n2985 , _f_permutation__n2984 ,
         _f_permutation__n2983 , _f_permutation__n2982 ,
         _f_permutation__n2981 , _f_permutation__n2980 ,
         _f_permutation__n2979 , _f_permutation__n2978 ,
         _f_permutation__n2977 , _f_permutation__n2976 ,
         _f_permutation__n2975 , _f_permutation__n2974 ,
         _f_permutation__n2973 , _f_permutation__n2972 ,
         _f_permutation__n2971 , _f_permutation__n2970 ,
         _f_permutation__n2969 , _f_permutation__n2968 ,
         _f_permutation__n2967 , _f_permutation__n2966 ,
         _f_permutation__n2965 , _f_permutation__n2964 ,
         _f_permutation__n2963 , _f_permutation__n2962 ,
         _f_permutation__n2961 , _f_permutation__n2960 ,
         _f_permutation__n2959 , _f_permutation__n2958 ,
         _f_permutation__n2957 , _f_permutation__n2956 ,
         _f_permutation__n2955 , _f_permutation__n2954 ,
         _f_permutation__n2953 , _f_permutation__n2952 ,
         _f_permutation__n2951 , _f_permutation__n2950 ,
         _f_permutation__n2949 , _f_permutation__n2948 ,
         _f_permutation__n2947 , _f_permutation__n2946 ,
         _f_permutation__n2945 , _f_permutation__n2944 ,
         _f_permutation__n2943 , _f_permutation__n2942 ,
         _f_permutation__n2941 , _f_permutation__n2940 ,
         _f_permutation__n2939 , _f_permutation__n2938 ,
         _f_permutation__n2937 , _f_permutation__n2936 ,
         _f_permutation__n2935 , _f_permutation__n2934 ,
         _f_permutation__n2933 , _f_permutation__n2932 ,
         _f_permutation__n2931 , _f_permutation__n2930 ,
         _f_permutation__n2929 , _f_permutation__n2928 ,
         _f_permutation__n2927 , _f_permutation__n2926 ,
         _f_permutation__n2925 , _f_permutation__n2924 ,
         _f_permutation__n2923 , _f_permutation__n2922 ,
         _f_permutation__n2921 , _f_permutation__n2920 ,
         _f_permutation__n2919 , _f_permutation__n2918 ,
         _f_permutation__n2917 , _f_permutation__n2916 ,
         _f_permutation__n2915 , _f_permutation__n2914 ,
         _f_permutation__n2913 , _f_permutation__n2912 ,
         _f_permutation__n2911 , _f_permutation__n2910 ,
         _f_permutation__n2909 , _f_permutation__n2908 ,
         _f_permutation__n2907 , _f_permutation__n2906 ,
         _f_permutation__n2905 , _f_permutation__n2904 ,
         _f_permutation__n2903 , _f_permutation__n2902 ,
         _f_permutation__n2901 , _f_permutation__n2900 ,
         _f_permutation__n2899 , _f_permutation__n2898 ,
         _f_permutation__n2897 , _f_permutation__n2896 ,
         _f_permutation__n2895 , _f_permutation__n2894 ,
         _f_permutation__n2893 , _f_permutation__n2892 ,
         _f_permutation__n2891 , _f_permutation__n2890 ,
         _f_permutation__n2889 , _f_permutation__n2888 ,
         _f_permutation__n2887 , _f_permutation__n2886 ,
         _f_permutation__n2885 , _f_permutation__n2884 ,
         _f_permutation__n2883 , _f_permutation__n2882 ,
         _f_permutation__n2881 , _f_permutation__n2880 ,
         _f_permutation__n2879 , _f_permutation__n2878 ,
         _f_permutation__n2877 , _f_permutation__n2876 ,
         _f_permutation__n2875 , _f_permutation__n2874 ,
         _f_permutation__n2873 , _f_permutation__n2872 ,
         _f_permutation__n2871 , _f_permutation__n2870 ,
         _f_permutation__n2869 , _f_permutation__n2868 ,
         _f_permutation__n2867 , _f_permutation__n2866 ,
         _f_permutation__n2865 , _f_permutation__n2864 ,
         _f_permutation__n2863 , _f_permutation__n2862 ,
         _f_permutation__n2861 , _f_permutation__n2860 ,
         _f_permutation__n2859 , _f_permutation__n2858 ,
         _f_permutation__n2857 , _f_permutation__n2856 ,
         _f_permutation__n2855 , _f_permutation__n2854 ,
         _f_permutation__n2853 , _f_permutation__n2852 ,
         _f_permutation__n2851 , _f_permutation__n2850 ,
         _f_permutation__n2849 , _f_permutation__n2848 ,
         _f_permutation__n2847 , _f_permutation__n2846 ,
         _f_permutation__n2845 , _f_permutation__n2844 ,
         _f_permutation__n2843 , _f_permutation__n2842 ,
         _f_permutation__n2841 , _f_permutation__n2840 ,
         _f_permutation__n2839 , _f_permutation__n2838 ,
         _f_permutation__n2837 , _f_permutation__n2836 ,
         _f_permutation__n2835 , _f_permutation__n2834 ,
         _f_permutation__n2833 , _f_permutation__n2832 ,
         _f_permutation__n2831 , _f_permutation__n2830 ,
         _f_permutation__n2829 , _f_permutation__n2828 ,
         _f_permutation__n2827 , _f_permutation__n2826 ,
         _f_permutation__n2825 , _f_permutation__n2824 ,
         _f_permutation__n2823 , _f_permutation__n2822 ,
         _f_permutation__n2821 , _f_permutation__n2820 ,
         _f_permutation__n2819 , _f_permutation__n2818 ,
         _f_permutation__n2817 , _f_permutation__n2816 ,
         _f_permutation__n2815 , _f_permutation__n2814 ,
         _f_permutation__n2813 , _f_permutation__n2812 ,
         _f_permutation__n2811 , _f_permutation__n2810 ,
         _f_permutation__n2809 , _f_permutation__n2808 ,
         _f_permutation__n2807 , _f_permutation__n2806 ,
         _f_permutation__n2805 , _f_permutation__n2804 ,
         _f_permutation__n2803 , _f_permutation__n2802 ,
         _f_permutation__n2801 , _f_permutation__n2800 ,
         _f_permutation__n2799 , _f_permutation__n2798 ,
         _f_permutation__n2797 , _f_permutation__n2796 ,
         _f_permutation__n2795 , _f_permutation__n2794 ,
         _f_permutation__n2793 , _f_permutation__n2792 ,
         _f_permutation__n2791 , _f_permutation__n2790 ,
         _f_permutation__n2789 , _f_permutation__n2788 ,
         _f_permutation__n2787 , _f_permutation__n2786 ,
         _f_permutation__n2785 , _f_permutation__n2784 ,
         _f_permutation__n2783 , _f_permutation__n2782 ,
         _f_permutation__n2781 , _f_permutation__n2780 ,
         _f_permutation__n2779 , _f_permutation__n2778 ,
         _f_permutation__n2777 , _f_permutation__n2776 ,
         _f_permutation__n2775 , _f_permutation__n2774 ,
         _f_permutation__n2773 , _f_permutation__n2772 ,
         _f_permutation__n2771 , _f_permutation__n2770 ,
         _f_permutation__n2769 , _f_permutation__n2768 ,
         _f_permutation__n2767 , _f_permutation__n2766 ,
         _f_permutation__n2765 , _f_permutation__n2764 ,
         _f_permutation__n2763 , _f_permutation__n2762 ,
         _f_permutation__n2761 , _f_permutation__n2760 ,
         _f_permutation__n2759 , _f_permutation__n2758 ,
         _f_permutation__n2757 , _f_permutation__n2756 ,
         _f_permutation__n2755 , _f_permutation__n2754 ,
         _f_permutation__n2753 , _f_permutation__n2752 ,
         _f_permutation__n2751 , _f_permutation__n2750 ,
         _f_permutation__n2749 , _f_permutation__n2748 ,
         _f_permutation__n2747 , _f_permutation__n2746 ,
         _f_permutation__n2745 , _f_permutation__n2744 ,
         _f_permutation__n2743 , _f_permutation__n2742 ,
         _f_permutation__n2741 , _f_permutation__n2740 ,
         _f_permutation__n2739 , _f_permutation__n2738 ,
         _f_permutation__n2737 , _f_permutation__n2736 ,
         _f_permutation__n2735 , _f_permutation__n2734 ,
         _f_permutation__n2733 , _f_permutation__n2732 ,
         _f_permutation__n2731 , _f_permutation__n2730 ,
         _f_permutation__n2729 , _f_permutation__n2728 ,
         _f_permutation__n2727 , _f_permutation__n2726 ,
         _f_permutation__n2725 , _f_permutation__n2724 ,
         _f_permutation__n2723 , _f_permutation__n2722 ,
         _f_permutation__n2721 , _f_permutation__n2720 ,
         _f_permutation__n2719 , _f_permutation__n2718 ,
         _f_permutation__n2717 , _f_permutation__n2716 ,
         _f_permutation__n2715 , _f_permutation__n2714 ,
         _f_permutation__n2713 , _f_permutation__n2712 ,
         _f_permutation__n2711 , _f_permutation__n2710 ,
         _f_permutation__n2709 , _f_permutation__n2708 ,
         _f_permutation__n2707 , _f_permutation__n2706 ,
         _f_permutation__n2705 , _f_permutation__n2704 ,
         _f_permutation__n2703 , _f_permutation__n2702 ,
         _f_permutation__n2701 , _f_permutation__n2700 ,
         _f_permutation__n2699 , _f_permutation__n2698 ,
         _f_permutation__n2697 , _f_permutation__n2696 ,
         _f_permutation__n2695 , _f_permutation__n2694 ,
         _f_permutation__n2693 , _f_permutation__n2692 ,
         _f_permutation__n2691 , _f_permutation__n2690 ,
         _f_permutation__n2689 , _f_permutation__n2688 ,
         _f_permutation__n2687 , _f_permutation__n2686 ,
         _f_permutation__n2685 , _f_permutation__n2684 ,
         _f_permutation__n2683 , _f_permutation__n2682 ,
         _f_permutation__n2681 , _f_permutation__n2680 ,
         _f_permutation__n2679 , _f_permutation__n2678 ,
         _f_permutation__n2677 , _f_permutation__n2676 ,
         _f_permutation__n2675 , _f_permutation__n2674 ,
         _f_permutation__n2673 , _f_permutation__n2672 ,
         _f_permutation__n2671 , _f_permutation__n2670 ,
         _f_permutation__n2669 , _f_permutation__n2668 ,
         _f_permutation__n2667 , _f_permutation__n2666 ,
         _f_permutation__n2665 , _f_permutation__n2664 ,
         _f_permutation__n2663 , _f_permutation__n2662 ,
         _f_permutation__n2661 , _f_permutation__n2660 ,
         _f_permutation__n2659 , _f_permutation__n2658 ,
         _f_permutation__n2657 , _f_permutation__n2656 ,
         _f_permutation__n2655 , _f_permutation__n2654 ,
         _f_permutation__n2653 , _f_permutation__n2652 ,
         _f_permutation__n2651 , _f_permutation__n2650 ,
         _f_permutation__n2649 , _f_permutation__n2648 ,
         _f_permutation__n2647 , _f_permutation__n2646 ,
         _f_permutation__n2645 , _f_permutation__n2644 ,
         _f_permutation__n2643 , _f_permutation__n2642 ,
         _f_permutation__n2641 , _f_permutation__n2640 ,
         _f_permutation__n2639 , _f_permutation__n2638 ,
         _f_permutation__n2637 , _f_permutation__n2636 ,
         _f_permutation__n2635 , _f_permutation__n2634 ,
         _f_permutation__n2633 , _f_permutation__n2632 ,
         _f_permutation__n2631 , _f_permutation__n2630 ,
         _f_permutation__n2629 , _f_permutation__n2628 ,
         _f_permutation__n2627 , _f_permutation__n2626 ,
         _f_permutation__n2625 , _f_permutation__n2624 ,
         _f_permutation__n2623 , _f_permutation__n2622 ,
         _f_permutation__n2621 , _f_permutation__n2620 ,
         _f_permutation__n2619 , _f_permutation__n2618 ,
         _f_permutation__n2617 , _f_permutation__n2616 ,
         _f_permutation__n2615 , _f_permutation__n2614 ,
         _f_permutation__n2613 , _f_permutation__n2612 ,
         _f_permutation__n2611 , _f_permutation__n2610 ,
         _f_permutation__n2609 , _f_permutation__n2608 ,
         _f_permutation__n2607 , _f_permutation__n2606 ,
         _f_permutation__n2605 , _f_permutation__n2604 ,
         _f_permutation__n2603 , _f_permutation__n2602 ,
         _f_permutation__n2601 , _f_permutation__n2600 ,
         _f_permutation__n2599 , _f_permutation__n2598 ,
         _f_permutation__n2597 , _f_permutation__n2596 ,
         _f_permutation__n2595 , _f_permutation__n2594 ,
         _f_permutation__n2593 , _f_permutation__n2592 ,
         _f_permutation__n2591 , _f_permutation__n2590 ,
         _f_permutation__n2589 , _f_permutation__n2588 ,
         _f_permutation__n2587 , _f_permutation__n2586 ,
         _f_permutation__n2585 , _f_permutation__n2584 ,
         _f_permutation__n2583 , _f_permutation__n2582 ,
         _f_permutation__n2581 , _f_permutation__n2580 ,
         _f_permutation__n2579 , _f_permutation__n2578 ,
         _f_permutation__n2577 , _f_permutation__n2576 ,
         _f_permutation__n2575 , _f_permutation__n2574 ,
         _f_permutation__n2573 , _f_permutation__n2572 ,
         _f_permutation__n2571 , _f_permutation__n2570 ,
         _f_permutation__n2569 , _f_permutation__n2568 ,
         _f_permutation__n2567 , _f_permutation__n2566 ,
         _f_permutation__n2565 , _f_permutation__n2564 ,
         _f_permutation__n2563 , _f_permutation__n2562 ,
         _f_permutation__n2561 , _f_permutation__n2560 ,
         _f_permutation__n2559 , _f_permutation__n2558 ,
         _f_permutation__n2557 , _f_permutation__n2556 ,
         _f_permutation__n2555 , _f_permutation__n2554 ,
         _f_permutation__n2553 , _f_permutation__n2552 ,
         _f_permutation__n2551 , _f_permutation__n2550 ,
         _f_permutation__n2549 , _f_permutation__n2548 ,
         _f_permutation__n2547 , _f_permutation__n2546 ,
         _f_permutation__n2545 , _f_permutation__n2544 ,
         _f_permutation__n2543 , _f_permutation__n2542 ,
         _f_permutation__n2541 , _f_permutation__n2540 ,
         _f_permutation__n2539 , _f_permutation__n2538 ,
         _f_permutation__n2537 , _f_permutation__n2536 ,
         _f_permutation__n2535 , _f_permutation__n2534 ,
         _f_permutation__n2533 , _f_permutation__n2532 ,
         _f_permutation__n2531 , _f_permutation__n2530 ,
         _f_permutation__n2529 , _f_permutation__n2528 ,
         _f_permutation__n2527 , _f_permutation__n2526 ,
         _f_permutation__n2525 , _f_permutation__n2524 ,
         _f_permutation__n2523 , _f_permutation__n2522 ,
         _f_permutation__n2521 , _f_permutation__n2520 ,
         _f_permutation__n2519 , _f_permutation__n2518 ,
         _f_permutation__n2517 , _f_permutation__n2516 ,
         _f_permutation__n2515 , _f_permutation__n2514 ,
         _f_permutation__n2513 , _f_permutation__n2512 ,
         _f_permutation__n2511 , _f_permutation__n2510 ,
         _f_permutation__n2509 , _f_permutation__n2508 ,
         _f_permutation__n2507 , _f_permutation__n2506 ,
         _f_permutation__n2505 , _f_permutation__n2504 ,
         _f_permutation__n2503 , _f_permutation__n2502 ,
         _f_permutation__n2501 , _f_permutation__n2500 ,
         _f_permutation__n2499 , _f_permutation__n2498 ,
         _f_permutation__n2497 , _f_permutation__n2496 ,
         _f_permutation__n2495 , _f_permutation__n2494 ,
         _f_permutation__n2493 , _f_permutation__n2492 ,
         _f_permutation__n2491 , _f_permutation__n2490 ,
         _f_permutation__n2489 , _f_permutation__n2488 ,
         _f_permutation__n2487 , _f_permutation__n2486 ,
         _f_permutation__n2485 , _f_permutation__n2484 ,
         _f_permutation__n2483 , _f_permutation__n2482 ,
         _f_permutation__n2481 , _f_permutation__n2480 ,
         _f_permutation__n2479 , _f_permutation__n2478 ,
         _f_permutation__n2477 , _f_permutation__n2476 ,
         _f_permutation__n2475 , _f_permutation__n2474 ,
         _f_permutation__n2473 , _f_permutation__n2472 ,
         _f_permutation__n2471 , _f_permutation__n2470 ,
         _f_permutation__n2469 , _f_permutation__n2468 ,
         _f_permutation__n2467 , _f_permutation__n2466 ,
         _f_permutation__n2465 , _f_permutation__n2464 ,
         _f_permutation__n2463 , _f_permutation__n2462 ,
         _f_permutation__n2461 , _f_permutation__n2460 ,
         _f_permutation__n2459 , _f_permutation__n2458 ,
         _f_permutation__n2457 , _f_permutation__n2456 ,
         _f_permutation__n2455 , _f_permutation__n2454 ,
         _f_permutation__n2453 , _f_permutation__n2452 ,
         _f_permutation__n2451 , _f_permutation__n2450 ,
         _f_permutation__n2449 , _f_permutation__n2448 ,
         _f_permutation__n2447 , _f_permutation__n2446 ,
         _f_permutation__n2445 , _f_permutation__n2444 ,
         _f_permutation__n2443 , _f_permutation__n2442 ,
         _f_permutation__n2441 , _f_permutation__n2440 ,
         _f_permutation__n2439 , _f_permutation__n2438 ,
         _f_permutation__n2437 , _f_permutation__n2436 ,
         _f_permutation__n2435 , _f_permutation__n2434 ,
         _f_permutation__n2433 , _f_permutation__n2432 ,
         _f_permutation__n2431 , _f_permutation__n2430 ,
         _f_permutation__n2429 , _f_permutation__n2428 ,
         _f_permutation__n2427 , _f_permutation__n2426 ,
         _f_permutation__n2425 , _f_permutation__n2424 ,
         _f_permutation__n2423 , _f_permutation__n2422 ,
         _f_permutation__n2421 , _f_permutation__n2420 ,
         _f_permutation__n2419 , _f_permutation__n2418 ,
         _f_permutation__n2417 , _f_permutation__n2416 ,
         _f_permutation__n2415 , _f_permutation__n2414 ,
         _f_permutation__n2413 , _f_permutation__n2412 ,
         _f_permutation__n2411 , _f_permutation__n2410 ,
         _f_permutation__n2409 , _f_permutation__n2408 ,
         _f_permutation__n2407 , _f_permutation__n2406 ,
         _f_permutation__n2405 , _f_permutation__n2404 ,
         _f_permutation__n2403 , _f_permutation__n2402 ,
         _f_permutation__n2401 , _f_permutation__n2400 ,
         _f_permutation__n2399 , _f_permutation__n2398 ,
         _f_permutation__n2397 , _f_permutation__n2396 ,
         _f_permutation__n2395 , _f_permutation__n2394 ,
         _f_permutation__n2393 , _f_permutation__n2392 ,
         _f_permutation__n2391 , _f_permutation__n2390 ,
         _f_permutation__n2389 , _f_permutation__n2388 ,
         _f_permutation__n2387 , _f_permutation__n2386 ,
         _f_permutation__n2385 , _f_permutation__n2384 ,
         _f_permutation__n2383 , _f_permutation__n2382 ,
         _f_permutation__n2381 , _f_permutation__n2380 ,
         _f_permutation__n2379 , _f_permutation__n2378 ,
         _f_permutation__n2377 , _f_permutation__n2376 ,
         _f_permutation__n2375 , _f_permutation__n2374 ,
         _f_permutation__n2373 , _f_permutation__n2372 ,
         _f_permutation__n2371 , _f_permutation__n2370 ,
         _f_permutation__n2369 , _f_permutation__n2368 ,
         _f_permutation__n2367 , _f_permutation__n2366 ,
         _f_permutation__n2365 , _f_permutation__n2364 ,
         _f_permutation__n2363 , _f_permutation__n2362 ,
         _f_permutation__n2361 , _f_permutation__n2360 ,
         _f_permutation__n2359 , _f_permutation__n2358 ,
         _f_permutation__n2357 , _f_permutation__n2356 ,
         _f_permutation__n2355 , _f_permutation__n2354 ,
         _f_permutation__n2353 , _f_permutation__n2352 ,
         _f_permutation__n2351 , _f_permutation__n2350 ,
         _f_permutation__n2349 , _f_permutation__n2348 ,
         _f_permutation__n2347 , _f_permutation__n2346 ,
         _f_permutation__n2345 , _f_permutation__n2344 ,
         _f_permutation__n2343 , _f_permutation__n2342 ,
         _f_permutation__n2341 , _f_permutation__n2340 ,
         _f_permutation__n2339 , _f_permutation__n2338 ,
         _f_permutation__n2337 , _f_permutation__n2336 ,
         _f_permutation__n2335 , _f_permutation__n2334 ,
         _f_permutation__n2333 , _f_permutation__n2332 ,
         _f_permutation__n2331 , _f_permutation__n2330 ,
         _f_permutation__n2329 , _f_permutation__n2328 ,
         _f_permutation__n2327 , _f_permutation__n2326 ,
         _f_permutation__n2325 , _f_permutation__n2324 ,
         _f_permutation__n2323 , _f_permutation__n2322 ,
         _f_permutation__n2321 , _f_permutation__n2320 ,
         _f_permutation__n2319 , _f_permutation__n2318 ,
         _f_permutation__n2317 , _f_permutation__n2316 ,
         _f_permutation__n2315 , _f_permutation__n2314 ,
         _f_permutation__n2313 , _f_permutation__n2312 ,
         _f_permutation__n2311 , _f_permutation__n2310 ,
         _f_permutation__n2309 , _f_permutation__n2308 ,
         _f_permutation__n2307 , _f_permutation__n2306 ,
         _f_permutation__n2305 , _f_permutation__n2304 ,
         _f_permutation__n2303 , _f_permutation__n2302 ,
         _f_permutation__n2301 , _f_permutation__n2300 ,
         _f_permutation__n2299 , _f_permutation__n2298 ,
         _f_permutation__n2297 , _f_permutation__n2296 ,
         _f_permutation__n2295 , _f_permutation__n2294 ,
         _f_permutation__n2293 , _f_permutation__n2292 ,
         _f_permutation__n2291 , _f_permutation__n2290 ,
         _f_permutation__n2289 , _f_permutation__n2288 ,
         _f_permutation__n2287 , _f_permutation__n2286 ,
         _f_permutation__n2285 , _f_permutation__n2284 ,
         _f_permutation__n2283 , _f_permutation__n2282 ,
         _f_permutation__n2281 , _f_permutation__n2280 ,
         _f_permutation__n2279 , _f_permutation__n2278 ,
         _f_permutation__n2277 , _f_permutation__n2276 ,
         _f_permutation__n2275 , _f_permutation__n2274 ,
         _f_permutation__n2273 , _f_permutation__n2272 ,
         _f_permutation__n2271 , _f_permutation__n2270 ,
         _f_permutation__n2269 , _f_permutation__n2268 ,
         _f_permutation__n2267 , _f_permutation__n2266 ,
         _f_permutation__n2265 , _f_permutation__n2264 ,
         _f_permutation__n2263 , _f_permutation__n2262 ,
         _f_permutation__n2261 , _f_permutation__n2260 ,
         _f_permutation__n2259 , _f_permutation__n2258 ,
         _f_permutation__n2257 , _f_permutation__n2256 ,
         _f_permutation__n2255 , _f_permutation__n2254 ,
         _f_permutation__n2253 , _f_permutation__n2252 ,
         _f_permutation__n2251 , _f_permutation__n2250 ,
         _f_permutation__n2249 , _f_permutation__n2248 ,
         _f_permutation__n2247 , _f_permutation__n2246 ,
         _f_permutation__n2245 , _f_permutation__n2244 ,
         _f_permutation__n2243 , _f_permutation__n2242 ,
         _f_permutation__n2241 , _f_permutation__n2240 ,
         _f_permutation__n2239 , _f_permutation__n2238 ,
         _f_permutation__n2237 , _f_permutation__n2236 ,
         _f_permutation__n2235 , _f_permutation__n2234 ,
         _f_permutation__n2233 , _f_permutation__n2232 ,
         _f_permutation__n2231 , _f_permutation__n2230 ,
         _f_permutation__n2229 , _f_permutation__n2228 ,
         _f_permutation__n2227 , _f_permutation__n2226 ,
         _f_permutation__n2225 , _f_permutation__n2224 ,
         _f_permutation__n2223 , _f_permutation__n2222 ,
         _f_permutation__n2221 , _f_permutation__n2220 ,
         _f_permutation__n2219 , _f_permutation__n2218 ,
         _f_permutation__n2217 , _f_permutation__n2216 ,
         _f_permutation__n2215 , _f_permutation__n2214 ,
         _f_permutation__n2211 , _f_permutation__n2210 ,
         _f_permutation__n2209 , _f_permutation__n2208 ,
         _f_permutation__n2207 , _f_permutation__n2206 ,
         _f_permutation__n2205 , _f_permutation__n2204 ,
         _f_permutation__n2203 , _f_permutation__n2202 ,
         _f_permutation__n2201 , _f_permutation__n2200 ,
         _f_permutation__n2199 , _f_permutation__n2198 ,
         _f_permutation__n2197 , _f_permutation__n2196 ,
         _f_permutation__n2195 , _f_permutation__n2194 ,
         _f_permutation__n2193 , _f_permutation__n2192 ,
         _f_permutation__n2191 , _f_permutation__n2190 ,
         _f_permutation__n2189 , _f_permutation__n2188 ,
         _f_permutation__n2187 , _f_permutation__n2186 ,
         _f_permutation__n2185 , _f_permutation__n2184 ,
         _f_permutation__n2183 , _f_permutation__n2182 ,
         _f_permutation__n2181 , _f_permutation__n2180 ,
         _f_permutation__n2179 , _f_permutation__n2178 ,
         _f_permutation__n2177 , _f_permutation__n2176 ,
         _f_permutation__n2175 , _f_permutation__n2174 ,
         _f_permutation__n2173 , _f_permutation__n2172 ,
         _f_permutation__n2171 , _f_permutation__n2170 ,
         _f_permutation__n2169 , _f_permutation__n2168 ,
         _f_permutation__n2167 , _f_permutation__n2166 ,
         _f_permutation__n2165 , _f_permutation__n2164 ,
         _f_permutation__n2163 , _f_permutation__n2162 ,
         _f_permutation__n2161 , _f_permutation__n2160 ,
         _f_permutation__n2159 , _f_permutation__n2158 ,
         _f_permutation__n2157 , _f_permutation__n2156 ,
         _f_permutation__n2155 , _f_permutation__n2154 ,
         _f_permutation__n2153 , _f_permutation__n2152 ,
         _f_permutation__n2151 , _f_permutation__n2150 ,
         _f_permutation__n2149 , _f_permutation__n2148 ,
         _f_permutation__n2147 , _f_permutation__n2146 ,
         _f_permutation__n2145 , _f_permutation__n2144 ,
         _f_permutation__n2143 , _f_permutation__n2142 ,
         _f_permutation__n2141 , _f_permutation__n2140 ,
         _f_permutation__n2139 , _f_permutation__n2138 ,
         _f_permutation__n2137 , _f_permutation__n2136 ,
         _f_permutation__n2135 , _f_permutation__n2134 ,
         _f_permutation__n2133 , _f_permutation__n2132 ,
         _f_permutation__n2131 , _f_permutation__n2130 ,
         _f_permutation__n2129 , _f_permutation__n2128 ,
         _f_permutation__n2127 , _f_permutation__n2126 ,
         _f_permutation__n2125 , _f_permutation__n2124 ,
         _f_permutation__n2123 , _f_permutation__n2122 ,
         _f_permutation__n2121 , _f_permutation__n2120 ,
         _f_permutation__n2119 , _f_permutation__n2118 ,
         _f_permutation__n2117 , _f_permutation__n2116 ,
         _f_permutation__n2115 , _f_permutation__n2114 ,
         _f_permutation__n2113 , _f_permutation__n2112 ,
         _f_permutation__n2111 , _f_permutation__n2110 ,
         _f_permutation__n2109 , _f_permutation__n2108 ,
         _f_permutation__n2107 , _f_permutation__n2106 ,
         _f_permutation__n2105 , _f_permutation__n2104 ,
         _f_permutation__n2103 , _f_permutation__n2102 ,
         _f_permutation__n2101 , _f_permutation__n2100 ,
         _f_permutation__n2099 , _f_permutation__n2098 ,
         _f_permutation__n2097 , _f_permutation__n2096 ,
         _f_permutation__n2095 , _f_permutation__n2094 ,
         _f_permutation__n2093 , _f_permutation__n2092 ,
         _f_permutation__n2091 , _f_permutation__n2090 ,
         _f_permutation__n2089 , _f_permutation__n2088 ,
         _f_permutation__n2087 , _f_permutation__n2086 ,
         _f_permutation__n2085 , _f_permutation__n2084 ,
         _f_permutation__n2083 , _f_permutation__n2082 ,
         _f_permutation__n2081 , _f_permutation__n2080 ,
         _f_permutation__n2079 , _f_permutation__n2078 ,
         _f_permutation__n2077 , _f_permutation__n2076 ,
         _f_permutation__n2075 , _f_permutation__n2074 ,
         _f_permutation__n2073 , _f_permutation__n2072 ,
         _f_permutation__n2071 , _f_permutation__n2070 ,
         _f_permutation__n2069 , _f_permutation__n2068 ,
         _f_permutation__n2067 , _f_permutation__n2066 ,
         _f_permutation__n2065 , _f_permutation__n2064 ,
         _f_permutation__n2063 , _f_permutation__n2062 ,
         _f_permutation__n2061 , _f_permutation__n2060 ,
         _f_permutation__n2059 , _f_permutation__n2058 ,
         _f_permutation__n2057 , _f_permutation__n2056 ,
         _f_permutation__n2055 , _f_permutation__n2054 ,
         _f_permutation__n2053 , _f_permutation__n2052 ,
         _f_permutation__n2051 , _f_permutation__n2050 ,
         _f_permutation__n2049 , _f_permutation__n2048 ,
         _f_permutation__n2047 , _f_permutation__n2046 ,
         _f_permutation__n2045 , _f_permutation__n2044 ,
         _f_permutation__n2043 , _f_permutation__n2042 ,
         _f_permutation__n2041 , _f_permutation__n2040 ,
         _f_permutation__n2039 , _f_permutation__n2038 ,
         _f_permutation__n2037 , _f_permutation__n2036 ,
         _f_permutation__n2035 , _f_permutation__n2034 ,
         _f_permutation__n2033 , _f_permutation__n2032 ,
         _f_permutation__n2031 , _f_permutation__n2030 ,
         _f_permutation__n2029 , _f_permutation__n2028 ,
         _f_permutation__n2027 , _f_permutation__n2026 ,
         _f_permutation__n2025 , _f_permutation__n2024 ,
         _f_permutation__n2023 , _f_permutation__n2022 ,
         _f_permutation__n2021 , _f_permutation__n2020 ,
         _f_permutation__n2019 , _f_permutation__n2018 ,
         _f_permutation__n2017 , _f_permutation__n2016 ,
         _f_permutation__n2015 , _f_permutation__n2014 ,
         _f_permutation__n2013 , _f_permutation__n2012 ,
         _f_permutation__n2011 , _f_permutation__n2010 ,
         _f_permutation__n2009 , _f_permutation__n2008 ,
         _f_permutation__n2007 , _f_permutation__n2006 ,
         _f_permutation__n2005 , _f_permutation__n2004 ,
         _f_permutation__n2003 , _f_permutation__n2002 ,
         _f_permutation__n2001 , _f_permutation__n2000 ,
         _f_permutation__n1999 , _f_permutation__n1998 ,
         _f_permutation__n1997 , _f_permutation__n1996 ,
         _f_permutation__n1995 , _f_permutation__n1994 ,
         _f_permutation__n1993 , _f_permutation__n1992 ,
         _f_permutation__n1991 , _f_permutation__n1990 ,
         _f_permutation__n1989 , _f_permutation__n1988 ,
         _f_permutation__n1987 , _f_permutation__n1986 ,
         _f_permutation__n1985 , _f_permutation__n1984 ,
         _f_permutation__n1983 , _f_permutation__n1982 ,
         _f_permutation__n1981 , _f_permutation__n1980 ,
         _f_permutation__n1979 , _f_permutation__n1978 ,
         _f_permutation__n1977 , _f_permutation__n1976 ,
         _f_permutation__n1975 , _f_permutation__n1974 ,
         _f_permutation__n1973 , _f_permutation__n1972 ,
         _f_permutation__n1971 , _f_permutation__n1970 ,
         _f_permutation__n1969 , _f_permutation__n1968 ,
         _f_permutation__n1967 , _f_permutation__n1966 ,
         _f_permutation__n1965 , _f_permutation__n1964 ,
         _f_permutation__n1963 , _f_permutation__n1962 ,
         _f_permutation__n1961 , _f_permutation__n1960 ,
         _f_permutation__n1959 , _f_permutation__n1958 ,
         _f_permutation__n1957 , _f_permutation__n1956 ,
         _f_permutation__n1955 , _f_permutation__n1954 ,
         _f_permutation__n1953 , _f_permutation__n1952 ,
         _f_permutation__n1951 , _f_permutation__n1950 ,
         _f_permutation__n1949 , _f_permutation__n1948 ,
         _f_permutation__n1947 , _f_permutation__n1946 ,
         _f_permutation__n1945 , _f_permutation__n1944 ,
         _f_permutation__n1943 , _f_permutation__n1942 ,
         _f_permutation__n1941 , _f_permutation__n1940 ,
         _f_permutation__n1939 , _f_permutation__n1938 ,
         _f_permutation__n1937 , _f_permutation__n1936 ,
         _f_permutation__n1935 , _f_permutation__n1934 ,
         _f_permutation__n1933 , _f_permutation__n1932 ,
         _f_permutation__n1931 , _f_permutation__n1930 ,
         _f_permutation__n1929 , _f_permutation__n1928 ,
         _f_permutation__n1927 , _f_permutation__n1926 ,
         _f_permutation__n1925 , _f_permutation__n1924 ,
         _f_permutation__n1923 , _f_permutation__n1922 ,
         _f_permutation__n1921 , _f_permutation__n1920 ,
         _f_permutation__n1919 , _f_permutation__n1918 ,
         _f_permutation__n1917 , _f_permutation__n1916 ,
         _f_permutation__n1915 , _f_permutation__n1914 ,
         _f_permutation__n1913 , _f_permutation__n1912 ,
         _f_permutation__n1911 , _f_permutation__n1910 ,
         _f_permutation__n1909 , _f_permutation__n1908 ,
         _f_permutation__n1907 , _f_permutation__n1906 ,
         _f_permutation__n1905 , _f_permutation__n1904 ,
         _f_permutation__n1903 , _f_permutation__n1902 ,
         _f_permutation__n1901 , _f_permutation__n1900 ,
         _f_permutation__n1899 , _f_permutation__n1898 ,
         _f_permutation__n1897 , _f_permutation__n1896 ,
         _f_permutation__n1895 , _f_permutation__n1894 ,
         _f_permutation__n1893 , _f_permutation__n1892 ,
         _f_permutation__n1891 , _f_permutation__n1890 ,
         _f_permutation__n1889 , _f_permutation__n1888 ,
         _f_permutation__n1887 , _f_permutation__n1886 ,
         _f_permutation__n1885 , _f_permutation__n1884 ,
         _f_permutation__n1883 , _f_permutation__n1882 ,
         _f_permutation__n1881 , _f_permutation__n1880 ,
         _f_permutation__n1879 , _f_permutation__n1878 ,
         _f_permutation__n1877 , _f_permutation__n1876 ,
         _f_permutation__n1875 , _f_permutation__n1874 ,
         _f_permutation__n1873 , _f_permutation__n1872 ,
         _f_permutation__n1871 , _f_permutation__n1870 ,
         _f_permutation__n1869 , _f_permutation__n1868 ,
         _f_permutation__n1867 , _f_permutation__n1866 ,
         _f_permutation__n1865 , _f_permutation__n1864 ,
         _f_permutation__n1863 , _f_permutation__n1862 ,
         _f_permutation__n1861 , _f_permutation__n1860 ,
         _f_permutation__n1859 , _f_permutation__n1858 ,
         _f_permutation__n1857 , _f_permutation__n1856 ,
         _f_permutation__n1855 , _f_permutation__n1854 ,
         _f_permutation__n1853 , _f_permutation__n1852 ,
         _f_permutation__n1851 , _f_permutation__n1850 ,
         _f_permutation__n1849 , _f_permutation__n1848 ,
         _f_permutation__n1847 , _f_permutation__n1846 ,
         _f_permutation__n1845 , _f_permutation__n1844 ,
         _f_permutation__n1843 , _f_permutation__n1842 ,
         _f_permutation__n1841 , _f_permutation__n1840 ,
         _f_permutation__n1839 , _f_permutation__n1838 ,
         _f_permutation__n1837 , _f_permutation__n1836 ,
         _f_permutation__n1835 , _f_permutation__n1834 ,
         _f_permutation__n1833 , _f_permutation__n1832 ,
         _f_permutation__n1831 , _f_permutation__n1830 ,
         _f_permutation__n1829 , _f_permutation__n1828 ,
         _f_permutation__n1827 , _f_permutation__n1826 ,
         _f_permutation__n1825 , _f_permutation__n1824 ,
         _f_permutation__n1823 , _f_permutation__n1822 ,
         _f_permutation__n1821 , _f_permutation__n1820 ,
         _f_permutation__n1819 , _f_permutation__n1818 ,
         _f_permutation__n1817 , _f_permutation__n1816 ,
         _f_permutation__n1815 , _f_permutation__n1814 ,
         _f_permutation__n1813 , _f_permutation__n1812 ,
         _f_permutation__n1811 , _f_permutation__n1810 ,
         _f_permutation__n1809 , _f_permutation__n1808 ,
         _f_permutation__n1807 , _f_permutation__n1806 ,
         _f_permutation__n1805 , _f_permutation__n1804 ,
         _f_permutation__n1803 , _f_permutation__n1802 ,
         _f_permutation__n1801 , _f_permutation__n1800 ,
         _f_permutation__n1799 , _f_permutation__n1798 ,
         _f_permutation__n1797 , _f_permutation__n1796 ,
         _f_permutation__n1795 , _f_permutation__n1794 ,
         _f_permutation__n1793 , _f_permutation__n1792 ,
         _f_permutation__n1791 , _f_permutation__n1790 ,
         _f_permutation__n1789 , _f_permutation__n1788 ,
         _f_permutation__n1787 , _f_permutation__n1786 ,
         _f_permutation__n1785 , _f_permutation__n1784 ,
         _f_permutation__n1783 , _f_permutation__n1782 ,
         _f_permutation__n1781 , _f_permutation__n1780 ,
         _f_permutation__n1779 , _f_permutation__n1778 ,
         _f_permutation__n1777 , _f_permutation__n1776 ,
         _f_permutation__n1775 , _f_permutation__n1774 ,
         _f_permutation__n1773 , _f_permutation__n1772 ,
         _f_permutation__n1771 , _f_permutation__n1770 ,
         _f_permutation__n1769 , _f_permutation__n1768 ,
         _f_permutation__n1767 , _f_permutation__n1766 ,
         _f_permutation__n1765 , _f_permutation__n1764 ,
         _f_permutation__n1763 , _f_permutation__n1762 ,
         _f_permutation__n1761 , _f_permutation__n1760 ,
         _f_permutation__n1759 , _f_permutation__n1758 ,
         _f_permutation__n1757 , _f_permutation__n1756 ,
         _f_permutation__n1755 , _f_permutation__n1754 ,
         _f_permutation__n1753 , _f_permutation__n1752 ,
         _f_permutation__n1751 , _f_permutation__n1750 ,
         _f_permutation__n1749 , _f_permutation__n1748 ,
         _f_permutation__n1747 , _f_permutation__n1746 ,
         _f_permutation__n1745 , _f_permutation__n1744 ,
         _f_permutation__n1743 , _f_permutation__n1742 ,
         _f_permutation__n1741 , _f_permutation__n1740 ,
         _f_permutation__n1739 , _f_permutation__n1738 ,
         _f_permutation__n1737 , _f_permutation__n1736 ,
         _f_permutation__n1735 , _f_permutation__n1734 ,
         _f_permutation__n1733 , _f_permutation__n1732 ,
         _f_permutation__n1731 , _f_permutation__n1730 ,
         _f_permutation__n1729 , _f_permutation__n1728 ,
         _f_permutation__n1727 , _f_permutation__n1726 ,
         _f_permutation__n1725 , _f_permutation__n1724 ,
         _f_permutation__n1723 , _f_permutation__n1722 ,
         _f_permutation__n1721 , _f_permutation__n1720 ,
         _f_permutation__n1719 , _f_permutation__n1718 ,
         _f_permutation__n1717 , _f_permutation__n1716 ,
         _f_permutation__n1715 , _f_permutation__n1714 ,
         _f_permutation__n1713 , _f_permutation__n1712 ,
         _f_permutation__n1711 , _f_permutation__n1710 ,
         _f_permutation__n1709 , _f_permutation__n1708 ,
         _f_permutation__n1707 , _f_permutation__n1706 ,
         _f_permutation__n1705 , _f_permutation__n1704 ,
         _f_permutation__n1703 , _f_permutation__n1702 ,
         _f_permutation__n1701 , _f_permutation__n1700 ,
         _f_permutation__n1699 , _f_permutation__n1698 ,
         _f_permutation__n1697 , _f_permutation__n1696 ,
         _f_permutation__n1695 , _f_permutation__n1694 ,
         _f_permutation__n1693 , _f_permutation__n1692 ,
         _f_permutation__n1691 , _f_permutation__n1690 ,
         _f_permutation__n1689 , _f_permutation__n1688 ,
         _f_permutation__n1687 , _f_permutation__n1686 ,
         _f_permutation__n1685 , _f_permutation__n1684 ,
         _f_permutation__n1683 , _f_permutation__n1682 ,
         _f_permutation__n1681 , _f_permutation__n1680 ,
         _f_permutation__n1679 , _f_permutation__n1678 ,
         _f_permutation__n1677 , _f_permutation__n1676 ,
         _f_permutation__n1675 , _f_permutation__n1674 ,
         _f_permutation__n1673 , _f_permutation__n1672 ,
         _f_permutation__n1671 , _f_permutation__n1670 ,
         _f_permutation__n1669 , _f_permutation__n1668 ,
         _f_permutation__n1667 , _f_permutation__n1666 ,
         _f_permutation__n1665 , _f_permutation__n1664 ,
         _f_permutation__n1663 , _f_permutation__n1662 ,
         _f_permutation__n1661 , _f_permutation__n1660 ,
         _f_permutation__n1659 , _f_permutation__n1658 ,
         _f_permutation__n1657 , _f_permutation__n1656 ,
         _f_permutation__n1655 , _f_permutation__n1654 ,
         _f_permutation__n1653 , _f_permutation__n1652 ,
         _f_permutation__n1651 , _f_permutation__n1650 ,
         _f_permutation__n1649 , _f_permutation__n1648 ,
         _f_permutation__n1647 , _f_permutation__n1646 ,
         _f_permutation__n1645 , _f_permutation__n1644 ,
         _f_permutation__n1643 , _f_permutation__n1642 ,
         _f_permutation__n1641 , _f_permutation__n1640 ,
         _f_permutation__n1639 , _f_permutation__n1638 ,
         _f_permutation__n1637 , _f_permutation__n1636 ,
         _f_permutation__n1635 , _f_permutation__n1634 ,
         _f_permutation__n1633 , _f_permutation__n1632 ,
         _f_permutation__n1628 , _f_permutation__n5804 ,
         _f_permutation__n5803 , _f_permutation__n5802 ,
         _f_permutation__n5801 , _f_permutation__n5800 ,
         _f_permutation__n5799 , _f_permutation__n5798 ,
         _f_permutation__n5797 , _f_permutation__n5796 ,
         _f_permutation__n5795 , _f_permutation__n5794 ,
         _f_permutation__n5793 , _f_permutation__n5792 ,
         _f_permutation__n5791 , _f_permutation__n5790 ,
         _f_permutation__n5789 , _f_permutation__n5788 ,
         _f_permutation__n5787 , _f_permutation__n5786 ,
         _f_permutation__n5785 , _f_permutation__n5784 ,
         _f_permutation__n5783 , _f_permutation__n5782 , _f_permutation__n3 ,
         _f_permutation__n5388 , _f_permutation__n5387 ,
         _f_permutation__n5386 , _f_permutation__n5385 ,
         _f_permutation__n5384 , _f_permutation__n5383 ,
         _f_permutation__n5382 , _f_permutation__n5381 ,
         _f_permutation__n5380 , _f_permutation__n5379 ,
         _f_permutation__n5378 , _f_permutation__n5377 ,
         _f_permutation__n5376 , _f_permutation__n5375 ,
         _f_permutation__n5374 , _f_permutation__n5373 ,
         _f_permutation__n5372 , _f_permutation__n5371 ,
         _f_permutation__n5370 , _f_permutation__n5369 ,
         _f_permutation__n5368 , _f_permutation__n5367 ,
         _f_permutation__n5366 , _f_permutation__n5365 ,
         _f_permutation__n5364 , _f_permutation__n5363 ,
         _f_permutation__n5362 , _f_permutation__n5361 ,
         _f_permutation__n5360 , _f_permutation__n5359 ,
         _f_permutation__n5358 , _f_permutation__n5357 ,
         _f_permutation__n5356 , _f_permutation__n5355 ,
         _f_permutation__n5354 , _f_permutation__n5353 ,
         _f_permutation__n5352 , _f_permutation__n5351 ,
         _f_permutation__n5350 , _f_permutation__n5349 ,
         _f_permutation__n5348 , _f_permutation__n5347 ,
         _f_permutation__n5346 , _f_permutation__n5345 ,
         _f_permutation__n5344 , _f_permutation__n5343 ,
         _f_permutation__n5342 , _f_permutation__n5341 ,
         _f_permutation__n5340 , _f_permutation__n5339 ,
         _f_permutation__n5338 , _f_permutation__n5337 ,
         _f_permutation__n5336 , _f_permutation__n5335 ,
         _f_permutation__n5334 , _f_permutation__n5333 ,
         _f_permutation__n5332 , _f_permutation__n5331 ,
         _f_permutation__n5330 , _f_permutation__n5329 ,
         _f_permutation__n5328 , _f_permutation__n5327 ,
         _f_permutation__n5326 , _f_permutation__n5325 ,
         _f_permutation__n5324 , _f_permutation__n5323 ,
         _f_permutation__n5322 , _f_permutation__n5321 ,
         _f_permutation__n5320 , _f_permutation__n5319 ,
         _f_permutation__n5318 , _f_permutation__n5317 ,
         _f_permutation__n5316 , _f_permutation__n5315 ,
         _f_permutation__n5314 , _f_permutation__n5313 ,
         _f_permutation__n5312 , _f_permutation__n5311 ,
         _f_permutation__n5310 , _f_permutation__n5309 ,
         _f_permutation__n5308 , _f_permutation__n5307 ,
         _f_permutation__n5306 , _f_permutation__n5305 ,
         _f_permutation__n5304 , _f_permutation__n5303 ,
         _f_permutation__n5302 , _f_permutation__n5301 ,
         _f_permutation__n5300 , _f_permutation__n5299 ,
         _f_permutation__n5298 , _f_permutation__n5297 ,
         _f_permutation__n5296 , _f_permutation__n5295 ,
         _f_permutation__n5294 , _f_permutation__n5293 ,
         _f_permutation__n5292 , _f_permutation__n5291 ,
         _f_permutation__n5290 , _f_permutation__n5289 ,
         _f_permutation__n5288 , _f_permutation__n5287 ,
         _f_permutation__n5286 , _f_permutation__n5285 ,
         _f_permutation__n5284 , _f_permutation__n5283 ,
         _f_permutation__n5282 , _f_permutation__n5281 ,
         _f_permutation__n5280 , _f_permutation__n5279 ,
         _f_permutation__n5278 , _f_permutation__n5277 ,
         _f_permutation__n5276 , _f_permutation__n5275 ,
         _f_permutation__n5274 , _f_permutation__n5273 ,
         _f_permutation__n5272 , _f_permutation__n5271 ,
         _f_permutation__n5270 , _f_permutation__n5269 ,
         _f_permutation__n5268 , _f_permutation__n5267 ,
         _f_permutation__n5266 , _f_permutation__n5265 ,
         _f_permutation__n5264 , _f_permutation__n5263 ,
         _f_permutation__n5262 , _f_permutation__n5261 ,
         _f_permutation__n5260 , _f_permutation__n5259 ,
         _f_permutation__n5258 , _f_permutation__n5257 ,
         _f_permutation__n5256 , _f_permutation__n5255 ,
         _f_permutation__n5254 , _f_permutation__n5253 ,
         _f_permutation__n5252 , _f_permutation__n5251 ,
         _f_permutation__n5250 , _f_permutation__n5249 ,
         _f_permutation__n5248 , _f_permutation__n5247 ,
         _f_permutation__n5246 , _f_permutation__n5245 ,
         _f_permutation__n5244 , _f_permutation__n5243 ,
         _f_permutation__n5242 , _f_permutation__n5241 ,
         _f_permutation__n5240 , _f_permutation__n5239 ,
         _f_permutation__n5238 , _f_permutation__n5237 ,
         _f_permutation__n5236 , _f_permutation__n5235 ,
         _f_permutation__n5234 , _f_permutation__n5233 ,
         _f_permutation__n5232 , _f_permutation__n5231 ,
         _f_permutation__n5230 , _f_permutation__n5229 ,
         _f_permutation__n5228 , _f_permutation__n5227 ,
         _f_permutation__n5226 , _f_permutation__n5225 ,
         _f_permutation__n5224 , _f_permutation__n5223 ,
         _f_permutation__n5222 , _f_permutation__n5221 ,
         _f_permutation__n5220 , _f_permutation__n5219 ,
         _f_permutation__n5218 , _f_permutation__n5217 ,
         _f_permutation__n5216 , _f_permutation__n5215 ,
         _f_permutation__n5214 , _f_permutation__n5213 ,
         _f_permutation__n5212 , _f_permutation__n5211 ,
         _f_permutation__n5210 , _f_permutation__n5209 ,
         _f_permutation__n5208 , _f_permutation__n5207 ,
         _f_permutation__n5206 , _f_permutation__n5205 ,
         _f_permutation__n5204 , _f_permutation__n5203 ,
         _f_permutation__n5202 , _f_permutation__n5201 ,
         _f_permutation__n5200 , _f_permutation__n5199 ,
         _f_permutation__n5198 , _f_permutation__n5197 ,
         _f_permutation__n5196 , _f_permutation__n5195 ,
         _f_permutation__n5194 , _f_permutation__n5193 ,
         _f_permutation__n5192 , _f_permutation__n5191 ,
         _f_permutation__n5190 , _f_permutation__n5189 ,
         _f_permutation__n5188 , _f_permutation__n5187 ,
         _f_permutation__n5186 , _f_permutation__n5185 ,
         _f_permutation__n5184 , _f_permutation__n5183 ,
         _f_permutation__n5182 , _f_permutation__n5181 ,
         _f_permutation__n5180 , _f_permutation__n5179 ,
         _f_permutation__n5178 , _f_permutation__n5177 ,
         _f_permutation__n5176 , _f_permutation__n5175 ,
         _f_permutation__n5174 , _f_permutation__n5173 ,
         _f_permutation__n5172 , _f_permutation__n5171 ,
         _f_permutation__n5170 , _f_permutation__n5169 ,
         _f_permutation__n5168 , _f_permutation__n5167 ,
         _f_permutation__n5166 , _f_permutation__n5165 ,
         _f_permutation__n5164 , _f_permutation__n5163 ,
         _f_permutation__n5162 , _f_permutation__n5161 ,
         _f_permutation__n5160 , _f_permutation__n5159 ,
         _f_permutation__n5158 , _f_permutation__n5157 ,
         _f_permutation__n5156 , _f_permutation__n5155 ,
         _f_permutation__n5154 , _f_permutation__n5153 ,
         _f_permutation__n5152 , _f_permutation__n5151 ,
         _f_permutation__n5150 , _f_permutation__n5149 ,
         _f_permutation__n5148 , _f_permutation__n5147 ,
         _f_permutation__n5146 , _f_permutation__n5145 ,
         _f_permutation__n5144 , _f_permutation__n5143 ,
         _f_permutation__n5142 , _f_permutation__n5141 ,
         _f_permutation__n5140 , _f_permutation__n5139 ,
         _f_permutation__n5138 , _f_permutation__n5137 ,
         _f_permutation__n5136 , _f_permutation__n5135 ,
         _f_permutation__n5134 , _f_permutation__n5133 ,
         _f_permutation__n5132 , _f_permutation__n5131 ,
         _f_permutation__n5130 , _f_permutation__n5129 ,
         _f_permutation__n5128 , _f_permutation__n5127 ,
         _f_permutation__n5126 , _f_permutation__n5125 ,
         _f_permutation__n5124 , _f_permutation__n5123 ,
         _f_permutation__n5122 , _f_permutation__n5121 ,
         _f_permutation__n5120 , _f_permutation__n5119 ,
         _f_permutation__n5118 , _f_permutation__n5117 ,
         _f_permutation__n5116 , _f_permutation__n5115 ,
         _f_permutation__n5114 , _f_permutation__n5113 ,
         _f_permutation__n5112 , _f_permutation__n5111 ,
         _f_permutation__n5110 , _f_permutation__n5109 ,
         _f_permutation__n5108 , _f_permutation__n5107 ,
         _f_permutation__n5106 , _f_permutation__n5105 ,
         _f_permutation__n5104 , _f_permutation__n5103 ,
         _f_permutation__n5102 , _f_permutation__n5101 ,
         _f_permutation__n5100 , _f_permutation__n5099 ,
         _f_permutation__n5098 , _f_permutation__n5097 ,
         _f_permutation__n5096 , _f_permutation__n5095 ,
         _f_permutation__n5094 , _f_permutation__n5093 ,
         _f_permutation__n5092 , _f_permutation__n5091 ,
         _f_permutation__n5090 , _f_permutation__n5089 ,
         _f_permutation__n5088 , _f_permutation__n5087 ,
         _f_permutation__n5086 , _f_permutation__n5085 ,
         _f_permutation__n5084 , _f_permutation__n5083 ,
         _f_permutation__n5082 , _f_permutation__n5081 ,
         _f_permutation__n5080 , _f_permutation__n5079 ,
         _f_permutation__n5078 , _f_permutation__n5077 ,
         _f_permutation__n5076 , _f_permutation__n5075 ,
         _f_permutation__n5074 , _f_permutation__n5073 ,
         _f_permutation__n5072 , _f_permutation__n5071 ,
         _f_permutation__n5070 , _f_permutation__n5069 ,
         _f_permutation__n5068 , _f_permutation__n5067 ,
         _f_permutation__n5066 , _f_permutation__n5065 ,
         _f_permutation__n5064 , _f_permutation__n5063 ,
         _f_permutation__n5062 , _f_permutation__n5061 ,
         _f_permutation__n5060 , _f_permutation__n5059 ,
         _f_permutation__n5058 , _f_permutation__n5057 ,
         _f_permutation__n5056 , _f_permutation__n5055 ,
         _f_permutation__n5054 , _f_permutation__n5053 ,
         _f_permutation__n5052 , _f_permutation__n5051 ,
         _f_permutation__n5050 , _f_permutation__n5049 ,
         _f_permutation__n5048 , _f_permutation__n5047 ,
         _f_permutation__n5046 , _f_permutation__n5045 ,
         _f_permutation__n5044 , _f_permutation__n5043 ,
         _f_permutation__n5042 , _f_permutation__n5041 ,
         _f_permutation__n5040 , _f_permutation__n5039 ,
         _f_permutation__n5038 , _f_permutation__n5037 ,
         _f_permutation__n5036 , _f_permutation__n5035 ,
         _f_permutation__n5034 , _f_permutation__n5033 ,
         _f_permutation__n5032 , _f_permutation__n5031 ,
         _f_permutation__n5030 , _f_permutation__n5029 ,
         _f_permutation__n5028 , _f_permutation__n5027 ,
         _f_permutation__n5026 , _f_permutation__n5025 ,
         _f_permutation__n5024 , _f_permutation__n5023 ,
         _f_permutation__n5022 , _f_permutation__n5021 ,
         _f_permutation__n5020 , _f_permutation__n5019 ,
         _f_permutation__n5018 , _f_permutation__n5017 ,
         _f_permutation__n5016 , _f_permutation__n5015 ,
         _f_permutation__n5014 , _f_permutation__n5013 ,
         _f_permutation__n5012 , _f_permutation__n5011 ,
         _f_permutation__n5010 , _f_permutation__n5009 ,
         _f_permutation__n5008 , _f_permutation__n5007 ,
         _f_permutation__n5006 , _f_permutation__n5005 ,
         _f_permutation__n5004 , _f_permutation__n5003 ,
         _f_permutation__n5002 , _f_permutation__n5001 ,
         _f_permutation__n5000 , _f_permutation__n4999 ,
         _f_permutation__n4998 , _f_permutation__n4997 ,
         _f_permutation__n4996 , _f_permutation__n4995 ,
         _f_permutation__n4994 , _f_permutation__n4993 ,
         _f_permutation__n4992 , _f_permutation__n4991 ,
         _f_permutation__n4990 , _f_permutation__n4989 ,
         _f_permutation__n4988 , _f_permutation__n4987 ,
         _f_permutation__n4986 , _f_permutation__n4985 ,
         _f_permutation__n4984 , _f_permutation__n4983 ,
         _f_permutation__n4982 , _f_permutation__n4981 ,
         _f_permutation__n4980 , _f_permutation__n4979 ,
         _f_permutation__n4978 , _f_permutation__n4977 ,
         _f_permutation__n4976 , _f_permutation__n4975 ,
         _f_permutation__n4974 , _f_permutation__n4973 ,
         _f_permutation__n4972 , _f_permutation__n4971 ,
         _f_permutation__n4970 , _f_permutation__n4969 ,
         _f_permutation__n4968 , _f_permutation__n4967 ,
         _f_permutation__n4966 , _f_permutation__n4965 ,
         _f_permutation__n4964 , _f_permutation__n4963 ,
         _f_permutation__n4962 , _f_permutation__n4961 ,
         _f_permutation__n4960 , _f_permutation__n4959 ,
         _f_permutation__n4958 , _f_permutation__n4957 ,
         _f_permutation__n4956 , _f_permutation__n4955 ,
         _f_permutation__n4954 , _f_permutation__n4953 ,
         _f_permutation__n4952 , _f_permutation__n4951 ,
         _f_permutation__n4950 , _f_permutation__n4949 ,
         _f_permutation__n4948 , _f_permutation__n4947 ,
         _f_permutation__n4946 , _f_permutation__n4945 ,
         _f_permutation__n4944 , _f_permutation__n4943 ,
         _f_permutation__n4942 , _f_permutation__n4941 ,
         _f_permutation__n4940 , _f_permutation__n4939 ,
         _f_permutation__n4938 , _f_permutation__n4937 ,
         _f_permutation__n4936 , _f_permutation__n4935 ,
         _f_permutation__n4934 , _f_permutation__n4933 ,
         _f_permutation__n4932 , _f_permutation__n4931 ,
         _f_permutation__n4930 , _f_permutation__n4929 ,
         _f_permutation__n4928 , _f_permutation__n4927 ,
         _f_permutation__n4926 , _f_permutation__n4925 ,
         _f_permutation__n4924 , _f_permutation__n4923 ,
         _f_permutation__n4922 , _f_permutation__n4921 ,
         _f_permutation__n4920 , _f_permutation__n4919 ,
         _f_permutation__n4918 , _f_permutation__n4917 ,
         _f_permutation__n4916 , _f_permutation__n4915 ,
         _f_permutation__n4914 , _f_permutation__n4913 ,
         _f_permutation__n4912 , _f_permutation__n4911 ,
         _f_permutation__n4910 , _f_permutation__n4909 ,
         _f_permutation__n4908 , _f_permutation__n4907 ,
         _f_permutation__n4906 , _f_permutation__n4905 ,
         _f_permutation__n4904 , _f_permutation__n4903 ,
         _f_permutation__n4902 , _f_permutation__n4901 ,
         _f_permutation__n4900 , _f_permutation__n4899 ,
         _f_permutation__n4898 , _f_permutation__n4897 ,
         _f_permutation__n4896 , _f_permutation__n4895 ,
         _f_permutation__n4894 , _f_permutation__n4893 ,
         _f_permutation__n4892 , _f_permutation__n4891 ,
         _f_permutation__n4890 , _f_permutation__n4889 ,
         _f_permutation__n4888 , _f_permutation__n4887 ,
         _f_permutation__n4886 , _f_permutation__n4885 ,
         _f_permutation__n4884 , _f_permutation__n4883 ,
         _f_permutation__n4882 , _f_permutation__n4881 ,
         _f_permutation__n4880 , _f_permutation__n4879 ,
         _f_permutation__n4878 , _f_permutation__n4877 ,
         _f_permutation__n4876 , _f_permutation__n4875 ,
         _f_permutation__n4874 , _f_permutation__n4873 ,
         _f_permutation__n4872 , _f_permutation__n4871 ,
         _f_permutation__n4870 , _f_permutation__n4869 ,
         _f_permutation__n4868 , _f_permutation__n4867 ,
         _f_permutation__n4866 , _f_permutation__n4865 ,
         _f_permutation__n4864 , _f_permutation__n4863 ,
         _f_permutation__n4862 , _f_permutation__n4861 ,
         _f_permutation__n4860 , _f_permutation__n4859 ,
         _f_permutation__n4858 , _f_permutation__n4857 ,
         _f_permutation__n4856 , _f_permutation__n4855 ,
         _f_permutation__n4854 , _f_permutation__n4853 ,
         _f_permutation__n4852 , _f_permutation__n4851 ,
         _f_permutation__n4850 , _f_permutation__n4849 ,
         _f_permutation__n4848 , _f_permutation__n4847 ,
         _f_permutation__n4846 , _f_permutation__n4845 ,
         _f_permutation__n4844 , _f_permutation__n4843 ,
         _f_permutation__n4842 , _f_permutation__n4841 ,
         _f_permutation__n4840 , _f_permutation__n4839 ,
         _f_permutation__n4838 , _f_permutation__n4837 ,
         _f_permutation__n4836 , _f_permutation__n4835 ,
         _f_permutation__n4834 , _f_permutation__n4833 ,
         _f_permutation__n4832 , _f_permutation__n4831 ,
         _f_permutation__n4830 , _f_permutation__n4829 ,
         _f_permutation__n4828 , _f_permutation__n4827 ,
         _f_permutation__n4826 , _f_permutation__n4825 ,
         _f_permutation__n4824 , _f_permutation__n4823 ,
         _f_permutation__n4822 , _f_permutation__n4821 ,
         _f_permutation__n4820 , _f_permutation__n4819 ,
         _f_permutation__n4818 , _f_permutation__n4817 ,
         _f_permutation__n4816 , _f_permutation__n4815 ,
         _f_permutation__n4814 , _f_permutation__n4813 ,
         _f_permutation__n4812 , _f_permutation__n4811 ,
         _f_permutation__n4810 , _f_permutation__n4809 ,
         _f_permutation__n4808 , _f_permutation__n4807 ,
         _f_permutation__n4806 , _f_permutation__n4805 ,
         _f_permutation__n4804 , _f_permutation__n4803 ,
         _f_permutation__n4802 , _f_permutation__n4801 ,
         _f_permutation__n4800 , _f_permutation__n4799 ,
         _f_permutation__n4798 , _f_permutation__n4797 ,
         _f_permutation__n4796 , _f_permutation__n4795 ,
         _f_permutation__n4794 , _f_permutation__n4793 ,
         _f_permutation__n4792 , _f_permutation__n4791 ,
         _f_permutation__n4790 , _f_permutation__n4789 ,
         _f_permutation__n4788 , _f_permutation__n4787 ,
         _f_permutation__n4786 , _f_permutation__n4785 ,
         _f_permutation__n4784 , _f_permutation__n4783 ,
         _f_permutation__n4782 , _f_permutation__n4781 ,
         _f_permutation__n4780 , _f_permutation__n4779 ,
         _f_permutation__n4778 , _f_permutation__n4777 ,
         _f_permutation__n4776 , _f_permutation__n4775 ,
         _f_permutation__n4774 , _f_permutation__n4773 ,
         _f_permutation__n4772 , _f_permutation__n4771 ,
         _f_permutation__n4770 , _f_permutation__n4769 ,
         _f_permutation__n4768 , _f_permutation__n4767 ,
         _f_permutation__n4766 , _f_permutation__n4765 ,
         _f_permutation__n4764 , _f_permutation__n4763 ,
         _f_permutation__n4762 , _f_permutation__n4761 ,
         _f_permutation__n4760 , _f_permutation__n4759 ,
         _f_permutation__n4758 , _f_permutation__n4757 ,
         _f_permutation__n4756 , _f_permutation__n4755 ,
         _f_permutation__n4754 , _f_permutation__n4753 ,
         _f_permutation__n4752 , _f_permutation__n4751 ,
         _f_permutation__n4750 , _f_permutation__n4749 ,
         _f_permutation__n4748 , _f_permutation__n4747 ,
         _f_permutation__n4746 , _f_permutation__n4745 ,
         _f_permutation__n4744 , _f_permutation__n4743 ,
         _f_permutation__n4742 , _f_permutation__n4741 ,
         _f_permutation__n4740 , _f_permutation__n4739 ,
         _f_permutation__n4738 , _f_permutation__n4737 ,
         _f_permutation__n4736 , _f_permutation__n4735 ,
         _f_permutation__n4734 , _f_permutation__n4733 ,
         _f_permutation__n4732 , _f_permutation__n4731 ,
         _f_permutation__n4730 , _f_permutation__n4729 ,
         _f_permutation__n4728 , _f_permutation__n4727 ,
         _f_permutation__n4726 , _f_permutation__n4725 ,
         _f_permutation__n4724 , _f_permutation__n4723 ,
         _f_permutation__n4722 , _f_permutation__n4721 ,
         _f_permutation__n4720 , _f_permutation__n4719 ,
         _f_permutation__n4718 , _f_permutation__n4717 ,
         _f_permutation__n4716 , _f_permutation__n4715 ,
         _f_permutation__n4714 , _f_permutation__n4713 ,
         _f_permutation__n4712 , _f_permutation__n4711 ,
         _f_permutation__n4710 , _f_permutation__n4709 ,
         _f_permutation__n4708 , _f_permutation__n4707 ,
         _f_permutation__n4706 , _f_permutation__n4705 ,
         _f_permutation__n4704 , _f_permutation__n4703 ,
         _f_permutation__n4702 , _f_permutation__n4701 ,
         _f_permutation__n4700 , _f_permutation__n4699 ,
         _f_permutation__n4698 , _f_permutation__n4697 ,
         _f_permutation__n4696 , _f_permutation__n4695 ,
         _f_permutation__n4694 , _f_permutation__n4693 ,
         _f_permutation__n4692 , _f_permutation__n4691 ,
         _f_permutation__n4690 , _f_permutation__n4689 ,
         _f_permutation__n4688 , _f_permutation__n4687 ,
         _f_permutation__n4686 , _f_permutation__n4685 ,
         _f_permutation__n4684 , _f_permutation__n4683 ,
         _f_permutation__n4682 , _f_permutation__n4681 ,
         _f_permutation__n4680 , _f_permutation__n4679 ,
         _f_permutation__n4678 , _f_permutation__n4677 ,
         _f_permutation__n4676 , _f_permutation__n4675 ,
         _f_permutation__n4674 , _f_permutation__n4673 ,
         _f_permutation__n4672 , _f_permutation__n4671 ,
         _f_permutation__n4670 , _f_permutation__n4669 ,
         _f_permutation__n4668 , _f_permutation__n4667 ,
         _f_permutation__n4666 , _f_permutation__n4665 ,
         _f_permutation__n4664 , _f_permutation__n4663 ,
         _f_permutation__n4662 , _f_permutation__n4661 ,
         _f_permutation__n4660 , _f_permutation__n4659 ,
         _f_permutation__n4658 , _f_permutation__n4657 ,
         _f_permutation__n4656 , _f_permutation__n4655 ,
         _f_permutation__n4654 , _f_permutation__n4653 ,
         _f_permutation__n4652 , _f_permutation__n4651 ,
         _f_permutation__n4650 , _f_permutation__n4649 ,
         _f_permutation__n4648 , _f_permutation__n4647 ,
         _f_permutation__n4646 , _f_permutation__n4645 ,
         _f_permutation__n4644 , _f_permutation__n4643 ,
         _f_permutation__n4642 , _f_permutation__n4641 ,
         _f_permutation__n4640 , _f_permutation__n4639 ,
         _f_permutation__n4638 , _f_permutation__n4637 ,
         _f_permutation__n4636 , _f_permutation__n4635 ,
         _f_permutation__n4634 , _f_permutation__n4633 ,
         _f_permutation__n4632 , _f_permutation__n4631 ,
         _f_permutation__n4630 , _f_permutation__n4629 ,
         _f_permutation__n4628 , _f_permutation__n4627 ,
         _f_permutation__n4626 , _f_permutation__n4625 ,
         _f_permutation__n4624 , _f_permutation__n4623 ,
         _f_permutation__n4622 , _f_permutation__n4621 ,
         _f_permutation__n4620 , _f_permutation__n4619 ,
         _f_permutation__n4618 , _f_permutation__n4617 ,
         _f_permutation__n4616 , _f_permutation__n4615 ,
         _f_permutation__n4614 , _f_permutation__n4613 ,
         _f_permutation__n4612 , _f_permutation__n4611 ,
         _f_permutation__n4610 , _f_permutation__n4609 ,
         _f_permutation__n4608 , _f_permutation__n4607 ,
         _f_permutation__n4606 , _f_permutation__n4605 ,
         _f_permutation__n4604 , _f_permutation__n4603 ,
         _f_permutation__n4602 , _f_permutation__n4601 ,
         _f_permutation__n4600 , _f_permutation__n4599 ,
         _f_permutation__n4598 , _f_permutation__n4597 ,
         _f_permutation__n4596 , _f_permutation__n4595 ,
         _f_permutation__n4594 , _f_permutation__n4593 ,
         _f_permutation__n4592 , _f_permutation__n4591 ,
         _f_permutation__n4590 , _f_permutation__n4589 ,
         _f_permutation__n4588 , _f_permutation__n4587 ,
         _f_permutation__n4586 , _f_permutation__n4585 ,
         _f_permutation__n4584 , _f_permutation__n4583 ,
         _f_permutation__n4582 , _f_permutation__n4581 ,
         _f_permutation__n4580 , _f_permutation__n4579 ,
         _f_permutation__n4578 , _f_permutation__n4577 ,
         _f_permutation__n4576 , _f_permutation__n4575 ,
         _f_permutation__n4574 , _f_permutation__n4573 ,
         _f_permutation__n4572 , _f_permutation__n4571 ,
         _f_permutation__n4570 , _f_permutation__n4569 ,
         _f_permutation__n4568 , _f_permutation__n4567 ,
         _f_permutation__n4566 , _f_permutation__n4565 ,
         _f_permutation__n4564 , _f_permutation__n4563 ,
         _f_permutation__n4562 , _f_permutation__n4561 ,
         _f_permutation__n4560 , _f_permutation__n4559 ,
         _f_permutation__n4558 , _f_permutation__n4557 ,
         _f_permutation__n4556 , _f_permutation__n4555 ,
         _f_permutation__n4554 , _f_permutation__n4553 ,
         _f_permutation__n4552 , _f_permutation__n4551 ,
         _f_permutation__n4550 , _f_permutation__n4549 ,
         _f_permutation__n4548 , _f_permutation__n4547 ,
         _f_permutation__n4546 , _f_permutation__n4545 ,
         _f_permutation__n4544 , _f_permutation__n4543 ,
         _f_permutation__n4542 , _f_permutation__n4541 ,
         _f_permutation__n4540 , _f_permutation__n4539 ,
         _f_permutation__n4538 , _f_permutation__n4537 ,
         _f_permutation__n4536 , _f_permutation__n4535 ,
         _f_permutation__n4534 , _f_permutation__n4533 ,
         _f_permutation__n4532 , _f_permutation__n4531 ,
         _f_permutation__n4530 , _f_permutation__n4529 ,
         _f_permutation__n4528 , _f_permutation__n4527 ,
         _f_permutation__n4526 , _f_permutation__n4525 ,
         _f_permutation__n4524 , _f_permutation__n4523 ,
         _f_permutation__n4522 , _f_permutation__n4521 ,
         _f_permutation__n4520 , _f_permutation__n4519 ,
         _f_permutation__n4518 , _f_permutation__n4517 ,
         _f_permutation__n4516 , _f_permutation__n4515 ,
         _f_permutation__n4514 , _f_permutation__n4513 ,
         _f_permutation__n4512 , _f_permutation__n4511 ,
         _f_permutation__n4510 , _f_permutation__n4509 ,
         _f_permutation__n4508 , _f_permutation__n4507 ,
         _f_permutation__n4506 , _f_permutation__n4505 ,
         _f_permutation__n4504 , _f_permutation__n4503 ,
         _f_permutation__n4502 , _f_permutation__n4501 ,
         _f_permutation__n4500 , _f_permutation__n4499 ,
         _f_permutation__n4498 , _f_permutation__n4497 ,
         _f_permutation__n4496 , _f_permutation__n4495 ,
         _f_permutation__n4494 , _f_permutation__n4493 ,
         _f_permutation__n4492 , _f_permutation__n4491 ,
         _f_permutation__n4490 , _f_permutation__n4489 ,
         _f_permutation__n4488 , _f_permutation__n4487 ,
         _f_permutation__n4486 , _f_permutation__n4485 ,
         _f_permutation__n4484 , _f_permutation__n4483 ,
         _f_permutation__n4482 , _f_permutation__n4481 ,
         _f_permutation__n4480 , _f_permutation__n4479 ,
         _f_permutation__n4478 , _f_permutation__n4477 ,
         _f_permutation__n4476 , _f_permutation__n4475 ,
         _f_permutation__n4474 , _f_permutation__n4473 ,
         _f_permutation__n4472 , _f_permutation__n4471 ,
         _f_permutation__n4470 , _f_permutation__n4469 ,
         _f_permutation__n4468 , _f_permutation__n4467 ,
         _f_permutation__n4466 , _f_permutation__n4465 ,
         _f_permutation__n4464 , _f_permutation__n4463 ,
         _f_permutation__n4462 , _f_permutation__n4461 ,
         _f_permutation__n4460 , _f_permutation__n4459 ,
         _f_permutation__n4458 , _f_permutation__n4457 ,
         _f_permutation__n4456 , _f_permutation__n4455 ,
         _f_permutation__n4454 , _f_permutation__n4453 ,
         _f_permutation__n4452 , _f_permutation__n4451 ,
         _f_permutation__n4450 , _f_permutation__n4449 ,
         _f_permutation__n4448 , _f_permutation__n4447 ,
         _f_permutation__n4446 , _f_permutation__n4445 ,
         _f_permutation__n4444 , _f_permutation__n4443 ,
         _f_permutation__n4442 , _f_permutation__n4441 ,
         _f_permutation__n4440 , _f_permutation__n4439 ,
         _f_permutation__n4438 , _f_permutation__n4437 ,
         _f_permutation__n4436 , _f_permutation__n4435 ,
         _f_permutation__n4434 , _f_permutation__n4433 ,
         _f_permutation__n4432 , _f_permutation__n4431 ,
         _f_permutation__n4430 , _f_permutation__n4429 ,
         _f_permutation__n4428 , _f_permutation__n4427 ,
         _f_permutation__n4426 , _f_permutation__n4425 ,
         _f_permutation__n4424 , _f_permutation__n4423 ,
         _f_permutation__n4422 , _f_permutation__n4421 ,
         _f_permutation__n4420 , _f_permutation__n4419 ,
         _f_permutation__n4418 , _f_permutation__n4417 ,
         _f_permutation__n4416 , _f_permutation__n4415 ,
         _f_permutation__n4414 , _f_permutation__n4413 ,
         _f_permutation__n4412 , _f_permutation__n4411 ,
         _f_permutation__n4410 , _f_permutation__n4409 ,
         _f_permutation__n4408 , _f_permutation__n4407 ,
         _f_permutation__n4406 , _f_permutation__n4405 ,
         _f_permutation__n4404 , _f_permutation__n4403 ,
         _f_permutation__n4402 , _f_permutation__n4401 ,
         _f_permutation__n4400 , _f_permutation__n4399 ,
         _f_permutation__n4398 , _f_permutation__n4397 ,
         _f_permutation__n4396 , _f_permutation__n4395 ,
         _f_permutation__n4394 , _f_permutation__n4393 ,
         _f_permutation__n4392 , _f_permutation__n4391 ,
         _f_permutation__n4390 , _f_permutation__n4389 ,
         _f_permutation__n4388 , _f_permutation__n4387 ,
         _f_permutation__n4386 , _f_permutation__n4385 ,
         _f_permutation__n4384 , _f_permutation__n4383 ,
         _f_permutation__n4382 , _f_permutation__n4381 ,
         _f_permutation__n4380 , _f_permutation__n4379 ,
         _f_permutation__n4378 , _f_permutation__n4377 ,
         _f_permutation__n4376 , _f_permutation__n4375 ,
         _f_permutation__n4374 , _f_permutation__n4373 ,
         _f_permutation__n4372 , _f_permutation__n4371 ,
         _f_permutation__n4370 , _f_permutation__n4369 ,
         _f_permutation__n4368 , _f_permutation__n4367 ,
         _f_permutation__n4366 , _f_permutation__n4365 ,
         _f_permutation__n4364 , _f_permutation__n4363 ,
         _f_permutation__n4362 , _f_permutation__n4361 ,
         _f_permutation__n4360 , _f_permutation__n4359 ,
         _f_permutation__n4358 , _f_permutation__n4357 ,
         _f_permutation__n4356 , _f_permutation__n4355 ,
         _f_permutation__n4354 , _f_permutation__n4353 ,
         _f_permutation__n4352 , _f_permutation__n4351 ,
         _f_permutation__n4350 , _f_permutation__n4349 ,
         _f_permutation__n4348 , _f_permutation__n4347 ,
         _f_permutation__n4346 , _f_permutation__n4345 ,
         _f_permutation__n4344 , _f_permutation__n4343 ,
         _f_permutation__n4342 , _f_permutation__n4341 ,
         _f_permutation__n4340 , _f_permutation__n4339 ,
         _f_permutation__n4338 , _f_permutation__n4337 ,
         _f_permutation__n4336 , _f_permutation__n4335 ,
         _f_permutation__n4334 , _f_permutation__n4333 ,
         _f_permutation__n4332 , _f_permutation__n4331 ,
         _f_permutation__n4330 , _f_permutation__n4329 ,
         _f_permutation__n4328 , _f_permutation__n4327 ,
         _f_permutation__n4326 , _f_permutation__n4325 ,
         _f_permutation__n4324 , _f_permutation__n4323 ,
         _f_permutation__n4322 , _f_permutation__n4321 ,
         _f_permutation__n4320 , _f_permutation__n4319 ,
         _f_permutation__n4318 , _f_permutation__n4317 ,
         _f_permutation__n4316 , _f_permutation__n4315 ,
         _f_permutation__n4314 , _f_permutation__n4313 ,
         _f_permutation__n4312 , _f_permutation__n4311 ,
         _f_permutation__n4310 , _f_permutation__n4309 ,
         _f_permutation__n4308 , _f_permutation__n4307 ,
         _f_permutation__n4306 , _f_permutation__n4305 ,
         _f_permutation__n4304 , _f_permutation__n4303 ,
         _f_permutation__n4302 , _f_permutation__n4301 ,
         _f_permutation__n4300 , _f_permutation__n4299 ,
         _f_permutation__n4298 , _f_permutation__n4297 ,
         _f_permutation__n4296 , _f_permutation__n4295 ,
         _f_permutation__n4294 , _f_permutation__n4293 ,
         _f_permutation__n4292 , _f_permutation__n4291 ,
         _f_permutation__n4290 , _f_permutation__n4289 ,
         _f_permutation__n4288 , _f_permutation__n4287 ,
         _f_permutation__n4286 , _f_permutation__n4285 ,
         _f_permutation__n4284 , _f_permutation__n4283 ,
         _f_permutation__n4282 , _f_permutation__n4281 ,
         _f_permutation__n4280 , _f_permutation__n4279 ,
         _f_permutation__n4278 , _f_permutation__n4277 ,
         _f_permutation__n4276 , _f_permutation__n4275 ,
         _f_permutation__n4274 , _f_permutation__n4273 ,
         _f_permutation__n4272 , _f_permutation__n4271 ,
         _f_permutation__n4270 , _f_permutation__n4269 ,
         _f_permutation__n4268 , _f_permutation__n4267 ,
         _f_permutation__n4266 , _f_permutation__n4265 ,
         _f_permutation__n4264 , _f_permutation__n4263 ,
         _f_permutation__n4262 , _f_permutation__n4261 ,
         _f_permutation__n4260 , _f_permutation__n4259 ,
         _f_permutation__n4258 , _f_permutation__n4257 ,
         _f_permutation__n4256 , _f_permutation__n4255 ,
         _f_permutation__n4254 , _f_permutation__n4253 ,
         _f_permutation__n4252 , _f_permutation__n4251 ,
         _f_permutation__n4250 , _f_permutation__n4249 ,
         _f_permutation__n4248 , _f_permutation__n4247 ,
         _f_permutation__n4246 , _f_permutation__n4245 ,
         _f_permutation__n4244 , _f_permutation__n4243 ,
         _f_permutation__n4242 , _f_permutation__n4241 ,
         _f_permutation__n4240 , _f_permutation__n4239 ,
         _f_permutation__n4238 , _f_permutation__n4237 ,
         _f_permutation__n4236 , _f_permutation__n4235 ,
         _f_permutation__n4234 , _f_permutation__n4233 ,
         _f_permutation__n4232 , _f_permutation__n4231 ,
         _f_permutation__n4230 , _f_permutation__n4229 ,
         _f_permutation__n4228 , _f_permutation__n4227 ,
         _f_permutation__n4226 , _f_permutation__n4225 ,
         _f_permutation__n4224 , _f_permutation__n4223 ,
         _f_permutation__n4222 , _f_permutation__n4221 ,
         _f_permutation__n4220 , _f_permutation__n4219 ,
         _f_permutation__n4218 , _f_permutation__n4217 ,
         _f_permutation__n4216 , _f_permutation__n4215 ,
         _f_permutation__n4214 , _f_permutation__n4213 ,
         _f_permutation__n4212 , _f_permutation__n4211 ,
         _f_permutation__n4210 , _f_permutation__n4209 ,
         _f_permutation__n4208 , _f_permutation__n4207 ,
         _f_permutation__n4206 , _f_permutation__n4205 ,
         _f_permutation__n4204 , _f_permutation__n4203 ,
         _f_permutation__n4202 , _f_permutation__n4201 ,
         _f_permutation__n4200 , _f_permutation__n4199 ,
         _f_permutation__n4198 , _f_permutation__n4197 ,
         _f_permutation__n4196 , _f_permutation__n4195 ,
         _f_permutation__n4194 , _f_permutation__n4193 ,
         _f_permutation__n4192 , _f_permutation__n4191 ,
         _f_permutation__n4190 , _f_permutation__n4189 ,
         _f_permutation__n4188 , _f_permutation__n4187 ,
         _f_permutation__n4186 , _f_permutation__n4185 ,
         _f_permutation__n4184 , _f_permutation__n4183 ,
         _f_permutation__n4182 , _f_permutation__n4181 ,
         _f_permutation__n4180 , _f_permutation__n4179 ,
         _f_permutation__n4178 , _f_permutation__n4177 ,
         _f_permutation__n4176 , _f_permutation__n4175 ,
         _f_permutation__n4174 , _f_permutation__n4173 ,
         _f_permutation__n4172 , _f_permutation__n4171 ,
         _f_permutation__n4170 , _f_permutation__n4169 ,
         _f_permutation__n4168 , _f_permutation__n4167 ,
         _f_permutation__n4166 , _f_permutation__n4165 ,
         _f_permutation__n4164 , _f_permutation__n4163 ,
         _f_permutation__n4162 , _f_permutation__n4161 ,
         _f_permutation__n4160 , _f_permutation__n4159 ,
         _f_permutation__n4158 , _f_permutation__n4157 ,
         _f_permutation__n4156 , _f_permutation__n4155 ,
         _f_permutation__n4154 , _f_permutation__n4153 ,
         _f_permutation__n4152 , _f_permutation__n4151 ,
         _f_permutation__n4150 , _f_permutation__n4149 ,
         _f_permutation__n4148 , _f_permutation__n4147 ,
         _f_permutation__n4146 , _f_permutation__n4145 ,
         _f_permutation__n4144 , _f_permutation__n4143 ,
         _f_permutation__n4142 , _f_permutation__n4141 ,
         _f_permutation__n4140 , _f_permutation__n4139 ,
         _f_permutation__n4138 , _f_permutation__n4137 ,
         _f_permutation__n4136 , _f_permutation__n4135 ,
         _f_permutation__n4134 , _f_permutation__n4133 ,
         _f_permutation__n4132 , _f_permutation__n4131 ,
         _f_permutation__n4130 , _f_permutation__n4129 ,
         _f_permutation__n4128 , _f_permutation__n4127 ,
         _f_permutation__n4126 , _f_permutation__n4125 ,
         _f_permutation__n4124 , _f_permutation__n4123 ,
         _f_permutation__n4122 , _f_permutation__n4121 ,
         _f_permutation__n4120 , _f_permutation__n4119 ,
         _f_permutation__n4118 , _f_permutation__n4117 ,
         _f_permutation__n4116 , _f_permutation__n4115 ,
         _f_permutation__n4114 , _f_permutation__n4113 ,
         _f_permutation__n4112 , _f_permutation__n4111 ,
         _f_permutation__n4110 , _f_permutation__n4109 ,
         _f_permutation__n4108 , _f_permutation__n4107 ,
         _f_permutation__n4106 , _f_permutation__n4105 ,
         _f_permutation__n4104 , _f_permutation__n4103 ,
         _f_permutation__n4102 , _f_permutation__n4101 ,
         _f_permutation__n4100 , _f_permutation__n4099 ,
         _f_permutation__n4098 , _f_permutation__n4097 ,
         _f_permutation__n4096 , _f_permutation__n4095 ,
         _f_permutation__n4094 , _f_permutation__n4093 ,
         _f_permutation__n4092 , _f_permutation__n4091 ,
         _f_permutation__n4090 , _f_permutation__n4089 ,
         _f_permutation__n4088 , _f_permutation__n4087 ,
         _f_permutation__n4086 , _f_permutation__n4085 ,
         _f_permutation__n4084 , _f_permutation__n4083 ,
         _f_permutation__n4082 , _f_permutation__n4081 ,
         _f_permutation__n4080 , _f_permutation__n4079 ,
         _f_permutation__n4078 , _f_permutation__n4077 ,
         _f_permutation__n4076 , _f_permutation__n4075 ,
         _f_permutation__n4074 , _f_permutation__n4073 ,
         _f_permutation__n4072 , _f_permutation__n4071 ,
         _f_permutation__n4070 , _f_permutation__n4069 ,
         _f_permutation__n4068 , _f_permutation__n4067 ,
         _f_permutation__n4066 , _f_permutation__n4065 ,
         _f_permutation__n4064 , _f_permutation__n4063 ,
         _f_permutation__n4062 , _f_permutation__n4061 ,
         _f_permutation__n4060 , _f_permutation__n4059 ,
         _f_permutation__n4058 , _f_permutation__n4057 ,
         _f_permutation__n4056 , _f_permutation__n4055 ,
         _f_permutation__n4054 , _f_permutation__n4053 ,
         _f_permutation__n4052 , _f_permutation__n4051 ,
         _f_permutation__n4050 , _f_permutation__n4049 ,
         _f_permutation__n4048 , _f_permutation__n4047 ,
         _f_permutation__n4046 , _f_permutation__n4045 ,
         _f_permutation__n4044 , _f_permutation__n4043 ,
         _f_permutation__n4042 , _f_permutation__n4041 ,
         _f_permutation__n4040 , _f_permutation__n4039 ,
         _f_permutation__n4038 , _f_permutation__n4037 ,
         _f_permutation__n4036 , _f_permutation__n4035 ,
         _f_permutation__n4034 , _f_permutation__n4033 ,
         _f_permutation__n4032 , _f_permutation__n4031 ,
         _f_permutation__n4030 , _f_permutation__n4029 ,
         _f_permutation__n4028 , _f_permutation__n4027 ,
         _f_permutation__n4026 , _f_permutation__n4025 ,
         _f_permutation__n4024 , _f_permutation__n4023 ,
         _f_permutation__n4022 , _f_permutation__n4021 ,
         _f_permutation__n4020 , _f_permutation__n4019 ,
         _f_permutation__n4018 , _f_permutation__n4017 ,
         _f_permutation__n4016 , _f_permutation__n4015 ,
         _f_permutation__n4014 , _f_permutation__n4013 ,
         _f_permutation__n4012 , _f_permutation__n4011 ,
         _f_permutation__n4010 , _f_permutation__n4009 ,
         _f_permutation__n4008 , _f_permutation__n4007 ,
         _f_permutation__n4006 , _f_permutation__n4005 ,
         _f_permutation__n4004 , _f_permutation__n4003 ,
         _f_permutation__n4002 , _f_permutation__n4001 ,
         _f_permutation__n4000 , _f_permutation__n3999 ,
         _f_permutation__n3998 , _f_permutation__n3997 ,
         _f_permutation__n3996 , _f_permutation__n3995 ,
         _f_permutation__n3994 , _f_permutation__n3993 ,
         _f_permutation__n3992 , _f_permutation__n3991 ,
         _f_permutation__n3990 , _f_permutation__n3989 ,
         _f_permutation__n3988 , _f_permutation__n3987 ,
         _f_permutation__n3986 , _f_permutation__n3985 ,
         _f_permutation__n3984 , _f_permutation__n3983 ,
         _f_permutation__n3982 , _f_permutation__n3981 ,
         _f_permutation__n3980 , _f_permutation__n3979 ,
         _f_permutation__n3978 , _f_permutation__n3977 ,
         _f_permutation__n3976 , _f_permutation__n3975 ,
         _f_permutation__n3974 , _f_permutation__n3973 ,
         _f_permutation__n3972 , _f_permutation__n3971 ,
         _f_permutation__n3970 , _f_permutation__n3969 ,
         _f_permutation__n3968 , _f_permutation__n3967 ,
         _f_permutation__n3966 , _f_permutation__n3965 ,
         _f_permutation__n3964 , _f_permutation__n3963 ,
         _f_permutation__n3962 , _f_permutation__n3961 ,
         _f_permutation__n3960 , _f_permutation__n3959 ,
         _f_permutation__n3958 , _f_permutation__n3957 ,
         _f_permutation__n3956 , _f_permutation__n3955 ,
         _f_permutation__n3954 , _f_permutation__n3953 ,
         _f_permutation__n3952 , _f_permutation__n3951 ,
         _f_permutation__n3950 , _f_permutation__n3949 ,
         _f_permutation__n3948 , _f_permutation__n3947 ,
         _f_permutation__n3946 , _f_permutation__n3945 ,
         _f_permutation__n3944 , _f_permutation__n3943 ,
         _f_permutation__n3942 , _f_permutation__n3941 ,
         _f_permutation__n3940 , _f_permutation__n3939 ,
         _f_permutation__n3938 , _f_permutation__n3937 ,
         _f_permutation__n3936 , _f_permutation__n3935 ,
         _f_permutation__n3934 , _f_permutation__n3933 ,
         _f_permutation__n3932 , _f_permutation__n3931 ,
         _f_permutation__n3930 , _f_permutation__n3929 ,
         _f_permutation__n3928 , _f_permutation__n3927 ,
         _f_permutation__n3926 , _f_permutation__n3925 ,
         _f_permutation__n3924 , _f_permutation__n3923 ,
         _f_permutation__n3922 , _f_permutation__n3921 ,
         _f_permutation__n3920 , _f_permutation__n3919 ,
         _f_permutation__n3918 , _f_permutation__n3917 ,
         _f_permutation__n3916 , _f_permutation__n3915 ,
         _f_permutation__n3914 , _f_permutation__n3913 ,
         _f_permutation__n3912 , _f_permutation__n3911 ,
         _f_permutation__n3910 , _f_permutation__n3909 ,
         _f_permutation__n3908 , _f_permutation__n3907 ,
         _f_permutation__n3906 , _f_permutation__n3905 ,
         _f_permutation__n3904 , _f_permutation__n3903 ,
         _f_permutation__n3902 , _f_permutation__n3901 ,
         _f_permutation__n3900 , _f_permutation__n3899 ,
         _f_permutation__n3898 , _f_permutation__n3897 ,
         _f_permutation__n3896 , _f_permutation__n3895 ,
         _f_permutation__n3894 , _f_permutation__n3893 ,
         _f_permutation__n3892 , _f_permutation__n3891 ,
         _f_permutation__n3890 , _f_permutation__n3889 ,
         _f_permutation__n3888 , _f_permutation__n3887 ,
         _f_permutation__n3886 , _f_permutation__n3885 ,
         _f_permutation__n3884 , _f_permutation__n3883 ,
         _f_permutation__n3882 , _f_permutation__n3881 ,
         _f_permutation__n3880 , _f_permutation__n3879 ,
         _f_permutation__n3878 , _f_permutation__n3877 ,
         _f_permutation__n3876 , _f_permutation__n3875 ,
         _f_permutation__n3874 , _f_permutation__n3873 ,
         _f_permutation__n3872 , _f_permutation__n3871 ,
         _f_permutation__n3870 , _f_permutation__n3869 ,
         _f_permutation__n3868 , _f_permutation__n3867 ,
         _f_permutation__n3866 , _f_permutation__n3865 ,
         _f_permutation__n3864 , _f_permutation__n3863 ,
         _f_permutation__n3862 , _f_permutation__n3861 ,
         _f_permutation__n3860 , _f_permutation__n3859 ,
         _f_permutation__n3858 , _f_permutation__n3857 ,
         _f_permutation__n3856 , _f_permutation__n3855 ,
         _f_permutation__n3854 , _f_permutation__n3853 ,
         _f_permutation__n3852 , _f_permutation__n3851 ,
         _f_permutation__n3850 , _f_permutation__n3849 ,
         _f_permutation__n3848 , _f_permutation__n3847 ,
         _f_permutation__n3846 , _f_permutation__n3845 ,
         _f_permutation__n3844 , _f_permutation__n3843 ,
         _f_permutation__n3842 , _f_permutation__n3841 ,
         _f_permutation__n3840 , _f_permutation__n3839 ,
         _f_permutation__n3838 , _f_permutation__n3837 ,
         _f_permutation__n3836 , _f_permutation__n3835 ,
         _f_permutation__n3834 , _f_permutation__n3833 ,
         _f_permutation__n3832 , _f_permutation__n3831 ,
         _f_permutation__n3830 , _f_permutation__n3829 ,
         _f_permutation__n3828 , _f_permutation__n3827 ,
         _f_permutation__n3826 , _f_permutation__n3825 ,
         _f_permutation__n3824 , _f_permutation__n3823 ,
         _f_permutation__n3822 , _f_permutation__n3821 ,
         _f_permutation__n3820 , _f_permutation__n3819 ,
         _f_permutation__n3818 , _f_permutation__n3817 ,
         _f_permutation__n3816 , _f_permutation__n3815 ,
         _f_permutation__n3814 , _f_permutation__n3813 ,
         _f_permutation__n3812 , _f_permutation__n3811 ,
         _f_permutation__n3810 , _f_permutation__n3809 ,
         _f_permutation__n3808 , _f_permutation__n3807 ,
         _f_permutation__n3806 , _f_permutation__n3805 ,
         _f_permutation__n3804 , _f_permutation__n3803 ,
         _f_permutation__n3802 , _f_permutation__n3801 ,
         _f_permutation__n3800 , _f_permutation__n3799 ,
         _f_permutation__n3798 , _f_permutation__n3797 ,
         _f_permutation__n3796 , _f_permutation__n3795 ,
         _f_permutation__n3794 , _f_permutation__n3793 ,
         _f_permutation__n3792 , _f_permutation__n3791 ,
         _f_permutation__n3790 , _f_permutation__n3789 ,
         _f_permutation__n3788 , _f_permutation__N29 , _f_permutation__N27 ,
         _f_permutation__N26 , _f_permutation__N25 , _f_permutation__N24 ,
         _f_permutation__N23 , _f_permutation__N22 , _f_permutation__N21 ,
         _f_permutation__N20 , _f_permutation__N19 , _f_permutation__N18 ,
         _f_permutation__N17 , _f_permutation__N16 , _f_permutation__N15 ,
         _f_permutation__N14 , _f_permutation__N13 , _f_permutation__N12 ,
         _f_permutation__N11 , _f_permutation__N10 , _f_permutation__N9 ,
         _f_permutation__N8 , _f_permutation__N7 , _f_permutation__N6 ,
         _f_permutation__i[0] , _f_permutation__i[1] , _f_permutation__i[2] ,
         _f_permutation__i[3] , _f_permutation__i[4] , _f_permutation__i[5] ,
         _f_permutation__i[6] , _f_permutation__i[7] , _f_permutation__i[8] ,
         _f_permutation__i[9] , _f_permutation__i[10] , _f_permutation__i[11] ,
         _f_permutation__i[12] , _f_permutation__i[13] ,
         _f_permutation__i[14] , _f_permutation__i[15] ,
         _f_permutation__i[16] , _f_permutation__i[17] ,
         _f_permutation__i[18] , _f_permutation__i[19] ,
         _f_permutation__i[20] , _f_permutation__i[21] ,
         _f_permutation__i[22] , _f_permutation__out_ready ,
         _f_permutation__rconst__rc[62] , _f_permutation__rconst__rc[61] ,
         _f_permutation__rconst__rc[60] , _f_permutation__rconst__rc[59] ,
         _f_permutation__rconst__rc[58] , _f_permutation__rconst__rc[57] ,
         _f_permutation__rconst__rc[56] , _f_permutation__rconst__rc[55] ,
         _f_permutation__rconst__rc[54] , _f_permutation__rconst__rc[53] ,
         _f_permutation__rconst__rc[52] , _f_permutation__rconst__rc[51] ,
         _f_permutation__rconst__rc[50] , _f_permutation__rconst__rc[49] ,
         _f_permutation__rconst__rc[48] , _f_permutation__rconst__rc[47] ,
         _f_permutation__rconst__rc[46] , _f_permutation__rconst__rc[45] ,
         _f_permutation__rconst__rc[44] , _f_permutation__rconst__rc[43] ,
         _f_permutation__rconst__rc[42] , _f_permutation__rconst__rc[41] ,
         _f_permutation__rconst__rc[40] , _f_permutation__rconst__rc[39] ,
         _f_permutation__rconst__rc[38] , _f_permutation__rconst__rc[37] ,
         _f_permutation__rconst__rc[36] , _f_permutation__rconst__rc[35] ,
         _f_permutation__rconst__rc[34] , _f_permutation__rconst__rc[33] ,
         _f_permutation__rconst__rc[32] , _f_permutation__rconst__rc[30] ,
         _f_permutation__rconst__rc[29] , _f_permutation__rconst__rc[28] ,
         _f_permutation__rconst__rc[27] , _f_permutation__rconst__rc[26] ,
         _f_permutation__rconst__rc[25] , _f_permutation__rconst__rc[24] ,
         _f_permutation__rconst__rc[23] , _f_permutation__rconst__rc[22] ,
         _f_permutation__rconst__rc[21] , _f_permutation__rconst__rc[20] ,
         _f_permutation__rconst__rc[19] , _f_permutation__rconst__rc[18] ,
         _f_permutation__rconst__rc[17] , _f_permutation__rconst__rc[16] ,
         _f_permutation__rconst__rc[14] , _f_permutation__rconst__rc[13] ,
         _f_permutation__rconst__rc[12] , _f_permutation__rconst__rc[11] ,
         _f_permutation__rconst__rc[10] , _f_permutation__rconst__rc[9] ,
         _f_permutation__rconst__rc[8] , _f_permutation__rconst__rc[6] ,
         _f_permutation__rconst__rc[5] , _f_permutation__rconst__rc[4] ,
         _f_permutation__rconst__rc[2] , _f_permutation__rconst__n23 ,
         _f_permutation__rconst__n22 , _f_permutation__rconst__n21 ,
         _f_permutation__rconst__n20 , _f_permutation__rconst__n19 ,
         _f_permutation__rconst__n18 , _f_permutation__rconst__n17 ,
         _f_permutation__rconst__n16 , _f_permutation__rconst__n15 ,
         _f_permutation__rconst__n14 , _f_permutation__rconst__n13 ,
         _f_permutation__rconst__n12 , _f_permutation__rconst__n11 ,
         _f_permutation__rconst__n10 , _f_permutation__rconst__n9 ,
         _f_permutation__rconst__n8 , _f_permutation__rconst__n7 ,
         _f_permutation__rconst__n6 , _f_permutation__rconst__n5 ,
         _f_permutation__rconst__n4 , _f_permutation__rconst__n3 ,
         _f_permutation__rconst__n2 , _f_permutation__rconst__n1 ,
         _f_permutation__round__n960 , _f_permutation__round__n959 ,
         _f_permutation__round__n958 , _f_permutation__round__n957 ,
         _f_permutation__round__n956 , _f_permutation__round__n955 ,
         _f_permutation__round__n954 , _f_permutation__round__n953 ,
         _f_permutation__round__n952 , _f_permutation__round__n951 ,
         _f_permutation__round__n950 , _f_permutation__round__n949 ,
         _f_permutation__round__n948 , _f_permutation__round__n947 ,
         _f_permutation__round__n946 , _f_permutation__round__n945 ,
         _f_permutation__round__n944 , _f_permutation__round__n943 ,
         _f_permutation__round__n942 , _f_permutation__round__n941 ,
         _f_permutation__round__n940 , _f_permutation__round__n939 ,
         _f_permutation__round__n938 , _f_permutation__round__n937 ,
         _f_permutation__round__n936 , _f_permutation__round__n935 ,
         _f_permutation__round__n934 , _f_permutation__round__n933 ,
         _f_permutation__round__n932 , _f_permutation__round__n931 ,
         _f_permutation__round__n930 , _f_permutation__round__n929 ,
         _f_permutation__round__n928 , _f_permutation__round__n927 ,
         _f_permutation__round__n926 , _f_permutation__round__n925 ,
         _f_permutation__round__n924 , _f_permutation__round__n923 ,
         _f_permutation__round__n922 , _f_permutation__round__n921 ,
         _f_permutation__round__n920 , _f_permutation__round__n919 ,
         _f_permutation__round__n918 , _f_permutation__round__n917 ,
         _f_permutation__round__n916 , _f_permutation__round__n915 ,
         _f_permutation__round__n914 , _f_permutation__round__n913 ,
         _f_permutation__round__n912 , _f_permutation__round__n911 ,
         _f_permutation__round__n910 , _f_permutation__round__n909 ,
         _f_permutation__round__n908 , _f_permutation__round__n907 ,
         _f_permutation__round__n906 , _f_permutation__round__n905 ,
         _f_permutation__round__n904 , _f_permutation__round__n903 ,
         _f_permutation__round__n902 , _f_permutation__round__n901 ,
         _f_permutation__round__n900 , _f_permutation__round__n899 ,
         _f_permutation__round__n898 , _f_permutation__round__n897 ,
         _f_permutation__round__n896 , _f_permutation__round__n895 ,
         _f_permutation__round__n894 , _f_permutation__round__n893 ,
         _f_permutation__round__n892 , _f_permutation__round__n891 ,
         _f_permutation__round__n890 , _f_permutation__round__n889 ,
         _f_permutation__round__n888 , _f_permutation__round__n887 ,
         _f_permutation__round__n886 , _f_permutation__round__n885 ,
         _f_permutation__round__n884 , _f_permutation__round__n883 ,
         _f_permutation__round__n882 , _f_permutation__round__n881 ,
         _f_permutation__round__n880 , _f_permutation__round__n879 ,
         _f_permutation__round__n878 , _f_permutation__round__n877 ,
         _f_permutation__round__n876 , _f_permutation__round__n875 ,
         _f_permutation__round__n874 , _f_permutation__round__n873 ,
         _f_permutation__round__n872 , _f_permutation__round__n871 ,
         _f_permutation__round__n870 , _f_permutation__round__n869 ,
         _f_permutation__round__n868 , _f_permutation__round__n867 ,
         _f_permutation__round__n866 , _f_permutation__round__n865 ,
         _f_permutation__round__n864 , _f_permutation__round__n863 ,
         _f_permutation__round__n862 , _f_permutation__round__n861 ,
         _f_permutation__round__n860 , _f_permutation__round__n859 ,
         _f_permutation__round__n858 , _f_permutation__round__n857 ,
         _f_permutation__round__n856 , _f_permutation__round__n855 ,
         _f_permutation__round__n854 , _f_permutation__round__n853 ,
         _f_permutation__round__n852 , _f_permutation__round__n851 ,
         _f_permutation__round__n850 , _f_permutation__round__n849 ,
         _f_permutation__round__n848 , _f_permutation__round__n847 ,
         _f_permutation__round__n846 , _f_permutation__round__n845 ,
         _f_permutation__round__n844 , _f_permutation__round__n843 ,
         _f_permutation__round__n842 , _f_permutation__round__n841 ,
         _f_permutation__round__n840 , _f_permutation__round__n839 ,
         _f_permutation__round__n838 , _f_permutation__round__n837 ,
         _f_permutation__round__n836 , _f_permutation__round__n835 ,
         _f_permutation__round__n834 , _f_permutation__round__n833 ,
         _f_permutation__round__n832 , _f_permutation__round__n831 ,
         _f_permutation__round__n830 , _f_permutation__round__n829 ,
         _f_permutation__round__n828 , _f_permutation__round__n827 ,
         _f_permutation__round__n826 , _f_permutation__round__n825 ,
         _f_permutation__round__n824 , _f_permutation__round__n823 ,
         _f_permutation__round__n822 , _f_permutation__round__n821 ,
         _f_permutation__round__n820 , _f_permutation__round__n819 ,
         _f_permutation__round__n818 , _f_permutation__round__n817 ,
         _f_permutation__round__n816 , _f_permutation__round__n815 ,
         _f_permutation__round__n814 , _f_permutation__round__n813 ,
         _f_permutation__round__n812 , _f_permutation__round__n811 ,
         _f_permutation__round__n810 , _f_permutation__round__n809 ,
         _f_permutation__round__n808 , _f_permutation__round__n807 ,
         _f_permutation__round__n806 , _f_permutation__round__n805 ,
         _f_permutation__round__n804 , _f_permutation__round__n803 ,
         _f_permutation__round__n802 , _f_permutation__round__n801 ,
         _f_permutation__round__n800 , _f_permutation__round__n799 ,
         _f_permutation__round__n798 , _f_permutation__round__n797 ,
         _f_permutation__round__n796 , _f_permutation__round__n795 ,
         _f_permutation__round__n794 , _f_permutation__round__n793 ,
         _f_permutation__round__n792 , _f_permutation__round__n791 ,
         _f_permutation__round__n790 , _f_permutation__round__n789 ,
         _f_permutation__round__n788 , _f_permutation__round__n787 ,
         _f_permutation__round__n786 , _f_permutation__round__n785 ,
         _f_permutation__round__n784 , _f_permutation__round__n783 ,
         _f_permutation__round__n782 , _f_permutation__round__n781 ,
         _f_permutation__round__n780 , _f_permutation__round__n779 ,
         _f_permutation__round__n778 , _f_permutation__round__n777 ,
         _f_permutation__round__n776 , _f_permutation__round__n775 ,
         _f_permutation__round__n774 , _f_permutation__round__n773 ,
         _f_permutation__round__n772 , _f_permutation__round__n771 ,
         _f_permutation__round__n770 , _f_permutation__round__n769 ,
         _f_permutation__round__n768 , _f_permutation__round__n767 ,
         _f_permutation__round__n766 , _f_permutation__round__n765 ,
         _f_permutation__round__n764 , _f_permutation__round__n763 ,
         _f_permutation__round__n762 , _f_permutation__round__n761 ,
         _f_permutation__round__n760 , _f_permutation__round__n759 ,
         _f_permutation__round__n758 , _f_permutation__round__n757 ,
         _f_permutation__round__n756 , _f_permutation__round__n755 ,
         _f_permutation__round__n754 , _f_permutation__round__n753 ,
         _f_permutation__round__n752 , _f_permutation__round__n751 ,
         _f_permutation__round__n750 , _f_permutation__round__n749 ,
         _f_permutation__round__n748 , _f_permutation__round__n747 ,
         _f_permutation__round__n746 , _f_permutation__round__n745 ,
         _f_permutation__round__n744 , _f_permutation__round__n743 ,
         _f_permutation__round__n742 , _f_permutation__round__n741 ,
         _f_permutation__round__n740 , _f_permutation__round__n739 ,
         _f_permutation__round__n738 , _f_permutation__round__n737 ,
         _f_permutation__round__n736 , _f_permutation__round__n735 ,
         _f_permutation__round__n734 , _f_permutation__round__n733 ,
         _f_permutation__round__n732 , _f_permutation__round__n731 ,
         _f_permutation__round__n730 , _f_permutation__round__n729 ,
         _f_permutation__round__n728 , _f_permutation__round__n727 ,
         _f_permutation__round__n726 , _f_permutation__round__n725 ,
         _f_permutation__round__n724 , _f_permutation__round__n723 ,
         _f_permutation__round__n722 , _f_permutation__round__n721 ,
         _f_permutation__round__n720 , _f_permutation__round__n719 ,
         _f_permutation__round__n718 , _f_permutation__round__n717 ,
         _f_permutation__round__n716 , _f_permutation__round__n715 ,
         _f_permutation__round__n714 , _f_permutation__round__n713 ,
         _f_permutation__round__n712 , _f_permutation__round__n711 ,
         _f_permutation__round__n710 , _f_permutation__round__n709 ,
         _f_permutation__round__n708 , _f_permutation__round__n707 ,
         _f_permutation__round__n706 , _f_permutation__round__n705 ,
         _f_permutation__round__n704 , _f_permutation__round__n703 ,
         _f_permutation__round__n702 , _f_permutation__round__n701 ,
         _f_permutation__round__n700 , _f_permutation__round__n699 ,
         _f_permutation__round__n698 , _f_permutation__round__n697 ,
         _f_permutation__round__n696 , _f_permutation__round__n695 ,
         _f_permutation__round__n694 , _f_permutation__round__n693 ,
         _f_permutation__round__n692 , _f_permutation__round__n691 ,
         _f_permutation__round__n690 , _f_permutation__round__n689 ,
         _f_permutation__round__n688 , _f_permutation__round__n687 ,
         _f_permutation__round__n686 , _f_permutation__round__n685 ,
         _f_permutation__round__n684 , _f_permutation__round__n683 ,
         _f_permutation__round__n682 , _f_permutation__round__n681 ,
         _f_permutation__round__n680 , _f_permutation__round__n679 ,
         _f_permutation__round__n678 , _f_permutation__round__n677 ,
         _f_permutation__round__n676 , _f_permutation__round__n675 ,
         _f_permutation__round__n674 , _f_permutation__round__n673 ,
         _f_permutation__round__n672 , _f_permutation__round__n671 ,
         _f_permutation__round__n670 , _f_permutation__round__n669 ,
         _f_permutation__round__n668 , _f_permutation__round__n667 ,
         _f_permutation__round__n666 , _f_permutation__round__n665 ,
         _f_permutation__round__n664 , _f_permutation__round__n663 ,
         _f_permutation__round__n662 , _f_permutation__round__n661 ,
         _f_permutation__round__n660 , _f_permutation__round__n659 ,
         _f_permutation__round__n658 , _f_permutation__round__n657 ,
         _f_permutation__round__n656 , _f_permutation__round__n655 ,
         _f_permutation__round__n654 , _f_permutation__round__n653 ,
         _f_permutation__round__n652 , _f_permutation__round__n651 ,
         _f_permutation__round__n650 , _f_permutation__round__n649 ,
         _f_permutation__round__n648 , _f_permutation__round__n647 ,
         _f_permutation__round__n646 , _f_permutation__round__n645 ,
         _f_permutation__round__n644 , _f_permutation__round__n643 ,
         _f_permutation__round__n642 , _f_permutation__round__n641 ,
         _f_permutation__round__n640 , _f_permutation__round__n639 ,
         _f_permutation__round__n638 , _f_permutation__round__n637 ,
         _f_permutation__round__n636 , _f_permutation__round__n635 ,
         _f_permutation__round__n634 , _f_permutation__round__n633 ,
         _f_permutation__round__n632 , _f_permutation__round__n631 ,
         _f_permutation__round__n630 , _f_permutation__round__n629 ,
         _f_permutation__round__n628 , _f_permutation__round__n627 ,
         _f_permutation__round__n626 , _f_permutation__round__n625 ,
         _f_permutation__round__n624 , _f_permutation__round__n623 ,
         _f_permutation__round__n622 , _f_permutation__round__n621 ,
         _f_permutation__round__n620 , _f_permutation__round__n619 ,
         _f_permutation__round__n618 , _f_permutation__round__n617 ,
         _f_permutation__round__n616 , _f_permutation__round__n615 ,
         _f_permutation__round__n614 , _f_permutation__round__n613 ,
         _f_permutation__round__n612 , _f_permutation__round__n611 ,
         _f_permutation__round__n610 , _f_permutation__round__n609 ,
         _f_permutation__round__n608 , _f_permutation__round__n607 ,
         _f_permutation__round__n606 , _f_permutation__round__n605 ,
         _f_permutation__round__n604 , _f_permutation__round__n603 ,
         _f_permutation__round__n602 , _f_permutation__round__n601 ,
         _f_permutation__round__n600 , _f_permutation__round__n599 ,
         _f_permutation__round__n598 , _f_permutation__round__n597 ,
         _f_permutation__round__n596 , _f_permutation__round__n595 ,
         _f_permutation__round__n594 , _f_permutation__round__n593 ,
         _f_permutation__round__n592 , _f_permutation__round__n591 ,
         _f_permutation__round__n590 , _f_permutation__round__n589 ,
         _f_permutation__round__n588 , _f_permutation__round__n587 ,
         _f_permutation__round__n586 , _f_permutation__round__n585 ,
         _f_permutation__round__n584 , _f_permutation__round__n583 ,
         _f_permutation__round__n582 , _f_permutation__round__n581 ,
         _f_permutation__round__n580 , _f_permutation__round__n579 ,
         _f_permutation__round__n578 , _f_permutation__round__n577 ,
         _f_permutation__round__n576 , _f_permutation__round__n575 ,
         _f_permutation__round__n574 , _f_permutation__round__n573 ,
         _f_permutation__round__n572 , _f_permutation__round__n571 ,
         _f_permutation__round__n570 , _f_permutation__round__n569 ,
         _f_permutation__round__n568 , _f_permutation__round__n567 ,
         _f_permutation__round__n566 , _f_permutation__round__n565 ,
         _f_permutation__round__n564 , _f_permutation__round__n563 ,
         _f_permutation__round__n562 , _f_permutation__round__n561 ,
         _f_permutation__round__n560 , _f_permutation__round__n559 ,
         _f_permutation__round__n558 , _f_permutation__round__n557 ,
         _f_permutation__round__n556 , _f_permutation__round__n555 ,
         _f_permutation__round__n554 , _f_permutation__round__n553 ,
         _f_permutation__round__n552 , _f_permutation__round__n551 ,
         _f_permutation__round__n550 , _f_permutation__round__n549 ,
         _f_permutation__round__n548 , _f_permutation__round__n547 ,
         _f_permutation__round__n546 , _f_permutation__round__n545 ,
         _f_permutation__round__n544 , _f_permutation__round__n543 ,
         _f_permutation__round__n542 , _f_permutation__round__n541 ,
         _f_permutation__round__n540 , _f_permutation__round__n539 ,
         _f_permutation__round__n538 , _f_permutation__round__n537 ,
         _f_permutation__round__n536 , _f_permutation__round__n535 ,
         _f_permutation__round__n534 , _f_permutation__round__n533 ,
         _f_permutation__round__n532 , _f_permutation__round__n531 ,
         _f_permutation__round__n530 , _f_permutation__round__n529 ,
         _f_permutation__round__n528 , _f_permutation__round__n527 ,
         _f_permutation__round__n526 , _f_permutation__round__n525 ,
         _f_permutation__round__n524 , _f_permutation__round__n523 ,
         _f_permutation__round__n522 , _f_permutation__round__n521 ,
         _f_permutation__round__n520 , _f_permutation__round__n519 ,
         _f_permutation__round__n518 , _f_permutation__round__n517 ,
         _f_permutation__round__n516 , _f_permutation__round__n515 ,
         _f_permutation__round__n514 , _f_permutation__round__n513 ,
         _f_permutation__round__n512 , _f_permutation__round__n511 ,
         _f_permutation__round__n510 , _f_permutation__round__n509 ,
         _f_permutation__round__n508 , _f_permutation__round__n507 ,
         _f_permutation__round__n506 , _f_permutation__round__n505 ,
         _f_permutation__round__n504 , _f_permutation__round__n503 ,
         _f_permutation__round__n502 , _f_permutation__round__n501 ,
         _f_permutation__round__n500 , _f_permutation__round__n499 ,
         _f_permutation__round__n498 , _f_permutation__round__n497 ,
         _f_permutation__round__n496 , _f_permutation__round__n495 ,
         _f_permutation__round__n494 , _f_permutation__round__n493 ,
         _f_permutation__round__n492 , _f_permutation__round__n491 ,
         _f_permutation__round__n490 , _f_permutation__round__n489 ,
         _f_permutation__round__n488 , _f_permutation__round__n487 ,
         _f_permutation__round__n486 , _f_permutation__round__n485 ,
         _f_permutation__round__n484 , _f_permutation__round__n483 ,
         _f_permutation__round__n482 , _f_permutation__round__n481 ,
         _f_permutation__round__n480 , _f_permutation__round__n479 ,
         _f_permutation__round__n478 , _f_permutation__round__n477 ,
         _f_permutation__round__n476 , _f_permutation__round__n475 ,
         _f_permutation__round__n474 , _f_permutation__round__n473 ,
         _f_permutation__round__n472 , _f_permutation__round__n471 ,
         _f_permutation__round__n470 , _f_permutation__round__n469 ,
         _f_permutation__round__n468 , _f_permutation__round__n467 ,
         _f_permutation__round__n466 , _f_permutation__round__n465 ,
         _f_permutation__round__n464 , _f_permutation__round__n463 ,
         _f_permutation__round__n462 , _f_permutation__round__n461 ,
         _f_permutation__round__n460 , _f_permutation__round__n459 ,
         _f_permutation__round__n458 , _f_permutation__round__n457 ,
         _f_permutation__round__n456 , _f_permutation__round__n455 ,
         _f_permutation__round__n454 , _f_permutation__round__n453 ,
         _f_permutation__round__n452 , _f_permutation__round__n451 ,
         _f_permutation__round__n450 , _f_permutation__round__n449 ,
         _f_permutation__round__n448 , _f_permutation__round__n447 ,
         _f_permutation__round__n446 , _f_permutation__round__n445 ,
         _f_permutation__round__n444 , _f_permutation__round__n443 ,
         _f_permutation__round__n442 , _f_permutation__round__n441 ,
         _f_permutation__round__n440 , _f_permutation__round__n439 ,
         _f_permutation__round__n438 , _f_permutation__round__n437 ,
         _f_permutation__round__n436 , _f_permutation__round__n435 ,
         _f_permutation__round__n434 , _f_permutation__round__n433 ,
         _f_permutation__round__n432 , _f_permutation__round__n431 ,
         _f_permutation__round__n430 , _f_permutation__round__n429 ,
         _f_permutation__round__n428 , _f_permutation__round__n427 ,
         _f_permutation__round__n426 , _f_permutation__round__n425 ,
         _f_permutation__round__n424 , _f_permutation__round__n423 ,
         _f_permutation__round__n422 , _f_permutation__round__n421 ,
         _f_permutation__round__n420 , _f_permutation__round__n419 ,
         _f_permutation__round__n418 , _f_permutation__round__n417 ,
         _f_permutation__round__n416 , _f_permutation__round__n415 ,
         _f_permutation__round__n414 , _f_permutation__round__n413 ,
         _f_permutation__round__n412 , _f_permutation__round__n411 ,
         _f_permutation__round__n410 , _f_permutation__round__n409 ,
         _f_permutation__round__n408 , _f_permutation__round__n407 ,
         _f_permutation__round__n406 , _f_permutation__round__n405 ,
         _f_permutation__round__n404 , _f_permutation__round__n403 ,
         _f_permutation__round__n402 , _f_permutation__round__n401 ,
         _f_permutation__round__n400 , _f_permutation__round__n399 ,
         _f_permutation__round__n398 , _f_permutation__round__n397 ,
         _f_permutation__round__n396 , _f_permutation__round__n395 ,
         _f_permutation__round__n394 , _f_permutation__round__n393 ,
         _f_permutation__round__n392 , _f_permutation__round__n391 ,
         _f_permutation__round__n390 , _f_permutation__round__n389 ,
         _f_permutation__round__n388 , _f_permutation__round__n387 ,
         _f_permutation__round__n386 , _f_permutation__round__n385 ,
         _f_permutation__round__n384 , _f_permutation__round__n383 ,
         _f_permutation__round__n382 , _f_permutation__round__n381 ,
         _f_permutation__round__n380 , _f_permutation__round__n379 ,
         _f_permutation__round__n378 , _f_permutation__round__n377 ,
         _f_permutation__round__n376 , _f_permutation__round__n375 ,
         _f_permutation__round__n374 , _f_permutation__round__n373 ,
         _f_permutation__round__n372 , _f_permutation__round__n371 ,
         _f_permutation__round__n370 , _f_permutation__round__n369 ,
         _f_permutation__round__n368 , _f_permutation__round__n367 ,
         _f_permutation__round__n366 , _f_permutation__round__n365 ,
         _f_permutation__round__n364 , _f_permutation__round__n363 ,
         _f_permutation__round__n362 , _f_permutation__round__n361 ,
         _f_permutation__round__n360 , _f_permutation__round__n359 ,
         _f_permutation__round__n358 , _f_permutation__round__n357 ,
         _f_permutation__round__n356 , _f_permutation__round__n355 ,
         _f_permutation__round__n354 , _f_permutation__round__n353 ,
         _f_permutation__round__n352 , _f_permutation__round__n351 ,
         _f_permutation__round__n350 , _f_permutation__round__n349 ,
         _f_permutation__round__n348 , _f_permutation__round__n347 ,
         _f_permutation__round__n346 , _f_permutation__round__n345 ,
         _f_permutation__round__n344 , _f_permutation__round__n343 ,
         _f_permutation__round__n342 , _f_permutation__round__n341 ,
         _f_permutation__round__n340 , _f_permutation__round__n339 ,
         _f_permutation__round__n338 , _f_permutation__round__n337 ,
         _f_permutation__round__n336 , _f_permutation__round__n335 ,
         _f_permutation__round__n334 , _f_permutation__round__n333 ,
         _f_permutation__round__n332 , _f_permutation__round__n331 ,
         _f_permutation__round__n330 , _f_permutation__round__n329 ,
         _f_permutation__round__n328 , _f_permutation__round__n327 ,
         _f_permutation__round__n326 , _f_permutation__round__n325 ,
         _f_permutation__round__n324 , _f_permutation__round__n323 ,
         _f_permutation__round__n322 , _f_permutation__round__n321 ,
         _f_permutation__round__n320 , _f_permutation__round__n319 ,
         _f_permutation__round__n318 , _f_permutation__round__n317 ,
         _f_permutation__round__n316 , _f_permutation__round__n315 ,
         _f_permutation__round__n314 , _f_permutation__round__n313 ,
         _f_permutation__round__n312 , _f_permutation__round__n311 ,
         _f_permutation__round__n310 , _f_permutation__round__n309 ,
         _f_permutation__round__n308 , _f_permutation__round__n307 ,
         _f_permutation__round__n306 , _f_permutation__round__n305 ,
         _f_permutation__round__n304 , _f_permutation__round__n303 ,
         _f_permutation__round__n302 , _f_permutation__round__n301 ,
         _f_permutation__round__n300 , _f_permutation__round__n299 ,
         _f_permutation__round__n298 , _f_permutation__round__n297 ,
         _f_permutation__round__n296 , _f_permutation__round__n295 ,
         _f_permutation__round__n294 , _f_permutation__round__n293 ,
         _f_permutation__round__n292 , _f_permutation__round__n291 ,
         _f_permutation__round__n290 , _f_permutation__round__n289 ,
         _f_permutation__round__n288 , _f_permutation__round__n287 ,
         _f_permutation__round__n286 , _f_permutation__round__n285 ,
         _f_permutation__round__n284 , _f_permutation__round__n283 ,
         _f_permutation__round__n282 , _f_permutation__round__n281 ,
         _f_permutation__round__n280 , _f_permutation__round__n279 ,
         _f_permutation__round__n278 , _f_permutation__round__n277 ,
         _f_permutation__round__n276 , _f_permutation__round__n275 ,
         _f_permutation__round__n274 , _f_permutation__round__n273 ,
         _f_permutation__round__n272 , _f_permutation__round__n271 ,
         _f_permutation__round__n270 , _f_permutation__round__n269 ,
         _f_permutation__round__n268 , _f_permutation__round__n267 ,
         _f_permutation__round__n266 , _f_permutation__round__n265 ,
         _f_permutation__round__n264 , _f_permutation__round__n263 ,
         _f_permutation__round__n262 , _f_permutation__round__n261 ,
         _f_permutation__round__n260 , _f_permutation__round__n259 ,
         _f_permutation__round__n258 , _f_permutation__round__n257 ,
         _f_permutation__round__n256 , _f_permutation__round__n255 ,
         _f_permutation__round__n254 , _f_permutation__round__n253 ,
         _f_permutation__round__n252 , _f_permutation__round__n251 ,
         _f_permutation__round__n250 , _f_permutation__round__n249 ,
         _f_permutation__round__n248 , _f_permutation__round__n247 ,
         _f_permutation__round__n246 , _f_permutation__round__n245 ,
         _f_permutation__round__n244 , _f_permutation__round__n243 ,
         _f_permutation__round__n242 , _f_permutation__round__n241 ,
         _f_permutation__round__n240 , _f_permutation__round__n239 ,
         _f_permutation__round__n238 , _f_permutation__round__n237 ,
         _f_permutation__round__n236 , _f_permutation__round__n235 ,
         _f_permutation__round__n234 , _f_permutation__round__n233 ,
         _f_permutation__round__n232 , _f_permutation__round__n231 ,
         _f_permutation__round__n230 , _f_permutation__round__n229 ,
         _f_permutation__round__n228 , _f_permutation__round__n227 ,
         _f_permutation__round__n226 , _f_permutation__round__n225 ,
         _f_permutation__round__n224 , _f_permutation__round__n223 ,
         _f_permutation__round__n222 , _f_permutation__round__n221 ,
         _f_permutation__round__n220 , _f_permutation__round__n219 ,
         _f_permutation__round__n218 , _f_permutation__round__n217 ,
         _f_permutation__round__n216 , _f_permutation__round__n215 ,
         _f_permutation__round__n214 , _f_permutation__round__n213 ,
         _f_permutation__round__n212 , _f_permutation__round__n211 ,
         _f_permutation__round__n210 , _f_permutation__round__n209 ,
         _f_permutation__round__n208 , _f_permutation__round__n207 ,
         _f_permutation__round__n206 , _f_permutation__round__n205 ,
         _f_permutation__round__n204 , _f_permutation__round__n203 ,
         _f_permutation__round__n202 , _f_permutation__round__n201 ,
         _f_permutation__round__n200 , _f_permutation__round__n199 ,
         _f_permutation__round__n198 , _f_permutation__round__n197 ,
         _f_permutation__round__n196 , _f_permutation__round__n195 ,
         _f_permutation__round__n194 , _f_permutation__round__n193 ,
         _f_permutation__round__n192 , _f_permutation__round__n191 ,
         _f_permutation__round__n190 , _f_permutation__round__n189 ,
         _f_permutation__round__n188 , _f_permutation__round__n187 ,
         _f_permutation__round__n186 , _f_permutation__round__n185 ,
         _f_permutation__round__n184 , _f_permutation__round__n183 ,
         _f_permutation__round__n182 , _f_permutation__round__n181 ,
         _f_permutation__round__n180 , _f_permutation__round__n179 ,
         _f_permutation__round__n178 , _f_permutation__round__n177 ,
         _f_permutation__round__n176 , _f_permutation__round__n175 ,
         _f_permutation__round__n174 , _f_permutation__round__n173 ,
         _f_permutation__round__n172 , _f_permutation__round__n171 ,
         _f_permutation__round__n170 , _f_permutation__round__n169 ,
         _f_permutation__round__n168 , _f_permutation__round__n167 ,
         _f_permutation__round__n166 , _f_permutation__round__n165 ,
         _f_permutation__round__n164 , _f_permutation__round__n163 ,
         _f_permutation__round__n162 , _f_permutation__round__n161 ,
         _f_permutation__round__n160 , _f_permutation__round__n159 ,
         _f_permutation__round__n158 , _f_permutation__round__n157 ,
         _f_permutation__round__n156 , _f_permutation__round__n155 ,
         _f_permutation__round__n154 , _f_permutation__round__n153 ,
         _f_permutation__round__n152 , _f_permutation__round__n151 ,
         _f_permutation__round__n150 , _f_permutation__round__n149 ,
         _f_permutation__round__n148 , _f_permutation__round__n147 ,
         _f_permutation__round__n146 , _f_permutation__round__n145 ,
         _f_permutation__round__n144 , _f_permutation__round__n143 ,
         _f_permutation__round__n142 , _f_permutation__round__n141 ,
         _f_permutation__round__n140 , _f_permutation__round__n139 ,
         _f_permutation__round__n138 , _f_permutation__round__n137 ,
         _f_permutation__round__n136 , _f_permutation__round__n135 ,
         _f_permutation__round__n134 , _f_permutation__round__n133 ,
         _f_permutation__round__n132 , _f_permutation__round__n131 ,
         _f_permutation__round__n130 , _f_permutation__round__n129 ,
         _f_permutation__round__n128 , _f_permutation__round__n127 ,
         _f_permutation__round__n126 , _f_permutation__round__n125 ,
         _f_permutation__round__n124 , _f_permutation__round__n123 ,
         _f_permutation__round__n122 , _f_permutation__round__n121 ,
         _f_permutation__round__n120 , _f_permutation__round__n119 ,
         _f_permutation__round__n118 , _f_permutation__round__n117 ,
         _f_permutation__round__n116 , _f_permutation__round__n115 ,
         _f_permutation__round__n114 , _f_permutation__round__n113 ,
         _f_permutation__round__n112 , _f_permutation__round__n111 ,
         _f_permutation__round__n110 , _f_permutation__round__n109 ,
         _f_permutation__round__n108 , _f_permutation__round__n107 ,
         _f_permutation__round__n106 , _f_permutation__round__n105 ,
         _f_permutation__round__n104 , _f_permutation__round__n103 ,
         _f_permutation__round__n102 , _f_permutation__round__n101 ,
         _f_permutation__round__n100 , _f_permutation__round__n99 ,
         _f_permutation__round__n98 , _f_permutation__round__n97 ,
         _f_permutation__round__n96 , _f_permutation__round__n95 ,
         _f_permutation__round__n94 , _f_permutation__round__n93 ,
         _f_permutation__round__n92 , _f_permutation__round__n91 ,
         _f_permutation__round__n90 , _f_permutation__round__n89 ,
         _f_permutation__round__n88 , _f_permutation__round__n87 ,
         _f_permutation__round__n86 , _f_permutation__round__n85 ,
         _f_permutation__round__n84 , _f_permutation__round__n83 ,
         _f_permutation__round__n82 , _f_permutation__round__n81 ,
         _f_permutation__round__n80 , _f_permutation__round__n79 ,
         _f_permutation__round__n78 , _f_permutation__round__n77 ,
         _f_permutation__round__n76 , _f_permutation__round__n75 ,
         _f_permutation__round__n74 , _f_permutation__round__n73 ,
         _f_permutation__round__n72 , _f_permutation__round__n71 ,
         _f_permutation__round__n70 , _f_permutation__round__n69 ,
         _f_permutation__round__n68 , _f_permutation__round__n67 ,
         _f_permutation__round__n66 , _f_permutation__round__n65 ,
         _f_permutation__round__n64 , _f_permutation__round__n63 ,
         _f_permutation__round__n62 , _f_permutation__round__n61 ,
         _f_permutation__round__n60 , _f_permutation__round__n59 ,
         _f_permutation__round__n58 , _f_permutation__round__n57 ,
         _f_permutation__round__n56 , _f_permutation__round__n55 ,
         _f_permutation__round__n54 , _f_permutation__round__n53 ,
         _f_permutation__round__n52 , _f_permutation__round__n51 ,
         _f_permutation__round__n50 , _f_permutation__round__n49 ,
         _f_permutation__round__n48 , _f_permutation__round__n47 ,
         _f_permutation__round__n46 , _f_permutation__round__n45 ,
         _f_permutation__round__n44 , _f_permutation__round__n43 ,
         _f_permutation__round__n42 , _f_permutation__round__n41 ,
         _f_permutation__round__n40 , _f_permutation__round__n39 ,
         _f_permutation__round__n38 , _f_permutation__round__n37 ,
         _f_permutation__round__n36 , _f_permutation__round__n35 ,
         _f_permutation__round__n34 , _f_permutation__round__n33 ,
         _f_permutation__round__n32 , _f_permutation__round__n31 ,
         _f_permutation__round__n30 , _f_permutation__round__n29 ,
         _f_permutation__round__n28 , _f_permutation__round__n27 ,
         _f_permutation__round__n26 , _f_permutation__round__n25 ,
         _f_permutation__round__n24 , _f_permutation__round__n23 ,
         _f_permutation__round__n22 , _f_permutation__round__n21 ,
         _f_permutation__round__n20 , _f_permutation__round__n19 ,
         _f_permutation__round__n18 , _f_permutation__round__n17 ,
         _f_permutation__round__n16 , _f_permutation__round__n15 ,
         _f_permutation__round__n14 , _f_permutation__round__n13 ,
         _f_permutation__round__n12 , _f_permutation__round__n11 ,
         _f_permutation__round__n10 , _f_permutation__round__n9 ,
         _f_permutation__round__n8 , _f_permutation__round__n7 ,
         _f_permutation__round__n6 , _f_permutation__round__n5 ,
         _f_permutation__round__n4 , _f_permutation__round__n3 ,
         _f_permutation__round__n2 , _f_permutation__round__n1 ,
         _f_permutation__round__n25670 , _f_permutation__round__n2566 ,
         _f_permutation__round__n25650 , _f_permutation__round__n2564 ,
         _f_permutation__round__n25630 , _f_permutation__round__n2562 ,
         _f_permutation__round__n25610 , _f_permutation__round__n2560 ,
         _f_permutation__round__n2559 , _f_permutation__round__n2558 ,
         _f_permutation__round__n2557 , _f_permutation__round__n2556 ,
         _f_permutation__round__n2555 , _f_permutation__round__n2554 ,
         _f_permutation__round__n2553 , _f_permutation__round__n2552 ,
         _f_permutation__round__n2551 , _f_permutation__round__n2550 ,
         _f_permutation__round__n2549 , _f_permutation__round__n2548 ,
         _f_permutation__round__n2547 , _f_permutation__round__n2546 ,
         _f_permutation__round__n2545 , _f_permutation__round__n2544 ,
         _f_permutation__round__n2543 , _f_permutation__round__n2542 ,
         _f_permutation__round__n2541 , _f_permutation__round__n2540 ,
         _f_permutation__round__n2539 , _f_permutation__round__n2538 ,
         _f_permutation__round__n2537 , _f_permutation__round__n2536 ,
         _f_permutation__round__n2535 , _f_permutation__round__n2534 ,
         _f_permutation__round__n2533 , _f_permutation__round__n2532 ,
         _f_permutation__round__n2531 , _f_permutation__round__n2530 ,
         _f_permutation__round__n2529 , _f_permutation__round__n2528 ,
         _f_permutation__round__n2527 , _f_permutation__round__n2526 ,
         _f_permutation__round__n2525 , _f_permutation__round__n2524 ,
         _f_permutation__round__n2523 , _f_permutation__round__n2522 ,
         _f_permutation__round__n2521 , _f_permutation__round__n2520 ,
         _f_permutation__round__n2519 , _f_permutation__round__n2518 ,
         _f_permutation__round__n2517 , _f_permutation__round__n2516 ,
         _f_permutation__round__n2515 , _f_permutation__round__n2514 ,
         _f_permutation__round__n2513 , _f_permutation__round__n2512 ,
         _f_permutation__round__n2511 , _f_permutation__round__n2510 ,
         _f_permutation__round__n2509 , _f_permutation__round__n2508 ,
         _f_permutation__round__n2507 , _f_permutation__round__n2506 ,
         _f_permutation__round__n2505 , _f_permutation__round__n2504 ,
         _f_permutation__round__n2503 , _f_permutation__round__n2502 ,
         _f_permutation__round__n2501 , _f_permutation__round__n2500 ,
         _f_permutation__round__n2499 , _f_permutation__round__n2498 ,
         _f_permutation__round__n2497 , _f_permutation__round__n2496 ,
         _f_permutation__round__n2495 , _f_permutation__round__n2494 ,
         _f_permutation__round__n2493 , _f_permutation__round__n2492 ,
         _f_permutation__round__n2491 , _f_permutation__round__n2490 ,
         _f_permutation__round__n2489 , _f_permutation__round__n2488 ,
         _f_permutation__round__n2487 , _f_permutation__round__n2486 ,
         _f_permutation__round__n2485 , _f_permutation__round__n2484 ,
         _f_permutation__round__n2483 , _f_permutation__round__n2482 ,
         _f_permutation__round__n2481 , _f_permutation__round__n2480 ,
         _f_permutation__round__n2479 , _f_permutation__round__n2478 ,
         _f_permutation__round__n2477 , _f_permutation__round__n2476 ,
         _f_permutation__round__n2475 , _f_permutation__round__n2474 ,
         _f_permutation__round__n2473 , _f_permutation__round__n2472 ,
         _f_permutation__round__n2471 , _f_permutation__round__n2470 ,
         _f_permutation__round__n2469 , _f_permutation__round__n2468 ,
         _f_permutation__round__n2467 , _f_permutation__round__n2466 ,
         _f_permutation__round__n2465 , _f_permutation__round__n2464 ,
         _f_permutation__round__n2463 , _f_permutation__round__n2462 ,
         _f_permutation__round__n2461 , _f_permutation__round__n2460 ,
         _f_permutation__round__n2459 , _f_permutation__round__n2458 ,
         _f_permutation__round__n2457 , _f_permutation__round__n2456 ,
         _f_permutation__round__n2455 , _f_permutation__round__n2454 ,
         _f_permutation__round__n2453 , _f_permutation__round__n2452 ,
         _f_permutation__round__n2451 , _f_permutation__round__n2450 ,
         _f_permutation__round__n2449 , _f_permutation__round__n2448 ,
         _f_permutation__round__n2447 , _f_permutation__round__n2446 ,
         _f_permutation__round__n2445 , _f_permutation__round__n2444 ,
         _f_permutation__round__n2443 , _f_permutation__round__n2442 ,
         _f_permutation__round__n2441 , _f_permutation__round__n2440 ,
         _f_permutation__round__n2439 , _f_permutation__round__n2438 ,
         _f_permutation__round__n2437 , _f_permutation__round__n2436 ,
         _f_permutation__round__n2435 , _f_permutation__round__n2434 ,
         _f_permutation__round__n2433 , _f_permutation__round__n2432 ,
         _f_permutation__round__n2431 , _f_permutation__round__n2430 ,
         _f_permutation__round__n2429 , _f_permutation__round__n2428 ,
         _f_permutation__round__n2427 , _f_permutation__round__n2426 ,
         _f_permutation__round__n2425 , _f_permutation__round__n2424 ,
         _f_permutation__round__n2423 , _f_permutation__round__n2422 ,
         _f_permutation__round__n2421 , _f_permutation__round__n2420 ,
         _f_permutation__round__n2419 , _f_permutation__round__n2418 ,
         _f_permutation__round__n2417 , _f_permutation__round__n2416 ,
         _f_permutation__round__n2415 , _f_permutation__round__n2414 ,
         _f_permutation__round__n2413 , _f_permutation__round__n2412 ,
         _f_permutation__round__n2411 , _f_permutation__round__n2410 ,
         _f_permutation__round__n2409 , _f_permutation__round__n2408 ,
         _f_permutation__round__n2407 , _f_permutation__round__n2406 ,
         _f_permutation__round__n2405 , _f_permutation__round__n2404 ,
         _f_permutation__round__n2403 , _f_permutation__round__n2402 ,
         _f_permutation__round__n2401 , _f_permutation__round__n2400 ,
         _f_permutation__round__n2399 , _f_permutation__round__n2398 ,
         _f_permutation__round__n2397 , _f_permutation__round__n2396 ,
         _f_permutation__round__n2395 , _f_permutation__round__n2394 ,
         _f_permutation__round__n2393 , _f_permutation__round__n2392 ,
         _f_permutation__round__n2391 , _f_permutation__round__n2390 ,
         _f_permutation__round__n2389 , _f_permutation__round__n2388 ,
         _f_permutation__round__n2387 , _f_permutation__round__n2386 ,
         _f_permutation__round__n2385 , _f_permutation__round__n2384 ,
         _f_permutation__round__n2383 , _f_permutation__round__n2382 ,
         _f_permutation__round__n2381 , _f_permutation__round__n2380 ,
         _f_permutation__round__n2379 , _f_permutation__round__n2378 ,
         _f_permutation__round__n2377 , _f_permutation__round__n2376 ,
         _f_permutation__round__n2375 , _f_permutation__round__n2374 ,
         _f_permutation__round__n2373 , _f_permutation__round__n2372 ,
         _f_permutation__round__n2371 , _f_permutation__round__n2370 ,
         _f_permutation__round__n2369 , _f_permutation__round__n2368 ,
         _f_permutation__round__n2367 , _f_permutation__round__n2366 ,
         _f_permutation__round__n2365 , _f_permutation__round__n2364 ,
         _f_permutation__round__n2363 , _f_permutation__round__n2362 ,
         _f_permutation__round__n2361 , _f_permutation__round__n2360 ,
         _f_permutation__round__n2359 , _f_permutation__round__n2358 ,
         _f_permutation__round__n2357 , _f_permutation__round__n2356 ,
         _f_permutation__round__n2355 , _f_permutation__round__n2354 ,
         _f_permutation__round__n2353 , _f_permutation__round__n2352 ,
         _f_permutation__round__n2351 , _f_permutation__round__n2350 ,
         _f_permutation__round__n2349 , _f_permutation__round__n2348 ,
         _f_permutation__round__n2347 , _f_permutation__round__n2346 ,
         _f_permutation__round__n2345 , _f_permutation__round__n2344 ,
         _f_permutation__round__n2343 , _f_permutation__round__n2342 ,
         _f_permutation__round__n2341 , _f_permutation__round__n2340 ,
         _f_permutation__round__n2339 , _f_permutation__round__n2338 ,
         _f_permutation__round__n2337 , _f_permutation__round__n2336 ,
         _f_permutation__round__n2335 , _f_permutation__round__n2334 ,
         _f_permutation__round__n2333 , _f_permutation__round__n2332 ,
         _f_permutation__round__n2331 , _f_permutation__round__n2330 ,
         _f_permutation__round__n2329 , _f_permutation__round__n2328 ,
         _f_permutation__round__n2327 , _f_permutation__round__n2326 ,
         _f_permutation__round__n2325 , _f_permutation__round__n2324 ,
         _f_permutation__round__n2323 , _f_permutation__round__n2322 ,
         _f_permutation__round__n2321 , _f_permutation__round__n2320 ,
         _f_permutation__round__n2319 , _f_permutation__round__n2318 ,
         _f_permutation__round__n2317 , _f_permutation__round__n2316 ,
         _f_permutation__round__n2315 , _f_permutation__round__n2314 ,
         _f_permutation__round__n2313 , _f_permutation__round__n2312 ,
         _f_permutation__round__n2311 , _f_permutation__round__n2310 ,
         _f_permutation__round__n2309 , _f_permutation__round__n2308 ,
         _f_permutation__round__n2307 , _f_permutation__round__n2306 ,
         _f_permutation__round__n2305 , _f_permutation__round__n2304 ,
         _f_permutation__round__n2303 , _f_permutation__round__n2302 ,
         _f_permutation__round__n2301 , _f_permutation__round__n2300 ,
         _f_permutation__round__n2299 , _f_permutation__round__n2298 ,
         _f_permutation__round__n2297 , _f_permutation__round__n2296 ,
         _f_permutation__round__n2295 , _f_permutation__round__n2294 ,
         _f_permutation__round__n2293 , _f_permutation__round__n2292 ,
         _f_permutation__round__n2291 , _f_permutation__round__n2290 ,
         _f_permutation__round__n2289 , _f_permutation__round__n2288 ,
         _f_permutation__round__n2287 , _f_permutation__round__n2286 ,
         _f_permutation__round__n2285 , _f_permutation__round__n2284 ,
         _f_permutation__round__n2283 , _f_permutation__round__n2282 ,
         _f_permutation__round__n2281 , _f_permutation__round__n2280 ,
         _f_permutation__round__n2279 , _f_permutation__round__n2278 ,
         _f_permutation__round__n2277 , _f_permutation__round__n2276 ,
         _f_permutation__round__n2275 , _f_permutation__round__n2274 ,
         _f_permutation__round__n2273 , _f_permutation__round__n2272 ,
         _f_permutation__round__n2271 , _f_permutation__round__n2270 ,
         _f_permutation__round__n2269 , _f_permutation__round__n2268 ,
         _f_permutation__round__n2267 , _f_permutation__round__n2266 ,
         _f_permutation__round__n2265 , _f_permutation__round__n2264 ,
         _f_permutation__round__n2263 , _f_permutation__round__n2262 ,
         _f_permutation__round__n2261 , _f_permutation__round__n2260 ,
         _f_permutation__round__n2259 , _f_permutation__round__n2258 ,
         _f_permutation__round__n2257 , _f_permutation__round__n2256 ,
         _f_permutation__round__n2255 , _f_permutation__round__n2254 ,
         _f_permutation__round__n2253 , _f_permutation__round__n2252 ,
         _f_permutation__round__n2251 , _f_permutation__round__n2250 ,
         _f_permutation__round__n2249 , _f_permutation__round__n2248 ,
         _f_permutation__round__n2247 , _f_permutation__round__n2246 ,
         _f_permutation__round__n2245 , _f_permutation__round__n2244 ,
         _f_permutation__round__n2243 , _f_permutation__round__n2242 ,
         _f_permutation__round__n2241 , _f_permutation__round__n2240 ,
         _f_permutation__round__n2239 , _f_permutation__round__n2238 ,
         _f_permutation__round__n2237 , _f_permutation__round__n2236 ,
         _f_permutation__round__n2235 , _f_permutation__round__n2234 ,
         _f_permutation__round__n2233 , _f_permutation__round__n2232 ,
         _f_permutation__round__n2231 , _f_permutation__round__n2230 ,
         _f_permutation__round__n2229 , _f_permutation__round__n2228 ,
         _f_permutation__round__n2227 , _f_permutation__round__n2226 ,
         _f_permutation__round__n2225 , _f_permutation__round__n2224 ,
         _f_permutation__round__n2223 , _f_permutation__round__n2222 ,
         _f_permutation__round__n2221 , _f_permutation__round__n2220 ,
         _f_permutation__round__n2219 , _f_permutation__round__n2218 ,
         _f_permutation__round__n2217 , _f_permutation__round__n2216 ,
         _f_permutation__round__n2215 , _f_permutation__round__n2214 ,
         _f_permutation__round__n2213 , _f_permutation__round__n2212 ,
         _f_permutation__round__n2211 , _f_permutation__round__n2210 ,
         _f_permutation__round__n2209 , _f_permutation__round__n2208 ,
         _f_permutation__round__n2207 , _f_permutation__round__n2206 ,
         _f_permutation__round__n2205 , _f_permutation__round__n2204 ,
         _f_permutation__round__n2203 , _f_permutation__round__n2202 ,
         _f_permutation__round__n2201 , _f_permutation__round__n2200 ,
         _f_permutation__round__n2199 , _f_permutation__round__n2198 ,
         _f_permutation__round__n2197 , _f_permutation__round__n2196 ,
         _f_permutation__round__n2195 , _f_permutation__round__n2194 ,
         _f_permutation__round__n2193 , _f_permutation__round__n2192 ,
         _f_permutation__round__n2191 , _f_permutation__round__n2190 ,
         _f_permutation__round__n2189 , _f_permutation__round__n2188 ,
         _f_permutation__round__n2187 , _f_permutation__round__n2186 ,
         _f_permutation__round__n2185 , _f_permutation__round__n2184 ,
         _f_permutation__round__n2183 , _f_permutation__round__n2182 ,
         _f_permutation__round__n2181 , _f_permutation__round__n2180 ,
         _f_permutation__round__n2179 , _f_permutation__round__n2178 ,
         _f_permutation__round__n2177 , _f_permutation__round__n2176 ,
         _f_permutation__round__n2175 , _f_permutation__round__n2174 ,
         _f_permutation__round__n2173 , _f_permutation__round__n2172 ,
         _f_permutation__round__n2171 , _f_permutation__round__n2170 ,
         _f_permutation__round__n2169 , _f_permutation__round__n2168 ,
         _f_permutation__round__n2167 , _f_permutation__round__n2166 ,
         _f_permutation__round__n2165 , _f_permutation__round__n2164 ,
         _f_permutation__round__n2163 , _f_permutation__round__n2162 ,
         _f_permutation__round__n2161 , _f_permutation__round__n2160 ,
         _f_permutation__round__n2159 , _f_permutation__round__n2158 ,
         _f_permutation__round__n2157 , _f_permutation__round__n2156 ,
         _f_permutation__round__n2155 , _f_permutation__round__n2154 ,
         _f_permutation__round__n2153 , _f_permutation__round__n2152 ,
         _f_permutation__round__n2151 , _f_permutation__round__n2150 ,
         _f_permutation__round__n2149 , _f_permutation__round__n2148 ,
         _f_permutation__round__n2147 , _f_permutation__round__n2146 ,
         _f_permutation__round__n2145 , _f_permutation__round__n2144 ,
         _f_permutation__round__n2143 , _f_permutation__round__n2142 ,
         _f_permutation__round__n2141 , _f_permutation__round__n2140 ,
         _f_permutation__round__n2139 , _f_permutation__round__n2138 ,
         _f_permutation__round__n2137 , _f_permutation__round__n2136 ,
         _f_permutation__round__n2135 , _f_permutation__round__n2134 ,
         _f_permutation__round__n2133 , _f_permutation__round__n2132 ,
         _f_permutation__round__n2131 , _f_permutation__round__n2130 ,
         _f_permutation__round__n2129 , _f_permutation__round__n2128 ,
         _f_permutation__round__n2127 , _f_permutation__round__n2126 ,
         _f_permutation__round__n2125 , _f_permutation__round__n2124 ,
         _f_permutation__round__n2123 , _f_permutation__round__n2122 ,
         _f_permutation__round__n2121 , _f_permutation__round__n2120 ,
         _f_permutation__round__n2119 , _f_permutation__round__n2118 ,
         _f_permutation__round__n2117 , _f_permutation__round__n2116 ,
         _f_permutation__round__n2115 , _f_permutation__round__n2114 ,
         _f_permutation__round__n2113 , _f_permutation__round__n2112 ,
         _f_permutation__round__n2111 , _f_permutation__round__n2110 ,
         _f_permutation__round__n2109 , _f_permutation__round__n2108 ,
         _f_permutation__round__n2107 , _f_permutation__round__n2106 ,
         _f_permutation__round__n2105 , _f_permutation__round__n2104 ,
         _f_permutation__round__n2103 , _f_permutation__round__n2102 ,
         _f_permutation__round__n2101 , _f_permutation__round__n2100 ,
         _f_permutation__round__n2099 , _f_permutation__round__n2098 ,
         _f_permutation__round__n2097 , _f_permutation__round__n2096 ,
         _f_permutation__round__n2095 , _f_permutation__round__n2094 ,
         _f_permutation__round__n2093 , _f_permutation__round__n2092 ,
         _f_permutation__round__n2091 , _f_permutation__round__n2090 ,
         _f_permutation__round__n2089 , _f_permutation__round__n2088 ,
         _f_permutation__round__n2087 , _f_permutation__round__n2086 ,
         _f_permutation__round__n2085 , _f_permutation__round__n2084 ,
         _f_permutation__round__n2083 , _f_permutation__round__n2082 ,
         _f_permutation__round__n2081 , _f_permutation__round__n2080 ,
         _f_permutation__round__n2079 , _f_permutation__round__n2078 ,
         _f_permutation__round__n2077 , _f_permutation__round__n2076 ,
         _f_permutation__round__n2075 , _f_permutation__round__n2074 ,
         _f_permutation__round__n2073 , _f_permutation__round__n2072 ,
         _f_permutation__round__n2071 , _f_permutation__round__n2070 ,
         _f_permutation__round__n2069 , _f_permutation__round__n2068 ,
         _f_permutation__round__n2067 , _f_permutation__round__n2066 ,
         _f_permutation__round__n2065 , _f_permutation__round__n2064 ,
         _f_permutation__round__n2063 , _f_permutation__round__n2062 ,
         _f_permutation__round__n2061 , _f_permutation__round__n2060 ,
         _f_permutation__round__n2059 , _f_permutation__round__n2058 ,
         _f_permutation__round__n2057 , _f_permutation__round__n2056 ,
         _f_permutation__round__n2055 , _f_permutation__round__n2054 ,
         _f_permutation__round__n2053 , _f_permutation__round__n2052 ,
         _f_permutation__round__n2051 , _f_permutation__round__n2050 ,
         _f_permutation__round__n2049 , _f_permutation__round__n2048 ,
         _f_permutation__round__n2047 , _f_permutation__round__n2046 ,
         _f_permutation__round__n2045 , _f_permutation__round__n2044 ,
         _f_permutation__round__n2043 , _f_permutation__round__n2042 ,
         _f_permutation__round__n2041 , _f_permutation__round__n2040 ,
         _f_permutation__round__n2039 , _f_permutation__round__n2038 ,
         _f_permutation__round__n2037 , _f_permutation__round__n2036 ,
         _f_permutation__round__n2035 , _f_permutation__round__n2034 ,
         _f_permutation__round__n2033 , _f_permutation__round__n2032 ,
         _f_permutation__round__n2031 , _f_permutation__round__n2030 ,
         _f_permutation__round__n2029 , _f_permutation__round__n2028 ,
         _f_permutation__round__n2027 , _f_permutation__round__n2026 ,
         _f_permutation__round__n2025 , _f_permutation__round__n2024 ,
         _f_permutation__round__n2023 , _f_permutation__round__n2022 ,
         _f_permutation__round__n2021 , _f_permutation__round__n2020 ,
         _f_permutation__round__n2019 , _f_permutation__round__n2018 ,
         _f_permutation__round__n2017 , _f_permutation__round__n2016 ,
         _f_permutation__round__n2015 , _f_permutation__round__n2014 ,
         _f_permutation__round__n2013 , _f_permutation__round__n2012 ,
         _f_permutation__round__n2011 , _f_permutation__round__n2010 ,
         _f_permutation__round__n2009 , _f_permutation__round__n2008 ,
         _f_permutation__round__n2007 , _f_permutation__round__n2006 ,
         _f_permutation__round__n2005 , _f_permutation__round__n2004 ,
         _f_permutation__round__n2003 , _f_permutation__round__n2002 ,
         _f_permutation__round__n2001 , _f_permutation__round__n2000 ,
         _f_permutation__round__n1999 , _f_permutation__round__n1998 ,
         _f_permutation__round__n1997 , _f_permutation__round__n1996 ,
         _f_permutation__round__n1995 , _f_permutation__round__n1994 ,
         _f_permutation__round__n1993 , _f_permutation__round__n1992 ,
         _f_permutation__round__n1991 , _f_permutation__round__n1990 ,
         _f_permutation__round__n1989 , _f_permutation__round__n1988 ,
         _f_permutation__round__n1987 , _f_permutation__round__n1986 ,
         _f_permutation__round__n1985 , _f_permutation__round__n1984 ,
         _f_permutation__round__n1983 , _f_permutation__round__n1982 ,
         _f_permutation__round__n1981 , _f_permutation__round__n1980 ,
         _f_permutation__round__n1979 , _f_permutation__round__n1978 ,
         _f_permutation__round__n1977 , _f_permutation__round__n1976 ,
         _f_permutation__round__n1975 , _f_permutation__round__n1974 ,
         _f_permutation__round__n1973 , _f_permutation__round__n1972 ,
         _f_permutation__round__n1971 , _f_permutation__round__n1970 ,
         _f_permutation__round__n1969 , _f_permutation__round__n1968 ,
         _f_permutation__round__n1967 , _f_permutation__round__n1966 ,
         _f_permutation__round__n1965 , _f_permutation__round__n1964 ,
         _f_permutation__round__n1963 , _f_permutation__round__n1962 ,
         _f_permutation__round__n1961 , _f_permutation__round__n1960 ,
         _f_permutation__round__n1959 , _f_permutation__round__n1958 ,
         _f_permutation__round__n1957 , _f_permutation__round__n1956 ,
         _f_permutation__round__n1955 , _f_permutation__round__n1954 ,
         _f_permutation__round__n1953 , _f_permutation__round__n1952 ,
         _f_permutation__round__n1951 , _f_permutation__round__n1950 ,
         _f_permutation__round__n1949 , _f_permutation__round__n1948 ,
         _f_permutation__round__n1947 , _f_permutation__round__n1946 ,
         _f_permutation__round__n1945 , _f_permutation__round__n1944 ,
         _f_permutation__round__n1943 , _f_permutation__round__n1942 ,
         _f_permutation__round__n1941 , _f_permutation__round__n1940 ,
         _f_permutation__round__n1939 , _f_permutation__round__n1938 ,
         _f_permutation__round__n1937 , _f_permutation__round__n1936 ,
         _f_permutation__round__n1935 , _f_permutation__round__n1934 ,
         _f_permutation__round__n1933 , _f_permutation__round__n1932 ,
         _f_permutation__round__n1931 , _f_permutation__round__n1930 ,
         _f_permutation__round__n1929 , _f_permutation__round__n1928 ,
         _f_permutation__round__n1927 , _f_permutation__round__n1926 ,
         _f_permutation__round__n1925 , _f_permutation__round__n1924 ,
         _f_permutation__round__n1923 , _f_permutation__round__n1922 ,
         _f_permutation__round__n1921 , _f_permutation__round__n1920 ,
         _f_permutation__round__n1919 , _f_permutation__round__n1918 ,
         _f_permutation__round__n1917 , _f_permutation__round__n1916 ,
         _f_permutation__round__n1915 , _f_permutation__round__n1914 ,
         _f_permutation__round__n1913 , _f_permutation__round__n1912 ,
         _f_permutation__round__n1911 , _f_permutation__round__n1910 ,
         _f_permutation__round__n1909 , _f_permutation__round__n1908 ,
         _f_permutation__round__n1907 , _f_permutation__round__n1906 ,
         _f_permutation__round__n1905 , _f_permutation__round__n1904 ,
         _f_permutation__round__n1903 , _f_permutation__round__n1902 ,
         _f_permutation__round__n1901 , _f_permutation__round__n1900 ,
         _f_permutation__round__n1899 , _f_permutation__round__n1898 ,
         _f_permutation__round__n1897 , _f_permutation__round__n1896 ,
         _f_permutation__round__n1895 , _f_permutation__round__n1894 ,
         _f_permutation__round__n1893 , _f_permutation__round__n1892 ,
         _f_permutation__round__n1891 , _f_permutation__round__n1890 ,
         _f_permutation__round__n1889 , _f_permutation__round__n1888 ,
         _f_permutation__round__n1887 , _f_permutation__round__n1886 ,
         _f_permutation__round__n1885 , _f_permutation__round__n1884 ,
         _f_permutation__round__n1883 , _f_permutation__round__n1882 ,
         _f_permutation__round__n1881 , _f_permutation__round__n1880 ,
         _f_permutation__round__n1879 , _f_permutation__round__n1878 ,
         _f_permutation__round__n1877 , _f_permutation__round__n1876 ,
         _f_permutation__round__n1875 , _f_permutation__round__n1874 ,
         _f_permutation__round__n1873 , _f_permutation__round__n1872 ,
         _f_permutation__round__n1871 , _f_permutation__round__n1870 ,
         _f_permutation__round__n1869 , _f_permutation__round__n1868 ,
         _f_permutation__round__n1867 , _f_permutation__round__n1866 ,
         _f_permutation__round__n1865 , _f_permutation__round__n1864 ,
         _f_permutation__round__n1863 , _f_permutation__round__n1862 ,
         _f_permutation__round__n1861 , _f_permutation__round__n1860 ,
         _f_permutation__round__n1859 , _f_permutation__round__n1858 ,
         _f_permutation__round__n1857 , _f_permutation__round__n1856 ,
         _f_permutation__round__n1855 , _f_permutation__round__n1854 ,
         _f_permutation__round__n1853 , _f_permutation__round__n1852 ,
         _f_permutation__round__n1851 , _f_permutation__round__n1850 ,
         _f_permutation__round__n1849 , _f_permutation__round__n1848 ,
         _f_permutation__round__n1847 , _f_permutation__round__n1846 ,
         _f_permutation__round__n1845 , _f_permutation__round__n1844 ,
         _f_permutation__round__n1843 , _f_permutation__round__n1842 ,
         _f_permutation__round__n1841 , _f_permutation__round__n1840 ,
         _f_permutation__round__n1839 , _f_permutation__round__n1838 ,
         _f_permutation__round__n1837 , _f_permutation__round__n1836 ,
         _f_permutation__round__n1835 , _f_permutation__round__n1834 ,
         _f_permutation__round__n1833 , _f_permutation__round__n1832 ,
         _f_permutation__round__n1831 , _f_permutation__round__n1830 ,
         _f_permutation__round__n1829 , _f_permutation__round__n1828 ,
         _f_permutation__round__n1827 , _f_permutation__round__n1826 ,
         _f_permutation__round__n1825 , _f_permutation__round__n1824 ,
         _f_permutation__round__n1823 , _f_permutation__round__n1822 ,
         _f_permutation__round__n1821 , _f_permutation__round__n1820 ,
         _f_permutation__round__n1819 , _f_permutation__round__n1818 ,
         _f_permutation__round__n1817 , _f_permutation__round__n1816 ,
         _f_permutation__round__n1815 , _f_permutation__round__n1814 ,
         _f_permutation__round__n1813 , _f_permutation__round__n1812 ,
         _f_permutation__round__n1811 , _f_permutation__round__n1810 ,
         _f_permutation__round__n1809 , _f_permutation__round__n1808 ,
         _f_permutation__round__n1807 , _f_permutation__round__n1806 ,
         _f_permutation__round__n1805 , _f_permutation__round__n1804 ,
         _f_permutation__round__n1803 , _f_permutation__round__n1802 ,
         _f_permutation__round__n1801 , _f_permutation__round__n1800 ,
         _f_permutation__round__n1799 , _f_permutation__round__n1798 ,
         _f_permutation__round__n1797 , _f_permutation__round__n1796 ,
         _f_permutation__round__n1795 , _f_permutation__round__n1794 ,
         _f_permutation__round__n1793 , _f_permutation__round__n1792 ,
         _f_permutation__round__n1791 , _f_permutation__round__n1790 ,
         _f_permutation__round__n1789 , _f_permutation__round__n1788 ,
         _f_permutation__round__n1787 , _f_permutation__round__n1786 ,
         _f_permutation__round__n1785 , _f_permutation__round__n1784 ,
         _f_permutation__round__n1783 , _f_permutation__round__n1782 ,
         _f_permutation__round__n1781 , _f_permutation__round__n1780 ,
         _f_permutation__round__n1779 , _f_permutation__round__n1778 ,
         _f_permutation__round__n1777 , _f_permutation__round__n1776 ,
         _f_permutation__round__n1775 , _f_permutation__round__n1774 ,
         _f_permutation__round__n1773 , _f_permutation__round__n1772 ,
         _f_permutation__round__n1771 , _f_permutation__round__n1770 ,
         _f_permutation__round__n1769 , _f_permutation__round__n1768 ,
         _f_permutation__round__n1767 , _f_permutation__round__n1766 ,
         _f_permutation__round__n1765 , _f_permutation__round__n1764 ,
         _f_permutation__round__n1763 , _f_permutation__round__n1762 ,
         _f_permutation__round__n1761 , _f_permutation__round__n1760 ,
         _f_permutation__round__n1759 , _f_permutation__round__n1758 ,
         _f_permutation__round__n1757 , _f_permutation__round__n1756 ,
         _f_permutation__round__n1755 , _f_permutation__round__n1754 ,
         _f_permutation__round__n1753 , _f_permutation__round__n1752 ,
         _f_permutation__round__n1751 , _f_permutation__round__n1750 ,
         _f_permutation__round__n1749 , _f_permutation__round__n1748 ,
         _f_permutation__round__n1747 , _f_permutation__round__n1746 ,
         _f_permutation__round__n1745 , _f_permutation__round__n1744 ,
         _f_permutation__round__n1743 , _f_permutation__round__n1742 ,
         _f_permutation__round__n1741 , _f_permutation__round__n1740 ,
         _f_permutation__round__n1739 , _f_permutation__round__n1738 ,
         _f_permutation__round__n1737 , _f_permutation__round__n1736 ,
         _f_permutation__round__n1735 , _f_permutation__round__n1734 ,
         _f_permutation__round__n1733 , _f_permutation__round__n1732 ,
         _f_permutation__round__n1731 , _f_permutation__round__n1730 ,
         _f_permutation__round__n1729 , _f_permutation__round__n1728 ,
         _f_permutation__round__n1727 , _f_permutation__round__n1726 ,
         _f_permutation__round__n1725 , _f_permutation__round__n1724 ,
         _f_permutation__round__n1723 , _f_permutation__round__n1722 ,
         _f_permutation__round__n1721 , _f_permutation__round__n1720 ,
         _f_permutation__round__n1719 , _f_permutation__round__n1718 ,
         _f_permutation__round__n1717 , _f_permutation__round__n1716 ,
         _f_permutation__round__n1715 , _f_permutation__round__n1714 ,
         _f_permutation__round__n1713 , _f_permutation__round__n1712 ,
         _f_permutation__round__n1711 , _f_permutation__round__n1710 ,
         _f_permutation__round__n1709 , _f_permutation__round__n1708 ,
         _f_permutation__round__n1707 , _f_permutation__round__n1706 ,
         _f_permutation__round__n1705 , _f_permutation__round__n1704 ,
         _f_permutation__round__n1703 , _f_permutation__round__n1702 ,
         _f_permutation__round__n1701 , _f_permutation__round__n1700 ,
         _f_permutation__round__n1699 , _f_permutation__round__n1698 ,
         _f_permutation__round__n1697 , _f_permutation__round__n1696 ,
         _f_permutation__round__n1695 , _f_permutation__round__n1694 ,
         _f_permutation__round__n1693 , _f_permutation__round__n1692 ,
         _f_permutation__round__n1691 , _f_permutation__round__n1690 ,
         _f_permutation__round__n1689 , _f_permutation__round__n1688 ,
         _f_permutation__round__n1687 , _f_permutation__round__n1686 ,
         _f_permutation__round__n1685 , _f_permutation__round__n1684 ,
         _f_permutation__round__n1683 , _f_permutation__round__n1682 ,
         _f_permutation__round__n1681 , _f_permutation__round__n1680 ,
         _f_permutation__round__n1679 , _f_permutation__round__n1678 ,
         _f_permutation__round__n1677 , _f_permutation__round__n1676 ,
         _f_permutation__round__n1675 , _f_permutation__round__n1674 ,
         _f_permutation__round__n1673 , _f_permutation__round__n1672 ,
         _f_permutation__round__n1671 , _f_permutation__round__n1670 ,
         _f_permutation__round__n1669 , _f_permutation__round__n1668 ,
         _f_permutation__round__n1667 , _f_permutation__round__n1666 ,
         _f_permutation__round__n1665 , _f_permutation__round__n1664 ,
         _f_permutation__round__n1663 , _f_permutation__round__n1662 ,
         _f_permutation__round__n1661 , _f_permutation__round__n1660 ,
         _f_permutation__round__n1659 , _f_permutation__round__n1658 ,
         _f_permutation__round__n1657 , _f_permutation__round__n1656 ,
         _f_permutation__round__n1655 , _f_permutation__round__n1654 ,
         _f_permutation__round__n1653 , _f_permutation__round__n1652 ,
         _f_permutation__round__n1651 , _f_permutation__round__n1650 ,
         _f_permutation__round__n1649 , _f_permutation__round__n1648 ,
         _f_permutation__round__n1647 , _f_permutation__round__n1646 ,
         _f_permutation__round__n1645 , _f_permutation__round__n1644 ,
         _f_permutation__round__n1643 , _f_permutation__round__n1642 ,
         _f_permutation__round__n1641 , _f_permutation__round__n1640 ,
         _f_permutation__round__n1639 , _f_permutation__round__n1638 ,
         _f_permutation__round__n1637 , _f_permutation__round__n1636 ,
         _f_permutation__round__n1635 , _f_permutation__round__n1634 ,
         _f_permutation__round__n1633 , _f_permutation__round__n1632 ,
         _f_permutation__round__n1631 , _f_permutation__round__n1630 ,
         _f_permutation__round__n1629 , _f_permutation__round__n1628 ,
         _f_permutation__round__n1627 , _f_permutation__round__n1626 ,
         _f_permutation__round__n1625 , _f_permutation__round__n1624 ,
         _f_permutation__round__n1623 , _f_permutation__round__n1622 ,
         _f_permutation__round__n1621 , _f_permutation__round__n1620 ,
         _f_permutation__round__n1619 , _f_permutation__round__n1618 ,
         _f_permutation__round__n1617 , _f_permutation__round__n1616 ,
         _f_permutation__round__n1615 , _f_permutation__round__n1614 ,
         _f_permutation__round__n1613 , _f_permutation__round__n1612 ,
         _f_permutation__round__n1611 , _f_permutation__round__n1610 ,
         _f_permutation__round__n1609 , _f_permutation__round__n1608 ,
         _f_permutation__round__n1607 , _f_permutation__round__n1606 ,
         _f_permutation__round__n1605 , _f_permutation__round__n1604 ,
         _f_permutation__round__n1603 , _f_permutation__round__n1602 ,
         _f_permutation__round__n1601 , _f_permutation__round__n1600 ,
         _f_permutation__round__n1599 , _f_permutation__round__n1598 ,
         _f_permutation__round__n1597 , _f_permutation__round__n1596 ,
         _f_permutation__round__n1595 , _f_permutation__round__n1594 ,
         _f_permutation__round__n1593 , _f_permutation__round__n1592 ,
         _f_permutation__round__n1591 , _f_permutation__round__n1590 ,
         _f_permutation__round__n1589 , _f_permutation__round__n1588 ,
         _f_permutation__round__n1587 , _f_permutation__round__n1586 ,
         _f_permutation__round__n1585 , _f_permutation__round__n1584 ,
         _f_permutation__round__n1583 , _f_permutation__round__n1582 ,
         _f_permutation__round__n1581 , _f_permutation__round__n1580 ,
         _f_permutation__round__n1579 , _f_permutation__round__n1578 ,
         _f_permutation__round__n1577 , _f_permutation__round__n1576 ,
         _f_permutation__round__n1575 , _f_permutation__round__n1574 ,
         _f_permutation__round__n1573 , _f_permutation__round__n1572 ,
         _f_permutation__round__n1571 , _f_permutation__round__n1570 ,
         _f_permutation__round__n1569 , _f_permutation__round__n1568 ,
         _f_permutation__round__n1567 , _f_permutation__round__n1566 ,
         _f_permutation__round__n1565 , _f_permutation__round__n1564 ,
         _f_permutation__round__n1563 , _f_permutation__round__n1562 ,
         _f_permutation__round__n1561 , _f_permutation__round__n1560 ,
         _f_permutation__round__n1559 , _f_permutation__round__n1558 ,
         _f_permutation__round__n1557 , _f_permutation__round__n1556 ,
         _f_permutation__round__n1555 , _f_permutation__round__n1554 ,
         _f_permutation__round__n1553 , _f_permutation__round__n1552 ,
         _f_permutation__round__n1551 , _f_permutation__round__n1550 ,
         _f_permutation__round__n1549 , _f_permutation__round__n1548 ,
         _f_permutation__round__n1547 , _f_permutation__round__n1546 ,
         _f_permutation__round__n1545 , _f_permutation__round__n1544 ,
         _f_permutation__round__n1543 , _f_permutation__round__n1542 ,
         _f_permutation__round__n1541 , _f_permutation__round__n1540 ,
         _f_permutation__round__n1539 , _f_permutation__round__n1538 ,
         _f_permutation__round__n1537 , _f_permutation__round__n1536 ,
         _f_permutation__round__n1535 , _f_permutation__round__n1534 ,
         _f_permutation__round__n1533 , _f_permutation__round__n1532 ,
         _f_permutation__round__n1531 , _f_permutation__round__n1530 ,
         _f_permutation__round__n1529 , _f_permutation__round__n1528 ,
         _f_permutation__round__n1527 , _f_permutation__round__n1526 ,
         _f_permutation__round__n1525 , _f_permutation__round__n1524 ,
         _f_permutation__round__n1523 , _f_permutation__round__n1522 ,
         _f_permutation__round__n1521 , _f_permutation__round__n1520 ,
         _f_permutation__round__n1519 , _f_permutation__round__n1518 ,
         _f_permutation__round__n1517 , _f_permutation__round__n1516 ,
         _f_permutation__round__n1515 , _f_permutation__round__n1514 ,
         _f_permutation__round__n1513 , _f_permutation__round__n1512 ,
         _f_permutation__round__n1511 , _f_permutation__round__n1510 ,
         _f_permutation__round__n1509 , _f_permutation__round__n1508 ,
         _f_permutation__round__n1507 , _f_permutation__round__n1506 ,
         _f_permutation__round__n1505 , _f_permutation__round__n1504 ,
         _f_permutation__round__n1503 , _f_permutation__round__n1502 ,
         _f_permutation__round__n1501 , _f_permutation__round__n1500 ,
         _f_permutation__round__n1499 , _f_permutation__round__n1498 ,
         _f_permutation__round__n1497 , _f_permutation__round__n1496 ,
         _f_permutation__round__n1495 , _f_permutation__round__n1494 ,
         _f_permutation__round__n1493 , _f_permutation__round__n1492 ,
         _f_permutation__round__n1491 , _f_permutation__round__n1490 ,
         _f_permutation__round__n1489 , _f_permutation__round__n1488 ,
         _f_permutation__round__n1487 , _f_permutation__round__n1486 ,
         _f_permutation__round__n1485 , _f_permutation__round__n1484 ,
         _f_permutation__round__n1483 , _f_permutation__round__n1482 ,
         _f_permutation__round__n1481 , _f_permutation__round__n1480 ,
         _f_permutation__round__n1479 , _f_permutation__round__n1478 ,
         _f_permutation__round__n1477 , _f_permutation__round__n1476 ,
         _f_permutation__round__n1475 , _f_permutation__round__n1474 ,
         _f_permutation__round__n1473 , _f_permutation__round__n1472 ,
         _f_permutation__round__n1471 , _f_permutation__round__n1470 ,
         _f_permutation__round__n1469 , _f_permutation__round__n1468 ,
         _f_permutation__round__n1467 , _f_permutation__round__n1466 ,
         _f_permutation__round__n1465 , _f_permutation__round__n1464 ,
         _f_permutation__round__n1463 , _f_permutation__round__n1462 ,
         _f_permutation__round__n1461 , _f_permutation__round__n1460 ,
         _f_permutation__round__n1459 , _f_permutation__round__n1458 ,
         _f_permutation__round__n1457 , _f_permutation__round__n1456 ,
         _f_permutation__round__n1455 , _f_permutation__round__n1454 ,
         _f_permutation__round__n1453 , _f_permutation__round__n1452 ,
         _f_permutation__round__n1451 , _f_permutation__round__n1450 ,
         _f_permutation__round__n1449 , _f_permutation__round__n1448 ,
         _f_permutation__round__n1447 , _f_permutation__round__n1446 ,
         _f_permutation__round__n1445 , _f_permutation__round__n1444 ,
         _f_permutation__round__n1443 , _f_permutation__round__n1442 ,
         _f_permutation__round__n1441 , _f_permutation__round__n1440 ,
         _f_permutation__round__n1439 , _f_permutation__round__n1438 ,
         _f_permutation__round__n1437 , _f_permutation__round__n1436 ,
         _f_permutation__round__n1435 , _f_permutation__round__n1434 ,
         _f_permutation__round__n1433 , _f_permutation__round__n1432 ,
         _f_permutation__round__n1431 , _f_permutation__round__n1430 ,
         _f_permutation__round__n1429 , _f_permutation__round__n1428 ,
         _f_permutation__round__n1427 , _f_permutation__round__n1426 ,
         _f_permutation__round__n1425 , _f_permutation__round__n1424 ,
         _f_permutation__round__n1423 , _f_permutation__round__n1422 ,
         _f_permutation__round__n1421 , _f_permutation__round__n1420 ,
         _f_permutation__round__n1419 , _f_permutation__round__n1418 ,
         _f_permutation__round__n1417 , _f_permutation__round__n1416 ,
         _f_permutation__round__n1415 , _f_permutation__round__n1414 ,
         _f_permutation__round__n1413 , _f_permutation__round__n1412 ,
         _f_permutation__round__n1411 , _f_permutation__round__n1410 ,
         _f_permutation__round__n1409 , _f_permutation__round__n1408 ,
         _f_permutation__round__n1407 , _f_permutation__round__n1406 ,
         _f_permutation__round__n1405 , _f_permutation__round__n1404 ,
         _f_permutation__round__n1403 , _f_permutation__round__n1402 ,
         _f_permutation__round__n1401 , _f_permutation__round__n1400 ,
         _f_permutation__round__n1399 , _f_permutation__round__n1398 ,
         _f_permutation__round__n1397 , _f_permutation__round__n1396 ,
         _f_permutation__round__n1395 , _f_permutation__round__n1394 ,
         _f_permutation__round__n1393 , _f_permutation__round__n1392 ,
         _f_permutation__round__n1391 , _f_permutation__round__n1390 ,
         _f_permutation__round__n1389 , _f_permutation__round__n1388 ,
         _f_permutation__round__n1387 , _f_permutation__round__n1386 ,
         _f_permutation__round__n1385 , _f_permutation__round__n1384 ,
         _f_permutation__round__n1383 , _f_permutation__round__n1382 ,
         _f_permutation__round__n1381 , _f_permutation__round__n1380 ,
         _f_permutation__round__n1379 , _f_permutation__round__n1378 ,
         _f_permutation__round__n1377 , _f_permutation__round__n1376 ,
         _f_permutation__round__n1375 , _f_permutation__round__n1374 ,
         _f_permutation__round__n1373 , _f_permutation__round__n1372 ,
         _f_permutation__round__n1371 , _f_permutation__round__n1370 ,
         _f_permutation__round__n1369 , _f_permutation__round__n1368 ,
         _f_permutation__round__n1367 , _f_permutation__round__n1366 ,
         _f_permutation__round__n1365 , _f_permutation__round__n1364 ,
         _f_permutation__round__n1363 , _f_permutation__round__n1362 ,
         _f_permutation__round__n1361 , _f_permutation__round__n1360 ,
         _f_permutation__round__n1359 , _f_permutation__round__n1358 ,
         _f_permutation__round__n1357 , _f_permutation__round__n1356 ,
         _f_permutation__round__n1355 , _f_permutation__round__n1354 ,
         _f_permutation__round__n1353 , _f_permutation__round__n1352 ,
         _f_permutation__round__n1351 , _f_permutation__round__n1350 ,
         _f_permutation__round__n1349 , _f_permutation__round__n1348 ,
         _f_permutation__round__n1347 , _f_permutation__round__n1346 ,
         _f_permutation__round__n1345 , _f_permutation__round__n1344 ,
         _f_permutation__round__n1343 , _f_permutation__round__n1342 ,
         _f_permutation__round__n1341 , _f_permutation__round__n1340 ,
         _f_permutation__round__n1339 , _f_permutation__round__n1338 ,
         _f_permutation__round__n1337 , _f_permutation__round__n1336 ,
         _f_permutation__round__n1335 , _f_permutation__round__n1334 ,
         _f_permutation__round__n1333 , _f_permutation__round__n1332 ,
         _f_permutation__round__n1331 , _f_permutation__round__n1330 ,
         _f_permutation__round__n1329 , _f_permutation__round__n1328 ,
         _f_permutation__round__n1327 , _f_permutation__round__n1326 ,
         _f_permutation__round__n1325 , _f_permutation__round__n1324 ,
         _f_permutation__round__n1323 , _f_permutation__round__n1322 ,
         _f_permutation__round__n1321 , _f_permutation__round__n1320 ,
         _f_permutation__round__n1319 , _f_permutation__round__n1318 ,
         _f_permutation__round__n1317 , _f_permutation__round__n1316 ,
         _f_permutation__round__n1315 , _f_permutation__round__n1314 ,
         _f_permutation__round__n1313 , _f_permutation__round__n1312 ,
         _f_permutation__round__n1311 , _f_permutation__round__n1310 ,
         _f_permutation__round__n1309 , _f_permutation__round__n1308 ,
         _f_permutation__round__n1307 , _f_permutation__round__n1306 ,
         _f_permutation__round__n1305 , _f_permutation__round__n1304 ,
         _f_permutation__round__n1303 , _f_permutation__round__n1302 ,
         _f_permutation__round__n1301 , _f_permutation__round__n1300 ,
         _f_permutation__round__n1299 , _f_permutation__round__n1298 ,
         _f_permutation__round__n1297 , _f_permutation__round__n1296 ,
         _f_permutation__round__n1295 , _f_permutation__round__n1294 ,
         _f_permutation__round__n1293 , _f_permutation__round__n1292 ,
         _f_permutation__round__n1291 , _f_permutation__round__n1290 ,
         _f_permutation__round__n1289 , _f_permutation__round__n1288 ,
         _f_permutation__round__n1287 , _f_permutation__round__n1286 ,
         _f_permutation__round__n1285 , _f_permutation__round__n1284 ,
         _f_permutation__round__n1283 , _f_permutation__round__n1282 ,
         _f_permutation__round__n1281 , _f_permutation__round__n1280 ,
         _f_permutation__round__n1279 , _f_permutation__round__n1278 ,
         _f_permutation__round__n1277 , _f_permutation__round__n1276 ,
         _f_permutation__round__n1275 , _f_permutation__round__n1274 ,
         _f_permutation__round__n1273 , _f_permutation__round__n1272 ,
         _f_permutation__round__n1271 , _f_permutation__round__n1270 ,
         _f_permutation__round__n1269 , _f_permutation__round__n1268 ,
         _f_permutation__round__n1267 , _f_permutation__round__n1266 ,
         _f_permutation__round__n1265 , _f_permutation__round__n1264 ,
         _f_permutation__round__n1263 , _f_permutation__round__n1262 ,
         _f_permutation__round__n1261 , _f_permutation__round__n1260 ,
         _f_permutation__round__n1259 , _f_permutation__round__n1258 ,
         _f_permutation__round__n1257 , _f_permutation__round__n1256 ,
         _f_permutation__round__n1255 , _f_permutation__round__n1254 ,
         _f_permutation__round__n1253 , _f_permutation__round__n1252 ,
         _f_permutation__round__n1251 , _f_permutation__round__n1250 ,
         _f_permutation__round__n1249 , _f_permutation__round__n1248 ,
         _f_permutation__round__n1247 , _f_permutation__round__n1246 ,
         _f_permutation__round__n1245 , _f_permutation__round__n1244 ,
         _f_permutation__round__n1243 , _f_permutation__round__n1242 ,
         _f_permutation__round__n1241 , _f_permutation__round__n1240 ,
         _f_permutation__round__n1239 , _f_permutation__round__n1238 ,
         _f_permutation__round__n1237 , _f_permutation__round__n1236 ,
         _f_permutation__round__n1235 , _f_permutation__round__n1234 ,
         _f_permutation__round__n1233 , _f_permutation__round__n1232 ,
         _f_permutation__round__n1231 , _f_permutation__round__n1230 ,
         _f_permutation__round__n1229 , _f_permutation__round__n1228 ,
         _f_permutation__round__n1227 , _f_permutation__round__n1226 ,
         _f_permutation__round__n1225 , _f_permutation__round__n1224 ,
         _f_permutation__round__n1223 , _f_permutation__round__n1222 ,
         _f_permutation__round__n1221 , _f_permutation__round__n1220 ,
         _f_permutation__round__n1219 , _f_permutation__round__n1218 ,
         _f_permutation__round__n1217 , _f_permutation__round__n1216 ,
         _f_permutation__round__n1215 , _f_permutation__round__n1214 ,
         _f_permutation__round__n1213 , _f_permutation__round__n1212 ,
         _f_permutation__round__n1211 , _f_permutation__round__n1210 ,
         _f_permutation__round__n1209 , _f_permutation__round__n1208 ,
         _f_permutation__round__n1207 , _f_permutation__round__n1206 ,
         _f_permutation__round__n1205 , _f_permutation__round__n1204 ,
         _f_permutation__round__n1203 , _f_permutation__round__n1202 ,
         _f_permutation__round__n1201 , _f_permutation__round__n1200 ,
         _f_permutation__round__n1199 , _f_permutation__round__n1198 ,
         _f_permutation__round__n1197 , _f_permutation__round__n1196 ,
         _f_permutation__round__n1195 , _f_permutation__round__n1194 ,
         _f_permutation__round__n1193 , _f_permutation__round__n1192 ,
         _f_permutation__round__n1191 , _f_permutation__round__n1190 ,
         _f_permutation__round__n1189 , _f_permutation__round__n1188 ,
         _f_permutation__round__n1187 , _f_permutation__round__n1186 ,
         _f_permutation__round__n1185 , _f_permutation__round__n1184 ,
         _f_permutation__round__n1183 , _f_permutation__round__n1182 ,
         _f_permutation__round__n1181 , _f_permutation__round__n1180 ,
         _f_permutation__round__n1179 , _f_permutation__round__n1178 ,
         _f_permutation__round__n1177 , _f_permutation__round__n1176 ,
         _f_permutation__round__n1175 , _f_permutation__round__n1174 ,
         _f_permutation__round__n1173 , _f_permutation__round__n1172 ,
         _f_permutation__round__n1171 , _f_permutation__round__n1170 ,
         _f_permutation__round__n1169 , _f_permutation__round__n1168 ,
         _f_permutation__round__n1167 , _f_permutation__round__n1166 ,
         _f_permutation__round__n1165 , _f_permutation__round__n1164 ,
         _f_permutation__round__n1163 , _f_permutation__round__n1162 ,
         _f_permutation__round__n1161 , _f_permutation__round__n1160 ,
         _f_permutation__round__n1159 , _f_permutation__round__n1158 ,
         _f_permutation__round__n1157 , _f_permutation__round__n1156 ,
         _f_permutation__round__n1155 , _f_permutation__round__n1154 ,
         _f_permutation__round__n1153 , _f_permutation__round__n1152 ,
         _f_permutation__round__n1151 , _f_permutation__round__n1150 ,
         _f_permutation__round__n1149 , _f_permutation__round__n1148 ,
         _f_permutation__round__n1147 , _f_permutation__round__n1146 ,
         _f_permutation__round__n1145 , _f_permutation__round__n1144 ,
         _f_permutation__round__n1143 , _f_permutation__round__n1142 ,
         _f_permutation__round__n1141 , _f_permutation__round__n1140 ,
         _f_permutation__round__n1139 , _f_permutation__round__n1138 ,
         _f_permutation__round__n1137 , _f_permutation__round__n1136 ,
         _f_permutation__round__n1135 , _f_permutation__round__n1134 ,
         _f_permutation__round__n1133 , _f_permutation__round__n1132 ,
         _f_permutation__round__n1131 , _f_permutation__round__n1130 ,
         _f_permutation__round__n1129 , _f_permutation__round__n1128 ,
         _f_permutation__round__n1127 , _f_permutation__round__n1126 ,
         _f_permutation__round__n1125 , _f_permutation__round__n1124 ,
         _f_permutation__round__n1123 , _f_permutation__round__n1122 ,
         _f_permutation__round__n1121 , _f_permutation__round__n1120 ,
         _f_permutation__round__n1119 , _f_permutation__round__n1118 ,
         _f_permutation__round__n1117 , _f_permutation__round__n1116 ,
         _f_permutation__round__n1115 , _f_permutation__round__n1114 ,
         _f_permutation__round__n1113 , _f_permutation__round__n1112 ,
         _f_permutation__round__n1111 , _f_permutation__round__n1110 ,
         _f_permutation__round__n1109 , _f_permutation__round__n1108 ,
         _f_permutation__round__n1107 , _f_permutation__round__n1106 ,
         _f_permutation__round__n1105 , _f_permutation__round__n1104 ,
         _f_permutation__round__n1103 , _f_permutation__round__n1102 ,
         _f_permutation__round__n1101 , _f_permutation__round__n1100 ,
         _f_permutation__round__n1099 , _f_permutation__round__n1098 ,
         _f_permutation__round__n1097 , _f_permutation__round__n1096 ,
         _f_permutation__round__n1095 , _f_permutation__round__n1094 ,
         _f_permutation__round__n1093 , _f_permutation__round__n1092 ,
         _f_permutation__round__n1091 , _f_permutation__round__n1090 ,
         _f_permutation__round__n1089 , _f_permutation__round__n1088 ,
         _f_permutation__round__n1087 , _f_permutation__round__n1086 ,
         _f_permutation__round__n1085 , _f_permutation__round__n1084 ,
         _f_permutation__round__n1083 , _f_permutation__round__n1082 ,
         _f_permutation__round__n1081 , _f_permutation__round__n1080 ,
         _f_permutation__round__n1079 , _f_permutation__round__n1078 ,
         _f_permutation__round__n1077 , _f_permutation__round__n1076 ,
         _f_permutation__round__n1075 , _f_permutation__round__n1074 ,
         _f_permutation__round__n1073 , _f_permutation__round__n1072 ,
         _f_permutation__round__n1071 , _f_permutation__round__n1070 ,
         _f_permutation__round__n1069 , _f_permutation__round__n1068 ,
         _f_permutation__round__n1067 , _f_permutation__round__n1066 ,
         _f_permutation__round__n1065 , _f_permutation__round__n1064 ,
         _f_permutation__round__n1063 , _f_permutation__round__n1062 ,
         _f_permutation__round__n1061 , _f_permutation__round__n1060 ,
         _f_permutation__round__n1059 , _f_permutation__round__n1058 ,
         _f_permutation__round__n1057 , _f_permutation__round__n1056 ,
         _f_permutation__round__n1055 , _f_permutation__round__n1054 ,
         _f_permutation__round__n1053 , _f_permutation__round__n1052 ,
         _f_permutation__round__n1051 , _f_permutation__round__n1050 ,
         _f_permutation__round__n1049 , _f_permutation__round__n1048 ,
         _f_permutation__round__n1047 , _f_permutation__round__n1046 ,
         _f_permutation__round__n1045 , _f_permutation__round__n1044 ,
         _f_permutation__round__n1043 , _f_permutation__round__n1042 ,
         _f_permutation__round__n1041 , _f_permutation__round__n1040 ,
         _f_permutation__round__n1039 , _f_permutation__round__n1038 ,
         _f_permutation__round__n1037 , _f_permutation__round__n1036 ,
         _f_permutation__round__n1035 , _f_permutation__round__n1034 ,
         _f_permutation__round__n1033 , _f_permutation__round__n1032 ,
         _f_permutation__round__n1031 , _f_permutation__round__n1030 ,
         _f_permutation__round__n1029 , _f_permutation__round__n1028 ,
         _f_permutation__round__n1027 , _f_permutation__round__n1026 ,
         _f_permutation__round__n1025 , _f_permutation__round__n1024 ,
         _f_permutation__round__n1023 , _f_permutation__round__n1022 ,
         _f_permutation__round__n1021 , _f_permutation__round__n1020 ,
         _f_permutation__round__n1019 , _f_permutation__round__n1018 ,
         _f_permutation__round__n1017 , _f_permutation__round__n1016 ,
         _f_permutation__round__n1015 , _f_permutation__round__n1014 ,
         _f_permutation__round__n1013 , _f_permutation__round__n1012 ,
         _f_permutation__round__n1011 , _f_permutation__round__n1010 ,
         _f_permutation__round__n1009 , _f_permutation__round__n1008 ,
         _f_permutation__round__n1007 , _f_permutation__round__n1006 ,
         _f_permutation__round__n1005 , _f_permutation__round__n1004 ,
         _f_permutation__round__n1003 , _f_permutation__round__n1002 ,
         _f_permutation__round__n1001 , _f_permutation__round__n1000 ,
         _f_permutation__round__n999 , _f_permutation__round__n998 ,
         _f_permutation__round__n997 , _f_permutation__round__n996 ,
         _f_permutation__round__n995 , _f_permutation__round__n994 ,
         _f_permutation__round__n993 , _f_permutation__round__n992 ,
         _f_permutation__round__n991 , _f_permutation__round__n990 ,
         _f_permutation__round__n989 , _f_permutation__round__n988 ,
         _f_permutation__round__n987 , _f_permutation__round__n986 ,
         _f_permutation__round__n985 , _f_permutation__round__n984 ,
         _f_permutation__round__n983 , _f_permutation__round__n982 ,
         _f_permutation__round__n981 , _f_permutation__round__n980 ,
         _f_permutation__round__n979 , _f_permutation__round__n978 ,
         _f_permutation__round__n977 , _f_permutation__round__n976 ,
         _f_permutation__round__n975 , _f_permutation__round__n974 ,
         _f_permutation__round__n973 , _f_permutation__round__n972 ,
         _f_permutation__round__n971 , _f_permutation__round__n970 ,
         _f_permutation__round__n969 , _f_permutation__round__n968 ,
         _f_permutation__round__n967 , _f_permutation__round__n966 ,
         _f_permutation__round__n965 , _f_permutation__round__n964 ,
         _f_permutation__round__n963 , _f_permutation__round__n962 ,
         _f_permutation__round__n961 , _f_permutation__round__N5759 ,
         _f_permutation__round__N5757 , _f_permutation__round__N5755 ,
         _f_permutation__round__N5753 , _f_permutation__round__N5751 ,
         _f_permutation__round__N5749 , _f_permutation__round__N5747 ,
         _f_permutation__round__N5745 , _f_permutation__round__N5743 ,
         _f_permutation__round__N5741 , _f_permutation__round__N5739 ,
         _f_permutation__round__N5737 , _f_permutation__round__N5735 ,
         _f_permutation__round__N5733 , _f_permutation__round__N5731 ,
         _f_permutation__round__N5729 , _f_permutation__round__N5727 ,
         _f_permutation__round__N5725 , _f_permutation__round__N5723 ,
         _f_permutation__round__N5721 , _f_permutation__round__N5719 ,
         _f_permutation__round__N5717 , _f_permutation__round__N5715 ,
         _f_permutation__round__N5713 , _f_permutation__round__N5711 ,
         _f_permutation__round__N5709 , _f_permutation__round__N5707 ,
         _f_permutation__round__N5705 , _f_permutation__round__N5703 ,
         _f_permutation__round__N5701 , _f_permutation__round__N5699 ,
         _f_permutation__round__N5697 , _f_permutation__round__N5695 ,
         _f_permutation__round__N5693 , _f_permutation__round__N5691 ,
         _f_permutation__round__N5689 , _f_permutation__round__N5687 ,
         _f_permutation__round__N5685 , _f_permutation__round__N5683 ,
         _f_permutation__round__N5681 , _f_permutation__round__N5679 ,
         _f_permutation__round__N5677 , _f_permutation__round__N5675 ,
         _f_permutation__round__N5673 , _f_permutation__round__N5671 ,
         _f_permutation__round__N5669 , _f_permutation__round__N5667 ,
         _f_permutation__round__N5665 , _f_permutation__round__N5663 ,
         _f_permutation__round__N5661 , _f_permutation__round__N5659 ,
         _f_permutation__round__N5657 , _f_permutation__round__N5655 ,
         _f_permutation__round__N5653 , _f_permutation__round__N5651 ,
         _f_permutation__round__N5649 , _f_permutation__round__N5647 ,
         _f_permutation__round__N5645 , _f_permutation__round__N5643 ,
         _f_permutation__round__N5641 , _f_permutation__round__N5639 ,
         _f_permutation__round__N5637 , _f_permutation__round__N5635 ,
         _f_permutation__round__N5633 , _f_permutation__round__N5631 ,
         _f_permutation__round__N5629 , _f_permutation__round__N5627 ,
         _f_permutation__round__N5625 , _f_permutation__round__N5623 ,
         _f_permutation__round__N5621 , _f_permutation__round__N5619 ,
         _f_permutation__round__N5617 , _f_permutation__round__N5615 ,
         _f_permutation__round__N5613 , _f_permutation__round__N5611 ,
         _f_permutation__round__N5609 , _f_permutation__round__N5607 ,
         _f_permutation__round__N5605 , _f_permutation__round__N5603 ,
         _f_permutation__round__N5601 , _f_permutation__round__N5599 ,
         _f_permutation__round__N5597 , _f_permutation__round__N5595 ,
         _f_permutation__round__N5593 , _f_permutation__round__N5591 ,
         _f_permutation__round__N5589 , _f_permutation__round__N5587 ,
         _f_permutation__round__N5585 , _f_permutation__round__N5583 ,
         _f_permutation__round__N5581 , _f_permutation__round__N5579 ,
         _f_permutation__round__N5577 , _f_permutation__round__N5575 ,
         _f_permutation__round__N5573 , _f_permutation__round__N5571 ,
         _f_permutation__round__N5569 , _f_permutation__round__N5567 ,
         _f_permutation__round__N5565 , _f_permutation__round__N5563 ,
         _f_permutation__round__N5561 , _f_permutation__round__N5559 ,
         _f_permutation__round__N5557 , _f_permutation__round__N5555 ,
         _f_permutation__round__N5553 , _f_permutation__round__N5551 ,
         _f_permutation__round__N5549 , _f_permutation__round__N5547 ,
         _f_permutation__round__N5545 , _f_permutation__round__N5543 ,
         _f_permutation__round__N5541 , _f_permutation__round__N5539 ,
         _f_permutation__round__N5537 , _f_permutation__round__N5535 ,
         _f_permutation__round__N5533 , _f_permutation__round__N5531 ,
         _f_permutation__round__N5529 , _f_permutation__round__N5527 ,
         _f_permutation__round__N5525 , _f_permutation__round__N5523 ,
         _f_permutation__round__N5521 , _f_permutation__round__N5519 ,
         _f_permutation__round__N5517 , _f_permutation__round__N5515 ,
         _f_permutation__round__N5513 , _f_permutation__round__N5511 ,
         _f_permutation__round__N5509 , _f_permutation__round__N5507 ,
         _f_permutation__round__N5505 , _f_permutation__round__N5503 ,
         _f_permutation__round__N5501 , _f_permutation__round__N5499 ,
         _f_permutation__round__N5497 , _f_permutation__round__N5495 ,
         _f_permutation__round__N5493 , _f_permutation__round__N5491 ,
         _f_permutation__round__N5489 , _f_permutation__round__N5487 ,
         _f_permutation__round__N5485 , _f_permutation__round__N5483 ,
         _f_permutation__round__N5481 , _f_permutation__round__N5479 ,
         _f_permutation__round__N5477 , _f_permutation__round__N5475 ,
         _f_permutation__round__N5473 , _f_permutation__round__N5471 ,
         _f_permutation__round__N5469 , _f_permutation__round__N5467 ,
         _f_permutation__round__N5465 , _f_permutation__round__N5463 ,
         _f_permutation__round__N5461 , _f_permutation__round__N5459 ,
         _f_permutation__round__N5457 , _f_permutation__round__N5455 ,
         _f_permutation__round__N5453 , _f_permutation__round__N5451 ,
         _f_permutation__round__N5449 , _f_permutation__round__N5447 ,
         _f_permutation__round__N5445 , _f_permutation__round__N5443 ,
         _f_permutation__round__N5441 , _f_permutation__round__N5439 ,
         _f_permutation__round__N5437 , _f_permutation__round__N5435 ,
         _f_permutation__round__N5433 , _f_permutation__round__N5431 ,
         _f_permutation__round__N5429 , _f_permutation__round__N5427 ,
         _f_permutation__round__N5425 , _f_permutation__round__N5423 ,
         _f_permutation__round__N5421 , _f_permutation__round__N5419 ,
         _f_permutation__round__N5417 , _f_permutation__round__N5415 ,
         _f_permutation__round__N5413 , _f_permutation__round__N5411 ,
         _f_permutation__round__N5409 , _f_permutation__round__N5407 ,
         _f_permutation__round__N5405 , _f_permutation__round__N5403 ,
         _f_permutation__round__N5401 , _f_permutation__round__N5399 ,
         _f_permutation__round__N5397 , _f_permutation__round__N5395 ,
         _f_permutation__round__N5393 , _f_permutation__round__N5391 ,
         _f_permutation__round__N5389 , _f_permutation__round__N5387 ,
         _f_permutation__round__N5385 , _f_permutation__round__N5383 ,
         _f_permutation__round__N5381 , _f_permutation__round__N5379 ,
         _f_permutation__round__N5377 , _f_permutation__round__N5375 ,
         _f_permutation__round__N5373 , _f_permutation__round__N5371 ,
         _f_permutation__round__N5369 , _f_permutation__round__N5367 ,
         _f_permutation__round__N5365 , _f_permutation__round__N5363 ,
         _f_permutation__round__N5361 , _f_permutation__round__N5359 ,
         _f_permutation__round__N5357 , _f_permutation__round__N5355 ,
         _f_permutation__round__N5353 , _f_permutation__round__N5351 ,
         _f_permutation__round__N5349 , _f_permutation__round__N5347 ,
         _f_permutation__round__N5345 , _f_permutation__round__N5343 ,
         _f_permutation__round__N5341 , _f_permutation__round__N5339 ,
         _f_permutation__round__N5337 , _f_permutation__round__N5335 ,
         _f_permutation__round__N5333 , _f_permutation__round__N5331 ,
         _f_permutation__round__N5329 , _f_permutation__round__N5327 ,
         _f_permutation__round__N5325 , _f_permutation__round__N5323 ,
         _f_permutation__round__N5321 , _f_permutation__round__N5319 ,
         _f_permutation__round__N5317 , _f_permutation__round__N5315 ,
         _f_permutation__round__N5313 , _f_permutation__round__N5311 ,
         _f_permutation__round__N5309 , _f_permutation__round__N5307 ,
         _f_permutation__round__N5305 , _f_permutation__round__N5303 ,
         _f_permutation__round__N5301 , _f_permutation__round__N5299 ,
         _f_permutation__round__N5297 , _f_permutation__round__N5295 ,
         _f_permutation__round__N5293 , _f_permutation__round__N5291 ,
         _f_permutation__round__N5289 , _f_permutation__round__N5287 ,
         _f_permutation__round__N5285 , _f_permutation__round__N5283 ,
         _f_permutation__round__N5281 , _f_permutation__round__N5279 ,
         _f_permutation__round__N5277 , _f_permutation__round__N5275 ,
         _f_permutation__round__N5273 , _f_permutation__round__N5271 ,
         _f_permutation__round__N5269 , _f_permutation__round__N5267 ,
         _f_permutation__round__N5265 , _f_permutation__round__N5263 ,
         _f_permutation__round__N5261 , _f_permutation__round__N5259 ,
         _f_permutation__round__N5257 , _f_permutation__round__N5255 ,
         _f_permutation__round__N5253 , _f_permutation__round__N5251 ,
         _f_permutation__round__N5249 , _f_permutation__round__N5247 ,
         _f_permutation__round__N5245 , _f_permutation__round__N5243 ,
         _f_permutation__round__N5241 , _f_permutation__round__N5239 ,
         _f_permutation__round__N5237 , _f_permutation__round__N5235 ,
         _f_permutation__round__N5233 , _f_permutation__round__N5231 ,
         _f_permutation__round__N5229 , _f_permutation__round__N5227 ,
         _f_permutation__round__N5225 , _f_permutation__round__N5223 ,
         _f_permutation__round__N5221 , _f_permutation__round__N5219 ,
         _f_permutation__round__N5217 , _f_permutation__round__N5215 ,
         _f_permutation__round__N5213 , _f_permutation__round__N5211 ,
         _f_permutation__round__N5209 , _f_permutation__round__N5207 ,
         _f_permutation__round__N5205 , _f_permutation__round__N5203 ,
         _f_permutation__round__N5201 , _f_permutation__round__N5199 ,
         _f_permutation__round__N5197 , _f_permutation__round__N5195 ,
         _f_permutation__round__N5193 , _f_permutation__round__N5191 ,
         _f_permutation__round__N5189 , _f_permutation__round__N5187 ,
         _f_permutation__round__N5185 , _f_permutation__round__N5183 ,
         _f_permutation__round__N5181 , _f_permutation__round__N5179 ,
         _f_permutation__round__N5177 , _f_permutation__round__N5175 ,
         _f_permutation__round__N5173 , _f_permutation__round__N5171 ,
         _f_permutation__round__N5169 , _f_permutation__round__N5167 ,
         _f_permutation__round__N5165 , _f_permutation__round__N5163 ,
         _f_permutation__round__N5161 , _f_permutation__round__N5159 ,
         _f_permutation__round__N5157 , _f_permutation__round__N5155 ,
         _f_permutation__round__N5153 , _f_permutation__round__N5151 ,
         _f_permutation__round__N5149 , _f_permutation__round__N5147 ,
         _f_permutation__round__N5145 , _f_permutation__round__N5143 ,
         _f_permutation__round__N5141 , _f_permutation__round__N5139 ,
         _f_permutation__round__N5137 , _f_permutation__round__N5135 ,
         _f_permutation__round__N5133 , _f_permutation__round__N5131 ,
         _f_permutation__round__N5129 , _f_permutation__round__N5127 ,
         _f_permutation__round__N5125 , _f_permutation__round__N5123 ,
         _f_permutation__round__N5121 , _f_permutation__round__N5119 ,
         _f_permutation__round__N5117 , _f_permutation__round__N5115 ,
         _f_permutation__round__N5113 , _f_permutation__round__N5111 ,
         _f_permutation__round__N5109 , _f_permutation__round__N5107 ,
         _f_permutation__round__N5105 , _f_permutation__round__N5103 ,
         _f_permutation__round__N5101 , _f_permutation__round__N5099 ,
         _f_permutation__round__N5097 , _f_permutation__round__N5095 ,
         _f_permutation__round__N5093 , _f_permutation__round__N5091 ,
         _f_permutation__round__N5089 , _f_permutation__round__N5087 ,
         _f_permutation__round__N5085 , _f_permutation__round__N5083 ,
         _f_permutation__round__N5081 , _f_permutation__round__N5079 ,
         _f_permutation__round__N5077 , _f_permutation__round__N5075 ,
         _f_permutation__round__N5073 , _f_permutation__round__N5071 ,
         _f_permutation__round__N5069 , _f_permutation__round__N5067 ,
         _f_permutation__round__N5065 , _f_permutation__round__N5063 ,
         _f_permutation__round__N5061 , _f_permutation__round__N5059 ,
         _f_permutation__round__N5057 , _f_permutation__round__N5055 ,
         _f_permutation__round__N5053 , _f_permutation__round__N5051 ,
         _f_permutation__round__N5049 , _f_permutation__round__N5047 ,
         _f_permutation__round__N5045 , _f_permutation__round__N5043 ,
         _f_permutation__round__N5041 , _f_permutation__round__N5039 ,
         _f_permutation__round__N5037 , _f_permutation__round__N5035 ,
         _f_permutation__round__N5033 , _f_permutation__round__N5031 ,
         _f_permutation__round__N5029 , _f_permutation__round__N5027 ,
         _f_permutation__round__N5025 , _f_permutation__round__N5023 ,
         _f_permutation__round__N5021 , _f_permutation__round__N5019 ,
         _f_permutation__round__N5017 , _f_permutation__round__N5015 ,
         _f_permutation__round__N5013 , _f_permutation__round__N5011 ,
         _f_permutation__round__N5009 , _f_permutation__round__N5007 ,
         _f_permutation__round__N5005 , _f_permutation__round__N5003 ,
         _f_permutation__round__N5001 , _f_permutation__round__N4999 ,
         _f_permutation__round__N4997 , _f_permutation__round__N4995 ,
         _f_permutation__round__N4993 , _f_permutation__round__N4991 ,
         _f_permutation__round__N4989 , _f_permutation__round__N4987 ,
         _f_permutation__round__N4985 , _f_permutation__round__N4983 ,
         _f_permutation__round__N4981 , _f_permutation__round__N4979 ,
         _f_permutation__round__N4977 , _f_permutation__round__N4975 ,
         _f_permutation__round__N4973 , _f_permutation__round__N4971 ,
         _f_permutation__round__N4969 , _f_permutation__round__N4967 ,
         _f_permutation__round__N4965 , _f_permutation__round__N4963 ,
         _f_permutation__round__N4961 , _f_permutation__round__N4959 ,
         _f_permutation__round__N4957 , _f_permutation__round__N4955 ,
         _f_permutation__round__N4953 , _f_permutation__round__N4951 ,
         _f_permutation__round__N4949 , _f_permutation__round__N4947 ,
         _f_permutation__round__N4945 , _f_permutation__round__N4943 ,
         _f_permutation__round__N4941 , _f_permutation__round__N4939 ,
         _f_permutation__round__N4937 , _f_permutation__round__N4935 ,
         _f_permutation__round__N4933 , _f_permutation__round__N4931 ,
         _f_permutation__round__N4929 , _f_permutation__round__N4927 ,
         _f_permutation__round__N4925 , _f_permutation__round__N4923 ,
         _f_permutation__round__N4921 , _f_permutation__round__N4919 ,
         _f_permutation__round__N4917 , _f_permutation__round__N4915 ,
         _f_permutation__round__N4913 , _f_permutation__round__N4911 ,
         _f_permutation__round__N4909 , _f_permutation__round__N4907 ,
         _f_permutation__round__N4905 , _f_permutation__round__N4903 ,
         _f_permutation__round__N4901 , _f_permutation__round__N4899 ,
         _f_permutation__round__N4897 , _f_permutation__round__N4895 ,
         _f_permutation__round__N4893 , _f_permutation__round__N4891 ,
         _f_permutation__round__N4889 , _f_permutation__round__N4887 ,
         _f_permutation__round__N4885 , _f_permutation__round__N4883 ,
         _f_permutation__round__N4881 , _f_permutation__round__N4879 ,
         _f_permutation__round__N4877 , _f_permutation__round__N4875 ,
         _f_permutation__round__N4873 , _f_permutation__round__N4871 ,
         _f_permutation__round__N4869 , _f_permutation__round__N4867 ,
         _f_permutation__round__N4865 , _f_permutation__round__N4863 ,
         _f_permutation__round__N4861 , _f_permutation__round__N4859 ,
         _f_permutation__round__N4857 , _f_permutation__round__N4855 ,
         _f_permutation__round__N4853 , _f_permutation__round__N4851 ,
         _f_permutation__round__N4849 , _f_permutation__round__N4847 ,
         _f_permutation__round__N4845 , _f_permutation__round__N4843 ,
         _f_permutation__round__N4841 , _f_permutation__round__N4839 ,
         _f_permutation__round__N4837 , _f_permutation__round__N4835 ,
         _f_permutation__round__N4833 , _f_permutation__round__N4831 ,
         _f_permutation__round__N4829 , _f_permutation__round__N4827 ,
         _f_permutation__round__N4825 , _f_permutation__round__N4823 ,
         _f_permutation__round__N4821 , _f_permutation__round__N4819 ,
         _f_permutation__round__N4817 , _f_permutation__round__N4815 ,
         _f_permutation__round__N4813 , _f_permutation__round__N4811 ,
         _f_permutation__round__N4809 , _f_permutation__round__N4807 ,
         _f_permutation__round__N4805 , _f_permutation__round__N4803 ,
         _f_permutation__round__N4801 , _f_permutation__round__N4799 ,
         _f_permutation__round__N4797 , _f_permutation__round__N4795 ,
         _f_permutation__round__N4793 , _f_permutation__round__N4791 ,
         _f_permutation__round__N4789 , _f_permutation__round__N4787 ,
         _f_permutation__round__N4785 , _f_permutation__round__N4783 ,
         _f_permutation__round__N4781 , _f_permutation__round__N4779 ,
         _f_permutation__round__N4777 , _f_permutation__round__N4775 ,
         _f_permutation__round__N4773 , _f_permutation__round__N4771 ,
         _f_permutation__round__N4769 , _f_permutation__round__N4767 ,
         _f_permutation__round__N4765 , _f_permutation__round__N4763 ,
         _f_permutation__round__N4761 , _f_permutation__round__N4759 ,
         _f_permutation__round__N4757 , _f_permutation__round__N4755 ,
         _f_permutation__round__N4753 , _f_permutation__round__N4751 ,
         _f_permutation__round__N4749 , _f_permutation__round__N4747 ,
         _f_permutation__round__N4745 , _f_permutation__round__N4743 ,
         _f_permutation__round__N4741 , _f_permutation__round__N4739 ,
         _f_permutation__round__N4737 , _f_permutation__round__N4735 ,
         _f_permutation__round__N4733 , _f_permutation__round__N4731 ,
         _f_permutation__round__N4729 , _f_permutation__round__N4727 ,
         _f_permutation__round__N4725 , _f_permutation__round__N4723 ,
         _f_permutation__round__N4721 , _f_permutation__round__N4719 ,
         _f_permutation__round__N4717 , _f_permutation__round__N4715 ,
         _f_permutation__round__N4713 , _f_permutation__round__N4711 ,
         _f_permutation__round__N4709 , _f_permutation__round__N4707 ,
         _f_permutation__round__N4705 , _f_permutation__round__N4703 ,
         _f_permutation__round__N4701 , _f_permutation__round__N4699 ,
         _f_permutation__round__N4697 , _f_permutation__round__N4695 ,
         _f_permutation__round__N4693 , _f_permutation__round__N4691 ,
         _f_permutation__round__N4689 , _f_permutation__round__N4687 ,
         _f_permutation__round__N4685 , _f_permutation__round__N4683 ,
         _f_permutation__round__N4681 , _f_permutation__round__N4679 ,
         _f_permutation__round__N4677 , _f_permutation__round__N4675 ,
         _f_permutation__round__N4673 , _f_permutation__round__N4671 ,
         _f_permutation__round__N4669 , _f_permutation__round__N4667 ,
         _f_permutation__round__N4665 , _f_permutation__round__N4663 ,
         _f_permutation__round__N4661 , _f_permutation__round__N4659 ,
         _f_permutation__round__N4657 , _f_permutation__round__N4655 ,
         _f_permutation__round__N4653 , _f_permutation__round__N4651 ,
         _f_permutation__round__N4649 , _f_permutation__round__N4647 ,
         _f_permutation__round__N4645 , _f_permutation__round__N4643 ,
         _f_permutation__round__N4641 , _f_permutation__round__N4639 ,
         _f_permutation__round__N4637 , _f_permutation__round__N4635 ,
         _f_permutation__round__N4633 , _f_permutation__round__N4631 ,
         _f_permutation__round__N4629 , _f_permutation__round__N4627 ,
         _f_permutation__round__N4625 , _f_permutation__round__N4623 ,
         _f_permutation__round__N4621 , _f_permutation__round__N4619 ,
         _f_permutation__round__N4617 , _f_permutation__round__N4615 ,
         _f_permutation__round__N4613 , _f_permutation__round__N4611 ,
         _f_permutation__round__N4609 , _f_permutation__round__N4607 ,
         _f_permutation__round__N4605 , _f_permutation__round__N4603 ,
         _f_permutation__round__N4601 , _f_permutation__round__N4599 ,
         _f_permutation__round__N4597 , _f_permutation__round__N4595 ,
         _f_permutation__round__N4593 , _f_permutation__round__N4591 ,
         _f_permutation__round__N4589 , _f_permutation__round__N4587 ,
         _f_permutation__round__N4585 , _f_permutation__round__N4583 ,
         _f_permutation__round__N4581 , _f_permutation__round__N4579 ,
         _f_permutation__round__N4577 , _f_permutation__round__N4575 ,
         _f_permutation__round__N4573 , _f_permutation__round__N4571 ,
         _f_permutation__round__N4569 , _f_permutation__round__N4567 ,
         _f_permutation__round__N4565 , _f_permutation__round__N4563 ,
         _f_permutation__round__N4561 , _f_permutation__round__N4559 ,
         _f_permutation__round__N4557 , _f_permutation__round__N4555 ,
         _f_permutation__round__N4553 , _f_permutation__round__N4551 ,
         _f_permutation__round__N4549 , _f_permutation__round__N4547 ,
         _f_permutation__round__N4545 , _f_permutation__round__N4543 ,
         _f_permutation__round__N4541 , _f_permutation__round__N4539 ,
         _f_permutation__round__N4537 , _f_permutation__round__N4535 ,
         _f_permutation__round__N4533 , _f_permutation__round__N4531 ,
         _f_permutation__round__N4529 , _f_permutation__round__N4527 ,
         _f_permutation__round__N4525 , _f_permutation__round__N4523 ,
         _f_permutation__round__N4521 , _f_permutation__round__N4519 ,
         _f_permutation__round__N4517 , _f_permutation__round__N4515 ,
         _f_permutation__round__N4513 , _f_permutation__round__N4511 ,
         _f_permutation__round__N4509 , _f_permutation__round__N4507 ,
         _f_permutation__round__N4505 , _f_permutation__round__N4503 ,
         _f_permutation__round__N4501 , _f_permutation__round__N4499 ,
         _f_permutation__round__N4497 , _f_permutation__round__N4495 ,
         _f_permutation__round__N4493 , _f_permutation__round__N4491 ,
         _f_permutation__round__N4489 , _f_permutation__round__N4487 ,
         _f_permutation__round__N4485 , _f_permutation__round__N4483 ,
         _f_permutation__round__N4481 , _f_permutation__round__N4479 ,
         _f_permutation__round__N4477 , _f_permutation__round__N4475 ,
         _f_permutation__round__N4473 , _f_permutation__round__N4471 ,
         _f_permutation__round__N4469 , _f_permutation__round__N4467 ,
         _f_permutation__round__N4465 , _f_permutation__round__N4463 ,
         _f_permutation__round__N4461 , _f_permutation__round__N4459 ,
         _f_permutation__round__N4457 , _f_permutation__round__N4455 ,
         _f_permutation__round__N4453 , _f_permutation__round__N4451 ,
         _f_permutation__round__N4449 , _f_permutation__round__N4447 ,
         _f_permutation__round__N4445 , _f_permutation__round__N4443 ,
         _f_permutation__round__N4441 , _f_permutation__round__N4439 ,
         _f_permutation__round__N4437 , _f_permutation__round__N4435 ,
         _f_permutation__round__N4433 , _f_permutation__round__N4431 ,
         _f_permutation__round__N4429 , _f_permutation__round__N4427 ,
         _f_permutation__round__N4425 , _f_permutation__round__N4423 ,
         _f_permutation__round__N4421 , _f_permutation__round__N4419 ,
         _f_permutation__round__N4417 , _f_permutation__round__N4415 ,
         _f_permutation__round__N4413 , _f_permutation__round__N4411 ,
         _f_permutation__round__N4409 , _f_permutation__round__N4407 ,
         _f_permutation__round__N4405 , _f_permutation__round__N4403 ,
         _f_permutation__round__N4401 , _f_permutation__round__N4399 ,
         _f_permutation__round__N4397 , _f_permutation__round__N4395 ,
         _f_permutation__round__N4393 , _f_permutation__round__N4391 ,
         _f_permutation__round__N4389 , _f_permutation__round__N4387 ,
         _f_permutation__round__N4385 , _f_permutation__round__N4383 ,
         _f_permutation__round__N4381 , _f_permutation__round__N4379 ,
         _f_permutation__round__N4377 , _f_permutation__round__N4375 ,
         _f_permutation__round__N4373 , _f_permutation__round__N4371 ,
         _f_permutation__round__N4369 , _f_permutation__round__N4367 ,
         _f_permutation__round__N4365 , _f_permutation__round__N4363 ,
         _f_permutation__round__N4361 , _f_permutation__round__N4359 ,
         _f_permutation__round__N4357 , _f_permutation__round__N4355 ,
         _f_permutation__round__N4353 , _f_permutation__round__N4351 ,
         _f_permutation__round__N4349 , _f_permutation__round__N4347 ,
         _f_permutation__round__N4345 , _f_permutation__round__N4343 ,
         _f_permutation__round__N4341 , _f_permutation__round__N4339 ,
         _f_permutation__round__N4337 , _f_permutation__round__N4335 ,
         _f_permutation__round__N4333 , _f_permutation__round__N4331 ,
         _f_permutation__round__N4329 , _f_permutation__round__N4327 ,
         _f_permutation__round__N4325 , _f_permutation__round__N4323 ,
         _f_permutation__round__N4321 , _f_permutation__round__N4319 ,
         _f_permutation__round__N4317 , _f_permutation__round__N4315 ,
         _f_permutation__round__N4313 , _f_permutation__round__N4311 ,
         _f_permutation__round__N4309 , _f_permutation__round__N4307 ,
         _f_permutation__round__N4305 , _f_permutation__round__N4303 ,
         _f_permutation__round__N4301 , _f_permutation__round__N4299 ,
         _f_permutation__round__N4297 , _f_permutation__round__N4295 ,
         _f_permutation__round__N4293 , _f_permutation__round__N4291 ,
         _f_permutation__round__N4289 , _f_permutation__round__N4287 ,
         _f_permutation__round__N4285 , _f_permutation__round__N4283 ,
         _f_permutation__round__N4281 , _f_permutation__round__N4279 ,
         _f_permutation__round__N4277 , _f_permutation__round__N4275 ,
         _f_permutation__round__N4273 , _f_permutation__round__N4271 ,
         _f_permutation__round__N4269 , _f_permutation__round__N4267 ,
         _f_permutation__round__N4265 , _f_permutation__round__N4263 ,
         _f_permutation__round__N4261 , _f_permutation__round__N4259 ,
         _f_permutation__round__N4257 , _f_permutation__round__N4255 ,
         _f_permutation__round__N4253 , _f_permutation__round__N4251 ,
         _f_permutation__round__N4249 , _f_permutation__round__N4247 ,
         _f_permutation__round__N4245 , _f_permutation__round__N4243 ,
         _f_permutation__round__N4241 , _f_permutation__round__N4239 ,
         _f_permutation__round__N4237 , _f_permutation__round__N4235 ,
         _f_permutation__round__N4233 , _f_permutation__round__N4231 ,
         _f_permutation__round__N4229 , _f_permutation__round__N4227 ,
         _f_permutation__round__N4225 , _f_permutation__round__N4223 ,
         _f_permutation__round__N4221 , _f_permutation__round__N4219 ,
         _f_permutation__round__N4217 , _f_permutation__round__N4215 ,
         _f_permutation__round__N4213 , _f_permutation__round__N4211 ,
         _f_permutation__round__N4209 , _f_permutation__round__N4207 ,
         _f_permutation__round__N4205 , _f_permutation__round__N4203 ,
         _f_permutation__round__N4201 , _f_permutation__round__N4199 ,
         _f_permutation__round__N4197 , _f_permutation__round__N4195 ,
         _f_permutation__round__N4193 , _f_permutation__round__N4191 ,
         _f_permutation__round__N4189 , _f_permutation__round__N4187 ,
         _f_permutation__round__N4185 , _f_permutation__round__N4183 ,
         _f_permutation__round__N4181 , _f_permutation__round__N4179 ,
         _f_permutation__round__N4177 , _f_permutation__round__N4175 ,
         _f_permutation__round__N4173 , _f_permutation__round__N4171 ,
         _f_permutation__round__N4169 , _f_permutation__round__N4167 ,
         _f_permutation__round__N4165 , _f_permutation__round__N4163 ,
         _f_permutation__round__N4161 , _f_permutation__round__N4159 ,
         _f_permutation__round__N4157 , _f_permutation__round__N4155 ,
         _f_permutation__round__N4153 , _f_permutation__round__N4151 ,
         _f_permutation__round__N4149 , _f_permutation__round__N4147 ,
         _f_permutation__round__N4145 , _f_permutation__round__N4143 ,
         _f_permutation__round__N4141 , _f_permutation__round__N4139 ,
         _f_permutation__round__N4137 , _f_permutation__round__N4135 ,
         _f_permutation__round__N4133 , _f_permutation__round__N4131 ,
         _f_permutation__round__N4129 , _f_permutation__round__N4127 ,
         _f_permutation__round__N4125 , _f_permutation__round__N4123 ,
         _f_permutation__round__N4121 , _f_permutation__round__N4119 ,
         _f_permutation__round__N4117 , _f_permutation__round__N4115 ,
         _f_permutation__round__N4113 , _f_permutation__round__N4111 ,
         _f_permutation__round__N4109 , _f_permutation__round__N4107 ,
         _f_permutation__round__N4105 , _f_permutation__round__N4103 ,
         _f_permutation__round__N4101 , _f_permutation__round__N4099 ,
         _f_permutation__round__N4097 , _f_permutation__round__N4095 ,
         _f_permutation__round__N4093 , _f_permutation__round__N4091 ,
         _f_permutation__round__N4089 , _f_permutation__round__N4087 ,
         _f_permutation__round__N4085 , _f_permutation__round__N4083 ,
         _f_permutation__round__N4081 , _f_permutation__round__N4079 ,
         _f_permutation__round__N4077 , _f_permutation__round__N4075 ,
         _f_permutation__round__N4073 , _f_permutation__round__N4071 ,
         _f_permutation__round__N4069 , _f_permutation__round__N4067 ,
         _f_permutation__round__N4065 , _f_permutation__round__N4063 ,
         _f_permutation__round__N4061 , _f_permutation__round__N4059 ,
         _f_permutation__round__N4057 , _f_permutation__round__N4055 ,
         _f_permutation__round__N4053 , _f_permutation__round__N4051 ,
         _f_permutation__round__N4049 , _f_permutation__round__N4047 ,
         _f_permutation__round__N4045 , _f_permutation__round__N4043 ,
         _f_permutation__round__N4041 , _f_permutation__round__N4039 ,
         _f_permutation__round__N4037 , _f_permutation__round__N4035 ,
         _f_permutation__round__N4033 , _f_permutation__round__N4031 ,
         _f_permutation__round__N4029 , _f_permutation__round__N4027 ,
         _f_permutation__round__N4025 , _f_permutation__round__N4023 ,
         _f_permutation__round__N4021 , _f_permutation__round__N4019 ,
         _f_permutation__round__N4017 , _f_permutation__round__N4015 ,
         _f_permutation__round__N4013 , _f_permutation__round__N4011 ,
         _f_permutation__round__N4009 , _f_permutation__round__N4007 ,
         _f_permutation__round__N4005 , _f_permutation__round__N4003 ,
         _f_permutation__round__N4001 , _f_permutation__round__N3999 ,
         _f_permutation__round__N3997 , _f_permutation__round__N3995 ,
         _f_permutation__round__N3993 , _f_permutation__round__N3991 ,
         _f_permutation__round__N3989 , _f_permutation__round__N3987 ,
         _f_permutation__round__N3985 , _f_permutation__round__N3983 ,
         _f_permutation__round__N3981 , _f_permutation__round__N3979 ,
         _f_permutation__round__N3977 , _f_permutation__round__N3975 ,
         _f_permutation__round__N3973 , _f_permutation__round__N3971 ,
         _f_permutation__round__N3969 , _f_permutation__round__N3967 ,
         _f_permutation__round__N3965 , _f_permutation__round__N3963 ,
         _f_permutation__round__N3961 , _f_permutation__round__N3959 ,
         _f_permutation__round__N3957 , _f_permutation__round__N3955 ,
         _f_permutation__round__N3953 , _f_permutation__round__N3951 ,
         _f_permutation__round__N3949 , _f_permutation__round__N3947 ,
         _f_permutation__round__N3945 , _f_permutation__round__N3943 ,
         _f_permutation__round__N3941 , _f_permutation__round__N3939 ,
         _f_permutation__round__N3937 , _f_permutation__round__N3935 ,
         _f_permutation__round__N3933 , _f_permutation__round__N3931 ,
         _f_permutation__round__N3929 , _f_permutation__round__N3927 ,
         _f_permutation__round__N3925 , _f_permutation__round__N3923 ,
         _f_permutation__round__N3921 , _f_permutation__round__N3919 ,
         _f_permutation__round__N3917 , _f_permutation__round__N3915 ,
         _f_permutation__round__N3913 , _f_permutation__round__N3911 ,
         _f_permutation__round__N3909 , _f_permutation__round__N3907 ,
         _f_permutation__round__N3905 , _f_permutation__round__N3903 ,
         _f_permutation__round__N3901 , _f_permutation__round__N3899 ,
         _f_permutation__round__N3897 , _f_permutation__round__N3895 ,
         _f_permutation__round__N3893 , _f_permutation__round__N3891 ,
         _f_permutation__round__N3889 , _f_permutation__round__N3887 ,
         _f_permutation__round__N3885 , _f_permutation__round__N3883 ,
         _f_permutation__round__N3881 , _f_permutation__round__N3879 ,
         _f_permutation__round__N3877 , _f_permutation__round__N3875 ,
         _f_permutation__round__N3873 , _f_permutation__round__N3871 ,
         _f_permutation__round__N3869 , _f_permutation__round__N3867 ,
         _f_permutation__round__N3865 , _f_permutation__round__N3863 ,
         _f_permutation__round__N3861 , _f_permutation__round__N3859 ,
         _f_permutation__round__N3857 , _f_permutation__round__N3855 ,
         _f_permutation__round__N3853 , _f_permutation__round__N3851 ,
         _f_permutation__round__N3849 , _f_permutation__round__N3847 ,
         _f_permutation__round__N3845 , _f_permutation__round__N3843 ,
         _f_permutation__round__N3841 , _f_permutation__round__N3839 ,
         _f_permutation__round__N3837 , _f_permutation__round__N3835 ,
         _f_permutation__round__N3833 , _f_permutation__round__N3831 ,
         _f_permutation__round__N3829 , _f_permutation__round__N3827 ,
         _f_permutation__round__N3825 , _f_permutation__round__N3823 ,
         _f_permutation__round__N3821 , _f_permutation__round__N3819 ,
         _f_permutation__round__N3817 , _f_permutation__round__N3815 ,
         _f_permutation__round__N3813 , _f_permutation__round__N3811 ,
         _f_permutation__round__N3809 , _f_permutation__round__N3807 ,
         _f_permutation__round__N3805 , _f_permutation__round__N3803 ,
         _f_permutation__round__N3801 , _f_permutation__round__N3799 ,
         _f_permutation__round__N3797 , _f_permutation__round__N3795 ,
         _f_permutation__round__N3793 , _f_permutation__round__N3791 ,
         _f_permutation__round__N3789 , _f_permutation__round__N3787 ,
         _f_permutation__round__N3785 , _f_permutation__round__N3783 ,
         _f_permutation__round__N3781 , _f_permutation__round__N3779 ,
         _f_permutation__round__N3777 , _f_permutation__round__N3775 ,
         _f_permutation__round__N3773 , _f_permutation__round__N3771 ,
         _f_permutation__round__N3769 , _f_permutation__round__N3767 ,
         _f_permutation__round__N3765 , _f_permutation__round__N3763 ,
         _f_permutation__round__N3761 , _f_permutation__round__N3759 ,
         _f_permutation__round__N3757 , _f_permutation__round__N3755 ,
         _f_permutation__round__N3753 , _f_permutation__round__N3751 ,
         _f_permutation__round__N3749 , _f_permutation__round__N3747 ,
         _f_permutation__round__N3745 , _f_permutation__round__N3743 ,
         _f_permutation__round__N3741 , _f_permutation__round__N3739 ,
         _f_permutation__round__N3737 , _f_permutation__round__N3735 ,
         _f_permutation__round__N3733 , _f_permutation__round__N3731 ,
         _f_permutation__round__N3729 , _f_permutation__round__N3727 ,
         _f_permutation__round__N3725 , _f_permutation__round__N3723 ,
         _f_permutation__round__N3721 , _f_permutation__round__N3719 ,
         _f_permutation__round__N3717 , _f_permutation__round__N3715 ,
         _f_permutation__round__N3713 , _f_permutation__round__N3711 ,
         _f_permutation__round__N3709 , _f_permutation__round__N3707 ,
         _f_permutation__round__N3705 , _f_permutation__round__N3703 ,
         _f_permutation__round__N3701 , _f_permutation__round__N3699 ,
         _f_permutation__round__N3697 , _f_permutation__round__N3695 ,
         _f_permutation__round__N3693 , _f_permutation__round__N3691 ,
         _f_permutation__round__N3689 , _f_permutation__round__N3687 ,
         _f_permutation__round__N3685 , _f_permutation__round__N3683 ,
         _f_permutation__round__N3681 , _f_permutation__round__N3679 ,
         _f_permutation__round__N3677 , _f_permutation__round__N3675 ,
         _f_permutation__round__N3673 , _f_permutation__round__N3671 ,
         _f_permutation__round__N3669 , _f_permutation__round__N3667 ,
         _f_permutation__round__N3665 , _f_permutation__round__N3663 ,
         _f_permutation__round__N3661 , _f_permutation__round__N3659 ,
         _f_permutation__round__N3657 , _f_permutation__round__N3655 ,
         _f_permutation__round__N3653 , _f_permutation__round__N3651 ,
         _f_permutation__round__N3649 , _f_permutation__round__N3647 ,
         _f_permutation__round__N3645 , _f_permutation__round__N3643 ,
         _f_permutation__round__N3641 , _f_permutation__round__N3639 ,
         _f_permutation__round__N3637 , _f_permutation__round__N3635 ,
         _f_permutation__round__N3633 , _f_permutation__round__N3631 ,
         _f_permutation__round__N3629 , _f_permutation__round__N3627 ,
         _f_permutation__round__N3625 , _f_permutation__round__N3623 ,
         _f_permutation__round__N3621 , _f_permutation__round__N3619 ,
         _f_permutation__round__N3617 , _f_permutation__round__N3615 ,
         _f_permutation__round__N3613 , _f_permutation__round__N3611 ,
         _f_permutation__round__N3609 , _f_permutation__round__N3607 ,
         _f_permutation__round__N3605 , _f_permutation__round__N3603 ,
         _f_permutation__round__N3601 , _f_permutation__round__N3599 ,
         _f_permutation__round__N3597 , _f_permutation__round__N3595 ,
         _f_permutation__round__N3593 , _f_permutation__round__N3591 ,
         _f_permutation__round__N3589 , _f_permutation__round__N3587 ,
         _f_permutation__round__N3585 , _f_permutation__round__N3583 ,
         _f_permutation__round__N3581 , _f_permutation__round__N3579 ,
         _f_permutation__round__N3577 , _f_permutation__round__N3575 ,
         _f_permutation__round__N3573 , _f_permutation__round__N3571 ,
         _f_permutation__round__N3569 , _f_permutation__round__N3567 ,
         _f_permutation__round__N3565 , _f_permutation__round__N3563 ,
         _f_permutation__round__N3561 , _f_permutation__round__N3559 ,
         _f_permutation__round__N3557 , _f_permutation__round__N3555 ,
         _f_permutation__round__N3553 , _f_permutation__round__N3551 ,
         _f_permutation__round__N3549 , _f_permutation__round__N3547 ,
         _f_permutation__round__N3545 , _f_permutation__round__N3543 ,
         _f_permutation__round__N3541 , _f_permutation__round__N3539 ,
         _f_permutation__round__N3537 , _f_permutation__round__N3535 ,
         _f_permutation__round__N3533 , _f_permutation__round__N3531 ,
         _f_permutation__round__N3529 , _f_permutation__round__N3527 ,
         _f_permutation__round__N3525 , _f_permutation__round__N3523 ,
         _f_permutation__round__N3521 , _f_permutation__round__N3519 ,
         _f_permutation__round__N3517 , _f_permutation__round__N3515 ,
         _f_permutation__round__N3513 , _f_permutation__round__N3511 ,
         _f_permutation__round__N3509 , _f_permutation__round__N3507 ,
         _f_permutation__round__N3505 , _f_permutation__round__N3503 ,
         _f_permutation__round__N3501 , _f_permutation__round__N3499 ,
         _f_permutation__round__N3497 , _f_permutation__round__N3495 ,
         _f_permutation__round__N3493 , _f_permutation__round__N3491 ,
         _f_permutation__round__N3489 , _f_permutation__round__N3487 ,
         _f_permutation__round__N3485 , _f_permutation__round__N3483 ,
         _f_permutation__round__N3481 , _f_permutation__round__N3479 ,
         _f_permutation__round__N3477 , _f_permutation__round__N3475 ,
         _f_permutation__round__N3473 , _f_permutation__round__N3471 ,
         _f_permutation__round__N3469 , _f_permutation__round__N3467 ,
         _f_permutation__round__N3465 , _f_permutation__round__N3463 ,
         _f_permutation__round__N3461 , _f_permutation__round__N3459 ,
         _f_permutation__round__N3457 , _f_permutation__round__N3455 ,
         _f_permutation__round__N3453 , _f_permutation__round__N3451 ,
         _f_permutation__round__N3449 , _f_permutation__round__N3447 ,
         _f_permutation__round__N3445 , _f_permutation__round__N3443 ,
         _f_permutation__round__N3441 , _f_permutation__round__N3439 ,
         _f_permutation__round__N3437 , _f_permutation__round__N3435 ,
         _f_permutation__round__N3433 , _f_permutation__round__N3431 ,
         _f_permutation__round__N3429 , _f_permutation__round__N3427 ,
         _f_permutation__round__N3425 , _f_permutation__round__N3423 ,
         _f_permutation__round__N3421 , _f_permutation__round__N3419 ,
         _f_permutation__round__N3417 , _f_permutation__round__N3415 ,
         _f_permutation__round__N3413 , _f_permutation__round__N3411 ,
         _f_permutation__round__N3409 , _f_permutation__round__N3407 ,
         _f_permutation__round__N3405 , _f_permutation__round__N3403 ,
         _f_permutation__round__N3401 , _f_permutation__round__N3399 ,
         _f_permutation__round__N3397 , _f_permutation__round__N3395 ,
         _f_permutation__round__N3393 , _f_permutation__round__N3391 ,
         _f_permutation__round__N3389 , _f_permutation__round__N3387 ,
         _f_permutation__round__N3385 , _f_permutation__round__N3383 ,
         _f_permutation__round__N3381 , _f_permutation__round__N3379 ,
         _f_permutation__round__N3377 , _f_permutation__round__N3375 ,
         _f_permutation__round__N3373 , _f_permutation__round__N3371 ,
         _f_permutation__round__N3369 , _f_permutation__round__N3367 ,
         _f_permutation__round__N3365 , _f_permutation__round__N3363 ,
         _f_permutation__round__N3361 , _f_permutation__round__N3359 ,
         _f_permutation__round__N3357 , _f_permutation__round__N3355 ,
         _f_permutation__round__N3353 , _f_permutation__round__N3351 ,
         _f_permutation__round__N3349 , _f_permutation__round__N3347 ,
         _f_permutation__round__N3345 , _f_permutation__round__N3343 ,
         _f_permutation__round__N3341 , _f_permutation__round__N3339 ,
         _f_permutation__round__N3337 , _f_permutation__round__N3335 ,
         _f_permutation__round__N3333 , _f_permutation__round__N3331 ,
         _f_permutation__round__N3329 , _f_permutation__round__N3327 ,
         _f_permutation__round__N3325 , _f_permutation__round__N3323 ,
         _f_permutation__round__N3321 , _f_permutation__round__N3319 ,
         _f_permutation__round__N3317 , _f_permutation__round__N3315 ,
         _f_permutation__round__N3313 , _f_permutation__round__N3311 ,
         _f_permutation__round__N3309 , _f_permutation__round__N3307 ,
         _f_permutation__round__N3305 , _f_permutation__round__N3303 ,
         _f_permutation__round__N3301 , _f_permutation__round__N3299 ,
         _f_permutation__round__N3297 , _f_permutation__round__N3295 ,
         _f_permutation__round__N3293 , _f_permutation__round__N3291 ,
         _f_permutation__round__N3289 , _f_permutation__round__N3287 ,
         _f_permutation__round__N3285 , _f_permutation__round__N3283 ,
         _f_permutation__round__N3281 , _f_permutation__round__N3279 ,
         _f_permutation__round__N3277 , _f_permutation__round__N3275 ,
         _f_permutation__round__N3273 , _f_permutation__round__N3271 ,
         _f_permutation__round__N3269 , _f_permutation__round__N3267 ,
         _f_permutation__round__N3265 , _f_permutation__round__N3263 ,
         _f_permutation__round__N3261 , _f_permutation__round__N3259 ,
         _f_permutation__round__N3257 , _f_permutation__round__N3255 ,
         _f_permutation__round__N3253 , _f_permutation__round__N3251 ,
         _f_permutation__round__N3249 , _f_permutation__round__N3247 ,
         _f_permutation__round__N3245 , _f_permutation__round__N3243 ,
         _f_permutation__round__N3241 , _f_permutation__round__N3239 ,
         _f_permutation__round__N3237 , _f_permutation__round__N3235 ,
         _f_permutation__round__N3233 , _f_permutation__round__N3231 ,
         _f_permutation__round__N3229 , _f_permutation__round__N3227 ,
         _f_permutation__round__N3225 , _f_permutation__round__N3223 ,
         _f_permutation__round__N3221 , _f_permutation__round__N3219 ,
         _f_permutation__round__N3217 , _f_permutation__round__N3215 ,
         _f_permutation__round__N3213 , _f_permutation__round__N3211 ,
         _f_permutation__round__N3209 , _f_permutation__round__N3207 ,
         _f_permutation__round__N3205 , _f_permutation__round__N3203 ,
         _f_permutation__round__N3201 , _f_permutation__round__N3199 ,
         _f_permutation__round__N3197 , _f_permutation__round__N3195 ,
         _f_permutation__round__N3193 , _f_permutation__round__N3191 ,
         _f_permutation__round__N3189 , _f_permutation__round__N3187 ,
         _f_permutation__round__N3185 , _f_permutation__round__N3183 ,
         _f_permutation__round__N3181 , _f_permutation__round__N3179 ,
         _f_permutation__round__N3177 , _f_permutation__round__N3175 ,
         _f_permutation__round__N3173 , _f_permutation__round__N3171 ,
         _f_permutation__round__N3169 , _f_permutation__round__N3167 ,
         _f_permutation__round__N3165 , _f_permutation__round__N3163 ,
         _f_permutation__round__N3161 , _f_permutation__round__N3159 ,
         _f_permutation__round__N3157 , _f_permutation__round__N3155 ,
         _f_permutation__round__N3153 , _f_permutation__round__N3151 ,
         _f_permutation__round__N3149 , _f_permutation__round__N3147 ,
         _f_permutation__round__N3145 , _f_permutation__round__N3143 ,
         _f_permutation__round__N3141 , _f_permutation__round__N3139 ,
         _f_permutation__round__N3137 , _f_permutation__round__N3135 ,
         _f_permutation__round__N3133 , _f_permutation__round__N3131 ,
         _f_permutation__round__N3129 , _f_permutation__round__N3127 ,
         _f_permutation__round__N3125 , _f_permutation__round__N3123 ,
         _f_permutation__round__N3121 , _f_permutation__round__N3119 ,
         _f_permutation__round__N3117 , _f_permutation__round__N3115 ,
         _f_permutation__round__N3113 , _f_permutation__round__N3111 ,
         _f_permutation__round__N3109 , _f_permutation__round__N3107 ,
         _f_permutation__round__N3105 , _f_permutation__round__N3103 ,
         _f_permutation__round__N3101 , _f_permutation__round__N3099 ,
         _f_permutation__round__N3097 , _f_permutation__round__N3095 ,
         _f_permutation__round__N3093 , _f_permutation__round__N3091 ,
         _f_permutation__round__N3089 , _f_permutation__round__N3087 ,
         _f_permutation__round__N3085 , _f_permutation__round__N3083 ,
         _f_permutation__round__N3081 , _f_permutation__round__N3079 ,
         _f_permutation__round__N3077 , _f_permutation__round__N3075 ,
         _f_permutation__round__N3073 , _f_permutation__round__N3071 ,
         _f_permutation__round__N3069 , _f_permutation__round__N3067 ,
         _f_permutation__round__N3065 , _f_permutation__round__N3063 ,
         _f_permutation__round__N3061 , _f_permutation__round__N3059 ,
         _f_permutation__round__N3057 , _f_permutation__round__N3055 ,
         _f_permutation__round__N3053 , _f_permutation__round__N3051 ,
         _f_permutation__round__N3049 , _f_permutation__round__N3047 ,
         _f_permutation__round__N3045 , _f_permutation__round__N3043 ,
         _f_permutation__round__N3041 , _f_permutation__round__N3039 ,
         _f_permutation__round__N3037 , _f_permutation__round__N3035 ,
         _f_permutation__round__N3033 , _f_permutation__round__N3031 ,
         _f_permutation__round__N3029 , _f_permutation__round__N3027 ,
         _f_permutation__round__N3025 , _f_permutation__round__N3023 ,
         _f_permutation__round__N3021 , _f_permutation__round__N3019 ,
         _f_permutation__round__N3017 , _f_permutation__round__N3015 ,
         _f_permutation__round__N3013 , _f_permutation__round__N3011 ,
         _f_permutation__round__N3009 , _f_permutation__round__N3007 ,
         _f_permutation__round__N3005 , _f_permutation__round__N3003 ,
         _f_permutation__round__N3001 , _f_permutation__round__N2999 ,
         _f_permutation__round__N2997 , _f_permutation__round__N2995 ,
         _f_permutation__round__N2993 , _f_permutation__round__N2991 ,
         _f_permutation__round__N2989 , _f_permutation__round__N2987 ,
         _f_permutation__round__N2985 , _f_permutation__round__N2983 ,
         _f_permutation__round__N2981 , _f_permutation__round__N2979 ,
         _f_permutation__round__N2977 , _f_permutation__round__N2975 ,
         _f_permutation__round__N2973 , _f_permutation__round__N2971 ,
         _f_permutation__round__N2969 , _f_permutation__round__N2967 ,
         _f_permutation__round__N2965 , _f_permutation__round__N2963 ,
         _f_permutation__round__N2961 , _f_permutation__round__N2959 ,
         _f_permutation__round__N2957 , _f_permutation__round__N2955 ,
         _f_permutation__round__N2953 , _f_permutation__round__N2951 ,
         _f_permutation__round__N2949 , _f_permutation__round__N2947 ,
         _f_permutation__round__N2945 , _f_permutation__round__N2943 ,
         _f_permutation__round__N2941 , _f_permutation__round__N2939 ,
         _f_permutation__round__N2937 , _f_permutation__round__N2935 ,
         _f_permutation__round__N2933 , _f_permutation__round__N2931 ,
         _f_permutation__round__N2929 , _f_permutation__round__N2927 ,
         _f_permutation__round__N2925 , _f_permutation__round__N2923 ,
         _f_permutation__round__N2921 , _f_permutation__round__N2919 ,
         _f_permutation__round__N2917 , _f_permutation__round__N2915 ,
         _f_permutation__round__N2913 , _f_permutation__round__N2911 ,
         _f_permutation__round__N2909 , _f_permutation__round__N2907 ,
         _f_permutation__round__N2905 , _f_permutation__round__N2903 ,
         _f_permutation__round__N2901 , _f_permutation__round__N2899 ,
         _f_permutation__round__N2897 , _f_permutation__round__N2895 ,
         _f_permutation__round__N2893 , _f_permutation__round__N2891 ,
         _f_permutation__round__N2889 , _f_permutation__round__N2887 ,
         _f_permutation__round__N2885 , _f_permutation__round__N2883 ,
         _f_permutation__round__N2881 , _f_permutation__round__N2879 ,
         _f_permutation__round__N2877 , _f_permutation__round__N2875 ,
         _f_permutation__round__N2873 , _f_permutation__round__N2871 ,
         _f_permutation__round__N2869 , _f_permutation__round__N2867 ,
         _f_permutation__round__N2865 , _f_permutation__round__N2863 ,
         _f_permutation__round__N2861 , _f_permutation__round__N2859 ,
         _f_permutation__round__N2857 , _f_permutation__round__N2855 ,
         _f_permutation__round__N2853 , _f_permutation__round__N2851 ,
         _f_permutation__round__N2849 , _f_permutation__round__N2847 ,
         _f_permutation__round__N2845 , _f_permutation__round__N2843 ,
         _f_permutation__round__N2841 , _f_permutation__round__N2839 ,
         _f_permutation__round__N2837 , _f_permutation__round__N2835 ,
         _f_permutation__round__N2833 , _f_permutation__round__N2831 ,
         _f_permutation__round__N2829 , _f_permutation__round__N2827 ,
         _f_permutation__round__N2825 , _f_permutation__round__N2823 ,
         _f_permutation__round__N2821 , _f_permutation__round__N2819 ,
         _f_permutation__round__N2817 , _f_permutation__round__N2815 ,
         _f_permutation__round__N2813 , _f_permutation__round__N2811 ,
         _f_permutation__round__N2809 , _f_permutation__round__N2807 ,
         _f_permutation__round__N2805 , _f_permutation__round__N2803 ,
         _f_permutation__round__N2801 , _f_permutation__round__N2799 ,
         _f_permutation__round__N2797 , _f_permutation__round__N2795 ,
         _f_permutation__round__N2793 , _f_permutation__round__N2791 ,
         _f_permutation__round__N2789 , _f_permutation__round__N2787 ,
         _f_permutation__round__N2785 , _f_permutation__round__N2783 ,
         _f_permutation__round__N2781 , _f_permutation__round__N2779 ,
         _f_permutation__round__N2777 , _f_permutation__round__N2775 ,
         _f_permutation__round__N2773 , _f_permutation__round__N2771 ,
         _f_permutation__round__N2769 , _f_permutation__round__N2767 ,
         _f_permutation__round__N2765 , _f_permutation__round__N2763 ,
         _f_permutation__round__N2761 , _f_permutation__round__N2759 ,
         _f_permutation__round__N2757 , _f_permutation__round__N2755 ,
         _f_permutation__round__N2753 , _f_permutation__round__N2751 ,
         _f_permutation__round__N2749 , _f_permutation__round__N2747 ,
         _f_permutation__round__N2745 , _f_permutation__round__N2743 ,
         _f_permutation__round__N2741 , _f_permutation__round__N2739 ,
         _f_permutation__round__N2737 , _f_permutation__round__N2735 ,
         _f_permutation__round__N2733 , _f_permutation__round__N2731 ,
         _f_permutation__round__N2729 , _f_permutation__round__N2727 ,
         _f_permutation__round__N2725 , _f_permutation__round__N2723 ,
         _f_permutation__round__N2721 , _f_permutation__round__N2719 ,
         _f_permutation__round__N2717 , _f_permutation__round__N2715 ,
         _f_permutation__round__N2713 , _f_permutation__round__N2711 ,
         _f_permutation__round__N2709 , _f_permutation__round__N2707 ,
         _f_permutation__round__N2705 , _f_permutation__round__N2703 ,
         _f_permutation__round__N2701 , _f_permutation__round__N2699 ,
         _f_permutation__round__N2697 , _f_permutation__round__N2695 ,
         _f_permutation__round__N2693 , _f_permutation__round__N2691 ,
         _f_permutation__round__N2689 , _f_permutation__round__N2687 ,
         _f_permutation__round__N2685 , _f_permutation__round__N2683 ,
         _f_permutation__round__N2681 , _f_permutation__round__N2679 ,
         _f_permutation__round__N2677 , _f_permutation__round__N2675 ,
         _f_permutation__round__N2673 , _f_permutation__round__N2671 ,
         _f_permutation__round__N2669 , _f_permutation__round__N2667 ,
         _f_permutation__round__N2665 , _f_permutation__round__N2663 ,
         _f_permutation__round__N2661 , _f_permutation__round__N2659 ,
         _f_permutation__round__N2657 , _f_permutation__round__N2655 ,
         _f_permutation__round__N2653 , _f_permutation__round__N2651 ,
         _f_permutation__round__N2649 , _f_permutation__round__N2647 ,
         _f_permutation__round__N2645 , _f_permutation__round__N2643 ,
         _f_permutation__round__N2641 , _f_permutation__round__N2639 ,
         _f_permutation__round__N2637 , _f_permutation__round__N2635 ,
         _f_permutation__round__N2633 , _f_permutation__round__N2631 ,
         _f_permutation__round__N2629 , _f_permutation__round__N2627 ,
         _f_permutation__round__N2625 , _f_permutation__round__N2623 ,
         _f_permutation__round__N2621 , _f_permutation__round__N2619 ,
         _f_permutation__round__N2617 , _f_permutation__round__N2615 ,
         _f_permutation__round__N2613 , _f_permutation__round__N2611 ,
         _f_permutation__round__N2609 , _f_permutation__round__N2607 ,
         _f_permutation__round__N2605 , _f_permutation__round__N2603 ,
         _f_permutation__round__N2601 , _f_permutation__round__N2599 ,
         _f_permutation__round__N2597 , _f_permutation__round__N2595 ,
         _f_permutation__round__N2593 , _f_permutation__round__N2591 ,
         _f_permutation__round__N2589 , _f_permutation__round__N2587 ,
         _f_permutation__round__N2585 , _f_permutation__round__N2583 ,
         _f_permutation__round__N2581 , _f_permutation__round__N2579 ,
         _f_permutation__round__N2577 , _f_permutation__round__N2575 ,
         _f_permutation__round__N2573 , _f_permutation__round__N2571 ,
         _f_permutation__round__N2569 , _f_permutation__round__N2567 ,
         _f_permutation__round__N2565 , _f_permutation__round__N2563 ,
         _f_permutation__round__N2561 , _f_permutation__round__c[64] ,
         _f_permutation__round__c[65] , _f_permutation__round__c[66] ,
         _f_permutation__round__c[67] , _f_permutation__round__c[68] ,
         _f_permutation__round__c[69] , _f_permutation__round__c[70] ,
         _f_permutation__round__c[71] , _f_permutation__round__c[72] ,
         _f_permutation__round__c[73] , _f_permutation__round__c[74] ,
         _f_permutation__round__c[75] , _f_permutation__round__c[76] ,
         _f_permutation__round__c[77] , _f_permutation__round__c[78] ,
         _f_permutation__round__c[79] , _f_permutation__round__c[80] ,
         _f_permutation__round__c[81] , _f_permutation__round__c[82] ,
         _f_permutation__round__c[83] , _f_permutation__round__c[84] ,
         _f_permutation__round__c[85] , _f_permutation__round__c[86] ,
         _f_permutation__round__c[87] , _f_permutation__round__c[88] ,
         _f_permutation__round__c[89] , _f_permutation__round__c[90] ,
         _f_permutation__round__c[91] , _f_permutation__round__c[92] ,
         _f_permutation__round__c[93] , _f_permutation__round__c[94] ,
         _f_permutation__round__c[95] , _f_permutation__round__c[96] ,
         _f_permutation__round__c[97] , _f_permutation__round__c[98] ,
         _f_permutation__round__c[99] , _f_permutation__round__c[100] ,
         _f_permutation__round__c[101] , _f_permutation__round__c[102] ,
         _f_permutation__round__c[103] , _f_permutation__round__c[104] ,
         _f_permutation__round__c[105] , _f_permutation__round__c[106] ,
         _f_permutation__round__c[107] , _f_permutation__round__c[108] ,
         _f_permutation__round__c[109] , _f_permutation__round__c[110] ,
         _f_permutation__round__c[111] , _f_permutation__round__c[112] ,
         _f_permutation__round__c[113] , _f_permutation__round__c[114] ,
         _f_permutation__round__c[115] , _f_permutation__round__c[116] ,
         _f_permutation__round__c[117] , _f_permutation__round__c[118] ,
         _f_permutation__round__c[119] , _f_permutation__round__c[120] ,
         _f_permutation__round__c[121] , _f_permutation__round__c[122] ,
         _f_permutation__round__c[123] , _f_permutation__round__c[124] ,
         _f_permutation__round__c[125] , _f_permutation__round__c[126] ,
         _f_permutation__round__c[127] , _f_permutation__round__c[128] ,
         _f_permutation__round__c[129] , _f_permutation__round__c[130] ,
         _f_permutation__round__c[131] , _f_permutation__round__c[132] ,
         _f_permutation__round__c[133] , _f_permutation__round__c[134] ,
         _f_permutation__round__c[135] , _f_permutation__round__c[136] ,
         _f_permutation__round__c[137] , _f_permutation__round__c[138] ,
         _f_permutation__round__c[139] , _f_permutation__round__c[140] ,
         _f_permutation__round__c[141] , _f_permutation__round__c[142] ,
         _f_permutation__round__c[143] , _f_permutation__round__c[144] ,
         _f_permutation__round__c[145] , _f_permutation__round__c[146] ,
         _f_permutation__round__c[147] , _f_permutation__round__c[148] ,
         _f_permutation__round__c[149] , _f_permutation__round__c[150] ,
         _f_permutation__round__c[151] , _f_permutation__round__c[152] ,
         _f_permutation__round__c[153] , _f_permutation__round__c[154] ,
         _f_permutation__round__c[155] , _f_permutation__round__c[156] ,
         _f_permutation__round__c[157] , _f_permutation__round__c[158] ,
         _f_permutation__round__c[159] , _f_permutation__round__c[160] ,
         _f_permutation__round__c[161] , _f_permutation__round__c[162] ,
         _f_permutation__round__c[163] , _f_permutation__round__c[164] ,
         _f_permutation__round__c[165] , _f_permutation__round__c[166] ,
         _f_permutation__round__c[167] , _f_permutation__round__c[168] ,
         _f_permutation__round__c[169] , _f_permutation__round__c[170] ,
         _f_permutation__round__c[171] , _f_permutation__round__c[172] ,
         _f_permutation__round__c[173] , _f_permutation__round__c[174] ,
         _f_permutation__round__c[175] , _f_permutation__round__c[176] ,
         _f_permutation__round__c[177] , _f_permutation__round__c[178] ,
         _f_permutation__round__c[179] , _f_permutation__round__c[180] ,
         _f_permutation__round__c[181] , _f_permutation__round__c[182] ,
         _f_permutation__round__c[183] , _f_permutation__round__c[184] ,
         _f_permutation__round__c[185] , _f_permutation__round__c[186] ,
         _f_permutation__round__c[187] , _f_permutation__round__c[188] ,
         _f_permutation__round__c[189] , _f_permutation__round__c[190] ,
         _f_permutation__round__c[191] , _f_permutation__round__c[192] ,
         _f_permutation__round__c[193] , _f_permutation__round__c[194] ,
         _f_permutation__round__c[195] , _f_permutation__round__c[196] ,
         _f_permutation__round__c[197] , _f_permutation__round__c[198] ,
         _f_permutation__round__c[199] , _f_permutation__round__c[200] ,
         _f_permutation__round__c[201] , _f_permutation__round__c[202] ,
         _f_permutation__round__c[203] , _f_permutation__round__c[204] ,
         _f_permutation__round__c[205] , _f_permutation__round__c[206] ,
         _f_permutation__round__c[207] , _f_permutation__round__c[208] ,
         _f_permutation__round__c[209] , _f_permutation__round__c[210] ,
         _f_permutation__round__c[211] , _f_permutation__round__c[212] ,
         _f_permutation__round__c[213] , _f_permutation__round__c[214] ,
         _f_permutation__round__c[215] , _f_permutation__round__c[216] ,
         _f_permutation__round__c[217] , _f_permutation__round__c[218] ,
         _f_permutation__round__c[219] , _f_permutation__round__c[220] ,
         _f_permutation__round__c[221] , _f_permutation__round__c[222] ,
         _f_permutation__round__c[223] , _f_permutation__round__c[224] ,
         _f_permutation__round__c[225] , _f_permutation__round__c[226] ,
         _f_permutation__round__c[227] , _f_permutation__round__c[228] ,
         _f_permutation__round__c[229] , _f_permutation__round__c[230] ,
         _f_permutation__round__c[231] , _f_permutation__round__c[232] ,
         _f_permutation__round__c[233] , _f_permutation__round__c[234] ,
         _f_permutation__round__c[235] , _f_permutation__round__c[236] ,
         _f_permutation__round__c[237] , _f_permutation__round__c[238] ,
         _f_permutation__round__c[239] , _f_permutation__round__c[240] ,
         _f_permutation__round__c[241] , _f_permutation__round__c[242] ,
         _f_permutation__round__c[243] , _f_permutation__round__c[244] ,
         _f_permutation__round__c[245] , _f_permutation__round__c[246] ,
         _f_permutation__round__c[247] , _f_permutation__round__c[248] ,
         _f_permutation__round__c[249] , _f_permutation__round__c[250] ,
         _f_permutation__round__c[251] , _f_permutation__round__c[252] ,
         _f_permutation__round__c[253] , _f_permutation__round__c[254] ,
         _f_permutation__round__c[255] , _f_permutation__round__c[256] ,
         _f_permutation__round__c[257] , _f_permutation__round__c[258] ,
         _f_permutation__round__c[259] , _f_permutation__round__c[260] ,
         _f_permutation__round__c[261] , _f_permutation__round__c[262] ,
         _f_permutation__round__c[263] , _f_permutation__round__c[264] ,
         _f_permutation__round__c[265] , _f_permutation__round__c[266] ,
         _f_permutation__round__c[267] , _f_permutation__round__c[268] ,
         _f_permutation__round__c[269] , _f_permutation__round__c[270] ,
         _f_permutation__round__c[271] , _f_permutation__round__c[272] ,
         _f_permutation__round__c[273] , _f_permutation__round__c[274] ,
         _f_permutation__round__c[275] , _f_permutation__round__c[276] ,
         _f_permutation__round__c[277] , _f_permutation__round__c[278] ,
         _f_permutation__round__c[279] , _f_permutation__round__c[280] ,
         _f_permutation__round__c[281] , _f_permutation__round__c[282] ,
         _f_permutation__round__c[283] , _f_permutation__round__c[284] ,
         _f_permutation__round__c[285] , _f_permutation__round__c[286] ,
         _f_permutation__round__c[287] , _f_permutation__round__c[288] ,
         _f_permutation__round__c[289] , _f_permutation__round__c[290] ,
         _f_permutation__round__c[291] , _f_permutation__round__c[292] ,
         _f_permutation__round__c[293] , _f_permutation__round__c[294] ,
         _f_permutation__round__c[295] , _f_permutation__round__c[296] ,
         _f_permutation__round__c[297] , _f_permutation__round__c[298] ,
         _f_permutation__round__c[299] , _f_permutation__round__c[300] ,
         _f_permutation__round__c[301] , _f_permutation__round__c[302] ,
         _f_permutation__round__c[303] , _f_permutation__round__c[304] ,
         _f_permutation__round__c[305] , _f_permutation__round__c[306] ,
         _f_permutation__round__c[307] , _f_permutation__round__c[308] ,
         _f_permutation__round__c[309] , _f_permutation__round__c[310] ,
         _f_permutation__round__c[311] , _f_permutation__round__c[312] ,
         _f_permutation__round__c[313] , _f_permutation__round__c[314] ,
         _f_permutation__round__c[315] , _f_permutation__round__c[316] ,
         _f_permutation__round__c[317] , _f_permutation__round__c[318] ,
         _f_permutation__round__c[319] , _f_permutation__round__c[320] ,
         _f_permutation__round__c[321] , _f_permutation__round__c[322] ,
         _f_permutation__round__c[323] , _f_permutation__round__c[324] ,
         _f_permutation__round__c[325] , _f_permutation__round__c[326] ,
         _f_permutation__round__c[327] , _f_permutation__round__c[328] ,
         _f_permutation__round__c[329] , _f_permutation__round__c[330] ,
         _f_permutation__round__c[331] , _f_permutation__round__c[332] ,
         _f_permutation__round__c[333] , _f_permutation__round__c[334] ,
         _f_permutation__round__c[335] , _f_permutation__round__c[336] ,
         _f_permutation__round__c[337] , _f_permutation__round__c[338] ,
         _f_permutation__round__c[339] , _f_permutation__round__c[340] ,
         _f_permutation__round__c[341] , _f_permutation__round__c[342] ,
         _f_permutation__round__c[343] , _f_permutation__round__c[344] ,
         _f_permutation__round__c[345] , _f_permutation__round__c[346] ,
         _f_permutation__round__c[347] , _f_permutation__round__c[348] ,
         _f_permutation__round__c[349] , _f_permutation__round__c[350] ,
         _f_permutation__round__c[351] , _f_permutation__round__c[352] ,
         _f_permutation__round__c[353] , _f_permutation__round__c[354] ,
         _f_permutation__round__c[355] , _f_permutation__round__c[356] ,
         _f_permutation__round__c[357] , _f_permutation__round__c[358] ,
         _f_permutation__round__c[359] , _f_permutation__round__c[360] ,
         _f_permutation__round__c[361] , _f_permutation__round__c[362] ,
         _f_permutation__round__c[363] , _f_permutation__round__c[364] ,
         _f_permutation__round__c[365] , _f_permutation__round__c[366] ,
         _f_permutation__round__c[367] , _f_permutation__round__c[368] ,
         _f_permutation__round__c[369] , _f_permutation__round__c[370] ,
         _f_permutation__round__c[371] , _f_permutation__round__c[372] ,
         _f_permutation__round__c[373] , _f_permutation__round__c[374] ,
         _f_permutation__round__c[375] , _f_permutation__round__c[376] ,
         _f_permutation__round__c[377] , _f_permutation__round__c[378] ,
         _f_permutation__round__c[379] , _f_permutation__round__c[380] ,
         _f_permutation__round__c[381] , _f_permutation__round__c[382] ,
         _f_permutation__round__c[383] , _f_permutation__round__c[384] ,
         _f_permutation__round__c[385] , _f_permutation__round__c[386] ,
         _f_permutation__round__c[387] , _f_permutation__round__c[388] ,
         _f_permutation__round__c[389] , _f_permutation__round__c[390] ,
         _f_permutation__round__c[391] , _f_permutation__round__c[392] ,
         _f_permutation__round__c[393] , _f_permutation__round__c[394] ,
         _f_permutation__round__c[395] , _f_permutation__round__c[396] ,
         _f_permutation__round__c[397] , _f_permutation__round__c[398] ,
         _f_permutation__round__c[399] , _f_permutation__round__c[400] ,
         _f_permutation__round__c[401] , _f_permutation__round__c[402] ,
         _f_permutation__round__c[403] , _f_permutation__round__c[404] ,
         _f_permutation__round__c[405] , _f_permutation__round__c[406] ,
         _f_permutation__round__c[407] , _f_permutation__round__c[408] ,
         _f_permutation__round__c[409] , _f_permutation__round__c[410] ,
         _f_permutation__round__c[411] , _f_permutation__round__c[412] ,
         _f_permutation__round__c[413] , _f_permutation__round__c[414] ,
         _f_permutation__round__c[415] , _f_permutation__round__c[416] ,
         _f_permutation__round__c[417] , _f_permutation__round__c[418] ,
         _f_permutation__round__c[419] , _f_permutation__round__c[420] ,
         _f_permutation__round__c[421] , _f_permutation__round__c[422] ,
         _f_permutation__round__c[423] , _f_permutation__round__c[424] ,
         _f_permutation__round__c[425] , _f_permutation__round__c[426] ,
         _f_permutation__round__c[427] , _f_permutation__round__c[428] ,
         _f_permutation__round__c[429] , _f_permutation__round__c[430] ,
         _f_permutation__round__c[431] , _f_permutation__round__c[432] ,
         _f_permutation__round__c[433] , _f_permutation__round__c[434] ,
         _f_permutation__round__c[435] , _f_permutation__round__c[436] ,
         _f_permutation__round__c[437] , _f_permutation__round__c[438] ,
         _f_permutation__round__c[439] , _f_permutation__round__c[440] ,
         _f_permutation__round__c[441] , _f_permutation__round__c[442] ,
         _f_permutation__round__c[443] , _f_permutation__round__c[444] ,
         _f_permutation__round__c[445] , _f_permutation__round__c[446] ,
         _f_permutation__round__c[447] , _f_permutation__round__c[448] ,
         _f_permutation__round__c[449] , _f_permutation__round__c[450] ,
         _f_permutation__round__c[451] , _f_permutation__round__c[452] ,
         _f_permutation__round__c[453] , _f_permutation__round__c[454] ,
         _f_permutation__round__c[455] , _f_permutation__round__c[456] ,
         _f_permutation__round__c[457] , _f_permutation__round__c[458] ,
         _f_permutation__round__c[459] , _f_permutation__round__c[460] ,
         _f_permutation__round__c[461] , _f_permutation__round__c[462] ,
         _f_permutation__round__c[463] , _f_permutation__round__c[464] ,
         _f_permutation__round__c[465] , _f_permutation__round__c[466] ,
         _f_permutation__round__c[467] , _f_permutation__round__c[468] ,
         _f_permutation__round__c[469] , _f_permutation__round__c[470] ,
         _f_permutation__round__c[471] , _f_permutation__round__c[472] ,
         _f_permutation__round__c[473] , _f_permutation__round__c[474] ,
         _f_permutation__round__c[475] , _f_permutation__round__c[476] ,
         _f_permutation__round__c[477] , _f_permutation__round__c[478] ,
         _f_permutation__round__c[479] , _f_permutation__round__c[480] ,
         _f_permutation__round__c[481] , _f_permutation__round__c[482] ,
         _f_permutation__round__c[483] , _f_permutation__round__c[484] ,
         _f_permutation__round__c[485] , _f_permutation__round__c[486] ,
         _f_permutation__round__c[487] , _f_permutation__round__c[488] ,
         _f_permutation__round__c[489] , _f_permutation__round__c[490] ,
         _f_permutation__round__c[491] , _f_permutation__round__c[492] ,
         _f_permutation__round__c[493] , _f_permutation__round__c[494] ,
         _f_permutation__round__c[495] , _f_permutation__round__c[496] ,
         _f_permutation__round__c[497] , _f_permutation__round__c[498] ,
         _f_permutation__round__c[499] , _f_permutation__round__c[500] ,
         _f_permutation__round__c[501] , _f_permutation__round__c[502] ,
         _f_permutation__round__c[503] , _f_permutation__round__c[504] ,
         _f_permutation__round__c[505] , _f_permutation__round__c[506] ,
         _f_permutation__round__c[507] , _f_permutation__round__c[508] ,
         _f_permutation__round__c[509] , _f_permutation__round__c[510] ,
         _f_permutation__round__c[511] , _f_permutation__round__c[512] ,
         _f_permutation__round__c[513] , _f_permutation__round__c[514] ,
         _f_permutation__round__c[515] , _f_permutation__round__c[516] ,
         _f_permutation__round__c[517] , _f_permutation__round__c[518] ,
         _f_permutation__round__c[519] , _f_permutation__round__c[520] ,
         _f_permutation__round__c[521] , _f_permutation__round__c[522] ,
         _f_permutation__round__c[523] , _f_permutation__round__c[524] ,
         _f_permutation__round__c[525] , _f_permutation__round__c[526] ,
         _f_permutation__round__c[527] , _f_permutation__round__c[528] ,
         _f_permutation__round__c[529] , _f_permutation__round__c[530] ,
         _f_permutation__round__c[531] , _f_permutation__round__c[532] ,
         _f_permutation__round__c[533] , _f_permutation__round__c[534] ,
         _f_permutation__round__c[535] , _f_permutation__round__c[536] ,
         _f_permutation__round__c[537] , _f_permutation__round__c[538] ,
         _f_permutation__round__c[539] , _f_permutation__round__c[540] ,
         _f_permutation__round__c[541] , _f_permutation__round__c[542] ,
         _f_permutation__round__c[543] , _f_permutation__round__c[544] ,
         _f_permutation__round__c[545] , _f_permutation__round__c[546] ,
         _f_permutation__round__c[547] , _f_permutation__round__c[548] ,
         _f_permutation__round__c[549] , _f_permutation__round__c[550] ,
         _f_permutation__round__c[551] , _f_permutation__round__c[552] ,
         _f_permutation__round__c[553] , _f_permutation__round__c[554] ,
         _f_permutation__round__c[555] , _f_permutation__round__c[556] ,
         _f_permutation__round__c[557] , _f_permutation__round__c[558] ,
         _f_permutation__round__c[559] , _f_permutation__round__c[560] ,
         _f_permutation__round__c[561] , _f_permutation__round__c[562] ,
         _f_permutation__round__c[563] , _f_permutation__round__c[564] ,
         _f_permutation__round__c[565] , _f_permutation__round__c[566] ,
         _f_permutation__round__c[567] , _f_permutation__round__c[568] ,
         _f_permutation__round__c[569] , _f_permutation__round__c[570] ,
         _f_permutation__round__c[571] , _f_permutation__round__c[572] ,
         _f_permutation__round__c[573] , _f_permutation__round__c[574] ,
         _f_permutation__round__c[575] , _f_permutation__round__c[576] ,
         _f_permutation__round__c[577] , _f_permutation__round__c[578] ,
         _f_permutation__round__c[579] , _f_permutation__round__c[580] ,
         _f_permutation__round__c[581] , _f_permutation__round__c[582] ,
         _f_permutation__round__c[583] , _f_permutation__round__c[584] ,
         _f_permutation__round__c[585] , _f_permutation__round__c[586] ,
         _f_permutation__round__c[587] , _f_permutation__round__c[588] ,
         _f_permutation__round__c[589] , _f_permutation__round__c[590] ,
         _f_permutation__round__c[591] , _f_permutation__round__c[592] ,
         _f_permutation__round__c[593] , _f_permutation__round__c[594] ,
         _f_permutation__round__c[595] , _f_permutation__round__c[596] ,
         _f_permutation__round__c[597] , _f_permutation__round__c[598] ,
         _f_permutation__round__c[599] , _f_permutation__round__c[600] ,
         _f_permutation__round__c[601] , _f_permutation__round__c[602] ,
         _f_permutation__round__c[603] , _f_permutation__round__c[604] ,
         _f_permutation__round__c[605] , _f_permutation__round__c[606] ,
         _f_permutation__round__c[607] , _f_permutation__round__c[608] ,
         _f_permutation__round__c[609] , _f_permutation__round__c[610] ,
         _f_permutation__round__c[611] , _f_permutation__round__c[612] ,
         _f_permutation__round__c[613] , _f_permutation__round__c[614] ,
         _f_permutation__round__c[615] , _f_permutation__round__c[616] ,
         _f_permutation__round__c[617] , _f_permutation__round__c[618] ,
         _f_permutation__round__c[619] , _f_permutation__round__c[620] ,
         _f_permutation__round__c[621] , _f_permutation__round__c[622] ,
         _f_permutation__round__c[623] , _f_permutation__round__c[624] ,
         _f_permutation__round__c[625] , _f_permutation__round__c[626] ,
         _f_permutation__round__c[627] , _f_permutation__round__c[628] ,
         _f_permutation__round__c[629] , _f_permutation__round__c[630] ,
         _f_permutation__round__c[631] , _f_permutation__round__c[632] ,
         _f_permutation__round__c[633] , _f_permutation__round__c[634] ,
         _f_permutation__round__c[635] , _f_permutation__round__c[636] ,
         _f_permutation__round__c[637] , _f_permutation__round__c[638] ,
         _f_permutation__round__c[639] , _f_permutation__round__c[640] ,
         _f_permutation__round__c[641] , _f_permutation__round__c[642] ,
         _f_permutation__round__c[643] , _f_permutation__round__c[644] ,
         _f_permutation__round__c[645] , _f_permutation__round__c[646] ,
         _f_permutation__round__c[647] , _f_permutation__round__c[648] ,
         _f_permutation__round__c[649] , _f_permutation__round__c[650] ,
         _f_permutation__round__c[651] , _f_permutation__round__c[652] ,
         _f_permutation__round__c[653] , _f_permutation__round__c[654] ,
         _f_permutation__round__c[655] , _f_permutation__round__c[656] ,
         _f_permutation__round__c[657] , _f_permutation__round__c[658] ,
         _f_permutation__round__c[659] , _f_permutation__round__c[660] ,
         _f_permutation__round__c[661] , _f_permutation__round__c[662] ,
         _f_permutation__round__c[663] , _f_permutation__round__c[664] ,
         _f_permutation__round__c[665] , _f_permutation__round__c[666] ,
         _f_permutation__round__c[667] , _f_permutation__round__c[668] ,
         _f_permutation__round__c[669] , _f_permutation__round__c[670] ,
         _f_permutation__round__c[671] , _f_permutation__round__c[672] ,
         _f_permutation__round__c[673] , _f_permutation__round__c[674] ,
         _f_permutation__round__c[675] , _f_permutation__round__c[676] ,
         _f_permutation__round__c[677] , _f_permutation__round__c[678] ,
         _f_permutation__round__c[679] , _f_permutation__round__c[680] ,
         _f_permutation__round__c[681] , _f_permutation__round__c[682] ,
         _f_permutation__round__c[683] , _f_permutation__round__c[684] ,
         _f_permutation__round__c[685] , _f_permutation__round__c[686] ,
         _f_permutation__round__c[687] , _f_permutation__round__c[688] ,
         _f_permutation__round__c[689] , _f_permutation__round__c[690] ,
         _f_permutation__round__c[691] , _f_permutation__round__c[692] ,
         _f_permutation__round__c[693] , _f_permutation__round__c[694] ,
         _f_permutation__round__c[695] , _f_permutation__round__c[696] ,
         _f_permutation__round__c[697] , _f_permutation__round__c[698] ,
         _f_permutation__round__c[699] , _f_permutation__round__c[700] ,
         _f_permutation__round__c[701] , _f_permutation__round__c[702] ,
         _f_permutation__round__c[703] , _f_permutation__round__c[704] ,
         _f_permutation__round__c[705] , _f_permutation__round__c[706] ,
         _f_permutation__round__c[707] , _f_permutation__round__c[708] ,
         _f_permutation__round__c[709] , _f_permutation__round__c[710] ,
         _f_permutation__round__c[711] , _f_permutation__round__c[712] ,
         _f_permutation__round__c[713] , _f_permutation__round__c[714] ,
         _f_permutation__round__c[715] , _f_permutation__round__c[716] ,
         _f_permutation__round__c[717] , _f_permutation__round__c[718] ,
         _f_permutation__round__c[719] , _f_permutation__round__c[720] ,
         _f_permutation__round__c[721] , _f_permutation__round__c[722] ,
         _f_permutation__round__c[723] , _f_permutation__round__c[724] ,
         _f_permutation__round__c[725] , _f_permutation__round__c[726] ,
         _f_permutation__round__c[727] , _f_permutation__round__c[728] ,
         _f_permutation__round__c[729] , _f_permutation__round__c[730] ,
         _f_permutation__round__c[731] , _f_permutation__round__c[732] ,
         _f_permutation__round__c[733] , _f_permutation__round__c[734] ,
         _f_permutation__round__c[735] , _f_permutation__round__c[736] ,
         _f_permutation__round__c[737] , _f_permutation__round__c[738] ,
         _f_permutation__round__c[739] , _f_permutation__round__c[740] ,
         _f_permutation__round__c[741] , _f_permutation__round__c[742] ,
         _f_permutation__round__c[743] , _f_permutation__round__c[744] ,
         _f_permutation__round__c[745] , _f_permutation__round__c[746] ,
         _f_permutation__round__c[747] , _f_permutation__round__c[748] ,
         _f_permutation__round__c[749] , _f_permutation__round__c[750] ,
         _f_permutation__round__c[751] , _f_permutation__round__c[752] ,
         _f_permutation__round__c[753] , _f_permutation__round__c[754] ,
         _f_permutation__round__c[755] , _f_permutation__round__c[756] ,
         _f_permutation__round__c[757] , _f_permutation__round__c[758] ,
         _f_permutation__round__c[759] , _f_permutation__round__c[760] ,
         _f_permutation__round__c[761] , _f_permutation__round__c[762] ,
         _f_permutation__round__c[763] , _f_permutation__round__c[764] ,
         _f_permutation__round__c[765] , _f_permutation__round__c[766] ,
         _f_permutation__round__c[767] , _f_permutation__round__c[768] ,
         _f_permutation__round__c[769] , _f_permutation__round__c[770] ,
         _f_permutation__round__c[771] , _f_permutation__round__c[772] ,
         _f_permutation__round__c[773] , _f_permutation__round__c[774] ,
         _f_permutation__round__c[775] , _f_permutation__round__c[776] ,
         _f_permutation__round__c[777] , _f_permutation__round__c[778] ,
         _f_permutation__round__c[779] , _f_permutation__round__c[780] ,
         _f_permutation__round__c[781] , _f_permutation__round__c[782] ,
         _f_permutation__round__c[783] , _f_permutation__round__c[784] ,
         _f_permutation__round__c[785] , _f_permutation__round__c[786] ,
         _f_permutation__round__c[787] , _f_permutation__round__c[788] ,
         _f_permutation__round__c[789] , _f_permutation__round__c[790] ,
         _f_permutation__round__c[791] , _f_permutation__round__c[792] ,
         _f_permutation__round__c[793] , _f_permutation__round__c[794] ,
         _f_permutation__round__c[795] , _f_permutation__round__c[796] ,
         _f_permutation__round__c[797] , _f_permutation__round__c[798] ,
         _f_permutation__round__c[799] , _f_permutation__round__c[800] ,
         _f_permutation__round__c[801] , _f_permutation__round__c[802] ,
         _f_permutation__round__c[803] , _f_permutation__round__c[804] ,
         _f_permutation__round__c[805] , _f_permutation__round__c[806] ,
         _f_permutation__round__c[807] , _f_permutation__round__c[808] ,
         _f_permutation__round__c[809] , _f_permutation__round__c[810] ,
         _f_permutation__round__c[811] , _f_permutation__round__c[812] ,
         _f_permutation__round__c[813] , _f_permutation__round__c[814] ,
         _f_permutation__round__c[815] , _f_permutation__round__c[816] ,
         _f_permutation__round__c[817] , _f_permutation__round__c[818] ,
         _f_permutation__round__c[819] , _f_permutation__round__c[820] ,
         _f_permutation__round__c[821] , _f_permutation__round__c[822] ,
         _f_permutation__round__c[823] , _f_permutation__round__c[824] ,
         _f_permutation__round__c[825] , _f_permutation__round__c[826] ,
         _f_permutation__round__c[827] , _f_permutation__round__c[828] ,
         _f_permutation__round__c[829] , _f_permutation__round__c[830] ,
         _f_permutation__round__c[831] , _f_permutation__round__c[832] ,
         _f_permutation__round__c[833] , _f_permutation__round__c[834] ,
         _f_permutation__round__c[835] , _f_permutation__round__c[836] ,
         _f_permutation__round__c[837] , _f_permutation__round__c[838] ,
         _f_permutation__round__c[839] , _f_permutation__round__c[840] ,
         _f_permutation__round__c[841] , _f_permutation__round__c[842] ,
         _f_permutation__round__c[843] , _f_permutation__round__c[844] ,
         _f_permutation__round__c[845] , _f_permutation__round__c[846] ,
         _f_permutation__round__c[847] , _f_permutation__round__c[848] ,
         _f_permutation__round__c[849] , _f_permutation__round__c[850] ,
         _f_permutation__round__c[851] , _f_permutation__round__c[852] ,
         _f_permutation__round__c[853] , _f_permutation__round__c[854] ,
         _f_permutation__round__c[855] , _f_permutation__round__c[856] ,
         _f_permutation__round__c[857] , _f_permutation__round__c[858] ,
         _f_permutation__round__c[859] , _f_permutation__round__c[860] ,
         _f_permutation__round__c[861] , _f_permutation__round__c[862] ,
         _f_permutation__round__c[863] , _f_permutation__round__c[864] ,
         _f_permutation__round__c[865] , _f_permutation__round__c[866] ,
         _f_permutation__round__c[867] , _f_permutation__round__c[868] ,
         _f_permutation__round__c[869] , _f_permutation__round__c[870] ,
         _f_permutation__round__c[871] , _f_permutation__round__c[872] ,
         _f_permutation__round__c[873] , _f_permutation__round__c[874] ,
         _f_permutation__round__c[875] , _f_permutation__round__c[876] ,
         _f_permutation__round__c[877] , _f_permutation__round__c[878] ,
         _f_permutation__round__c[879] , _f_permutation__round__c[880] ,
         _f_permutation__round__c[881] , _f_permutation__round__c[882] ,
         _f_permutation__round__c[883] , _f_permutation__round__c[884] ,
         _f_permutation__round__c[885] , _f_permutation__round__c[886] ,
         _f_permutation__round__c[887] , _f_permutation__round__c[888] ,
         _f_permutation__round__c[889] , _f_permutation__round__c[890] ,
         _f_permutation__round__c[891] , _f_permutation__round__c[892] ,
         _f_permutation__round__c[893] , _f_permutation__round__c[894] ,
         _f_permutation__round__c[895] , _f_permutation__round__c[896] ,
         _f_permutation__round__c[897] , _f_permutation__round__c[898] ,
         _f_permutation__round__c[899] , _f_permutation__round__c[900] ,
         _f_permutation__round__c[901] , _f_permutation__round__c[902] ,
         _f_permutation__round__c[903] , _f_permutation__round__c[904] ,
         _f_permutation__round__c[905] , _f_permutation__round__c[906] ,
         _f_permutation__round__c[907] , _f_permutation__round__c[908] ,
         _f_permutation__round__c[909] , _f_permutation__round__c[910] ,
         _f_permutation__round__c[911] , _f_permutation__round__c[912] ,
         _f_permutation__round__c[913] , _f_permutation__round__c[914] ,
         _f_permutation__round__c[915] , _f_permutation__round__c[916] ,
         _f_permutation__round__c[917] , _f_permutation__round__c[918] ,
         _f_permutation__round__c[919] , _f_permutation__round__c[920] ,
         _f_permutation__round__c[921] , _f_permutation__round__c[922] ,
         _f_permutation__round__c[923] , _f_permutation__round__c[924] ,
         _f_permutation__round__c[925] , _f_permutation__round__c[926] ,
         _f_permutation__round__c[927] , _f_permutation__round__c[928] ,
         _f_permutation__round__c[929] , _f_permutation__round__c[930] ,
         _f_permutation__round__c[931] , _f_permutation__round__c[932] ,
         _f_permutation__round__c[933] , _f_permutation__round__c[934] ,
         _f_permutation__round__c[935] , _f_permutation__round__c[936] ,
         _f_permutation__round__c[937] , _f_permutation__round__c[938] ,
         _f_permutation__round__c[939] , _f_permutation__round__c[940] ,
         _f_permutation__round__c[941] , _f_permutation__round__c[942] ,
         _f_permutation__round__c[943] , _f_permutation__round__c[944] ,
         _f_permutation__round__c[945] , _f_permutation__round__c[946] ,
         _f_permutation__round__c[947] , _f_permutation__round__c[948] ,
         _f_permutation__round__c[949] , _f_permutation__round__c[950] ,
         _f_permutation__round__c[951] , _f_permutation__round__c[952] ,
         _f_permutation__round__c[953] , _f_permutation__round__c[954] ,
         _f_permutation__round__c[955] , _f_permutation__round__c[956] ,
         _f_permutation__round__c[957] , _f_permutation__round__c[958] ,
         _f_permutation__round__c[959] , _f_permutation__round__c[960] ,
         _f_permutation__round__c[961] , _f_permutation__round__c[962] ,
         _f_permutation__round__c[963] , _f_permutation__round__c[964] ,
         _f_permutation__round__c[965] , _f_permutation__round__c[966] ,
         _f_permutation__round__c[967] , _f_permutation__round__c[968] ,
         _f_permutation__round__c[969] , _f_permutation__round__c[970] ,
         _f_permutation__round__c[971] , _f_permutation__round__c[972] ,
         _f_permutation__round__c[973] , _f_permutation__round__c[974] ,
         _f_permutation__round__c[975] , _f_permutation__round__c[976] ,
         _f_permutation__round__c[977] , _f_permutation__round__c[978] ,
         _f_permutation__round__c[979] , _f_permutation__round__c[980] ,
         _f_permutation__round__c[981] , _f_permutation__round__c[982] ,
         _f_permutation__round__c[983] , _f_permutation__round__c[984] ,
         _f_permutation__round__c[985] , _f_permutation__round__c[986] ,
         _f_permutation__round__c[987] , _f_permutation__round__c[988] ,
         _f_permutation__round__c[989] , _f_permutation__round__c[990] ,
         _f_permutation__round__c[991] , _f_permutation__round__c[992] ,
         _f_permutation__round__c[993] , _f_permutation__round__c[994] ,
         _f_permutation__round__c[995] , _f_permutation__round__c[996] ,
         _f_permutation__round__c[997] , _f_permutation__round__c[998] ,
         _f_permutation__round__c[999] , _f_permutation__round__c[1000] ,
         _f_permutation__round__c[1001] , _f_permutation__round__c[1002] ,
         _f_permutation__round__c[1003] , _f_permutation__round__c[1004] ,
         _f_permutation__round__c[1005] , _f_permutation__round__c[1006] ,
         _f_permutation__round__c[1007] , _f_permutation__round__c[1008] ,
         _f_permutation__round__c[1009] , _f_permutation__round__c[1010] ,
         _f_permutation__round__c[1011] , _f_permutation__round__c[1012] ,
         _f_permutation__round__c[1013] , _f_permutation__round__c[1014] ,
         _f_permutation__round__c[1015] , _f_permutation__round__c[1016] ,
         _f_permutation__round__c[1017] , _f_permutation__round__c[1018] ,
         _f_permutation__round__c[1019] , _f_permutation__round__c[1020] ,
         _f_permutation__round__c[1021] , _f_permutation__round__c[1022] ,
         _f_permutation__round__c[1023] , _f_permutation__round__c[1024] ,
         _f_permutation__round__c[1025] , _f_permutation__round__c[1026] ,
         _f_permutation__round__c[1027] , _f_permutation__round__c[1028] ,
         _f_permutation__round__c[1029] , _f_permutation__round__c[1030] ,
         _f_permutation__round__c[1031] , _f_permutation__round__c[1032] ,
         _f_permutation__round__c[1033] , _f_permutation__round__c[1034] ,
         _f_permutation__round__c[1035] , _f_permutation__round__c[1036] ,
         _f_permutation__round__c[1037] , _f_permutation__round__c[1038] ,
         _f_permutation__round__c[1039] , _f_permutation__round__c[1040] ,
         _f_permutation__round__c[1041] , _f_permutation__round__c[1042] ,
         _f_permutation__round__c[1043] , _f_permutation__round__c[1044] ,
         _f_permutation__round__c[1045] , _f_permutation__round__c[1046] ,
         _f_permutation__round__c[1047] , _f_permutation__round__c[1048] ,
         _f_permutation__round__c[1049] , _f_permutation__round__c[1050] ,
         _f_permutation__round__c[1051] , _f_permutation__round__c[1052] ,
         _f_permutation__round__c[1053] , _f_permutation__round__c[1054] ,
         _f_permutation__round__c[1055] , _f_permutation__round__c[1056] ,
         _f_permutation__round__c[1057] , _f_permutation__round__c[1058] ,
         _f_permutation__round__c[1059] , _f_permutation__round__c[1060] ,
         _f_permutation__round__c[1061] , _f_permutation__round__c[1062] ,
         _f_permutation__round__c[1063] , _f_permutation__round__c[1064] ,
         _f_permutation__round__c[1065] , _f_permutation__round__c[1066] ,
         _f_permutation__round__c[1067] , _f_permutation__round__c[1068] ,
         _f_permutation__round__c[1069] , _f_permutation__round__c[1070] ,
         _f_permutation__round__c[1071] , _f_permutation__round__c[1072] ,
         _f_permutation__round__c[1073] , _f_permutation__round__c[1074] ,
         _f_permutation__round__c[1075] , _f_permutation__round__c[1076] ,
         _f_permutation__round__c[1077] , _f_permutation__round__c[1078] ,
         _f_permutation__round__c[1079] , _f_permutation__round__c[1080] ,
         _f_permutation__round__c[1081] , _f_permutation__round__c[1082] ,
         _f_permutation__round__c[1083] , _f_permutation__round__c[1084] ,
         _f_permutation__round__c[1085] , _f_permutation__round__c[1086] ,
         _f_permutation__round__c[1087] , _f_permutation__round__c[1088] ,
         _f_permutation__round__c[1089] , _f_permutation__round__c[1090] ,
         _f_permutation__round__c[1091] , _f_permutation__round__c[1092] ,
         _f_permutation__round__c[1093] , _f_permutation__round__c[1094] ,
         _f_permutation__round__c[1095] , _f_permutation__round__c[1096] ,
         _f_permutation__round__c[1097] , _f_permutation__round__c[1098] ,
         _f_permutation__round__c[1099] , _f_permutation__round__c[1100] ,
         _f_permutation__round__c[1101] , _f_permutation__round__c[1102] ,
         _f_permutation__round__c[1103] , _f_permutation__round__c[1104] ,
         _f_permutation__round__c[1105] , _f_permutation__round__c[1106] ,
         _f_permutation__round__c[1107] , _f_permutation__round__c[1108] ,
         _f_permutation__round__c[1109] , _f_permutation__round__c[1110] ,
         _f_permutation__round__c[1111] , _f_permutation__round__c[1112] ,
         _f_permutation__round__c[1113] , _f_permutation__round__c[1114] ,
         _f_permutation__round__c[1115] , _f_permutation__round__c[1116] ,
         _f_permutation__round__c[1117] , _f_permutation__round__c[1118] ,
         _f_permutation__round__c[1119] , _f_permutation__round__c[1120] ,
         _f_permutation__round__c[1121] , _f_permutation__round__c[1122] ,
         _f_permutation__round__c[1123] , _f_permutation__round__c[1124] ,
         _f_permutation__round__c[1125] , _f_permutation__round__c[1126] ,
         _f_permutation__round__c[1127] , _f_permutation__round__c[1128] ,
         _f_permutation__round__c[1129] , _f_permutation__round__c[1130] ,
         _f_permutation__round__c[1131] , _f_permutation__round__c[1132] ,
         _f_permutation__round__c[1133] , _f_permutation__round__c[1134] ,
         _f_permutation__round__c[1135] , _f_permutation__round__c[1136] ,
         _f_permutation__round__c[1137] , _f_permutation__round__c[1138] ,
         _f_permutation__round__c[1139] , _f_permutation__round__c[1140] ,
         _f_permutation__round__c[1141] , _f_permutation__round__c[1142] ,
         _f_permutation__round__c[1143] , _f_permutation__round__c[1144] ,
         _f_permutation__round__c[1145] , _f_permutation__round__c[1146] ,
         _f_permutation__round__c[1147] , _f_permutation__round__c[1148] ,
         _f_permutation__round__c[1149] , _f_permutation__round__c[1150] ,
         _f_permutation__round__c[1151] , _f_permutation__round__c[1152] ,
         _f_permutation__round__c[1153] , _f_permutation__round__c[1154] ,
         _f_permutation__round__c[1155] , _f_permutation__round__c[1156] ,
         _f_permutation__round__c[1157] , _f_permutation__round__c[1158] ,
         _f_permutation__round__c[1159] , _f_permutation__round__c[1160] ,
         _f_permutation__round__c[1161] , _f_permutation__round__c[1162] ,
         _f_permutation__round__c[1163] , _f_permutation__round__c[1164] ,
         _f_permutation__round__c[1165] , _f_permutation__round__c[1166] ,
         _f_permutation__round__c[1167] , _f_permutation__round__c[1168] ,
         _f_permutation__round__c[1169] , _f_permutation__round__c[1170] ,
         _f_permutation__round__c[1171] , _f_permutation__round__c[1172] ,
         _f_permutation__round__c[1173] , _f_permutation__round__c[1174] ,
         _f_permutation__round__c[1175] , _f_permutation__round__c[1176] ,
         _f_permutation__round__c[1177] , _f_permutation__round__c[1178] ,
         _f_permutation__round__c[1179] , _f_permutation__round__c[1180] ,
         _f_permutation__round__c[1181] , _f_permutation__round__c[1182] ,
         _f_permutation__round__c[1183] , _f_permutation__round__c[1184] ,
         _f_permutation__round__c[1185] , _f_permutation__round__c[1186] ,
         _f_permutation__round__c[1187] , _f_permutation__round__c[1188] ,
         _f_permutation__round__c[1189] , _f_permutation__round__c[1190] ,
         _f_permutation__round__c[1191] , _f_permutation__round__c[1192] ,
         _f_permutation__round__c[1193] , _f_permutation__round__c[1194] ,
         _f_permutation__round__c[1195] , _f_permutation__round__c[1196] ,
         _f_permutation__round__c[1197] , _f_permutation__round__c[1198] ,
         _f_permutation__round__c[1199] , _f_permutation__round__c[1200] ,
         _f_permutation__round__c[1201] , _f_permutation__round__c[1202] ,
         _f_permutation__round__c[1203] , _f_permutation__round__c[1204] ,
         _f_permutation__round__c[1205] , _f_permutation__round__c[1206] ,
         _f_permutation__round__c[1207] , _f_permutation__round__c[1208] ,
         _f_permutation__round__c[1209] , _f_permutation__round__c[1210] ,
         _f_permutation__round__c[1211] , _f_permutation__round__c[1212] ,
         _f_permutation__round__c[1213] , _f_permutation__round__c[1214] ,
         _f_permutation__round__c[1215] , _f_permutation__round__c[1216] ,
         _f_permutation__round__c[1217] , _f_permutation__round__c[1218] ,
         _f_permutation__round__c[1219] , _f_permutation__round__c[1220] ,
         _f_permutation__round__c[1221] , _f_permutation__round__c[1222] ,
         _f_permutation__round__c[1223] , _f_permutation__round__c[1224] ,
         _f_permutation__round__c[1225] , _f_permutation__round__c[1226] ,
         _f_permutation__round__c[1227] , _f_permutation__round__c[1228] ,
         _f_permutation__round__c[1229] , _f_permutation__round__c[1230] ,
         _f_permutation__round__c[1231] , _f_permutation__round__c[1232] ,
         _f_permutation__round__c[1233] , _f_permutation__round__c[1234] ,
         _f_permutation__round__c[1235] , _f_permutation__round__c[1236] ,
         _f_permutation__round__c[1237] , _f_permutation__round__c[1238] ,
         _f_permutation__round__c[1239] , _f_permutation__round__c[1240] ,
         _f_permutation__round__c[1241] , _f_permutation__round__c[1242] ,
         _f_permutation__round__c[1243] , _f_permutation__round__c[1244] ,
         _f_permutation__round__c[1245] , _f_permutation__round__c[1246] ,
         _f_permutation__round__c[1247] , _f_permutation__round__c[1248] ,
         _f_permutation__round__c[1249] , _f_permutation__round__c[1250] ,
         _f_permutation__round__c[1251] , _f_permutation__round__c[1252] ,
         _f_permutation__round__c[1253] , _f_permutation__round__c[1254] ,
         _f_permutation__round__c[1255] , _f_permutation__round__c[1256] ,
         _f_permutation__round__c[1257] , _f_permutation__round__c[1258] ,
         _f_permutation__round__c[1259] , _f_permutation__round__c[1260] ,
         _f_permutation__round__c[1261] , _f_permutation__round__c[1262] ,
         _f_permutation__round__c[1263] , _f_permutation__round__c[1264] ,
         _f_permutation__round__c[1265] , _f_permutation__round__c[1266] ,
         _f_permutation__round__c[1267] , _f_permutation__round__c[1268] ,
         _f_permutation__round__c[1269] , _f_permutation__round__c[1270] ,
         _f_permutation__round__c[1271] , _f_permutation__round__c[1272] ,
         _f_permutation__round__c[1273] , _f_permutation__round__c[1274] ,
         _f_permutation__round__c[1275] , _f_permutation__round__c[1276] ,
         _f_permutation__round__c[1277] , _f_permutation__round__c[1278] ,
         _f_permutation__round__c[1279] , _f_permutation__round__c[1280] ,
         _f_permutation__round__c[1281] , _f_permutation__round__c[1282] ,
         _f_permutation__round__c[1283] , _f_permutation__round__c[1284] ,
         _f_permutation__round__c[1285] , _f_permutation__round__c[1286] ,
         _f_permutation__round__c[1287] , _f_permutation__round__c[1288] ,
         _f_permutation__round__c[1289] , _f_permutation__round__c[1290] ,
         _f_permutation__round__c[1291] , _f_permutation__round__c[1292] ,
         _f_permutation__round__c[1293] , _f_permutation__round__c[1294] ,
         _f_permutation__round__c[1295] , _f_permutation__round__c[1296] ,
         _f_permutation__round__c[1297] , _f_permutation__round__c[1298] ,
         _f_permutation__round__c[1299] , _f_permutation__round__c[1300] ,
         _f_permutation__round__c[1301] , _f_permutation__round__c[1302] ,
         _f_permutation__round__c[1303] , _f_permutation__round__c[1304] ,
         _f_permutation__round__c[1305] , _f_permutation__round__c[1306] ,
         _f_permutation__round__c[1307] , _f_permutation__round__c[1308] ,
         _f_permutation__round__c[1309] , _f_permutation__round__c[1310] ,
         _f_permutation__round__c[1311] , _f_permutation__round__c[1312] ,
         _f_permutation__round__c[1313] , _f_permutation__round__c[1314] ,
         _f_permutation__round__c[1315] , _f_permutation__round__c[1316] ,
         _f_permutation__round__c[1317] , _f_permutation__round__c[1318] ,
         _f_permutation__round__c[1319] , _f_permutation__round__c[1320] ,
         _f_permutation__round__c[1321] , _f_permutation__round__c[1322] ,
         _f_permutation__round__c[1323] , _f_permutation__round__c[1324] ,
         _f_permutation__round__c[1325] , _f_permutation__round__c[1326] ,
         _f_permutation__round__c[1327] , _f_permutation__round__c[1328] ,
         _f_permutation__round__c[1329] , _f_permutation__round__c[1330] ,
         _f_permutation__round__c[1331] , _f_permutation__round__c[1332] ,
         _f_permutation__round__c[1333] , _f_permutation__round__c[1334] ,
         _f_permutation__round__c[1335] , _f_permutation__round__c[1336] ,
         _f_permutation__round__c[1337] , _f_permutation__round__c[1338] ,
         _f_permutation__round__c[1339] , _f_permutation__round__c[1340] ,
         _f_permutation__round__c[1341] , _f_permutation__round__c[1342] ,
         _f_permutation__round__c[1343] , _f_permutation__round__c[1344] ,
         _f_permutation__round__c[1345] , _f_permutation__round__c[1346] ,
         _f_permutation__round__c[1347] , _f_permutation__round__c[1348] ,
         _f_permutation__round__c[1349] , _f_permutation__round__c[1350] ,
         _f_permutation__round__c[1351] , _f_permutation__round__c[1352] ,
         _f_permutation__round__c[1353] , _f_permutation__round__c[1354] ,
         _f_permutation__round__c[1355] , _f_permutation__round__c[1356] ,
         _f_permutation__round__c[1357] , _f_permutation__round__c[1358] ,
         _f_permutation__round__c[1359] , _f_permutation__round__c[1360] ,
         _f_permutation__round__c[1361] , _f_permutation__round__c[1362] ,
         _f_permutation__round__c[1363] , _f_permutation__round__c[1364] ,
         _f_permutation__round__c[1365] , _f_permutation__round__c[1366] ,
         _f_permutation__round__c[1367] , _f_permutation__round__c[1368] ,
         _f_permutation__round__c[1369] , _f_permutation__round__c[1370] ,
         _f_permutation__round__c[1371] , _f_permutation__round__c[1372] ,
         _f_permutation__round__c[1373] , _f_permutation__round__c[1374] ,
         _f_permutation__round__c[1375] , _f_permutation__round__c[1376] ,
         _f_permutation__round__c[1377] , _f_permutation__round__c[1378] ,
         _f_permutation__round__c[1379] , _f_permutation__round__c[1380] ,
         _f_permutation__round__c[1381] , _f_permutation__round__c[1382] ,
         _f_permutation__round__c[1383] , _f_permutation__round__c[1384] ,
         _f_permutation__round__c[1385] , _f_permutation__round__c[1386] ,
         _f_permutation__round__c[1387] , _f_permutation__round__c[1388] ,
         _f_permutation__round__c[1389] , _f_permutation__round__c[1390] ,
         _f_permutation__round__c[1391] , _f_permutation__round__c[1392] ,
         _f_permutation__round__c[1393] , _f_permutation__round__c[1394] ,
         _f_permutation__round__c[1395] , _f_permutation__round__c[1396] ,
         _f_permutation__round__c[1397] , _f_permutation__round__c[1398] ,
         _f_permutation__round__c[1399] , _f_permutation__round__c[1400] ,
         _f_permutation__round__c[1401] , _f_permutation__round__c[1402] ,
         _f_permutation__round__c[1403] , _f_permutation__round__c[1404] ,
         _f_permutation__round__c[1405] , _f_permutation__round__c[1406] ,
         _f_permutation__round__c[1407] , _f_permutation__round__c[1408] ,
         _f_permutation__round__c[1409] , _f_permutation__round__c[1410] ,
         _f_permutation__round__c[1411] , _f_permutation__round__c[1412] ,
         _f_permutation__round__c[1413] , _f_permutation__round__c[1414] ,
         _f_permutation__round__c[1415] , _f_permutation__round__c[1416] ,
         _f_permutation__round__c[1417] , _f_permutation__round__c[1418] ,
         _f_permutation__round__c[1419] , _f_permutation__round__c[1420] ,
         _f_permutation__round__c[1421] , _f_permutation__round__c[1422] ,
         _f_permutation__round__c[1423] , _f_permutation__round__c[1424] ,
         _f_permutation__round__c[1425] , _f_permutation__round__c[1426] ,
         _f_permutation__round__c[1427] , _f_permutation__round__c[1428] ,
         _f_permutation__round__c[1429] , _f_permutation__round__c[1430] ,
         _f_permutation__round__c[1431] , _f_permutation__round__c[1432] ,
         _f_permutation__round__c[1433] , _f_permutation__round__c[1434] ,
         _f_permutation__round__c[1435] , _f_permutation__round__c[1436] ,
         _f_permutation__round__c[1437] , _f_permutation__round__c[1438] ,
         _f_permutation__round__c[1439] , _f_permutation__round__c[1440] ,
         _f_permutation__round__c[1441] , _f_permutation__round__c[1442] ,
         _f_permutation__round__c[1443] , _f_permutation__round__c[1444] ,
         _f_permutation__round__c[1445] , _f_permutation__round__c[1446] ,
         _f_permutation__round__c[1447] , _f_permutation__round__c[1448] ,
         _f_permutation__round__c[1449] , _f_permutation__round__c[1450] ,
         _f_permutation__round__c[1451] , _f_permutation__round__c[1452] ,
         _f_permutation__round__c[1453] , _f_permutation__round__c[1454] ,
         _f_permutation__round__c[1455] , _f_permutation__round__c[1456] ,
         _f_permutation__round__c[1457] , _f_permutation__round__c[1458] ,
         _f_permutation__round__c[1459] , _f_permutation__round__c[1460] ,
         _f_permutation__round__c[1461] , _f_permutation__round__c[1462] ,
         _f_permutation__round__c[1463] , _f_permutation__round__c[1464] ,
         _f_permutation__round__c[1465] , _f_permutation__round__c[1466] ,
         _f_permutation__round__c[1467] , _f_permutation__round__c[1468] ,
         _f_permutation__round__c[1469] , _f_permutation__round__c[1470] ,
         _f_permutation__round__c[1471] , _f_permutation__round__c[1472] ,
         _f_permutation__round__c[1473] , _f_permutation__round__c[1474] ,
         _f_permutation__round__c[1475] , _f_permutation__round__c[1476] ,
         _f_permutation__round__c[1477] , _f_permutation__round__c[1478] ,
         _f_permutation__round__c[1479] , _f_permutation__round__c[1480] ,
         _f_permutation__round__c[1481] , _f_permutation__round__c[1482] ,
         _f_permutation__round__c[1483] , _f_permutation__round__c[1484] ,
         _f_permutation__round__c[1485] , _f_permutation__round__c[1486] ,
         _f_permutation__round__c[1487] , _f_permutation__round__c[1488] ,
         _f_permutation__round__c[1489] , _f_permutation__round__c[1490] ,
         _f_permutation__round__c[1491] , _f_permutation__round__c[1492] ,
         _f_permutation__round__c[1493] , _f_permutation__round__c[1494] ,
         _f_permutation__round__c[1495] , _f_permutation__round__c[1496] ,
         _f_permutation__round__c[1497] , _f_permutation__round__c[1498] ,
         _f_permutation__round__c[1499] , _f_permutation__round__c[1500] ,
         _f_permutation__round__c[1501] , _f_permutation__round__c[1502] ,
         _f_permutation__round__c[1503] , _f_permutation__round__c[1504] ,
         _f_permutation__round__c[1505] , _f_permutation__round__c[1506] ,
         _f_permutation__round__c[1507] , _f_permutation__round__c[1508] ,
         _f_permutation__round__c[1509] , _f_permutation__round__c[1510] ,
         _f_permutation__round__c[1511] , _f_permutation__round__c[1512] ,
         _f_permutation__round__c[1513] , _f_permutation__round__c[1514] ,
         _f_permutation__round__c[1515] , _f_permutation__round__c[1516] ,
         _f_permutation__round__c[1517] , _f_permutation__round__c[1518] ,
         _f_permutation__round__c[1519] , _f_permutation__round__c[1520] ,
         _f_permutation__round__c[1521] , _f_permutation__round__c[1522] ,
         _f_permutation__round__c[1523] , _f_permutation__round__c[1524] ,
         _f_permutation__round__c[1525] , _f_permutation__round__c[1526] ,
         _f_permutation__round__c[1527] , _f_permutation__round__c[1528] ,
         _f_permutation__round__c[1529] , _f_permutation__round__c[1530] ,
         _f_permutation__round__c[1531] , _f_permutation__round__c[1532] ,
         _f_permutation__round__c[1533] , _f_permutation__round__c[1534] ,
         _f_permutation__round__c[1535] , _f_permutation__round__c[1536] ,
         _f_permutation__round__c[1537] , _f_permutation__round__c[1538] ,
         _f_permutation__round__c[1539] , _f_permutation__round__c[1540] ,
         _f_permutation__round__c[1541] , _f_permutation__round__c[1542] ,
         _f_permutation__round__c[1543] , _f_permutation__round__c[1544] ,
         _f_permutation__round__c[1545] , _f_permutation__round__c[1546] ,
         _f_permutation__round__c[1547] , _f_permutation__round__c[1548] ,
         _f_permutation__round__c[1549] , _f_permutation__round__c[1550] ,
         _f_permutation__round__c[1551] , _f_permutation__round__c[1552] ,
         _f_permutation__round__c[1553] , _f_permutation__round__c[1554] ,
         _f_permutation__round__c[1555] , _f_permutation__round__c[1556] ,
         _f_permutation__round__c[1557] , _f_permutation__round__c[1558] ,
         _f_permutation__round__c[1559] , _f_permutation__round__c[1560] ,
         _f_permutation__round__c[1561] , _f_permutation__round__c[1562] ,
         _f_permutation__round__c[1563] , _f_permutation__round__c[1564] ,
         _f_permutation__round__c[1565] , _f_permutation__round__c[1566] ,
         _f_permutation__round__c[1567] , _f_permutation__round__c[1568] ,
         _f_permutation__round__c[1569] , _f_permutation__round__c[1570] ,
         _f_permutation__round__c[1571] , _f_permutation__round__c[1572] ,
         _f_permutation__round__c[1573] , _f_permutation__round__c[1574] ,
         _f_permutation__round__c[1575] , _f_permutation__round__c[1576] ,
         _f_permutation__round__c[1577] , _f_permutation__round__c[1578] ,
         _f_permutation__round__c[1579] , _f_permutation__round__c[1580] ,
         _f_permutation__round__c[1581] , _f_permutation__round__c[1582] ,
         _f_permutation__round__c[1583] , _f_permutation__round__c[1584] ,
         _f_permutation__round__c[1585] , _f_permutation__round__c[1586] ,
         _f_permutation__round__c[1587] , _f_permutation__round__c[1588] ,
         _f_permutation__round__c[1589] , _f_permutation__round__c[1590] ,
         _f_permutation__round__c[1591] , _f_permutation__round__c[1592] ,
         _f_permutation__round__c[1593] , _f_permutation__round__c[1594] ,
         _f_permutation__round__c[1595] , _f_permutation__round__c[1596] ,
         _f_permutation__round__c[1597] , _f_permutation__round__c[1598] ,
         _f_permutation__round__c[1599] , _f_permutation__round__c[0] ,
         _f_permutation__round__c[1] , _f_permutation__round__c[2] ,
         _f_permutation__round__c[3] , _f_permutation__round__c[4] ,
         _f_permutation__round__c[5] , _f_permutation__round__c[6] ,
         _f_permutation__round__c[7] , _f_permutation__round__c[8] ,
         _f_permutation__round__c[9] , _f_permutation__round__c[10] ,
         _f_permutation__round__c[11] , _f_permutation__round__c[12] ,
         _f_permutation__round__c[13] , _f_permutation__round__c[14] ,
         _f_permutation__round__c[15] , _f_permutation__round__c[16] ,
         _f_permutation__round__c[17] , _f_permutation__round__c[18] ,
         _f_permutation__round__c[19] , _f_permutation__round__c[20] ,
         _f_permutation__round__c[21] , _f_permutation__round__c[22] ,
         _f_permutation__round__c[23] , _f_permutation__round__c[24] ,
         _f_permutation__round__c[25] , _f_permutation__round__c[26] ,
         _f_permutation__round__c[27] , _f_permutation__round__c[28] ,
         _f_permutation__round__c[29] , _f_permutation__round__c[30] ,
         _f_permutation__round__c[31] , _f_permutation__round__c[32] ,
         _f_permutation__round__c[33] , _f_permutation__round__c[34] ,
         _f_permutation__round__c[35] , _f_permutation__round__c[36] ,
         _f_permutation__round__c[37] , _f_permutation__round__c[38] ,
         _f_permutation__round__c[39] , _f_permutation__round__c[40] ,
         _f_permutation__round__c[41] , _f_permutation__round__c[42] ,
         _f_permutation__round__c[43] , _f_permutation__round__c[44] ,
         _f_permutation__round__c[45] , _f_permutation__round__c[46] ,
         _f_permutation__round__c[47] , _f_permutation__round__c[48] ,
         _f_permutation__round__c[49] , _f_permutation__round__c[50] ,
         _f_permutation__round__c[51] , _f_permutation__round__c[52] ,
         _f_permutation__round__c[53] , _f_permutation__round__c[54] ,
         _f_permutation__round__c[55] , _f_permutation__round__c[56] ,
         _f_permutation__round__c[57] , _f_permutation__round__c[58] ,
         _f_permutation__round__c[59] , _f_permutation__round__c[60] ,
         _f_permutation__round__c[61] , _f_permutation__round__c[62] ,
         _f_permutation__round__c[63] ;
  wire   [575:0] padder_out;
  wire   [31:0] _padder__v0;
  wire   [1599:0] _f_permutation__round_out;
  wire   [63:0] _f_permutation__rc;
  wire   [1599:1024] _f_permutation__round_in;

  DFF_X2 i_reg_0_ ( .D(n104), .CK(clk), .Q(), .QN(n120) );
  DFF_X2 i_reg_1_ ( .D(n103), .CK(clk), .Q(), .QN(n1100) );
  DFF_X2 i_reg_2_ ( .D(n102), .CK(clk), .Q(), .QN(n1000) );
  DFF_X2 i_reg_3_ ( .D(n101), .CK(clk), .Q(), .QN(n900) );
  DFF_X2 i_reg_4_ ( .D(n1001), .CK(clk), .Q(), .QN(n30) );
  DFF_X2 i_reg_5_ ( .D(n99), .CK(clk), .Q(), .QN(n29) );
  DFF_X2 i_reg_6_ ( .D(n98), .CK(clk), .Q(), .QN(n28) );
  DFF_X2 i_reg_7_ ( .D(n97), .CK(clk), .Q(), .QN(n270) );
  DFF_X2 i_reg_8_ ( .D(n96), .CK(clk), .Q(), .QN(n260) );
  DFF_X2 i_reg_9_ ( .D(n95), .CK(clk), .Q(), .QN(n250) );
  DFF_X2 i_reg_10_ ( .D(n94), .CK(clk), .Q(), .QN(n240) );
  DFF_X2 i_reg_11_ ( .D(n93), .CK(clk), .Q(), .QN(n230) );
  DFF_X2 i_reg_12_ ( .D(n92), .CK(clk), .Q(), .QN(n220) );
  DFF_X2 i_reg_13_ ( .D(n91), .CK(clk), .Q(), .QN(n210) );
  DFF_X2 i_reg_14_ ( .D(n901), .CK(clk), .Q(), .QN(n200) );
  DFF_X2 i_reg_15_ ( .D(n89), .CK(clk), .Q(), .QN(n190) );
  DFF_X2 i_reg_16_ ( .D(n88), .CK(clk), .Q(), .QN(n180) );
  DFF_X2 i_reg_17_ ( .D(n87), .CK(clk), .Q(), .QN(n170) );
  DFF_X2 i_reg_18_ ( .D(n86), .CK(clk), .Q(), .QN(n160) );
  DFF_X2 i_reg_19_ ( .D(n85), .CK(clk), .Q(), .QN(n150) );
  DFF_X2 i_reg_20_ ( .D(n84), .CK(clk), .Q(), .QN(n140) );
  DFF_X2 i_reg_21_ ( .D(n83), .CK(clk), .Q(), .QN(n130) );
  DFF_X1 i_reg_22_ ( .D(n114), .CK(clk), .Q(i_22_), .QN() );
  DFF_X1 out_ready_reg ( .D(n4), .CK(clk), .Q(out_ready), .QN() );
  DFF_X1 state_reg ( .D(n50), .CK(clk), .Q(state), .QN() );
  CLKBUF_X2 U59 ( .A(in[4]), .Z(n59) );
  CLKBUF_X1 U60 ( .A(in[7]), .Z(n60) );
  CLKBUF_X2 U61 ( .A(in[9]), .Z(n61) );
  CLKBUF_X2 U62 ( .A(in[10]), .Z(n62) );
  CLKBUF_X2 U63 ( .A(in[11]), .Z(n63) );
  CLKBUF_X2 U64 ( .A(in[12]), .Z(n64) );
  CLKBUF_X2 U65 ( .A(in[13]), .Z(n65) );
  CLKBUF_X2 U66 ( .A(in[14]), .Z(n66) );
  CLKBUF_X2 U67 ( .A(in[15]), .Z(n67) );
  CLKBUF_X2 U68 ( .A(in[17]), .Z(n68) );
  CLKBUF_X2 U69 ( .A(in[18]), .Z(n69) );
  CLKBUF_X2 U70 ( .A(in[19]), .Z(n70) );
  CLKBUF_X2 U71 ( .A(in[20]), .Z(n71) );
  CLKBUF_X2 U72 ( .A(in[21]), .Z(n72) );
  CLKBUF_X2 U73 ( .A(in[22]), .Z(n73) );
  CLKBUF_X2 U74 ( .A(in[23]), .Z(n74) );
  CLKBUF_X2 U75 ( .A(in[24]), .Z(n75) );
  CLKBUF_X2 U76 ( .A(in[25]), .Z(n76) );
  CLKBUF_X2 U77 ( .A(in[26]), .Z(n77) );
  CLKBUF_X2 U78 ( .A(in[27]), .Z(n78) );
  CLKBUF_X2 U79 ( .A(in[28]), .Z(n79) );
  CLKBUF_X2 U80 ( .A(in[29]), .Z(n80) );
  CLKBUF_X2 U81 ( .A(in[30]), .Z(n81) );
  CLKBUF_X2 U82 ( .A(in[31]), .Z(n82) );
  CLKBUF_X2 U83 ( .A(N26), .Z(n83) );
  CLKBUF_X2 U84 ( .A(N25), .Z(n84) );
  CLKBUF_X2 U85 ( .A(N24), .Z(n85) );
  CLKBUF_X2 U86 ( .A(N23), .Z(n86) );
  CLKBUF_X2 U87 ( .A(N22), .Z(n87) );
  CLKBUF_X2 U88 ( .A(N21), .Z(n88) );
  CLKBUF_X2 U89 ( .A(N20), .Z(n89) );
  CLKBUF_X2 U90 ( .A(N19), .Z(n901) );
  CLKBUF_X2 U91 ( .A(N18), .Z(n91) );
  CLKBUF_X2 U92 ( .A(N17), .Z(n92) );
  CLKBUF_X2 U93 ( .A(N16), .Z(n93) );
  CLKBUF_X2 U94 ( .A(N15), .Z(n94) );
  CLKBUF_X2 U95 ( .A(N14), .Z(n95) );
  CLKBUF_X2 U96 ( .A(N13), .Z(n96) );
  CLKBUF_X2 U97 ( .A(N12), .Z(n97) );
  CLKBUF_X2 U98 ( .A(N11), .Z(n98) );
  CLKBUF_X2 U99 ( .A(N10), .Z(n99) );
  CLKBUF_X2 U100 ( .A(N9), .Z(n1001) );
  CLKBUF_X2 U101 ( .A(N8), .Z(n101) );
  CLKBUF_X2 U102 ( .A(N7), .Z(n102) );
  CLKBUF_X2 U103 ( .A(N6), .Z(n103) );
  CLKBUF_X2 U104 ( .A(N5), .Z(n104) );
  CLKBUF_X1 U105 ( .A(n116), .Z(n105) );
  AND3_X4 U106 ( .A1(f_ack), .A2(n105), .A3(state), .ZN(N5) );
  CLKBUF_X2 U107 ( .A(in[5]), .Z(n106) );
  CLKBUF_X2 U108 ( .A(in[6]), .Z(n107) );
  CLKBUF_X1 U109 ( .A(in[0]), .Z(n108) );
  CLKBUF_X2 U110 ( .A(in[1]), .Z(n109) );
  CLKBUF_X2 U111 ( .A(in[2]), .Z(n1101) );
  CLKBUF_X2 U112 ( .A(in[3]), .Z(n111) );
  CLKBUF_X1 U113 ( .A(is_last), .Z(n113) );
  CLKBUF_X2 U114 ( .A(n113), .Z(n112) );
  NOR2_X1 U115 ( .A1(n112), .A2(state), .ZN(n57) );
  CLKBUF_X2 U116 ( .A(N27), .Z(n114) );
  INV_X1 U117 ( .A(reset), .ZN(n116) );
  INV_X4 U118 ( .A(n116), .ZN(n115) );
  NOR2_X2 U119 ( .A1(n115), .A2(n57), .ZN(n50) );
  NOR2_X2 U120 ( .A1(n115), .A2(n58), .ZN(n4) );
  NOR2_X2 U121 ( .A1(out_ready), .A2(i_22_), .ZN(n58) );
  NOR2_X2 U122 ( .A1(n115), .A2(n130), .ZN(N27) );
  NOR2_X2 U123 ( .A1(n115), .A2(n140), .ZN(N26) );
  NOR2_X2 U124 ( .A1(n115), .A2(n150), .ZN(N25) );
  NOR2_X2 U125 ( .A1(n115), .A2(n160), .ZN(N24) );
  NOR2_X2 U126 ( .A1(n115), .A2(n170), .ZN(N23) );
  NOR2_X2 U127 ( .A1(n115), .A2(n180), .ZN(N22) );
  NOR2_X2 U128 ( .A1(n115), .A2(n190), .ZN(N21) );
  NOR2_X2 U129 ( .A1(n115), .A2(n200), .ZN(N20) );
  NOR2_X2 U130 ( .A1(n115), .A2(n210), .ZN(N19) );
  NOR2_X2 U131 ( .A1(n115), .A2(n220), .ZN(N18) );
  NOR2_X2 U132 ( .A1(n115), .A2(n230), .ZN(N17) );
  NOR2_X2 U133 ( .A1(n115), .A2(n240), .ZN(N16) );
  NOR2_X2 U134 ( .A1(n115), .A2(n250), .ZN(N15) );
  NOR2_X2 U135 ( .A1(n115), .A2(n260), .ZN(N14) );
  NOR2_X2 U136 ( .A1(n115), .A2(n270), .ZN(N13) );
  NOR2_X2 U137 ( .A1(n115), .A2(n28), .ZN(N12) );
  NOR2_X2 U138 ( .A1(n115), .A2(n29), .ZN(N11) );
  NOR2_X2 U139 ( .A1(n115), .A2(n30), .ZN(N10) );
  NOR2_X2 U140 ( .A1(n115), .A2(n900), .ZN(N9) );
  NOR2_X2 U141 ( .A1(n115), .A2(n1000), .ZN(N8) );
  NOR2_X2 U142 ( .A1(n115), .A2(n1100), .ZN(N7) );
  NOR2_X2 U143 ( .A1(n115), .A2(n120), .ZN(N6) );
  BUF_X4 _padder__U1945  ( .A(padder_out_ready), .Z(buffer_full) );
  NOR2_X2 _padder__U1944  ( .A1(_padder__n1961 ), .A2(_padder__n598 ), .ZN(
        _padder__n623 ) );
  NOR2_X2 _padder__U1943  ( .A1(_padder__n623 ), .A2(_padder__n602 ), .ZN(
        _padder__n622 ) );
  NOR2_X2 _padder__U1942  ( .A1(n115), .A2(_padder__n622 ), .ZN(
        _padder__n1835 ) );
  NAND3_X2 _padder__U1941  ( .A1(_padder__n2484 ), .A2(_padder__n598 ), .A3(
        n112), .ZN(_padder__n682 ) );
  NOR2_X2 _padder__U1940  ( .A1(n112), .A2(_padder__state ), .ZN(
        _padder__n621 ) );
  NOR2_X2 _padder__U1939  ( .A1(n115), .A2(_padder__n621 ), .ZN(
        _padder__n1836 ) );
  NOR2_X2 _padder__U1938  ( .A1(in_ready), .A2(_padder__state ), .ZN(
        _padder__n2442 ) );
  OR3_X2 _padder__U1937  ( .A1(n112), .A2(_padder__state ), .A3(
        _padder__n2444 ), .ZN(_padder__n2480 ) );
  INV_X4 _padder__U1936  ( .A(_padder__n2480 ), .ZN(_padder__n2510 ) );
  INV_X4 _padder__U1935  ( .A(_padder__n2480 ), .ZN(_padder__n2509 ) );
  INV_X4 _padder__U1934  ( .A(_padder__n2480 ), .ZN(_padder__n2508 ) );
  INV_X4 _padder__U1933  ( .A(_padder__n2444 ), .ZN(_padder__n2483 ) );
  INV_X4 _padder__U1932  ( .A(_padder__n682 ), .ZN(_padder__n2571 ) );
  INV_X4 _padder__U1931  ( .A(_padder__n682 ), .ZN(_padder__n2570 ) );
  INV_X4 _padder__U1930  ( .A(_padder__n2483 ), .ZN(_padder__n2506 ) );
  INV_X4 _padder__U1929  ( .A(_padder__n2483 ), .ZN(_padder__n2507 ) );
  INV_X4 _padder__U1928  ( .A(_padder__n2479 ), .ZN(_padder__n2482 ) );
  INV_X4 _padder__U1927  ( .A(_padder__n2506 ), .ZN(_padder__n2505 ) );
  INV_X4 _padder__U1926  ( .A(_padder__n2444 ), .ZN(_padder__n2484 ) );
  INV_X4 _padder__U1925  ( .A(_padder__n2507 ), .ZN(_padder__n2485 ) );
  INV_X4 _padder__U1924  ( .A(_padder__n2507 ), .ZN(_padder__n2486 ) );
  INV_X4 _padder__U1923  ( .A(_padder__n2506 ), .ZN(_padder__n2487 ) );
  INV_X4 _padder__U1922  ( .A(_padder__n2506 ), .ZN(_padder__n2490 ) );
  INV_X4 _padder__U1921  ( .A(_padder__n2506 ), .ZN(_padder__n2491 ) );
  INV_X4 _padder__U1920  ( .A(_padder__n2506 ), .ZN(_padder__n2492 ) );
  INV_X4 _padder__U1919  ( .A(_padder__n2506 ), .ZN(_padder__n2494 ) );
  INV_X4 _padder__U1918  ( .A(_padder__n2506 ), .ZN(_padder__n2488 ) );
  INV_X4 _padder__U1917  ( .A(_padder__n2507 ), .ZN(_padder__n2500 ) );
  INV_X4 _padder__U1916  ( .A(_padder__n2507 ), .ZN(_padder__n2502 ) );
  INV_X4 _padder__U1915  ( .A(_padder__n2506 ), .ZN(_padder__n2503 ) );
  INV_X4 _padder__U1914  ( .A(_padder__n2506 ), .ZN(_padder__n2504 ) );
  INV_X4 _padder__U1913  ( .A(_padder__n2507 ), .ZN(_padder__n2496 ) );
  INV_X4 _padder__U1912  ( .A(_padder__n2507 ), .ZN(_padder__n2497 ) );
  INV_X4 _padder__U1911  ( .A(_padder__n2507 ), .ZN(_padder__n2498 ) );
  INV_X4 _padder__U1910  ( .A(_padder__n2507 ), .ZN(_padder__n2489 ) );
  INV_X4 _padder__U1909  ( .A(_padder__n2507 ), .ZN(_padder__n2493 ) );
  INV_X4 _padder__U1908  ( .A(_padder__n2506 ), .ZN(_padder__n2501 ) );
  INV_X4 _padder__U1907  ( .A(_padder__n2506 ), .ZN(_padder__n2495 ) );
  INV_X4 _padder__U1906  ( .A(_padder__n2507 ), .ZN(_padder__n2499 ) );
  INV_X4 _padder__U1905  ( .A(_padder__n2443 ), .ZN(_padder__n2569 ) );
  INV_X4 _padder__U1904  ( .A(_padder__n2569 ), .ZN(_padder__n2563 ) );
  INV_X4 _padder__U1903  ( .A(_padder__n2569 ), .ZN(_padder__n2564 ) );
  INV_X4 _padder__U1902  ( .A(_padder__n2517 ), .ZN(_padder__n2565 ) );
  INV_X4 _padder__U1901  ( .A(_padder__n2569 ), .ZN(_padder__n2566 ) );
  INV_X4 _padder__U1900  ( .A(_padder__n2518 ), .ZN(_padder__n2567 ) );
  INV_X4 _padder__U1899  ( .A(_padder__n2539 ), .ZN(_padder__n2568 ) );
  INV_X4 _padder__U1898  ( .A(_padder__n2564 ), .ZN(_padder__n2511 ) );
  INV_X4 _padder__U1897  ( .A(_padder__n2564 ), .ZN(_padder__n2512 ) );
  INV_X4 _padder__U1896  ( .A(_padder__n2566 ), .ZN(_padder__n2560 ) );
  INV_X4 _padder__U1895  ( .A(_padder__n2563 ), .ZN(_padder__n2557 ) );
  INV_X4 _padder__U1894  ( .A(_padder__n2565 ), .ZN(_padder__n2554 ) );
  INV_X4 _padder__U1893  ( .A(_padder__n2563 ), .ZN(_padder__n2551 ) );
  INV_X4 _padder__U1892  ( .A(_padder__n2564 ), .ZN(_padder__n2548 ) );
  INV_X4 _padder__U1891  ( .A(_padder__n2563 ), .ZN(_padder__n2545 ) );
  INV_X4 _padder__U1890  ( .A(_padder__n2568 ), .ZN(_padder__n2543 ) );
  INV_X4 _padder__U1889  ( .A(_padder__n2565 ), .ZN(_padder__n2540 ) );
  INV_X4 _padder__U1888  ( .A(_padder__n2563 ), .ZN(_padder__n2537 ) );
  INV_X4 _padder__U1887  ( .A(_padder__n2567 ), .ZN(_padder__n2534 ) );
  INV_X4 _padder__U1886  ( .A(_padder__n2566 ), .ZN(_padder__n2531 ) );
  INV_X4 _padder__U1885  ( .A(_padder__n2567 ), .ZN(_padder__n2528 ) );
  INV_X4 _padder__U1884  ( .A(_padder__n2563 ), .ZN(_padder__n2525 ) );
  INV_X4 _padder__U1883  ( .A(_padder__n2568 ), .ZN(_padder__n2522 ) );
  INV_X4 _padder__U1882  ( .A(_padder__n2564 ), .ZN(_padder__n2519 ) );
  INV_X4 _padder__U1881  ( .A(_padder__n2563 ), .ZN(_padder__n2516 ) );
  INV_X4 _padder__U1880  ( .A(_padder__n2564 ), .ZN(_padder__n2513 ) );
  INV_X4 _padder__U1879  ( .A(_padder__n2564 ), .ZN(_padder__n2546 ) );
  INV_X4 _padder__U1878  ( .A(_padder__n2564 ), .ZN(_padder__n2514 ) );
  INV_X4 _padder__U1877  ( .A(_padder__n2563 ), .ZN(_padder__n2549 ) );
  INV_X4 _padder__U1876  ( .A(_padder__n2566 ), .ZN(_padder__n2517 ) );
  INV_X4 _padder__U1875  ( .A(_padder__n2563 ), .ZN(_padder__n2552 ) );
  INV_X4 _padder__U1874  ( .A(_padder__n2563 ), .ZN(_padder__n2520 ) );
  INV_X4 _padder__U1873  ( .A(_padder__n2564 ), .ZN(_padder__n2555 ) );
  INV_X4 _padder__U1872  ( .A(_padder__n2568 ), .ZN(_padder__n2523 ) );
  INV_X4 _padder__U1871  ( .A(_padder__n2565 ), .ZN(_padder__n2558 ) );
  INV_X4 _padder__U1870  ( .A(_padder__n2568 ), .ZN(_padder__n2526 ) );
  INV_X4 _padder__U1869  ( .A(_padder__n2443 ), .ZN(_padder__n2561 ) );
  INV_X4 _padder__U1868  ( .A(_padder__n2567 ), .ZN(_padder__n2529 ) );
  INV_X4 _padder__U1867  ( .A(_padder__n2566 ), .ZN(_padder__n2532 ) );
  INV_X4 _padder__U1866  ( .A(_padder__n2566 ), .ZN(_padder__n2535 ) );
  INV_X4 _padder__U1865  ( .A(_padder__n2566 ), .ZN(_padder__n2538 ) );
  INV_X4 _padder__U1864  ( .A(_padder__n2565 ), .ZN(_padder__n2541 ) );
  INV_X4 _padder__U1863  ( .A(_padder__n2568 ), .ZN(_padder__n2544 ) );
  INV_X4 _padder__U1862  ( .A(_padder__n2564 ), .ZN(_padder__n2547 ) );
  INV_X4 _padder__U1861  ( .A(_padder__n2563 ), .ZN(_padder__n2515 ) );
  INV_X4 _padder__U1860  ( .A(_padder__n2563 ), .ZN(_padder__n2550 ) );
  INV_X4 _padder__U1859  ( .A(_padder__n2566 ), .ZN(_padder__n2518 ) );
  INV_X4 _padder__U1858  ( .A(_padder__n2564 ), .ZN(_padder__n2553 ) );
  INV_X4 _padder__U1857  ( .A(_padder__n2564 ), .ZN(_padder__n2521 ) );
  INV_X4 _padder__U1856  ( .A(_padder__n2563 ), .ZN(_padder__n2556 ) );
  INV_X4 _padder__U1855  ( .A(_padder__n2568 ), .ZN(_padder__n2524 ) );
  INV_X4 _padder__U1854  ( .A(_padder__n2564 ), .ZN(_padder__n2559 ) );
  INV_X4 _padder__U1853  ( .A(_padder__n2564 ), .ZN(_padder__n2527 ) );
  INV_X4 _padder__U1852  ( .A(_padder__n2443 ), .ZN(_padder__n2562 ) );
  INV_X4 _padder__U1851  ( .A(_padder__n2567 ), .ZN(_padder__n2530 ) );
  INV_X4 _padder__U1850  ( .A(_padder__n2566 ), .ZN(_padder__n2533 ) );
  INV_X4 _padder__U1849  ( .A(_padder__n2567 ), .ZN(_padder__n2536 ) );
  INV_X4 _padder__U1848  ( .A(_padder__n2566 ), .ZN(_padder__n2539 ) );
  INV_X4 _padder__U1847  ( .A(_padder__n2565 ), .ZN(_padder__n2542 ) );
  OR2_X2 _padder__U1846  ( .A1(_padder__n2444 ), .A2(f_ack), .ZN(
        _padder__n2479 ) );
  NAND2_X1 _padder__U1845  ( .A1(n111), .A2(_padder__n2508 ), .ZN(
        _padder__n671 ) );
  BUF_X16 _padder__U1844  ( .A(_padder__n671 ), .Z(_padder__n2478 ) );
  NAND2_X1 _padder__U1843  ( .A1(n1101), .A2(_padder__n2508 ), .ZN(
        _padder__n669 ) );
  BUF_X16 _padder__U1842  ( .A(_padder__n669 ), .Z(_padder__n2477 ) );
  NAND2_X1 _padder__U1841  ( .A1(n109), .A2(_padder__n2508 ), .ZN(
        _padder__n667 ) );
  BUF_X16 _padder__U1840  ( .A(_padder__n667 ), .Z(_padder__n2476 ) );
  NAND2_X1 _padder__U1839  ( .A1(n108), .A2(_padder__n2508 ), .ZN(
        _padder__n663 ) );
  NAND3_X1 _padder__U1838  ( .A1(_padder__n662 ), .A2(_padder__n663 ), .A3(
        _padder__n664 ), .ZN(_padder__n1816 ) );
  CLKBUF_X1 _padder__U1837  ( .A(_padder__n1816 ), .Z(_padder__n2475 ) );
  NAND2_X1 _padder__U1836  ( .A1(n107), .A2(_padder__n2508 ), .ZN(
        _padder__n677 ) );
  BUF_X16 _padder__U1835  ( .A(_padder__n677 ), .Z(_padder__n2474 ) );
  NAND2_X1 _padder__U1834  ( .A1(n106), .A2(_padder__n2508 ), .ZN(
        _padder__n675 ) );
  BUF_X16 _padder__U1833  ( .A(_padder__n675 ), .Z(_padder__n2473 ) );
  NAND2_X1 _padder__U1832  ( .A1(n82), .A2(_padder__n2510 ), .ZN(
        _padder__n755 ) );
  NAND3_X1 _padder__U1831  ( .A1(_padder__n754 ), .A2(_padder__n755 ), .A3(
        _padder__n756 ), .ZN(_padder__n1785 ) );
  CLKBUF_X1 _padder__U1830  ( .A(_padder__n1785 ), .Z(_padder__n2472 ) );
  NAND2_X1 _padder__U1829  ( .A1(n81), .A2(_padder__n2510 ), .ZN(
        _padder__n752 ) );
  NAND3_X1 _padder__U1828  ( .A1(_padder__n751 ), .A2(_padder__n752 ), .A3(
        _padder__n753 ), .ZN(_padder__n1786 ) );
  CLKBUF_X1 _padder__U1827  ( .A(_padder__n1786 ), .Z(_padder__n2471 ) );
  NAND2_X1 _padder__U1826  ( .A1(n80), .A2(_padder__n2510 ), .ZN(
        _padder__n749 ) );
  NAND3_X1 _padder__U1825  ( .A1(_padder__n748 ), .A2(_padder__n749 ), .A3(
        _padder__n750 ), .ZN(_padder__n1787 ) );
  CLKBUF_X1 _padder__U1824  ( .A(_padder__n1787 ), .Z(_padder__n2470 ) );
  NAND2_X1 _padder__U1823  ( .A1(n79), .A2(_padder__n2510 ), .ZN(
        _padder__n746 ) );
  NAND3_X1 _padder__U1822  ( .A1(_padder__n745 ), .A2(_padder__n746 ), .A3(
        _padder__n747 ), .ZN(_padder__n1788 ) );
  CLKBUF_X1 _padder__U1821  ( .A(_padder__n1788 ), .Z(_padder__n2469 ) );
  NAND2_X1 _padder__U1819  ( .A1(n78), .A2(_padder__n2510 ), .ZN(
        _padder__n743 ) );
  NAND3_X1 _padder__U187  ( .A1(_padder__n742 ), .A2(_padder__n743 ), .A3(
        _padder__n744 ), .ZN(_padder__n1789 ) );
  CLKBUF_X1 _padder__U185  ( .A(_padder__n1789 ), .Z(_padder__n2468 ) );
  NAND2_X1 _padder__U184  ( .A1(n77), .A2(_padder__n2510 ), .ZN(_padder__n740 ) );
  NAND3_X1 _padder__U182  ( .A1(_padder__n739 ), .A2(_padder__n740 ), .A3(
        _padder__n741 ), .ZN(_padder__n1790 ) );
  CLKBUF_X1 _padder__U180  ( .A(_padder__n1790 ), .Z(_padder__n2467 ) );
  NAND2_X1 _padder__U178  ( .A1(n76), .A2(_padder__n2510 ), .ZN(_padder__n737 ) );
  NAND3_X1 _padder__U176  ( .A1(_padder__n736 ), .A2(_padder__n737 ), .A3(
        _padder__n738 ), .ZN(_padder__n1791 ) );
  CLKBUF_X1 _padder__U174  ( .A(_padder__n1791 ), .Z(_padder__n2466 ) );
  NAND2_X1 _padder__U172  ( .A1(n75), .A2(_padder__n2510 ), .ZN(_padder__n734 ) );
  CLKBUF_X2 _padder__U170  ( .A(_padder__n1792 ), .Z(_padder__n2465 ) );
  NAND3_X1 _padder__U168  ( .A1(_padder__n733 ), .A2(_padder__n734 ), .A3(
        _padder__n735 ), .ZN(_padder__n1792 ) );
  NAND2_X1 _padder__U166  ( .A1(n74), .A2(_padder__n2510 ), .ZN(_padder__n731 ) );
  CLKBUF_X2 _padder__U164  ( .A(_padder__n1793 ), .Z(_padder__n2464 ) );
  NAND3_X1 _padder__U162  ( .A1(_padder__n730 ), .A2(_padder__n731 ), .A3(
        _padder__n732 ), .ZN(_padder__n1793 ) );
  NAND2_X1 _padder__U160  ( .A1(n73), .A2(_padder__n2510 ), .ZN(_padder__n728 ) );
  CLKBUF_X2 _padder__U158  ( .A(_padder__n1794 ), .Z(_padder__n2463 ) );
  NAND3_X1 _padder__U156  ( .A1(_padder__n727 ), .A2(_padder__n728 ), .A3(
        _padder__n729 ), .ZN(_padder__n1794 ) );
  NAND2_X1 _padder__U154  ( .A1(n72), .A2(_padder__n2509 ), .ZN(_padder__n725 ) );
  CLKBUF_X2 _padder__U152  ( .A(_padder__n1795 ), .Z(_padder__n2462 ) );
  NAND3_X1 _padder__U150  ( .A1(_padder__n724 ), .A2(_padder__n725 ), .A3(
        _padder__n726 ), .ZN(_padder__n1795 ) );
  NAND2_X1 _padder__U148  ( .A1(n71), .A2(_padder__n2509 ), .ZN(_padder__n722 ) );
  CLKBUF_X2 _padder__U146  ( .A(_padder__n1796 ), .Z(_padder__n2461 ) );
  NAND3_X1 _padder__U144  ( .A1(_padder__n721 ), .A2(_padder__n722 ), .A3(
        _padder__n723 ), .ZN(_padder__n1796 ) );
  NAND2_X1 _padder__U142  ( .A1(n70), .A2(_padder__n2509 ), .ZN(_padder__n719 ) );
  CLKBUF_X2 _padder__U140  ( .A(_padder__n1797 ), .Z(_padder__n2460 ) );
  NAND3_X1 _padder__U138  ( .A1(_padder__n718 ), .A2(_padder__n719 ), .A3(
        _padder__n720 ), .ZN(_padder__n1797 ) );
  NAND2_X1 _padder__U136  ( .A1(n69), .A2(_padder__n2509 ), .ZN(_padder__n716 ) );
  CLKBUF_X2 _padder__U134  ( .A(_padder__n1798 ), .Z(_padder__n2459 ) );
  NAND3_X1 _padder__U132  ( .A1(_padder__n715 ), .A2(_padder__n716 ), .A3(
        _padder__n717 ), .ZN(_padder__n1798 ) );
  NAND2_X1 _padder__U130  ( .A1(n68), .A2(_padder__n2509 ), .ZN(_padder__n713 ) );
  CLKBUF_X2 _padder__U128  ( .A(_padder__n1799 ), .Z(_padder__n2458 ) );
  NAND3_X1 _padder__U126  ( .A1(_padder__n712 ), .A2(_padder__n713 ), .A3(
        _padder__n714 ), .ZN(_padder__n1799 ) );
  NAND2_X1 _padder__U124  ( .A1(in[16]), .A2(_padder__n2509 ), .ZN(
        _padder__n710 ) );
  NAND3_X1 _padder__U122  ( .A1(_padder__n709 ), .A2(_padder__n710 ), .A3(
        _padder__n711 ), .ZN(_padder__n1800 ) );
  BUF_X32 _padder__U120  ( .A(_padder__n1800 ), .Z(_padder__n2457 ) );
  NAND2_X1 _padder__U118  ( .A1(n67), .A2(_padder__n2509 ), .ZN(_padder__n707 ) );
  NAND3_X1 _padder__U116  ( .A1(_padder__n706 ), .A2(_padder__n707 ), .A3(
        _padder__n708 ), .ZN(_padder__n1801 ) );
  CLKBUF_X1 _padder__U114  ( .A(_padder__n1801 ), .Z(_padder__n2456 ) );
  NAND2_X1 _padder__U112  ( .A1(n66), .A2(_padder__n2509 ), .ZN(_padder__n704 ) );
  NAND3_X1 _padder__U110  ( .A1(_padder__n703 ), .A2(_padder__n704 ), .A3(
        _padder__n705 ), .ZN(_padder__n1802 ) );
  CLKBUF_X1 _padder__U108  ( .A(_padder__n1802 ), .Z(_padder__n2455 ) );
  NAND2_X1 _padder__U106  ( .A1(n65), .A2(_padder__n2509 ), .ZN(_padder__n701 ) );
  NAND3_X1 _padder__U104  ( .A1(_padder__n700 ), .A2(_padder__n701 ), .A3(
        _padder__n702 ), .ZN(_padder__n1803 ) );
  CLKBUF_X1 _padder__U102  ( .A(_padder__n1803 ), .Z(_padder__n2454 ) );
  NAND2_X1 _padder__U100  ( .A1(n64), .A2(_padder__n2509 ), .ZN(_padder__n698 ) );
  NAND3_X1 _padder__U98  ( .A1(_padder__n697 ), .A2(_padder__n698 ), .A3(
        _padder__n699 ), .ZN(_padder__n1804 ) );
  CLKBUF_X1 _padder__U96  ( .A(_padder__n1804 ), .Z(_padder__n2453 ) );
  NAND2_X1 _padder__U94  ( .A1(n63), .A2(_padder__n2509 ), .ZN(_padder__n695 )
         );
  NAND3_X1 _padder__U92  ( .A1(_padder__n694 ), .A2(_padder__n695 ), .A3(
        _padder__n696 ), .ZN(_padder__n1805 ) );
  CLKBUF_X1 _padder__U90  ( .A(_padder__n1805 ), .Z(_padder__n2452 ) );
  NAND2_X1 _padder__U89  ( .A1(n62), .A2(_padder__n2508 ), .ZN(_padder__n692 )
         );
  NAND3_X1 _padder__U84  ( .A1(_padder__n691 ), .A2(_padder__n692 ), .A3(
        _padder__n693 ), .ZN(_padder__n1806 ) );
  CLKBUF_X1 _padder__U82  ( .A(_padder__n1806 ), .Z(_padder__n2451 ) );
  NAND2_X1 _padder__U79  ( .A1(n61), .A2(_padder__n2508 ), .ZN(_padder__n689 )
         );
  NAND3_X1 _padder__U76  ( .A1(_padder__n688 ), .A2(_padder__n689 ), .A3(
        _padder__n690 ), .ZN(_padder__n1807 ) );
  CLKBUF_X1 _padder__U73  ( .A(_padder__n1807 ), .Z(_padder__n2450 ) );
  NAND2_X1 _padder__U70  ( .A1(in[8]), .A2(_padder__n2508 ), .ZN(
        _padder__n686 ) );
  NAND3_X1 _padder__U67  ( .A1(_padder__n685 ), .A2(_padder__n686 ), .A3(
        _padder__n687 ), .ZN(_padder__n1808 ) );
  BUF_X32 _padder__U64  ( .A(_padder__n1808 ), .Z(_padder__n2449 ) );
  NAND2_X1 _padder__U62  ( .A1(n60), .A2(_padder__n2508 ), .ZN(_padder__n678 )
         );
  INV_X4 _padder__U61  ( .A(_padder__n2446 ), .ZN(_padder__n2448 ) );
  NAND2_X1 _padder__U59  ( .A1(n59), .A2(_padder__n2508 ), .ZN(_padder__n673 )
         );
  BUF_X16 _padder__U6  ( .A(_padder__n673 ), .Z(_padder__n2447 ) );
  AND3_X4 _padder__U5  ( .A1(_padder__n678 ), .A2(_padder__n679 ), .A3(
        _padder__n680 ), .ZN(_padder__n2446 ) );
  NOR2_X2 _padder__U4  ( .A1(_padder__n2443 ), .A2(f_ack), .ZN(_padder__n2445 ) );
  OR4_X4 _padder__U3  ( .A1(_padder__n602 ), .A2(padder_out_ready), .A3(n115), 
        .A4(_padder__n2442 ), .ZN(_padder__n2444 ) );
  OR2_X4 _padder__U2  ( .A1(_padder__n2484 ), .A2(n115), .ZN(_padder__n2443 )
         );
  DFF_X1 _padder__out_reg_524_  ( .D(_padder__n1292 ), .CK(clk), .Q(
        padder_out[564]), .QN() );
  DFF_X1 _padder__out_reg_525_  ( .D(_padder__n1291 ), .CK(clk), .Q(
        padder_out[565]), .QN() );
  DFF_X1 _padder__out_reg_526_  ( .D(_padder__n1290 ), .CK(clk), .Q(
        padder_out[566]), .QN() );
  DFF_X1 _padder__out_reg_527_  ( .D(_padder__n1289 ), .CK(clk), .Q(
        padder_out[567]), .QN() );
  DFF_X1 _padder__out_reg_528_  ( .D(_padder__n1288 ), .CK(clk), .Q(
        padder_out[552]), .QN() );
  DFF_X1 _padder__out_reg_529_  ( .D(_padder__n1287 ), .CK(clk), .Q(
        padder_out[553]), .QN() );
  DFF_X1 _padder__out_reg_530_  ( .D(_padder__n1286 ), .CK(clk), .Q(
        padder_out[554]), .QN() );
  DFF_X1 _padder__out_reg_531_  ( .D(_padder__n1285 ), .CK(clk), .Q(
        padder_out[555]), .QN() );
  DFF_X1 _padder__out_reg_532_  ( .D(_padder__n1284 ), .CK(clk), .Q(
        padder_out[556]), .QN() );
  DFF_X1 _padder__out_reg_533_  ( .D(_padder__n1283 ), .CK(clk), .Q(
        padder_out[557]), .QN() );
  DFF_X1 _padder__out_reg_534_  ( .D(_padder__n1282 ), .CK(clk), .Q(
        padder_out[558]), .QN() );
  DFF_X1 _padder__out_reg_535_  ( .D(_padder__n1281 ), .CK(clk), .Q(
        padder_out[559]), .QN() );
  DFF_X1 _padder__out_reg_536_  ( .D(_padder__n1280 ), .CK(clk), .Q(
        padder_out[544]), .QN() );
  DFF_X1 _padder__out_reg_537_  ( .D(_padder__n1279 ), .CK(clk), .Q(
        padder_out[545]), .QN() );
  DFF_X1 _padder__out_reg_538_  ( .D(_padder__n1278 ), .CK(clk), .Q(
        padder_out[546]), .QN() );
  DFF_X1 _padder__out_reg_539_  ( .D(_padder__n1277 ), .CK(clk), .Q(
        padder_out[547]), .QN() );
  DFF_X1 _padder__out_reg_540_  ( .D(_padder__n1276 ), .CK(clk), .Q(
        padder_out[548]), .QN() );
  DFF_X1 _padder__out_reg_541_  ( .D(_padder__n1275 ), .CK(clk), .Q(
        padder_out[549]), .QN() );
  DFF_X1 _padder__out_reg_542_  ( .D(_padder__n1274 ), .CK(clk), .Q(
        padder_out[550]), .QN() );
  DFF_X1 _padder__out_reg_543_  ( .D(_padder__n1273 ), .CK(clk), .Q(
        padder_out[551]), .QN() );
  DFF_X1 _padder__out_reg_544_  ( .D(_padder__n1272 ), .CK(clk), .Q(
        padder_out[536]), .QN() );
  DFF_X1 _padder__out_reg_545_  ( .D(_padder__n1271 ), .CK(clk), .Q(
        padder_out[537]), .QN() );
  DFF_X1 _padder__out_reg_546_  ( .D(_padder__n1270 ), .CK(clk), .Q(
        padder_out[538]), .QN() );
  DFF_X1 _padder__out_reg_547_  ( .D(_padder__n1269 ), .CK(clk), .Q(
        padder_out[539]), .QN() );
  DFF_X1 _padder__out_reg_548_  ( .D(_padder__n1268 ), .CK(clk), .Q(
        padder_out[540]), .QN() );
  DFF_X1 _padder__out_reg_549_  ( .D(_padder__n1267 ), .CK(clk), .Q(
        padder_out[541]), .QN() );
  DFF_X1 _padder__out_reg_550_  ( .D(_padder__n1266 ), .CK(clk), .Q(
        padder_out[542]), .QN() );
  DFF_X1 _padder__out_reg_551_  ( .D(_padder__n1265 ), .CK(clk), .Q(
        padder_out[543]), .QN() );
  DFF_X1 _padder__out_reg_552_  ( .D(_padder__n1264 ), .CK(clk), .Q(
        padder_out[528]), .QN() );
  DFF_X1 _padder__out_reg_553_  ( .D(_padder__n1263 ), .CK(clk), .Q(
        padder_out[529]), .QN() );
  DFF_X1 _padder__out_reg_554_  ( .D(_padder__n1262 ), .CK(clk), .Q(
        padder_out[530]), .QN() );
  DFF_X1 _padder__out_reg_555_  ( .D(_padder__n1261 ), .CK(clk), .Q(
        padder_out[531]), .QN() );
  DFF_X1 _padder__out_reg_556_  ( .D(_padder__n1260 ), .CK(clk), .Q(
        padder_out[532]), .QN() );
  DFF_X1 _padder__out_reg_557_  ( .D(_padder__n1259 ), .CK(clk), .Q(
        padder_out[533]), .QN() );
  DFF_X1 _padder__out_reg_558_  ( .D(_padder__n1258 ), .CK(clk), .Q(
        padder_out[534]), .QN() );
  DFF_X1 _padder__out_reg_559_  ( .D(_padder__n1257 ), .CK(clk), .Q(
        padder_out[535]), .QN() );
  DFF_X1 _padder__out_reg_560_  ( .D(_padder__n1256 ), .CK(clk), .Q(
        padder_out[520]), .QN() );
  DFF_X1 _padder__out_reg_561_  ( .D(_padder__n1255 ), .CK(clk), .Q(
        padder_out[521]), .QN() );
  DFF_X1 _padder__out_reg_562_  ( .D(_padder__n1254 ), .CK(clk), .Q(
        padder_out[522]), .QN() );
  DFF_X1 _padder__out_reg_563_  ( .D(_padder__n1253 ), .CK(clk), .Q(
        padder_out[523]), .QN() );
  DFF_X1 _padder__out_reg_564_  ( .D(_padder__n1252 ), .CK(clk), .Q(
        padder_out[524]), .QN() );
  DFF_X1 _padder__out_reg_565_  ( .D(_padder__n1251 ), .CK(clk), .Q(
        padder_out[525]), .QN() );
  DFF_X1 _padder__out_reg_566_  ( .D(_padder__n1250 ), .CK(clk), .Q(
        padder_out[526]), .QN() );
  DFF_X1 _padder__out_reg_567_  ( .D(_padder__n1249 ), .CK(clk), .Q(
        padder_out[527]), .QN() );
  DFF_X1 _padder__out_reg_568_  ( .D(_padder__n1248 ), .CK(clk), .Q(
        padder_out[512]), .QN() );
  DFF_X1 _padder__out_reg_569_  ( .D(_padder__n1247 ), .CK(clk), .Q(
        padder_out[513]), .QN() );
  DFF_X1 _padder__out_reg_570_  ( .D(_padder__n1246 ), .CK(clk), .Q(
        padder_out[514]), .QN() );
  DFF_X1 _padder__out_reg_571_  ( .D(_padder__n1245 ), .CK(clk), .Q(
        padder_out[515]), .QN() );
  DFF_X1 _padder__out_reg_572_  ( .D(_padder__n1244 ), .CK(clk), .Q(
        padder_out[516]), .QN() );
  DFF_X1 _padder__out_reg_573_  ( .D(_padder__n1243 ), .CK(clk), .Q(
        padder_out[517]), .QN() );
  DFF_X1 _padder__out_reg_574_  ( .D(_padder__n1242 ), .CK(clk), .Q(
        padder_out[518]), .QN() );
  DFF_X1 _padder__out_reg_575_  ( .D(_padder__n1241 ), .CK(clk), .Q(
        padder_out[519]), .QN() );
  DFF_X1 _padder__out_reg_4_  ( .D(_padder__n1812 ), .CK(clk), .Q(
        padder_out[60]), .QN() );
  DFF_X1 _padder__out_reg_5_  ( .D(_padder__n1811 ), .CK(clk), .Q(
        padder_out[61]), .QN() );
  DFF_X1 _padder__out_reg_6_  ( .D(_padder__n1810 ), .CK(clk), .Q(
        padder_out[62]), .QN() );
  DFF_X1 _padder__out_reg_0_  ( .D(_padder__n2475 ), .CK(clk), .Q(
        padder_out[56]), .QN() );
  DFF_X1 _padder__out_reg_1_  ( .D(_padder__n1815 ), .CK(clk), .Q(
        padder_out[57]), .QN() );
  DFF_X1 _padder__out_reg_2_  ( .D(_padder__n1814 ), .CK(clk), .Q(
        padder_out[58]), .QN() );
  DFF_X1 _padder__out_reg_3_  ( .D(_padder__n1813 ), .CK(clk), .Q(
        padder_out[59]), .QN() );
  DFF_X1 _padder__state_reg  ( .D(_padder__n1836 ), .CK(clk), .Q(
        _padder__state ), .QN(_padder__n598 ) );
  DFF_X1 _padder__i_reg_17_  ( .D(_padder__n1817 ), .CK(clk), .Q(
        padder_out_ready), .QN(_padder__n1961 ) );
  NAND2_X2 _padder__U1820  ( .A1(padder_out[551]), .A2(_padder__n2484 ), .ZN(
        _padder__n2440 ) );
  NAND2_X2 _padder__U1818  ( .A1(padder_out[519]), .A2(_padder__n2511 ), .ZN(
        _padder__n2441 ) );
  NAND2_X2 _padder__U1817  ( .A1(_padder__n2440 ), .A2(_padder__n2441 ), .ZN(
        _padder__n1241 ) );
  NAND2_X2 _padder__U1816  ( .A1(padder_out[550]), .A2(_padder__n2500 ), .ZN(
        _padder__n2438 ) );
  NAND2_X2 _padder__U1815  ( .A1(padder_out[518]), .A2(_padder__n2511 ), .ZN(
        _padder__n2439 ) );
  NAND2_X2 _padder__U1814  ( .A1(_padder__n2438 ), .A2(_padder__n2439 ), .ZN(
        _padder__n1242 ) );
  NAND2_X2 _padder__U1813  ( .A1(padder_out[549]), .A2(_padder__n2500 ), .ZN(
        _padder__n2436 ) );
  NAND2_X2 _padder__U1812  ( .A1(padder_out[517]), .A2(_padder__n2511 ), .ZN(
        _padder__n2437 ) );
  NAND2_X2 _padder__U1811  ( .A1(_padder__n2436 ), .A2(_padder__n2437 ), .ZN(
        _padder__n1243 ) );
  NAND2_X2 _padder__U1810  ( .A1(padder_out[548]), .A2(_padder__n2500 ), .ZN(
        _padder__n2434 ) );
  NAND2_X2 _padder__U1809  ( .A1(padder_out[516]), .A2(_padder__n2511 ), .ZN(
        _padder__n2435 ) );
  NAND2_X2 _padder__U1808  ( .A1(_padder__n2434 ), .A2(_padder__n2435 ), .ZN(
        _padder__n1244 ) );
  NAND2_X2 _padder__U1807  ( .A1(padder_out[547]), .A2(_padder__n2500 ), .ZN(
        _padder__n2432 ) );
  NAND2_X2 _padder__U1806  ( .A1(padder_out[515]), .A2(_padder__n2511 ), .ZN(
        _padder__n2433 ) );
  NAND2_X2 _padder__U1805  ( .A1(_padder__n2432 ), .A2(_padder__n2433 ), .ZN(
        _padder__n1245 ) );
  NAND2_X2 _padder__U1804  ( .A1(padder_out[546]), .A2(_padder__n2500 ), .ZN(
        _padder__n2430 ) );
  NAND2_X2 _padder__U1803  ( .A1(padder_out[514]), .A2(_padder__n2511 ), .ZN(
        _padder__n2431 ) );
  NAND2_X2 _padder__U1802  ( .A1(_padder__n2430 ), .A2(_padder__n2431 ), .ZN(
        _padder__n1246 ) );
  NAND2_X2 _padder__U1801  ( .A1(padder_out[545]), .A2(_padder__n2499 ), .ZN(
        _padder__n2428 ) );
  NAND2_X2 _padder__U1800  ( .A1(padder_out[513]), .A2(_padder__n2511 ), .ZN(
        _padder__n2429 ) );
  NAND2_X2 _padder__U1799  ( .A1(_padder__n2428 ), .A2(_padder__n2429 ), .ZN(
        _padder__n1247 ) );
  NAND2_X2 _padder__U1798  ( .A1(padder_out[544]), .A2(_padder__n2499 ), .ZN(
        _padder__n2426 ) );
  NAND2_X2 _padder__U1797  ( .A1(padder_out[512]), .A2(_padder__n2511 ), .ZN(
        _padder__n2427 ) );
  NAND2_X2 _padder__U1796  ( .A1(_padder__n2426 ), .A2(_padder__n2427 ), .ZN(
        _padder__n1248 ) );
  NAND2_X2 _padder__U1795  ( .A1(padder_out[559]), .A2(_padder__n2499 ), .ZN(
        _padder__n2424 ) );
  NAND2_X2 _padder__U1794  ( .A1(padder_out[527]), .A2(_padder__n2511 ), .ZN(
        _padder__n2425 ) );
  NAND2_X2 _padder__U1793  ( .A1(_padder__n2424 ), .A2(_padder__n2425 ), .ZN(
        _padder__n1249 ) );
  NAND2_X2 _padder__U1792  ( .A1(padder_out[558]), .A2(_padder__n2499 ), .ZN(
        _padder__n2422 ) );
  NAND2_X2 _padder__U1791  ( .A1(padder_out[526]), .A2(_padder__n2511 ), .ZN(
        _padder__n2423 ) );
  NAND2_X2 _padder__U1790  ( .A1(_padder__n2422 ), .A2(_padder__n2423 ), .ZN(
        _padder__n1250 ) );
  NAND2_X2 _padder__U1789  ( .A1(padder_out[557]), .A2(_padder__n2499 ), .ZN(
        _padder__n2420 ) );
  NAND2_X2 _padder__U1788  ( .A1(padder_out[525]), .A2(_padder__n2511 ), .ZN(
        _padder__n2421 ) );
  NAND2_X2 _padder__U1787  ( .A1(_padder__n2420 ), .A2(_padder__n2421 ), .ZN(
        _padder__n1251 ) );
  NAND2_X2 _padder__U1786  ( .A1(padder_out[556]), .A2(_padder__n2499 ), .ZN(
        _padder__n2418 ) );
  NAND2_X2 _padder__U1785  ( .A1(padder_out[524]), .A2(_padder__n2512 ), .ZN(
        _padder__n2419 ) );
  NAND2_X2 _padder__U1784  ( .A1(_padder__n2418 ), .A2(_padder__n2419 ), .ZN(
        _padder__n1252 ) );
  NAND2_X2 _padder__U1783  ( .A1(padder_out[555]), .A2(_padder__n2499 ), .ZN(
        _padder__n2416 ) );
  NAND2_X2 _padder__U1782  ( .A1(padder_out[523]), .A2(_padder__n2512 ), .ZN(
        _padder__n2417 ) );
  NAND2_X2 _padder__U1781  ( .A1(_padder__n2416 ), .A2(_padder__n2417 ), .ZN(
        _padder__n1253 ) );
  NAND2_X2 _padder__U1780  ( .A1(padder_out[554]), .A2(_padder__n2499 ), .ZN(
        _padder__n2414 ) );
  NAND2_X2 _padder__U1779  ( .A1(padder_out[522]), .A2(_padder__n2512 ), .ZN(
        _padder__n2415 ) );
  NAND2_X2 _padder__U1778  ( .A1(_padder__n2414 ), .A2(_padder__n2415 ), .ZN(
        _padder__n1254 ) );
  NAND2_X2 _padder__U1777  ( .A1(padder_out[553]), .A2(_padder__n2499 ), .ZN(
        _padder__n2412 ) );
  NAND2_X2 _padder__U1776  ( .A1(padder_out[521]), .A2(_padder__n2512 ), .ZN(
        _padder__n2413 ) );
  NAND2_X2 _padder__U1775  ( .A1(_padder__n2412 ), .A2(_padder__n2413 ), .ZN(
        _padder__n1255 ) );
  NAND2_X2 _padder__U1774  ( .A1(padder_out[552]), .A2(_padder__n2499 ), .ZN(
        _padder__n2410 ) );
  NAND2_X2 _padder__U1773  ( .A1(padder_out[520]), .A2(_padder__n2512 ), .ZN(
        _padder__n2411 ) );
  NAND2_X2 _padder__U1772  ( .A1(_padder__n2410 ), .A2(_padder__n2411 ), .ZN(
        _padder__n1256 ) );
  NAND2_X2 _padder__U1771  ( .A1(padder_out[567]), .A2(_padder__n2499 ), .ZN(
        _padder__n2408 ) );
  NAND2_X2 _padder__U1770  ( .A1(padder_out[535]), .A2(_padder__n2512 ), .ZN(
        _padder__n2409 ) );
  NAND2_X2 _padder__U1769  ( .A1(_padder__n2408 ), .A2(_padder__n2409 ), .ZN(
        _padder__n1257 ) );
  NAND2_X2 _padder__U1768  ( .A1(padder_out[566]), .A2(_padder__n2499 ), .ZN(
        _padder__n2406 ) );
  NAND2_X2 _padder__U1767  ( .A1(padder_out[534]), .A2(_padder__n2512 ), .ZN(
        _padder__n2407 ) );
  NAND2_X2 _padder__U1766  ( .A1(_padder__n2406 ), .A2(_padder__n2407 ), .ZN(
        _padder__n1258 ) );
  NAND2_X2 _padder__U1765  ( .A1(padder_out[565]), .A2(_padder__n2499 ), .ZN(
        _padder__n2404 ) );
  NAND2_X2 _padder__U1764  ( .A1(padder_out[533]), .A2(_padder__n2512 ), .ZN(
        _padder__n2405 ) );
  NAND2_X2 _padder__U1763  ( .A1(_padder__n2404 ), .A2(_padder__n2405 ), .ZN(
        _padder__n1259 ) );
  NAND2_X2 _padder__U1762  ( .A1(padder_out[564]), .A2(_padder__n2499 ), .ZN(
        _padder__n2402 ) );
  NAND2_X2 _padder__U1761  ( .A1(padder_out[532]), .A2(_padder__n2512 ), .ZN(
        _padder__n2403 ) );
  NAND2_X2 _padder__U1760  ( .A1(_padder__n2402 ), .A2(_padder__n2403 ), .ZN(
        _padder__n1260 ) );
  NAND2_X2 _padder__U1759  ( .A1(padder_out[563]), .A2(_padder__n2499 ), .ZN(
        _padder__n2400 ) );
  NAND2_X2 _padder__U1758  ( .A1(padder_out[531]), .A2(_padder__n2512 ), .ZN(
        _padder__n2401 ) );
  NAND2_X2 _padder__U1757  ( .A1(_padder__n2400 ), .A2(_padder__n2401 ), .ZN(
        _padder__n1261 ) );
  NAND2_X2 _padder__U1756  ( .A1(padder_out[562]), .A2(_padder__n2499 ), .ZN(
        _padder__n2398 ) );
  NAND2_X2 _padder__U1755  ( .A1(padder_out[530]), .A2(_padder__n2512 ), .ZN(
        _padder__n2399 ) );
  NAND2_X2 _padder__U1754  ( .A1(_padder__n2398 ), .A2(_padder__n2399 ), .ZN(
        _padder__n1262 ) );
  NAND2_X2 _padder__U1753  ( .A1(padder_out[561]), .A2(_padder__n2499 ), .ZN(
        _padder__n2396 ) );
  NAND2_X2 _padder__U1752  ( .A1(padder_out[529]), .A2(_padder__n2513 ), .ZN(
        _padder__n2397 ) );
  NAND2_X2 _padder__U1751  ( .A1(_padder__n2396 ), .A2(_padder__n2397 ), .ZN(
        _padder__n1263 ) );
  NAND2_X2 _padder__U1750  ( .A1(padder_out[560]), .A2(_padder__n2499 ), .ZN(
        _padder__n2394 ) );
  NAND2_X2 _padder__U1749  ( .A1(padder_out[528]), .A2(_padder__n2513 ), .ZN(
        _padder__n2395 ) );
  NAND2_X2 _padder__U1748  ( .A1(_padder__n2394 ), .A2(_padder__n2395 ), .ZN(
        _padder__n1264 ) );
  NAND2_X2 _padder__U1747  ( .A1(padder_out[575]), .A2(_padder__n2499 ), .ZN(
        _padder__n2392 ) );
  NAND2_X2 _padder__U1746  ( .A1(padder_out[543]), .A2(_padder__n2513 ), .ZN(
        _padder__n2393 ) );
  NAND2_X2 _padder__U1745  ( .A1(_padder__n2392 ), .A2(_padder__n2393 ), .ZN(
        _padder__n1265 ) );
  NAND2_X2 _padder__U1744  ( .A1(padder_out[574]), .A2(_padder__n2499 ), .ZN(
        _padder__n2390 ) );
  NAND2_X2 _padder__U1743  ( .A1(padder_out[542]), .A2(_padder__n2513 ), .ZN(
        _padder__n2391 ) );
  NAND2_X2 _padder__U1742  ( .A1(_padder__n2390 ), .A2(_padder__n2391 ), .ZN(
        _padder__n1266 ) );
  NAND2_X2 _padder__U1741  ( .A1(padder_out[573]), .A2(_padder__n2499 ), .ZN(
        _padder__n2388 ) );
  NAND2_X2 _padder__U1740  ( .A1(padder_out[541]), .A2(_padder__n2513 ), .ZN(
        _padder__n2389 ) );
  NAND2_X2 _padder__U1739  ( .A1(_padder__n2388 ), .A2(_padder__n2389 ), .ZN(
        _padder__n1267 ) );
  NAND2_X2 _padder__U1738  ( .A1(padder_out[572]), .A2(_padder__n2499 ), .ZN(
        _padder__n2386 ) );
  NAND2_X2 _padder__U1737  ( .A1(padder_out[540]), .A2(_padder__n2513 ), .ZN(
        _padder__n2387 ) );
  NAND2_X2 _padder__U1736  ( .A1(_padder__n2386 ), .A2(_padder__n2387 ), .ZN(
        _padder__n1268 ) );
  NAND2_X2 _padder__U1735  ( .A1(padder_out[571]), .A2(_padder__n2499 ), .ZN(
        _padder__n2384 ) );
  NAND2_X2 _padder__U1734  ( .A1(padder_out[539]), .A2(_padder__n2513 ), .ZN(
        _padder__n2385 ) );
  NAND2_X2 _padder__U1733  ( .A1(_padder__n2384 ), .A2(_padder__n2385 ), .ZN(
        _padder__n1269 ) );
  NAND2_X2 _padder__U1732  ( .A1(padder_out[570]), .A2(_padder__n2499 ), .ZN(
        _padder__n2382 ) );
  NAND2_X2 _padder__U1731  ( .A1(padder_out[538]), .A2(_padder__n2513 ), .ZN(
        _padder__n2383 ) );
  NAND2_X2 _padder__U1730  ( .A1(_padder__n2382 ), .A2(_padder__n2383 ), .ZN(
        _padder__n1270 ) );
  NAND2_X2 _padder__U1729  ( .A1(padder_out[569]), .A2(_padder__n2498 ), .ZN(
        _padder__n2380 ) );
  NAND2_X2 _padder__U1728  ( .A1(padder_out[537]), .A2(_padder__n2513 ), .ZN(
        _padder__n2381 ) );
  NAND2_X2 _padder__U1727  ( .A1(_padder__n2380 ), .A2(_padder__n2381 ), .ZN(
        _padder__n1271 ) );
  NAND2_X2 _padder__U1726  ( .A1(padder_out[568]), .A2(_padder__n2498 ), .ZN(
        _padder__n2378 ) );
  NAND2_X2 _padder__U1725  ( .A1(padder_out[536]), .A2(_padder__n2513 ), .ZN(
        _padder__n2379 ) );
  NAND2_X2 _padder__U1724  ( .A1(_padder__n2378 ), .A2(_padder__n2379 ), .ZN(
        _padder__n1272 ) );
  NAND2_X2 _padder__U1723  ( .A1(padder_out[455]), .A2(_padder__n2498 ), .ZN(
        _padder__n2376 ) );
  NAND2_X2 _padder__U1722  ( .A1(padder_out[551]), .A2(_padder__n2513 ), .ZN(
        _padder__n2377 ) );
  NAND2_X2 _padder__U1721  ( .A1(_padder__n2376 ), .A2(_padder__n2377 ), .ZN(
        _padder__n1273 ) );
  NAND2_X2 _padder__U1720  ( .A1(padder_out[454]), .A2(_padder__n2498 ), .ZN(
        _padder__n2374 ) );
  NAND2_X2 _padder__U1719  ( .A1(padder_out[550]), .A2(_padder__n2514 ), .ZN(
        _padder__n2375 ) );
  NAND2_X2 _padder__U1718  ( .A1(_padder__n2374 ), .A2(_padder__n2375 ), .ZN(
        _padder__n1274 ) );
  NAND2_X2 _padder__U1717  ( .A1(padder_out[453]), .A2(_padder__n2498 ), .ZN(
        _padder__n2372 ) );
  NAND2_X2 _padder__U1716  ( .A1(padder_out[549]), .A2(_padder__n2514 ), .ZN(
        _padder__n2373 ) );
  NAND2_X2 _padder__U1715  ( .A1(_padder__n2372 ), .A2(_padder__n2373 ), .ZN(
        _padder__n1275 ) );
  NAND2_X2 _padder__U1714  ( .A1(padder_out[452]), .A2(_padder__n2498 ), .ZN(
        _padder__n2370 ) );
  NAND2_X2 _padder__U1713  ( .A1(padder_out[548]), .A2(_padder__n2514 ), .ZN(
        _padder__n2371 ) );
  NAND2_X2 _padder__U1712  ( .A1(_padder__n2370 ), .A2(_padder__n2371 ), .ZN(
        _padder__n1276 ) );
  NAND2_X2 _padder__U1711  ( .A1(padder_out[451]), .A2(_padder__n2498 ), .ZN(
        _padder__n2368 ) );
  NAND2_X2 _padder__U1710  ( .A1(padder_out[547]), .A2(_padder__n2514 ), .ZN(
        _padder__n2369 ) );
  NAND2_X2 _padder__U1709  ( .A1(_padder__n2368 ), .A2(_padder__n2369 ), .ZN(
        _padder__n1277 ) );
  NAND2_X2 _padder__U1708  ( .A1(padder_out[450]), .A2(_padder__n2498 ), .ZN(
        _padder__n2366 ) );
  NAND2_X2 _padder__U1707  ( .A1(padder_out[546]), .A2(_padder__n2514 ), .ZN(
        _padder__n2367 ) );
  NAND2_X2 _padder__U1706  ( .A1(_padder__n2366 ), .A2(_padder__n2367 ), .ZN(
        _padder__n1278 ) );
  NAND2_X2 _padder__U1705  ( .A1(padder_out[449]), .A2(_padder__n2498 ), .ZN(
        _padder__n2364 ) );
  NAND2_X2 _padder__U1704  ( .A1(padder_out[545]), .A2(_padder__n2514 ), .ZN(
        _padder__n2365 ) );
  NAND2_X2 _padder__U1703  ( .A1(_padder__n2364 ), .A2(_padder__n2365 ), .ZN(
        _padder__n1279 ) );
  NAND2_X2 _padder__U1702  ( .A1(padder_out[448]), .A2(_padder__n2498 ), .ZN(
        _padder__n2362 ) );
  NAND2_X2 _padder__U1701  ( .A1(padder_out[544]), .A2(_padder__n2514 ), .ZN(
        _padder__n2363 ) );
  NAND2_X2 _padder__U1700  ( .A1(_padder__n2362 ), .A2(_padder__n2363 ), .ZN(
        _padder__n1280 ) );
  NAND2_X2 _padder__U1699  ( .A1(padder_out[463]), .A2(_padder__n2498 ), .ZN(
        _padder__n2360 ) );
  NAND2_X2 _padder__U1698  ( .A1(padder_out[559]), .A2(_padder__n2514 ), .ZN(
        _padder__n2361 ) );
  NAND2_X2 _padder__U1697  ( .A1(_padder__n2360 ), .A2(_padder__n2361 ), .ZN(
        _padder__n1281 ) );
  NAND2_X2 _padder__U1696  ( .A1(padder_out[462]), .A2(_padder__n2498 ), .ZN(
        _padder__n2358 ) );
  NAND2_X2 _padder__U1695  ( .A1(padder_out[558]), .A2(_padder__n2514 ), .ZN(
        _padder__n2359 ) );
  NAND2_X2 _padder__U1694  ( .A1(_padder__n2358 ), .A2(_padder__n2359 ), .ZN(
        _padder__n1282 ) );
  NAND2_X2 _padder__U1693  ( .A1(padder_out[461]), .A2(_padder__n2498 ), .ZN(
        _padder__n2356 ) );
  NAND2_X2 _padder__U1692  ( .A1(padder_out[557]), .A2(_padder__n2514 ), .ZN(
        _padder__n2357 ) );
  NAND2_X2 _padder__U1691  ( .A1(_padder__n2356 ), .A2(_padder__n2357 ), .ZN(
        _padder__n1283 ) );
  NAND2_X2 _padder__U1690  ( .A1(padder_out[460]), .A2(_padder__n2498 ), .ZN(
        _padder__n2354 ) );
  NAND2_X2 _padder__U1689  ( .A1(padder_out[556]), .A2(_padder__n2514 ), .ZN(
        _padder__n2355 ) );
  NAND2_X2 _padder__U1688  ( .A1(_padder__n2354 ), .A2(_padder__n2355 ), .ZN(
        _padder__n1284 ) );
  NAND2_X2 _padder__U1687  ( .A1(padder_out[459]), .A2(_padder__n2498 ), .ZN(
        _padder__n2352 ) );
  NAND2_X2 _padder__U1686  ( .A1(padder_out[555]), .A2(_padder__n2515 ), .ZN(
        _padder__n2353 ) );
  NAND2_X2 _padder__U1685  ( .A1(_padder__n2352 ), .A2(_padder__n2353 ), .ZN(
        _padder__n1285 ) );
  NAND2_X2 _padder__U1684  ( .A1(padder_out[458]), .A2(_padder__n2498 ), .ZN(
        _padder__n2350 ) );
  NAND2_X2 _padder__U1683  ( .A1(padder_out[554]), .A2(_padder__n2515 ), .ZN(
        _padder__n2351 ) );
  NAND2_X2 _padder__U1682  ( .A1(_padder__n2350 ), .A2(_padder__n2351 ), .ZN(
        _padder__n1286 ) );
  NAND2_X2 _padder__U1681  ( .A1(padder_out[457]), .A2(_padder__n2498 ), .ZN(
        _padder__n2348 ) );
  NAND2_X2 _padder__U1680  ( .A1(padder_out[553]), .A2(_padder__n2515 ), .ZN(
        _padder__n2349 ) );
  NAND2_X2 _padder__U1679  ( .A1(_padder__n2348 ), .A2(_padder__n2349 ), .ZN(
        _padder__n1287 ) );
  NAND2_X2 _padder__U1678  ( .A1(padder_out[456]), .A2(_padder__n2498 ), .ZN(
        _padder__n2346 ) );
  NAND2_X2 _padder__U1677  ( .A1(padder_out[552]), .A2(_padder__n2515 ), .ZN(
        _padder__n2347 ) );
  NAND2_X2 _padder__U1676  ( .A1(_padder__n2346 ), .A2(_padder__n2347 ), .ZN(
        _padder__n1288 ) );
  NAND2_X2 _padder__U1675  ( .A1(padder_out[471]), .A2(_padder__n2498 ), .ZN(
        _padder__n2344 ) );
  NAND2_X2 _padder__U1674  ( .A1(padder_out[567]), .A2(_padder__n2515 ), .ZN(
        _padder__n2345 ) );
  NAND2_X2 _padder__U1673  ( .A1(_padder__n2344 ), .A2(_padder__n2345 ), .ZN(
        _padder__n1289 ) );
  NAND2_X2 _padder__U1672  ( .A1(padder_out[470]), .A2(_padder__n2498 ), .ZN(
        _padder__n2342 ) );
  NAND2_X2 _padder__U1671  ( .A1(padder_out[566]), .A2(_padder__n2515 ), .ZN(
        _padder__n2343 ) );
  NAND2_X2 _padder__U1670  ( .A1(_padder__n2342 ), .A2(_padder__n2343 ), .ZN(
        _padder__n1290 ) );
  NAND2_X2 _padder__U1669  ( .A1(padder_out[469]), .A2(_padder__n2498 ), .ZN(
        _padder__n2340 ) );
  NAND2_X2 _padder__U1668  ( .A1(padder_out[565]), .A2(_padder__n2515 ), .ZN(
        _padder__n2341 ) );
  NAND2_X2 _padder__U1667  ( .A1(_padder__n2340 ), .A2(_padder__n2341 ), .ZN(
        _padder__n1291 ) );
  NAND2_X2 _padder__U1666  ( .A1(padder_out[468]), .A2(_padder__n2498 ), .ZN(
        _padder__n2338 ) );
  NAND2_X2 _padder__U1665  ( .A1(padder_out[564]), .A2(_padder__n2515 ), .ZN(
        _padder__n2339 ) );
  NAND2_X2 _padder__U1664  ( .A1(_padder__n2338 ), .A2(_padder__n2339 ), .ZN(
        _padder__n1292 ) );
  NAND2_X2 _padder__U1663  ( .A1(padder_out[467]), .A2(_padder__n2498 ), .ZN(
        _padder__n2336 ) );
  NAND2_X2 _padder__U1662  ( .A1(padder_out[563]), .A2(_padder__n2515 ), .ZN(
        _padder__n2337 ) );
  NAND2_X2 _padder__U1661  ( .A1(_padder__n2336 ), .A2(_padder__n2337 ), .ZN(
        _padder__n1293 ) );
  NAND2_X2 _padder__U1660  ( .A1(padder_out[466]), .A2(_padder__n2498 ), .ZN(
        _padder__n2334 ) );
  NAND2_X2 _padder__U1659  ( .A1(padder_out[562]), .A2(_padder__n2515 ), .ZN(
        _padder__n2335 ) );
  NAND2_X2 _padder__U1658  ( .A1(_padder__n2334 ), .A2(_padder__n2335 ), .ZN(
        _padder__n1294 ) );
  NAND2_X2 _padder__U1657  ( .A1(padder_out[465]), .A2(_padder__n2497 ), .ZN(
        _padder__n2332 ) );
  NAND2_X2 _padder__U1656  ( .A1(padder_out[561]), .A2(_padder__n2515 ), .ZN(
        _padder__n2333 ) );
  NAND2_X2 _padder__U1655  ( .A1(_padder__n2332 ), .A2(_padder__n2333 ), .ZN(
        _padder__n1295 ) );
  NAND2_X2 _padder__U1654  ( .A1(padder_out[464]), .A2(_padder__n2497 ), .ZN(
        _padder__n2330 ) );
  NAND2_X2 _padder__U1653  ( .A1(padder_out[560]), .A2(_padder__n2516 ), .ZN(
        _padder__n2331 ) );
  NAND2_X2 _padder__U1652  ( .A1(_padder__n2330 ), .A2(_padder__n2331 ), .ZN(
        _padder__n1296 ) );
  NAND2_X2 _padder__U1651  ( .A1(padder_out[479]), .A2(_padder__n2497 ), .ZN(
        _padder__n2328 ) );
  NAND2_X2 _padder__U1650  ( .A1(padder_out[575]), .A2(_padder__n2516 ), .ZN(
        _padder__n2329 ) );
  NAND2_X2 _padder__U1649  ( .A1(_padder__n2328 ), .A2(_padder__n2329 ), .ZN(
        _padder__n1297 ) );
  NAND2_X2 _padder__U1648  ( .A1(padder_out[478]), .A2(_padder__n2497 ), .ZN(
        _padder__n2326 ) );
  NAND2_X2 _padder__U1647  ( .A1(padder_out[574]), .A2(_padder__n2516 ), .ZN(
        _padder__n2327 ) );
  NAND2_X2 _padder__U1646  ( .A1(_padder__n2326 ), .A2(_padder__n2327 ), .ZN(
        _padder__n1298 ) );
  NAND2_X2 _padder__U1645  ( .A1(padder_out[477]), .A2(_padder__n2497 ), .ZN(
        _padder__n2324 ) );
  NAND2_X2 _padder__U1644  ( .A1(padder_out[573]), .A2(_padder__n2516 ), .ZN(
        _padder__n2325 ) );
  NAND2_X2 _padder__U1643  ( .A1(_padder__n2324 ), .A2(_padder__n2325 ), .ZN(
        _padder__n1299 ) );
  NAND2_X2 _padder__U1642  ( .A1(padder_out[476]), .A2(_padder__n2497 ), .ZN(
        _padder__n2322 ) );
  NAND2_X2 _padder__U1641  ( .A1(padder_out[572]), .A2(_padder__n2516 ), .ZN(
        _padder__n2323 ) );
  NAND2_X2 _padder__U1640  ( .A1(_padder__n2322 ), .A2(_padder__n2323 ), .ZN(
        _padder__n1300 ) );
  NAND2_X2 _padder__U1639  ( .A1(padder_out[475]), .A2(_padder__n2497 ), .ZN(
        _padder__n2320 ) );
  NAND2_X2 _padder__U1638  ( .A1(padder_out[571]), .A2(_padder__n2516 ), .ZN(
        _padder__n2321 ) );
  NAND2_X2 _padder__U1637  ( .A1(_padder__n2320 ), .A2(_padder__n2321 ), .ZN(
        _padder__n1301 ) );
  NAND2_X2 _padder__U1636  ( .A1(padder_out[474]), .A2(_padder__n2497 ), .ZN(
        _padder__n2318 ) );
  NAND2_X2 _padder__U1635  ( .A1(padder_out[570]), .A2(_padder__n2516 ), .ZN(
        _padder__n2319 ) );
  NAND2_X2 _padder__U1634  ( .A1(_padder__n2318 ), .A2(_padder__n2319 ), .ZN(
        _padder__n1302 ) );
  NAND2_X2 _padder__U1633  ( .A1(padder_out[473]), .A2(_padder__n2497 ), .ZN(
        _padder__n2316 ) );
  NAND2_X2 _padder__U1632  ( .A1(padder_out[569]), .A2(_padder__n2516 ), .ZN(
        _padder__n2317 ) );
  NAND2_X2 _padder__U1631  ( .A1(_padder__n2316 ), .A2(_padder__n2317 ), .ZN(
        _padder__n1303 ) );
  NAND2_X2 _padder__U1630  ( .A1(padder_out[472]), .A2(_padder__n2497 ), .ZN(
        _padder__n2314 ) );
  NAND2_X2 _padder__U1629  ( .A1(padder_out[568]), .A2(_padder__n2516 ), .ZN(
        _padder__n2315 ) );
  NAND2_X2 _padder__U1628  ( .A1(_padder__n2314 ), .A2(_padder__n2315 ), .ZN(
        _padder__n1304 ) );
  NAND2_X2 _padder__U1627  ( .A1(padder_out[487]), .A2(_padder__n2497 ), .ZN(
        _padder__n2312 ) );
  NAND2_X2 _padder__U1626  ( .A1(padder_out[455]), .A2(_padder__n2516 ), .ZN(
        _padder__n2313 ) );
  NAND2_X2 _padder__U1625  ( .A1(_padder__n2312 ), .A2(_padder__n2313 ), .ZN(
        _padder__n1305 ) );
  NAND2_X2 _padder__U1624  ( .A1(padder_out[486]), .A2(_padder__n2497 ), .ZN(
        _padder__n2310 ) );
  NAND2_X2 _padder__U1623  ( .A1(padder_out[454]), .A2(_padder__n2516 ), .ZN(
        _padder__n2311 ) );
  NAND2_X2 _padder__U1622  ( .A1(_padder__n2310 ), .A2(_padder__n2311 ), .ZN(
        _padder__n1306 ) );
  NAND2_X2 _padder__U1621  ( .A1(padder_out[485]), .A2(_padder__n2497 ), .ZN(
        _padder__n2308 ) );
  NAND2_X2 _padder__U1620  ( .A1(padder_out[453]), .A2(_padder__n2517 ), .ZN(
        _padder__n2309 ) );
  NAND2_X2 _padder__U1619  ( .A1(_padder__n2308 ), .A2(_padder__n2309 ), .ZN(
        _padder__n1307 ) );
  NAND2_X2 _padder__U1618  ( .A1(padder_out[484]), .A2(_padder__n2497 ), .ZN(
        _padder__n2306 ) );
  NAND2_X2 _padder__U1617  ( .A1(padder_out[452]), .A2(_padder__n2517 ), .ZN(
        _padder__n2307 ) );
  NAND2_X2 _padder__U1616  ( .A1(_padder__n2306 ), .A2(_padder__n2307 ), .ZN(
        _padder__n1308 ) );
  NAND2_X2 _padder__U1615  ( .A1(padder_out[483]), .A2(_padder__n2497 ), .ZN(
        _padder__n2304 ) );
  NAND2_X2 _padder__U1614  ( .A1(padder_out[451]), .A2(_padder__n2517 ), .ZN(
        _padder__n2305 ) );
  NAND2_X2 _padder__U1613  ( .A1(_padder__n2304 ), .A2(_padder__n2305 ), .ZN(
        _padder__n1309 ) );
  NAND2_X2 _padder__U1612  ( .A1(padder_out[482]), .A2(_padder__n2497 ), .ZN(
        _padder__n2302 ) );
  NAND2_X2 _padder__U1611  ( .A1(padder_out[450]), .A2(_padder__n2517 ), .ZN(
        _padder__n2303 ) );
  NAND2_X2 _padder__U1610  ( .A1(_padder__n2302 ), .A2(_padder__n2303 ), .ZN(
        _padder__n1310 ) );
  NAND2_X2 _padder__U1609  ( .A1(padder_out[481]), .A2(_padder__n2497 ), .ZN(
        _padder__n2300 ) );
  NAND2_X2 _padder__U1608  ( .A1(padder_out[449]), .A2(_padder__n2517 ), .ZN(
        _padder__n2301 ) );
  NAND2_X2 _padder__U1607  ( .A1(_padder__n2300 ), .A2(_padder__n2301 ), .ZN(
        _padder__n1311 ) );
  NAND2_X2 _padder__U1606  ( .A1(padder_out[480]), .A2(_padder__n2497 ), .ZN(
        _padder__n2298 ) );
  NAND2_X2 _padder__U1605  ( .A1(padder_out[448]), .A2(_padder__n2517 ), .ZN(
        _padder__n2299 ) );
  NAND2_X2 _padder__U1604  ( .A1(_padder__n2298 ), .A2(_padder__n2299 ), .ZN(
        _padder__n1312 ) );
  NAND2_X2 _padder__U1603  ( .A1(padder_out[495]), .A2(_padder__n2497 ), .ZN(
        _padder__n2296 ) );
  NAND2_X2 _padder__U1602  ( .A1(padder_out[463]), .A2(_padder__n2517 ), .ZN(
        _padder__n2297 ) );
  NAND2_X2 _padder__U1601  ( .A1(_padder__n2296 ), .A2(_padder__n2297 ), .ZN(
        _padder__n1313 ) );
  NAND2_X2 _padder__U1600  ( .A1(padder_out[494]), .A2(_padder__n2497 ), .ZN(
        _padder__n2294 ) );
  NAND2_X2 _padder__U1599  ( .A1(padder_out[462]), .A2(_padder__n2517 ), .ZN(
        _padder__n2295 ) );
  NAND2_X2 _padder__U1598  ( .A1(_padder__n2294 ), .A2(_padder__n2295 ), .ZN(
        _padder__n1314 ) );
  NAND2_X2 _padder__U1597  ( .A1(padder_out[493]), .A2(_padder__n2497 ), .ZN(
        _padder__n2292 ) );
  NAND2_X2 _padder__U1596  ( .A1(padder_out[461]), .A2(_padder__n2517 ), .ZN(
        _padder__n2293 ) );
  NAND2_X2 _padder__U1595  ( .A1(_padder__n2292 ), .A2(_padder__n2293 ), .ZN(
        _padder__n1315 ) );
  NAND2_X2 _padder__U1594  ( .A1(padder_out[492]), .A2(_padder__n2497 ), .ZN(
        _padder__n2290 ) );
  NAND2_X2 _padder__U1593  ( .A1(padder_out[460]), .A2(_padder__n2517 ), .ZN(
        _padder__n2291 ) );
  NAND2_X2 _padder__U1592  ( .A1(_padder__n2290 ), .A2(_padder__n2291 ), .ZN(
        _padder__n1316 ) );
  NAND2_X2 _padder__U1591  ( .A1(padder_out[491]), .A2(_padder__n2497 ), .ZN(
        _padder__n2288 ) );
  NAND2_X2 _padder__U1590  ( .A1(padder_out[459]), .A2(_padder__n2517 ), .ZN(
        _padder__n2289 ) );
  NAND2_X2 _padder__U1589  ( .A1(_padder__n2288 ), .A2(_padder__n2289 ), .ZN(
        _padder__n1317 ) );
  NAND2_X2 _padder__U1588  ( .A1(padder_out[490]), .A2(_padder__n2496 ), .ZN(
        _padder__n2286 ) );
  NAND2_X2 _padder__U1587  ( .A1(padder_out[458]), .A2(_padder__n2518 ), .ZN(
        _padder__n2287 ) );
  NAND2_X2 _padder__U1586  ( .A1(_padder__n2286 ), .A2(_padder__n2287 ), .ZN(
        _padder__n1318 ) );
  NAND2_X2 _padder__U1585  ( .A1(padder_out[489]), .A2(_padder__n2496 ), .ZN(
        _padder__n2284 ) );
  NAND2_X2 _padder__U1584  ( .A1(padder_out[457]), .A2(_padder__n2518 ), .ZN(
        _padder__n2285 ) );
  NAND2_X2 _padder__U1583  ( .A1(_padder__n2284 ), .A2(_padder__n2285 ), .ZN(
        _padder__n1319 ) );
  NAND2_X2 _padder__U1582  ( .A1(padder_out[488]), .A2(_padder__n2496 ), .ZN(
        _padder__n2282 ) );
  NAND2_X2 _padder__U1581  ( .A1(padder_out[456]), .A2(_padder__n2518 ), .ZN(
        _padder__n2283 ) );
  NAND2_X2 _padder__U1580  ( .A1(_padder__n2282 ), .A2(_padder__n2283 ), .ZN(
        _padder__n1320 ) );
  NAND2_X2 _padder__U1579  ( .A1(padder_out[503]), .A2(_padder__n2496 ), .ZN(
        _padder__n2280 ) );
  NAND2_X2 _padder__U1578  ( .A1(padder_out[471]), .A2(_padder__n2518 ), .ZN(
        _padder__n2281 ) );
  NAND2_X2 _padder__U1577  ( .A1(_padder__n2280 ), .A2(_padder__n2281 ), .ZN(
        _padder__n1321 ) );
  NAND2_X2 _padder__U1576  ( .A1(padder_out[502]), .A2(_padder__n2496 ), .ZN(
        _padder__n2278 ) );
  NAND2_X2 _padder__U1575  ( .A1(padder_out[470]), .A2(_padder__n2518 ), .ZN(
        _padder__n2279 ) );
  NAND2_X2 _padder__U1574  ( .A1(_padder__n2278 ), .A2(_padder__n2279 ), .ZN(
        _padder__n1322 ) );
  NAND2_X2 _padder__U1573  ( .A1(padder_out[501]), .A2(_padder__n2496 ), .ZN(
        _padder__n2276 ) );
  NAND2_X2 _padder__U1572  ( .A1(padder_out[469]), .A2(_padder__n2518 ), .ZN(
        _padder__n2277 ) );
  NAND2_X2 _padder__U1571  ( .A1(_padder__n2276 ), .A2(_padder__n2277 ), .ZN(
        _padder__n1323 ) );
  NAND2_X2 _padder__U1570  ( .A1(padder_out[500]), .A2(_padder__n2496 ), .ZN(
        _padder__n2274 ) );
  NAND2_X2 _padder__U1569  ( .A1(padder_out[468]), .A2(_padder__n2518 ), .ZN(
        _padder__n2275 ) );
  NAND2_X2 _padder__U1568  ( .A1(_padder__n2274 ), .A2(_padder__n2275 ), .ZN(
        _padder__n1324 ) );
  NAND2_X2 _padder__U1567  ( .A1(padder_out[499]), .A2(_padder__n2496 ), .ZN(
        _padder__n2272 ) );
  NAND2_X2 _padder__U1566  ( .A1(padder_out[467]), .A2(_padder__n2518 ), .ZN(
        _padder__n2273 ) );
  NAND2_X2 _padder__U1565  ( .A1(_padder__n2272 ), .A2(_padder__n2273 ), .ZN(
        _padder__n1325 ) );
  NAND2_X2 _padder__U1564  ( .A1(padder_out[498]), .A2(_padder__n2496 ), .ZN(
        _padder__n2270 ) );
  NAND2_X2 _padder__U1563  ( .A1(padder_out[466]), .A2(_padder__n2518 ), .ZN(
        _padder__n2271 ) );
  NAND2_X2 _padder__U1562  ( .A1(_padder__n2270 ), .A2(_padder__n2271 ), .ZN(
        _padder__n1326 ) );
  NAND2_X2 _padder__U1561  ( .A1(padder_out[497]), .A2(_padder__n2496 ), .ZN(
        _padder__n2268 ) );
  NAND2_X2 _padder__U1560  ( .A1(padder_out[465]), .A2(_padder__n2518 ), .ZN(
        _padder__n2269 ) );
  NAND2_X2 _padder__U1559  ( .A1(_padder__n2268 ), .A2(_padder__n2269 ), .ZN(
        _padder__n1327 ) );
  NAND2_X2 _padder__U1558  ( .A1(padder_out[496]), .A2(_padder__n2496 ), .ZN(
        _padder__n2266 ) );
  NAND2_X2 _padder__U1557  ( .A1(padder_out[464]), .A2(_padder__n2518 ), .ZN(
        _padder__n2267 ) );
  NAND2_X2 _padder__U1556  ( .A1(_padder__n2266 ), .A2(_padder__n2267 ), .ZN(
        _padder__n1328 ) );
  NAND2_X2 _padder__U1555  ( .A1(padder_out[511]), .A2(_padder__n2496 ), .ZN(
        _padder__n2264 ) );
  NAND2_X2 _padder__U1554  ( .A1(padder_out[479]), .A2(_padder__n2519 ), .ZN(
        _padder__n2265 ) );
  NAND2_X2 _padder__U1553  ( .A1(_padder__n2264 ), .A2(_padder__n2265 ), .ZN(
        _padder__n1329 ) );
  NAND2_X2 _padder__U1552  ( .A1(padder_out[510]), .A2(_padder__n2496 ), .ZN(
        _padder__n2262 ) );
  NAND2_X2 _padder__U1551  ( .A1(padder_out[478]), .A2(_padder__n2519 ), .ZN(
        _padder__n2263 ) );
  NAND2_X2 _padder__U1550  ( .A1(_padder__n2262 ), .A2(_padder__n2263 ), .ZN(
        _padder__n1330 ) );
  NAND2_X2 _padder__U1549  ( .A1(padder_out[509]), .A2(_padder__n2496 ), .ZN(
        _padder__n2260 ) );
  NAND2_X2 _padder__U1548  ( .A1(padder_out[477]), .A2(_padder__n2519 ), .ZN(
        _padder__n2261 ) );
  NAND2_X2 _padder__U1547  ( .A1(_padder__n2260 ), .A2(_padder__n2261 ), .ZN(
        _padder__n1331 ) );
  NAND2_X2 _padder__U1546  ( .A1(padder_out[508]), .A2(_padder__n2496 ), .ZN(
        _padder__n2258 ) );
  NAND2_X2 _padder__U1545  ( .A1(padder_out[476]), .A2(_padder__n2519 ), .ZN(
        _padder__n2259 ) );
  NAND2_X2 _padder__U1544  ( .A1(_padder__n2258 ), .A2(_padder__n2259 ), .ZN(
        _padder__n1332 ) );
  NAND2_X2 _padder__U1543  ( .A1(padder_out[507]), .A2(_padder__n2496 ), .ZN(
        _padder__n2256 ) );
  NAND2_X2 _padder__U1542  ( .A1(padder_out[475]), .A2(_padder__n2519 ), .ZN(
        _padder__n2257 ) );
  NAND2_X2 _padder__U1541  ( .A1(_padder__n2256 ), .A2(_padder__n2257 ), .ZN(
        _padder__n1333 ) );
  NAND2_X2 _padder__U1540  ( .A1(padder_out[506]), .A2(_padder__n2496 ), .ZN(
        _padder__n2254 ) );
  NAND2_X2 _padder__U1539  ( .A1(padder_out[474]), .A2(_padder__n2519 ), .ZN(
        _padder__n2255 ) );
  NAND2_X2 _padder__U1538  ( .A1(_padder__n2254 ), .A2(_padder__n2255 ), .ZN(
        _padder__n1334 ) );
  NAND2_X2 _padder__U1537  ( .A1(padder_out[505]), .A2(_padder__n2496 ), .ZN(
        _padder__n2252 ) );
  NAND2_X2 _padder__U1536  ( .A1(padder_out[473]), .A2(_padder__n2519 ), .ZN(
        _padder__n2253 ) );
  NAND2_X2 _padder__U1535  ( .A1(_padder__n2252 ), .A2(_padder__n2253 ), .ZN(
        _padder__n1335 ) );
  NAND2_X2 _padder__U1534  ( .A1(padder_out[504]), .A2(_padder__n2496 ), .ZN(
        _padder__n2250 ) );
  NAND2_X2 _padder__U1533  ( .A1(padder_out[472]), .A2(_padder__n2519 ), .ZN(
        _padder__n2251 ) );
  NAND2_X2 _padder__U1532  ( .A1(_padder__n2250 ), .A2(_padder__n2251 ), .ZN(
        _padder__n1336 ) );
  NAND2_X2 _padder__U1531  ( .A1(padder_out[391]), .A2(_padder__n2496 ), .ZN(
        _padder__n2248 ) );
  NAND2_X2 _padder__U1530  ( .A1(padder_out[487]), .A2(_padder__n2519 ), .ZN(
        _padder__n2249 ) );
  NAND2_X2 _padder__U1529  ( .A1(_padder__n2248 ), .A2(_padder__n2249 ), .ZN(
        _padder__n1337 ) );
  NAND2_X2 _padder__U1528  ( .A1(padder_out[390]), .A2(_padder__n2496 ), .ZN(
        _padder__n2246 ) );
  NAND2_X2 _padder__U1527  ( .A1(padder_out[486]), .A2(_padder__n2519 ), .ZN(
        _padder__n2247 ) );
  NAND2_X2 _padder__U1526  ( .A1(_padder__n2246 ), .A2(_padder__n2247 ), .ZN(
        _padder__n1338 ) );
  NAND2_X2 _padder__U1525  ( .A1(padder_out[389]), .A2(_padder__n2496 ), .ZN(
        _padder__n2244 ) );
  NAND2_X2 _padder__U1524  ( .A1(padder_out[485]), .A2(_padder__n2519 ), .ZN(
        _padder__n2245 ) );
  NAND2_X2 _padder__U1523  ( .A1(_padder__n2244 ), .A2(_padder__n2245 ), .ZN(
        _padder__n1339 ) );
  NAND2_X2 _padder__U1522  ( .A1(padder_out[388]), .A2(_padder__n2496 ), .ZN(
        _padder__n2242 ) );
  NAND2_X2 _padder__U1521  ( .A1(padder_out[484]), .A2(_padder__n2520 ), .ZN(
        _padder__n2243 ) );
  NAND2_X2 _padder__U1520  ( .A1(_padder__n2242 ), .A2(_padder__n2243 ), .ZN(
        _padder__n1340 ) );
  NAND2_X2 _padder__U1519  ( .A1(padder_out[387]), .A2(_padder__n2496 ), .ZN(
        _padder__n2240 ) );
  NAND2_X2 _padder__U1518  ( .A1(padder_out[483]), .A2(_padder__n2520 ), .ZN(
        _padder__n2241 ) );
  NAND2_X2 _padder__U1517  ( .A1(_padder__n2240 ), .A2(_padder__n2241 ), .ZN(
        _padder__n1341 ) );
  NAND2_X2 _padder__U1516  ( .A1(padder_out[386]), .A2(_padder__n2495 ), .ZN(
        _padder__n2238 ) );
  NAND2_X2 _padder__U1515  ( .A1(padder_out[482]), .A2(_padder__n2520 ), .ZN(
        _padder__n2239 ) );
  NAND2_X2 _padder__U1514  ( .A1(_padder__n2238 ), .A2(_padder__n2239 ), .ZN(
        _padder__n1342 ) );
  NAND2_X2 _padder__U1513  ( .A1(padder_out[385]), .A2(_padder__n2495 ), .ZN(
        _padder__n2236 ) );
  NAND2_X2 _padder__U1512  ( .A1(padder_out[481]), .A2(_padder__n2520 ), .ZN(
        _padder__n2237 ) );
  NAND2_X2 _padder__U1511  ( .A1(_padder__n2236 ), .A2(_padder__n2237 ), .ZN(
        _padder__n1343 ) );
  NAND2_X2 _padder__U1510  ( .A1(padder_out[384]), .A2(_padder__n2495 ), .ZN(
        _padder__n2234 ) );
  NAND2_X2 _padder__U1509  ( .A1(padder_out[480]), .A2(_padder__n2520 ), .ZN(
        _padder__n2235 ) );
  NAND2_X2 _padder__U1508  ( .A1(_padder__n2234 ), .A2(_padder__n2235 ), .ZN(
        _padder__n1344 ) );
  NAND2_X2 _padder__U1507  ( .A1(padder_out[399]), .A2(_padder__n2495 ), .ZN(
        _padder__n2232 ) );
  NAND2_X2 _padder__U1506  ( .A1(padder_out[495]), .A2(_padder__n2520 ), .ZN(
        _padder__n2233 ) );
  NAND2_X2 _padder__U1505  ( .A1(_padder__n2232 ), .A2(_padder__n2233 ), .ZN(
        _padder__n1345 ) );
  NAND2_X2 _padder__U1504  ( .A1(padder_out[398]), .A2(_padder__n2495 ), .ZN(
        _padder__n2230 ) );
  NAND2_X2 _padder__U1503  ( .A1(padder_out[494]), .A2(_padder__n2520 ), .ZN(
        _padder__n2231 ) );
  NAND2_X2 _padder__U1502  ( .A1(_padder__n2230 ), .A2(_padder__n2231 ), .ZN(
        _padder__n1346 ) );
  NAND2_X2 _padder__U1501  ( .A1(padder_out[397]), .A2(_padder__n2495 ), .ZN(
        _padder__n2228 ) );
  NAND2_X2 _padder__U1500  ( .A1(padder_out[493]), .A2(_padder__n2520 ), .ZN(
        _padder__n2229 ) );
  NAND2_X2 _padder__U1499  ( .A1(_padder__n2228 ), .A2(_padder__n2229 ), .ZN(
        _padder__n1347 ) );
  NAND2_X2 _padder__U1498  ( .A1(padder_out[396]), .A2(_padder__n2495 ), .ZN(
        _padder__n2226 ) );
  NAND2_X2 _padder__U1497  ( .A1(padder_out[492]), .A2(_padder__n2520 ), .ZN(
        _padder__n2227 ) );
  NAND2_X2 _padder__U1496  ( .A1(_padder__n2226 ), .A2(_padder__n2227 ), .ZN(
        _padder__n1348 ) );
  NAND2_X2 _padder__U1495  ( .A1(padder_out[395]), .A2(_padder__n2495 ), .ZN(
        _padder__n2224 ) );
  NAND2_X2 _padder__U1494  ( .A1(padder_out[491]), .A2(_padder__n2520 ), .ZN(
        _padder__n2225 ) );
  NAND2_X2 _padder__U1493  ( .A1(_padder__n2224 ), .A2(_padder__n2225 ), .ZN(
        _padder__n1349 ) );
  NAND2_X2 _padder__U1492  ( .A1(padder_out[394]), .A2(_padder__n2495 ), .ZN(
        _padder__n2222 ) );
  NAND2_X2 _padder__U1491  ( .A1(padder_out[490]), .A2(_padder__n2520 ), .ZN(
        _padder__n2223 ) );
  NAND2_X2 _padder__U1490  ( .A1(_padder__n2222 ), .A2(_padder__n2223 ), .ZN(
        _padder__n1350 ) );
  NAND2_X2 _padder__U1489  ( .A1(padder_out[393]), .A2(_padder__n2495 ), .ZN(
        _padder__n2220 ) );
  NAND2_X2 _padder__U1488  ( .A1(padder_out[489]), .A2(_padder__n2521 ), .ZN(
        _padder__n2221 ) );
  NAND2_X2 _padder__U1487  ( .A1(_padder__n2220 ), .A2(_padder__n2221 ), .ZN(
        _padder__n1351 ) );
  NAND2_X2 _padder__U1486  ( .A1(padder_out[392]), .A2(_padder__n2495 ), .ZN(
        _padder__n2218 ) );
  NAND2_X2 _padder__U1485  ( .A1(padder_out[488]), .A2(_padder__n2521 ), .ZN(
        _padder__n2219 ) );
  NAND2_X2 _padder__U1484  ( .A1(_padder__n2218 ), .A2(_padder__n2219 ), .ZN(
        _padder__n1352 ) );
  NAND2_X2 _padder__U1483  ( .A1(padder_out[407]), .A2(_padder__n2495 ), .ZN(
        _padder__n2216 ) );
  NAND2_X2 _padder__U1482  ( .A1(padder_out[503]), .A2(_padder__n2521 ), .ZN(
        _padder__n2217 ) );
  NAND2_X2 _padder__U1481  ( .A1(_padder__n2216 ), .A2(_padder__n2217 ), .ZN(
        _padder__n1353 ) );
  NAND2_X2 _padder__U1480  ( .A1(padder_out[406]), .A2(_padder__n2495 ), .ZN(
        _padder__n2214 ) );
  NAND2_X2 _padder__U1479  ( .A1(padder_out[502]), .A2(_padder__n2521 ), .ZN(
        _padder__n2215 ) );
  NAND2_X2 _padder__U1478  ( .A1(_padder__n2214 ), .A2(_padder__n2215 ), .ZN(
        _padder__n1354 ) );
  NAND2_X2 _padder__U1477  ( .A1(padder_out[405]), .A2(_padder__n2495 ), .ZN(
        _padder__n2212 ) );
  NAND2_X2 _padder__U1476  ( .A1(padder_out[501]), .A2(_padder__n2521 ), .ZN(
        _padder__n2213 ) );
  NAND2_X2 _padder__U1475  ( .A1(_padder__n2212 ), .A2(_padder__n2213 ), .ZN(
        _padder__n1355 ) );
  NAND2_X2 _padder__U1474  ( .A1(padder_out[404]), .A2(_padder__n2495 ), .ZN(
        _padder__n2210 ) );
  NAND2_X2 _padder__U1473  ( .A1(padder_out[500]), .A2(_padder__n2521 ), .ZN(
        _padder__n2211 ) );
  NAND2_X2 _padder__U1472  ( .A1(_padder__n2210 ), .A2(_padder__n2211 ), .ZN(
        _padder__n1356 ) );
  NAND2_X2 _padder__U1471  ( .A1(padder_out[403]), .A2(_padder__n2495 ), .ZN(
        _padder__n2208 ) );
  NAND2_X2 _padder__U1470  ( .A1(padder_out[499]), .A2(_padder__n2521 ), .ZN(
        _padder__n2209 ) );
  NAND2_X2 _padder__U1469  ( .A1(_padder__n2208 ), .A2(_padder__n2209 ), .ZN(
        _padder__n1357 ) );
  NAND2_X2 _padder__U1468  ( .A1(padder_out[402]), .A2(_padder__n2495 ), .ZN(
        _padder__n2206 ) );
  NAND2_X2 _padder__U1467  ( .A1(padder_out[498]), .A2(_padder__n2521 ), .ZN(
        _padder__n2207 ) );
  NAND2_X2 _padder__U1466  ( .A1(_padder__n2206 ), .A2(_padder__n2207 ), .ZN(
        _padder__n1358 ) );
  NAND2_X2 _padder__U1465  ( .A1(padder_out[401]), .A2(_padder__n2495 ), .ZN(
        _padder__n2204 ) );
  NAND2_X2 _padder__U1464  ( .A1(padder_out[497]), .A2(_padder__n2521 ), .ZN(
        _padder__n2205 ) );
  NAND2_X2 _padder__U1463  ( .A1(_padder__n2204 ), .A2(_padder__n2205 ), .ZN(
        _padder__n1359 ) );
  NAND2_X2 _padder__U1462  ( .A1(padder_out[400]), .A2(_padder__n2495 ), .ZN(
        _padder__n2202 ) );
  NAND2_X2 _padder__U1461  ( .A1(padder_out[496]), .A2(_padder__n2521 ), .ZN(
        _padder__n2203 ) );
  NAND2_X2 _padder__U1460  ( .A1(_padder__n2202 ), .A2(_padder__n2203 ), .ZN(
        _padder__n1360 ) );
  NAND2_X2 _padder__U1459  ( .A1(padder_out[415]), .A2(_padder__n2495 ), .ZN(
        _padder__n2200 ) );
  NAND2_X2 _padder__U1458  ( .A1(padder_out[511]), .A2(_padder__n2521 ), .ZN(
        _padder__n2201 ) );
  NAND2_X2 _padder__U1457  ( .A1(_padder__n2200 ), .A2(_padder__n2201 ), .ZN(
        _padder__n1361 ) );
  NAND2_X2 _padder__U1456  ( .A1(padder_out[414]), .A2(_padder__n2495 ), .ZN(
        _padder__n2198 ) );
  NAND2_X2 _padder__U1455  ( .A1(padder_out[510]), .A2(_padder__n2522 ), .ZN(
        _padder__n2199 ) );
  NAND2_X2 _padder__U1454  ( .A1(_padder__n2198 ), .A2(_padder__n2199 ), .ZN(
        _padder__n1362 ) );
  NAND2_X2 _padder__U1453  ( .A1(padder_out[413]), .A2(_padder__n2495 ), .ZN(
        _padder__n2196 ) );
  NAND2_X2 _padder__U1452  ( .A1(padder_out[509]), .A2(_padder__n2522 ), .ZN(
        _padder__n2197 ) );
  NAND2_X2 _padder__U1451  ( .A1(_padder__n2196 ), .A2(_padder__n2197 ), .ZN(
        _padder__n1363 ) );
  NAND2_X2 _padder__U1450  ( .A1(padder_out[412]), .A2(_padder__n2495 ), .ZN(
        _padder__n2194 ) );
  NAND2_X2 _padder__U1449  ( .A1(padder_out[508]), .A2(_padder__n2522 ), .ZN(
        _padder__n2195 ) );
  NAND2_X2 _padder__U1448  ( .A1(_padder__n2194 ), .A2(_padder__n2195 ), .ZN(
        _padder__n1364 ) );
  NAND2_X2 _padder__U1447  ( .A1(padder_out[411]), .A2(_padder__n2495 ), .ZN(
        _padder__n2192 ) );
  NAND2_X2 _padder__U1446  ( .A1(padder_out[507]), .A2(_padder__n2522 ), .ZN(
        _padder__n2193 ) );
  NAND2_X2 _padder__U1445  ( .A1(_padder__n2192 ), .A2(_padder__n2193 ), .ZN(
        _padder__n1365 ) );
  NAND2_X2 _padder__U1444  ( .A1(padder_out[410]), .A2(_padder__n2494 ), .ZN(
        _padder__n2190 ) );
  NAND2_X2 _padder__U1443  ( .A1(padder_out[506]), .A2(_padder__n2522 ), .ZN(
        _padder__n2191 ) );
  NAND2_X2 _padder__U1442  ( .A1(_padder__n2190 ), .A2(_padder__n2191 ), .ZN(
        _padder__n1366 ) );
  NAND2_X2 _padder__U1441  ( .A1(padder_out[409]), .A2(_padder__n2494 ), .ZN(
        _padder__n2188 ) );
  NAND2_X2 _padder__U1440  ( .A1(padder_out[505]), .A2(_padder__n2522 ), .ZN(
        _padder__n2189 ) );
  NAND2_X2 _padder__U1439  ( .A1(_padder__n2188 ), .A2(_padder__n2189 ), .ZN(
        _padder__n1367 ) );
  NAND2_X2 _padder__U1438  ( .A1(padder_out[408]), .A2(_padder__n2494 ), .ZN(
        _padder__n2186 ) );
  NAND2_X2 _padder__U1437  ( .A1(padder_out[504]), .A2(_padder__n2522 ), .ZN(
        _padder__n2187 ) );
  NAND2_X2 _padder__U1436  ( .A1(_padder__n2186 ), .A2(_padder__n2187 ), .ZN(
        _padder__n1368 ) );
  NAND2_X2 _padder__U1435  ( .A1(padder_out[423]), .A2(_padder__n2494 ), .ZN(
        _padder__n2184 ) );
  NAND2_X2 _padder__U1434  ( .A1(padder_out[391]), .A2(_padder__n2522 ), .ZN(
        _padder__n2185 ) );
  NAND2_X2 _padder__U1433  ( .A1(_padder__n2184 ), .A2(_padder__n2185 ), .ZN(
        _padder__n1369 ) );
  NAND2_X2 _padder__U1432  ( .A1(padder_out[422]), .A2(_padder__n2494 ), .ZN(
        _padder__n2182 ) );
  NAND2_X2 _padder__U1431  ( .A1(padder_out[390]), .A2(_padder__n2522 ), .ZN(
        _padder__n2183 ) );
  NAND2_X2 _padder__U1430  ( .A1(_padder__n2182 ), .A2(_padder__n2183 ), .ZN(
        _padder__n1370 ) );
  NAND2_X2 _padder__U1429  ( .A1(padder_out[421]), .A2(_padder__n2494 ), .ZN(
        _padder__n2180 ) );
  NAND2_X2 _padder__U1428  ( .A1(padder_out[389]), .A2(_padder__n2522 ), .ZN(
        _padder__n2181 ) );
  NAND2_X2 _padder__U1427  ( .A1(_padder__n2180 ), .A2(_padder__n2181 ), .ZN(
        _padder__n1371 ) );
  NAND2_X2 _padder__U1426  ( .A1(padder_out[420]), .A2(_padder__n2494 ), .ZN(
        _padder__n2178 ) );
  NAND2_X2 _padder__U1425  ( .A1(padder_out[388]), .A2(_padder__n2522 ), .ZN(
        _padder__n2179 ) );
  NAND2_X2 _padder__U1424  ( .A1(_padder__n2178 ), .A2(_padder__n2179 ), .ZN(
        _padder__n1372 ) );
  NAND2_X2 _padder__U1423  ( .A1(padder_out[419]), .A2(_padder__n2494 ), .ZN(
        _padder__n2176 ) );
  NAND2_X2 _padder__U1422  ( .A1(padder_out[387]), .A2(_padder__n2523 ), .ZN(
        _padder__n2177 ) );
  NAND2_X2 _padder__U1421  ( .A1(_padder__n2176 ), .A2(_padder__n2177 ), .ZN(
        _padder__n1373 ) );
  NAND2_X2 _padder__U1420  ( .A1(padder_out[418]), .A2(_padder__n2494 ), .ZN(
        _padder__n2174 ) );
  NAND2_X2 _padder__U1419  ( .A1(padder_out[386]), .A2(_padder__n2523 ), .ZN(
        _padder__n2175 ) );
  NAND2_X2 _padder__U1418  ( .A1(_padder__n2174 ), .A2(_padder__n2175 ), .ZN(
        _padder__n1374 ) );
  NAND2_X2 _padder__U1417  ( .A1(padder_out[417]), .A2(_padder__n2494 ), .ZN(
        _padder__n2172 ) );
  NAND2_X2 _padder__U1416  ( .A1(padder_out[385]), .A2(_padder__n2523 ), .ZN(
        _padder__n2173 ) );
  NAND2_X2 _padder__U1415  ( .A1(_padder__n2172 ), .A2(_padder__n2173 ), .ZN(
        _padder__n1375 ) );
  NAND2_X2 _padder__U1414  ( .A1(padder_out[416]), .A2(_padder__n2494 ), .ZN(
        _padder__n2170 ) );
  NAND2_X2 _padder__U1413  ( .A1(padder_out[384]), .A2(_padder__n2523 ), .ZN(
        _padder__n2171 ) );
  NAND2_X2 _padder__U1412  ( .A1(_padder__n2170 ), .A2(_padder__n2171 ), .ZN(
        _padder__n1376 ) );
  NAND2_X2 _padder__U1411  ( .A1(padder_out[431]), .A2(_padder__n2497 ), .ZN(
        _padder__n2168 ) );
  NAND2_X2 _padder__U1410  ( .A1(padder_out[399]), .A2(_padder__n2523 ), .ZN(
        _padder__n2169 ) );
  NAND2_X2 _padder__U1409  ( .A1(_padder__n2168 ), .A2(_padder__n2169 ), .ZN(
        _padder__n1377 ) );
  NAND2_X2 _padder__U1408  ( .A1(padder_out[430]), .A2(_padder__n2505 ), .ZN(
        _padder__n2166 ) );
  NAND2_X2 _padder__U1407  ( .A1(padder_out[398]), .A2(_padder__n2523 ), .ZN(
        _padder__n2167 ) );
  NAND2_X2 _padder__U1406  ( .A1(_padder__n2166 ), .A2(_padder__n2167 ), .ZN(
        _padder__n1378 ) );
  NAND2_X2 _padder__U1405  ( .A1(padder_out[429]), .A2(_padder__n2505 ), .ZN(
        _padder__n2164 ) );
  NAND2_X2 _padder__U1404  ( .A1(padder_out[397]), .A2(_padder__n2523 ), .ZN(
        _padder__n2165 ) );
  NAND2_X2 _padder__U1403  ( .A1(_padder__n2164 ), .A2(_padder__n2165 ), .ZN(
        _padder__n1379 ) );
  NAND2_X2 _padder__U1402  ( .A1(padder_out[428]), .A2(_padder__n2505 ), .ZN(
        _padder__n2162 ) );
  NAND2_X2 _padder__U1401  ( .A1(padder_out[396]), .A2(_padder__n2523 ), .ZN(
        _padder__n2163 ) );
  NAND2_X2 _padder__U1400  ( .A1(_padder__n2162 ), .A2(_padder__n2163 ), .ZN(
        _padder__n1380 ) );
  NAND2_X2 _padder__U1399  ( .A1(padder_out[427]), .A2(_padder__n2505 ), .ZN(
        _padder__n2160 ) );
  NAND2_X2 _padder__U1398  ( .A1(padder_out[395]), .A2(_padder__n2523 ), .ZN(
        _padder__n2161 ) );
  NAND2_X2 _padder__U1397  ( .A1(_padder__n2160 ), .A2(_padder__n2161 ), .ZN(
        _padder__n1381 ) );
  NAND2_X2 _padder__U1396  ( .A1(padder_out[426]), .A2(_padder__n2505 ), .ZN(
        _padder__n2158 ) );
  NAND2_X2 _padder__U1395  ( .A1(padder_out[394]), .A2(_padder__n2523 ), .ZN(
        _padder__n2159 ) );
  NAND2_X2 _padder__U1394  ( .A1(_padder__n2158 ), .A2(_padder__n2159 ), .ZN(
        _padder__n1382 ) );
  NAND2_X2 _padder__U1393  ( .A1(padder_out[425]), .A2(_padder__n2505 ), .ZN(
        _padder__n2156 ) );
  NAND2_X2 _padder__U1392  ( .A1(padder_out[393]), .A2(_padder__n2523 ), .ZN(
        _padder__n2157 ) );
  NAND2_X2 _padder__U1391  ( .A1(_padder__n2156 ), .A2(_padder__n2157 ), .ZN(
        _padder__n1383 ) );
  NAND2_X2 _padder__U1390  ( .A1(padder_out[424]), .A2(_padder__n2505 ), .ZN(
        _padder__n2154 ) );
  NAND2_X2 _padder__U1389  ( .A1(padder_out[392]), .A2(_padder__n2524 ), .ZN(
        _padder__n2155 ) );
  NAND2_X2 _padder__U1388  ( .A1(_padder__n2154 ), .A2(_padder__n2155 ), .ZN(
        _padder__n1384 ) );
  NAND2_X2 _padder__U1387  ( .A1(padder_out[439]), .A2(_padder__n2505 ), .ZN(
        _padder__n2152 ) );
  NAND2_X2 _padder__U1386  ( .A1(padder_out[407]), .A2(_padder__n2524 ), .ZN(
        _padder__n2153 ) );
  NAND2_X2 _padder__U1385  ( .A1(_padder__n2152 ), .A2(_padder__n2153 ), .ZN(
        _padder__n1385 ) );
  NAND2_X2 _padder__U1384  ( .A1(padder_out[438]), .A2(_padder__n2505 ), .ZN(
        _padder__n2150 ) );
  NAND2_X2 _padder__U1383  ( .A1(padder_out[406]), .A2(_padder__n2524 ), .ZN(
        _padder__n2151 ) );
  NAND2_X2 _padder__U1382  ( .A1(_padder__n2150 ), .A2(_padder__n2151 ), .ZN(
        _padder__n1386 ) );
  NAND2_X2 _padder__U1381  ( .A1(padder_out[437]), .A2(_padder__n2505 ), .ZN(
        _padder__n2148 ) );
  NAND2_X2 _padder__U1380  ( .A1(padder_out[405]), .A2(_padder__n2524 ), .ZN(
        _padder__n2149 ) );
  NAND2_X2 _padder__U1379  ( .A1(_padder__n2148 ), .A2(_padder__n2149 ), .ZN(
        _padder__n1387 ) );
  NAND2_X2 _padder__U1378  ( .A1(padder_out[436]), .A2(_padder__n2505 ), .ZN(
        _padder__n2146 ) );
  NAND2_X2 _padder__U1377  ( .A1(padder_out[404]), .A2(_padder__n2524 ), .ZN(
        _padder__n2147 ) );
  NAND2_X2 _padder__U1376  ( .A1(_padder__n2146 ), .A2(_padder__n2147 ), .ZN(
        _padder__n1388 ) );
  NAND2_X2 _padder__U1375  ( .A1(padder_out[435]), .A2(_padder__n2505 ), .ZN(
        _padder__n2144 ) );
  NAND2_X2 _padder__U1374  ( .A1(padder_out[403]), .A2(_padder__n2524 ), .ZN(
        _padder__n2145 ) );
  NAND2_X2 _padder__U1373  ( .A1(_padder__n2144 ), .A2(_padder__n2145 ), .ZN(
        _padder__n1389 ) );
  NAND2_X2 _padder__U1372  ( .A1(padder_out[434]), .A2(_padder__n2505 ), .ZN(
        _padder__n2142 ) );
  NAND2_X2 _padder__U1371  ( .A1(padder_out[402]), .A2(_padder__n2524 ), .ZN(
        _padder__n2143 ) );
  NAND2_X2 _padder__U1370  ( .A1(_padder__n2142 ), .A2(_padder__n2143 ), .ZN(
        _padder__n1390 ) );
  NAND2_X2 _padder__U1369  ( .A1(padder_out[433]), .A2(_padder__n2505 ), .ZN(
        _padder__n2140 ) );
  NAND2_X2 _padder__U1368  ( .A1(padder_out[401]), .A2(_padder__n2524 ), .ZN(
        _padder__n2141 ) );
  NAND2_X2 _padder__U1367  ( .A1(_padder__n2140 ), .A2(_padder__n2141 ), .ZN(
        _padder__n1391 ) );
  NAND2_X2 _padder__U1366  ( .A1(padder_out[432]), .A2(_padder__n2505 ), .ZN(
        _padder__n2138 ) );
  NAND2_X2 _padder__U1365  ( .A1(padder_out[400]), .A2(_padder__n2524 ), .ZN(
        _padder__n2139 ) );
  NAND2_X2 _padder__U1364  ( .A1(_padder__n2138 ), .A2(_padder__n2139 ), .ZN(
        _padder__n1392 ) );
  NAND2_X2 _padder__U1363  ( .A1(padder_out[447]), .A2(_padder__n2505 ), .ZN(
        _padder__n2136 ) );
  NAND2_X2 _padder__U1362  ( .A1(padder_out[415]), .A2(_padder__n2524 ), .ZN(
        _padder__n2137 ) );
  NAND2_X2 _padder__U1361  ( .A1(_padder__n2136 ), .A2(_padder__n2137 ), .ZN(
        _padder__n1393 ) );
  NAND2_X2 _padder__U1360  ( .A1(padder_out[446]), .A2(_padder__n2505 ), .ZN(
        _padder__n2134 ) );
  NAND2_X2 _padder__U1359  ( .A1(padder_out[414]), .A2(_padder__n2524 ), .ZN(
        _padder__n2135 ) );
  NAND2_X2 _padder__U1358  ( .A1(_padder__n2134 ), .A2(_padder__n2135 ), .ZN(
        _padder__n1394 ) );
  NAND2_X2 _padder__U1357  ( .A1(padder_out[445]), .A2(_padder__n2505 ), .ZN(
        _padder__n2132 ) );
  NAND2_X2 _padder__U1356  ( .A1(padder_out[413]), .A2(_padder__n2525 ), .ZN(
        _padder__n2133 ) );
  NAND2_X2 _padder__U1355  ( .A1(_padder__n2132 ), .A2(_padder__n2133 ), .ZN(
        _padder__n1395 ) );
  NAND2_X2 _padder__U1354  ( .A1(padder_out[444]), .A2(_padder__n2505 ), .ZN(
        _padder__n2130 ) );
  NAND2_X2 _padder__U1353  ( .A1(padder_out[412]), .A2(_padder__n2525 ), .ZN(
        _padder__n2131 ) );
  NAND2_X2 _padder__U1352  ( .A1(_padder__n2130 ), .A2(_padder__n2131 ), .ZN(
        _padder__n1396 ) );
  NAND2_X2 _padder__U1351  ( .A1(padder_out[443]), .A2(_padder__n2505 ), .ZN(
        _padder__n2128 ) );
  NAND2_X2 _padder__U1350  ( .A1(padder_out[411]), .A2(_padder__n2525 ), .ZN(
        _padder__n2129 ) );
  NAND2_X2 _padder__U1349  ( .A1(_padder__n2128 ), .A2(_padder__n2129 ), .ZN(
        _padder__n1397 ) );
  NAND2_X2 _padder__U1348  ( .A1(padder_out[442]), .A2(_padder__n2505 ), .ZN(
        _padder__n2126 ) );
  NAND2_X2 _padder__U1347  ( .A1(padder_out[410]), .A2(_padder__n2525 ), .ZN(
        _padder__n2127 ) );
  NAND2_X2 _padder__U1346  ( .A1(_padder__n2126 ), .A2(_padder__n2127 ), .ZN(
        _padder__n1398 ) );
  NAND2_X2 _padder__U1345  ( .A1(padder_out[441]), .A2(_padder__n2504 ), .ZN(
        _padder__n2124 ) );
  NAND2_X2 _padder__U1344  ( .A1(padder_out[409]), .A2(_padder__n2525 ), .ZN(
        _padder__n2125 ) );
  NAND2_X2 _padder__U1343  ( .A1(_padder__n2124 ), .A2(_padder__n2125 ), .ZN(
        _padder__n1399 ) );
  NAND2_X2 _padder__U1342  ( .A1(padder_out[440]), .A2(_padder__n2504 ), .ZN(
        _padder__n2122 ) );
  NAND2_X2 _padder__U1341  ( .A1(padder_out[408]), .A2(_padder__n2525 ), .ZN(
        _padder__n2123 ) );
  NAND2_X2 _padder__U1340  ( .A1(_padder__n2122 ), .A2(_padder__n2123 ), .ZN(
        _padder__n1400 ) );
  NAND2_X2 _padder__U1339  ( .A1(padder_out[327]), .A2(_padder__n2504 ), .ZN(
        _padder__n2120 ) );
  NAND2_X2 _padder__U1338  ( .A1(padder_out[423]), .A2(_padder__n2525 ), .ZN(
        _padder__n2121 ) );
  NAND2_X2 _padder__U1337  ( .A1(_padder__n2120 ), .A2(_padder__n2121 ), .ZN(
        _padder__n1401 ) );
  NAND2_X2 _padder__U1336  ( .A1(padder_out[326]), .A2(_padder__n2504 ), .ZN(
        _padder__n2118 ) );
  NAND2_X2 _padder__U1335  ( .A1(padder_out[422]), .A2(_padder__n2525 ), .ZN(
        _padder__n2119 ) );
  NAND2_X2 _padder__U1334  ( .A1(_padder__n2118 ), .A2(_padder__n2119 ), .ZN(
        _padder__n1402 ) );
  NAND2_X2 _padder__U1333  ( .A1(padder_out[325]), .A2(_padder__n2504 ), .ZN(
        _padder__n2116 ) );
  NAND2_X2 _padder__U1332  ( .A1(padder_out[421]), .A2(_padder__n2525 ), .ZN(
        _padder__n2117 ) );
  NAND2_X2 _padder__U1331  ( .A1(_padder__n2116 ), .A2(_padder__n2117 ), .ZN(
        _padder__n1403 ) );
  NAND2_X2 _padder__U1330  ( .A1(padder_out[324]), .A2(_padder__n2504 ), .ZN(
        _padder__n2114 ) );
  NAND2_X2 _padder__U1329  ( .A1(padder_out[420]), .A2(_padder__n2525 ), .ZN(
        _padder__n2115 ) );
  NAND2_X2 _padder__U1328  ( .A1(_padder__n2114 ), .A2(_padder__n2115 ), .ZN(
        _padder__n1404 ) );
  NAND2_X2 _padder__U1327  ( .A1(padder_out[323]), .A2(_padder__n2504 ), .ZN(
        _padder__n2112 ) );
  NAND2_X2 _padder__U1326  ( .A1(padder_out[419]), .A2(_padder__n2525 ), .ZN(
        _padder__n2113 ) );
  NAND2_X2 _padder__U1325  ( .A1(_padder__n2112 ), .A2(_padder__n2113 ), .ZN(
        _padder__n1405 ) );
  NAND2_X2 _padder__U1324  ( .A1(padder_out[322]), .A2(_padder__n2504 ), .ZN(
        _padder__n2110 ) );
  NAND2_X2 _padder__U1323  ( .A1(padder_out[418]), .A2(_padder__n2526 ), .ZN(
        _padder__n2111 ) );
  NAND2_X2 _padder__U1322  ( .A1(_padder__n2110 ), .A2(_padder__n2111 ), .ZN(
        _padder__n1406 ) );
  NAND2_X2 _padder__U1321  ( .A1(padder_out[321]), .A2(_padder__n2504 ), .ZN(
        _padder__n2108 ) );
  NAND2_X2 _padder__U1320  ( .A1(padder_out[417]), .A2(_padder__n2526 ), .ZN(
        _padder__n2109 ) );
  NAND2_X2 _padder__U1319  ( .A1(_padder__n2108 ), .A2(_padder__n2109 ), .ZN(
        _padder__n1407 ) );
  NAND2_X2 _padder__U1318  ( .A1(padder_out[320]), .A2(_padder__n2504 ), .ZN(
        _padder__n2106 ) );
  NAND2_X2 _padder__U1317  ( .A1(padder_out[416]), .A2(_padder__n2526 ), .ZN(
        _padder__n2107 ) );
  NAND2_X2 _padder__U1316  ( .A1(_padder__n2106 ), .A2(_padder__n2107 ), .ZN(
        _padder__n1408 ) );
  NAND2_X2 _padder__U1315  ( .A1(padder_out[335]), .A2(_padder__n2504 ), .ZN(
        _padder__n2104 ) );
  NAND2_X2 _padder__U1314  ( .A1(padder_out[431]), .A2(_padder__n2526 ), .ZN(
        _padder__n2105 ) );
  NAND2_X2 _padder__U1313  ( .A1(_padder__n2104 ), .A2(_padder__n2105 ), .ZN(
        _padder__n1409 ) );
  NAND2_X2 _padder__U1312  ( .A1(padder_out[334]), .A2(_padder__n2504 ), .ZN(
        _padder__n2102 ) );
  NAND2_X2 _padder__U1311  ( .A1(padder_out[430]), .A2(_padder__n2526 ), .ZN(
        _padder__n2103 ) );
  NAND2_X2 _padder__U1310  ( .A1(_padder__n2102 ), .A2(_padder__n2103 ), .ZN(
        _padder__n1410 ) );
  NAND2_X2 _padder__U1309  ( .A1(padder_out[333]), .A2(_padder__n2504 ), .ZN(
        _padder__n2100 ) );
  NAND2_X2 _padder__U1308  ( .A1(padder_out[429]), .A2(_padder__n2526 ), .ZN(
        _padder__n2101 ) );
  NAND2_X2 _padder__U1307  ( .A1(_padder__n2100 ), .A2(_padder__n2101 ), .ZN(
        _padder__n1411 ) );
  NAND2_X2 _padder__U1306  ( .A1(padder_out[332]), .A2(_padder__n2504 ), .ZN(
        _padder__n2098 ) );
  NAND2_X2 _padder__U1305  ( .A1(padder_out[428]), .A2(_padder__n2526 ), .ZN(
        _padder__n2099 ) );
  NAND2_X2 _padder__U1304  ( .A1(_padder__n2098 ), .A2(_padder__n2099 ), .ZN(
        _padder__n1412 ) );
  NAND2_X2 _padder__U1303  ( .A1(padder_out[331]), .A2(_padder__n2504 ), .ZN(
        _padder__n2096 ) );
  NAND2_X2 _padder__U1302  ( .A1(padder_out[427]), .A2(_padder__n2526 ), .ZN(
        _padder__n2097 ) );
  NAND2_X2 _padder__U1301  ( .A1(_padder__n2096 ), .A2(_padder__n2097 ), .ZN(
        _padder__n1413 ) );
  NAND2_X2 _padder__U1300  ( .A1(padder_out[330]), .A2(_padder__n2504 ), .ZN(
        _padder__n2094 ) );
  NAND2_X2 _padder__U1299  ( .A1(padder_out[426]), .A2(_padder__n2526 ), .ZN(
        _padder__n2095 ) );
  NAND2_X2 _padder__U1298  ( .A1(_padder__n2094 ), .A2(_padder__n2095 ), .ZN(
        _padder__n1414 ) );
  NAND2_X2 _padder__U1297  ( .A1(padder_out[329]), .A2(_padder__n2504 ), .ZN(
        _padder__n2092 ) );
  NAND2_X2 _padder__U1296  ( .A1(padder_out[425]), .A2(_padder__n2526 ), .ZN(
        _padder__n2093 ) );
  NAND2_X2 _padder__U1295  ( .A1(_padder__n2092 ), .A2(_padder__n2093 ), .ZN(
        _padder__n1415 ) );
  NAND2_X2 _padder__U1294  ( .A1(padder_out[328]), .A2(_padder__n2504 ), .ZN(
        _padder__n2090 ) );
  NAND2_X2 _padder__U1293  ( .A1(padder_out[424]), .A2(_padder__n2526 ), .ZN(
        _padder__n2091 ) );
  NAND2_X2 _padder__U1292  ( .A1(_padder__n2090 ), .A2(_padder__n2091 ), .ZN(
        _padder__n1416 ) );
  NAND2_X2 _padder__U1291  ( .A1(padder_out[343]), .A2(_padder__n2504 ), .ZN(
        _padder__n2088 ) );
  NAND2_X2 _padder__U1290  ( .A1(padder_out[439]), .A2(_padder__n2527 ), .ZN(
        _padder__n2089 ) );
  NAND2_X2 _padder__U1289  ( .A1(_padder__n2088 ), .A2(_padder__n2089 ), .ZN(
        _padder__n1417 ) );
  NAND2_X2 _padder__U1288  ( .A1(padder_out[342]), .A2(_padder__n2504 ), .ZN(
        _padder__n2086 ) );
  NAND2_X2 _padder__U1287  ( .A1(padder_out[438]), .A2(_padder__n2527 ), .ZN(
        _padder__n2087 ) );
  NAND2_X2 _padder__U1286  ( .A1(_padder__n2086 ), .A2(_padder__n2087 ), .ZN(
        _padder__n1418 ) );
  NAND2_X2 _padder__U1285  ( .A1(padder_out[341]), .A2(_padder__n2504 ), .ZN(
        _padder__n2084 ) );
  NAND2_X2 _padder__U1284  ( .A1(padder_out[437]), .A2(_padder__n2527 ), .ZN(
        _padder__n2085 ) );
  NAND2_X2 _padder__U1283  ( .A1(_padder__n2084 ), .A2(_padder__n2085 ), .ZN(
        _padder__n1419 ) );
  NAND2_X2 _padder__U1282  ( .A1(padder_out[340]), .A2(_padder__n2504 ), .ZN(
        _padder__n2082 ) );
  NAND2_X2 _padder__U1281  ( .A1(padder_out[436]), .A2(_padder__n2527 ), .ZN(
        _padder__n2083 ) );
  NAND2_X2 _padder__U1280  ( .A1(_padder__n2082 ), .A2(_padder__n2083 ), .ZN(
        _padder__n1420 ) );
  NAND2_X2 _padder__U1279  ( .A1(padder_out[339]), .A2(_padder__n2504 ), .ZN(
        _padder__n2080 ) );
  NAND2_X2 _padder__U1278  ( .A1(padder_out[435]), .A2(_padder__n2527 ), .ZN(
        _padder__n2081 ) );
  NAND2_X2 _padder__U1277  ( .A1(_padder__n2080 ), .A2(_padder__n2081 ), .ZN(
        _padder__n1421 ) );
  NAND2_X2 _padder__U1276  ( .A1(padder_out[338]), .A2(_padder__n2504 ), .ZN(
        _padder__n2078 ) );
  NAND2_X2 _padder__U1275  ( .A1(padder_out[434]), .A2(_padder__n2527 ), .ZN(
        _padder__n2079 ) );
  NAND2_X2 _padder__U1274  ( .A1(_padder__n2078 ), .A2(_padder__n2079 ), .ZN(
        _padder__n1422 ) );
  NAND2_X2 _padder__U1273  ( .A1(padder_out[337]), .A2(_padder__n2503 ), .ZN(
        _padder__n2076 ) );
  NAND2_X2 _padder__U1272  ( .A1(padder_out[433]), .A2(_padder__n2527 ), .ZN(
        _padder__n2077 ) );
  NAND2_X2 _padder__U1271  ( .A1(_padder__n2076 ), .A2(_padder__n2077 ), .ZN(
        _padder__n1423 ) );
  NAND2_X2 _padder__U1270  ( .A1(padder_out[336]), .A2(_padder__n2503 ), .ZN(
        _padder__n2074 ) );
  NAND2_X2 _padder__U1269  ( .A1(padder_out[432]), .A2(_padder__n2527 ), .ZN(
        _padder__n2075 ) );
  NAND2_X2 _padder__U1268  ( .A1(_padder__n2074 ), .A2(_padder__n2075 ), .ZN(
        _padder__n1424 ) );
  NAND2_X2 _padder__U1267  ( .A1(padder_out[351]), .A2(_padder__n2503 ), .ZN(
        _padder__n2072 ) );
  NAND2_X2 _padder__U1266  ( .A1(padder_out[447]), .A2(_padder__n2527 ), .ZN(
        _padder__n2073 ) );
  NAND2_X2 _padder__U1265  ( .A1(_padder__n2072 ), .A2(_padder__n2073 ), .ZN(
        _padder__n1425 ) );
  NAND2_X2 _padder__U1264  ( .A1(padder_out[350]), .A2(_padder__n2503 ), .ZN(
        _padder__n2070 ) );
  NAND2_X2 _padder__U1263  ( .A1(padder_out[446]), .A2(_padder__n2527 ), .ZN(
        _padder__n2071 ) );
  NAND2_X2 _padder__U1262  ( .A1(_padder__n2070 ), .A2(_padder__n2071 ), .ZN(
        _padder__n1426 ) );
  NAND2_X2 _padder__U1261  ( .A1(padder_out[349]), .A2(_padder__n2503 ), .ZN(
        _padder__n2068 ) );
  NAND2_X2 _padder__U1260  ( .A1(padder_out[445]), .A2(_padder__n2527 ), .ZN(
        _padder__n2069 ) );
  NAND2_X2 _padder__U1259  ( .A1(_padder__n2068 ), .A2(_padder__n2069 ), .ZN(
        _padder__n1427 ) );
  NAND2_X2 _padder__U1258  ( .A1(padder_out[348]), .A2(_padder__n2503 ), .ZN(
        _padder__n2066 ) );
  NAND2_X2 _padder__U1257  ( .A1(padder_out[444]), .A2(_padder__n2528 ), .ZN(
        _padder__n2067 ) );
  NAND2_X2 _padder__U1256  ( .A1(_padder__n2066 ), .A2(_padder__n2067 ), .ZN(
        _padder__n1428 ) );
  NAND2_X2 _padder__U1255  ( .A1(padder_out[347]), .A2(_padder__n2503 ), .ZN(
        _padder__n2064 ) );
  NAND2_X2 _padder__U1254  ( .A1(padder_out[443]), .A2(_padder__n2528 ), .ZN(
        _padder__n2065 ) );
  NAND2_X2 _padder__U1253  ( .A1(_padder__n2064 ), .A2(_padder__n2065 ), .ZN(
        _padder__n1429 ) );
  NAND2_X2 _padder__U1252  ( .A1(padder_out[346]), .A2(_padder__n2503 ), .ZN(
        _padder__n2062 ) );
  NAND2_X2 _padder__U1251  ( .A1(padder_out[442]), .A2(_padder__n2528 ), .ZN(
        _padder__n2063 ) );
  NAND2_X2 _padder__U1250  ( .A1(_padder__n2062 ), .A2(_padder__n2063 ), .ZN(
        _padder__n1430 ) );
  NAND2_X2 _padder__U1249  ( .A1(padder_out[345]), .A2(_padder__n2503 ), .ZN(
        _padder__n2060 ) );
  NAND2_X2 _padder__U1248  ( .A1(padder_out[441]), .A2(_padder__n2528 ), .ZN(
        _padder__n2061 ) );
  NAND2_X2 _padder__U1247  ( .A1(_padder__n2060 ), .A2(_padder__n2061 ), .ZN(
        _padder__n1431 ) );
  NAND2_X2 _padder__U1246  ( .A1(padder_out[344]), .A2(_padder__n2503 ), .ZN(
        _padder__n2058 ) );
  NAND2_X2 _padder__U1245  ( .A1(padder_out[440]), .A2(_padder__n2528 ), .ZN(
        _padder__n2059 ) );
  NAND2_X2 _padder__U1244  ( .A1(_padder__n2058 ), .A2(_padder__n2059 ), .ZN(
        _padder__n1432 ) );
  NAND2_X2 _padder__U1243  ( .A1(padder_out[359]), .A2(_padder__n2503 ), .ZN(
        _padder__n2056 ) );
  NAND2_X2 _padder__U1242  ( .A1(padder_out[327]), .A2(_padder__n2528 ), .ZN(
        _padder__n2057 ) );
  NAND2_X2 _padder__U1241  ( .A1(_padder__n2056 ), .A2(_padder__n2057 ), .ZN(
        _padder__n1433 ) );
  NAND2_X2 _padder__U1240  ( .A1(padder_out[358]), .A2(_padder__n2503 ), .ZN(
        _padder__n2054 ) );
  NAND2_X2 _padder__U1239  ( .A1(padder_out[326]), .A2(_padder__n2528 ), .ZN(
        _padder__n2055 ) );
  NAND2_X2 _padder__U1238  ( .A1(_padder__n2054 ), .A2(_padder__n2055 ), .ZN(
        _padder__n1434 ) );
  NAND2_X2 _padder__U1237  ( .A1(padder_out[357]), .A2(_padder__n2503 ), .ZN(
        _padder__n2052 ) );
  NAND2_X2 _padder__U1236  ( .A1(padder_out[325]), .A2(_padder__n2528 ), .ZN(
        _padder__n2053 ) );
  NAND2_X2 _padder__U1235  ( .A1(_padder__n2052 ), .A2(_padder__n2053 ), .ZN(
        _padder__n1435 ) );
  NAND2_X2 _padder__U1234  ( .A1(padder_out[356]), .A2(_padder__n2503 ), .ZN(
        _padder__n2050 ) );
  NAND2_X2 _padder__U1233  ( .A1(padder_out[324]), .A2(_padder__n2528 ), .ZN(
        _padder__n2051 ) );
  NAND2_X2 _padder__U1232  ( .A1(_padder__n2050 ), .A2(_padder__n2051 ), .ZN(
        _padder__n1436 ) );
  NAND2_X2 _padder__U1231  ( .A1(padder_out[355]), .A2(_padder__n2503 ), .ZN(
        _padder__n2048 ) );
  NAND2_X2 _padder__U1230  ( .A1(padder_out[323]), .A2(_padder__n2528 ), .ZN(
        _padder__n2049 ) );
  NAND2_X2 _padder__U1229  ( .A1(_padder__n2048 ), .A2(_padder__n2049 ), .ZN(
        _padder__n1437 ) );
  NAND2_X2 _padder__U1228  ( .A1(padder_out[354]), .A2(_padder__n2503 ), .ZN(
        _padder__n2046 ) );
  NAND2_X2 _padder__U1227  ( .A1(padder_out[322]), .A2(_padder__n2528 ), .ZN(
        _padder__n2047 ) );
  NAND2_X2 _padder__U1226  ( .A1(_padder__n2046 ), .A2(_padder__n2047 ), .ZN(
        _padder__n1438 ) );
  NAND2_X2 _padder__U1225  ( .A1(padder_out[353]), .A2(_padder__n2503 ), .ZN(
        _padder__n2044 ) );
  NAND2_X2 _padder__U1224  ( .A1(padder_out[321]), .A2(_padder__n2529 ), .ZN(
        _padder__n2045 ) );
  NAND2_X2 _padder__U1223  ( .A1(_padder__n2044 ), .A2(_padder__n2045 ), .ZN(
        _padder__n1439 ) );
  NAND2_X2 _padder__U1222  ( .A1(padder_out[352]), .A2(_padder__n2503 ), .ZN(
        _padder__n2042 ) );
  NAND2_X2 _padder__U1221  ( .A1(padder_out[320]), .A2(_padder__n2529 ), .ZN(
        _padder__n2043 ) );
  NAND2_X2 _padder__U1220  ( .A1(_padder__n2042 ), .A2(_padder__n2043 ), .ZN(
        _padder__n1440 ) );
  NAND2_X2 _padder__U1219  ( .A1(padder_out[367]), .A2(_padder__n2503 ), .ZN(
        _padder__n2040 ) );
  NAND2_X2 _padder__U1218  ( .A1(padder_out[335]), .A2(_padder__n2529 ), .ZN(
        _padder__n2041 ) );
  NAND2_X2 _padder__U1217  ( .A1(_padder__n2040 ), .A2(_padder__n2041 ), .ZN(
        _padder__n1441 ) );
  NAND2_X2 _padder__U1216  ( .A1(padder_out[366]), .A2(_padder__n2503 ), .ZN(
        _padder__n2038 ) );
  NAND2_X2 _padder__U1215  ( .A1(padder_out[334]), .A2(_padder__n2529 ), .ZN(
        _padder__n2039 ) );
  NAND2_X2 _padder__U1214  ( .A1(_padder__n2038 ), .A2(_padder__n2039 ), .ZN(
        _padder__n1442 ) );
  NAND2_X2 _padder__U1213  ( .A1(padder_out[365]), .A2(_padder__n2503 ), .ZN(
        _padder__n2036 ) );
  NAND2_X2 _padder__U1212  ( .A1(padder_out[333]), .A2(_padder__n2529 ), .ZN(
        _padder__n2037 ) );
  NAND2_X2 _padder__U1211  ( .A1(_padder__n2036 ), .A2(_padder__n2037 ), .ZN(
        _padder__n1443 ) );
  NAND2_X2 _padder__U1210  ( .A1(padder_out[364]), .A2(_padder__n2503 ), .ZN(
        _padder__n2034 ) );
  NAND2_X2 _padder__U1209  ( .A1(padder_out[332]), .A2(_padder__n2529 ), .ZN(
        _padder__n2035 ) );
  NAND2_X2 _padder__U1208  ( .A1(_padder__n2034 ), .A2(_padder__n2035 ), .ZN(
        _padder__n1444 ) );
  NAND2_X2 _padder__U1207  ( .A1(padder_out[363]), .A2(_padder__n2503 ), .ZN(
        _padder__n2032 ) );
  NAND2_X2 _padder__U1206  ( .A1(padder_out[331]), .A2(_padder__n2529 ), .ZN(
        _padder__n2033 ) );
  NAND2_X2 _padder__U1205  ( .A1(_padder__n2032 ), .A2(_padder__n2033 ), .ZN(
        _padder__n1445 ) );
  NAND2_X2 _padder__U1204  ( .A1(padder_out[362]), .A2(_padder__n2502 ), .ZN(
        _padder__n2030 ) );
  NAND2_X2 _padder__U1203  ( .A1(padder_out[330]), .A2(_padder__n2529 ), .ZN(
        _padder__n2031 ) );
  NAND2_X2 _padder__U1202  ( .A1(_padder__n2030 ), .A2(_padder__n2031 ), .ZN(
        _padder__n1446 ) );
  NAND2_X2 _padder__U1201  ( .A1(padder_out[361]), .A2(_padder__n2502 ), .ZN(
        _padder__n2028 ) );
  NAND2_X2 _padder__U1200  ( .A1(padder_out[329]), .A2(_padder__n2529 ), .ZN(
        _padder__n2029 ) );
  NAND2_X2 _padder__U1199  ( .A1(_padder__n2028 ), .A2(_padder__n2029 ), .ZN(
        _padder__n1447 ) );
  NAND2_X2 _padder__U1198  ( .A1(padder_out[360]), .A2(_padder__n2502 ), .ZN(
        _padder__n2026 ) );
  NAND2_X2 _padder__U1197  ( .A1(padder_out[328]), .A2(_padder__n2529 ), .ZN(
        _padder__n2027 ) );
  NAND2_X2 _padder__U1196  ( .A1(_padder__n2026 ), .A2(_padder__n2027 ), .ZN(
        _padder__n1448 ) );
  NAND2_X2 _padder__U1195  ( .A1(padder_out[375]), .A2(_padder__n2502 ), .ZN(
        _padder__n2024 ) );
  NAND2_X2 _padder__U1194  ( .A1(padder_out[343]), .A2(_padder__n2529 ), .ZN(
        _padder__n2025 ) );
  NAND2_X2 _padder__U1193  ( .A1(_padder__n2024 ), .A2(_padder__n2025 ), .ZN(
        _padder__n1449 ) );
  NAND2_X2 _padder__U1192  ( .A1(padder_out[374]), .A2(_padder__n2502 ), .ZN(
        _padder__n2022 ) );
  NAND2_X2 _padder__U1191  ( .A1(padder_out[342]), .A2(_padder__n2530 ), .ZN(
        _padder__n2023 ) );
  NAND2_X2 _padder__U1190  ( .A1(_padder__n2022 ), .A2(_padder__n2023 ), .ZN(
        _padder__n1450 ) );
  NAND2_X2 _padder__U1189  ( .A1(padder_out[373]), .A2(_padder__n2502 ), .ZN(
        _padder__n2020 ) );
  NAND2_X2 _padder__U1188  ( .A1(padder_out[341]), .A2(_padder__n2530 ), .ZN(
        _padder__n2021 ) );
  NAND2_X2 _padder__U1187  ( .A1(_padder__n2020 ), .A2(_padder__n2021 ), .ZN(
        _padder__n1451 ) );
  NAND2_X2 _padder__U1186  ( .A1(padder_out[372]), .A2(_padder__n2502 ), .ZN(
        _padder__n2018 ) );
  NAND2_X2 _padder__U1185  ( .A1(padder_out[340]), .A2(_padder__n2530 ), .ZN(
        _padder__n2019 ) );
  NAND2_X2 _padder__U1184  ( .A1(_padder__n2018 ), .A2(_padder__n2019 ), .ZN(
        _padder__n1452 ) );
  NAND2_X2 _padder__U1183  ( .A1(padder_out[371]), .A2(_padder__n2502 ), .ZN(
        _padder__n2016 ) );
  NAND2_X2 _padder__U1182  ( .A1(padder_out[339]), .A2(_padder__n2530 ), .ZN(
        _padder__n2017 ) );
  NAND2_X2 _padder__U1181  ( .A1(_padder__n2016 ), .A2(_padder__n2017 ), .ZN(
        _padder__n1453 ) );
  NAND2_X2 _padder__U1180  ( .A1(padder_out[370]), .A2(_padder__n2502 ), .ZN(
        _padder__n2014 ) );
  NAND2_X2 _padder__U1179  ( .A1(padder_out[338]), .A2(_padder__n2530 ), .ZN(
        _padder__n2015 ) );
  NAND2_X2 _padder__U1178  ( .A1(_padder__n2014 ), .A2(_padder__n2015 ), .ZN(
        _padder__n1454 ) );
  NAND2_X2 _padder__U1177  ( .A1(padder_out[369]), .A2(_padder__n2502 ), .ZN(
        _padder__n2012 ) );
  NAND2_X2 _padder__U1176  ( .A1(padder_out[337]), .A2(_padder__n2530 ), .ZN(
        _padder__n2013 ) );
  NAND2_X2 _padder__U1175  ( .A1(_padder__n2012 ), .A2(_padder__n2013 ), .ZN(
        _padder__n1455 ) );
  NAND2_X2 _padder__U1174  ( .A1(padder_out[368]), .A2(_padder__n2502 ), .ZN(
        _padder__n2010 ) );
  NAND2_X2 _padder__U1173  ( .A1(padder_out[336]), .A2(_padder__n2530 ), .ZN(
        _padder__n2011 ) );
  NAND2_X2 _padder__U1172  ( .A1(_padder__n2010 ), .A2(_padder__n2011 ), .ZN(
        _padder__n1456 ) );
  NAND2_X2 _padder__U1171  ( .A1(padder_out[383]), .A2(_padder__n2502 ), .ZN(
        _padder__n2008 ) );
  NAND2_X2 _padder__U1170  ( .A1(padder_out[351]), .A2(_padder__n2530 ), .ZN(
        _padder__n2009 ) );
  NAND2_X2 _padder__U1169  ( .A1(_padder__n2008 ), .A2(_padder__n2009 ), .ZN(
        _padder__n1457 ) );
  NAND2_X2 _padder__U1168  ( .A1(padder_out[382]), .A2(_padder__n2502 ), .ZN(
        _padder__n2006 ) );
  NAND2_X2 _padder__U1167  ( .A1(padder_out[350]), .A2(_padder__n2530 ), .ZN(
        _padder__n2007 ) );
  NAND2_X2 _padder__U1166  ( .A1(_padder__n2006 ), .A2(_padder__n2007 ), .ZN(
        _padder__n1458 ) );
  NAND2_X2 _padder__U1165  ( .A1(padder_out[381]), .A2(_padder__n2502 ), .ZN(
        _padder__n2004 ) );
  NAND2_X2 _padder__U1164  ( .A1(padder_out[349]), .A2(_padder__n2530 ), .ZN(
        _padder__n2005 ) );
  NAND2_X2 _padder__U1163  ( .A1(_padder__n2004 ), .A2(_padder__n2005 ), .ZN(
        _padder__n1459 ) );
  NAND2_X2 _padder__U1162  ( .A1(padder_out[380]), .A2(_padder__n2502 ), .ZN(
        _padder__n2002 ) );
  NAND2_X2 _padder__U1161  ( .A1(padder_out[348]), .A2(_padder__n2530 ), .ZN(
        _padder__n2003 ) );
  NAND2_X2 _padder__U1160  ( .A1(_padder__n2002 ), .A2(_padder__n2003 ), .ZN(
        _padder__n1460 ) );
  NAND2_X2 _padder__U1159  ( .A1(padder_out[379]), .A2(_padder__n2502 ), .ZN(
        _padder__n2000 ) );
  NAND2_X2 _padder__U1158  ( .A1(padder_out[347]), .A2(_padder__n2531 ), .ZN(
        _padder__n2001 ) );
  NAND2_X2 _padder__U1157  ( .A1(_padder__n2000 ), .A2(_padder__n2001 ), .ZN(
        _padder__n1461 ) );
  NAND2_X2 _padder__U1156  ( .A1(padder_out[378]), .A2(_padder__n2502 ), .ZN(
        _padder__n1998 ) );
  NAND2_X2 _padder__U1155  ( .A1(padder_out[346]), .A2(_padder__n2531 ), .ZN(
        _padder__n1999 ) );
  NAND2_X2 _padder__U1154  ( .A1(_padder__n1998 ), .A2(_padder__n1999 ), .ZN(
        _padder__n1462 ) );
  NAND2_X2 _padder__U1153  ( .A1(padder_out[377]), .A2(_padder__n2502 ), .ZN(
        _padder__n1996 ) );
  NAND2_X2 _padder__U1152  ( .A1(padder_out[345]), .A2(_padder__n2531 ), .ZN(
        _padder__n1997 ) );
  NAND2_X2 _padder__U1151  ( .A1(_padder__n1996 ), .A2(_padder__n1997 ), .ZN(
        _padder__n1463 ) );
  NAND2_X2 _padder__U1150  ( .A1(padder_out[376]), .A2(_padder__n2502 ), .ZN(
        _padder__n1994 ) );
  NAND2_X2 _padder__U1149  ( .A1(padder_out[344]), .A2(_padder__n2531 ), .ZN(
        _padder__n1995 ) );
  NAND2_X2 _padder__U1148  ( .A1(_padder__n1994 ), .A2(_padder__n1995 ), .ZN(
        _padder__n1464 ) );
  NAND2_X2 _padder__U1147  ( .A1(padder_out[263]), .A2(_padder__n2502 ), .ZN(
        _padder__n1992 ) );
  NAND2_X2 _padder__U1146  ( .A1(padder_out[359]), .A2(_padder__n2531 ), .ZN(
        _padder__n1993 ) );
  NAND2_X2 _padder__U1145  ( .A1(_padder__n1992 ), .A2(_padder__n1993 ), .ZN(
        _padder__n1465 ) );
  NAND2_X2 _padder__U1144  ( .A1(padder_out[262]), .A2(_padder__n2502 ), .ZN(
        _padder__n1990 ) );
  NAND2_X2 _padder__U1143  ( .A1(padder_out[358]), .A2(_padder__n2531 ), .ZN(
        _padder__n1991 ) );
  NAND2_X2 _padder__U1142  ( .A1(_padder__n1990 ), .A2(_padder__n1991 ), .ZN(
        _padder__n1466 ) );
  NAND2_X2 _padder__U1141  ( .A1(padder_out[261]), .A2(_padder__n2502 ), .ZN(
        _padder__n1988 ) );
  NAND2_X2 _padder__U1140  ( .A1(padder_out[357]), .A2(_padder__n2531 ), .ZN(
        _padder__n1989 ) );
  NAND2_X2 _padder__U1139  ( .A1(_padder__n1988 ), .A2(_padder__n1989 ), .ZN(
        _padder__n1467 ) );
  NAND2_X2 _padder__U1138  ( .A1(padder_out[260]), .A2(_padder__n2502 ), .ZN(
        _padder__n1986 ) );
  NAND2_X2 _padder__U1137  ( .A1(padder_out[356]), .A2(_padder__n2531 ), .ZN(
        _padder__n1987 ) );
  NAND2_X2 _padder__U1136  ( .A1(_padder__n1986 ), .A2(_padder__n1987 ), .ZN(
        _padder__n1468 ) );
  NAND2_X2 _padder__U1135  ( .A1(padder_out[259]), .A2(_padder__n2502 ), .ZN(
        _padder__n1984 ) );
  NAND2_X2 _padder__U1134  ( .A1(padder_out[355]), .A2(_padder__n2531 ), .ZN(
        _padder__n1985 ) );
  NAND2_X2 _padder__U1133  ( .A1(_padder__n1984 ), .A2(_padder__n1985 ), .ZN(
        _padder__n1469 ) );
  NAND2_X2 _padder__U1132  ( .A1(padder_out[258]), .A2(_padder__n2501 ), .ZN(
        _padder__n1982 ) );
  NAND2_X2 _padder__U1131  ( .A1(padder_out[354]), .A2(_padder__n2531 ), .ZN(
        _padder__n1983 ) );
  NAND2_X2 _padder__U1130  ( .A1(_padder__n1982 ), .A2(_padder__n1983 ), .ZN(
        _padder__n1470 ) );
  NAND2_X2 _padder__U1129  ( .A1(padder_out[257]), .A2(_padder__n2501 ), .ZN(
        _padder__n1980 ) );
  NAND2_X2 _padder__U1128  ( .A1(padder_out[353]), .A2(_padder__n2531 ), .ZN(
        _padder__n1981 ) );
  NAND2_X2 _padder__U1127  ( .A1(_padder__n1980 ), .A2(_padder__n1981 ), .ZN(
        _padder__n1471 ) );
  NAND2_X2 _padder__U1126  ( .A1(padder_out[256]), .A2(_padder__n2501 ), .ZN(
        _padder__n1978 ) );
  NAND2_X2 _padder__U1125  ( .A1(padder_out[352]), .A2(_padder__n2532 ), .ZN(
        _padder__n1979 ) );
  NAND2_X2 _padder__U1124  ( .A1(_padder__n1978 ), .A2(_padder__n1979 ), .ZN(
        _padder__n1472 ) );
  NAND2_X2 _padder__U1123  ( .A1(padder_out[271]), .A2(_padder__n2501 ), .ZN(
        _padder__n1976 ) );
  NAND2_X2 _padder__U1122  ( .A1(padder_out[367]), .A2(_padder__n2532 ), .ZN(
        _padder__n1977 ) );
  NAND2_X2 _padder__U1121  ( .A1(_padder__n1976 ), .A2(_padder__n1977 ), .ZN(
        _padder__n1473 ) );
  NAND2_X2 _padder__U1120  ( .A1(padder_out[270]), .A2(_padder__n2501 ), .ZN(
        _padder__n1974 ) );
  NAND2_X2 _padder__U1119  ( .A1(padder_out[366]), .A2(_padder__n2532 ), .ZN(
        _padder__n1975 ) );
  NAND2_X2 _padder__U1118  ( .A1(_padder__n1974 ), .A2(_padder__n1975 ), .ZN(
        _padder__n1474 ) );
  NAND2_X2 _padder__U1117  ( .A1(padder_out[269]), .A2(_padder__n2501 ), .ZN(
        _padder__n1972 ) );
  NAND2_X2 _padder__U1116  ( .A1(padder_out[365]), .A2(_padder__n2532 ), .ZN(
        _padder__n1973 ) );
  NAND2_X2 _padder__U1115  ( .A1(_padder__n1972 ), .A2(_padder__n1973 ), .ZN(
        _padder__n1475 ) );
  NAND2_X2 _padder__U1114  ( .A1(padder_out[268]), .A2(_padder__n2501 ), .ZN(
        _padder__n1970 ) );
  NAND2_X2 _padder__U1113  ( .A1(padder_out[364]), .A2(_padder__n2532 ), .ZN(
        _padder__n1971 ) );
  NAND2_X2 _padder__U1112  ( .A1(_padder__n1970 ), .A2(_padder__n1971 ), .ZN(
        _padder__n1476 ) );
  NAND2_X2 _padder__U1111  ( .A1(padder_out[267]), .A2(_padder__n2501 ), .ZN(
        _padder__n1968 ) );
  NAND2_X2 _padder__U1110  ( .A1(padder_out[363]), .A2(_padder__n2532 ), .ZN(
        _padder__n1969 ) );
  NAND2_X2 _padder__U1109  ( .A1(_padder__n1968 ), .A2(_padder__n1969 ), .ZN(
        _padder__n1477 ) );
  NAND2_X2 _padder__U1108  ( .A1(padder_out[266]), .A2(_padder__n2501 ), .ZN(
        _padder__n1966 ) );
  NAND2_X2 _padder__U1107  ( .A1(padder_out[362]), .A2(_padder__n2532 ), .ZN(
        _padder__n1967 ) );
  NAND2_X2 _padder__U1106  ( .A1(_padder__n1966 ), .A2(_padder__n1967 ), .ZN(
        _padder__n1478 ) );
  NAND2_X2 _padder__U1105  ( .A1(padder_out[265]), .A2(_padder__n2501 ), .ZN(
        _padder__n1964 ) );
  NAND2_X2 _padder__U1104  ( .A1(padder_out[361]), .A2(_padder__n2532 ), .ZN(
        _padder__n1965 ) );
  NAND2_X2 _padder__U1103  ( .A1(_padder__n1964 ), .A2(_padder__n1965 ), .ZN(
        _padder__n1479 ) );
  NAND2_X2 _padder__U1102  ( .A1(padder_out[264]), .A2(_padder__n2501 ), .ZN(
        _padder__n1962 ) );
  NAND2_X2 _padder__U1101  ( .A1(padder_out[360]), .A2(_padder__n2532 ), .ZN(
        _padder__n1963 ) );
  NAND2_X2 _padder__U1100  ( .A1(_padder__n1962 ), .A2(_padder__n1963 ), .ZN(
        _padder__n1480 ) );
  NAND2_X2 _padder__U1099  ( .A1(padder_out[279]), .A2(_padder__n2501 ), .ZN(
        _padder__n1959 ) );
  NAND2_X2 _padder__U1098  ( .A1(padder_out[375]), .A2(_padder__n2532 ), .ZN(
        _padder__n1960 ) );
  NAND2_X2 _padder__U1097  ( .A1(_padder__n1959 ), .A2(_padder__n1960 ), .ZN(
        _padder__n1481 ) );
  NAND2_X2 _padder__U1096  ( .A1(padder_out[278]), .A2(_padder__n2501 ), .ZN(
        _padder__n1957 ) );
  NAND2_X2 _padder__U1095  ( .A1(padder_out[374]), .A2(_padder__n2532 ), .ZN(
        _padder__n1958 ) );
  NAND2_X2 _padder__U1094  ( .A1(_padder__n1957 ), .A2(_padder__n1958 ), .ZN(
        _padder__n1482 ) );
  NAND2_X2 _padder__U1093  ( .A1(padder_out[277]), .A2(_padder__n2501 ), .ZN(
        _padder__n1955 ) );
  NAND2_X2 _padder__U1092  ( .A1(padder_out[373]), .A2(_padder__n2533 ), .ZN(
        _padder__n1956 ) );
  NAND2_X2 _padder__U1091  ( .A1(_padder__n1955 ), .A2(_padder__n1956 ), .ZN(
        _padder__n1483 ) );
  NAND2_X2 _padder__U1090  ( .A1(padder_out[276]), .A2(_padder__n2501 ), .ZN(
        _padder__n1953 ) );
  NAND2_X2 _padder__U1089  ( .A1(padder_out[372]), .A2(_padder__n2533 ), .ZN(
        _padder__n1954 ) );
  NAND2_X2 _padder__U1088  ( .A1(_padder__n1953 ), .A2(_padder__n1954 ), .ZN(
        _padder__n1484 ) );
  NAND2_X2 _padder__U1087  ( .A1(padder_out[275]), .A2(_padder__n2501 ), .ZN(
        _padder__n1951 ) );
  NAND2_X2 _padder__U1086  ( .A1(padder_out[371]), .A2(_padder__n2533 ), .ZN(
        _padder__n1952 ) );
  NAND2_X2 _padder__U1085  ( .A1(_padder__n1951 ), .A2(_padder__n1952 ), .ZN(
        _padder__n1485 ) );
  NAND2_X2 _padder__U1084  ( .A1(padder_out[274]), .A2(_padder__n2501 ), .ZN(
        _padder__n1949 ) );
  NAND2_X2 _padder__U1083  ( .A1(padder_out[370]), .A2(_padder__n2533 ), .ZN(
        _padder__n1950 ) );
  NAND2_X2 _padder__U1082  ( .A1(_padder__n1949 ), .A2(_padder__n1950 ), .ZN(
        _padder__n1486 ) );
  NAND2_X2 _padder__U1081  ( .A1(padder_out[273]), .A2(_padder__n2501 ), .ZN(
        _padder__n1947 ) );
  NAND2_X2 _padder__U1080  ( .A1(padder_out[369]), .A2(_padder__n2533 ), .ZN(
        _padder__n1948 ) );
  NAND2_X2 _padder__U1079  ( .A1(_padder__n1947 ), .A2(_padder__n1948 ), .ZN(
        _padder__n1487 ) );
  NAND2_X2 _padder__U1078  ( .A1(padder_out[272]), .A2(_padder__n2501 ), .ZN(
        _padder__n1945 ) );
  NAND2_X2 _padder__U1077  ( .A1(padder_out[368]), .A2(_padder__n2533 ), .ZN(
        _padder__n1946 ) );
  NAND2_X2 _padder__U1076  ( .A1(_padder__n1945 ), .A2(_padder__n1946 ), .ZN(
        _padder__n1488 ) );
  NAND2_X2 _padder__U1075  ( .A1(padder_out[287]), .A2(_padder__n2501 ), .ZN(
        _padder__n1943 ) );
  NAND2_X2 _padder__U1074  ( .A1(padder_out[383]), .A2(_padder__n2533 ), .ZN(
        _padder__n1944 ) );
  NAND2_X2 _padder__U1073  ( .A1(_padder__n1943 ), .A2(_padder__n1944 ), .ZN(
        _padder__n1489 ) );
  NAND2_X2 _padder__U1072  ( .A1(padder_out[286]), .A2(_padder__n2501 ), .ZN(
        _padder__n1941 ) );
  NAND2_X2 _padder__U1071  ( .A1(padder_out[382]), .A2(_padder__n2533 ), .ZN(
        _padder__n1942 ) );
  NAND2_X2 _padder__U1070  ( .A1(_padder__n1941 ), .A2(_padder__n1942 ), .ZN(
        _padder__n1490 ) );
  NAND2_X2 _padder__U1069  ( .A1(padder_out[285]), .A2(_padder__n2501 ), .ZN(
        _padder__n1939 ) );
  NAND2_X2 _padder__U1068  ( .A1(padder_out[381]), .A2(_padder__n2533 ), .ZN(
        _padder__n1940 ) );
  NAND2_X2 _padder__U1067  ( .A1(_padder__n1939 ), .A2(_padder__n1940 ), .ZN(
        _padder__n1491 ) );
  NAND2_X2 _padder__U1066  ( .A1(padder_out[284]), .A2(_padder__n2501 ), .ZN(
        _padder__n1937 ) );
  NAND2_X2 _padder__U1065  ( .A1(padder_out[380]), .A2(_padder__n2533 ), .ZN(
        _padder__n1938 ) );
  NAND2_X2 _padder__U1064  ( .A1(_padder__n1937 ), .A2(_padder__n1938 ), .ZN(
        _padder__n1492 ) );
  NAND2_X2 _padder__U1063  ( .A1(padder_out[283]), .A2(_padder__n2501 ), .ZN(
        _padder__n1935 ) );
  NAND2_X2 _padder__U1062  ( .A1(padder_out[379]), .A2(_padder__n2533 ), .ZN(
        _padder__n1936 ) );
  NAND2_X2 _padder__U1061  ( .A1(_padder__n1935 ), .A2(_padder__n1936 ), .ZN(
        _padder__n1493 ) );
  NAND2_X2 _padder__U1060  ( .A1(padder_out[282]), .A2(_padder__n2500 ), .ZN(
        _padder__n1933 ) );
  NAND2_X2 _padder__U1059  ( .A1(padder_out[378]), .A2(_padder__n2534 ), .ZN(
        _padder__n1934 ) );
  NAND2_X2 _padder__U1058  ( .A1(_padder__n1933 ), .A2(_padder__n1934 ), .ZN(
        _padder__n1494 ) );
  NAND2_X2 _padder__U1057  ( .A1(padder_out[281]), .A2(_padder__n2500 ), .ZN(
        _padder__n1931 ) );
  NAND2_X2 _padder__U1056  ( .A1(padder_out[377]), .A2(_padder__n2534 ), .ZN(
        _padder__n1932 ) );
  NAND2_X2 _padder__U1055  ( .A1(_padder__n1931 ), .A2(_padder__n1932 ), .ZN(
        _padder__n1495 ) );
  NAND2_X2 _padder__U1054  ( .A1(padder_out[280]), .A2(_padder__n2500 ), .ZN(
        _padder__n1929 ) );
  NAND2_X2 _padder__U1053  ( .A1(padder_out[376]), .A2(_padder__n2534 ), .ZN(
        _padder__n1930 ) );
  NAND2_X2 _padder__U1052  ( .A1(_padder__n1929 ), .A2(_padder__n1930 ), .ZN(
        _padder__n1496 ) );
  NAND2_X2 _padder__U1051  ( .A1(padder_out[295]), .A2(_padder__n2500 ), .ZN(
        _padder__n1927 ) );
  NAND2_X2 _padder__U1050  ( .A1(padder_out[263]), .A2(_padder__n2534 ), .ZN(
        _padder__n1928 ) );
  NAND2_X2 _padder__U1049  ( .A1(_padder__n1927 ), .A2(_padder__n1928 ), .ZN(
        _padder__n1497 ) );
  NAND2_X2 _padder__U1048  ( .A1(padder_out[294]), .A2(_padder__n2500 ), .ZN(
        _padder__n1925 ) );
  NAND2_X2 _padder__U1047  ( .A1(padder_out[262]), .A2(_padder__n2534 ), .ZN(
        _padder__n1926 ) );
  NAND2_X2 _padder__U1046  ( .A1(_padder__n1925 ), .A2(_padder__n1926 ), .ZN(
        _padder__n1498 ) );
  NAND2_X2 _padder__U1045  ( .A1(padder_out[293]), .A2(_padder__n2500 ), .ZN(
        _padder__n1923 ) );
  NAND2_X2 _padder__U1044  ( .A1(padder_out[261]), .A2(_padder__n2534 ), .ZN(
        _padder__n1924 ) );
  NAND2_X2 _padder__U1043  ( .A1(_padder__n1923 ), .A2(_padder__n1924 ), .ZN(
        _padder__n1499 ) );
  NAND2_X2 _padder__U1042  ( .A1(padder_out[292]), .A2(_padder__n2500 ), .ZN(
        _padder__n1921 ) );
  NAND2_X2 _padder__U1041  ( .A1(padder_out[260]), .A2(_padder__n2534 ), .ZN(
        _padder__n1922 ) );
  NAND2_X2 _padder__U1040  ( .A1(_padder__n1921 ), .A2(_padder__n1922 ), .ZN(
        _padder__n1500 ) );
  NAND2_X2 _padder__U1039  ( .A1(padder_out[291]), .A2(_padder__n2500 ), .ZN(
        _padder__n1919 ) );
  NAND2_X2 _padder__U1038  ( .A1(padder_out[259]), .A2(_padder__n2534 ), .ZN(
        _padder__n1920 ) );
  NAND2_X2 _padder__U1037  ( .A1(_padder__n1919 ), .A2(_padder__n1920 ), .ZN(
        _padder__n1501 ) );
  NAND2_X2 _padder__U1036  ( .A1(padder_out[290]), .A2(_padder__n2500 ), .ZN(
        _padder__n1917 ) );
  NAND2_X2 _padder__U1035  ( .A1(padder_out[258]), .A2(_padder__n2534 ), .ZN(
        _padder__n1918 ) );
  NAND2_X2 _padder__U1034  ( .A1(_padder__n1917 ), .A2(_padder__n1918 ), .ZN(
        _padder__n1502 ) );
  NAND2_X2 _padder__U1033  ( .A1(padder_out[289]), .A2(_padder__n2500 ), .ZN(
        _padder__n1915 ) );
  NAND2_X2 _padder__U1032  ( .A1(padder_out[257]), .A2(_padder__n2534 ), .ZN(
        _padder__n1916 ) );
  NAND2_X2 _padder__U1031  ( .A1(_padder__n1915 ), .A2(_padder__n1916 ), .ZN(
        _padder__n1503 ) );
  NAND2_X2 _padder__U1030  ( .A1(padder_out[288]), .A2(_padder__n2500 ), .ZN(
        _padder__n1913 ) );
  NAND2_X2 _padder__U1029  ( .A1(padder_out[256]), .A2(_padder__n2534 ), .ZN(
        _padder__n1914 ) );
  NAND2_X2 _padder__U1028  ( .A1(_padder__n1913 ), .A2(_padder__n1914 ), .ZN(
        _padder__n1504 ) );
  NAND2_X2 _padder__U1027  ( .A1(padder_out[303]), .A2(_padder__n2500 ), .ZN(
        _padder__n1911 ) );
  NAND2_X2 _padder__U1026  ( .A1(padder_out[271]), .A2(_padder__n2535 ), .ZN(
        _padder__n1912 ) );
  NAND2_X2 _padder__U1025  ( .A1(_padder__n1911 ), .A2(_padder__n1912 ), .ZN(
        _padder__n1505 ) );
  NAND2_X2 _padder__U1024  ( .A1(padder_out[302]), .A2(_padder__n2500 ), .ZN(
        _padder__n1909 ) );
  NAND2_X2 _padder__U1023  ( .A1(padder_out[270]), .A2(_padder__n2535 ), .ZN(
        _padder__n1910 ) );
  NAND2_X2 _padder__U1022  ( .A1(_padder__n1909 ), .A2(_padder__n1910 ), .ZN(
        _padder__n1506 ) );
  NAND2_X2 _padder__U1021  ( .A1(padder_out[301]), .A2(_padder__n2500 ), .ZN(
        _padder__n1907 ) );
  NAND2_X2 _padder__U1020  ( .A1(padder_out[269]), .A2(_padder__n2535 ), .ZN(
        _padder__n1908 ) );
  NAND2_X2 _padder__U1019  ( .A1(_padder__n1907 ), .A2(_padder__n1908 ), .ZN(
        _padder__n1507 ) );
  NAND2_X2 _padder__U1018  ( .A1(padder_out[300]), .A2(_padder__n2500 ), .ZN(
        _padder__n1905 ) );
  NAND2_X2 _padder__U1017  ( .A1(padder_out[268]), .A2(_padder__n2535 ), .ZN(
        _padder__n1906 ) );
  NAND2_X2 _padder__U1016  ( .A1(_padder__n1905 ), .A2(_padder__n1906 ), .ZN(
        _padder__n1508 ) );
  NAND2_X2 _padder__U1015  ( .A1(padder_out[299]), .A2(_padder__n2500 ), .ZN(
        _padder__n1903 ) );
  NAND2_X2 _padder__U1014  ( .A1(padder_out[267]), .A2(_padder__n2535 ), .ZN(
        _padder__n1904 ) );
  NAND2_X2 _padder__U1013  ( .A1(_padder__n1903 ), .A2(_padder__n1904 ), .ZN(
        _padder__n1509 ) );
  NAND2_X2 _padder__U1012  ( .A1(padder_out[298]), .A2(_padder__n2500 ), .ZN(
        _padder__n1901 ) );
  NAND2_X2 _padder__U1011  ( .A1(padder_out[266]), .A2(_padder__n2535 ), .ZN(
        _padder__n1902 ) );
  NAND2_X2 _padder__U1010  ( .A1(_padder__n1901 ), .A2(_padder__n1902 ), .ZN(
        _padder__n1510 ) );
  NAND2_X2 _padder__U1009  ( .A1(padder_out[297]), .A2(_padder__n2500 ), .ZN(
        _padder__n1899 ) );
  NAND2_X2 _padder__U1008  ( .A1(padder_out[265]), .A2(_padder__n2535 ), .ZN(
        _padder__n1900 ) );
  NAND2_X2 _padder__U1007  ( .A1(_padder__n1899 ), .A2(_padder__n1900 ), .ZN(
        _padder__n1511 ) );
  NAND2_X2 _padder__U1006  ( .A1(padder_out[296]), .A2(_padder__n2500 ), .ZN(
        _padder__n1897 ) );
  NAND2_X2 _padder__U1005  ( .A1(padder_out[264]), .A2(_padder__n2535 ), .ZN(
        _padder__n1898 ) );
  NAND2_X2 _padder__U1004  ( .A1(_padder__n1897 ), .A2(_padder__n1898 ), .ZN(
        _padder__n1512 ) );
  NAND2_X2 _padder__U1003  ( .A1(padder_out[311]), .A2(_padder__n2503 ), .ZN(
        _padder__n1895 ) );
  NAND2_X2 _padder__U1002  ( .A1(padder_out[279]), .A2(_padder__n2535 ), .ZN(
        _padder__n1896 ) );
  NAND2_X2 _padder__U1001  ( .A1(_padder__n1895 ), .A2(_padder__n1896 ), .ZN(
        _padder__n1513 ) );
  NAND2_X2 _padder__U1000  ( .A1(padder_out[310]), .A2(_padder__n2488 ), .ZN(
        _padder__n1893 ) );
  NAND2_X2 _padder__U999  ( .A1(padder_out[278]), .A2(_padder__n2535 ), .ZN(
        _padder__n1894 ) );
  NAND2_X2 _padder__U998  ( .A1(_padder__n1893 ), .A2(_padder__n1894 ), .ZN(
        _padder__n1514 ) );
  NAND2_X2 _padder__U997  ( .A1(padder_out[309]), .A2(_padder__n2488 ), .ZN(
        _padder__n1891 ) );
  NAND2_X2 _padder__U996  ( .A1(padder_out[277]), .A2(_padder__n2535 ), .ZN(
        _padder__n1892 ) );
  NAND2_X2 _padder__U995  ( .A1(_padder__n1891 ), .A2(_padder__n1892 ), .ZN(
        _padder__n1515 ) );
  NAND2_X2 _padder__U994  ( .A1(padder_out[308]), .A2(_padder__n2488 ), .ZN(
        _padder__n1889 ) );
  NAND2_X2 _padder__U993  ( .A1(padder_out[276]), .A2(_padder__n2536 ), .ZN(
        _padder__n1890 ) );
  NAND2_X2 _padder__U992  ( .A1(_padder__n1889 ), .A2(_padder__n1890 ), .ZN(
        _padder__n1516 ) );
  NAND2_X2 _padder__U991  ( .A1(padder_out[307]), .A2(_padder__n2488 ), .ZN(
        _padder__n1887 ) );
  NAND2_X2 _padder__U990  ( .A1(padder_out[275]), .A2(_padder__n2536 ), .ZN(
        _padder__n1888 ) );
  NAND2_X2 _padder__U989  ( .A1(_padder__n1887 ), .A2(_padder__n1888 ), .ZN(
        _padder__n1517 ) );
  NAND2_X2 _padder__U988  ( .A1(padder_out[306]), .A2(_padder__n2488 ), .ZN(
        _padder__n1885 ) );
  NAND2_X2 _padder__U987  ( .A1(padder_out[274]), .A2(_padder__n2536 ), .ZN(
        _padder__n1886 ) );
  NAND2_X2 _padder__U986  ( .A1(_padder__n1885 ), .A2(_padder__n1886 ), .ZN(
        _padder__n1518 ) );
  NAND2_X2 _padder__U985  ( .A1(padder_out[305]), .A2(_padder__n2488 ), .ZN(
        _padder__n1883 ) );
  NAND2_X2 _padder__U984  ( .A1(padder_out[273]), .A2(_padder__n2536 ), .ZN(
        _padder__n1884 ) );
  NAND2_X2 _padder__U983  ( .A1(_padder__n1883 ), .A2(_padder__n1884 ), .ZN(
        _padder__n1519 ) );
  NAND2_X2 _padder__U982  ( .A1(padder_out[304]), .A2(_padder__n2488 ), .ZN(
        _padder__n1881 ) );
  NAND2_X2 _padder__U981  ( .A1(padder_out[272]), .A2(_padder__n2536 ), .ZN(
        _padder__n1882 ) );
  NAND2_X2 _padder__U980  ( .A1(_padder__n1881 ), .A2(_padder__n1882 ), .ZN(
        _padder__n1520 ) );
  NAND2_X2 _padder__U979  ( .A1(padder_out[319]), .A2(_padder__n2488 ), .ZN(
        _padder__n1879 ) );
  NAND2_X2 _padder__U978  ( .A1(padder_out[287]), .A2(_padder__n2536 ), .ZN(
        _padder__n1880 ) );
  NAND2_X2 _padder__U977  ( .A1(_padder__n1879 ), .A2(_padder__n1880 ), .ZN(
        _padder__n1521 ) );
  NAND2_X2 _padder__U976  ( .A1(padder_out[318]), .A2(_padder__n2488 ), .ZN(
        _padder__n1877 ) );
  NAND2_X2 _padder__U975  ( .A1(padder_out[286]), .A2(_padder__n2536 ), .ZN(
        _padder__n1878 ) );
  NAND2_X2 _padder__U974  ( .A1(_padder__n1877 ), .A2(_padder__n1878 ), .ZN(
        _padder__n1522 ) );
  NAND2_X2 _padder__U973  ( .A1(padder_out[317]), .A2(_padder__n2488 ), .ZN(
        _padder__n1875 ) );
  NAND2_X2 _padder__U972  ( .A1(padder_out[285]), .A2(_padder__n2536 ), .ZN(
        _padder__n1876 ) );
  NAND2_X2 _padder__U971  ( .A1(_padder__n1875 ), .A2(_padder__n1876 ), .ZN(
        _padder__n1523 ) );
  NAND2_X2 _padder__U970  ( .A1(padder_out[316]), .A2(_padder__n2488 ), .ZN(
        _padder__n1873 ) );
  NAND2_X2 _padder__U969  ( .A1(padder_out[284]), .A2(_padder__n2536 ), .ZN(
        _padder__n1874 ) );
  NAND2_X2 _padder__U968  ( .A1(_padder__n1873 ), .A2(_padder__n1874 ), .ZN(
        _padder__n1524 ) );
  NAND2_X2 _padder__U967  ( .A1(padder_out[315]), .A2(_padder__n2488 ), .ZN(
        _padder__n1871 ) );
  NAND2_X2 _padder__U966  ( .A1(padder_out[283]), .A2(_padder__n2536 ), .ZN(
        _padder__n1872 ) );
  NAND2_X2 _padder__U965  ( .A1(_padder__n1871 ), .A2(_padder__n1872 ), .ZN(
        _padder__n1525 ) );
  NAND2_X2 _padder__U964  ( .A1(padder_out[314]), .A2(_padder__n2488 ), .ZN(
        _padder__n1869 ) );
  NAND2_X2 _padder__U963  ( .A1(padder_out[282]), .A2(_padder__n2536 ), .ZN(
        _padder__n1870 ) );
  NAND2_X2 _padder__U962  ( .A1(_padder__n1869 ), .A2(_padder__n1870 ), .ZN(
        _padder__n1526 ) );
  NAND2_X2 _padder__U961  ( .A1(padder_out[313]), .A2(_padder__n2488 ), .ZN(
        _padder__n1867 ) );
  NAND2_X2 _padder__U960  ( .A1(padder_out[281]), .A2(_padder__n2537 ), .ZN(
        _padder__n1868 ) );
  NAND2_X2 _padder__U959  ( .A1(_padder__n1867 ), .A2(_padder__n1868 ), .ZN(
        _padder__n1527 ) );
  NAND2_X2 _padder__U958  ( .A1(padder_out[312]), .A2(_padder__n2488 ), .ZN(
        _padder__n1865 ) );
  NAND2_X2 _padder__U957  ( .A1(padder_out[280]), .A2(_padder__n2537 ), .ZN(
        _padder__n1866 ) );
  NAND2_X2 _padder__U956  ( .A1(_padder__n1865 ), .A2(_padder__n1866 ), .ZN(
        _padder__n1528 ) );
  NAND2_X2 _padder__U955  ( .A1(padder_out[199]), .A2(_padder__n2488 ), .ZN(
        _padder__n1863 ) );
  NAND2_X2 _padder__U954  ( .A1(padder_out[295]), .A2(_padder__n2537 ), .ZN(
        _padder__n1864 ) );
  NAND2_X2 _padder__U953  ( .A1(_padder__n1863 ), .A2(_padder__n1864 ), .ZN(
        _padder__n1529 ) );
  NAND2_X2 _padder__U952  ( .A1(padder_out[198]), .A2(_padder__n2488 ), .ZN(
        _padder__n1861 ) );
  NAND2_X2 _padder__U951  ( .A1(padder_out[294]), .A2(_padder__n2537 ), .ZN(
        _padder__n1862 ) );
  NAND2_X2 _padder__U950  ( .A1(_padder__n1861 ), .A2(_padder__n1862 ), .ZN(
        _padder__n1530 ) );
  NAND2_X2 _padder__U949  ( .A1(padder_out[197]), .A2(_padder__n2488 ), .ZN(
        _padder__n1859 ) );
  NAND2_X2 _padder__U948  ( .A1(padder_out[293]), .A2(_padder__n2537 ), .ZN(
        _padder__n1860 ) );
  NAND2_X2 _padder__U947  ( .A1(_padder__n1859 ), .A2(_padder__n1860 ), .ZN(
        _padder__n1531 ) );
  NAND2_X2 _padder__U946  ( .A1(padder_out[196]), .A2(_padder__n2488 ), .ZN(
        _padder__n1857 ) );
  NAND2_X2 _padder__U945  ( .A1(padder_out[292]), .A2(_padder__n2537 ), .ZN(
        _padder__n1858 ) );
  NAND2_X2 _padder__U944  ( .A1(_padder__n1857 ), .A2(_padder__n1858 ), .ZN(
        _padder__n1532 ) );
  NAND2_X2 _padder__U943  ( .A1(padder_out[195]), .A2(_padder__n2488 ), .ZN(
        _padder__n1855 ) );
  NAND2_X2 _padder__U942  ( .A1(padder_out[291]), .A2(_padder__n2537 ), .ZN(
        _padder__n1856 ) );
  NAND2_X2 _padder__U941  ( .A1(_padder__n1855 ), .A2(_padder__n1856 ), .ZN(
        _padder__n1533 ) );
  NAND2_X2 _padder__U940  ( .A1(padder_out[194]), .A2(_padder__n2488 ), .ZN(
        _padder__n1853 ) );
  NAND2_X2 _padder__U939  ( .A1(padder_out[290]), .A2(_padder__n2537 ), .ZN(
        _padder__n1854 ) );
  NAND2_X2 _padder__U938  ( .A1(_padder__n1853 ), .A2(_padder__n1854 ), .ZN(
        _padder__n1534 ) );
  NAND2_X2 _padder__U937  ( .A1(padder_out[193]), .A2(_padder__n2487 ), .ZN(
        _padder__n1851 ) );
  NAND2_X2 _padder__U936  ( .A1(padder_out[289]), .A2(_padder__n2537 ), .ZN(
        _padder__n1852 ) );
  NAND2_X2 _padder__U935  ( .A1(_padder__n1851 ), .A2(_padder__n1852 ), .ZN(
        _padder__n1535 ) );
  NAND2_X2 _padder__U934  ( .A1(padder_out[192]), .A2(_padder__n2487 ), .ZN(
        _padder__n1849 ) );
  NAND2_X2 _padder__U933  ( .A1(padder_out[288]), .A2(_padder__n2537 ), .ZN(
        _padder__n1850 ) );
  NAND2_X2 _padder__U932  ( .A1(_padder__n1849 ), .A2(_padder__n1850 ), .ZN(
        _padder__n1536 ) );
  NAND2_X2 _padder__U931  ( .A1(padder_out[207]), .A2(_padder__n2487 ), .ZN(
        _padder__n1847 ) );
  NAND2_X2 _padder__U930  ( .A1(padder_out[303]), .A2(_padder__n2537 ), .ZN(
        _padder__n1848 ) );
  NAND2_X2 _padder__U929  ( .A1(_padder__n1847 ), .A2(_padder__n1848 ), .ZN(
        _padder__n1537 ) );
  NAND2_X2 _padder__U928  ( .A1(padder_out[206]), .A2(_padder__n2487 ), .ZN(
        _padder__n1845 ) );
  NAND2_X2 _padder__U927  ( .A1(padder_out[302]), .A2(_padder__n2538 ), .ZN(
        _padder__n1846 ) );
  NAND2_X2 _padder__U926  ( .A1(_padder__n1845 ), .A2(_padder__n1846 ), .ZN(
        _padder__n1538 ) );
  NAND2_X2 _padder__U925  ( .A1(padder_out[205]), .A2(_padder__n2487 ), .ZN(
        _padder__n1843 ) );
  NAND2_X2 _padder__U924  ( .A1(padder_out[301]), .A2(_padder__n2538 ), .ZN(
        _padder__n1844 ) );
  NAND2_X2 _padder__U923  ( .A1(_padder__n1843 ), .A2(_padder__n1844 ), .ZN(
        _padder__n1539 ) );
  NAND2_X2 _padder__U922  ( .A1(padder_out[204]), .A2(_padder__n2487 ), .ZN(
        _padder__n1841 ) );
  NAND2_X2 _padder__U921  ( .A1(padder_out[300]), .A2(_padder__n2538 ), .ZN(
        _padder__n1842 ) );
  NAND2_X2 _padder__U920  ( .A1(_padder__n1841 ), .A2(_padder__n1842 ), .ZN(
        _padder__n1540 ) );
  NAND2_X2 _padder__U919  ( .A1(padder_out[203]), .A2(_padder__n2487 ), .ZN(
        _padder__n1839 ) );
  NAND2_X2 _padder__U918  ( .A1(padder_out[299]), .A2(_padder__n2538 ), .ZN(
        _padder__n1840 ) );
  NAND2_X2 _padder__U917  ( .A1(_padder__n1839 ), .A2(_padder__n1840 ), .ZN(
        _padder__n1541 ) );
  NAND2_X2 _padder__U916  ( .A1(padder_out[202]), .A2(_padder__n2487 ), .ZN(
        _padder__n1837 ) );
  NAND2_X2 _padder__U915  ( .A1(padder_out[298]), .A2(_padder__n2538 ), .ZN(
        _padder__n1838 ) );
  NAND2_X2 _padder__U914  ( .A1(_padder__n1837 ), .A2(_padder__n1838 ), .ZN(
        _padder__n1542 ) );
  NAND2_X2 _padder__U913  ( .A1(padder_out[201]), .A2(_padder__n2487 ), .ZN(
        _padder__n1239 ) );
  NAND2_X2 _padder__U912  ( .A1(padder_out[297]), .A2(_padder__n2538 ), .ZN(
        _padder__n1240 ) );
  NAND2_X2 _padder__U911  ( .A1(_padder__n1239 ), .A2(_padder__n1240 ), .ZN(
        _padder__n1543 ) );
  NAND2_X2 _padder__U910  ( .A1(padder_out[200]), .A2(_padder__n2487 ), .ZN(
        _padder__n1237 ) );
  NAND2_X2 _padder__U909  ( .A1(padder_out[296]), .A2(_padder__n2538 ), .ZN(
        _padder__n1238 ) );
  NAND2_X2 _padder__U908  ( .A1(_padder__n1237 ), .A2(_padder__n1238 ), .ZN(
        _padder__n1544 ) );
  NAND2_X2 _padder__U907  ( .A1(padder_out[215]), .A2(_padder__n2487 ), .ZN(
        _padder__n1235 ) );
  NAND2_X2 _padder__U906  ( .A1(padder_out[311]), .A2(_padder__n2538 ), .ZN(
        _padder__n1236 ) );
  NAND2_X2 _padder__U905  ( .A1(_padder__n1235 ), .A2(_padder__n1236 ), .ZN(
        _padder__n1545 ) );
  NAND2_X2 _padder__U904  ( .A1(padder_out[214]), .A2(_padder__n2487 ), .ZN(
        _padder__n1233 ) );
  NAND2_X2 _padder__U903  ( .A1(padder_out[310]), .A2(_padder__n2538 ), .ZN(
        _padder__n1234 ) );
  NAND2_X2 _padder__U902  ( .A1(_padder__n1233 ), .A2(_padder__n1234 ), .ZN(
        _padder__n1546 ) );
  NAND2_X2 _padder__U901  ( .A1(padder_out[213]), .A2(_padder__n2487 ), .ZN(
        _padder__n1231 ) );
  NAND2_X2 _padder__U900  ( .A1(padder_out[309]), .A2(_padder__n2538 ), .ZN(
        _padder__n1232 ) );
  NAND2_X2 _padder__U899  ( .A1(_padder__n1231 ), .A2(_padder__n1232 ), .ZN(
        _padder__n1547 ) );
  NAND2_X2 _padder__U898  ( .A1(padder_out[212]), .A2(_padder__n2487 ), .ZN(
        _padder__n1229 ) );
  NAND2_X2 _padder__U897  ( .A1(padder_out[308]), .A2(_padder__n2538 ), .ZN(
        _padder__n1230 ) );
  NAND2_X2 _padder__U896  ( .A1(_padder__n1229 ), .A2(_padder__n1230 ), .ZN(
        _padder__n1548 ) );
  NAND2_X2 _padder__U895  ( .A1(padder_out[211]), .A2(_padder__n2487 ), .ZN(
        _padder__n1227 ) );
  NAND2_X2 _padder__U894  ( .A1(padder_out[307]), .A2(_padder__n2539 ), .ZN(
        _padder__n1228 ) );
  NAND2_X2 _padder__U893  ( .A1(_padder__n1227 ), .A2(_padder__n1228 ), .ZN(
        _padder__n1549 ) );
  NAND2_X2 _padder__U892  ( .A1(padder_out[210]), .A2(_padder__n2487 ), .ZN(
        _padder__n1225 ) );
  NAND2_X2 _padder__U891  ( .A1(padder_out[306]), .A2(_padder__n2539 ), .ZN(
        _padder__n1226 ) );
  NAND2_X2 _padder__U890  ( .A1(_padder__n1225 ), .A2(_padder__n1226 ), .ZN(
        _padder__n1550 ) );
  NAND2_X2 _padder__U889  ( .A1(padder_out[209]), .A2(_padder__n2487 ), .ZN(
        _padder__n1223 ) );
  NAND2_X2 _padder__U888  ( .A1(padder_out[305]), .A2(_padder__n2539 ), .ZN(
        _padder__n1224 ) );
  NAND2_X2 _padder__U887  ( .A1(_padder__n1223 ), .A2(_padder__n1224 ), .ZN(
        _padder__n1551 ) );
  NAND2_X2 _padder__U886  ( .A1(padder_out[208]), .A2(_padder__n2487 ), .ZN(
        _padder__n1221 ) );
  NAND2_X2 _padder__U885  ( .A1(padder_out[304]), .A2(_padder__n2539 ), .ZN(
        _padder__n1222 ) );
  NAND2_X2 _padder__U884  ( .A1(_padder__n1221 ), .A2(_padder__n1222 ), .ZN(
        _padder__n1552 ) );
  NAND2_X2 _padder__U883  ( .A1(padder_out[223]), .A2(_padder__n2487 ), .ZN(
        _padder__n1219 ) );
  NAND2_X2 _padder__U882  ( .A1(padder_out[319]), .A2(_padder__n2539 ), .ZN(
        _padder__n1220 ) );
  NAND2_X2 _padder__U881  ( .A1(_padder__n1219 ), .A2(_padder__n1220 ), .ZN(
        _padder__n1553 ) );
  NAND2_X2 _padder__U880  ( .A1(padder_out[222]), .A2(_padder__n2487 ), .ZN(
        _padder__n1217 ) );
  NAND2_X2 _padder__U879  ( .A1(padder_out[318]), .A2(_padder__n2539 ), .ZN(
        _padder__n1218 ) );
  NAND2_X2 _padder__U878  ( .A1(_padder__n1217 ), .A2(_padder__n1218 ), .ZN(
        _padder__n1554 ) );
  NAND2_X2 _padder__U877  ( .A1(padder_out[221]), .A2(_padder__n2487 ), .ZN(
        _padder__n1215 ) );
  NAND2_X2 _padder__U876  ( .A1(padder_out[317]), .A2(_padder__n2539 ), .ZN(
        _padder__n1216 ) );
  NAND2_X2 _padder__U875  ( .A1(_padder__n1215 ), .A2(_padder__n1216 ), .ZN(
        _padder__n1555 ) );
  NAND2_X2 _padder__U874  ( .A1(padder_out[220]), .A2(_padder__n2487 ), .ZN(
        _padder__n1213 ) );
  NAND2_X2 _padder__U873  ( .A1(padder_out[316]), .A2(_padder__n2539 ), .ZN(
        _padder__n1214 ) );
  NAND2_X2 _padder__U872  ( .A1(_padder__n1213 ), .A2(_padder__n1214 ), .ZN(
        _padder__n1556 ) );
  NAND2_X2 _padder__U871  ( .A1(padder_out[219]), .A2(_padder__n2487 ), .ZN(
        _padder__n1211 ) );
  NAND2_X2 _padder__U870  ( .A1(padder_out[315]), .A2(_padder__n2539 ), .ZN(
        _padder__n1212 ) );
  NAND2_X2 _padder__U869  ( .A1(_padder__n1211 ), .A2(_padder__n1212 ), .ZN(
        _padder__n1557 ) );
  NAND2_X2 _padder__U868  ( .A1(padder_out[218]), .A2(_padder__n2487 ), .ZN(
        _padder__n1209 ) );
  NAND2_X2 _padder__U867  ( .A1(padder_out[314]), .A2(_padder__n2539 ), .ZN(
        _padder__n1210 ) );
  NAND2_X2 _padder__U866  ( .A1(_padder__n1209 ), .A2(_padder__n1210 ), .ZN(
        _padder__n1558 ) );
  NAND2_X2 _padder__U865  ( .A1(padder_out[217]), .A2(_padder__n2486 ), .ZN(
        _padder__n1207 ) );
  NAND2_X2 _padder__U864  ( .A1(padder_out[313]), .A2(_padder__n2539 ), .ZN(
        _padder__n1208 ) );
  NAND2_X2 _padder__U863  ( .A1(_padder__n1207 ), .A2(_padder__n1208 ), .ZN(
        _padder__n1559 ) );
  NAND2_X2 _padder__U862  ( .A1(padder_out[216]), .A2(_padder__n2486 ), .ZN(
        _padder__n1205 ) );
  NAND2_X2 _padder__U861  ( .A1(padder_out[312]), .A2(_padder__n2540 ), .ZN(
        _padder__n1206 ) );
  NAND2_X2 _padder__U860  ( .A1(_padder__n1205 ), .A2(_padder__n1206 ), .ZN(
        _padder__n1560 ) );
  NAND2_X2 _padder__U859  ( .A1(padder_out[231]), .A2(_padder__n2486 ), .ZN(
        _padder__n1203 ) );
  NAND2_X2 _padder__U858  ( .A1(padder_out[199]), .A2(_padder__n2540 ), .ZN(
        _padder__n1204 ) );
  NAND2_X2 _padder__U857  ( .A1(_padder__n1203 ), .A2(_padder__n1204 ), .ZN(
        _padder__n1561 ) );
  NAND2_X2 _padder__U856  ( .A1(padder_out[230]), .A2(_padder__n2486 ), .ZN(
        _padder__n1201 ) );
  NAND2_X2 _padder__U855  ( .A1(padder_out[198]), .A2(_padder__n2540 ), .ZN(
        _padder__n1202 ) );
  NAND2_X2 _padder__U854  ( .A1(_padder__n1201 ), .A2(_padder__n1202 ), .ZN(
        _padder__n1562 ) );
  NAND2_X2 _padder__U853  ( .A1(padder_out[229]), .A2(_padder__n2486 ), .ZN(
        _padder__n1199 ) );
  NAND2_X2 _padder__U852  ( .A1(padder_out[197]), .A2(_padder__n2540 ), .ZN(
        _padder__n1200 ) );
  NAND2_X2 _padder__U851  ( .A1(_padder__n1199 ), .A2(_padder__n1200 ), .ZN(
        _padder__n1563 ) );
  NAND2_X2 _padder__U850  ( .A1(padder_out[228]), .A2(_padder__n2486 ), .ZN(
        _padder__n1197 ) );
  NAND2_X2 _padder__U849  ( .A1(padder_out[196]), .A2(_padder__n2540 ), .ZN(
        _padder__n1198 ) );
  NAND2_X2 _padder__U848  ( .A1(_padder__n1197 ), .A2(_padder__n1198 ), .ZN(
        _padder__n1564 ) );
  NAND2_X2 _padder__U847  ( .A1(padder_out[227]), .A2(_padder__n2486 ), .ZN(
        _padder__n1195 ) );
  NAND2_X2 _padder__U846  ( .A1(padder_out[195]), .A2(_padder__n2540 ), .ZN(
        _padder__n1196 ) );
  NAND2_X2 _padder__U845  ( .A1(_padder__n1195 ), .A2(_padder__n1196 ), .ZN(
        _padder__n1565 ) );
  NAND2_X2 _padder__U844  ( .A1(padder_out[226]), .A2(_padder__n2486 ), .ZN(
        _padder__n1193 ) );
  NAND2_X2 _padder__U843  ( .A1(padder_out[194]), .A2(_padder__n2540 ), .ZN(
        _padder__n1194 ) );
  NAND2_X2 _padder__U842  ( .A1(_padder__n1193 ), .A2(_padder__n1194 ), .ZN(
        _padder__n1566 ) );
  NAND2_X2 _padder__U841  ( .A1(padder_out[225]), .A2(_padder__n2486 ), .ZN(
        _padder__n1191 ) );
  NAND2_X2 _padder__U840  ( .A1(padder_out[193]), .A2(_padder__n2540 ), .ZN(
        _padder__n1192 ) );
  NAND2_X2 _padder__U839  ( .A1(_padder__n1191 ), .A2(_padder__n1192 ), .ZN(
        _padder__n1567 ) );
  NAND2_X2 _padder__U838  ( .A1(padder_out[224]), .A2(_padder__n2486 ), .ZN(
        _padder__n1189 ) );
  NAND2_X2 _padder__U837  ( .A1(padder_out[192]), .A2(_padder__n2540 ), .ZN(
        _padder__n1190 ) );
  NAND2_X2 _padder__U836  ( .A1(_padder__n1189 ), .A2(_padder__n1190 ), .ZN(
        _padder__n1568 ) );
  NAND2_X2 _padder__U835  ( .A1(padder_out[239]), .A2(_padder__n2486 ), .ZN(
        _padder__n1187 ) );
  NAND2_X2 _padder__U834  ( .A1(padder_out[207]), .A2(_padder__n2540 ), .ZN(
        _padder__n1188 ) );
  NAND2_X2 _padder__U833  ( .A1(_padder__n1187 ), .A2(_padder__n1188 ), .ZN(
        _padder__n1569 ) );
  NAND2_X2 _padder__U832  ( .A1(padder_out[238]), .A2(_padder__n2486 ), .ZN(
        _padder__n1185 ) );
  NAND2_X2 _padder__U831  ( .A1(padder_out[206]), .A2(_padder__n2540 ), .ZN(
        _padder__n1186 ) );
  NAND2_X2 _padder__U830  ( .A1(_padder__n1185 ), .A2(_padder__n1186 ), .ZN(
        _padder__n1570 ) );
  NAND2_X2 _padder__U829  ( .A1(padder_out[237]), .A2(_padder__n2486 ), .ZN(
        _padder__n1183 ) );
  NAND2_X2 _padder__U828  ( .A1(padder_out[205]), .A2(_padder__n2541 ), .ZN(
        _padder__n1184 ) );
  NAND2_X2 _padder__U827  ( .A1(_padder__n1183 ), .A2(_padder__n1184 ), .ZN(
        _padder__n1571 ) );
  NAND2_X2 _padder__U826  ( .A1(padder_out[236]), .A2(_padder__n2486 ), .ZN(
        _padder__n1181 ) );
  NAND2_X2 _padder__U825  ( .A1(padder_out[204]), .A2(_padder__n2541 ), .ZN(
        _padder__n1182 ) );
  NAND2_X2 _padder__U824  ( .A1(_padder__n1181 ), .A2(_padder__n1182 ), .ZN(
        _padder__n1572 ) );
  NAND2_X2 _padder__U823  ( .A1(padder_out[235]), .A2(_padder__n2486 ), .ZN(
        _padder__n1179 ) );
  NAND2_X2 _padder__U822  ( .A1(padder_out[203]), .A2(_padder__n2541 ), .ZN(
        _padder__n1180 ) );
  NAND2_X2 _padder__U821  ( .A1(_padder__n1179 ), .A2(_padder__n1180 ), .ZN(
        _padder__n1573 ) );
  NAND2_X2 _padder__U820  ( .A1(padder_out[234]), .A2(_padder__n2486 ), .ZN(
        _padder__n1177 ) );
  NAND2_X2 _padder__U819  ( .A1(padder_out[202]), .A2(_padder__n2541 ), .ZN(
        _padder__n1178 ) );
  NAND2_X2 _padder__U818  ( .A1(_padder__n1177 ), .A2(_padder__n1178 ), .ZN(
        _padder__n1574 ) );
  NAND2_X2 _padder__U817  ( .A1(padder_out[233]), .A2(_padder__n2486 ), .ZN(
        _padder__n1175 ) );
  NAND2_X2 _padder__U816  ( .A1(padder_out[201]), .A2(_padder__n2541 ), .ZN(
        _padder__n1176 ) );
  NAND2_X2 _padder__U815  ( .A1(_padder__n1175 ), .A2(_padder__n1176 ), .ZN(
        _padder__n1575 ) );
  NAND2_X2 _padder__U814  ( .A1(padder_out[232]), .A2(_padder__n2486 ), .ZN(
        _padder__n1173 ) );
  NAND2_X2 _padder__U813  ( .A1(padder_out[200]), .A2(_padder__n2541 ), .ZN(
        _padder__n1174 ) );
  NAND2_X2 _padder__U812  ( .A1(_padder__n1173 ), .A2(_padder__n1174 ), .ZN(
        _padder__n1576 ) );
  NAND2_X2 _padder__U811  ( .A1(padder_out[247]), .A2(_padder__n2486 ), .ZN(
        _padder__n1171 ) );
  NAND2_X2 _padder__U810  ( .A1(padder_out[215]), .A2(_padder__n2541 ), .ZN(
        _padder__n1172 ) );
  NAND2_X2 _padder__U809  ( .A1(_padder__n1171 ), .A2(_padder__n1172 ), .ZN(
        _padder__n1577 ) );
  NAND2_X2 _padder__U808  ( .A1(padder_out[246]), .A2(_padder__n2486 ), .ZN(
        _padder__n1169 ) );
  NAND2_X2 _padder__U807  ( .A1(padder_out[214]), .A2(_padder__n2541 ), .ZN(
        _padder__n1170 ) );
  NAND2_X2 _padder__U806  ( .A1(_padder__n1169 ), .A2(_padder__n1170 ), .ZN(
        _padder__n1578 ) );
  NAND2_X2 _padder__U805  ( .A1(padder_out[245]), .A2(_padder__n2486 ), .ZN(
        _padder__n1167 ) );
  NAND2_X2 _padder__U804  ( .A1(padder_out[213]), .A2(_padder__n2541 ), .ZN(
        _padder__n1168 ) );
  NAND2_X2 _padder__U803  ( .A1(_padder__n1167 ), .A2(_padder__n1168 ), .ZN(
        _padder__n1579 ) );
  NAND2_X2 _padder__U802  ( .A1(padder_out[244]), .A2(_padder__n2486 ), .ZN(
        _padder__n1165 ) );
  NAND2_X2 _padder__U801  ( .A1(padder_out[212]), .A2(_padder__n2541 ), .ZN(
        _padder__n1166 ) );
  NAND2_X2 _padder__U800  ( .A1(_padder__n1165 ), .A2(_padder__n1166 ), .ZN(
        _padder__n1580 ) );
  NAND2_X2 _padder__U799  ( .A1(padder_out[243]), .A2(_padder__n2486 ), .ZN(
        _padder__n1163 ) );
  NAND2_X2 _padder__U798  ( .A1(padder_out[211]), .A2(_padder__n2541 ), .ZN(
        _padder__n1164 ) );
  NAND2_X2 _padder__U797  ( .A1(_padder__n1163 ), .A2(_padder__n1164 ), .ZN(
        _padder__n1581 ) );
  NAND2_X2 _padder__U796  ( .A1(padder_out[242]), .A2(_padder__n2485 ), .ZN(
        _padder__n1161 ) );
  NAND2_X2 _padder__U795  ( .A1(padder_out[210]), .A2(_padder__n2542 ), .ZN(
        _padder__n1162 ) );
  NAND2_X2 _padder__U794  ( .A1(_padder__n1161 ), .A2(_padder__n1162 ), .ZN(
        _padder__n1582 ) );
  NAND2_X2 _padder__U793  ( .A1(padder_out[241]), .A2(_padder__n2485 ), .ZN(
        _padder__n1159 ) );
  NAND2_X2 _padder__U792  ( .A1(padder_out[209]), .A2(_padder__n2542 ), .ZN(
        _padder__n1160 ) );
  NAND2_X2 _padder__U791  ( .A1(_padder__n1159 ), .A2(_padder__n1160 ), .ZN(
        _padder__n1583 ) );
  NAND2_X2 _padder__U790  ( .A1(padder_out[240]), .A2(_padder__n2485 ), .ZN(
        _padder__n1157 ) );
  NAND2_X2 _padder__U789  ( .A1(padder_out[208]), .A2(_padder__n2542 ), .ZN(
        _padder__n1158 ) );
  NAND2_X2 _padder__U788  ( .A1(_padder__n1157 ), .A2(_padder__n1158 ), .ZN(
        _padder__n1584 ) );
  NAND2_X2 _padder__U787  ( .A1(padder_out[255]), .A2(_padder__n2485 ), .ZN(
        _padder__n1155 ) );
  NAND2_X2 _padder__U786  ( .A1(padder_out[223]), .A2(_padder__n2542 ), .ZN(
        _padder__n1156 ) );
  NAND2_X2 _padder__U785  ( .A1(_padder__n1155 ), .A2(_padder__n1156 ), .ZN(
        _padder__n1585 ) );
  NAND2_X2 _padder__U784  ( .A1(padder_out[254]), .A2(_padder__n2485 ), .ZN(
        _padder__n1153 ) );
  NAND2_X2 _padder__U783  ( .A1(padder_out[222]), .A2(_padder__n2542 ), .ZN(
        _padder__n1154 ) );
  NAND2_X2 _padder__U782  ( .A1(_padder__n1153 ), .A2(_padder__n1154 ), .ZN(
        _padder__n1586 ) );
  NAND2_X2 _padder__U781  ( .A1(padder_out[253]), .A2(_padder__n2485 ), .ZN(
        _padder__n1151 ) );
  NAND2_X2 _padder__U780  ( .A1(padder_out[221]), .A2(_padder__n2542 ), .ZN(
        _padder__n1152 ) );
  NAND2_X2 _padder__U779  ( .A1(_padder__n1151 ), .A2(_padder__n1152 ), .ZN(
        _padder__n1587 ) );
  NAND2_X2 _padder__U778  ( .A1(padder_out[252]), .A2(_padder__n2485 ), .ZN(
        _padder__n1149 ) );
  NAND2_X2 _padder__U777  ( .A1(padder_out[220]), .A2(_padder__n2542 ), .ZN(
        _padder__n1150 ) );
  NAND2_X2 _padder__U776  ( .A1(_padder__n1149 ), .A2(_padder__n1150 ), .ZN(
        _padder__n1588 ) );
  NAND2_X2 _padder__U775  ( .A1(padder_out[251]), .A2(_padder__n2485 ), .ZN(
        _padder__n1147 ) );
  NAND2_X2 _padder__U774  ( .A1(padder_out[219]), .A2(_padder__n2542 ), .ZN(
        _padder__n1148 ) );
  NAND2_X2 _padder__U773  ( .A1(_padder__n1147 ), .A2(_padder__n1148 ), .ZN(
        _padder__n1589 ) );
  NAND2_X2 _padder__U772  ( .A1(padder_out[250]), .A2(_padder__n2485 ), .ZN(
        _padder__n1145 ) );
  NAND2_X2 _padder__U771  ( .A1(padder_out[218]), .A2(_padder__n2542 ), .ZN(
        _padder__n1146 ) );
  NAND2_X2 _padder__U770  ( .A1(_padder__n1145 ), .A2(_padder__n1146 ), .ZN(
        _padder__n1590 ) );
  NAND2_X2 _padder__U769  ( .A1(padder_out[249]), .A2(_padder__n2485 ), .ZN(
        _padder__n1143 ) );
  NAND2_X2 _padder__U768  ( .A1(padder_out[217]), .A2(_padder__n2542 ), .ZN(
        _padder__n1144 ) );
  NAND2_X2 _padder__U767  ( .A1(_padder__n1143 ), .A2(_padder__n1144 ), .ZN(
        _padder__n1591 ) );
  NAND2_X2 _padder__U766  ( .A1(padder_out[248]), .A2(_padder__n2485 ), .ZN(
        _padder__n1141 ) );
  NAND2_X2 _padder__U765  ( .A1(padder_out[216]), .A2(_padder__n2542 ), .ZN(
        _padder__n1142 ) );
  NAND2_X2 _padder__U764  ( .A1(_padder__n1141 ), .A2(_padder__n1142 ), .ZN(
        _padder__n1592 ) );
  NAND2_X2 _padder__U763  ( .A1(padder_out[135]), .A2(_padder__n2485 ), .ZN(
        _padder__n1139 ) );
  NAND2_X2 _padder__U762  ( .A1(padder_out[231]), .A2(_padder__n2543 ), .ZN(
        _padder__n1140 ) );
  NAND2_X2 _padder__U761  ( .A1(_padder__n1139 ), .A2(_padder__n1140 ), .ZN(
        _padder__n1593 ) );
  NAND2_X2 _padder__U760  ( .A1(padder_out[134]), .A2(_padder__n2485 ), .ZN(
        _padder__n1137 ) );
  NAND2_X2 _padder__U759  ( .A1(padder_out[230]), .A2(_padder__n2543 ), .ZN(
        _padder__n1138 ) );
  NAND2_X2 _padder__U758  ( .A1(_padder__n1137 ), .A2(_padder__n1138 ), .ZN(
        _padder__n1594 ) );
  NAND2_X2 _padder__U757  ( .A1(padder_out[133]), .A2(_padder__n2485 ), .ZN(
        _padder__n1135 ) );
  NAND2_X2 _padder__U756  ( .A1(padder_out[229]), .A2(_padder__n2543 ), .ZN(
        _padder__n1136 ) );
  NAND2_X2 _padder__U755  ( .A1(_padder__n1135 ), .A2(_padder__n1136 ), .ZN(
        _padder__n1595 ) );
  NAND2_X2 _padder__U754  ( .A1(padder_out[132]), .A2(_padder__n2485 ), .ZN(
        _padder__n1133 ) );
  NAND2_X2 _padder__U753  ( .A1(padder_out[228]), .A2(_padder__n2543 ), .ZN(
        _padder__n1134 ) );
  NAND2_X2 _padder__U752  ( .A1(_padder__n1133 ), .A2(_padder__n1134 ), .ZN(
        _padder__n1596 ) );
  NAND2_X2 _padder__U751  ( .A1(padder_out[131]), .A2(_padder__n2485 ), .ZN(
        _padder__n1131 ) );
  NAND2_X2 _padder__U750  ( .A1(padder_out[227]), .A2(_padder__n2543 ), .ZN(
        _padder__n1132 ) );
  NAND2_X2 _padder__U749  ( .A1(_padder__n1131 ), .A2(_padder__n1132 ), .ZN(
        _padder__n1597 ) );
  NAND2_X2 _padder__U748  ( .A1(padder_out[130]), .A2(_padder__n2485 ), .ZN(
        _padder__n1129 ) );
  NAND2_X2 _padder__U747  ( .A1(padder_out[226]), .A2(_padder__n2543 ), .ZN(
        _padder__n1130 ) );
  NAND2_X2 _padder__U746  ( .A1(_padder__n1129 ), .A2(_padder__n1130 ), .ZN(
        _padder__n1598 ) );
  NAND2_X2 _padder__U745  ( .A1(padder_out[129]), .A2(_padder__n2485 ), .ZN(
        _padder__n1127 ) );
  NAND2_X2 _padder__U744  ( .A1(padder_out[225]), .A2(_padder__n2543 ), .ZN(
        _padder__n1128 ) );
  NAND2_X2 _padder__U743  ( .A1(_padder__n1127 ), .A2(_padder__n1128 ), .ZN(
        _padder__n1599 ) );
  NAND2_X2 _padder__U742  ( .A1(padder_out[128]), .A2(_padder__n2485 ), .ZN(
        _padder__n1125 ) );
  NAND2_X2 _padder__U741  ( .A1(padder_out[224]), .A2(_padder__n2543 ), .ZN(
        _padder__n1126 ) );
  NAND2_X2 _padder__U740  ( .A1(_padder__n1125 ), .A2(_padder__n1126 ), .ZN(
        _padder__n1600 ) );
  NAND2_X2 _padder__U739  ( .A1(padder_out[143]), .A2(_padder__n2485 ), .ZN(
        _padder__n1123 ) );
  NAND2_X2 _padder__U738  ( .A1(padder_out[239]), .A2(_padder__n2543 ), .ZN(
        _padder__n1124 ) );
  NAND2_X2 _padder__U737  ( .A1(_padder__n1123 ), .A2(_padder__n1124 ), .ZN(
        _padder__n1601 ) );
  NAND2_X2 _padder__U736  ( .A1(padder_out[142]), .A2(_padder__n2485 ), .ZN(
        _padder__n1121 ) );
  NAND2_X2 _padder__U735  ( .A1(padder_out[238]), .A2(_padder__n2543 ), .ZN(
        _padder__n1122 ) );
  NAND2_X2 _padder__U734  ( .A1(_padder__n1121 ), .A2(_padder__n1122 ), .ZN(
        _padder__n1602 ) );
  NAND2_X2 _padder__U733  ( .A1(padder_out[141]), .A2(_padder__n2485 ), .ZN(
        _padder__n1119 ) );
  NAND2_X2 _padder__U732  ( .A1(padder_out[237]), .A2(_padder__n2543 ), .ZN(
        _padder__n1120 ) );
  NAND2_X2 _padder__U731  ( .A1(_padder__n1119 ), .A2(_padder__n1120 ), .ZN(
        _padder__n1603 ) );
  NAND2_X2 _padder__U730  ( .A1(padder_out[140]), .A2(_padder__n2485 ), .ZN(
        _padder__n1117 ) );
  NAND2_X2 _padder__U729  ( .A1(padder_out[236]), .A2(_padder__n2544 ), .ZN(
        _padder__n1118 ) );
  NAND2_X2 _padder__U728  ( .A1(_padder__n1117 ), .A2(_padder__n1118 ), .ZN(
        _padder__n1604 ) );
  NAND2_X2 _padder__U727  ( .A1(padder_out[139]), .A2(_padder__n2485 ), .ZN(
        _padder__n1115 ) );
  NAND2_X2 _padder__U726  ( .A1(padder_out[235]), .A2(_padder__n2544 ), .ZN(
        _padder__n1116 ) );
  NAND2_X2 _padder__U725  ( .A1(_padder__n1115 ), .A2(_padder__n1116 ), .ZN(
        _padder__n1605 ) );
  NAND2_X2 _padder__U724  ( .A1(padder_out[138]), .A2(_padder__n2505 ), .ZN(
        _padder__n1113 ) );
  NAND2_X2 _padder__U723  ( .A1(padder_out[234]), .A2(_padder__n2544 ), .ZN(
        _padder__n1114 ) );
  NAND2_X2 _padder__U722  ( .A1(_padder__n1113 ), .A2(_padder__n1114 ), .ZN(
        _padder__n1606 ) );
  NAND2_X2 _padder__U721  ( .A1(padder_out[137]), .A2(_padder__n2505 ), .ZN(
        _padder__n1111 ) );
  NAND2_X2 _padder__U720  ( .A1(padder_out[233]), .A2(_padder__n2544 ), .ZN(
        _padder__n1112 ) );
  NAND2_X2 _padder__U719  ( .A1(_padder__n1111 ), .A2(_padder__n1112 ), .ZN(
        _padder__n1607 ) );
  NAND2_X2 _padder__U718  ( .A1(padder_out[136]), .A2(_padder__n2505 ), .ZN(
        _padder__n1109 ) );
  NAND2_X2 _padder__U717  ( .A1(padder_out[232]), .A2(_padder__n2544 ), .ZN(
        _padder__n1110 ) );
  NAND2_X2 _padder__U716  ( .A1(_padder__n1109 ), .A2(_padder__n1110 ), .ZN(
        _padder__n1608 ) );
  NAND2_X2 _padder__U715  ( .A1(padder_out[151]), .A2(_padder__n2489 ), .ZN(
        _padder__n1107 ) );
  NAND2_X2 _padder__U714  ( .A1(padder_out[247]), .A2(_padder__n2544 ), .ZN(
        _padder__n1108 ) );
  NAND2_X2 _padder__U713  ( .A1(_padder__n1107 ), .A2(_padder__n1108 ), .ZN(
        _padder__n1609 ) );
  NAND2_X2 _padder__U712  ( .A1(padder_out[150]), .A2(_padder__n2486 ), .ZN(
        _padder__n1105 ) );
  NAND2_X2 _padder__U711  ( .A1(padder_out[246]), .A2(_padder__n2544 ), .ZN(
        _padder__n1106 ) );
  NAND2_X2 _padder__U710  ( .A1(_padder__n1105 ), .A2(_padder__n1106 ), .ZN(
        _padder__n1610 ) );
  NAND2_X2 _padder__U709  ( .A1(padder_out[149]), .A2(_padder__n2496 ), .ZN(
        _padder__n1103 ) );
  NAND2_X2 _padder__U708  ( .A1(padder_out[245]), .A2(_padder__n2544 ), .ZN(
        _padder__n1104 ) );
  NAND2_X2 _padder__U707  ( .A1(_padder__n1103 ), .A2(_padder__n1104 ), .ZN(
        _padder__n1611 ) );
  NAND2_X2 _padder__U706  ( .A1(padder_out[148]), .A2(_padder__n2485 ), .ZN(
        _padder__n1101 ) );
  NAND2_X2 _padder__U705  ( .A1(padder_out[244]), .A2(_padder__n2544 ), .ZN(
        _padder__n1102 ) );
  NAND2_X2 _padder__U704  ( .A1(_padder__n1101 ), .A2(_padder__n1102 ), .ZN(
        _padder__n1612 ) );
  NAND2_X2 _padder__U703  ( .A1(padder_out[147]), .A2(_padder__n2493 ), .ZN(
        _padder__n1099 ) );
  NAND2_X2 _padder__U702  ( .A1(padder_out[243]), .A2(_padder__n2544 ), .ZN(
        _padder__n1100 ) );
  NAND2_X2 _padder__U701  ( .A1(_padder__n1099 ), .A2(_padder__n1100 ), .ZN(
        _padder__n1613 ) );
  NAND2_X2 _padder__U700  ( .A1(padder_out[146]), .A2(_padder__n2502 ), .ZN(
        _padder__n1097 ) );
  NAND2_X2 _padder__U699  ( .A1(padder_out[242]), .A2(_padder__n2544 ), .ZN(
        _padder__n1098 ) );
  NAND2_X2 _padder__U698  ( .A1(_padder__n1097 ), .A2(_padder__n1098 ), .ZN(
        _padder__n1614 ) );
  NAND2_X2 _padder__U697  ( .A1(padder_out[145]), .A2(_padder__n2486 ), .ZN(
        _padder__n1095 ) );
  NAND2_X2 _padder__U696  ( .A1(padder_out[241]), .A2(_padder__n2545 ), .ZN(
        _padder__n1096 ) );
  NAND2_X2 _padder__U695  ( .A1(_padder__n1095 ), .A2(_padder__n1096 ), .ZN(
        _padder__n1615 ) );
  NAND2_X2 _padder__U694  ( .A1(padder_out[144]), .A2(_padder__n2497 ), .ZN(
        _padder__n1093 ) );
  NAND2_X2 _padder__U693  ( .A1(padder_out[240]), .A2(_padder__n2545 ), .ZN(
        _padder__n1094 ) );
  NAND2_X2 _padder__U692  ( .A1(_padder__n1093 ), .A2(_padder__n1094 ), .ZN(
        _padder__n1616 ) );
  NAND2_X2 _padder__U691  ( .A1(padder_out[159]), .A2(_padder__n2500 ), .ZN(
        _padder__n1091 ) );
  NAND2_X2 _padder__U690  ( .A1(padder_out[255]), .A2(_padder__n2545 ), .ZN(
        _padder__n1092 ) );
  NAND2_X2 _padder__U689  ( .A1(_padder__n1091 ), .A2(_padder__n1092 ), .ZN(
        _padder__n1617 ) );
  NAND2_X2 _padder__U688  ( .A1(padder_out[158]), .A2(_padder__n2499 ), .ZN(
        _padder__n1089 ) );
  NAND2_X2 _padder__U687  ( .A1(padder_out[254]), .A2(_padder__n2545 ), .ZN(
        _padder__n1090 ) );
  NAND2_X2 _padder__U686  ( .A1(_padder__n1089 ), .A2(_padder__n1090 ), .ZN(
        _padder__n1618 ) );
  NAND2_X2 _padder__U685  ( .A1(padder_out[157]), .A2(_padder__n2498 ), .ZN(
        _padder__n1087 ) );
  NAND2_X2 _padder__U684  ( .A1(padder_out[253]), .A2(_padder__n2545 ), .ZN(
        _padder__n1088 ) );
  NAND2_X2 _padder__U683  ( .A1(_padder__n1087 ), .A2(_padder__n1088 ), .ZN(
        _padder__n1619 ) );
  NAND2_X2 _padder__U682  ( .A1(padder_out[156]), .A2(_padder__n2483 ), .ZN(
        _padder__n1085 ) );
  NAND2_X2 _padder__U681  ( .A1(padder_out[252]), .A2(_padder__n2545 ), .ZN(
        _padder__n1086 ) );
  NAND2_X2 _padder__U680  ( .A1(_padder__n1085 ), .A2(_padder__n1086 ), .ZN(
        _padder__n1620 ) );
  NAND2_X2 _padder__U679  ( .A1(padder_out[155]), .A2(_padder__n2483 ), .ZN(
        _padder__n1083 ) );
  NAND2_X2 _padder__U678  ( .A1(padder_out[251]), .A2(_padder__n2545 ), .ZN(
        _padder__n1084 ) );
  NAND2_X2 _padder__U677  ( .A1(_padder__n1083 ), .A2(_padder__n1084 ), .ZN(
        _padder__n1621 ) );
  NAND2_X2 _padder__U676  ( .A1(padder_out[154]), .A2(_padder__n2483 ), .ZN(
        _padder__n1081 ) );
  NAND2_X2 _padder__U675  ( .A1(padder_out[250]), .A2(_padder__n2545 ), .ZN(
        _padder__n1082 ) );
  NAND2_X2 _padder__U674  ( .A1(_padder__n1081 ), .A2(_padder__n1082 ), .ZN(
        _padder__n1622 ) );
  NAND2_X2 _padder__U673  ( .A1(padder_out[153]), .A2(_padder__n2483 ), .ZN(
        _padder__n1079 ) );
  NAND2_X2 _padder__U672  ( .A1(padder_out[249]), .A2(_padder__n2545 ), .ZN(
        _padder__n1080 ) );
  NAND2_X2 _padder__U671  ( .A1(_padder__n1079 ), .A2(_padder__n1080 ), .ZN(
        _padder__n1623 ) );
  NAND2_X2 _padder__U670  ( .A1(padder_out[152]), .A2(_padder__n2483 ), .ZN(
        _padder__n1077 ) );
  NAND2_X2 _padder__U669  ( .A1(padder_out[248]), .A2(_padder__n2545 ), .ZN(
        _padder__n1078 ) );
  NAND2_X2 _padder__U668  ( .A1(_padder__n1077 ), .A2(_padder__n1078 ), .ZN(
        _padder__n1624 ) );
  NAND2_X2 _padder__U667  ( .A1(padder_out[167]), .A2(_padder__n2483 ), .ZN(
        _padder__n1075 ) );
  NAND2_X2 _padder__U666  ( .A1(padder_out[135]), .A2(_padder__n2545 ), .ZN(
        _padder__n1076 ) );
  NAND2_X2 _padder__U665  ( .A1(_padder__n1075 ), .A2(_padder__n1076 ), .ZN(
        _padder__n1625 ) );
  NAND2_X2 _padder__U664  ( .A1(padder_out[166]), .A2(_padder__n2483 ), .ZN(
        _padder__n1073 ) );
  NAND2_X2 _padder__U663  ( .A1(padder_out[134]), .A2(_padder__n2546 ), .ZN(
        _padder__n1074 ) );
  NAND2_X2 _padder__U662  ( .A1(_padder__n1073 ), .A2(_padder__n1074 ), .ZN(
        _padder__n1626 ) );
  NAND2_X2 _padder__U661  ( .A1(padder_out[165]), .A2(_padder__n2483 ), .ZN(
        _padder__n1071 ) );
  NAND2_X2 _padder__U660  ( .A1(padder_out[133]), .A2(_padder__n2546 ), .ZN(
        _padder__n1072 ) );
  NAND2_X2 _padder__U659  ( .A1(_padder__n1071 ), .A2(_padder__n1072 ), .ZN(
        _padder__n1627 ) );
  NAND2_X2 _padder__U658  ( .A1(padder_out[164]), .A2(_padder__n2483 ), .ZN(
        _padder__n1069 ) );
  NAND2_X2 _padder__U657  ( .A1(padder_out[132]), .A2(_padder__n2546 ), .ZN(
        _padder__n1070 ) );
  NAND2_X2 _padder__U656  ( .A1(_padder__n1069 ), .A2(_padder__n1070 ), .ZN(
        _padder__n1628 ) );
  NAND2_X2 _padder__U655  ( .A1(padder_out[163]), .A2(_padder__n2483 ), .ZN(
        _padder__n1067 ) );
  NAND2_X2 _padder__U654  ( .A1(padder_out[131]), .A2(_padder__n2546 ), .ZN(
        _padder__n1068 ) );
  NAND2_X2 _padder__U653  ( .A1(_padder__n1067 ), .A2(_padder__n1068 ), .ZN(
        _padder__n1629 ) );
  NAND2_X2 _padder__U652  ( .A1(padder_out[162]), .A2(_padder__n2483 ), .ZN(
        _padder__n1065 ) );
  NAND2_X2 _padder__U651  ( .A1(padder_out[130]), .A2(_padder__n2546 ), .ZN(
        _padder__n1066 ) );
  NAND2_X2 _padder__U650  ( .A1(_padder__n1065 ), .A2(_padder__n1066 ), .ZN(
        _padder__n1630 ) );
  NAND2_X2 _padder__U649  ( .A1(padder_out[161]), .A2(_padder__n2484 ), .ZN(
        _padder__n1063 ) );
  NAND2_X2 _padder__U648  ( .A1(padder_out[129]), .A2(_padder__n2546 ), .ZN(
        _padder__n1064 ) );
  NAND2_X2 _padder__U647  ( .A1(_padder__n1063 ), .A2(_padder__n1064 ), .ZN(
        _padder__n1631 ) );
  NAND2_X2 _padder__U646  ( .A1(padder_out[160]), .A2(_padder__n2484 ), .ZN(
        _padder__n1061 ) );
  NAND2_X2 _padder__U645  ( .A1(padder_out[128]), .A2(_padder__n2546 ), .ZN(
        _padder__n1062 ) );
  NAND2_X2 _padder__U644  ( .A1(_padder__n1061 ), .A2(_padder__n1062 ), .ZN(
        _padder__n1632 ) );
  NAND2_X2 _padder__U643  ( .A1(padder_out[175]), .A2(_padder__n2484 ), .ZN(
        _padder__n1059 ) );
  NAND2_X2 _padder__U642  ( .A1(padder_out[143]), .A2(_padder__n2546 ), .ZN(
        _padder__n1060 ) );
  NAND2_X2 _padder__U641  ( .A1(_padder__n1059 ), .A2(_padder__n1060 ), .ZN(
        _padder__n1633 ) );
  NAND2_X2 _padder__U640  ( .A1(padder_out[174]), .A2(_padder__n2484 ), .ZN(
        _padder__n1057 ) );
  NAND2_X2 _padder__U639  ( .A1(padder_out[142]), .A2(_padder__n2546 ), .ZN(
        _padder__n1058 ) );
  NAND2_X2 _padder__U638  ( .A1(_padder__n1057 ), .A2(_padder__n1058 ), .ZN(
        _padder__n1634 ) );
  NAND2_X2 _padder__U637  ( .A1(padder_out[173]), .A2(_padder__n2484 ), .ZN(
        _padder__n1055 ) );
  NAND2_X2 _padder__U636  ( .A1(padder_out[141]), .A2(_padder__n2546 ), .ZN(
        _padder__n1056 ) );
  NAND2_X2 _padder__U635  ( .A1(_padder__n1055 ), .A2(_padder__n1056 ), .ZN(
        _padder__n1635 ) );
  NAND2_X2 _padder__U634  ( .A1(padder_out[172]), .A2(_padder__n2484 ), .ZN(
        _padder__n1053 ) );
  NAND2_X2 _padder__U633  ( .A1(padder_out[140]), .A2(_padder__n2546 ), .ZN(
        _padder__n1054 ) );
  NAND2_X2 _padder__U632  ( .A1(_padder__n1053 ), .A2(_padder__n1054 ), .ZN(
        _padder__n1636 ) );
  NAND2_X2 _padder__U631  ( .A1(padder_out[171]), .A2(_padder__n2484 ), .ZN(
        _padder__n1051 ) );
  NAND2_X2 _padder__U630  ( .A1(padder_out[139]), .A2(_padder__n2547 ), .ZN(
        _padder__n1052 ) );
  NAND2_X2 _padder__U629  ( .A1(_padder__n1051 ), .A2(_padder__n1052 ), .ZN(
        _padder__n1637 ) );
  NAND2_X2 _padder__U628  ( .A1(padder_out[170]), .A2(_padder__n2484 ), .ZN(
        _padder__n1049 ) );
  NAND2_X2 _padder__U627  ( .A1(padder_out[138]), .A2(_padder__n2547 ), .ZN(
        _padder__n1050 ) );
  NAND2_X2 _padder__U626  ( .A1(_padder__n1049 ), .A2(_padder__n1050 ), .ZN(
        _padder__n1638 ) );
  NAND2_X2 _padder__U625  ( .A1(padder_out[169]), .A2(_padder__n2484 ), .ZN(
        _padder__n1047 ) );
  NAND2_X2 _padder__U624  ( .A1(padder_out[137]), .A2(_padder__n2547 ), .ZN(
        _padder__n1048 ) );
  NAND2_X2 _padder__U623  ( .A1(_padder__n1047 ), .A2(_padder__n1048 ), .ZN(
        _padder__n1639 ) );
  NAND2_X2 _padder__U622  ( .A1(padder_out[168]), .A2(_padder__n2484 ), .ZN(
        _padder__n1045 ) );
  NAND2_X2 _padder__U621  ( .A1(padder_out[136]), .A2(_padder__n2547 ), .ZN(
        _padder__n1046 ) );
  NAND2_X2 _padder__U620  ( .A1(_padder__n1045 ), .A2(_padder__n1046 ), .ZN(
        _padder__n1640 ) );
  NAND2_X2 _padder__U619  ( .A1(padder_out[183]), .A2(_padder__n2484 ), .ZN(
        _padder__n1043 ) );
  NAND2_X2 _padder__U618  ( .A1(padder_out[151]), .A2(_padder__n2547 ), .ZN(
        _padder__n1044 ) );
  NAND2_X2 _padder__U617  ( .A1(_padder__n1043 ), .A2(_padder__n1044 ), .ZN(
        _padder__n1641 ) );
  NAND2_X2 _padder__U616  ( .A1(padder_out[182]), .A2(_padder__n2484 ), .ZN(
        _padder__n1041 ) );
  NAND2_X2 _padder__U615  ( .A1(padder_out[150]), .A2(_padder__n2547 ), .ZN(
        _padder__n1042 ) );
  NAND2_X2 _padder__U614  ( .A1(_padder__n1041 ), .A2(_padder__n1042 ), .ZN(
        _padder__n1642 ) );
  NAND2_X2 _padder__U613  ( .A1(padder_out[181]), .A2(_padder__n2484 ), .ZN(
        _padder__n1039 ) );
  NAND2_X2 _padder__U612  ( .A1(padder_out[149]), .A2(_padder__n2547 ), .ZN(
        _padder__n1040 ) );
  NAND2_X2 _padder__U611  ( .A1(_padder__n1039 ), .A2(_padder__n1040 ), .ZN(
        _padder__n1643 ) );
  NAND2_X2 _padder__U610  ( .A1(padder_out[180]), .A2(_padder__n2484 ), .ZN(
        _padder__n1037 ) );
  NAND2_X2 _padder__U609  ( .A1(padder_out[148]), .A2(_padder__n2547 ), .ZN(
        _padder__n1038 ) );
  NAND2_X2 _padder__U608  ( .A1(_padder__n1037 ), .A2(_padder__n1038 ), .ZN(
        _padder__n1644 ) );
  NAND2_X2 _padder__U607  ( .A1(padder_out[179]), .A2(_padder__n2484 ), .ZN(
        _padder__n1035 ) );
  NAND2_X2 _padder__U606  ( .A1(padder_out[147]), .A2(_padder__n2547 ), .ZN(
        _padder__n1036 ) );
  NAND2_X2 _padder__U605  ( .A1(_padder__n1035 ), .A2(_padder__n1036 ), .ZN(
        _padder__n1645 ) );
  NAND2_X2 _padder__U604  ( .A1(padder_out[178]), .A2(_padder__n2484 ), .ZN(
        _padder__n1033 ) );
  NAND2_X2 _padder__U603  ( .A1(padder_out[146]), .A2(_padder__n2547 ), .ZN(
        _padder__n1034 ) );
  NAND2_X2 _padder__U602  ( .A1(_padder__n1033 ), .A2(_padder__n1034 ), .ZN(
        _padder__n1646 ) );
  NAND2_X2 _padder__U601  ( .A1(padder_out[177]), .A2(_padder__n2484 ), .ZN(
        _padder__n1031 ) );
  NAND2_X2 _padder__U600  ( .A1(padder_out[145]), .A2(_padder__n2547 ), .ZN(
        _padder__n1032 ) );
  NAND2_X2 _padder__U599  ( .A1(_padder__n1031 ), .A2(_padder__n1032 ), .ZN(
        _padder__n1647 ) );
  NAND2_X2 _padder__U598  ( .A1(padder_out[176]), .A2(_padder__n2484 ), .ZN(
        _padder__n1029 ) );
  NAND2_X2 _padder__U597  ( .A1(padder_out[144]), .A2(_padder__n2548 ), .ZN(
        _padder__n1030 ) );
  NAND2_X2 _padder__U596  ( .A1(_padder__n1029 ), .A2(_padder__n1030 ), .ZN(
        _padder__n1648 ) );
  NAND2_X2 _padder__U595  ( .A1(padder_out[191]), .A2(_padder__n2494 ), .ZN(
        _padder__n1027 ) );
  NAND2_X2 _padder__U594  ( .A1(padder_out[159]), .A2(_padder__n2548 ), .ZN(
        _padder__n1028 ) );
  NAND2_X2 _padder__U593  ( .A1(_padder__n1027 ), .A2(_padder__n1028 ), .ZN(
        _padder__n1649 ) );
  NAND2_X2 _padder__U592  ( .A1(padder_out[190]), .A2(_padder__n2494 ), .ZN(
        _padder__n1025 ) );
  NAND2_X2 _padder__U591  ( .A1(padder_out[158]), .A2(_padder__n2548 ), .ZN(
        _padder__n1026 ) );
  NAND2_X2 _padder__U590  ( .A1(_padder__n1025 ), .A2(_padder__n1026 ), .ZN(
        _padder__n1650 ) );
  NAND2_X2 _padder__U589  ( .A1(padder_out[189]), .A2(_padder__n2494 ), .ZN(
        _padder__n1023 ) );
  NAND2_X2 _padder__U588  ( .A1(padder_out[157]), .A2(_padder__n2548 ), .ZN(
        _padder__n1024 ) );
  NAND2_X2 _padder__U587  ( .A1(_padder__n1023 ), .A2(_padder__n1024 ), .ZN(
        _padder__n1651 ) );
  NAND2_X2 _padder__U586  ( .A1(padder_out[188]), .A2(_padder__n2494 ), .ZN(
        _padder__n1021 ) );
  NAND2_X2 _padder__U585  ( .A1(padder_out[156]), .A2(_padder__n2548 ), .ZN(
        _padder__n1022 ) );
  NAND2_X2 _padder__U584  ( .A1(_padder__n1021 ), .A2(_padder__n1022 ), .ZN(
        _padder__n1652 ) );
  NAND2_X2 _padder__U583  ( .A1(padder_out[187]), .A2(_padder__n2494 ), .ZN(
        _padder__n1019 ) );
  NAND2_X2 _padder__U582  ( .A1(padder_out[155]), .A2(_padder__n2548 ), .ZN(
        _padder__n1020 ) );
  NAND2_X2 _padder__U581  ( .A1(_padder__n1019 ), .A2(_padder__n1020 ), .ZN(
        _padder__n1653 ) );
  NAND2_X2 _padder__U580  ( .A1(padder_out[186]), .A2(_padder__n2494 ), .ZN(
        _padder__n1017 ) );
  NAND2_X2 _padder__U579  ( .A1(padder_out[154]), .A2(_padder__n2548 ), .ZN(
        _padder__n1018 ) );
  NAND2_X2 _padder__U578  ( .A1(_padder__n1017 ), .A2(_padder__n1018 ), .ZN(
        _padder__n1654 ) );
  NAND2_X2 _padder__U577  ( .A1(padder_out[185]), .A2(_padder__n2494 ), .ZN(
        _padder__n1015 ) );
  NAND2_X2 _padder__U576  ( .A1(padder_out[153]), .A2(_padder__n2548 ), .ZN(
        _padder__n1016 ) );
  NAND2_X2 _padder__U575  ( .A1(_padder__n1015 ), .A2(_padder__n1016 ), .ZN(
        _padder__n1655 ) );
  NAND2_X2 _padder__U574  ( .A1(padder_out[184]), .A2(_padder__n2494 ), .ZN(
        _padder__n1013 ) );
  NAND2_X2 _padder__U573  ( .A1(padder_out[152]), .A2(_padder__n2548 ), .ZN(
        _padder__n1014 ) );
  NAND2_X2 _padder__U572  ( .A1(_padder__n1013 ), .A2(_padder__n1014 ), .ZN(
        _padder__n1656 ) );
  NAND2_X2 _padder__U571  ( .A1(padder_out[71]), .A2(_padder__n2494 ), .ZN(
        _padder__n1011 ) );
  NAND2_X2 _padder__U570  ( .A1(padder_out[167]), .A2(_padder__n2548 ), .ZN(
        _padder__n1012 ) );
  NAND2_X2 _padder__U569  ( .A1(_padder__n1011 ), .A2(_padder__n1012 ), .ZN(
        _padder__n1657 ) );
  NAND2_X2 _padder__U568  ( .A1(padder_out[70]), .A2(_padder__n2494 ), .ZN(
        _padder__n1009 ) );
  NAND2_X2 _padder__U567  ( .A1(padder_out[166]), .A2(_padder__n2548 ), .ZN(
        _padder__n1010 ) );
  NAND2_X2 _padder__U566  ( .A1(_padder__n1009 ), .A2(_padder__n1010 ), .ZN(
        _padder__n1658 ) );
  NAND2_X2 _padder__U565  ( .A1(padder_out[69]), .A2(_padder__n2494 ), .ZN(
        _padder__n1007 ) );
  NAND2_X2 _padder__U564  ( .A1(padder_out[165]), .A2(_padder__n2549 ), .ZN(
        _padder__n1008 ) );
  NAND2_X2 _padder__U563  ( .A1(_padder__n1007 ), .A2(_padder__n1008 ), .ZN(
        _padder__n1659 ) );
  NAND2_X2 _padder__U562  ( .A1(padder_out[68]), .A2(_padder__n2494 ), .ZN(
        _padder__n1005 ) );
  NAND2_X2 _padder__U561  ( .A1(padder_out[164]), .A2(_padder__n2549 ), .ZN(
        _padder__n1006 ) );
  NAND2_X2 _padder__U560  ( .A1(_padder__n1005 ), .A2(_padder__n1006 ), .ZN(
        _padder__n1660 ) );
  NAND2_X2 _padder__U559  ( .A1(padder_out[67]), .A2(_padder__n2494 ), .ZN(
        _padder__n1003 ) );
  NAND2_X2 _padder__U558  ( .A1(padder_out[163]), .A2(_padder__n2549 ), .ZN(
        _padder__n1004 ) );
  NAND2_X2 _padder__U557  ( .A1(_padder__n1003 ), .A2(_padder__n1004 ), .ZN(
        _padder__n1661 ) );
  NAND2_X2 _padder__U556  ( .A1(padder_out[66]), .A2(_padder__n2493 ), .ZN(
        _padder__n1001 ) );
  NAND2_X2 _padder__U555  ( .A1(padder_out[162]), .A2(_padder__n2549 ), .ZN(
        _padder__n1002 ) );
  NAND2_X2 _padder__U554  ( .A1(_padder__n1001 ), .A2(_padder__n1002 ), .ZN(
        _padder__n1662 ) );
  NAND2_X2 _padder__U553  ( .A1(padder_out[65]), .A2(_padder__n2493 ), .ZN(
        _padder__n999 ) );
  NAND2_X2 _padder__U552  ( .A1(padder_out[161]), .A2(_padder__n2549 ), .ZN(
        _padder__n1000 ) );
  NAND2_X2 _padder__U551  ( .A1(_padder__n999 ), .A2(_padder__n1000 ), .ZN(
        _padder__n1663 ) );
  NAND2_X2 _padder__U550  ( .A1(padder_out[64]), .A2(_padder__n2493 ), .ZN(
        _padder__n997 ) );
  NAND2_X2 _padder__U549  ( .A1(padder_out[160]), .A2(_padder__n2549 ), .ZN(
        _padder__n998 ) );
  NAND2_X2 _padder__U548  ( .A1(_padder__n997 ), .A2(_padder__n998 ), .ZN(
        _padder__n1664 ) );
  NAND2_X2 _padder__U547  ( .A1(padder_out[79]), .A2(_padder__n2493 ), .ZN(
        _padder__n995 ) );
  NAND2_X2 _padder__U546  ( .A1(padder_out[175]), .A2(_padder__n2549 ), .ZN(
        _padder__n996 ) );
  NAND2_X2 _padder__U545  ( .A1(_padder__n995 ), .A2(_padder__n996 ), .ZN(
        _padder__n1665 ) );
  NAND2_X2 _padder__U544  ( .A1(padder_out[78]), .A2(_padder__n2493 ), .ZN(
        _padder__n993 ) );
  NAND2_X2 _padder__U543  ( .A1(padder_out[174]), .A2(_padder__n2549 ), .ZN(
        _padder__n994 ) );
  NAND2_X2 _padder__U542  ( .A1(_padder__n993 ), .A2(_padder__n994 ), .ZN(
        _padder__n1666 ) );
  NAND2_X2 _padder__U541  ( .A1(padder_out[77]), .A2(_padder__n2493 ), .ZN(
        _padder__n991 ) );
  NAND2_X2 _padder__U540  ( .A1(padder_out[173]), .A2(_padder__n2549 ), .ZN(
        _padder__n992 ) );
  NAND2_X2 _padder__U539  ( .A1(_padder__n991 ), .A2(_padder__n992 ), .ZN(
        _padder__n1667 ) );
  NAND2_X2 _padder__U538  ( .A1(padder_out[76]), .A2(_padder__n2493 ), .ZN(
        _padder__n989 ) );
  NAND2_X2 _padder__U537  ( .A1(padder_out[172]), .A2(_padder__n2549 ), .ZN(
        _padder__n990 ) );
  NAND2_X2 _padder__U536  ( .A1(_padder__n989 ), .A2(_padder__n990 ), .ZN(
        _padder__n1668 ) );
  NAND2_X2 _padder__U535  ( .A1(padder_out[75]), .A2(_padder__n2493 ), .ZN(
        _padder__n987 ) );
  NAND2_X2 _padder__U534  ( .A1(padder_out[171]), .A2(_padder__n2549 ), .ZN(
        _padder__n988 ) );
  NAND2_X2 _padder__U533  ( .A1(_padder__n987 ), .A2(_padder__n988 ), .ZN(
        _padder__n1669 ) );
  NAND2_X2 _padder__U532  ( .A1(padder_out[74]), .A2(_padder__n2493 ), .ZN(
        _padder__n985 ) );
  NAND2_X2 _padder__U531  ( .A1(padder_out[170]), .A2(_padder__n2550 ), .ZN(
        _padder__n986 ) );
  NAND2_X2 _padder__U530  ( .A1(_padder__n985 ), .A2(_padder__n986 ), .ZN(
        _padder__n1670 ) );
  NAND2_X2 _padder__U529  ( .A1(padder_out[73]), .A2(_padder__n2493 ), .ZN(
        _padder__n983 ) );
  NAND2_X2 _padder__U528  ( .A1(padder_out[169]), .A2(_padder__n2550 ), .ZN(
        _padder__n984 ) );
  NAND2_X2 _padder__U527  ( .A1(_padder__n983 ), .A2(_padder__n984 ), .ZN(
        _padder__n1671 ) );
  NAND2_X2 _padder__U526  ( .A1(padder_out[72]), .A2(_padder__n2493 ), .ZN(
        _padder__n981 ) );
  NAND2_X2 _padder__U525  ( .A1(padder_out[168]), .A2(_padder__n2550 ), .ZN(
        _padder__n982 ) );
  NAND2_X2 _padder__U524  ( .A1(_padder__n981 ), .A2(_padder__n982 ), .ZN(
        _padder__n1672 ) );
  NAND2_X2 _padder__U523  ( .A1(padder_out[87]), .A2(_padder__n2493 ), .ZN(
        _padder__n979 ) );
  NAND2_X2 _padder__U522  ( .A1(padder_out[183]), .A2(_padder__n2550 ), .ZN(
        _padder__n980 ) );
  NAND2_X2 _padder__U521  ( .A1(_padder__n979 ), .A2(_padder__n980 ), .ZN(
        _padder__n1673 ) );
  NAND2_X2 _padder__U520  ( .A1(padder_out[86]), .A2(_padder__n2493 ), .ZN(
        _padder__n977 ) );
  NAND2_X2 _padder__U519  ( .A1(padder_out[182]), .A2(_padder__n2550 ), .ZN(
        _padder__n978 ) );
  NAND2_X2 _padder__U518  ( .A1(_padder__n977 ), .A2(_padder__n978 ), .ZN(
        _padder__n1674 ) );
  NAND2_X2 _padder__U517  ( .A1(padder_out[85]), .A2(_padder__n2493 ), .ZN(
        _padder__n975 ) );
  NAND2_X2 _padder__U516  ( .A1(padder_out[181]), .A2(_padder__n2550 ), .ZN(
        _padder__n976 ) );
  NAND2_X2 _padder__U515  ( .A1(_padder__n975 ), .A2(_padder__n976 ), .ZN(
        _padder__n1675 ) );
  NAND2_X2 _padder__U514  ( .A1(padder_out[84]), .A2(_padder__n2493 ), .ZN(
        _padder__n973 ) );
  NAND2_X2 _padder__U513  ( .A1(padder_out[180]), .A2(_padder__n2550 ), .ZN(
        _padder__n974 ) );
  NAND2_X2 _padder__U512  ( .A1(_padder__n973 ), .A2(_padder__n974 ), .ZN(
        _padder__n1676 ) );
  NAND2_X2 _padder__U511  ( .A1(padder_out[83]), .A2(_padder__n2493 ), .ZN(
        _padder__n971 ) );
  NAND2_X2 _padder__U510  ( .A1(padder_out[179]), .A2(_padder__n2550 ), .ZN(
        _padder__n972 ) );
  NAND2_X2 _padder__U509  ( .A1(_padder__n971 ), .A2(_padder__n972 ), .ZN(
        _padder__n1677 ) );
  NAND2_X2 _padder__U508  ( .A1(padder_out[82]), .A2(_padder__n2493 ), .ZN(
        _padder__n969 ) );
  NAND2_X2 _padder__U507  ( .A1(padder_out[178]), .A2(_padder__n2550 ), .ZN(
        _padder__n970 ) );
  NAND2_X2 _padder__U506  ( .A1(_padder__n969 ), .A2(_padder__n970 ), .ZN(
        _padder__n1678 ) );
  NAND2_X2 _padder__U505  ( .A1(padder_out[81]), .A2(_padder__n2493 ), .ZN(
        _padder__n967 ) );
  NAND2_X2 _padder__U504  ( .A1(padder_out[177]), .A2(_padder__n2550 ), .ZN(
        _padder__n968 ) );
  NAND2_X2 _padder__U503  ( .A1(_padder__n967 ), .A2(_padder__n968 ), .ZN(
        _padder__n1679 ) );
  NAND2_X2 _padder__U502  ( .A1(padder_out[80]), .A2(_padder__n2493 ), .ZN(
        _padder__n965 ) );
  NAND2_X2 _padder__U501  ( .A1(padder_out[176]), .A2(_padder__n2550 ), .ZN(
        _padder__n966 ) );
  NAND2_X2 _padder__U500  ( .A1(_padder__n965 ), .A2(_padder__n966 ), .ZN(
        _padder__n1680 ) );
  NAND2_X2 _padder__U499  ( .A1(padder_out[95]), .A2(_padder__n2493 ), .ZN(
        _padder__n963 ) );
  NAND2_X2 _padder__U498  ( .A1(padder_out[191]), .A2(_padder__n2551 ), .ZN(
        _padder__n964 ) );
  NAND2_X2 _padder__U497  ( .A1(_padder__n963 ), .A2(_padder__n964 ), .ZN(
        _padder__n1681 ) );
  NAND2_X2 _padder__U496  ( .A1(padder_out[94]), .A2(_padder__n2493 ), .ZN(
        _padder__n961 ) );
  NAND2_X2 _padder__U495  ( .A1(padder_out[190]), .A2(_padder__n2551 ), .ZN(
        _padder__n962 ) );
  NAND2_X2 _padder__U494  ( .A1(_padder__n961 ), .A2(_padder__n962 ), .ZN(
        _padder__n1682 ) );
  NAND2_X2 _padder__U493  ( .A1(padder_out[93]), .A2(_padder__n2493 ), .ZN(
        _padder__n959 ) );
  NAND2_X2 _padder__U492  ( .A1(padder_out[189]), .A2(_padder__n2551 ), .ZN(
        _padder__n960 ) );
  NAND2_X2 _padder__U491  ( .A1(_padder__n959 ), .A2(_padder__n960 ), .ZN(
        _padder__n1683 ) );
  NAND2_X2 _padder__U490  ( .A1(padder_out[92]), .A2(_padder__n2493 ), .ZN(
        _padder__n957 ) );
  NAND2_X2 _padder__U489  ( .A1(padder_out[188]), .A2(_padder__n2551 ), .ZN(
        _padder__n958 ) );
  NAND2_X2 _padder__U488  ( .A1(_padder__n957 ), .A2(_padder__n958 ), .ZN(
        _padder__n1684 ) );
  NAND2_X2 _padder__U487  ( .A1(padder_out[91]), .A2(_padder__n2493 ), .ZN(
        _padder__n955 ) );
  NAND2_X2 _padder__U486  ( .A1(padder_out[187]), .A2(_padder__n2551 ), .ZN(
        _padder__n956 ) );
  NAND2_X2 _padder__U485  ( .A1(_padder__n955 ), .A2(_padder__n956 ), .ZN(
        _padder__n1685 ) );
  NAND2_X2 _padder__U484  ( .A1(padder_out[90]), .A2(_padder__n2492 ), .ZN(
        _padder__n953 ) );
  NAND2_X2 _padder__U483  ( .A1(padder_out[186]), .A2(_padder__n2551 ), .ZN(
        _padder__n954 ) );
  NAND2_X2 _padder__U482  ( .A1(_padder__n953 ), .A2(_padder__n954 ), .ZN(
        _padder__n1686 ) );
  NAND2_X2 _padder__U481  ( .A1(padder_out[89]), .A2(_padder__n2492 ), .ZN(
        _padder__n951 ) );
  NAND2_X2 _padder__U480  ( .A1(padder_out[185]), .A2(_padder__n2551 ), .ZN(
        _padder__n952 ) );
  NAND2_X2 _padder__U479  ( .A1(_padder__n951 ), .A2(_padder__n952 ), .ZN(
        _padder__n1687 ) );
  NAND2_X2 _padder__U478  ( .A1(padder_out[88]), .A2(_padder__n2492 ), .ZN(
        _padder__n949 ) );
  NAND2_X2 _padder__U477  ( .A1(padder_out[184]), .A2(_padder__n2551 ), .ZN(
        _padder__n950 ) );
  NAND2_X2 _padder__U476  ( .A1(_padder__n949 ), .A2(_padder__n950 ), .ZN(
        _padder__n1688 ) );
  NAND2_X2 _padder__U475  ( .A1(padder_out[103]), .A2(_padder__n2492 ), .ZN(
        _padder__n947 ) );
  NAND2_X2 _padder__U474  ( .A1(padder_out[71]), .A2(_padder__n2551 ), .ZN(
        _padder__n948 ) );
  NAND2_X2 _padder__U473  ( .A1(_padder__n947 ), .A2(_padder__n948 ), .ZN(
        _padder__n1689 ) );
  NAND2_X2 _padder__U472  ( .A1(padder_out[102]), .A2(_padder__n2492 ), .ZN(
        _padder__n945 ) );
  NAND2_X2 _padder__U471  ( .A1(padder_out[70]), .A2(_padder__n2551 ), .ZN(
        _padder__n946 ) );
  NAND2_X2 _padder__U470  ( .A1(_padder__n945 ), .A2(_padder__n946 ), .ZN(
        _padder__n1690 ) );
  NAND2_X2 _padder__U469  ( .A1(padder_out[101]), .A2(_padder__n2492 ), .ZN(
        _padder__n943 ) );
  NAND2_X2 _padder__U468  ( .A1(padder_out[69]), .A2(_padder__n2551 ), .ZN(
        _padder__n944 ) );
  NAND2_X2 _padder__U467  ( .A1(_padder__n943 ), .A2(_padder__n944 ), .ZN(
        _padder__n1691 ) );
  NAND2_X2 _padder__U466  ( .A1(padder_out[100]), .A2(_padder__n2492 ), .ZN(
        _padder__n941 ) );
  NAND2_X2 _padder__U465  ( .A1(padder_out[68]), .A2(_padder__n2552 ), .ZN(
        _padder__n942 ) );
  NAND2_X2 _padder__U464  ( .A1(_padder__n941 ), .A2(_padder__n942 ), .ZN(
        _padder__n1692 ) );
  NAND2_X2 _padder__U463  ( .A1(padder_out[99]), .A2(_padder__n2492 ), .ZN(
        _padder__n939 ) );
  NAND2_X2 _padder__U462  ( .A1(padder_out[67]), .A2(_padder__n2552 ), .ZN(
        _padder__n940 ) );
  NAND2_X2 _padder__U461  ( .A1(_padder__n939 ), .A2(_padder__n940 ), .ZN(
        _padder__n1693 ) );
  NAND2_X2 _padder__U460  ( .A1(padder_out[98]), .A2(_padder__n2492 ), .ZN(
        _padder__n937 ) );
  NAND2_X2 _padder__U459  ( .A1(padder_out[66]), .A2(_padder__n2552 ), .ZN(
        _padder__n938 ) );
  NAND2_X2 _padder__U458  ( .A1(_padder__n937 ), .A2(_padder__n938 ), .ZN(
        _padder__n1694 ) );
  NAND2_X2 _padder__U457  ( .A1(padder_out[97]), .A2(_padder__n2492 ), .ZN(
        _padder__n935 ) );
  NAND2_X2 _padder__U456  ( .A1(padder_out[65]), .A2(_padder__n2552 ), .ZN(
        _padder__n936 ) );
  NAND2_X2 _padder__U455  ( .A1(_padder__n935 ), .A2(_padder__n936 ), .ZN(
        _padder__n1695 ) );
  NAND2_X2 _padder__U454  ( .A1(padder_out[96]), .A2(_padder__n2492 ), .ZN(
        _padder__n933 ) );
  NAND2_X2 _padder__U453  ( .A1(padder_out[64]), .A2(_padder__n2552 ), .ZN(
        _padder__n934 ) );
  NAND2_X2 _padder__U452  ( .A1(_padder__n933 ), .A2(_padder__n934 ), .ZN(
        _padder__n1696 ) );
  NAND2_X2 _padder__U451  ( .A1(padder_out[111]), .A2(_padder__n2492 ), .ZN(
        _padder__n931 ) );
  NAND2_X2 _padder__U450  ( .A1(padder_out[79]), .A2(_padder__n2552 ), .ZN(
        _padder__n932 ) );
  NAND2_X2 _padder__U449  ( .A1(_padder__n931 ), .A2(_padder__n932 ), .ZN(
        _padder__n1697 ) );
  NAND2_X2 _padder__U448  ( .A1(padder_out[110]), .A2(_padder__n2492 ), .ZN(
        _padder__n929 ) );
  NAND2_X2 _padder__U447  ( .A1(padder_out[78]), .A2(_padder__n2552 ), .ZN(
        _padder__n930 ) );
  NAND2_X2 _padder__U446  ( .A1(_padder__n929 ), .A2(_padder__n930 ), .ZN(
        _padder__n1698 ) );
  NAND2_X2 _padder__U445  ( .A1(padder_out[109]), .A2(_padder__n2492 ), .ZN(
        _padder__n927 ) );
  NAND2_X2 _padder__U444  ( .A1(padder_out[77]), .A2(_padder__n2552 ), .ZN(
        _padder__n928 ) );
  NAND2_X2 _padder__U443  ( .A1(_padder__n927 ), .A2(_padder__n928 ), .ZN(
        _padder__n1699 ) );
  NAND2_X2 _padder__U442  ( .A1(padder_out[108]), .A2(_padder__n2492 ), .ZN(
        _padder__n925 ) );
  NAND2_X2 _padder__U441  ( .A1(padder_out[76]), .A2(_padder__n2552 ), .ZN(
        _padder__n926 ) );
  NAND2_X2 _padder__U440  ( .A1(_padder__n925 ), .A2(_padder__n926 ), .ZN(
        _padder__n1700 ) );
  NAND2_X2 _padder__U439  ( .A1(padder_out[107]), .A2(_padder__n2492 ), .ZN(
        _padder__n923 ) );
  NAND2_X2 _padder__U438  ( .A1(padder_out[75]), .A2(_padder__n2552 ), .ZN(
        _padder__n924 ) );
  NAND2_X2 _padder__U437  ( .A1(_padder__n923 ), .A2(_padder__n924 ), .ZN(
        _padder__n1701 ) );
  NAND2_X2 _padder__U436  ( .A1(padder_out[106]), .A2(_padder__n2492 ), .ZN(
        _padder__n921 ) );
  NAND2_X2 _padder__U435  ( .A1(padder_out[74]), .A2(_padder__n2552 ), .ZN(
        _padder__n922 ) );
  NAND2_X2 _padder__U434  ( .A1(_padder__n921 ), .A2(_padder__n922 ), .ZN(
        _padder__n1702 ) );
  NAND2_X2 _padder__U433  ( .A1(padder_out[105]), .A2(_padder__n2492 ), .ZN(
        _padder__n919 ) );
  NAND2_X2 _padder__U432  ( .A1(padder_out[73]), .A2(_padder__n2553 ), .ZN(
        _padder__n920 ) );
  NAND2_X2 _padder__U431  ( .A1(_padder__n919 ), .A2(_padder__n920 ), .ZN(
        _padder__n1703 ) );
  NAND2_X2 _padder__U430  ( .A1(padder_out[104]), .A2(_padder__n2492 ), .ZN(
        _padder__n917 ) );
  NAND2_X2 _padder__U429  ( .A1(padder_out[72]), .A2(_padder__n2553 ), .ZN(
        _padder__n918 ) );
  NAND2_X2 _padder__U428  ( .A1(_padder__n917 ), .A2(_padder__n918 ), .ZN(
        _padder__n1704 ) );
  NAND2_X2 _padder__U427  ( .A1(padder_out[119]), .A2(_padder__n2492 ), .ZN(
        _padder__n915 ) );
  NAND2_X2 _padder__U426  ( .A1(padder_out[87]), .A2(_padder__n2553 ), .ZN(
        _padder__n916 ) );
  NAND2_X2 _padder__U425  ( .A1(_padder__n915 ), .A2(_padder__n916 ), .ZN(
        _padder__n1705 ) );
  NAND2_X2 _padder__U424  ( .A1(padder_out[118]), .A2(_padder__n2492 ), .ZN(
        _padder__n913 ) );
  NAND2_X2 _padder__U423  ( .A1(padder_out[86]), .A2(_padder__n2553 ), .ZN(
        _padder__n914 ) );
  NAND2_X2 _padder__U422  ( .A1(_padder__n913 ), .A2(_padder__n914 ), .ZN(
        _padder__n1706 ) );
  NAND2_X2 _padder__U421  ( .A1(padder_out[117]), .A2(_padder__n2492 ), .ZN(
        _padder__n911 ) );
  NAND2_X2 _padder__U420  ( .A1(padder_out[85]), .A2(_padder__n2553 ), .ZN(
        _padder__n912 ) );
  NAND2_X2 _padder__U419  ( .A1(_padder__n911 ), .A2(_padder__n912 ), .ZN(
        _padder__n1707 ) );
  NAND2_X2 _padder__U418  ( .A1(padder_out[116]), .A2(_padder__n2492 ), .ZN(
        _padder__n909 ) );
  NAND2_X2 _padder__U417  ( .A1(padder_out[84]), .A2(_padder__n2553 ), .ZN(
        _padder__n910 ) );
  NAND2_X2 _padder__U416  ( .A1(_padder__n909 ), .A2(_padder__n910 ), .ZN(
        _padder__n1708 ) );
  NAND2_X2 _padder__U415  ( .A1(padder_out[115]), .A2(_padder__n2492 ), .ZN(
        _padder__n907 ) );
  NAND2_X2 _padder__U414  ( .A1(padder_out[83]), .A2(_padder__n2553 ), .ZN(
        _padder__n908 ) );
  NAND2_X2 _padder__U413  ( .A1(_padder__n907 ), .A2(_padder__n908 ), .ZN(
        _padder__n1709 ) );
  NAND2_X2 _padder__U412  ( .A1(padder_out[114]), .A2(_padder__n2491 ), .ZN(
        _padder__n905 ) );
  NAND2_X2 _padder__U411  ( .A1(padder_out[82]), .A2(_padder__n2553 ), .ZN(
        _padder__n906 ) );
  NAND2_X2 _padder__U410  ( .A1(_padder__n905 ), .A2(_padder__n906 ), .ZN(
        _padder__n1710 ) );
  NAND2_X2 _padder__U409  ( .A1(padder_out[113]), .A2(_padder__n2491 ), .ZN(
        _padder__n903 ) );
  NAND2_X2 _padder__U408  ( .A1(padder_out[81]), .A2(_padder__n2553 ), .ZN(
        _padder__n904 ) );
  NAND2_X2 _padder__U407  ( .A1(_padder__n903 ), .A2(_padder__n904 ), .ZN(
        _padder__n1711 ) );
  NAND2_X2 _padder__U406  ( .A1(padder_out[112]), .A2(_padder__n2491 ), .ZN(
        _padder__n901 ) );
  NAND2_X2 _padder__U405  ( .A1(padder_out[80]), .A2(_padder__n2553 ), .ZN(
        _padder__n902 ) );
  NAND2_X2 _padder__U404  ( .A1(_padder__n901 ), .A2(_padder__n902 ), .ZN(
        _padder__n1712 ) );
  NAND2_X2 _padder__U403  ( .A1(padder_out[127]), .A2(_padder__n2491 ), .ZN(
        _padder__n899 ) );
  NAND2_X2 _padder__U402  ( .A1(padder_out[95]), .A2(_padder__n2553 ), .ZN(
        _padder__n900 ) );
  NAND2_X2 _padder__U401  ( .A1(_padder__n899 ), .A2(_padder__n900 ), .ZN(
        _padder__n1713 ) );
  NAND2_X2 _padder__U400  ( .A1(padder_out[126]), .A2(_padder__n2491 ), .ZN(
        _padder__n897 ) );
  NAND2_X2 _padder__U399  ( .A1(padder_out[94]), .A2(_padder__n2554 ), .ZN(
        _padder__n898 ) );
  NAND2_X2 _padder__U398  ( .A1(_padder__n897 ), .A2(_padder__n898 ), .ZN(
        _padder__n1714 ) );
  NAND2_X2 _padder__U397  ( .A1(padder_out[125]), .A2(_padder__n2491 ), .ZN(
        _padder__n895 ) );
  NAND2_X2 _padder__U396  ( .A1(padder_out[93]), .A2(_padder__n2554 ), .ZN(
        _padder__n896 ) );
  NAND2_X2 _padder__U395  ( .A1(_padder__n895 ), .A2(_padder__n896 ), .ZN(
        _padder__n1715 ) );
  NAND2_X2 _padder__U394  ( .A1(padder_out[124]), .A2(_padder__n2491 ), .ZN(
        _padder__n893 ) );
  NAND2_X2 _padder__U393  ( .A1(padder_out[92]), .A2(_padder__n2554 ), .ZN(
        _padder__n894 ) );
  NAND2_X2 _padder__U392  ( .A1(_padder__n893 ), .A2(_padder__n894 ), .ZN(
        _padder__n1716 ) );
  NAND2_X2 _padder__U391  ( .A1(padder_out[123]), .A2(_padder__n2491 ), .ZN(
        _padder__n891 ) );
  NAND2_X2 _padder__U390  ( .A1(padder_out[91]), .A2(_padder__n2554 ), .ZN(
        _padder__n892 ) );
  NAND2_X2 _padder__U389  ( .A1(_padder__n891 ), .A2(_padder__n892 ), .ZN(
        _padder__n1717 ) );
  NAND2_X2 _padder__U388  ( .A1(padder_out[122]), .A2(_padder__n2491 ), .ZN(
        _padder__n889 ) );
  NAND2_X2 _padder__U387  ( .A1(padder_out[90]), .A2(_padder__n2554 ), .ZN(
        _padder__n890 ) );
  NAND2_X2 _padder__U386  ( .A1(_padder__n889 ), .A2(_padder__n890 ), .ZN(
        _padder__n1718 ) );
  NAND2_X2 _padder__U385  ( .A1(padder_out[121]), .A2(_padder__n2491 ), .ZN(
        _padder__n887 ) );
  NAND2_X2 _padder__U384  ( .A1(padder_out[89]), .A2(_padder__n2554 ), .ZN(
        _padder__n888 ) );
  NAND2_X2 _padder__U383  ( .A1(_padder__n887 ), .A2(_padder__n888 ), .ZN(
        _padder__n1719 ) );
  NAND2_X2 _padder__U382  ( .A1(padder_out[120]), .A2(_padder__n2491 ), .ZN(
        _padder__n885 ) );
  NAND2_X2 _padder__U381  ( .A1(padder_out[88]), .A2(_padder__n2554 ), .ZN(
        _padder__n886 ) );
  NAND2_X2 _padder__U380  ( .A1(_padder__n885 ), .A2(_padder__n886 ), .ZN(
        _padder__n1720 ) );
  NAND2_X2 _padder__U379  ( .A1(padder_out[7]), .A2(_padder__n2491 ), .ZN(
        _padder__n883 ) );
  NAND2_X2 _padder__U378  ( .A1(padder_out[103]), .A2(_padder__n2554 ), .ZN(
        _padder__n884 ) );
  NAND2_X2 _padder__U377  ( .A1(_padder__n883 ), .A2(_padder__n884 ), .ZN(
        _padder__n1721 ) );
  NAND2_X2 _padder__U376  ( .A1(padder_out[6]), .A2(_padder__n2491 ), .ZN(
        _padder__n881 ) );
  NAND2_X2 _padder__U375  ( .A1(padder_out[102]), .A2(_padder__n2554 ), .ZN(
        _padder__n882 ) );
  NAND2_X2 _padder__U374  ( .A1(_padder__n881 ), .A2(_padder__n882 ), .ZN(
        _padder__n1722 ) );
  NAND2_X2 _padder__U373  ( .A1(padder_out[5]), .A2(_padder__n2491 ), .ZN(
        _padder__n879 ) );
  NAND2_X2 _padder__U372  ( .A1(padder_out[101]), .A2(_padder__n2554 ), .ZN(
        _padder__n880 ) );
  NAND2_X2 _padder__U371  ( .A1(_padder__n879 ), .A2(_padder__n880 ), .ZN(
        _padder__n1723 ) );
  NAND2_X2 _padder__U370  ( .A1(padder_out[4]), .A2(_padder__n2491 ), .ZN(
        _padder__n877 ) );
  NAND2_X2 _padder__U369  ( .A1(padder_out[100]), .A2(_padder__n2554 ), .ZN(
        _padder__n878 ) );
  NAND2_X2 _padder__U368  ( .A1(_padder__n877 ), .A2(_padder__n878 ), .ZN(
        _padder__n1724 ) );
  NAND2_X2 _padder__U367  ( .A1(padder_out[3]), .A2(_padder__n2491 ), .ZN(
        _padder__n875 ) );
  NAND2_X2 _padder__U366  ( .A1(padder_out[99]), .A2(_padder__n2555 ), .ZN(
        _padder__n876 ) );
  NAND2_X2 _padder__U365  ( .A1(_padder__n875 ), .A2(_padder__n876 ), .ZN(
        _padder__n1725 ) );
  NAND2_X2 _padder__U364  ( .A1(padder_out[2]), .A2(_padder__n2491 ), .ZN(
        _padder__n873 ) );
  NAND2_X2 _padder__U363  ( .A1(padder_out[98]), .A2(_padder__n2555 ), .ZN(
        _padder__n874 ) );
  NAND2_X2 _padder__U362  ( .A1(_padder__n873 ), .A2(_padder__n874 ), .ZN(
        _padder__n1726 ) );
  NAND2_X2 _padder__U361  ( .A1(padder_out[1]), .A2(_padder__n2491 ), .ZN(
        _padder__n871 ) );
  NAND2_X2 _padder__U360  ( .A1(padder_out[97]), .A2(_padder__n2555 ), .ZN(
        _padder__n872 ) );
  NAND2_X2 _padder__U359  ( .A1(_padder__n871 ), .A2(_padder__n872 ), .ZN(
        _padder__n1727 ) );
  NAND2_X2 _padder__U358  ( .A1(padder_out[0]), .A2(_padder__n2491 ), .ZN(
        _padder__n869 ) );
  NAND2_X2 _padder__U357  ( .A1(padder_out[96]), .A2(_padder__n2555 ), .ZN(
        _padder__n870 ) );
  NAND2_X2 _padder__U356  ( .A1(_padder__n869 ), .A2(_padder__n870 ), .ZN(
        _padder__n1728 ) );
  NAND2_X2 _padder__U355  ( .A1(padder_out[15]), .A2(_padder__n2491 ), .ZN(
        _padder__n867 ) );
  NAND2_X2 _padder__U354  ( .A1(padder_out[111]), .A2(_padder__n2555 ), .ZN(
        _padder__n868 ) );
  NAND2_X2 _padder__U353  ( .A1(_padder__n867 ), .A2(_padder__n868 ), .ZN(
        _padder__n1729 ) );
  NAND2_X2 _padder__U352  ( .A1(padder_out[14]), .A2(_padder__n2491 ), .ZN(
        _padder__n865 ) );
  NAND2_X2 _padder__U351  ( .A1(padder_out[110]), .A2(_padder__n2555 ), .ZN(
        _padder__n866 ) );
  NAND2_X2 _padder__U350  ( .A1(_padder__n865 ), .A2(_padder__n866 ), .ZN(
        _padder__n1730 ) );
  NAND2_X2 _padder__U349  ( .A1(padder_out[13]), .A2(_padder__n2491 ), .ZN(
        _padder__n863 ) );
  NAND2_X2 _padder__U348  ( .A1(padder_out[109]), .A2(_padder__n2555 ), .ZN(
        _padder__n864 ) );
  NAND2_X2 _padder__U347  ( .A1(_padder__n863 ), .A2(_padder__n864 ), .ZN(
        _padder__n1731 ) );
  NAND2_X2 _padder__U346  ( .A1(padder_out[12]), .A2(_padder__n2491 ), .ZN(
        _padder__n861 ) );
  NAND2_X2 _padder__U345  ( .A1(padder_out[108]), .A2(_padder__n2555 ), .ZN(
        _padder__n862 ) );
  NAND2_X2 _padder__U344  ( .A1(_padder__n861 ), .A2(_padder__n862 ), .ZN(
        _padder__n1732 ) );
  NAND2_X2 _padder__U343  ( .A1(padder_out[11]), .A2(_padder__n2490 ), .ZN(
        _padder__n859 ) );
  NAND2_X2 _padder__U342  ( .A1(padder_out[107]), .A2(_padder__n2555 ), .ZN(
        _padder__n860 ) );
  NAND2_X2 _padder__U341  ( .A1(_padder__n859 ), .A2(_padder__n860 ), .ZN(
        _padder__n1733 ) );
  NAND2_X2 _padder__U340  ( .A1(padder_out[10]), .A2(_padder__n2490 ), .ZN(
        _padder__n857 ) );
  NAND2_X2 _padder__U339  ( .A1(padder_out[106]), .A2(_padder__n2555 ), .ZN(
        _padder__n858 ) );
  NAND2_X2 _padder__U338  ( .A1(_padder__n857 ), .A2(_padder__n858 ), .ZN(
        _padder__n1734 ) );
  NAND2_X2 _padder__U337  ( .A1(padder_out[9]), .A2(_padder__n2490 ), .ZN(
        _padder__n855 ) );
  NAND2_X2 _padder__U336  ( .A1(padder_out[105]), .A2(_padder__n2555 ), .ZN(
        _padder__n856 ) );
  NAND2_X2 _padder__U335  ( .A1(_padder__n855 ), .A2(_padder__n856 ), .ZN(
        _padder__n1735 ) );
  NAND2_X2 _padder__U334  ( .A1(padder_out[8]), .A2(_padder__n2490 ), .ZN(
        _padder__n853 ) );
  NAND2_X2 _padder__U333  ( .A1(padder_out[104]), .A2(_padder__n2556 ), .ZN(
        _padder__n854 ) );
  NAND2_X2 _padder__U332  ( .A1(_padder__n853 ), .A2(_padder__n854 ), .ZN(
        _padder__n1736 ) );
  NAND2_X2 _padder__U331  ( .A1(padder_out[23]), .A2(_padder__n2490 ), .ZN(
        _padder__n851 ) );
  NAND2_X2 _padder__U330  ( .A1(padder_out[119]), .A2(_padder__n2556 ), .ZN(
        _padder__n852 ) );
  NAND2_X2 _padder__U329  ( .A1(_padder__n851 ), .A2(_padder__n852 ), .ZN(
        _padder__n1737 ) );
  NAND2_X2 _padder__U328  ( .A1(padder_out[22]), .A2(_padder__n2490 ), .ZN(
        _padder__n849 ) );
  NAND2_X2 _padder__U327  ( .A1(padder_out[118]), .A2(_padder__n2556 ), .ZN(
        _padder__n850 ) );
  NAND2_X2 _padder__U326  ( .A1(_padder__n849 ), .A2(_padder__n850 ), .ZN(
        _padder__n1738 ) );
  NAND2_X2 _padder__U325  ( .A1(padder_out[21]), .A2(_padder__n2490 ), .ZN(
        _padder__n847 ) );
  NAND2_X2 _padder__U324  ( .A1(padder_out[117]), .A2(_padder__n2556 ), .ZN(
        _padder__n848 ) );
  NAND2_X2 _padder__U323  ( .A1(_padder__n847 ), .A2(_padder__n848 ), .ZN(
        _padder__n1739 ) );
  NAND2_X2 _padder__U322  ( .A1(padder_out[20]), .A2(_padder__n2490 ), .ZN(
        _padder__n845 ) );
  NAND2_X2 _padder__U321  ( .A1(padder_out[116]), .A2(_padder__n2556 ), .ZN(
        _padder__n846 ) );
  NAND2_X2 _padder__U320  ( .A1(_padder__n845 ), .A2(_padder__n846 ), .ZN(
        _padder__n1740 ) );
  NAND2_X2 _padder__U319  ( .A1(padder_out[19]), .A2(_padder__n2490 ), .ZN(
        _padder__n843 ) );
  NAND2_X2 _padder__U318  ( .A1(padder_out[115]), .A2(_padder__n2556 ), .ZN(
        _padder__n844 ) );
  NAND2_X2 _padder__U317  ( .A1(_padder__n843 ), .A2(_padder__n844 ), .ZN(
        _padder__n1741 ) );
  NAND2_X2 _padder__U316  ( .A1(padder_out[18]), .A2(_padder__n2490 ), .ZN(
        _padder__n841 ) );
  NAND2_X2 _padder__U315  ( .A1(padder_out[114]), .A2(_padder__n2556 ), .ZN(
        _padder__n842 ) );
  NAND2_X2 _padder__U314  ( .A1(_padder__n841 ), .A2(_padder__n842 ), .ZN(
        _padder__n1742 ) );
  NAND2_X2 _padder__U313  ( .A1(padder_out[17]), .A2(_padder__n2490 ), .ZN(
        _padder__n839 ) );
  NAND2_X2 _padder__U312  ( .A1(padder_out[113]), .A2(_padder__n2556 ), .ZN(
        _padder__n840 ) );
  NAND2_X2 _padder__U311  ( .A1(_padder__n839 ), .A2(_padder__n840 ), .ZN(
        _padder__n1743 ) );
  NAND2_X2 _padder__U310  ( .A1(padder_out[16]), .A2(_padder__n2490 ), .ZN(
        _padder__n837 ) );
  NAND2_X2 _padder__U309  ( .A1(padder_out[112]), .A2(_padder__n2556 ), .ZN(
        _padder__n838 ) );
  NAND2_X2 _padder__U308  ( .A1(_padder__n837 ), .A2(_padder__n838 ), .ZN(
        _padder__n1744 ) );
  NAND2_X2 _padder__U307  ( .A1(padder_out[31]), .A2(_padder__n2490 ), .ZN(
        _padder__n835 ) );
  NAND2_X2 _padder__U306  ( .A1(padder_out[127]), .A2(_padder__n2556 ), .ZN(
        _padder__n836 ) );
  NAND2_X2 _padder__U305  ( .A1(_padder__n835 ), .A2(_padder__n836 ), .ZN(
        _padder__n1745 ) );
  NAND2_X2 _padder__U304  ( .A1(padder_out[30]), .A2(_padder__n2490 ), .ZN(
        _padder__n833 ) );
  NAND2_X2 _padder__U303  ( .A1(padder_out[126]), .A2(_padder__n2556 ), .ZN(
        _padder__n834 ) );
  NAND2_X2 _padder__U302  ( .A1(_padder__n833 ), .A2(_padder__n834 ), .ZN(
        _padder__n1746 ) );
  NAND2_X2 _padder__U301  ( .A1(padder_out[29]), .A2(_padder__n2490 ), .ZN(
        _padder__n831 ) );
  NAND2_X2 _padder__U300  ( .A1(padder_out[125]), .A2(_padder__n2557 ), .ZN(
        _padder__n832 ) );
  NAND2_X2 _padder__U299  ( .A1(_padder__n831 ), .A2(_padder__n832 ), .ZN(
        _padder__n1747 ) );
  NAND2_X2 _padder__U298  ( .A1(padder_out[28]), .A2(_padder__n2490 ), .ZN(
        _padder__n829 ) );
  NAND2_X2 _padder__U297  ( .A1(padder_out[124]), .A2(_padder__n2557 ), .ZN(
        _padder__n830 ) );
  NAND2_X2 _padder__U296  ( .A1(_padder__n829 ), .A2(_padder__n830 ), .ZN(
        _padder__n1748 ) );
  NAND2_X2 _padder__U295  ( .A1(padder_out[27]), .A2(_padder__n2490 ), .ZN(
        _padder__n827 ) );
  NAND2_X2 _padder__U294  ( .A1(padder_out[123]), .A2(_padder__n2557 ), .ZN(
        _padder__n828 ) );
  NAND2_X2 _padder__U293  ( .A1(_padder__n827 ), .A2(_padder__n828 ), .ZN(
        _padder__n1749 ) );
  NAND2_X2 _padder__U292  ( .A1(padder_out[26]), .A2(_padder__n2490 ), .ZN(
        _padder__n825 ) );
  NAND2_X2 _padder__U291  ( .A1(padder_out[122]), .A2(_padder__n2557 ), .ZN(
        _padder__n826 ) );
  NAND2_X2 _padder__U290  ( .A1(_padder__n825 ), .A2(_padder__n826 ), .ZN(
        _padder__n1750 ) );
  NAND2_X2 _padder__U289  ( .A1(padder_out[25]), .A2(_padder__n2490 ), .ZN(
        _padder__n823 ) );
  NAND2_X2 _padder__U288  ( .A1(padder_out[121]), .A2(_padder__n2557 ), .ZN(
        _padder__n824 ) );
  NAND2_X2 _padder__U287  ( .A1(_padder__n823 ), .A2(_padder__n824 ), .ZN(
        _padder__n1751 ) );
  NAND2_X2 _padder__U286  ( .A1(padder_out[24]), .A2(_padder__n2490 ), .ZN(
        _padder__n821 ) );
  NAND2_X2 _padder__U285  ( .A1(padder_out[120]), .A2(_padder__n2557 ), .ZN(
        _padder__n822 ) );
  NAND2_X2 _padder__U284  ( .A1(_padder__n821 ), .A2(_padder__n822 ), .ZN(
        _padder__n1752 ) );
  NAND2_X2 _padder__U283  ( .A1(padder_out[39]), .A2(_padder__n2490 ), .ZN(
        _padder__n819 ) );
  NAND2_X2 _padder__U282  ( .A1(padder_out[7]), .A2(_padder__n2557 ), .ZN(
        _padder__n820 ) );
  NAND2_X2 _padder__U281  ( .A1(_padder__n819 ), .A2(_padder__n820 ), .ZN(
        _padder__n1753 ) );
  NAND2_X2 _padder__U280  ( .A1(padder_out[38]), .A2(_padder__n2490 ), .ZN(
        _padder__n817 ) );
  NAND2_X2 _padder__U279  ( .A1(padder_out[6]), .A2(_padder__n2557 ), .ZN(
        _padder__n818 ) );
  NAND2_X2 _padder__U278  ( .A1(_padder__n817 ), .A2(_padder__n818 ), .ZN(
        _padder__n1754 ) );
  NAND2_X2 _padder__U277  ( .A1(padder_out[37]), .A2(_padder__n2490 ), .ZN(
        _padder__n815 ) );
  NAND2_X2 _padder__U276  ( .A1(padder_out[5]), .A2(_padder__n2557 ), .ZN(
        _padder__n816 ) );
  NAND2_X2 _padder__U275  ( .A1(_padder__n815 ), .A2(_padder__n816 ), .ZN(
        _padder__n1755 ) );
  NAND2_X2 _padder__U274  ( .A1(padder_out[36]), .A2(_padder__n2490 ), .ZN(
        _padder__n813 ) );
  NAND2_X2 _padder__U273  ( .A1(padder_out[4]), .A2(_padder__n2557 ), .ZN(
        _padder__n814 ) );
  NAND2_X2 _padder__U272  ( .A1(_padder__n813 ), .A2(_padder__n814 ), .ZN(
        _padder__n1756 ) );
  NAND2_X2 _padder__U271  ( .A1(padder_out[35]), .A2(_padder__n2489 ), .ZN(
        _padder__n811 ) );
  NAND2_X2 _padder__U270  ( .A1(padder_out[3]), .A2(_padder__n2557 ), .ZN(
        _padder__n812 ) );
  NAND2_X2 _padder__U269  ( .A1(_padder__n811 ), .A2(_padder__n812 ), .ZN(
        _padder__n1757 ) );
  NAND2_X2 _padder__U268  ( .A1(padder_out[34]), .A2(_padder__n2489 ), .ZN(
        _padder__n809 ) );
  NAND2_X2 _padder__U267  ( .A1(padder_out[2]), .A2(_padder__n2558 ), .ZN(
        _padder__n810 ) );
  NAND2_X2 _padder__U266  ( .A1(_padder__n809 ), .A2(_padder__n810 ), .ZN(
        _padder__n1758 ) );
  NAND2_X2 _padder__U265  ( .A1(padder_out[33]), .A2(_padder__n2489 ), .ZN(
        _padder__n807 ) );
  NAND2_X2 _padder__U264  ( .A1(padder_out[1]), .A2(_padder__n2558 ), .ZN(
        _padder__n808 ) );
  NAND2_X2 _padder__U263  ( .A1(_padder__n807 ), .A2(_padder__n808 ), .ZN(
        _padder__n1759 ) );
  NAND2_X2 _padder__U262  ( .A1(padder_out[32]), .A2(_padder__n2489 ), .ZN(
        _padder__n805 ) );
  NAND2_X2 _padder__U261  ( .A1(padder_out[0]), .A2(_padder__n2558 ), .ZN(
        _padder__n806 ) );
  NAND2_X2 _padder__U260  ( .A1(_padder__n805 ), .A2(_padder__n806 ), .ZN(
        _padder__n1760 ) );
  NAND2_X2 _padder__U259  ( .A1(padder_out[47]), .A2(_padder__n2489 ), .ZN(
        _padder__n803 ) );
  NAND2_X2 _padder__U258  ( .A1(padder_out[15]), .A2(_padder__n2558 ), .ZN(
        _padder__n804 ) );
  NAND2_X2 _padder__U257  ( .A1(_padder__n803 ), .A2(_padder__n804 ), .ZN(
        _padder__n1761 ) );
  NAND2_X2 _padder__U256  ( .A1(padder_out[46]), .A2(_padder__n2489 ), .ZN(
        _padder__n801 ) );
  NAND2_X2 _padder__U255  ( .A1(padder_out[14]), .A2(_padder__n2558 ), .ZN(
        _padder__n802 ) );
  NAND2_X2 _padder__U254  ( .A1(_padder__n801 ), .A2(_padder__n802 ), .ZN(
        _padder__n1762 ) );
  NAND2_X2 _padder__U253  ( .A1(padder_out[45]), .A2(_padder__n2489 ), .ZN(
        _padder__n799 ) );
  NAND2_X2 _padder__U252  ( .A1(padder_out[13]), .A2(_padder__n2558 ), .ZN(
        _padder__n800 ) );
  NAND2_X2 _padder__U251  ( .A1(_padder__n799 ), .A2(_padder__n800 ), .ZN(
        _padder__n1763 ) );
  NAND2_X2 _padder__U250  ( .A1(padder_out[44]), .A2(_padder__n2489 ), .ZN(
        _padder__n797 ) );
  NAND2_X2 _padder__U249  ( .A1(padder_out[12]), .A2(_padder__n2558 ), .ZN(
        _padder__n798 ) );
  NAND2_X2 _padder__U248  ( .A1(_padder__n797 ), .A2(_padder__n798 ), .ZN(
        _padder__n1764 ) );
  NAND2_X2 _padder__U247  ( .A1(padder_out[43]), .A2(_padder__n2489 ), .ZN(
        _padder__n795 ) );
  NAND2_X2 _padder__U246  ( .A1(padder_out[11]), .A2(_padder__n2558 ), .ZN(
        _padder__n796 ) );
  NAND2_X2 _padder__U245  ( .A1(_padder__n795 ), .A2(_padder__n796 ), .ZN(
        _padder__n1765 ) );
  NAND2_X2 _padder__U244  ( .A1(padder_out[42]), .A2(_padder__n2489 ), .ZN(
        _padder__n793 ) );
  NAND2_X2 _padder__U243  ( .A1(padder_out[10]), .A2(_padder__n2558 ), .ZN(
        _padder__n794 ) );
  NAND2_X2 _padder__U242  ( .A1(_padder__n793 ), .A2(_padder__n794 ), .ZN(
        _padder__n1766 ) );
  NAND2_X2 _padder__U241  ( .A1(padder_out[41]), .A2(_padder__n2489 ), .ZN(
        _padder__n791 ) );
  NAND2_X2 _padder__U240  ( .A1(padder_out[9]), .A2(_padder__n2558 ), .ZN(
        _padder__n792 ) );
  NAND2_X2 _padder__U239  ( .A1(_padder__n791 ), .A2(_padder__n792 ), .ZN(
        _padder__n1767 ) );
  NAND2_X2 _padder__U238  ( .A1(padder_out[40]), .A2(_padder__n2489 ), .ZN(
        _padder__n789 ) );
  NAND2_X2 _padder__U237  ( .A1(padder_out[8]), .A2(_padder__n2558 ), .ZN(
        _padder__n790 ) );
  NAND2_X2 _padder__U236  ( .A1(_padder__n789 ), .A2(_padder__n790 ), .ZN(
        _padder__n1768 ) );
  NAND2_X2 _padder__U235  ( .A1(padder_out[55]), .A2(_padder__n2489 ), .ZN(
        _padder__n787 ) );
  NAND2_X2 _padder__U234  ( .A1(padder_out[23]), .A2(_padder__n2559 ), .ZN(
        _padder__n788 ) );
  NAND2_X2 _padder__U233  ( .A1(_padder__n787 ), .A2(_padder__n788 ), .ZN(
        _padder__n1769 ) );
  NAND2_X2 _padder__U232  ( .A1(padder_out[54]), .A2(_padder__n2489 ), .ZN(
        _padder__n785 ) );
  NAND2_X2 _padder__U231  ( .A1(padder_out[22]), .A2(_padder__n2559 ), .ZN(
        _padder__n786 ) );
  NAND2_X2 _padder__U230  ( .A1(_padder__n785 ), .A2(_padder__n786 ), .ZN(
        _padder__n1770 ) );
  NAND2_X2 _padder__U229  ( .A1(padder_out[53]), .A2(_padder__n2489 ), .ZN(
        _padder__n783 ) );
  NAND2_X2 _padder__U228  ( .A1(padder_out[21]), .A2(_padder__n2559 ), .ZN(
        _padder__n784 ) );
  NAND2_X2 _padder__U227  ( .A1(_padder__n783 ), .A2(_padder__n784 ), .ZN(
        _padder__n1771 ) );
  NAND2_X2 _padder__U226  ( .A1(padder_out[52]), .A2(_padder__n2489 ), .ZN(
        _padder__n781 ) );
  NAND2_X2 _padder__U225  ( .A1(padder_out[20]), .A2(_padder__n2559 ), .ZN(
        _padder__n782 ) );
  NAND2_X2 _padder__U224  ( .A1(_padder__n781 ), .A2(_padder__n782 ), .ZN(
        _padder__n1772 ) );
  NAND2_X2 _padder__U223  ( .A1(padder_out[51]), .A2(_padder__n2489 ), .ZN(
        _padder__n779 ) );
  NAND2_X2 _padder__U222  ( .A1(padder_out[19]), .A2(_padder__n2559 ), .ZN(
        _padder__n780 ) );
  NAND2_X2 _padder__U221  ( .A1(_padder__n779 ), .A2(_padder__n780 ), .ZN(
        _padder__n1773 ) );
  NAND2_X2 _padder__U220  ( .A1(padder_out[50]), .A2(_padder__n2489 ), .ZN(
        _padder__n777 ) );
  NAND2_X2 _padder__U219  ( .A1(padder_out[18]), .A2(_padder__n2559 ), .ZN(
        _padder__n778 ) );
  NAND2_X2 _padder__U218  ( .A1(_padder__n777 ), .A2(_padder__n778 ), .ZN(
        _padder__n1774 ) );
  NAND2_X2 _padder__U217  ( .A1(padder_out[49]), .A2(_padder__n2489 ), .ZN(
        _padder__n775 ) );
  NAND2_X2 _padder__U216  ( .A1(padder_out[17]), .A2(_padder__n2559 ), .ZN(
        _padder__n776 ) );
  NAND2_X2 _padder__U215  ( .A1(_padder__n775 ), .A2(_padder__n776 ), .ZN(
        _padder__n1775 ) );
  NAND2_X2 _padder__U214  ( .A1(padder_out[48]), .A2(_padder__n2489 ), .ZN(
        _padder__n773 ) );
  NAND2_X2 _padder__U213  ( .A1(padder_out[16]), .A2(_padder__n2559 ), .ZN(
        _padder__n774 ) );
  NAND2_X2 _padder__U212  ( .A1(_padder__n773 ), .A2(_padder__n774 ), .ZN(
        _padder__n1776 ) );
  NAND2_X2 _padder__U211  ( .A1(padder_out[63]), .A2(_padder__n2489 ), .ZN(
        _padder__n771 ) );
  NAND2_X2 _padder__U210  ( .A1(padder_out[31]), .A2(_padder__n2559 ), .ZN(
        _padder__n772 ) );
  NAND2_X2 _padder__U209  ( .A1(_padder__n771 ), .A2(_padder__n772 ), .ZN(
        _padder__n1777 ) );
  NAND2_X2 _padder__U208  ( .A1(padder_out[62]), .A2(_padder__n2489 ), .ZN(
        _padder__n769 ) );
  NAND2_X2 _padder__U207  ( .A1(padder_out[30]), .A2(_padder__n2559 ), .ZN(
        _padder__n770 ) );
  NAND2_X2 _padder__U206  ( .A1(_padder__n769 ), .A2(_padder__n770 ), .ZN(
        _padder__n1778 ) );
  NAND2_X2 _padder__U205  ( .A1(padder_out[61]), .A2(_padder__n2489 ), .ZN(
        _padder__n767 ) );
  NAND2_X2 _padder__U204  ( .A1(padder_out[29]), .A2(_padder__n2559 ), .ZN(
        _padder__n768 ) );
  NAND2_X2 _padder__U203  ( .A1(_padder__n767 ), .A2(_padder__n768 ), .ZN(
        _padder__n1779 ) );
  NAND2_X2 _padder__U202  ( .A1(padder_out[60]), .A2(_padder__n2489 ), .ZN(
        _padder__n765 ) );
  NAND2_X2 _padder__U201  ( .A1(padder_out[28]), .A2(_padder__n2560 ), .ZN(
        _padder__n766 ) );
  NAND2_X2 _padder__U200  ( .A1(_padder__n765 ), .A2(_padder__n766 ), .ZN(
        _padder__n1780 ) );
  NAND2_X2 _padder__U199  ( .A1(padder_out[59]), .A2(_padder__n2488 ), .ZN(
        _padder__n763 ) );
  NAND2_X2 _padder__U198  ( .A1(padder_out[27]), .A2(_padder__n2560 ), .ZN(
        _padder__n764 ) );
  NAND2_X2 _padder__U197  ( .A1(_padder__n763 ), .A2(_padder__n764 ), .ZN(
        _padder__n1781 ) );
  NAND2_X2 _padder__U196  ( .A1(padder_out[58]), .A2(_padder__n2488 ), .ZN(
        _padder__n761 ) );
  NAND2_X2 _padder__U195  ( .A1(padder_out[26]), .A2(_padder__n2560 ), .ZN(
        _padder__n762 ) );
  NAND2_X2 _padder__U194  ( .A1(_padder__n761 ), .A2(_padder__n762 ), .ZN(
        _padder__n1782 ) );
  NAND2_X2 _padder__U193  ( .A1(padder_out[57]), .A2(_padder__n2488 ), .ZN(
        _padder__n759 ) );
  NAND2_X2 _padder__U192  ( .A1(padder_out[25]), .A2(_padder__n2560 ), .ZN(
        _padder__n760 ) );
  NAND2_X2 _padder__U191  ( .A1(_padder__n759 ), .A2(_padder__n760 ), .ZN(
        _padder__n1783 ) );
  NAND2_X2 _padder__U190  ( .A1(padder_out[56]), .A2(_padder__n2491 ), .ZN(
        _padder__n757 ) );
  NAND2_X2 _padder__U189  ( .A1(padder_out[24]), .A2(_padder__n2560 ), .ZN(
        _padder__n758 ) );
  NAND2_X2 _padder__U188  ( .A1(_padder__n757 ), .A2(_padder__n758 ), .ZN(
        _padder__n1784 ) );
  NAND2_X2 _padder__U186  ( .A1(_padder__v0[31]), .A2(_padder__n2571 ), .ZN(
        _padder__n754 ) );
  NAND2_X2 _padder__U183  ( .A1(padder_out[39]), .A2(_padder__n2560 ), .ZN(
        _padder__n756 ) );
  NAND2_X2 _padder__U181  ( .A1(_padder__v0[30]), .A2(_padder__n2571 ), .ZN(
        _padder__n751 ) );
  NAND2_X2 _padder__U179  ( .A1(padder_out[38]), .A2(_padder__n2560 ), .ZN(
        _padder__n753 ) );
  NAND2_X2 _padder__U177  ( .A1(_padder__v0[29]), .A2(_padder__n2571 ), .ZN(
        _padder__n748 ) );
  NAND2_X2 _padder__U175  ( .A1(padder_out[37]), .A2(_padder__n2560 ), .ZN(
        _padder__n750 ) );
  NAND2_X2 _padder__U173  ( .A1(_padder__v0[28]), .A2(_padder__n2571 ), .ZN(
        _padder__n745 ) );
  NAND2_X2 _padder__U171  ( .A1(padder_out[36]), .A2(_padder__n2560 ), .ZN(
        _padder__n747 ) );
  NAND2_X2 _padder__U169  ( .A1(_padder__v0[27]), .A2(_padder__n2571 ), .ZN(
        _padder__n742 ) );
  NAND2_X2 _padder__U167  ( .A1(padder_out[35]), .A2(_padder__n2560 ), .ZN(
        _padder__n744 ) );
  NAND2_X2 _padder__U165  ( .A1(_padder__v0[26]), .A2(_padder__n2571 ), .ZN(
        _padder__n739 ) );
  NAND2_X2 _padder__U163  ( .A1(padder_out[34]), .A2(_padder__n2560 ), .ZN(
        _padder__n741 ) );
  NAND2_X2 _padder__U161  ( .A1(_padder__v0[25]), .A2(_padder__n2571 ), .ZN(
        _padder__n736 ) );
  NAND2_X2 _padder__U159  ( .A1(padder_out[33]), .A2(_padder__n2561 ), .ZN(
        _padder__n738 ) );
  NAND2_X2 _padder__U157  ( .A1(_padder__v0[24]), .A2(_padder__n2571 ), .ZN(
        _padder__n733 ) );
  NAND2_X2 _padder__U155  ( .A1(padder_out[32]), .A2(_padder__n2561 ), .ZN(
        _padder__n735 ) );
  NAND2_X2 _padder__U153  ( .A1(_padder__v0[23]), .A2(_padder__n2571 ), .ZN(
        _padder__n730 ) );
  NAND2_X2 _padder__U151  ( .A1(padder_out[47]), .A2(_padder__n2561 ), .ZN(
        _padder__n732 ) );
  NAND2_X2 _padder__U149  ( .A1(_padder__v0[22]), .A2(_padder__n2571 ), .ZN(
        _padder__n727 ) );
  NAND2_X2 _padder__U147  ( .A1(padder_out[46]), .A2(_padder__n2561 ), .ZN(
        _padder__n729 ) );
  NAND2_X2 _padder__U145  ( .A1(_padder__v0[21]), .A2(_padder__n2571 ), .ZN(
        _padder__n724 ) );
  NAND2_X2 _padder__U143  ( .A1(padder_out[45]), .A2(_padder__n2561 ), .ZN(
        _padder__n726 ) );
  NAND2_X2 _padder__U141  ( .A1(_padder__v0[20]), .A2(_padder__n2571 ), .ZN(
        _padder__n721 ) );
  NAND2_X2 _padder__U139  ( .A1(padder_out[44]), .A2(_padder__n2561 ), .ZN(
        _padder__n723 ) );
  NAND2_X2 _padder__U137  ( .A1(_padder__v0[19]), .A2(_padder__n2571 ), .ZN(
        _padder__n718 ) );
  NAND2_X2 _padder__U135  ( .A1(padder_out[43]), .A2(_padder__n2561 ), .ZN(
        _padder__n720 ) );
  NAND2_X2 _padder__U133  ( .A1(_padder__v0[18]), .A2(_padder__n2571 ), .ZN(
        _padder__n715 ) );
  NAND2_X2 _padder__U131  ( .A1(padder_out[42]), .A2(_padder__n2561 ), .ZN(
        _padder__n717 ) );
  NAND2_X2 _padder__U129  ( .A1(_padder__v0[17]), .A2(_padder__n2570 ), .ZN(
        _padder__n712 ) );
  NAND2_X2 _padder__U127  ( .A1(padder_out[41]), .A2(_padder__n2561 ), .ZN(
        _padder__n714 ) );
  NAND2_X2 _padder__U125  ( .A1(_padder__v0[16]), .A2(_padder__n2570 ), .ZN(
        _padder__n709 ) );
  NAND2_X2 _padder__U123  ( .A1(padder_out[40]), .A2(_padder__n2561 ), .ZN(
        _padder__n711 ) );
  NAND2_X2 _padder__U121  ( .A1(_padder__v0[15]), .A2(_padder__n2570 ), .ZN(
        _padder__n706 ) );
  NAND2_X2 _padder__U119  ( .A1(padder_out[55]), .A2(_padder__n2561 ), .ZN(
        _padder__n708 ) );
  NAND2_X2 _padder__U117  ( .A1(_padder__v0[14]), .A2(_padder__n2570 ), .ZN(
        _padder__n703 ) );
  NAND2_X2 _padder__U115  ( .A1(padder_out[54]), .A2(_padder__n2562 ), .ZN(
        _padder__n705 ) );
  NAND2_X2 _padder__U113  ( .A1(_padder__v0[13]), .A2(_padder__n2570 ), .ZN(
        _padder__n700 ) );
  NAND2_X2 _padder__U111  ( .A1(padder_out[53]), .A2(_padder__n2562 ), .ZN(
        _padder__n702 ) );
  NAND2_X2 _padder__U109  ( .A1(_padder__v0[12]), .A2(_padder__n2570 ), .ZN(
        _padder__n697 ) );
  NAND2_X2 _padder__U107  ( .A1(padder_out[52]), .A2(_padder__n2562 ), .ZN(
        _padder__n699 ) );
  NAND2_X2 _padder__U105  ( .A1(_padder__v0[11]), .A2(_padder__n2570 ), .ZN(
        _padder__n694 ) );
  NAND2_X2 _padder__U103  ( .A1(padder_out[51]), .A2(_padder__n2562 ), .ZN(
        _padder__n696 ) );
  NAND2_X2 _padder__U101  ( .A1(_padder__v0[10]), .A2(_padder__n2570 ), .ZN(
        _padder__n691 ) );
  NAND2_X2 _padder__U99  ( .A1(padder_out[50]), .A2(_padder__n2562 ), .ZN(
        _padder__n693 ) );
  NAND2_X2 _padder__U97  ( .A1(_padder__v0[9]), .A2(_padder__n2570 ), .ZN(
        _padder__n688 ) );
  NAND2_X2 _padder__U95  ( .A1(padder_out[49]), .A2(_padder__n2562 ), .ZN(
        _padder__n690 ) );
  NAND2_X2 _padder__U93  ( .A1(_padder__v0[8]), .A2(_padder__n2570 ), .ZN(
        _padder__n685 ) );
  NAND2_X2 _padder__U91  ( .A1(padder_out[48]), .A2(_padder__n2562 ), .ZN(
        _padder__n687 ) );
  NAND2_X2 _padder__U88  ( .A1(_padder__n2484 ), .A2(_padder__state ), .ZN(
        _padder__n683 ) );
  NAND2_X2 _padder__U87  ( .A1(_padder__n682 ), .A2(_padder__n683 ), .ZN(
        _padder__n681 ) );
  NAND2_X2 _padder__U86  ( .A1(_padder__n681 ), .A2(_padder__n619 ), .ZN(
        _padder__n679 ) );
  NAND2_X2 _padder__U85  ( .A1(padder_out[63]), .A2(_padder__n2562 ), .ZN(
        _padder__n680 ) );
  NAND2_X2 _padder__U83  ( .A1(padder_out[62]), .A2(_padder__n2562 ), .ZN(
        _padder__n676 ) );
  NAND2_X2 _padder__U81  ( .A1(_padder__n676 ), .A2(_padder__n2474 ), .ZN(
        _padder__n1810 ) );
  NAND2_X2 _padder__U80  ( .A1(padder_out[61]), .A2(_padder__n2562 ), .ZN(
        _padder__n674 ) );
  NAND2_X2 _padder__U78  ( .A1(_padder__n674 ), .A2(_padder__n2473 ), .ZN(
        _padder__n1811 ) );
  NAND2_X2 _padder__U77  ( .A1(padder_out[60]), .A2(_padder__n2562 ), .ZN(
        _padder__n672 ) );
  NAND2_X2 _padder__U75  ( .A1(_padder__n672 ), .A2(_padder__n2447 ), .ZN(
        _padder__n1812 ) );
  NAND2_X2 _padder__U74  ( .A1(padder_out[59]), .A2(_padder__n2555 ), .ZN(
        _padder__n670 ) );
  NAND2_X2 _padder__U72  ( .A1(_padder__n670 ), .A2(_padder__n2478 ), .ZN(
        _padder__n1813 ) );
  NAND2_X2 _padder__U71  ( .A1(padder_out[58]), .A2(_padder__n2556 ), .ZN(
        _padder__n668 ) );
  NAND2_X2 _padder__U69  ( .A1(_padder__n668 ), .A2(_padder__n2477 ), .ZN(
        _padder__n1814 ) );
  NAND2_X2 _padder__U68  ( .A1(padder_out[57]), .A2(_padder__n2569 ), .ZN(
        _padder__n666 ) );
  NAND2_X2 _padder__U66  ( .A1(_padder__n666 ), .A2(_padder__n2476 ), .ZN(
        _padder__n1815 ) );
  NAND2_X2 _padder__U65  ( .A1(_padder__v0[0]), .A2(_padder__n2570 ), .ZN(
        _padder__n662 ) );
  NAND2_X2 _padder__U63  ( .A1(padder_out[56]), .A2(_padder__n2516 ), .ZN(
        _padder__n664 ) );
  NAND2_X2 _padder__U60  ( .A1(_padder__n2445 ), .A2(padder_out_ready), .ZN(
        _padder__n659 ) );
  NAND2_X2 _padder__U58  ( .A1(_padder__n2482 ), .A2(_padder__n619 ), .ZN(
        _padder__n660 ) );
  NAND2_X2 _padder__U57  ( .A1(_padder__n659 ), .A2(_padder__n660 ), .ZN(
        _padder__n1817 ) );
  NAND2_X2 _padder__U56  ( .A1(_padder__n2445 ), .A2(_padder__n619 ), .ZN(
        _padder__n657 ) );
  NAND2_X2 _padder__U55  ( .A1(_padder__n2482 ), .A2(_padder__n618 ), .ZN(
        _padder__n658 ) );
  NAND2_X2 _padder__U54  ( .A1(_padder__n657 ), .A2(_padder__n658 ), .ZN(
        _padder__n1818 ) );
  NAND2_X2 _padder__U53  ( .A1(_padder__n2445 ), .A2(_padder__n618 ), .ZN(
        _padder__n655 ) );
  NAND2_X2 _padder__U52  ( .A1(_padder__n2482 ), .A2(_padder__n617 ), .ZN(
        _padder__n656 ) );
  NAND2_X2 _padder__U51  ( .A1(_padder__n655 ), .A2(_padder__n656 ), .ZN(
        _padder__n1819 ) );
  NAND2_X2 _padder__U50  ( .A1(_padder__n2445 ), .A2(_padder__n617 ), .ZN(
        _padder__n653 ) );
  NAND2_X2 _padder__U49  ( .A1(_padder__n2482 ), .A2(_padder__n616 ), .ZN(
        _padder__n654 ) );
  NAND2_X2 _padder__U48  ( .A1(_padder__n653 ), .A2(_padder__n654 ), .ZN(
        _padder__n1820 ) );
  NAND2_X2 _padder__U47  ( .A1(_padder__n2445 ), .A2(_padder__n616 ), .ZN(
        _padder__n651 ) );
  NAND2_X2 _padder__U46  ( .A1(_padder__n2482 ), .A2(_padder__n615 ), .ZN(
        _padder__n652 ) );
  NAND2_X2 _padder__U45  ( .A1(_padder__n651 ), .A2(_padder__n652 ), .ZN(
        _padder__n1821 ) );
  NAND2_X2 _padder__U44  ( .A1(_padder__n2445 ), .A2(_padder__n615 ), .ZN(
        _padder__n649 ) );
  NAND2_X2 _padder__U43  ( .A1(_padder__n2482 ), .A2(_padder__n614 ), .ZN(
        _padder__n650 ) );
  NAND2_X2 _padder__U42  ( .A1(_padder__n649 ), .A2(_padder__n650 ), .ZN(
        _padder__n1822 ) );
  NAND2_X2 _padder__U41  ( .A1(_padder__n2445 ), .A2(_padder__n614 ), .ZN(
        _padder__n647 ) );
  NAND2_X2 _padder__U40  ( .A1(_padder__n2482 ), .A2(_padder__n613 ), .ZN(
        _padder__n648 ) );
  NAND2_X2 _padder__U39  ( .A1(_padder__n647 ), .A2(_padder__n648 ), .ZN(
        _padder__n1823 ) );
  NAND2_X2 _padder__U38  ( .A1(_padder__n2445 ), .A2(_padder__n613 ), .ZN(
        _padder__n645 ) );
  NAND2_X2 _padder__U37  ( .A1(_padder__n2482 ), .A2(_padder__n612 ), .ZN(
        _padder__n646 ) );
  NAND2_X2 _padder__U36  ( .A1(_padder__n645 ), .A2(_padder__n646 ), .ZN(
        _padder__n1824 ) );
  NAND2_X2 _padder__U35  ( .A1(_padder__n2445 ), .A2(_padder__n612 ), .ZN(
        _padder__n643 ) );
  NAND2_X2 _padder__U34  ( .A1(_padder__n2482 ), .A2(_padder__n611 ), .ZN(
        _padder__n644 ) );
  NAND2_X2 _padder__U33  ( .A1(_padder__n643 ), .A2(_padder__n644 ), .ZN(
        _padder__n1825 ) );
  NAND2_X2 _padder__U32  ( .A1(_padder__n2445 ), .A2(_padder__n611 ), .ZN(
        _padder__n641 ) );
  NAND2_X2 _padder__U31  ( .A1(_padder__n2482 ), .A2(_padder__n610 ), .ZN(
        _padder__n642 ) );
  NAND2_X2 _padder__U30  ( .A1(_padder__n641 ), .A2(_padder__n642 ), .ZN(
        _padder__n1826 ) );
  NAND2_X2 _padder__U29  ( .A1(_padder__n2445 ), .A2(_padder__n610 ), .ZN(
        _padder__n639 ) );
  NAND2_X2 _padder__U28  ( .A1(_padder__n2482 ), .A2(_padder__n609 ), .ZN(
        _padder__n640 ) );
  NAND2_X2 _padder__U27  ( .A1(_padder__n639 ), .A2(_padder__n640 ), .ZN(
        _padder__n1827 ) );
  NAND2_X2 _padder__U26  ( .A1(_padder__n2445 ), .A2(_padder__n609 ), .ZN(
        _padder__n637 ) );
  NAND2_X2 _padder__U25  ( .A1(_padder__n2482 ), .A2(_padder__n608 ), .ZN(
        _padder__n638 ) );
  NAND2_X2 _padder__U24  ( .A1(_padder__n637 ), .A2(_padder__n638 ), .ZN(
        _padder__n1828 ) );
  NAND2_X2 _padder__U23  ( .A1(_padder__n2445 ), .A2(_padder__n608 ), .ZN(
        _padder__n635 ) );
  NAND2_X2 _padder__U22  ( .A1(_padder__n2482 ), .A2(_padder__n607 ), .ZN(
        _padder__n636 ) );
  NAND2_X2 _padder__U21  ( .A1(_padder__n635 ), .A2(_padder__n636 ), .ZN(
        _padder__n1829 ) );
  NAND2_X2 _padder__U20  ( .A1(_padder__n2445 ), .A2(_padder__n607 ), .ZN(
        _padder__n633 ) );
  NAND2_X2 _padder__U19  ( .A1(_padder__n2482 ), .A2(_padder__n606 ), .ZN(
        _padder__n634 ) );
  NAND2_X2 _padder__U18  ( .A1(_padder__n633 ), .A2(_padder__n634 ), .ZN(
        _padder__n1830 ) );
  NAND2_X2 _padder__U17  ( .A1(_padder__n2445 ), .A2(_padder__n606 ), .ZN(
        _padder__n631 ) );
  NAND2_X2 _padder__U16  ( .A1(_padder__n2482 ), .A2(_padder__n605 ), .ZN(
        _padder__n632 ) );
  NAND2_X2 _padder__U15  ( .A1(_padder__n631 ), .A2(_padder__n632 ), .ZN(
        _padder__n1831 ) );
  NAND2_X2 _padder__U14  ( .A1(_padder__n2445 ), .A2(_padder__n605 ), .ZN(
        _padder__n629 ) );
  NAND2_X2 _padder__U13  ( .A1(_padder__n2482 ), .A2(_padder__n604 ), .ZN(
        _padder__n630 ) );
  NAND2_X2 _padder__U12  ( .A1(_padder__n629 ), .A2(_padder__n630 ), .ZN(
        _padder__n1832 ) );
  NAND2_X2 _padder__U11  ( .A1(_padder__n2445 ), .A2(_padder__n604 ), .ZN(
        _padder__n627 ) );
  NAND2_X2 _padder__U10  ( .A1(_padder__n2482 ), .A2(_padder__n603 ), .ZN(
        _padder__n628 ) );
  NAND2_X2 _padder__U9  ( .A1(_padder__n627 ), .A2(_padder__n628 ), .ZN(
        _padder__n1833 ) );
  NAND2_X2 _padder__U8  ( .A1(_padder__n2445 ), .A2(_padder__n603 ), .ZN(
        _padder__n624 ) );
  NAND2_X2 _padder__U7  ( .A1(_padder__n2479 ), .A2(_padder__n624 ), .ZN(
        _padder__n1834 ) );
  DFF_X2 _padder__out_reg_519_  ( .D(_padder__n1297 ), .CK(clk), .Q(
        padder_out[575]), .QN() );
  DFF_X2 _padder__out_reg_487_  ( .D(_padder__n1329 ), .CK(clk), .Q(
        padder_out[479]), .QN() );
  DFF_X2 _padder__out_reg_455_  ( .D(_padder__n1361 ), .CK(clk), .Q(
        padder_out[511]), .QN() );
  DFF_X2 _padder__out_reg_423_  ( .D(_padder__n1393 ), .CK(clk), .Q(
        padder_out[415]), .QN() );
  DFF_X2 _padder__out_reg_391_  ( .D(_padder__n1425 ), .CK(clk), .Q(
        padder_out[447]), .QN() );
  DFF_X2 _padder__out_reg_359_  ( .D(_padder__n1457 ), .CK(clk), .Q(
        padder_out[351]), .QN() );
  DFF_X2 _padder__out_reg_327_  ( .D(_padder__n1489 ), .CK(clk), .Q(
        padder_out[383]), .QN() );
  DFF_X2 _padder__out_reg_295_  ( .D(_padder__n1521 ), .CK(clk), .Q(
        padder_out[287]), .QN() );
  DFF_X2 _padder__out_reg_263_  ( .D(_padder__n1553 ), .CK(clk), .Q(
        padder_out[319]), .QN() );
  DFF_X2 _padder__out_reg_231_  ( .D(_padder__n1585 ), .CK(clk), .Q(
        padder_out[223]), .QN() );
  DFF_X2 _padder__out_reg_199_  ( .D(_padder__n1617 ), .CK(clk), .Q(
        padder_out[255]), .QN() );
  DFF_X2 _padder__out_reg_167_  ( .D(_padder__n1649 ), .CK(clk), .Q(
        padder_out[159]), .QN() );
  DFF_X2 _padder__out_reg_135_  ( .D(_padder__n1681 ), .CK(clk), .Q(
        padder_out[191]), .QN() );
  DFF_X2 _padder__out_reg_103_  ( .D(_padder__n1713 ), .CK(clk), .Q(
        padder_out[95]), .QN() );
  DFF_X2 _padder__out_reg_71_  ( .D(_padder__n1745 ), .CK(clk), .Q(
        padder_out[127]), .QN() );
  DFF_X2 _padder__out_reg_39_  ( .D(_padder__n1777 ), .CK(clk), .Q(
        padder_out[31]), .QN() );
  DFF_X2 _padder__out_reg_7_  ( .D(_padder__n2448 ), .CK(clk), .Q(
        padder_out[63]), .QN() );
  DFF_X2 _padder__i_reg_16_  ( .D(_padder__n1818 ), .CK(clk), .Q(
        _padder__n619 ), .QN() );
  DFF_X2 _padder__i_reg_15_  ( .D(_padder__n1819 ), .CK(clk), .Q(
        _padder__n618 ), .QN() );
  DFF_X2 _padder__i_reg_14_  ( .D(_padder__n1820 ), .CK(clk), .Q(
        _padder__n617 ), .QN() );
  DFF_X2 _padder__i_reg_13_  ( .D(_padder__n1821 ), .CK(clk), .Q(
        _padder__n616 ), .QN() );
  DFF_X2 _padder__i_reg_12_  ( .D(_padder__n1822 ), .CK(clk), .Q(
        _padder__n615 ), .QN() );
  DFF_X2 _padder__i_reg_11_  ( .D(_padder__n1823 ), .CK(clk), .Q(
        _padder__n614 ), .QN() );
  DFF_X2 _padder__i_reg_10_  ( .D(_padder__n1824 ), .CK(clk), .Q(
        _padder__n613 ), .QN() );
  DFF_X2 _padder__i_reg_9_  ( .D(_padder__n1825 ), .CK(clk), .Q(_padder__n612 ), .QN() );
  DFF_X2 _padder__i_reg_8_  ( .D(_padder__n1826 ), .CK(clk), .Q(_padder__n611 ), .QN() );
  DFF_X2 _padder__i_reg_7_  ( .D(_padder__n1827 ), .CK(clk), .Q(_padder__n610 ), .QN() );
  DFF_X2 _padder__i_reg_6_  ( .D(_padder__n1828 ), .CK(clk), .Q(_padder__n609 ), .QN() );
  DFF_X2 _padder__i_reg_5_  ( .D(_padder__n1829 ), .CK(clk), .Q(_padder__n608 ), .QN() );
  DFF_X2 _padder__i_reg_4_  ( .D(_padder__n1830 ), .CK(clk), .Q(_padder__n607 ), .QN() );
  DFF_X2 _padder__i_reg_3_  ( .D(_padder__n1831 ), .CK(clk), .Q(_padder__n606 ), .QN() );
  DFF_X2 _padder__i_reg_2_  ( .D(_padder__n1832 ), .CK(clk), .Q(_padder__n605 ), .QN() );
  DFF_X2 _padder__i_reg_1_  ( .D(_padder__n1833 ), .CK(clk), .Q(_padder__n604 ), .QN() );
  DFF_X2 _padder__i_reg_0_  ( .D(_padder__n1834 ), .CK(clk), .Q(_padder__n603 ), .QN() );
  DFF_X2 _padder__out_reg_512_  ( .D(_padder__n1304 ), .CK(clk), .Q(
        padder_out[568]), .QN() );
  DFF_X2 _padder__out_reg_480_  ( .D(_padder__n1336 ), .CK(clk), .Q(
        padder_out[472]), .QN() );
  DFF_X2 _padder__out_reg_448_  ( .D(_padder__n1368 ), .CK(clk), .Q(
        padder_out[504]), .QN() );
  DFF_X2 _padder__out_reg_416_  ( .D(_padder__n1400 ), .CK(clk), .Q(
        padder_out[408]), .QN() );
  DFF_X2 _padder__out_reg_384_  ( .D(_padder__n1432 ), .CK(clk), .Q(
        padder_out[440]), .QN() );
  DFF_X2 _padder__out_reg_352_  ( .D(_padder__n1464 ), .CK(clk), .Q(
        padder_out[344]), .QN() );
  DFF_X2 _padder__out_reg_320_  ( .D(_padder__n1496 ), .CK(clk), .Q(
        padder_out[376]), .QN() );
  DFF_X2 _padder__out_reg_288_  ( .D(_padder__n1528 ), .CK(clk), .Q(
        padder_out[280]), .QN() );
  DFF_X2 _padder__out_reg_256_  ( .D(_padder__n1560 ), .CK(clk), .Q(
        padder_out[312]), .QN() );
  DFF_X2 _padder__out_reg_224_  ( .D(_padder__n1592 ), .CK(clk), .Q(
        padder_out[216]), .QN() );
  DFF_X2 _padder__out_reg_192_  ( .D(_padder__n1624 ), .CK(clk), .Q(
        padder_out[248]), .QN() );
  DFF_X2 _padder__out_reg_160_  ( .D(_padder__n1656 ), .CK(clk), .Q(
        padder_out[152]), .QN() );
  DFF_X2 _padder__out_reg_128_  ( .D(_padder__n1688 ), .CK(clk), .Q(
        padder_out[184]), .QN() );
  DFF_X2 _padder__out_reg_96_  ( .D(_padder__n1720 ), .CK(clk), .Q(
        padder_out[88]), .QN() );
  DFF_X2 _padder__out_reg_64_  ( .D(_padder__n1752 ), .CK(clk), .Q(
        padder_out[120]), .QN() );
  DFF_X2 _padder__out_reg_32_  ( .D(_padder__n1784 ), .CK(clk), .Q(
        padder_out[24]), .QN() );
  DFF_X2 _padder__out_reg_513_  ( .D(_padder__n1303 ), .CK(clk), .Q(
        padder_out[569]), .QN() );
  DFF_X2 _padder__out_reg_481_  ( .D(_padder__n1335 ), .CK(clk), .Q(
        padder_out[473]), .QN() );
  DFF_X2 _padder__out_reg_449_  ( .D(_padder__n1367 ), .CK(clk), .Q(
        padder_out[505]), .QN() );
  DFF_X2 _padder__out_reg_417_  ( .D(_padder__n1399 ), .CK(clk), .Q(
        padder_out[409]), .QN() );
  DFF_X2 _padder__out_reg_385_  ( .D(_padder__n1431 ), .CK(clk), .Q(
        padder_out[441]), .QN() );
  DFF_X2 _padder__out_reg_353_  ( .D(_padder__n1463 ), .CK(clk), .Q(
        padder_out[345]), .QN() );
  DFF_X2 _padder__out_reg_321_  ( .D(_padder__n1495 ), .CK(clk), .Q(
        padder_out[377]), .QN() );
  DFF_X2 _padder__out_reg_289_  ( .D(_padder__n1527 ), .CK(clk), .Q(
        padder_out[281]), .QN() );
  DFF_X2 _padder__out_reg_257_  ( .D(_padder__n1559 ), .CK(clk), .Q(
        padder_out[313]), .QN() );
  DFF_X2 _padder__out_reg_225_  ( .D(_padder__n1591 ), .CK(clk), .Q(
        padder_out[217]), .QN() );
  DFF_X2 _padder__out_reg_193_  ( .D(_padder__n1623 ), .CK(clk), .Q(
        padder_out[249]), .QN() );
  DFF_X2 _padder__out_reg_161_  ( .D(_padder__n1655 ), .CK(clk), .Q(
        padder_out[153]), .QN() );
  DFF_X2 _padder__out_reg_129_  ( .D(_padder__n1687 ), .CK(clk), .Q(
        padder_out[185]), .QN() );
  DFF_X2 _padder__out_reg_97_  ( .D(_padder__n1719 ), .CK(clk), .Q(
        padder_out[89]), .QN() );
  DFF_X2 _padder__out_reg_65_  ( .D(_padder__n1751 ), .CK(clk), .Q(
        padder_out[121]), .QN() );
  DFF_X2 _padder__out_reg_33_  ( .D(_padder__n1783 ), .CK(clk), .Q(
        padder_out[25]), .QN() );
  DFF_X2 _padder__out_reg_514_  ( .D(_padder__n1302 ), .CK(clk), .Q(
        padder_out[570]), .QN() );
  DFF_X2 _padder__out_reg_482_  ( .D(_padder__n1334 ), .CK(clk), .Q(
        padder_out[474]), .QN() );
  DFF_X2 _padder__out_reg_450_  ( .D(_padder__n1366 ), .CK(clk), .Q(
        padder_out[506]), .QN() );
  DFF_X2 _padder__out_reg_418_  ( .D(_padder__n1398 ), .CK(clk), .Q(
        padder_out[410]), .QN() );
  DFF_X2 _padder__out_reg_386_  ( .D(_padder__n1430 ), .CK(clk), .Q(
        padder_out[442]), .QN() );
  DFF_X2 _padder__out_reg_354_  ( .D(_padder__n1462 ), .CK(clk), .Q(
        padder_out[346]), .QN() );
  DFF_X2 _padder__out_reg_322_  ( .D(_padder__n1494 ), .CK(clk), .Q(
        padder_out[378]), .QN() );
  DFF_X2 _padder__out_reg_290_  ( .D(_padder__n1526 ), .CK(clk), .Q(
        padder_out[282]), .QN() );
  DFF_X2 _padder__out_reg_258_  ( .D(_padder__n1558 ), .CK(clk), .Q(
        padder_out[314]), .QN() );
  DFF_X2 _padder__out_reg_226_  ( .D(_padder__n1590 ), .CK(clk), .Q(
        padder_out[218]), .QN() );
  DFF_X2 _padder__out_reg_194_  ( .D(_padder__n1622 ), .CK(clk), .Q(
        padder_out[250]), .QN() );
  DFF_X2 _padder__out_reg_162_  ( .D(_padder__n1654 ), .CK(clk), .Q(
        padder_out[154]), .QN() );
  DFF_X2 _padder__out_reg_130_  ( .D(_padder__n1686 ), .CK(clk), .Q(
        padder_out[186]), .QN() );
  DFF_X2 _padder__out_reg_98_  ( .D(_padder__n1718 ), .CK(clk), .Q(
        padder_out[90]), .QN() );
  DFF_X2 _padder__out_reg_66_  ( .D(_padder__n1750 ), .CK(clk), .Q(
        padder_out[122]), .QN() );
  DFF_X2 _padder__out_reg_34_  ( .D(_padder__n1782 ), .CK(clk), .Q(
        padder_out[26]), .QN() );
  DFF_X2 _padder__out_reg_515_  ( .D(_padder__n1301 ), .CK(clk), .Q(
        padder_out[571]), .QN() );
  DFF_X2 _padder__out_reg_483_  ( .D(_padder__n1333 ), .CK(clk), .Q(
        padder_out[475]), .QN() );
  DFF_X2 _padder__out_reg_451_  ( .D(_padder__n1365 ), .CK(clk), .Q(
        padder_out[507]), .QN() );
  DFF_X2 _padder__out_reg_419_  ( .D(_padder__n1397 ), .CK(clk), .Q(
        padder_out[411]), .QN() );
  DFF_X2 _padder__out_reg_387_  ( .D(_padder__n1429 ), .CK(clk), .Q(
        padder_out[443]), .QN() );
  DFF_X2 _padder__out_reg_355_  ( .D(_padder__n1461 ), .CK(clk), .Q(
        padder_out[347]), .QN() );
  DFF_X2 _padder__out_reg_323_  ( .D(_padder__n1493 ), .CK(clk), .Q(
        padder_out[379]), .QN() );
  DFF_X2 _padder__out_reg_291_  ( .D(_padder__n1525 ), .CK(clk), .Q(
        padder_out[283]), .QN() );
  DFF_X2 _padder__out_reg_259_  ( .D(_padder__n1557 ), .CK(clk), .Q(
        padder_out[315]), .QN() );
  DFF_X2 _padder__out_reg_227_  ( .D(_padder__n1589 ), .CK(clk), .Q(
        padder_out[219]), .QN() );
  DFF_X2 _padder__out_reg_195_  ( .D(_padder__n1621 ), .CK(clk), .Q(
        padder_out[251]), .QN() );
  DFF_X2 _padder__out_reg_163_  ( .D(_padder__n1653 ), .CK(clk), .Q(
        padder_out[155]), .QN() );
  DFF_X2 _padder__out_reg_131_  ( .D(_padder__n1685 ), .CK(clk), .Q(
        padder_out[187]), .QN() );
  DFF_X2 _padder__out_reg_99_  ( .D(_padder__n1717 ), .CK(clk), .Q(
        padder_out[91]), .QN() );
  DFF_X2 _padder__out_reg_67_  ( .D(_padder__n1749 ), .CK(clk), .Q(
        padder_out[123]), .QN() );
  DFF_X2 _padder__out_reg_35_  ( .D(_padder__n1781 ), .CK(clk), .Q(
        padder_out[27]), .QN() );
  DFF_X2 _padder__out_reg_516_  ( .D(_padder__n1300 ), .CK(clk), .Q(
        padder_out[572]), .QN() );
  DFF_X2 _padder__out_reg_484_  ( .D(_padder__n1332 ), .CK(clk), .Q(
        padder_out[476]), .QN() );
  DFF_X2 _padder__out_reg_452_  ( .D(_padder__n1364 ), .CK(clk), .Q(
        padder_out[508]), .QN() );
  DFF_X2 _padder__out_reg_420_  ( .D(_padder__n1396 ), .CK(clk), .Q(
        padder_out[412]), .QN() );
  DFF_X2 _padder__out_reg_388_  ( .D(_padder__n1428 ), .CK(clk), .Q(
        padder_out[444]), .QN() );
  DFF_X2 _padder__out_reg_356_  ( .D(_padder__n1460 ), .CK(clk), .Q(
        padder_out[348]), .QN() );
  DFF_X2 _padder__out_reg_324_  ( .D(_padder__n1492 ), .CK(clk), .Q(
        padder_out[380]), .QN() );
  DFF_X2 _padder__out_reg_292_  ( .D(_padder__n1524 ), .CK(clk), .Q(
        padder_out[284]), .QN() );
  DFF_X2 _padder__out_reg_260_  ( .D(_padder__n1556 ), .CK(clk), .Q(
        padder_out[316]), .QN() );
  DFF_X2 _padder__out_reg_228_  ( .D(_padder__n1588 ), .CK(clk), .Q(
        padder_out[220]), .QN() );
  DFF_X2 _padder__out_reg_196_  ( .D(_padder__n1620 ), .CK(clk), .Q(
        padder_out[252]), .QN() );
  DFF_X2 _padder__out_reg_164_  ( .D(_padder__n1652 ), .CK(clk), .Q(
        padder_out[156]), .QN() );
  DFF_X2 _padder__out_reg_132_  ( .D(_padder__n1684 ), .CK(clk), .Q(
        padder_out[188]), .QN() );
  DFF_X2 _padder__out_reg_100_  ( .D(_padder__n1716 ), .CK(clk), .Q(
        padder_out[92]), .QN() );
  DFF_X2 _padder__out_reg_68_  ( .D(_padder__n1748 ), .CK(clk), .Q(
        padder_out[124]), .QN() );
  DFF_X2 _padder__out_reg_36_  ( .D(_padder__n1780 ), .CK(clk), .Q(
        padder_out[28]), .QN() );
  DFF_X2 _padder__out_reg_517_  ( .D(_padder__n1299 ), .CK(clk), .Q(
        padder_out[573]), .QN() );
  DFF_X2 _padder__out_reg_485_  ( .D(_padder__n1331 ), .CK(clk), .Q(
        padder_out[477]), .QN() );
  DFF_X2 _padder__out_reg_453_  ( .D(_padder__n1363 ), .CK(clk), .Q(
        padder_out[509]), .QN() );
  DFF_X2 _padder__out_reg_421_  ( .D(_padder__n1395 ), .CK(clk), .Q(
        padder_out[413]), .QN() );
  DFF_X2 _padder__out_reg_389_  ( .D(_padder__n1427 ), .CK(clk), .Q(
        padder_out[445]), .QN() );
  DFF_X2 _padder__out_reg_357_  ( .D(_padder__n1459 ), .CK(clk), .Q(
        padder_out[349]), .QN() );
  DFF_X2 _padder__out_reg_325_  ( .D(_padder__n1491 ), .CK(clk), .Q(
        padder_out[381]), .QN() );
  DFF_X2 _padder__out_reg_293_  ( .D(_padder__n1523 ), .CK(clk), .Q(
        padder_out[285]), .QN() );
  DFF_X2 _padder__out_reg_261_  ( .D(_padder__n1555 ), .CK(clk), .Q(
        padder_out[317]), .QN() );
  DFF_X2 _padder__out_reg_229_  ( .D(_padder__n1587 ), .CK(clk), .Q(
        padder_out[221]), .QN() );
  DFF_X2 _padder__out_reg_197_  ( .D(_padder__n1619 ), .CK(clk), .Q(
        padder_out[253]), .QN() );
  DFF_X2 _padder__out_reg_165_  ( .D(_padder__n1651 ), .CK(clk), .Q(
        padder_out[157]), .QN() );
  DFF_X2 _padder__out_reg_133_  ( .D(_padder__n1683 ), .CK(clk), .Q(
        padder_out[189]), .QN() );
  DFF_X2 _padder__out_reg_101_  ( .D(_padder__n1715 ), .CK(clk), .Q(
        padder_out[93]), .QN() );
  DFF_X2 _padder__out_reg_69_  ( .D(_padder__n1747 ), .CK(clk), .Q(
        padder_out[125]), .QN() );
  DFF_X2 _padder__out_reg_37_  ( .D(_padder__n1779 ), .CK(clk), .Q(
        padder_out[29]), .QN() );
  DFF_X2 _padder__out_reg_518_  ( .D(_padder__n1298 ), .CK(clk), .Q(
        padder_out[574]), .QN() );
  DFF_X2 _padder__out_reg_486_  ( .D(_padder__n1330 ), .CK(clk), .Q(
        padder_out[478]), .QN() );
  DFF_X2 _padder__out_reg_454_  ( .D(_padder__n1362 ), .CK(clk), .Q(
        padder_out[510]), .QN() );
  DFF_X2 _padder__out_reg_422_  ( .D(_padder__n1394 ), .CK(clk), .Q(
        padder_out[414]), .QN() );
  DFF_X2 _padder__out_reg_390_  ( .D(_padder__n1426 ), .CK(clk), .Q(
        padder_out[446]), .QN() );
  DFF_X2 _padder__out_reg_358_  ( .D(_padder__n1458 ), .CK(clk), .Q(
        padder_out[350]), .QN() );
  DFF_X2 _padder__out_reg_326_  ( .D(_padder__n1490 ), .CK(clk), .Q(
        padder_out[382]), .QN() );
  DFF_X2 _padder__out_reg_294_  ( .D(_padder__n1522 ), .CK(clk), .Q(
        padder_out[286]), .QN() );
  DFF_X2 _padder__out_reg_262_  ( .D(_padder__n1554 ), .CK(clk), .Q(
        padder_out[318]), .QN() );
  DFF_X2 _padder__out_reg_230_  ( .D(_padder__n1586 ), .CK(clk), .Q(
        padder_out[222]), .QN() );
  DFF_X2 _padder__out_reg_198_  ( .D(_padder__n1618 ), .CK(clk), .Q(
        padder_out[254]), .QN() );
  DFF_X2 _padder__out_reg_166_  ( .D(_padder__n1650 ), .CK(clk), .Q(
        padder_out[158]), .QN() );
  DFF_X2 _padder__out_reg_134_  ( .D(_padder__n1682 ), .CK(clk), .Q(
        padder_out[190]), .QN() );
  DFF_X2 _padder__out_reg_102_  ( .D(_padder__n1714 ), .CK(clk), .Q(
        padder_out[94]), .QN() );
  DFF_X2 _padder__out_reg_70_  ( .D(_padder__n1746 ), .CK(clk), .Q(
        padder_out[126]), .QN() );
  DFF_X2 _padder__out_reg_38_  ( .D(_padder__n1778 ), .CK(clk), .Q(
        padder_out[30]), .QN() );
  DFF_X2 _padder__out_reg_520_  ( .D(_padder__n1296 ), .CK(clk), .Q(
        padder_out[560]), .QN() );
  DFF_X2 _padder__out_reg_488_  ( .D(_padder__n1328 ), .CK(clk), .Q(
        padder_out[464]), .QN() );
  DFF_X2 _padder__out_reg_456_  ( .D(_padder__n1360 ), .CK(clk), .Q(
        padder_out[496]), .QN() );
  DFF_X2 _padder__out_reg_424_  ( .D(_padder__n1392 ), .CK(clk), .Q(
        padder_out[400]), .QN() );
  DFF_X2 _padder__out_reg_392_  ( .D(_padder__n1424 ), .CK(clk), .Q(
        padder_out[432]), .QN() );
  DFF_X2 _padder__out_reg_360_  ( .D(_padder__n1456 ), .CK(clk), .Q(
        padder_out[336]), .QN() );
  DFF_X2 _padder__out_reg_328_  ( .D(_padder__n1488 ), .CK(clk), .Q(
        padder_out[368]), .QN() );
  DFF_X2 _padder__out_reg_296_  ( .D(_padder__n1520 ), .CK(clk), .Q(
        padder_out[272]), .QN() );
  DFF_X2 _padder__out_reg_264_  ( .D(_padder__n1552 ), .CK(clk), .Q(
        padder_out[304]), .QN() );
  DFF_X2 _padder__out_reg_232_  ( .D(_padder__n1584 ), .CK(clk), .Q(
        padder_out[208]), .QN() );
  DFF_X2 _padder__out_reg_200_  ( .D(_padder__n1616 ), .CK(clk), .Q(
        padder_out[240]), .QN() );
  DFF_X2 _padder__out_reg_168_  ( .D(_padder__n1648 ), .CK(clk), .Q(
        padder_out[144]), .QN() );
  DFF_X2 _padder__out_reg_136_  ( .D(_padder__n1680 ), .CK(clk), .Q(
        padder_out[176]), .QN() );
  DFF_X2 _padder__out_reg_104_  ( .D(_padder__n1712 ), .CK(clk), .Q(
        padder_out[80]), .QN() );
  DFF_X2 _padder__out_reg_72_  ( .D(_padder__n1744 ), .CK(clk), .Q(
        padder_out[112]), .QN() );
  DFF_X2 _padder__out_reg_40_  ( .D(_padder__n1776 ), .CK(clk), .Q(
        padder_out[16]), .QN() );
  DFF_X2 _padder__out_reg_8_  ( .D(_padder__n2449 ), .CK(clk), .Q(
        padder_out[48]), .QN() );
  DFF_X2 _padder__out_reg_521_  ( .D(_padder__n1295 ), .CK(clk), .Q(
        padder_out[561]), .QN() );
  DFF_X2 _padder__out_reg_489_  ( .D(_padder__n1327 ), .CK(clk), .Q(
        padder_out[465]), .QN() );
  DFF_X2 _padder__out_reg_457_  ( .D(_padder__n1359 ), .CK(clk), .Q(
        padder_out[497]), .QN() );
  DFF_X2 _padder__out_reg_425_  ( .D(_padder__n1391 ), .CK(clk), .Q(
        padder_out[401]), .QN() );
  DFF_X2 _padder__out_reg_393_  ( .D(_padder__n1423 ), .CK(clk), .Q(
        padder_out[433]), .QN() );
  DFF_X2 _padder__out_reg_361_  ( .D(_padder__n1455 ), .CK(clk), .Q(
        padder_out[337]), .QN() );
  DFF_X2 _padder__out_reg_329_  ( .D(_padder__n1487 ), .CK(clk), .Q(
        padder_out[369]), .QN() );
  DFF_X2 _padder__out_reg_297_  ( .D(_padder__n1519 ), .CK(clk), .Q(
        padder_out[273]), .QN() );
  DFF_X2 _padder__out_reg_265_  ( .D(_padder__n1551 ), .CK(clk), .Q(
        padder_out[305]), .QN() );
  DFF_X2 _padder__out_reg_233_  ( .D(_padder__n1583 ), .CK(clk), .Q(
        padder_out[209]), .QN() );
  DFF_X2 _padder__out_reg_201_  ( .D(_padder__n1615 ), .CK(clk), .Q(
        padder_out[241]), .QN() );
  DFF_X2 _padder__out_reg_169_  ( .D(_padder__n1647 ), .CK(clk), .Q(
        padder_out[145]), .QN() );
  DFF_X2 _padder__out_reg_137_  ( .D(_padder__n1679 ), .CK(clk), .Q(
        padder_out[177]), .QN() );
  DFF_X2 _padder__out_reg_105_  ( .D(_padder__n1711 ), .CK(clk), .Q(
        padder_out[81]), .QN() );
  DFF_X2 _padder__out_reg_73_  ( .D(_padder__n1743 ), .CK(clk), .Q(
        padder_out[113]), .QN() );
  DFF_X2 _padder__out_reg_41_  ( .D(_padder__n1775 ), .CK(clk), .Q(
        padder_out[17]), .QN() );
  DFF_X2 _padder__out_reg_9_  ( .D(_padder__n2450 ), .CK(clk), .Q(
        padder_out[49]), .QN() );
  DFF_X2 _padder__out_reg_522_  ( .D(_padder__n1294 ), .CK(clk), .Q(
        padder_out[562]), .QN() );
  DFF_X2 _padder__out_reg_490_  ( .D(_padder__n1326 ), .CK(clk), .Q(
        padder_out[466]), .QN() );
  DFF_X2 _padder__out_reg_458_  ( .D(_padder__n1358 ), .CK(clk), .Q(
        padder_out[498]), .QN() );
  DFF_X2 _padder__out_reg_426_  ( .D(_padder__n1390 ), .CK(clk), .Q(
        padder_out[402]), .QN() );
  DFF_X2 _padder__out_reg_394_  ( .D(_padder__n1422 ), .CK(clk), .Q(
        padder_out[434]), .QN() );
  DFF_X2 _padder__out_reg_362_  ( .D(_padder__n1454 ), .CK(clk), .Q(
        padder_out[338]), .QN() );
  DFF_X2 _padder__out_reg_330_  ( .D(_padder__n1486 ), .CK(clk), .Q(
        padder_out[370]), .QN() );
  DFF_X2 _padder__out_reg_298_  ( .D(_padder__n1518 ), .CK(clk), .Q(
        padder_out[274]), .QN() );
  DFF_X2 _padder__out_reg_266_  ( .D(_padder__n1550 ), .CK(clk), .Q(
        padder_out[306]), .QN() );
  DFF_X2 _padder__out_reg_234_  ( .D(_padder__n1582 ), .CK(clk), .Q(
        padder_out[210]), .QN() );
  DFF_X2 _padder__out_reg_202_  ( .D(_padder__n1614 ), .CK(clk), .Q(
        padder_out[242]), .QN() );
  DFF_X2 _padder__out_reg_170_  ( .D(_padder__n1646 ), .CK(clk), .Q(
        padder_out[146]), .QN() );
  DFF_X2 _padder__out_reg_138_  ( .D(_padder__n1678 ), .CK(clk), .Q(
        padder_out[178]), .QN() );
  DFF_X2 _padder__out_reg_106_  ( .D(_padder__n1710 ), .CK(clk), .Q(
        padder_out[82]), .QN() );
  DFF_X2 _padder__out_reg_74_  ( .D(_padder__n1742 ), .CK(clk), .Q(
        padder_out[114]), .QN() );
  DFF_X2 _padder__out_reg_42_  ( .D(_padder__n1774 ), .CK(clk), .Q(
        padder_out[18]), .QN() );
  DFF_X2 _padder__out_reg_10_  ( .D(_padder__n2451 ), .CK(clk), .Q(
        padder_out[50]), .QN() );
  DFF_X2 _padder__out_reg_523_  ( .D(_padder__n1293 ), .CK(clk), .Q(
        padder_out[563]), .QN() );
  DFF_X2 _padder__out_reg_491_  ( .D(_padder__n1325 ), .CK(clk), .Q(
        padder_out[467]), .QN() );
  DFF_X2 _padder__out_reg_459_  ( .D(_padder__n1357 ), .CK(clk), .Q(
        padder_out[499]), .QN() );
  DFF_X2 _padder__out_reg_427_  ( .D(_padder__n1389 ), .CK(clk), .Q(
        padder_out[403]), .QN() );
  DFF_X2 _padder__out_reg_395_  ( .D(_padder__n1421 ), .CK(clk), .Q(
        padder_out[435]), .QN() );
  DFF_X2 _padder__out_reg_363_  ( .D(_padder__n1453 ), .CK(clk), .Q(
        padder_out[339]), .QN() );
  DFF_X2 _padder__out_reg_331_  ( .D(_padder__n1485 ), .CK(clk), .Q(
        padder_out[371]), .QN() );
  DFF_X2 _padder__out_reg_299_  ( .D(_padder__n1517 ), .CK(clk), .Q(
        padder_out[275]), .QN() );
  DFF_X2 _padder__out_reg_267_  ( .D(_padder__n1549 ), .CK(clk), .Q(
        padder_out[307]), .QN() );
  DFF_X2 _padder__out_reg_235_  ( .D(_padder__n1581 ), .CK(clk), .Q(
        padder_out[211]), .QN() );
  DFF_X2 _padder__out_reg_203_  ( .D(_padder__n1613 ), .CK(clk), .Q(
        padder_out[243]), .QN() );
  DFF_X2 _padder__out_reg_171_  ( .D(_padder__n1645 ), .CK(clk), .Q(
        padder_out[147]), .QN() );
  DFF_X2 _padder__out_reg_139_  ( .D(_padder__n1677 ), .CK(clk), .Q(
        padder_out[179]), .QN() );
  DFF_X2 _padder__out_reg_107_  ( .D(_padder__n1709 ), .CK(clk), .Q(
        padder_out[83]), .QN() );
  DFF_X2 _padder__out_reg_75_  ( .D(_padder__n1741 ), .CK(clk), .Q(
        padder_out[115]), .QN() );
  DFF_X2 _padder__out_reg_43_  ( .D(_padder__n1773 ), .CK(clk), .Q(
        padder_out[19]), .QN() );
  DFF_X2 _padder__out_reg_11_  ( .D(_padder__n2452 ), .CK(clk), .Q(
        padder_out[51]), .QN() );
  DFF_X2 _padder__out_reg_492_  ( .D(_padder__n1324 ), .CK(clk), .Q(
        padder_out[468]), .QN() );
  DFF_X2 _padder__out_reg_460_  ( .D(_padder__n1356 ), .CK(clk), .Q(
        padder_out[500]), .QN() );
  DFF_X2 _padder__out_reg_428_  ( .D(_padder__n1388 ), .CK(clk), .Q(
        padder_out[404]), .QN() );
  DFF_X2 _padder__out_reg_396_  ( .D(_padder__n1420 ), .CK(clk), .Q(
        padder_out[436]), .QN() );
  DFF_X2 _padder__out_reg_364_  ( .D(_padder__n1452 ), .CK(clk), .Q(
        padder_out[340]), .QN() );
  DFF_X2 _padder__out_reg_332_  ( .D(_padder__n1484 ), .CK(clk), .Q(
        padder_out[372]), .QN() );
  DFF_X2 _padder__out_reg_300_  ( .D(_padder__n1516 ), .CK(clk), .Q(
        padder_out[276]), .QN() );
  DFF_X2 _padder__out_reg_268_  ( .D(_padder__n1548 ), .CK(clk), .Q(
        padder_out[308]), .QN() );
  DFF_X2 _padder__out_reg_236_  ( .D(_padder__n1580 ), .CK(clk), .Q(
        padder_out[212]), .QN() );
  DFF_X2 _padder__out_reg_204_  ( .D(_padder__n1612 ), .CK(clk), .Q(
        padder_out[244]), .QN() );
  DFF_X2 _padder__out_reg_172_  ( .D(_padder__n1644 ), .CK(clk), .Q(
        padder_out[148]), .QN() );
  DFF_X2 _padder__out_reg_140_  ( .D(_padder__n1676 ), .CK(clk), .Q(
        padder_out[180]), .QN() );
  DFF_X2 _padder__out_reg_108_  ( .D(_padder__n1708 ), .CK(clk), .Q(
        padder_out[84]), .QN() );
  DFF_X2 _padder__out_reg_76_  ( .D(_padder__n1740 ), .CK(clk), .Q(
        padder_out[116]), .QN() );
  DFF_X2 _padder__out_reg_44_  ( .D(_padder__n1772 ), .CK(clk), .Q(
        padder_out[20]), .QN() );
  DFF_X2 _padder__out_reg_12_  ( .D(_padder__n2453 ), .CK(clk), .Q(
        padder_out[52]), .QN() );
  DFF_X2 _padder__out_reg_493_  ( .D(_padder__n1323 ), .CK(clk), .Q(
        padder_out[469]), .QN() );
  DFF_X2 _padder__out_reg_461_  ( .D(_padder__n1355 ), .CK(clk), .Q(
        padder_out[501]), .QN() );
  DFF_X2 _padder__out_reg_429_  ( .D(_padder__n1387 ), .CK(clk), .Q(
        padder_out[405]), .QN() );
  DFF_X2 _padder__out_reg_397_  ( .D(_padder__n1419 ), .CK(clk), .Q(
        padder_out[437]), .QN() );
  DFF_X2 _padder__out_reg_365_  ( .D(_padder__n1451 ), .CK(clk), .Q(
        padder_out[341]), .QN() );
  DFF_X2 _padder__out_reg_333_  ( .D(_padder__n1483 ), .CK(clk), .Q(
        padder_out[373]), .QN() );
  DFF_X2 _padder__out_reg_301_  ( .D(_padder__n1515 ), .CK(clk), .Q(
        padder_out[277]), .QN() );
  DFF_X2 _padder__out_reg_269_  ( .D(_padder__n1547 ), .CK(clk), .Q(
        padder_out[309]), .QN() );
  DFF_X2 _padder__out_reg_237_  ( .D(_padder__n1579 ), .CK(clk), .Q(
        padder_out[213]), .QN() );
  DFF_X2 _padder__out_reg_205_  ( .D(_padder__n1611 ), .CK(clk), .Q(
        padder_out[245]), .QN() );
  DFF_X2 _padder__out_reg_173_  ( .D(_padder__n1643 ), .CK(clk), .Q(
        padder_out[149]), .QN() );
  DFF_X2 _padder__out_reg_141_  ( .D(_padder__n1675 ), .CK(clk), .Q(
        padder_out[181]), .QN() );
  DFF_X2 _padder__out_reg_109_  ( .D(_padder__n1707 ), .CK(clk), .Q(
        padder_out[85]), .QN() );
  DFF_X2 _padder__out_reg_77_  ( .D(_padder__n1739 ), .CK(clk), .Q(
        padder_out[117]), .QN() );
  DFF_X2 _padder__out_reg_45_  ( .D(_padder__n1771 ), .CK(clk), .Q(
        padder_out[21]), .QN() );
  DFF_X2 _padder__out_reg_13_  ( .D(_padder__n2454 ), .CK(clk), .Q(
        padder_out[53]), .QN() );
  DFF_X2 _padder__out_reg_494_  ( .D(_padder__n1322 ), .CK(clk), .Q(
        padder_out[470]), .QN() );
  DFF_X2 _padder__out_reg_462_  ( .D(_padder__n1354 ), .CK(clk), .Q(
        padder_out[502]), .QN() );
  DFF_X2 _padder__out_reg_430_  ( .D(_padder__n1386 ), .CK(clk), .Q(
        padder_out[406]), .QN() );
  DFF_X2 _padder__out_reg_398_  ( .D(_padder__n1418 ), .CK(clk), .Q(
        padder_out[438]), .QN() );
  DFF_X2 _padder__out_reg_366_  ( .D(_padder__n1450 ), .CK(clk), .Q(
        padder_out[342]), .QN() );
  DFF_X2 _padder__out_reg_334_  ( .D(_padder__n1482 ), .CK(clk), .Q(
        padder_out[374]), .QN() );
  DFF_X2 _padder__out_reg_302_  ( .D(_padder__n1514 ), .CK(clk), .Q(
        padder_out[278]), .QN() );
  DFF_X2 _padder__out_reg_270_  ( .D(_padder__n1546 ), .CK(clk), .Q(
        padder_out[310]), .QN() );
  DFF_X2 _padder__out_reg_238_  ( .D(_padder__n1578 ), .CK(clk), .Q(
        padder_out[214]), .QN() );
  DFF_X2 _padder__out_reg_206_  ( .D(_padder__n1610 ), .CK(clk), .Q(
        padder_out[246]), .QN() );
  DFF_X2 _padder__out_reg_174_  ( .D(_padder__n1642 ), .CK(clk), .Q(
        padder_out[150]), .QN() );
  DFF_X2 _padder__out_reg_142_  ( .D(_padder__n1674 ), .CK(clk), .Q(
        padder_out[182]), .QN() );
  DFF_X2 _padder__out_reg_110_  ( .D(_padder__n1706 ), .CK(clk), .Q(
        padder_out[86]), .QN() );
  DFF_X2 _padder__out_reg_78_  ( .D(_padder__n1738 ), .CK(clk), .Q(
        padder_out[118]), .QN() );
  DFF_X2 _padder__out_reg_46_  ( .D(_padder__n1770 ), .CK(clk), .Q(
        padder_out[22]), .QN() );
  DFF_X2 _padder__out_reg_14_  ( .D(_padder__n2455 ), .CK(clk), .Q(
        padder_out[54]), .QN() );
  DFF_X2 _padder__out_reg_495_  ( .D(_padder__n1321 ), .CK(clk), .Q(
        padder_out[471]), .QN() );
  DFF_X2 _padder__out_reg_463_  ( .D(_padder__n1353 ), .CK(clk), .Q(
        padder_out[503]), .QN() );
  DFF_X2 _padder__out_reg_431_  ( .D(_padder__n1385 ), .CK(clk), .Q(
        padder_out[407]), .QN() );
  DFF_X2 _padder__out_reg_399_  ( .D(_padder__n1417 ), .CK(clk), .Q(
        padder_out[439]), .QN() );
  DFF_X2 _padder__out_reg_367_  ( .D(_padder__n1449 ), .CK(clk), .Q(
        padder_out[343]), .QN() );
  DFF_X2 _padder__out_reg_335_  ( .D(_padder__n1481 ), .CK(clk), .Q(
        padder_out[375]), .QN() );
  DFF_X2 _padder__out_reg_303_  ( .D(_padder__n1513 ), .CK(clk), .Q(
        padder_out[279]), .QN() );
  DFF_X2 _padder__out_reg_271_  ( .D(_padder__n1545 ), .CK(clk), .Q(
        padder_out[311]), .QN() );
  DFF_X2 _padder__out_reg_239_  ( .D(_padder__n1577 ), .CK(clk), .Q(
        padder_out[215]), .QN() );
  DFF_X2 _padder__out_reg_207_  ( .D(_padder__n1609 ), .CK(clk), .Q(
        padder_out[247]), .QN() );
  DFF_X2 _padder__out_reg_175_  ( .D(_padder__n1641 ), .CK(clk), .Q(
        padder_out[151]), .QN() );
  DFF_X2 _padder__out_reg_143_  ( .D(_padder__n1673 ), .CK(clk), .Q(
        padder_out[183]), .QN() );
  DFF_X2 _padder__out_reg_111_  ( .D(_padder__n1705 ), .CK(clk), .Q(
        padder_out[87]), .QN() );
  DFF_X2 _padder__out_reg_79_  ( .D(_padder__n1737 ), .CK(clk), .Q(
        padder_out[119]), .QN() );
  DFF_X2 _padder__out_reg_47_  ( .D(_padder__n1769 ), .CK(clk), .Q(
        padder_out[23]), .QN() );
  DFF_X2 _padder__out_reg_15_  ( .D(_padder__n2456 ), .CK(clk), .Q(
        padder_out[55]), .QN() );
  DFF_X2 _padder__out_reg_496_  ( .D(_padder__n1320 ), .CK(clk), .Q(
        padder_out[456]), .QN() );
  DFF_X2 _padder__out_reg_464_  ( .D(_padder__n1352 ), .CK(clk), .Q(
        padder_out[488]), .QN() );
  DFF_X2 _padder__out_reg_432_  ( .D(_padder__n1384 ), .CK(clk), .Q(
        padder_out[392]), .QN() );
  DFF_X2 _padder__out_reg_400_  ( .D(_padder__n1416 ), .CK(clk), .Q(
        padder_out[424]), .QN() );
  DFF_X2 _padder__out_reg_368_  ( .D(_padder__n1448 ), .CK(clk), .Q(
        padder_out[328]), .QN() );
  DFF_X2 _padder__out_reg_336_  ( .D(_padder__n1480 ), .CK(clk), .Q(
        padder_out[360]), .QN() );
  DFF_X2 _padder__out_reg_304_  ( .D(_padder__n1512 ), .CK(clk), .Q(
        padder_out[264]), .QN() );
  DFF_X2 _padder__out_reg_272_  ( .D(_padder__n1544 ), .CK(clk), .Q(
        padder_out[296]), .QN() );
  DFF_X2 _padder__out_reg_240_  ( .D(_padder__n1576 ), .CK(clk), .Q(
        padder_out[200]), .QN() );
  DFF_X2 _padder__out_reg_208_  ( .D(_padder__n1608 ), .CK(clk), .Q(
        padder_out[232]), .QN() );
  DFF_X2 _padder__out_reg_176_  ( .D(_padder__n1640 ), .CK(clk), .Q(
        padder_out[136]), .QN() );
  DFF_X2 _padder__out_reg_144_  ( .D(_padder__n1672 ), .CK(clk), .Q(
        padder_out[168]), .QN() );
  DFF_X2 _padder__out_reg_112_  ( .D(_padder__n1704 ), .CK(clk), .Q(
        padder_out[72]), .QN() );
  DFF_X2 _padder__out_reg_80_  ( .D(_padder__n1736 ), .CK(clk), .Q(
        padder_out[104]), .QN() );
  DFF_X2 _padder__out_reg_48_  ( .D(_padder__n1768 ), .CK(clk), .Q(
        padder_out[8]), .QN() );
  DFF_X2 _padder__out_reg_16_  ( .D(_padder__n2457 ), .CK(clk), .Q(
        padder_out[40]), .QN() );
  DFF_X2 _padder__out_reg_497_  ( .D(_padder__n1319 ), .CK(clk), .Q(
        padder_out[457]), .QN() );
  DFF_X2 _padder__out_reg_465_  ( .D(_padder__n1351 ), .CK(clk), .Q(
        padder_out[489]), .QN() );
  DFF_X2 _padder__out_reg_433_  ( .D(_padder__n1383 ), .CK(clk), .Q(
        padder_out[393]), .QN() );
  DFF_X2 _padder__out_reg_401_  ( .D(_padder__n1415 ), .CK(clk), .Q(
        padder_out[425]), .QN() );
  DFF_X2 _padder__out_reg_369_  ( .D(_padder__n1447 ), .CK(clk), .Q(
        padder_out[329]), .QN() );
  DFF_X2 _padder__out_reg_337_  ( .D(_padder__n1479 ), .CK(clk), .Q(
        padder_out[361]), .QN() );
  DFF_X2 _padder__out_reg_305_  ( .D(_padder__n1511 ), .CK(clk), .Q(
        padder_out[265]), .QN() );
  DFF_X2 _padder__out_reg_273_  ( .D(_padder__n1543 ), .CK(clk), .Q(
        padder_out[297]), .QN() );
  DFF_X2 _padder__out_reg_241_  ( .D(_padder__n1575 ), .CK(clk), .Q(
        padder_out[201]), .QN() );
  DFF_X2 _padder__out_reg_209_  ( .D(_padder__n1607 ), .CK(clk), .Q(
        padder_out[233]), .QN() );
  DFF_X2 _padder__out_reg_177_  ( .D(_padder__n1639 ), .CK(clk), .Q(
        padder_out[137]), .QN() );
  DFF_X2 _padder__out_reg_145_  ( .D(_padder__n1671 ), .CK(clk), .Q(
        padder_out[169]), .QN() );
  DFF_X2 _padder__out_reg_113_  ( .D(_padder__n1703 ), .CK(clk), .Q(
        padder_out[73]), .QN() );
  DFF_X2 _padder__out_reg_81_  ( .D(_padder__n1735 ), .CK(clk), .Q(
        padder_out[105]), .QN() );
  DFF_X2 _padder__out_reg_49_  ( .D(_padder__n1767 ), .CK(clk), .Q(
        padder_out[9]), .QN() );
  DFF_X2 _padder__out_reg_17_  ( .D(_padder__n2458 ), .CK(clk), .Q(
        padder_out[41]), .QN() );
  DFF_X2 _padder__out_reg_498_  ( .D(_padder__n1318 ), .CK(clk), .Q(
        padder_out[458]), .QN() );
  DFF_X2 _padder__out_reg_466_  ( .D(_padder__n1350 ), .CK(clk), .Q(
        padder_out[490]), .QN() );
  DFF_X2 _padder__out_reg_434_  ( .D(_padder__n1382 ), .CK(clk), .Q(
        padder_out[394]), .QN() );
  DFF_X2 _padder__out_reg_402_  ( .D(_padder__n1414 ), .CK(clk), .Q(
        padder_out[426]), .QN() );
  DFF_X2 _padder__out_reg_370_  ( .D(_padder__n1446 ), .CK(clk), .Q(
        padder_out[330]), .QN() );
  DFF_X2 _padder__out_reg_338_  ( .D(_padder__n1478 ), .CK(clk), .Q(
        padder_out[362]), .QN() );
  DFF_X2 _padder__out_reg_306_  ( .D(_padder__n1510 ), .CK(clk), .Q(
        padder_out[266]), .QN() );
  DFF_X2 _padder__out_reg_274_  ( .D(_padder__n1542 ), .CK(clk), .Q(
        padder_out[298]), .QN() );
  DFF_X2 _padder__out_reg_242_  ( .D(_padder__n1574 ), .CK(clk), .Q(
        padder_out[202]), .QN() );
  DFF_X2 _padder__out_reg_210_  ( .D(_padder__n1606 ), .CK(clk), .Q(
        padder_out[234]), .QN() );
  DFF_X2 _padder__out_reg_178_  ( .D(_padder__n1638 ), .CK(clk), .Q(
        padder_out[138]), .QN() );
  DFF_X2 _padder__out_reg_146_  ( .D(_padder__n1670 ), .CK(clk), .Q(
        padder_out[170]), .QN() );
  DFF_X2 _padder__out_reg_114_  ( .D(_padder__n1702 ), .CK(clk), .Q(
        padder_out[74]), .QN() );
  DFF_X2 _padder__out_reg_82_  ( .D(_padder__n1734 ), .CK(clk), .Q(
        padder_out[106]), .QN() );
  DFF_X2 _padder__out_reg_50_  ( .D(_padder__n1766 ), .CK(clk), .Q(
        padder_out[10]), .QN() );
  DFF_X2 _padder__out_reg_18_  ( .D(_padder__n2459 ), .CK(clk), .Q(
        padder_out[42]), .QN() );
  DFF_X2 _padder__out_reg_499_  ( .D(_padder__n1317 ), .CK(clk), .Q(
        padder_out[459]), .QN() );
  DFF_X2 _padder__out_reg_467_  ( .D(_padder__n1349 ), .CK(clk), .Q(
        padder_out[491]), .QN() );
  DFF_X2 _padder__out_reg_435_  ( .D(_padder__n1381 ), .CK(clk), .Q(
        padder_out[395]), .QN() );
  DFF_X2 _padder__out_reg_403_  ( .D(_padder__n1413 ), .CK(clk), .Q(
        padder_out[427]), .QN() );
  DFF_X2 _padder__out_reg_371_  ( .D(_padder__n1445 ), .CK(clk), .Q(
        padder_out[331]), .QN() );
  DFF_X2 _padder__out_reg_339_  ( .D(_padder__n1477 ), .CK(clk), .Q(
        padder_out[363]), .QN() );
  DFF_X2 _padder__out_reg_307_  ( .D(_padder__n1509 ), .CK(clk), .Q(
        padder_out[267]), .QN() );
  DFF_X2 _padder__out_reg_275_  ( .D(_padder__n1541 ), .CK(clk), .Q(
        padder_out[299]), .QN() );
  DFF_X2 _padder__out_reg_243_  ( .D(_padder__n1573 ), .CK(clk), .Q(
        padder_out[203]), .QN() );
  DFF_X2 _padder__out_reg_211_  ( .D(_padder__n1605 ), .CK(clk), .Q(
        padder_out[235]), .QN() );
  DFF_X2 _padder__out_reg_179_  ( .D(_padder__n1637 ), .CK(clk), .Q(
        padder_out[139]), .QN() );
  DFF_X2 _padder__out_reg_147_  ( .D(_padder__n1669 ), .CK(clk), .Q(
        padder_out[171]), .QN() );
  DFF_X2 _padder__out_reg_115_  ( .D(_padder__n1701 ), .CK(clk), .Q(
        padder_out[75]), .QN() );
  DFF_X2 _padder__out_reg_83_  ( .D(_padder__n1733 ), .CK(clk), .Q(
        padder_out[107]), .QN() );
  DFF_X2 _padder__out_reg_51_  ( .D(_padder__n1765 ), .CK(clk), .Q(
        padder_out[11]), .QN() );
  DFF_X2 _padder__out_reg_19_  ( .D(_padder__n2460 ), .CK(clk), .Q(
        padder_out[43]), .QN() );
  DFF_X2 _padder__out_reg_500_  ( .D(_padder__n1316 ), .CK(clk), .Q(
        padder_out[460]), .QN() );
  DFF_X2 _padder__out_reg_468_  ( .D(_padder__n1348 ), .CK(clk), .Q(
        padder_out[492]), .QN() );
  DFF_X2 _padder__out_reg_436_  ( .D(_padder__n1380 ), .CK(clk), .Q(
        padder_out[396]), .QN() );
  DFF_X2 _padder__out_reg_404_  ( .D(_padder__n1412 ), .CK(clk), .Q(
        padder_out[428]), .QN() );
  DFF_X2 _padder__out_reg_372_  ( .D(_padder__n1444 ), .CK(clk), .Q(
        padder_out[332]), .QN() );
  DFF_X2 _padder__out_reg_340_  ( .D(_padder__n1476 ), .CK(clk), .Q(
        padder_out[364]), .QN() );
  DFF_X2 _padder__out_reg_308_  ( .D(_padder__n1508 ), .CK(clk), .Q(
        padder_out[268]), .QN() );
  DFF_X2 _padder__out_reg_276_  ( .D(_padder__n1540 ), .CK(clk), .Q(
        padder_out[300]), .QN() );
  DFF_X2 _padder__out_reg_244_  ( .D(_padder__n1572 ), .CK(clk), .Q(
        padder_out[204]), .QN() );
  DFF_X2 _padder__out_reg_212_  ( .D(_padder__n1604 ), .CK(clk), .Q(
        padder_out[236]), .QN() );
  DFF_X2 _padder__out_reg_180_  ( .D(_padder__n1636 ), .CK(clk), .Q(
        padder_out[140]), .QN() );
  DFF_X2 _padder__out_reg_148_  ( .D(_padder__n1668 ), .CK(clk), .Q(
        padder_out[172]), .QN() );
  DFF_X2 _padder__out_reg_116_  ( .D(_padder__n1700 ), .CK(clk), .Q(
        padder_out[76]), .QN() );
  DFF_X2 _padder__out_reg_84_  ( .D(_padder__n1732 ), .CK(clk), .Q(
        padder_out[108]), .QN() );
  DFF_X2 _padder__out_reg_52_  ( .D(_padder__n1764 ), .CK(clk), .Q(
        padder_out[12]), .QN() );
  DFF_X2 _padder__out_reg_20_  ( .D(_padder__n2461 ), .CK(clk), .Q(
        padder_out[44]), .QN() );
  DFF_X2 _padder__out_reg_501_  ( .D(_padder__n1315 ), .CK(clk), .Q(
        padder_out[461]), .QN() );
  DFF_X2 _padder__out_reg_469_  ( .D(_padder__n1347 ), .CK(clk), .Q(
        padder_out[493]), .QN() );
  DFF_X2 _padder__out_reg_437_  ( .D(_padder__n1379 ), .CK(clk), .Q(
        padder_out[397]), .QN() );
  DFF_X2 _padder__out_reg_405_  ( .D(_padder__n1411 ), .CK(clk), .Q(
        padder_out[429]), .QN() );
  DFF_X2 _padder__out_reg_373_  ( .D(_padder__n1443 ), .CK(clk), .Q(
        padder_out[333]), .QN() );
  DFF_X2 _padder__out_reg_341_  ( .D(_padder__n1475 ), .CK(clk), .Q(
        padder_out[365]), .QN() );
  DFF_X2 _padder__out_reg_309_  ( .D(_padder__n1507 ), .CK(clk), .Q(
        padder_out[269]), .QN() );
  DFF_X2 _padder__out_reg_277_  ( .D(_padder__n1539 ), .CK(clk), .Q(
        padder_out[301]), .QN() );
  DFF_X2 _padder__out_reg_245_  ( .D(_padder__n1571 ), .CK(clk), .Q(
        padder_out[205]), .QN() );
  DFF_X2 _padder__out_reg_213_  ( .D(_padder__n1603 ), .CK(clk), .Q(
        padder_out[237]), .QN() );
  DFF_X2 _padder__out_reg_181_  ( .D(_padder__n1635 ), .CK(clk), .Q(
        padder_out[141]), .QN() );
  DFF_X2 _padder__out_reg_149_  ( .D(_padder__n1667 ), .CK(clk), .Q(
        padder_out[173]), .QN() );
  DFF_X2 _padder__out_reg_117_  ( .D(_padder__n1699 ), .CK(clk), .Q(
        padder_out[77]), .QN() );
  DFF_X2 _padder__out_reg_85_  ( .D(_padder__n1731 ), .CK(clk), .Q(
        padder_out[109]), .QN() );
  DFF_X2 _padder__out_reg_53_  ( .D(_padder__n1763 ), .CK(clk), .Q(
        padder_out[13]), .QN() );
  DFF_X2 _padder__out_reg_21_  ( .D(_padder__n2462 ), .CK(clk), .Q(
        padder_out[45]), .QN() );
  DFF_X2 _padder__out_reg_502_  ( .D(_padder__n1314 ), .CK(clk), .Q(
        padder_out[462]), .QN() );
  DFF_X2 _padder__out_reg_470_  ( .D(_padder__n1346 ), .CK(clk), .Q(
        padder_out[494]), .QN() );
  DFF_X2 _padder__out_reg_438_  ( .D(_padder__n1378 ), .CK(clk), .Q(
        padder_out[398]), .QN() );
  DFF_X2 _padder__out_reg_406_  ( .D(_padder__n1410 ), .CK(clk), .Q(
        padder_out[430]), .QN() );
  DFF_X2 _padder__out_reg_374_  ( .D(_padder__n1442 ), .CK(clk), .Q(
        padder_out[334]), .QN() );
  DFF_X2 _padder__out_reg_342_  ( .D(_padder__n1474 ), .CK(clk), .Q(
        padder_out[366]), .QN() );
  DFF_X2 _padder__out_reg_310_  ( .D(_padder__n1506 ), .CK(clk), .Q(
        padder_out[270]), .QN() );
  DFF_X2 _padder__out_reg_278_  ( .D(_padder__n1538 ), .CK(clk), .Q(
        padder_out[302]), .QN() );
  DFF_X2 _padder__out_reg_246_  ( .D(_padder__n1570 ), .CK(clk), .Q(
        padder_out[206]), .QN() );
  DFF_X2 _padder__out_reg_214_  ( .D(_padder__n1602 ), .CK(clk), .Q(
        padder_out[238]), .QN() );
  DFF_X2 _padder__out_reg_182_  ( .D(_padder__n1634 ), .CK(clk), .Q(
        padder_out[142]), .QN() );
  DFF_X2 _padder__out_reg_150_  ( .D(_padder__n1666 ), .CK(clk), .Q(
        padder_out[174]), .QN() );
  DFF_X2 _padder__out_reg_118_  ( .D(_padder__n1698 ), .CK(clk), .Q(
        padder_out[78]), .QN() );
  DFF_X2 _padder__out_reg_86_  ( .D(_padder__n1730 ), .CK(clk), .Q(
        padder_out[110]), .QN() );
  DFF_X2 _padder__out_reg_54_  ( .D(_padder__n1762 ), .CK(clk), .Q(
        padder_out[14]), .QN() );
  DFF_X2 _padder__out_reg_22_  ( .D(_padder__n2463 ), .CK(clk), .Q(
        padder_out[46]), .QN() );
  DFF_X2 _padder__out_reg_503_  ( .D(_padder__n1313 ), .CK(clk), .Q(
        padder_out[463]), .QN() );
  DFF_X2 _padder__out_reg_471_  ( .D(_padder__n1345 ), .CK(clk), .Q(
        padder_out[495]), .QN() );
  DFF_X2 _padder__out_reg_439_  ( .D(_padder__n1377 ), .CK(clk), .Q(
        padder_out[399]), .QN() );
  DFF_X2 _padder__out_reg_407_  ( .D(_padder__n1409 ), .CK(clk), .Q(
        padder_out[431]), .QN() );
  DFF_X2 _padder__out_reg_375_  ( .D(_padder__n1441 ), .CK(clk), .Q(
        padder_out[335]), .QN() );
  DFF_X2 _padder__out_reg_343_  ( .D(_padder__n1473 ), .CK(clk), .Q(
        padder_out[367]), .QN() );
  DFF_X2 _padder__out_reg_311_  ( .D(_padder__n1505 ), .CK(clk), .Q(
        padder_out[271]), .QN() );
  DFF_X2 _padder__out_reg_279_  ( .D(_padder__n1537 ), .CK(clk), .Q(
        padder_out[303]), .QN() );
  DFF_X2 _padder__out_reg_247_  ( .D(_padder__n1569 ), .CK(clk), .Q(
        padder_out[207]), .QN() );
  DFF_X2 _padder__out_reg_215_  ( .D(_padder__n1601 ), .CK(clk), .Q(
        padder_out[239]), .QN() );
  DFF_X2 _padder__out_reg_183_  ( .D(_padder__n1633 ), .CK(clk), .Q(
        padder_out[143]), .QN() );
  DFF_X2 _padder__out_reg_151_  ( .D(_padder__n1665 ), .CK(clk), .Q(
        padder_out[175]), .QN() );
  DFF_X2 _padder__out_reg_119_  ( .D(_padder__n1697 ), .CK(clk), .Q(
        padder_out[79]), .QN() );
  DFF_X2 _padder__out_reg_87_  ( .D(_padder__n1729 ), .CK(clk), .Q(
        padder_out[111]), .QN() );
  DFF_X2 _padder__out_reg_55_  ( .D(_padder__n1761 ), .CK(clk), .Q(
        padder_out[15]), .QN() );
  DFF_X2 _padder__out_reg_23_  ( .D(_padder__n2464 ), .CK(clk), .Q(
        padder_out[47]), .QN() );
  DFF_X2 _padder__out_reg_504_  ( .D(_padder__n1312 ), .CK(clk), .Q(
        padder_out[448]), .QN() );
  DFF_X2 _padder__out_reg_472_  ( .D(_padder__n1344 ), .CK(clk), .Q(
        padder_out[480]), .QN() );
  DFF_X2 _padder__out_reg_440_  ( .D(_padder__n1376 ), .CK(clk), .Q(
        padder_out[384]), .QN() );
  DFF_X2 _padder__out_reg_408_  ( .D(_padder__n1408 ), .CK(clk), .Q(
        padder_out[416]), .QN() );
  DFF_X2 _padder__out_reg_376_  ( .D(_padder__n1440 ), .CK(clk), .Q(
        padder_out[320]), .QN() );
  DFF_X2 _padder__out_reg_344_  ( .D(_padder__n1472 ), .CK(clk), .Q(
        padder_out[352]), .QN() );
  DFF_X2 _padder__out_reg_312_  ( .D(_padder__n1504 ), .CK(clk), .Q(
        padder_out[256]), .QN() );
  DFF_X2 _padder__out_reg_280_  ( .D(_padder__n1536 ), .CK(clk), .Q(
        padder_out[288]), .QN() );
  DFF_X2 _padder__out_reg_248_  ( .D(_padder__n1568 ), .CK(clk), .Q(
        padder_out[192]), .QN() );
  DFF_X2 _padder__out_reg_216_  ( .D(_padder__n1600 ), .CK(clk), .Q(
        padder_out[224]), .QN() );
  DFF_X2 _padder__out_reg_184_  ( .D(_padder__n1632 ), .CK(clk), .Q(
        padder_out[128]), .QN() );
  DFF_X2 _padder__out_reg_152_  ( .D(_padder__n1664 ), .CK(clk), .Q(
        padder_out[160]), .QN() );
  DFF_X2 _padder__out_reg_120_  ( .D(_padder__n1696 ), .CK(clk), .Q(
        padder_out[64]), .QN() );
  DFF_X2 _padder__out_reg_88_  ( .D(_padder__n1728 ), .CK(clk), .Q(
        padder_out[96]), .QN() );
  DFF_X2 _padder__out_reg_56_  ( .D(_padder__n1760 ), .CK(clk), .Q(
        padder_out[0]), .QN() );
  DFF_X2 _padder__out_reg_24_  ( .D(_padder__n2465 ), .CK(clk), .Q(
        padder_out[32]), .QN() );
  DFF_X2 _padder__out_reg_505_  ( .D(_padder__n1311 ), .CK(clk), .Q(
        padder_out[449]), .QN() );
  DFF_X2 _padder__out_reg_473_  ( .D(_padder__n1343 ), .CK(clk), .Q(
        padder_out[481]), .QN() );
  DFF_X2 _padder__out_reg_441_  ( .D(_padder__n1375 ), .CK(clk), .Q(
        padder_out[385]), .QN() );
  DFF_X2 _padder__out_reg_409_  ( .D(_padder__n1407 ), .CK(clk), .Q(
        padder_out[417]), .QN() );
  DFF_X2 _padder__out_reg_377_  ( .D(_padder__n1439 ), .CK(clk), .Q(
        padder_out[321]), .QN() );
  DFF_X2 _padder__out_reg_345_  ( .D(_padder__n1471 ), .CK(clk), .Q(
        padder_out[353]), .QN() );
  DFF_X2 _padder__out_reg_313_  ( .D(_padder__n1503 ), .CK(clk), .Q(
        padder_out[257]), .QN() );
  DFF_X2 _padder__out_reg_281_  ( .D(_padder__n1535 ), .CK(clk), .Q(
        padder_out[289]), .QN() );
  DFF_X2 _padder__out_reg_249_  ( .D(_padder__n1567 ), .CK(clk), .Q(
        padder_out[193]), .QN() );
  DFF_X2 _padder__out_reg_217_  ( .D(_padder__n1599 ), .CK(clk), .Q(
        padder_out[225]), .QN() );
  DFF_X2 _padder__out_reg_185_  ( .D(_padder__n1631 ), .CK(clk), .Q(
        padder_out[129]), .QN() );
  DFF_X2 _padder__out_reg_153_  ( .D(_padder__n1663 ), .CK(clk), .Q(
        padder_out[161]), .QN() );
  DFF_X2 _padder__out_reg_121_  ( .D(_padder__n1695 ), .CK(clk), .Q(
        padder_out[65]), .QN() );
  DFF_X2 _padder__out_reg_89_  ( .D(_padder__n1727 ), .CK(clk), .Q(
        padder_out[97]), .QN() );
  DFF_X2 _padder__out_reg_57_  ( .D(_padder__n1759 ), .CK(clk), .Q(
        padder_out[1]), .QN() );
  DFF_X2 _padder__out_reg_25_  ( .D(_padder__n2466 ), .CK(clk), .Q(
        padder_out[33]), .QN() );
  DFF_X2 _padder__out_reg_506_  ( .D(_padder__n1310 ), .CK(clk), .Q(
        padder_out[450]), .QN() );
  DFF_X2 _padder__out_reg_474_  ( .D(_padder__n1342 ), .CK(clk), .Q(
        padder_out[482]), .QN() );
  DFF_X2 _padder__out_reg_442_  ( .D(_padder__n1374 ), .CK(clk), .Q(
        padder_out[386]), .QN() );
  DFF_X2 _padder__out_reg_410_  ( .D(_padder__n1406 ), .CK(clk), .Q(
        padder_out[418]), .QN() );
  DFF_X2 _padder__out_reg_378_  ( .D(_padder__n1438 ), .CK(clk), .Q(
        padder_out[322]), .QN() );
  DFF_X2 _padder__out_reg_346_  ( .D(_padder__n1470 ), .CK(clk), .Q(
        padder_out[354]), .QN() );
  DFF_X2 _padder__out_reg_314_  ( .D(_padder__n1502 ), .CK(clk), .Q(
        padder_out[258]), .QN() );
  DFF_X2 _padder__out_reg_282_  ( .D(_padder__n1534 ), .CK(clk), .Q(
        padder_out[290]), .QN() );
  DFF_X2 _padder__out_reg_250_  ( .D(_padder__n1566 ), .CK(clk), .Q(
        padder_out[194]), .QN() );
  DFF_X2 _padder__out_reg_218_  ( .D(_padder__n1598 ), .CK(clk), .Q(
        padder_out[226]), .QN() );
  DFF_X2 _padder__out_reg_186_  ( .D(_padder__n1630 ), .CK(clk), .Q(
        padder_out[130]), .QN() );
  DFF_X2 _padder__out_reg_154_  ( .D(_padder__n1662 ), .CK(clk), .Q(
        padder_out[162]), .QN() );
  DFF_X2 _padder__out_reg_122_  ( .D(_padder__n1694 ), .CK(clk), .Q(
        padder_out[66]), .QN() );
  DFF_X2 _padder__out_reg_90_  ( .D(_padder__n1726 ), .CK(clk), .Q(
        padder_out[98]), .QN() );
  DFF_X2 _padder__out_reg_58_  ( .D(_padder__n1758 ), .CK(clk), .Q(
        padder_out[2]), .QN() );
  DFF_X2 _padder__out_reg_26_  ( .D(_padder__n2467 ), .CK(clk), .Q(
        padder_out[34]), .QN() );
  DFF_X2 _padder__out_reg_507_  ( .D(_padder__n1309 ), .CK(clk), .Q(
        padder_out[451]), .QN() );
  DFF_X2 _padder__out_reg_475_  ( .D(_padder__n1341 ), .CK(clk), .Q(
        padder_out[483]), .QN() );
  DFF_X2 _padder__out_reg_443_  ( .D(_padder__n1373 ), .CK(clk), .Q(
        padder_out[387]), .QN() );
  DFF_X2 _padder__out_reg_411_  ( .D(_padder__n1405 ), .CK(clk), .Q(
        padder_out[419]), .QN() );
  DFF_X2 _padder__out_reg_379_  ( .D(_padder__n1437 ), .CK(clk), .Q(
        padder_out[323]), .QN() );
  DFF_X2 _padder__out_reg_347_  ( .D(_padder__n1469 ), .CK(clk), .Q(
        padder_out[355]), .QN() );
  DFF_X2 _padder__out_reg_315_  ( .D(_padder__n1501 ), .CK(clk), .Q(
        padder_out[259]), .QN() );
  DFF_X2 _padder__out_reg_283_  ( .D(_padder__n1533 ), .CK(clk), .Q(
        padder_out[291]), .QN() );
  DFF_X2 _padder__out_reg_251_  ( .D(_padder__n1565 ), .CK(clk), .Q(
        padder_out[195]), .QN() );
  DFF_X2 _padder__out_reg_219_  ( .D(_padder__n1597 ), .CK(clk), .Q(
        padder_out[227]), .QN() );
  DFF_X2 _padder__out_reg_187_  ( .D(_padder__n1629 ), .CK(clk), .Q(
        padder_out[131]), .QN() );
  DFF_X2 _padder__out_reg_155_  ( .D(_padder__n1661 ), .CK(clk), .Q(
        padder_out[163]), .QN() );
  DFF_X2 _padder__out_reg_123_  ( .D(_padder__n1693 ), .CK(clk), .Q(
        padder_out[67]), .QN() );
  DFF_X2 _padder__out_reg_91_  ( .D(_padder__n1725 ), .CK(clk), .Q(
        padder_out[99]), .QN() );
  DFF_X2 _padder__out_reg_59_  ( .D(_padder__n1757 ), .CK(clk), .Q(
        padder_out[3]), .QN() );
  DFF_X2 _padder__out_reg_27_  ( .D(_padder__n2468 ), .CK(clk), .Q(
        padder_out[35]), .QN() );
  DFF_X2 _padder__out_reg_508_  ( .D(_padder__n1308 ), .CK(clk), .Q(
        padder_out[452]), .QN() );
  DFF_X2 _padder__out_reg_476_  ( .D(_padder__n1340 ), .CK(clk), .Q(
        padder_out[484]), .QN() );
  DFF_X2 _padder__out_reg_444_  ( .D(_padder__n1372 ), .CK(clk), .Q(
        padder_out[388]), .QN() );
  DFF_X2 _padder__out_reg_412_  ( .D(_padder__n1404 ), .CK(clk), .Q(
        padder_out[420]), .QN() );
  DFF_X2 _padder__out_reg_380_  ( .D(_padder__n1436 ), .CK(clk), .Q(
        padder_out[324]), .QN() );
  DFF_X2 _padder__out_reg_348_  ( .D(_padder__n1468 ), .CK(clk), .Q(
        padder_out[356]), .QN() );
  DFF_X2 _padder__out_reg_316_  ( .D(_padder__n1500 ), .CK(clk), .Q(
        padder_out[260]), .QN() );
  DFF_X2 _padder__out_reg_284_  ( .D(_padder__n1532 ), .CK(clk), .Q(
        padder_out[292]), .QN() );
  DFF_X2 _padder__out_reg_252_  ( .D(_padder__n1564 ), .CK(clk), .Q(
        padder_out[196]), .QN() );
  DFF_X2 _padder__out_reg_220_  ( .D(_padder__n1596 ), .CK(clk), .Q(
        padder_out[228]), .QN() );
  DFF_X2 _padder__out_reg_188_  ( .D(_padder__n1628 ), .CK(clk), .Q(
        padder_out[132]), .QN() );
  DFF_X2 _padder__out_reg_156_  ( .D(_padder__n1660 ), .CK(clk), .Q(
        padder_out[164]), .QN() );
  DFF_X2 _padder__out_reg_124_  ( .D(_padder__n1692 ), .CK(clk), .Q(
        padder_out[68]), .QN() );
  DFF_X2 _padder__out_reg_92_  ( .D(_padder__n1724 ), .CK(clk), .Q(
        padder_out[100]), .QN() );
  DFF_X2 _padder__out_reg_60_  ( .D(_padder__n1756 ), .CK(clk), .Q(
        padder_out[4]), .QN() );
  DFF_X2 _padder__out_reg_28_  ( .D(_padder__n2469 ), .CK(clk), .Q(
        padder_out[36]), .QN() );
  DFF_X2 _padder__out_reg_509_  ( .D(_padder__n1307 ), .CK(clk), .Q(
        padder_out[453]), .QN() );
  DFF_X2 _padder__out_reg_477_  ( .D(_padder__n1339 ), .CK(clk), .Q(
        padder_out[485]), .QN() );
  DFF_X2 _padder__out_reg_445_  ( .D(_padder__n1371 ), .CK(clk), .Q(
        padder_out[389]), .QN() );
  DFF_X2 _padder__out_reg_413_  ( .D(_padder__n1403 ), .CK(clk), .Q(
        padder_out[421]), .QN() );
  DFF_X2 _padder__out_reg_381_  ( .D(_padder__n1435 ), .CK(clk), .Q(
        padder_out[325]), .QN() );
  DFF_X2 _padder__out_reg_349_  ( .D(_padder__n1467 ), .CK(clk), .Q(
        padder_out[357]), .QN() );
  DFF_X2 _padder__out_reg_317_  ( .D(_padder__n1499 ), .CK(clk), .Q(
        padder_out[261]), .QN() );
  DFF_X2 _padder__out_reg_285_  ( .D(_padder__n1531 ), .CK(clk), .Q(
        padder_out[293]), .QN() );
  DFF_X2 _padder__out_reg_253_  ( .D(_padder__n1563 ), .CK(clk), .Q(
        padder_out[197]), .QN() );
  DFF_X2 _padder__out_reg_221_  ( .D(_padder__n1595 ), .CK(clk), .Q(
        padder_out[229]), .QN() );
  DFF_X2 _padder__out_reg_189_  ( .D(_padder__n1627 ), .CK(clk), .Q(
        padder_out[133]), .QN() );
  DFF_X2 _padder__out_reg_157_  ( .D(_padder__n1659 ), .CK(clk), .Q(
        padder_out[165]), .QN() );
  DFF_X2 _padder__out_reg_125_  ( .D(_padder__n1691 ), .CK(clk), .Q(
        padder_out[69]), .QN() );
  DFF_X2 _padder__out_reg_93_  ( .D(_padder__n1723 ), .CK(clk), .Q(
        padder_out[101]), .QN() );
  DFF_X2 _padder__out_reg_61_  ( .D(_padder__n1755 ), .CK(clk), .Q(
        padder_out[5]), .QN() );
  DFF_X2 _padder__out_reg_29_  ( .D(_padder__n2470 ), .CK(clk), .Q(
        padder_out[37]), .QN() );
  DFF_X2 _padder__out_reg_510_  ( .D(_padder__n1306 ), .CK(clk), .Q(
        padder_out[454]), .QN() );
  DFF_X2 _padder__out_reg_478_  ( .D(_padder__n1338 ), .CK(clk), .Q(
        padder_out[486]), .QN() );
  DFF_X2 _padder__out_reg_446_  ( .D(_padder__n1370 ), .CK(clk), .Q(
        padder_out[390]), .QN() );
  DFF_X2 _padder__out_reg_414_  ( .D(_padder__n1402 ), .CK(clk), .Q(
        padder_out[422]), .QN() );
  DFF_X2 _padder__out_reg_382_  ( .D(_padder__n1434 ), .CK(clk), .Q(
        padder_out[326]), .QN() );
  DFF_X2 _padder__out_reg_350_  ( .D(_padder__n1466 ), .CK(clk), .Q(
        padder_out[358]), .QN() );
  DFF_X2 _padder__out_reg_318_  ( .D(_padder__n1498 ), .CK(clk), .Q(
        padder_out[262]), .QN() );
  DFF_X2 _padder__out_reg_286_  ( .D(_padder__n1530 ), .CK(clk), .Q(
        padder_out[294]), .QN() );
  DFF_X2 _padder__out_reg_254_  ( .D(_padder__n1562 ), .CK(clk), .Q(
        padder_out[198]), .QN() );
  DFF_X2 _padder__out_reg_222_  ( .D(_padder__n1594 ), .CK(clk), .Q(
        padder_out[230]), .QN() );
  DFF_X2 _padder__out_reg_190_  ( .D(_padder__n1626 ), .CK(clk), .Q(
        padder_out[134]), .QN() );
  DFF_X2 _padder__out_reg_158_  ( .D(_padder__n1658 ), .CK(clk), .Q(
        padder_out[166]), .QN() );
  DFF_X2 _padder__out_reg_126_  ( .D(_padder__n1690 ), .CK(clk), .Q(
        padder_out[70]), .QN() );
  DFF_X2 _padder__out_reg_94_  ( .D(_padder__n1722 ), .CK(clk), .Q(
        padder_out[102]), .QN() );
  DFF_X2 _padder__out_reg_62_  ( .D(_padder__n1754 ), .CK(clk), .Q(
        padder_out[6]), .QN() );
  DFF_X2 _padder__out_reg_30_  ( .D(_padder__n2471 ), .CK(clk), .Q(
        padder_out[38]), .QN() );
  DFF_X2 _padder__out_reg_511_  ( .D(_padder__n1305 ), .CK(clk), .Q(
        padder_out[455]), .QN() );
  DFF_X2 _padder__out_reg_479_  ( .D(_padder__n1337 ), .CK(clk), .Q(
        padder_out[487]), .QN() );
  DFF_X2 _padder__out_reg_447_  ( .D(_padder__n1369 ), .CK(clk), .Q(
        padder_out[391]), .QN() );
  DFF_X2 _padder__out_reg_415_  ( .D(_padder__n1401 ), .CK(clk), .Q(
        padder_out[423]), .QN() );
  DFF_X2 _padder__out_reg_383_  ( .D(_padder__n1433 ), .CK(clk), .Q(
        padder_out[327]), .QN() );
  DFF_X2 _padder__out_reg_351_  ( .D(_padder__n1465 ), .CK(clk), .Q(
        padder_out[359]), .QN() );
  DFF_X2 _padder__out_reg_319_  ( .D(_padder__n1497 ), .CK(clk), .Q(
        padder_out[263]), .QN() );
  DFF_X2 _padder__out_reg_287_  ( .D(_padder__n1529 ), .CK(clk), .Q(
        padder_out[295]), .QN() );
  DFF_X2 _padder__out_reg_255_  ( .D(_padder__n1561 ), .CK(clk), .Q(
        padder_out[199]), .QN() );
  DFF_X2 _padder__out_reg_223_  ( .D(_padder__n1593 ), .CK(clk), .Q(
        padder_out[231]), .QN() );
  DFF_X2 _padder__out_reg_191_  ( .D(_padder__n1625 ), .CK(clk), .Q(
        padder_out[135]), .QN() );
  DFF_X2 _padder__out_reg_159_  ( .D(_padder__n1657 ), .CK(clk), .Q(
        padder_out[167]), .QN() );
  DFF_X2 _padder__out_reg_127_  ( .D(_padder__n1689 ), .CK(clk), .Q(
        padder_out[71]), .QN() );
  DFF_X2 _padder__out_reg_95_  ( .D(_padder__n1721 ), .CK(clk), .Q(
        padder_out[103]), .QN() );
  DFF_X2 _padder__out_reg_63_  ( .D(_padder__n1753 ), .CK(clk), .Q(
        padder_out[7]), .QN() );
  DFF_X2 _padder__out_reg_31_  ( .D(_padder__n2472 ), .CK(clk), .Q(
        padder_out[39]), .QN() );
  DFF_X2 _padder__done_reg  ( .D(_padder__n1835 ), .CK(clk), .Q(_padder__n602 ), .QN() );
  NOR2_X2 _padder__p0_U49  ( .A1(_padder__p0_n2 ), .A2(_padder__p0_n3 ), .ZN(
        _padder__v0[0]) );
  AND2_X1 _padder__p0_U48  ( .A1(n74), .A2(byte_num[1]), .ZN(_padder__v0[23])
         );
  AND2_X1 _padder__p0_U47  ( .A1(n73), .A2(byte_num[1]), .ZN(_padder__v0[22])
         );
  AND2_X1 _padder__p0_U46  ( .A1(n72), .A2(byte_num[1]), .ZN(_padder__v0[21])
         );
  AND2_X1 _padder__p0_U45  ( .A1(n71), .A2(byte_num[1]), .ZN(_padder__v0[20])
         );
  AND2_X1 _padder__p0_U44  ( .A1(n70), .A2(byte_num[1]), .ZN(_padder__v0[19])
         );
  AND2_X1 _padder__p0_U43  ( .A1(n69), .A2(byte_num[1]), .ZN(_padder__v0[18])
         );
  AND2_X1 _padder__p0_U42  ( .A1(n68), .A2(byte_num[1]), .ZN(_padder__v0[17])
         );
  INV_X4 _padder__p0_U40  ( .A(1'b1), .ZN(_padder__p0_out[7] ) );
  INV_X4 _padder__p0_U38  ( .A(1'b1), .ZN(_padder__p0_out[6] ) );
  INV_X4 _padder__p0_U36  ( .A(1'b1), .ZN(_padder__p0_out[5] ) );
  INV_X4 _padder__p0_U22  ( .A(1'b1), .ZN(_padder__p0_out[4] ) );
  INV_X4 _padder__p0_U20  ( .A(1'b1), .ZN(_padder__p0_out[3] ) );
  INV_X4 _padder__p0_U18  ( .A(1'b1), .ZN(_padder__p0_out[2] ) );
  INV_X4 _padder__p0_U16  ( .A(1'b1), .ZN(_padder__p0_out[1] ) );
  INV_X4 _padder__p0_U35  ( .A(byte_num[0]), .ZN(_padder__p0_n3 ) );
  INV_X4 _padder__p0_U34  ( .A(byte_num[1]), .ZN(_padder__p0_n2 ) );
  INV_X4 _padder__p0_U33  ( .A(n75), .ZN(_padder__p0_n1 ) );
  AND2_X2 _padder__p0_U31  ( .A1(n62), .A2(_padder__v0[0]), .ZN(
        _padder__v0[10]) );
  AND2_X2 _padder__p0_U30  ( .A1(n63), .A2(_padder__v0[0]), .ZN(
        _padder__v0[11]) );
  AND2_X2 _padder__p0_U29  ( .A1(n64), .A2(_padder__v0[0]), .ZN(
        _padder__v0[12]) );
  AND2_X2 _padder__p0_U28  ( .A1(n65), .A2(_padder__v0[0]), .ZN(
        _padder__v0[13]) );
  AND2_X2 _padder__p0_U27  ( .A1(n66), .A2(_padder__v0[0]), .ZN(
        _padder__v0[14]) );
  AND2_X2 _padder__p0_U26  ( .A1(n67), .A2(_padder__v0[0]), .ZN(
        _padder__v0[15]) );
  NAND2_X2 _padder__p0_U25  ( .A1(in[16]), .A2(byte_num[1]), .ZN(
        _padder__p0_n7 ) );
  NAND2_X2 _padder__p0_U24  ( .A1(byte_num[0]), .A2(_padder__p0_n2 ), .ZN(
        _padder__p0_n8 ) );
  NAND2_X2 _padder__p0_U23  ( .A1(_padder__p0_n7 ), .A2(_padder__p0_n8 ), .ZN(
        _padder__v0[16]) );
  NAND2_X2 _padder__p0_U15  ( .A1(_padder__p0_n2 ), .A2(_padder__p0_n3 ), .ZN(
        _padder__p0_n6 ) );
  NAND2_X2 _padder__p0_U14  ( .A1(_padder__p0_n6 ), .A2(_padder__p0_n1 ), .ZN(
        _padder__v0[24]) );
  AND2_X2 _padder__p0_U13  ( .A1(n76), .A2(_padder__p0_n6 ), .ZN(
        _padder__v0[25]) );
  AND2_X2 _padder__p0_U12  ( .A1(n77), .A2(_padder__p0_n6 ), .ZN(
        _padder__v0[26]) );
  AND2_X2 _padder__p0_U11  ( .A1(n78), .A2(_padder__p0_n6 ), .ZN(
        _padder__v0[27]) );
  AND2_X2 _padder__p0_U10  ( .A1(n79), .A2(_padder__p0_n6 ), .ZN(
        _padder__v0[28]) );
  AND2_X2 _padder__p0_U9  ( .A1(n80), .A2(_padder__p0_n6 ), .ZN(
        _padder__v0[29]) );
  AND2_X2 _padder__p0_U8  ( .A1(n81), .A2(_padder__p0_n6 ), .ZN(
        _padder__v0[30]) );
  AND2_X2 _padder__p0_U7  ( .A1(n82), .A2(_padder__p0_n6 ), .ZN(
        _padder__v0[31]) );
  NAND2_X2 _padder__p0_U6  ( .A1(byte_num[1]), .A2(_padder__p0_n3 ), .ZN(
        _padder__p0_n4 ) );
  NAND2_X2 _padder__p0_U5  ( .A1(in[8]), .A2(_padder__v0[0]), .ZN(
        _padder__p0_n5 ) );
  NAND2_X2 _padder__p0_U4  ( .A1(_padder__p0_n4 ), .A2(_padder__p0_n5 ), .ZN(
        _padder__v0[8]) );
  AND2_X2 _padder__p0_U3  ( .A1(n61), .A2(_padder__v0[0]), .ZN(
        _padder__v0[9]) );
  NOR2_X2 _f_permutation__U6271  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5785 ), .ZN(_f_permutation__N6 ) );
  NOR2_X2 _f_permutation__U6270  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5784 ), .ZN(_f_permutation__N7 ) );
  NOR2_X2 _f_permutation__U6269  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5783 ), .ZN(_f_permutation__N8 ) );
  NOR2_X2 _f_permutation__U6268  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5782 ), .ZN(_f_permutation__N9 ) );
  NOR2_X2 _f_permutation__U6267  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5804 ), .ZN(_f_permutation__N10 ) );
  NOR2_X2 _f_permutation__U6266  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5803 ), .ZN(_f_permutation__N11 ) );
  NOR2_X2 _f_permutation__U6265  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5802 ), .ZN(_f_permutation__N12 ) );
  NOR2_X2 _f_permutation__U6264  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5801 ), .ZN(_f_permutation__N13 ) );
  NOR2_X2 _f_permutation__U6263  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5800 ), .ZN(_f_permutation__N14 ) );
  NOR2_X2 _f_permutation__U6262  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5799 ), .ZN(_f_permutation__N15 ) );
  NOR2_X2 _f_permutation__U6261  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5798 ), .ZN(_f_permutation__N16 ) );
  NOR2_X2 _f_permutation__U6260  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5797 ), .ZN(_f_permutation__N17 ) );
  NOR2_X2 _f_permutation__U6259  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5796 ), .ZN(_f_permutation__N18 ) );
  NOR2_X2 _f_permutation__U6258  ( .A1(_f_permutation__n7325 ), .A2(
        _f_permutation__n5795 ), .ZN(_f_permutation__N19 ) );
  NOR2_X2 _f_permutation__U6257  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5794 ), .ZN(_f_permutation__N20 ) );
  NOR2_X2 _f_permutation__U6256  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5793 ), .ZN(_f_permutation__N21 ) );
  NOR2_X2 _f_permutation__U6255  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5792 ), .ZN(_f_permutation__N22 ) );
  NOR2_X2 _f_permutation__U6254  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5791 ), .ZN(_f_permutation__N23 ) );
  NOR2_X2 _f_permutation__U6253  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5790 ), .ZN(_f_permutation__N24 ) );
  NOR2_X2 _f_permutation__U6252  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5789 ), .ZN(_f_permutation__N25 ) );
  NOR2_X2 _f_permutation__U6251  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5788 ), .ZN(_f_permutation__N26 ) );
  NOR2_X2 _f_permutation__U6250  ( .A1(_f_permutation__n7324 ), .A2(
        _f_permutation__n5787 ), .ZN(_f_permutation__N27 ) );
  NAND3_X2 _f_permutation__U6249  ( .A1(_f_permutation__n5786 ), .A2(
        _f_permutation__n7326 ), .A3(_f_permutation__n3 ), .ZN(
        _f_permutation__n7038 ) );
  NOR2_X2 _f_permutation__U6248  ( .A1(_f_permutation__out_ready ), .A2(
        _f_permutation__i[22] ), .ZN(_f_permutation__n2209 ) );
  NOR3_X2 _f_permutation__U6247  ( .A1(_f_permutation__n2209 ), .A2(
        _f_permutation__n7324 ), .A3(f_ack), .ZN(_f_permutation__n5388 ) );
  BUF_X4 _f_permutation__U6246  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7153 ) );
  BUF_X4 _f_permutation__U6245  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7157 ) );
  BUF_X4 _f_permutation__U6244  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7158 ) );
  BUF_X4 _f_permutation__U6243  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7159 ) );
  BUF_X4 _f_permutation__U6242  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7160 ) );
  BUF_X4 _f_permutation__U6241  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7161 ) );
  BUF_X4 _f_permutation__U6240  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7154 ) );
  BUF_X4 _f_permutation__U6239  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7155 ) );
  BUF_X4 _f_permutation__U6238  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7156 ) );
  BUF_X4 _f_permutation__U6237  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7164 ) );
  BUF_X4 _f_permutation__U6236  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7165 ) );
  BUF_X4 _f_permutation__U6235  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7166 ) );
  BUF_X4 _f_permutation__U6234  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7167 ) );
  BUF_X4 _f_permutation__U6233  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7162 ) );
  BUF_X4 _f_permutation__U6232  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7163 ) );
  BUF_X4 _f_permutation__U6231  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7142 ) );
  BUF_X4 _f_permutation__U6230  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7143 ) );
  BUF_X4 _f_permutation__U6229  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7144 ) );
  BUF_X4 _f_permutation__U6228  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7145 ) );
  BUF_X4 _f_permutation__U6227  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7146 ) );
  BUF_X4 _f_permutation__U6226  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7139 ) );
  BUF_X4 _f_permutation__U6225  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7140 ) );
  BUF_X4 _f_permutation__U6224  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7141 ) );
  BUF_X4 _f_permutation__U6223  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7150 ) );
  BUF_X4 _f_permutation__U6222  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7151 ) );
  BUF_X4 _f_permutation__U6221  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7152 ) );
  BUF_X4 _f_permutation__U6220  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7147 ) );
  BUF_X4 _f_permutation__U6219  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7148 ) );
  BUF_X4 _f_permutation__U6218  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7149 ) );
  BUF_X4 _f_permutation__U6217  ( .A(_f_permutation__n7039 ), .Z(
        _f_permutation__n7168 ) );
  BUF_X4 _f_permutation__U6216  ( .A(_f_permutation__n7158 ), .Z(
        _f_permutation__n7087 ) );
  BUF_X4 _f_permutation__U6215  ( .A(_f_permutation__n7160 ), .Z(
        _f_permutation__n7085 ) );
  BUF_X4 _f_permutation__U6214  ( .A(_f_permutation__n7159 ), .Z(
        _f_permutation__n7086 ) );
  BUF_X4 _f_permutation__U6213  ( .A(_f_permutation__n7154 ), .Z(
        _f_permutation__n7093 ) );
  BUF_X4 _f_permutation__U6212  ( .A(_f_permutation__n7154 ), .Z(
        _f_permutation__n7094 ) );
  BUF_X4 _f_permutation__U6211  ( .A(_f_permutation__n7156 ), .Z(
        _f_permutation__n7090 ) );
  BUF_X4 _f_permutation__U6210  ( .A(_f_permutation__n7157 ), .Z(
        _f_permutation__n7088 ) );
  BUF_X4 _f_permutation__U6209  ( .A(_f_permutation__n7156 ), .Z(
        _f_permutation__n7089 ) );
  BUF_X4 _f_permutation__U6208  ( .A(_f_permutation__n7156 ), .Z(
        _f_permutation__n7091 ) );
  BUF_X4 _f_permutation__U6207  ( .A(_f_permutation__n7155 ), .Z(
        _f_permutation__n7092 ) );
  BUF_X4 _f_permutation__U6206  ( .A(_f_permutation__n7165 ), .Z(
        _f_permutation__n7072 ) );
  BUF_X4 _f_permutation__U6205  ( .A(_f_permutation__n7166 ), .Z(
        _f_permutation__n7069 ) );
  BUF_X4 _f_permutation__U6204  ( .A(_f_permutation__n7166 ), .Z(
        _f_permutation__n7070 ) );
  BUF_X4 _f_permutation__U6203  ( .A(_f_permutation__n7166 ), .Z(
        _f_permutation__n7071 ) );
  BUF_X4 _f_permutation__U6202  ( .A(_f_permutation__n7165 ), .Z(
        _f_permutation__n7073 ) );
  BUF_X4 _f_permutation__U6201  ( .A(_f_permutation__n7165 ), .Z(
        _f_permutation__n7074 ) );
  BUF_X4 _f_permutation__U6200  ( .A(_f_permutation__n7167 ), .Z(
        _f_permutation__n7066 ) );
  BUF_X4 _f_permutation__U6199  ( .A(_f_permutation__n7168 ), .Z(
        _f_permutation__n7065 ) );
  BUF_X4 _f_permutation__U6198  ( .A(_f_permutation__n7167 ), .Z(
        _f_permutation__n7067 ) );
  BUF_X4 _f_permutation__U6197  ( .A(_f_permutation__n7167 ), .Z(
        _f_permutation__n7068 ) );
  BUF_X4 _f_permutation__U6196  ( .A(_f_permutation__n7162 ), .Z(
        _f_permutation__n7082 ) );
  BUF_X4 _f_permutation__U6195  ( .A(_f_permutation__n7163 ), .Z(
        _f_permutation__n7079 ) );
  BUF_X4 _f_permutation__U6194  ( .A(_f_permutation__n7162 ), .Z(
        _f_permutation__n7080 ) );
  BUF_X4 _f_permutation__U6193  ( .A(_f_permutation__n7162 ), .Z(
        _f_permutation__n7081 ) );
  BUF_X4 _f_permutation__U6192  ( .A(_f_permutation__n7161 ), .Z(
        _f_permutation__n7083 ) );
  BUF_X4 _f_permutation__U6191  ( .A(_f_permutation__n7161 ), .Z(
        _f_permutation__n7084 ) );
  BUF_X4 _f_permutation__U6190  ( .A(_f_permutation__n7163 ), .Z(
        _f_permutation__n7077 ) );
  BUF_X4 _f_permutation__U6189  ( .A(_f_permutation__n7164 ), .Z(
        _f_permutation__n7075 ) );
  BUF_X4 _f_permutation__U6188  ( .A(_f_permutation__n7164 ), .Z(
        _f_permutation__n7076 ) );
  BUF_X4 _f_permutation__U6187  ( .A(_f_permutation__n7163 ), .Z(
        _f_permutation__n7078 ) );
  BUF_X4 _f_permutation__U6186  ( .A(_f_permutation__n7142 ), .Z(
        _f_permutation__n7127 ) );
  BUF_X4 _f_permutation__U6185  ( .A(_f_permutation__n7143 ), .Z(
        _f_permutation__n7125 ) );
  BUF_X4 _f_permutation__U6184  ( .A(_f_permutation__n7144 ), .Z(
        _f_permutation__n7122 ) );
  BUF_X4 _f_permutation__U6183  ( .A(_f_permutation__n7144 ), .Z(
        _f_permutation__n7123 ) );
  BUF_X4 _f_permutation__U6182  ( .A(_f_permutation__n7143 ), .Z(
        _f_permutation__n7124 ) );
  BUF_X4 _f_permutation__U6181  ( .A(_f_permutation__n7143 ), .Z(
        _f_permutation__n7126 ) );
  BUF_X4 _f_permutation__U6180  ( .A(_f_permutation__n7145 ), .Z(
        _f_permutation__n7119 ) );
  BUF_X4 _f_permutation__U6179  ( .A(_f_permutation__n7146 ), .Z(
        _f_permutation__n7116 ) );
  BUF_X4 _f_permutation__U6178  ( .A(_f_permutation__n7146 ), .Z(
        _f_permutation__n7117 ) );
  BUF_X4 _f_permutation__U6177  ( .A(_f_permutation__n7145 ), .Z(
        _f_permutation__n7118 ) );
  BUF_X4 _f_permutation__U6176  ( .A(_f_permutation__n7145 ), .Z(
        _f_permutation__n7120 ) );
  BUF_X4 _f_permutation__U6175  ( .A(_f_permutation__n7144 ), .Z(
        _f_permutation__n7121 ) );
  BUF_X4 _f_permutation__U6174  ( .A(_f_permutation__n7139 ), .Z(
        _f_permutation__n7136 ) );
  BUF_X4 _f_permutation__U6173  ( .A(_f_permutation__n7140 ), .Z(
        _f_permutation__n7133 ) );
  BUF_X4 _f_permutation__U6172  ( .A(_f_permutation__n7140 ), .Z(
        _f_permutation__n7134 ) );
  BUF_X4 _f_permutation__U6171  ( .A(_f_permutation__n7140 ), .Z(
        _f_permutation__n7135 ) );
  BUF_X4 _f_permutation__U6170  ( .A(_f_permutation__n7139 ), .Z(
        _f_permutation__n7137 ) );
  BUF_X4 _f_permutation__U6169  ( .A(_f_permutation__n7139 ), .Z(
        _f_permutation__n7138 ) );
  BUF_X4 _f_permutation__U6168  ( .A(_f_permutation__n7141 ), .Z(
        _f_permutation__n7130 ) );
  BUF_X4 _f_permutation__U6167  ( .A(_f_permutation__n7142 ), .Z(
        _f_permutation__n7128 ) );
  BUF_X4 _f_permutation__U6166  ( .A(_f_permutation__n7142 ), .Z(
        _f_permutation__n7129 ) );
  BUF_X4 _f_permutation__U6165  ( .A(_f_permutation__n7141 ), .Z(
        _f_permutation__n7131 ) );
  BUF_X4 _f_permutation__U6164  ( .A(_f_permutation__n7141 ), .Z(
        _f_permutation__n7132 ) );
  BUF_X4 _f_permutation__U6163  ( .A(_f_permutation__n7150 ), .Z(
        _f_permutation__n7105 ) );
  BUF_X4 _f_permutation__U6162  ( .A(_f_permutation__n7151 ), .Z(
        _f_permutation__n7102 ) );
  BUF_X4 _f_permutation__U6161  ( .A(_f_permutation__n7151 ), .Z(
        _f_permutation__n7100 ) );
  BUF_X4 _f_permutation__U6160  ( .A(_f_permutation__n7151 ), .Z(
        _f_permutation__n7101 ) );
  BUF_X4 _f_permutation__U6159  ( .A(_f_permutation__n7150 ), .Z(
        _f_permutation__n7103 ) );
  BUF_X4 _f_permutation__U6158  ( .A(_f_permutation__n7150 ), .Z(
        _f_permutation__n7104 ) );
  BUF_X4 _f_permutation__U6157  ( .A(_f_permutation__n7152 ), .Z(
        _f_permutation__n7097 ) );
  BUF_X4 _f_permutation__U6156  ( .A(_f_permutation__n7153 ), .Z(
        _f_permutation__n7095 ) );
  BUF_X4 _f_permutation__U6155  ( .A(_f_permutation__n7153 ), .Z(
        _f_permutation__n7096 ) );
  BUF_X4 _f_permutation__U6154  ( .A(_f_permutation__n7152 ), .Z(
        _f_permutation__n7098 ) );
  BUF_X4 _f_permutation__U6153  ( .A(_f_permutation__n7152 ), .Z(
        _f_permutation__n7099 ) );
  BUF_X4 _f_permutation__U6152  ( .A(_f_permutation__n7147 ), .Z(
        _f_permutation__n7114 ) );
  BUF_X4 _f_permutation__U6151  ( .A(_f_permutation__n7148 ), .Z(
        _f_permutation__n7111 ) );
  BUF_X4 _f_permutation__U6150  ( .A(_f_permutation__n7147 ), .Z(
        _f_permutation__n7112 ) );
  BUF_X4 _f_permutation__U6149  ( .A(_f_permutation__n7147 ), .Z(
        _f_permutation__n7113 ) );
  BUF_X4 _f_permutation__U6148  ( .A(_f_permutation__n7146 ), .Z(
        _f_permutation__n7115 ) );
  BUF_X4 _f_permutation__U6147  ( .A(_f_permutation__n7149 ), .Z(
        _f_permutation__n7108 ) );
  BUF_X4 _f_permutation__U6146  ( .A(_f_permutation__n7149 ), .Z(
        _f_permutation__n7106 ) );
  BUF_X4 _f_permutation__U6145  ( .A(_f_permutation__n7149 ), .Z(
        _f_permutation__n7107 ) );
  BUF_X4 _f_permutation__U6144  ( .A(_f_permutation__n7148 ), .Z(
        _f_permutation__n7109 ) );
  BUF_X4 _f_permutation__U6143  ( .A(_f_permutation__n7148 ), .Z(
        _f_permutation__n7110 ) );
  INV_X4 _f_permutation__U6142  ( .A(n115), .ZN(_f_permutation__n7326 ) );
  INV_X4 _f_permutation__U6141  ( .A(_f_permutation__n7040 ), .ZN(f_ack) );
  INV_X4 _f_permutation__U6140  ( .A(_f_permutation__n7326 ), .ZN(
        _f_permutation__n7325 ) );
  INV_X4 _f_permutation__U6139  ( .A(_f_permutation__n7326 ), .ZN(
        _f_permutation__n7324 ) );
  INV_X4 _f_permutation__U6138  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7316 ) );
  INV_X4 _f_permutation__U6137  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7321 ) );
  INV_X4 _f_permutation__U6136  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7317 ) );
  INV_X4 _f_permutation__U6135  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7318 ) );
  INV_X4 _f_permutation__U6134  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7315 ) );
  INV_X4 _f_permutation__U6133  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7322 ) );
  INV_X4 _f_permutation__U6132  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7312 ) );
  INV_X4 _f_permutation__U6131  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7319 ) );
  INV_X4 _f_permutation__U6130  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7314 ) );
  INV_X4 _f_permutation__U6129  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7320 ) );
  INV_X4 _f_permutation__U6128  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7323 ) );
  INV_X4 _f_permutation__U6127  ( .A(_f_permutation__n7040 ), .ZN(
        _f_permutation__n7313 ) );
  BUF_X4 _f_permutation__U6126  ( .A(_f_permutation__n7041 ), .Z(
        _f_permutation__n7310 ) );
  BUF_X4 _f_permutation__U6125  ( .A(_f_permutation__n7310 ), .Z(
        _f_permutation__n7308 ) );
  BUF_X4 _f_permutation__U6124  ( .A(_f_permutation__n7310 ), .Z(
        _f_permutation__n7307 ) );
  BUF_X4 _f_permutation__U6123  ( .A(_f_permutation__n7310 ), .Z(
        _f_permutation__n7306 ) );
  BUF_X4 _f_permutation__U6122  ( .A(_f_permutation__n7310 ), .Z(
        _f_permutation__n7309 ) );
  BUF_X4 _f_permutation__U6121  ( .A(_f_permutation__n7041 ), .Z(
        _f_permutation__n7305 ) );
  BUF_X4 _f_permutation__U6120  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7177 ) );
  BUF_X4 _f_permutation__U6119  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7176 ) );
  BUF_X4 _f_permutation__U6118  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7175 ) );
  BUF_X4 _f_permutation__U6117  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7174 ) );
  BUF_X4 _f_permutation__U6116  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7173 ) );
  BUF_X4 _f_permutation__U6115  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7172 ) );
  BUF_X4 _f_permutation__U6114  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7171 ) );
  BUF_X4 _f_permutation__U6113  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7170 ) );
  BUF_X4 _f_permutation__U6112  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7169 ) );
  BUF_X4 _f_permutation__U6111  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7304 ) );
  BUF_X4 _f_permutation__U6110  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7303 ) );
  BUF_X4 _f_permutation__U6109  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7220 ) );
  BUF_X4 _f_permutation__U6108  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7219 ) );
  BUF_X4 _f_permutation__U6107  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7218 ) );
  BUF_X4 _f_permutation__U6106  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7217 ) );
  BUF_X4 _f_permutation__U6105  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7216 ) );
  BUF_X4 _f_permutation__U6104  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7215 ) );
  BUF_X4 _f_permutation__U6103  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7214 ) );
  BUF_X4 _f_permutation__U6102  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7213 ) );
  BUF_X4 _f_permutation__U6101  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7212 ) );
  BUF_X4 _f_permutation__U6100  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7211 ) );
  BUF_X4 _f_permutation__U6099  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7210 ) );
  BUF_X4 _f_permutation__U6098  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7209 ) );
  BUF_X4 _f_permutation__U6097  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7208 ) );
  BUF_X4 _f_permutation__U6096  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7207 ) );
  BUF_X4 _f_permutation__U6095  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7206 ) );
  BUF_X4 _f_permutation__U6094  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7205 ) );
  BUF_X4 _f_permutation__U6093  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7204 ) );
  BUF_X4 _f_permutation__U6092  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7203 ) );
  BUF_X4 _f_permutation__U6091  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7202 ) );
  BUF_X4 _f_permutation__U6090  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7201 ) );
  BUF_X4 _f_permutation__U6089  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7200 ) );
  BUF_X4 _f_permutation__U6088  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7199 ) );
  BUF_X4 _f_permutation__U6087  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7198 ) );
  BUF_X4 _f_permutation__U6086  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7197 ) );
  BUF_X4 _f_permutation__U6085  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7196 ) );
  BUF_X4 _f_permutation__U6084  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7195 ) );
  BUF_X4 _f_permutation__U6083  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7194 ) );
  BUF_X4 _f_permutation__U6082  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7193 ) );
  BUF_X4 _f_permutation__U6081  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7192 ) );
  BUF_X4 _f_permutation__U6080  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7191 ) );
  BUF_X4 _f_permutation__U6079  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7190 ) );
  BUF_X4 _f_permutation__U6078  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7189 ) );
  BUF_X4 _f_permutation__U6077  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7188 ) );
  BUF_X4 _f_permutation__U6076  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7187 ) );
  BUF_X4 _f_permutation__U6075  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7186 ) );
  BUF_X4 _f_permutation__U6074  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7185 ) );
  BUF_X4 _f_permutation__U6073  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7184 ) );
  BUF_X4 _f_permutation__U6072  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7183 ) );
  BUF_X4 _f_permutation__U6071  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7182 ) );
  BUF_X4 _f_permutation__U6070  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7181 ) );
  BUF_X4 _f_permutation__U6069  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7180 ) );
  BUF_X4 _f_permutation__U6068  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7179 ) );
  BUF_X4 _f_permutation__U6067  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7178 ) );
  BUF_X4 _f_permutation__U6066  ( .A(_f_permutation__n7041 ), .Z(
        _f_permutation__n7302 ) );
  BUF_X4 _f_permutation__U6065  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7301 ) );
  BUF_X4 _f_permutation__U6064  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7300 ) );
  BUF_X4 _f_permutation__U6063  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7299 ) );
  BUF_X4 _f_permutation__U6062  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7298 ) );
  BUF_X4 _f_permutation__U6061  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7297 ) );
  BUF_X4 _f_permutation__U6060  ( .A(_f_permutation__n7041 ), .Z(
        _f_permutation__n7296 ) );
  BUF_X4 _f_permutation__U6059  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7295 ) );
  BUF_X4 _f_permutation__U6058  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7294 ) );
  BUF_X4 _f_permutation__U6057  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7293 ) );
  BUF_X4 _f_permutation__U6056  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7292 ) );
  BUF_X4 _f_permutation__U6055  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7291 ) );
  BUF_X4 _f_permutation__U6054  ( .A(_f_permutation__n7283 ), .Z(
        _f_permutation__n7290 ) );
  BUF_X4 _f_permutation__U6053  ( .A(_f_permutation__n7284 ), .Z(
        _f_permutation__n7289 ) );
  BUF_X4 _f_permutation__U6052  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7288 ) );
  BUF_X4 _f_permutation__U6051  ( .A(_f_permutation__n7248 ), .Z(
        _f_permutation__n7287 ) );
  BUF_X4 _f_permutation__U6050  ( .A(_f_permutation__n7259 ), .Z(
        _f_permutation__n7286 ) );
  BUF_X4 _f_permutation__U6049  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7285 ) );
  BUF_X4 _f_permutation__U6048  ( .A(_f_permutation__n7041 ), .Z(
        _f_permutation__n7284 ) );
  BUF_X4 _f_permutation__U6047  ( .A(_f_permutation__n7310 ), .Z(
        _f_permutation__n7283 ) );
  BUF_X4 _f_permutation__U6046  ( .A(_f_permutation__n7041 ), .Z(
        _f_permutation__n7282 ) );
  BUF_X4 _f_permutation__U6045  ( .A(_f_permutation__n7284 ), .Z(
        _f_permutation__n7281 ) );
  BUF_X4 _f_permutation__U6044  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7280 ) );
  BUF_X4 _f_permutation__U6043  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7279 ) );
  BUF_X4 _f_permutation__U6042  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7278 ) );
  BUF_X4 _f_permutation__U6041  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7277 ) );
  BUF_X4 _f_permutation__U6040  ( .A(_f_permutation__n7284 ), .Z(
        _f_permutation__n7276 ) );
  BUF_X4 _f_permutation__U6039  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7275 ) );
  BUF_X4 _f_permutation__U6038  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7274 ) );
  BUF_X4 _f_permutation__U6037  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7273 ) );
  BUF_X4 _f_permutation__U6036  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7272 ) );
  BUF_X4 _f_permutation__U6035  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7271 ) );
  BUF_X4 _f_permutation__U6034  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7270 ) );
  BUF_X4 _f_permutation__U6033  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7269 ) );
  BUF_X4 _f_permutation__U6032  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7268 ) );
  BUF_X4 _f_permutation__U6031  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7267 ) );
  BUF_X4 _f_permutation__U6030  ( .A(_f_permutation__n7230 ), .Z(
        _f_permutation__n7266 ) );
  BUF_X4 _f_permutation__U6029  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7265 ) );
  BUF_X4 _f_permutation__U6028  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7264 ) );
  BUF_X4 _f_permutation__U6027  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7263 ) );
  BUF_X4 _f_permutation__U6026  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7262 ) );
  BUF_X4 _f_permutation__U6025  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7261 ) );
  BUF_X4 _f_permutation__U6024  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7260 ) );
  BUF_X4 _f_permutation__U6023  ( .A(_f_permutation__n7310 ), .Z(
        _f_permutation__n7259 ) );
  BUF_X4 _f_permutation__U6022  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7258 ) );
  BUF_X4 _f_permutation__U6021  ( .A(_f_permutation__n7284 ), .Z(
        _f_permutation__n7257 ) );
  BUF_X4 _f_permutation__U6020  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7256 ) );
  BUF_X4 _f_permutation__U6019  ( .A(_f_permutation__n7283 ), .Z(
        _f_permutation__n7255 ) );
  BUF_X4 _f_permutation__U6018  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7254 ) );
  BUF_X4 _f_permutation__U6017  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7253 ) );
  BUF_X4 _f_permutation__U6016  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7252 ) );
  BUF_X4 _f_permutation__U6015  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7251 ) );
  BUF_X4 _f_permutation__U6014  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7250 ) );
  BUF_X4 _f_permutation__U6013  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7249 ) );
  BUF_X4 _f_permutation__U6012  ( .A(_f_permutation__n7310 ), .Z(
        _f_permutation__n7248 ) );
  BUF_X4 _f_permutation__U6011  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7247 ) );
  BUF_X4 _f_permutation__U6010  ( .A(_f_permutation__n7284 ), .Z(
        _f_permutation__n7246 ) );
  BUF_X4 _f_permutation__U6009  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7245 ) );
  BUF_X4 _f_permutation__U6008  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7244 ) );
  BUF_X4 _f_permutation__U6007  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7243 ) );
  BUF_X4 _f_permutation__U6006  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7242 ) );
  BUF_X4 _f_permutation__U6005  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7241 ) );
  BUF_X4 _f_permutation__U6004  ( .A(_f_permutation__n7308 ), .Z(
        _f_permutation__n7240 ) );
  BUF_X4 _f_permutation__U6003  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7239 ) );
  BUF_X4 _f_permutation__U6002  ( .A(_f_permutation__n7306 ), .Z(
        _f_permutation__n7238 ) );
  BUF_X4 _f_permutation__U6001  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7237 ) );
  BUF_X4 _f_permutation__U6000  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7236 ) );
  BUF_X4 _f_permutation__U5999  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7235 ) );
  BUF_X4 _f_permutation__U5998  ( .A(_f_permutation__n7307 ), .Z(
        _f_permutation__n7234 ) );
  BUF_X4 _f_permutation__U5997  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7233 ) );
  BUF_X4 _f_permutation__U5996  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7232 ) );
  BUF_X4 _f_permutation__U5995  ( .A(_f_permutation__n7284 ), .Z(
        _f_permutation__n7231 ) );
  BUF_X4 _f_permutation__U5994  ( .A(_f_permutation__n7310 ), .Z(
        _f_permutation__n7230 ) );
  BUF_X4 _f_permutation__U5993  ( .A(_f_permutation__n7302 ), .Z(
        _f_permutation__n7229 ) );
  BUF_X4 _f_permutation__U5992  ( .A(_f_permutation__n7296 ), .Z(
        _f_permutation__n7228 ) );
  BUF_X4 _f_permutation__U5991  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7227 ) );
  BUF_X4 _f_permutation__U5990  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7226 ) );
  BUF_X4 _f_permutation__U5989  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7225 ) );
  BUF_X4 _f_permutation__U5988  ( .A(_f_permutation__n7282 ), .Z(
        _f_permutation__n7224 ) );
  BUF_X4 _f_permutation__U5986  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7223 ) );
  BUF_X4 _f_permutation__U5985  ( .A(_f_permutation__n7309 ), .Z(
        _f_permutation__n7222 ) );
  BUF_X4 _f_permutation__U5984  ( .A(_f_permutation__n7305 ), .Z(
        _f_permutation__n7221 ) );
  CLKBUF_X2 _f_permutation__U5983  ( .A(_f_permutation__N6 ), .Z(
        _f_permutation__n7063 ) );
  CLKBUF_X2 _f_permutation__U5982  ( .A(_f_permutation__N7 ), .Z(
        _f_permutation__n7062 ) );
  CLKBUF_X2 _f_permutation__U5981  ( .A(_f_permutation__N8 ), .Z(
        _f_permutation__n7061 ) );
  CLKBUF_X2 _f_permutation__U5980  ( .A(_f_permutation__N9 ), .Z(
        _f_permutation__n7060 ) );
  CLKBUF_X2 _f_permutation__U5979  ( .A(_f_permutation__N20 ), .Z(
        _f_permutation__n7059 ) );
  CLKBUF_X2 _f_permutation__U5978  ( .A(_f_permutation__N21 ), .Z(
        _f_permutation__n7058 ) );
  CLKBUF_X2 _f_permutation__U5977  ( .A(_f_permutation__N22 ), .Z(
        _f_permutation__n7057 ) );
  CLKBUF_X2 _f_permutation__U5976  ( .A(_f_permutation__N23 ), .Z(
        _f_permutation__n7056 ) );
  CLKBUF_X2 _f_permutation__U5975  ( .A(_f_permutation__N24 ), .Z(
        _f_permutation__n7055 ) );
  CLKBUF_X2 _f_permutation__U5974  ( .A(_f_permutation__N25 ), .Z(
        _f_permutation__n7054 ) );
  CLKBUF_X2 _f_permutation__U5973  ( .A(_f_permutation__N26 ), .Z(
        _f_permutation__n7053 ) );
  CLKBUF_X2 _f_permutation__U5972  ( .A(_f_permutation__N27 ), .Z(
        _f_permutation__n7052 ) );
  CLKBUF_X2 _f_permutation__U5971  ( .A(_f_permutation__N10 ), .Z(
        _f_permutation__n7051 ) );
  CLKBUF_X2 _f_permutation__U5970  ( .A(_f_permutation__N11 ), .Z(
        _f_permutation__n7050 ) );
  CLKBUF_X2 _f_permutation__U5969  ( .A(_f_permutation__N12 ), .Z(
        _f_permutation__n7049 ) );
  CLKBUF_X2 _f_permutation__U5968  ( .A(_f_permutation__N13 ), .Z(
        _f_permutation__n7048 ) );
  CLKBUF_X2 _f_permutation__U5966  ( .A(_f_permutation__N14 ), .Z(
        _f_permutation__n7047 ) );
  CLKBUF_X2 _f_permutation__U5964  ( .A(_f_permutation__N15 ), .Z(
        _f_permutation__n7046 ) );
  CLKBUF_X2 _f_permutation__U5963  ( .A(_f_permutation__N19 ), .Z(
        _f_permutation__n7045 ) );
  CLKBUF_X2 _f_permutation__U5962  ( .A(_f_permutation__N18 ), .Z(
        _f_permutation__n7044 ) );
  CLKBUF_X2 _f_permutation__U5961  ( .A(_f_permutation__N17 ), .Z(
        _f_permutation__n7043 ) );
  CLKBUF_X2 _f_permutation__U5959  ( .A(_f_permutation__N16 ), .Z(
        _f_permutation__n7042 ) );
  NOR2_X2 _f_permutation__U5957  ( .A1(_f_permutation__n7039 ), .A2(
        _f_permutation__n7324 ), .ZN(_f_permutation__n7041 ) );
  NAND2_X2 _f_permutation__U1157  ( .A1(padder_out_ready), .A2(
        _f_permutation__n7064 ), .ZN(_f_permutation__n7040 ) );
  NAND2_X2 _f_permutation__U1156  ( .A1(_f_permutation__n2208 ), .A2(
        _f_permutation__n7037 ), .ZN(_f_permutation__n7039 ) );
  DFF_X1 _f_permutation__out_ready_reg  ( .D(_f_permutation__n5388 ), .CK(clk), 
        .Q(_f_permutation__out_ready ), .QN() );
  DFF_X1 _f_permutation__calc_reg  ( .D(_f_permutation__N29 ), .CK(clk), .Q(
        _f_permutation__n3 ), .QN(_f_permutation__n7064 ) );
  DFF_X1 _f_permutation__i_reg_0_  ( .D(_f_permutation__n1628 ), .CK(clk), .Q(
        _f_permutation__i[0] ), .QN(_f_permutation__n5785 ) );
  DFF_X1 _f_permutation__i_reg_1_  ( .D(_f_permutation__n7063 ), .CK(clk), .Q(
        _f_permutation__i[1] ), .QN(_f_permutation__n5784 ) );
  DFF_X1 _f_permutation__i_reg_2_  ( .D(_f_permutation__n7062 ), .CK(clk), .Q(
        _f_permutation__i[2] ), .QN(_f_permutation__n5783 ) );
  DFF_X1 _f_permutation__i_reg_3_  ( .D(_f_permutation__n7061 ), .CK(clk), .Q(
        _f_permutation__i[3] ), .QN(_f_permutation__n5782 ) );
  DFF_X1 _f_permutation__i_reg_4_  ( .D(_f_permutation__n7060 ), .CK(clk), .Q(
        _f_permutation__i[4] ), .QN(_f_permutation__n5804 ) );
  DFF_X1 _f_permutation__i_reg_15_  ( .D(_f_permutation__n7059 ), .CK(clk), 
        .Q(_f_permutation__i[15] ), .QN(_f_permutation__n5793 ) );
  DFF_X1 _f_permutation__i_reg_16_  ( .D(_f_permutation__n7058 ), .CK(clk), 
        .Q(_f_permutation__i[16] ), .QN(_f_permutation__n5792 ) );
  DFF_X1 _f_permutation__i_reg_17_  ( .D(_f_permutation__n7057 ), .CK(clk), 
        .Q(_f_permutation__i[17] ), .QN(_f_permutation__n5791 ) );
  DFF_X1 _f_permutation__i_reg_18_  ( .D(_f_permutation__n7056 ), .CK(clk), 
        .Q(_f_permutation__i[18] ), .QN(_f_permutation__n5790 ) );
  DFF_X1 _f_permutation__i_reg_19_  ( .D(_f_permutation__n7055 ), .CK(clk), 
        .Q(_f_permutation__i[19] ), .QN(_f_permutation__n5789 ) );
  DFF_X1 _f_permutation__i_reg_20_  ( .D(_f_permutation__n7054 ), .CK(clk), 
        .Q(_f_permutation__i[20] ), .QN(_f_permutation__n5788 ) );
  DFF_X1 _f_permutation__i_reg_21_  ( .D(_f_permutation__n7053 ), .CK(clk), 
        .Q(_f_permutation__i[21] ), .QN(_f_permutation__n5787 ) );
  DFF_X1 _f_permutation__i_reg_22_  ( .D(_f_permutation__n7052 ), .CK(clk), 
        .Q(_f_permutation__i[22] ), .QN(_f_permutation__n5786 ) );
  DFF_X1 _f_permutation__i_reg_5_  ( .D(_f_permutation__n7051 ), .CK(clk), .Q(
        _f_permutation__i[5] ), .QN(_f_permutation__n5803 ) );
  DFF_X1 _f_permutation__i_reg_6_  ( .D(_f_permutation__n7050 ), .CK(clk), .Q(
        _f_permutation__i[6] ), .QN(_f_permutation__n5802 ) );
  DFF_X1 _f_permutation__i_reg_7_  ( .D(_f_permutation__n7049 ), .CK(clk), .Q(
        _f_permutation__i[7] ), .QN(_f_permutation__n5801 ) );
  DFF_X1 _f_permutation__i_reg_8_  ( .D(_f_permutation__n7048 ), .CK(clk), .Q(
        _f_permutation__i[8] ), .QN(_f_permutation__n5800 ) );
  DFF_X1 _f_permutation__i_reg_9_  ( .D(_f_permutation__n7047 ), .CK(clk), .Q(
        _f_permutation__i[9] ), .QN(_f_permutation__n5799 ) );
  DFF_X1 _f_permutation__i_reg_10_  ( .D(_f_permutation__n7046 ), .CK(clk), 
        .Q(_f_permutation__i[10] ), .QN(_f_permutation__n5798 ) );
  DFF_X1 _f_permutation__i_reg_11_  ( .D(_f_permutation__n7042 ), .CK(clk), 
        .Q(_f_permutation__i[11] ), .QN(_f_permutation__n5797 ) );
  DFF_X1 _f_permutation__i_reg_12_  ( .D(_f_permutation__n7043 ), .CK(clk), 
        .Q(_f_permutation__i[12] ), .QN(_f_permutation__n5796 ) );
  DFF_X1 _f_permutation__i_reg_13_  ( .D(_f_permutation__n7044 ), .CK(clk), 
        .Q(_f_permutation__i[13] ), .QN(_f_permutation__n5795 ) );
  DFF_X1 _f_permutation__i_reg_14_  ( .D(_f_permutation__n7045 ), .CK(clk), 
        .Q(_f_permutation__i[14] ), .QN(_f_permutation__n5794 ) );
  INV_X4 _f_permutation__U5987  ( .A(_f_permutation__n2208 ), .ZN(
        _f_permutation__n1628 ) );
  NAND2_X2 _f_permutation__U5967  ( .A1(f_ack), .A2(_f_permutation__n7326 ), 
        .ZN(_f_permutation__n2208 ) );
  NAND2_X2 _f_permutation__U5965  ( .A1(_f_permutation__n2208 ), .A2(
        _f_permutation__n7038 ), .ZN(_f_permutation__N29 ) );
  NAND2_X2 _f_permutation__U5960  ( .A1(_f_permutation__n3 ), .A2(
        _f_permutation__n7326 ), .ZN(_f_permutation__n7037 ) );
  NAND2_X2 _f_permutation__U5958  ( .A1(_f_permutation__round_out[1599]), 
        .A2(_f_permutation__n7168 ), .ZN(_f_permutation__n7035 ) );
  NAND2_X2 _f_permutation__U5956  ( .A1(_f_permutation__n7169 ), .A2(out[455]), 
        .ZN(_f_permutation__n7036 ) );
  NAND2_X2 _f_permutation__U5955  ( .A1(_f_permutation__n7035 ), .A2(
        _f_permutation__n7036 ), .ZN(_f_permutation__n3788 ) );
  NAND2_X2 _f_permutation__U5954  ( .A1(_f_permutation__round_out[1598]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n7033 ) );
  NAND2_X2 _f_permutation__U5953  ( .A1(_f_permutation__n7169 ), .A2(out[454]), 
        .ZN(_f_permutation__n7034 ) );
  NAND2_X2 _f_permutation__U5952  ( .A1(_f_permutation__n7033 ), .A2(
        _f_permutation__n7034 ), .ZN(_f_permutation__n3789 ) );
  NAND2_X2 _f_permutation__U5951  ( .A1(_f_permutation__round_out[1597]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n7031 ) );
  NAND2_X2 _f_permutation__U5950  ( .A1(_f_permutation__n7169 ), .A2(out[453]), 
        .ZN(_f_permutation__n7032 ) );
  NAND2_X2 _f_permutation__U5949  ( .A1(_f_permutation__n7031 ), .A2(
        _f_permutation__n7032 ), .ZN(_f_permutation__n3790 ) );
  NAND2_X2 _f_permutation__U5948  ( .A1(_f_permutation__round_out[1596]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n7029 ) );
  NAND2_X2 _f_permutation__U5947  ( .A1(_f_permutation__n7169 ), .A2(out[452]), 
        .ZN(_f_permutation__n7030 ) );
  NAND2_X2 _f_permutation__U5946  ( .A1(_f_permutation__n7029 ), .A2(
        _f_permutation__n7030 ), .ZN(_f_permutation__n3791 ) );
  NAND2_X2 _f_permutation__U5945  ( .A1(_f_permutation__round_out[1595]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n7027 ) );
  NAND2_X2 _f_permutation__U5944  ( .A1(_f_permutation__n7169 ), .A2(out[451]), 
        .ZN(_f_permutation__n7028 ) );
  NAND2_X2 _f_permutation__U5943  ( .A1(_f_permutation__n7027 ), .A2(
        _f_permutation__n7028 ), .ZN(_f_permutation__n3792 ) );
  NAND2_X2 _f_permutation__U5942  ( .A1(_f_permutation__round_out[1594]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n7025 ) );
  NAND2_X2 _f_permutation__U5941  ( .A1(_f_permutation__n7169 ), .A2(out[450]), 
        .ZN(_f_permutation__n7026 ) );
  NAND2_X2 _f_permutation__U5940  ( .A1(_f_permutation__n7025 ), .A2(
        _f_permutation__n7026 ), .ZN(_f_permutation__n3793 ) );
  NAND2_X2 _f_permutation__U5939  ( .A1(_f_permutation__round_out[1593]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n7023 ) );
  NAND2_X2 _f_permutation__U5938  ( .A1(_f_permutation__n7169 ), .A2(out[449]), 
        .ZN(_f_permutation__n7024 ) );
  NAND2_X2 _f_permutation__U5937  ( .A1(_f_permutation__n7023 ), .A2(
        _f_permutation__n7024 ), .ZN(_f_permutation__n3794 ) );
  NAND2_X2 _f_permutation__U5936  ( .A1(_f_permutation__round_out[1592]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7021 ) );
  NAND2_X2 _f_permutation__U5935  ( .A1(_f_permutation__n7169 ), .A2(out[448]), 
        .ZN(_f_permutation__n7022 ) );
  NAND2_X2 _f_permutation__U5934  ( .A1(_f_permutation__n7021 ), .A2(
        _f_permutation__n7022 ), .ZN(_f_permutation__n3795 ) );
  NAND2_X2 _f_permutation__U5933  ( .A1(_f_permutation__round_out[1591]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7019 ) );
  NAND2_X2 _f_permutation__U5932  ( .A1(_f_permutation__n7169 ), .A2(out[463]), 
        .ZN(_f_permutation__n7020 ) );
  NAND2_X2 _f_permutation__U5931  ( .A1(_f_permutation__n7019 ), .A2(
        _f_permutation__n7020 ), .ZN(_f_permutation__n3796 ) );
  NAND2_X2 _f_permutation__U5930  ( .A1(_f_permutation__round_out[1590]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7017 ) );
  NAND2_X2 _f_permutation__U5929  ( .A1(_f_permutation__n7169 ), .A2(out[462]), 
        .ZN(_f_permutation__n7018 ) );
  NAND2_X2 _f_permutation__U5928  ( .A1(_f_permutation__n7017 ), .A2(
        _f_permutation__n7018 ), .ZN(_f_permutation__n3797 ) );
  NAND2_X2 _f_permutation__U5927  ( .A1(_f_permutation__round_out[1589]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7015 ) );
  NAND2_X2 _f_permutation__U5926  ( .A1(_f_permutation__n7169 ), .A2(out[461]), 
        .ZN(_f_permutation__n7016 ) );
  NAND2_X2 _f_permutation__U5925  ( .A1(_f_permutation__n7015 ), .A2(
        _f_permutation__n7016 ), .ZN(_f_permutation__n3798 ) );
  NAND2_X2 _f_permutation__U5924  ( .A1(_f_permutation__round_out[1588]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7013 ) );
  NAND2_X2 _f_permutation__U5923  ( .A1(_f_permutation__n7170 ), .A2(out[460]), 
        .ZN(_f_permutation__n7014 ) );
  NAND2_X2 _f_permutation__U5922  ( .A1(_f_permutation__n7013 ), .A2(
        _f_permutation__n7014 ), .ZN(_f_permutation__n3799 ) );
  NAND2_X2 _f_permutation__U5921  ( .A1(_f_permutation__round_out[1587]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7011 ) );
  NAND2_X2 _f_permutation__U5920  ( .A1(_f_permutation__n7170 ), .A2(out[459]), 
        .ZN(_f_permutation__n7012 ) );
  NAND2_X2 _f_permutation__U5919  ( .A1(_f_permutation__n7011 ), .A2(
        _f_permutation__n7012 ), .ZN(_f_permutation__n3800 ) );
  NAND2_X2 _f_permutation__U5918  ( .A1(_f_permutation__round_out[1586]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7009 ) );
  NAND2_X2 _f_permutation__U5917  ( .A1(_f_permutation__n7170 ), .A2(out[458]), 
        .ZN(_f_permutation__n7010 ) );
  NAND2_X2 _f_permutation__U5916  ( .A1(_f_permutation__n7009 ), .A2(
        _f_permutation__n7010 ), .ZN(_f_permutation__n3801 ) );
  NAND2_X2 _f_permutation__U5915  ( .A1(_f_permutation__round_out[1585]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7007 ) );
  NAND2_X2 _f_permutation__U5914  ( .A1(_f_permutation__n7170 ), .A2(out[457]), 
        .ZN(_f_permutation__n7008 ) );
  NAND2_X2 _f_permutation__U5913  ( .A1(_f_permutation__n7007 ), .A2(
        _f_permutation__n7008 ), .ZN(_f_permutation__n3802 ) );
  NAND2_X2 _f_permutation__U5912  ( .A1(_f_permutation__round_out[1584]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7005 ) );
  NAND2_X2 _f_permutation__U5911  ( .A1(_f_permutation__n7170 ), .A2(out[456]), 
        .ZN(_f_permutation__n7006 ) );
  NAND2_X2 _f_permutation__U5910  ( .A1(_f_permutation__n7005 ), .A2(
        _f_permutation__n7006 ), .ZN(_f_permutation__n3803 ) );
  NAND2_X2 _f_permutation__U5909  ( .A1(_f_permutation__round_out[1583]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7003 ) );
  NAND2_X2 _f_permutation__U5908  ( .A1(_f_permutation__n7170 ), .A2(out[471]), 
        .ZN(_f_permutation__n7004 ) );
  NAND2_X2 _f_permutation__U5907  ( .A1(_f_permutation__n7003 ), .A2(
        _f_permutation__n7004 ), .ZN(_f_permutation__n3804 ) );
  NAND2_X2 _f_permutation__U5906  ( .A1(_f_permutation__round_out[1582]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n7001 ) );
  NAND2_X2 _f_permutation__U5905  ( .A1(_f_permutation__n7170 ), .A2(out[470]), 
        .ZN(_f_permutation__n7002 ) );
  NAND2_X2 _f_permutation__U5904  ( .A1(_f_permutation__n7001 ), .A2(
        _f_permutation__n7002 ), .ZN(_f_permutation__n3805 ) );
  NAND2_X2 _f_permutation__U5903  ( .A1(_f_permutation__round_out[1581]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n6999 ) );
  NAND2_X2 _f_permutation__U5902  ( .A1(_f_permutation__n7170 ), .A2(out[469]), 
        .ZN(_f_permutation__n7000 ) );
  NAND2_X2 _f_permutation__U5901  ( .A1(_f_permutation__n6999 ), .A2(
        _f_permutation__n7000 ), .ZN(_f_permutation__n3806 ) );
  NAND2_X2 _f_permutation__U5900  ( .A1(_f_permutation__round_out[1580]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n6997 ) );
  NAND2_X2 _f_permutation__U5899  ( .A1(_f_permutation__n7170 ), .A2(out[468]), 
        .ZN(_f_permutation__n6998 ) );
  NAND2_X2 _f_permutation__U5898  ( .A1(_f_permutation__n6997 ), .A2(
        _f_permutation__n6998 ), .ZN(_f_permutation__n3807 ) );
  NAND2_X2 _f_permutation__U5897  ( .A1(_f_permutation__round_out[1579]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n6995 ) );
  NAND2_X2 _f_permutation__U5896  ( .A1(_f_permutation__n7170 ), .A2(out[467]), 
        .ZN(_f_permutation__n6996 ) );
  NAND2_X2 _f_permutation__U5895  ( .A1(_f_permutation__n6995 ), .A2(
        _f_permutation__n6996 ), .ZN(_f_permutation__n3808 ) );
  NAND2_X2 _f_permutation__U5894  ( .A1(_f_permutation__round_out[1578]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n6993 ) );
  NAND2_X2 _f_permutation__U5893  ( .A1(_f_permutation__n7170 ), .A2(out[466]), 
        .ZN(_f_permutation__n6994 ) );
  NAND2_X2 _f_permutation__U5892  ( .A1(_f_permutation__n6993 ), .A2(
        _f_permutation__n6994 ), .ZN(_f_permutation__n3809 ) );
  NAND2_X2 _f_permutation__U5891  ( .A1(_f_permutation__round_out[1577]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n6991 ) );
  NAND2_X2 _f_permutation__U5890  ( .A1(_f_permutation__n7171 ), .A2(out[465]), 
        .ZN(_f_permutation__n6992 ) );
  NAND2_X2 _f_permutation__U5889  ( .A1(_f_permutation__n6991 ), .A2(
        _f_permutation__n6992 ), .ZN(_f_permutation__n3810 ) );
  NAND2_X2 _f_permutation__U5888  ( .A1(_f_permutation__round_out[1576]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n6989 ) );
  NAND2_X2 _f_permutation__U5887  ( .A1(_f_permutation__n7171 ), .A2(out[464]), 
        .ZN(_f_permutation__n6990 ) );
  NAND2_X2 _f_permutation__U5886  ( .A1(_f_permutation__n6989 ), .A2(
        _f_permutation__n6990 ), .ZN(_f_permutation__n3811 ) );
  NAND2_X2 _f_permutation__U5885  ( .A1(_f_permutation__round_out[1575]), 
        .A2(_f_permutation__n7110 ), .ZN(_f_permutation__n6987 ) );
  NAND2_X2 _f_permutation__U5884  ( .A1(_f_permutation__n7171 ), .A2(out[479]), 
        .ZN(_f_permutation__n6988 ) );
  NAND2_X2 _f_permutation__U5883  ( .A1(_f_permutation__n6987 ), .A2(
        _f_permutation__n6988 ), .ZN(_f_permutation__n3812 ) );
  NAND2_X2 _f_permutation__U5882  ( .A1(_f_permutation__round_out[1574]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6985 ) );
  NAND2_X2 _f_permutation__U5881  ( .A1(_f_permutation__n7171 ), .A2(out[478]), 
        .ZN(_f_permutation__n6986 ) );
  NAND2_X2 _f_permutation__U5880  ( .A1(_f_permutation__n6985 ), .A2(
        _f_permutation__n6986 ), .ZN(_f_permutation__n3813 ) );
  NAND2_X2 _f_permutation__U5879  ( .A1(_f_permutation__round_out[1573]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6983 ) );
  NAND2_X2 _f_permutation__U5878  ( .A1(_f_permutation__n7171 ), .A2(out[477]), 
        .ZN(_f_permutation__n6984 ) );
  NAND2_X2 _f_permutation__U5877  ( .A1(_f_permutation__n6983 ), .A2(
        _f_permutation__n6984 ), .ZN(_f_permutation__n3814 ) );
  NAND2_X2 _f_permutation__U5876  ( .A1(_f_permutation__round_out[1572]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6981 ) );
  NAND2_X2 _f_permutation__U5875  ( .A1(_f_permutation__n7171 ), .A2(out[476]), 
        .ZN(_f_permutation__n6982 ) );
  NAND2_X2 _f_permutation__U5874  ( .A1(_f_permutation__n6981 ), .A2(
        _f_permutation__n6982 ), .ZN(_f_permutation__n3815 ) );
  NAND2_X2 _f_permutation__U5873  ( .A1(_f_permutation__round_out[1571]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6979 ) );
  NAND2_X2 _f_permutation__U5872  ( .A1(_f_permutation__n7171 ), .A2(out[475]), 
        .ZN(_f_permutation__n6980 ) );
  NAND2_X2 _f_permutation__U5871  ( .A1(_f_permutation__n6979 ), .A2(
        _f_permutation__n6980 ), .ZN(_f_permutation__n3816 ) );
  NAND2_X2 _f_permutation__U5870  ( .A1(_f_permutation__round_out[1570]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6977 ) );
  NAND2_X2 _f_permutation__U5869  ( .A1(_f_permutation__n7171 ), .A2(out[474]), 
        .ZN(_f_permutation__n6978 ) );
  NAND2_X2 _f_permutation__U5868  ( .A1(_f_permutation__n6977 ), .A2(
        _f_permutation__n6978 ), .ZN(_f_permutation__n3817 ) );
  NAND2_X2 _f_permutation__U5867  ( .A1(_f_permutation__round_out[1569]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6975 ) );
  NAND2_X2 _f_permutation__U5866  ( .A1(_f_permutation__n7171 ), .A2(out[473]), 
        .ZN(_f_permutation__n6976 ) );
  NAND2_X2 _f_permutation__U5865  ( .A1(_f_permutation__n6975 ), .A2(
        _f_permutation__n6976 ), .ZN(_f_permutation__n3818 ) );
  NAND2_X2 _f_permutation__U5864  ( .A1(_f_permutation__round_out[1568]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6973 ) );
  NAND2_X2 _f_permutation__U5863  ( .A1(_f_permutation__n7171 ), .A2(out[472]), 
        .ZN(_f_permutation__n6974 ) );
  NAND2_X2 _f_permutation__U5862  ( .A1(_f_permutation__n6973 ), .A2(
        _f_permutation__n6974 ), .ZN(_f_permutation__n3819 ) );
  NAND2_X2 _f_permutation__U5861  ( .A1(_f_permutation__round_out[1567]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6971 ) );
  NAND2_X2 _f_permutation__U5860  ( .A1(_f_permutation__n7171 ), .A2(out[487]), 
        .ZN(_f_permutation__n6972 ) );
  NAND2_X2 _f_permutation__U5859  ( .A1(_f_permutation__n6971 ), .A2(
        _f_permutation__n6972 ), .ZN(_f_permutation__n3820 ) );
  NAND2_X2 _f_permutation__U5858  ( .A1(_f_permutation__round_out[1566]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6969 ) );
  NAND2_X2 _f_permutation__U5857  ( .A1(_f_permutation__n7172 ), .A2(out[486]), 
        .ZN(_f_permutation__n6970 ) );
  NAND2_X2 _f_permutation__U5856  ( .A1(_f_permutation__n6969 ), .A2(
        _f_permutation__n6970 ), .ZN(_f_permutation__n3821 ) );
  NAND2_X2 _f_permutation__U5855  ( .A1(_f_permutation__round_out[1565]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6967 ) );
  NAND2_X2 _f_permutation__U5854  ( .A1(_f_permutation__n7172 ), .A2(out[485]), 
        .ZN(_f_permutation__n6968 ) );
  NAND2_X2 _f_permutation__U5853  ( .A1(_f_permutation__n6967 ), .A2(
        _f_permutation__n6968 ), .ZN(_f_permutation__n3822 ) );
  NAND2_X2 _f_permutation__U5852  ( .A1(_f_permutation__round_out[1564]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6965 ) );
  NAND2_X2 _f_permutation__U5851  ( .A1(_f_permutation__n7172 ), .A2(out[484]), 
        .ZN(_f_permutation__n6966 ) );
  NAND2_X2 _f_permutation__U5850  ( .A1(_f_permutation__n6965 ), .A2(
        _f_permutation__n6966 ), .ZN(_f_permutation__n3823 ) );
  NAND2_X2 _f_permutation__U5849  ( .A1(_f_permutation__round_out[1563]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6963 ) );
  NAND2_X2 _f_permutation__U5848  ( .A1(_f_permutation__n7172 ), .A2(out[483]), 
        .ZN(_f_permutation__n6964 ) );
  NAND2_X2 _f_permutation__U5847  ( .A1(_f_permutation__n6963 ), .A2(
        _f_permutation__n6964 ), .ZN(_f_permutation__n3824 ) );
  NAND2_X2 _f_permutation__U5846  ( .A1(_f_permutation__round_out[1562]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6961 ) );
  NAND2_X2 _f_permutation__U5845  ( .A1(_f_permutation__n7172 ), .A2(out[482]), 
        .ZN(_f_permutation__n6962 ) );
  NAND2_X2 _f_permutation__U5844  ( .A1(_f_permutation__n6961 ), .A2(
        _f_permutation__n6962 ), .ZN(_f_permutation__n3825 ) );
  NAND2_X2 _f_permutation__U5843  ( .A1(_f_permutation__round_out[1561]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6959 ) );
  NAND2_X2 _f_permutation__U5842  ( .A1(_f_permutation__n7172 ), .A2(out[481]), 
        .ZN(_f_permutation__n6960 ) );
  NAND2_X2 _f_permutation__U5841  ( .A1(_f_permutation__n6959 ), .A2(
        _f_permutation__n6960 ), .ZN(_f_permutation__n3826 ) );
  NAND2_X2 _f_permutation__U5840  ( .A1(_f_permutation__round_out[1560]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6957 ) );
  NAND2_X2 _f_permutation__U5839  ( .A1(_f_permutation__n7172 ), .A2(out[480]), 
        .ZN(_f_permutation__n6958 ) );
  NAND2_X2 _f_permutation__U5838  ( .A1(_f_permutation__n6957 ), .A2(
        _f_permutation__n6958 ), .ZN(_f_permutation__n3827 ) );
  NAND2_X2 _f_permutation__U5837  ( .A1(_f_permutation__round_out[1559]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6955 ) );
  NAND2_X2 _f_permutation__U5836  ( .A1(_f_permutation__n7172 ), .A2(out[495]), 
        .ZN(_f_permutation__n6956 ) );
  NAND2_X2 _f_permutation__U5835  ( .A1(_f_permutation__n6955 ), .A2(
        _f_permutation__n6956 ), .ZN(_f_permutation__n3828 ) );
  NAND2_X2 _f_permutation__U5834  ( .A1(_f_permutation__round_out[1558]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6953 ) );
  NAND2_X2 _f_permutation__U5833  ( .A1(_f_permutation__n7172 ), .A2(out[494]), 
        .ZN(_f_permutation__n6954 ) );
  NAND2_X2 _f_permutation__U5832  ( .A1(_f_permutation__n6953 ), .A2(
        _f_permutation__n6954 ), .ZN(_f_permutation__n3829 ) );
  NAND2_X2 _f_permutation__U5831  ( .A1(_f_permutation__round_out[1557]), 
        .A2(_f_permutation__n7109 ), .ZN(_f_permutation__n6951 ) );
  NAND2_X2 _f_permutation__U5830  ( .A1(_f_permutation__n7172 ), .A2(out[493]), 
        .ZN(_f_permutation__n6952 ) );
  NAND2_X2 _f_permutation__U5829  ( .A1(_f_permutation__n6951 ), .A2(
        _f_permutation__n6952 ), .ZN(_f_permutation__n3830 ) );
  NAND2_X2 _f_permutation__U5828  ( .A1(_f_permutation__round_out[1556]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6949 ) );
  NAND2_X2 _f_permutation__U5827  ( .A1(_f_permutation__n7172 ), .A2(out[492]), 
        .ZN(_f_permutation__n6950 ) );
  NAND2_X2 _f_permutation__U5826  ( .A1(_f_permutation__n6949 ), .A2(
        _f_permutation__n6950 ), .ZN(_f_permutation__n3831 ) );
  NAND2_X2 _f_permutation__U5825  ( .A1(_f_permutation__round_out[1555]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6947 ) );
  NAND2_X2 _f_permutation__U5824  ( .A1(_f_permutation__n7173 ), .A2(out[491]), 
        .ZN(_f_permutation__n6948 ) );
  NAND2_X2 _f_permutation__U5823  ( .A1(_f_permutation__n6947 ), .A2(
        _f_permutation__n6948 ), .ZN(_f_permutation__n3832 ) );
  NAND2_X2 _f_permutation__U5822  ( .A1(_f_permutation__round_out[1554]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6945 ) );
  NAND2_X2 _f_permutation__U5821  ( .A1(_f_permutation__n7173 ), .A2(out[490]), 
        .ZN(_f_permutation__n6946 ) );
  NAND2_X2 _f_permutation__U5820  ( .A1(_f_permutation__n6945 ), .A2(
        _f_permutation__n6946 ), .ZN(_f_permutation__n3833 ) );
  NAND2_X2 _f_permutation__U5819  ( .A1(_f_permutation__round_out[1553]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6943 ) );
  NAND2_X2 _f_permutation__U5818  ( .A1(_f_permutation__n7173 ), .A2(out[489]), 
        .ZN(_f_permutation__n6944 ) );
  NAND2_X2 _f_permutation__U5817  ( .A1(_f_permutation__n6943 ), .A2(
        _f_permutation__n6944 ), .ZN(_f_permutation__n3834 ) );
  NAND2_X2 _f_permutation__U5816  ( .A1(_f_permutation__round_out[1552]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6941 ) );
  NAND2_X2 _f_permutation__U5815  ( .A1(_f_permutation__n7173 ), .A2(out[488]), 
        .ZN(_f_permutation__n6942 ) );
  NAND2_X2 _f_permutation__U5814  ( .A1(_f_permutation__n6941 ), .A2(
        _f_permutation__n6942 ), .ZN(_f_permutation__n3835 ) );
  NAND2_X2 _f_permutation__U5813  ( .A1(_f_permutation__round_out[1551]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6939 ) );
  NAND2_X2 _f_permutation__U5812  ( .A1(_f_permutation__n7173 ), .A2(out[503]), 
        .ZN(_f_permutation__n6940 ) );
  NAND2_X2 _f_permutation__U5811  ( .A1(_f_permutation__n6939 ), .A2(
        _f_permutation__n6940 ), .ZN(_f_permutation__n3836 ) );
  NAND2_X2 _f_permutation__U5810  ( .A1(_f_permutation__round_out[1550]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6937 ) );
  NAND2_X2 _f_permutation__U5809  ( .A1(_f_permutation__n7173 ), .A2(out[502]), 
        .ZN(_f_permutation__n6938 ) );
  NAND2_X2 _f_permutation__U5808  ( .A1(_f_permutation__n6937 ), .A2(
        _f_permutation__n6938 ), .ZN(_f_permutation__n3837 ) );
  NAND2_X2 _f_permutation__U5807  ( .A1(_f_permutation__round_out[1549]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6935 ) );
  NAND2_X2 _f_permutation__U5806  ( .A1(_f_permutation__n7173 ), .A2(out[501]), 
        .ZN(_f_permutation__n6936 ) );
  NAND2_X2 _f_permutation__U5805  ( .A1(_f_permutation__n6935 ), .A2(
        _f_permutation__n6936 ), .ZN(_f_permutation__n3838 ) );
  NAND2_X2 _f_permutation__U5804  ( .A1(_f_permutation__round_out[1548]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6933 ) );
  NAND2_X2 _f_permutation__U5803  ( .A1(_f_permutation__n7173 ), .A2(out[500]), 
        .ZN(_f_permutation__n6934 ) );
  NAND2_X2 _f_permutation__U5802  ( .A1(_f_permutation__n6933 ), .A2(
        _f_permutation__n6934 ), .ZN(_f_permutation__n3839 ) );
  NAND2_X2 _f_permutation__U5801  ( .A1(_f_permutation__round_out[1547]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6931 ) );
  NAND2_X2 _f_permutation__U5800  ( .A1(_f_permutation__n7173 ), .A2(out[499]), 
        .ZN(_f_permutation__n6932 ) );
  NAND2_X2 _f_permutation__U5799  ( .A1(_f_permutation__n6931 ), .A2(
        _f_permutation__n6932 ), .ZN(_f_permutation__n3840 ) );
  NAND2_X2 _f_permutation__U5798  ( .A1(_f_permutation__round_out[1546]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6929 ) );
  NAND2_X2 _f_permutation__U5797  ( .A1(_f_permutation__n7173 ), .A2(out[498]), 
        .ZN(_f_permutation__n6930 ) );
  NAND2_X2 _f_permutation__U5796  ( .A1(_f_permutation__n6929 ), .A2(
        _f_permutation__n6930 ), .ZN(_f_permutation__n3841 ) );
  NAND2_X2 _f_permutation__U5795  ( .A1(_f_permutation__round_out[1545]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6927 ) );
  NAND2_X2 _f_permutation__U5794  ( .A1(_f_permutation__n7173 ), .A2(out[497]), 
        .ZN(_f_permutation__n6928 ) );
  NAND2_X2 _f_permutation__U5793  ( .A1(_f_permutation__n6927 ), .A2(
        _f_permutation__n6928 ), .ZN(_f_permutation__n3842 ) );
  NAND2_X2 _f_permutation__U5792  ( .A1(_f_permutation__round_out[1544]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6925 ) );
  NAND2_X2 _f_permutation__U5791  ( .A1(_f_permutation__n7174 ), .A2(out[496]), 
        .ZN(_f_permutation__n6926 ) );
  NAND2_X2 _f_permutation__U5790  ( .A1(_f_permutation__n6925 ), .A2(
        _f_permutation__n6926 ), .ZN(_f_permutation__n3843 ) );
  NAND2_X2 _f_permutation__U5789  ( .A1(_f_permutation__round_out[1543]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6923 ) );
  NAND2_X2 _f_permutation__U5788  ( .A1(_f_permutation__n7174 ), .A2(out[511]), 
        .ZN(_f_permutation__n6924 ) );
  NAND2_X2 _f_permutation__U5787  ( .A1(_f_permutation__n6923 ), .A2(
        _f_permutation__n6924 ), .ZN(_f_permutation__n3844 ) );
  NAND2_X2 _f_permutation__U5786  ( .A1(_f_permutation__round_out[1542]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6921 ) );
  NAND2_X2 _f_permutation__U5785  ( .A1(_f_permutation__n7174 ), .A2(out[510]), 
        .ZN(_f_permutation__n6922 ) );
  NAND2_X2 _f_permutation__U5784  ( .A1(_f_permutation__n6921 ), .A2(
        _f_permutation__n6922 ), .ZN(_f_permutation__n3845 ) );
  NAND2_X2 _f_permutation__U5783  ( .A1(_f_permutation__round_out[1541]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6919 ) );
  NAND2_X2 _f_permutation__U5782  ( .A1(_f_permutation__n7174 ), .A2(out[509]), 
        .ZN(_f_permutation__n6920 ) );
  NAND2_X2 _f_permutation__U5781  ( .A1(_f_permutation__n6919 ), .A2(
        _f_permutation__n6920 ), .ZN(_f_permutation__n3846 ) );
  NAND2_X2 _f_permutation__U5780  ( .A1(_f_permutation__round_out[1540]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6917 ) );
  NAND2_X2 _f_permutation__U5779  ( .A1(_f_permutation__n7174 ), .A2(out[508]), 
        .ZN(_f_permutation__n6918 ) );
  NAND2_X2 _f_permutation__U5778  ( .A1(_f_permutation__n6917 ), .A2(
        _f_permutation__n6918 ), .ZN(_f_permutation__n3847 ) );
  NAND2_X2 _f_permutation__U5777  ( .A1(_f_permutation__round_out[1539]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6915 ) );
  NAND2_X2 _f_permutation__U5776  ( .A1(_f_permutation__n7174 ), .A2(out[507]), 
        .ZN(_f_permutation__n6916 ) );
  NAND2_X2 _f_permutation__U5775  ( .A1(_f_permutation__n6915 ), .A2(
        _f_permutation__n6916 ), .ZN(_f_permutation__n3848 ) );
  NAND2_X2 _f_permutation__U5774  ( .A1(_f_permutation__round_out[1538]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6913 ) );
  NAND2_X2 _f_permutation__U5773  ( .A1(_f_permutation__n7174 ), .A2(out[506]), 
        .ZN(_f_permutation__n6914 ) );
  NAND2_X2 _f_permutation__U5772  ( .A1(_f_permutation__n6913 ), .A2(
        _f_permutation__n6914 ), .ZN(_f_permutation__n3849 ) );
  NAND2_X2 _f_permutation__U5771  ( .A1(_f_permutation__round_out[1537]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6911 ) );
  NAND2_X2 _f_permutation__U5770  ( .A1(_f_permutation__n7174 ), .A2(out[505]), 
        .ZN(_f_permutation__n6912 ) );
  NAND2_X2 _f_permutation__U5769  ( .A1(_f_permutation__n6911 ), .A2(
        _f_permutation__n6912 ), .ZN(_f_permutation__n3850 ) );
  NAND2_X2 _f_permutation__U5768  ( .A1(_f_permutation__round_out[1536]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6909 ) );
  NAND2_X2 _f_permutation__U5767  ( .A1(_f_permutation__n7174 ), .A2(out[504]), 
        .ZN(_f_permutation__n6910 ) );
  NAND2_X2 _f_permutation__U5766  ( .A1(_f_permutation__n6909 ), .A2(
        _f_permutation__n6910 ), .ZN(_f_permutation__n3851 ) );
  NAND2_X2 _f_permutation__U5765  ( .A1(_f_permutation__round_out[1535]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6907 ) );
  NAND2_X2 _f_permutation__U5764  ( .A1(_f_permutation__n7174 ), .A2(out[391]), 
        .ZN(_f_permutation__n6908 ) );
  NAND2_X2 _f_permutation__U5763  ( .A1(_f_permutation__n6907 ), .A2(
        _f_permutation__n6908 ), .ZN(_f_permutation__n3852 ) );
  NAND2_X2 _f_permutation__U5762  ( .A1(_f_permutation__round_out[1534]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6905 ) );
  NAND2_X2 _f_permutation__U5761  ( .A1(_f_permutation__n7174 ), .A2(out[390]), 
        .ZN(_f_permutation__n6906 ) );
  NAND2_X2 _f_permutation__U5760  ( .A1(_f_permutation__n6905 ), .A2(
        _f_permutation__n6906 ), .ZN(_f_permutation__n3853 ) );
  NAND2_X2 _f_permutation__U5759  ( .A1(_f_permutation__round_out[1533]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6903 ) );
  NAND2_X2 _f_permutation__U5758  ( .A1(_f_permutation__n7175 ), .A2(out[389]), 
        .ZN(_f_permutation__n6904 ) );
  NAND2_X2 _f_permutation__U5757  ( .A1(_f_permutation__n6903 ), .A2(
        _f_permutation__n6904 ), .ZN(_f_permutation__n3854 ) );
  NAND2_X2 _f_permutation__U5756  ( .A1(_f_permutation__round_out[1532]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6901 ) );
  NAND2_X2 _f_permutation__U5755  ( .A1(_f_permutation__n7175 ), .A2(out[388]), 
        .ZN(_f_permutation__n6902 ) );
  NAND2_X2 _f_permutation__U5754  ( .A1(_f_permutation__n6901 ), .A2(
        _f_permutation__n6902 ), .ZN(_f_permutation__n3855 ) );
  NAND2_X2 _f_permutation__U5753  ( .A1(_f_permutation__round_out[1531]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6899 ) );
  NAND2_X2 _f_permutation__U5752  ( .A1(_f_permutation__n7175 ), .A2(out[387]), 
        .ZN(_f_permutation__n6900 ) );
  NAND2_X2 _f_permutation__U5751  ( .A1(_f_permutation__n6899 ), .A2(
        _f_permutation__n6900 ), .ZN(_f_permutation__n3856 ) );
  NAND2_X2 _f_permutation__U5750  ( .A1(_f_permutation__round_out[1530]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6897 ) );
  NAND2_X2 _f_permutation__U5749  ( .A1(_f_permutation__n7175 ), .A2(out[386]), 
        .ZN(_f_permutation__n6898 ) );
  NAND2_X2 _f_permutation__U5748  ( .A1(_f_permutation__n6897 ), .A2(
        _f_permutation__n6898 ), .ZN(_f_permutation__n3857 ) );
  NAND2_X2 _f_permutation__U5747  ( .A1(_f_permutation__round_out[1529]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6895 ) );
  NAND2_X2 _f_permutation__U5746  ( .A1(_f_permutation__n7175 ), .A2(out[385]), 
        .ZN(_f_permutation__n6896 ) );
  NAND2_X2 _f_permutation__U5745  ( .A1(_f_permutation__n6895 ), .A2(
        _f_permutation__n6896 ), .ZN(_f_permutation__n3858 ) );
  NAND2_X2 _f_permutation__U5744  ( .A1(_f_permutation__round_out[1528]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6893 ) );
  NAND2_X2 _f_permutation__U5743  ( .A1(_f_permutation__n7175 ), .A2(out[384]), 
        .ZN(_f_permutation__n6894 ) );
  NAND2_X2 _f_permutation__U5742  ( .A1(_f_permutation__n6893 ), .A2(
        _f_permutation__n6894 ), .ZN(_f_permutation__n3859 ) );
  NAND2_X2 _f_permutation__U5741  ( .A1(_f_permutation__round_out[1527]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6891 ) );
  NAND2_X2 _f_permutation__U5740  ( .A1(_f_permutation__n7175 ), .A2(out[399]), 
        .ZN(_f_permutation__n6892 ) );
  NAND2_X2 _f_permutation__U5739  ( .A1(_f_permutation__n6891 ), .A2(
        _f_permutation__n6892 ), .ZN(_f_permutation__n3860 ) );
  NAND2_X2 _f_permutation__U5738  ( .A1(_f_permutation__round_out[1526]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6889 ) );
  NAND2_X2 _f_permutation__U5737  ( .A1(_f_permutation__n7175 ), .A2(out[398]), 
        .ZN(_f_permutation__n6890 ) );
  NAND2_X2 _f_permutation__U5736  ( .A1(_f_permutation__n6889 ), .A2(
        _f_permutation__n6890 ), .ZN(_f_permutation__n3861 ) );
  NAND2_X2 _f_permutation__U5735  ( .A1(_f_permutation__round_out[1525]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6887 ) );
  NAND2_X2 _f_permutation__U5734  ( .A1(_f_permutation__n7175 ), .A2(out[397]), 
        .ZN(_f_permutation__n6888 ) );
  NAND2_X2 _f_permutation__U5733  ( .A1(_f_permutation__n6887 ), .A2(
        _f_permutation__n6888 ), .ZN(_f_permutation__n3862 ) );
  NAND2_X2 _f_permutation__U5732  ( .A1(_f_permutation__round_out[1524]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6885 ) );
  NAND2_X2 _f_permutation__U5731  ( .A1(_f_permutation__n7175 ), .A2(out[396]), 
        .ZN(_f_permutation__n6886 ) );
  NAND2_X2 _f_permutation__U5730  ( .A1(_f_permutation__n6885 ), .A2(
        _f_permutation__n6886 ), .ZN(_f_permutation__n3863 ) );
  NAND2_X2 _f_permutation__U5729  ( .A1(_f_permutation__round_out[1523]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6883 ) );
  NAND2_X2 _f_permutation__U5728  ( .A1(_f_permutation__n7175 ), .A2(out[395]), 
        .ZN(_f_permutation__n6884 ) );
  NAND2_X2 _f_permutation__U5727  ( .A1(_f_permutation__n6883 ), .A2(
        _f_permutation__n6884 ), .ZN(_f_permutation__n3864 ) );
  NAND2_X2 _f_permutation__U5726  ( .A1(_f_permutation__round_out[1522]), 
        .A2(_f_permutation__n7107 ), .ZN(_f_permutation__n6881 ) );
  NAND2_X2 _f_permutation__U5725  ( .A1(_f_permutation__n7176 ), .A2(out[394]), 
        .ZN(_f_permutation__n6882 ) );
  NAND2_X2 _f_permutation__U5724  ( .A1(_f_permutation__n6881 ), .A2(
        _f_permutation__n6882 ), .ZN(_f_permutation__n3865 ) );
  NAND2_X2 _f_permutation__U5723  ( .A1(_f_permutation__round_out[1521]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6879 ) );
  NAND2_X2 _f_permutation__U5722  ( .A1(_f_permutation__n7176 ), .A2(out[393]), 
        .ZN(_f_permutation__n6880 ) );
  NAND2_X2 _f_permutation__U5721  ( .A1(_f_permutation__n6879 ), .A2(
        _f_permutation__n6880 ), .ZN(_f_permutation__n3866 ) );
  NAND2_X2 _f_permutation__U5720  ( .A1(_f_permutation__round_out[1520]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6877 ) );
  NAND2_X2 _f_permutation__U5719  ( .A1(_f_permutation__n7176 ), .A2(out[392]), 
        .ZN(_f_permutation__n6878 ) );
  NAND2_X2 _f_permutation__U5718  ( .A1(_f_permutation__n6877 ), .A2(
        _f_permutation__n6878 ), .ZN(_f_permutation__n3867 ) );
  NAND2_X2 _f_permutation__U5717  ( .A1(_f_permutation__round_out[1519]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6875 ) );
  NAND2_X2 _f_permutation__U5716  ( .A1(_f_permutation__n7176 ), .A2(out[407]), 
        .ZN(_f_permutation__n6876 ) );
  NAND2_X2 _f_permutation__U5715  ( .A1(_f_permutation__n6875 ), .A2(
        _f_permutation__n6876 ), .ZN(_f_permutation__n3868 ) );
  NAND2_X2 _f_permutation__U5714  ( .A1(_f_permutation__round_out[1518]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6873 ) );
  NAND2_X2 _f_permutation__U5713  ( .A1(_f_permutation__n7176 ), .A2(out[406]), 
        .ZN(_f_permutation__n6874 ) );
  NAND2_X2 _f_permutation__U5712  ( .A1(_f_permutation__n6873 ), .A2(
        _f_permutation__n6874 ), .ZN(_f_permutation__n3869 ) );
  NAND2_X2 _f_permutation__U5711  ( .A1(_f_permutation__round_out[1517]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6871 ) );
  NAND2_X2 _f_permutation__U5710  ( .A1(_f_permutation__n7176 ), .A2(out[405]), 
        .ZN(_f_permutation__n6872 ) );
  NAND2_X2 _f_permutation__U5709  ( .A1(_f_permutation__n6871 ), .A2(
        _f_permutation__n6872 ), .ZN(_f_permutation__n3870 ) );
  NAND2_X2 _f_permutation__U5708  ( .A1(_f_permutation__round_out[1516]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6869 ) );
  NAND2_X2 _f_permutation__U5707  ( .A1(_f_permutation__n7176 ), .A2(out[404]), 
        .ZN(_f_permutation__n6870 ) );
  NAND2_X2 _f_permutation__U5706  ( .A1(_f_permutation__n6869 ), .A2(
        _f_permutation__n6870 ), .ZN(_f_permutation__n3871 ) );
  NAND2_X2 _f_permutation__U5705  ( .A1(_f_permutation__round_out[1515]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6867 ) );
  NAND2_X2 _f_permutation__U5704  ( .A1(_f_permutation__n7176 ), .A2(out[403]), 
        .ZN(_f_permutation__n6868 ) );
  NAND2_X2 _f_permutation__U5703  ( .A1(_f_permutation__n6867 ), .A2(
        _f_permutation__n6868 ), .ZN(_f_permutation__n3872 ) );
  NAND2_X2 _f_permutation__U5702  ( .A1(_f_permutation__round_out[1514]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6865 ) );
  NAND2_X2 _f_permutation__U5701  ( .A1(_f_permutation__n7176 ), .A2(out[402]), 
        .ZN(_f_permutation__n6866 ) );
  NAND2_X2 _f_permutation__U5700  ( .A1(_f_permutation__n6865 ), .A2(
        _f_permutation__n6866 ), .ZN(_f_permutation__n3873 ) );
  NAND2_X2 _f_permutation__U5699  ( .A1(_f_permutation__round_out[1513]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6863 ) );
  NAND2_X2 _f_permutation__U5698  ( .A1(_f_permutation__n7176 ), .A2(out[401]), 
        .ZN(_f_permutation__n6864 ) );
  NAND2_X2 _f_permutation__U5697  ( .A1(_f_permutation__n6863 ), .A2(
        _f_permutation__n6864 ), .ZN(_f_permutation__n3874 ) );
  NAND2_X2 _f_permutation__U5696  ( .A1(_f_permutation__round_out[1512]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6861 ) );
  NAND2_X2 _f_permutation__U5695  ( .A1(_f_permutation__n7176 ), .A2(out[400]), 
        .ZN(_f_permutation__n6862 ) );
  NAND2_X2 _f_permutation__U5694  ( .A1(_f_permutation__n6861 ), .A2(
        _f_permutation__n6862 ), .ZN(_f_permutation__n3875 ) );
  NAND2_X2 _f_permutation__U5693  ( .A1(_f_permutation__round_out[1511]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6859 ) );
  NAND2_X2 _f_permutation__U5692  ( .A1(_f_permutation__n7177 ), .A2(out[415]), 
        .ZN(_f_permutation__n6860 ) );
  NAND2_X2 _f_permutation__U5691  ( .A1(_f_permutation__n6859 ), .A2(
        _f_permutation__n6860 ), .ZN(_f_permutation__n3876 ) );
  NAND2_X2 _f_permutation__U5690  ( .A1(_f_permutation__round_out[1510]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6857 ) );
  NAND2_X2 _f_permutation__U5689  ( .A1(_f_permutation__n7177 ), .A2(out[414]), 
        .ZN(_f_permutation__n6858 ) );
  NAND2_X2 _f_permutation__U5688  ( .A1(_f_permutation__n6857 ), .A2(
        _f_permutation__n6858 ), .ZN(_f_permutation__n3877 ) );
  NAND2_X2 _f_permutation__U5687  ( .A1(_f_permutation__round_out[1509]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6855 ) );
  NAND2_X2 _f_permutation__U5686  ( .A1(_f_permutation__n7177 ), .A2(out[413]), 
        .ZN(_f_permutation__n6856 ) );
  NAND2_X2 _f_permutation__U5685  ( .A1(_f_permutation__n6855 ), .A2(
        _f_permutation__n6856 ), .ZN(_f_permutation__n3878 ) );
  NAND2_X2 _f_permutation__U5684  ( .A1(_f_permutation__round_out[1508]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6853 ) );
  NAND2_X2 _f_permutation__U5683  ( .A1(_f_permutation__n7177 ), .A2(out[412]), 
        .ZN(_f_permutation__n6854 ) );
  NAND2_X2 _f_permutation__U5682  ( .A1(_f_permutation__n6853 ), .A2(
        _f_permutation__n6854 ), .ZN(_f_permutation__n3879 ) );
  NAND2_X2 _f_permutation__U5681  ( .A1(_f_permutation__round_out[1507]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6851 ) );
  NAND2_X2 _f_permutation__U5680  ( .A1(_f_permutation__n7177 ), .A2(out[411]), 
        .ZN(_f_permutation__n6852 ) );
  NAND2_X2 _f_permutation__U5679  ( .A1(_f_permutation__n6851 ), .A2(
        _f_permutation__n6852 ), .ZN(_f_permutation__n3880 ) );
  NAND2_X2 _f_permutation__U5678  ( .A1(_f_permutation__round_out[1506]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6849 ) );
  NAND2_X2 _f_permutation__U5677  ( .A1(_f_permutation__n7177 ), .A2(out[410]), 
        .ZN(_f_permutation__n6850 ) );
  NAND2_X2 _f_permutation__U5676  ( .A1(_f_permutation__n6849 ), .A2(
        _f_permutation__n6850 ), .ZN(_f_permutation__n3881 ) );
  NAND2_X2 _f_permutation__U5675  ( .A1(_f_permutation__round_out[1505]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6847 ) );
  NAND2_X2 _f_permutation__U5674  ( .A1(_f_permutation__n7177 ), .A2(out[409]), 
        .ZN(_f_permutation__n6848 ) );
  NAND2_X2 _f_permutation__U5673  ( .A1(_f_permutation__n6847 ), .A2(
        _f_permutation__n6848 ), .ZN(_f_permutation__n3882 ) );
  NAND2_X2 _f_permutation__U5672  ( .A1(_f_permutation__round_out[1504]), 
        .A2(_f_permutation__n7106 ), .ZN(_f_permutation__n6845 ) );
  NAND2_X2 _f_permutation__U5671  ( .A1(_f_permutation__n7177 ), .A2(out[408]), 
        .ZN(_f_permutation__n6846 ) );
  NAND2_X2 _f_permutation__U5670  ( .A1(_f_permutation__n6845 ), .A2(
        _f_permutation__n6846 ), .ZN(_f_permutation__n3883 ) );
  NAND2_X2 _f_permutation__U5669  ( .A1(_f_permutation__round_out[1503]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6843 ) );
  NAND2_X2 _f_permutation__U5668  ( .A1(_f_permutation__n7177 ), .A2(out[423]), 
        .ZN(_f_permutation__n6844 ) );
  NAND2_X2 _f_permutation__U5667  ( .A1(_f_permutation__n6843 ), .A2(
        _f_permutation__n6844 ), .ZN(_f_permutation__n3884 ) );
  NAND2_X2 _f_permutation__U5666  ( .A1(_f_permutation__round_out[1502]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6841 ) );
  NAND2_X2 _f_permutation__U5665  ( .A1(_f_permutation__n7177 ), .A2(out[422]), 
        .ZN(_f_permutation__n6842 ) );
  NAND2_X2 _f_permutation__U5664  ( .A1(_f_permutation__n6841 ), .A2(
        _f_permutation__n6842 ), .ZN(_f_permutation__n3885 ) );
  NAND2_X2 _f_permutation__U5663  ( .A1(_f_permutation__round_out[1501]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6839 ) );
  NAND2_X2 _f_permutation__U5662  ( .A1(_f_permutation__n7177 ), .A2(out[421]), 
        .ZN(_f_permutation__n6840 ) );
  NAND2_X2 _f_permutation__U5661  ( .A1(_f_permutation__n6839 ), .A2(
        _f_permutation__n6840 ), .ZN(_f_permutation__n3886 ) );
  NAND2_X2 _f_permutation__U5660  ( .A1(_f_permutation__round_out[1500]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6837 ) );
  NAND2_X2 _f_permutation__U5659  ( .A1(_f_permutation__n7178 ), .A2(out[420]), 
        .ZN(_f_permutation__n6838 ) );
  NAND2_X2 _f_permutation__U5658  ( .A1(_f_permutation__n6837 ), .A2(
        _f_permutation__n6838 ), .ZN(_f_permutation__n3887 ) );
  NAND2_X2 _f_permutation__U5657  ( .A1(_f_permutation__round_out[1499]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6835 ) );
  NAND2_X2 _f_permutation__U5656  ( .A1(_f_permutation__n7178 ), .A2(out[419]), 
        .ZN(_f_permutation__n6836 ) );
  NAND2_X2 _f_permutation__U5655  ( .A1(_f_permutation__n6835 ), .A2(
        _f_permutation__n6836 ), .ZN(_f_permutation__n3888 ) );
  NAND2_X2 _f_permutation__U5654  ( .A1(_f_permutation__round_out[1498]), 
        .A2(_f_permutation__n7108 ), .ZN(_f_permutation__n6833 ) );
  NAND2_X2 _f_permutation__U5653  ( .A1(_f_permutation__n7178 ), .A2(out[418]), 
        .ZN(_f_permutation__n6834 ) );
  NAND2_X2 _f_permutation__U5652  ( .A1(_f_permutation__n6833 ), .A2(
        _f_permutation__n6834 ), .ZN(_f_permutation__n3889 ) );
  NAND2_X2 _f_permutation__U5651  ( .A1(_f_permutation__round_out[1497]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6831 ) );
  NAND2_X2 _f_permutation__U5650  ( .A1(_f_permutation__n7178 ), .A2(out[417]), 
        .ZN(_f_permutation__n6832 ) );
  NAND2_X2 _f_permutation__U5649  ( .A1(_f_permutation__n6831 ), .A2(
        _f_permutation__n6832 ), .ZN(_f_permutation__n3890 ) );
  NAND2_X2 _f_permutation__U5648  ( .A1(_f_permutation__round_out[1496]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6829 ) );
  NAND2_X2 _f_permutation__U5647  ( .A1(_f_permutation__n7178 ), .A2(out[416]), 
        .ZN(_f_permutation__n6830 ) );
  NAND2_X2 _f_permutation__U5646  ( .A1(_f_permutation__n6829 ), .A2(
        _f_permutation__n6830 ), .ZN(_f_permutation__n3891 ) );
  NAND2_X2 _f_permutation__U5645  ( .A1(_f_permutation__round_out[1495]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6827 ) );
  NAND2_X2 _f_permutation__U5644  ( .A1(_f_permutation__n7178 ), .A2(out[431]), 
        .ZN(_f_permutation__n6828 ) );
  NAND2_X2 _f_permutation__U5643  ( .A1(_f_permutation__n6827 ), .A2(
        _f_permutation__n6828 ), .ZN(_f_permutation__n3892 ) );
  NAND2_X2 _f_permutation__U5642  ( .A1(_f_permutation__round_out[1494]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6825 ) );
  NAND2_X2 _f_permutation__U5641  ( .A1(_f_permutation__n7178 ), .A2(out[430]), 
        .ZN(_f_permutation__n6826 ) );
  NAND2_X2 _f_permutation__U5640  ( .A1(_f_permutation__n6825 ), .A2(
        _f_permutation__n6826 ), .ZN(_f_permutation__n3893 ) );
  NAND2_X2 _f_permutation__U5639  ( .A1(_f_permutation__round_out[1493]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6823 ) );
  NAND2_X2 _f_permutation__U5638  ( .A1(_f_permutation__n7178 ), .A2(out[429]), 
        .ZN(_f_permutation__n6824 ) );
  NAND2_X2 _f_permutation__U5637  ( .A1(_f_permutation__n6823 ), .A2(
        _f_permutation__n6824 ), .ZN(_f_permutation__n3894 ) );
  NAND2_X2 _f_permutation__U5636  ( .A1(_f_permutation__round_out[1492]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6821 ) );
  NAND2_X2 _f_permutation__U5635  ( .A1(_f_permutation__n7178 ), .A2(out[428]), 
        .ZN(_f_permutation__n6822 ) );
  NAND2_X2 _f_permutation__U5634  ( .A1(_f_permutation__n6821 ), .A2(
        _f_permutation__n6822 ), .ZN(_f_permutation__n3895 ) );
  NAND2_X2 _f_permutation__U5633  ( .A1(_f_permutation__round_out[1491]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6819 ) );
  NAND2_X2 _f_permutation__U5632  ( .A1(_f_permutation__n7178 ), .A2(out[427]), 
        .ZN(_f_permutation__n6820 ) );
  NAND2_X2 _f_permutation__U5631  ( .A1(_f_permutation__n6819 ), .A2(
        _f_permutation__n6820 ), .ZN(_f_permutation__n3896 ) );
  NAND2_X2 _f_permutation__U5630  ( .A1(_f_permutation__round_out[1490]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6817 ) );
  NAND2_X2 _f_permutation__U5629  ( .A1(_f_permutation__n7178 ), .A2(out[426]), 
        .ZN(_f_permutation__n6818 ) );
  NAND2_X2 _f_permutation__U5628  ( .A1(_f_permutation__n6817 ), .A2(
        _f_permutation__n6818 ), .ZN(_f_permutation__n3897 ) );
  NAND2_X2 _f_permutation__U5627  ( .A1(_f_permutation__round_out[1489]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6815 ) );
  NAND2_X2 _f_permutation__U5626  ( .A1(_f_permutation__n7179 ), .A2(out[425]), 
        .ZN(_f_permutation__n6816 ) );
  NAND2_X2 _f_permutation__U5625  ( .A1(_f_permutation__n6815 ), .A2(
        _f_permutation__n6816 ), .ZN(_f_permutation__n3898 ) );
  NAND2_X2 _f_permutation__U5624  ( .A1(_f_permutation__round_out[1488]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6813 ) );
  NAND2_X2 _f_permutation__U5623  ( .A1(_f_permutation__n7179 ), .A2(out[424]), 
        .ZN(_f_permutation__n6814 ) );
  NAND2_X2 _f_permutation__U5622  ( .A1(_f_permutation__n6813 ), .A2(
        _f_permutation__n6814 ), .ZN(_f_permutation__n3899 ) );
  NAND2_X2 _f_permutation__U5621  ( .A1(_f_permutation__round_out[1487]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6811 ) );
  NAND2_X2 _f_permutation__U5620  ( .A1(_f_permutation__n7179 ), .A2(out[439]), 
        .ZN(_f_permutation__n6812 ) );
  NAND2_X2 _f_permutation__U5619  ( .A1(_f_permutation__n6811 ), .A2(
        _f_permutation__n6812 ), .ZN(_f_permutation__n3900 ) );
  NAND2_X2 _f_permutation__U5618  ( .A1(_f_permutation__round_out[1486]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6809 ) );
  NAND2_X2 _f_permutation__U5617  ( .A1(_f_permutation__n7179 ), .A2(out[438]), 
        .ZN(_f_permutation__n6810 ) );
  NAND2_X2 _f_permutation__U5616  ( .A1(_f_permutation__n6809 ), .A2(
        _f_permutation__n6810 ), .ZN(_f_permutation__n3901 ) );
  NAND2_X2 _f_permutation__U5615  ( .A1(_f_permutation__round_out[1485]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6807 ) );
  NAND2_X2 _f_permutation__U5614  ( .A1(_f_permutation__n7179 ), .A2(out[437]), 
        .ZN(_f_permutation__n6808 ) );
  NAND2_X2 _f_permutation__U5613  ( .A1(_f_permutation__n6807 ), .A2(
        _f_permutation__n6808 ), .ZN(_f_permutation__n3902 ) );
  NAND2_X2 _f_permutation__U5612  ( .A1(_f_permutation__round_out[1484]), 
        .A2(_f_permutation__n7116 ), .ZN(_f_permutation__n6805 ) );
  NAND2_X2 _f_permutation__U5611  ( .A1(_f_permutation__n7179 ), .A2(out[436]), 
        .ZN(_f_permutation__n6806 ) );
  NAND2_X2 _f_permutation__U5610  ( .A1(_f_permutation__n6805 ), .A2(
        _f_permutation__n6806 ), .ZN(_f_permutation__n3903 ) );
  NAND2_X2 _f_permutation__U5609  ( .A1(_f_permutation__round_out[1483]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6803 ) );
  NAND2_X2 _f_permutation__U5608  ( .A1(_f_permutation__n7179 ), .A2(out[435]), 
        .ZN(_f_permutation__n6804 ) );
  NAND2_X2 _f_permutation__U5607  ( .A1(_f_permutation__n6803 ), .A2(
        _f_permutation__n6804 ), .ZN(_f_permutation__n3904 ) );
  NAND2_X2 _f_permutation__U5606  ( .A1(_f_permutation__round_out[1482]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6801 ) );
  NAND2_X2 _f_permutation__U5605  ( .A1(_f_permutation__n7179 ), .A2(out[434]), 
        .ZN(_f_permutation__n6802 ) );
  NAND2_X2 _f_permutation__U5604  ( .A1(_f_permutation__n6801 ), .A2(
        _f_permutation__n6802 ), .ZN(_f_permutation__n3905 ) );
  NAND2_X2 _f_permutation__U5603  ( .A1(_f_permutation__round_out[1481]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6799 ) );
  NAND2_X2 _f_permutation__U5602  ( .A1(_f_permutation__n7179 ), .A2(out[433]), 
        .ZN(_f_permutation__n6800 ) );
  NAND2_X2 _f_permutation__U5601  ( .A1(_f_permutation__n6799 ), .A2(
        _f_permutation__n6800 ), .ZN(_f_permutation__n3906 ) );
  NAND2_X2 _f_permutation__U5600  ( .A1(_f_permutation__round_out[1480]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6797 ) );
  NAND2_X2 _f_permutation__U5599  ( .A1(_f_permutation__n7179 ), .A2(out[432]), 
        .ZN(_f_permutation__n6798 ) );
  NAND2_X2 _f_permutation__U5598  ( .A1(_f_permutation__n6797 ), .A2(
        _f_permutation__n6798 ), .ZN(_f_permutation__n3907 ) );
  NAND2_X2 _f_permutation__U5597  ( .A1(_f_permutation__round_out[1479]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6795 ) );
  NAND2_X2 _f_permutation__U5596  ( .A1(_f_permutation__n7179 ), .A2(out[447]), 
        .ZN(_f_permutation__n6796 ) );
  NAND2_X2 _f_permutation__U5595  ( .A1(_f_permutation__n6795 ), .A2(
        _f_permutation__n6796 ), .ZN(_f_permutation__n3908 ) );
  NAND2_X2 _f_permutation__U5594  ( .A1(_f_permutation__round_out[1478]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6793 ) );
  NAND2_X2 _f_permutation__U5593  ( .A1(_f_permutation__n7180 ), .A2(out[446]), 
        .ZN(_f_permutation__n6794 ) );
  NAND2_X2 _f_permutation__U5592  ( .A1(_f_permutation__n6793 ), .A2(
        _f_permutation__n6794 ), .ZN(_f_permutation__n3909 ) );
  NAND2_X2 _f_permutation__U5591  ( .A1(_f_permutation__round_out[1477]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6791 ) );
  NAND2_X2 _f_permutation__U5590  ( .A1(_f_permutation__n7180 ), .A2(out[445]), 
        .ZN(_f_permutation__n6792 ) );
  NAND2_X2 _f_permutation__U5589  ( .A1(_f_permutation__n6791 ), .A2(
        _f_permutation__n6792 ), .ZN(_f_permutation__n3910 ) );
  NAND2_X2 _f_permutation__U5588  ( .A1(_f_permutation__round_out[1476]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6789 ) );
  NAND2_X2 _f_permutation__U5587  ( .A1(_f_permutation__n7180 ), .A2(out[444]), 
        .ZN(_f_permutation__n6790 ) );
  NAND2_X2 _f_permutation__U5586  ( .A1(_f_permutation__n6789 ), .A2(
        _f_permutation__n6790 ), .ZN(_f_permutation__n3911 ) );
  NAND2_X2 _f_permutation__U5585  ( .A1(_f_permutation__round_out[1475]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6787 ) );
  NAND2_X2 _f_permutation__U5584  ( .A1(_f_permutation__n7180 ), .A2(out[443]), 
        .ZN(_f_permutation__n6788 ) );
  NAND2_X2 _f_permutation__U5583  ( .A1(_f_permutation__n6787 ), .A2(
        _f_permutation__n6788 ), .ZN(_f_permutation__n3912 ) );
  NAND2_X2 _f_permutation__U5582  ( .A1(_f_permutation__round_out[1474]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6785 ) );
  NAND2_X2 _f_permutation__U5581  ( .A1(_f_permutation__n7180 ), .A2(out[442]), 
        .ZN(_f_permutation__n6786 ) );
  NAND2_X2 _f_permutation__U5580  ( .A1(_f_permutation__n6785 ), .A2(
        _f_permutation__n6786 ), .ZN(_f_permutation__n3913 ) );
  NAND2_X2 _f_permutation__U5579  ( .A1(_f_permutation__round_out[1473]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6783 ) );
  NAND2_X2 _f_permutation__U5578  ( .A1(_f_permutation__n7180 ), .A2(out[441]), 
        .ZN(_f_permutation__n6784 ) );
  NAND2_X2 _f_permutation__U5577  ( .A1(_f_permutation__n6783 ), .A2(
        _f_permutation__n6784 ), .ZN(_f_permutation__n3914 ) );
  NAND2_X2 _f_permutation__U5576  ( .A1(_f_permutation__round_out[1472]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6781 ) );
  NAND2_X2 _f_permutation__U5575  ( .A1(_f_permutation__n7180 ), .A2(out[440]), 
        .ZN(_f_permutation__n6782 ) );
  NAND2_X2 _f_permutation__U5574  ( .A1(_f_permutation__n6781 ), .A2(
        _f_permutation__n6782 ), .ZN(_f_permutation__n3915 ) );
  NAND2_X2 _f_permutation__U5573  ( .A1(_f_permutation__round_out[1471]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6779 ) );
  NAND2_X2 _f_permutation__U5572  ( .A1(_f_permutation__n7180 ), .A2(out[327]), 
        .ZN(_f_permutation__n6780 ) );
  NAND2_X2 _f_permutation__U5571  ( .A1(_f_permutation__n6779 ), .A2(
        _f_permutation__n6780 ), .ZN(_f_permutation__n3916 ) );
  NAND2_X2 _f_permutation__U5570  ( .A1(_f_permutation__round_out[1470]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6777 ) );
  NAND2_X2 _f_permutation__U5569  ( .A1(_f_permutation__n7180 ), .A2(out[326]), 
        .ZN(_f_permutation__n6778 ) );
  NAND2_X2 _f_permutation__U5568  ( .A1(_f_permutation__n6777 ), .A2(
        _f_permutation__n6778 ), .ZN(_f_permutation__n3917 ) );
  NAND2_X2 _f_permutation__U5567  ( .A1(_f_permutation__round_out[1469]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6775 ) );
  NAND2_X2 _f_permutation__U5566  ( .A1(_f_permutation__n7180 ), .A2(out[325]), 
        .ZN(_f_permutation__n6776 ) );
  NAND2_X2 _f_permutation__U5565  ( .A1(_f_permutation__n6775 ), .A2(
        _f_permutation__n6776 ), .ZN(_f_permutation__n3918 ) );
  NAND2_X2 _f_permutation__U5564  ( .A1(_f_permutation__round_out[1468]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6773 ) );
  NAND2_X2 _f_permutation__U5563  ( .A1(_f_permutation__n7180 ), .A2(out[324]), 
        .ZN(_f_permutation__n6774 ) );
  NAND2_X2 _f_permutation__U5562  ( .A1(_f_permutation__n6773 ), .A2(
        _f_permutation__n6774 ), .ZN(_f_permutation__n3919 ) );
  NAND2_X2 _f_permutation__U5561  ( .A1(_f_permutation__round_out[1467]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6771 ) );
  NAND2_X2 _f_permutation__U5560  ( .A1(_f_permutation__n7181 ), .A2(out[323]), 
        .ZN(_f_permutation__n6772 ) );
  NAND2_X2 _f_permutation__U5559  ( .A1(_f_permutation__n6771 ), .A2(
        _f_permutation__n6772 ), .ZN(_f_permutation__n3920 ) );
  NAND2_X2 _f_permutation__U5558  ( .A1(_f_permutation__round_out[1466]), 
        .A2(_f_permutation__n7115 ), .ZN(_f_permutation__n6769 ) );
  NAND2_X2 _f_permutation__U5557  ( .A1(_f_permutation__n7181 ), .A2(out[322]), 
        .ZN(_f_permutation__n6770 ) );
  NAND2_X2 _f_permutation__U5556  ( .A1(_f_permutation__n6769 ), .A2(
        _f_permutation__n6770 ), .ZN(_f_permutation__n3921 ) );
  NAND2_X2 _f_permutation__U5555  ( .A1(_f_permutation__round_out[1465]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6767 ) );
  NAND2_X2 _f_permutation__U5554  ( .A1(_f_permutation__n7181 ), .A2(out[321]), 
        .ZN(_f_permutation__n6768 ) );
  NAND2_X2 _f_permutation__U5553  ( .A1(_f_permutation__n6767 ), .A2(
        _f_permutation__n6768 ), .ZN(_f_permutation__n3922 ) );
  NAND2_X2 _f_permutation__U5552  ( .A1(_f_permutation__round_out[1464]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6765 ) );
  NAND2_X2 _f_permutation__U5551  ( .A1(_f_permutation__n7181 ), .A2(out[320]), 
        .ZN(_f_permutation__n6766 ) );
  NAND2_X2 _f_permutation__U5550  ( .A1(_f_permutation__n6765 ), .A2(
        _f_permutation__n6766 ), .ZN(_f_permutation__n3923 ) );
  NAND2_X2 _f_permutation__U5549  ( .A1(_f_permutation__round_out[1463]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6763 ) );
  NAND2_X2 _f_permutation__U5548  ( .A1(_f_permutation__n7181 ), .A2(out[335]), 
        .ZN(_f_permutation__n6764 ) );
  NAND2_X2 _f_permutation__U5547  ( .A1(_f_permutation__n6763 ), .A2(
        _f_permutation__n6764 ), .ZN(_f_permutation__n3924 ) );
  NAND2_X2 _f_permutation__U5546  ( .A1(_f_permutation__round_out[1462]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6761 ) );
  NAND2_X2 _f_permutation__U5545  ( .A1(_f_permutation__n7181 ), .A2(out[334]), 
        .ZN(_f_permutation__n6762 ) );
  NAND2_X2 _f_permutation__U5544  ( .A1(_f_permutation__n6761 ), .A2(
        _f_permutation__n6762 ), .ZN(_f_permutation__n3925 ) );
  NAND2_X2 _f_permutation__U5543  ( .A1(_f_permutation__round_out[1461]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6759 ) );
  NAND2_X2 _f_permutation__U5542  ( .A1(_f_permutation__n7181 ), .A2(out[333]), 
        .ZN(_f_permutation__n6760 ) );
  NAND2_X2 _f_permutation__U5541  ( .A1(_f_permutation__n6759 ), .A2(
        _f_permutation__n6760 ), .ZN(_f_permutation__n3926 ) );
  NAND2_X2 _f_permutation__U5540  ( .A1(_f_permutation__round_out[1460]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6757 ) );
  NAND2_X2 _f_permutation__U5539  ( .A1(_f_permutation__n7181 ), .A2(out[332]), 
        .ZN(_f_permutation__n6758 ) );
  NAND2_X2 _f_permutation__U5538  ( .A1(_f_permutation__n6757 ), .A2(
        _f_permutation__n6758 ), .ZN(_f_permutation__n3927 ) );
  NAND2_X2 _f_permutation__U5537  ( .A1(_f_permutation__round_out[1459]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6755 ) );
  NAND2_X2 _f_permutation__U5536  ( .A1(_f_permutation__n7181 ), .A2(out[331]), 
        .ZN(_f_permutation__n6756 ) );
  NAND2_X2 _f_permutation__U5535  ( .A1(_f_permutation__n6755 ), .A2(
        _f_permutation__n6756 ), .ZN(_f_permutation__n3928 ) );
  NAND2_X2 _f_permutation__U5534  ( .A1(_f_permutation__round_out[1458]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6753 ) );
  NAND2_X2 _f_permutation__U5533  ( .A1(_f_permutation__n7181 ), .A2(out[330]), 
        .ZN(_f_permutation__n6754 ) );
  NAND2_X2 _f_permutation__U5532  ( .A1(_f_permutation__n6753 ), .A2(
        _f_permutation__n6754 ), .ZN(_f_permutation__n3929 ) );
  NAND2_X2 _f_permutation__U5531  ( .A1(_f_permutation__round_out[1457]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6751 ) );
  NAND2_X2 _f_permutation__U5530  ( .A1(_f_permutation__n7181 ), .A2(out[329]), 
        .ZN(_f_permutation__n6752 ) );
  NAND2_X2 _f_permutation__U5529  ( .A1(_f_permutation__n6751 ), .A2(
        _f_permutation__n6752 ), .ZN(_f_permutation__n3930 ) );
  NAND2_X2 _f_permutation__U5528  ( .A1(_f_permutation__round_out[1456]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6749 ) );
  NAND2_X2 _f_permutation__U5527  ( .A1(_f_permutation__n7182 ), .A2(out[328]), 
        .ZN(_f_permutation__n6750 ) );
  NAND2_X2 _f_permutation__U5526  ( .A1(_f_permutation__n6749 ), .A2(
        _f_permutation__n6750 ), .ZN(_f_permutation__n3931 ) );
  NAND2_X2 _f_permutation__U5525  ( .A1(_f_permutation__round_out[1455]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6747 ) );
  NAND2_X2 _f_permutation__U5524  ( .A1(_f_permutation__n7182 ), .A2(out[343]), 
        .ZN(_f_permutation__n6748 ) );
  NAND2_X2 _f_permutation__U5523  ( .A1(_f_permutation__n6747 ), .A2(
        _f_permutation__n6748 ), .ZN(_f_permutation__n3932 ) );
  NAND2_X2 _f_permutation__U5522  ( .A1(_f_permutation__round_out[1454]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6745 ) );
  NAND2_X2 _f_permutation__U5521  ( .A1(_f_permutation__n7182 ), .A2(out[342]), 
        .ZN(_f_permutation__n6746 ) );
  NAND2_X2 _f_permutation__U5520  ( .A1(_f_permutation__n6745 ), .A2(
        _f_permutation__n6746 ), .ZN(_f_permutation__n3933 ) );
  NAND2_X2 _f_permutation__U5519  ( .A1(_f_permutation__round_out[1453]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6743 ) );
  NAND2_X2 _f_permutation__U5518  ( .A1(_f_permutation__n7182 ), .A2(out[341]), 
        .ZN(_f_permutation__n6744 ) );
  NAND2_X2 _f_permutation__U5517  ( .A1(_f_permutation__n6743 ), .A2(
        _f_permutation__n6744 ), .ZN(_f_permutation__n3934 ) );
  NAND2_X2 _f_permutation__U5516  ( .A1(_f_permutation__round_out[1452]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6741 ) );
  NAND2_X2 _f_permutation__U5515  ( .A1(_f_permutation__n7182 ), .A2(out[340]), 
        .ZN(_f_permutation__n6742 ) );
  NAND2_X2 _f_permutation__U5514  ( .A1(_f_permutation__n6741 ), .A2(
        _f_permutation__n6742 ), .ZN(_f_permutation__n3935 ) );
  NAND2_X2 _f_permutation__U5513  ( .A1(_f_permutation__round_out[1451]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6739 ) );
  NAND2_X2 _f_permutation__U5512  ( .A1(_f_permutation__n7182 ), .A2(out[339]), 
        .ZN(_f_permutation__n6740 ) );
  NAND2_X2 _f_permutation__U5511  ( .A1(_f_permutation__n6739 ), .A2(
        _f_permutation__n6740 ), .ZN(_f_permutation__n3936 ) );
  NAND2_X2 _f_permutation__U5510  ( .A1(_f_permutation__round_out[1450]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6737 ) );
  NAND2_X2 _f_permutation__U5509  ( .A1(_f_permutation__n7182 ), .A2(out[338]), 
        .ZN(_f_permutation__n6738 ) );
  NAND2_X2 _f_permutation__U5508  ( .A1(_f_permutation__n6737 ), .A2(
        _f_permutation__n6738 ), .ZN(_f_permutation__n3937 ) );
  NAND2_X2 _f_permutation__U5507  ( .A1(_f_permutation__round_out[1449]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6735 ) );
  NAND2_X2 _f_permutation__U5506  ( .A1(_f_permutation__n7182 ), .A2(out[337]), 
        .ZN(_f_permutation__n6736 ) );
  NAND2_X2 _f_permutation__U5505  ( .A1(_f_permutation__n6735 ), .A2(
        _f_permutation__n6736 ), .ZN(_f_permutation__n3938 ) );
  NAND2_X2 _f_permutation__U5504  ( .A1(_f_permutation__round_out[1448]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6733 ) );
  NAND2_X2 _f_permutation__U5503  ( .A1(_f_permutation__n7182 ), .A2(out[336]), 
        .ZN(_f_permutation__n6734 ) );
  NAND2_X2 _f_permutation__U5502  ( .A1(_f_permutation__n6733 ), .A2(
        _f_permutation__n6734 ), .ZN(_f_permutation__n3939 ) );
  NAND2_X2 _f_permutation__U5501  ( .A1(_f_permutation__round_out[1447]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6731 ) );
  NAND2_X2 _f_permutation__U5500  ( .A1(_f_permutation__n7182 ), .A2(out[351]), 
        .ZN(_f_permutation__n6732 ) );
  NAND2_X2 _f_permutation__U5499  ( .A1(_f_permutation__n6731 ), .A2(
        _f_permutation__n6732 ), .ZN(_f_permutation__n3940 ) );
  NAND2_X2 _f_permutation__U5498  ( .A1(_f_permutation__round_out[1446]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6729 ) );
  NAND2_X2 _f_permutation__U5497  ( .A1(_f_permutation__n7182 ), .A2(out[350]), 
        .ZN(_f_permutation__n6730 ) );
  NAND2_X2 _f_permutation__U5496  ( .A1(_f_permutation__n6729 ), .A2(
        _f_permutation__n6730 ), .ZN(_f_permutation__n3941 ) );
  NAND2_X2 _f_permutation__U5495  ( .A1(_f_permutation__round_out[1445]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6727 ) );
  NAND2_X2 _f_permutation__U5494  ( .A1(_f_permutation__n7183 ), .A2(out[349]), 
        .ZN(_f_permutation__n6728 ) );
  NAND2_X2 _f_permutation__U5493  ( .A1(_f_permutation__n6727 ), .A2(
        _f_permutation__n6728 ), .ZN(_f_permutation__n3942 ) );
  NAND2_X2 _f_permutation__U5492  ( .A1(_f_permutation__round_out[1444]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6725 ) );
  NAND2_X2 _f_permutation__U5491  ( .A1(_f_permutation__n7183 ), .A2(out[348]), 
        .ZN(_f_permutation__n6726 ) );
  NAND2_X2 _f_permutation__U5490  ( .A1(_f_permutation__n6725 ), .A2(
        _f_permutation__n6726 ), .ZN(_f_permutation__n3943 ) );
  NAND2_X2 _f_permutation__U5489  ( .A1(_f_permutation__round_out[1443]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6723 ) );
  NAND2_X2 _f_permutation__U5488  ( .A1(_f_permutation__n7183 ), .A2(out[347]), 
        .ZN(_f_permutation__n6724 ) );
  NAND2_X2 _f_permutation__U5487  ( .A1(_f_permutation__n6723 ), .A2(
        _f_permutation__n6724 ), .ZN(_f_permutation__n3944 ) );
  NAND2_X2 _f_permutation__U5486  ( .A1(_f_permutation__round_out[1442]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6721 ) );
  NAND2_X2 _f_permutation__U5485  ( .A1(_f_permutation__n7183 ), .A2(out[346]), 
        .ZN(_f_permutation__n6722 ) );
  NAND2_X2 _f_permutation__U5484  ( .A1(_f_permutation__n6721 ), .A2(
        _f_permutation__n6722 ), .ZN(_f_permutation__n3945 ) );
  NAND2_X2 _f_permutation__U5483  ( .A1(_f_permutation__round_out[1441]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6719 ) );
  NAND2_X2 _f_permutation__U5482  ( .A1(_f_permutation__n7183 ), .A2(out[345]), 
        .ZN(_f_permutation__n6720 ) );
  NAND2_X2 _f_permutation__U5481  ( .A1(_f_permutation__n6719 ), .A2(
        _f_permutation__n6720 ), .ZN(_f_permutation__n3946 ) );
  NAND2_X2 _f_permutation__U5480  ( .A1(_f_permutation__round_out[1440]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6717 ) );
  NAND2_X2 _f_permutation__U5479  ( .A1(_f_permutation__n7183 ), .A2(out[344]), 
        .ZN(_f_permutation__n6718 ) );
  NAND2_X2 _f_permutation__U5478  ( .A1(_f_permutation__n6717 ), .A2(
        _f_permutation__n6718 ), .ZN(_f_permutation__n3947 ) );
  NAND2_X2 _f_permutation__U5477  ( .A1(_f_permutation__round_out[1439]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6715 ) );
  NAND2_X2 _f_permutation__U5476  ( .A1(_f_permutation__n7183 ), .A2(out[359]), 
        .ZN(_f_permutation__n6716 ) );
  NAND2_X2 _f_permutation__U5475  ( .A1(_f_permutation__n6715 ), .A2(
        _f_permutation__n6716 ), .ZN(_f_permutation__n3948 ) );
  NAND2_X2 _f_permutation__U5474  ( .A1(_f_permutation__round_out[1438]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6713 ) );
  NAND2_X2 _f_permutation__U5473  ( .A1(_f_permutation__n7183 ), .A2(out[358]), 
        .ZN(_f_permutation__n6714 ) );
  NAND2_X2 _f_permutation__U5472  ( .A1(_f_permutation__n6713 ), .A2(
        _f_permutation__n6714 ), .ZN(_f_permutation__n3949 ) );
  NAND2_X2 _f_permutation__U5471  ( .A1(_f_permutation__round_out[1437]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6711 ) );
  NAND2_X2 _f_permutation__U5470  ( .A1(_f_permutation__n7183 ), .A2(out[357]), 
        .ZN(_f_permutation__n6712 ) );
  NAND2_X2 _f_permutation__U5469  ( .A1(_f_permutation__n6711 ), .A2(
        _f_permutation__n6712 ), .ZN(_f_permutation__n3950 ) );
  NAND2_X2 _f_permutation__U5468  ( .A1(_f_permutation__round_out[1436]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6709 ) );
  NAND2_X2 _f_permutation__U5467  ( .A1(_f_permutation__n7183 ), .A2(out[356]), 
        .ZN(_f_permutation__n6710 ) );
  NAND2_X2 _f_permutation__U5466  ( .A1(_f_permutation__n6709 ), .A2(
        _f_permutation__n6710 ), .ZN(_f_permutation__n3951 ) );
  NAND2_X2 _f_permutation__U5465  ( .A1(_f_permutation__round_out[1435]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6707 ) );
  NAND2_X2 _f_permutation__U5464  ( .A1(_f_permutation__n7183 ), .A2(out[355]), 
        .ZN(_f_permutation__n6708 ) );
  NAND2_X2 _f_permutation__U5463  ( .A1(_f_permutation__n6707 ), .A2(
        _f_permutation__n6708 ), .ZN(_f_permutation__n3952 ) );
  NAND2_X2 _f_permutation__U5462  ( .A1(_f_permutation__round_out[1434]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6705 ) );
  NAND2_X2 _f_permutation__U5461  ( .A1(_f_permutation__n7184 ), .A2(out[354]), 
        .ZN(_f_permutation__n6706 ) );
  NAND2_X2 _f_permutation__U5460  ( .A1(_f_permutation__n6705 ), .A2(
        _f_permutation__n6706 ), .ZN(_f_permutation__n3953 ) );
  NAND2_X2 _f_permutation__U5459  ( .A1(_f_permutation__round_out[1433]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6703 ) );
  NAND2_X2 _f_permutation__U5458  ( .A1(_f_permutation__n7184 ), .A2(out[353]), 
        .ZN(_f_permutation__n6704 ) );
  NAND2_X2 _f_permutation__U5457  ( .A1(_f_permutation__n6703 ), .A2(
        _f_permutation__n6704 ), .ZN(_f_permutation__n3954 ) );
  NAND2_X2 _f_permutation__U5456  ( .A1(_f_permutation__round_out[1432]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6701 ) );
  NAND2_X2 _f_permutation__U5455  ( .A1(_f_permutation__n7184 ), .A2(out[352]), 
        .ZN(_f_permutation__n6702 ) );
  NAND2_X2 _f_permutation__U5454  ( .A1(_f_permutation__n6701 ), .A2(
        _f_permutation__n6702 ), .ZN(_f_permutation__n3955 ) );
  NAND2_X2 _f_permutation__U5453  ( .A1(_f_permutation__round_out[1431]), 
        .A2(_f_permutation__n7113 ), .ZN(_f_permutation__n6699 ) );
  NAND2_X2 _f_permutation__U5452  ( .A1(_f_permutation__n7184 ), .A2(out[367]), 
        .ZN(_f_permutation__n6700 ) );
  NAND2_X2 _f_permutation__U5451  ( .A1(_f_permutation__n6699 ), .A2(
        _f_permutation__n6700 ), .ZN(_f_permutation__n3956 ) );
  NAND2_X2 _f_permutation__U5450  ( .A1(_f_permutation__round_out[1430]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6697 ) );
  NAND2_X2 _f_permutation__U5449  ( .A1(_f_permutation__n7184 ), .A2(out[366]), 
        .ZN(_f_permutation__n6698 ) );
  NAND2_X2 _f_permutation__U5448  ( .A1(_f_permutation__n6697 ), .A2(
        _f_permutation__n6698 ), .ZN(_f_permutation__n3957 ) );
  NAND2_X2 _f_permutation__U5447  ( .A1(_f_permutation__round_out[1429]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6695 ) );
  NAND2_X2 _f_permutation__U5446  ( .A1(_f_permutation__n7184 ), .A2(out[365]), 
        .ZN(_f_permutation__n6696 ) );
  NAND2_X2 _f_permutation__U5445  ( .A1(_f_permutation__n6695 ), .A2(
        _f_permutation__n6696 ), .ZN(_f_permutation__n3958 ) );
  NAND2_X2 _f_permutation__U5444  ( .A1(_f_permutation__round_out[1428]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6693 ) );
  NAND2_X2 _f_permutation__U5443  ( .A1(_f_permutation__n7184 ), .A2(out[364]), 
        .ZN(_f_permutation__n6694 ) );
  NAND2_X2 _f_permutation__U5442  ( .A1(_f_permutation__n6693 ), .A2(
        _f_permutation__n6694 ), .ZN(_f_permutation__n3959 ) );
  NAND2_X2 _f_permutation__U5441  ( .A1(_f_permutation__round_out[1427]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6691 ) );
  NAND2_X2 _f_permutation__U5440  ( .A1(_f_permutation__n7184 ), .A2(out[363]), 
        .ZN(_f_permutation__n6692 ) );
  NAND2_X2 _f_permutation__U5439  ( .A1(_f_permutation__n6691 ), .A2(
        _f_permutation__n6692 ), .ZN(_f_permutation__n3960 ) );
  NAND2_X2 _f_permutation__U5438  ( .A1(_f_permutation__round_out[1426]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6689 ) );
  NAND2_X2 _f_permutation__U5437  ( .A1(_f_permutation__n7184 ), .A2(out[362]), 
        .ZN(_f_permutation__n6690 ) );
  NAND2_X2 _f_permutation__U5436  ( .A1(_f_permutation__n6689 ), .A2(
        _f_permutation__n6690 ), .ZN(_f_permutation__n3961 ) );
  NAND2_X2 _f_permutation__U5435  ( .A1(_f_permutation__round_out[1425]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6687 ) );
  NAND2_X2 _f_permutation__U5434  ( .A1(_f_permutation__n7184 ), .A2(out[361]), 
        .ZN(_f_permutation__n6688 ) );
  NAND2_X2 _f_permutation__U5433  ( .A1(_f_permutation__n6687 ), .A2(
        _f_permutation__n6688 ), .ZN(_f_permutation__n3962 ) );
  NAND2_X2 _f_permutation__U5432  ( .A1(_f_permutation__round_out[1424]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6685 ) );
  NAND2_X2 _f_permutation__U5431  ( .A1(_f_permutation__n7184 ), .A2(out[360]), 
        .ZN(_f_permutation__n6686 ) );
  NAND2_X2 _f_permutation__U5430  ( .A1(_f_permutation__n6685 ), .A2(
        _f_permutation__n6686 ), .ZN(_f_permutation__n3963 ) );
  NAND2_X2 _f_permutation__U5429  ( .A1(_f_permutation__round_out[1423]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6683 ) );
  NAND2_X2 _f_permutation__U5428  ( .A1(_f_permutation__n7185 ), .A2(out[375]), 
        .ZN(_f_permutation__n6684 ) );
  NAND2_X2 _f_permutation__U5427  ( .A1(_f_permutation__n6683 ), .A2(
        _f_permutation__n6684 ), .ZN(_f_permutation__n3964 ) );
  NAND2_X2 _f_permutation__U5426  ( .A1(_f_permutation__round_out[1422]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6681 ) );
  NAND2_X2 _f_permutation__U5425  ( .A1(_f_permutation__n7185 ), .A2(out[374]), 
        .ZN(_f_permutation__n6682 ) );
  NAND2_X2 _f_permutation__U5424  ( .A1(_f_permutation__n6681 ), .A2(
        _f_permutation__n6682 ), .ZN(_f_permutation__n3965 ) );
  NAND2_X2 _f_permutation__U5423  ( .A1(_f_permutation__round_out[1421]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6679 ) );
  NAND2_X2 _f_permutation__U5422  ( .A1(_f_permutation__n7185 ), .A2(out[373]), 
        .ZN(_f_permutation__n6680 ) );
  NAND2_X2 _f_permutation__U5421  ( .A1(_f_permutation__n6679 ), .A2(
        _f_permutation__n6680 ), .ZN(_f_permutation__n3966 ) );
  NAND2_X2 _f_permutation__U5420  ( .A1(_f_permutation__round_out[1420]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6677 ) );
  NAND2_X2 _f_permutation__U5419  ( .A1(_f_permutation__n7185 ), .A2(out[372]), 
        .ZN(_f_permutation__n6678 ) );
  NAND2_X2 _f_permutation__U5418  ( .A1(_f_permutation__n6677 ), .A2(
        _f_permutation__n6678 ), .ZN(_f_permutation__n3967 ) );
  NAND2_X2 _f_permutation__U5417  ( .A1(_f_permutation__round_out[1419]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6675 ) );
  NAND2_X2 _f_permutation__U5416  ( .A1(_f_permutation__n7185 ), .A2(out[371]), 
        .ZN(_f_permutation__n6676 ) );
  NAND2_X2 _f_permutation__U5415  ( .A1(_f_permutation__n6675 ), .A2(
        _f_permutation__n6676 ), .ZN(_f_permutation__n3968 ) );
  NAND2_X2 _f_permutation__U5414  ( .A1(_f_permutation__round_out[1418]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6673 ) );
  NAND2_X2 _f_permutation__U5413  ( .A1(_f_permutation__n7185 ), .A2(out[370]), 
        .ZN(_f_permutation__n6674 ) );
  NAND2_X2 _f_permutation__U5412  ( .A1(_f_permutation__n6673 ), .A2(
        _f_permutation__n6674 ), .ZN(_f_permutation__n3969 ) );
  NAND2_X2 _f_permutation__U5411  ( .A1(_f_permutation__round_out[1417]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6671 ) );
  NAND2_X2 _f_permutation__U5410  ( .A1(_f_permutation__n7185 ), .A2(out[369]), 
        .ZN(_f_permutation__n6672 ) );
  NAND2_X2 _f_permutation__U5409  ( .A1(_f_permutation__n6671 ), .A2(
        _f_permutation__n6672 ), .ZN(_f_permutation__n3970 ) );
  NAND2_X2 _f_permutation__U5408  ( .A1(_f_permutation__round_out[1416]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6669 ) );
  NAND2_X2 _f_permutation__U5407  ( .A1(_f_permutation__n7185 ), .A2(out[368]), 
        .ZN(_f_permutation__n6670 ) );
  NAND2_X2 _f_permutation__U5406  ( .A1(_f_permutation__n6669 ), .A2(
        _f_permutation__n6670 ), .ZN(_f_permutation__n3971 ) );
  NAND2_X2 _f_permutation__U5405  ( .A1(_f_permutation__round_out[1415]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6667 ) );
  NAND2_X2 _f_permutation__U5404  ( .A1(_f_permutation__n7185 ), .A2(out[383]), 
        .ZN(_f_permutation__n6668 ) );
  NAND2_X2 _f_permutation__U5403  ( .A1(_f_permutation__n6667 ), .A2(
        _f_permutation__n6668 ), .ZN(_f_permutation__n3972 ) );
  NAND2_X2 _f_permutation__U5402  ( .A1(_f_permutation__round_out[1414]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6665 ) );
  NAND2_X2 _f_permutation__U5401  ( .A1(_f_permutation__n7185 ), .A2(out[382]), 
        .ZN(_f_permutation__n6666 ) );
  NAND2_X2 _f_permutation__U5400  ( .A1(_f_permutation__n6665 ), .A2(
        _f_permutation__n6666 ), .ZN(_f_permutation__n3973 ) );
  NAND2_X2 _f_permutation__U5399  ( .A1(_f_permutation__round_out[1413]), 
        .A2(_f_permutation__n7112 ), .ZN(_f_permutation__n6663 ) );
  NAND2_X2 _f_permutation__U5398  ( .A1(_f_permutation__n7185 ), .A2(out[381]), 
        .ZN(_f_permutation__n6664 ) );
  NAND2_X2 _f_permutation__U5397  ( .A1(_f_permutation__n6663 ), .A2(
        _f_permutation__n6664 ), .ZN(_f_permutation__n3974 ) );
  NAND2_X2 _f_permutation__U5396  ( .A1(_f_permutation__round_out[1412]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6661 ) );
  NAND2_X2 _f_permutation__U5395  ( .A1(_f_permutation__n7186 ), .A2(out[380]), 
        .ZN(_f_permutation__n6662 ) );
  NAND2_X2 _f_permutation__U5394  ( .A1(_f_permutation__n6661 ), .A2(
        _f_permutation__n6662 ), .ZN(_f_permutation__n3975 ) );
  NAND2_X2 _f_permutation__U5393  ( .A1(_f_permutation__round_out[1411]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6659 ) );
  NAND2_X2 _f_permutation__U5392  ( .A1(_f_permutation__n7186 ), .A2(out[379]), 
        .ZN(_f_permutation__n6660 ) );
  NAND2_X2 _f_permutation__U5391  ( .A1(_f_permutation__n6659 ), .A2(
        _f_permutation__n6660 ), .ZN(_f_permutation__n3976 ) );
  NAND2_X2 _f_permutation__U5390  ( .A1(_f_permutation__round_out[1410]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6657 ) );
  NAND2_X2 _f_permutation__U5389  ( .A1(_f_permutation__n7186 ), .A2(out[378]), 
        .ZN(_f_permutation__n6658 ) );
  NAND2_X2 _f_permutation__U5388  ( .A1(_f_permutation__n6657 ), .A2(
        _f_permutation__n6658 ), .ZN(_f_permutation__n3977 ) );
  NAND2_X2 _f_permutation__U5387  ( .A1(_f_permutation__round_out[1409]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6655 ) );
  NAND2_X2 _f_permutation__U5386  ( .A1(_f_permutation__n7186 ), .A2(out[377]), 
        .ZN(_f_permutation__n6656 ) );
  NAND2_X2 _f_permutation__U5385  ( .A1(_f_permutation__n6655 ), .A2(
        _f_permutation__n6656 ), .ZN(_f_permutation__n3978 ) );
  NAND2_X2 _f_permutation__U5384  ( .A1(_f_permutation__round_out[1408]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6653 ) );
  NAND2_X2 _f_permutation__U5383  ( .A1(_f_permutation__n7186 ), .A2(out[376]), 
        .ZN(_f_permutation__n6654 ) );
  NAND2_X2 _f_permutation__U5382  ( .A1(_f_permutation__n6653 ), .A2(
        _f_permutation__n6654 ), .ZN(_f_permutation__n3979 ) );
  NAND2_X2 _f_permutation__U5381  ( .A1(_f_permutation__round_out[1407]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6651 ) );
  NAND2_X2 _f_permutation__U5380  ( .A1(_f_permutation__n7186 ), .A2(out[263]), 
        .ZN(_f_permutation__n6652 ) );
  NAND2_X2 _f_permutation__U5379  ( .A1(_f_permutation__n6651 ), .A2(
        _f_permutation__n6652 ), .ZN(_f_permutation__n3980 ) );
  NAND2_X2 _f_permutation__U5378  ( .A1(_f_permutation__round_out[1406]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6649 ) );
  NAND2_X2 _f_permutation__U5377  ( .A1(_f_permutation__n7186 ), .A2(out[262]), 
        .ZN(_f_permutation__n6650 ) );
  NAND2_X2 _f_permutation__U5376  ( .A1(_f_permutation__n6649 ), .A2(
        _f_permutation__n6650 ), .ZN(_f_permutation__n3981 ) );
  NAND2_X2 _f_permutation__U5375  ( .A1(_f_permutation__round_out[1405]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6647 ) );
  NAND2_X2 _f_permutation__U5374  ( .A1(_f_permutation__n7186 ), .A2(out[261]), 
        .ZN(_f_permutation__n6648 ) );
  NAND2_X2 _f_permutation__U5373  ( .A1(_f_permutation__n6647 ), .A2(
        _f_permutation__n6648 ), .ZN(_f_permutation__n3982 ) );
  NAND2_X2 _f_permutation__U5372  ( .A1(_f_permutation__round_out[1404]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6645 ) );
  NAND2_X2 _f_permutation__U5371  ( .A1(_f_permutation__n7186 ), .A2(out[260]), 
        .ZN(_f_permutation__n6646 ) );
  NAND2_X2 _f_permutation__U5370  ( .A1(_f_permutation__n6645 ), .A2(
        _f_permutation__n6646 ), .ZN(_f_permutation__n3983 ) );
  NAND2_X2 _f_permutation__U5369  ( .A1(_f_permutation__round_out[1403]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6643 ) );
  NAND2_X2 _f_permutation__U5368  ( .A1(_f_permutation__n7186 ), .A2(out[259]), 
        .ZN(_f_permutation__n6644 ) );
  NAND2_X2 _f_permutation__U5367  ( .A1(_f_permutation__n6643 ), .A2(
        _f_permutation__n6644 ), .ZN(_f_permutation__n3984 ) );
  NAND2_X2 _f_permutation__U5366  ( .A1(_f_permutation__round_out[1402]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6641 ) );
  NAND2_X2 _f_permutation__U5365  ( .A1(_f_permutation__n7186 ), .A2(out[258]), 
        .ZN(_f_permutation__n6642 ) );
  NAND2_X2 _f_permutation__U5364  ( .A1(_f_permutation__n6641 ), .A2(
        _f_permutation__n6642 ), .ZN(_f_permutation__n3985 ) );
  NAND2_X2 _f_permutation__U5363  ( .A1(_f_permutation__round_out[1401]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6639 ) );
  NAND2_X2 _f_permutation__U5362  ( .A1(_f_permutation__n7187 ), .A2(out[257]), 
        .ZN(_f_permutation__n6640 ) );
  NAND2_X2 _f_permutation__U5361  ( .A1(_f_permutation__n6639 ), .A2(
        _f_permutation__n6640 ), .ZN(_f_permutation__n3986 ) );
  NAND2_X2 _f_permutation__U5360  ( .A1(_f_permutation__round_out[1400]), 
        .A2(_f_permutation__n7111 ), .ZN(_f_permutation__n6637 ) );
  NAND2_X2 _f_permutation__U5359  ( .A1(_f_permutation__n7187 ), .A2(out[256]), 
        .ZN(_f_permutation__n6638 ) );
  NAND2_X2 _f_permutation__U5358  ( .A1(_f_permutation__n6637 ), .A2(
        _f_permutation__n6638 ), .ZN(_f_permutation__n3987 ) );
  NAND2_X2 _f_permutation__U5357  ( .A1(_f_permutation__round_out[1399]), 
        .A2(_f_permutation__n7114 ), .ZN(_f_permutation__n6635 ) );
  NAND2_X2 _f_permutation__U5356  ( .A1(_f_permutation__n7187 ), .A2(out[271]), 
        .ZN(_f_permutation__n6636 ) );
  NAND2_X2 _f_permutation__U5355  ( .A1(_f_permutation__n6635 ), .A2(
        _f_permutation__n6636 ), .ZN(_f_permutation__n3988 ) );
  NAND2_X2 _f_permutation__U5354  ( .A1(_f_permutation__round_out[1398]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6633 ) );
  NAND2_X2 _f_permutation__U5353  ( .A1(_f_permutation__n7187 ), .A2(out[270]), 
        .ZN(_f_permutation__n6634 ) );
  NAND2_X2 _f_permutation__U5352  ( .A1(_f_permutation__n6633 ), .A2(
        _f_permutation__n6634 ), .ZN(_f_permutation__n3989 ) );
  NAND2_X2 _f_permutation__U5351  ( .A1(_f_permutation__round_out[1397]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6631 ) );
  NAND2_X2 _f_permutation__U5350  ( .A1(_f_permutation__n7187 ), .A2(out[269]), 
        .ZN(_f_permutation__n6632 ) );
  NAND2_X2 _f_permutation__U5349  ( .A1(_f_permutation__n6631 ), .A2(
        _f_permutation__n6632 ), .ZN(_f_permutation__n3990 ) );
  NAND2_X2 _f_permutation__U5348  ( .A1(_f_permutation__round_out[1396]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6629 ) );
  NAND2_X2 _f_permutation__U5347  ( .A1(_f_permutation__n7187 ), .A2(out[268]), 
        .ZN(_f_permutation__n6630 ) );
  NAND2_X2 _f_permutation__U5346  ( .A1(_f_permutation__n6629 ), .A2(
        _f_permutation__n6630 ), .ZN(_f_permutation__n3991 ) );
  NAND2_X2 _f_permutation__U5345  ( .A1(_f_permutation__round_out[1395]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6627 ) );
  NAND2_X2 _f_permutation__U5344  ( .A1(_f_permutation__n7187 ), .A2(out[267]), 
        .ZN(_f_permutation__n6628 ) );
  NAND2_X2 _f_permutation__U5343  ( .A1(_f_permutation__n6627 ), .A2(
        _f_permutation__n6628 ), .ZN(_f_permutation__n3992 ) );
  NAND2_X2 _f_permutation__U5342  ( .A1(_f_permutation__round_out[1394]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6625 ) );
  NAND2_X2 _f_permutation__U5341  ( .A1(_f_permutation__n7187 ), .A2(out[266]), 
        .ZN(_f_permutation__n6626 ) );
  NAND2_X2 _f_permutation__U5340  ( .A1(_f_permutation__n6625 ), .A2(
        _f_permutation__n6626 ), .ZN(_f_permutation__n3993 ) );
  NAND2_X2 _f_permutation__U5339  ( .A1(_f_permutation__round_out[1393]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6623 ) );
  NAND2_X2 _f_permutation__U5338  ( .A1(_f_permutation__n7187 ), .A2(out[265]), 
        .ZN(_f_permutation__n6624 ) );
  NAND2_X2 _f_permutation__U5337  ( .A1(_f_permutation__n6623 ), .A2(
        _f_permutation__n6624 ), .ZN(_f_permutation__n3994 ) );
  NAND2_X2 _f_permutation__U5336  ( .A1(_f_permutation__round_out[1392]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6621 ) );
  NAND2_X2 _f_permutation__U5335  ( .A1(_f_permutation__n7187 ), .A2(out[264]), 
        .ZN(_f_permutation__n6622 ) );
  NAND2_X2 _f_permutation__U5334  ( .A1(_f_permutation__n6621 ), .A2(
        _f_permutation__n6622 ), .ZN(_f_permutation__n3995 ) );
  NAND2_X2 _f_permutation__U5333  ( .A1(_f_permutation__round_out[1391]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6619 ) );
  NAND2_X2 _f_permutation__U5332  ( .A1(_f_permutation__n7187 ), .A2(out[279]), 
        .ZN(_f_permutation__n6620 ) );
  NAND2_X2 _f_permutation__U5331  ( .A1(_f_permutation__n6619 ), .A2(
        _f_permutation__n6620 ), .ZN(_f_permutation__n3996 ) );
  NAND2_X2 _f_permutation__U5330  ( .A1(_f_permutation__round_out[1390]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6617 ) );
  NAND2_X2 _f_permutation__U5329  ( .A1(_f_permutation__n7188 ), .A2(out[278]), 
        .ZN(_f_permutation__n6618 ) );
  NAND2_X2 _f_permutation__U5328  ( .A1(_f_permutation__n6617 ), .A2(
        _f_permutation__n6618 ), .ZN(_f_permutation__n3997 ) );
  NAND2_X2 _f_permutation__U5327  ( .A1(_f_permutation__round_out[1389]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6615 ) );
  NAND2_X2 _f_permutation__U5326  ( .A1(_f_permutation__n7188 ), .A2(out[277]), 
        .ZN(_f_permutation__n6616 ) );
  NAND2_X2 _f_permutation__U5325  ( .A1(_f_permutation__n6615 ), .A2(
        _f_permutation__n6616 ), .ZN(_f_permutation__n3998 ) );
  NAND2_X2 _f_permutation__U5324  ( .A1(_f_permutation__round_out[1388]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6613 ) );
  NAND2_X2 _f_permutation__U5323  ( .A1(_f_permutation__n7188 ), .A2(out[276]), 
        .ZN(_f_permutation__n6614 ) );
  NAND2_X2 _f_permutation__U5322  ( .A1(_f_permutation__n6613 ), .A2(
        _f_permutation__n6614 ), .ZN(_f_permutation__n3999 ) );
  NAND2_X2 _f_permutation__U5321  ( .A1(_f_permutation__round_out[1387]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6611 ) );
  NAND2_X2 _f_permutation__U5320  ( .A1(_f_permutation__n7188 ), .A2(out[275]), 
        .ZN(_f_permutation__n6612 ) );
  NAND2_X2 _f_permutation__U5319  ( .A1(_f_permutation__n6611 ), .A2(
        _f_permutation__n6612 ), .ZN(_f_permutation__n4000 ) );
  NAND2_X2 _f_permutation__U5318  ( .A1(_f_permutation__round_out[1386]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6609 ) );
  NAND2_X2 _f_permutation__U5317  ( .A1(_f_permutation__n7188 ), .A2(out[274]), 
        .ZN(_f_permutation__n6610 ) );
  NAND2_X2 _f_permutation__U5316  ( .A1(_f_permutation__n6609 ), .A2(
        _f_permutation__n6610 ), .ZN(_f_permutation__n4001 ) );
  NAND2_X2 _f_permutation__U5315  ( .A1(_f_permutation__round_out[1385]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6607 ) );
  NAND2_X2 _f_permutation__U5314  ( .A1(_f_permutation__n7188 ), .A2(out[273]), 
        .ZN(_f_permutation__n6608 ) );
  NAND2_X2 _f_permutation__U5313  ( .A1(_f_permutation__n6607 ), .A2(
        _f_permutation__n6608 ), .ZN(_f_permutation__n4002 ) );
  NAND2_X2 _f_permutation__U5312  ( .A1(_f_permutation__round_out[1384]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6605 ) );
  NAND2_X2 _f_permutation__U5311  ( .A1(_f_permutation__n7188 ), .A2(out[272]), 
        .ZN(_f_permutation__n6606 ) );
  NAND2_X2 _f_permutation__U5310  ( .A1(_f_permutation__n6605 ), .A2(
        _f_permutation__n6606 ), .ZN(_f_permutation__n4003 ) );
  NAND2_X2 _f_permutation__U5309  ( .A1(_f_permutation__round_out[1383]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6603 ) );
  NAND2_X2 _f_permutation__U5308  ( .A1(_f_permutation__n7188 ), .A2(out[287]), 
        .ZN(_f_permutation__n6604 ) );
  NAND2_X2 _f_permutation__U5307  ( .A1(_f_permutation__n6603 ), .A2(
        _f_permutation__n6604 ), .ZN(_f_permutation__n4004 ) );
  NAND2_X2 _f_permutation__U5306  ( .A1(_f_permutation__round_out[1382]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6601 ) );
  NAND2_X2 _f_permutation__U5305  ( .A1(_f_permutation__n7188 ), .A2(out[286]), 
        .ZN(_f_permutation__n6602 ) );
  NAND2_X2 _f_permutation__U5304  ( .A1(_f_permutation__n6601 ), .A2(
        _f_permutation__n6602 ), .ZN(_f_permutation__n4005 ) );
  NAND2_X2 _f_permutation__U5303  ( .A1(_f_permutation__round_out[1381]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6599 ) );
  NAND2_X2 _f_permutation__U5302  ( .A1(_f_permutation__n7188 ), .A2(out[285]), 
        .ZN(_f_permutation__n6600 ) );
  NAND2_X2 _f_permutation__U5301  ( .A1(_f_permutation__n6599 ), .A2(
        _f_permutation__n6600 ), .ZN(_f_permutation__n4006 ) );
  NAND2_X2 _f_permutation__U5300  ( .A1(_f_permutation__round_out[1380]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6597 ) );
  NAND2_X2 _f_permutation__U5299  ( .A1(_f_permutation__n7188 ), .A2(out[284]), 
        .ZN(_f_permutation__n6598 ) );
  NAND2_X2 _f_permutation__U5298  ( .A1(_f_permutation__n6597 ), .A2(
        _f_permutation__n6598 ), .ZN(_f_permutation__n4007 ) );
  NAND2_X2 _f_permutation__U5297  ( .A1(_f_permutation__round_out[1379]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6595 ) );
  NAND2_X2 _f_permutation__U5296  ( .A1(_f_permutation__n7189 ), .A2(out[283]), 
        .ZN(_f_permutation__n6596 ) );
  NAND2_X2 _f_permutation__U5295  ( .A1(_f_permutation__n6595 ), .A2(
        _f_permutation__n6596 ), .ZN(_f_permutation__n4008 ) );
  NAND2_X2 _f_permutation__U5294  ( .A1(_f_permutation__round_out[1378]), 
        .A2(_f_permutation__n7099 ), .ZN(_f_permutation__n6593 ) );
  NAND2_X2 _f_permutation__U5293  ( .A1(_f_permutation__n7189 ), .A2(out[282]), 
        .ZN(_f_permutation__n6594 ) );
  NAND2_X2 _f_permutation__U5292  ( .A1(_f_permutation__n6593 ), .A2(
        _f_permutation__n6594 ), .ZN(_f_permutation__n4009 ) );
  NAND2_X2 _f_permutation__U5291  ( .A1(_f_permutation__round_out[1377]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6591 ) );
  NAND2_X2 _f_permutation__U5290  ( .A1(_f_permutation__n7189 ), .A2(out[281]), 
        .ZN(_f_permutation__n6592 ) );
  NAND2_X2 _f_permutation__U5289  ( .A1(_f_permutation__n6591 ), .A2(
        _f_permutation__n6592 ), .ZN(_f_permutation__n4010 ) );
  NAND2_X2 _f_permutation__U5288  ( .A1(_f_permutation__round_out[1376]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6589 ) );
  NAND2_X2 _f_permutation__U5287  ( .A1(_f_permutation__n7189 ), .A2(out[280]), 
        .ZN(_f_permutation__n6590 ) );
  NAND2_X2 _f_permutation__U5286  ( .A1(_f_permutation__n6589 ), .A2(
        _f_permutation__n6590 ), .ZN(_f_permutation__n4011 ) );
  NAND2_X2 _f_permutation__U5285  ( .A1(_f_permutation__round_out[1375]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6587 ) );
  NAND2_X2 _f_permutation__U5284  ( .A1(_f_permutation__n7189 ), .A2(out[295]), 
        .ZN(_f_permutation__n6588 ) );
  NAND2_X2 _f_permutation__U5283  ( .A1(_f_permutation__n6587 ), .A2(
        _f_permutation__n6588 ), .ZN(_f_permutation__n4012 ) );
  NAND2_X2 _f_permutation__U5282  ( .A1(_f_permutation__round_out[1374]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6585 ) );
  NAND2_X2 _f_permutation__U5281  ( .A1(_f_permutation__n7189 ), .A2(out[294]), 
        .ZN(_f_permutation__n6586 ) );
  NAND2_X2 _f_permutation__U5280  ( .A1(_f_permutation__n6585 ), .A2(
        _f_permutation__n6586 ), .ZN(_f_permutation__n4013 ) );
  NAND2_X2 _f_permutation__U5279  ( .A1(_f_permutation__round_out[1373]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6583 ) );
  NAND2_X2 _f_permutation__U5278  ( .A1(_f_permutation__n7189 ), .A2(out[293]), 
        .ZN(_f_permutation__n6584 ) );
  NAND2_X2 _f_permutation__U5277  ( .A1(_f_permutation__n6583 ), .A2(
        _f_permutation__n6584 ), .ZN(_f_permutation__n4014 ) );
  NAND2_X2 _f_permutation__U5276  ( .A1(_f_permutation__round_out[1372]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6581 ) );
  NAND2_X2 _f_permutation__U5275  ( .A1(_f_permutation__n7189 ), .A2(out[292]), 
        .ZN(_f_permutation__n6582 ) );
  NAND2_X2 _f_permutation__U5274  ( .A1(_f_permutation__n6581 ), .A2(
        _f_permutation__n6582 ), .ZN(_f_permutation__n4015 ) );
  NAND2_X2 _f_permutation__U5273  ( .A1(_f_permutation__round_out[1371]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6579 ) );
  NAND2_X2 _f_permutation__U5272  ( .A1(_f_permutation__n7189 ), .A2(out[291]), 
        .ZN(_f_permutation__n6580 ) );
  NAND2_X2 _f_permutation__U5271  ( .A1(_f_permutation__n6579 ), .A2(
        _f_permutation__n6580 ), .ZN(_f_permutation__n4016 ) );
  NAND2_X2 _f_permutation__U5270  ( .A1(_f_permutation__round_out[1370]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6577 ) );
  NAND2_X2 _f_permutation__U5269  ( .A1(_f_permutation__n7189 ), .A2(out[290]), 
        .ZN(_f_permutation__n6578 ) );
  NAND2_X2 _f_permutation__U5268  ( .A1(_f_permutation__n6577 ), .A2(
        _f_permutation__n6578 ), .ZN(_f_permutation__n4017 ) );
  NAND2_X2 _f_permutation__U5267  ( .A1(_f_permutation__round_out[1369]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6575 ) );
  NAND2_X2 _f_permutation__U5266  ( .A1(_f_permutation__n7189 ), .A2(out[289]), 
        .ZN(_f_permutation__n6576 ) );
  NAND2_X2 _f_permutation__U5265  ( .A1(_f_permutation__n6575 ), .A2(
        _f_permutation__n6576 ), .ZN(_f_permutation__n4018 ) );
  NAND2_X2 _f_permutation__U5264  ( .A1(_f_permutation__round_out[1368]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6573 ) );
  NAND2_X2 _f_permutation__U5263  ( .A1(_f_permutation__n7190 ), .A2(out[288]), 
        .ZN(_f_permutation__n6574 ) );
  NAND2_X2 _f_permutation__U5262  ( .A1(_f_permutation__n6573 ), .A2(
        _f_permutation__n6574 ), .ZN(_f_permutation__n4019 ) );
  NAND2_X2 _f_permutation__U5261  ( .A1(_f_permutation__round_out[1367]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6571 ) );
  NAND2_X2 _f_permutation__U5260  ( .A1(_f_permutation__n7190 ), .A2(out[303]), 
        .ZN(_f_permutation__n6572 ) );
  NAND2_X2 _f_permutation__U5259  ( .A1(_f_permutation__n6571 ), .A2(
        _f_permutation__n6572 ), .ZN(_f_permutation__n4020 ) );
  NAND2_X2 _f_permutation__U5258  ( .A1(_f_permutation__round_out[1366]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6569 ) );
  NAND2_X2 _f_permutation__U5257  ( .A1(_f_permutation__n7190 ), .A2(out[302]), 
        .ZN(_f_permutation__n6570 ) );
  NAND2_X2 _f_permutation__U5256  ( .A1(_f_permutation__n6569 ), .A2(
        _f_permutation__n6570 ), .ZN(_f_permutation__n4021 ) );
  NAND2_X2 _f_permutation__U5255  ( .A1(_f_permutation__round_out[1365]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6567 ) );
  NAND2_X2 _f_permutation__U5254  ( .A1(_f_permutation__n7190 ), .A2(out[301]), 
        .ZN(_f_permutation__n6568 ) );
  NAND2_X2 _f_permutation__U5253  ( .A1(_f_permutation__n6567 ), .A2(
        _f_permutation__n6568 ), .ZN(_f_permutation__n4022 ) );
  NAND2_X2 _f_permutation__U5252  ( .A1(_f_permutation__round_out[1364]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6565 ) );
  NAND2_X2 _f_permutation__U5251  ( .A1(_f_permutation__n7190 ), .A2(out[300]), 
        .ZN(_f_permutation__n6566 ) );
  NAND2_X2 _f_permutation__U5250  ( .A1(_f_permutation__n6565 ), .A2(
        _f_permutation__n6566 ), .ZN(_f_permutation__n4023 ) );
  NAND2_X2 _f_permutation__U5249  ( .A1(_f_permutation__round_out[1363]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6563 ) );
  NAND2_X2 _f_permutation__U5248  ( .A1(_f_permutation__n7190 ), .A2(out[299]), 
        .ZN(_f_permutation__n6564 ) );
  NAND2_X2 _f_permutation__U5247  ( .A1(_f_permutation__n6563 ), .A2(
        _f_permutation__n6564 ), .ZN(_f_permutation__n4024 ) );
  NAND2_X2 _f_permutation__U5246  ( .A1(_f_permutation__round_out[1362]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6561 ) );
  NAND2_X2 _f_permutation__U5245  ( .A1(_f_permutation__n7190 ), .A2(out[298]), 
        .ZN(_f_permutation__n6562 ) );
  NAND2_X2 _f_permutation__U5244  ( .A1(_f_permutation__n6561 ), .A2(
        _f_permutation__n6562 ), .ZN(_f_permutation__n4025 ) );
  NAND2_X2 _f_permutation__U5243  ( .A1(_f_permutation__round_out[1361]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6559 ) );
  NAND2_X2 _f_permutation__U5242  ( .A1(_f_permutation__n7190 ), .A2(out[297]), 
        .ZN(_f_permutation__n6560 ) );
  NAND2_X2 _f_permutation__U5241  ( .A1(_f_permutation__n6559 ), .A2(
        _f_permutation__n6560 ), .ZN(_f_permutation__n4026 ) );
  NAND2_X2 _f_permutation__U5240  ( .A1(_f_permutation__round_out[1360]), 
        .A2(_f_permutation__n7098 ), .ZN(_f_permutation__n6557 ) );
  NAND2_X2 _f_permutation__U5239  ( .A1(_f_permutation__n7190 ), .A2(out[296]), 
        .ZN(_f_permutation__n6558 ) );
  NAND2_X2 _f_permutation__U5238  ( .A1(_f_permutation__n6557 ), .A2(
        _f_permutation__n6558 ), .ZN(_f_permutation__n4027 ) );
  NAND2_X2 _f_permutation__U5237  ( .A1(_f_permutation__round_out[1359]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6555 ) );
  NAND2_X2 _f_permutation__U5236  ( .A1(_f_permutation__n7190 ), .A2(out[311]), 
        .ZN(_f_permutation__n6556 ) );
  NAND2_X2 _f_permutation__U5235  ( .A1(_f_permutation__n6555 ), .A2(
        _f_permutation__n6556 ), .ZN(_f_permutation__n4028 ) );
  NAND2_X2 _f_permutation__U5234  ( .A1(_f_permutation__round_out[1358]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6553 ) );
  NAND2_X2 _f_permutation__U5233  ( .A1(_f_permutation__n7190 ), .A2(out[310]), 
        .ZN(_f_permutation__n6554 ) );
  NAND2_X2 _f_permutation__U5232  ( .A1(_f_permutation__n6553 ), .A2(
        _f_permutation__n6554 ), .ZN(_f_permutation__n4029 ) );
  NAND2_X2 _f_permutation__U5231  ( .A1(_f_permutation__round_out[1357]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6551 ) );
  NAND2_X2 _f_permutation__U5230  ( .A1(_f_permutation__n7191 ), .A2(out[309]), 
        .ZN(_f_permutation__n6552 ) );
  NAND2_X2 _f_permutation__U5229  ( .A1(_f_permutation__n6551 ), .A2(
        _f_permutation__n6552 ), .ZN(_f_permutation__n4030 ) );
  NAND2_X2 _f_permutation__U5228  ( .A1(_f_permutation__round_out[1356]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6549 ) );
  NAND2_X2 _f_permutation__U5227  ( .A1(_f_permutation__n7191 ), .A2(out[308]), 
        .ZN(_f_permutation__n6550 ) );
  NAND2_X2 _f_permutation__U5226  ( .A1(_f_permutation__n6549 ), .A2(
        _f_permutation__n6550 ), .ZN(_f_permutation__n4031 ) );
  NAND2_X2 _f_permutation__U5225  ( .A1(_f_permutation__round_out[1355]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6547 ) );
  NAND2_X2 _f_permutation__U5224  ( .A1(_f_permutation__n7191 ), .A2(out[307]), 
        .ZN(_f_permutation__n6548 ) );
  NAND2_X2 _f_permutation__U5223  ( .A1(_f_permutation__n6547 ), .A2(
        _f_permutation__n6548 ), .ZN(_f_permutation__n4032 ) );
  NAND2_X2 _f_permutation__U5222  ( .A1(_f_permutation__round_out[1354]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6545 ) );
  NAND2_X2 _f_permutation__U5221  ( .A1(_f_permutation__n7191 ), .A2(out[306]), 
        .ZN(_f_permutation__n6546 ) );
  NAND2_X2 _f_permutation__U5220  ( .A1(_f_permutation__n6545 ), .A2(
        _f_permutation__n6546 ), .ZN(_f_permutation__n4033 ) );
  NAND2_X2 _f_permutation__U5219  ( .A1(_f_permutation__round_out[1353]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6543 ) );
  NAND2_X2 _f_permutation__U5218  ( .A1(_f_permutation__n7191 ), .A2(out[305]), 
        .ZN(_f_permutation__n6544 ) );
  NAND2_X2 _f_permutation__U5217  ( .A1(_f_permutation__n6543 ), .A2(
        _f_permutation__n6544 ), .ZN(_f_permutation__n4034 ) );
  NAND2_X2 _f_permutation__U5216  ( .A1(_f_permutation__round_out[1352]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6541 ) );
  NAND2_X2 _f_permutation__U5215  ( .A1(_f_permutation__n7191 ), .A2(out[304]), 
        .ZN(_f_permutation__n6542 ) );
  NAND2_X2 _f_permutation__U5214  ( .A1(_f_permutation__n6541 ), .A2(
        _f_permutation__n6542 ), .ZN(_f_permutation__n4035 ) );
  NAND2_X2 _f_permutation__U5213  ( .A1(_f_permutation__round_out[1351]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6539 ) );
  NAND2_X2 _f_permutation__U5212  ( .A1(_f_permutation__n7191 ), .A2(out[319]), 
        .ZN(_f_permutation__n6540 ) );
  NAND2_X2 _f_permutation__U5211  ( .A1(_f_permutation__n6539 ), .A2(
        _f_permutation__n6540 ), .ZN(_f_permutation__n4036 ) );
  NAND2_X2 _f_permutation__U5210  ( .A1(_f_permutation__round_out[1350]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6537 ) );
  NAND2_X2 _f_permutation__U5209  ( .A1(_f_permutation__n7191 ), .A2(out[318]), 
        .ZN(_f_permutation__n6538 ) );
  NAND2_X2 _f_permutation__U5208  ( .A1(_f_permutation__n6537 ), .A2(
        _f_permutation__n6538 ), .ZN(_f_permutation__n4037 ) );
  NAND2_X2 _f_permutation__U5207  ( .A1(_f_permutation__round_out[1349]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6535 ) );
  NAND2_X2 _f_permutation__U5206  ( .A1(_f_permutation__n7191 ), .A2(out[317]), 
        .ZN(_f_permutation__n6536 ) );
  NAND2_X2 _f_permutation__U5205  ( .A1(_f_permutation__n6535 ), .A2(
        _f_permutation__n6536 ), .ZN(_f_permutation__n4038 ) );
  NAND2_X2 _f_permutation__U5204  ( .A1(_f_permutation__round_out[1348]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6533 ) );
  NAND2_X2 _f_permutation__U5203  ( .A1(_f_permutation__n7191 ), .A2(out[316]), 
        .ZN(_f_permutation__n6534 ) );
  NAND2_X2 _f_permutation__U5202  ( .A1(_f_permutation__n6533 ), .A2(
        _f_permutation__n6534 ), .ZN(_f_permutation__n4039 ) );
  NAND2_X2 _f_permutation__U5201  ( .A1(_f_permutation__round_out[1347]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6531 ) );
  NAND2_X2 _f_permutation__U5200  ( .A1(_f_permutation__n7191 ), .A2(out[315]), 
        .ZN(_f_permutation__n6532 ) );
  NAND2_X2 _f_permutation__U5199  ( .A1(_f_permutation__n6531 ), .A2(
        _f_permutation__n6532 ), .ZN(_f_permutation__n4040 ) );
  NAND2_X2 _f_permutation__U5198  ( .A1(_f_permutation__round_out[1346]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6529 ) );
  NAND2_X2 _f_permutation__U5197  ( .A1(_f_permutation__n7192 ), .A2(out[314]), 
        .ZN(_f_permutation__n6530 ) );
  NAND2_X2 _f_permutation__U5196  ( .A1(_f_permutation__n6529 ), .A2(
        _f_permutation__n6530 ), .ZN(_f_permutation__n4041 ) );
  NAND2_X2 _f_permutation__U5195  ( .A1(_f_permutation__round_out[1345]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6527 ) );
  NAND2_X2 _f_permutation__U5194  ( .A1(_f_permutation__n7192 ), .A2(out[313]), 
        .ZN(_f_permutation__n6528 ) );
  NAND2_X2 _f_permutation__U5193  ( .A1(_f_permutation__n6527 ), .A2(
        _f_permutation__n6528 ), .ZN(_f_permutation__n4042 ) );
  NAND2_X2 _f_permutation__U5192  ( .A1(_f_permutation__round_out[1344]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6525 ) );
  NAND2_X2 _f_permutation__U5191  ( .A1(_f_permutation__n7192 ), .A2(out[312]), 
        .ZN(_f_permutation__n6526 ) );
  NAND2_X2 _f_permutation__U5190  ( .A1(_f_permutation__n6525 ), .A2(
        _f_permutation__n6526 ), .ZN(_f_permutation__n4043 ) );
  NAND2_X2 _f_permutation__U5189  ( .A1(_f_permutation__round_out[1343]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6523 ) );
  NAND2_X2 _f_permutation__U5188  ( .A1(_f_permutation__n7192 ), .A2(out[199]), 
        .ZN(_f_permutation__n6524 ) );
  NAND2_X2 _f_permutation__U5187  ( .A1(_f_permutation__n6523 ), .A2(
        _f_permutation__n6524 ), .ZN(_f_permutation__n4044 ) );
  NAND2_X2 _f_permutation__U5186  ( .A1(_f_permutation__round_out[1342]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6521 ) );
  NAND2_X2 _f_permutation__U5185  ( .A1(_f_permutation__n7192 ), .A2(out[198]), 
        .ZN(_f_permutation__n6522 ) );
  NAND2_X2 _f_permutation__U5184  ( .A1(_f_permutation__n6521 ), .A2(
        _f_permutation__n6522 ), .ZN(_f_permutation__n4045 ) );
  NAND2_X2 _f_permutation__U5183  ( .A1(_f_permutation__round_out[1341]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6519 ) );
  NAND2_X2 _f_permutation__U5182  ( .A1(_f_permutation__n7192 ), .A2(out[197]), 
        .ZN(_f_permutation__n6520 ) );
  NAND2_X2 _f_permutation__U5181  ( .A1(_f_permutation__n6519 ), .A2(
        _f_permutation__n6520 ), .ZN(_f_permutation__n4046 ) );
  NAND2_X2 _f_permutation__U5180  ( .A1(_f_permutation__round_out[1340]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6517 ) );
  NAND2_X2 _f_permutation__U5179  ( .A1(_f_permutation__n7192 ), .A2(out[196]), 
        .ZN(_f_permutation__n6518 ) );
  NAND2_X2 _f_permutation__U5178  ( .A1(_f_permutation__n6517 ), .A2(
        _f_permutation__n6518 ), .ZN(_f_permutation__n4047 ) );
  NAND2_X2 _f_permutation__U5177  ( .A1(_f_permutation__round_out[1339]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6515 ) );
  NAND2_X2 _f_permutation__U5176  ( .A1(_f_permutation__n7192 ), .A2(out[195]), 
        .ZN(_f_permutation__n6516 ) );
  NAND2_X2 _f_permutation__U5175  ( .A1(_f_permutation__n6515 ), .A2(
        _f_permutation__n6516 ), .ZN(_f_permutation__n4048 ) );
  NAND2_X2 _f_permutation__U5174  ( .A1(_f_permutation__round_out[1338]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6513 ) );
  NAND2_X2 _f_permutation__U5173  ( .A1(_f_permutation__n7192 ), .A2(out[194]), 
        .ZN(_f_permutation__n6514 ) );
  NAND2_X2 _f_permutation__U5172  ( .A1(_f_permutation__n6513 ), .A2(
        _f_permutation__n6514 ), .ZN(_f_permutation__n4049 ) );
  NAND2_X2 _f_permutation__U5171  ( .A1(_f_permutation__round_out[1337]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6511 ) );
  NAND2_X2 _f_permutation__U5170  ( .A1(_f_permutation__n7192 ), .A2(out[193]), 
        .ZN(_f_permutation__n6512 ) );
  NAND2_X2 _f_permutation__U5169  ( .A1(_f_permutation__n6511 ), .A2(
        _f_permutation__n6512 ), .ZN(_f_permutation__n4050 ) );
  NAND2_X2 _f_permutation__U5168  ( .A1(_f_permutation__round_out[1336]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6509 ) );
  NAND2_X2 _f_permutation__U5167  ( .A1(_f_permutation__n7192 ), .A2(out[192]), 
        .ZN(_f_permutation__n6510 ) );
  NAND2_X2 _f_permutation__U5166  ( .A1(_f_permutation__n6509 ), .A2(
        _f_permutation__n6510 ), .ZN(_f_permutation__n4051 ) );
  NAND2_X2 _f_permutation__U5165  ( .A1(_f_permutation__round_out[1335]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6507 ) );
  NAND2_X2 _f_permutation__U5164  ( .A1(_f_permutation__n7193 ), .A2(out[207]), 
        .ZN(_f_permutation__n6508 ) );
  NAND2_X2 _f_permutation__U5163  ( .A1(_f_permutation__n6507 ), .A2(
        _f_permutation__n6508 ), .ZN(_f_permutation__n4052 ) );
  NAND2_X2 _f_permutation__U5162  ( .A1(_f_permutation__round_out[1334]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6505 ) );
  NAND2_X2 _f_permutation__U5161  ( .A1(_f_permutation__n7193 ), .A2(out[206]), 
        .ZN(_f_permutation__n6506 ) );
  NAND2_X2 _f_permutation__U5160  ( .A1(_f_permutation__n6505 ), .A2(
        _f_permutation__n6506 ), .ZN(_f_permutation__n4053 ) );
  NAND2_X2 _f_permutation__U5159  ( .A1(_f_permutation__round_out[1333]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6503 ) );
  NAND2_X2 _f_permutation__U5158  ( .A1(_f_permutation__n7193 ), .A2(out[205]), 
        .ZN(_f_permutation__n6504 ) );
  NAND2_X2 _f_permutation__U5157  ( .A1(_f_permutation__n6503 ), .A2(
        _f_permutation__n6504 ), .ZN(_f_permutation__n4054 ) );
  NAND2_X2 _f_permutation__U5156  ( .A1(_f_permutation__round_out[1332]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6501 ) );
  NAND2_X2 _f_permutation__U5155  ( .A1(_f_permutation__n7193 ), .A2(out[204]), 
        .ZN(_f_permutation__n6502 ) );
  NAND2_X2 _f_permutation__U5154  ( .A1(_f_permutation__n6501 ), .A2(
        _f_permutation__n6502 ), .ZN(_f_permutation__n4055 ) );
  NAND2_X2 _f_permutation__U5153  ( .A1(_f_permutation__round_out[1331]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6499 ) );
  NAND2_X2 _f_permutation__U5152  ( .A1(_f_permutation__n7193 ), .A2(out[203]), 
        .ZN(_f_permutation__n6500 ) );
  NAND2_X2 _f_permutation__U5151  ( .A1(_f_permutation__n6499 ), .A2(
        _f_permutation__n6500 ), .ZN(_f_permutation__n4056 ) );
  NAND2_X2 _f_permutation__U5150  ( .A1(_f_permutation__round_out[1330]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6497 ) );
  NAND2_X2 _f_permutation__U5149  ( .A1(_f_permutation__n7193 ), .A2(out[202]), 
        .ZN(_f_permutation__n6498 ) );
  NAND2_X2 _f_permutation__U5148  ( .A1(_f_permutation__n6497 ), .A2(
        _f_permutation__n6498 ), .ZN(_f_permutation__n4057 ) );
  NAND2_X2 _f_permutation__U5147  ( .A1(_f_permutation__round_out[1329]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6495 ) );
  NAND2_X2 _f_permutation__U5146  ( .A1(_f_permutation__n7193 ), .A2(out[201]), 
        .ZN(_f_permutation__n6496 ) );
  NAND2_X2 _f_permutation__U5145  ( .A1(_f_permutation__n6495 ), .A2(
        _f_permutation__n6496 ), .ZN(_f_permutation__n4058 ) );
  NAND2_X2 _f_permutation__U5144  ( .A1(_f_permutation__round_out[1328]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6493 ) );
  NAND2_X2 _f_permutation__U5143  ( .A1(_f_permutation__n7193 ), .A2(out[200]), 
        .ZN(_f_permutation__n6494 ) );
  NAND2_X2 _f_permutation__U5142  ( .A1(_f_permutation__n6493 ), .A2(
        _f_permutation__n6494 ), .ZN(_f_permutation__n4059 ) );
  NAND2_X2 _f_permutation__U5141  ( .A1(_f_permutation__round_out[1327]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6491 ) );
  NAND2_X2 _f_permutation__U5140  ( .A1(_f_permutation__n7193 ), .A2(out[215]), 
        .ZN(_f_permutation__n6492 ) );
  NAND2_X2 _f_permutation__U5139  ( .A1(_f_permutation__n6491 ), .A2(
        _f_permutation__n6492 ), .ZN(_f_permutation__n4060 ) );
  NAND2_X2 _f_permutation__U5138  ( .A1(_f_permutation__round_out[1326]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6489 ) );
  NAND2_X2 _f_permutation__U5137  ( .A1(_f_permutation__n7193 ), .A2(out[214]), 
        .ZN(_f_permutation__n6490 ) );
  NAND2_X2 _f_permutation__U5136  ( .A1(_f_permutation__n6489 ), .A2(
        _f_permutation__n6490 ), .ZN(_f_permutation__n4061 ) );
  NAND2_X2 _f_permutation__U5135  ( .A1(_f_permutation__round_out[1325]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6487 ) );
  NAND2_X2 _f_permutation__U5134  ( .A1(_f_permutation__n7193 ), .A2(out[213]), 
        .ZN(_f_permutation__n6488 ) );
  NAND2_X2 _f_permutation__U5133  ( .A1(_f_permutation__n6487 ), .A2(
        _f_permutation__n6488 ), .ZN(_f_permutation__n4062 ) );
  NAND2_X2 _f_permutation__U5132  ( .A1(_f_permutation__round_out[1324]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6485 ) );
  NAND2_X2 _f_permutation__U5131  ( .A1(_f_permutation__n7194 ), .A2(out[212]), 
        .ZN(_f_permutation__n6486 ) );
  NAND2_X2 _f_permutation__U5130  ( .A1(_f_permutation__n6485 ), .A2(
        _f_permutation__n6486 ), .ZN(_f_permutation__n4063 ) );
  NAND2_X2 _f_permutation__U5129  ( .A1(_f_permutation__round_out[1323]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6483 ) );
  NAND2_X2 _f_permutation__U5128  ( .A1(_f_permutation__n7194 ), .A2(out[211]), 
        .ZN(_f_permutation__n6484 ) );
  NAND2_X2 _f_permutation__U5127  ( .A1(_f_permutation__n6483 ), .A2(
        _f_permutation__n6484 ), .ZN(_f_permutation__n4064 ) );
  NAND2_X2 _f_permutation__U5126  ( .A1(_f_permutation__round_out[1322]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6481 ) );
  NAND2_X2 _f_permutation__U5125  ( .A1(_f_permutation__n7194 ), .A2(out[210]), 
        .ZN(_f_permutation__n6482 ) );
  NAND2_X2 _f_permutation__U5124  ( .A1(_f_permutation__n6481 ), .A2(
        _f_permutation__n6482 ), .ZN(_f_permutation__n4065 ) );
  NAND2_X2 _f_permutation__U5123  ( .A1(_f_permutation__round_out[1321]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6479 ) );
  NAND2_X2 _f_permutation__U5122  ( .A1(_f_permutation__n7194 ), .A2(out[209]), 
        .ZN(_f_permutation__n6480 ) );
  NAND2_X2 _f_permutation__U5121  ( .A1(_f_permutation__n6479 ), .A2(
        _f_permutation__n6480 ), .ZN(_f_permutation__n4066 ) );
  NAND2_X2 _f_permutation__U5120  ( .A1(_f_permutation__round_out[1320]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6477 ) );
  NAND2_X2 _f_permutation__U5119  ( .A1(_f_permutation__n7194 ), .A2(out[208]), 
        .ZN(_f_permutation__n6478 ) );
  NAND2_X2 _f_permutation__U5118  ( .A1(_f_permutation__n6477 ), .A2(
        _f_permutation__n6478 ), .ZN(_f_permutation__n4067 ) );
  NAND2_X2 _f_permutation__U5117  ( .A1(_f_permutation__round_out[1319]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6475 ) );
  NAND2_X2 _f_permutation__U5116  ( .A1(_f_permutation__n7194 ), .A2(out[223]), 
        .ZN(_f_permutation__n6476 ) );
  NAND2_X2 _f_permutation__U5115  ( .A1(_f_permutation__n6475 ), .A2(
        _f_permutation__n6476 ), .ZN(_f_permutation__n4068 ) );
  NAND2_X2 _f_permutation__U5114  ( .A1(_f_permutation__round_out[1318]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6473 ) );
  NAND2_X2 _f_permutation__U5113  ( .A1(_f_permutation__n7194 ), .A2(out[222]), 
        .ZN(_f_permutation__n6474 ) );
  NAND2_X2 _f_permutation__U5112  ( .A1(_f_permutation__n6473 ), .A2(
        _f_permutation__n6474 ), .ZN(_f_permutation__n4069 ) );
  NAND2_X2 _f_permutation__U5111  ( .A1(_f_permutation__round_out[1317]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6471 ) );
  NAND2_X2 _f_permutation__U5110  ( .A1(_f_permutation__n7194 ), .A2(out[221]), 
        .ZN(_f_permutation__n6472 ) );
  NAND2_X2 _f_permutation__U5109  ( .A1(_f_permutation__n6471 ), .A2(
        _f_permutation__n6472 ), .ZN(_f_permutation__n4070 ) );
  NAND2_X2 _f_permutation__U5108  ( .A1(_f_permutation__round_out[1316]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6469 ) );
  NAND2_X2 _f_permutation__U5107  ( .A1(_f_permutation__n7194 ), .A2(out[220]), 
        .ZN(_f_permutation__n6470 ) );
  NAND2_X2 _f_permutation__U5106  ( .A1(_f_permutation__n6469 ), .A2(
        _f_permutation__n6470 ), .ZN(_f_permutation__n4071 ) );
  NAND2_X2 _f_permutation__U5105  ( .A1(_f_permutation__round_out[1315]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6467 ) );
  NAND2_X2 _f_permutation__U5104  ( .A1(_f_permutation__n7194 ), .A2(out[219]), 
        .ZN(_f_permutation__n6468 ) );
  NAND2_X2 _f_permutation__U5103  ( .A1(_f_permutation__n6467 ), .A2(
        _f_permutation__n6468 ), .ZN(_f_permutation__n4072 ) );
  NAND2_X2 _f_permutation__U5102  ( .A1(_f_permutation__round_out[1314]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6465 ) );
  NAND2_X2 _f_permutation__U5101  ( .A1(_f_permutation__n7194 ), .A2(out[218]), 
        .ZN(_f_permutation__n6466 ) );
  NAND2_X2 _f_permutation__U5100  ( .A1(_f_permutation__n6465 ), .A2(
        _f_permutation__n6466 ), .ZN(_f_permutation__n4073 ) );
  NAND2_X2 _f_permutation__U5099  ( .A1(_f_permutation__round_out[1313]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6463 ) );
  NAND2_X2 _f_permutation__U5098  ( .A1(_f_permutation__n7195 ), .A2(out[217]), 
        .ZN(_f_permutation__n6464 ) );
  NAND2_X2 _f_permutation__U5097  ( .A1(_f_permutation__n6463 ), .A2(
        _f_permutation__n6464 ), .ZN(_f_permutation__n4074 ) );
  NAND2_X2 _f_permutation__U5096  ( .A1(_f_permutation__round_out[1312]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6461 ) );
  NAND2_X2 _f_permutation__U5095  ( .A1(_f_permutation__n7195 ), .A2(out[216]), 
        .ZN(_f_permutation__n6462 ) );
  NAND2_X2 _f_permutation__U5094  ( .A1(_f_permutation__n6461 ), .A2(
        _f_permutation__n6462 ), .ZN(_f_permutation__n4075 ) );
  NAND2_X2 _f_permutation__U5093  ( .A1(_f_permutation__round_out[1311]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6459 ) );
  NAND2_X2 _f_permutation__U5092  ( .A1(_f_permutation__n7195 ), .A2(out[231]), 
        .ZN(_f_permutation__n6460 ) );
  NAND2_X2 _f_permutation__U5091  ( .A1(_f_permutation__n6459 ), .A2(
        _f_permutation__n6460 ), .ZN(_f_permutation__n4076 ) );
  NAND2_X2 _f_permutation__U5090  ( .A1(_f_permutation__round_out[1310]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6457 ) );
  NAND2_X2 _f_permutation__U5089  ( .A1(_f_permutation__n7195 ), .A2(out[230]), 
        .ZN(_f_permutation__n6458 ) );
  NAND2_X2 _f_permutation__U5088  ( .A1(_f_permutation__n6457 ), .A2(
        _f_permutation__n6458 ), .ZN(_f_permutation__n4077 ) );
  NAND2_X2 _f_permutation__U5087  ( .A1(_f_permutation__round_out[1309]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6455 ) );
  NAND2_X2 _f_permutation__U5086  ( .A1(_f_permutation__n7195 ), .A2(out[229]), 
        .ZN(_f_permutation__n6456 ) );
  NAND2_X2 _f_permutation__U5085  ( .A1(_f_permutation__n6455 ), .A2(
        _f_permutation__n6456 ), .ZN(_f_permutation__n4078 ) );
  NAND2_X2 _f_permutation__U5084  ( .A1(_f_permutation__round_out[1308]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6453 ) );
  NAND2_X2 _f_permutation__U5083  ( .A1(_f_permutation__n7195 ), .A2(out[228]), 
        .ZN(_f_permutation__n6454 ) );
  NAND2_X2 _f_permutation__U5082  ( .A1(_f_permutation__n6453 ), .A2(
        _f_permutation__n6454 ), .ZN(_f_permutation__n4079 ) );
  NAND2_X2 _f_permutation__U5081  ( .A1(_f_permutation__round_out[1307]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6451 ) );
  NAND2_X2 _f_permutation__U5080  ( .A1(_f_permutation__n7195 ), .A2(out[227]), 
        .ZN(_f_permutation__n6452 ) );
  NAND2_X2 _f_permutation__U5079  ( .A1(_f_permutation__n6451 ), .A2(
        _f_permutation__n6452 ), .ZN(_f_permutation__n4080 ) );
  NAND2_X2 _f_permutation__U5078  ( .A1(_f_permutation__round_out[1306]), 
        .A2(_f_permutation__n7096 ), .ZN(_f_permutation__n6449 ) );
  NAND2_X2 _f_permutation__U5077  ( .A1(_f_permutation__n7195 ), .A2(out[226]), 
        .ZN(_f_permutation__n6450 ) );
  NAND2_X2 _f_permutation__U5076  ( .A1(_f_permutation__n6449 ), .A2(
        _f_permutation__n6450 ), .ZN(_f_permutation__n4081 ) );
  NAND2_X2 _f_permutation__U5075  ( .A1(_f_permutation__round_out[1305]), 
        .A2(_f_permutation__n7095 ), .ZN(_f_permutation__n6447 ) );
  NAND2_X2 _f_permutation__U5074  ( .A1(_f_permutation__n7195 ), .A2(out[225]), 
        .ZN(_f_permutation__n6448 ) );
  NAND2_X2 _f_permutation__U5073  ( .A1(_f_permutation__n6447 ), .A2(
        _f_permutation__n6448 ), .ZN(_f_permutation__n4082 ) );
  NAND2_X2 _f_permutation__U5072  ( .A1(_f_permutation__round_out[1304]), 
        .A2(_f_permutation__n7153 ), .ZN(_f_permutation__n6445 ) );
  NAND2_X2 _f_permutation__U5071  ( .A1(_f_permutation__n7195 ), .A2(out[224]), 
        .ZN(_f_permutation__n6446 ) );
  NAND2_X2 _f_permutation__U5070  ( .A1(_f_permutation__n6445 ), .A2(
        _f_permutation__n6446 ), .ZN(_f_permutation__n4083 ) );
  NAND2_X2 _f_permutation__U5069  ( .A1(_f_permutation__round_out[1303]), 
        .A2(_f_permutation__n7163 ), .ZN(_f_permutation__n6443 ) );
  NAND2_X2 _f_permutation__U5068  ( .A1(_f_permutation__n7195 ), .A2(out[239]), 
        .ZN(_f_permutation__n6444 ) );
  NAND2_X2 _f_permutation__U5067  ( .A1(_f_permutation__n6443 ), .A2(
        _f_permutation__n6444 ), .ZN(_f_permutation__n4084 ) );
  NAND2_X2 _f_permutation__U5066  ( .A1(_f_permutation__round_out[1302]), 
        .A2(_f_permutation__n7162 ), .ZN(_f_permutation__n6441 ) );
  NAND2_X2 _f_permutation__U5065  ( .A1(_f_permutation__n7196 ), .A2(out[238]), 
        .ZN(_f_permutation__n6442 ) );
  NAND2_X2 _f_permutation__U5064  ( .A1(_f_permutation__n6441 ), .A2(
        _f_permutation__n6442 ), .ZN(_f_permutation__n4085 ) );
  NAND2_X2 _f_permutation__U5063  ( .A1(_f_permutation__round_out[1301]), 
        .A2(_f_permutation__n7167 ), .ZN(_f_permutation__n6439 ) );
  NAND2_X2 _f_permutation__U5062  ( .A1(_f_permutation__n7196 ), .A2(out[237]), 
        .ZN(_f_permutation__n6440 ) );
  NAND2_X2 _f_permutation__U5061  ( .A1(_f_permutation__n6439 ), .A2(
        _f_permutation__n6440 ), .ZN(_f_permutation__n4086 ) );
  NAND2_X2 _f_permutation__U5060  ( .A1(_f_permutation__round_out[1300]), 
        .A2(_f_permutation__n7166 ), .ZN(_f_permutation__n6437 ) );
  NAND2_X2 _f_permutation__U5059  ( .A1(_f_permutation__n7196 ), .A2(out[236]), 
        .ZN(_f_permutation__n6438 ) );
  NAND2_X2 _f_permutation__U5058  ( .A1(_f_permutation__n6437 ), .A2(
        _f_permutation__n6438 ), .ZN(_f_permutation__n4087 ) );
  NAND2_X2 _f_permutation__U5057  ( .A1(_f_permutation__round_out[1299]), 
        .A2(_f_permutation__n7097 ), .ZN(_f_permutation__n6435 ) );
  NAND2_X2 _f_permutation__U5056  ( .A1(_f_permutation__n7196 ), .A2(out[235]), 
        .ZN(_f_permutation__n6436 ) );
  NAND2_X2 _f_permutation__U5055  ( .A1(_f_permutation__n6435 ), .A2(
        _f_permutation__n6436 ), .ZN(_f_permutation__n4088 ) );
  NAND2_X2 _f_permutation__U5054  ( .A1(_f_permutation__round_out[1298]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6433 ) );
  NAND2_X2 _f_permutation__U5053  ( .A1(_f_permutation__n7196 ), .A2(out[234]), 
        .ZN(_f_permutation__n6434 ) );
  NAND2_X2 _f_permutation__U5052  ( .A1(_f_permutation__n6433 ), .A2(
        _f_permutation__n6434 ), .ZN(_f_permutation__n4089 ) );
  NAND2_X2 _f_permutation__U5051  ( .A1(_f_permutation__round_out[1297]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6431 ) );
  NAND2_X2 _f_permutation__U5050  ( .A1(_f_permutation__n7196 ), .A2(out[233]), 
        .ZN(_f_permutation__n6432 ) );
  NAND2_X2 _f_permutation__U5049  ( .A1(_f_permutation__n6431 ), .A2(
        _f_permutation__n6432 ), .ZN(_f_permutation__n4090 ) );
  NAND2_X2 _f_permutation__U5048  ( .A1(_f_permutation__round_out[1296]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6429 ) );
  NAND2_X2 _f_permutation__U5047  ( .A1(_f_permutation__n7196 ), .A2(out[232]), 
        .ZN(_f_permutation__n6430 ) );
  NAND2_X2 _f_permutation__U5046  ( .A1(_f_permutation__n6429 ), .A2(
        _f_permutation__n6430 ), .ZN(_f_permutation__n4091 ) );
  NAND2_X2 _f_permutation__U5045  ( .A1(_f_permutation__round_out[1295]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6427 ) );
  NAND2_X2 _f_permutation__U5044  ( .A1(_f_permutation__n7196 ), .A2(out[247]), 
        .ZN(_f_permutation__n6428 ) );
  NAND2_X2 _f_permutation__U5043  ( .A1(_f_permutation__n6427 ), .A2(
        _f_permutation__n6428 ), .ZN(_f_permutation__n4092 ) );
  NAND2_X2 _f_permutation__U5042  ( .A1(_f_permutation__round_out[1294]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6425 ) );
  NAND2_X2 _f_permutation__U5041  ( .A1(_f_permutation__n7196 ), .A2(out[246]), 
        .ZN(_f_permutation__n6426 ) );
  NAND2_X2 _f_permutation__U5040  ( .A1(_f_permutation__n6425 ), .A2(
        _f_permutation__n6426 ), .ZN(_f_permutation__n4093 ) );
  NAND2_X2 _f_permutation__U5039  ( .A1(_f_permutation__round_out[1293]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6423 ) );
  NAND2_X2 _f_permutation__U5038  ( .A1(_f_permutation__n7196 ), .A2(out[245]), 
        .ZN(_f_permutation__n6424 ) );
  NAND2_X2 _f_permutation__U5037  ( .A1(_f_permutation__n6423 ), .A2(
        _f_permutation__n6424 ), .ZN(_f_permutation__n4094 ) );
  NAND2_X2 _f_permutation__U5036  ( .A1(_f_permutation__round_out[1292]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6421 ) );
  NAND2_X2 _f_permutation__U5035  ( .A1(_f_permutation__n7196 ), .A2(out[244]), 
        .ZN(_f_permutation__n6422 ) );
  NAND2_X2 _f_permutation__U5034  ( .A1(_f_permutation__n6421 ), .A2(
        _f_permutation__n6422 ), .ZN(_f_permutation__n4095 ) );
  NAND2_X2 _f_permutation__U5033  ( .A1(_f_permutation__round_out[1291]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6419 ) );
  NAND2_X2 _f_permutation__U5032  ( .A1(_f_permutation__n7197 ), .A2(out[243]), 
        .ZN(_f_permutation__n6420 ) );
  NAND2_X2 _f_permutation__U5031  ( .A1(_f_permutation__n6419 ), .A2(
        _f_permutation__n6420 ), .ZN(_f_permutation__n4096 ) );
  NAND2_X2 _f_permutation__U5030  ( .A1(_f_permutation__round_out[1290]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6417 ) );
  NAND2_X2 _f_permutation__U5029  ( .A1(_f_permutation__n7197 ), .A2(out[242]), 
        .ZN(_f_permutation__n6418 ) );
  NAND2_X2 _f_permutation__U5028  ( .A1(_f_permutation__n6417 ), .A2(
        _f_permutation__n6418 ), .ZN(_f_permutation__n4097 ) );
  NAND2_X2 _f_permutation__U5027  ( .A1(_f_permutation__round_out[1289]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6415 ) );
  NAND2_X2 _f_permutation__U5026  ( .A1(_f_permutation__n7197 ), .A2(out[241]), 
        .ZN(_f_permutation__n6416 ) );
  NAND2_X2 _f_permutation__U5025  ( .A1(_f_permutation__n6415 ), .A2(
        _f_permutation__n6416 ), .ZN(_f_permutation__n4098 ) );
  NAND2_X2 _f_permutation__U5024  ( .A1(_f_permutation__round_out[1288]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6413 ) );
  NAND2_X2 _f_permutation__U5023  ( .A1(_f_permutation__n7197 ), .A2(out[240]), 
        .ZN(_f_permutation__n6414 ) );
  NAND2_X2 _f_permutation__U5022  ( .A1(_f_permutation__n6413 ), .A2(
        _f_permutation__n6414 ), .ZN(_f_permutation__n4099 ) );
  NAND2_X2 _f_permutation__U5021  ( .A1(_f_permutation__round_out[1287]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6411 ) );
  NAND2_X2 _f_permutation__U5020  ( .A1(_f_permutation__n7197 ), .A2(out[255]), 
        .ZN(_f_permutation__n6412 ) );
  NAND2_X2 _f_permutation__U5019  ( .A1(_f_permutation__n6411 ), .A2(
        _f_permutation__n6412 ), .ZN(_f_permutation__n4100 ) );
  NAND2_X2 _f_permutation__U5018  ( .A1(_f_permutation__round_out[1286]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6409 ) );
  NAND2_X2 _f_permutation__U5017  ( .A1(_f_permutation__n7197 ), .A2(out[254]), 
        .ZN(_f_permutation__n6410 ) );
  NAND2_X2 _f_permutation__U5016  ( .A1(_f_permutation__n6409 ), .A2(
        _f_permutation__n6410 ), .ZN(_f_permutation__n4101 ) );
  NAND2_X2 _f_permutation__U5015  ( .A1(_f_permutation__round_out[1285]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6407 ) );
  NAND2_X2 _f_permutation__U5014  ( .A1(_f_permutation__n7197 ), .A2(out[253]), 
        .ZN(_f_permutation__n6408 ) );
  NAND2_X2 _f_permutation__U5013  ( .A1(_f_permutation__n6407 ), .A2(
        _f_permutation__n6408 ), .ZN(_f_permutation__n4102 ) );
  NAND2_X2 _f_permutation__U5012  ( .A1(_f_permutation__round_out[1284]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6405 ) );
  NAND2_X2 _f_permutation__U5011  ( .A1(_f_permutation__n7197 ), .A2(out[252]), 
        .ZN(_f_permutation__n6406 ) );
  NAND2_X2 _f_permutation__U5010  ( .A1(_f_permutation__n6405 ), .A2(
        _f_permutation__n6406 ), .ZN(_f_permutation__n4103 ) );
  NAND2_X2 _f_permutation__U5009  ( .A1(_f_permutation__round_out[1283]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6403 ) );
  NAND2_X2 _f_permutation__U5008  ( .A1(_f_permutation__n7197 ), .A2(out[251]), 
        .ZN(_f_permutation__n6404 ) );
  NAND2_X2 _f_permutation__U5007  ( .A1(_f_permutation__n6403 ), .A2(
        _f_permutation__n6404 ), .ZN(_f_permutation__n4104 ) );
  NAND2_X2 _f_permutation__U5006  ( .A1(_f_permutation__round_out[1282]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6401 ) );
  NAND2_X2 _f_permutation__U5005  ( .A1(_f_permutation__n7197 ), .A2(out[250]), 
        .ZN(_f_permutation__n6402 ) );
  NAND2_X2 _f_permutation__U5004  ( .A1(_f_permutation__n6401 ), .A2(
        _f_permutation__n6402 ), .ZN(_f_permutation__n4105 ) );
  NAND2_X2 _f_permutation__U5003  ( .A1(_f_permutation__round_out[1281]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6399 ) );
  NAND2_X2 _f_permutation__U5002  ( .A1(_f_permutation__n7197 ), .A2(out[249]), 
        .ZN(_f_permutation__n6400 ) );
  NAND2_X2 _f_permutation__U5001  ( .A1(_f_permutation__n6399 ), .A2(
        _f_permutation__n6400 ), .ZN(_f_permutation__n4106 ) );
  NAND2_X2 _f_permutation__U5000  ( .A1(_f_permutation__round_out[1280]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6397 ) );
  NAND2_X2 _f_permutation__U4999  ( .A1(_f_permutation__n7198 ), .A2(out[248]), 
        .ZN(_f_permutation__n6398 ) );
  NAND2_X2 _f_permutation__U4998  ( .A1(_f_permutation__n6397 ), .A2(
        _f_permutation__n6398 ), .ZN(_f_permutation__n4107 ) );
  NAND2_X2 _f_permutation__U4997  ( .A1(_f_permutation__round_out[1279]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6395 ) );
  NAND2_X2 _f_permutation__U4996  ( .A1(_f_permutation__n7198 ), .A2(out[135]), 
        .ZN(_f_permutation__n6396 ) );
  NAND2_X2 _f_permutation__U4995  ( .A1(_f_permutation__n6395 ), .A2(
        _f_permutation__n6396 ), .ZN(_f_permutation__n4108 ) );
  NAND2_X2 _f_permutation__U4994  ( .A1(_f_permutation__round_out[1278]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6393 ) );
  NAND2_X2 _f_permutation__U4993  ( .A1(_f_permutation__n7198 ), .A2(out[134]), 
        .ZN(_f_permutation__n6394 ) );
  NAND2_X2 _f_permutation__U4992  ( .A1(_f_permutation__n6393 ), .A2(
        _f_permutation__n6394 ), .ZN(_f_permutation__n4109 ) );
  NAND2_X2 _f_permutation__U4991  ( .A1(_f_permutation__round_out[1277]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6391 ) );
  NAND2_X2 _f_permutation__U4990  ( .A1(_f_permutation__n7198 ), .A2(out[133]), 
        .ZN(_f_permutation__n6392 ) );
  NAND2_X2 _f_permutation__U4989  ( .A1(_f_permutation__n6391 ), .A2(
        _f_permutation__n6392 ), .ZN(_f_permutation__n4110 ) );
  NAND2_X2 _f_permutation__U4988  ( .A1(_f_permutation__round_out[1276]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6389 ) );
  NAND2_X2 _f_permutation__U4987  ( .A1(_f_permutation__n7198 ), .A2(out[132]), 
        .ZN(_f_permutation__n6390 ) );
  NAND2_X2 _f_permutation__U4986  ( .A1(_f_permutation__n6389 ), .A2(
        _f_permutation__n6390 ), .ZN(_f_permutation__n4111 ) );
  NAND2_X2 _f_permutation__U4985  ( .A1(_f_permutation__round_out[1275]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6387 ) );
  NAND2_X2 _f_permutation__U4984  ( .A1(_f_permutation__n7198 ), .A2(out[131]), 
        .ZN(_f_permutation__n6388 ) );
  NAND2_X2 _f_permutation__U4983  ( .A1(_f_permutation__n6387 ), .A2(
        _f_permutation__n6388 ), .ZN(_f_permutation__n4112 ) );
  NAND2_X2 _f_permutation__U4982  ( .A1(_f_permutation__round_out[1274]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6385 ) );
  NAND2_X2 _f_permutation__U4981  ( .A1(_f_permutation__n7198 ), .A2(out[130]), 
        .ZN(_f_permutation__n6386 ) );
  NAND2_X2 _f_permutation__U4980  ( .A1(_f_permutation__n6385 ), .A2(
        _f_permutation__n6386 ), .ZN(_f_permutation__n4113 ) );
  NAND2_X2 _f_permutation__U4979  ( .A1(_f_permutation__round_out[1273]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6383 ) );
  NAND2_X2 _f_permutation__U4978  ( .A1(_f_permutation__n7198 ), .A2(out[129]), 
        .ZN(_f_permutation__n6384 ) );
  NAND2_X2 _f_permutation__U4977  ( .A1(_f_permutation__n6383 ), .A2(
        _f_permutation__n6384 ), .ZN(_f_permutation__n4114 ) );
  NAND2_X2 _f_permutation__U4976  ( .A1(_f_permutation__round_out[1272]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6381 ) );
  NAND2_X2 _f_permutation__U4975  ( .A1(_f_permutation__n7198 ), .A2(out[128]), 
        .ZN(_f_permutation__n6382 ) );
  NAND2_X2 _f_permutation__U4974  ( .A1(_f_permutation__n6381 ), .A2(
        _f_permutation__n6382 ), .ZN(_f_permutation__n4115 ) );
  NAND2_X2 _f_permutation__U4973  ( .A1(_f_permutation__round_out[1271]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6379 ) );
  NAND2_X2 _f_permutation__U4972  ( .A1(_f_permutation__n7198 ), .A2(out[143]), 
        .ZN(_f_permutation__n6380 ) );
  NAND2_X2 _f_permutation__U4971  ( .A1(_f_permutation__n6379 ), .A2(
        _f_permutation__n6380 ), .ZN(_f_permutation__n4116 ) );
  NAND2_X2 _f_permutation__U4970  ( .A1(_f_permutation__round_out[1270]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6377 ) );
  NAND2_X2 _f_permutation__U4969  ( .A1(_f_permutation__n7198 ), .A2(out[142]), 
        .ZN(_f_permutation__n6378 ) );
  NAND2_X2 _f_permutation__U4968  ( .A1(_f_permutation__n6377 ), .A2(
        _f_permutation__n6378 ), .ZN(_f_permutation__n4117 ) );
  NAND2_X2 _f_permutation__U4967  ( .A1(_f_permutation__round_out[1269]), 
        .A2(_f_permutation__n7104 ), .ZN(_f_permutation__n6375 ) );
  NAND2_X2 _f_permutation__U4966  ( .A1(_f_permutation__n7199 ), .A2(out[141]), 
        .ZN(_f_permutation__n6376 ) );
  NAND2_X2 _f_permutation__U4965  ( .A1(_f_permutation__n6375 ), .A2(
        _f_permutation__n6376 ), .ZN(_f_permutation__n4118 ) );
  NAND2_X2 _f_permutation__U4964  ( .A1(_f_permutation__round_out[1268]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6373 ) );
  NAND2_X2 _f_permutation__U4963  ( .A1(_f_permutation__n7199 ), .A2(out[140]), 
        .ZN(_f_permutation__n6374 ) );
  NAND2_X2 _f_permutation__U4962  ( .A1(_f_permutation__n6373 ), .A2(
        _f_permutation__n6374 ), .ZN(_f_permutation__n4119 ) );
  NAND2_X2 _f_permutation__U4961  ( .A1(_f_permutation__round_out[1267]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6371 ) );
  NAND2_X2 _f_permutation__U4960  ( .A1(_f_permutation__n7199 ), .A2(out[139]), 
        .ZN(_f_permutation__n6372 ) );
  NAND2_X2 _f_permutation__U4959  ( .A1(_f_permutation__n6371 ), .A2(
        _f_permutation__n6372 ), .ZN(_f_permutation__n4120 ) );
  NAND2_X2 _f_permutation__U4958  ( .A1(_f_permutation__round_out[1266]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6369 ) );
  NAND2_X2 _f_permutation__U4957  ( .A1(_f_permutation__n7199 ), .A2(out[138]), 
        .ZN(_f_permutation__n6370 ) );
  NAND2_X2 _f_permutation__U4956  ( .A1(_f_permutation__n6369 ), .A2(
        _f_permutation__n6370 ), .ZN(_f_permutation__n4121 ) );
  NAND2_X2 _f_permutation__U4955  ( .A1(_f_permutation__round_out[1265]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6367 ) );
  NAND2_X2 _f_permutation__U4954  ( .A1(_f_permutation__n7199 ), .A2(out[137]), 
        .ZN(_f_permutation__n6368 ) );
  NAND2_X2 _f_permutation__U4953  ( .A1(_f_permutation__n6367 ), .A2(
        _f_permutation__n6368 ), .ZN(_f_permutation__n4122 ) );
  NAND2_X2 _f_permutation__U4952  ( .A1(_f_permutation__round_out[1264]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6365 ) );
  NAND2_X2 _f_permutation__U4951  ( .A1(_f_permutation__n7199 ), .A2(out[136]), 
        .ZN(_f_permutation__n6366 ) );
  NAND2_X2 _f_permutation__U4950  ( .A1(_f_permutation__n6365 ), .A2(
        _f_permutation__n6366 ), .ZN(_f_permutation__n4123 ) );
  NAND2_X2 _f_permutation__U4949  ( .A1(_f_permutation__round_out[1263]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6363 ) );
  NAND2_X2 _f_permutation__U4948  ( .A1(_f_permutation__n7199 ), .A2(out[151]), 
        .ZN(_f_permutation__n6364 ) );
  NAND2_X2 _f_permutation__U4947  ( .A1(_f_permutation__n6363 ), .A2(
        _f_permutation__n6364 ), .ZN(_f_permutation__n4124 ) );
  NAND2_X2 _f_permutation__U4946  ( .A1(_f_permutation__round_out[1262]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6361 ) );
  NAND2_X2 _f_permutation__U4945  ( .A1(_f_permutation__n7199 ), .A2(out[150]), 
        .ZN(_f_permutation__n6362 ) );
  NAND2_X2 _f_permutation__U4944  ( .A1(_f_permutation__n6361 ), .A2(
        _f_permutation__n6362 ), .ZN(_f_permutation__n4125 ) );
  NAND2_X2 _f_permutation__U4943  ( .A1(_f_permutation__round_out[1261]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6359 ) );
  NAND2_X2 _f_permutation__U4942  ( .A1(_f_permutation__n7199 ), .A2(out[149]), 
        .ZN(_f_permutation__n6360 ) );
  NAND2_X2 _f_permutation__U4941  ( .A1(_f_permutation__n6359 ), .A2(
        _f_permutation__n6360 ), .ZN(_f_permutation__n4126 ) );
  NAND2_X2 _f_permutation__U4940  ( .A1(_f_permutation__round_out[1260]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6357 ) );
  NAND2_X2 _f_permutation__U4939  ( .A1(_f_permutation__n7199 ), .A2(out[148]), 
        .ZN(_f_permutation__n6358 ) );
  NAND2_X2 _f_permutation__U4938  ( .A1(_f_permutation__n6357 ), .A2(
        _f_permutation__n6358 ), .ZN(_f_permutation__n4127 ) );
  NAND2_X2 _f_permutation__U4937  ( .A1(_f_permutation__round_out[1259]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6355 ) );
  NAND2_X2 _f_permutation__U4936  ( .A1(_f_permutation__n7199 ), .A2(out[147]), 
        .ZN(_f_permutation__n6356 ) );
  NAND2_X2 _f_permutation__U4935  ( .A1(_f_permutation__n6355 ), .A2(
        _f_permutation__n6356 ), .ZN(_f_permutation__n4128 ) );
  NAND2_X2 _f_permutation__U4934  ( .A1(_f_permutation__round_out[1258]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6353 ) );
  NAND2_X2 _f_permutation__U4933  ( .A1(_f_permutation__n7200 ), .A2(out[146]), 
        .ZN(_f_permutation__n6354 ) );
  NAND2_X2 _f_permutation__U4932  ( .A1(_f_permutation__n6353 ), .A2(
        _f_permutation__n6354 ), .ZN(_f_permutation__n4129 ) );
  NAND2_X2 _f_permutation__U4931  ( .A1(_f_permutation__round_out[1257]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6351 ) );
  NAND2_X2 _f_permutation__U4930  ( .A1(_f_permutation__n7200 ), .A2(out[145]), 
        .ZN(_f_permutation__n6352 ) );
  NAND2_X2 _f_permutation__U4929  ( .A1(_f_permutation__n6351 ), .A2(
        _f_permutation__n6352 ), .ZN(_f_permutation__n4130 ) );
  NAND2_X2 _f_permutation__U4928  ( .A1(_f_permutation__round_out[1256]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6349 ) );
  NAND2_X2 _f_permutation__U4927  ( .A1(_f_permutation__n7200 ), .A2(out[144]), 
        .ZN(_f_permutation__n6350 ) );
  NAND2_X2 _f_permutation__U4926  ( .A1(_f_permutation__n6349 ), .A2(
        _f_permutation__n6350 ), .ZN(_f_permutation__n4131 ) );
  NAND2_X2 _f_permutation__U4925  ( .A1(_f_permutation__round_out[1255]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6347 ) );
  NAND2_X2 _f_permutation__U4924  ( .A1(_f_permutation__n7200 ), .A2(out[159]), 
        .ZN(_f_permutation__n6348 ) );
  NAND2_X2 _f_permutation__U4923  ( .A1(_f_permutation__n6347 ), .A2(
        _f_permutation__n6348 ), .ZN(_f_permutation__n4132 ) );
  NAND2_X2 _f_permutation__U4922  ( .A1(_f_permutation__round_out[1254]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6345 ) );
  NAND2_X2 _f_permutation__U4921  ( .A1(_f_permutation__n7200 ), .A2(out[158]), 
        .ZN(_f_permutation__n6346 ) );
  NAND2_X2 _f_permutation__U4920  ( .A1(_f_permutation__n6345 ), .A2(
        _f_permutation__n6346 ), .ZN(_f_permutation__n4133 ) );
  NAND2_X2 _f_permutation__U4919  ( .A1(_f_permutation__round_out[1253]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6343 ) );
  NAND2_X2 _f_permutation__U4918  ( .A1(_f_permutation__n7200 ), .A2(out[157]), 
        .ZN(_f_permutation__n6344 ) );
  NAND2_X2 _f_permutation__U4917  ( .A1(_f_permutation__n6343 ), .A2(
        _f_permutation__n6344 ), .ZN(_f_permutation__n4134 ) );
  NAND2_X2 _f_permutation__U4916  ( .A1(_f_permutation__round_out[1252]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6341 ) );
  NAND2_X2 _f_permutation__U4915  ( .A1(_f_permutation__n7200 ), .A2(out[156]), 
        .ZN(_f_permutation__n6342 ) );
  NAND2_X2 _f_permutation__U4914  ( .A1(_f_permutation__n6341 ), .A2(
        _f_permutation__n6342 ), .ZN(_f_permutation__n4135 ) );
  NAND2_X2 _f_permutation__U4913  ( .A1(_f_permutation__round_out[1251]), 
        .A2(_f_permutation__n7103 ), .ZN(_f_permutation__n6339 ) );
  NAND2_X2 _f_permutation__U4912  ( .A1(_f_permutation__n7200 ), .A2(out[155]), 
        .ZN(_f_permutation__n6340 ) );
  NAND2_X2 _f_permutation__U4911  ( .A1(_f_permutation__n6339 ), .A2(
        _f_permutation__n6340 ), .ZN(_f_permutation__n4136 ) );
  NAND2_X2 _f_permutation__U4910  ( .A1(_f_permutation__round_out[1250]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6337 ) );
  NAND2_X2 _f_permutation__U4909  ( .A1(_f_permutation__n7200 ), .A2(out[154]), 
        .ZN(_f_permutation__n6338 ) );
  NAND2_X2 _f_permutation__U4908  ( .A1(_f_permutation__n6337 ), .A2(
        _f_permutation__n6338 ), .ZN(_f_permutation__n4137 ) );
  NAND2_X2 _f_permutation__U4907  ( .A1(_f_permutation__round_out[1249]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6335 ) );
  NAND2_X2 _f_permutation__U4906  ( .A1(_f_permutation__n7200 ), .A2(out[153]), 
        .ZN(_f_permutation__n6336 ) );
  NAND2_X2 _f_permutation__U4905  ( .A1(_f_permutation__n6335 ), .A2(
        _f_permutation__n6336 ), .ZN(_f_permutation__n4138 ) );
  NAND2_X2 _f_permutation__U4904  ( .A1(_f_permutation__round_out[1248]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6333 ) );
  NAND2_X2 _f_permutation__U4903  ( .A1(_f_permutation__n7200 ), .A2(out[152]), 
        .ZN(_f_permutation__n6334 ) );
  NAND2_X2 _f_permutation__U4902  ( .A1(_f_permutation__n6333 ), .A2(
        _f_permutation__n6334 ), .ZN(_f_permutation__n4139 ) );
  NAND2_X2 _f_permutation__U4901  ( .A1(_f_permutation__round_out[1247]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6331 ) );
  NAND2_X2 _f_permutation__U4900  ( .A1(_f_permutation__n7201 ), .A2(out[167]), 
        .ZN(_f_permutation__n6332 ) );
  NAND2_X2 _f_permutation__U4899  ( .A1(_f_permutation__n6331 ), .A2(
        _f_permutation__n6332 ), .ZN(_f_permutation__n4140 ) );
  NAND2_X2 _f_permutation__U4898  ( .A1(_f_permutation__round_out[1246]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6329 ) );
  NAND2_X2 _f_permutation__U4897  ( .A1(_f_permutation__n7201 ), .A2(out[166]), 
        .ZN(_f_permutation__n6330 ) );
  NAND2_X2 _f_permutation__U4896  ( .A1(_f_permutation__n6329 ), .A2(
        _f_permutation__n6330 ), .ZN(_f_permutation__n4141 ) );
  NAND2_X2 _f_permutation__U4895  ( .A1(_f_permutation__round_out[1245]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6327 ) );
  NAND2_X2 _f_permutation__U4894  ( .A1(_f_permutation__n7201 ), .A2(out[165]), 
        .ZN(_f_permutation__n6328 ) );
  NAND2_X2 _f_permutation__U4893  ( .A1(_f_permutation__n6327 ), .A2(
        _f_permutation__n6328 ), .ZN(_f_permutation__n4142 ) );
  NAND2_X2 _f_permutation__U4892  ( .A1(_f_permutation__round_out[1244]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6325 ) );
  NAND2_X2 _f_permutation__U4891  ( .A1(_f_permutation__n7201 ), .A2(out[164]), 
        .ZN(_f_permutation__n6326 ) );
  NAND2_X2 _f_permutation__U4890  ( .A1(_f_permutation__n6325 ), .A2(
        _f_permutation__n6326 ), .ZN(_f_permutation__n4143 ) );
  NAND2_X2 _f_permutation__U4889  ( .A1(_f_permutation__round_out[1243]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6323 ) );
  NAND2_X2 _f_permutation__U4888  ( .A1(_f_permutation__n7201 ), .A2(out[163]), 
        .ZN(_f_permutation__n6324 ) );
  NAND2_X2 _f_permutation__U4887  ( .A1(_f_permutation__n6323 ), .A2(
        _f_permutation__n6324 ), .ZN(_f_permutation__n4144 ) );
  NAND2_X2 _f_permutation__U4886  ( .A1(_f_permutation__round_out[1242]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6321 ) );
  NAND2_X2 _f_permutation__U4885  ( .A1(_f_permutation__n7201 ), .A2(out[162]), 
        .ZN(_f_permutation__n6322 ) );
  NAND2_X2 _f_permutation__U4884  ( .A1(_f_permutation__n6321 ), .A2(
        _f_permutation__n6322 ), .ZN(_f_permutation__n4145 ) );
  NAND2_X2 _f_permutation__U4883  ( .A1(_f_permutation__round_out[1241]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6319 ) );
  NAND2_X2 _f_permutation__U4882  ( .A1(_f_permutation__n7201 ), .A2(out[161]), 
        .ZN(_f_permutation__n6320 ) );
  NAND2_X2 _f_permutation__U4881  ( .A1(_f_permutation__n6319 ), .A2(
        _f_permutation__n6320 ), .ZN(_f_permutation__n4146 ) );
  NAND2_X2 _f_permutation__U4880  ( .A1(_f_permutation__round_out[1240]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6317 ) );
  NAND2_X2 _f_permutation__U4879  ( .A1(_f_permutation__n7201 ), .A2(out[160]), 
        .ZN(_f_permutation__n6318 ) );
  NAND2_X2 _f_permutation__U4878  ( .A1(_f_permutation__n6317 ), .A2(
        _f_permutation__n6318 ), .ZN(_f_permutation__n4147 ) );
  NAND2_X2 _f_permutation__U4877  ( .A1(_f_permutation__round_out[1239]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6315 ) );
  NAND2_X2 _f_permutation__U4876  ( .A1(_f_permutation__n7201 ), .A2(out[175]), 
        .ZN(_f_permutation__n6316 ) );
  NAND2_X2 _f_permutation__U4875  ( .A1(_f_permutation__n6315 ), .A2(
        _f_permutation__n6316 ), .ZN(_f_permutation__n4148 ) );
  NAND2_X2 _f_permutation__U4874  ( .A1(_f_permutation__round_out[1238]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6313 ) );
  NAND2_X2 _f_permutation__U4873  ( .A1(_f_permutation__n7201 ), .A2(out[174]), 
        .ZN(_f_permutation__n6314 ) );
  NAND2_X2 _f_permutation__U4872  ( .A1(_f_permutation__n6313 ), .A2(
        _f_permutation__n6314 ), .ZN(_f_permutation__n4149 ) );
  NAND2_X2 _f_permutation__U4871  ( .A1(_f_permutation__round_out[1237]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6311 ) );
  NAND2_X2 _f_permutation__U4870  ( .A1(_f_permutation__n7201 ), .A2(out[173]), 
        .ZN(_f_permutation__n6312 ) );
  NAND2_X2 _f_permutation__U4869  ( .A1(_f_permutation__n6311 ), .A2(
        _f_permutation__n6312 ), .ZN(_f_permutation__n4150 ) );
  NAND2_X2 _f_permutation__U4868  ( .A1(_f_permutation__round_out[1236]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6309 ) );
  NAND2_X2 _f_permutation__U4867  ( .A1(_f_permutation__n7202 ), .A2(out[172]), 
        .ZN(_f_permutation__n6310 ) );
  NAND2_X2 _f_permutation__U4866  ( .A1(_f_permutation__n6309 ), .A2(
        _f_permutation__n6310 ), .ZN(_f_permutation__n4151 ) );
  NAND2_X2 _f_permutation__U4865  ( .A1(_f_permutation__round_out[1235]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6307 ) );
  NAND2_X2 _f_permutation__U4864  ( .A1(_f_permutation__n7202 ), .A2(out[171]), 
        .ZN(_f_permutation__n6308 ) );
  NAND2_X2 _f_permutation__U4863  ( .A1(_f_permutation__n6307 ), .A2(
        _f_permutation__n6308 ), .ZN(_f_permutation__n4152 ) );
  NAND2_X2 _f_permutation__U4862  ( .A1(_f_permutation__round_out[1234]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6305 ) );
  NAND2_X2 _f_permutation__U4861  ( .A1(_f_permutation__n7202 ), .A2(out[170]), 
        .ZN(_f_permutation__n6306 ) );
  NAND2_X2 _f_permutation__U4860  ( .A1(_f_permutation__n6305 ), .A2(
        _f_permutation__n6306 ), .ZN(_f_permutation__n4153 ) );
  NAND2_X2 _f_permutation__U4859  ( .A1(_f_permutation__round_out[1233]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6303 ) );
  NAND2_X2 _f_permutation__U4858  ( .A1(_f_permutation__n7202 ), .A2(out[169]), 
        .ZN(_f_permutation__n6304 ) );
  NAND2_X2 _f_permutation__U4857  ( .A1(_f_permutation__n6303 ), .A2(
        _f_permutation__n6304 ), .ZN(_f_permutation__n4154 ) );
  NAND2_X2 _f_permutation__U4856  ( .A1(_f_permutation__round_out[1232]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6301 ) );
  NAND2_X2 _f_permutation__U4855  ( .A1(_f_permutation__n7202 ), .A2(out[168]), 
        .ZN(_f_permutation__n6302 ) );
  NAND2_X2 _f_permutation__U4854  ( .A1(_f_permutation__n6301 ), .A2(
        _f_permutation__n6302 ), .ZN(_f_permutation__n4155 ) );
  NAND2_X2 _f_permutation__U4853  ( .A1(_f_permutation__round_out[1231]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6299 ) );
  NAND2_X2 _f_permutation__U4852  ( .A1(_f_permutation__n7202 ), .A2(out[183]), 
        .ZN(_f_permutation__n6300 ) );
  NAND2_X2 _f_permutation__U4851  ( .A1(_f_permutation__n6299 ), .A2(
        _f_permutation__n6300 ), .ZN(_f_permutation__n4156 ) );
  NAND2_X2 _f_permutation__U4850  ( .A1(_f_permutation__round_out[1230]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6297 ) );
  NAND2_X2 _f_permutation__U4849  ( .A1(_f_permutation__n7202 ), .A2(out[182]), 
        .ZN(_f_permutation__n6298 ) );
  NAND2_X2 _f_permutation__U4848  ( .A1(_f_permutation__n6297 ), .A2(
        _f_permutation__n6298 ), .ZN(_f_permutation__n4157 ) );
  NAND2_X2 _f_permutation__U4847  ( .A1(_f_permutation__round_out[1229]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6295 ) );
  NAND2_X2 _f_permutation__U4846  ( .A1(_f_permutation__n7202 ), .A2(out[181]), 
        .ZN(_f_permutation__n6296 ) );
  NAND2_X2 _f_permutation__U4845  ( .A1(_f_permutation__n6295 ), .A2(
        _f_permutation__n6296 ), .ZN(_f_permutation__n4158 ) );
  NAND2_X2 _f_permutation__U4844  ( .A1(_f_permutation__round_out[1228]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6293 ) );
  NAND2_X2 _f_permutation__U4843  ( .A1(_f_permutation__n7202 ), .A2(out[180]), 
        .ZN(_f_permutation__n6294 ) );
  NAND2_X2 _f_permutation__U4842  ( .A1(_f_permutation__n6293 ), .A2(
        _f_permutation__n6294 ), .ZN(_f_permutation__n4159 ) );
  NAND2_X2 _f_permutation__U4841  ( .A1(_f_permutation__round_out[1227]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6291 ) );
  NAND2_X2 _f_permutation__U4840  ( .A1(_f_permutation__n7202 ), .A2(out[179]), 
        .ZN(_f_permutation__n6292 ) );
  NAND2_X2 _f_permutation__U4839  ( .A1(_f_permutation__n6291 ), .A2(
        _f_permutation__n6292 ), .ZN(_f_permutation__n4160 ) );
  NAND2_X2 _f_permutation__U4838  ( .A1(_f_permutation__round_out[1226]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6289 ) );
  NAND2_X2 _f_permutation__U4837  ( .A1(_f_permutation__n7202 ), .A2(out[178]), 
        .ZN(_f_permutation__n6290 ) );
  NAND2_X2 _f_permutation__U4836  ( .A1(_f_permutation__n6289 ), .A2(
        _f_permutation__n6290 ), .ZN(_f_permutation__n4161 ) );
  NAND2_X2 _f_permutation__U4835  ( .A1(_f_permutation__round_out[1225]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6287 ) );
  NAND2_X2 _f_permutation__U4834  ( .A1(_f_permutation__n7203 ), .A2(out[177]), 
        .ZN(_f_permutation__n6288 ) );
  NAND2_X2 _f_permutation__U4833  ( .A1(_f_permutation__n6287 ), .A2(
        _f_permutation__n6288 ), .ZN(_f_permutation__n4162 ) );
  NAND2_X2 _f_permutation__U4832  ( .A1(_f_permutation__round_out[1224]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6285 ) );
  NAND2_X2 _f_permutation__U4831  ( .A1(_f_permutation__n7203 ), .A2(out[176]), 
        .ZN(_f_permutation__n6286 ) );
  NAND2_X2 _f_permutation__U4830  ( .A1(_f_permutation__n6285 ), .A2(
        _f_permutation__n6286 ), .ZN(_f_permutation__n4163 ) );
  NAND2_X2 _f_permutation__U4829  ( .A1(_f_permutation__round_out[1223]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6283 ) );
  NAND2_X2 _f_permutation__U4828  ( .A1(_f_permutation__n7203 ), .A2(out[191]), 
        .ZN(_f_permutation__n6284 ) );
  NAND2_X2 _f_permutation__U4827  ( .A1(_f_permutation__n6283 ), .A2(
        _f_permutation__n6284 ), .ZN(_f_permutation__n4164 ) );
  NAND2_X2 _f_permutation__U4826  ( .A1(_f_permutation__round_out[1222]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6281 ) );
  NAND2_X2 _f_permutation__U4825  ( .A1(_f_permutation__n7203 ), .A2(out[190]), 
        .ZN(_f_permutation__n6282 ) );
  NAND2_X2 _f_permutation__U4824  ( .A1(_f_permutation__n6281 ), .A2(
        _f_permutation__n6282 ), .ZN(_f_permutation__n4165 ) );
  NAND2_X2 _f_permutation__U4823  ( .A1(_f_permutation__round_out[1221]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6279 ) );
  NAND2_X2 _f_permutation__U4822  ( .A1(_f_permutation__n7203 ), .A2(out[189]), 
        .ZN(_f_permutation__n6280 ) );
  NAND2_X2 _f_permutation__U4821  ( .A1(_f_permutation__n6279 ), .A2(
        _f_permutation__n6280 ), .ZN(_f_permutation__n4166 ) );
  NAND2_X2 _f_permutation__U4820  ( .A1(_f_permutation__round_out[1220]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6277 ) );
  NAND2_X2 _f_permutation__U4819  ( .A1(_f_permutation__n7203 ), .A2(out[188]), 
        .ZN(_f_permutation__n6278 ) );
  NAND2_X2 _f_permutation__U4818  ( .A1(_f_permutation__n6277 ), .A2(
        _f_permutation__n6278 ), .ZN(_f_permutation__n4167 ) );
  NAND2_X2 _f_permutation__U4817  ( .A1(_f_permutation__round_out[1219]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6275 ) );
  NAND2_X2 _f_permutation__U4816  ( .A1(_f_permutation__n7203 ), .A2(out[187]), 
        .ZN(_f_permutation__n6276 ) );
  NAND2_X2 _f_permutation__U4815  ( .A1(_f_permutation__n6275 ), .A2(
        _f_permutation__n6276 ), .ZN(_f_permutation__n4168 ) );
  NAND2_X2 _f_permutation__U4814  ( .A1(_f_permutation__round_out[1218]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6273 ) );
  NAND2_X2 _f_permutation__U4813  ( .A1(_f_permutation__n7203 ), .A2(out[186]), 
        .ZN(_f_permutation__n6274 ) );
  NAND2_X2 _f_permutation__U4812  ( .A1(_f_permutation__n6273 ), .A2(
        _f_permutation__n6274 ), .ZN(_f_permutation__n4169 ) );
  NAND2_X2 _f_permutation__U4811  ( .A1(_f_permutation__round_out[1217]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6271 ) );
  NAND2_X2 _f_permutation__U4810  ( .A1(_f_permutation__n7203 ), .A2(out[185]), 
        .ZN(_f_permutation__n6272 ) );
  NAND2_X2 _f_permutation__U4809  ( .A1(_f_permutation__n6271 ), .A2(
        _f_permutation__n6272 ), .ZN(_f_permutation__n4170 ) );
  NAND2_X2 _f_permutation__U4808  ( .A1(_f_permutation__round_out[1216]), 
        .A2(_f_permutation__n7101 ), .ZN(_f_permutation__n6269 ) );
  NAND2_X2 _f_permutation__U4807  ( .A1(_f_permutation__n7203 ), .A2(out[184]), 
        .ZN(_f_permutation__n6270 ) );
  NAND2_X2 _f_permutation__U4806  ( .A1(_f_permutation__n6269 ), .A2(
        _f_permutation__n6270 ), .ZN(_f_permutation__n4171 ) );
  NAND2_X2 _f_permutation__U4805  ( .A1(_f_permutation__round_out[1215]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6267 ) );
  NAND2_X2 _f_permutation__U4804  ( .A1(_f_permutation__n7203 ), .A2(out[71]), 
        .ZN(_f_permutation__n6268 ) );
  NAND2_X2 _f_permutation__U4803  ( .A1(_f_permutation__n6267 ), .A2(
        _f_permutation__n6268 ), .ZN(_f_permutation__n4172 ) );
  NAND2_X2 _f_permutation__U4802  ( .A1(_f_permutation__round_out[1214]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6265 ) );
  NAND2_X2 _f_permutation__U4801  ( .A1(_f_permutation__n7204 ), .A2(out[70]), 
        .ZN(_f_permutation__n6266 ) );
  NAND2_X2 _f_permutation__U4800  ( .A1(_f_permutation__n6265 ), .A2(
        _f_permutation__n6266 ), .ZN(_f_permutation__n4173 ) );
  NAND2_X2 _f_permutation__U4799  ( .A1(_f_permutation__round_out[1213]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6263 ) );
  NAND2_X2 _f_permutation__U4798  ( .A1(_f_permutation__n7204 ), .A2(out[69]), 
        .ZN(_f_permutation__n6264 ) );
  NAND2_X2 _f_permutation__U4797  ( .A1(_f_permutation__n6263 ), .A2(
        _f_permutation__n6264 ), .ZN(_f_permutation__n4174 ) );
  NAND2_X2 _f_permutation__U4796  ( .A1(_f_permutation__round_out[1212]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6261 ) );
  NAND2_X2 _f_permutation__U4795  ( .A1(_f_permutation__n7204 ), .A2(out[68]), 
        .ZN(_f_permutation__n6262 ) );
  NAND2_X2 _f_permutation__U4794  ( .A1(_f_permutation__n6261 ), .A2(
        _f_permutation__n6262 ), .ZN(_f_permutation__n4175 ) );
  NAND2_X2 _f_permutation__U4793  ( .A1(_f_permutation__round_out[1211]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6259 ) );
  NAND2_X2 _f_permutation__U4792  ( .A1(_f_permutation__n7204 ), .A2(out[67]), 
        .ZN(_f_permutation__n6260 ) );
  NAND2_X2 _f_permutation__U4791  ( .A1(_f_permutation__n6259 ), .A2(
        _f_permutation__n6260 ), .ZN(_f_permutation__n4176 ) );
  NAND2_X2 _f_permutation__U4790  ( .A1(_f_permutation__round_out[1210]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6257 ) );
  NAND2_X2 _f_permutation__U4789  ( .A1(_f_permutation__n7204 ), .A2(out[66]), 
        .ZN(_f_permutation__n6258 ) );
  NAND2_X2 _f_permutation__U4788  ( .A1(_f_permutation__n6257 ), .A2(
        _f_permutation__n6258 ), .ZN(_f_permutation__n4177 ) );
  NAND2_X2 _f_permutation__U4787  ( .A1(_f_permutation__round_out[1209]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6255 ) );
  NAND2_X2 _f_permutation__U4786  ( .A1(_f_permutation__n7204 ), .A2(out[65]), 
        .ZN(_f_permutation__n6256 ) );
  NAND2_X2 _f_permutation__U4785  ( .A1(_f_permutation__n6255 ), .A2(
        _f_permutation__n6256 ), .ZN(_f_permutation__n4178 ) );
  NAND2_X2 _f_permutation__U4784  ( .A1(_f_permutation__round_out[1208]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6253 ) );
  NAND2_X2 _f_permutation__U4783  ( .A1(_f_permutation__n7204 ), .A2(out[64]), 
        .ZN(_f_permutation__n6254 ) );
  NAND2_X2 _f_permutation__U4782  ( .A1(_f_permutation__n6253 ), .A2(
        _f_permutation__n6254 ), .ZN(_f_permutation__n4179 ) );
  NAND2_X2 _f_permutation__U4781  ( .A1(_f_permutation__round_out[1207]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6251 ) );
  NAND2_X2 _f_permutation__U4780  ( .A1(_f_permutation__n7204 ), .A2(out[79]), 
        .ZN(_f_permutation__n6252 ) );
  NAND2_X2 _f_permutation__U4779  ( .A1(_f_permutation__n6251 ), .A2(
        _f_permutation__n6252 ), .ZN(_f_permutation__n4180 ) );
  NAND2_X2 _f_permutation__U4778  ( .A1(_f_permutation__round_out[1206]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6249 ) );
  NAND2_X2 _f_permutation__U4777  ( .A1(_f_permutation__n7204 ), .A2(out[78]), 
        .ZN(_f_permutation__n6250 ) );
  NAND2_X2 _f_permutation__U4776  ( .A1(_f_permutation__n6249 ), .A2(
        _f_permutation__n6250 ), .ZN(_f_permutation__n4181 ) );
  NAND2_X2 _f_permutation__U4775  ( .A1(_f_permutation__round_out[1205]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6247 ) );
  NAND2_X2 _f_permutation__U4774  ( .A1(_f_permutation__n7204 ), .A2(out[77]), 
        .ZN(_f_permutation__n6248 ) );
  NAND2_X2 _f_permutation__U4773  ( .A1(_f_permutation__n6247 ), .A2(
        _f_permutation__n6248 ), .ZN(_f_permutation__n4182 ) );
  NAND2_X2 _f_permutation__U4772  ( .A1(_f_permutation__round_out[1204]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6245 ) );
  NAND2_X2 _f_permutation__U4771  ( .A1(_f_permutation__n7204 ), .A2(out[76]), 
        .ZN(_f_permutation__n6246 ) );
  NAND2_X2 _f_permutation__U4770  ( .A1(_f_permutation__n6245 ), .A2(
        _f_permutation__n6246 ), .ZN(_f_permutation__n4183 ) );
  NAND2_X2 _f_permutation__U4769  ( .A1(_f_permutation__round_out[1203]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6243 ) );
  NAND2_X2 _f_permutation__U4768  ( .A1(_f_permutation__n7205 ), .A2(out[75]), 
        .ZN(_f_permutation__n6244 ) );
  NAND2_X2 _f_permutation__U4767  ( .A1(_f_permutation__n6243 ), .A2(
        _f_permutation__n6244 ), .ZN(_f_permutation__n4184 ) );
  NAND2_X2 _f_permutation__U4766  ( .A1(_f_permutation__round_out[1202]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6241 ) );
  NAND2_X2 _f_permutation__U4765  ( .A1(_f_permutation__n7205 ), .A2(out[74]), 
        .ZN(_f_permutation__n6242 ) );
  NAND2_X2 _f_permutation__U4764  ( .A1(_f_permutation__n6241 ), .A2(
        _f_permutation__n6242 ), .ZN(_f_permutation__n4185 ) );
  NAND2_X2 _f_permutation__U4763  ( .A1(_f_permutation__round_out[1201]), 
        .A2(_f_permutation__n7100 ), .ZN(_f_permutation__n6239 ) );
  NAND2_X2 _f_permutation__U4762  ( .A1(_f_permutation__n7205 ), .A2(out[73]), 
        .ZN(_f_permutation__n6240 ) );
  NAND2_X2 _f_permutation__U4761  ( .A1(_f_permutation__n6239 ), .A2(
        _f_permutation__n6240 ), .ZN(_f_permutation__n4186 ) );
  NAND2_X2 _f_permutation__U4760  ( .A1(_f_permutation__round_out[1200]), 
        .A2(_f_permutation__n7102 ), .ZN(_f_permutation__n6237 ) );
  NAND2_X2 _f_permutation__U4759  ( .A1(_f_permutation__n7205 ), .A2(out[72]), 
        .ZN(_f_permutation__n6238 ) );
  NAND2_X2 _f_permutation__U4758  ( .A1(_f_permutation__n6237 ), .A2(
        _f_permutation__n6238 ), .ZN(_f_permutation__n4187 ) );
  NAND2_X2 _f_permutation__U4757  ( .A1(_f_permutation__round_out[1199]), 
        .A2(_f_permutation__n7105 ), .ZN(_f_permutation__n6235 ) );
  NAND2_X2 _f_permutation__U4756  ( .A1(_f_permutation__n7205 ), .A2(out[87]), 
        .ZN(_f_permutation__n6236 ) );
  NAND2_X2 _f_permutation__U4755  ( .A1(_f_permutation__n6235 ), .A2(
        _f_permutation__n6236 ), .ZN(_f_permutation__n4188 ) );
  NAND2_X2 _f_permutation__U4754  ( .A1(_f_permutation__round_out[1198]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n6233 ) );
  NAND2_X2 _f_permutation__U4753  ( .A1(_f_permutation__n7205 ), .A2(out[86]), 
        .ZN(_f_permutation__n6234 ) );
  NAND2_X2 _f_permutation__U4752  ( .A1(_f_permutation__n6233 ), .A2(
        _f_permutation__n6234 ), .ZN(_f_permutation__n4189 ) );
  NAND2_X2 _f_permutation__U4751  ( .A1(_f_permutation__round_out[1197]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n6231 ) );
  NAND2_X2 _f_permutation__U4750  ( .A1(_f_permutation__n7205 ), .A2(out[85]), 
        .ZN(_f_permutation__n6232 ) );
  NAND2_X2 _f_permutation__U4749  ( .A1(_f_permutation__n6231 ), .A2(
        _f_permutation__n6232 ), .ZN(_f_permutation__n4190 ) );
  NAND2_X2 _f_permutation__U4748  ( .A1(_f_permutation__round_out[1196]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n6229 ) );
  NAND2_X2 _f_permutation__U4747  ( .A1(_f_permutation__n7205 ), .A2(out[84]), 
        .ZN(_f_permutation__n6230 ) );
  NAND2_X2 _f_permutation__U4746  ( .A1(_f_permutation__n6229 ), .A2(
        _f_permutation__n6230 ), .ZN(_f_permutation__n4191 ) );
  NAND2_X2 _f_permutation__U4745  ( .A1(_f_permutation__round_out[1195]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n6227 ) );
  NAND2_X2 _f_permutation__U4744  ( .A1(_f_permutation__n7205 ), .A2(out[83]), 
        .ZN(_f_permutation__n6228 ) );
  NAND2_X2 _f_permutation__U4743  ( .A1(_f_permutation__n6227 ), .A2(
        _f_permutation__n6228 ), .ZN(_f_permutation__n4192 ) );
  NAND2_X2 _f_permutation__U4742  ( .A1(_f_permutation__round_out[1194]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n6225 ) );
  NAND2_X2 _f_permutation__U4741  ( .A1(_f_permutation__n7205 ), .A2(out[82]), 
        .ZN(_f_permutation__n6226 ) );
  NAND2_X2 _f_permutation__U4740  ( .A1(_f_permutation__n6225 ), .A2(
        _f_permutation__n6226 ), .ZN(_f_permutation__n4193 ) );
  NAND2_X2 _f_permutation__U4739  ( .A1(_f_permutation__round_out[1193]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n6223 ) );
  NAND2_X2 _f_permutation__U4738  ( .A1(_f_permutation__n7205 ), .A2(out[81]), 
        .ZN(_f_permutation__n6224 ) );
  NAND2_X2 _f_permutation__U4737  ( .A1(_f_permutation__n6223 ), .A2(
        _f_permutation__n6224 ), .ZN(_f_permutation__n4194 ) );
  NAND2_X2 _f_permutation__U4736  ( .A1(_f_permutation__round_out[1192]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n6221 ) );
  NAND2_X2 _f_permutation__U4735  ( .A1(_f_permutation__n7206 ), .A2(out[80]), 
        .ZN(_f_permutation__n6222 ) );
  NAND2_X2 _f_permutation__U4734  ( .A1(_f_permutation__n6221 ), .A2(
        _f_permutation__n6222 ), .ZN(_f_permutation__n4195 ) );
  NAND2_X2 _f_permutation__U4733  ( .A1(_f_permutation__round_out[1191]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n6219 ) );
  NAND2_X2 _f_permutation__U4732  ( .A1(_f_permutation__n7206 ), .A2(out[95]), 
        .ZN(_f_permutation__n6220 ) );
  NAND2_X2 _f_permutation__U4731  ( .A1(_f_permutation__n6219 ), .A2(
        _f_permutation__n6220 ), .ZN(_f_permutation__n4196 ) );
  NAND2_X2 _f_permutation__U4730  ( .A1(_f_permutation__round_out[1190]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n6217 ) );
  NAND2_X2 _f_permutation__U4729  ( .A1(_f_permutation__n7206 ), .A2(out[94]), 
        .ZN(_f_permutation__n6218 ) );
  NAND2_X2 _f_permutation__U4728  ( .A1(_f_permutation__n6217 ), .A2(
        _f_permutation__n6218 ), .ZN(_f_permutation__n4197 ) );
  NAND2_X2 _f_permutation__U4727  ( .A1(_f_permutation__round_out[1189]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6215 ) );
  NAND2_X2 _f_permutation__U4726  ( .A1(_f_permutation__n7206 ), .A2(out[93]), 
        .ZN(_f_permutation__n6216 ) );
  NAND2_X2 _f_permutation__U4725  ( .A1(_f_permutation__n6215 ), .A2(
        _f_permutation__n6216 ), .ZN(_f_permutation__n4198 ) );
  NAND2_X2 _f_permutation__U4724  ( .A1(_f_permutation__round_out[1188]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6213 ) );
  NAND2_X2 _f_permutation__U4723  ( .A1(_f_permutation__n7206 ), .A2(out[92]), 
        .ZN(_f_permutation__n6214 ) );
  NAND2_X2 _f_permutation__U4722  ( .A1(_f_permutation__n6213 ), .A2(
        _f_permutation__n6214 ), .ZN(_f_permutation__n4199 ) );
  NAND2_X2 _f_permutation__U4721  ( .A1(_f_permutation__round_out[1187]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6211 ) );
  NAND2_X2 _f_permutation__U4720  ( .A1(_f_permutation__n7206 ), .A2(out[91]), 
        .ZN(_f_permutation__n6212 ) );
  NAND2_X2 _f_permutation__U4719  ( .A1(_f_permutation__n6211 ), .A2(
        _f_permutation__n6212 ), .ZN(_f_permutation__n4200 ) );
  NAND2_X2 _f_permutation__U4718  ( .A1(_f_permutation__round_out[1186]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6209 ) );
  NAND2_X2 _f_permutation__U4717  ( .A1(_f_permutation__n7206 ), .A2(out[90]), 
        .ZN(_f_permutation__n6210 ) );
  NAND2_X2 _f_permutation__U4716  ( .A1(_f_permutation__n6209 ), .A2(
        _f_permutation__n6210 ), .ZN(_f_permutation__n4201 ) );
  NAND2_X2 _f_permutation__U4715  ( .A1(_f_permutation__round_out[1185]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6207 ) );
  NAND2_X2 _f_permutation__U4714  ( .A1(_f_permutation__n7206 ), .A2(out[89]), 
        .ZN(_f_permutation__n6208 ) );
  NAND2_X2 _f_permutation__U4713  ( .A1(_f_permutation__n6207 ), .A2(
        _f_permutation__n6208 ), .ZN(_f_permutation__n4202 ) );
  NAND2_X2 _f_permutation__U4712  ( .A1(_f_permutation__round_out[1184]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6205 ) );
  NAND2_X2 _f_permutation__U4711  ( .A1(_f_permutation__n7206 ), .A2(out[88]), 
        .ZN(_f_permutation__n6206 ) );
  NAND2_X2 _f_permutation__U4710  ( .A1(_f_permutation__n6205 ), .A2(
        _f_permutation__n6206 ), .ZN(_f_permutation__n4203 ) );
  NAND2_X2 _f_permutation__U4709  ( .A1(_f_permutation__round_out[1183]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6203 ) );
  NAND2_X2 _f_permutation__U4708  ( .A1(_f_permutation__n7206 ), .A2(out[103]), 
        .ZN(_f_permutation__n6204 ) );
  NAND2_X2 _f_permutation__U4707  ( .A1(_f_permutation__n6203 ), .A2(
        _f_permutation__n6204 ), .ZN(_f_permutation__n4204 ) );
  NAND2_X2 _f_permutation__U4706  ( .A1(_f_permutation__round_out[1182]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6201 ) );
  NAND2_X2 _f_permutation__U4705  ( .A1(_f_permutation__n7206 ), .A2(out[102]), 
        .ZN(_f_permutation__n6202 ) );
  NAND2_X2 _f_permutation__U4704  ( .A1(_f_permutation__n6201 ), .A2(
        _f_permutation__n6202 ), .ZN(_f_permutation__n4205 ) );
  NAND2_X2 _f_permutation__U4703  ( .A1(_f_permutation__round_out[1181]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6199 ) );
  NAND2_X2 _f_permutation__U4702  ( .A1(_f_permutation__n7207 ), .A2(out[101]), 
        .ZN(_f_permutation__n6200 ) );
  NAND2_X2 _f_permutation__U4701  ( .A1(_f_permutation__n6199 ), .A2(
        _f_permutation__n6200 ), .ZN(_f_permutation__n4206 ) );
  NAND2_X2 _f_permutation__U4700  ( .A1(_f_permutation__round_out[1180]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6197 ) );
  NAND2_X2 _f_permutation__U4699  ( .A1(_f_permutation__n7207 ), .A2(out[100]), 
        .ZN(_f_permutation__n6198 ) );
  NAND2_X2 _f_permutation__U4698  ( .A1(_f_permutation__n6197 ), .A2(
        _f_permutation__n6198 ), .ZN(_f_permutation__n4207 ) );
  NAND2_X2 _f_permutation__U4697  ( .A1(_f_permutation__round_out[1179]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6195 ) );
  NAND2_X2 _f_permutation__U4696  ( .A1(_f_permutation__n7207 ), .A2(out[99]), 
        .ZN(_f_permutation__n6196 ) );
  NAND2_X2 _f_permutation__U4695  ( .A1(_f_permutation__n6195 ), .A2(
        _f_permutation__n6196 ), .ZN(_f_permutation__n4208 ) );
  NAND2_X2 _f_permutation__U4694  ( .A1(_f_permutation__round_out[1178]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6193 ) );
  NAND2_X2 _f_permutation__U4693  ( .A1(_f_permutation__n7207 ), .A2(out[98]), 
        .ZN(_f_permutation__n6194 ) );
  NAND2_X2 _f_permutation__U4692  ( .A1(_f_permutation__n6193 ), .A2(
        _f_permutation__n6194 ), .ZN(_f_permutation__n4209 ) );
  NAND2_X2 _f_permutation__U4691  ( .A1(_f_permutation__round_out[1177]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6191 ) );
  NAND2_X2 _f_permutation__U4690  ( .A1(_f_permutation__n7207 ), .A2(out[97]), 
        .ZN(_f_permutation__n6192 ) );
  NAND2_X2 _f_permutation__U4689  ( .A1(_f_permutation__n6191 ), .A2(
        _f_permutation__n6192 ), .ZN(_f_permutation__n4210 ) );
  NAND2_X2 _f_permutation__U4688  ( .A1(_f_permutation__round_out[1176]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6189 ) );
  NAND2_X2 _f_permutation__U4687  ( .A1(_f_permutation__n7207 ), .A2(out[96]), 
        .ZN(_f_permutation__n6190 ) );
  NAND2_X2 _f_permutation__U4686  ( .A1(_f_permutation__n6189 ), .A2(
        _f_permutation__n6190 ), .ZN(_f_permutation__n4211 ) );
  NAND2_X2 _f_permutation__U4685  ( .A1(_f_permutation__round_out[1175]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6187 ) );
  NAND2_X2 _f_permutation__U4684  ( .A1(_f_permutation__n7207 ), .A2(out[111]), 
        .ZN(_f_permutation__n6188 ) );
  NAND2_X2 _f_permutation__U4683  ( .A1(_f_permutation__n6187 ), .A2(
        _f_permutation__n6188 ), .ZN(_f_permutation__n4212 ) );
  NAND2_X2 _f_permutation__U4682  ( .A1(_f_permutation__round_out[1174]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6185 ) );
  NAND2_X2 _f_permutation__U4681  ( .A1(_f_permutation__n7207 ), .A2(out[110]), 
        .ZN(_f_permutation__n6186 ) );
  NAND2_X2 _f_permutation__U4680  ( .A1(_f_permutation__n6185 ), .A2(
        _f_permutation__n6186 ), .ZN(_f_permutation__n4213 ) );
  NAND2_X2 _f_permutation__U4679  ( .A1(_f_permutation__round_out[1173]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6183 ) );
  NAND2_X2 _f_permutation__U4678  ( .A1(_f_permutation__n7207 ), .A2(out[109]), 
        .ZN(_f_permutation__n6184 ) );
  NAND2_X2 _f_permutation__U4677  ( .A1(_f_permutation__n6183 ), .A2(
        _f_permutation__n6184 ), .ZN(_f_permutation__n4214 ) );
  NAND2_X2 _f_permutation__U4676  ( .A1(_f_permutation__round_out[1172]), 
        .A2(_f_permutation__n7132 ), .ZN(_f_permutation__n6181 ) );
  NAND2_X2 _f_permutation__U4675  ( .A1(_f_permutation__n7207 ), .A2(out[108]), 
        .ZN(_f_permutation__n6182 ) );
  NAND2_X2 _f_permutation__U4674  ( .A1(_f_permutation__n6181 ), .A2(
        _f_permutation__n6182 ), .ZN(_f_permutation__n4215 ) );
  NAND2_X2 _f_permutation__U4673  ( .A1(_f_permutation__round_out[1171]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6179 ) );
  NAND2_X2 _f_permutation__U4672  ( .A1(_f_permutation__n7207 ), .A2(out[107]), 
        .ZN(_f_permutation__n6180 ) );
  NAND2_X2 _f_permutation__U4671  ( .A1(_f_permutation__n6179 ), .A2(
        _f_permutation__n6180 ), .ZN(_f_permutation__n4216 ) );
  NAND2_X2 _f_permutation__U4670  ( .A1(_f_permutation__round_out[1170]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6177 ) );
  NAND2_X2 _f_permutation__U4669  ( .A1(_f_permutation__n7208 ), .A2(out[106]), 
        .ZN(_f_permutation__n6178 ) );
  NAND2_X2 _f_permutation__U4668  ( .A1(_f_permutation__n6177 ), .A2(
        _f_permutation__n6178 ), .ZN(_f_permutation__n4217 ) );
  NAND2_X2 _f_permutation__U4667  ( .A1(_f_permutation__round_out[1169]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6175 ) );
  NAND2_X2 _f_permutation__U4666  ( .A1(_f_permutation__n7208 ), .A2(out[105]), 
        .ZN(_f_permutation__n6176 ) );
  NAND2_X2 _f_permutation__U4665  ( .A1(_f_permutation__n6175 ), .A2(
        _f_permutation__n6176 ), .ZN(_f_permutation__n4218 ) );
  NAND2_X2 _f_permutation__U4664  ( .A1(_f_permutation__round_out[1168]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6173 ) );
  NAND2_X2 _f_permutation__U4663  ( .A1(_f_permutation__n7208 ), .A2(out[104]), 
        .ZN(_f_permutation__n6174 ) );
  NAND2_X2 _f_permutation__U4662  ( .A1(_f_permutation__n6173 ), .A2(
        _f_permutation__n6174 ), .ZN(_f_permutation__n4219 ) );
  NAND2_X2 _f_permutation__U4661  ( .A1(_f_permutation__round_out[1167]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6171 ) );
  NAND2_X2 _f_permutation__U4660  ( .A1(_f_permutation__n7208 ), .A2(out[119]), 
        .ZN(_f_permutation__n6172 ) );
  NAND2_X2 _f_permutation__U4659  ( .A1(_f_permutation__n6171 ), .A2(
        _f_permutation__n6172 ), .ZN(_f_permutation__n4220 ) );
  NAND2_X2 _f_permutation__U4658  ( .A1(_f_permutation__round_out[1166]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6169 ) );
  NAND2_X2 _f_permutation__U4657  ( .A1(_f_permutation__n7208 ), .A2(out[118]), 
        .ZN(_f_permutation__n6170 ) );
  NAND2_X2 _f_permutation__U4656  ( .A1(_f_permutation__n6169 ), .A2(
        _f_permutation__n6170 ), .ZN(_f_permutation__n4221 ) );
  NAND2_X2 _f_permutation__U4655  ( .A1(_f_permutation__round_out[1165]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6167 ) );
  NAND2_X2 _f_permutation__U4654  ( .A1(_f_permutation__n7208 ), .A2(out[117]), 
        .ZN(_f_permutation__n6168 ) );
  NAND2_X2 _f_permutation__U4653  ( .A1(_f_permutation__n6167 ), .A2(
        _f_permutation__n6168 ), .ZN(_f_permutation__n4222 ) );
  NAND2_X2 _f_permutation__U4652  ( .A1(_f_permutation__round_out[1164]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6165 ) );
  NAND2_X2 _f_permutation__U4651  ( .A1(_f_permutation__n7208 ), .A2(out[116]), 
        .ZN(_f_permutation__n6166 ) );
  NAND2_X2 _f_permutation__U4650  ( .A1(_f_permutation__n6165 ), .A2(
        _f_permutation__n6166 ), .ZN(_f_permutation__n4223 ) );
  NAND2_X2 _f_permutation__U4649  ( .A1(_f_permutation__round_out[1163]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6163 ) );
  NAND2_X2 _f_permutation__U4648  ( .A1(_f_permutation__n7208 ), .A2(out[115]), 
        .ZN(_f_permutation__n6164 ) );
  NAND2_X2 _f_permutation__U4647  ( .A1(_f_permutation__n6163 ), .A2(
        _f_permutation__n6164 ), .ZN(_f_permutation__n4224 ) );
  NAND2_X2 _f_permutation__U4646  ( .A1(_f_permutation__round_out[1162]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6161 ) );
  NAND2_X2 _f_permutation__U4645  ( .A1(_f_permutation__n7208 ), .A2(out[114]), 
        .ZN(_f_permutation__n6162 ) );
  NAND2_X2 _f_permutation__U4644  ( .A1(_f_permutation__n6161 ), .A2(
        _f_permutation__n6162 ), .ZN(_f_permutation__n4225 ) );
  NAND2_X2 _f_permutation__U4643  ( .A1(_f_permutation__round_out[1161]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6159 ) );
  NAND2_X2 _f_permutation__U4642  ( .A1(_f_permutation__n7208 ), .A2(out[113]), 
        .ZN(_f_permutation__n6160 ) );
  NAND2_X2 _f_permutation__U4641  ( .A1(_f_permutation__n6159 ), .A2(
        _f_permutation__n6160 ), .ZN(_f_permutation__n4226 ) );
  NAND2_X2 _f_permutation__U4640  ( .A1(_f_permutation__round_out[1160]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6157 ) );
  NAND2_X2 _f_permutation__U4639  ( .A1(_f_permutation__n7208 ), .A2(out[112]), 
        .ZN(_f_permutation__n6158 ) );
  NAND2_X2 _f_permutation__U4638  ( .A1(_f_permutation__n6157 ), .A2(
        _f_permutation__n6158 ), .ZN(_f_permutation__n4227 ) );
  NAND2_X2 _f_permutation__U4637  ( .A1(_f_permutation__round_out[1159]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6155 ) );
  NAND2_X2 _f_permutation__U4636  ( .A1(_f_permutation__n7209 ), .A2(out[127]), 
        .ZN(_f_permutation__n6156 ) );
  NAND2_X2 _f_permutation__U4635  ( .A1(_f_permutation__n6155 ), .A2(
        _f_permutation__n6156 ), .ZN(_f_permutation__n4228 ) );
  NAND2_X2 _f_permutation__U4634  ( .A1(_f_permutation__round_out[1158]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6153 ) );
  NAND2_X2 _f_permutation__U4633  ( .A1(_f_permutation__n7209 ), .A2(out[126]), 
        .ZN(_f_permutation__n6154 ) );
  NAND2_X2 _f_permutation__U4632  ( .A1(_f_permutation__n6153 ), .A2(
        _f_permutation__n6154 ), .ZN(_f_permutation__n4229 ) );
  NAND2_X2 _f_permutation__U4631  ( .A1(_f_permutation__round_out[1157]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6151 ) );
  NAND2_X2 _f_permutation__U4630  ( .A1(_f_permutation__n7209 ), .A2(out[125]), 
        .ZN(_f_permutation__n6152 ) );
  NAND2_X2 _f_permutation__U4629  ( .A1(_f_permutation__n6151 ), .A2(
        _f_permutation__n6152 ), .ZN(_f_permutation__n4230 ) );
  NAND2_X2 _f_permutation__U4628  ( .A1(_f_permutation__round_out[1156]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6149 ) );
  NAND2_X2 _f_permutation__U4627  ( .A1(_f_permutation__n7209 ), .A2(out[124]), 
        .ZN(_f_permutation__n6150 ) );
  NAND2_X2 _f_permutation__U4626  ( .A1(_f_permutation__n6149 ), .A2(
        _f_permutation__n6150 ), .ZN(_f_permutation__n4231 ) );
  NAND2_X2 _f_permutation__U4625  ( .A1(_f_permutation__round_out[1155]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6147 ) );
  NAND2_X2 _f_permutation__U4624  ( .A1(_f_permutation__n7209 ), .A2(out[123]), 
        .ZN(_f_permutation__n6148 ) );
  NAND2_X2 _f_permutation__U4623  ( .A1(_f_permutation__n6147 ), .A2(
        _f_permutation__n6148 ), .ZN(_f_permutation__n4232 ) );
  NAND2_X2 _f_permutation__U4622  ( .A1(_f_permutation__round_out[1154]), 
        .A2(_f_permutation__n7131 ), .ZN(_f_permutation__n6145 ) );
  NAND2_X2 _f_permutation__U4621  ( .A1(_f_permutation__n7209 ), .A2(out[122]), 
        .ZN(_f_permutation__n6146 ) );
  NAND2_X2 _f_permutation__U4620  ( .A1(_f_permutation__n6145 ), .A2(
        _f_permutation__n6146 ), .ZN(_f_permutation__n4233 ) );
  NAND2_X2 _f_permutation__U4619  ( .A1(_f_permutation__round_out[1153]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6143 ) );
  NAND2_X2 _f_permutation__U4618  ( .A1(_f_permutation__n7209 ), .A2(out[121]), 
        .ZN(_f_permutation__n6144 ) );
  NAND2_X2 _f_permutation__U4617  ( .A1(_f_permutation__n6143 ), .A2(
        _f_permutation__n6144 ), .ZN(_f_permutation__n4234 ) );
  NAND2_X2 _f_permutation__U4616  ( .A1(_f_permutation__round_out[1152]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6141 ) );
  NAND2_X2 _f_permutation__U4615  ( .A1(_f_permutation__n7209 ), .A2(out[120]), 
        .ZN(_f_permutation__n6142 ) );
  NAND2_X2 _f_permutation__U4614  ( .A1(_f_permutation__n6141 ), .A2(
        _f_permutation__n6142 ), .ZN(_f_permutation__n4235 ) );
  NAND2_X2 _f_permutation__U4613  ( .A1(_f_permutation__round_out[1151]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6139 ) );
  NAND2_X2 _f_permutation__U4612  ( .A1(_f_permutation__n7209 ), .A2(out[7]), 
        .ZN(_f_permutation__n6140 ) );
  NAND2_X2 _f_permutation__U4611  ( .A1(_f_permutation__n6139 ), .A2(
        _f_permutation__n6140 ), .ZN(_f_permutation__n4236 ) );
  NAND2_X2 _f_permutation__U4610  ( .A1(_f_permutation__round_out[1150]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6137 ) );
  NAND2_X2 _f_permutation__U4609  ( .A1(_f_permutation__n7209 ), .A2(out[6]), 
        .ZN(_f_permutation__n6138 ) );
  NAND2_X2 _f_permutation__U4608  ( .A1(_f_permutation__n6137 ), .A2(
        _f_permutation__n6138 ), .ZN(_f_permutation__n4237 ) );
  NAND2_X2 _f_permutation__U4607  ( .A1(_f_permutation__round_out[1149]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6135 ) );
  NAND2_X2 _f_permutation__U4606  ( .A1(_f_permutation__n7209 ), .A2(out[5]), 
        .ZN(_f_permutation__n6136 ) );
  NAND2_X2 _f_permutation__U4605  ( .A1(_f_permutation__n6135 ), .A2(
        _f_permutation__n6136 ), .ZN(_f_permutation__n4238 ) );
  NAND2_X2 _f_permutation__U4604  ( .A1(_f_permutation__round_out[1148]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6133 ) );
  NAND2_X2 _f_permutation__U4603  ( .A1(_f_permutation__n7210 ), .A2(out[4]), 
        .ZN(_f_permutation__n6134 ) );
  NAND2_X2 _f_permutation__U4602  ( .A1(_f_permutation__n6133 ), .A2(
        _f_permutation__n6134 ), .ZN(_f_permutation__n4239 ) );
  NAND2_X2 _f_permutation__U4601  ( .A1(_f_permutation__round_out[1147]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6131 ) );
  NAND2_X2 _f_permutation__U4600  ( .A1(_f_permutation__n7210 ), .A2(out[3]), 
        .ZN(_f_permutation__n6132 ) );
  NAND2_X2 _f_permutation__U4599  ( .A1(_f_permutation__n6131 ), .A2(
        _f_permutation__n6132 ), .ZN(_f_permutation__n4240 ) );
  NAND2_X2 _f_permutation__U4598  ( .A1(_f_permutation__round_out[1146]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6129 ) );
  NAND2_X2 _f_permutation__U4597  ( .A1(_f_permutation__n7210 ), .A2(out[2]), 
        .ZN(_f_permutation__n6130 ) );
  NAND2_X2 _f_permutation__U4596  ( .A1(_f_permutation__n6129 ), .A2(
        _f_permutation__n6130 ), .ZN(_f_permutation__n4241 ) );
  NAND2_X2 _f_permutation__U4595  ( .A1(_f_permutation__round_out[1145]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6127 ) );
  NAND2_X2 _f_permutation__U4594  ( .A1(_f_permutation__n7210 ), .A2(out[1]), 
        .ZN(_f_permutation__n6128 ) );
  NAND2_X2 _f_permutation__U4593  ( .A1(_f_permutation__n6127 ), .A2(
        _f_permutation__n6128 ), .ZN(_f_permutation__n4242 ) );
  NAND2_X2 _f_permutation__U4592  ( .A1(_f_permutation__round_out[1144]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6125 ) );
  NAND2_X2 _f_permutation__U4591  ( .A1(_f_permutation__n7210 ), .A2(out[0]), 
        .ZN(_f_permutation__n6126 ) );
  NAND2_X2 _f_permutation__U4590  ( .A1(_f_permutation__n6125 ), .A2(
        _f_permutation__n6126 ), .ZN(_f_permutation__n4243 ) );
  NAND2_X2 _f_permutation__U4589  ( .A1(_f_permutation__round_out[1143]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6123 ) );
  NAND2_X2 _f_permutation__U4588  ( .A1(_f_permutation__n7210 ), .A2(out[15]), 
        .ZN(_f_permutation__n6124 ) );
  NAND2_X2 _f_permutation__U4587  ( .A1(_f_permutation__n6123 ), .A2(
        _f_permutation__n6124 ), .ZN(_f_permutation__n4244 ) );
  NAND2_X2 _f_permutation__U4586  ( .A1(_f_permutation__round_out[1142]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6121 ) );
  NAND2_X2 _f_permutation__U4585  ( .A1(_f_permutation__n7210 ), .A2(out[14]), 
        .ZN(_f_permutation__n6122 ) );
  NAND2_X2 _f_permutation__U4584  ( .A1(_f_permutation__n6121 ), .A2(
        _f_permutation__n6122 ), .ZN(_f_permutation__n4245 ) );
  NAND2_X2 _f_permutation__U4583  ( .A1(_f_permutation__round_out[1141]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6119 ) );
  NAND2_X2 _f_permutation__U4582  ( .A1(_f_permutation__n7210 ), .A2(out[13]), 
        .ZN(_f_permutation__n6120 ) );
  NAND2_X2 _f_permutation__U4581  ( .A1(_f_permutation__n6119 ), .A2(
        _f_permutation__n6120 ), .ZN(_f_permutation__n4246 ) );
  NAND2_X2 _f_permutation__U4580  ( .A1(_f_permutation__round_out[1140]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6117 ) );
  NAND2_X2 _f_permutation__U4579  ( .A1(_f_permutation__n7210 ), .A2(out[12]), 
        .ZN(_f_permutation__n6118 ) );
  NAND2_X2 _f_permutation__U4578  ( .A1(_f_permutation__n6117 ), .A2(
        _f_permutation__n6118 ), .ZN(_f_permutation__n4247 ) );
  NAND2_X2 _f_permutation__U4577  ( .A1(_f_permutation__round_out[1139]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6115 ) );
  NAND2_X2 _f_permutation__U4576  ( .A1(_f_permutation__n7210 ), .A2(out[11]), 
        .ZN(_f_permutation__n6116 ) );
  NAND2_X2 _f_permutation__U4575  ( .A1(_f_permutation__n6115 ), .A2(
        _f_permutation__n6116 ), .ZN(_f_permutation__n4248 ) );
  NAND2_X2 _f_permutation__U4574  ( .A1(_f_permutation__round_out[1138]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6113 ) );
  NAND2_X2 _f_permutation__U4573  ( .A1(_f_permutation__n7210 ), .A2(out[10]), 
        .ZN(_f_permutation__n6114 ) );
  NAND2_X2 _f_permutation__U4572  ( .A1(_f_permutation__n6113 ), .A2(
        _f_permutation__n6114 ), .ZN(_f_permutation__n4249 ) );
  NAND2_X2 _f_permutation__U4571  ( .A1(_f_permutation__round_out[1137]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6111 ) );
  NAND2_X2 _f_permutation__U4570  ( .A1(_f_permutation__n7211 ), .A2(out[9]), 
        .ZN(_f_permutation__n6112 ) );
  NAND2_X2 _f_permutation__U4569  ( .A1(_f_permutation__n6111 ), .A2(
        _f_permutation__n6112 ), .ZN(_f_permutation__n4250 ) );
  NAND2_X2 _f_permutation__U4568  ( .A1(_f_permutation__round_out[1136]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6109 ) );
  NAND2_X2 _f_permutation__U4567  ( .A1(_f_permutation__n7211 ), .A2(out[8]), 
        .ZN(_f_permutation__n6110 ) );
  NAND2_X2 _f_permutation__U4566  ( .A1(_f_permutation__n6109 ), .A2(
        _f_permutation__n6110 ), .ZN(_f_permutation__n4251 ) );
  NAND2_X2 _f_permutation__U4565  ( .A1(_f_permutation__round_out[1135]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6107 ) );
  NAND2_X2 _f_permutation__U4564  ( .A1(_f_permutation__n7211 ), .A2(out[23]), 
        .ZN(_f_permutation__n6108 ) );
  NAND2_X2 _f_permutation__U4563  ( .A1(_f_permutation__n6107 ), .A2(
        _f_permutation__n6108 ), .ZN(_f_permutation__n4252 ) );
  NAND2_X2 _f_permutation__U4562  ( .A1(_f_permutation__round_out[1134]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6105 ) );
  NAND2_X2 _f_permutation__U4561  ( .A1(_f_permutation__n7211 ), .A2(out[22]), 
        .ZN(_f_permutation__n6106 ) );
  NAND2_X2 _f_permutation__U4560  ( .A1(_f_permutation__n6105 ), .A2(
        _f_permutation__n6106 ), .ZN(_f_permutation__n4253 ) );
  NAND2_X2 _f_permutation__U4559  ( .A1(_f_permutation__round_out[1133]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6103 ) );
  NAND2_X2 _f_permutation__U4558  ( .A1(_f_permutation__n7211 ), .A2(out[21]), 
        .ZN(_f_permutation__n6104 ) );
  NAND2_X2 _f_permutation__U4557  ( .A1(_f_permutation__n6103 ), .A2(
        _f_permutation__n6104 ), .ZN(_f_permutation__n4254 ) );
  NAND2_X2 _f_permutation__U4556  ( .A1(_f_permutation__round_out[1132]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6101 ) );
  NAND2_X2 _f_permutation__U4555  ( .A1(_f_permutation__n7211 ), .A2(out[20]), 
        .ZN(_f_permutation__n6102 ) );
  NAND2_X2 _f_permutation__U4554  ( .A1(_f_permutation__n6101 ), .A2(
        _f_permutation__n6102 ), .ZN(_f_permutation__n4255 ) );
  NAND2_X2 _f_permutation__U4553  ( .A1(_f_permutation__round_out[1131]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6099 ) );
  NAND2_X2 _f_permutation__U4552  ( .A1(_f_permutation__n7211 ), .A2(out[19]), 
        .ZN(_f_permutation__n6100 ) );
  NAND2_X2 _f_permutation__U4551  ( .A1(_f_permutation__n6099 ), .A2(
        _f_permutation__n6100 ), .ZN(_f_permutation__n4256 ) );
  NAND2_X2 _f_permutation__U4550  ( .A1(_f_permutation__round_out[1130]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6097 ) );
  NAND2_X2 _f_permutation__U4549  ( .A1(_f_permutation__n7211 ), .A2(out[18]), 
        .ZN(_f_permutation__n6098 ) );
  NAND2_X2 _f_permutation__U4548  ( .A1(_f_permutation__n6097 ), .A2(
        _f_permutation__n6098 ), .ZN(_f_permutation__n4257 ) );
  NAND2_X2 _f_permutation__U4547  ( .A1(_f_permutation__round_out[1129]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6095 ) );
  NAND2_X2 _f_permutation__U4546  ( .A1(_f_permutation__n7211 ), .A2(out[17]), 
        .ZN(_f_permutation__n6096 ) );
  NAND2_X2 _f_permutation__U4545  ( .A1(_f_permutation__n6095 ), .A2(
        _f_permutation__n6096 ), .ZN(_f_permutation__n4258 ) );
  NAND2_X2 _f_permutation__U4544  ( .A1(_f_permutation__round_out[1128]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6093 ) );
  NAND2_X2 _f_permutation__U4543  ( .A1(_f_permutation__n7211 ), .A2(out[16]), 
        .ZN(_f_permutation__n6094 ) );
  NAND2_X2 _f_permutation__U4542  ( .A1(_f_permutation__n6093 ), .A2(
        _f_permutation__n6094 ), .ZN(_f_permutation__n4259 ) );
  NAND2_X2 _f_permutation__U4541  ( .A1(_f_permutation__round_out[1127]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6091 ) );
  NAND2_X2 _f_permutation__U4540  ( .A1(_f_permutation__n7211 ), .A2(out[31]), 
        .ZN(_f_permutation__n6092 ) );
  NAND2_X2 _f_permutation__U4539  ( .A1(_f_permutation__n6091 ), .A2(
        _f_permutation__n6092 ), .ZN(_f_permutation__n4260 ) );
  NAND2_X2 _f_permutation__U4538  ( .A1(_f_permutation__round_out[1126]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6089 ) );
  NAND2_X2 _f_permutation__U4537  ( .A1(_f_permutation__n7212 ), .A2(out[30]), 
        .ZN(_f_permutation__n6090 ) );
  NAND2_X2 _f_permutation__U4536  ( .A1(_f_permutation__n6089 ), .A2(
        _f_permutation__n6090 ), .ZN(_f_permutation__n4261 ) );
  NAND2_X2 _f_permutation__U4535  ( .A1(_f_permutation__round_out[1125]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6087 ) );
  NAND2_X2 _f_permutation__U4534  ( .A1(_f_permutation__n7212 ), .A2(out[29]), 
        .ZN(_f_permutation__n6088 ) );
  NAND2_X2 _f_permutation__U4533  ( .A1(_f_permutation__n6087 ), .A2(
        _f_permutation__n6088 ), .ZN(_f_permutation__n4262 ) );
  NAND2_X2 _f_permutation__U4532  ( .A1(_f_permutation__round_out[1124]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6085 ) );
  NAND2_X2 _f_permutation__U4531  ( .A1(_f_permutation__n7212 ), .A2(out[28]), 
        .ZN(_f_permutation__n6086 ) );
  NAND2_X2 _f_permutation__U4530  ( .A1(_f_permutation__n6085 ), .A2(
        _f_permutation__n6086 ), .ZN(_f_permutation__n4263 ) );
  NAND2_X2 _f_permutation__U4529  ( .A1(_f_permutation__round_out[1123]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6083 ) );
  NAND2_X2 _f_permutation__U4528  ( .A1(_f_permutation__n7212 ), .A2(out[27]), 
        .ZN(_f_permutation__n6084 ) );
  NAND2_X2 _f_permutation__U4527  ( .A1(_f_permutation__n6083 ), .A2(
        _f_permutation__n6084 ), .ZN(_f_permutation__n4264 ) );
  NAND2_X2 _f_permutation__U4526  ( .A1(_f_permutation__round_out[1122]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6081 ) );
  NAND2_X2 _f_permutation__U4525  ( .A1(_f_permutation__n7212 ), .A2(out[26]), 
        .ZN(_f_permutation__n6082 ) );
  NAND2_X2 _f_permutation__U4524  ( .A1(_f_permutation__n6081 ), .A2(
        _f_permutation__n6082 ), .ZN(_f_permutation__n4265 ) );
  NAND2_X2 _f_permutation__U4523  ( .A1(_f_permutation__round_out[1121]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6079 ) );
  NAND2_X2 _f_permutation__U4522  ( .A1(_f_permutation__n7212 ), .A2(out[25]), 
        .ZN(_f_permutation__n6080 ) );
  NAND2_X2 _f_permutation__U4521  ( .A1(_f_permutation__n6079 ), .A2(
        _f_permutation__n6080 ), .ZN(_f_permutation__n4266 ) );
  NAND2_X2 _f_permutation__U4520  ( .A1(_f_permutation__round_out[1120]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6077 ) );
  NAND2_X2 _f_permutation__U4519  ( .A1(_f_permutation__n7212 ), .A2(out[24]), 
        .ZN(_f_permutation__n6078 ) );
  NAND2_X2 _f_permutation__U4518  ( .A1(_f_permutation__n6077 ), .A2(
        _f_permutation__n6078 ), .ZN(_f_permutation__n4267 ) );
  NAND2_X2 _f_permutation__U4517  ( .A1(_f_permutation__round_out[1119]), 
        .A2(_f_permutation__n7129 ), .ZN(_f_permutation__n6075 ) );
  NAND2_X2 _f_permutation__U4516  ( .A1(_f_permutation__n7212 ), .A2(out[39]), 
        .ZN(_f_permutation__n6076 ) );
  NAND2_X2 _f_permutation__U4515  ( .A1(_f_permutation__n6075 ), .A2(
        _f_permutation__n6076 ), .ZN(_f_permutation__n4268 ) );
  NAND2_X2 _f_permutation__U4514  ( .A1(_f_permutation__round_out[1118]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6073 ) );
  NAND2_X2 _f_permutation__U4513  ( .A1(_f_permutation__n7212 ), .A2(out[38]), 
        .ZN(_f_permutation__n6074 ) );
  NAND2_X2 _f_permutation__U4512  ( .A1(_f_permutation__n6073 ), .A2(
        _f_permutation__n6074 ), .ZN(_f_permutation__n4269 ) );
  NAND2_X2 _f_permutation__U4511  ( .A1(_f_permutation__round_out[1117]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6071 ) );
  NAND2_X2 _f_permutation__U4510  ( .A1(_f_permutation__n7212 ), .A2(out[37]), 
        .ZN(_f_permutation__n6072 ) );
  NAND2_X2 _f_permutation__U4509  ( .A1(_f_permutation__n6071 ), .A2(
        _f_permutation__n6072 ), .ZN(_f_permutation__n4270 ) );
  NAND2_X2 _f_permutation__U4508  ( .A1(_f_permutation__round_out[1116]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6069 ) );
  NAND2_X2 _f_permutation__U4507  ( .A1(_f_permutation__n7212 ), .A2(out[36]), 
        .ZN(_f_permutation__n6070 ) );
  NAND2_X2 _f_permutation__U4506  ( .A1(_f_permutation__n6069 ), .A2(
        _f_permutation__n6070 ), .ZN(_f_permutation__n4271 ) );
  NAND2_X2 _f_permutation__U4505  ( .A1(_f_permutation__round_out[1115]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6067 ) );
  NAND2_X2 _f_permutation__U4504  ( .A1(_f_permutation__n7213 ), .A2(out[35]), 
        .ZN(_f_permutation__n6068 ) );
  NAND2_X2 _f_permutation__U4503  ( .A1(_f_permutation__n6067 ), .A2(
        _f_permutation__n6068 ), .ZN(_f_permutation__n4272 ) );
  NAND2_X2 _f_permutation__U4502  ( .A1(_f_permutation__round_out[1114]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6065 ) );
  NAND2_X2 _f_permutation__U4501  ( .A1(_f_permutation__n7213 ), .A2(out[34]), 
        .ZN(_f_permutation__n6066 ) );
  NAND2_X2 _f_permutation__U4500  ( .A1(_f_permutation__n6065 ), .A2(
        _f_permutation__n6066 ), .ZN(_f_permutation__n4273 ) );
  NAND2_X2 _f_permutation__U4499  ( .A1(_f_permutation__round_out[1113]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6063 ) );
  NAND2_X2 _f_permutation__U4498  ( .A1(_f_permutation__n7213 ), .A2(out[33]), 
        .ZN(_f_permutation__n6064 ) );
  NAND2_X2 _f_permutation__U4497  ( .A1(_f_permutation__n6063 ), .A2(
        _f_permutation__n6064 ), .ZN(_f_permutation__n4274 ) );
  NAND2_X2 _f_permutation__U4496  ( .A1(_f_permutation__round_out[1112]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6061 ) );
  NAND2_X2 _f_permutation__U4495  ( .A1(_f_permutation__n7213 ), .A2(out[32]), 
        .ZN(_f_permutation__n6062 ) );
  NAND2_X2 _f_permutation__U4494  ( .A1(_f_permutation__n6061 ), .A2(
        _f_permutation__n6062 ), .ZN(_f_permutation__n4275 ) );
  NAND2_X2 _f_permutation__U4493  ( .A1(_f_permutation__round_out[1111]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6059 ) );
  NAND2_X2 _f_permutation__U4492  ( .A1(_f_permutation__n7213 ), .A2(out[47]), 
        .ZN(_f_permutation__n6060 ) );
  NAND2_X2 _f_permutation__U4491  ( .A1(_f_permutation__n6059 ), .A2(
        _f_permutation__n6060 ), .ZN(_f_permutation__n4276 ) );
  NAND2_X2 _f_permutation__U4490  ( .A1(_f_permutation__round_out[1110]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6057 ) );
  NAND2_X2 _f_permutation__U4489  ( .A1(_f_permutation__n7213 ), .A2(out[46]), 
        .ZN(_f_permutation__n6058 ) );
  NAND2_X2 _f_permutation__U4488  ( .A1(_f_permutation__n6057 ), .A2(
        _f_permutation__n6058 ), .ZN(_f_permutation__n4277 ) );
  NAND2_X2 _f_permutation__U4487  ( .A1(_f_permutation__round_out[1109]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6055 ) );
  NAND2_X2 _f_permutation__U4486  ( .A1(_f_permutation__n7213 ), .A2(out[45]), 
        .ZN(_f_permutation__n6056 ) );
  NAND2_X2 _f_permutation__U4485  ( .A1(_f_permutation__n6055 ), .A2(
        _f_permutation__n6056 ), .ZN(_f_permutation__n4278 ) );
  NAND2_X2 _f_permutation__U4484  ( .A1(_f_permutation__round_out[1108]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6053 ) );
  NAND2_X2 _f_permutation__U4483  ( .A1(_f_permutation__n7213 ), .A2(out[44]), 
        .ZN(_f_permutation__n6054 ) );
  NAND2_X2 _f_permutation__U4482  ( .A1(_f_permutation__n6053 ), .A2(
        _f_permutation__n6054 ), .ZN(_f_permutation__n4279 ) );
  NAND2_X2 _f_permutation__U4481  ( .A1(_f_permutation__round_out[1107]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6051 ) );
  NAND2_X2 _f_permutation__U4480  ( .A1(_f_permutation__n7213 ), .A2(out[43]), 
        .ZN(_f_permutation__n6052 ) );
  NAND2_X2 _f_permutation__U4479  ( .A1(_f_permutation__n6051 ), .A2(
        _f_permutation__n6052 ), .ZN(_f_permutation__n4280 ) );
  NAND2_X2 _f_permutation__U4478  ( .A1(_f_permutation__round_out[1106]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6049 ) );
  NAND2_X2 _f_permutation__U4477  ( .A1(_f_permutation__n7213 ), .A2(out[42]), 
        .ZN(_f_permutation__n6050 ) );
  NAND2_X2 _f_permutation__U4476  ( .A1(_f_permutation__n6049 ), .A2(
        _f_permutation__n6050 ), .ZN(_f_permutation__n4281 ) );
  NAND2_X2 _f_permutation__U4475  ( .A1(_f_permutation__round_out[1105]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6047 ) );
  NAND2_X2 _f_permutation__U4474  ( .A1(_f_permutation__n7213 ), .A2(out[41]), 
        .ZN(_f_permutation__n6048 ) );
  NAND2_X2 _f_permutation__U4473  ( .A1(_f_permutation__n6047 ), .A2(
        _f_permutation__n6048 ), .ZN(_f_permutation__n4282 ) );
  NAND2_X2 _f_permutation__U4472  ( .A1(_f_permutation__round_out[1104]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6045 ) );
  NAND2_X2 _f_permutation__U4471  ( .A1(_f_permutation__n7214 ), .A2(out[40]), 
        .ZN(_f_permutation__n6046 ) );
  NAND2_X2 _f_permutation__U4470  ( .A1(_f_permutation__n6045 ), .A2(
        _f_permutation__n6046 ), .ZN(_f_permutation__n4283 ) );
  NAND2_X2 _f_permutation__U4469  ( .A1(_f_permutation__round_out[1103]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6043 ) );
  NAND2_X2 _f_permutation__U4468  ( .A1(_f_permutation__n7214 ), .A2(out[55]), 
        .ZN(_f_permutation__n6044 ) );
  NAND2_X2 _f_permutation__U4467  ( .A1(_f_permutation__n6043 ), .A2(
        _f_permutation__n6044 ), .ZN(_f_permutation__n4284 ) );
  NAND2_X2 _f_permutation__U4466  ( .A1(_f_permutation__round_out[1102]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6041 ) );
  NAND2_X2 _f_permutation__U4465  ( .A1(_f_permutation__n7214 ), .A2(out[54]), 
        .ZN(_f_permutation__n6042 ) );
  NAND2_X2 _f_permutation__U4464  ( .A1(_f_permutation__n6041 ), .A2(
        _f_permutation__n6042 ), .ZN(_f_permutation__n4285 ) );
  NAND2_X2 _f_permutation__U4463  ( .A1(_f_permutation__round_out[1101]), 
        .A2(_f_permutation__n7128 ), .ZN(_f_permutation__n6039 ) );
  NAND2_X2 _f_permutation__U4462  ( .A1(_f_permutation__n7214 ), .A2(out[53]), 
        .ZN(_f_permutation__n6040 ) );
  NAND2_X2 _f_permutation__U4461  ( .A1(_f_permutation__n6039 ), .A2(
        _f_permutation__n6040 ), .ZN(_f_permutation__n4286 ) );
  NAND2_X2 _f_permutation__U4460  ( .A1(_f_permutation__round_out[1100]), 
        .A2(_f_permutation__n7127 ), .ZN(_f_permutation__n6037 ) );
  NAND2_X2 _f_permutation__U4459  ( .A1(_f_permutation__n7214 ), .A2(out[52]), 
        .ZN(_f_permutation__n6038 ) );
  NAND2_X2 _f_permutation__U4458  ( .A1(_f_permutation__n6037 ), .A2(
        _f_permutation__n6038 ), .ZN(_f_permutation__n4287 ) );
  NAND2_X2 _f_permutation__U4457  ( .A1(_f_permutation__round_out[1099]), 
        .A2(_f_permutation__n7130 ), .ZN(_f_permutation__n6035 ) );
  NAND2_X2 _f_permutation__U4456  ( .A1(_f_permutation__n7214 ), .A2(out[51]), 
        .ZN(_f_permutation__n6036 ) );
  NAND2_X2 _f_permutation__U4455  ( .A1(_f_permutation__n6035 ), .A2(
        _f_permutation__n6036 ), .ZN(_f_permutation__n4288 ) );
  NAND2_X2 _f_permutation__U4454  ( .A1(_f_permutation__round_out[1098]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6033 ) );
  NAND2_X2 _f_permutation__U4453  ( .A1(_f_permutation__n7214 ), .A2(out[50]), 
        .ZN(_f_permutation__n6034 ) );
  NAND2_X2 _f_permutation__U4452  ( .A1(_f_permutation__n6033 ), .A2(
        _f_permutation__n6034 ), .ZN(_f_permutation__n4289 ) );
  NAND2_X2 _f_permutation__U4451  ( .A1(_f_permutation__round_out[1097]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6031 ) );
  NAND2_X2 _f_permutation__U4450  ( .A1(_f_permutation__n7214 ), .A2(out[49]), 
        .ZN(_f_permutation__n6032 ) );
  NAND2_X2 _f_permutation__U4449  ( .A1(_f_permutation__n6031 ), .A2(
        _f_permutation__n6032 ), .ZN(_f_permutation__n4290 ) );
  NAND2_X2 _f_permutation__U4448  ( .A1(_f_permutation__round_out[1096]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6029 ) );
  NAND2_X2 _f_permutation__U4447  ( .A1(_f_permutation__n7214 ), .A2(out[48]), 
        .ZN(_f_permutation__n6030 ) );
  NAND2_X2 _f_permutation__U4446  ( .A1(_f_permutation__n6029 ), .A2(
        _f_permutation__n6030 ), .ZN(_f_permutation__n4291 ) );
  NAND2_X2 _f_permutation__U4445  ( .A1(_f_permutation__round_out[1095]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6027 ) );
  NAND2_X2 _f_permutation__U4444  ( .A1(_f_permutation__n7214 ), .A2(out[63]), 
        .ZN(_f_permutation__n6028 ) );
  NAND2_X2 _f_permutation__U4443  ( .A1(_f_permutation__n6027 ), .A2(
        _f_permutation__n6028 ), .ZN(_f_permutation__n4292 ) );
  NAND2_X2 _f_permutation__U4442  ( .A1(_f_permutation__round_out[1094]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6025 ) );
  NAND2_X2 _f_permutation__U4441  ( .A1(_f_permutation__n7214 ), .A2(out[62]), 
        .ZN(_f_permutation__n6026 ) );
  NAND2_X2 _f_permutation__U4440  ( .A1(_f_permutation__n6025 ), .A2(
        _f_permutation__n6026 ), .ZN(_f_permutation__n4293 ) );
  NAND2_X2 _f_permutation__U4439  ( .A1(_f_permutation__round_out[1093]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6023 ) );
  NAND2_X2 _f_permutation__U4438  ( .A1(_f_permutation__n7215 ), .A2(out[61]), 
        .ZN(_f_permutation__n6024 ) );
  NAND2_X2 _f_permutation__U4437  ( .A1(_f_permutation__n6023 ), .A2(
        _f_permutation__n6024 ), .ZN(_f_permutation__n4294 ) );
  NAND2_X2 _f_permutation__U4436  ( .A1(_f_permutation__round_out[1092]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6021 ) );
  NAND2_X2 _f_permutation__U4435  ( .A1(_f_permutation__n7215 ), .A2(out[60]), 
        .ZN(_f_permutation__n6022 ) );
  NAND2_X2 _f_permutation__U4434  ( .A1(_f_permutation__n6021 ), .A2(
        _f_permutation__n6022 ), .ZN(_f_permutation__n4295 ) );
  NAND2_X2 _f_permutation__U4433  ( .A1(_f_permutation__round_out[1091]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6019 ) );
  NAND2_X2 _f_permutation__U4432  ( .A1(_f_permutation__n7215 ), .A2(out[59]), 
        .ZN(_f_permutation__n6020 ) );
  NAND2_X2 _f_permutation__U4431  ( .A1(_f_permutation__n6019 ), .A2(
        _f_permutation__n6020 ), .ZN(_f_permutation__n4296 ) );
  NAND2_X2 _f_permutation__U4430  ( .A1(_f_permutation__round_out[1090]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6017 ) );
  NAND2_X2 _f_permutation__U4429  ( .A1(_f_permutation__n7215 ), .A2(out[58]), 
        .ZN(_f_permutation__n6018 ) );
  NAND2_X2 _f_permutation__U4428  ( .A1(_f_permutation__n6017 ), .A2(
        _f_permutation__n6018 ), .ZN(_f_permutation__n4297 ) );
  NAND2_X2 _f_permutation__U4427  ( .A1(_f_permutation__round_out[1089]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6015 ) );
  NAND2_X2 _f_permutation__U4426  ( .A1(_f_permutation__n7215 ), .A2(out[57]), 
        .ZN(_f_permutation__n6016 ) );
  NAND2_X2 _f_permutation__U4425  ( .A1(_f_permutation__n6015 ), .A2(
        _f_permutation__n6016 ), .ZN(_f_permutation__n4298 ) );
  NAND2_X2 _f_permutation__U4424  ( .A1(_f_permutation__round_out[1088]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6013 ) );
  NAND2_X2 _f_permutation__U4423  ( .A1(_f_permutation__n7215 ), .A2(out[56]), 
        .ZN(_f_permutation__n6014 ) );
  NAND2_X2 _f_permutation__U4422  ( .A1(_f_permutation__n6013 ), .A2(
        _f_permutation__n6014 ), .ZN(_f_permutation__n4299 ) );
  NAND2_X2 _f_permutation__U4421  ( .A1(_f_permutation__round_out[1087]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6011 ) );
  NAND2_X2 _f_permutation__U4420  ( .A1(_f_permutation__n7215 ), .A2(
        SYNOPSYS_UNCONNECTED_1), .ZN(_f_permutation__n6012 ) );
  NAND2_X2 _f_permutation__U4419  ( .A1(_f_permutation__n6011 ), .A2(
        _f_permutation__n6012 ), .ZN(_f_permutation__n4300 ) );
  NAND2_X2 _f_permutation__U4418  ( .A1(_f_permutation__round_out[1086]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6009 ) );
  NAND2_X2 _f_permutation__U4417  ( .A1(_f_permutation__n7215 ), .A2(
        SYNOPSYS_UNCONNECTED_2), .ZN(_f_permutation__n6010 ) );
  NAND2_X2 _f_permutation__U4416  ( .A1(_f_permutation__n6009 ), .A2(
        _f_permutation__n6010 ), .ZN(_f_permutation__n4301 ) );
  NAND2_X2 _f_permutation__U4415  ( .A1(_f_permutation__round_out[1085]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6007 ) );
  NAND2_X2 _f_permutation__U4414  ( .A1(_f_permutation__n7215 ), .A2(
        SYNOPSYS_UNCONNECTED_3), .ZN(_f_permutation__n6008 ) );
  NAND2_X2 _f_permutation__U4413  ( .A1(_f_permutation__n6007 ), .A2(
        _f_permutation__n6008 ), .ZN(_f_permutation__n4302 ) );
  NAND2_X2 _f_permutation__U4412  ( .A1(_f_permutation__round_out[1084]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6005 ) );
  NAND2_X2 _f_permutation__U4411  ( .A1(_f_permutation__n7215 ), .A2(
        SYNOPSYS_UNCONNECTED_4), .ZN(_f_permutation__n6006 ) );
  NAND2_X2 _f_permutation__U4410  ( .A1(_f_permutation__n6005 ), .A2(
        _f_permutation__n6006 ), .ZN(_f_permutation__n4303 ) );
  NAND2_X2 _f_permutation__U4409  ( .A1(_f_permutation__round_out[1083]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6003 ) );
  NAND2_X2 _f_permutation__U4408  ( .A1(_f_permutation__n7215 ), .A2(
        SYNOPSYS_UNCONNECTED_5), .ZN(_f_permutation__n6004 ) );
  NAND2_X2 _f_permutation__U4407  ( .A1(_f_permutation__n6003 ), .A2(
        _f_permutation__n6004 ), .ZN(_f_permutation__n4304 ) );
  NAND2_X2 _f_permutation__U4406  ( .A1(_f_permutation__round_out[1082]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n6001 ) );
  NAND2_X2 _f_permutation__U4405  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_6), .ZN(_f_permutation__n6002 ) );
  NAND2_X2 _f_permutation__U4404  ( .A1(_f_permutation__n6001 ), .A2(
        _f_permutation__n6002 ), .ZN(_f_permutation__n4305 ) );
  NAND2_X2 _f_permutation__U4403  ( .A1(_f_permutation__round_out[1081]), 
        .A2(_f_permutation__n7138 ), .ZN(_f_permutation__n5999 ) );
  NAND2_X2 _f_permutation__U4402  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_7), .ZN(_f_permutation__n6000 ) );
  NAND2_X2 _f_permutation__U4401  ( .A1(_f_permutation__n5999 ), .A2(
        _f_permutation__n6000 ), .ZN(_f_permutation__n4306 ) );
  NAND2_X2 _f_permutation__U4400  ( .A1(_f_permutation__round_out[1080]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5997 ) );
  NAND2_X2 _f_permutation__U4399  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_8), .ZN(_f_permutation__n5998 ) );
  NAND2_X2 _f_permutation__U4398  ( .A1(_f_permutation__n5997 ), .A2(
        _f_permutation__n5998 ), .ZN(_f_permutation__n4307 ) );
  NAND2_X2 _f_permutation__U4397  ( .A1(_f_permutation__round_out[1079]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5995 ) );
  NAND2_X2 _f_permutation__U4396  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_9), .ZN(_f_permutation__n5996 ) );
  NAND2_X2 _f_permutation__U4395  ( .A1(_f_permutation__n5995 ), .A2(
        _f_permutation__n5996 ), .ZN(_f_permutation__n4308 ) );
  NAND2_X2 _f_permutation__U4394  ( .A1(_f_permutation__round_out[1078]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5993 ) );
  NAND2_X2 _f_permutation__U4393  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_10), .ZN(_f_permutation__n5994 ) );
  NAND2_X2 _f_permutation__U4392  ( .A1(_f_permutation__n5993 ), .A2(
        _f_permutation__n5994 ), .ZN(_f_permutation__n4309 ) );
  NAND2_X2 _f_permutation__U4391  ( .A1(_f_permutation__round_out[1077]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5991 ) );
  NAND2_X2 _f_permutation__U4390  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_11), .ZN(_f_permutation__n5992 ) );
  NAND2_X2 _f_permutation__U4389  ( .A1(_f_permutation__n5991 ), .A2(
        _f_permutation__n5992 ), .ZN(_f_permutation__n4310 ) );
  NAND2_X2 _f_permutation__U4388  ( .A1(_f_permutation__round_out[1076]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5989 ) );
  NAND2_X2 _f_permutation__U4387  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_12), .ZN(_f_permutation__n5990 ) );
  NAND2_X2 _f_permutation__U4386  ( .A1(_f_permutation__n5989 ), .A2(
        _f_permutation__n5990 ), .ZN(_f_permutation__n4311 ) );
  NAND2_X2 _f_permutation__U4385  ( .A1(_f_permutation__round_out[1075]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5987 ) );
  NAND2_X2 _f_permutation__U4384  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_13), .ZN(_f_permutation__n5988 ) );
  NAND2_X2 _f_permutation__U4383  ( .A1(_f_permutation__n5987 ), .A2(
        _f_permutation__n5988 ), .ZN(_f_permutation__n4312 ) );
  NAND2_X2 _f_permutation__U4382  ( .A1(_f_permutation__round_out[1074]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5985 ) );
  NAND2_X2 _f_permutation__U4381  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_14), .ZN(_f_permutation__n5986 ) );
  NAND2_X2 _f_permutation__U4380  ( .A1(_f_permutation__n5985 ), .A2(
        _f_permutation__n5986 ), .ZN(_f_permutation__n4313 ) );
  NAND2_X2 _f_permutation__U4379  ( .A1(_f_permutation__round_out[1073]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5983 ) );
  NAND2_X2 _f_permutation__U4378  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_15), .ZN(_f_permutation__n5984 ) );
  NAND2_X2 _f_permutation__U4377  ( .A1(_f_permutation__n5983 ), .A2(
        _f_permutation__n5984 ), .ZN(_f_permutation__n4314 ) );
  NAND2_X2 _f_permutation__U4376  ( .A1(_f_permutation__round_out[1072]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5981 ) );
  NAND2_X2 _f_permutation__U4375  ( .A1(_f_permutation__n7216 ), .A2(
        SYNOPSYS_UNCONNECTED_16), .ZN(_f_permutation__n5982 ) );
  NAND2_X2 _f_permutation__U4374  ( .A1(_f_permutation__n5981 ), .A2(
        _f_permutation__n5982 ), .ZN(_f_permutation__n4315 ) );
  NAND2_X2 _f_permutation__U4373  ( .A1(_f_permutation__round_out[1071]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5979 ) );
  NAND2_X2 _f_permutation__U4372  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_17), .ZN(_f_permutation__n5980 ) );
  NAND2_X2 _f_permutation__U4371  ( .A1(_f_permutation__n5979 ), .A2(
        _f_permutation__n5980 ), .ZN(_f_permutation__n4316 ) );
  NAND2_X2 _f_permutation__U4370  ( .A1(_f_permutation__round_out[1070]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5977 ) );
  NAND2_X2 _f_permutation__U4369  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_18), .ZN(_f_permutation__n5978 ) );
  NAND2_X2 _f_permutation__U4368  ( .A1(_f_permutation__n5977 ), .A2(
        _f_permutation__n5978 ), .ZN(_f_permutation__n4317 ) );
  NAND2_X2 _f_permutation__U4367  ( .A1(_f_permutation__round_out[1069]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5975 ) );
  NAND2_X2 _f_permutation__U4366  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_19), .ZN(_f_permutation__n5976 ) );
  NAND2_X2 _f_permutation__U4365  ( .A1(_f_permutation__n5975 ), .A2(
        _f_permutation__n5976 ), .ZN(_f_permutation__n4318 ) );
  NAND2_X2 _f_permutation__U4364  ( .A1(_f_permutation__round_out[1068]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5973 ) );
  NAND2_X2 _f_permutation__U4363  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_20), .ZN(_f_permutation__n5974 ) );
  NAND2_X2 _f_permutation__U4362  ( .A1(_f_permutation__n5973 ), .A2(
        _f_permutation__n5974 ), .ZN(_f_permutation__n4319 ) );
  NAND2_X2 _f_permutation__U4361  ( .A1(_f_permutation__round_out[1067]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5971 ) );
  NAND2_X2 _f_permutation__U4360  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_21), .ZN(_f_permutation__n5972 ) );
  NAND2_X2 _f_permutation__U4359  ( .A1(_f_permutation__n5971 ), .A2(
        _f_permutation__n5972 ), .ZN(_f_permutation__n4320 ) );
  NAND2_X2 _f_permutation__U4358  ( .A1(_f_permutation__round_out[1066]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5969 ) );
  NAND2_X2 _f_permutation__U4357  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_22), .ZN(_f_permutation__n5970 ) );
  NAND2_X2 _f_permutation__U4356  ( .A1(_f_permutation__n5969 ), .A2(
        _f_permutation__n5970 ), .ZN(_f_permutation__n4321 ) );
  NAND2_X2 _f_permutation__U4355  ( .A1(_f_permutation__round_out[1065]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5967 ) );
  NAND2_X2 _f_permutation__U4354  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_23), .ZN(_f_permutation__n5968 ) );
  NAND2_X2 _f_permutation__U4353  ( .A1(_f_permutation__n5967 ), .A2(
        _f_permutation__n5968 ), .ZN(_f_permutation__n4322 ) );
  NAND2_X2 _f_permutation__U4352  ( .A1(_f_permutation__round_out[1064]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5965 ) );
  NAND2_X2 _f_permutation__U4351  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_24), .ZN(_f_permutation__n5966 ) );
  NAND2_X2 _f_permutation__U4350  ( .A1(_f_permutation__n5965 ), .A2(
        _f_permutation__n5966 ), .ZN(_f_permutation__n4323 ) );
  NAND2_X2 _f_permutation__U4349  ( .A1(_f_permutation__round_out[1063]), 
        .A2(_f_permutation__n7137 ), .ZN(_f_permutation__n5963 ) );
  NAND2_X2 _f_permutation__U4348  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_25), .ZN(_f_permutation__n5964 ) );
  NAND2_X2 _f_permutation__U4347  ( .A1(_f_permutation__n5963 ), .A2(
        _f_permutation__n5964 ), .ZN(_f_permutation__n4324 ) );
  NAND2_X2 _f_permutation__U4346  ( .A1(_f_permutation__round_out[1062]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5961 ) );
  NAND2_X2 _f_permutation__U4345  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_26), .ZN(_f_permutation__n5962 ) );
  NAND2_X2 _f_permutation__U4344  ( .A1(_f_permutation__n5961 ), .A2(
        _f_permutation__n5962 ), .ZN(_f_permutation__n4325 ) );
  NAND2_X2 _f_permutation__U4343  ( .A1(_f_permutation__round_out[1061]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5959 ) );
  NAND2_X2 _f_permutation__U4342  ( .A1(_f_permutation__n7217 ), .A2(
        SYNOPSYS_UNCONNECTED_27), .ZN(_f_permutation__n5960 ) );
  NAND2_X2 _f_permutation__U4341  ( .A1(_f_permutation__n5959 ), .A2(
        _f_permutation__n5960 ), .ZN(_f_permutation__n4326 ) );
  NAND2_X2 _f_permutation__U4340  ( .A1(_f_permutation__round_out[1060]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5957 ) );
  NAND2_X2 _f_permutation__U4339  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_28), .ZN(_f_permutation__n5958 ) );
  NAND2_X2 _f_permutation__U4338  ( .A1(_f_permutation__n5957 ), .A2(
        _f_permutation__n5958 ), .ZN(_f_permutation__n4327 ) );
  NAND2_X2 _f_permutation__U4337  ( .A1(_f_permutation__round_out[1059]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5955 ) );
  NAND2_X2 _f_permutation__U4336  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_29), .ZN(_f_permutation__n5956 ) );
  NAND2_X2 _f_permutation__U4335  ( .A1(_f_permutation__n5955 ), .A2(
        _f_permutation__n5956 ), .ZN(_f_permutation__n4328 ) );
  NAND2_X2 _f_permutation__U4334  ( .A1(_f_permutation__round_out[1058]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5953 ) );
  NAND2_X2 _f_permutation__U4333  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_30), .ZN(_f_permutation__n5954 ) );
  NAND2_X2 _f_permutation__U4332  ( .A1(_f_permutation__n5953 ), .A2(
        _f_permutation__n5954 ), .ZN(_f_permutation__n4329 ) );
  NAND2_X2 _f_permutation__U4331  ( .A1(_f_permutation__round_out[1057]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5951 ) );
  NAND2_X2 _f_permutation__U4330  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_31), .ZN(_f_permutation__n5952 ) );
  NAND2_X2 _f_permutation__U4329  ( .A1(_f_permutation__n5951 ), .A2(
        _f_permutation__n5952 ), .ZN(_f_permutation__n4330 ) );
  NAND2_X2 _f_permutation__U4328  ( .A1(_f_permutation__round_out[1056]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5949 ) );
  NAND2_X2 _f_permutation__U4327  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_32), .ZN(_f_permutation__n5950 ) );
  NAND2_X2 _f_permutation__U4326  ( .A1(_f_permutation__n5949 ), .A2(
        _f_permutation__n5950 ), .ZN(_f_permutation__n4331 ) );
  NAND2_X2 _f_permutation__U4325  ( .A1(_f_permutation__round_out[1055]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5947 ) );
  NAND2_X2 _f_permutation__U4324  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_33), .ZN(_f_permutation__n5948 ) );
  NAND2_X2 _f_permutation__U4323  ( .A1(_f_permutation__n5947 ), .A2(
        _f_permutation__n5948 ), .ZN(_f_permutation__n4332 ) );
  NAND2_X2 _f_permutation__U4322  ( .A1(_f_permutation__round_out[1054]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5945 ) );
  NAND2_X2 _f_permutation__U4321  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_34), .ZN(_f_permutation__n5946 ) );
  NAND2_X2 _f_permutation__U4320  ( .A1(_f_permutation__n5945 ), .A2(
        _f_permutation__n5946 ), .ZN(_f_permutation__n4333 ) );
  NAND2_X2 _f_permutation__U4319  ( .A1(_f_permutation__round_out[1053]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5943 ) );
  NAND2_X2 _f_permutation__U4318  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_35), .ZN(_f_permutation__n5944 ) );
  NAND2_X2 _f_permutation__U4317  ( .A1(_f_permutation__n5943 ), .A2(
        _f_permutation__n5944 ), .ZN(_f_permutation__n4334 ) );
  NAND2_X2 _f_permutation__U4316  ( .A1(_f_permutation__round_out[1052]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5941 ) );
  NAND2_X2 _f_permutation__U4315  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_36), .ZN(_f_permutation__n5942 ) );
  NAND2_X2 _f_permutation__U4314  ( .A1(_f_permutation__n5941 ), .A2(
        _f_permutation__n5942 ), .ZN(_f_permutation__n4335 ) );
  NAND2_X2 _f_permutation__U4313  ( .A1(_f_permutation__round_out[1051]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5939 ) );
  NAND2_X2 _f_permutation__U4312  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_37), .ZN(_f_permutation__n5940 ) );
  NAND2_X2 _f_permutation__U4311  ( .A1(_f_permutation__n5939 ), .A2(
        _f_permutation__n5940 ), .ZN(_f_permutation__n4336 ) );
  NAND2_X2 _f_permutation__U4310  ( .A1(_f_permutation__round_out[1050]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5937 ) );
  NAND2_X2 _f_permutation__U4309  ( .A1(_f_permutation__n7218 ), .A2(
        SYNOPSYS_UNCONNECTED_38), .ZN(_f_permutation__n5938 ) );
  NAND2_X2 _f_permutation__U4308  ( .A1(_f_permutation__n5937 ), .A2(
        _f_permutation__n5938 ), .ZN(_f_permutation__n4337 ) );
  NAND2_X2 _f_permutation__U4307  ( .A1(_f_permutation__round_out[1049]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5935 ) );
  NAND2_X2 _f_permutation__U4306  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_39), .ZN(_f_permutation__n5936 ) );
  NAND2_X2 _f_permutation__U4305  ( .A1(_f_permutation__n5935 ), .A2(
        _f_permutation__n5936 ), .ZN(_f_permutation__n4338 ) );
  NAND2_X2 _f_permutation__U4304  ( .A1(_f_permutation__round_out[1048]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5933 ) );
  NAND2_X2 _f_permutation__U4303  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_40), .ZN(_f_permutation__n5934 ) );
  NAND2_X2 _f_permutation__U4302  ( .A1(_f_permutation__n5933 ), .A2(
        _f_permutation__n5934 ), .ZN(_f_permutation__n4339 ) );
  NAND2_X2 _f_permutation__U4301  ( .A1(_f_permutation__round_out[1047]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5931 ) );
  NAND2_X2 _f_permutation__U4300  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_41), .ZN(_f_permutation__n5932 ) );
  NAND2_X2 _f_permutation__U4299  ( .A1(_f_permutation__n5931 ), .A2(
        _f_permutation__n5932 ), .ZN(_f_permutation__n4340 ) );
  NAND2_X2 _f_permutation__U4298  ( .A1(_f_permutation__round_out[1046]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5929 ) );
  NAND2_X2 _f_permutation__U4297  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_42), .ZN(_f_permutation__n5930 ) );
  NAND2_X2 _f_permutation__U4296  ( .A1(_f_permutation__n5929 ), .A2(
        _f_permutation__n5930 ), .ZN(_f_permutation__n4341 ) );
  NAND2_X2 _f_permutation__U4295  ( .A1(_f_permutation__round_out[1045]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5927 ) );
  NAND2_X2 _f_permutation__U4294  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_43), .ZN(_f_permutation__n5928 ) );
  NAND2_X2 _f_permutation__U4293  ( .A1(_f_permutation__n5927 ), .A2(
        _f_permutation__n5928 ), .ZN(_f_permutation__n4342 ) );
  NAND2_X2 _f_permutation__U4292  ( .A1(_f_permutation__round_out[1044]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5925 ) );
  NAND2_X2 _f_permutation__U4291  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_44), .ZN(_f_permutation__n5926 ) );
  NAND2_X2 _f_permutation__U4290  ( .A1(_f_permutation__n5925 ), .A2(
        _f_permutation__n5926 ), .ZN(_f_permutation__n4343 ) );
  NAND2_X2 _f_permutation__U4289  ( .A1(_f_permutation__round_out[1043]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5923 ) );
  NAND2_X2 _f_permutation__U4288  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_45), .ZN(_f_permutation__n5924 ) );
  NAND2_X2 _f_permutation__U4287  ( .A1(_f_permutation__n5923 ), .A2(
        _f_permutation__n5924 ), .ZN(_f_permutation__n4344 ) );
  NAND2_X2 _f_permutation__U4286  ( .A1(_f_permutation__round_out[1042]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5921 ) );
  NAND2_X2 _f_permutation__U4285  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_46), .ZN(_f_permutation__n5922 ) );
  NAND2_X2 _f_permutation__U4284  ( .A1(_f_permutation__n5921 ), .A2(
        _f_permutation__n5922 ), .ZN(_f_permutation__n4345 ) );
  NAND2_X2 _f_permutation__U4283  ( .A1(_f_permutation__round_out[1041]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5919 ) );
  NAND2_X2 _f_permutation__U4282  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_47), .ZN(_f_permutation__n5920 ) );
  NAND2_X2 _f_permutation__U4281  ( .A1(_f_permutation__n5919 ), .A2(
        _f_permutation__n5920 ), .ZN(_f_permutation__n4346 ) );
  NAND2_X2 _f_permutation__U4280  ( .A1(_f_permutation__round_out[1040]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5917 ) );
  NAND2_X2 _f_permutation__U4279  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_48), .ZN(_f_permutation__n5918 ) );
  NAND2_X2 _f_permutation__U4278  ( .A1(_f_permutation__n5917 ), .A2(
        _f_permutation__n5918 ), .ZN(_f_permutation__n4347 ) );
  NAND2_X2 _f_permutation__U4277  ( .A1(_f_permutation__round_out[1039]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5915 ) );
  NAND2_X2 _f_permutation__U4276  ( .A1(_f_permutation__n7219 ), .A2(
        SYNOPSYS_UNCONNECTED_49), .ZN(_f_permutation__n5916 ) );
  NAND2_X2 _f_permutation__U4275  ( .A1(_f_permutation__n5915 ), .A2(
        _f_permutation__n5916 ), .ZN(_f_permutation__n4348 ) );
  NAND2_X2 _f_permutation__U4274  ( .A1(_f_permutation__round_out[1038]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5913 ) );
  NAND2_X2 _f_permutation__U4273  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_50), .ZN(_f_permutation__n5914 ) );
  NAND2_X2 _f_permutation__U4272  ( .A1(_f_permutation__n5913 ), .A2(
        _f_permutation__n5914 ), .ZN(_f_permutation__n4349 ) );
  NAND2_X2 _f_permutation__U4271  ( .A1(_f_permutation__round_out[1037]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5911 ) );
  NAND2_X2 _f_permutation__U4270  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_51), .ZN(_f_permutation__n5912 ) );
  NAND2_X2 _f_permutation__U4269  ( .A1(_f_permutation__n5911 ), .A2(
        _f_permutation__n5912 ), .ZN(_f_permutation__n4350 ) );
  NAND2_X2 _f_permutation__U4268  ( .A1(_f_permutation__round_out[1036]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5909 ) );
  NAND2_X2 _f_permutation__U4267  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_52), .ZN(_f_permutation__n5910 ) );
  NAND2_X2 _f_permutation__U4266  ( .A1(_f_permutation__n5909 ), .A2(
        _f_permutation__n5910 ), .ZN(_f_permutation__n4351 ) );
  NAND2_X2 _f_permutation__U4265  ( .A1(_f_permutation__round_out[1035]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5907 ) );
  NAND2_X2 _f_permutation__U4264  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_53), .ZN(_f_permutation__n5908 ) );
  NAND2_X2 _f_permutation__U4263  ( .A1(_f_permutation__n5907 ), .A2(
        _f_permutation__n5908 ), .ZN(_f_permutation__n4352 ) );
  NAND2_X2 _f_permutation__U4262  ( .A1(_f_permutation__round_out[1034]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5905 ) );
  NAND2_X2 _f_permutation__U4261  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_54), .ZN(_f_permutation__n5906 ) );
  NAND2_X2 _f_permutation__U4260  ( .A1(_f_permutation__n5905 ), .A2(
        _f_permutation__n5906 ), .ZN(_f_permutation__n4353 ) );
  NAND2_X2 _f_permutation__U4259  ( .A1(_f_permutation__round_out[1033]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5903 ) );
  NAND2_X2 _f_permutation__U4258  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_55), .ZN(_f_permutation__n5904 ) );
  NAND2_X2 _f_permutation__U4257  ( .A1(_f_permutation__n5903 ), .A2(
        _f_permutation__n5904 ), .ZN(_f_permutation__n4354 ) );
  NAND2_X2 _f_permutation__U4256  ( .A1(_f_permutation__round_out[1032]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5901 ) );
  NAND2_X2 _f_permutation__U4255  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_56), .ZN(_f_permutation__n5902 ) );
  NAND2_X2 _f_permutation__U4254  ( .A1(_f_permutation__n5901 ), .A2(
        _f_permutation__n5902 ), .ZN(_f_permutation__n4355 ) );
  NAND2_X2 _f_permutation__U4253  ( .A1(_f_permutation__round_out[1031]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5899 ) );
  NAND2_X2 _f_permutation__U4252  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_57), .ZN(_f_permutation__n5900 ) );
  NAND2_X2 _f_permutation__U4251  ( .A1(_f_permutation__n5899 ), .A2(
        _f_permutation__n5900 ), .ZN(_f_permutation__n4356 ) );
  NAND2_X2 _f_permutation__U4250  ( .A1(_f_permutation__round_out[1030]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5897 ) );
  NAND2_X2 _f_permutation__U4249  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_58), .ZN(_f_permutation__n5898 ) );
  NAND2_X2 _f_permutation__U4248  ( .A1(_f_permutation__n5897 ), .A2(
        _f_permutation__n5898 ), .ZN(_f_permutation__n4357 ) );
  NAND2_X2 _f_permutation__U4247  ( .A1(_f_permutation__round_out[1029]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5895 ) );
  NAND2_X2 _f_permutation__U4246  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_59), .ZN(_f_permutation__n5896 ) );
  NAND2_X2 _f_permutation__U4245  ( .A1(_f_permutation__n5895 ), .A2(
        _f_permutation__n5896 ), .ZN(_f_permutation__n4358 ) );
  NAND2_X2 _f_permutation__U4244  ( .A1(_f_permutation__round_out[1028]), 
        .A2(_f_permutation__n7135 ), .ZN(_f_permutation__n5893 ) );
  NAND2_X2 _f_permutation__U4243  ( .A1(_f_permutation__n7220 ), .A2(
        SYNOPSYS_UNCONNECTED_60), .ZN(_f_permutation__n5894 ) );
  NAND2_X2 _f_permutation__U4242  ( .A1(_f_permutation__n5893 ), .A2(
        _f_permutation__n5894 ), .ZN(_f_permutation__n4359 ) );
  NAND2_X2 _f_permutation__U4241  ( .A1(_f_permutation__round_out[1027]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5891 ) );
  NAND2_X2 _f_permutation__U4240  ( .A1(_f_permutation__n7231 ), .A2(
        SYNOPSYS_UNCONNECTED_61), .ZN(_f_permutation__n5892 ) );
  NAND2_X2 _f_permutation__U4239  ( .A1(_f_permutation__n5891 ), .A2(
        _f_permutation__n5892 ), .ZN(_f_permutation__n4360 ) );
  NAND2_X2 _f_permutation__U4238  ( .A1(_f_permutation__round_out[1026]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5889 ) );
  NAND2_X2 _f_permutation__U4237  ( .A1(_f_permutation__n7308 ), .A2(
        SYNOPSYS_UNCONNECTED_62), .ZN(_f_permutation__n5890 ) );
  NAND2_X2 _f_permutation__U4236  ( .A1(_f_permutation__n5889 ), .A2(
        _f_permutation__n5890 ), .ZN(_f_permutation__n4361 ) );
  NAND2_X2 _f_permutation__U4235  ( .A1(_f_permutation__round_out[1025]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5887 ) );
  NAND2_X2 _f_permutation__U4234  ( .A1(_f_permutation__n7214 ), .A2(
        SYNOPSYS_UNCONNECTED_63), .ZN(_f_permutation__n5888 ) );
  NAND2_X2 _f_permutation__U4233  ( .A1(_f_permutation__n5887 ), .A2(
        _f_permutation__n5888 ), .ZN(_f_permutation__n4362 ) );
  NAND2_X2 _f_permutation__U4232  ( .A1(_f_permutation__round_out[1024]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5885 ) );
  NAND2_X2 _f_permutation__U4231  ( .A1(_f_permutation__n7214 ), .A2(
        SYNOPSYS_UNCONNECTED_64), .ZN(_f_permutation__n5886 ) );
  NAND2_X2 _f_permutation__U4230  ( .A1(_f_permutation__n5885 ), .A2(
        _f_permutation__n5886 ), .ZN(_f_permutation__n4363 ) );
  NAND2_X2 _f_permutation__U4229  ( .A1(_f_permutation__round_out[1023]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5883 ) );
  NAND2_X2 _f_permutation__U4228  ( .A1(SYNOPSYS_UNCONNECTED_65), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n5884 ) );
  NAND2_X2 _f_permutation__U4227  ( .A1(_f_permutation__n5883 ), .A2(
        _f_permutation__n5884 ), .ZN(_f_permutation__n4364 ) );
  NAND2_X2 _f_permutation__U4226  ( .A1(_f_permutation__round_out[1022]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5881 ) );
  NAND2_X2 _f_permutation__U4225  ( .A1(SYNOPSYS_UNCONNECTED_66), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5882 ) );
  NAND2_X2 _f_permutation__U4224  ( .A1(_f_permutation__n5881 ), .A2(
        _f_permutation__n5882 ), .ZN(_f_permutation__n4365 ) );
  NAND2_X2 _f_permutation__U4223  ( .A1(_f_permutation__round_out[1021]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5879 ) );
  NAND2_X2 _f_permutation__U4222  ( .A1(SYNOPSYS_UNCONNECTED_67), .A2(
        _f_permutation__n7308 ), .ZN(_f_permutation__n5880 ) );
  NAND2_X2 _f_permutation__U4221  ( .A1(_f_permutation__n5879 ), .A2(
        _f_permutation__n5880 ), .ZN(_f_permutation__n4366 ) );
  NAND2_X2 _f_permutation__U4220  ( .A1(_f_permutation__round_out[1020]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5877 ) );
  NAND2_X2 _f_permutation__U4219  ( .A1(SYNOPSYS_UNCONNECTED_68), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n5878 ) );
  NAND2_X2 _f_permutation__U4218  ( .A1(_f_permutation__n5877 ), .A2(
        _f_permutation__n5878 ), .ZN(_f_permutation__n4367 ) );
  NAND2_X2 _f_permutation__U4217  ( .A1(_f_permutation__round_out[1019]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5875 ) );
  NAND2_X2 _f_permutation__U4216  ( .A1(SYNOPSYS_UNCONNECTED_69), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n5876 ) );
  NAND2_X2 _f_permutation__U4215  ( .A1(_f_permutation__n5875 ), .A2(
        _f_permutation__n5876 ), .ZN(_f_permutation__n4368 ) );
  NAND2_X2 _f_permutation__U4214  ( .A1(_f_permutation__round_out[1018]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5873 ) );
  NAND2_X2 _f_permutation__U4213  ( .A1(SYNOPSYS_UNCONNECTED_70), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n5874 ) );
  NAND2_X2 _f_permutation__U4212  ( .A1(_f_permutation__n5873 ), .A2(
        _f_permutation__n5874 ), .ZN(_f_permutation__n4369 ) );
  NAND2_X2 _f_permutation__U4211  ( .A1(_f_permutation__round_out[1017]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5871 ) );
  NAND2_X2 _f_permutation__U4210  ( .A1(SYNOPSYS_UNCONNECTED_71), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n5872 ) );
  NAND2_X2 _f_permutation__U4209  ( .A1(_f_permutation__n5871 ), .A2(
        _f_permutation__n5872 ), .ZN(_f_permutation__n4370 ) );
  NAND2_X2 _f_permutation__U4208  ( .A1(_f_permutation__round_out[1016]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5869 ) );
  NAND2_X2 _f_permutation__U4207  ( .A1(SYNOPSYS_UNCONNECTED_72), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5870 ) );
  NAND2_X2 _f_permutation__U4206  ( .A1(_f_permutation__n5869 ), .A2(
        _f_permutation__n5870 ), .ZN(_f_permutation__n4371 ) );
  NAND2_X2 _f_permutation__U4205  ( .A1(_f_permutation__round_out[1015]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5867 ) );
  NAND2_X2 _f_permutation__U4204  ( .A1(SYNOPSYS_UNCONNECTED_73), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5868 ) );
  NAND2_X2 _f_permutation__U4203  ( .A1(_f_permutation__n5867 ), .A2(
        _f_permutation__n5868 ), .ZN(_f_permutation__n4372 ) );
  NAND2_X2 _f_permutation__U4202  ( .A1(_f_permutation__round_out[1014]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5865 ) );
  NAND2_X2 _f_permutation__U4201  ( .A1(SYNOPSYS_UNCONNECTED_74), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5866 ) );
  NAND2_X2 _f_permutation__U4200  ( .A1(_f_permutation__n5865 ), .A2(
        _f_permutation__n5866 ), .ZN(_f_permutation__n4373 ) );
  NAND2_X2 _f_permutation__U4199  ( .A1(_f_permutation__round_out[1013]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5863 ) );
  NAND2_X2 _f_permutation__U4198  ( .A1(SYNOPSYS_UNCONNECTED_75), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5864 ) );
  NAND2_X2 _f_permutation__U4197  ( .A1(_f_permutation__n5863 ), .A2(
        _f_permutation__n5864 ), .ZN(_f_permutation__n4374 ) );
  NAND2_X2 _f_permutation__U4196  ( .A1(_f_permutation__round_out[1012]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5861 ) );
  NAND2_X2 _f_permutation__U4195  ( .A1(SYNOPSYS_UNCONNECTED_76), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5862 ) );
  NAND2_X2 _f_permutation__U4194  ( .A1(_f_permutation__n5861 ), .A2(
        _f_permutation__n5862 ), .ZN(_f_permutation__n4375 ) );
  NAND2_X2 _f_permutation__U4193  ( .A1(_f_permutation__round_out[1011]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5859 ) );
  NAND2_X2 _f_permutation__U4192  ( .A1(SYNOPSYS_UNCONNECTED_77), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5860 ) );
  NAND2_X2 _f_permutation__U4191  ( .A1(_f_permutation__n5859 ), .A2(
        _f_permutation__n5860 ), .ZN(_f_permutation__n4376 ) );
  NAND2_X2 _f_permutation__U4190  ( .A1(_f_permutation__round_out[1010]), 
        .A2(_f_permutation__n7134 ), .ZN(_f_permutation__n5857 ) );
  NAND2_X2 _f_permutation__U4189  ( .A1(SYNOPSYS_UNCONNECTED_78), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5858 ) );
  NAND2_X2 _f_permutation__U4188  ( .A1(_f_permutation__n5857 ), .A2(
        _f_permutation__n5858 ), .ZN(_f_permutation__n4377 ) );
  NAND2_X2 _f_permutation__U4187  ( .A1(_f_permutation__round_out[1009]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n5855 ) );
  NAND2_X2 _f_permutation__U4186  ( .A1(SYNOPSYS_UNCONNECTED_79), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5856 ) );
  NAND2_X2 _f_permutation__U4185  ( .A1(_f_permutation__n5855 ), .A2(
        _f_permutation__n5856 ), .ZN(_f_permutation__n4378 ) );
  NAND2_X2 _f_permutation__U4184  ( .A1(_f_permutation__round_out[1008]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n5853 ) );
  NAND2_X2 _f_permutation__U4183  ( .A1(SYNOPSYS_UNCONNECTED_80), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5854 ) );
  NAND2_X2 _f_permutation__U4182  ( .A1(_f_permutation__n5853 ), .A2(
        _f_permutation__n5854 ), .ZN(_f_permutation__n4379 ) );
  NAND2_X2 _f_permutation__U4181  ( .A1(_f_permutation__round_out[1007]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n5851 ) );
  NAND2_X2 _f_permutation__U4180  ( .A1(SYNOPSYS_UNCONNECTED_81), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5852 ) );
  NAND2_X2 _f_permutation__U4179  ( .A1(_f_permutation__n5851 ), .A2(
        _f_permutation__n5852 ), .ZN(_f_permutation__n4380 ) );
  NAND2_X2 _f_permutation__U4178  ( .A1(_f_permutation__round_out[1006]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n5849 ) );
  NAND2_X2 _f_permutation__U4177  ( .A1(SYNOPSYS_UNCONNECTED_82), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5850 ) );
  NAND2_X2 _f_permutation__U4176  ( .A1(_f_permutation__n5849 ), .A2(
        _f_permutation__n5850 ), .ZN(_f_permutation__n4381 ) );
  NAND2_X2 _f_permutation__U4175  ( .A1(_f_permutation__round_out[1005]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n5847 ) );
  NAND2_X2 _f_permutation__U4174  ( .A1(SYNOPSYS_UNCONNECTED_83), .A2(
        _f_permutation__n7221 ), .ZN(_f_permutation__n5848 ) );
  NAND2_X2 _f_permutation__U4173  ( .A1(_f_permutation__n5847 ), .A2(
        _f_permutation__n5848 ), .ZN(_f_permutation__n4382 ) );
  NAND2_X2 _f_permutation__U4172  ( .A1(_f_permutation__round_out[1004]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n5845 ) );
  NAND2_X2 _f_permutation__U4171  ( .A1(SYNOPSYS_UNCONNECTED_84), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5846 ) );
  NAND2_X2 _f_permutation__U4170  ( .A1(_f_permutation__n5845 ), .A2(
        _f_permutation__n5846 ), .ZN(_f_permutation__n4383 ) );
  NAND2_X2 _f_permutation__U4169  ( .A1(_f_permutation__round_out[1003]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n5843 ) );
  NAND2_X2 _f_permutation__U4168  ( .A1(SYNOPSYS_UNCONNECTED_85), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5844 ) );
  NAND2_X2 _f_permutation__U4167  ( .A1(_f_permutation__n5843 ), .A2(
        _f_permutation__n5844 ), .ZN(_f_permutation__n4384 ) );
  NAND2_X2 _f_permutation__U4166  ( .A1(_f_permutation__round_out[1002]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n5841 ) );
  NAND2_X2 _f_permutation__U4165  ( .A1(SYNOPSYS_UNCONNECTED_86), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5842 ) );
  NAND2_X2 _f_permutation__U4164  ( .A1(_f_permutation__n5841 ), .A2(
        _f_permutation__n5842 ), .ZN(_f_permutation__n4385 ) );
  NAND2_X2 _f_permutation__U4163  ( .A1(_f_permutation__round_out[1001]), 
        .A2(_f_permutation__n7133 ), .ZN(_f_permutation__n5839 ) );
  NAND2_X2 _f_permutation__U4162  ( .A1(SYNOPSYS_UNCONNECTED_87), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5840 ) );
  NAND2_X2 _f_permutation__U4161  ( .A1(_f_permutation__n5839 ), .A2(
        _f_permutation__n5840 ), .ZN(_f_permutation__n4386 ) );
  NAND2_X2 _f_permutation__U4160  ( .A1(_f_permutation__round_out[1000]), 
        .A2(_f_permutation__n7136 ), .ZN(_f_permutation__n5837 ) );
  NAND2_X2 _f_permutation__U4159  ( .A1(SYNOPSYS_UNCONNECTED_88), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5838 ) );
  NAND2_X2 _f_permutation__U4158  ( .A1(_f_permutation__n5837 ), .A2(
        _f_permutation__n5838 ), .ZN(_f_permutation__n4387 ) );
  NAND2_X2 _f_permutation__U4157  ( .A1(_f_permutation__round_out[999]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5835 ) );
  NAND2_X2 _f_permutation__U4156  ( .A1(SYNOPSYS_UNCONNECTED_89), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5836 ) );
  NAND2_X2 _f_permutation__U4155  ( .A1(_f_permutation__n5835 ), .A2(
        _f_permutation__n5836 ), .ZN(_f_permutation__n4388 ) );
  NAND2_X2 _f_permutation__U4154  ( .A1(_f_permutation__round_out[998]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5833 ) );
  NAND2_X2 _f_permutation__U4153  ( .A1(SYNOPSYS_UNCONNECTED_90), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5834 ) );
  NAND2_X2 _f_permutation__U4152  ( .A1(_f_permutation__n5833 ), .A2(
        _f_permutation__n5834 ), .ZN(_f_permutation__n4389 ) );
  NAND2_X2 _f_permutation__U4151  ( .A1(_f_permutation__round_out[997]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5831 ) );
  NAND2_X2 _f_permutation__U4150  ( .A1(SYNOPSYS_UNCONNECTED_91), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5832 ) );
  NAND2_X2 _f_permutation__U4149  ( .A1(_f_permutation__n5831 ), .A2(
        _f_permutation__n5832 ), .ZN(_f_permutation__n4390 ) );
  NAND2_X2 _f_permutation__U4148  ( .A1(_f_permutation__round_out[996]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5829 ) );
  NAND2_X2 _f_permutation__U4147  ( .A1(SYNOPSYS_UNCONNECTED_92), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5830 ) );
  NAND2_X2 _f_permutation__U4146  ( .A1(_f_permutation__n5829 ), .A2(
        _f_permutation__n5830 ), .ZN(_f_permutation__n4391 ) );
  NAND2_X2 _f_permutation__U4145  ( .A1(_f_permutation__round_out[995]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5827 ) );
  NAND2_X2 _f_permutation__U4144  ( .A1(SYNOPSYS_UNCONNECTED_93), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5828 ) );
  NAND2_X2 _f_permutation__U4143  ( .A1(_f_permutation__n5827 ), .A2(
        _f_permutation__n5828 ), .ZN(_f_permutation__n4392 ) );
  NAND2_X2 _f_permutation__U4142  ( .A1(_f_permutation__round_out[994]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5825 ) );
  NAND2_X2 _f_permutation__U4141  ( .A1(SYNOPSYS_UNCONNECTED_94), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5826 ) );
  NAND2_X2 _f_permutation__U4140  ( .A1(_f_permutation__n5825 ), .A2(
        _f_permutation__n5826 ), .ZN(_f_permutation__n4393 ) );
  NAND2_X2 _f_permutation__U4139  ( .A1(_f_permutation__round_out[993]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5823 ) );
  NAND2_X2 _f_permutation__U4138  ( .A1(SYNOPSYS_UNCONNECTED_95), .A2(
        _f_permutation__n7222 ), .ZN(_f_permutation__n5824 ) );
  NAND2_X2 _f_permutation__U4137  ( .A1(_f_permutation__n5823 ), .A2(
        _f_permutation__n5824 ), .ZN(_f_permutation__n4394 ) );
  NAND2_X2 _f_permutation__U4136  ( .A1(_f_permutation__round_out[992]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5821 ) );
  NAND2_X2 _f_permutation__U4135  ( .A1(SYNOPSYS_UNCONNECTED_96), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5822 ) );
  NAND2_X2 _f_permutation__U4134  ( .A1(_f_permutation__n5821 ), .A2(
        _f_permutation__n5822 ), .ZN(_f_permutation__n4395 ) );
  NAND2_X2 _f_permutation__U4133  ( .A1(_f_permutation__round_out[991]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5819 ) );
  NAND2_X2 _f_permutation__U4132  ( .A1(SYNOPSYS_UNCONNECTED_97), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5820 ) );
  NAND2_X2 _f_permutation__U4131  ( .A1(_f_permutation__n5819 ), .A2(
        _f_permutation__n5820 ), .ZN(_f_permutation__n4396 ) );
  NAND2_X2 _f_permutation__U4130  ( .A1(_f_permutation__round_out[990]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5817 ) );
  NAND2_X2 _f_permutation__U4129  ( .A1(SYNOPSYS_UNCONNECTED_98), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5818 ) );
  NAND2_X2 _f_permutation__U4128  ( .A1(_f_permutation__n5817 ), .A2(
        _f_permutation__n5818 ), .ZN(_f_permutation__n4397 ) );
  NAND2_X2 _f_permutation__U4127  ( .A1(_f_permutation__round_out[989]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5815 ) );
  NAND2_X2 _f_permutation__U4126  ( .A1(SYNOPSYS_UNCONNECTED_99), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5816 ) );
  NAND2_X2 _f_permutation__U4125  ( .A1(_f_permutation__n5815 ), .A2(
        _f_permutation__n5816 ), .ZN(_f_permutation__n4398 ) );
  NAND2_X2 _f_permutation__U4124  ( .A1(_f_permutation__round_out[988]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5813 ) );
  NAND2_X2 _f_permutation__U4123  ( .A1(SYNOPSYS_UNCONNECTED_100), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5814 ) );
  NAND2_X2 _f_permutation__U4122  ( .A1(_f_permutation__n5813 ), .A2(
        _f_permutation__n5814 ), .ZN(_f_permutation__n4399 ) );
  NAND2_X2 _f_permutation__U4121  ( .A1(_f_permutation__round_out[987]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5811 ) );
  NAND2_X2 _f_permutation__U4120  ( .A1(SYNOPSYS_UNCONNECTED_101), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5812 ) );
  NAND2_X2 _f_permutation__U4119  ( .A1(_f_permutation__n5811 ), .A2(
        _f_permutation__n5812 ), .ZN(_f_permutation__n4400 ) );
  NAND2_X2 _f_permutation__U4118  ( .A1(_f_permutation__round_out[986]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5809 ) );
  NAND2_X2 _f_permutation__U4117  ( .A1(SYNOPSYS_UNCONNECTED_102), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5810 ) );
  NAND2_X2 _f_permutation__U4116  ( .A1(_f_permutation__n5809 ), .A2(
        _f_permutation__n5810 ), .ZN(_f_permutation__n4401 ) );
  NAND2_X2 _f_permutation__U4115  ( .A1(_f_permutation__round_out[985]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5807 ) );
  NAND2_X2 _f_permutation__U4114  ( .A1(SYNOPSYS_UNCONNECTED_103), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5808 ) );
  NAND2_X2 _f_permutation__U4113  ( .A1(_f_permutation__n5807 ), .A2(
        _f_permutation__n5808 ), .ZN(_f_permutation__n4402 ) );
  NAND2_X2 _f_permutation__U4112  ( .A1(_f_permutation__round_out[984]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5781 ) );
  NAND2_X2 _f_permutation__U4111  ( .A1(SYNOPSYS_UNCONNECTED_104), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5806 ) );
  NAND2_X2 _f_permutation__U4110  ( .A1(_f_permutation__n5781 ), .A2(
        _f_permutation__n5806 ), .ZN(_f_permutation__n4403 ) );
  NAND2_X2 _f_permutation__U4109  ( .A1(_f_permutation__round_out[983]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5779 ) );
  NAND2_X2 _f_permutation__U4108  ( .A1(SYNOPSYS_UNCONNECTED_105), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5780 ) );
  NAND2_X2 _f_permutation__U4107  ( .A1(_f_permutation__n5779 ), .A2(
        _f_permutation__n5780 ), .ZN(_f_permutation__n4404 ) );
  NAND2_X2 _f_permutation__U4106  ( .A1(_f_permutation__round_out[982]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5777 ) );
  NAND2_X2 _f_permutation__U4105  ( .A1(SYNOPSYS_UNCONNECTED_106), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5778 ) );
  NAND2_X2 _f_permutation__U4104  ( .A1(_f_permutation__n5777 ), .A2(
        _f_permutation__n5778 ), .ZN(_f_permutation__n4405 ) );
  NAND2_X2 _f_permutation__U4103  ( .A1(_f_permutation__round_out[981]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5775 ) );
  NAND2_X2 _f_permutation__U4102  ( .A1(SYNOPSYS_UNCONNECTED_107), .A2(
        _f_permutation__n7223 ), .ZN(_f_permutation__n5776 ) );
  NAND2_X2 _f_permutation__U4101  ( .A1(_f_permutation__n5775 ), .A2(
        _f_permutation__n5776 ), .ZN(_f_permutation__n4406 ) );
  NAND2_X2 _f_permutation__U4100  ( .A1(_f_permutation__round_out[980]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5773 ) );
  NAND2_X2 _f_permutation__U4099  ( .A1(SYNOPSYS_UNCONNECTED_108), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5774 ) );
  NAND2_X2 _f_permutation__U4098  ( .A1(_f_permutation__n5773 ), .A2(
        _f_permutation__n5774 ), .ZN(_f_permutation__n4407 ) );
  NAND2_X2 _f_permutation__U4097  ( .A1(_f_permutation__round_out[979]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5771 ) );
  NAND2_X2 _f_permutation__U4096  ( .A1(SYNOPSYS_UNCONNECTED_109), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5772 ) );
  NAND2_X2 _f_permutation__U4095  ( .A1(_f_permutation__n5771 ), .A2(
        _f_permutation__n5772 ), .ZN(_f_permutation__n4408 ) );
  NAND2_X2 _f_permutation__U4094  ( .A1(_f_permutation__round_out[978]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5769 ) );
  NAND2_X2 _f_permutation__U4093  ( .A1(SYNOPSYS_UNCONNECTED_110), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5770 ) );
  NAND2_X2 _f_permutation__U4092  ( .A1(_f_permutation__n5769 ), .A2(
        _f_permutation__n5770 ), .ZN(_f_permutation__n4409 ) );
  NAND2_X2 _f_permutation__U4091  ( .A1(_f_permutation__round_out[977]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5767 ) );
  NAND2_X2 _f_permutation__U4090  ( .A1(SYNOPSYS_UNCONNECTED_111), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5768 ) );
  NAND2_X2 _f_permutation__U4089  ( .A1(_f_permutation__n5767 ), .A2(
        _f_permutation__n5768 ), .ZN(_f_permutation__n4410 ) );
  NAND2_X2 _f_permutation__U4088  ( .A1(_f_permutation__round_out[976]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5765 ) );
  NAND2_X2 _f_permutation__U4087  ( .A1(SYNOPSYS_UNCONNECTED_112), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5766 ) );
  NAND2_X2 _f_permutation__U4086  ( .A1(_f_permutation__n5765 ), .A2(
        _f_permutation__n5766 ), .ZN(_f_permutation__n4411 ) );
  NAND2_X2 _f_permutation__U4085  ( .A1(_f_permutation__round_out[975]), .A2(
        _f_permutation__n7121 ), .ZN(_f_permutation__n5763 ) );
  NAND2_X2 _f_permutation__U4084  ( .A1(SYNOPSYS_UNCONNECTED_113), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5764 ) );
  NAND2_X2 _f_permutation__U4083  ( .A1(_f_permutation__n5763 ), .A2(
        _f_permutation__n5764 ), .ZN(_f_permutation__n4412 ) );
  NAND2_X2 _f_permutation__U4082  ( .A1(_f_permutation__round_out[974]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5761 ) );
  NAND2_X2 _f_permutation__U4081  ( .A1(SYNOPSYS_UNCONNECTED_114), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5762 ) );
  NAND2_X2 _f_permutation__U4080  ( .A1(_f_permutation__n5761 ), .A2(
        _f_permutation__n5762 ), .ZN(_f_permutation__n4413 ) );
  NAND2_X2 _f_permutation__U4079  ( .A1(_f_permutation__round_out[973]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5759 ) );
  NAND2_X2 _f_permutation__U4078  ( .A1(SYNOPSYS_UNCONNECTED_115), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5760 ) );
  NAND2_X2 _f_permutation__U4077  ( .A1(_f_permutation__n5759 ), .A2(
        _f_permutation__n5760 ), .ZN(_f_permutation__n4414 ) );
  NAND2_X2 _f_permutation__U4076  ( .A1(_f_permutation__round_out[972]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5757 ) );
  NAND2_X2 _f_permutation__U4075  ( .A1(SYNOPSYS_UNCONNECTED_116), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5758 ) );
  NAND2_X2 _f_permutation__U4074  ( .A1(_f_permutation__n5757 ), .A2(
        _f_permutation__n5758 ), .ZN(_f_permutation__n4415 ) );
  NAND2_X2 _f_permutation__U4073  ( .A1(_f_permutation__round_out[971]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5755 ) );
  NAND2_X2 _f_permutation__U4072  ( .A1(SYNOPSYS_UNCONNECTED_117), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5756 ) );
  NAND2_X2 _f_permutation__U4071  ( .A1(_f_permutation__n5755 ), .A2(
        _f_permutation__n5756 ), .ZN(_f_permutation__n4416 ) );
  NAND2_X2 _f_permutation__U4070  ( .A1(_f_permutation__round_out[970]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5753 ) );
  NAND2_X2 _f_permutation__U4069  ( .A1(SYNOPSYS_UNCONNECTED_118), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5754 ) );
  NAND2_X2 _f_permutation__U4068  ( .A1(_f_permutation__n5753 ), .A2(
        _f_permutation__n5754 ), .ZN(_f_permutation__n4417 ) );
  NAND2_X2 _f_permutation__U4067  ( .A1(_f_permutation__round_out[969]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5751 ) );
  NAND2_X2 _f_permutation__U4066  ( .A1(SYNOPSYS_UNCONNECTED_119), .A2(
        _f_permutation__n7224 ), .ZN(_f_permutation__n5752 ) );
  NAND2_X2 _f_permutation__U4065  ( .A1(_f_permutation__n5751 ), .A2(
        _f_permutation__n5752 ), .ZN(_f_permutation__n4418 ) );
  NAND2_X2 _f_permutation__U4064  ( .A1(_f_permutation__round_out[968]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5749 ) );
  NAND2_X2 _f_permutation__U4063  ( .A1(SYNOPSYS_UNCONNECTED_120), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5750 ) );
  NAND2_X2 _f_permutation__U4062  ( .A1(_f_permutation__n5749 ), .A2(
        _f_permutation__n5750 ), .ZN(_f_permutation__n4419 ) );
  NAND2_X2 _f_permutation__U4061  ( .A1(_f_permutation__round_out[967]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5747 ) );
  NAND2_X2 _f_permutation__U4060  ( .A1(SYNOPSYS_UNCONNECTED_121), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5748 ) );
  NAND2_X2 _f_permutation__U4059  ( .A1(_f_permutation__n5747 ), .A2(
        _f_permutation__n5748 ), .ZN(_f_permutation__n4420 ) );
  NAND2_X2 _f_permutation__U4058  ( .A1(_f_permutation__round_out[966]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5745 ) );
  NAND2_X2 _f_permutation__U4057  ( .A1(SYNOPSYS_UNCONNECTED_122), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5746 ) );
  NAND2_X2 _f_permutation__U4056  ( .A1(_f_permutation__n5745 ), .A2(
        _f_permutation__n5746 ), .ZN(_f_permutation__n4421 ) );
  NAND2_X2 _f_permutation__U4055  ( .A1(_f_permutation__round_out[965]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5743 ) );
  NAND2_X2 _f_permutation__U4054  ( .A1(SYNOPSYS_UNCONNECTED_123), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5744 ) );
  NAND2_X2 _f_permutation__U4053  ( .A1(_f_permutation__n5743 ), .A2(
        _f_permutation__n5744 ), .ZN(_f_permutation__n4422 ) );
  NAND2_X2 _f_permutation__U4052  ( .A1(_f_permutation__round_out[964]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5741 ) );
  NAND2_X2 _f_permutation__U4051  ( .A1(SYNOPSYS_UNCONNECTED_124), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5742 ) );
  NAND2_X2 _f_permutation__U4050  ( .A1(_f_permutation__n5741 ), .A2(
        _f_permutation__n5742 ), .ZN(_f_permutation__n4423 ) );
  NAND2_X2 _f_permutation__U4049  ( .A1(_f_permutation__round_out[963]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5739 ) );
  NAND2_X2 _f_permutation__U4048  ( .A1(SYNOPSYS_UNCONNECTED_125), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5740 ) );
  NAND2_X2 _f_permutation__U4047  ( .A1(_f_permutation__n5739 ), .A2(
        _f_permutation__n5740 ), .ZN(_f_permutation__n4424 ) );
  NAND2_X2 _f_permutation__U4046  ( .A1(_f_permutation__round_out[962]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5737 ) );
  NAND2_X2 _f_permutation__U4045  ( .A1(SYNOPSYS_UNCONNECTED_126), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5738 ) );
  NAND2_X2 _f_permutation__U4044  ( .A1(_f_permutation__n5737 ), .A2(
        _f_permutation__n5738 ), .ZN(_f_permutation__n4425 ) );
  NAND2_X2 _f_permutation__U4043  ( .A1(_f_permutation__round_out[961]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5735 ) );
  NAND2_X2 _f_permutation__U4042  ( .A1(SYNOPSYS_UNCONNECTED_127), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5736 ) );
  NAND2_X2 _f_permutation__U4041  ( .A1(_f_permutation__n5735 ), .A2(
        _f_permutation__n5736 ), .ZN(_f_permutation__n4426 ) );
  NAND2_X2 _f_permutation__U4040  ( .A1(_f_permutation__round_out[960]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5733 ) );
  NAND2_X2 _f_permutation__U4039  ( .A1(SYNOPSYS_UNCONNECTED_128), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5734 ) );
  NAND2_X2 _f_permutation__U4038  ( .A1(_f_permutation__n5733 ), .A2(
        _f_permutation__n5734 ), .ZN(_f_permutation__n4427 ) );
  NAND2_X2 _f_permutation__U4037  ( .A1(_f_permutation__round_out[959]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5731 ) );
  NAND2_X2 _f_permutation__U4036  ( .A1(SYNOPSYS_UNCONNECTED_129), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5732 ) );
  NAND2_X2 _f_permutation__U4035  ( .A1(_f_permutation__n5731 ), .A2(
        _f_permutation__n5732 ), .ZN(_f_permutation__n4428 ) );
  NAND2_X2 _f_permutation__U4034  ( .A1(_f_permutation__round_out[958]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5729 ) );
  NAND2_X2 _f_permutation__U4033  ( .A1(SYNOPSYS_UNCONNECTED_130), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5730 ) );
  NAND2_X2 _f_permutation__U4032  ( .A1(_f_permutation__n5729 ), .A2(
        _f_permutation__n5730 ), .ZN(_f_permutation__n4429 ) );
  NAND2_X2 _f_permutation__U4031  ( .A1(_f_permutation__round_out[957]), .A2(
        _f_permutation__n7120 ), .ZN(_f_permutation__n5727 ) );
  NAND2_X2 _f_permutation__U4030  ( .A1(SYNOPSYS_UNCONNECTED_131), .A2(
        _f_permutation__n7225 ), .ZN(_f_permutation__n5728 ) );
  NAND2_X2 _f_permutation__U4029  ( .A1(_f_permutation__n5727 ), .A2(
        _f_permutation__n5728 ), .ZN(_f_permutation__n4430 ) );
  NAND2_X2 _f_permutation__U4028  ( .A1(_f_permutation__round_out[956]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5725 ) );
  NAND2_X2 _f_permutation__U4027  ( .A1(SYNOPSYS_UNCONNECTED_132), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5726 ) );
  NAND2_X2 _f_permutation__U4026  ( .A1(_f_permutation__n5725 ), .A2(
        _f_permutation__n5726 ), .ZN(_f_permutation__n4431 ) );
  NAND2_X2 _f_permutation__U4025  ( .A1(_f_permutation__round_out[955]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5723 ) );
  NAND2_X2 _f_permutation__U4024  ( .A1(SYNOPSYS_UNCONNECTED_133), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5724 ) );
  NAND2_X2 _f_permutation__U4023  ( .A1(_f_permutation__n5723 ), .A2(
        _f_permutation__n5724 ), .ZN(_f_permutation__n4432 ) );
  NAND2_X2 _f_permutation__U4022  ( .A1(_f_permutation__round_out[954]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5721 ) );
  NAND2_X2 _f_permutation__U4021  ( .A1(SYNOPSYS_UNCONNECTED_134), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5722 ) );
  NAND2_X2 _f_permutation__U4020  ( .A1(_f_permutation__n5721 ), .A2(
        _f_permutation__n5722 ), .ZN(_f_permutation__n4433 ) );
  NAND2_X2 _f_permutation__U4019  ( .A1(_f_permutation__round_out[953]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5719 ) );
  NAND2_X2 _f_permutation__U4018  ( .A1(SYNOPSYS_UNCONNECTED_135), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5720 ) );
  NAND2_X2 _f_permutation__U4017  ( .A1(_f_permutation__n5719 ), .A2(
        _f_permutation__n5720 ), .ZN(_f_permutation__n4434 ) );
  NAND2_X2 _f_permutation__U4016  ( .A1(_f_permutation__round_out[952]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5717 ) );
  NAND2_X2 _f_permutation__U4015  ( .A1(SYNOPSYS_UNCONNECTED_136), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5718 ) );
  NAND2_X2 _f_permutation__U4014  ( .A1(_f_permutation__n5717 ), .A2(
        _f_permutation__n5718 ), .ZN(_f_permutation__n4435 ) );
  NAND2_X2 _f_permutation__U4013  ( .A1(_f_permutation__round_out[951]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5715 ) );
  NAND2_X2 _f_permutation__U4012  ( .A1(SYNOPSYS_UNCONNECTED_137), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5716 ) );
  NAND2_X2 _f_permutation__U4011  ( .A1(_f_permutation__n5715 ), .A2(
        _f_permutation__n5716 ), .ZN(_f_permutation__n4436 ) );
  NAND2_X2 _f_permutation__U4010  ( .A1(_f_permutation__round_out[950]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5713 ) );
  NAND2_X2 _f_permutation__U4009  ( .A1(SYNOPSYS_UNCONNECTED_138), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5714 ) );
  NAND2_X2 _f_permutation__U4008  ( .A1(_f_permutation__n5713 ), .A2(
        _f_permutation__n5714 ), .ZN(_f_permutation__n4437 ) );
  NAND2_X2 _f_permutation__U4007  ( .A1(_f_permutation__round_out[949]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5711 ) );
  NAND2_X2 _f_permutation__U4006  ( .A1(SYNOPSYS_UNCONNECTED_139), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5712 ) );
  NAND2_X2 _f_permutation__U4005  ( .A1(_f_permutation__n5711 ), .A2(
        _f_permutation__n5712 ), .ZN(_f_permutation__n4438 ) );
  NAND2_X2 _f_permutation__U4004  ( .A1(_f_permutation__round_out[948]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5709 ) );
  NAND2_X2 _f_permutation__U4003  ( .A1(SYNOPSYS_UNCONNECTED_140), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5710 ) );
  NAND2_X2 _f_permutation__U4002  ( .A1(_f_permutation__n5709 ), .A2(
        _f_permutation__n5710 ), .ZN(_f_permutation__n4439 ) );
  NAND2_X2 _f_permutation__U4001  ( .A1(_f_permutation__round_out[947]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5707 ) );
  NAND2_X2 _f_permutation__U4000  ( .A1(SYNOPSYS_UNCONNECTED_141), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5708 ) );
  NAND2_X2 _f_permutation__U3999  ( .A1(_f_permutation__n5707 ), .A2(
        _f_permutation__n5708 ), .ZN(_f_permutation__n4440 ) );
  NAND2_X2 _f_permutation__U3998  ( .A1(_f_permutation__round_out[946]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5705 ) );
  NAND2_X2 _f_permutation__U3997  ( .A1(SYNOPSYS_UNCONNECTED_142), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5706 ) );
  NAND2_X2 _f_permutation__U3996  ( .A1(_f_permutation__n5705 ), .A2(
        _f_permutation__n5706 ), .ZN(_f_permutation__n4441 ) );
  NAND2_X2 _f_permutation__U3995  ( .A1(_f_permutation__round_out[945]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5703 ) );
  NAND2_X2 _f_permutation__U3994  ( .A1(SYNOPSYS_UNCONNECTED_143), .A2(
        _f_permutation__n7226 ), .ZN(_f_permutation__n5704 ) );
  NAND2_X2 _f_permutation__U3993  ( .A1(_f_permutation__n5703 ), .A2(
        _f_permutation__n5704 ), .ZN(_f_permutation__n4442 ) );
  NAND2_X2 _f_permutation__U3992  ( .A1(_f_permutation__round_out[944]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5701 ) );
  NAND2_X2 _f_permutation__U3991  ( .A1(SYNOPSYS_UNCONNECTED_144), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5702 ) );
  NAND2_X2 _f_permutation__U3990  ( .A1(_f_permutation__n5701 ), .A2(
        _f_permutation__n5702 ), .ZN(_f_permutation__n4443 ) );
  NAND2_X2 _f_permutation__U3989  ( .A1(_f_permutation__round_out[943]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5699 ) );
  NAND2_X2 _f_permutation__U3988  ( .A1(SYNOPSYS_UNCONNECTED_145), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5700 ) );
  NAND2_X2 _f_permutation__U3987  ( .A1(_f_permutation__n5699 ), .A2(
        _f_permutation__n5700 ), .ZN(_f_permutation__n4444 ) );
  NAND2_X2 _f_permutation__U3986  ( .A1(_f_permutation__round_out[942]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5697 ) );
  NAND2_X2 _f_permutation__U3985  ( .A1(SYNOPSYS_UNCONNECTED_146), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5698 ) );
  NAND2_X2 _f_permutation__U3984  ( .A1(_f_permutation__n5697 ), .A2(
        _f_permutation__n5698 ), .ZN(_f_permutation__n4445 ) );
  NAND2_X2 _f_permutation__U3983  ( .A1(_f_permutation__round_out[941]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5695 ) );
  NAND2_X2 _f_permutation__U3982  ( .A1(SYNOPSYS_UNCONNECTED_147), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5696 ) );
  NAND2_X2 _f_permutation__U3981  ( .A1(_f_permutation__n5695 ), .A2(
        _f_permutation__n5696 ), .ZN(_f_permutation__n4446 ) );
  NAND2_X2 _f_permutation__U3980  ( .A1(_f_permutation__round_out[940]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5693 ) );
  NAND2_X2 _f_permutation__U3979  ( .A1(SYNOPSYS_UNCONNECTED_148), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5694 ) );
  NAND2_X2 _f_permutation__U3978  ( .A1(_f_permutation__n5693 ), .A2(
        _f_permutation__n5694 ), .ZN(_f_permutation__n4447 ) );
  NAND2_X2 _f_permutation__U3977  ( .A1(_f_permutation__round_out[939]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5691 ) );
  NAND2_X2 _f_permutation__U3976  ( .A1(SYNOPSYS_UNCONNECTED_149), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5692 ) );
  NAND2_X2 _f_permutation__U3975  ( .A1(_f_permutation__n5691 ), .A2(
        _f_permutation__n5692 ), .ZN(_f_permutation__n4448 ) );
  NAND2_X2 _f_permutation__U3974  ( .A1(_f_permutation__round_out[938]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5689 ) );
  NAND2_X2 _f_permutation__U3973  ( .A1(SYNOPSYS_UNCONNECTED_150), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5690 ) );
  NAND2_X2 _f_permutation__U3972  ( .A1(_f_permutation__n5689 ), .A2(
        _f_permutation__n5690 ), .ZN(_f_permutation__n4449 ) );
  NAND2_X2 _f_permutation__U3971  ( .A1(_f_permutation__round_out[937]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5687 ) );
  NAND2_X2 _f_permutation__U3970  ( .A1(SYNOPSYS_UNCONNECTED_151), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5688 ) );
  NAND2_X2 _f_permutation__U3969  ( .A1(_f_permutation__n5687 ), .A2(
        _f_permutation__n5688 ), .ZN(_f_permutation__n4450 ) );
  NAND2_X2 _f_permutation__U3968  ( .A1(_f_permutation__round_out[936]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5685 ) );
  NAND2_X2 _f_permutation__U3967  ( .A1(SYNOPSYS_UNCONNECTED_152), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5686 ) );
  NAND2_X2 _f_permutation__U3966  ( .A1(_f_permutation__n5685 ), .A2(
        _f_permutation__n5686 ), .ZN(_f_permutation__n4451 ) );
  NAND2_X2 _f_permutation__U3965  ( .A1(_f_permutation__round_out[935]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5683 ) );
  NAND2_X2 _f_permutation__U3964  ( .A1(SYNOPSYS_UNCONNECTED_153), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5684 ) );
  NAND2_X2 _f_permutation__U3963  ( .A1(_f_permutation__n5683 ), .A2(
        _f_permutation__n5684 ), .ZN(_f_permutation__n4452 ) );
  NAND2_X2 _f_permutation__U3962  ( .A1(_f_permutation__round_out[934]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5681 ) );
  NAND2_X2 _f_permutation__U3961  ( .A1(SYNOPSYS_UNCONNECTED_154), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5682 ) );
  NAND2_X2 _f_permutation__U3960  ( .A1(_f_permutation__n5681 ), .A2(
        _f_permutation__n5682 ), .ZN(_f_permutation__n4453 ) );
  NAND2_X2 _f_permutation__U3959  ( .A1(_f_permutation__round_out[933]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5679 ) );
  NAND2_X2 _f_permutation__U3958  ( .A1(SYNOPSYS_UNCONNECTED_155), .A2(
        _f_permutation__n7227 ), .ZN(_f_permutation__n5680 ) );
  NAND2_X2 _f_permutation__U3957  ( .A1(_f_permutation__n5679 ), .A2(
        _f_permutation__n5680 ), .ZN(_f_permutation__n4454 ) );
  NAND2_X2 _f_permutation__U3956  ( .A1(_f_permutation__round_out[932]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5677 ) );
  NAND2_X2 _f_permutation__U3955  ( .A1(SYNOPSYS_UNCONNECTED_156), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5678 ) );
  NAND2_X2 _f_permutation__U3954  ( .A1(_f_permutation__n5677 ), .A2(
        _f_permutation__n5678 ), .ZN(_f_permutation__n4455 ) );
  NAND2_X2 _f_permutation__U3953  ( .A1(_f_permutation__round_out[931]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5675 ) );
  NAND2_X2 _f_permutation__U3952  ( .A1(SYNOPSYS_UNCONNECTED_157), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5676 ) );
  NAND2_X2 _f_permutation__U3951  ( .A1(_f_permutation__n5675 ), .A2(
        _f_permutation__n5676 ), .ZN(_f_permutation__n4456 ) );
  NAND2_X2 _f_permutation__U3950  ( .A1(_f_permutation__round_out[930]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5673 ) );
  NAND2_X2 _f_permutation__U3949  ( .A1(SYNOPSYS_UNCONNECTED_158), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5674 ) );
  NAND2_X2 _f_permutation__U3948  ( .A1(_f_permutation__n5673 ), .A2(
        _f_permutation__n5674 ), .ZN(_f_permutation__n4457 ) );
  NAND2_X2 _f_permutation__U3947  ( .A1(_f_permutation__round_out[929]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5671 ) );
  NAND2_X2 _f_permutation__U3946  ( .A1(SYNOPSYS_UNCONNECTED_159), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5672 ) );
  NAND2_X2 _f_permutation__U3945  ( .A1(_f_permutation__n5671 ), .A2(
        _f_permutation__n5672 ), .ZN(_f_permutation__n4458 ) );
  NAND2_X2 _f_permutation__U3944  ( .A1(_f_permutation__round_out[928]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5669 ) );
  NAND2_X2 _f_permutation__U3943  ( .A1(SYNOPSYS_UNCONNECTED_160), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5670 ) );
  NAND2_X2 _f_permutation__U3942  ( .A1(_f_permutation__n5669 ), .A2(
        _f_permutation__n5670 ), .ZN(_f_permutation__n4459 ) );
  NAND2_X2 _f_permutation__U3941  ( .A1(_f_permutation__round_out[927]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5667 ) );
  NAND2_X2 _f_permutation__U3940  ( .A1(SYNOPSYS_UNCONNECTED_161), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5668 ) );
  NAND2_X2 _f_permutation__U3939  ( .A1(_f_permutation__n5667 ), .A2(
        _f_permutation__n5668 ), .ZN(_f_permutation__n4460 ) );
  NAND2_X2 _f_permutation__U3938  ( .A1(_f_permutation__round_out[926]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5665 ) );
  NAND2_X2 _f_permutation__U3937  ( .A1(SYNOPSYS_UNCONNECTED_162), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5666 ) );
  NAND2_X2 _f_permutation__U3936  ( .A1(_f_permutation__n5665 ), .A2(
        _f_permutation__n5666 ), .ZN(_f_permutation__n4461 ) );
  NAND2_X2 _f_permutation__U3935  ( .A1(_f_permutation__round_out[925]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5663 ) );
  NAND2_X2 _f_permutation__U3934  ( .A1(SYNOPSYS_UNCONNECTED_163), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5664 ) );
  NAND2_X2 _f_permutation__U3933  ( .A1(_f_permutation__n5663 ), .A2(
        _f_permutation__n5664 ), .ZN(_f_permutation__n4462 ) );
  NAND2_X2 _f_permutation__U3932  ( .A1(_f_permutation__round_out[924]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5661 ) );
  NAND2_X2 _f_permutation__U3931  ( .A1(SYNOPSYS_UNCONNECTED_164), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5662 ) );
  NAND2_X2 _f_permutation__U3930  ( .A1(_f_permutation__n5661 ), .A2(
        _f_permutation__n5662 ), .ZN(_f_permutation__n4463 ) );
  NAND2_X2 _f_permutation__U3929  ( .A1(_f_permutation__round_out[923]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5659 ) );
  NAND2_X2 _f_permutation__U3928  ( .A1(SYNOPSYS_UNCONNECTED_165), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5660 ) );
  NAND2_X2 _f_permutation__U3927  ( .A1(_f_permutation__n5659 ), .A2(
        _f_permutation__n5660 ), .ZN(_f_permutation__n4464 ) );
  NAND2_X2 _f_permutation__U3926  ( .A1(_f_permutation__round_out[922]), .A2(
        _f_permutation__n7118 ), .ZN(_f_permutation__n5657 ) );
  NAND2_X2 _f_permutation__U3925  ( .A1(SYNOPSYS_UNCONNECTED_166), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5658 ) );
  NAND2_X2 _f_permutation__U3924  ( .A1(_f_permutation__n5657 ), .A2(
        _f_permutation__n5658 ), .ZN(_f_permutation__n4465 ) );
  NAND2_X2 _f_permutation__U3923  ( .A1(_f_permutation__round_out[921]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5655 ) );
  NAND2_X2 _f_permutation__U3922  ( .A1(SYNOPSYS_UNCONNECTED_167), .A2(
        _f_permutation__n7228 ), .ZN(_f_permutation__n5656 ) );
  NAND2_X2 _f_permutation__U3921  ( .A1(_f_permutation__n5655 ), .A2(
        _f_permutation__n5656 ), .ZN(_f_permutation__n4466 ) );
  NAND2_X2 _f_permutation__U3920  ( .A1(_f_permutation__round_out[920]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5653 ) );
  NAND2_X2 _f_permutation__U3919  ( .A1(SYNOPSYS_UNCONNECTED_168), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5654 ) );
  NAND2_X2 _f_permutation__U3918  ( .A1(_f_permutation__n5653 ), .A2(
        _f_permutation__n5654 ), .ZN(_f_permutation__n4467 ) );
  NAND2_X2 _f_permutation__U3917  ( .A1(_f_permutation__round_out[919]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5651 ) );
  NAND2_X2 _f_permutation__U3916  ( .A1(SYNOPSYS_UNCONNECTED_169), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5652 ) );
  NAND2_X2 _f_permutation__U3915  ( .A1(_f_permutation__n5651 ), .A2(
        _f_permutation__n5652 ), .ZN(_f_permutation__n4468 ) );
  NAND2_X2 _f_permutation__U3914  ( .A1(_f_permutation__round_out[918]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5649 ) );
  NAND2_X2 _f_permutation__U3913  ( .A1(SYNOPSYS_UNCONNECTED_170), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5650 ) );
  NAND2_X2 _f_permutation__U3912  ( .A1(_f_permutation__n5649 ), .A2(
        _f_permutation__n5650 ), .ZN(_f_permutation__n4469 ) );
  NAND2_X2 _f_permutation__U3911  ( .A1(_f_permutation__round_out[917]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5647 ) );
  NAND2_X2 _f_permutation__U3910  ( .A1(SYNOPSYS_UNCONNECTED_171), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5648 ) );
  NAND2_X2 _f_permutation__U3909  ( .A1(_f_permutation__n5647 ), .A2(
        _f_permutation__n5648 ), .ZN(_f_permutation__n4470 ) );
  NAND2_X2 _f_permutation__U3908  ( .A1(_f_permutation__round_out[916]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5645 ) );
  NAND2_X2 _f_permutation__U3907  ( .A1(SYNOPSYS_UNCONNECTED_172), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5646 ) );
  NAND2_X2 _f_permutation__U3906  ( .A1(_f_permutation__n5645 ), .A2(
        _f_permutation__n5646 ), .ZN(_f_permutation__n4471 ) );
  NAND2_X2 _f_permutation__U3905  ( .A1(_f_permutation__round_out[915]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5643 ) );
  NAND2_X2 _f_permutation__U3904  ( .A1(SYNOPSYS_UNCONNECTED_173), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5644 ) );
  NAND2_X2 _f_permutation__U3903  ( .A1(_f_permutation__n5643 ), .A2(
        _f_permutation__n5644 ), .ZN(_f_permutation__n4472 ) );
  NAND2_X2 _f_permutation__U3902  ( .A1(_f_permutation__round_out[914]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5641 ) );
  NAND2_X2 _f_permutation__U3901  ( .A1(SYNOPSYS_UNCONNECTED_174), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5642 ) );
  NAND2_X2 _f_permutation__U3900  ( .A1(_f_permutation__n5641 ), .A2(
        _f_permutation__n5642 ), .ZN(_f_permutation__n4473 ) );
  NAND2_X2 _f_permutation__U3899  ( .A1(_f_permutation__round_out[913]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5639 ) );
  NAND2_X2 _f_permutation__U3898  ( .A1(SYNOPSYS_UNCONNECTED_175), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5640 ) );
  NAND2_X2 _f_permutation__U3897  ( .A1(_f_permutation__n5639 ), .A2(
        _f_permutation__n5640 ), .ZN(_f_permutation__n4474 ) );
  NAND2_X2 _f_permutation__U3896  ( .A1(_f_permutation__round_out[912]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5637 ) );
  NAND2_X2 _f_permutation__U3895  ( .A1(SYNOPSYS_UNCONNECTED_176), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5638 ) );
  NAND2_X2 _f_permutation__U3894  ( .A1(_f_permutation__n5637 ), .A2(
        _f_permutation__n5638 ), .ZN(_f_permutation__n4475 ) );
  NAND2_X2 _f_permutation__U3893  ( .A1(_f_permutation__round_out[911]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5635 ) );
  NAND2_X2 _f_permutation__U3892  ( .A1(SYNOPSYS_UNCONNECTED_177), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5636 ) );
  NAND2_X2 _f_permutation__U3891  ( .A1(_f_permutation__n5635 ), .A2(
        _f_permutation__n5636 ), .ZN(_f_permutation__n4476 ) );
  NAND2_X2 _f_permutation__U3890  ( .A1(_f_permutation__round_out[910]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5633 ) );
  NAND2_X2 _f_permutation__U3889  ( .A1(SYNOPSYS_UNCONNECTED_178), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5634 ) );
  NAND2_X2 _f_permutation__U3888  ( .A1(_f_permutation__n5633 ), .A2(
        _f_permutation__n5634 ), .ZN(_f_permutation__n4477 ) );
  NAND2_X2 _f_permutation__U3887  ( .A1(_f_permutation__round_out[909]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5631 ) );
  NAND2_X2 _f_permutation__U3886  ( .A1(SYNOPSYS_UNCONNECTED_179), .A2(
        _f_permutation__n7229 ), .ZN(_f_permutation__n5632 ) );
  NAND2_X2 _f_permutation__U3885  ( .A1(_f_permutation__n5631 ), .A2(
        _f_permutation__n5632 ), .ZN(_f_permutation__n4478 ) );
  NAND2_X2 _f_permutation__U3884  ( .A1(_f_permutation__round_out[908]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5629 ) );
  NAND2_X2 _f_permutation__U3883  ( .A1(SYNOPSYS_UNCONNECTED_180), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5630 ) );
  NAND2_X2 _f_permutation__U3882  ( .A1(_f_permutation__n5629 ), .A2(
        _f_permutation__n5630 ), .ZN(_f_permutation__n4479 ) );
  NAND2_X2 _f_permutation__U3881  ( .A1(_f_permutation__round_out[907]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5627 ) );
  NAND2_X2 _f_permutation__U3880  ( .A1(SYNOPSYS_UNCONNECTED_181), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5628 ) );
  NAND2_X2 _f_permutation__U3879  ( .A1(_f_permutation__n5627 ), .A2(
        _f_permutation__n5628 ), .ZN(_f_permutation__n4480 ) );
  NAND2_X2 _f_permutation__U3878  ( .A1(_f_permutation__round_out[906]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5625 ) );
  NAND2_X2 _f_permutation__U3877  ( .A1(SYNOPSYS_UNCONNECTED_182), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5626 ) );
  NAND2_X2 _f_permutation__U3876  ( .A1(_f_permutation__n5625 ), .A2(
        _f_permutation__n5626 ), .ZN(_f_permutation__n4481 ) );
  NAND2_X2 _f_permutation__U3875  ( .A1(_f_permutation__round_out[905]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5623 ) );
  NAND2_X2 _f_permutation__U3874  ( .A1(SYNOPSYS_UNCONNECTED_183), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5624 ) );
  NAND2_X2 _f_permutation__U3873  ( .A1(_f_permutation__n5623 ), .A2(
        _f_permutation__n5624 ), .ZN(_f_permutation__n4482 ) );
  NAND2_X2 _f_permutation__U3872  ( .A1(_f_permutation__round_out[904]), .A2(
        _f_permutation__n7117 ), .ZN(_f_permutation__n5621 ) );
  NAND2_X2 _f_permutation__U3871  ( .A1(SYNOPSYS_UNCONNECTED_184), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5622 ) );
  NAND2_X2 _f_permutation__U3870  ( .A1(_f_permutation__n5621 ), .A2(
        _f_permutation__n5622 ), .ZN(_f_permutation__n4483 ) );
  NAND2_X2 _f_permutation__U3869  ( .A1(_f_permutation__round_out[903]), .A2(
        _f_permutation__n7116 ), .ZN(_f_permutation__n5619 ) );
  NAND2_X2 _f_permutation__U3868  ( .A1(SYNOPSYS_UNCONNECTED_185), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5620 ) );
  NAND2_X2 _f_permutation__U3867  ( .A1(_f_permutation__n5619 ), .A2(
        _f_permutation__n5620 ), .ZN(_f_permutation__n4484 ) );
  NAND2_X2 _f_permutation__U3866  ( .A1(_f_permutation__round_out[902]), .A2(
        _f_permutation__n7116 ), .ZN(_f_permutation__n5617 ) );
  NAND2_X2 _f_permutation__U3865  ( .A1(SYNOPSYS_UNCONNECTED_186), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5618 ) );
  NAND2_X2 _f_permutation__U3864  ( .A1(_f_permutation__n5617 ), .A2(
        _f_permutation__n5618 ), .ZN(_f_permutation__n4485 ) );
  NAND2_X2 _f_permutation__U3863  ( .A1(_f_permutation__round_out[901]), .A2(
        _f_permutation__n7116 ), .ZN(_f_permutation__n5615 ) );
  NAND2_X2 _f_permutation__U3862  ( .A1(SYNOPSYS_UNCONNECTED_187), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5616 ) );
  NAND2_X2 _f_permutation__U3861  ( .A1(_f_permutation__n5615 ), .A2(
        _f_permutation__n5616 ), .ZN(_f_permutation__n4486 ) );
  NAND2_X2 _f_permutation__U3860  ( .A1(_f_permutation__round_out[900]), .A2(
        _f_permutation__n7119 ), .ZN(_f_permutation__n5613 ) );
  NAND2_X2 _f_permutation__U3859  ( .A1(SYNOPSYS_UNCONNECTED_188), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5614 ) );
  NAND2_X2 _f_permutation__U3858  ( .A1(_f_permutation__n5613 ), .A2(
        _f_permutation__n5614 ), .ZN(_f_permutation__n4487 ) );
  NAND2_X2 _f_permutation__U3857  ( .A1(_f_permutation__round_out[899]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5611 ) );
  NAND2_X2 _f_permutation__U3856  ( .A1(SYNOPSYS_UNCONNECTED_189), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5612 ) );
  NAND2_X2 _f_permutation__U3855  ( .A1(_f_permutation__n5611 ), .A2(
        _f_permutation__n5612 ), .ZN(_f_permutation__n4488 ) );
  NAND2_X2 _f_permutation__U3854  ( .A1(_f_permutation__round_out[898]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5609 ) );
  NAND2_X2 _f_permutation__U3853  ( .A1(SYNOPSYS_UNCONNECTED_190), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5610 ) );
  NAND2_X2 _f_permutation__U3852  ( .A1(_f_permutation__n5609 ), .A2(
        _f_permutation__n5610 ), .ZN(_f_permutation__n4489 ) );
  NAND2_X2 _f_permutation__U3851  ( .A1(_f_permutation__round_out[897]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5607 ) );
  NAND2_X2 _f_permutation__U3850  ( .A1(SYNOPSYS_UNCONNECTED_191), .A2(
        _f_permutation__n7230 ), .ZN(_f_permutation__n5608 ) );
  NAND2_X2 _f_permutation__U3849  ( .A1(_f_permutation__n5607 ), .A2(
        _f_permutation__n5608 ), .ZN(_f_permutation__n4490 ) );
  NAND2_X2 _f_permutation__U3848  ( .A1(_f_permutation__round_out[896]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5605 ) );
  NAND2_X2 _f_permutation__U3847  ( .A1(SYNOPSYS_UNCONNECTED_192), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5606 ) );
  NAND2_X2 _f_permutation__U3846  ( .A1(_f_permutation__n5605 ), .A2(
        _f_permutation__n5606 ), .ZN(_f_permutation__n4491 ) );
  NAND2_X2 _f_permutation__U3845  ( .A1(_f_permutation__round_out[895]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5603 ) );
  NAND2_X2 _f_permutation__U3844  ( .A1(SYNOPSYS_UNCONNECTED_193), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5604 ) );
  NAND2_X2 _f_permutation__U3843  ( .A1(_f_permutation__n5603 ), .A2(
        _f_permutation__n5604 ), .ZN(_f_permutation__n4492 ) );
  NAND2_X2 _f_permutation__U3842  ( .A1(_f_permutation__round_out[894]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5601 ) );
  NAND2_X2 _f_permutation__U3841  ( .A1(SYNOPSYS_UNCONNECTED_194), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5602 ) );
  NAND2_X2 _f_permutation__U3840  ( .A1(_f_permutation__n5601 ), .A2(
        _f_permutation__n5602 ), .ZN(_f_permutation__n4493 ) );
  NAND2_X2 _f_permutation__U3839  ( .A1(_f_permutation__round_out[893]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5599 ) );
  NAND2_X2 _f_permutation__U3838  ( .A1(SYNOPSYS_UNCONNECTED_195), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5600 ) );
  NAND2_X2 _f_permutation__U3837  ( .A1(_f_permutation__n5599 ), .A2(
        _f_permutation__n5600 ), .ZN(_f_permutation__n4494 ) );
  NAND2_X2 _f_permutation__U3836  ( .A1(_f_permutation__round_out[892]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5597 ) );
  NAND2_X2 _f_permutation__U3835  ( .A1(SYNOPSYS_UNCONNECTED_196), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5598 ) );
  NAND2_X2 _f_permutation__U3834  ( .A1(_f_permutation__n5597 ), .A2(
        _f_permutation__n5598 ), .ZN(_f_permutation__n4495 ) );
  NAND2_X2 _f_permutation__U3833  ( .A1(_f_permutation__round_out[891]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5595 ) );
  NAND2_X2 _f_permutation__U3832  ( .A1(SYNOPSYS_UNCONNECTED_197), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5596 ) );
  NAND2_X2 _f_permutation__U3831  ( .A1(_f_permutation__n5595 ), .A2(
        _f_permutation__n5596 ), .ZN(_f_permutation__n4496 ) );
  NAND2_X2 _f_permutation__U3830  ( .A1(_f_permutation__round_out[890]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5593 ) );
  NAND2_X2 _f_permutation__U3829  ( .A1(SYNOPSYS_UNCONNECTED_198), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5594 ) );
  NAND2_X2 _f_permutation__U3828  ( .A1(_f_permutation__n5593 ), .A2(
        _f_permutation__n5594 ), .ZN(_f_permutation__n4497 ) );
  NAND2_X2 _f_permutation__U3827  ( .A1(_f_permutation__round_out[889]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5591 ) );
  NAND2_X2 _f_permutation__U3826  ( .A1(SYNOPSYS_UNCONNECTED_199), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5592 ) );
  NAND2_X2 _f_permutation__U3825  ( .A1(_f_permutation__n5591 ), .A2(
        _f_permutation__n5592 ), .ZN(_f_permutation__n4498 ) );
  NAND2_X2 _f_permutation__U3824  ( .A1(_f_permutation__round_out[888]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5589 ) );
  NAND2_X2 _f_permutation__U3823  ( .A1(SYNOPSYS_UNCONNECTED_200), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5590 ) );
  NAND2_X2 _f_permutation__U3822  ( .A1(_f_permutation__n5589 ), .A2(
        _f_permutation__n5590 ), .ZN(_f_permutation__n4499 ) );
  NAND2_X2 _f_permutation__U3821  ( .A1(_f_permutation__round_out[887]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5587 ) );
  NAND2_X2 _f_permutation__U3820  ( .A1(SYNOPSYS_UNCONNECTED_201), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5588 ) );
  NAND2_X2 _f_permutation__U3819  ( .A1(_f_permutation__n5587 ), .A2(
        _f_permutation__n5588 ), .ZN(_f_permutation__n4500 ) );
  NAND2_X2 _f_permutation__U3818  ( .A1(_f_permutation__round_out[886]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5585 ) );
  NAND2_X2 _f_permutation__U3817  ( .A1(SYNOPSYS_UNCONNECTED_202), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5586 ) );
  NAND2_X2 _f_permutation__U3816  ( .A1(_f_permutation__n5585 ), .A2(
        _f_permutation__n5586 ), .ZN(_f_permutation__n4501 ) );
  NAND2_X2 _f_permutation__U3815  ( .A1(_f_permutation__round_out[885]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5583 ) );
  NAND2_X2 _f_permutation__U3814  ( .A1(SYNOPSYS_UNCONNECTED_203), .A2(
        _f_permutation__n7231 ), .ZN(_f_permutation__n5584 ) );
  NAND2_X2 _f_permutation__U3813  ( .A1(_f_permutation__n5583 ), .A2(
        _f_permutation__n5584 ), .ZN(_f_permutation__n4502 ) );
  NAND2_X2 _f_permutation__U3812  ( .A1(_f_permutation__round_out[884]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5581 ) );
  NAND2_X2 _f_permutation__U3811  ( .A1(SYNOPSYS_UNCONNECTED_204), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5582 ) );
  NAND2_X2 _f_permutation__U3810  ( .A1(_f_permutation__n5581 ), .A2(
        _f_permutation__n5582 ), .ZN(_f_permutation__n4503 ) );
  NAND2_X2 _f_permutation__U3809  ( .A1(_f_permutation__round_out[883]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5579 ) );
  NAND2_X2 _f_permutation__U3808  ( .A1(SYNOPSYS_UNCONNECTED_205), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5580 ) );
  NAND2_X2 _f_permutation__U3807  ( .A1(_f_permutation__n5579 ), .A2(
        _f_permutation__n5580 ), .ZN(_f_permutation__n4504 ) );
  NAND2_X2 _f_permutation__U3806  ( .A1(_f_permutation__round_out[882]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5577 ) );
  NAND2_X2 _f_permutation__U3805  ( .A1(SYNOPSYS_UNCONNECTED_206), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5578 ) );
  NAND2_X2 _f_permutation__U3804  ( .A1(_f_permutation__n5577 ), .A2(
        _f_permutation__n5578 ), .ZN(_f_permutation__n4505 ) );
  NAND2_X2 _f_permutation__U3803  ( .A1(_f_permutation__round_out[881]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5575 ) );
  NAND2_X2 _f_permutation__U3802  ( .A1(SYNOPSYS_UNCONNECTED_207), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5576 ) );
  NAND2_X2 _f_permutation__U3801  ( .A1(_f_permutation__n5575 ), .A2(
        _f_permutation__n5576 ), .ZN(_f_permutation__n4506 ) );
  NAND2_X2 _f_permutation__U3800  ( .A1(_f_permutation__round_out[880]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5573 ) );
  NAND2_X2 _f_permutation__U3799  ( .A1(SYNOPSYS_UNCONNECTED_208), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5574 ) );
  NAND2_X2 _f_permutation__U3798  ( .A1(_f_permutation__n5573 ), .A2(
        _f_permutation__n5574 ), .ZN(_f_permutation__n4507 ) );
  NAND2_X2 _f_permutation__U3797  ( .A1(_f_permutation__round_out[879]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5571 ) );
  NAND2_X2 _f_permutation__U3796  ( .A1(SYNOPSYS_UNCONNECTED_209), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5572 ) );
  NAND2_X2 _f_permutation__U3795  ( .A1(_f_permutation__n5571 ), .A2(
        _f_permutation__n5572 ), .ZN(_f_permutation__n4508 ) );
  NAND2_X2 _f_permutation__U3794  ( .A1(_f_permutation__round_out[878]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5569 ) );
  NAND2_X2 _f_permutation__U3793  ( .A1(SYNOPSYS_UNCONNECTED_210), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5570 ) );
  NAND2_X2 _f_permutation__U3792  ( .A1(_f_permutation__n5569 ), .A2(
        _f_permutation__n5570 ), .ZN(_f_permutation__n4509 ) );
  NAND2_X2 _f_permutation__U3791  ( .A1(_f_permutation__round_out[877]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5567 ) );
  NAND2_X2 _f_permutation__U3790  ( .A1(SYNOPSYS_UNCONNECTED_211), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5568 ) );
  NAND2_X2 _f_permutation__U3789  ( .A1(_f_permutation__n5567 ), .A2(
        _f_permutation__n5568 ), .ZN(_f_permutation__n4510 ) );
  NAND2_X2 _f_permutation__U3788  ( .A1(_f_permutation__round_out[876]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5565 ) );
  NAND2_X2 _f_permutation__U3787  ( .A1(SYNOPSYS_UNCONNECTED_212), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5566 ) );
  NAND2_X2 _f_permutation__U3786  ( .A1(_f_permutation__n5565 ), .A2(
        _f_permutation__n5566 ), .ZN(_f_permutation__n4511 ) );
  NAND2_X2 _f_permutation__U3785  ( .A1(_f_permutation__round_out[875]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5563 ) );
  NAND2_X2 _f_permutation__U3784  ( .A1(SYNOPSYS_UNCONNECTED_213), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5564 ) );
  NAND2_X2 _f_permutation__U3783  ( .A1(_f_permutation__n5563 ), .A2(
        _f_permutation__n5564 ), .ZN(_f_permutation__n4512 ) );
  NAND2_X2 _f_permutation__U3782  ( .A1(_f_permutation__round_out[874]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5561 ) );
  NAND2_X2 _f_permutation__U3781  ( .A1(SYNOPSYS_UNCONNECTED_214), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5562 ) );
  NAND2_X2 _f_permutation__U3780  ( .A1(_f_permutation__n5561 ), .A2(
        _f_permutation__n5562 ), .ZN(_f_permutation__n4513 ) );
  NAND2_X2 _f_permutation__U3779  ( .A1(_f_permutation__round_out[873]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5559 ) );
  NAND2_X2 _f_permutation__U3778  ( .A1(SYNOPSYS_UNCONNECTED_215), .A2(
        _f_permutation__n7232 ), .ZN(_f_permutation__n5560 ) );
  NAND2_X2 _f_permutation__U3777  ( .A1(_f_permutation__n5559 ), .A2(
        _f_permutation__n5560 ), .ZN(_f_permutation__n4514 ) );
  NAND2_X2 _f_permutation__U3776  ( .A1(_f_permutation__round_out[872]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5557 ) );
  NAND2_X2 _f_permutation__U3775  ( .A1(SYNOPSYS_UNCONNECTED_216), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5558 ) );
  NAND2_X2 _f_permutation__U3774  ( .A1(_f_permutation__n5557 ), .A2(
        _f_permutation__n5558 ), .ZN(_f_permutation__n4515 ) );
  NAND2_X2 _f_permutation__U3773  ( .A1(_f_permutation__round_out[871]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5555 ) );
  NAND2_X2 _f_permutation__U3772  ( .A1(SYNOPSYS_UNCONNECTED_217), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5556 ) );
  NAND2_X2 _f_permutation__U3771  ( .A1(_f_permutation__n5555 ), .A2(
        _f_permutation__n5556 ), .ZN(_f_permutation__n4516 ) );
  NAND2_X2 _f_permutation__U3770  ( .A1(_f_permutation__round_out[870]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5553 ) );
  NAND2_X2 _f_permutation__U3769  ( .A1(SYNOPSYS_UNCONNECTED_218), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5554 ) );
  NAND2_X2 _f_permutation__U3768  ( .A1(_f_permutation__n5553 ), .A2(
        _f_permutation__n5554 ), .ZN(_f_permutation__n4517 ) );
  NAND2_X2 _f_permutation__U3767  ( .A1(_f_permutation__round_out[869]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5551 ) );
  NAND2_X2 _f_permutation__U3766  ( .A1(SYNOPSYS_UNCONNECTED_219), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5552 ) );
  NAND2_X2 _f_permutation__U3765  ( .A1(_f_permutation__n5551 ), .A2(
        _f_permutation__n5552 ), .ZN(_f_permutation__n4518 ) );
  NAND2_X2 _f_permutation__U3764  ( .A1(_f_permutation__round_out[868]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5549 ) );
  NAND2_X2 _f_permutation__U3763  ( .A1(SYNOPSYS_UNCONNECTED_220), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5550 ) );
  NAND2_X2 _f_permutation__U3762  ( .A1(_f_permutation__n5549 ), .A2(
        _f_permutation__n5550 ), .ZN(_f_permutation__n4519 ) );
  NAND2_X2 _f_permutation__U3761  ( .A1(_f_permutation__round_out[867]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5547 ) );
  NAND2_X2 _f_permutation__U3760  ( .A1(SYNOPSYS_UNCONNECTED_221), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5548 ) );
  NAND2_X2 _f_permutation__U3759  ( .A1(_f_permutation__n5547 ), .A2(
        _f_permutation__n5548 ), .ZN(_f_permutation__n4520 ) );
  NAND2_X2 _f_permutation__U3758  ( .A1(_f_permutation__round_out[866]), .A2(
        _f_permutation__n7126 ), .ZN(_f_permutation__n5545 ) );
  NAND2_X2 _f_permutation__U3757  ( .A1(SYNOPSYS_UNCONNECTED_222), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5546 ) );
  NAND2_X2 _f_permutation__U3756  ( .A1(_f_permutation__n5545 ), .A2(
        _f_permutation__n5546 ), .ZN(_f_permutation__n4521 ) );
  NAND2_X2 _f_permutation__U3755  ( .A1(_f_permutation__round_out[865]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5543 ) );
  NAND2_X2 _f_permutation__U3754  ( .A1(SYNOPSYS_UNCONNECTED_223), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5544 ) );
  NAND2_X2 _f_permutation__U3753  ( .A1(_f_permutation__n5543 ), .A2(
        _f_permutation__n5544 ), .ZN(_f_permutation__n4522 ) );
  NAND2_X2 _f_permutation__U3752  ( .A1(_f_permutation__round_out[864]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5541 ) );
  NAND2_X2 _f_permutation__U3751  ( .A1(SYNOPSYS_UNCONNECTED_224), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5542 ) );
  NAND2_X2 _f_permutation__U3750  ( .A1(_f_permutation__n5541 ), .A2(
        _f_permutation__n5542 ), .ZN(_f_permutation__n4523 ) );
  NAND2_X2 _f_permutation__U3749  ( .A1(_f_permutation__round_out[863]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5539 ) );
  NAND2_X2 _f_permutation__U3748  ( .A1(SYNOPSYS_UNCONNECTED_225), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5540 ) );
  NAND2_X2 _f_permutation__U3747  ( .A1(_f_permutation__n5539 ), .A2(
        _f_permutation__n5540 ), .ZN(_f_permutation__n4524 ) );
  NAND2_X2 _f_permutation__U3746  ( .A1(_f_permutation__round_out[862]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5537 ) );
  NAND2_X2 _f_permutation__U3745  ( .A1(SYNOPSYS_UNCONNECTED_226), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5538 ) );
  NAND2_X2 _f_permutation__U3744  ( .A1(_f_permutation__n5537 ), .A2(
        _f_permutation__n5538 ), .ZN(_f_permutation__n4525 ) );
  NAND2_X2 _f_permutation__U3743  ( .A1(_f_permutation__round_out[861]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5535 ) );
  NAND2_X2 _f_permutation__U3742  ( .A1(SYNOPSYS_UNCONNECTED_227), .A2(
        _f_permutation__n7233 ), .ZN(_f_permutation__n5536 ) );
  NAND2_X2 _f_permutation__U3741  ( .A1(_f_permutation__n5535 ), .A2(
        _f_permutation__n5536 ), .ZN(_f_permutation__n4526 ) );
  NAND2_X2 _f_permutation__U3740  ( .A1(_f_permutation__round_out[860]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5533 ) );
  NAND2_X2 _f_permutation__U3739  ( .A1(SYNOPSYS_UNCONNECTED_228), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5534 ) );
  NAND2_X2 _f_permutation__U3738  ( .A1(_f_permutation__n5533 ), .A2(
        _f_permutation__n5534 ), .ZN(_f_permutation__n4527 ) );
  NAND2_X2 _f_permutation__U3737  ( .A1(_f_permutation__round_out[859]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5531 ) );
  NAND2_X2 _f_permutation__U3736  ( .A1(SYNOPSYS_UNCONNECTED_229), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5532 ) );
  NAND2_X2 _f_permutation__U3735  ( .A1(_f_permutation__n5531 ), .A2(
        _f_permutation__n5532 ), .ZN(_f_permutation__n4528 ) );
  NAND2_X2 _f_permutation__U3734  ( .A1(_f_permutation__round_out[858]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5529 ) );
  NAND2_X2 _f_permutation__U3733  ( .A1(SYNOPSYS_UNCONNECTED_230), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5530 ) );
  NAND2_X2 _f_permutation__U3732  ( .A1(_f_permutation__n5529 ), .A2(
        _f_permutation__n5530 ), .ZN(_f_permutation__n4529 ) );
  NAND2_X2 _f_permutation__U3731  ( .A1(_f_permutation__round_out[857]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5527 ) );
  NAND2_X2 _f_permutation__U3730  ( .A1(SYNOPSYS_UNCONNECTED_231), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5528 ) );
  NAND2_X2 _f_permutation__U3729  ( .A1(_f_permutation__n5527 ), .A2(
        _f_permutation__n5528 ), .ZN(_f_permutation__n4530 ) );
  NAND2_X2 _f_permutation__U3728  ( .A1(_f_permutation__round_out[856]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5525 ) );
  NAND2_X2 _f_permutation__U3727  ( .A1(SYNOPSYS_UNCONNECTED_232), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5526 ) );
  NAND2_X2 _f_permutation__U3726  ( .A1(_f_permutation__n5525 ), .A2(
        _f_permutation__n5526 ), .ZN(_f_permutation__n4531 ) );
  NAND2_X2 _f_permutation__U3725  ( .A1(_f_permutation__round_out[855]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5523 ) );
  NAND2_X2 _f_permutation__U3724  ( .A1(SYNOPSYS_UNCONNECTED_233), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5524 ) );
  NAND2_X2 _f_permutation__U3723  ( .A1(_f_permutation__n5523 ), .A2(
        _f_permutation__n5524 ), .ZN(_f_permutation__n4532 ) );
  NAND2_X2 _f_permutation__U3722  ( .A1(_f_permutation__round_out[854]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5521 ) );
  NAND2_X2 _f_permutation__U3721  ( .A1(SYNOPSYS_UNCONNECTED_234), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5522 ) );
  NAND2_X2 _f_permutation__U3720  ( .A1(_f_permutation__n5521 ), .A2(
        _f_permutation__n5522 ), .ZN(_f_permutation__n4533 ) );
  NAND2_X2 _f_permutation__U3719  ( .A1(_f_permutation__round_out[853]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5519 ) );
  NAND2_X2 _f_permutation__U3718  ( .A1(SYNOPSYS_UNCONNECTED_235), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5520 ) );
  NAND2_X2 _f_permutation__U3717  ( .A1(_f_permutation__n5519 ), .A2(
        _f_permutation__n5520 ), .ZN(_f_permutation__n4534 ) );
  NAND2_X2 _f_permutation__U3716  ( .A1(_f_permutation__round_out[852]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5517 ) );
  NAND2_X2 _f_permutation__U3715  ( .A1(SYNOPSYS_UNCONNECTED_236), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5518 ) );
  NAND2_X2 _f_permutation__U3714  ( .A1(_f_permutation__n5517 ), .A2(
        _f_permutation__n5518 ), .ZN(_f_permutation__n4535 ) );
  NAND2_X2 _f_permutation__U3713  ( .A1(_f_permutation__round_out[851]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5515 ) );
  NAND2_X2 _f_permutation__U3712  ( .A1(SYNOPSYS_UNCONNECTED_237), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5516 ) );
  NAND2_X2 _f_permutation__U3711  ( .A1(_f_permutation__n5515 ), .A2(
        _f_permutation__n5516 ), .ZN(_f_permutation__n4536 ) );
  NAND2_X2 _f_permutation__U3710  ( .A1(_f_permutation__round_out[850]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5513 ) );
  NAND2_X2 _f_permutation__U3709  ( .A1(SYNOPSYS_UNCONNECTED_238), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5514 ) );
  NAND2_X2 _f_permutation__U3708  ( .A1(_f_permutation__n5513 ), .A2(
        _f_permutation__n5514 ), .ZN(_f_permutation__n4537 ) );
  NAND2_X2 _f_permutation__U3707  ( .A1(_f_permutation__round_out[849]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5511 ) );
  NAND2_X2 _f_permutation__U3706  ( .A1(SYNOPSYS_UNCONNECTED_239), .A2(
        _f_permutation__n7234 ), .ZN(_f_permutation__n5512 ) );
  NAND2_X2 _f_permutation__U3705  ( .A1(_f_permutation__n5511 ), .A2(
        _f_permutation__n5512 ), .ZN(_f_permutation__n4538 ) );
  NAND2_X2 _f_permutation__U3704  ( .A1(_f_permutation__round_out[848]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5509 ) );
  NAND2_X2 _f_permutation__U3703  ( .A1(SYNOPSYS_UNCONNECTED_240), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5510 ) );
  NAND2_X2 _f_permutation__U3702  ( .A1(_f_permutation__n5509 ), .A2(
        _f_permutation__n5510 ), .ZN(_f_permutation__n4539 ) );
  NAND2_X2 _f_permutation__U3701  ( .A1(_f_permutation__round_out[847]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5507 ) );
  NAND2_X2 _f_permutation__U3700  ( .A1(SYNOPSYS_UNCONNECTED_241), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5508 ) );
  NAND2_X2 _f_permutation__U3699  ( .A1(_f_permutation__n5507 ), .A2(
        _f_permutation__n5508 ), .ZN(_f_permutation__n4540 ) );
  NAND2_X2 _f_permutation__U3698  ( .A1(_f_permutation__round_out[846]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5505 ) );
  NAND2_X2 _f_permutation__U3697  ( .A1(SYNOPSYS_UNCONNECTED_242), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5506 ) );
  NAND2_X2 _f_permutation__U3696  ( .A1(_f_permutation__n5505 ), .A2(
        _f_permutation__n5506 ), .ZN(_f_permutation__n4541 ) );
  NAND2_X2 _f_permutation__U3695  ( .A1(_f_permutation__round_out[845]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5503 ) );
  NAND2_X2 _f_permutation__U3694  ( .A1(SYNOPSYS_UNCONNECTED_243), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5504 ) );
  NAND2_X2 _f_permutation__U3693  ( .A1(_f_permutation__n5503 ), .A2(
        _f_permutation__n5504 ), .ZN(_f_permutation__n4542 ) );
  NAND2_X2 _f_permutation__U3692  ( .A1(_f_permutation__round_out[844]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5501 ) );
  NAND2_X2 _f_permutation__U3691  ( .A1(SYNOPSYS_UNCONNECTED_244), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5502 ) );
  NAND2_X2 _f_permutation__U3690  ( .A1(_f_permutation__n5501 ), .A2(
        _f_permutation__n5502 ), .ZN(_f_permutation__n4543 ) );
  NAND2_X2 _f_permutation__U3689  ( .A1(_f_permutation__round_out[843]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5499 ) );
  NAND2_X2 _f_permutation__U3688  ( .A1(SYNOPSYS_UNCONNECTED_245), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5500 ) );
  NAND2_X2 _f_permutation__U3687  ( .A1(_f_permutation__n5499 ), .A2(
        _f_permutation__n5500 ), .ZN(_f_permutation__n4544 ) );
  NAND2_X2 _f_permutation__U3686  ( .A1(_f_permutation__round_out[842]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5497 ) );
  NAND2_X2 _f_permutation__U3685  ( .A1(SYNOPSYS_UNCONNECTED_246), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5498 ) );
  NAND2_X2 _f_permutation__U3684  ( .A1(_f_permutation__n5497 ), .A2(
        _f_permutation__n5498 ), .ZN(_f_permutation__n4545 ) );
  NAND2_X2 _f_permutation__U3683  ( .A1(_f_permutation__round_out[841]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5495 ) );
  NAND2_X2 _f_permutation__U3682  ( .A1(SYNOPSYS_UNCONNECTED_247), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5496 ) );
  NAND2_X2 _f_permutation__U3681  ( .A1(_f_permutation__n5495 ), .A2(
        _f_permutation__n5496 ), .ZN(_f_permutation__n4546 ) );
  NAND2_X2 _f_permutation__U3680  ( .A1(_f_permutation__round_out[840]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5493 ) );
  NAND2_X2 _f_permutation__U3679  ( .A1(SYNOPSYS_UNCONNECTED_248), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5494 ) );
  NAND2_X2 _f_permutation__U3678  ( .A1(_f_permutation__n5493 ), .A2(
        _f_permutation__n5494 ), .ZN(_f_permutation__n4547 ) );
  NAND2_X2 _f_permutation__U3677  ( .A1(_f_permutation__round_out[839]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5491 ) );
  NAND2_X2 _f_permutation__U3676  ( .A1(SYNOPSYS_UNCONNECTED_249), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5492 ) );
  NAND2_X2 _f_permutation__U3675  ( .A1(_f_permutation__n5491 ), .A2(
        _f_permutation__n5492 ), .ZN(_f_permutation__n4548 ) );
  NAND2_X2 _f_permutation__U3674  ( .A1(_f_permutation__round_out[838]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5489 ) );
  NAND2_X2 _f_permutation__U3673  ( .A1(SYNOPSYS_UNCONNECTED_250), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5490 ) );
  NAND2_X2 _f_permutation__U3672  ( .A1(_f_permutation__n5489 ), .A2(
        _f_permutation__n5490 ), .ZN(_f_permutation__n4549 ) );
  NAND2_X2 _f_permutation__U3671  ( .A1(_f_permutation__round_out[837]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5487 ) );
  NAND2_X2 _f_permutation__U3670  ( .A1(SYNOPSYS_UNCONNECTED_251), .A2(
        _f_permutation__n7235 ), .ZN(_f_permutation__n5488 ) );
  NAND2_X2 _f_permutation__U3669  ( .A1(_f_permutation__n5487 ), .A2(
        _f_permutation__n5488 ), .ZN(_f_permutation__n4550 ) );
  NAND2_X2 _f_permutation__U3668  ( .A1(_f_permutation__round_out[836]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5485 ) );
  NAND2_X2 _f_permutation__U3667  ( .A1(SYNOPSYS_UNCONNECTED_252), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5486 ) );
  NAND2_X2 _f_permutation__U3666  ( .A1(_f_permutation__n5485 ), .A2(
        _f_permutation__n5486 ), .ZN(_f_permutation__n4551 ) );
  NAND2_X2 _f_permutation__U3665  ( .A1(_f_permutation__round_out[835]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5483 ) );
  NAND2_X2 _f_permutation__U3664  ( .A1(SYNOPSYS_UNCONNECTED_253), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5484 ) );
  NAND2_X2 _f_permutation__U3663  ( .A1(_f_permutation__n5483 ), .A2(
        _f_permutation__n5484 ), .ZN(_f_permutation__n4552 ) );
  NAND2_X2 _f_permutation__U3662  ( .A1(_f_permutation__round_out[834]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5481 ) );
  NAND2_X2 _f_permutation__U3661  ( .A1(SYNOPSYS_UNCONNECTED_254), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5482 ) );
  NAND2_X2 _f_permutation__U3660  ( .A1(_f_permutation__n5481 ), .A2(
        _f_permutation__n5482 ), .ZN(_f_permutation__n4553 ) );
  NAND2_X2 _f_permutation__U3659  ( .A1(_f_permutation__round_out[833]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5479 ) );
  NAND2_X2 _f_permutation__U3658  ( .A1(SYNOPSYS_UNCONNECTED_255), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5480 ) );
  NAND2_X2 _f_permutation__U3657  ( .A1(_f_permutation__n5479 ), .A2(
        _f_permutation__n5480 ), .ZN(_f_permutation__n4554 ) );
  NAND2_X2 _f_permutation__U3656  ( .A1(_f_permutation__round_out[832]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5477 ) );
  NAND2_X2 _f_permutation__U3655  ( .A1(SYNOPSYS_UNCONNECTED_256), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5478 ) );
  NAND2_X2 _f_permutation__U3654  ( .A1(_f_permutation__n5477 ), .A2(
        _f_permutation__n5478 ), .ZN(_f_permutation__n4555 ) );
  NAND2_X2 _f_permutation__U3653  ( .A1(_f_permutation__round_out[831]), .A2(
        _f_permutation__n7124 ), .ZN(_f_permutation__n5475 ) );
  NAND2_X2 _f_permutation__U3652  ( .A1(SYNOPSYS_UNCONNECTED_257), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5476 ) );
  NAND2_X2 _f_permutation__U3651  ( .A1(_f_permutation__n5475 ), .A2(
        _f_permutation__n5476 ), .ZN(_f_permutation__n4556 ) );
  NAND2_X2 _f_permutation__U3650  ( .A1(_f_permutation__round_out[830]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5473 ) );
  NAND2_X2 _f_permutation__U3649  ( .A1(SYNOPSYS_UNCONNECTED_258), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5474 ) );
  NAND2_X2 _f_permutation__U3648  ( .A1(_f_permutation__n5473 ), .A2(
        _f_permutation__n5474 ), .ZN(_f_permutation__n4557 ) );
  NAND2_X2 _f_permutation__U3647  ( .A1(_f_permutation__round_out[829]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5471 ) );
  NAND2_X2 _f_permutation__U3646  ( .A1(SYNOPSYS_UNCONNECTED_259), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5472 ) );
  NAND2_X2 _f_permutation__U3645  ( .A1(_f_permutation__n5471 ), .A2(
        _f_permutation__n5472 ), .ZN(_f_permutation__n4558 ) );
  NAND2_X2 _f_permutation__U3644  ( .A1(_f_permutation__round_out[828]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5469 ) );
  NAND2_X2 _f_permutation__U3643  ( .A1(SYNOPSYS_UNCONNECTED_260), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5470 ) );
  NAND2_X2 _f_permutation__U3642  ( .A1(_f_permutation__n5469 ), .A2(
        _f_permutation__n5470 ), .ZN(_f_permutation__n4559 ) );
  NAND2_X2 _f_permutation__U3641  ( .A1(_f_permutation__round_out[827]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5467 ) );
  NAND2_X2 _f_permutation__U3640  ( .A1(SYNOPSYS_UNCONNECTED_261), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5468 ) );
  NAND2_X2 _f_permutation__U3639  ( .A1(_f_permutation__n5467 ), .A2(
        _f_permutation__n5468 ), .ZN(_f_permutation__n4560 ) );
  NAND2_X2 _f_permutation__U3638  ( .A1(_f_permutation__round_out[826]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5465 ) );
  NAND2_X2 _f_permutation__U3637  ( .A1(SYNOPSYS_UNCONNECTED_262), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5466 ) );
  NAND2_X2 _f_permutation__U3636  ( .A1(_f_permutation__n5465 ), .A2(
        _f_permutation__n5466 ), .ZN(_f_permutation__n4561 ) );
  NAND2_X2 _f_permutation__U3635  ( .A1(_f_permutation__round_out[825]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5463 ) );
  NAND2_X2 _f_permutation__U3634  ( .A1(SYNOPSYS_UNCONNECTED_263), .A2(
        _f_permutation__n7236 ), .ZN(_f_permutation__n5464 ) );
  NAND2_X2 _f_permutation__U3633  ( .A1(_f_permutation__n5463 ), .A2(
        _f_permutation__n5464 ), .ZN(_f_permutation__n4562 ) );
  NAND2_X2 _f_permutation__U3632  ( .A1(_f_permutation__round_out[824]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5461 ) );
  NAND2_X2 _f_permutation__U3631  ( .A1(SYNOPSYS_UNCONNECTED_264), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5462 ) );
  NAND2_X2 _f_permutation__U3630  ( .A1(_f_permutation__n5461 ), .A2(
        _f_permutation__n5462 ), .ZN(_f_permutation__n4563 ) );
  NAND2_X2 _f_permutation__U3629  ( .A1(_f_permutation__round_out[823]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5459 ) );
  NAND2_X2 _f_permutation__U3628  ( .A1(SYNOPSYS_UNCONNECTED_265), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5460 ) );
  NAND2_X2 _f_permutation__U3627  ( .A1(_f_permutation__n5459 ), .A2(
        _f_permutation__n5460 ), .ZN(_f_permutation__n4564 ) );
  NAND2_X2 _f_permutation__U3626  ( .A1(_f_permutation__round_out[822]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5457 ) );
  NAND2_X2 _f_permutation__U3625  ( .A1(SYNOPSYS_UNCONNECTED_266), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5458 ) );
  NAND2_X2 _f_permutation__U3624  ( .A1(_f_permutation__n5457 ), .A2(
        _f_permutation__n5458 ), .ZN(_f_permutation__n4565 ) );
  NAND2_X2 _f_permutation__U3623  ( .A1(_f_permutation__round_out[821]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5455 ) );
  NAND2_X2 _f_permutation__U3622  ( .A1(SYNOPSYS_UNCONNECTED_267), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5456 ) );
  NAND2_X2 _f_permutation__U3621  ( .A1(_f_permutation__n5455 ), .A2(
        _f_permutation__n5456 ), .ZN(_f_permutation__n4566 ) );
  NAND2_X2 _f_permutation__U3620  ( .A1(_f_permutation__round_out[820]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5453 ) );
  NAND2_X2 _f_permutation__U3619  ( .A1(SYNOPSYS_UNCONNECTED_268), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5454 ) );
  NAND2_X2 _f_permutation__U3618  ( .A1(_f_permutation__n5453 ), .A2(
        _f_permutation__n5454 ), .ZN(_f_permutation__n4567 ) );
  NAND2_X2 _f_permutation__U3617  ( .A1(_f_permutation__round_out[819]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5451 ) );
  NAND2_X2 _f_permutation__U3616  ( .A1(SYNOPSYS_UNCONNECTED_269), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5452 ) );
  NAND2_X2 _f_permutation__U3615  ( .A1(_f_permutation__n5451 ), .A2(
        _f_permutation__n5452 ), .ZN(_f_permutation__n4568 ) );
  NAND2_X2 _f_permutation__U3614  ( .A1(_f_permutation__round_out[818]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5449 ) );
  NAND2_X2 _f_permutation__U3613  ( .A1(SYNOPSYS_UNCONNECTED_270), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5450 ) );
  NAND2_X2 _f_permutation__U3612  ( .A1(_f_permutation__n5449 ), .A2(
        _f_permutation__n5450 ), .ZN(_f_permutation__n4569 ) );
  NAND2_X2 _f_permutation__U3611  ( .A1(_f_permutation__round_out[817]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5447 ) );
  NAND2_X2 _f_permutation__U3610  ( .A1(SYNOPSYS_UNCONNECTED_271), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5448 ) );
  NAND2_X2 _f_permutation__U3609  ( .A1(_f_permutation__n5447 ), .A2(
        _f_permutation__n5448 ), .ZN(_f_permutation__n4570 ) );
  NAND2_X2 _f_permutation__U3608  ( .A1(_f_permutation__round_out[816]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5445 ) );
  NAND2_X2 _f_permutation__U3607  ( .A1(SYNOPSYS_UNCONNECTED_272), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5446 ) );
  NAND2_X2 _f_permutation__U3606  ( .A1(_f_permutation__n5445 ), .A2(
        _f_permutation__n5446 ), .ZN(_f_permutation__n4571 ) );
  NAND2_X2 _f_permutation__U3605  ( .A1(_f_permutation__round_out[815]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5443 ) );
  NAND2_X2 _f_permutation__U3604  ( .A1(SYNOPSYS_UNCONNECTED_273), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5444 ) );
  NAND2_X2 _f_permutation__U3603  ( .A1(_f_permutation__n5443 ), .A2(
        _f_permutation__n5444 ), .ZN(_f_permutation__n4572 ) );
  NAND2_X2 _f_permutation__U3602  ( .A1(_f_permutation__round_out[814]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5441 ) );
  NAND2_X2 _f_permutation__U3601  ( .A1(SYNOPSYS_UNCONNECTED_274), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5442 ) );
  NAND2_X2 _f_permutation__U3600  ( .A1(_f_permutation__n5441 ), .A2(
        _f_permutation__n5442 ), .ZN(_f_permutation__n4573 ) );
  NAND2_X2 _f_permutation__U3599  ( .A1(_f_permutation__round_out[813]), .A2(
        _f_permutation__n7123 ), .ZN(_f_permutation__n5439 ) );
  NAND2_X2 _f_permutation__U3598  ( .A1(SYNOPSYS_UNCONNECTED_275), .A2(
        _f_permutation__n7237 ), .ZN(_f_permutation__n5440 ) );
  NAND2_X2 _f_permutation__U3597  ( .A1(_f_permutation__n5439 ), .A2(
        _f_permutation__n5440 ), .ZN(_f_permutation__n4574 ) );
  NAND2_X2 _f_permutation__U3596  ( .A1(_f_permutation__round_out[812]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5437 ) );
  NAND2_X2 _f_permutation__U3595  ( .A1(SYNOPSYS_UNCONNECTED_276), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5438 ) );
  NAND2_X2 _f_permutation__U3594  ( .A1(_f_permutation__n5437 ), .A2(
        _f_permutation__n5438 ), .ZN(_f_permutation__n4575 ) );
  NAND2_X2 _f_permutation__U3593  ( .A1(_f_permutation__round_out[811]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5435 ) );
  NAND2_X2 _f_permutation__U3592  ( .A1(SYNOPSYS_UNCONNECTED_277), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5436 ) );
  NAND2_X2 _f_permutation__U3591  ( .A1(_f_permutation__n5435 ), .A2(
        _f_permutation__n5436 ), .ZN(_f_permutation__n4576 ) );
  NAND2_X2 _f_permutation__U3590  ( .A1(_f_permutation__round_out[810]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5433 ) );
  NAND2_X2 _f_permutation__U3589  ( .A1(SYNOPSYS_UNCONNECTED_278), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5434 ) );
  NAND2_X2 _f_permutation__U3588  ( .A1(_f_permutation__n5433 ), .A2(
        _f_permutation__n5434 ), .ZN(_f_permutation__n4577 ) );
  NAND2_X2 _f_permutation__U3587  ( .A1(_f_permutation__round_out[809]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5431 ) );
  NAND2_X2 _f_permutation__U3586  ( .A1(SYNOPSYS_UNCONNECTED_279), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5432 ) );
  NAND2_X2 _f_permutation__U3585  ( .A1(_f_permutation__n5431 ), .A2(
        _f_permutation__n5432 ), .ZN(_f_permutation__n4578 ) );
  NAND2_X2 _f_permutation__U3584  ( .A1(_f_permutation__round_out[808]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5429 ) );
  NAND2_X2 _f_permutation__U3583  ( .A1(SYNOPSYS_UNCONNECTED_280), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5430 ) );
  NAND2_X2 _f_permutation__U3582  ( .A1(_f_permutation__n5429 ), .A2(
        _f_permutation__n5430 ), .ZN(_f_permutation__n4579 ) );
  NAND2_X2 _f_permutation__U3581  ( .A1(_f_permutation__round_out[807]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5427 ) );
  NAND2_X2 _f_permutation__U3580  ( .A1(SYNOPSYS_UNCONNECTED_281), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5428 ) );
  NAND2_X2 _f_permutation__U3579  ( .A1(_f_permutation__n5427 ), .A2(
        _f_permutation__n5428 ), .ZN(_f_permutation__n4580 ) );
  NAND2_X2 _f_permutation__U3578  ( .A1(_f_permutation__round_out[806]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5425 ) );
  NAND2_X2 _f_permutation__U3577  ( .A1(SYNOPSYS_UNCONNECTED_282), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5426 ) );
  NAND2_X2 _f_permutation__U3576  ( .A1(_f_permutation__n5425 ), .A2(
        _f_permutation__n5426 ), .ZN(_f_permutation__n4581 ) );
  NAND2_X2 _f_permutation__U3575  ( .A1(_f_permutation__round_out[805]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5423 ) );
  NAND2_X2 _f_permutation__U3574  ( .A1(SYNOPSYS_UNCONNECTED_283), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5424 ) );
  NAND2_X2 _f_permutation__U3573  ( .A1(_f_permutation__n5423 ), .A2(
        _f_permutation__n5424 ), .ZN(_f_permutation__n4582 ) );
  NAND2_X2 _f_permutation__U3572  ( .A1(_f_permutation__round_out[804]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5421 ) );
  NAND2_X2 _f_permutation__U3571  ( .A1(SYNOPSYS_UNCONNECTED_284), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5422 ) );
  NAND2_X2 _f_permutation__U3570  ( .A1(_f_permutation__n5421 ), .A2(
        _f_permutation__n5422 ), .ZN(_f_permutation__n4583 ) );
  NAND2_X2 _f_permutation__U3569  ( .A1(_f_permutation__round_out[803]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5419 ) );
  NAND2_X2 _f_permutation__U3568  ( .A1(SYNOPSYS_UNCONNECTED_285), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5420 ) );
  NAND2_X2 _f_permutation__U3567  ( .A1(_f_permutation__n5419 ), .A2(
        _f_permutation__n5420 ), .ZN(_f_permutation__n4584 ) );
  NAND2_X2 _f_permutation__U3566  ( .A1(_f_permutation__round_out[802]), .A2(
        _f_permutation__n7122 ), .ZN(_f_permutation__n5417 ) );
  NAND2_X2 _f_permutation__U3565  ( .A1(SYNOPSYS_UNCONNECTED_286), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5418 ) );
  NAND2_X2 _f_permutation__U3564  ( .A1(_f_permutation__n5417 ), .A2(
        _f_permutation__n5418 ), .ZN(_f_permutation__n4585 ) );
  NAND2_X2 _f_permutation__U3563  ( .A1(_f_permutation__round_out[801]), .A2(
        _f_permutation__n7125 ), .ZN(_f_permutation__n5415 ) );
  NAND2_X2 _f_permutation__U3562  ( .A1(SYNOPSYS_UNCONNECTED_287), .A2(
        _f_permutation__n7238 ), .ZN(_f_permutation__n5416 ) );
  NAND2_X2 _f_permutation__U3561  ( .A1(_f_permutation__n5415 ), .A2(
        _f_permutation__n5416 ), .ZN(_f_permutation__n4586 ) );
  NAND2_X2 _f_permutation__U3560  ( .A1(_f_permutation__round_out[800]), .A2(
        _f_permutation__n7127 ), .ZN(_f_permutation__n5413 ) );
  NAND2_X2 _f_permutation__U3559  ( .A1(SYNOPSYS_UNCONNECTED_288), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5414 ) );
  NAND2_X2 _f_permutation__U3558  ( .A1(_f_permutation__n5413 ), .A2(
        _f_permutation__n5414 ), .ZN(_f_permutation__n4587 ) );
  NAND2_X2 _f_permutation__U3557  ( .A1(_f_permutation__round_out[799]), .A2(
        _f_permutation__n7139 ), .ZN(_f_permutation__n5411 ) );
  NAND2_X2 _f_permutation__U3556  ( .A1(SYNOPSYS_UNCONNECTED_289), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5412 ) );
  NAND2_X2 _f_permutation__U3555  ( .A1(_f_permutation__n5411 ), .A2(
        _f_permutation__n5412 ), .ZN(_f_permutation__n4588 ) );
  NAND2_X2 _f_permutation__U3554  ( .A1(_f_permutation__round_out[798]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5409 ) );
  NAND2_X2 _f_permutation__U3553  ( .A1(SYNOPSYS_UNCONNECTED_290), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5410 ) );
  NAND2_X2 _f_permutation__U3552  ( .A1(_f_permutation__n5409 ), .A2(
        _f_permutation__n5410 ), .ZN(_f_permutation__n4589 ) );
  NAND2_X2 _f_permutation__U3551  ( .A1(_f_permutation__round_out[797]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5407 ) );
  NAND2_X2 _f_permutation__U3550  ( .A1(SYNOPSYS_UNCONNECTED_291), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5408 ) );
  NAND2_X2 _f_permutation__U3549  ( .A1(_f_permutation__n5407 ), .A2(
        _f_permutation__n5408 ), .ZN(_f_permutation__n4590 ) );
  NAND2_X2 _f_permutation__U3548  ( .A1(_f_permutation__round_out[796]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5405 ) );
  NAND2_X2 _f_permutation__U3547  ( .A1(SYNOPSYS_UNCONNECTED_292), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5406 ) );
  NAND2_X2 _f_permutation__U3546  ( .A1(_f_permutation__n5405 ), .A2(
        _f_permutation__n5406 ), .ZN(_f_permutation__n4591 ) );
  NAND2_X2 _f_permutation__U3545  ( .A1(_f_permutation__round_out[795]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5403 ) );
  NAND2_X2 _f_permutation__U3544  ( .A1(SYNOPSYS_UNCONNECTED_293), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5404 ) );
  NAND2_X2 _f_permutation__U3543  ( .A1(_f_permutation__n5403 ), .A2(
        _f_permutation__n5404 ), .ZN(_f_permutation__n4592 ) );
  NAND2_X2 _f_permutation__U3542  ( .A1(_f_permutation__round_out[794]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5401 ) );
  NAND2_X2 _f_permutation__U3541  ( .A1(SYNOPSYS_UNCONNECTED_294), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5402 ) );
  NAND2_X2 _f_permutation__U3540  ( .A1(_f_permutation__n5401 ), .A2(
        _f_permutation__n5402 ), .ZN(_f_permutation__n4593 ) );
  NAND2_X2 _f_permutation__U3539  ( .A1(_f_permutation__round_out[793]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5399 ) );
  NAND2_X2 _f_permutation__U3538  ( .A1(SYNOPSYS_UNCONNECTED_295), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5400 ) );
  NAND2_X2 _f_permutation__U3537  ( .A1(_f_permutation__n5399 ), .A2(
        _f_permutation__n5400 ), .ZN(_f_permutation__n4594 ) );
  NAND2_X2 _f_permutation__U3536  ( .A1(_f_permutation__round_out[792]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5397 ) );
  NAND2_X2 _f_permutation__U3535  ( .A1(SYNOPSYS_UNCONNECTED_296), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5398 ) );
  NAND2_X2 _f_permutation__U3534  ( .A1(_f_permutation__n5397 ), .A2(
        _f_permutation__n5398 ), .ZN(_f_permutation__n4595 ) );
  NAND2_X2 _f_permutation__U3533  ( .A1(_f_permutation__round_out[791]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5395 ) );
  NAND2_X2 _f_permutation__U3532  ( .A1(SYNOPSYS_UNCONNECTED_297), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5396 ) );
  NAND2_X2 _f_permutation__U3531  ( .A1(_f_permutation__n5395 ), .A2(
        _f_permutation__n5396 ), .ZN(_f_permutation__n4596 ) );
  NAND2_X2 _f_permutation__U3530  ( .A1(_f_permutation__round_out[790]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5393 ) );
  NAND2_X2 _f_permutation__U3529  ( .A1(SYNOPSYS_UNCONNECTED_298), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5394 ) );
  NAND2_X2 _f_permutation__U3528  ( .A1(_f_permutation__n5393 ), .A2(
        _f_permutation__n5394 ), .ZN(_f_permutation__n4597 ) );
  NAND2_X2 _f_permutation__U3527  ( .A1(_f_permutation__round_out[789]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5391 ) );
  NAND2_X2 _f_permutation__U3526  ( .A1(SYNOPSYS_UNCONNECTED_299), .A2(
        _f_permutation__n7239 ), .ZN(_f_permutation__n5392 ) );
  NAND2_X2 _f_permutation__U3525  ( .A1(_f_permutation__n5391 ), .A2(
        _f_permutation__n5392 ), .ZN(_f_permutation__n4598 ) );
  NAND2_X2 _f_permutation__U3524  ( .A1(_f_permutation__round_out[788]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n5389 ) );
  NAND2_X2 _f_permutation__U3523  ( .A1(SYNOPSYS_UNCONNECTED_300), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n5390 ) );
  NAND2_X2 _f_permutation__U3522  ( .A1(_f_permutation__n5389 ), .A2(
        _f_permutation__n5390 ), .ZN(_f_permutation__n4599 ) );
  NAND2_X2 _f_permutation__U3521  ( .A1(_f_permutation__round_out[787]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n3786 ) );
  NAND2_X2 _f_permutation__U3520  ( .A1(SYNOPSYS_UNCONNECTED_301), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3787 ) );
  NAND2_X2 _f_permutation__U3519  ( .A1(_f_permutation__n3786 ), .A2(
        _f_permutation__n3787 ), .ZN(_f_permutation__n4600 ) );
  NAND2_X2 _f_permutation__U3518  ( .A1(_f_permutation__round_out[786]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n3784 ) );
  NAND2_X2 _f_permutation__U3517  ( .A1(SYNOPSYS_UNCONNECTED_302), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3785 ) );
  NAND2_X2 _f_permutation__U3516  ( .A1(_f_permutation__n3784 ), .A2(
        _f_permutation__n3785 ), .ZN(_f_permutation__n4601 ) );
  NAND2_X2 _f_permutation__U3515  ( .A1(_f_permutation__round_out[785]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n3782 ) );
  NAND2_X2 _f_permutation__U3514  ( .A1(SYNOPSYS_UNCONNECTED_303), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3783 ) );
  NAND2_X2 _f_permutation__U3513  ( .A1(_f_permutation__n3782 ), .A2(
        _f_permutation__n3783 ), .ZN(_f_permutation__n4602 ) );
  NAND2_X2 _f_permutation__U3512  ( .A1(_f_permutation__round_out[784]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n3780 ) );
  NAND2_X2 _f_permutation__U3511  ( .A1(SYNOPSYS_UNCONNECTED_304), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3781 ) );
  NAND2_X2 _f_permutation__U3510  ( .A1(_f_permutation__n3780 ), .A2(
        _f_permutation__n3781 ), .ZN(_f_permutation__n4603 ) );
  NAND2_X2 _f_permutation__U3509  ( .A1(_f_permutation__round_out[783]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3778 ) );
  NAND2_X2 _f_permutation__U3508  ( .A1(SYNOPSYS_UNCONNECTED_305), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3779 ) );
  NAND2_X2 _f_permutation__U3507  ( .A1(_f_permutation__n3778 ), .A2(
        _f_permutation__n3779 ), .ZN(_f_permutation__n4604 ) );
  NAND2_X2 _f_permutation__U3506  ( .A1(_f_permutation__round_out[782]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3776 ) );
  NAND2_X2 _f_permutation__U3505  ( .A1(SYNOPSYS_UNCONNECTED_306), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3777 ) );
  NAND2_X2 _f_permutation__U3504  ( .A1(_f_permutation__n3776 ), .A2(
        _f_permutation__n3777 ), .ZN(_f_permutation__n4605 ) );
  NAND2_X2 _f_permutation__U3503  ( .A1(_f_permutation__round_out[781]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3774 ) );
  NAND2_X2 _f_permutation__U3502  ( .A1(SYNOPSYS_UNCONNECTED_307), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3775 ) );
  NAND2_X2 _f_permutation__U3501  ( .A1(_f_permutation__n3774 ), .A2(
        _f_permutation__n3775 ), .ZN(_f_permutation__n4606 ) );
  NAND2_X2 _f_permutation__U3500  ( .A1(_f_permutation__round_out[780]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3772 ) );
  NAND2_X2 _f_permutation__U3499  ( .A1(SYNOPSYS_UNCONNECTED_308), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3773 ) );
  NAND2_X2 _f_permutation__U3498  ( .A1(_f_permutation__n3772 ), .A2(
        _f_permutation__n3773 ), .ZN(_f_permutation__n4607 ) );
  NAND2_X2 _f_permutation__U3497  ( .A1(_f_permutation__round_out[779]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3770 ) );
  NAND2_X2 _f_permutation__U3496  ( .A1(SYNOPSYS_UNCONNECTED_309), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3771 ) );
  NAND2_X2 _f_permutation__U3495  ( .A1(_f_permutation__n3770 ), .A2(
        _f_permutation__n3771 ), .ZN(_f_permutation__n4608 ) );
  NAND2_X2 _f_permutation__U3494  ( .A1(_f_permutation__round_out[778]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3768 ) );
  NAND2_X2 _f_permutation__U3493  ( .A1(SYNOPSYS_UNCONNECTED_310), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3769 ) );
  NAND2_X2 _f_permutation__U3492  ( .A1(_f_permutation__n3768 ), .A2(
        _f_permutation__n3769 ), .ZN(_f_permutation__n4609 ) );
  NAND2_X2 _f_permutation__U3491  ( .A1(_f_permutation__round_out[777]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3766 ) );
  NAND2_X2 _f_permutation__U3490  ( .A1(SYNOPSYS_UNCONNECTED_311), .A2(
        _f_permutation__n7240 ), .ZN(_f_permutation__n3767 ) );
  NAND2_X2 _f_permutation__U3489  ( .A1(_f_permutation__n3766 ), .A2(
        _f_permutation__n3767 ), .ZN(_f_permutation__n4610 ) );
  NAND2_X2 _f_permutation__U3488  ( .A1(_f_permutation__round_out[776]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3764 ) );
  NAND2_X2 _f_permutation__U3487  ( .A1(SYNOPSYS_UNCONNECTED_312), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3765 ) );
  NAND2_X2 _f_permutation__U3486  ( .A1(_f_permutation__n3764 ), .A2(
        _f_permutation__n3765 ), .ZN(_f_permutation__n4611 ) );
  NAND2_X2 _f_permutation__U3485  ( .A1(_f_permutation__round_out[775]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3762 ) );
  NAND2_X2 _f_permutation__U3484  ( .A1(SYNOPSYS_UNCONNECTED_313), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3763 ) );
  NAND2_X2 _f_permutation__U3483  ( .A1(_f_permutation__n3762 ), .A2(
        _f_permutation__n3763 ), .ZN(_f_permutation__n4612 ) );
  NAND2_X2 _f_permutation__U3482  ( .A1(_f_permutation__round_out[774]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3760 ) );
  NAND2_X2 _f_permutation__U3481  ( .A1(SYNOPSYS_UNCONNECTED_314), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3761 ) );
  NAND2_X2 _f_permutation__U3480  ( .A1(_f_permutation__n3760 ), .A2(
        _f_permutation__n3761 ), .ZN(_f_permutation__n4613 ) );
  NAND2_X2 _f_permutation__U3479  ( .A1(_f_permutation__round_out[773]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3758 ) );
  NAND2_X2 _f_permutation__U3478  ( .A1(SYNOPSYS_UNCONNECTED_315), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3759 ) );
  NAND2_X2 _f_permutation__U3477  ( .A1(_f_permutation__n3758 ), .A2(
        _f_permutation__n3759 ), .ZN(_f_permutation__n4614 ) );
  NAND2_X2 _f_permutation__U3476  ( .A1(_f_permutation__round_out[772]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3756 ) );
  NAND2_X2 _f_permutation__U3475  ( .A1(SYNOPSYS_UNCONNECTED_316), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3757 ) );
  NAND2_X2 _f_permutation__U3474  ( .A1(_f_permutation__n3756 ), .A2(
        _f_permutation__n3757 ), .ZN(_f_permutation__n4615 ) );
  NAND2_X2 _f_permutation__U3473  ( .A1(_f_permutation__round_out[771]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3754 ) );
  NAND2_X2 _f_permutation__U3472  ( .A1(SYNOPSYS_UNCONNECTED_317), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3755 ) );
  NAND2_X2 _f_permutation__U3471  ( .A1(_f_permutation__n3754 ), .A2(
        _f_permutation__n3755 ), .ZN(_f_permutation__n4616 ) );
  NAND2_X2 _f_permutation__U3470  ( .A1(_f_permutation__round_out[770]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3752 ) );
  NAND2_X2 _f_permutation__U3469  ( .A1(SYNOPSYS_UNCONNECTED_318), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3753 ) );
  NAND2_X2 _f_permutation__U3468  ( .A1(_f_permutation__n3752 ), .A2(
        _f_permutation__n3753 ), .ZN(_f_permutation__n4617 ) );
  NAND2_X2 _f_permutation__U3467  ( .A1(_f_permutation__round_out[769]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3750 ) );
  NAND2_X2 _f_permutation__U3466  ( .A1(SYNOPSYS_UNCONNECTED_319), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3751 ) );
  NAND2_X2 _f_permutation__U3465  ( .A1(_f_permutation__n3750 ), .A2(
        _f_permutation__n3751 ), .ZN(_f_permutation__n4618 ) );
  NAND2_X2 _f_permutation__U3464  ( .A1(_f_permutation__round_out[768]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3748 ) );
  NAND2_X2 _f_permutation__U3463  ( .A1(SYNOPSYS_UNCONNECTED_320), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3749 ) );
  NAND2_X2 _f_permutation__U3462  ( .A1(_f_permutation__n3748 ), .A2(
        _f_permutation__n3749 ), .ZN(_f_permutation__n4619 ) );
  NAND2_X2 _f_permutation__U3461  ( .A1(_f_permutation__round_out[767]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3746 ) );
  NAND2_X2 _f_permutation__U3460  ( .A1(SYNOPSYS_UNCONNECTED_321), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3747 ) );
  NAND2_X2 _f_permutation__U3459  ( .A1(_f_permutation__n3746 ), .A2(
        _f_permutation__n3747 ), .ZN(_f_permutation__n4620 ) );
  NAND2_X2 _f_permutation__U3458  ( .A1(_f_permutation__round_out[766]), .A2(
        _f_permutation__n7078 ), .ZN(_f_permutation__n3744 ) );
  NAND2_X2 _f_permutation__U3457  ( .A1(SYNOPSYS_UNCONNECTED_322), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3745 ) );
  NAND2_X2 _f_permutation__U3456  ( .A1(_f_permutation__n3744 ), .A2(
        _f_permutation__n3745 ), .ZN(_f_permutation__n4621 ) );
  NAND2_X2 _f_permutation__U3455  ( .A1(_f_permutation__round_out[765]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3742 ) );
  NAND2_X2 _f_permutation__U3454  ( .A1(SYNOPSYS_UNCONNECTED_323), .A2(
        _f_permutation__n7241 ), .ZN(_f_permutation__n3743 ) );
  NAND2_X2 _f_permutation__U3453  ( .A1(_f_permutation__n3742 ), .A2(
        _f_permutation__n3743 ), .ZN(_f_permutation__n4622 ) );
  NAND2_X2 _f_permutation__U3452  ( .A1(_f_permutation__round_out[764]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3740 ) );
  NAND2_X2 _f_permutation__U3451  ( .A1(SYNOPSYS_UNCONNECTED_324), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3741 ) );
  NAND2_X2 _f_permutation__U3450  ( .A1(_f_permutation__n3740 ), .A2(
        _f_permutation__n3741 ), .ZN(_f_permutation__n4623 ) );
  NAND2_X2 _f_permutation__U3449  ( .A1(_f_permutation__round_out[763]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3738 ) );
  NAND2_X2 _f_permutation__U3448  ( .A1(SYNOPSYS_UNCONNECTED_325), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3739 ) );
  NAND2_X2 _f_permutation__U3447  ( .A1(_f_permutation__n3738 ), .A2(
        _f_permutation__n3739 ), .ZN(_f_permutation__n4624 ) );
  NAND2_X2 _f_permutation__U3446  ( .A1(_f_permutation__round_out[762]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3736 ) );
  NAND2_X2 _f_permutation__U3445  ( .A1(SYNOPSYS_UNCONNECTED_326), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3737 ) );
  NAND2_X2 _f_permutation__U3444  ( .A1(_f_permutation__n3736 ), .A2(
        _f_permutation__n3737 ), .ZN(_f_permutation__n4625 ) );
  NAND2_X2 _f_permutation__U3443  ( .A1(_f_permutation__round_out[761]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3734 ) );
  NAND2_X2 _f_permutation__U3442  ( .A1(SYNOPSYS_UNCONNECTED_327), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3735 ) );
  NAND2_X2 _f_permutation__U3441  ( .A1(_f_permutation__n3734 ), .A2(
        _f_permutation__n3735 ), .ZN(_f_permutation__n4626 ) );
  NAND2_X2 _f_permutation__U3440  ( .A1(_f_permutation__round_out[760]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3732 ) );
  NAND2_X2 _f_permutation__U3439  ( .A1(SYNOPSYS_UNCONNECTED_328), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3733 ) );
  NAND2_X2 _f_permutation__U3438  ( .A1(_f_permutation__n3732 ), .A2(
        _f_permutation__n3733 ), .ZN(_f_permutation__n4627 ) );
  NAND2_X2 _f_permutation__U3437  ( .A1(_f_permutation__round_out[759]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3730 ) );
  NAND2_X2 _f_permutation__U3436  ( .A1(SYNOPSYS_UNCONNECTED_329), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3731 ) );
  NAND2_X2 _f_permutation__U3435  ( .A1(_f_permutation__n3730 ), .A2(
        _f_permutation__n3731 ), .ZN(_f_permutation__n4628 ) );
  NAND2_X2 _f_permutation__U3434  ( .A1(_f_permutation__round_out[758]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3728 ) );
  NAND2_X2 _f_permutation__U3433  ( .A1(SYNOPSYS_UNCONNECTED_330), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3729 ) );
  NAND2_X2 _f_permutation__U3432  ( .A1(_f_permutation__n3728 ), .A2(
        _f_permutation__n3729 ), .ZN(_f_permutation__n4629 ) );
  NAND2_X2 _f_permutation__U3431  ( .A1(_f_permutation__round_out[757]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3726 ) );
  NAND2_X2 _f_permutation__U3430  ( .A1(SYNOPSYS_UNCONNECTED_331), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3727 ) );
  NAND2_X2 _f_permutation__U3429  ( .A1(_f_permutation__n3726 ), .A2(
        _f_permutation__n3727 ), .ZN(_f_permutation__n4630 ) );
  NAND2_X2 _f_permutation__U3428  ( .A1(_f_permutation__round_out[756]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3724 ) );
  NAND2_X2 _f_permutation__U3427  ( .A1(SYNOPSYS_UNCONNECTED_332), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3725 ) );
  NAND2_X2 _f_permutation__U3426  ( .A1(_f_permutation__n3724 ), .A2(
        _f_permutation__n3725 ), .ZN(_f_permutation__n4631 ) );
  NAND2_X2 _f_permutation__U3425  ( .A1(_f_permutation__round_out[755]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3722 ) );
  NAND2_X2 _f_permutation__U3424  ( .A1(SYNOPSYS_UNCONNECTED_333), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3723 ) );
  NAND2_X2 _f_permutation__U3423  ( .A1(_f_permutation__n3722 ), .A2(
        _f_permutation__n3723 ), .ZN(_f_permutation__n4632 ) );
  NAND2_X2 _f_permutation__U3422  ( .A1(_f_permutation__round_out[754]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3720 ) );
  NAND2_X2 _f_permutation__U3421  ( .A1(SYNOPSYS_UNCONNECTED_334), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3721 ) );
  NAND2_X2 _f_permutation__U3420  ( .A1(_f_permutation__n3720 ), .A2(
        _f_permutation__n3721 ), .ZN(_f_permutation__n4633 ) );
  NAND2_X2 _f_permutation__U3419  ( .A1(_f_permutation__round_out[753]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3718 ) );
  NAND2_X2 _f_permutation__U3418  ( .A1(SYNOPSYS_UNCONNECTED_335), .A2(
        _f_permutation__n7242 ), .ZN(_f_permutation__n3719 ) );
  NAND2_X2 _f_permutation__U3417  ( .A1(_f_permutation__n3718 ), .A2(
        _f_permutation__n3719 ), .ZN(_f_permutation__n4634 ) );
  NAND2_X2 _f_permutation__U3416  ( .A1(_f_permutation__round_out[752]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3716 ) );
  NAND2_X2 _f_permutation__U3415  ( .A1(SYNOPSYS_UNCONNECTED_336), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3717 ) );
  NAND2_X2 _f_permutation__U3414  ( .A1(_f_permutation__n3716 ), .A2(
        _f_permutation__n3717 ), .ZN(_f_permutation__n4635 ) );
  NAND2_X2 _f_permutation__U3413  ( .A1(_f_permutation__round_out[751]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3714 ) );
  NAND2_X2 _f_permutation__U3412  ( .A1(SYNOPSYS_UNCONNECTED_337), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3715 ) );
  NAND2_X2 _f_permutation__U3411  ( .A1(_f_permutation__n3714 ), .A2(
        _f_permutation__n3715 ), .ZN(_f_permutation__n4636 ) );
  NAND2_X2 _f_permutation__U3410  ( .A1(_f_permutation__round_out[750]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3712 ) );
  NAND2_X2 _f_permutation__U3409  ( .A1(SYNOPSYS_UNCONNECTED_338), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3713 ) );
  NAND2_X2 _f_permutation__U3408  ( .A1(_f_permutation__n3712 ), .A2(
        _f_permutation__n3713 ), .ZN(_f_permutation__n4637 ) );
  NAND2_X2 _f_permutation__U3407  ( .A1(_f_permutation__round_out[749]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3710 ) );
  NAND2_X2 _f_permutation__U3406  ( .A1(SYNOPSYS_UNCONNECTED_339), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3711 ) );
  NAND2_X2 _f_permutation__U3405  ( .A1(_f_permutation__n3710 ), .A2(
        _f_permutation__n3711 ), .ZN(_f_permutation__n4638 ) );
  NAND2_X2 _f_permutation__U3404  ( .A1(_f_permutation__round_out[748]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3708 ) );
  NAND2_X2 _f_permutation__U3403  ( .A1(SYNOPSYS_UNCONNECTED_340), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3709 ) );
  NAND2_X2 _f_permutation__U3402  ( .A1(_f_permutation__n3708 ), .A2(
        _f_permutation__n3709 ), .ZN(_f_permutation__n4639 ) );
  NAND2_X2 _f_permutation__U3401  ( .A1(_f_permutation__round_out[747]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3706 ) );
  NAND2_X2 _f_permutation__U3400  ( .A1(SYNOPSYS_UNCONNECTED_341), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3707 ) );
  NAND2_X2 _f_permutation__U3399  ( .A1(_f_permutation__n3706 ), .A2(
        _f_permutation__n3707 ), .ZN(_f_permutation__n4640 ) );
  NAND2_X2 _f_permutation__U3398  ( .A1(_f_permutation__round_out[746]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3704 ) );
  NAND2_X2 _f_permutation__U3397  ( .A1(SYNOPSYS_UNCONNECTED_342), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3705 ) );
  NAND2_X2 _f_permutation__U3396  ( .A1(_f_permutation__n3704 ), .A2(
        _f_permutation__n3705 ), .ZN(_f_permutation__n4641 ) );
  NAND2_X2 _f_permutation__U3395  ( .A1(_f_permutation__round_out[745]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3702 ) );
  NAND2_X2 _f_permutation__U3394  ( .A1(SYNOPSYS_UNCONNECTED_343), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3703 ) );
  NAND2_X2 _f_permutation__U3393  ( .A1(_f_permutation__n3702 ), .A2(
        _f_permutation__n3703 ), .ZN(_f_permutation__n4642 ) );
  NAND2_X2 _f_permutation__U3392  ( .A1(_f_permutation__round_out[744]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3700 ) );
  NAND2_X2 _f_permutation__U3391  ( .A1(SYNOPSYS_UNCONNECTED_344), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3701 ) );
  NAND2_X2 _f_permutation__U3390  ( .A1(_f_permutation__n3700 ), .A2(
        _f_permutation__n3701 ), .ZN(_f_permutation__n4643 ) );
  NAND2_X2 _f_permutation__U3389  ( .A1(_f_permutation__round_out[743]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3698 ) );
  NAND2_X2 _f_permutation__U3388  ( .A1(SYNOPSYS_UNCONNECTED_345), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3699 ) );
  NAND2_X2 _f_permutation__U3387  ( .A1(_f_permutation__n3698 ), .A2(
        _f_permutation__n3699 ), .ZN(_f_permutation__n4644 ) );
  NAND2_X2 _f_permutation__U3386  ( .A1(_f_permutation__round_out[742]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3696 ) );
  NAND2_X2 _f_permutation__U3385  ( .A1(SYNOPSYS_UNCONNECTED_346), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3697 ) );
  NAND2_X2 _f_permutation__U3384  ( .A1(_f_permutation__n3696 ), .A2(
        _f_permutation__n3697 ), .ZN(_f_permutation__n4645 ) );
  NAND2_X2 _f_permutation__U3383  ( .A1(_f_permutation__round_out[741]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3694 ) );
  NAND2_X2 _f_permutation__U3382  ( .A1(SYNOPSYS_UNCONNECTED_347), .A2(
        _f_permutation__n7243 ), .ZN(_f_permutation__n3695 ) );
  NAND2_X2 _f_permutation__U3381  ( .A1(_f_permutation__n3694 ), .A2(
        _f_permutation__n3695 ), .ZN(_f_permutation__n4646 ) );
  NAND2_X2 _f_permutation__U3380  ( .A1(_f_permutation__round_out[740]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3692 ) );
  NAND2_X2 _f_permutation__U3379  ( .A1(SYNOPSYS_UNCONNECTED_348), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3693 ) );
  NAND2_X2 _f_permutation__U3378  ( .A1(_f_permutation__n3692 ), .A2(
        _f_permutation__n3693 ), .ZN(_f_permutation__n4647 ) );
  NAND2_X2 _f_permutation__U3377  ( .A1(_f_permutation__round_out[739]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3690 ) );
  NAND2_X2 _f_permutation__U3376  ( .A1(SYNOPSYS_UNCONNECTED_349), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3691 ) );
  NAND2_X2 _f_permutation__U3375  ( .A1(_f_permutation__n3690 ), .A2(
        _f_permutation__n3691 ), .ZN(_f_permutation__n4648 ) );
  NAND2_X2 _f_permutation__U3374  ( .A1(_f_permutation__round_out[738]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3688 ) );
  NAND2_X2 _f_permutation__U3373  ( .A1(SYNOPSYS_UNCONNECTED_350), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3689 ) );
  NAND2_X2 _f_permutation__U3372  ( .A1(_f_permutation__n3688 ), .A2(
        _f_permutation__n3689 ), .ZN(_f_permutation__n4649 ) );
  NAND2_X2 _f_permutation__U3371  ( .A1(_f_permutation__round_out[737]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3686 ) );
  NAND2_X2 _f_permutation__U3370  ( .A1(SYNOPSYS_UNCONNECTED_351), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3687 ) );
  NAND2_X2 _f_permutation__U3369  ( .A1(_f_permutation__n3686 ), .A2(
        _f_permutation__n3687 ), .ZN(_f_permutation__n4650 ) );
  NAND2_X2 _f_permutation__U3368  ( .A1(_f_permutation__round_out[736]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3684 ) );
  NAND2_X2 _f_permutation__U3367  ( .A1(SYNOPSYS_UNCONNECTED_352), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3685 ) );
  NAND2_X2 _f_permutation__U3366  ( .A1(_f_permutation__n3684 ), .A2(
        _f_permutation__n3685 ), .ZN(_f_permutation__n4651 ) );
  NAND2_X2 _f_permutation__U3365  ( .A1(_f_permutation__round_out[735]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3682 ) );
  NAND2_X2 _f_permutation__U3364  ( .A1(SYNOPSYS_UNCONNECTED_353), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3683 ) );
  NAND2_X2 _f_permutation__U3363  ( .A1(_f_permutation__n3682 ), .A2(
        _f_permutation__n3683 ), .ZN(_f_permutation__n4652 ) );
  NAND2_X2 _f_permutation__U3362  ( .A1(_f_permutation__round_out[734]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3680 ) );
  NAND2_X2 _f_permutation__U3361  ( .A1(SYNOPSYS_UNCONNECTED_354), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3681 ) );
  NAND2_X2 _f_permutation__U3360  ( .A1(_f_permutation__n3680 ), .A2(
        _f_permutation__n3681 ), .ZN(_f_permutation__n4653 ) );
  NAND2_X2 _f_permutation__U3359  ( .A1(_f_permutation__round_out[733]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3678 ) );
  NAND2_X2 _f_permutation__U3358  ( .A1(SYNOPSYS_UNCONNECTED_355), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3679 ) );
  NAND2_X2 _f_permutation__U3357  ( .A1(_f_permutation__n3678 ), .A2(
        _f_permutation__n3679 ), .ZN(_f_permutation__n4654 ) );
  NAND2_X2 _f_permutation__U3356  ( .A1(_f_permutation__round_out[732]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3676 ) );
  NAND2_X2 _f_permutation__U3355  ( .A1(SYNOPSYS_UNCONNECTED_356), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3677 ) );
  NAND2_X2 _f_permutation__U3354  ( .A1(_f_permutation__n3676 ), .A2(
        _f_permutation__n3677 ), .ZN(_f_permutation__n4655 ) );
  NAND2_X2 _f_permutation__U3353  ( .A1(_f_permutation__round_out[731]), .A2(
        _f_permutation__n7076 ), .ZN(_f_permutation__n3674 ) );
  NAND2_X2 _f_permutation__U3352  ( .A1(SYNOPSYS_UNCONNECTED_357), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3675 ) );
  NAND2_X2 _f_permutation__U3351  ( .A1(_f_permutation__n3674 ), .A2(
        _f_permutation__n3675 ), .ZN(_f_permutation__n4656 ) );
  NAND2_X2 _f_permutation__U3350  ( .A1(_f_permutation__round_out[730]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3672 ) );
  NAND2_X2 _f_permutation__U3349  ( .A1(SYNOPSYS_UNCONNECTED_358), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3673 ) );
  NAND2_X2 _f_permutation__U3348  ( .A1(_f_permutation__n3672 ), .A2(
        _f_permutation__n3673 ), .ZN(_f_permutation__n4657 ) );
  NAND2_X2 _f_permutation__U3347  ( .A1(_f_permutation__round_out[729]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3670 ) );
  NAND2_X2 _f_permutation__U3346  ( .A1(SYNOPSYS_UNCONNECTED_359), .A2(
        _f_permutation__n7244 ), .ZN(_f_permutation__n3671 ) );
  NAND2_X2 _f_permutation__U3345  ( .A1(_f_permutation__n3670 ), .A2(
        _f_permutation__n3671 ), .ZN(_f_permutation__n4658 ) );
  NAND2_X2 _f_permutation__U3344  ( .A1(_f_permutation__round_out[728]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3668 ) );
  NAND2_X2 _f_permutation__U3343  ( .A1(SYNOPSYS_UNCONNECTED_360), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3669 ) );
  NAND2_X2 _f_permutation__U3342  ( .A1(_f_permutation__n3668 ), .A2(
        _f_permutation__n3669 ), .ZN(_f_permutation__n4659 ) );
  NAND2_X2 _f_permutation__U3341  ( .A1(_f_permutation__round_out[727]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3666 ) );
  NAND2_X2 _f_permutation__U3340  ( .A1(SYNOPSYS_UNCONNECTED_361), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3667 ) );
  NAND2_X2 _f_permutation__U3339  ( .A1(_f_permutation__n3666 ), .A2(
        _f_permutation__n3667 ), .ZN(_f_permutation__n4660 ) );
  NAND2_X2 _f_permutation__U3338  ( .A1(_f_permutation__round_out[726]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3664 ) );
  NAND2_X2 _f_permutation__U3337  ( .A1(SYNOPSYS_UNCONNECTED_362), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3665 ) );
  NAND2_X2 _f_permutation__U3336  ( .A1(_f_permutation__n3664 ), .A2(
        _f_permutation__n3665 ), .ZN(_f_permutation__n4661 ) );
  NAND2_X2 _f_permutation__U3335  ( .A1(_f_permutation__round_out[725]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3662 ) );
  NAND2_X2 _f_permutation__U3334  ( .A1(SYNOPSYS_UNCONNECTED_363), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3663 ) );
  NAND2_X2 _f_permutation__U3333  ( .A1(_f_permutation__n3662 ), .A2(
        _f_permutation__n3663 ), .ZN(_f_permutation__n4662 ) );
  NAND2_X2 _f_permutation__U3332  ( .A1(_f_permutation__round_out[724]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3660 ) );
  NAND2_X2 _f_permutation__U3331  ( .A1(SYNOPSYS_UNCONNECTED_364), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3661 ) );
  NAND2_X2 _f_permutation__U3330  ( .A1(_f_permutation__n3660 ), .A2(
        _f_permutation__n3661 ), .ZN(_f_permutation__n4663 ) );
  NAND2_X2 _f_permutation__U3329  ( .A1(_f_permutation__round_out[723]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3658 ) );
  NAND2_X2 _f_permutation__U3328  ( .A1(SYNOPSYS_UNCONNECTED_365), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3659 ) );
  NAND2_X2 _f_permutation__U3327  ( .A1(_f_permutation__n3658 ), .A2(
        _f_permutation__n3659 ), .ZN(_f_permutation__n4664 ) );
  NAND2_X2 _f_permutation__U3326  ( .A1(_f_permutation__round_out[722]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3656 ) );
  NAND2_X2 _f_permutation__U3325  ( .A1(SYNOPSYS_UNCONNECTED_366), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3657 ) );
  NAND2_X2 _f_permutation__U3324  ( .A1(_f_permutation__n3656 ), .A2(
        _f_permutation__n3657 ), .ZN(_f_permutation__n4665 ) );
  NAND2_X2 _f_permutation__U3323  ( .A1(_f_permutation__round_out[721]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3654 ) );
  NAND2_X2 _f_permutation__U3322  ( .A1(SYNOPSYS_UNCONNECTED_367), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3655 ) );
  NAND2_X2 _f_permutation__U3321  ( .A1(_f_permutation__n3654 ), .A2(
        _f_permutation__n3655 ), .ZN(_f_permutation__n4666 ) );
  NAND2_X2 _f_permutation__U3320  ( .A1(_f_permutation__round_out[720]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3652 ) );
  NAND2_X2 _f_permutation__U3319  ( .A1(SYNOPSYS_UNCONNECTED_368), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3653 ) );
  NAND2_X2 _f_permutation__U3318  ( .A1(_f_permutation__n3652 ), .A2(
        _f_permutation__n3653 ), .ZN(_f_permutation__n4667 ) );
  NAND2_X2 _f_permutation__U3317  ( .A1(_f_permutation__round_out[719]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3650 ) );
  NAND2_X2 _f_permutation__U3316  ( .A1(SYNOPSYS_UNCONNECTED_369), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3651 ) );
  NAND2_X2 _f_permutation__U3315  ( .A1(_f_permutation__n3650 ), .A2(
        _f_permutation__n3651 ), .ZN(_f_permutation__n4668 ) );
  NAND2_X2 _f_permutation__U3314  ( .A1(_f_permutation__round_out[718]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3648 ) );
  NAND2_X2 _f_permutation__U3313  ( .A1(SYNOPSYS_UNCONNECTED_370), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3649 ) );
  NAND2_X2 _f_permutation__U3312  ( .A1(_f_permutation__n3648 ), .A2(
        _f_permutation__n3649 ), .ZN(_f_permutation__n4669 ) );
  NAND2_X2 _f_permutation__U3311  ( .A1(_f_permutation__round_out[717]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3646 ) );
  NAND2_X2 _f_permutation__U3310  ( .A1(SYNOPSYS_UNCONNECTED_371), .A2(
        _f_permutation__n7245 ), .ZN(_f_permutation__n3647 ) );
  NAND2_X2 _f_permutation__U3309  ( .A1(_f_permutation__n3646 ), .A2(
        _f_permutation__n3647 ), .ZN(_f_permutation__n4670 ) );
  NAND2_X2 _f_permutation__U3308  ( .A1(_f_permutation__round_out[716]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3644 ) );
  NAND2_X2 _f_permutation__U3307  ( .A1(SYNOPSYS_UNCONNECTED_372), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3645 ) );
  NAND2_X2 _f_permutation__U3306  ( .A1(_f_permutation__n3644 ), .A2(
        _f_permutation__n3645 ), .ZN(_f_permutation__n4671 ) );
  NAND2_X2 _f_permutation__U3305  ( .A1(_f_permutation__round_out[715]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3642 ) );
  NAND2_X2 _f_permutation__U3304  ( .A1(SYNOPSYS_UNCONNECTED_373), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3643 ) );
  NAND2_X2 _f_permutation__U3303  ( .A1(_f_permutation__n3642 ), .A2(
        _f_permutation__n3643 ), .ZN(_f_permutation__n4672 ) );
  NAND2_X2 _f_permutation__U3302  ( .A1(_f_permutation__round_out[714]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3640 ) );
  NAND2_X2 _f_permutation__U3301  ( .A1(SYNOPSYS_UNCONNECTED_374), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3641 ) );
  NAND2_X2 _f_permutation__U3300  ( .A1(_f_permutation__n3640 ), .A2(
        _f_permutation__n3641 ), .ZN(_f_permutation__n4673 ) );
  NAND2_X2 _f_permutation__U3299  ( .A1(_f_permutation__round_out[713]), .A2(
        _f_permutation__n7075 ), .ZN(_f_permutation__n3638 ) );
  NAND2_X2 _f_permutation__U3298  ( .A1(SYNOPSYS_UNCONNECTED_375), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3639 ) );
  NAND2_X2 _f_permutation__U3297  ( .A1(_f_permutation__n3638 ), .A2(
        _f_permutation__n3639 ), .ZN(_f_permutation__n4674 ) );
  NAND2_X2 _f_permutation__U3296  ( .A1(_f_permutation__round_out[712]), .A2(
        _f_permutation__n7148 ), .ZN(_f_permutation__n3636 ) );
  NAND2_X2 _f_permutation__U3295  ( .A1(SYNOPSYS_UNCONNECTED_376), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3637 ) );
  NAND2_X2 _f_permutation__U3294  ( .A1(_f_permutation__n3636 ), .A2(
        _f_permutation__n3637 ), .ZN(_f_permutation__n4675 ) );
  NAND2_X2 _f_permutation__U3293  ( .A1(_f_permutation__round_out[711]), .A2(
        _f_permutation__n7147 ), .ZN(_f_permutation__n3634 ) );
  NAND2_X2 _f_permutation__U3292  ( .A1(SYNOPSYS_UNCONNECTED_377), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3635 ) );
  NAND2_X2 _f_permutation__U3291  ( .A1(_f_permutation__n3634 ), .A2(
        _f_permutation__n3635 ), .ZN(_f_permutation__n4676 ) );
  NAND2_X2 _f_permutation__U3290  ( .A1(_f_permutation__round_out[710]), .A2(
        _f_permutation__n7152 ), .ZN(_f_permutation__n3632 ) );
  NAND2_X2 _f_permutation__U3289  ( .A1(SYNOPSYS_UNCONNECTED_378), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3633 ) );
  NAND2_X2 _f_permutation__U3288  ( .A1(_f_permutation__n3632 ), .A2(
        _f_permutation__n3633 ), .ZN(_f_permutation__n4677 ) );
  NAND2_X2 _f_permutation__U3287  ( .A1(_f_permutation__round_out[709]), .A2(
        _f_permutation__n7151 ), .ZN(_f_permutation__n3630 ) );
  NAND2_X2 _f_permutation__U3286  ( .A1(SYNOPSYS_UNCONNECTED_379), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3631 ) );
  NAND2_X2 _f_permutation__U3285  ( .A1(_f_permutation__n3630 ), .A2(
        _f_permutation__n3631 ), .ZN(_f_permutation__n4678 ) );
  NAND2_X2 _f_permutation__U3284  ( .A1(_f_permutation__round_out[708]), .A2(
        _f_permutation__n7150 ), .ZN(_f_permutation__n3628 ) );
  NAND2_X2 _f_permutation__U3283  ( .A1(SYNOPSYS_UNCONNECTED_380), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3629 ) );
  NAND2_X2 _f_permutation__U3282  ( .A1(_f_permutation__n3628 ), .A2(
        _f_permutation__n3629 ), .ZN(_f_permutation__n4679 ) );
  NAND2_X2 _f_permutation__U3281  ( .A1(_f_permutation__round_out[707]), .A2(
        _f_permutation__n7146 ), .ZN(_f_permutation__n3626 ) );
  NAND2_X2 _f_permutation__U3280  ( .A1(SYNOPSYS_UNCONNECTED_381), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3627 ) );
  NAND2_X2 _f_permutation__U3279  ( .A1(_f_permutation__n3626 ), .A2(
        _f_permutation__n3627 ), .ZN(_f_permutation__n4680 ) );
  NAND2_X2 _f_permutation__U3278  ( .A1(_f_permutation__round_out[706]), .A2(
        _f_permutation__n7145 ), .ZN(_f_permutation__n3624 ) );
  NAND2_X2 _f_permutation__U3277  ( .A1(SYNOPSYS_UNCONNECTED_382), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3625 ) );
  NAND2_X2 _f_permutation__U3276  ( .A1(_f_permutation__n3624 ), .A2(
        _f_permutation__n3625 ), .ZN(_f_permutation__n4681 ) );
  NAND2_X2 _f_permutation__U3275  ( .A1(_f_permutation__round_out[705]), .A2(
        _f_permutation__n7144 ), .ZN(_f_permutation__n3622 ) );
  NAND2_X2 _f_permutation__U3274  ( .A1(SYNOPSYS_UNCONNECTED_383), .A2(
        _f_permutation__n7246 ), .ZN(_f_permutation__n3623 ) );
  NAND2_X2 _f_permutation__U3273  ( .A1(_f_permutation__n3622 ), .A2(
        _f_permutation__n3623 ), .ZN(_f_permutation__n4682 ) );
  NAND2_X2 _f_permutation__U3272  ( .A1(_f_permutation__round_out[704]), .A2(
        _f_permutation__n7143 ), .ZN(_f_permutation__n3620 ) );
  NAND2_X2 _f_permutation__U3271  ( .A1(SYNOPSYS_UNCONNECTED_384), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3621 ) );
  NAND2_X2 _f_permutation__U3270  ( .A1(_f_permutation__n3620 ), .A2(
        _f_permutation__n3621 ), .ZN(_f_permutation__n4683 ) );
  NAND2_X2 _f_permutation__U3269  ( .A1(_f_permutation__round_out[703]), .A2(
        _f_permutation__n7163 ), .ZN(_f_permutation__n3618 ) );
  NAND2_X2 _f_permutation__U3268  ( .A1(SYNOPSYS_UNCONNECTED_385), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3619 ) );
  NAND2_X2 _f_permutation__U3267  ( .A1(_f_permutation__n3618 ), .A2(
        _f_permutation__n3619 ), .ZN(_f_permutation__n4684 ) );
  NAND2_X2 _f_permutation__U3266  ( .A1(_f_permutation__round_out[702]), .A2(
        _f_permutation__n7162 ), .ZN(_f_permutation__n3616 ) );
  NAND2_X2 _f_permutation__U3265  ( .A1(SYNOPSYS_UNCONNECTED_386), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3617 ) );
  NAND2_X2 _f_permutation__U3264  ( .A1(_f_permutation__n3616 ), .A2(
        _f_permutation__n3617 ), .ZN(_f_permutation__n4685 ) );
  NAND2_X2 _f_permutation__U3263  ( .A1(_f_permutation__round_out[701]), .A2(
        _f_permutation__n7167 ), .ZN(_f_permutation__n3614 ) );
  NAND2_X2 _f_permutation__U3262  ( .A1(SYNOPSYS_UNCONNECTED_387), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3615 ) );
  NAND2_X2 _f_permutation__U3261  ( .A1(_f_permutation__n3614 ), .A2(
        _f_permutation__n3615 ), .ZN(_f_permutation__n4686 ) );
  NAND2_X2 _f_permutation__U3260  ( .A1(_f_permutation__round_out[700]), .A2(
        _f_permutation__n7166 ), .ZN(_f_permutation__n3612 ) );
  NAND2_X2 _f_permutation__U3259  ( .A1(SYNOPSYS_UNCONNECTED_388), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3613 ) );
  NAND2_X2 _f_permutation__U3258  ( .A1(_f_permutation__n3612 ), .A2(
        _f_permutation__n3613 ), .ZN(_f_permutation__n4687 ) );
  NAND2_X2 _f_permutation__U3257  ( .A1(_f_permutation__round_out[699]), .A2(
        _f_permutation__n7077 ), .ZN(_f_permutation__n3610 ) );
  NAND2_X2 _f_permutation__U3256  ( .A1(SYNOPSYS_UNCONNECTED_389), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3611 ) );
  NAND2_X2 _f_permutation__U3255  ( .A1(_f_permutation__n3610 ), .A2(
        _f_permutation__n3611 ), .ZN(_f_permutation__n4688 ) );
  NAND2_X2 _f_permutation__U3254  ( .A1(_f_permutation__round_out[698]), .A2(
        _f_permutation__n7142 ), .ZN(_f_permutation__n3608 ) );
  NAND2_X2 _f_permutation__U3253  ( .A1(SYNOPSYS_UNCONNECTED_390), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3609 ) );
  NAND2_X2 _f_permutation__U3252  ( .A1(_f_permutation__n3608 ), .A2(
        _f_permutation__n3609 ), .ZN(_f_permutation__n4689 ) );
  NAND2_X2 _f_permutation__U3251  ( .A1(_f_permutation__round_out[697]), .A2(
        _f_permutation__n7161 ), .ZN(_f_permutation__n3606 ) );
  NAND2_X2 _f_permutation__U3250  ( .A1(SYNOPSYS_UNCONNECTED_391), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3607 ) );
  NAND2_X2 _f_permutation__U3249  ( .A1(_f_permutation__n3606 ), .A2(
        _f_permutation__n3607 ), .ZN(_f_permutation__n4690 ) );
  NAND2_X2 _f_permutation__U3248  ( .A1(_f_permutation__round_out[696]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n3604 ) );
  NAND2_X2 _f_permutation__U3247  ( .A1(SYNOPSYS_UNCONNECTED_392), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3605 ) );
  NAND2_X2 _f_permutation__U3246  ( .A1(_f_permutation__n3604 ), .A2(
        _f_permutation__n3605 ), .ZN(_f_permutation__n4691 ) );
  NAND2_X2 _f_permutation__U3245  ( .A1(_f_permutation__round_out[695]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n3602 ) );
  NAND2_X2 _f_permutation__U3244  ( .A1(SYNOPSYS_UNCONNECTED_393), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3603 ) );
  NAND2_X2 _f_permutation__U3243  ( .A1(_f_permutation__n3602 ), .A2(
        _f_permutation__n3603 ), .ZN(_f_permutation__n4692 ) );
  NAND2_X2 _f_permutation__U3242  ( .A1(_f_permutation__round_out[694]), .A2(
        _f_permutation__n7168 ), .ZN(_f_permutation__n3600 ) );
  NAND2_X2 _f_permutation__U3241  ( .A1(SYNOPSYS_UNCONNECTED_394), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3601 ) );
  NAND2_X2 _f_permutation__U3240  ( .A1(_f_permutation__n3600 ), .A2(
        _f_permutation__n3601 ), .ZN(_f_permutation__n4693 ) );
  NAND2_X2 _f_permutation__U3239  ( .A1(_f_permutation__round_out[693]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n3598 ) );
  NAND2_X2 _f_permutation__U3238  ( .A1(SYNOPSYS_UNCONNECTED_395), .A2(
        _f_permutation__n7247 ), .ZN(_f_permutation__n3599 ) );
  NAND2_X2 _f_permutation__U3237  ( .A1(_f_permutation__n3598 ), .A2(
        _f_permutation__n3599 ), .ZN(_f_permutation__n4694 ) );
  NAND2_X2 _f_permutation__U3236  ( .A1(_f_permutation__round_out[692]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3596 ) );
  NAND2_X2 _f_permutation__U3235  ( .A1(SYNOPSYS_UNCONNECTED_396), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3597 ) );
  NAND2_X2 _f_permutation__U3234  ( .A1(_f_permutation__n3596 ), .A2(
        _f_permutation__n3597 ), .ZN(_f_permutation__n4695 ) );
  NAND2_X2 _f_permutation__U3233  ( .A1(_f_permutation__round_out[691]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3594 ) );
  NAND2_X2 _f_permutation__U3232  ( .A1(SYNOPSYS_UNCONNECTED_397), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3595 ) );
  NAND2_X2 _f_permutation__U3231  ( .A1(_f_permutation__n3594 ), .A2(
        _f_permutation__n3595 ), .ZN(_f_permutation__n4696 ) );
  NAND2_X2 _f_permutation__U3230  ( .A1(_f_permutation__round_out[690]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3592 ) );
  NAND2_X2 _f_permutation__U3229  ( .A1(SYNOPSYS_UNCONNECTED_398), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3593 ) );
  NAND2_X2 _f_permutation__U3228  ( .A1(_f_permutation__n3592 ), .A2(
        _f_permutation__n3593 ), .ZN(_f_permutation__n4697 ) );
  NAND2_X2 _f_permutation__U3227  ( .A1(_f_permutation__round_out[689]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3590 ) );
  NAND2_X2 _f_permutation__U3226  ( .A1(SYNOPSYS_UNCONNECTED_399), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3591 ) );
  NAND2_X2 _f_permutation__U3225  ( .A1(_f_permutation__n3590 ), .A2(
        _f_permutation__n3591 ), .ZN(_f_permutation__n4698 ) );
  NAND2_X2 _f_permutation__U3224  ( .A1(_f_permutation__round_out[688]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3588 ) );
  NAND2_X2 _f_permutation__U3223  ( .A1(SYNOPSYS_UNCONNECTED_400), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3589 ) );
  NAND2_X2 _f_permutation__U3222  ( .A1(_f_permutation__n3588 ), .A2(
        _f_permutation__n3589 ), .ZN(_f_permutation__n4699 ) );
  NAND2_X2 _f_permutation__U3221  ( .A1(_f_permutation__round_out[687]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3586 ) );
  NAND2_X2 _f_permutation__U3220  ( .A1(SYNOPSYS_UNCONNECTED_401), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3587 ) );
  NAND2_X2 _f_permutation__U3219  ( .A1(_f_permutation__n3586 ), .A2(
        _f_permutation__n3587 ), .ZN(_f_permutation__n4700 ) );
  NAND2_X2 _f_permutation__U3218  ( .A1(_f_permutation__round_out[686]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3584 ) );
  NAND2_X2 _f_permutation__U3217  ( .A1(SYNOPSYS_UNCONNECTED_402), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3585 ) );
  NAND2_X2 _f_permutation__U3216  ( .A1(_f_permutation__n3584 ), .A2(
        _f_permutation__n3585 ), .ZN(_f_permutation__n4701 ) );
  NAND2_X2 _f_permutation__U3215  ( .A1(_f_permutation__round_out[685]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3582 ) );
  NAND2_X2 _f_permutation__U3214  ( .A1(SYNOPSYS_UNCONNECTED_403), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3583 ) );
  NAND2_X2 _f_permutation__U3213  ( .A1(_f_permutation__n3582 ), .A2(
        _f_permutation__n3583 ), .ZN(_f_permutation__n4702 ) );
  NAND2_X2 _f_permutation__U3212  ( .A1(_f_permutation__round_out[684]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3580 ) );
  NAND2_X2 _f_permutation__U3211  ( .A1(SYNOPSYS_UNCONNECTED_404), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3581 ) );
  NAND2_X2 _f_permutation__U3210  ( .A1(_f_permutation__n3580 ), .A2(
        _f_permutation__n3581 ), .ZN(_f_permutation__n4703 ) );
  NAND2_X2 _f_permutation__U3209  ( .A1(_f_permutation__round_out[683]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3578 ) );
  NAND2_X2 _f_permutation__U3208  ( .A1(SYNOPSYS_UNCONNECTED_405), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3579 ) );
  NAND2_X2 _f_permutation__U3207  ( .A1(_f_permutation__n3578 ), .A2(
        _f_permutation__n3579 ), .ZN(_f_permutation__n4704 ) );
  NAND2_X2 _f_permutation__U3206  ( .A1(_f_permutation__round_out[682]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3576 ) );
  NAND2_X2 _f_permutation__U3205  ( .A1(SYNOPSYS_UNCONNECTED_406), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3577 ) );
  NAND2_X2 _f_permutation__U3204  ( .A1(_f_permutation__n3576 ), .A2(
        _f_permutation__n3577 ), .ZN(_f_permutation__n4705 ) );
  NAND2_X2 _f_permutation__U3203  ( .A1(_f_permutation__round_out[681]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3574 ) );
  NAND2_X2 _f_permutation__U3202  ( .A1(SYNOPSYS_UNCONNECTED_407), .A2(
        _f_permutation__n7248 ), .ZN(_f_permutation__n3575 ) );
  NAND2_X2 _f_permutation__U3201  ( .A1(_f_permutation__n3574 ), .A2(
        _f_permutation__n3575 ), .ZN(_f_permutation__n4706 ) );
  NAND2_X2 _f_permutation__U3200  ( .A1(_f_permutation__round_out[680]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3572 ) );
  NAND2_X2 _f_permutation__U3199  ( .A1(SYNOPSYS_UNCONNECTED_408), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3573 ) );
  NAND2_X2 _f_permutation__U3198  ( .A1(_f_permutation__n3572 ), .A2(
        _f_permutation__n3573 ), .ZN(_f_permutation__n4707 ) );
  NAND2_X2 _f_permutation__U3197  ( .A1(_f_permutation__round_out[679]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3570 ) );
  NAND2_X2 _f_permutation__U3196  ( .A1(SYNOPSYS_UNCONNECTED_409), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3571 ) );
  NAND2_X2 _f_permutation__U3195  ( .A1(_f_permutation__n3570 ), .A2(
        _f_permutation__n3571 ), .ZN(_f_permutation__n4708 ) );
  NAND2_X2 _f_permutation__U3194  ( .A1(_f_permutation__round_out[678]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3568 ) );
  NAND2_X2 _f_permutation__U3193  ( .A1(SYNOPSYS_UNCONNECTED_410), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3569 ) );
  NAND2_X2 _f_permutation__U3192  ( .A1(_f_permutation__n3568 ), .A2(
        _f_permutation__n3569 ), .ZN(_f_permutation__n4709 ) );
  NAND2_X2 _f_permutation__U3191  ( .A1(_f_permutation__round_out[677]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3566 ) );
  NAND2_X2 _f_permutation__U3190  ( .A1(SYNOPSYS_UNCONNECTED_411), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3567 ) );
  NAND2_X2 _f_permutation__U3189  ( .A1(_f_permutation__n3566 ), .A2(
        _f_permutation__n3567 ), .ZN(_f_permutation__n4710 ) );
  NAND2_X2 _f_permutation__U3188  ( .A1(_f_permutation__round_out[676]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3564 ) );
  NAND2_X2 _f_permutation__U3187  ( .A1(SYNOPSYS_UNCONNECTED_412), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3565 ) );
  NAND2_X2 _f_permutation__U3186  ( .A1(_f_permutation__n3564 ), .A2(
        _f_permutation__n3565 ), .ZN(_f_permutation__n4711 ) );
  NAND2_X2 _f_permutation__U3185  ( .A1(_f_permutation__round_out[675]), .A2(
        _f_permutation__n7084 ), .ZN(_f_permutation__n3562 ) );
  NAND2_X2 _f_permutation__U3184  ( .A1(SYNOPSYS_UNCONNECTED_413), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3563 ) );
  NAND2_X2 _f_permutation__U3183  ( .A1(_f_permutation__n3562 ), .A2(
        _f_permutation__n3563 ), .ZN(_f_permutation__n4712 ) );
  NAND2_X2 _f_permutation__U3182  ( .A1(_f_permutation__round_out[674]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3560 ) );
  NAND2_X2 _f_permutation__U3181  ( .A1(SYNOPSYS_UNCONNECTED_414), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3561 ) );
  NAND2_X2 _f_permutation__U3180  ( .A1(_f_permutation__n3560 ), .A2(
        _f_permutation__n3561 ), .ZN(_f_permutation__n4713 ) );
  NAND2_X2 _f_permutation__U3179  ( .A1(_f_permutation__round_out[673]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3558 ) );
  NAND2_X2 _f_permutation__U3178  ( .A1(SYNOPSYS_UNCONNECTED_415), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3559 ) );
  NAND2_X2 _f_permutation__U3177  ( .A1(_f_permutation__n3558 ), .A2(
        _f_permutation__n3559 ), .ZN(_f_permutation__n4714 ) );
  NAND2_X2 _f_permutation__U3176  ( .A1(_f_permutation__round_out[672]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3556 ) );
  NAND2_X2 _f_permutation__U3175  ( .A1(SYNOPSYS_UNCONNECTED_416), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3557 ) );
  NAND2_X2 _f_permutation__U3174  ( .A1(_f_permutation__n3556 ), .A2(
        _f_permutation__n3557 ), .ZN(_f_permutation__n4715 ) );
  NAND2_X2 _f_permutation__U3173  ( .A1(_f_permutation__round_out[671]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3554 ) );
  NAND2_X2 _f_permutation__U3172  ( .A1(SYNOPSYS_UNCONNECTED_417), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3555 ) );
  NAND2_X2 _f_permutation__U3171  ( .A1(_f_permutation__n3554 ), .A2(
        _f_permutation__n3555 ), .ZN(_f_permutation__n4716 ) );
  NAND2_X2 _f_permutation__U3170  ( .A1(_f_permutation__round_out[670]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3552 ) );
  NAND2_X2 _f_permutation__U3169  ( .A1(SYNOPSYS_UNCONNECTED_418), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3553 ) );
  NAND2_X2 _f_permutation__U3168  ( .A1(_f_permutation__n3552 ), .A2(
        _f_permutation__n3553 ), .ZN(_f_permutation__n4717 ) );
  NAND2_X2 _f_permutation__U3167  ( .A1(_f_permutation__round_out[669]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3550 ) );
  NAND2_X2 _f_permutation__U3166  ( .A1(SYNOPSYS_UNCONNECTED_419), .A2(
        _f_permutation__n7249 ), .ZN(_f_permutation__n3551 ) );
  NAND2_X2 _f_permutation__U3165  ( .A1(_f_permutation__n3550 ), .A2(
        _f_permutation__n3551 ), .ZN(_f_permutation__n4718 ) );
  NAND2_X2 _f_permutation__U3164  ( .A1(_f_permutation__round_out[668]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3548 ) );
  NAND2_X2 _f_permutation__U3163  ( .A1(SYNOPSYS_UNCONNECTED_420), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3549 ) );
  NAND2_X2 _f_permutation__U3162  ( .A1(_f_permutation__n3548 ), .A2(
        _f_permutation__n3549 ), .ZN(_f_permutation__n4719 ) );
  NAND2_X2 _f_permutation__U3161  ( .A1(_f_permutation__round_out[667]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3546 ) );
  NAND2_X2 _f_permutation__U3160  ( .A1(SYNOPSYS_UNCONNECTED_421), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3547 ) );
  NAND2_X2 _f_permutation__U3159  ( .A1(_f_permutation__n3546 ), .A2(
        _f_permutation__n3547 ), .ZN(_f_permutation__n4720 ) );
  NAND2_X2 _f_permutation__U3158  ( .A1(_f_permutation__round_out[666]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3544 ) );
  NAND2_X2 _f_permutation__U3157  ( .A1(SYNOPSYS_UNCONNECTED_422), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3545 ) );
  NAND2_X2 _f_permutation__U3156  ( .A1(_f_permutation__n3544 ), .A2(
        _f_permutation__n3545 ), .ZN(_f_permutation__n4721 ) );
  NAND2_X2 _f_permutation__U3155  ( .A1(_f_permutation__round_out[665]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3542 ) );
  NAND2_X2 _f_permutation__U3154  ( .A1(SYNOPSYS_UNCONNECTED_423), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3543 ) );
  NAND2_X2 _f_permutation__U3153  ( .A1(_f_permutation__n3542 ), .A2(
        _f_permutation__n3543 ), .ZN(_f_permutation__n4722 ) );
  NAND2_X2 _f_permutation__U3152  ( .A1(_f_permutation__round_out[664]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3540 ) );
  NAND2_X2 _f_permutation__U3151  ( .A1(SYNOPSYS_UNCONNECTED_424), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3541 ) );
  NAND2_X2 _f_permutation__U3150  ( .A1(_f_permutation__n3540 ), .A2(
        _f_permutation__n3541 ), .ZN(_f_permutation__n4723 ) );
  NAND2_X2 _f_permutation__U3149  ( .A1(_f_permutation__round_out[663]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3538 ) );
  NAND2_X2 _f_permutation__U3148  ( .A1(SYNOPSYS_UNCONNECTED_425), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3539 ) );
  NAND2_X2 _f_permutation__U3147  ( .A1(_f_permutation__n3538 ), .A2(
        _f_permutation__n3539 ), .ZN(_f_permutation__n4724 ) );
  NAND2_X2 _f_permutation__U3146  ( .A1(_f_permutation__round_out[662]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3536 ) );
  NAND2_X2 _f_permutation__U3145  ( .A1(SYNOPSYS_UNCONNECTED_426), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3537 ) );
  NAND2_X2 _f_permutation__U3144  ( .A1(_f_permutation__n3536 ), .A2(
        _f_permutation__n3537 ), .ZN(_f_permutation__n4725 ) );
  NAND2_X2 _f_permutation__U3143  ( .A1(_f_permutation__round_out[661]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3534 ) );
  NAND2_X2 _f_permutation__U3142  ( .A1(SYNOPSYS_UNCONNECTED_427), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3535 ) );
  NAND2_X2 _f_permutation__U3141  ( .A1(_f_permutation__n3534 ), .A2(
        _f_permutation__n3535 ), .ZN(_f_permutation__n4726 ) );
  NAND2_X2 _f_permutation__U3140  ( .A1(_f_permutation__round_out[660]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3532 ) );
  NAND2_X2 _f_permutation__U3139  ( .A1(SYNOPSYS_UNCONNECTED_428), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3533 ) );
  NAND2_X2 _f_permutation__U3138  ( .A1(_f_permutation__n3532 ), .A2(
        _f_permutation__n3533 ), .ZN(_f_permutation__n4727 ) );
  NAND2_X2 _f_permutation__U3137  ( .A1(_f_permutation__round_out[659]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3530 ) );
  NAND2_X2 _f_permutation__U3136  ( .A1(SYNOPSYS_UNCONNECTED_429), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3531 ) );
  NAND2_X2 _f_permutation__U3135  ( .A1(_f_permutation__n3530 ), .A2(
        _f_permutation__n3531 ), .ZN(_f_permutation__n4728 ) );
  NAND2_X2 _f_permutation__U3134  ( .A1(_f_permutation__round_out[658]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3528 ) );
  NAND2_X2 _f_permutation__U3133  ( .A1(SYNOPSYS_UNCONNECTED_430), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3529 ) );
  NAND2_X2 _f_permutation__U3132  ( .A1(_f_permutation__n3528 ), .A2(
        _f_permutation__n3529 ), .ZN(_f_permutation__n4729 ) );
  NAND2_X2 _f_permutation__U3131  ( .A1(_f_permutation__round_out[657]), .A2(
        _f_permutation__n7083 ), .ZN(_f_permutation__n3526 ) );
  NAND2_X2 _f_permutation__U3130  ( .A1(SYNOPSYS_UNCONNECTED_431), .A2(
        _f_permutation__n7250 ), .ZN(_f_permutation__n3527 ) );
  NAND2_X2 _f_permutation__U3129  ( .A1(_f_permutation__n3526 ), .A2(
        _f_permutation__n3527 ), .ZN(_f_permutation__n4730 ) );
  NAND2_X2 _f_permutation__U3128  ( .A1(_f_permutation__round_out[656]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3524 ) );
  NAND2_X2 _f_permutation__U3127  ( .A1(SYNOPSYS_UNCONNECTED_432), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3525 ) );
  NAND2_X2 _f_permutation__U3126  ( .A1(_f_permutation__n3524 ), .A2(
        _f_permutation__n3525 ), .ZN(_f_permutation__n4731 ) );
  NAND2_X2 _f_permutation__U3125  ( .A1(_f_permutation__round_out[655]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3522 ) );
  NAND2_X2 _f_permutation__U3124  ( .A1(SYNOPSYS_UNCONNECTED_433), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3523 ) );
  NAND2_X2 _f_permutation__U3123  ( .A1(_f_permutation__n3522 ), .A2(
        _f_permutation__n3523 ), .ZN(_f_permutation__n4732 ) );
  NAND2_X2 _f_permutation__U3122  ( .A1(_f_permutation__round_out[654]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3520 ) );
  NAND2_X2 _f_permutation__U3121  ( .A1(SYNOPSYS_UNCONNECTED_434), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3521 ) );
  NAND2_X2 _f_permutation__U3120  ( .A1(_f_permutation__n3520 ), .A2(
        _f_permutation__n3521 ), .ZN(_f_permutation__n4733 ) );
  NAND2_X2 _f_permutation__U3119  ( .A1(_f_permutation__round_out[653]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3518 ) );
  NAND2_X2 _f_permutation__U3118  ( .A1(SYNOPSYS_UNCONNECTED_435), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3519 ) );
  NAND2_X2 _f_permutation__U3117  ( .A1(_f_permutation__n3518 ), .A2(
        _f_permutation__n3519 ), .ZN(_f_permutation__n4734 ) );
  NAND2_X2 _f_permutation__U3116  ( .A1(_f_permutation__round_out[652]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3516 ) );
  NAND2_X2 _f_permutation__U3115  ( .A1(SYNOPSYS_UNCONNECTED_436), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3517 ) );
  NAND2_X2 _f_permutation__U3114  ( .A1(_f_permutation__n3516 ), .A2(
        _f_permutation__n3517 ), .ZN(_f_permutation__n4735 ) );
  NAND2_X2 _f_permutation__U3113  ( .A1(_f_permutation__round_out[651]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3514 ) );
  NAND2_X2 _f_permutation__U3112  ( .A1(SYNOPSYS_UNCONNECTED_437), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3515 ) );
  NAND2_X2 _f_permutation__U3111  ( .A1(_f_permutation__n3514 ), .A2(
        _f_permutation__n3515 ), .ZN(_f_permutation__n4736 ) );
  NAND2_X2 _f_permutation__U3110  ( .A1(_f_permutation__round_out[650]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3512 ) );
  NAND2_X2 _f_permutation__U3109  ( .A1(SYNOPSYS_UNCONNECTED_438), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3513 ) );
  NAND2_X2 _f_permutation__U3108  ( .A1(_f_permutation__n3512 ), .A2(
        _f_permutation__n3513 ), .ZN(_f_permutation__n4737 ) );
  NAND2_X2 _f_permutation__U3107  ( .A1(_f_permutation__round_out[649]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3510 ) );
  NAND2_X2 _f_permutation__U3106  ( .A1(SYNOPSYS_UNCONNECTED_439), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3511 ) );
  NAND2_X2 _f_permutation__U3105  ( .A1(_f_permutation__n3510 ), .A2(
        _f_permutation__n3511 ), .ZN(_f_permutation__n4738 ) );
  NAND2_X2 _f_permutation__U3104  ( .A1(_f_permutation__round_out[648]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3508 ) );
  NAND2_X2 _f_permutation__U3103  ( .A1(SYNOPSYS_UNCONNECTED_440), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3509 ) );
  NAND2_X2 _f_permutation__U3102  ( .A1(_f_permutation__n3508 ), .A2(
        _f_permutation__n3509 ), .ZN(_f_permutation__n4739 ) );
  NAND2_X2 _f_permutation__U3101  ( .A1(_f_permutation__round_out[647]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3506 ) );
  NAND2_X2 _f_permutation__U3100  ( .A1(SYNOPSYS_UNCONNECTED_441), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3507 ) );
  NAND2_X2 _f_permutation__U3099  ( .A1(_f_permutation__n3506 ), .A2(
        _f_permutation__n3507 ), .ZN(_f_permutation__n4740 ) );
  NAND2_X2 _f_permutation__U3098  ( .A1(_f_permutation__round_out[646]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3504 ) );
  NAND2_X2 _f_permutation__U3097  ( .A1(SYNOPSYS_UNCONNECTED_442), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3505 ) );
  NAND2_X2 _f_permutation__U3096  ( .A1(_f_permutation__n3504 ), .A2(
        _f_permutation__n3505 ), .ZN(_f_permutation__n4741 ) );
  NAND2_X2 _f_permutation__U3095  ( .A1(_f_permutation__round_out[645]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3502 ) );
  NAND2_X2 _f_permutation__U3094  ( .A1(SYNOPSYS_UNCONNECTED_443), .A2(
        _f_permutation__n7251 ), .ZN(_f_permutation__n3503 ) );
  NAND2_X2 _f_permutation__U3093  ( .A1(_f_permutation__n3502 ), .A2(
        _f_permutation__n3503 ), .ZN(_f_permutation__n4742 ) );
  NAND2_X2 _f_permutation__U3092  ( .A1(_f_permutation__round_out[644]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3500 ) );
  NAND2_X2 _f_permutation__U3091  ( .A1(SYNOPSYS_UNCONNECTED_444), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3501 ) );
  NAND2_X2 _f_permutation__U3090  ( .A1(_f_permutation__n3500 ), .A2(
        _f_permutation__n3501 ), .ZN(_f_permutation__n4743 ) );
  NAND2_X2 _f_permutation__U3089  ( .A1(_f_permutation__round_out[643]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3498 ) );
  NAND2_X2 _f_permutation__U3088  ( .A1(SYNOPSYS_UNCONNECTED_445), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3499 ) );
  NAND2_X2 _f_permutation__U3087  ( .A1(_f_permutation__n3498 ), .A2(
        _f_permutation__n3499 ), .ZN(_f_permutation__n4744 ) );
  NAND2_X2 _f_permutation__U3086  ( .A1(_f_permutation__round_out[642]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3496 ) );
  NAND2_X2 _f_permutation__U3085  ( .A1(SYNOPSYS_UNCONNECTED_446), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3497 ) );
  NAND2_X2 _f_permutation__U3084  ( .A1(_f_permutation__n3496 ), .A2(
        _f_permutation__n3497 ), .ZN(_f_permutation__n4745 ) );
  NAND2_X2 _f_permutation__U3083  ( .A1(_f_permutation__round_out[641]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3494 ) );
  NAND2_X2 _f_permutation__U3082  ( .A1(SYNOPSYS_UNCONNECTED_447), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3495 ) );
  NAND2_X2 _f_permutation__U3081  ( .A1(_f_permutation__n3494 ), .A2(
        _f_permutation__n3495 ), .ZN(_f_permutation__n4746 ) );
  NAND2_X2 _f_permutation__U3080  ( .A1(_f_permutation__round_out[640]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3492 ) );
  NAND2_X2 _f_permutation__U3079  ( .A1(SYNOPSYS_UNCONNECTED_448), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3493 ) );
  NAND2_X2 _f_permutation__U3078  ( .A1(_f_permutation__n3492 ), .A2(
        _f_permutation__n3493 ), .ZN(_f_permutation__n4747 ) );
  NAND2_X2 _f_permutation__U3077  ( .A1(_f_permutation__round_out[639]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3490 ) );
  NAND2_X2 _f_permutation__U3076  ( .A1(SYNOPSYS_UNCONNECTED_449), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3491 ) );
  NAND2_X2 _f_permutation__U3075  ( .A1(_f_permutation__n3490 ), .A2(
        _f_permutation__n3491 ), .ZN(_f_permutation__n4748 ) );
  NAND2_X2 _f_permutation__U3074  ( .A1(_f_permutation__round_out[638]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3488 ) );
  NAND2_X2 _f_permutation__U3073  ( .A1(SYNOPSYS_UNCONNECTED_450), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3489 ) );
  NAND2_X2 _f_permutation__U3072  ( .A1(_f_permutation__n3488 ), .A2(
        _f_permutation__n3489 ), .ZN(_f_permutation__n4749 ) );
  NAND2_X2 _f_permutation__U3071  ( .A1(_f_permutation__round_out[637]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3486 ) );
  NAND2_X2 _f_permutation__U3070  ( .A1(SYNOPSYS_UNCONNECTED_451), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3487 ) );
  NAND2_X2 _f_permutation__U3069  ( .A1(_f_permutation__n3486 ), .A2(
        _f_permutation__n3487 ), .ZN(_f_permutation__n4750 ) );
  NAND2_X2 _f_permutation__U3068  ( .A1(_f_permutation__round_out[636]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3484 ) );
  NAND2_X2 _f_permutation__U3067  ( .A1(SYNOPSYS_UNCONNECTED_452), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3485 ) );
  NAND2_X2 _f_permutation__U3066  ( .A1(_f_permutation__n3484 ), .A2(
        _f_permutation__n3485 ), .ZN(_f_permutation__n4751 ) );
  NAND2_X2 _f_permutation__U3065  ( .A1(_f_permutation__round_out[635]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3482 ) );
  NAND2_X2 _f_permutation__U3064  ( .A1(SYNOPSYS_UNCONNECTED_453), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3483 ) );
  NAND2_X2 _f_permutation__U3063  ( .A1(_f_permutation__n3482 ), .A2(
        _f_permutation__n3483 ), .ZN(_f_permutation__n4752 ) );
  NAND2_X2 _f_permutation__U3062  ( .A1(_f_permutation__round_out[634]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3480 ) );
  NAND2_X2 _f_permutation__U3061  ( .A1(SYNOPSYS_UNCONNECTED_454), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3481 ) );
  NAND2_X2 _f_permutation__U3060  ( .A1(_f_permutation__n3480 ), .A2(
        _f_permutation__n3481 ), .ZN(_f_permutation__n4753 ) );
  NAND2_X2 _f_permutation__U3059  ( .A1(_f_permutation__round_out[633]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3478 ) );
  NAND2_X2 _f_permutation__U3058  ( .A1(SYNOPSYS_UNCONNECTED_455), .A2(
        _f_permutation__n7252 ), .ZN(_f_permutation__n3479 ) );
  NAND2_X2 _f_permutation__U3057  ( .A1(_f_permutation__n3478 ), .A2(
        _f_permutation__n3479 ), .ZN(_f_permutation__n4754 ) );
  NAND2_X2 _f_permutation__U3056  ( .A1(_f_permutation__round_out[632]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3476 ) );
  NAND2_X2 _f_permutation__U3055  ( .A1(SYNOPSYS_UNCONNECTED_456), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3477 ) );
  NAND2_X2 _f_permutation__U3054  ( .A1(_f_permutation__n3476 ), .A2(
        _f_permutation__n3477 ), .ZN(_f_permutation__n4755 ) );
  NAND2_X2 _f_permutation__U3053  ( .A1(_f_permutation__round_out[631]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3474 ) );
  NAND2_X2 _f_permutation__U3052  ( .A1(SYNOPSYS_UNCONNECTED_457), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3475 ) );
  NAND2_X2 _f_permutation__U3051  ( .A1(_f_permutation__n3474 ), .A2(
        _f_permutation__n3475 ), .ZN(_f_permutation__n4756 ) );
  NAND2_X2 _f_permutation__U3050  ( .A1(_f_permutation__round_out[630]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3472 ) );
  NAND2_X2 _f_permutation__U3049  ( .A1(SYNOPSYS_UNCONNECTED_458), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3473 ) );
  NAND2_X2 _f_permutation__U3048  ( .A1(_f_permutation__n3472 ), .A2(
        _f_permutation__n3473 ), .ZN(_f_permutation__n4757 ) );
  NAND2_X2 _f_permutation__U3047  ( .A1(_f_permutation__round_out[629]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3470 ) );
  NAND2_X2 _f_permutation__U3046  ( .A1(SYNOPSYS_UNCONNECTED_459), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3471 ) );
  NAND2_X2 _f_permutation__U3045  ( .A1(_f_permutation__n3470 ), .A2(
        _f_permutation__n3471 ), .ZN(_f_permutation__n4758 ) );
  NAND2_X2 _f_permutation__U3044  ( .A1(_f_permutation__round_out[628]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3468 ) );
  NAND2_X2 _f_permutation__U3043  ( .A1(SYNOPSYS_UNCONNECTED_460), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3469 ) );
  NAND2_X2 _f_permutation__U3042  ( .A1(_f_permutation__n3468 ), .A2(
        _f_permutation__n3469 ), .ZN(_f_permutation__n4759 ) );
  NAND2_X2 _f_permutation__U3041  ( .A1(_f_permutation__round_out[627]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3466 ) );
  NAND2_X2 _f_permutation__U3040  ( .A1(SYNOPSYS_UNCONNECTED_461), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3467 ) );
  NAND2_X2 _f_permutation__U3039  ( .A1(_f_permutation__n3466 ), .A2(
        _f_permutation__n3467 ), .ZN(_f_permutation__n4760 ) );
  NAND2_X2 _f_permutation__U3038  ( .A1(_f_permutation__round_out[626]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3464 ) );
  NAND2_X2 _f_permutation__U3037  ( .A1(SYNOPSYS_UNCONNECTED_462), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3465 ) );
  NAND2_X2 _f_permutation__U3036  ( .A1(_f_permutation__n3464 ), .A2(
        _f_permutation__n3465 ), .ZN(_f_permutation__n4761 ) );
  NAND2_X2 _f_permutation__U3035  ( .A1(_f_permutation__round_out[625]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3462 ) );
  NAND2_X2 _f_permutation__U3034  ( .A1(SYNOPSYS_UNCONNECTED_463), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3463 ) );
  NAND2_X2 _f_permutation__U3033  ( .A1(_f_permutation__n3462 ), .A2(
        _f_permutation__n3463 ), .ZN(_f_permutation__n4762 ) );
  NAND2_X2 _f_permutation__U3032  ( .A1(_f_permutation__round_out[624]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3460 ) );
  NAND2_X2 _f_permutation__U3031  ( .A1(SYNOPSYS_UNCONNECTED_464), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3461 ) );
  NAND2_X2 _f_permutation__U3030  ( .A1(_f_permutation__n3460 ), .A2(
        _f_permutation__n3461 ), .ZN(_f_permutation__n4763 ) );
  NAND2_X2 _f_permutation__U3029  ( .A1(_f_permutation__round_out[623]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3458 ) );
  NAND2_X2 _f_permutation__U3028  ( .A1(SYNOPSYS_UNCONNECTED_465), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3459 ) );
  NAND2_X2 _f_permutation__U3027  ( .A1(_f_permutation__n3458 ), .A2(
        _f_permutation__n3459 ), .ZN(_f_permutation__n4764 ) );
  NAND2_X2 _f_permutation__U3026  ( .A1(_f_permutation__round_out[622]), .A2(
        _f_permutation__n7081 ), .ZN(_f_permutation__n3456 ) );
  NAND2_X2 _f_permutation__U3025  ( .A1(SYNOPSYS_UNCONNECTED_466), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3457 ) );
  NAND2_X2 _f_permutation__U3024  ( .A1(_f_permutation__n3456 ), .A2(
        _f_permutation__n3457 ), .ZN(_f_permutation__n4765 ) );
  NAND2_X2 _f_permutation__U3023  ( .A1(_f_permutation__round_out[621]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3454 ) );
  NAND2_X2 _f_permutation__U3022  ( .A1(SYNOPSYS_UNCONNECTED_467), .A2(
        _f_permutation__n7253 ), .ZN(_f_permutation__n3455 ) );
  NAND2_X2 _f_permutation__U3021  ( .A1(_f_permutation__n3454 ), .A2(
        _f_permutation__n3455 ), .ZN(_f_permutation__n4766 ) );
  NAND2_X2 _f_permutation__U3020  ( .A1(_f_permutation__round_out[620]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3452 ) );
  NAND2_X2 _f_permutation__U3019  ( .A1(SYNOPSYS_UNCONNECTED_468), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3453 ) );
  NAND2_X2 _f_permutation__U3018  ( .A1(_f_permutation__n3452 ), .A2(
        _f_permutation__n3453 ), .ZN(_f_permutation__n4767 ) );
  NAND2_X2 _f_permutation__U3017  ( .A1(_f_permutation__round_out[619]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3450 ) );
  NAND2_X2 _f_permutation__U3016  ( .A1(SYNOPSYS_UNCONNECTED_469), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3451 ) );
  NAND2_X2 _f_permutation__U3015  ( .A1(_f_permutation__n3450 ), .A2(
        _f_permutation__n3451 ), .ZN(_f_permutation__n4768 ) );
  NAND2_X2 _f_permutation__U3014  ( .A1(_f_permutation__round_out[618]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3448 ) );
  NAND2_X2 _f_permutation__U3013  ( .A1(SYNOPSYS_UNCONNECTED_470), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3449 ) );
  NAND2_X2 _f_permutation__U3012  ( .A1(_f_permutation__n3448 ), .A2(
        _f_permutation__n3449 ), .ZN(_f_permutation__n4769 ) );
  NAND2_X2 _f_permutation__U3011  ( .A1(_f_permutation__round_out[617]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3446 ) );
  NAND2_X2 _f_permutation__U3010  ( .A1(SYNOPSYS_UNCONNECTED_471), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3447 ) );
  NAND2_X2 _f_permutation__U3009  ( .A1(_f_permutation__n3446 ), .A2(
        _f_permutation__n3447 ), .ZN(_f_permutation__n4770 ) );
  NAND2_X2 _f_permutation__U3008  ( .A1(_f_permutation__round_out[616]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3444 ) );
  NAND2_X2 _f_permutation__U3007  ( .A1(SYNOPSYS_UNCONNECTED_472), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3445 ) );
  NAND2_X2 _f_permutation__U3006  ( .A1(_f_permutation__n3444 ), .A2(
        _f_permutation__n3445 ), .ZN(_f_permutation__n4771 ) );
  NAND2_X2 _f_permutation__U3005  ( .A1(_f_permutation__round_out[615]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3442 ) );
  NAND2_X2 _f_permutation__U3004  ( .A1(SYNOPSYS_UNCONNECTED_473), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3443 ) );
  NAND2_X2 _f_permutation__U3003  ( .A1(_f_permutation__n3442 ), .A2(
        _f_permutation__n3443 ), .ZN(_f_permutation__n4772 ) );
  NAND2_X2 _f_permutation__U3002  ( .A1(_f_permutation__round_out[614]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3440 ) );
  NAND2_X2 _f_permutation__U3001  ( .A1(SYNOPSYS_UNCONNECTED_474), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3441 ) );
  NAND2_X2 _f_permutation__U3000  ( .A1(_f_permutation__n3440 ), .A2(
        _f_permutation__n3441 ), .ZN(_f_permutation__n4773 ) );
  NAND2_X2 _f_permutation__U2999  ( .A1(_f_permutation__round_out[613]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3438 ) );
  NAND2_X2 _f_permutation__U2998  ( .A1(SYNOPSYS_UNCONNECTED_475), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3439 ) );
  NAND2_X2 _f_permutation__U2997  ( .A1(_f_permutation__n3438 ), .A2(
        _f_permutation__n3439 ), .ZN(_f_permutation__n4774 ) );
  NAND2_X2 _f_permutation__U2996  ( .A1(_f_permutation__round_out[612]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3436 ) );
  NAND2_X2 _f_permutation__U2995  ( .A1(SYNOPSYS_UNCONNECTED_476), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3437 ) );
  NAND2_X2 _f_permutation__U2994  ( .A1(_f_permutation__n3436 ), .A2(
        _f_permutation__n3437 ), .ZN(_f_permutation__n4775 ) );
  NAND2_X2 _f_permutation__U2993  ( .A1(_f_permutation__round_out[611]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3434 ) );
  NAND2_X2 _f_permutation__U2992  ( .A1(SYNOPSYS_UNCONNECTED_477), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3435 ) );
  NAND2_X2 _f_permutation__U2991  ( .A1(_f_permutation__n3434 ), .A2(
        _f_permutation__n3435 ), .ZN(_f_permutation__n4776 ) );
  NAND2_X2 _f_permutation__U2990  ( .A1(_f_permutation__round_out[610]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3432 ) );
  NAND2_X2 _f_permutation__U2989  ( .A1(SYNOPSYS_UNCONNECTED_478), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3433 ) );
  NAND2_X2 _f_permutation__U2988  ( .A1(_f_permutation__n3432 ), .A2(
        _f_permutation__n3433 ), .ZN(_f_permutation__n4777 ) );
  NAND2_X2 _f_permutation__U2987  ( .A1(_f_permutation__round_out[609]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3430 ) );
  NAND2_X2 _f_permutation__U2986  ( .A1(SYNOPSYS_UNCONNECTED_479), .A2(
        _f_permutation__n7254 ), .ZN(_f_permutation__n3431 ) );
  NAND2_X2 _f_permutation__U2985  ( .A1(_f_permutation__n3430 ), .A2(
        _f_permutation__n3431 ), .ZN(_f_permutation__n4778 ) );
  NAND2_X2 _f_permutation__U2984  ( .A1(_f_permutation__round_out[608]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3428 ) );
  NAND2_X2 _f_permutation__U2983  ( .A1(SYNOPSYS_UNCONNECTED_480), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3429 ) );
  NAND2_X2 _f_permutation__U2982  ( .A1(_f_permutation__n3428 ), .A2(
        _f_permutation__n3429 ), .ZN(_f_permutation__n4779 ) );
  NAND2_X2 _f_permutation__U2981  ( .A1(_f_permutation__round_out[607]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3426 ) );
  NAND2_X2 _f_permutation__U2980  ( .A1(SYNOPSYS_UNCONNECTED_481), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3427 ) );
  NAND2_X2 _f_permutation__U2979  ( .A1(_f_permutation__n3426 ), .A2(
        _f_permutation__n3427 ), .ZN(_f_permutation__n4780 ) );
  NAND2_X2 _f_permutation__U2978  ( .A1(_f_permutation__round_out[606]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3424 ) );
  NAND2_X2 _f_permutation__U2977  ( .A1(SYNOPSYS_UNCONNECTED_482), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3425 ) );
  NAND2_X2 _f_permutation__U2976  ( .A1(_f_permutation__n3424 ), .A2(
        _f_permutation__n3425 ), .ZN(_f_permutation__n4781 ) );
  NAND2_X2 _f_permutation__U2975  ( .A1(_f_permutation__round_out[605]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3422 ) );
  NAND2_X2 _f_permutation__U2974  ( .A1(SYNOPSYS_UNCONNECTED_483), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3423 ) );
  NAND2_X2 _f_permutation__U2973  ( .A1(_f_permutation__n3422 ), .A2(
        _f_permutation__n3423 ), .ZN(_f_permutation__n4782 ) );
  NAND2_X2 _f_permutation__U2972  ( .A1(_f_permutation__round_out[604]), .A2(
        _f_permutation__n7080 ), .ZN(_f_permutation__n3420 ) );
  NAND2_X2 _f_permutation__U2971  ( .A1(SYNOPSYS_UNCONNECTED_484), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3421 ) );
  NAND2_X2 _f_permutation__U2970  ( .A1(_f_permutation__n3420 ), .A2(
        _f_permutation__n3421 ), .ZN(_f_permutation__n4783 ) );
  NAND2_X2 _f_permutation__U2969  ( .A1(_f_permutation__round_out[603]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n3418 ) );
  NAND2_X2 _f_permutation__U2968  ( .A1(SYNOPSYS_UNCONNECTED_485), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3419 ) );
  NAND2_X2 _f_permutation__U2967  ( .A1(_f_permutation__n3418 ), .A2(
        _f_permutation__n3419 ), .ZN(_f_permutation__n4784 ) );
  NAND2_X2 _f_permutation__U2966  ( .A1(_f_permutation__round_out[602]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n3416 ) );
  NAND2_X2 _f_permutation__U2965  ( .A1(SYNOPSYS_UNCONNECTED_486), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3417 ) );
  NAND2_X2 _f_permutation__U2964  ( .A1(_f_permutation__n3416 ), .A2(
        _f_permutation__n3417 ), .ZN(_f_permutation__n4785 ) );
  NAND2_X2 _f_permutation__U2963  ( .A1(_f_permutation__round_out[601]), .A2(
        _f_permutation__n7079 ), .ZN(_f_permutation__n3414 ) );
  NAND2_X2 _f_permutation__U2962  ( .A1(SYNOPSYS_UNCONNECTED_487), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3415 ) );
  NAND2_X2 _f_permutation__U2961  ( .A1(_f_permutation__n3414 ), .A2(
        _f_permutation__n3415 ), .ZN(_f_permutation__n4786 ) );
  NAND2_X2 _f_permutation__U2960  ( .A1(_f_permutation__round_out[600]), .A2(
        _f_permutation__n7082 ), .ZN(_f_permutation__n3412 ) );
  NAND2_X2 _f_permutation__U2959  ( .A1(SYNOPSYS_UNCONNECTED_488), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3413 ) );
  NAND2_X2 _f_permutation__U2958  ( .A1(_f_permutation__n3412 ), .A2(
        _f_permutation__n3413 ), .ZN(_f_permutation__n4787 ) );
  NAND2_X2 _f_permutation__U2957  ( .A1(_f_permutation__round_out[599]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3410 ) );
  NAND2_X2 _f_permutation__U2956  ( .A1(SYNOPSYS_UNCONNECTED_489), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3411 ) );
  NAND2_X2 _f_permutation__U2955  ( .A1(_f_permutation__n3410 ), .A2(
        _f_permutation__n3411 ), .ZN(_f_permutation__n4788 ) );
  NAND2_X2 _f_permutation__U2954  ( .A1(_f_permutation__round_out[598]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3408 ) );
  NAND2_X2 _f_permutation__U2953  ( .A1(SYNOPSYS_UNCONNECTED_490), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3409 ) );
  NAND2_X2 _f_permutation__U2952  ( .A1(_f_permutation__n3408 ), .A2(
        _f_permutation__n3409 ), .ZN(_f_permutation__n4789 ) );
  NAND2_X2 _f_permutation__U2951  ( .A1(_f_permutation__round_out[597]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3406 ) );
  NAND2_X2 _f_permutation__U2950  ( .A1(SYNOPSYS_UNCONNECTED_491), .A2(
        _f_permutation__n7255 ), .ZN(_f_permutation__n3407 ) );
  NAND2_X2 _f_permutation__U2949  ( .A1(_f_permutation__n3406 ), .A2(
        _f_permutation__n3407 ), .ZN(_f_permutation__n4790 ) );
  NAND2_X2 _f_permutation__U2948  ( .A1(_f_permutation__round_out[596]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3404 ) );
  NAND2_X2 _f_permutation__U2947  ( .A1(SYNOPSYS_UNCONNECTED_492), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3405 ) );
  NAND2_X2 _f_permutation__U2946  ( .A1(_f_permutation__n3404 ), .A2(
        _f_permutation__n3405 ), .ZN(_f_permutation__n4791 ) );
  NAND2_X2 _f_permutation__U2945  ( .A1(_f_permutation__round_out[595]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3402 ) );
  NAND2_X2 _f_permutation__U2944  ( .A1(SYNOPSYS_UNCONNECTED_493), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3403 ) );
  NAND2_X2 _f_permutation__U2943  ( .A1(_f_permutation__n3402 ), .A2(
        _f_permutation__n3403 ), .ZN(_f_permutation__n4792 ) );
  NAND2_X2 _f_permutation__U2942  ( .A1(_f_permutation__round_out[594]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3400 ) );
  NAND2_X2 _f_permutation__U2941  ( .A1(SYNOPSYS_UNCONNECTED_494), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3401 ) );
  NAND2_X2 _f_permutation__U2940  ( .A1(_f_permutation__n3400 ), .A2(
        _f_permutation__n3401 ), .ZN(_f_permutation__n4793 ) );
  NAND2_X2 _f_permutation__U2939  ( .A1(_f_permutation__round_out[593]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3398 ) );
  NAND2_X2 _f_permutation__U2938  ( .A1(SYNOPSYS_UNCONNECTED_495), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3399 ) );
  NAND2_X2 _f_permutation__U2937  ( .A1(_f_permutation__n3398 ), .A2(
        _f_permutation__n3399 ), .ZN(_f_permutation__n4794 ) );
  NAND2_X2 _f_permutation__U2936  ( .A1(_f_permutation__round_out[592]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3396 ) );
  NAND2_X2 _f_permutation__U2935  ( .A1(SYNOPSYS_UNCONNECTED_496), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3397 ) );
  NAND2_X2 _f_permutation__U2934  ( .A1(_f_permutation__n3396 ), .A2(
        _f_permutation__n3397 ), .ZN(_f_permutation__n4795 ) );
  NAND2_X2 _f_permutation__U2933  ( .A1(_f_permutation__round_out[591]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3394 ) );
  NAND2_X2 _f_permutation__U2932  ( .A1(SYNOPSYS_UNCONNECTED_497), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3395 ) );
  NAND2_X2 _f_permutation__U2931  ( .A1(_f_permutation__n3394 ), .A2(
        _f_permutation__n3395 ), .ZN(_f_permutation__n4796 ) );
  NAND2_X2 _f_permutation__U2930  ( .A1(_f_permutation__round_out[590]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3392 ) );
  NAND2_X2 _f_permutation__U2929  ( .A1(SYNOPSYS_UNCONNECTED_498), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3393 ) );
  NAND2_X2 _f_permutation__U2928  ( .A1(_f_permutation__n3392 ), .A2(
        _f_permutation__n3393 ), .ZN(_f_permutation__n4797 ) );
  NAND2_X2 _f_permutation__U2927  ( .A1(_f_permutation__round_out[589]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3390 ) );
  NAND2_X2 _f_permutation__U2926  ( .A1(SYNOPSYS_UNCONNECTED_499), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3391 ) );
  NAND2_X2 _f_permutation__U2925  ( .A1(_f_permutation__n3390 ), .A2(
        _f_permutation__n3391 ), .ZN(_f_permutation__n4798 ) );
  NAND2_X2 _f_permutation__U2924  ( .A1(_f_permutation__round_out[588]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3388 ) );
  NAND2_X2 _f_permutation__U2923  ( .A1(SYNOPSYS_UNCONNECTED_500), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3389 ) );
  NAND2_X2 _f_permutation__U2922  ( .A1(_f_permutation__n3388 ), .A2(
        _f_permutation__n3389 ), .ZN(_f_permutation__n4799 ) );
  NAND2_X2 _f_permutation__U2921  ( .A1(_f_permutation__round_out[587]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3386 ) );
  NAND2_X2 _f_permutation__U2920  ( .A1(SYNOPSYS_UNCONNECTED_501), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3387 ) );
  NAND2_X2 _f_permutation__U2919  ( .A1(_f_permutation__n3386 ), .A2(
        _f_permutation__n3387 ), .ZN(_f_permutation__n4800 ) );
  NAND2_X2 _f_permutation__U2918  ( .A1(_f_permutation__round_out[586]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3384 ) );
  NAND2_X2 _f_permutation__U2917  ( .A1(SYNOPSYS_UNCONNECTED_502), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3385 ) );
  NAND2_X2 _f_permutation__U2916  ( .A1(_f_permutation__n3384 ), .A2(
        _f_permutation__n3385 ), .ZN(_f_permutation__n4801 ) );
  NAND2_X2 _f_permutation__U2915  ( .A1(_f_permutation__round_out[585]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3382 ) );
  NAND2_X2 _f_permutation__U2914  ( .A1(SYNOPSYS_UNCONNECTED_503), .A2(
        _f_permutation__n7256 ), .ZN(_f_permutation__n3383 ) );
  NAND2_X2 _f_permutation__U2913  ( .A1(_f_permutation__n3382 ), .A2(
        _f_permutation__n3383 ), .ZN(_f_permutation__n4802 ) );
  NAND2_X2 _f_permutation__U2912  ( .A1(_f_permutation__round_out[584]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3380 ) );
  NAND2_X2 _f_permutation__U2911  ( .A1(SYNOPSYS_UNCONNECTED_504), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3381 ) );
  NAND2_X2 _f_permutation__U2910  ( .A1(_f_permutation__n3380 ), .A2(
        _f_permutation__n3381 ), .ZN(_f_permutation__n4803 ) );
  NAND2_X2 _f_permutation__U2909  ( .A1(_f_permutation__round_out[583]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3378 ) );
  NAND2_X2 _f_permutation__U2908  ( .A1(SYNOPSYS_UNCONNECTED_505), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3379 ) );
  NAND2_X2 _f_permutation__U2907  ( .A1(_f_permutation__n3378 ), .A2(
        _f_permutation__n3379 ), .ZN(_f_permutation__n4804 ) );
  NAND2_X2 _f_permutation__U2906  ( .A1(_f_permutation__round_out[582]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3376 ) );
  NAND2_X2 _f_permutation__U2905  ( .A1(SYNOPSYS_UNCONNECTED_506), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3377 ) );
  NAND2_X2 _f_permutation__U2904  ( .A1(_f_permutation__n3376 ), .A2(
        _f_permutation__n3377 ), .ZN(_f_permutation__n4805 ) );
  NAND2_X2 _f_permutation__U2903  ( .A1(_f_permutation__round_out[581]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3374 ) );
  NAND2_X2 _f_permutation__U2902  ( .A1(SYNOPSYS_UNCONNECTED_507), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3375 ) );
  NAND2_X2 _f_permutation__U2901  ( .A1(_f_permutation__n3374 ), .A2(
        _f_permutation__n3375 ), .ZN(_f_permutation__n4806 ) );
  NAND2_X2 _f_permutation__U2900  ( .A1(_f_permutation__round_out[580]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3372 ) );
  NAND2_X2 _f_permutation__U2899  ( .A1(SYNOPSYS_UNCONNECTED_508), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3373 ) );
  NAND2_X2 _f_permutation__U2898  ( .A1(_f_permutation__n3372 ), .A2(
        _f_permutation__n3373 ), .ZN(_f_permutation__n4807 ) );
  NAND2_X2 _f_permutation__U2897  ( .A1(_f_permutation__round_out[579]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3370 ) );
  NAND2_X2 _f_permutation__U2896  ( .A1(SYNOPSYS_UNCONNECTED_509), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3371 ) );
  NAND2_X2 _f_permutation__U2895  ( .A1(_f_permutation__n3370 ), .A2(
        _f_permutation__n3371 ), .ZN(_f_permutation__n4808 ) );
  NAND2_X2 _f_permutation__U2894  ( .A1(_f_permutation__round_out[578]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3368 ) );
  NAND2_X2 _f_permutation__U2893  ( .A1(SYNOPSYS_UNCONNECTED_510), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3369 ) );
  NAND2_X2 _f_permutation__U2892  ( .A1(_f_permutation__n3368 ), .A2(
        _f_permutation__n3369 ), .ZN(_f_permutation__n4809 ) );
  NAND2_X2 _f_permutation__U2891  ( .A1(_f_permutation__round_out[577]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3366 ) );
  NAND2_X2 _f_permutation__U2890  ( .A1(SYNOPSYS_UNCONNECTED_511), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3367 ) );
  NAND2_X2 _f_permutation__U2889  ( .A1(_f_permutation__n3366 ), .A2(
        _f_permutation__n3367 ), .ZN(_f_permutation__n4810 ) );
  NAND2_X2 _f_permutation__U2888  ( .A1(_f_permutation__round_out[576]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3364 ) );
  NAND2_X2 _f_permutation__U2887  ( .A1(SYNOPSYS_UNCONNECTED_512), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3365 ) );
  NAND2_X2 _f_permutation__U2886  ( .A1(_f_permutation__n3364 ), .A2(
        _f_permutation__n3365 ), .ZN(_f_permutation__n4811 ) );
  NAND2_X2 _f_permutation__U2885  ( .A1(_f_permutation__round_out[575]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3362 ) );
  NAND2_X2 _f_permutation__U2884  ( .A1(SYNOPSYS_UNCONNECTED_513), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3363 ) );
  NAND2_X2 _f_permutation__U2883  ( .A1(_f_permutation__n3362 ), .A2(
        _f_permutation__n3363 ), .ZN(_f_permutation__n4812 ) );
  NAND2_X2 _f_permutation__U2882  ( .A1(_f_permutation__round_out[574]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3360 ) );
  NAND2_X2 _f_permutation__U2881  ( .A1(SYNOPSYS_UNCONNECTED_514), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3361 ) );
  NAND2_X2 _f_permutation__U2880  ( .A1(_f_permutation__n3360 ), .A2(
        _f_permutation__n3361 ), .ZN(_f_permutation__n4813 ) );
  NAND2_X2 _f_permutation__U2879  ( .A1(_f_permutation__round_out[573]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3358 ) );
  NAND2_X2 _f_permutation__U2878  ( .A1(SYNOPSYS_UNCONNECTED_515), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n3359 ) );
  NAND2_X2 _f_permutation__U2877  ( .A1(_f_permutation__n3358 ), .A2(
        _f_permutation__n3359 ), .ZN(_f_permutation__n4814 ) );
  NAND2_X2 _f_permutation__U2876  ( .A1(_f_permutation__round_out[572]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3356 ) );
  NAND2_X2 _f_permutation__U2875  ( .A1(SYNOPSYS_UNCONNECTED_516), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3357 ) );
  NAND2_X2 _f_permutation__U2874  ( .A1(_f_permutation__n3356 ), .A2(
        _f_permutation__n3357 ), .ZN(_f_permutation__n4815 ) );
  NAND2_X2 _f_permutation__U2873  ( .A1(_f_permutation__round_out[571]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3354 ) );
  NAND2_X2 _f_permutation__U2872  ( .A1(SYNOPSYS_UNCONNECTED_517), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3355 ) );
  NAND2_X2 _f_permutation__U2871  ( .A1(_f_permutation__n3354 ), .A2(
        _f_permutation__n3355 ), .ZN(_f_permutation__n4816 ) );
  NAND2_X2 _f_permutation__U2870  ( .A1(_f_permutation__round_out[570]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3352 ) );
  NAND2_X2 _f_permutation__U2869  ( .A1(SYNOPSYS_UNCONNECTED_518), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3353 ) );
  NAND2_X2 _f_permutation__U2868  ( .A1(_f_permutation__n3352 ), .A2(
        _f_permutation__n3353 ), .ZN(_f_permutation__n4817 ) );
  NAND2_X2 _f_permutation__U2867  ( .A1(_f_permutation__round_out[569]), .A2(
        _f_permutation__n7068 ), .ZN(_f_permutation__n3350 ) );
  NAND2_X2 _f_permutation__U2866  ( .A1(SYNOPSYS_UNCONNECTED_519), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3351 ) );
  NAND2_X2 _f_permutation__U2865  ( .A1(_f_permutation__n3350 ), .A2(
        _f_permutation__n3351 ), .ZN(_f_permutation__n4818 ) );
  NAND2_X2 _f_permutation__U2864  ( .A1(_f_permutation__round_out[568]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3348 ) );
  NAND2_X2 _f_permutation__U2863  ( .A1(SYNOPSYS_UNCONNECTED_520), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3349 ) );
  NAND2_X2 _f_permutation__U2862  ( .A1(_f_permutation__n3348 ), .A2(
        _f_permutation__n3349 ), .ZN(_f_permutation__n4819 ) );
  NAND2_X2 _f_permutation__U2861  ( .A1(_f_permutation__round_out[567]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3346 ) );
  NAND2_X2 _f_permutation__U2860  ( .A1(SYNOPSYS_UNCONNECTED_521), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3347 ) );
  NAND2_X2 _f_permutation__U2859  ( .A1(_f_permutation__n3346 ), .A2(
        _f_permutation__n3347 ), .ZN(_f_permutation__n4820 ) );
  NAND2_X2 _f_permutation__U2858  ( .A1(_f_permutation__round_out[566]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3344 ) );
  NAND2_X2 _f_permutation__U2857  ( .A1(SYNOPSYS_UNCONNECTED_522), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3345 ) );
  NAND2_X2 _f_permutation__U2856  ( .A1(_f_permutation__n3344 ), .A2(
        _f_permutation__n3345 ), .ZN(_f_permutation__n4821 ) );
  NAND2_X2 _f_permutation__U2855  ( .A1(_f_permutation__round_out[565]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3342 ) );
  NAND2_X2 _f_permutation__U2854  ( .A1(SYNOPSYS_UNCONNECTED_523), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3343 ) );
  NAND2_X2 _f_permutation__U2853  ( .A1(_f_permutation__n3342 ), .A2(
        _f_permutation__n3343 ), .ZN(_f_permutation__n4822 ) );
  NAND2_X2 _f_permutation__U2852  ( .A1(_f_permutation__round_out[564]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3340 ) );
  NAND2_X2 _f_permutation__U2851  ( .A1(SYNOPSYS_UNCONNECTED_524), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3341 ) );
  NAND2_X2 _f_permutation__U2850  ( .A1(_f_permutation__n3340 ), .A2(
        _f_permutation__n3341 ), .ZN(_f_permutation__n4823 ) );
  NAND2_X2 _f_permutation__U2849  ( .A1(_f_permutation__round_out[563]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3338 ) );
  NAND2_X2 _f_permutation__U2848  ( .A1(SYNOPSYS_UNCONNECTED_525), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3339 ) );
  NAND2_X2 _f_permutation__U2847  ( .A1(_f_permutation__n3338 ), .A2(
        _f_permutation__n3339 ), .ZN(_f_permutation__n4824 ) );
  NAND2_X2 _f_permutation__U2846  ( .A1(_f_permutation__round_out[562]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3336 ) );
  NAND2_X2 _f_permutation__U2845  ( .A1(SYNOPSYS_UNCONNECTED_526), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3337 ) );
  NAND2_X2 _f_permutation__U2844  ( .A1(_f_permutation__n3336 ), .A2(
        _f_permutation__n3337 ), .ZN(_f_permutation__n4825 ) );
  NAND2_X2 _f_permutation__U2843  ( .A1(_f_permutation__round_out[561]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3334 ) );
  NAND2_X2 _f_permutation__U2842  ( .A1(SYNOPSYS_UNCONNECTED_527), .A2(
        _f_permutation__n7258 ), .ZN(_f_permutation__n3335 ) );
  NAND2_X2 _f_permutation__U2841  ( .A1(_f_permutation__n3334 ), .A2(
        _f_permutation__n3335 ), .ZN(_f_permutation__n4826 ) );
  NAND2_X2 _f_permutation__U2840  ( .A1(_f_permutation__round_out[560]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3332 ) );
  NAND2_X2 _f_permutation__U2839  ( .A1(SYNOPSYS_UNCONNECTED_528), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3333 ) );
  NAND2_X2 _f_permutation__U2838  ( .A1(_f_permutation__n3332 ), .A2(
        _f_permutation__n3333 ), .ZN(_f_permutation__n4827 ) );
  NAND2_X2 _f_permutation__U2837  ( .A1(_f_permutation__round_out[559]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3330 ) );
  NAND2_X2 _f_permutation__U2836  ( .A1(SYNOPSYS_UNCONNECTED_529), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3331 ) );
  NAND2_X2 _f_permutation__U2835  ( .A1(_f_permutation__n3330 ), .A2(
        _f_permutation__n3331 ), .ZN(_f_permutation__n4828 ) );
  NAND2_X2 _f_permutation__U2834  ( .A1(_f_permutation__round_out[558]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3328 ) );
  NAND2_X2 _f_permutation__U2833  ( .A1(SYNOPSYS_UNCONNECTED_530), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3329 ) );
  NAND2_X2 _f_permutation__U2832  ( .A1(_f_permutation__n3328 ), .A2(
        _f_permutation__n3329 ), .ZN(_f_permutation__n4829 ) );
  NAND2_X2 _f_permutation__U2831  ( .A1(_f_permutation__round_out[557]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3326 ) );
  NAND2_X2 _f_permutation__U2830  ( .A1(SYNOPSYS_UNCONNECTED_531), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3327 ) );
  NAND2_X2 _f_permutation__U2829  ( .A1(_f_permutation__n3326 ), .A2(
        _f_permutation__n3327 ), .ZN(_f_permutation__n4830 ) );
  NAND2_X2 _f_permutation__U2828  ( .A1(_f_permutation__round_out[556]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3324 ) );
  NAND2_X2 _f_permutation__U2827  ( .A1(SYNOPSYS_UNCONNECTED_532), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3325 ) );
  NAND2_X2 _f_permutation__U2826  ( .A1(_f_permutation__n3324 ), .A2(
        _f_permutation__n3325 ), .ZN(_f_permutation__n4831 ) );
  NAND2_X2 _f_permutation__U2825  ( .A1(_f_permutation__round_out[555]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3322 ) );
  NAND2_X2 _f_permutation__U2824  ( .A1(SYNOPSYS_UNCONNECTED_533), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3323 ) );
  NAND2_X2 _f_permutation__U2823  ( .A1(_f_permutation__n3322 ), .A2(
        _f_permutation__n3323 ), .ZN(_f_permutation__n4832 ) );
  NAND2_X2 _f_permutation__U2822  ( .A1(_f_permutation__round_out[554]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3320 ) );
  NAND2_X2 _f_permutation__U2821  ( .A1(SYNOPSYS_UNCONNECTED_534), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3321 ) );
  NAND2_X2 _f_permutation__U2820  ( .A1(_f_permutation__n3320 ), .A2(
        _f_permutation__n3321 ), .ZN(_f_permutation__n4833 ) );
  NAND2_X2 _f_permutation__U2819  ( .A1(_f_permutation__round_out[553]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3318 ) );
  NAND2_X2 _f_permutation__U2818  ( .A1(SYNOPSYS_UNCONNECTED_535), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3319 ) );
  NAND2_X2 _f_permutation__U2817  ( .A1(_f_permutation__n3318 ), .A2(
        _f_permutation__n3319 ), .ZN(_f_permutation__n4834 ) );
  NAND2_X2 _f_permutation__U2816  ( .A1(_f_permutation__round_out[552]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3316 ) );
  NAND2_X2 _f_permutation__U2815  ( .A1(SYNOPSYS_UNCONNECTED_536), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3317 ) );
  NAND2_X2 _f_permutation__U2814  ( .A1(_f_permutation__n3316 ), .A2(
        _f_permutation__n3317 ), .ZN(_f_permutation__n4835 ) );
  NAND2_X2 _f_permutation__U2813  ( .A1(_f_permutation__round_out[551]), .A2(
        _f_permutation__n7067 ), .ZN(_f_permutation__n3314 ) );
  NAND2_X2 _f_permutation__U2812  ( .A1(SYNOPSYS_UNCONNECTED_537), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3315 ) );
  NAND2_X2 _f_permutation__U2811  ( .A1(_f_permutation__n3314 ), .A2(
        _f_permutation__n3315 ), .ZN(_f_permutation__n4836 ) );
  NAND2_X2 _f_permutation__U2810  ( .A1(_f_permutation__round_out[550]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3312 ) );
  NAND2_X2 _f_permutation__U2809  ( .A1(SYNOPSYS_UNCONNECTED_538), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3313 ) );
  NAND2_X2 _f_permutation__U2808  ( .A1(_f_permutation__n3312 ), .A2(
        _f_permutation__n3313 ), .ZN(_f_permutation__n4837 ) );
  NAND2_X2 _f_permutation__U2807  ( .A1(_f_permutation__round_out[549]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3310 ) );
  NAND2_X2 _f_permutation__U2806  ( .A1(SYNOPSYS_UNCONNECTED_539), .A2(
        _f_permutation__n7259 ), .ZN(_f_permutation__n3311 ) );
  NAND2_X2 _f_permutation__U2805  ( .A1(_f_permutation__n3310 ), .A2(
        _f_permutation__n3311 ), .ZN(_f_permutation__n4838 ) );
  NAND2_X2 _f_permutation__U2804  ( .A1(_f_permutation__round_out[548]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3308 ) );
  NAND2_X2 _f_permutation__U2803  ( .A1(SYNOPSYS_UNCONNECTED_540), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3309 ) );
  NAND2_X2 _f_permutation__U2802  ( .A1(_f_permutation__n3308 ), .A2(
        _f_permutation__n3309 ), .ZN(_f_permutation__n4839 ) );
  NAND2_X2 _f_permutation__U2801  ( .A1(_f_permutation__round_out[547]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3306 ) );
  NAND2_X2 _f_permutation__U2800  ( .A1(SYNOPSYS_UNCONNECTED_541), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3307 ) );
  NAND2_X2 _f_permutation__U2799  ( .A1(_f_permutation__n3306 ), .A2(
        _f_permutation__n3307 ), .ZN(_f_permutation__n4840 ) );
  NAND2_X2 _f_permutation__U2798  ( .A1(_f_permutation__round_out[546]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3304 ) );
  NAND2_X2 _f_permutation__U2797  ( .A1(SYNOPSYS_UNCONNECTED_542), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3305 ) );
  NAND2_X2 _f_permutation__U2796  ( .A1(_f_permutation__n3304 ), .A2(
        _f_permutation__n3305 ), .ZN(_f_permutation__n4841 ) );
  NAND2_X2 _f_permutation__U2795  ( .A1(_f_permutation__round_out[545]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3302 ) );
  NAND2_X2 _f_permutation__U2794  ( .A1(SYNOPSYS_UNCONNECTED_543), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3303 ) );
  NAND2_X2 _f_permutation__U2793  ( .A1(_f_permutation__n3302 ), .A2(
        _f_permutation__n3303 ), .ZN(_f_permutation__n4842 ) );
  NAND2_X2 _f_permutation__U2792  ( .A1(_f_permutation__round_out[544]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3300 ) );
  NAND2_X2 _f_permutation__U2791  ( .A1(SYNOPSYS_UNCONNECTED_544), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3301 ) );
  NAND2_X2 _f_permutation__U2790  ( .A1(_f_permutation__n3300 ), .A2(
        _f_permutation__n3301 ), .ZN(_f_permutation__n4843 ) );
  NAND2_X2 _f_permutation__U2789  ( .A1(_f_permutation__round_out[543]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3298 ) );
  NAND2_X2 _f_permutation__U2788  ( .A1(SYNOPSYS_UNCONNECTED_545), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3299 ) );
  NAND2_X2 _f_permutation__U2787  ( .A1(_f_permutation__n3298 ), .A2(
        _f_permutation__n3299 ), .ZN(_f_permutation__n4844 ) );
  NAND2_X2 _f_permutation__U2786  ( .A1(_f_permutation__round_out[542]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3296 ) );
  NAND2_X2 _f_permutation__U2785  ( .A1(SYNOPSYS_UNCONNECTED_546), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3297 ) );
  NAND2_X2 _f_permutation__U2784  ( .A1(_f_permutation__n3296 ), .A2(
        _f_permutation__n3297 ), .ZN(_f_permutation__n4845 ) );
  NAND2_X2 _f_permutation__U2783  ( .A1(_f_permutation__round_out[541]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3294 ) );
  NAND2_X2 _f_permutation__U2782  ( .A1(SYNOPSYS_UNCONNECTED_547), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3295 ) );
  NAND2_X2 _f_permutation__U2781  ( .A1(_f_permutation__n3294 ), .A2(
        _f_permutation__n3295 ), .ZN(_f_permutation__n4846 ) );
  NAND2_X2 _f_permutation__U2780  ( .A1(_f_permutation__round_out[540]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3292 ) );
  NAND2_X2 _f_permutation__U2779  ( .A1(SYNOPSYS_UNCONNECTED_548), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3293 ) );
  NAND2_X2 _f_permutation__U2778  ( .A1(_f_permutation__n3292 ), .A2(
        _f_permutation__n3293 ), .ZN(_f_permutation__n4847 ) );
  NAND2_X2 _f_permutation__U2777  ( .A1(_f_permutation__round_out[539]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3290 ) );
  NAND2_X2 _f_permutation__U2776  ( .A1(SYNOPSYS_UNCONNECTED_549), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3291 ) );
  NAND2_X2 _f_permutation__U2775  ( .A1(_f_permutation__n3290 ), .A2(
        _f_permutation__n3291 ), .ZN(_f_permutation__n4848 ) );
  NAND2_X2 _f_permutation__U2774  ( .A1(_f_permutation__round_out[538]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3288 ) );
  NAND2_X2 _f_permutation__U2773  ( .A1(SYNOPSYS_UNCONNECTED_550), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3289 ) );
  NAND2_X2 _f_permutation__U2772  ( .A1(_f_permutation__n3288 ), .A2(
        _f_permutation__n3289 ), .ZN(_f_permutation__n4849 ) );
  NAND2_X2 _f_permutation__U2771  ( .A1(_f_permutation__round_out[537]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3286 ) );
  NAND2_X2 _f_permutation__U2770  ( .A1(SYNOPSYS_UNCONNECTED_551), .A2(
        _f_permutation__n7260 ), .ZN(_f_permutation__n3287 ) );
  NAND2_X2 _f_permutation__U2769  ( .A1(_f_permutation__n3286 ), .A2(
        _f_permutation__n3287 ), .ZN(_f_permutation__n4850 ) );
  NAND2_X2 _f_permutation__U2768  ( .A1(_f_permutation__round_out[536]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3284 ) );
  NAND2_X2 _f_permutation__U2767  ( .A1(SYNOPSYS_UNCONNECTED_552), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3285 ) );
  NAND2_X2 _f_permutation__U2766  ( .A1(_f_permutation__n3284 ), .A2(
        _f_permutation__n3285 ), .ZN(_f_permutation__n4851 ) );
  NAND2_X2 _f_permutation__U2765  ( .A1(_f_permutation__round_out[535]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3282 ) );
  NAND2_X2 _f_permutation__U2764  ( .A1(SYNOPSYS_UNCONNECTED_553), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3283 ) );
  NAND2_X2 _f_permutation__U2763  ( .A1(_f_permutation__n3282 ), .A2(
        _f_permutation__n3283 ), .ZN(_f_permutation__n4852 ) );
  NAND2_X2 _f_permutation__U2762  ( .A1(_f_permutation__round_out[534]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3280 ) );
  NAND2_X2 _f_permutation__U2761  ( .A1(SYNOPSYS_UNCONNECTED_554), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3281 ) );
  NAND2_X2 _f_permutation__U2760  ( .A1(_f_permutation__n3280 ), .A2(
        _f_permutation__n3281 ), .ZN(_f_permutation__n4853 ) );
  NAND2_X2 _f_permutation__U2759  ( .A1(_f_permutation__round_out[533]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3278 ) );
  NAND2_X2 _f_permutation__U2758  ( .A1(SYNOPSYS_UNCONNECTED_555), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3279 ) );
  NAND2_X2 _f_permutation__U2757  ( .A1(_f_permutation__n3278 ), .A2(
        _f_permutation__n3279 ), .ZN(_f_permutation__n4854 ) );
  NAND2_X2 _f_permutation__U2756  ( .A1(_f_permutation__round_out[532]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3276 ) );
  NAND2_X2 _f_permutation__U2755  ( .A1(SYNOPSYS_UNCONNECTED_556), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3277 ) );
  NAND2_X2 _f_permutation__U2754  ( .A1(_f_permutation__n3276 ), .A2(
        _f_permutation__n3277 ), .ZN(_f_permutation__n4855 ) );
  NAND2_X2 _f_permutation__U2753  ( .A1(_f_permutation__round_out[531]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3274 ) );
  NAND2_X2 _f_permutation__U2752  ( .A1(SYNOPSYS_UNCONNECTED_557), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3275 ) );
  NAND2_X2 _f_permutation__U2751  ( .A1(_f_permutation__n3274 ), .A2(
        _f_permutation__n3275 ), .ZN(_f_permutation__n4856 ) );
  NAND2_X2 _f_permutation__U2750  ( .A1(_f_permutation__round_out[530]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3272 ) );
  NAND2_X2 _f_permutation__U2749  ( .A1(SYNOPSYS_UNCONNECTED_558), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3273 ) );
  NAND2_X2 _f_permutation__U2748  ( .A1(_f_permutation__n3272 ), .A2(
        _f_permutation__n3273 ), .ZN(_f_permutation__n4857 ) );
  NAND2_X2 _f_permutation__U2747  ( .A1(_f_permutation__round_out[529]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3270 ) );
  NAND2_X2 _f_permutation__U2746  ( .A1(SYNOPSYS_UNCONNECTED_559), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3271 ) );
  NAND2_X2 _f_permutation__U2745  ( .A1(_f_permutation__n3270 ), .A2(
        _f_permutation__n3271 ), .ZN(_f_permutation__n4858 ) );
  NAND2_X2 _f_permutation__U2744  ( .A1(_f_permutation__round_out[528]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3268 ) );
  NAND2_X2 _f_permutation__U2743  ( .A1(SYNOPSYS_UNCONNECTED_560), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3269 ) );
  NAND2_X2 _f_permutation__U2742  ( .A1(_f_permutation__n3268 ), .A2(
        _f_permutation__n3269 ), .ZN(_f_permutation__n4859 ) );
  NAND2_X2 _f_permutation__U2741  ( .A1(_f_permutation__round_out[527]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3266 ) );
  NAND2_X2 _f_permutation__U2740  ( .A1(SYNOPSYS_UNCONNECTED_561), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3267 ) );
  NAND2_X2 _f_permutation__U2739  ( .A1(_f_permutation__n3266 ), .A2(
        _f_permutation__n3267 ), .ZN(_f_permutation__n4860 ) );
  NAND2_X2 _f_permutation__U2738  ( .A1(_f_permutation__round_out[526]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3264 ) );
  NAND2_X2 _f_permutation__U2737  ( .A1(SYNOPSYS_UNCONNECTED_562), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3265 ) );
  NAND2_X2 _f_permutation__U2736  ( .A1(_f_permutation__n3264 ), .A2(
        _f_permutation__n3265 ), .ZN(_f_permutation__n4861 ) );
  NAND2_X2 _f_permutation__U2735  ( .A1(_f_permutation__round_out[525]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3262 ) );
  NAND2_X2 _f_permutation__U2734  ( .A1(SYNOPSYS_UNCONNECTED_563), .A2(
        _f_permutation__n7261 ), .ZN(_f_permutation__n3263 ) );
  NAND2_X2 _f_permutation__U2733  ( .A1(_f_permutation__n3262 ), .A2(
        _f_permutation__n3263 ), .ZN(_f_permutation__n4862 ) );
  NAND2_X2 _f_permutation__U2732  ( .A1(_f_permutation__round_out[524]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3260 ) );
  NAND2_X2 _f_permutation__U2731  ( .A1(SYNOPSYS_UNCONNECTED_564), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3261 ) );
  NAND2_X2 _f_permutation__U2730  ( .A1(_f_permutation__n3260 ), .A2(
        _f_permutation__n3261 ), .ZN(_f_permutation__n4863 ) );
  NAND2_X2 _f_permutation__U2729  ( .A1(_f_permutation__round_out[523]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3258 ) );
  NAND2_X2 _f_permutation__U2728  ( .A1(SYNOPSYS_UNCONNECTED_565), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3259 ) );
  NAND2_X2 _f_permutation__U2727  ( .A1(_f_permutation__n3258 ), .A2(
        _f_permutation__n3259 ), .ZN(_f_permutation__n4864 ) );
  NAND2_X2 _f_permutation__U2726  ( .A1(_f_permutation__round_out[522]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3256 ) );
  NAND2_X2 _f_permutation__U2725  ( .A1(SYNOPSYS_UNCONNECTED_566), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3257 ) );
  NAND2_X2 _f_permutation__U2724  ( .A1(_f_permutation__n3256 ), .A2(
        _f_permutation__n3257 ), .ZN(_f_permutation__n4865 ) );
  NAND2_X2 _f_permutation__U2723  ( .A1(_f_permutation__round_out[521]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3254 ) );
  NAND2_X2 _f_permutation__U2722  ( .A1(SYNOPSYS_UNCONNECTED_567), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3255 ) );
  NAND2_X2 _f_permutation__U2721  ( .A1(_f_permutation__n3254 ), .A2(
        _f_permutation__n3255 ), .ZN(_f_permutation__n4866 ) );
  NAND2_X2 _f_permutation__U2720  ( .A1(_f_permutation__round_out[520]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3252 ) );
  NAND2_X2 _f_permutation__U2719  ( .A1(SYNOPSYS_UNCONNECTED_568), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3253 ) );
  NAND2_X2 _f_permutation__U2718  ( .A1(_f_permutation__n3252 ), .A2(
        _f_permutation__n3253 ), .ZN(_f_permutation__n4867 ) );
  NAND2_X2 _f_permutation__U2717  ( .A1(_f_permutation__round_out[519]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3250 ) );
  NAND2_X2 _f_permutation__U2716  ( .A1(SYNOPSYS_UNCONNECTED_569), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3251 ) );
  NAND2_X2 _f_permutation__U2715  ( .A1(_f_permutation__n3250 ), .A2(
        _f_permutation__n3251 ), .ZN(_f_permutation__n4868 ) );
  NAND2_X2 _f_permutation__U2714  ( .A1(_f_permutation__round_out[518]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3248 ) );
  NAND2_X2 _f_permutation__U2713  ( .A1(SYNOPSYS_UNCONNECTED_570), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3249 ) );
  NAND2_X2 _f_permutation__U2712  ( .A1(_f_permutation__n3248 ), .A2(
        _f_permutation__n3249 ), .ZN(_f_permutation__n4869 ) );
  NAND2_X2 _f_permutation__U2711  ( .A1(_f_permutation__round_out[517]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3246 ) );
  NAND2_X2 _f_permutation__U2710  ( .A1(SYNOPSYS_UNCONNECTED_571), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3247 ) );
  NAND2_X2 _f_permutation__U2709  ( .A1(_f_permutation__n3246 ), .A2(
        _f_permutation__n3247 ), .ZN(_f_permutation__n4870 ) );
  NAND2_X2 _f_permutation__U2708  ( .A1(_f_permutation__round_out[516]), .A2(
        _f_permutation__n7065 ), .ZN(_f_permutation__n3244 ) );
  NAND2_X2 _f_permutation__U2707  ( .A1(SYNOPSYS_UNCONNECTED_572), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3245 ) );
  NAND2_X2 _f_permutation__U2706  ( .A1(_f_permutation__n3244 ), .A2(
        _f_permutation__n3245 ), .ZN(_f_permutation__n4871 ) );
  NAND2_X2 _f_permutation__U2705  ( .A1(_f_permutation__round_out[515]), .A2(
        _f_permutation__n7168 ), .ZN(_f_permutation__n3242 ) );
  NAND2_X2 _f_permutation__U2704  ( .A1(SYNOPSYS_UNCONNECTED_573), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3243 ) );
  NAND2_X2 _f_permutation__U2703  ( .A1(_f_permutation__n3242 ), .A2(
        _f_permutation__n3243 ), .ZN(_f_permutation__n4872 ) );
  NAND2_X2 _f_permutation__U2702  ( .A1(_f_permutation__round_out[514]), .A2(
        _f_permutation__n7149 ), .ZN(_f_permutation__n3240 ) );
  NAND2_X2 _f_permutation__U2701  ( .A1(SYNOPSYS_UNCONNECTED_574), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3241 ) );
  NAND2_X2 _f_permutation__U2700  ( .A1(_f_permutation__n3240 ), .A2(
        _f_permutation__n3241 ), .ZN(_f_permutation__n4873 ) );
  NAND2_X2 _f_permutation__U2699  ( .A1(_f_permutation__round_out[513]), .A2(
        _f_permutation__n7148 ), .ZN(_f_permutation__n3238 ) );
  NAND2_X2 _f_permutation__U2698  ( .A1(SYNOPSYS_UNCONNECTED_575), .A2(
        _f_permutation__n7262 ), .ZN(_f_permutation__n3239 ) );
  NAND2_X2 _f_permutation__U2697  ( .A1(_f_permutation__n3238 ), .A2(
        _f_permutation__n3239 ), .ZN(_f_permutation__n4874 ) );
  NAND2_X2 _f_permutation__U2696  ( .A1(_f_permutation__round_out[512]), .A2(
        _f_permutation__n7147 ), .ZN(_f_permutation__n3236 ) );
  NAND2_X2 _f_permutation__U2695  ( .A1(SYNOPSYS_UNCONNECTED_576), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3237 ) );
  NAND2_X2 _f_permutation__U2694  ( .A1(_f_permutation__n3236 ), .A2(
        _f_permutation__n3237 ), .ZN(_f_permutation__n4875 ) );
  NAND2_X2 _f_permutation__U2693  ( .A1(_f_permutation__round_out[511]), .A2(
        _f_permutation__n7152 ), .ZN(_f_permutation__n3234 ) );
  NAND2_X2 _f_permutation__U2692  ( .A1(SYNOPSYS_UNCONNECTED_577), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3235 ) );
  NAND2_X2 _f_permutation__U2691  ( .A1(_f_permutation__n3234 ), .A2(
        _f_permutation__n3235 ), .ZN(_f_permutation__n4876 ) );
  NAND2_X2 _f_permutation__U2690  ( .A1(_f_permutation__round_out[510]), .A2(
        _f_permutation__n7151 ), .ZN(_f_permutation__n3232 ) );
  NAND2_X2 _f_permutation__U2689  ( .A1(SYNOPSYS_UNCONNECTED_578), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3233 ) );
  NAND2_X2 _f_permutation__U2688  ( .A1(_f_permutation__n3232 ), .A2(
        _f_permutation__n3233 ), .ZN(_f_permutation__n4877 ) );
  NAND2_X2 _f_permutation__U2687  ( .A1(_f_permutation__round_out[509]), .A2(
        _f_permutation__n7150 ), .ZN(_f_permutation__n3230 ) );
  NAND2_X2 _f_permutation__U2686  ( .A1(SYNOPSYS_UNCONNECTED_579), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3231 ) );
  NAND2_X2 _f_permutation__U2685  ( .A1(_f_permutation__n3230 ), .A2(
        _f_permutation__n3231 ), .ZN(_f_permutation__n4878 ) );
  NAND2_X2 _f_permutation__U2684  ( .A1(_f_permutation__round_out[508]), .A2(
        _f_permutation__n7141 ), .ZN(_f_permutation__n3228 ) );
  NAND2_X2 _f_permutation__U2683  ( .A1(SYNOPSYS_UNCONNECTED_580), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3229 ) );
  NAND2_X2 _f_permutation__U2682  ( .A1(_f_permutation__n3228 ), .A2(
        _f_permutation__n3229 ), .ZN(_f_permutation__n4879 ) );
  NAND2_X2 _f_permutation__U2681  ( .A1(_f_permutation__round_out[507]), .A2(
        _f_permutation__n7140 ), .ZN(_f_permutation__n3226 ) );
  NAND2_X2 _f_permutation__U2680  ( .A1(SYNOPSYS_UNCONNECTED_581), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3227 ) );
  NAND2_X2 _f_permutation__U2679  ( .A1(_f_permutation__n3226 ), .A2(
        _f_permutation__n3227 ), .ZN(_f_permutation__n4880 ) );
  NAND2_X2 _f_permutation__U2678  ( .A1(_f_permutation__round_out[506]), .A2(
        _f_permutation__n7139 ), .ZN(_f_permutation__n3224 ) );
  NAND2_X2 _f_permutation__U2677  ( .A1(SYNOPSYS_UNCONNECTED_582), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3225 ) );
  NAND2_X2 _f_permutation__U2676  ( .A1(_f_permutation__n3224 ), .A2(
        _f_permutation__n3225 ), .ZN(_f_permutation__n4881 ) );
  NAND2_X2 _f_permutation__U2675  ( .A1(_f_permutation__round_out[505]), .A2(
        _f_permutation__n7146 ), .ZN(_f_permutation__n3222 ) );
  NAND2_X2 _f_permutation__U2674  ( .A1(SYNOPSYS_UNCONNECTED_583), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3223 ) );
  NAND2_X2 _f_permutation__U2673  ( .A1(_f_permutation__n3222 ), .A2(
        _f_permutation__n3223 ), .ZN(_f_permutation__n4882 ) );
  NAND2_X2 _f_permutation__U2672  ( .A1(_f_permutation__round_out[504]), .A2(
        _f_permutation__n7145 ), .ZN(_f_permutation__n3220 ) );
  NAND2_X2 _f_permutation__U2671  ( .A1(SYNOPSYS_UNCONNECTED_584), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3221 ) );
  NAND2_X2 _f_permutation__U2670  ( .A1(_f_permutation__n3220 ), .A2(
        _f_permutation__n3221 ), .ZN(_f_permutation__n4883 ) );
  NAND2_X2 _f_permutation__U2669  ( .A1(_f_permutation__round_out[503]), .A2(
        _f_permutation__n7144 ), .ZN(_f_permutation__n3218 ) );
  NAND2_X2 _f_permutation__U2668  ( .A1(SYNOPSYS_UNCONNECTED_585), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3219 ) );
  NAND2_X2 _f_permutation__U2667  ( .A1(_f_permutation__n3218 ), .A2(
        _f_permutation__n3219 ), .ZN(_f_permutation__n4884 ) );
  NAND2_X2 _f_permutation__U2666  ( .A1(_f_permutation__round_out[502]), .A2(
        _f_permutation__n7143 ), .ZN(_f_permutation__n3216 ) );
  NAND2_X2 _f_permutation__U2665  ( .A1(SYNOPSYS_UNCONNECTED_586), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3217 ) );
  NAND2_X2 _f_permutation__U2664  ( .A1(_f_permutation__n3216 ), .A2(
        _f_permutation__n3217 ), .ZN(_f_permutation__n4885 ) );
  NAND2_X2 _f_permutation__U2663  ( .A1(_f_permutation__round_out[501]), .A2(
        _f_permutation__n7142 ), .ZN(_f_permutation__n3214 ) );
  NAND2_X2 _f_permutation__U2662  ( .A1(SYNOPSYS_UNCONNECTED_587), .A2(
        _f_permutation__n7263 ), .ZN(_f_permutation__n3215 ) );
  NAND2_X2 _f_permutation__U2661  ( .A1(_f_permutation__n3214 ), .A2(
        _f_permutation__n3215 ), .ZN(_f_permutation__n4886 ) );
  NAND2_X2 _f_permutation__U2660  ( .A1(_f_permutation__round_out[500]), .A2(
        _f_permutation__n7066 ), .ZN(_f_permutation__n3212 ) );
  NAND2_X2 _f_permutation__U2659  ( .A1(SYNOPSYS_UNCONNECTED_588), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3213 ) );
  NAND2_X2 _f_permutation__U2658  ( .A1(_f_permutation__n3212 ), .A2(
        _f_permutation__n3213 ), .ZN(_f_permutation__n4887 ) );
  NAND2_X2 _f_permutation__U2657  ( .A1(_f_permutation__round_out[499]), .A2(
        _f_permutation__n7168 ), .ZN(_f_permutation__n3210 ) );
  NAND2_X2 _f_permutation__U2656  ( .A1(SYNOPSYS_UNCONNECTED_589), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3211 ) );
  NAND2_X2 _f_permutation__U2655  ( .A1(_f_permutation__n3210 ), .A2(
        _f_permutation__n3211 ), .ZN(_f_permutation__n4888 ) );
  NAND2_X2 _f_permutation__U2654  ( .A1(_f_permutation__round_out[498]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n3208 ) );
  NAND2_X2 _f_permutation__U2653  ( .A1(SYNOPSYS_UNCONNECTED_590), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3209 ) );
  NAND2_X2 _f_permutation__U2652  ( .A1(_f_permutation__n3208 ), .A2(
        _f_permutation__n3209 ), .ZN(_f_permutation__n4889 ) );
  NAND2_X2 _f_permutation__U2651  ( .A1(_f_permutation__round_out[497]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n3206 ) );
  NAND2_X2 _f_permutation__U2650  ( .A1(SYNOPSYS_UNCONNECTED_591), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3207 ) );
  NAND2_X2 _f_permutation__U2649  ( .A1(_f_permutation__n3206 ), .A2(
        _f_permutation__n3207 ), .ZN(_f_permutation__n4890 ) );
  NAND2_X2 _f_permutation__U2648  ( .A1(_f_permutation__round_out[496]), .A2(
        _f_permutation__n7149 ), .ZN(_f_permutation__n3204 ) );
  NAND2_X2 _f_permutation__U2647  ( .A1(SYNOPSYS_UNCONNECTED_592), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3205 ) );
  NAND2_X2 _f_permutation__U2646  ( .A1(_f_permutation__n3204 ), .A2(
        _f_permutation__n3205 ), .ZN(_f_permutation__n4891 ) );
  NAND2_X2 _f_permutation__U2645  ( .A1(_f_permutation__round_out[495]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3202 ) );
  NAND2_X2 _f_permutation__U2644  ( .A1(SYNOPSYS_UNCONNECTED_593), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3203 ) );
  NAND2_X2 _f_permutation__U2643  ( .A1(_f_permutation__n3202 ), .A2(
        _f_permutation__n3203 ), .ZN(_f_permutation__n4892 ) );
  NAND2_X2 _f_permutation__U2642  ( .A1(_f_permutation__round_out[494]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3200 ) );
  NAND2_X2 _f_permutation__U2641  ( .A1(SYNOPSYS_UNCONNECTED_594), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3201 ) );
  NAND2_X2 _f_permutation__U2640  ( .A1(_f_permutation__n3200 ), .A2(
        _f_permutation__n3201 ), .ZN(_f_permutation__n4893 ) );
  NAND2_X2 _f_permutation__U2639  ( .A1(_f_permutation__round_out[493]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3198 ) );
  NAND2_X2 _f_permutation__U2638  ( .A1(SYNOPSYS_UNCONNECTED_595), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3199 ) );
  NAND2_X2 _f_permutation__U2637  ( .A1(_f_permutation__n3198 ), .A2(
        _f_permutation__n3199 ), .ZN(_f_permutation__n4894 ) );
  NAND2_X2 _f_permutation__U2636  ( .A1(_f_permutation__round_out[492]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3196 ) );
  NAND2_X2 _f_permutation__U2635  ( .A1(SYNOPSYS_UNCONNECTED_596), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3197 ) );
  NAND2_X2 _f_permutation__U2634  ( .A1(_f_permutation__n3196 ), .A2(
        _f_permutation__n3197 ), .ZN(_f_permutation__n4895 ) );
  NAND2_X2 _f_permutation__U2633  ( .A1(_f_permutation__round_out[491]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3194 ) );
  NAND2_X2 _f_permutation__U2632  ( .A1(SYNOPSYS_UNCONNECTED_597), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3195 ) );
  NAND2_X2 _f_permutation__U2631  ( .A1(_f_permutation__n3194 ), .A2(
        _f_permutation__n3195 ), .ZN(_f_permutation__n4896 ) );
  NAND2_X2 _f_permutation__U2630  ( .A1(_f_permutation__round_out[490]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3192 ) );
  NAND2_X2 _f_permutation__U2629  ( .A1(SYNOPSYS_UNCONNECTED_598), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3193 ) );
  NAND2_X2 _f_permutation__U2628  ( .A1(_f_permutation__n3192 ), .A2(
        _f_permutation__n3193 ), .ZN(_f_permutation__n4897 ) );
  NAND2_X2 _f_permutation__U2627  ( .A1(_f_permutation__round_out[489]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3190 ) );
  NAND2_X2 _f_permutation__U2626  ( .A1(SYNOPSYS_UNCONNECTED_599), .A2(
        _f_permutation__n7264 ), .ZN(_f_permutation__n3191 ) );
  NAND2_X2 _f_permutation__U2625  ( .A1(_f_permutation__n3190 ), .A2(
        _f_permutation__n3191 ), .ZN(_f_permutation__n4898 ) );
  NAND2_X2 _f_permutation__U2624  ( .A1(_f_permutation__round_out[488]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3188 ) );
  NAND2_X2 _f_permutation__U2623  ( .A1(SYNOPSYS_UNCONNECTED_600), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3189 ) );
  NAND2_X2 _f_permutation__U2622  ( .A1(_f_permutation__n3188 ), .A2(
        _f_permutation__n3189 ), .ZN(_f_permutation__n4899 ) );
  NAND2_X2 _f_permutation__U2621  ( .A1(_f_permutation__round_out[487]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3186 ) );
  NAND2_X2 _f_permutation__U2620  ( .A1(SYNOPSYS_UNCONNECTED_601), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3187 ) );
  NAND2_X2 _f_permutation__U2619  ( .A1(_f_permutation__n3186 ), .A2(
        _f_permutation__n3187 ), .ZN(_f_permutation__n4900 ) );
  NAND2_X2 _f_permutation__U2618  ( .A1(_f_permutation__round_out[486]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3184 ) );
  NAND2_X2 _f_permutation__U2617  ( .A1(SYNOPSYS_UNCONNECTED_602), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3185 ) );
  NAND2_X2 _f_permutation__U2616  ( .A1(_f_permutation__n3184 ), .A2(
        _f_permutation__n3185 ), .ZN(_f_permutation__n4901 ) );
  NAND2_X2 _f_permutation__U2615  ( .A1(_f_permutation__round_out[485]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3182 ) );
  NAND2_X2 _f_permutation__U2614  ( .A1(SYNOPSYS_UNCONNECTED_603), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3183 ) );
  NAND2_X2 _f_permutation__U2613  ( .A1(_f_permutation__n3182 ), .A2(
        _f_permutation__n3183 ), .ZN(_f_permutation__n4902 ) );
  NAND2_X2 _f_permutation__U2612  ( .A1(_f_permutation__round_out[484]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3180 ) );
  NAND2_X2 _f_permutation__U2611  ( .A1(SYNOPSYS_UNCONNECTED_604), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3181 ) );
  NAND2_X2 _f_permutation__U2610  ( .A1(_f_permutation__n3180 ), .A2(
        _f_permutation__n3181 ), .ZN(_f_permutation__n4903 ) );
  NAND2_X2 _f_permutation__U2609  ( .A1(_f_permutation__round_out[483]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3178 ) );
  NAND2_X2 _f_permutation__U2608  ( .A1(SYNOPSYS_UNCONNECTED_605), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3179 ) );
  NAND2_X2 _f_permutation__U2607  ( .A1(_f_permutation__n3178 ), .A2(
        _f_permutation__n3179 ), .ZN(_f_permutation__n4904 ) );
  NAND2_X2 _f_permutation__U2606  ( .A1(_f_permutation__round_out[482]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3176 ) );
  NAND2_X2 _f_permutation__U2605  ( .A1(SYNOPSYS_UNCONNECTED_606), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3177 ) );
  NAND2_X2 _f_permutation__U2604  ( .A1(_f_permutation__n3176 ), .A2(
        _f_permutation__n3177 ), .ZN(_f_permutation__n4905 ) );
  NAND2_X2 _f_permutation__U2603  ( .A1(_f_permutation__round_out[481]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3174 ) );
  NAND2_X2 _f_permutation__U2602  ( .A1(SYNOPSYS_UNCONNECTED_607), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3175 ) );
  NAND2_X2 _f_permutation__U2601  ( .A1(_f_permutation__n3174 ), .A2(
        _f_permutation__n3175 ), .ZN(_f_permutation__n4906 ) );
  NAND2_X2 _f_permutation__U2600  ( .A1(_f_permutation__round_out[480]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3172 ) );
  NAND2_X2 _f_permutation__U2599  ( .A1(SYNOPSYS_UNCONNECTED_608), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3173 ) );
  NAND2_X2 _f_permutation__U2598  ( .A1(_f_permutation__n3172 ), .A2(
        _f_permutation__n3173 ), .ZN(_f_permutation__n4907 ) );
  NAND2_X2 _f_permutation__U2597  ( .A1(_f_permutation__round_out[479]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3170 ) );
  NAND2_X2 _f_permutation__U2596  ( .A1(SYNOPSYS_UNCONNECTED_609), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3171 ) );
  NAND2_X2 _f_permutation__U2595  ( .A1(_f_permutation__n3170 ), .A2(
        _f_permutation__n3171 ), .ZN(_f_permutation__n4908 ) );
  NAND2_X2 _f_permutation__U2594  ( .A1(_f_permutation__round_out[478]), .A2(
        _f_permutation__n7074 ), .ZN(_f_permutation__n3168 ) );
  NAND2_X2 _f_permutation__U2593  ( .A1(SYNOPSYS_UNCONNECTED_610), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3169 ) );
  NAND2_X2 _f_permutation__U2592  ( .A1(_f_permutation__n3168 ), .A2(
        _f_permutation__n3169 ), .ZN(_f_permutation__n4909 ) );
  NAND2_X2 _f_permutation__U2591  ( .A1(_f_permutation__round_out[477]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3166 ) );
  NAND2_X2 _f_permutation__U2590  ( .A1(SYNOPSYS_UNCONNECTED_611), .A2(
        _f_permutation__n7265 ), .ZN(_f_permutation__n3167 ) );
  NAND2_X2 _f_permutation__U2589  ( .A1(_f_permutation__n3166 ), .A2(
        _f_permutation__n3167 ), .ZN(_f_permutation__n4910 ) );
  NAND2_X2 _f_permutation__U2588  ( .A1(_f_permutation__round_out[476]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3164 ) );
  NAND2_X2 _f_permutation__U2587  ( .A1(SYNOPSYS_UNCONNECTED_612), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3165 ) );
  NAND2_X2 _f_permutation__U2586  ( .A1(_f_permutation__n3164 ), .A2(
        _f_permutation__n3165 ), .ZN(_f_permutation__n4911 ) );
  NAND2_X2 _f_permutation__U2585  ( .A1(_f_permutation__round_out[475]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3162 ) );
  NAND2_X2 _f_permutation__U2584  ( .A1(SYNOPSYS_UNCONNECTED_613), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3163 ) );
  NAND2_X2 _f_permutation__U2583  ( .A1(_f_permutation__n3162 ), .A2(
        _f_permutation__n3163 ), .ZN(_f_permutation__n4912 ) );
  NAND2_X2 _f_permutation__U2582  ( .A1(_f_permutation__round_out[474]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3160 ) );
  NAND2_X2 _f_permutation__U2581  ( .A1(SYNOPSYS_UNCONNECTED_614), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3161 ) );
  NAND2_X2 _f_permutation__U2580  ( .A1(_f_permutation__n3160 ), .A2(
        _f_permutation__n3161 ), .ZN(_f_permutation__n4913 ) );
  NAND2_X2 _f_permutation__U2579  ( .A1(_f_permutation__round_out[473]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3158 ) );
  NAND2_X2 _f_permutation__U2578  ( .A1(SYNOPSYS_UNCONNECTED_615), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3159 ) );
  NAND2_X2 _f_permutation__U2577  ( .A1(_f_permutation__n3158 ), .A2(
        _f_permutation__n3159 ), .ZN(_f_permutation__n4914 ) );
  NAND2_X2 _f_permutation__U2576  ( .A1(_f_permutation__round_out[472]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3156 ) );
  NAND2_X2 _f_permutation__U2575  ( .A1(SYNOPSYS_UNCONNECTED_616), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3157 ) );
  NAND2_X2 _f_permutation__U2574  ( .A1(_f_permutation__n3156 ), .A2(
        _f_permutation__n3157 ), .ZN(_f_permutation__n4915 ) );
  NAND2_X2 _f_permutation__U2573  ( .A1(_f_permutation__round_out[471]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3154 ) );
  NAND2_X2 _f_permutation__U2572  ( .A1(SYNOPSYS_UNCONNECTED_617), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3155 ) );
  NAND2_X2 _f_permutation__U2571  ( .A1(_f_permutation__n3154 ), .A2(
        _f_permutation__n3155 ), .ZN(_f_permutation__n4916 ) );
  NAND2_X2 _f_permutation__U2570  ( .A1(_f_permutation__round_out[470]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3152 ) );
  NAND2_X2 _f_permutation__U2569  ( .A1(SYNOPSYS_UNCONNECTED_618), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3153 ) );
  NAND2_X2 _f_permutation__U2568  ( .A1(_f_permutation__n3152 ), .A2(
        _f_permutation__n3153 ), .ZN(_f_permutation__n4917 ) );
  NAND2_X2 _f_permutation__U2567  ( .A1(_f_permutation__round_out[469]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3150 ) );
  NAND2_X2 _f_permutation__U2566  ( .A1(SYNOPSYS_UNCONNECTED_619), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3151 ) );
  NAND2_X2 _f_permutation__U2565  ( .A1(_f_permutation__n3150 ), .A2(
        _f_permutation__n3151 ), .ZN(_f_permutation__n4918 ) );
  NAND2_X2 _f_permutation__U2564  ( .A1(_f_permutation__round_out[468]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3148 ) );
  NAND2_X2 _f_permutation__U2563  ( .A1(SYNOPSYS_UNCONNECTED_620), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3149 ) );
  NAND2_X2 _f_permutation__U2562  ( .A1(_f_permutation__n3148 ), .A2(
        _f_permutation__n3149 ), .ZN(_f_permutation__n4919 ) );
  NAND2_X2 _f_permutation__U2561  ( .A1(_f_permutation__round_out[467]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3146 ) );
  NAND2_X2 _f_permutation__U2560  ( .A1(SYNOPSYS_UNCONNECTED_621), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3147 ) );
  NAND2_X2 _f_permutation__U2559  ( .A1(_f_permutation__n3146 ), .A2(
        _f_permutation__n3147 ), .ZN(_f_permutation__n4920 ) );
  NAND2_X2 _f_permutation__U2558  ( .A1(_f_permutation__round_out[466]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3144 ) );
  NAND2_X2 _f_permutation__U2557  ( .A1(SYNOPSYS_UNCONNECTED_622), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3145 ) );
  NAND2_X2 _f_permutation__U2556  ( .A1(_f_permutation__n3144 ), .A2(
        _f_permutation__n3145 ), .ZN(_f_permutation__n4921 ) );
  NAND2_X2 _f_permutation__U2555  ( .A1(_f_permutation__round_out[465]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3142 ) );
  NAND2_X2 _f_permutation__U2554  ( .A1(SYNOPSYS_UNCONNECTED_623), .A2(
        _f_permutation__n7266 ), .ZN(_f_permutation__n3143 ) );
  NAND2_X2 _f_permutation__U2553  ( .A1(_f_permutation__n3142 ), .A2(
        _f_permutation__n3143 ), .ZN(_f_permutation__n4922 ) );
  NAND2_X2 _f_permutation__U2552  ( .A1(_f_permutation__round_out[464]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3140 ) );
  NAND2_X2 _f_permutation__U2551  ( .A1(SYNOPSYS_UNCONNECTED_624), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3141 ) );
  NAND2_X2 _f_permutation__U2550  ( .A1(_f_permutation__n3140 ), .A2(
        _f_permutation__n3141 ), .ZN(_f_permutation__n4923 ) );
  NAND2_X2 _f_permutation__U2549  ( .A1(_f_permutation__round_out[463]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3138 ) );
  NAND2_X2 _f_permutation__U2548  ( .A1(SYNOPSYS_UNCONNECTED_625), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3139 ) );
  NAND2_X2 _f_permutation__U2547  ( .A1(_f_permutation__n3138 ), .A2(
        _f_permutation__n3139 ), .ZN(_f_permutation__n4924 ) );
  NAND2_X2 _f_permutation__U2546  ( .A1(_f_permutation__round_out[462]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3136 ) );
  NAND2_X2 _f_permutation__U2545  ( .A1(SYNOPSYS_UNCONNECTED_626), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3137 ) );
  NAND2_X2 _f_permutation__U2544  ( .A1(_f_permutation__n3136 ), .A2(
        _f_permutation__n3137 ), .ZN(_f_permutation__n4925 ) );
  NAND2_X2 _f_permutation__U2543  ( .A1(_f_permutation__round_out[461]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3134 ) );
  NAND2_X2 _f_permutation__U2542  ( .A1(SYNOPSYS_UNCONNECTED_627), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3135 ) );
  NAND2_X2 _f_permutation__U2541  ( .A1(_f_permutation__n3134 ), .A2(
        _f_permutation__n3135 ), .ZN(_f_permutation__n4926 ) );
  NAND2_X2 _f_permutation__U2540  ( .A1(_f_permutation__round_out[460]), .A2(
        _f_permutation__n7073 ), .ZN(_f_permutation__n3132 ) );
  NAND2_X2 _f_permutation__U2539  ( .A1(SYNOPSYS_UNCONNECTED_628), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3133 ) );
  NAND2_X2 _f_permutation__U2538  ( .A1(_f_permutation__n3132 ), .A2(
        _f_permutation__n3133 ), .ZN(_f_permutation__n4927 ) );
  NAND2_X2 _f_permutation__U2537  ( .A1(_f_permutation__round_out[459]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3130 ) );
  NAND2_X2 _f_permutation__U2536  ( .A1(SYNOPSYS_UNCONNECTED_629), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3131 ) );
  NAND2_X2 _f_permutation__U2535  ( .A1(_f_permutation__n3130 ), .A2(
        _f_permutation__n3131 ), .ZN(_f_permutation__n4928 ) );
  NAND2_X2 _f_permutation__U2534  ( .A1(_f_permutation__round_out[458]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3128 ) );
  NAND2_X2 _f_permutation__U2533  ( .A1(SYNOPSYS_UNCONNECTED_630), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3129 ) );
  NAND2_X2 _f_permutation__U2532  ( .A1(_f_permutation__n3128 ), .A2(
        _f_permutation__n3129 ), .ZN(_f_permutation__n4929 ) );
  NAND2_X2 _f_permutation__U2531  ( .A1(_f_permutation__round_out[457]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3126 ) );
  NAND2_X2 _f_permutation__U2530  ( .A1(SYNOPSYS_UNCONNECTED_631), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3127 ) );
  NAND2_X2 _f_permutation__U2529  ( .A1(_f_permutation__n3126 ), .A2(
        _f_permutation__n3127 ), .ZN(_f_permutation__n4930 ) );
  NAND2_X2 _f_permutation__U2528  ( .A1(_f_permutation__round_out[456]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3124 ) );
  NAND2_X2 _f_permutation__U2527  ( .A1(SYNOPSYS_UNCONNECTED_632), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3125 ) );
  NAND2_X2 _f_permutation__U2526  ( .A1(_f_permutation__n3124 ), .A2(
        _f_permutation__n3125 ), .ZN(_f_permutation__n4931 ) );
  NAND2_X2 _f_permutation__U2525  ( .A1(_f_permutation__round_out[455]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3122 ) );
  NAND2_X2 _f_permutation__U2524  ( .A1(SYNOPSYS_UNCONNECTED_633), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3123 ) );
  NAND2_X2 _f_permutation__U2523  ( .A1(_f_permutation__n3122 ), .A2(
        _f_permutation__n3123 ), .ZN(_f_permutation__n4932 ) );
  NAND2_X2 _f_permutation__U2522  ( .A1(_f_permutation__round_out[454]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3120 ) );
  NAND2_X2 _f_permutation__U2521  ( .A1(SYNOPSYS_UNCONNECTED_634), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3121 ) );
  NAND2_X2 _f_permutation__U2520  ( .A1(_f_permutation__n3120 ), .A2(
        _f_permutation__n3121 ), .ZN(_f_permutation__n4933 ) );
  NAND2_X2 _f_permutation__U2519  ( .A1(_f_permutation__round_out[453]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3118 ) );
  NAND2_X2 _f_permutation__U2518  ( .A1(SYNOPSYS_UNCONNECTED_635), .A2(
        _f_permutation__n7267 ), .ZN(_f_permutation__n3119 ) );
  NAND2_X2 _f_permutation__U2517  ( .A1(_f_permutation__n3118 ), .A2(
        _f_permutation__n3119 ), .ZN(_f_permutation__n4934 ) );
  NAND2_X2 _f_permutation__U2516  ( .A1(_f_permutation__round_out[452]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3116 ) );
  NAND2_X2 _f_permutation__U2515  ( .A1(SYNOPSYS_UNCONNECTED_636), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3117 ) );
  NAND2_X2 _f_permutation__U2514  ( .A1(_f_permutation__n3116 ), .A2(
        _f_permutation__n3117 ), .ZN(_f_permutation__n4935 ) );
  NAND2_X2 _f_permutation__U2513  ( .A1(_f_permutation__round_out[451]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3114 ) );
  NAND2_X2 _f_permutation__U2512  ( .A1(SYNOPSYS_UNCONNECTED_637), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3115 ) );
  NAND2_X2 _f_permutation__U2511  ( .A1(_f_permutation__n3114 ), .A2(
        _f_permutation__n3115 ), .ZN(_f_permutation__n4936 ) );
  NAND2_X2 _f_permutation__U2510  ( .A1(_f_permutation__round_out[450]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3112 ) );
  NAND2_X2 _f_permutation__U2509  ( .A1(SYNOPSYS_UNCONNECTED_638), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3113 ) );
  NAND2_X2 _f_permutation__U2508  ( .A1(_f_permutation__n3112 ), .A2(
        _f_permutation__n3113 ), .ZN(_f_permutation__n4937 ) );
  NAND2_X2 _f_permutation__U2507  ( .A1(_f_permutation__round_out[449]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3110 ) );
  NAND2_X2 _f_permutation__U2506  ( .A1(SYNOPSYS_UNCONNECTED_639), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3111 ) );
  NAND2_X2 _f_permutation__U2505  ( .A1(_f_permutation__n3110 ), .A2(
        _f_permutation__n3111 ), .ZN(_f_permutation__n4938 ) );
  NAND2_X2 _f_permutation__U2504  ( .A1(_f_permutation__round_out[448]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3108 ) );
  NAND2_X2 _f_permutation__U2503  ( .A1(SYNOPSYS_UNCONNECTED_640), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3109 ) );
  NAND2_X2 _f_permutation__U2502  ( .A1(_f_permutation__n3108 ), .A2(
        _f_permutation__n3109 ), .ZN(_f_permutation__n4939 ) );
  NAND2_X2 _f_permutation__U2501  ( .A1(_f_permutation__round_out[447]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3106 ) );
  NAND2_X2 _f_permutation__U2500  ( .A1(SYNOPSYS_UNCONNECTED_641), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3107 ) );
  NAND2_X2 _f_permutation__U2499  ( .A1(_f_permutation__n3106 ), .A2(
        _f_permutation__n3107 ), .ZN(_f_permutation__n4940 ) );
  NAND2_X2 _f_permutation__U2498  ( .A1(_f_permutation__round_out[446]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3104 ) );
  NAND2_X2 _f_permutation__U2497  ( .A1(SYNOPSYS_UNCONNECTED_642), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3105 ) );
  NAND2_X2 _f_permutation__U2496  ( .A1(_f_permutation__n3104 ), .A2(
        _f_permutation__n3105 ), .ZN(_f_permutation__n4941 ) );
  NAND2_X2 _f_permutation__U2495  ( .A1(_f_permutation__round_out[445]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3102 ) );
  NAND2_X2 _f_permutation__U2494  ( .A1(SYNOPSYS_UNCONNECTED_643), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3103 ) );
  NAND2_X2 _f_permutation__U2493  ( .A1(_f_permutation__n3102 ), .A2(
        _f_permutation__n3103 ), .ZN(_f_permutation__n4942 ) );
  NAND2_X2 _f_permutation__U2492  ( .A1(_f_permutation__round_out[444]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3100 ) );
  NAND2_X2 _f_permutation__U2491  ( .A1(SYNOPSYS_UNCONNECTED_644), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3101 ) );
  NAND2_X2 _f_permutation__U2490  ( .A1(_f_permutation__n3100 ), .A2(
        _f_permutation__n3101 ), .ZN(_f_permutation__n4943 ) );
  NAND2_X2 _f_permutation__U2489  ( .A1(_f_permutation__round_out[443]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3098 ) );
  NAND2_X2 _f_permutation__U2488  ( .A1(SYNOPSYS_UNCONNECTED_645), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3099 ) );
  NAND2_X2 _f_permutation__U2487  ( .A1(_f_permutation__n3098 ), .A2(
        _f_permutation__n3099 ), .ZN(_f_permutation__n4944 ) );
  NAND2_X2 _f_permutation__U2486  ( .A1(_f_permutation__round_out[442]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3096 ) );
  NAND2_X2 _f_permutation__U2485  ( .A1(SYNOPSYS_UNCONNECTED_646), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3097 ) );
  NAND2_X2 _f_permutation__U2484  ( .A1(_f_permutation__n3096 ), .A2(
        _f_permutation__n3097 ), .ZN(_f_permutation__n4945 ) );
  NAND2_X2 _f_permutation__U2483  ( .A1(_f_permutation__round_out[441]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3094 ) );
  NAND2_X2 _f_permutation__U2482  ( .A1(SYNOPSYS_UNCONNECTED_647), .A2(
        _f_permutation__n7268 ), .ZN(_f_permutation__n3095 ) );
  NAND2_X2 _f_permutation__U2481  ( .A1(_f_permutation__n3094 ), .A2(
        _f_permutation__n3095 ), .ZN(_f_permutation__n4946 ) );
  NAND2_X2 _f_permutation__U2480  ( .A1(_f_permutation__round_out[440]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3092 ) );
  NAND2_X2 _f_permutation__U2479  ( .A1(SYNOPSYS_UNCONNECTED_648), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3093 ) );
  NAND2_X2 _f_permutation__U2478  ( .A1(_f_permutation__n3092 ), .A2(
        _f_permutation__n3093 ), .ZN(_f_permutation__n4947 ) );
  NAND2_X2 _f_permutation__U2477  ( .A1(_f_permutation__round_out[439]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3090 ) );
  NAND2_X2 _f_permutation__U2476  ( .A1(SYNOPSYS_UNCONNECTED_649), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3091 ) );
  NAND2_X2 _f_permutation__U2475  ( .A1(_f_permutation__n3090 ), .A2(
        _f_permutation__n3091 ), .ZN(_f_permutation__n4948 ) );
  NAND2_X2 _f_permutation__U2474  ( .A1(_f_permutation__round_out[438]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3088 ) );
  NAND2_X2 _f_permutation__U2473  ( .A1(SYNOPSYS_UNCONNECTED_650), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3089 ) );
  NAND2_X2 _f_permutation__U2472  ( .A1(_f_permutation__n3088 ), .A2(
        _f_permutation__n3089 ), .ZN(_f_permutation__n4949 ) );
  NAND2_X2 _f_permutation__U2471  ( .A1(_f_permutation__round_out[437]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3086 ) );
  NAND2_X2 _f_permutation__U2470  ( .A1(SYNOPSYS_UNCONNECTED_651), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3087 ) );
  NAND2_X2 _f_permutation__U2469  ( .A1(_f_permutation__n3086 ), .A2(
        _f_permutation__n3087 ), .ZN(_f_permutation__n4950 ) );
  NAND2_X2 _f_permutation__U2468  ( .A1(_f_permutation__round_out[436]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3084 ) );
  NAND2_X2 _f_permutation__U2467  ( .A1(SYNOPSYS_UNCONNECTED_652), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3085 ) );
  NAND2_X2 _f_permutation__U2466  ( .A1(_f_permutation__n3084 ), .A2(
        _f_permutation__n3085 ), .ZN(_f_permutation__n4951 ) );
  NAND2_X2 _f_permutation__U2465  ( .A1(_f_permutation__round_out[435]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3082 ) );
  NAND2_X2 _f_permutation__U2464  ( .A1(SYNOPSYS_UNCONNECTED_653), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3083 ) );
  NAND2_X2 _f_permutation__U2463  ( .A1(_f_permutation__n3082 ), .A2(
        _f_permutation__n3083 ), .ZN(_f_permutation__n4952 ) );
  NAND2_X2 _f_permutation__U2462  ( .A1(_f_permutation__round_out[434]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3080 ) );
  NAND2_X2 _f_permutation__U2461  ( .A1(SYNOPSYS_UNCONNECTED_654), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3081 ) );
  NAND2_X2 _f_permutation__U2460  ( .A1(_f_permutation__n3080 ), .A2(
        _f_permutation__n3081 ), .ZN(_f_permutation__n4953 ) );
  NAND2_X2 _f_permutation__U2459  ( .A1(_f_permutation__round_out[433]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3078 ) );
  NAND2_X2 _f_permutation__U2458  ( .A1(SYNOPSYS_UNCONNECTED_655), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3079 ) );
  NAND2_X2 _f_permutation__U2457  ( .A1(_f_permutation__n3078 ), .A2(
        _f_permutation__n3079 ), .ZN(_f_permutation__n4954 ) );
  NAND2_X2 _f_permutation__U2456  ( .A1(_f_permutation__round_out[432]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3076 ) );
  NAND2_X2 _f_permutation__U2455  ( .A1(SYNOPSYS_UNCONNECTED_656), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3077 ) );
  NAND2_X2 _f_permutation__U2454  ( .A1(_f_permutation__n3076 ), .A2(
        _f_permutation__n3077 ), .ZN(_f_permutation__n4955 ) );
  NAND2_X2 _f_permutation__U2453  ( .A1(_f_permutation__round_out[431]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3074 ) );
  NAND2_X2 _f_permutation__U2452  ( .A1(SYNOPSYS_UNCONNECTED_657), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3075 ) );
  NAND2_X2 _f_permutation__U2451  ( .A1(_f_permutation__n3074 ), .A2(
        _f_permutation__n3075 ), .ZN(_f_permutation__n4956 ) );
  NAND2_X2 _f_permutation__U2450  ( .A1(_f_permutation__round_out[430]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3072 ) );
  NAND2_X2 _f_permutation__U2449  ( .A1(SYNOPSYS_UNCONNECTED_658), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3073 ) );
  NAND2_X2 _f_permutation__U2448  ( .A1(_f_permutation__n3072 ), .A2(
        _f_permutation__n3073 ), .ZN(_f_permutation__n4957 ) );
  NAND2_X2 _f_permutation__U2447  ( .A1(_f_permutation__round_out[429]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3070 ) );
  NAND2_X2 _f_permutation__U2446  ( .A1(SYNOPSYS_UNCONNECTED_659), .A2(
        _f_permutation__n7269 ), .ZN(_f_permutation__n3071 ) );
  NAND2_X2 _f_permutation__U2445  ( .A1(_f_permutation__n3070 ), .A2(
        _f_permutation__n3071 ), .ZN(_f_permutation__n4958 ) );
  NAND2_X2 _f_permutation__U2444  ( .A1(_f_permutation__round_out[428]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3068 ) );
  NAND2_X2 _f_permutation__U2443  ( .A1(SYNOPSYS_UNCONNECTED_660), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3069 ) );
  NAND2_X2 _f_permutation__U2442  ( .A1(_f_permutation__n3068 ), .A2(
        _f_permutation__n3069 ), .ZN(_f_permutation__n4959 ) );
  NAND2_X2 _f_permutation__U2441  ( .A1(_f_permutation__round_out[427]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3066 ) );
  NAND2_X2 _f_permutation__U2440  ( .A1(SYNOPSYS_UNCONNECTED_661), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3067 ) );
  NAND2_X2 _f_permutation__U2439  ( .A1(_f_permutation__n3066 ), .A2(
        _f_permutation__n3067 ), .ZN(_f_permutation__n4960 ) );
  NAND2_X2 _f_permutation__U2438  ( .A1(_f_permutation__round_out[426]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3064 ) );
  NAND2_X2 _f_permutation__U2437  ( .A1(SYNOPSYS_UNCONNECTED_662), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3065 ) );
  NAND2_X2 _f_permutation__U2436  ( .A1(_f_permutation__n3064 ), .A2(
        _f_permutation__n3065 ), .ZN(_f_permutation__n4961 ) );
  NAND2_X2 _f_permutation__U2435  ( .A1(_f_permutation__round_out[425]), .A2(
        _f_permutation__n7071 ), .ZN(_f_permutation__n3062 ) );
  NAND2_X2 _f_permutation__U2434  ( .A1(SYNOPSYS_UNCONNECTED_663), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3063 ) );
  NAND2_X2 _f_permutation__U2433  ( .A1(_f_permutation__n3062 ), .A2(
        _f_permutation__n3063 ), .ZN(_f_permutation__n4962 ) );
  NAND2_X2 _f_permutation__U2432  ( .A1(_f_permutation__round_out[424]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3060 ) );
  NAND2_X2 _f_permutation__U2431  ( .A1(SYNOPSYS_UNCONNECTED_664), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3061 ) );
  NAND2_X2 _f_permutation__U2430  ( .A1(_f_permutation__n3060 ), .A2(
        _f_permutation__n3061 ), .ZN(_f_permutation__n4963 ) );
  NAND2_X2 _f_permutation__U2429  ( .A1(_f_permutation__round_out[423]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3058 ) );
  NAND2_X2 _f_permutation__U2428  ( .A1(SYNOPSYS_UNCONNECTED_665), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3059 ) );
  NAND2_X2 _f_permutation__U2427  ( .A1(_f_permutation__n3058 ), .A2(
        _f_permutation__n3059 ), .ZN(_f_permutation__n4964 ) );
  NAND2_X2 _f_permutation__U2426  ( .A1(_f_permutation__round_out[422]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3056 ) );
  NAND2_X2 _f_permutation__U2425  ( .A1(SYNOPSYS_UNCONNECTED_666), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3057 ) );
  NAND2_X2 _f_permutation__U2424  ( .A1(_f_permutation__n3056 ), .A2(
        _f_permutation__n3057 ), .ZN(_f_permutation__n4965 ) );
  NAND2_X2 _f_permutation__U2423  ( .A1(_f_permutation__round_out[421]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3054 ) );
  NAND2_X2 _f_permutation__U2422  ( .A1(SYNOPSYS_UNCONNECTED_667), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3055 ) );
  NAND2_X2 _f_permutation__U2421  ( .A1(_f_permutation__n3054 ), .A2(
        _f_permutation__n3055 ), .ZN(_f_permutation__n4966 ) );
  NAND2_X2 _f_permutation__U2420  ( .A1(_f_permutation__round_out[420]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3052 ) );
  NAND2_X2 _f_permutation__U2419  ( .A1(SYNOPSYS_UNCONNECTED_668), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3053 ) );
  NAND2_X2 _f_permutation__U2418  ( .A1(_f_permutation__n3052 ), .A2(
        _f_permutation__n3053 ), .ZN(_f_permutation__n4967 ) );
  NAND2_X2 _f_permutation__U2417  ( .A1(_f_permutation__round_out[419]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3050 ) );
  NAND2_X2 _f_permutation__U2416  ( .A1(SYNOPSYS_UNCONNECTED_669), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3051 ) );
  NAND2_X2 _f_permutation__U2415  ( .A1(_f_permutation__n3050 ), .A2(
        _f_permutation__n3051 ), .ZN(_f_permutation__n4968 ) );
  NAND2_X2 _f_permutation__U2414  ( .A1(_f_permutation__round_out[418]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3048 ) );
  NAND2_X2 _f_permutation__U2413  ( .A1(SYNOPSYS_UNCONNECTED_670), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3049 ) );
  NAND2_X2 _f_permutation__U2412  ( .A1(_f_permutation__n3048 ), .A2(
        _f_permutation__n3049 ), .ZN(_f_permutation__n4969 ) );
  NAND2_X2 _f_permutation__U2411  ( .A1(_f_permutation__round_out[417]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3046 ) );
  NAND2_X2 _f_permutation__U2410  ( .A1(SYNOPSYS_UNCONNECTED_671), .A2(
        _f_permutation__n7270 ), .ZN(_f_permutation__n3047 ) );
  NAND2_X2 _f_permutation__U2409  ( .A1(_f_permutation__n3046 ), .A2(
        _f_permutation__n3047 ), .ZN(_f_permutation__n4970 ) );
  NAND2_X2 _f_permutation__U2408  ( .A1(_f_permutation__round_out[416]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3044 ) );
  NAND2_X2 _f_permutation__U2407  ( .A1(SYNOPSYS_UNCONNECTED_672), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3045 ) );
  NAND2_X2 _f_permutation__U2406  ( .A1(_f_permutation__n3044 ), .A2(
        _f_permutation__n3045 ), .ZN(_f_permutation__n4971 ) );
  NAND2_X2 _f_permutation__U2405  ( .A1(_f_permutation__round_out[415]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3042 ) );
  NAND2_X2 _f_permutation__U2404  ( .A1(SYNOPSYS_UNCONNECTED_673), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3043 ) );
  NAND2_X2 _f_permutation__U2403  ( .A1(_f_permutation__n3042 ), .A2(
        _f_permutation__n3043 ), .ZN(_f_permutation__n4972 ) );
  NAND2_X2 _f_permutation__U2402  ( .A1(_f_permutation__round_out[414]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3040 ) );
  NAND2_X2 _f_permutation__U2401  ( .A1(SYNOPSYS_UNCONNECTED_674), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3041 ) );
  NAND2_X2 _f_permutation__U2400  ( .A1(_f_permutation__n3040 ), .A2(
        _f_permutation__n3041 ), .ZN(_f_permutation__n4973 ) );
  NAND2_X2 _f_permutation__U2399  ( .A1(_f_permutation__round_out[413]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3038 ) );
  NAND2_X2 _f_permutation__U2398  ( .A1(SYNOPSYS_UNCONNECTED_675), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3039 ) );
  NAND2_X2 _f_permutation__U2397  ( .A1(_f_permutation__n3038 ), .A2(
        _f_permutation__n3039 ), .ZN(_f_permutation__n4974 ) );
  NAND2_X2 _f_permutation__U2396  ( .A1(_f_permutation__round_out[412]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3036 ) );
  NAND2_X2 _f_permutation__U2395  ( .A1(SYNOPSYS_UNCONNECTED_676), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3037 ) );
  NAND2_X2 _f_permutation__U2394  ( .A1(_f_permutation__n3036 ), .A2(
        _f_permutation__n3037 ), .ZN(_f_permutation__n4975 ) );
  NAND2_X2 _f_permutation__U2393  ( .A1(_f_permutation__round_out[411]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3034 ) );
  NAND2_X2 _f_permutation__U2392  ( .A1(SYNOPSYS_UNCONNECTED_677), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3035 ) );
  NAND2_X2 _f_permutation__U2391  ( .A1(_f_permutation__n3034 ), .A2(
        _f_permutation__n3035 ), .ZN(_f_permutation__n4976 ) );
  NAND2_X2 _f_permutation__U2390  ( .A1(_f_permutation__round_out[410]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3032 ) );
  NAND2_X2 _f_permutation__U2389  ( .A1(SYNOPSYS_UNCONNECTED_678), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3033 ) );
  NAND2_X2 _f_permutation__U2388  ( .A1(_f_permutation__n3032 ), .A2(
        _f_permutation__n3033 ), .ZN(_f_permutation__n4977 ) );
  NAND2_X2 _f_permutation__U2387  ( .A1(_f_permutation__round_out[409]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3030 ) );
  NAND2_X2 _f_permutation__U2386  ( .A1(SYNOPSYS_UNCONNECTED_679), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3031 ) );
  NAND2_X2 _f_permutation__U2385  ( .A1(_f_permutation__n3030 ), .A2(
        _f_permutation__n3031 ), .ZN(_f_permutation__n4978 ) );
  NAND2_X2 _f_permutation__U2384  ( .A1(_f_permutation__round_out[408]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3028 ) );
  NAND2_X2 _f_permutation__U2383  ( .A1(SYNOPSYS_UNCONNECTED_680), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3029 ) );
  NAND2_X2 _f_permutation__U2382  ( .A1(_f_permutation__n3028 ), .A2(
        _f_permutation__n3029 ), .ZN(_f_permutation__n4979 ) );
  NAND2_X2 _f_permutation__U2381  ( .A1(_f_permutation__round_out[407]), .A2(
        _f_permutation__n7070 ), .ZN(_f_permutation__n3026 ) );
  NAND2_X2 _f_permutation__U2380  ( .A1(SYNOPSYS_UNCONNECTED_681), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3027 ) );
  NAND2_X2 _f_permutation__U2379  ( .A1(_f_permutation__n3026 ), .A2(
        _f_permutation__n3027 ), .ZN(_f_permutation__n4980 ) );
  NAND2_X2 _f_permutation__U2378  ( .A1(_f_permutation__round_out[406]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3024 ) );
  NAND2_X2 _f_permutation__U2377  ( .A1(SYNOPSYS_UNCONNECTED_682), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3025 ) );
  NAND2_X2 _f_permutation__U2376  ( .A1(_f_permutation__n3024 ), .A2(
        _f_permutation__n3025 ), .ZN(_f_permutation__n4981 ) );
  NAND2_X2 _f_permutation__U2375  ( .A1(_f_permutation__round_out[405]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3022 ) );
  NAND2_X2 _f_permutation__U2374  ( .A1(SYNOPSYS_UNCONNECTED_683), .A2(
        _f_permutation__n7271 ), .ZN(_f_permutation__n3023 ) );
  NAND2_X2 _f_permutation__U2373  ( .A1(_f_permutation__n3022 ), .A2(
        _f_permutation__n3023 ), .ZN(_f_permutation__n4982 ) );
  NAND2_X2 _f_permutation__U2372  ( .A1(_f_permutation__round_out[404]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3020 ) );
  NAND2_X2 _f_permutation__U2371  ( .A1(SYNOPSYS_UNCONNECTED_684), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3021 ) );
  NAND2_X2 _f_permutation__U2370  ( .A1(_f_permutation__n3020 ), .A2(
        _f_permutation__n3021 ), .ZN(_f_permutation__n4983 ) );
  NAND2_X2 _f_permutation__U2369  ( .A1(_f_permutation__round_out[403]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3018 ) );
  NAND2_X2 _f_permutation__U2368  ( .A1(SYNOPSYS_UNCONNECTED_685), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3019 ) );
  NAND2_X2 _f_permutation__U2367  ( .A1(_f_permutation__n3018 ), .A2(
        _f_permutation__n3019 ), .ZN(_f_permutation__n4984 ) );
  NAND2_X2 _f_permutation__U2366  ( .A1(_f_permutation__round_out[402]), .A2(
        _f_permutation__n7069 ), .ZN(_f_permutation__n3016 ) );
  NAND2_X2 _f_permutation__U2365  ( .A1(SYNOPSYS_UNCONNECTED_686), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3017 ) );
  NAND2_X2 _f_permutation__U2364  ( .A1(_f_permutation__n3016 ), .A2(
        _f_permutation__n3017 ), .ZN(_f_permutation__n4985 ) );
  NAND2_X2 _f_permutation__U2363  ( .A1(_f_permutation__round_out[401]), .A2(
        _f_permutation__n7072 ), .ZN(_f_permutation__n3014 ) );
  NAND2_X2 _f_permutation__U2362  ( .A1(SYNOPSYS_UNCONNECTED_687), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3015 ) );
  NAND2_X2 _f_permutation__U2361  ( .A1(_f_permutation__n3014 ), .A2(
        _f_permutation__n3015 ), .ZN(_f_permutation__n4986 ) );
  NAND2_X2 _f_permutation__U2360  ( .A1(_f_permutation__round_out[400]), .A2(
        _f_permutation__n7164 ), .ZN(_f_permutation__n3012 ) );
  NAND2_X2 _f_permutation__U2359  ( .A1(SYNOPSYS_UNCONNECTED_688), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3013 ) );
  NAND2_X2 _f_permutation__U2358  ( .A1(_f_permutation__n3012 ), .A2(
        _f_permutation__n3013 ), .ZN(_f_permutation__n4987 ) );
  NAND2_X2 _f_permutation__U2357  ( .A1(_f_permutation__round_out[399]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n3010 ) );
  NAND2_X2 _f_permutation__U2356  ( .A1(SYNOPSYS_UNCONNECTED_689), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3011 ) );
  NAND2_X2 _f_permutation__U2355  ( .A1(_f_permutation__n3010 ), .A2(
        _f_permutation__n3011 ), .ZN(_f_permutation__n4988 ) );
  NAND2_X2 _f_permutation__U2354  ( .A1(_f_permutation__round_out[398]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n3008 ) );
  NAND2_X2 _f_permutation__U2353  ( .A1(SYNOPSYS_UNCONNECTED_690), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3009 ) );
  NAND2_X2 _f_permutation__U2352  ( .A1(_f_permutation__n3008 ), .A2(
        _f_permutation__n3009 ), .ZN(_f_permutation__n4989 ) );
  NAND2_X2 _f_permutation__U2351  ( .A1(_f_permutation__round_out[397]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n3006 ) );
  NAND2_X2 _f_permutation__U2350  ( .A1(SYNOPSYS_UNCONNECTED_691), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3007 ) );
  NAND2_X2 _f_permutation__U2349  ( .A1(_f_permutation__n3006 ), .A2(
        _f_permutation__n3007 ), .ZN(_f_permutation__n4990 ) );
  NAND2_X2 _f_permutation__U2348  ( .A1(_f_permutation__round_out[396]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n3004 ) );
  NAND2_X2 _f_permutation__U2347  ( .A1(SYNOPSYS_UNCONNECTED_692), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3005 ) );
  NAND2_X2 _f_permutation__U2346  ( .A1(_f_permutation__n3004 ), .A2(
        _f_permutation__n3005 ), .ZN(_f_permutation__n4991 ) );
  NAND2_X2 _f_permutation__U2345  ( .A1(_f_permutation__round_out[395]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n3002 ) );
  NAND2_X2 _f_permutation__U2344  ( .A1(SYNOPSYS_UNCONNECTED_693), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3003 ) );
  NAND2_X2 _f_permutation__U2343  ( .A1(_f_permutation__n3002 ), .A2(
        _f_permutation__n3003 ), .ZN(_f_permutation__n4992 ) );
  NAND2_X2 _f_permutation__U2342  ( .A1(_f_permutation__round_out[394]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n3000 ) );
  NAND2_X2 _f_permutation__U2341  ( .A1(SYNOPSYS_UNCONNECTED_694), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n3001 ) );
  NAND2_X2 _f_permutation__U2340  ( .A1(_f_permutation__n3000 ), .A2(
        _f_permutation__n3001 ), .ZN(_f_permutation__n4993 ) );
  NAND2_X2 _f_permutation__U2339  ( .A1(_f_permutation__round_out[393]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2998 ) );
  NAND2_X2 _f_permutation__U2338  ( .A1(SYNOPSYS_UNCONNECTED_695), .A2(
        _f_permutation__n7272 ), .ZN(_f_permutation__n2999 ) );
  NAND2_X2 _f_permutation__U2337  ( .A1(_f_permutation__n2998 ), .A2(
        _f_permutation__n2999 ), .ZN(_f_permutation__n4994 ) );
  NAND2_X2 _f_permutation__U2336  ( .A1(_f_permutation__round_out[392]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2996 ) );
  NAND2_X2 _f_permutation__U2335  ( .A1(SYNOPSYS_UNCONNECTED_696), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2997 ) );
  NAND2_X2 _f_permutation__U2334  ( .A1(_f_permutation__n2996 ), .A2(
        _f_permutation__n2997 ), .ZN(_f_permutation__n4995 ) );
  NAND2_X2 _f_permutation__U2333  ( .A1(_f_permutation__round_out[391]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2994 ) );
  NAND2_X2 _f_permutation__U2332  ( .A1(SYNOPSYS_UNCONNECTED_697), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2995 ) );
  NAND2_X2 _f_permutation__U2331  ( .A1(_f_permutation__n2994 ), .A2(
        _f_permutation__n2995 ), .ZN(_f_permutation__n4996 ) );
  NAND2_X2 _f_permutation__U2330  ( .A1(_f_permutation__round_out[390]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2992 ) );
  NAND2_X2 _f_permutation__U2329  ( .A1(SYNOPSYS_UNCONNECTED_698), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2993 ) );
  NAND2_X2 _f_permutation__U2328  ( .A1(_f_permutation__n2992 ), .A2(
        _f_permutation__n2993 ), .ZN(_f_permutation__n4997 ) );
  NAND2_X2 _f_permutation__U2327  ( .A1(_f_permutation__round_out[389]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2990 ) );
  NAND2_X2 _f_permutation__U2326  ( .A1(SYNOPSYS_UNCONNECTED_699), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2991 ) );
  NAND2_X2 _f_permutation__U2325  ( .A1(_f_permutation__n2990 ), .A2(
        _f_permutation__n2991 ), .ZN(_f_permutation__n4998 ) );
  NAND2_X2 _f_permutation__U2324  ( .A1(_f_permutation__round_out[388]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2988 ) );
  NAND2_X2 _f_permutation__U2323  ( .A1(SYNOPSYS_UNCONNECTED_700), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2989 ) );
  NAND2_X2 _f_permutation__U2322  ( .A1(_f_permutation__n2988 ), .A2(
        _f_permutation__n2989 ), .ZN(_f_permutation__n4999 ) );
  NAND2_X2 _f_permutation__U2321  ( .A1(_f_permutation__round_out[387]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2986 ) );
  NAND2_X2 _f_permutation__U2320  ( .A1(SYNOPSYS_UNCONNECTED_701), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2987 ) );
  NAND2_X2 _f_permutation__U2319  ( .A1(_f_permutation__n2986 ), .A2(
        _f_permutation__n2987 ), .ZN(_f_permutation__n5000 ) );
  NAND2_X2 _f_permutation__U2318  ( .A1(_f_permutation__round_out[386]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2984 ) );
  NAND2_X2 _f_permutation__U2317  ( .A1(SYNOPSYS_UNCONNECTED_702), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2985 ) );
  NAND2_X2 _f_permutation__U2316  ( .A1(_f_permutation__n2984 ), .A2(
        _f_permutation__n2985 ), .ZN(_f_permutation__n5001 ) );
  NAND2_X2 _f_permutation__U2315  ( .A1(_f_permutation__round_out[385]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2982 ) );
  NAND2_X2 _f_permutation__U2314  ( .A1(SYNOPSYS_UNCONNECTED_703), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2983 ) );
  NAND2_X2 _f_permutation__U2313  ( .A1(_f_permutation__n2982 ), .A2(
        _f_permutation__n2983 ), .ZN(_f_permutation__n5002 ) );
  NAND2_X2 _f_permutation__U2312  ( .A1(_f_permutation__round_out[384]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2980 ) );
  NAND2_X2 _f_permutation__U2311  ( .A1(SYNOPSYS_UNCONNECTED_704), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2981 ) );
  NAND2_X2 _f_permutation__U2310  ( .A1(_f_permutation__n2980 ), .A2(
        _f_permutation__n2981 ), .ZN(_f_permutation__n5003 ) );
  NAND2_X2 _f_permutation__U2309  ( .A1(_f_permutation__round_out[383]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2978 ) );
  NAND2_X2 _f_permutation__U2308  ( .A1(SYNOPSYS_UNCONNECTED_705), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2979 ) );
  NAND2_X2 _f_permutation__U2307  ( .A1(_f_permutation__n2978 ), .A2(
        _f_permutation__n2979 ), .ZN(_f_permutation__n5004 ) );
  NAND2_X2 _f_permutation__U2306  ( .A1(_f_permutation__round_out[382]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2976 ) );
  NAND2_X2 _f_permutation__U2305  ( .A1(SYNOPSYS_UNCONNECTED_706), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2977 ) );
  NAND2_X2 _f_permutation__U2304  ( .A1(_f_permutation__n2976 ), .A2(
        _f_permutation__n2977 ), .ZN(_f_permutation__n5005 ) );
  NAND2_X2 _f_permutation__U2303  ( .A1(_f_permutation__round_out[381]), .A2(
        _f_permutation__n7092 ), .ZN(_f_permutation__n2974 ) );
  NAND2_X2 _f_permutation__U2302  ( .A1(SYNOPSYS_UNCONNECTED_707), .A2(
        _f_permutation__n7273 ), .ZN(_f_permutation__n2975 ) );
  NAND2_X2 _f_permutation__U2301  ( .A1(_f_permutation__n2974 ), .A2(
        _f_permutation__n2975 ), .ZN(_f_permutation__n5006 ) );
  NAND2_X2 _f_permutation__U2300  ( .A1(_f_permutation__round_out[380]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2972 ) );
  NAND2_X2 _f_permutation__U2299  ( .A1(SYNOPSYS_UNCONNECTED_708), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2973 ) );
  NAND2_X2 _f_permutation__U2298  ( .A1(_f_permutation__n2972 ), .A2(
        _f_permutation__n2973 ), .ZN(_f_permutation__n5007 ) );
  NAND2_X2 _f_permutation__U2297  ( .A1(_f_permutation__round_out[379]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2970 ) );
  NAND2_X2 _f_permutation__U2296  ( .A1(SYNOPSYS_UNCONNECTED_709), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2971 ) );
  NAND2_X2 _f_permutation__U2295  ( .A1(_f_permutation__n2970 ), .A2(
        _f_permutation__n2971 ), .ZN(_f_permutation__n5008 ) );
  NAND2_X2 _f_permutation__U2294  ( .A1(_f_permutation__round_out[378]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2968 ) );
  NAND2_X2 _f_permutation__U2293  ( .A1(SYNOPSYS_UNCONNECTED_710), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2969 ) );
  NAND2_X2 _f_permutation__U2292  ( .A1(_f_permutation__n2968 ), .A2(
        _f_permutation__n2969 ), .ZN(_f_permutation__n5009 ) );
  NAND2_X2 _f_permutation__U2291  ( .A1(_f_permutation__round_out[377]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2966 ) );
  NAND2_X2 _f_permutation__U2290  ( .A1(SYNOPSYS_UNCONNECTED_711), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2967 ) );
  NAND2_X2 _f_permutation__U2289  ( .A1(_f_permutation__n2966 ), .A2(
        _f_permutation__n2967 ), .ZN(_f_permutation__n5010 ) );
  NAND2_X2 _f_permutation__U2288  ( .A1(_f_permutation__round_out[376]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2964 ) );
  NAND2_X2 _f_permutation__U2287  ( .A1(SYNOPSYS_UNCONNECTED_712), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2965 ) );
  NAND2_X2 _f_permutation__U2286  ( .A1(_f_permutation__n2964 ), .A2(
        _f_permutation__n2965 ), .ZN(_f_permutation__n5011 ) );
  NAND2_X2 _f_permutation__U2285  ( .A1(_f_permutation__round_out[375]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2962 ) );
  NAND2_X2 _f_permutation__U2284  ( .A1(SYNOPSYS_UNCONNECTED_713), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2963 ) );
  NAND2_X2 _f_permutation__U2283  ( .A1(_f_permutation__n2962 ), .A2(
        _f_permutation__n2963 ), .ZN(_f_permutation__n5012 ) );
  NAND2_X2 _f_permutation__U2282  ( .A1(_f_permutation__round_out[374]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2960 ) );
  NAND2_X2 _f_permutation__U2281  ( .A1(SYNOPSYS_UNCONNECTED_714), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2961 ) );
  NAND2_X2 _f_permutation__U2280  ( .A1(_f_permutation__n2960 ), .A2(
        _f_permutation__n2961 ), .ZN(_f_permutation__n5013 ) );
  NAND2_X2 _f_permutation__U2279  ( .A1(_f_permutation__round_out[373]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2958 ) );
  NAND2_X2 _f_permutation__U2278  ( .A1(SYNOPSYS_UNCONNECTED_715), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2959 ) );
  NAND2_X2 _f_permutation__U2277  ( .A1(_f_permutation__n2958 ), .A2(
        _f_permutation__n2959 ), .ZN(_f_permutation__n5014 ) );
  NAND2_X2 _f_permutation__U2276  ( .A1(_f_permutation__round_out[372]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2956 ) );
  NAND2_X2 _f_permutation__U2275  ( .A1(SYNOPSYS_UNCONNECTED_716), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2957 ) );
  NAND2_X2 _f_permutation__U2274  ( .A1(_f_permutation__n2956 ), .A2(
        _f_permutation__n2957 ), .ZN(_f_permutation__n5015 ) );
  NAND2_X2 _f_permutation__U2273  ( .A1(_f_permutation__round_out[371]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2954 ) );
  NAND2_X2 _f_permutation__U2272  ( .A1(SYNOPSYS_UNCONNECTED_717), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2955 ) );
  NAND2_X2 _f_permutation__U2271  ( .A1(_f_permutation__n2954 ), .A2(
        _f_permutation__n2955 ), .ZN(_f_permutation__n5016 ) );
  NAND2_X2 _f_permutation__U2270  ( .A1(_f_permutation__round_out[370]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2952 ) );
  NAND2_X2 _f_permutation__U2269  ( .A1(SYNOPSYS_UNCONNECTED_718), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2953 ) );
  NAND2_X2 _f_permutation__U2268  ( .A1(_f_permutation__n2952 ), .A2(
        _f_permutation__n2953 ), .ZN(_f_permutation__n5017 ) );
  NAND2_X2 _f_permutation__U2267  ( .A1(_f_permutation__round_out[369]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2950 ) );
  NAND2_X2 _f_permutation__U2266  ( .A1(SYNOPSYS_UNCONNECTED_719), .A2(
        _f_permutation__n7274 ), .ZN(_f_permutation__n2951 ) );
  NAND2_X2 _f_permutation__U2265  ( .A1(_f_permutation__n2950 ), .A2(
        _f_permutation__n2951 ), .ZN(_f_permutation__n5018 ) );
  NAND2_X2 _f_permutation__U2264  ( .A1(_f_permutation__round_out[368]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2948 ) );
  NAND2_X2 _f_permutation__U2263  ( .A1(SYNOPSYS_UNCONNECTED_720), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2949 ) );
  NAND2_X2 _f_permutation__U2262  ( .A1(_f_permutation__n2948 ), .A2(
        _f_permutation__n2949 ), .ZN(_f_permutation__n5019 ) );
  NAND2_X2 _f_permutation__U2261  ( .A1(_f_permutation__round_out[367]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2946 ) );
  NAND2_X2 _f_permutation__U2260  ( .A1(SYNOPSYS_UNCONNECTED_721), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2947 ) );
  NAND2_X2 _f_permutation__U2259  ( .A1(_f_permutation__n2946 ), .A2(
        _f_permutation__n2947 ), .ZN(_f_permutation__n5020 ) );
  NAND2_X2 _f_permutation__U2258  ( .A1(_f_permutation__round_out[366]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2944 ) );
  NAND2_X2 _f_permutation__U2257  ( .A1(SYNOPSYS_UNCONNECTED_722), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2945 ) );
  NAND2_X2 _f_permutation__U2256  ( .A1(_f_permutation__n2944 ), .A2(
        _f_permutation__n2945 ), .ZN(_f_permutation__n5021 ) );
  NAND2_X2 _f_permutation__U2255  ( .A1(_f_permutation__round_out[365]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2942 ) );
  NAND2_X2 _f_permutation__U2254  ( .A1(SYNOPSYS_UNCONNECTED_723), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2943 ) );
  NAND2_X2 _f_permutation__U2253  ( .A1(_f_permutation__n2942 ), .A2(
        _f_permutation__n2943 ), .ZN(_f_permutation__n5022 ) );
  NAND2_X2 _f_permutation__U2252  ( .A1(_f_permutation__round_out[364]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2940 ) );
  NAND2_X2 _f_permutation__U2251  ( .A1(SYNOPSYS_UNCONNECTED_724), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2941 ) );
  NAND2_X2 _f_permutation__U2250  ( .A1(_f_permutation__n2940 ), .A2(
        _f_permutation__n2941 ), .ZN(_f_permutation__n5023 ) );
  NAND2_X2 _f_permutation__U2249  ( .A1(_f_permutation__round_out[363]), .A2(
        _f_permutation__n7091 ), .ZN(_f_permutation__n2938 ) );
  NAND2_X2 _f_permutation__U2248  ( .A1(SYNOPSYS_UNCONNECTED_725), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2939 ) );
  NAND2_X2 _f_permutation__U2247  ( .A1(_f_permutation__n2938 ), .A2(
        _f_permutation__n2939 ), .ZN(_f_permutation__n5024 ) );
  NAND2_X2 _f_permutation__U2246  ( .A1(_f_permutation__round_out[362]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2936 ) );
  NAND2_X2 _f_permutation__U2245  ( .A1(SYNOPSYS_UNCONNECTED_726), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2937 ) );
  NAND2_X2 _f_permutation__U2244  ( .A1(_f_permutation__n2936 ), .A2(
        _f_permutation__n2937 ), .ZN(_f_permutation__n5025 ) );
  NAND2_X2 _f_permutation__U2243  ( .A1(_f_permutation__round_out[361]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2934 ) );
  NAND2_X2 _f_permutation__U2242  ( .A1(SYNOPSYS_UNCONNECTED_727), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2935 ) );
  NAND2_X2 _f_permutation__U2241  ( .A1(_f_permutation__n2934 ), .A2(
        _f_permutation__n2935 ), .ZN(_f_permutation__n5026 ) );
  NAND2_X2 _f_permutation__U2240  ( .A1(_f_permutation__round_out[360]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2932 ) );
  NAND2_X2 _f_permutation__U2239  ( .A1(SYNOPSYS_UNCONNECTED_728), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2933 ) );
  NAND2_X2 _f_permutation__U2238  ( .A1(_f_permutation__n2932 ), .A2(
        _f_permutation__n2933 ), .ZN(_f_permutation__n5027 ) );
  NAND2_X2 _f_permutation__U2237  ( .A1(_f_permutation__round_out[359]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2930 ) );
  NAND2_X2 _f_permutation__U2236  ( .A1(SYNOPSYS_UNCONNECTED_729), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2931 ) );
  NAND2_X2 _f_permutation__U2235  ( .A1(_f_permutation__n2930 ), .A2(
        _f_permutation__n2931 ), .ZN(_f_permutation__n5028 ) );
  NAND2_X2 _f_permutation__U2234  ( .A1(_f_permutation__round_out[358]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2928 ) );
  NAND2_X2 _f_permutation__U2233  ( .A1(SYNOPSYS_UNCONNECTED_730), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2929 ) );
  NAND2_X2 _f_permutation__U2232  ( .A1(_f_permutation__n2928 ), .A2(
        _f_permutation__n2929 ), .ZN(_f_permutation__n5029 ) );
  NAND2_X2 _f_permutation__U2231  ( .A1(_f_permutation__round_out[357]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2926 ) );
  NAND2_X2 _f_permutation__U2230  ( .A1(SYNOPSYS_UNCONNECTED_731), .A2(
        _f_permutation__n7275 ), .ZN(_f_permutation__n2927 ) );
  NAND2_X2 _f_permutation__U2229  ( .A1(_f_permutation__n2926 ), .A2(
        _f_permutation__n2927 ), .ZN(_f_permutation__n5030 ) );
  NAND2_X2 _f_permutation__U2228  ( .A1(_f_permutation__round_out[356]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2924 ) );
  NAND2_X2 _f_permutation__U2227  ( .A1(SYNOPSYS_UNCONNECTED_732), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2925 ) );
  NAND2_X2 _f_permutation__U2226  ( .A1(_f_permutation__n2924 ), .A2(
        _f_permutation__n2925 ), .ZN(_f_permutation__n5031 ) );
  NAND2_X2 _f_permutation__U2225  ( .A1(_f_permutation__round_out[355]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2922 ) );
  NAND2_X2 _f_permutation__U2224  ( .A1(SYNOPSYS_UNCONNECTED_733), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2923 ) );
  NAND2_X2 _f_permutation__U2223  ( .A1(_f_permutation__n2922 ), .A2(
        _f_permutation__n2923 ), .ZN(_f_permutation__n5032 ) );
  NAND2_X2 _f_permutation__U2222  ( .A1(_f_permutation__round_out[354]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2920 ) );
  NAND2_X2 _f_permutation__U2221  ( .A1(SYNOPSYS_UNCONNECTED_734), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2921 ) );
  NAND2_X2 _f_permutation__U2220  ( .A1(_f_permutation__n2920 ), .A2(
        _f_permutation__n2921 ), .ZN(_f_permutation__n5033 ) );
  NAND2_X2 _f_permutation__U2219  ( .A1(_f_permutation__round_out[353]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2918 ) );
  NAND2_X2 _f_permutation__U2218  ( .A1(SYNOPSYS_UNCONNECTED_735), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2919 ) );
  NAND2_X2 _f_permutation__U2217  ( .A1(_f_permutation__n2918 ), .A2(
        _f_permutation__n2919 ), .ZN(_f_permutation__n5034 ) );
  NAND2_X2 _f_permutation__U2216  ( .A1(_f_permutation__round_out[352]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2916 ) );
  NAND2_X2 _f_permutation__U2215  ( .A1(SYNOPSYS_UNCONNECTED_736), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2917 ) );
  NAND2_X2 _f_permutation__U2214  ( .A1(_f_permutation__n2916 ), .A2(
        _f_permutation__n2917 ), .ZN(_f_permutation__n5035 ) );
  NAND2_X2 _f_permutation__U2213  ( .A1(_f_permutation__round_out[351]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2914 ) );
  NAND2_X2 _f_permutation__U2212  ( .A1(SYNOPSYS_UNCONNECTED_737), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2915 ) );
  NAND2_X2 _f_permutation__U2211  ( .A1(_f_permutation__n2914 ), .A2(
        _f_permutation__n2915 ), .ZN(_f_permutation__n5036 ) );
  NAND2_X2 _f_permutation__U2210  ( .A1(_f_permutation__round_out[350]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2912 ) );
  NAND2_X2 _f_permutation__U2209  ( .A1(SYNOPSYS_UNCONNECTED_738), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2913 ) );
  NAND2_X2 _f_permutation__U2208  ( .A1(_f_permutation__n2912 ), .A2(
        _f_permutation__n2913 ), .ZN(_f_permutation__n5037 ) );
  NAND2_X2 _f_permutation__U2207  ( .A1(_f_permutation__round_out[349]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2910 ) );
  NAND2_X2 _f_permutation__U2206  ( .A1(SYNOPSYS_UNCONNECTED_739), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2911 ) );
  NAND2_X2 _f_permutation__U2205  ( .A1(_f_permutation__n2910 ), .A2(
        _f_permutation__n2911 ), .ZN(_f_permutation__n5038 ) );
  NAND2_X2 _f_permutation__U2204  ( .A1(_f_permutation__round_out[348]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2908 ) );
  NAND2_X2 _f_permutation__U2203  ( .A1(SYNOPSYS_UNCONNECTED_740), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2909 ) );
  NAND2_X2 _f_permutation__U2202  ( .A1(_f_permutation__n2908 ), .A2(
        _f_permutation__n2909 ), .ZN(_f_permutation__n5039 ) );
  NAND2_X2 _f_permutation__U2201  ( .A1(_f_permutation__round_out[347]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2906 ) );
  NAND2_X2 _f_permutation__U2200  ( .A1(SYNOPSYS_UNCONNECTED_741), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2907 ) );
  NAND2_X2 _f_permutation__U2199  ( .A1(_f_permutation__n2906 ), .A2(
        _f_permutation__n2907 ), .ZN(_f_permutation__n5040 ) );
  NAND2_X2 _f_permutation__U2198  ( .A1(_f_permutation__round_out[346]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2904 ) );
  NAND2_X2 _f_permutation__U2197  ( .A1(SYNOPSYS_UNCONNECTED_742), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2905 ) );
  NAND2_X2 _f_permutation__U2196  ( .A1(_f_permutation__n2904 ), .A2(
        _f_permutation__n2905 ), .ZN(_f_permutation__n5041 ) );
  NAND2_X2 _f_permutation__U2195  ( .A1(_f_permutation__round_out[345]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2902 ) );
  NAND2_X2 _f_permutation__U2194  ( .A1(SYNOPSYS_UNCONNECTED_743), .A2(
        _f_permutation__n7276 ), .ZN(_f_permutation__n2903 ) );
  NAND2_X2 _f_permutation__U2193  ( .A1(_f_permutation__n2902 ), .A2(
        _f_permutation__n2903 ), .ZN(_f_permutation__n5042 ) );
  NAND2_X2 _f_permutation__U2192  ( .A1(_f_permutation__round_out[344]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2900 ) );
  NAND2_X2 _f_permutation__U2191  ( .A1(SYNOPSYS_UNCONNECTED_744), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2901 ) );
  NAND2_X2 _f_permutation__U2190  ( .A1(_f_permutation__n2900 ), .A2(
        _f_permutation__n2901 ), .ZN(_f_permutation__n5043 ) );
  NAND2_X2 _f_permutation__U2189  ( .A1(_f_permutation__round_out[343]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2898 ) );
  NAND2_X2 _f_permutation__U2188  ( .A1(SYNOPSYS_UNCONNECTED_745), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2899 ) );
  NAND2_X2 _f_permutation__U2187  ( .A1(_f_permutation__n2898 ), .A2(
        _f_permutation__n2899 ), .ZN(_f_permutation__n5044 ) );
  NAND2_X2 _f_permutation__U2186  ( .A1(_f_permutation__round_out[342]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2896 ) );
  NAND2_X2 _f_permutation__U2185  ( .A1(SYNOPSYS_UNCONNECTED_746), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2897 ) );
  NAND2_X2 _f_permutation__U2184  ( .A1(_f_permutation__n2896 ), .A2(
        _f_permutation__n2897 ), .ZN(_f_permutation__n5045 ) );
  NAND2_X2 _f_permutation__U2183  ( .A1(_f_permutation__round_out[341]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2894 ) );
  NAND2_X2 _f_permutation__U2182  ( .A1(SYNOPSYS_UNCONNECTED_747), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2895 ) );
  NAND2_X2 _f_permutation__U2181  ( .A1(_f_permutation__n2894 ), .A2(
        _f_permutation__n2895 ), .ZN(_f_permutation__n5046 ) );
  NAND2_X2 _f_permutation__U2180  ( .A1(_f_permutation__round_out[340]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2892 ) );
  NAND2_X2 _f_permutation__U2179  ( .A1(SYNOPSYS_UNCONNECTED_748), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2893 ) );
  NAND2_X2 _f_permutation__U2178  ( .A1(_f_permutation__n2892 ), .A2(
        _f_permutation__n2893 ), .ZN(_f_permutation__n5047 ) );
  NAND2_X2 _f_permutation__U2177  ( .A1(_f_permutation__round_out[339]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2890 ) );
  NAND2_X2 _f_permutation__U2176  ( .A1(SYNOPSYS_UNCONNECTED_749), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2891 ) );
  NAND2_X2 _f_permutation__U2175  ( .A1(_f_permutation__n2890 ), .A2(
        _f_permutation__n2891 ), .ZN(_f_permutation__n5048 ) );
  NAND2_X2 _f_permutation__U2174  ( .A1(_f_permutation__round_out[338]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2888 ) );
  NAND2_X2 _f_permutation__U2173  ( .A1(SYNOPSYS_UNCONNECTED_750), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2889 ) );
  NAND2_X2 _f_permutation__U2172  ( .A1(_f_permutation__n2888 ), .A2(
        _f_permutation__n2889 ), .ZN(_f_permutation__n5049 ) );
  NAND2_X2 _f_permutation__U2171  ( .A1(_f_permutation__round_out[337]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2886 ) );
  NAND2_X2 _f_permutation__U2170  ( .A1(SYNOPSYS_UNCONNECTED_751), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2887 ) );
  NAND2_X2 _f_permutation__U2169  ( .A1(_f_permutation__n2886 ), .A2(
        _f_permutation__n2887 ), .ZN(_f_permutation__n5050 ) );
  NAND2_X2 _f_permutation__U2168  ( .A1(_f_permutation__round_out[336]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2884 ) );
  NAND2_X2 _f_permutation__U2167  ( .A1(SYNOPSYS_UNCONNECTED_752), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2885 ) );
  NAND2_X2 _f_permutation__U2166  ( .A1(_f_permutation__n2884 ), .A2(
        _f_permutation__n2885 ), .ZN(_f_permutation__n5051 ) );
  NAND2_X2 _f_permutation__U2165  ( .A1(_f_permutation__round_out[335]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2882 ) );
  NAND2_X2 _f_permutation__U2164  ( .A1(SYNOPSYS_UNCONNECTED_753), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2883 ) );
  NAND2_X2 _f_permutation__U2163  ( .A1(_f_permutation__n2882 ), .A2(
        _f_permutation__n2883 ), .ZN(_f_permutation__n5052 ) );
  NAND2_X2 _f_permutation__U2162  ( .A1(_f_permutation__round_out[334]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2880 ) );
  NAND2_X2 _f_permutation__U2161  ( .A1(SYNOPSYS_UNCONNECTED_754), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2881 ) );
  NAND2_X2 _f_permutation__U2160  ( .A1(_f_permutation__n2880 ), .A2(
        _f_permutation__n2881 ), .ZN(_f_permutation__n5053 ) );
  NAND2_X2 _f_permutation__U2159  ( .A1(_f_permutation__round_out[333]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2878 ) );
  NAND2_X2 _f_permutation__U2158  ( .A1(SYNOPSYS_UNCONNECTED_755), .A2(
        _f_permutation__n7277 ), .ZN(_f_permutation__n2879 ) );
  NAND2_X2 _f_permutation__U2157  ( .A1(_f_permutation__n2878 ), .A2(
        _f_permutation__n2879 ), .ZN(_f_permutation__n5054 ) );
  NAND2_X2 _f_permutation__U2156  ( .A1(_f_permutation__round_out[332]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2876 ) );
  NAND2_X2 _f_permutation__U2155  ( .A1(SYNOPSYS_UNCONNECTED_756), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2877 ) );
  NAND2_X2 _f_permutation__U2154  ( .A1(_f_permutation__n2876 ), .A2(
        _f_permutation__n2877 ), .ZN(_f_permutation__n5055 ) );
  NAND2_X2 _f_permutation__U2153  ( .A1(_f_permutation__round_out[331]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2874 ) );
  NAND2_X2 _f_permutation__U2152  ( .A1(SYNOPSYS_UNCONNECTED_757), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2875 ) );
  NAND2_X2 _f_permutation__U2151  ( .A1(_f_permutation__n2874 ), .A2(
        _f_permutation__n2875 ), .ZN(_f_permutation__n5056 ) );
  NAND2_X2 _f_permutation__U2150  ( .A1(_f_permutation__round_out[330]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2872 ) );
  NAND2_X2 _f_permutation__U2149  ( .A1(SYNOPSYS_UNCONNECTED_758), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2873 ) );
  NAND2_X2 _f_permutation__U2148  ( .A1(_f_permutation__n2872 ), .A2(
        _f_permutation__n2873 ), .ZN(_f_permutation__n5057 ) );
  NAND2_X2 _f_permutation__U2147  ( .A1(_f_permutation__round_out[329]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2870 ) );
  NAND2_X2 _f_permutation__U2146  ( .A1(SYNOPSYS_UNCONNECTED_759), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2871 ) );
  NAND2_X2 _f_permutation__U2145  ( .A1(_f_permutation__n2870 ), .A2(
        _f_permutation__n2871 ), .ZN(_f_permutation__n5058 ) );
  NAND2_X2 _f_permutation__U2144  ( .A1(_f_permutation__round_out[328]), .A2(
        _f_permutation__n7089 ), .ZN(_f_permutation__n2868 ) );
  NAND2_X2 _f_permutation__U2143  ( .A1(SYNOPSYS_UNCONNECTED_760), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2869 ) );
  NAND2_X2 _f_permutation__U2142  ( .A1(_f_permutation__n2868 ), .A2(
        _f_permutation__n2869 ), .ZN(_f_permutation__n5059 ) );
  NAND2_X2 _f_permutation__U2141  ( .A1(_f_permutation__round_out[327]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2866 ) );
  NAND2_X2 _f_permutation__U2140  ( .A1(SYNOPSYS_UNCONNECTED_761), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2867 ) );
  NAND2_X2 _f_permutation__U2139  ( .A1(_f_permutation__n2866 ), .A2(
        _f_permutation__n2867 ), .ZN(_f_permutation__n5060 ) );
  NAND2_X2 _f_permutation__U2138  ( .A1(_f_permutation__round_out[326]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2864 ) );
  NAND2_X2 _f_permutation__U2137  ( .A1(SYNOPSYS_UNCONNECTED_762), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2865 ) );
  NAND2_X2 _f_permutation__U2136  ( .A1(_f_permutation__n2864 ), .A2(
        _f_permutation__n2865 ), .ZN(_f_permutation__n5061 ) );
  NAND2_X2 _f_permutation__U2135  ( .A1(_f_permutation__round_out[325]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2862 ) );
  NAND2_X2 _f_permutation__U2134  ( .A1(SYNOPSYS_UNCONNECTED_763), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2863 ) );
  NAND2_X2 _f_permutation__U2133  ( .A1(_f_permutation__n2862 ), .A2(
        _f_permutation__n2863 ), .ZN(_f_permutation__n5062 ) );
  NAND2_X2 _f_permutation__U2132  ( .A1(_f_permutation__round_out[324]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2860 ) );
  NAND2_X2 _f_permutation__U2131  ( .A1(SYNOPSYS_UNCONNECTED_764), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2861 ) );
  NAND2_X2 _f_permutation__U2130  ( .A1(_f_permutation__n2860 ), .A2(
        _f_permutation__n2861 ), .ZN(_f_permutation__n5063 ) );
  NAND2_X2 _f_permutation__U2129  ( .A1(_f_permutation__round_out[323]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2858 ) );
  NAND2_X2 _f_permutation__U2128  ( .A1(SYNOPSYS_UNCONNECTED_765), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2859 ) );
  NAND2_X2 _f_permutation__U2127  ( .A1(_f_permutation__n2858 ), .A2(
        _f_permutation__n2859 ), .ZN(_f_permutation__n5064 ) );
  NAND2_X2 _f_permutation__U2126  ( .A1(_f_permutation__round_out[322]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2856 ) );
  NAND2_X2 _f_permutation__U2125  ( .A1(SYNOPSYS_UNCONNECTED_766), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2857 ) );
  NAND2_X2 _f_permutation__U2124  ( .A1(_f_permutation__n2856 ), .A2(
        _f_permutation__n2857 ), .ZN(_f_permutation__n5065 ) );
  NAND2_X2 _f_permutation__U2123  ( .A1(_f_permutation__round_out[321]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2854 ) );
  NAND2_X2 _f_permutation__U2122  ( .A1(SYNOPSYS_UNCONNECTED_767), .A2(
        _f_permutation__n7278 ), .ZN(_f_permutation__n2855 ) );
  NAND2_X2 _f_permutation__U2121  ( .A1(_f_permutation__n2854 ), .A2(
        _f_permutation__n2855 ), .ZN(_f_permutation__n5066 ) );
  NAND2_X2 _f_permutation__U2120  ( .A1(_f_permutation__round_out[320]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2852 ) );
  NAND2_X2 _f_permutation__U2119  ( .A1(SYNOPSYS_UNCONNECTED_768), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2853 ) );
  NAND2_X2 _f_permutation__U2118  ( .A1(_f_permutation__n2852 ), .A2(
        _f_permutation__n2853 ), .ZN(_f_permutation__n5067 ) );
  NAND2_X2 _f_permutation__U2117  ( .A1(_f_permutation__round_out[319]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2850 ) );
  NAND2_X2 _f_permutation__U2116  ( .A1(SYNOPSYS_UNCONNECTED_769), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2851 ) );
  NAND2_X2 _f_permutation__U2115  ( .A1(_f_permutation__n2850 ), .A2(
        _f_permutation__n2851 ), .ZN(_f_permutation__n5068 ) );
  NAND2_X2 _f_permutation__U2114  ( .A1(_f_permutation__round_out[318]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2848 ) );
  NAND2_X2 _f_permutation__U2113  ( .A1(SYNOPSYS_UNCONNECTED_770), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2849 ) );
  NAND2_X2 _f_permutation__U2112  ( .A1(_f_permutation__n2848 ), .A2(
        _f_permutation__n2849 ), .ZN(_f_permutation__n5069 ) );
  NAND2_X2 _f_permutation__U2111  ( .A1(_f_permutation__round_out[317]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2846 ) );
  NAND2_X2 _f_permutation__U2110  ( .A1(SYNOPSYS_UNCONNECTED_771), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2847 ) );
  NAND2_X2 _f_permutation__U2109  ( .A1(_f_permutation__n2846 ), .A2(
        _f_permutation__n2847 ), .ZN(_f_permutation__n5070 ) );
  NAND2_X2 _f_permutation__U2108  ( .A1(_f_permutation__round_out[316]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2844 ) );
  NAND2_X2 _f_permutation__U2107  ( .A1(SYNOPSYS_UNCONNECTED_772), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2845 ) );
  NAND2_X2 _f_permutation__U2106  ( .A1(_f_permutation__n2844 ), .A2(
        _f_permutation__n2845 ), .ZN(_f_permutation__n5071 ) );
  NAND2_X2 _f_permutation__U2105  ( .A1(_f_permutation__round_out[315]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2842 ) );
  NAND2_X2 _f_permutation__U2104  ( .A1(SYNOPSYS_UNCONNECTED_773), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2843 ) );
  NAND2_X2 _f_permutation__U2103  ( .A1(_f_permutation__n2842 ), .A2(
        _f_permutation__n2843 ), .ZN(_f_permutation__n5072 ) );
  NAND2_X2 _f_permutation__U2102  ( .A1(_f_permutation__round_out[314]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2840 ) );
  NAND2_X2 _f_permutation__U2101  ( .A1(SYNOPSYS_UNCONNECTED_774), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2841 ) );
  NAND2_X2 _f_permutation__U2100  ( .A1(_f_permutation__n2840 ), .A2(
        _f_permutation__n2841 ), .ZN(_f_permutation__n5073 ) );
  NAND2_X2 _f_permutation__U2099  ( .A1(_f_permutation__round_out[313]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2838 ) );
  NAND2_X2 _f_permutation__U2098  ( .A1(SYNOPSYS_UNCONNECTED_775), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2839 ) );
  NAND2_X2 _f_permutation__U2097  ( .A1(_f_permutation__n2838 ), .A2(
        _f_permutation__n2839 ), .ZN(_f_permutation__n5074 ) );
  NAND2_X2 _f_permutation__U2096  ( .A1(_f_permutation__round_out[312]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2836 ) );
  NAND2_X2 _f_permutation__U2095  ( .A1(SYNOPSYS_UNCONNECTED_776), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2837 ) );
  NAND2_X2 _f_permutation__U2094  ( .A1(_f_permutation__n2836 ), .A2(
        _f_permutation__n2837 ), .ZN(_f_permutation__n5075 ) );
  NAND2_X2 _f_permutation__U2093  ( .A1(_f_permutation__round_out[311]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2834 ) );
  NAND2_X2 _f_permutation__U2092  ( .A1(SYNOPSYS_UNCONNECTED_777), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2835 ) );
  NAND2_X2 _f_permutation__U2091  ( .A1(_f_permutation__n2834 ), .A2(
        _f_permutation__n2835 ), .ZN(_f_permutation__n5076 ) );
  NAND2_X2 _f_permutation__U2090  ( .A1(_f_permutation__round_out[310]), .A2(
        _f_permutation__n7088 ), .ZN(_f_permutation__n2832 ) );
  NAND2_X2 _f_permutation__U2089  ( .A1(SYNOPSYS_UNCONNECTED_778), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2833 ) );
  NAND2_X2 _f_permutation__U2088  ( .A1(_f_permutation__n2832 ), .A2(
        _f_permutation__n2833 ), .ZN(_f_permutation__n5077 ) );
  NAND2_X2 _f_permutation__U2087  ( .A1(_f_permutation__round_out[309]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n2830 ) );
  NAND2_X2 _f_permutation__U2086  ( .A1(SYNOPSYS_UNCONNECTED_779), .A2(
        _f_permutation__n7279 ), .ZN(_f_permutation__n2831 ) );
  NAND2_X2 _f_permutation__U2085  ( .A1(_f_permutation__n2830 ), .A2(
        _f_permutation__n2831 ), .ZN(_f_permutation__n5078 ) );
  NAND2_X2 _f_permutation__U2084  ( .A1(_f_permutation__round_out[308]), .A2(
        _f_permutation__n7168 ), .ZN(_f_permutation__n2828 ) );
  NAND2_X2 _f_permutation__U2083  ( .A1(SYNOPSYS_UNCONNECTED_780), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2829 ) );
  NAND2_X2 _f_permutation__U2082  ( .A1(_f_permutation__n2828 ), .A2(
        _f_permutation__n2829 ), .ZN(_f_permutation__n5079 ) );
  NAND2_X2 _f_permutation__U2081  ( .A1(_f_permutation__round_out[307]), .A2(
        _f_permutation__n7140 ), .ZN(_f_permutation__n2826 ) );
  NAND2_X2 _f_permutation__U2080  ( .A1(SYNOPSYS_UNCONNECTED_781), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2827 ) );
  NAND2_X2 _f_permutation__U2079  ( .A1(_f_permutation__n2826 ), .A2(
        _f_permutation__n2827 ), .ZN(_f_permutation__n5080 ) );
  NAND2_X2 _f_permutation__U2078  ( .A1(_f_permutation__round_out[306]), .A2(
        _f_permutation__n7149 ), .ZN(_f_permutation__n2824 ) );
  NAND2_X2 _f_permutation__U2077  ( .A1(SYNOPSYS_UNCONNECTED_782), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2825 ) );
  NAND2_X2 _f_permutation__U2076  ( .A1(_f_permutation__n2824 ), .A2(
        _f_permutation__n2825 ), .ZN(_f_permutation__n5081 ) );
  NAND2_X2 _f_permutation__U2075  ( .A1(_f_permutation__round_out[305]), .A2(
        _f_permutation__n7148 ), .ZN(_f_permutation__n2822 ) );
  NAND2_X2 _f_permutation__U2074  ( .A1(SYNOPSYS_UNCONNECTED_783), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2823 ) );
  NAND2_X2 _f_permutation__U2073  ( .A1(_f_permutation__n2822 ), .A2(
        _f_permutation__n2823 ), .ZN(_f_permutation__n5082 ) );
  NAND2_X2 _f_permutation__U2072  ( .A1(_f_permutation__round_out[304]), .A2(
        _f_permutation__n7147 ), .ZN(_f_permutation__n2820 ) );
  NAND2_X2 _f_permutation__U2071  ( .A1(SYNOPSYS_UNCONNECTED_784), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2821 ) );
  NAND2_X2 _f_permutation__U2070  ( .A1(_f_permutation__n2820 ), .A2(
        _f_permutation__n2821 ), .ZN(_f_permutation__n5083 ) );
  NAND2_X2 _f_permutation__U2069  ( .A1(_f_permutation__round_out[303]), .A2(
        _f_permutation__n7152 ), .ZN(_f_permutation__n2818 ) );
  NAND2_X2 _f_permutation__U2068  ( .A1(SYNOPSYS_UNCONNECTED_785), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2819 ) );
  NAND2_X2 _f_permutation__U2067  ( .A1(_f_permutation__n2818 ), .A2(
        _f_permutation__n2819 ), .ZN(_f_permutation__n5084 ) );
  NAND2_X2 _f_permutation__U2066  ( .A1(_f_permutation__round_out[302]), .A2(
        _f_permutation__n7151 ), .ZN(_f_permutation__n2816 ) );
  NAND2_X2 _f_permutation__U2065  ( .A1(SYNOPSYS_UNCONNECTED_786), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2817 ) );
  NAND2_X2 _f_permutation__U2064  ( .A1(_f_permutation__n2816 ), .A2(
        _f_permutation__n2817 ), .ZN(_f_permutation__n5085 ) );
  NAND2_X2 _f_permutation__U2063  ( .A1(_f_permutation__round_out[301]), .A2(
        _f_permutation__n7150 ), .ZN(_f_permutation__n2814 ) );
  NAND2_X2 _f_permutation__U2062  ( .A1(SYNOPSYS_UNCONNECTED_787), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2815 ) );
  NAND2_X2 _f_permutation__U2061  ( .A1(_f_permutation__n2814 ), .A2(
        _f_permutation__n2815 ), .ZN(_f_permutation__n5086 ) );
  NAND2_X2 _f_permutation__U2060  ( .A1(_f_permutation__round_out[300]), .A2(
        _f_permutation__n7090 ), .ZN(_f_permutation__n2812 ) );
  NAND2_X2 _f_permutation__U2059  ( .A1(SYNOPSYS_UNCONNECTED_788), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2813 ) );
  NAND2_X2 _f_permutation__U2058  ( .A1(_f_permutation__n2812 ), .A2(
        _f_permutation__n2813 ), .ZN(_f_permutation__n5087 ) );
  NAND2_X2 _f_permutation__U2057  ( .A1(_f_permutation__round_out[299]), .A2(
        _f_permutation__n7164 ), .ZN(_f_permutation__n2810 ) );
  NAND2_X2 _f_permutation__U2056  ( .A1(SYNOPSYS_UNCONNECTED_789), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2811 ) );
  NAND2_X2 _f_permutation__U2055  ( .A1(_f_permutation__n2810 ), .A2(
        _f_permutation__n2811 ), .ZN(_f_permutation__n5088 ) );
  NAND2_X2 _f_permutation__U2054  ( .A1(_f_permutation__round_out[298]), .A2(
        _f_permutation__n7156 ), .ZN(_f_permutation__n2808 ) );
  NAND2_X2 _f_permutation__U2053  ( .A1(SYNOPSYS_UNCONNECTED_790), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2809 ) );
  NAND2_X2 _f_permutation__U2052  ( .A1(_f_permutation__n2808 ), .A2(
        _f_permutation__n2809 ), .ZN(_f_permutation__n5089 ) );
  NAND2_X2 _f_permutation__U2051  ( .A1(_f_permutation__round_out[297]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n2806 ) );
  NAND2_X2 _f_permutation__U2050  ( .A1(SYNOPSYS_UNCONNECTED_791), .A2(
        _f_permutation__n7280 ), .ZN(_f_permutation__n2807 ) );
  NAND2_X2 _f_permutation__U2049  ( .A1(_f_permutation__n2806 ), .A2(
        _f_permutation__n2807 ), .ZN(_f_permutation__n5090 ) );
  NAND2_X2 _f_permutation__U2048  ( .A1(_f_permutation__round_out[296]), .A2(
        _f_permutation__n7154 ), .ZN(_f_permutation__n2804 ) );
  NAND2_X2 _f_permutation__U2047  ( .A1(SYNOPSYS_UNCONNECTED_792), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2805 ) );
  NAND2_X2 _f_permutation__U2046  ( .A1(_f_permutation__n2804 ), .A2(
        _f_permutation__n2805 ), .ZN(_f_permutation__n5091 ) );
  NAND2_X2 _f_permutation__U2045  ( .A1(_f_permutation__round_out[295]), .A2(
        _f_permutation__n7161 ), .ZN(_f_permutation__n2802 ) );
  NAND2_X2 _f_permutation__U2044  ( .A1(SYNOPSYS_UNCONNECTED_793), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2803 ) );
  NAND2_X2 _f_permutation__U2043  ( .A1(_f_permutation__n2802 ), .A2(
        _f_permutation__n2803 ), .ZN(_f_permutation__n5092 ) );
  NAND2_X2 _f_permutation__U2042  ( .A1(_f_permutation__round_out[294]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n2800 ) );
  NAND2_X2 _f_permutation__U2041  ( .A1(SYNOPSYS_UNCONNECTED_794), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2801 ) );
  NAND2_X2 _f_permutation__U2040  ( .A1(_f_permutation__n2800 ), .A2(
        _f_permutation__n2801 ), .ZN(_f_permutation__n5093 ) );
  NAND2_X2 _f_permutation__U2039  ( .A1(_f_permutation__round_out[293]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n2798 ) );
  NAND2_X2 _f_permutation__U2038  ( .A1(SYNOPSYS_UNCONNECTED_795), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2799 ) );
  NAND2_X2 _f_permutation__U2037  ( .A1(_f_permutation__n2798 ), .A2(
        _f_permutation__n2799 ), .ZN(_f_permutation__n5094 ) );
  NAND2_X2 _f_permutation__U2036  ( .A1(_f_permutation__round_out[292]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n2796 ) );
  NAND2_X2 _f_permutation__U2035  ( .A1(SYNOPSYS_UNCONNECTED_796), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2797 ) );
  NAND2_X2 _f_permutation__U2034  ( .A1(_f_permutation__n2796 ), .A2(
        _f_permutation__n2797 ), .ZN(_f_permutation__n5095 ) );
  NAND2_X2 _f_permutation__U2033  ( .A1(_f_permutation__round_out[291]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n2794 ) );
  NAND2_X2 _f_permutation__U2032  ( .A1(SYNOPSYS_UNCONNECTED_797), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2795 ) );
  NAND2_X2 _f_permutation__U2031  ( .A1(_f_permutation__n2794 ), .A2(
        _f_permutation__n2795 ), .ZN(_f_permutation__n5096 ) );
  NAND2_X2 _f_permutation__U2030  ( .A1(_f_permutation__round_out[290]), .A2(
        _f_permutation__n7153 ), .ZN(_f_permutation__n2792 ) );
  NAND2_X2 _f_permutation__U2029  ( .A1(SYNOPSYS_UNCONNECTED_798), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2793 ) );
  NAND2_X2 _f_permutation__U2028  ( .A1(_f_permutation__n2792 ), .A2(
        _f_permutation__n2793 ), .ZN(_f_permutation__n5097 ) );
  NAND2_X2 _f_permutation__U2027  ( .A1(_f_permutation__round_out[289]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2790 ) );
  NAND2_X2 _f_permutation__U2026  ( .A1(SYNOPSYS_UNCONNECTED_799), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2791 ) );
  NAND2_X2 _f_permutation__U2025  ( .A1(_f_permutation__n2790 ), .A2(
        _f_permutation__n2791 ), .ZN(_f_permutation__n5098 ) );
  NAND2_X2 _f_permutation__U2024  ( .A1(_f_permutation__round_out[288]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2788 ) );
  NAND2_X2 _f_permutation__U2023  ( .A1(SYNOPSYS_UNCONNECTED_800), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2789 ) );
  NAND2_X2 _f_permutation__U2022  ( .A1(_f_permutation__n2788 ), .A2(
        _f_permutation__n2789 ), .ZN(_f_permutation__n5099 ) );
  NAND2_X2 _f_permutation__U2021  ( .A1(_f_permutation__round_out[287]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2786 ) );
  NAND2_X2 _f_permutation__U2020  ( .A1(SYNOPSYS_UNCONNECTED_801), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2787 ) );
  NAND2_X2 _f_permutation__U2019  ( .A1(_f_permutation__n2786 ), .A2(
        _f_permutation__n2787 ), .ZN(_f_permutation__n5100 ) );
  NAND2_X2 _f_permutation__U2018  ( .A1(_f_permutation__round_out[286]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2784 ) );
  NAND2_X2 _f_permutation__U2017  ( .A1(SYNOPSYS_UNCONNECTED_802), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2785 ) );
  NAND2_X2 _f_permutation__U2016  ( .A1(_f_permutation__n2784 ), .A2(
        _f_permutation__n2785 ), .ZN(_f_permutation__n5101 ) );
  NAND2_X2 _f_permutation__U2015  ( .A1(_f_permutation__round_out[285]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2782 ) );
  NAND2_X2 _f_permutation__U2014  ( .A1(SYNOPSYS_UNCONNECTED_803), .A2(
        _f_permutation__n7281 ), .ZN(_f_permutation__n2783 ) );
  NAND2_X2 _f_permutation__U2013  ( .A1(_f_permutation__n2782 ), .A2(
        _f_permutation__n2783 ), .ZN(_f_permutation__n5102 ) );
  NAND2_X2 _f_permutation__U2012  ( .A1(_f_permutation__round_out[284]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2780 ) );
  NAND2_X2 _f_permutation__U2011  ( .A1(SYNOPSYS_UNCONNECTED_804), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2781 ) );
  NAND2_X2 _f_permutation__U2010  ( .A1(_f_permutation__n2780 ), .A2(
        _f_permutation__n2781 ), .ZN(_f_permutation__n5103 ) );
  NAND2_X2 _f_permutation__U2009  ( .A1(_f_permutation__round_out[283]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2778 ) );
  NAND2_X2 _f_permutation__U2008  ( .A1(SYNOPSYS_UNCONNECTED_805), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2779 ) );
  NAND2_X2 _f_permutation__U2007  ( .A1(_f_permutation__n2778 ), .A2(
        _f_permutation__n2779 ), .ZN(_f_permutation__n5104 ) );
  NAND2_X2 _f_permutation__U2006  ( .A1(_f_permutation__round_out[282]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2776 ) );
  NAND2_X2 _f_permutation__U2005  ( .A1(SYNOPSYS_UNCONNECTED_806), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2777 ) );
  NAND2_X2 _f_permutation__U2004  ( .A1(_f_permutation__n2776 ), .A2(
        _f_permutation__n2777 ), .ZN(_f_permutation__n5105 ) );
  NAND2_X2 _f_permutation__U2003  ( .A1(_f_permutation__round_out[281]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2774 ) );
  NAND2_X2 _f_permutation__U2002  ( .A1(SYNOPSYS_UNCONNECTED_807), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2775 ) );
  NAND2_X2 _f_permutation__U2001  ( .A1(_f_permutation__n2774 ), .A2(
        _f_permutation__n2775 ), .ZN(_f_permutation__n5106 ) );
  NAND2_X2 _f_permutation__U2000  ( .A1(_f_permutation__round_out[280]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2772 ) );
  NAND2_X2 _f_permutation__U1999  ( .A1(SYNOPSYS_UNCONNECTED_808), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2773 ) );
  NAND2_X2 _f_permutation__U1998  ( .A1(_f_permutation__n2772 ), .A2(
        _f_permutation__n2773 ), .ZN(_f_permutation__n5107 ) );
  NAND2_X2 _f_permutation__U1997  ( .A1(_f_permutation__round_out[279]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2770 ) );
  NAND2_X2 _f_permutation__U1996  ( .A1(SYNOPSYS_UNCONNECTED_809), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2771 ) );
  NAND2_X2 _f_permutation__U1995  ( .A1(_f_permutation__n2770 ), .A2(
        _f_permutation__n2771 ), .ZN(_f_permutation__n5108 ) );
  NAND2_X2 _f_permutation__U1994  ( .A1(_f_permutation__round_out[278]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2768 ) );
  NAND2_X2 _f_permutation__U1993  ( .A1(SYNOPSYS_UNCONNECTED_810), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2769 ) );
  NAND2_X2 _f_permutation__U1992  ( .A1(_f_permutation__n2768 ), .A2(
        _f_permutation__n2769 ), .ZN(_f_permutation__n5109 ) );
  NAND2_X2 _f_permutation__U1991  ( .A1(_f_permutation__round_out[277]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2766 ) );
  NAND2_X2 _f_permutation__U1990  ( .A1(SYNOPSYS_UNCONNECTED_811), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2767 ) );
  NAND2_X2 _f_permutation__U1989  ( .A1(_f_permutation__n2766 ), .A2(
        _f_permutation__n2767 ), .ZN(_f_permutation__n5110 ) );
  NAND2_X2 _f_permutation__U1988  ( .A1(_f_permutation__round_out[276]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2764 ) );
  NAND2_X2 _f_permutation__U1987  ( .A1(SYNOPSYS_UNCONNECTED_812), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2765 ) );
  NAND2_X2 _f_permutation__U1986  ( .A1(_f_permutation__n2764 ), .A2(
        _f_permutation__n2765 ), .ZN(_f_permutation__n5111 ) );
  NAND2_X2 _f_permutation__U1985  ( .A1(_f_permutation__round_out[275]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2762 ) );
  NAND2_X2 _f_permutation__U1984  ( .A1(SYNOPSYS_UNCONNECTED_813), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2763 ) );
  NAND2_X2 _f_permutation__U1983  ( .A1(_f_permutation__n2762 ), .A2(
        _f_permutation__n2763 ), .ZN(_f_permutation__n5112 ) );
  NAND2_X2 _f_permutation__U1982  ( .A1(_f_permutation__round_out[274]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2760 ) );
  NAND2_X2 _f_permutation__U1981  ( .A1(SYNOPSYS_UNCONNECTED_814), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2761 ) );
  NAND2_X2 _f_permutation__U1980  ( .A1(_f_permutation__n2760 ), .A2(
        _f_permutation__n2761 ), .ZN(_f_permutation__n5113 ) );
  NAND2_X2 _f_permutation__U1979  ( .A1(_f_permutation__round_out[273]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2758 ) );
  NAND2_X2 _f_permutation__U1978  ( .A1(SYNOPSYS_UNCONNECTED_815), .A2(
        _f_permutation__n7282 ), .ZN(_f_permutation__n2759 ) );
  NAND2_X2 _f_permutation__U1977  ( .A1(_f_permutation__n2758 ), .A2(
        _f_permutation__n2759 ), .ZN(_f_permutation__n5114 ) );
  NAND2_X2 _f_permutation__U1976  ( .A1(_f_permutation__round_out[272]), .A2(
        _f_permutation__n7094 ), .ZN(_f_permutation__n2756 ) );
  NAND2_X2 _f_permutation__U1975  ( .A1(SYNOPSYS_UNCONNECTED_816), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2757 ) );
  NAND2_X2 _f_permutation__U1974  ( .A1(_f_permutation__n2756 ), .A2(
        _f_permutation__n2757 ), .ZN(_f_permutation__n5115 ) );
  NAND2_X2 _f_permutation__U1973  ( .A1(_f_permutation__round_out[271]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2754 ) );
  NAND2_X2 _f_permutation__U1972  ( .A1(SYNOPSYS_UNCONNECTED_817), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2755 ) );
  NAND2_X2 _f_permutation__U1971  ( .A1(_f_permutation__n2754 ), .A2(
        _f_permutation__n2755 ), .ZN(_f_permutation__n5116 ) );
  NAND2_X2 _f_permutation__U1970  ( .A1(_f_permutation__round_out[270]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2752 ) );
  NAND2_X2 _f_permutation__U1969  ( .A1(SYNOPSYS_UNCONNECTED_818), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2753 ) );
  NAND2_X2 _f_permutation__U1968  ( .A1(_f_permutation__n2752 ), .A2(
        _f_permutation__n2753 ), .ZN(_f_permutation__n5117 ) );
  NAND2_X2 _f_permutation__U1967  ( .A1(_f_permutation__round_out[269]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2750 ) );
  NAND2_X2 _f_permutation__U1966  ( .A1(SYNOPSYS_UNCONNECTED_819), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2751 ) );
  NAND2_X2 _f_permutation__U1965  ( .A1(_f_permutation__n2750 ), .A2(
        _f_permutation__n2751 ), .ZN(_f_permutation__n5118 ) );
  NAND2_X2 _f_permutation__U1964  ( .A1(_f_permutation__round_out[268]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2748 ) );
  NAND2_X2 _f_permutation__U1963  ( .A1(SYNOPSYS_UNCONNECTED_820), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2749 ) );
  NAND2_X2 _f_permutation__U1962  ( .A1(_f_permutation__n2748 ), .A2(
        _f_permutation__n2749 ), .ZN(_f_permutation__n5119 ) );
  NAND2_X2 _f_permutation__U1961  ( .A1(_f_permutation__round_out[267]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2746 ) );
  NAND2_X2 _f_permutation__U1960  ( .A1(SYNOPSYS_UNCONNECTED_821), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2747 ) );
  NAND2_X2 _f_permutation__U1959  ( .A1(_f_permutation__n2746 ), .A2(
        _f_permutation__n2747 ), .ZN(_f_permutation__n5120 ) );
  NAND2_X2 _f_permutation__U1958  ( .A1(_f_permutation__round_out[266]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2744 ) );
  NAND2_X2 _f_permutation__U1957  ( .A1(SYNOPSYS_UNCONNECTED_822), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2745 ) );
  NAND2_X2 _f_permutation__U1956  ( .A1(_f_permutation__n2744 ), .A2(
        _f_permutation__n2745 ), .ZN(_f_permutation__n5121 ) );
  NAND2_X2 _f_permutation__U1955  ( .A1(_f_permutation__round_out[265]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2742 ) );
  NAND2_X2 _f_permutation__U1954  ( .A1(SYNOPSYS_UNCONNECTED_823), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2743 ) );
  NAND2_X2 _f_permutation__U1953  ( .A1(_f_permutation__n2742 ), .A2(
        _f_permutation__n2743 ), .ZN(_f_permutation__n5122 ) );
  NAND2_X2 _f_permutation__U1952  ( .A1(_f_permutation__round_out[264]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2740 ) );
  NAND2_X2 _f_permutation__U1951  ( .A1(SYNOPSYS_UNCONNECTED_824), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2741 ) );
  NAND2_X2 _f_permutation__U1950  ( .A1(_f_permutation__n2740 ), .A2(
        _f_permutation__n2741 ), .ZN(_f_permutation__n5123 ) );
  NAND2_X2 _f_permutation__U1949  ( .A1(_f_permutation__round_out[263]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2738 ) );
  NAND2_X2 _f_permutation__U1948  ( .A1(SYNOPSYS_UNCONNECTED_825), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2739 ) );
  NAND2_X2 _f_permutation__U1947  ( .A1(_f_permutation__n2738 ), .A2(
        _f_permutation__n2739 ), .ZN(_f_permutation__n5124 ) );
  NAND2_X2 _f_permutation__U1946  ( .A1(_f_permutation__round_out[262]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2736 ) );
  NAND2_X2 _f_permutation__U1945  ( .A1(SYNOPSYS_UNCONNECTED_826), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2737 ) );
  NAND2_X2 _f_permutation__U1944  ( .A1(_f_permutation__n2736 ), .A2(
        _f_permutation__n2737 ), .ZN(_f_permutation__n5125 ) );
  NAND2_X2 _f_permutation__U1943  ( .A1(_f_permutation__round_out[261]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2734 ) );
  NAND2_X2 _f_permutation__U1942  ( .A1(SYNOPSYS_UNCONNECTED_827), .A2(
        _f_permutation__n7283 ), .ZN(_f_permutation__n2735 ) );
  NAND2_X2 _f_permutation__U1941  ( .A1(_f_permutation__n2734 ), .A2(
        _f_permutation__n2735 ), .ZN(_f_permutation__n5126 ) );
  NAND2_X2 _f_permutation__U1940  ( .A1(_f_permutation__round_out[260]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2732 ) );
  NAND2_X2 _f_permutation__U1939  ( .A1(SYNOPSYS_UNCONNECTED_828), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2733 ) );
  NAND2_X2 _f_permutation__U1938  ( .A1(_f_permutation__n2732 ), .A2(
        _f_permutation__n2733 ), .ZN(_f_permutation__n5127 ) );
  NAND2_X2 _f_permutation__U1937  ( .A1(_f_permutation__round_out[259]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2730 ) );
  NAND2_X2 _f_permutation__U1936  ( .A1(SYNOPSYS_UNCONNECTED_829), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2731 ) );
  NAND2_X2 _f_permutation__U1935  ( .A1(_f_permutation__n2730 ), .A2(
        _f_permutation__n2731 ), .ZN(_f_permutation__n5128 ) );
  NAND2_X2 _f_permutation__U1934  ( .A1(_f_permutation__round_out[258]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2728 ) );
  NAND2_X2 _f_permutation__U1933  ( .A1(SYNOPSYS_UNCONNECTED_830), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2729 ) );
  NAND2_X2 _f_permutation__U1932  ( .A1(_f_permutation__n2728 ), .A2(
        _f_permutation__n2729 ), .ZN(_f_permutation__n5129 ) );
  NAND2_X2 _f_permutation__U1931  ( .A1(_f_permutation__round_out[257]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2726 ) );
  NAND2_X2 _f_permutation__U1930  ( .A1(SYNOPSYS_UNCONNECTED_831), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2727 ) );
  NAND2_X2 _f_permutation__U1929  ( .A1(_f_permutation__n2726 ), .A2(
        _f_permutation__n2727 ), .ZN(_f_permutation__n5130 ) );
  NAND2_X2 _f_permutation__U1928  ( .A1(_f_permutation__round_out[256]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2724 ) );
  NAND2_X2 _f_permutation__U1927  ( .A1(SYNOPSYS_UNCONNECTED_832), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2725 ) );
  NAND2_X2 _f_permutation__U1926  ( .A1(_f_permutation__n2724 ), .A2(
        _f_permutation__n2725 ), .ZN(_f_permutation__n5131 ) );
  NAND2_X2 _f_permutation__U1925  ( .A1(_f_permutation__round_out[255]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2722 ) );
  NAND2_X2 _f_permutation__U1924  ( .A1(SYNOPSYS_UNCONNECTED_833), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2723 ) );
  NAND2_X2 _f_permutation__U1923  ( .A1(_f_permutation__n2722 ), .A2(
        _f_permutation__n2723 ), .ZN(_f_permutation__n5132 ) );
  NAND2_X2 _f_permutation__U1922  ( .A1(_f_permutation__round_out[254]), .A2(
        _f_permutation__n7093 ), .ZN(_f_permutation__n2720 ) );
  NAND2_X2 _f_permutation__U1921  ( .A1(SYNOPSYS_UNCONNECTED_834), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2721 ) );
  NAND2_X2 _f_permutation__U1920  ( .A1(_f_permutation__n2720 ), .A2(
        _f_permutation__n2721 ), .ZN(_f_permutation__n5133 ) );
  NAND2_X2 _f_permutation__U1919  ( .A1(_f_permutation__round_out[253]), .A2(
        _f_permutation__n7154 ), .ZN(_f_permutation__n2718 ) );
  NAND2_X2 _f_permutation__U1918  ( .A1(SYNOPSYS_UNCONNECTED_835), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2719 ) );
  NAND2_X2 _f_permutation__U1917  ( .A1(_f_permutation__n2718 ), .A2(
        _f_permutation__n2719 ), .ZN(_f_permutation__n5134 ) );
  NAND2_X2 _f_permutation__U1916  ( .A1(_f_permutation__round_out[252]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n2716 ) );
  NAND2_X2 _f_permutation__U1915  ( .A1(SYNOPSYS_UNCONNECTED_836), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2717 ) );
  NAND2_X2 _f_permutation__U1914  ( .A1(_f_permutation__n2716 ), .A2(
        _f_permutation__n2717 ), .ZN(_f_permutation__n5135 ) );
  NAND2_X2 _f_permutation__U1913  ( .A1(_f_permutation__round_out[251]), .A2(
        _f_permutation__n7149 ), .ZN(_f_permutation__n2714 ) );
  NAND2_X2 _f_permutation__U1912  ( .A1(SYNOPSYS_UNCONNECTED_837), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2715 ) );
  NAND2_X2 _f_permutation__U1911  ( .A1(_f_permutation__n2714 ), .A2(
        _f_permutation__n2715 ), .ZN(_f_permutation__n5136 ) );
  NAND2_X2 _f_permutation__U1910  ( .A1(_f_permutation__round_out[250]), .A2(
        _f_permutation__n7147 ), .ZN(_f_permutation__n2712 ) );
  NAND2_X2 _f_permutation__U1909  ( .A1(SYNOPSYS_UNCONNECTED_838), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2713 ) );
  NAND2_X2 _f_permutation__U1908  ( .A1(_f_permutation__n2712 ), .A2(
        _f_permutation__n2713 ), .ZN(_f_permutation__n5137 ) );
  NAND2_X2 _f_permutation__U1907  ( .A1(_f_permutation__round_out[249]), .A2(
        _f_permutation__n7152 ), .ZN(_f_permutation__n2710 ) );
  NAND2_X2 _f_permutation__U1906  ( .A1(SYNOPSYS_UNCONNECTED_839), .A2(
        _f_permutation__n7284 ), .ZN(_f_permutation__n2711 ) );
  NAND2_X2 _f_permutation__U1905  ( .A1(_f_permutation__n2710 ), .A2(
        _f_permutation__n2711 ), .ZN(_f_permutation__n5138 ) );
  NAND2_X2 _f_permutation__U1904  ( .A1(_f_permutation__round_out[248]), .A2(
        _f_permutation__n7151 ), .ZN(_f_permutation__n2708 ) );
  NAND2_X2 _f_permutation__U1903  ( .A1(SYNOPSYS_UNCONNECTED_840), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2709 ) );
  NAND2_X2 _f_permutation__U1902  ( .A1(_f_permutation__n2708 ), .A2(
        _f_permutation__n2709 ), .ZN(_f_permutation__n5139 ) );
  NAND2_X2 _f_permutation__U1901  ( .A1(_f_permutation__round_out[247]), .A2(
        _f_permutation__n7150 ), .ZN(_f_permutation__n2706 ) );
  NAND2_X2 _f_permutation__U1900  ( .A1(SYNOPSYS_UNCONNECTED_841), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2707 ) );
  NAND2_X2 _f_permutation__U1899  ( .A1(_f_permutation__n2706 ), .A2(
        _f_permutation__n2707 ), .ZN(_f_permutation__n5140 ) );
  NAND2_X2 _f_permutation__U1898  ( .A1(_f_permutation__round_out[246]), .A2(
        _f_permutation__n7146 ), .ZN(_f_permutation__n2704 ) );
  NAND2_X2 _f_permutation__U1897  ( .A1(SYNOPSYS_UNCONNECTED_842), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2705 ) );
  NAND2_X2 _f_permutation__U1896  ( .A1(_f_permutation__n2704 ), .A2(
        _f_permutation__n2705 ), .ZN(_f_permutation__n5141 ) );
  NAND2_X2 _f_permutation__U1895  ( .A1(_f_permutation__round_out[245]), .A2(
        _f_permutation__n7145 ), .ZN(_f_permutation__n2702 ) );
  NAND2_X2 _f_permutation__U1894  ( .A1(SYNOPSYS_UNCONNECTED_843), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2703 ) );
  NAND2_X2 _f_permutation__U1893  ( .A1(_f_permutation__n2702 ), .A2(
        _f_permutation__n2703 ), .ZN(_f_permutation__n5142 ) );
  NAND2_X2 _f_permutation__U1892  ( .A1(_f_permutation__round_out[244]), .A2(
        _f_permutation__n7144 ), .ZN(_f_permutation__n2700 ) );
  NAND2_X2 _f_permutation__U1891  ( .A1(SYNOPSYS_UNCONNECTED_844), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2701 ) );
  NAND2_X2 _f_permutation__U1890  ( .A1(_f_permutation__n2700 ), .A2(
        _f_permutation__n2701 ), .ZN(_f_permutation__n5143 ) );
  NAND2_X2 _f_permutation__U1889  ( .A1(_f_permutation__round_out[243]), .A2(
        _f_permutation__n7143 ), .ZN(_f_permutation__n2698 ) );
  NAND2_X2 _f_permutation__U1888  ( .A1(SYNOPSYS_UNCONNECTED_845), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2699 ) );
  NAND2_X2 _f_permutation__U1887  ( .A1(_f_permutation__n2698 ), .A2(
        _f_permutation__n2699 ), .ZN(_f_permutation__n5144 ) );
  NAND2_X2 _f_permutation__U1886  ( .A1(_f_permutation__round_out[242]), .A2(
        _f_permutation__n7163 ), .ZN(_f_permutation__n2696 ) );
  NAND2_X2 _f_permutation__U1885  ( .A1(SYNOPSYS_UNCONNECTED_846), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2697 ) );
  NAND2_X2 _f_permutation__U1884  ( .A1(_f_permutation__n2696 ), .A2(
        _f_permutation__n2697 ), .ZN(_f_permutation__n5145 ) );
  NAND2_X2 _f_permutation__U1883  ( .A1(_f_permutation__round_out[241]), .A2(
        _f_permutation__n7162 ), .ZN(_f_permutation__n2694 ) );
  NAND2_X2 _f_permutation__U1882  ( .A1(SYNOPSYS_UNCONNECTED_847), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2695 ) );
  NAND2_X2 _f_permutation__U1881  ( .A1(_f_permutation__n2694 ), .A2(
        _f_permutation__n2695 ), .ZN(_f_permutation__n5146 ) );
  NAND2_X2 _f_permutation__U1880  ( .A1(_f_permutation__round_out[240]), .A2(
        _f_permutation__n7167 ), .ZN(_f_permutation__n2692 ) );
  NAND2_X2 _f_permutation__U1879  ( .A1(SYNOPSYS_UNCONNECTED_848), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2693 ) );
  NAND2_X2 _f_permutation__U1878  ( .A1(_f_permutation__n2692 ), .A2(
        _f_permutation__n2693 ), .ZN(_f_permutation__n5147 ) );
  NAND2_X2 _f_permutation__U1877  ( .A1(_f_permutation__round_out[239]), .A2(
        _f_permutation__n7166 ), .ZN(_f_permutation__n2690 ) );
  NAND2_X2 _f_permutation__U1876  ( .A1(SYNOPSYS_UNCONNECTED_849), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2691 ) );
  NAND2_X2 _f_permutation__U1875  ( .A1(_f_permutation__n2690 ), .A2(
        _f_permutation__n2691 ), .ZN(_f_permutation__n5148 ) );
  NAND2_X2 _f_permutation__U1874  ( .A1(_f_permutation__round_out[238]), .A2(
        _f_permutation__n7165 ), .ZN(_f_permutation__n2688 ) );
  NAND2_X2 _f_permutation__U1873  ( .A1(SYNOPSYS_UNCONNECTED_850), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2689 ) );
  NAND2_X2 _f_permutation__U1872  ( .A1(_f_permutation__n2688 ), .A2(
        _f_permutation__n2689 ), .ZN(_f_permutation__n5149 ) );
  NAND2_X2 _f_permutation__U1871  ( .A1(_f_permutation__round_out[237]), .A2(
        _f_permutation__n7164 ), .ZN(_f_permutation__n2686 ) );
  NAND2_X2 _f_permutation__U1870  ( .A1(SYNOPSYS_UNCONNECTED_851), .A2(
        _f_permutation__n7285 ), .ZN(_f_permutation__n2687 ) );
  NAND2_X2 _f_permutation__U1869  ( .A1(_f_permutation__n2686 ), .A2(
        _f_permutation__n2687 ), .ZN(_f_permutation__n5150 ) );
  NAND2_X2 _f_permutation__U1868  ( .A1(_f_permutation__round_out[236]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n2684 ) );
  NAND2_X2 _f_permutation__U1867  ( .A1(SYNOPSYS_UNCONNECTED_852), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2685 ) );
  NAND2_X2 _f_permutation__U1866  ( .A1(_f_permutation__n2684 ), .A2(
        _f_permutation__n2685 ), .ZN(_f_permutation__n5151 ) );
  NAND2_X2 _f_permutation__U1865  ( .A1(_f_permutation__round_out[235]), .A2(
        _f_permutation__n7168 ), .ZN(_f_permutation__n2682 ) );
  NAND2_X2 _f_permutation__U1864  ( .A1(SYNOPSYS_UNCONNECTED_853), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2683 ) );
  NAND2_X2 _f_permutation__U1863  ( .A1(_f_permutation__n2682 ), .A2(
        _f_permutation__n2683 ), .ZN(_f_permutation__n5152 ) );
  NAND2_X2 _f_permutation__U1862  ( .A1(_f_permutation__round_out[234]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n2680 ) );
  NAND2_X2 _f_permutation__U1861  ( .A1(SYNOPSYS_UNCONNECTED_854), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2681 ) );
  NAND2_X2 _f_permutation__U1860  ( .A1(_f_permutation__n2680 ), .A2(
        _f_permutation__n2681 ), .ZN(_f_permutation__n5153 ) );
  NAND2_X2 _f_permutation__U1859  ( .A1(_f_permutation__round_out[233]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n2678 ) );
  NAND2_X2 _f_permutation__U1858  ( .A1(SYNOPSYS_UNCONNECTED_855), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2679 ) );
  NAND2_X2 _f_permutation__U1857  ( .A1(_f_permutation__n2678 ), .A2(
        _f_permutation__n2679 ), .ZN(_f_permutation__n5154 ) );
  NAND2_X2 _f_permutation__U1856  ( .A1(_f_permutation__round_out[232]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n2676 ) );
  NAND2_X2 _f_permutation__U1855  ( .A1(SYNOPSYS_UNCONNECTED_856), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2677 ) );
  NAND2_X2 _f_permutation__U1854  ( .A1(_f_permutation__n2676 ), .A2(
        _f_permutation__n2677 ), .ZN(_f_permutation__n5155 ) );
  NAND2_X2 _f_permutation__U1853  ( .A1(_f_permutation__round_out[231]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n2674 ) );
  NAND2_X2 _f_permutation__U1852  ( .A1(SYNOPSYS_UNCONNECTED_857), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2675 ) );
  NAND2_X2 _f_permutation__U1851  ( .A1(_f_permutation__n2674 ), .A2(
        _f_permutation__n2675 ), .ZN(_f_permutation__n5156 ) );
  NAND2_X2 _f_permutation__U1850  ( .A1(_f_permutation__round_out[230]), .A2(
        _f_permutation__n7153 ), .ZN(_f_permutation__n2672 ) );
  NAND2_X2 _f_permutation__U1849  ( .A1(SYNOPSYS_UNCONNECTED_858), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2673 ) );
  NAND2_X2 _f_permutation__U1848  ( .A1(_f_permutation__n2672 ), .A2(
        _f_permutation__n2673 ), .ZN(_f_permutation__n5157 ) );
  NAND2_X2 _f_permutation__U1847  ( .A1(_f_permutation__round_out[229]), .A2(
        _f_permutation__n7149 ), .ZN(_f_permutation__n2670 ) );
  NAND2_X2 _f_permutation__U1846  ( .A1(SYNOPSYS_UNCONNECTED_859), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2671 ) );
  NAND2_X2 _f_permutation__U1845  ( .A1(_f_permutation__n2670 ), .A2(
        _f_permutation__n2671 ), .ZN(_f_permutation__n5158 ) );
  NAND2_X2 _f_permutation__U1844  ( .A1(_f_permutation__round_out[228]), .A2(
        _f_permutation__n7148 ), .ZN(_f_permutation__n2668 ) );
  NAND2_X2 _f_permutation__U1843  ( .A1(SYNOPSYS_UNCONNECTED_860), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2669 ) );
  NAND2_X2 _f_permutation__U1842  ( .A1(_f_permutation__n2668 ), .A2(
        _f_permutation__n2669 ), .ZN(_f_permutation__n5159 ) );
  NAND2_X2 _f_permutation__U1841  ( .A1(_f_permutation__round_out[227]), .A2(
        _f_permutation__n7147 ), .ZN(_f_permutation__n2666 ) );
  NAND2_X2 _f_permutation__U1840  ( .A1(SYNOPSYS_UNCONNECTED_861), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2667 ) );
  NAND2_X2 _f_permutation__U1839  ( .A1(_f_permutation__n2666 ), .A2(
        _f_permutation__n2667 ), .ZN(_f_permutation__n5160 ) );
  NAND2_X2 _f_permutation__U1838  ( .A1(_f_permutation__round_out[226]), .A2(
        _f_permutation__n7152 ), .ZN(_f_permutation__n2664 ) );
  NAND2_X2 _f_permutation__U1837  ( .A1(SYNOPSYS_UNCONNECTED_862), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2665 ) );
  NAND2_X2 _f_permutation__U1836  ( .A1(_f_permutation__n2664 ), .A2(
        _f_permutation__n2665 ), .ZN(_f_permutation__n5161 ) );
  NAND2_X2 _f_permutation__U1835  ( .A1(_f_permutation__round_out[225]), .A2(
        _f_permutation__n7151 ), .ZN(_f_permutation__n2662 ) );
  NAND2_X2 _f_permutation__U1834  ( .A1(SYNOPSYS_UNCONNECTED_863), .A2(
        _f_permutation__n7286 ), .ZN(_f_permutation__n2663 ) );
  NAND2_X2 _f_permutation__U1833  ( .A1(_f_permutation__n2662 ), .A2(
        _f_permutation__n2663 ), .ZN(_f_permutation__n5162 ) );
  NAND2_X2 _f_permutation__U1832  ( .A1(_f_permutation__round_out[224]), .A2(
        _f_permutation__n7150 ), .ZN(_f_permutation__n2660 ) );
  NAND2_X2 _f_permutation__U1831  ( .A1(SYNOPSYS_UNCONNECTED_864), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2661 ) );
  NAND2_X2 _f_permutation__U1830  ( .A1(_f_permutation__n2660 ), .A2(
        _f_permutation__n2661 ), .ZN(_f_permutation__n5163 ) );
  NAND2_X2 _f_permutation__U1829  ( .A1(_f_permutation__round_out[223]), .A2(
        _f_permutation__n7146 ), .ZN(_f_permutation__n2658 ) );
  NAND2_X2 _f_permutation__U1828  ( .A1(SYNOPSYS_UNCONNECTED_865), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2659 ) );
  NAND2_X2 _f_permutation__U1827  ( .A1(_f_permutation__n2658 ), .A2(
        _f_permutation__n2659 ), .ZN(_f_permutation__n5164 ) );
  NAND2_X2 _f_permutation__U1826  ( .A1(_f_permutation__round_out[222]), .A2(
        _f_permutation__n7145 ), .ZN(_f_permutation__n2656 ) );
  NAND2_X2 _f_permutation__U1825  ( .A1(SYNOPSYS_UNCONNECTED_866), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2657 ) );
  NAND2_X2 _f_permutation__U1824  ( .A1(_f_permutation__n2656 ), .A2(
        _f_permutation__n2657 ), .ZN(_f_permutation__n5165 ) );
  NAND2_X2 _f_permutation__U1823  ( .A1(_f_permutation__round_out[221]), .A2(
        _f_permutation__n7144 ), .ZN(_f_permutation__n2654 ) );
  NAND2_X2 _f_permutation__U1822  ( .A1(SYNOPSYS_UNCONNECTED_867), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2655 ) );
  NAND2_X2 _f_permutation__U1821  ( .A1(_f_permutation__n2654 ), .A2(
        _f_permutation__n2655 ), .ZN(_f_permutation__n5166 ) );
  NAND2_X2 _f_permutation__U1820  ( .A1(_f_permutation__round_out[220]), .A2(
        _f_permutation__n7143 ), .ZN(_f_permutation__n2652 ) );
  NAND2_X2 _f_permutation__U1819  ( .A1(SYNOPSYS_UNCONNECTED_868), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2653 ) );
  NAND2_X2 _f_permutation__U1818  ( .A1(_f_permutation__n2652 ), .A2(
        _f_permutation__n2653 ), .ZN(_f_permutation__n5167 ) );
  NAND2_X2 _f_permutation__U1817  ( .A1(_f_permutation__round_out[219]), .A2(
        _f_permutation__n7163 ), .ZN(_f_permutation__n2650 ) );
  NAND2_X2 _f_permutation__U1816  ( .A1(SYNOPSYS_UNCONNECTED_869), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2651 ) );
  NAND2_X2 _f_permutation__U1815  ( .A1(_f_permutation__n2650 ), .A2(
        _f_permutation__n2651 ), .ZN(_f_permutation__n5168 ) );
  NAND2_X2 _f_permutation__U1814  ( .A1(_f_permutation__round_out[218]), .A2(
        _f_permutation__n7156 ), .ZN(_f_permutation__n2648 ) );
  NAND2_X2 _f_permutation__U1813  ( .A1(SYNOPSYS_UNCONNECTED_870), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2649 ) );
  NAND2_X2 _f_permutation__U1812  ( .A1(_f_permutation__n2648 ), .A2(
        _f_permutation__n2649 ), .ZN(_f_permutation__n5169 ) );
  NAND2_X2 _f_permutation__U1811  ( .A1(_f_permutation__round_out[217]), .A2(
        _f_permutation__n7141 ), .ZN(_f_permutation__n2646 ) );
  NAND2_X2 _f_permutation__U1810  ( .A1(SYNOPSYS_UNCONNECTED_871), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2647 ) );
  NAND2_X2 _f_permutation__U1809  ( .A1(_f_permutation__n2646 ), .A2(
        _f_permutation__n2647 ), .ZN(_f_permutation__n5170 ) );
  NAND2_X2 _f_permutation__U1808  ( .A1(_f_permutation__round_out[216]), .A2(
        _f_permutation__n7140 ), .ZN(_f_permutation__n2644 ) );
  NAND2_X2 _f_permutation__U1807  ( .A1(SYNOPSYS_UNCONNECTED_872), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2645 ) );
  NAND2_X2 _f_permutation__U1806  ( .A1(_f_permutation__n2644 ), .A2(
        _f_permutation__n2645 ), .ZN(_f_permutation__n5171 ) );
  NAND2_X2 _f_permutation__U1805  ( .A1(_f_permutation__round_out[215]), .A2(
        _f_permutation__n7139 ), .ZN(_f_permutation__n2642 ) );
  NAND2_X2 _f_permutation__U1804  ( .A1(SYNOPSYS_UNCONNECTED_873), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2643 ) );
  NAND2_X2 _f_permutation__U1803  ( .A1(_f_permutation__n2642 ), .A2(
        _f_permutation__n2643 ), .ZN(_f_permutation__n5172 ) );
  NAND2_X2 _f_permutation__U1802  ( .A1(_f_permutation__round_out[214]), .A2(
        _f_permutation__n7142 ), .ZN(_f_permutation__n2640 ) );
  NAND2_X2 _f_permutation__U1801  ( .A1(SYNOPSYS_UNCONNECTED_874), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2641 ) );
  NAND2_X2 _f_permutation__U1800  ( .A1(_f_permutation__n2640 ), .A2(
        _f_permutation__n2641 ), .ZN(_f_permutation__n5173 ) );
  NAND2_X2 _f_permutation__U1799  ( .A1(_f_permutation__round_out[213]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n2638 ) );
  NAND2_X2 _f_permutation__U1798  ( .A1(SYNOPSYS_UNCONNECTED_875), .A2(
        _f_permutation__n7287 ), .ZN(_f_permutation__n2639 ) );
  NAND2_X2 _f_permutation__U1797  ( .A1(_f_permutation__n2638 ), .A2(
        _f_permutation__n2639 ), .ZN(_f_permutation__n5174 ) );
  NAND2_X2 _f_permutation__U1796  ( .A1(_f_permutation__round_out[212]), .A2(
        _f_permutation__n7153 ), .ZN(_f_permutation__n2636 ) );
  NAND2_X2 _f_permutation__U1795  ( .A1(SYNOPSYS_UNCONNECTED_876), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2637 ) );
  NAND2_X2 _f_permutation__U1794  ( .A1(_f_permutation__n2636 ), .A2(
        _f_permutation__n2637 ), .ZN(_f_permutation__n5175 ) );
  NAND2_X2 _f_permutation__U1793  ( .A1(_f_permutation__round_out[211]), .A2(
        _f_permutation__n7161 ), .ZN(_f_permutation__n2634 ) );
  NAND2_X2 _f_permutation__U1792  ( .A1(SYNOPSYS_UNCONNECTED_877), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2635 ) );
  NAND2_X2 _f_permutation__U1791  ( .A1(_f_permutation__n2634 ), .A2(
        _f_permutation__n2635 ), .ZN(_f_permutation__n5176 ) );
  NAND2_X2 _f_permutation__U1790  ( .A1(_f_permutation__round_out[210]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n2632 ) );
  NAND2_X2 _f_permutation__U1789  ( .A1(SYNOPSYS_UNCONNECTED_878), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2633 ) );
  NAND2_X2 _f_permutation__U1788  ( .A1(_f_permutation__n2632 ), .A2(
        _f_permutation__n2633 ), .ZN(_f_permutation__n5177 ) );
  NAND2_X2 _f_permutation__U1787  ( .A1(_f_permutation__round_out[209]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n2630 ) );
  NAND2_X2 _f_permutation__U1786  ( .A1(SYNOPSYS_UNCONNECTED_879), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2631 ) );
  NAND2_X2 _f_permutation__U1785  ( .A1(_f_permutation__n2630 ), .A2(
        _f_permutation__n2631 ), .ZN(_f_permutation__n5178 ) );
  NAND2_X2 _f_permutation__U1784  ( .A1(_f_permutation__round_out[208]), .A2(
        _f_permutation__n7154 ), .ZN(_f_permutation__n2628 ) );
  NAND2_X2 _f_permutation__U1783  ( .A1(SYNOPSYS_UNCONNECTED_880), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2629 ) );
  NAND2_X2 _f_permutation__U1782  ( .A1(_f_permutation__n2628 ), .A2(
        _f_permutation__n2629 ), .ZN(_f_permutation__n5179 ) );
  NAND2_X2 _f_permutation__U1781  ( .A1(_f_permutation__round_out[207]), .A2(
        _f_permutation__n7156 ), .ZN(_f_permutation__n2626 ) );
  NAND2_X2 _f_permutation__U1780  ( .A1(SYNOPSYS_UNCONNECTED_881), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2627 ) );
  NAND2_X2 _f_permutation__U1779  ( .A1(_f_permutation__n2626 ), .A2(
        _f_permutation__n2627 ), .ZN(_f_permutation__n5180 ) );
  NAND2_X2 _f_permutation__U1778  ( .A1(_f_permutation__round_out[206]), .A2(
        _f_permutation__n7141 ), .ZN(_f_permutation__n2624 ) );
  NAND2_X2 _f_permutation__U1777  ( .A1(SYNOPSYS_UNCONNECTED_882), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2625 ) );
  NAND2_X2 _f_permutation__U1776  ( .A1(_f_permutation__n2624 ), .A2(
        _f_permutation__n2625 ), .ZN(_f_permutation__n5181 ) );
  NAND2_X2 _f_permutation__U1775  ( .A1(_f_permutation__round_out[205]), .A2(
        _f_permutation__n7140 ), .ZN(_f_permutation__n2622 ) );
  NAND2_X2 _f_permutation__U1774  ( .A1(SYNOPSYS_UNCONNECTED_883), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2623 ) );
  NAND2_X2 _f_permutation__U1773  ( .A1(_f_permutation__n2622 ), .A2(
        _f_permutation__n2623 ), .ZN(_f_permutation__n5182 ) );
  NAND2_X2 _f_permutation__U1772  ( .A1(_f_permutation__round_out[204]), .A2(
        _f_permutation__n7139 ), .ZN(_f_permutation__n2620 ) );
  NAND2_X2 _f_permutation__U1771  ( .A1(SYNOPSYS_UNCONNECTED_884), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2621 ) );
  NAND2_X2 _f_permutation__U1770  ( .A1(_f_permutation__n2620 ), .A2(
        _f_permutation__n2621 ), .ZN(_f_permutation__n5183 ) );
  NAND2_X2 _f_permutation__U1769  ( .A1(_f_permutation__round_out[203]), .A2(
        _f_permutation__n7142 ), .ZN(_f_permutation__n2618 ) );
  NAND2_X2 _f_permutation__U1768  ( .A1(SYNOPSYS_UNCONNECTED_885), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2619 ) );
  NAND2_X2 _f_permutation__U1767  ( .A1(_f_permutation__n2618 ), .A2(
        _f_permutation__n2619 ), .ZN(_f_permutation__n5184 ) );
  NAND2_X2 _f_permutation__U1766  ( .A1(_f_permutation__round_out[202]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n2616 ) );
  NAND2_X2 _f_permutation__U1765  ( .A1(SYNOPSYS_UNCONNECTED_886), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2617 ) );
  NAND2_X2 _f_permutation__U1764  ( .A1(_f_permutation__n2616 ), .A2(
        _f_permutation__n2617 ), .ZN(_f_permutation__n5185 ) );
  NAND2_X2 _f_permutation__U1763  ( .A1(_f_permutation__round_out[201]), .A2(
        _f_permutation__n7148 ), .ZN(_f_permutation__n2614 ) );
  NAND2_X2 _f_permutation__U1762  ( .A1(SYNOPSYS_UNCONNECTED_887), .A2(
        _f_permutation__n7288 ), .ZN(_f_permutation__n2615 ) );
  NAND2_X2 _f_permutation__U1761  ( .A1(_f_permutation__n2614 ), .A2(
        _f_permutation__n2615 ), .ZN(_f_permutation__n5186 ) );
  NAND2_X2 _f_permutation__U1760  ( .A1(_f_permutation__round_out[200]), .A2(
        _f_permutation__n7149 ), .ZN(_f_permutation__n2612 ) );
  NAND2_X2 _f_permutation__U1759  ( .A1(SYNOPSYS_UNCONNECTED_888), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2613 ) );
  NAND2_X2 _f_permutation__U1758  ( .A1(_f_permutation__n2612 ), .A2(
        _f_permutation__n2613 ), .ZN(_f_permutation__n5187 ) );
  NAND2_X2 _f_permutation__U1757  ( .A1(_f_permutation__round_out[199]), .A2(
        _f_permutation__n7148 ), .ZN(_f_permutation__n2610 ) );
  NAND2_X2 _f_permutation__U1756  ( .A1(SYNOPSYS_UNCONNECTED_889), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2611 ) );
  NAND2_X2 _f_permutation__U1755  ( .A1(_f_permutation__n2610 ), .A2(
        _f_permutation__n2611 ), .ZN(_f_permutation__n5188 ) );
  NAND2_X2 _f_permutation__U1754  ( .A1(_f_permutation__round_out[198]), .A2(
        _f_permutation__n7147 ), .ZN(_f_permutation__n2608 ) );
  NAND2_X2 _f_permutation__U1753  ( .A1(SYNOPSYS_UNCONNECTED_890), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2609 ) );
  NAND2_X2 _f_permutation__U1752  ( .A1(_f_permutation__n2608 ), .A2(
        _f_permutation__n2609 ), .ZN(_f_permutation__n5189 ) );
  NAND2_X2 _f_permutation__U1751  ( .A1(_f_permutation__round_out[197]), .A2(
        _f_permutation__n7152 ), .ZN(_f_permutation__n2606 ) );
  NAND2_X2 _f_permutation__U1750  ( .A1(SYNOPSYS_UNCONNECTED_891), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2607 ) );
  NAND2_X2 _f_permutation__U1749  ( .A1(_f_permutation__n2606 ), .A2(
        _f_permutation__n2607 ), .ZN(_f_permutation__n5190 ) );
  NAND2_X2 _f_permutation__U1748  ( .A1(_f_permutation__round_out[196]), .A2(
        _f_permutation__n7151 ), .ZN(_f_permutation__n2604 ) );
  NAND2_X2 _f_permutation__U1747  ( .A1(SYNOPSYS_UNCONNECTED_892), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2605 ) );
  NAND2_X2 _f_permutation__U1746  ( .A1(_f_permutation__n2604 ), .A2(
        _f_permutation__n2605 ), .ZN(_f_permutation__n5191 ) );
  NAND2_X2 _f_permutation__U1745  ( .A1(_f_permutation__round_out[195]), .A2(
        _f_permutation__n7150 ), .ZN(_f_permutation__n2602 ) );
  NAND2_X2 _f_permutation__U1744  ( .A1(SYNOPSYS_UNCONNECTED_893), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2603 ) );
  NAND2_X2 _f_permutation__U1743  ( .A1(_f_permutation__n2602 ), .A2(
        _f_permutation__n2603 ), .ZN(_f_permutation__n5192 ) );
  NAND2_X2 _f_permutation__U1742  ( .A1(_f_permutation__round_out[194]), .A2(
        _f_permutation__n7146 ), .ZN(_f_permutation__n2600 ) );
  NAND2_X2 _f_permutation__U1741  ( .A1(SYNOPSYS_UNCONNECTED_894), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2601 ) );
  NAND2_X2 _f_permutation__U1740  ( .A1(_f_permutation__n2600 ), .A2(
        _f_permutation__n2601 ), .ZN(_f_permutation__n5193 ) );
  NAND2_X2 _f_permutation__U1739  ( .A1(_f_permutation__round_out[193]), .A2(
        _f_permutation__n7145 ), .ZN(_f_permutation__n2598 ) );
  NAND2_X2 _f_permutation__U1738  ( .A1(SYNOPSYS_UNCONNECTED_895), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2599 ) );
  NAND2_X2 _f_permutation__U1737  ( .A1(_f_permutation__n2598 ), .A2(
        _f_permutation__n2599 ), .ZN(_f_permutation__n5194 ) );
  NAND2_X2 _f_permutation__U1736  ( .A1(_f_permutation__round_out[192]), .A2(
        _f_permutation__n7144 ), .ZN(_f_permutation__n2596 ) );
  NAND2_X2 _f_permutation__U1735  ( .A1(SYNOPSYS_UNCONNECTED_896), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2597 ) );
  NAND2_X2 _f_permutation__U1734  ( .A1(_f_permutation__n2596 ), .A2(
        _f_permutation__n2597 ), .ZN(_f_permutation__n5195 ) );
  NAND2_X2 _f_permutation__U1733  ( .A1(_f_permutation__round_out[191]), .A2(
        _f_permutation__n7143 ), .ZN(_f_permutation__n2594 ) );
  NAND2_X2 _f_permutation__U1732  ( .A1(SYNOPSYS_UNCONNECTED_897), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2595 ) );
  NAND2_X2 _f_permutation__U1731  ( .A1(_f_permutation__n2594 ), .A2(
        _f_permutation__n2595 ), .ZN(_f_permutation__n5196 ) );
  NAND2_X2 _f_permutation__U1730  ( .A1(_f_permutation__round_out[190]), .A2(
        _f_permutation__n7163 ), .ZN(_f_permutation__n2592 ) );
  NAND2_X2 _f_permutation__U1729  ( .A1(SYNOPSYS_UNCONNECTED_898), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2593 ) );
  NAND2_X2 _f_permutation__U1728  ( .A1(_f_permutation__n2592 ), .A2(
        _f_permutation__n2593 ), .ZN(_f_permutation__n5197 ) );
  NAND2_X2 _f_permutation__U1727  ( .A1(_f_permutation__round_out[189]), .A2(
        _f_permutation__n7162 ), .ZN(_f_permutation__n2590 ) );
  NAND2_X2 _f_permutation__U1726  ( .A1(SYNOPSYS_UNCONNECTED_899), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2591 ) );
  NAND2_X2 _f_permutation__U1725  ( .A1(_f_permutation__n2590 ), .A2(
        _f_permutation__n2591 ), .ZN(_f_permutation__n5198 ) );
  NAND2_X2 _f_permutation__U1724  ( .A1(_f_permutation__round_out[188]), .A2(
        _f_permutation__n7156 ), .ZN(_f_permutation__n2588 ) );
  NAND2_X2 _f_permutation__U1723  ( .A1(SYNOPSYS_UNCONNECTED_900), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2589 ) );
  NAND2_X2 _f_permutation__U1722  ( .A1(_f_permutation__n2588 ), .A2(
        _f_permutation__n2589 ), .ZN(_f_permutation__n5199 ) );
  NAND2_X2 _f_permutation__U1721  ( .A1(_f_permutation__round_out[187]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n2586 ) );
  NAND2_X2 _f_permutation__U1720  ( .A1(SYNOPSYS_UNCONNECTED_901), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2587 ) );
  NAND2_X2 _f_permutation__U1719  ( .A1(_f_permutation__n2586 ), .A2(
        _f_permutation__n2587 ), .ZN(_f_permutation__n5200 ) );
  NAND2_X2 _f_permutation__U1718  ( .A1(_f_permutation__round_out[186]), .A2(
        _f_permutation__n7154 ), .ZN(_f_permutation__n2584 ) );
  NAND2_X2 _f_permutation__U1717  ( .A1(SYNOPSYS_UNCONNECTED_902), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2585 ) );
  NAND2_X2 _f_permutation__U1716  ( .A1(_f_permutation__n2584 ), .A2(
        _f_permutation__n2585 ), .ZN(_f_permutation__n5201 ) );
  NAND2_X2 _f_permutation__U1715  ( .A1(_f_permutation__round_out[185]), .A2(
        _f_permutation__n7161 ), .ZN(_f_permutation__n2582 ) );
  NAND2_X2 _f_permutation__U1714  ( .A1(SYNOPSYS_UNCONNECTED_903), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2583 ) );
  NAND2_X2 _f_permutation__U1713  ( .A1(_f_permutation__n2582 ), .A2(
        _f_permutation__n2583 ), .ZN(_f_permutation__n5202 ) );
  NAND2_X2 _f_permutation__U1712  ( .A1(_f_permutation__round_out[184]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n2580 ) );
  NAND2_X2 _f_permutation__U1711  ( .A1(SYNOPSYS_UNCONNECTED_904), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2581 ) );
  NAND2_X2 _f_permutation__U1710  ( .A1(_f_permutation__n2580 ), .A2(
        _f_permutation__n2581 ), .ZN(_f_permutation__n5203 ) );
  NAND2_X2 _f_permutation__U1709  ( .A1(_f_permutation__round_out[183]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2578 ) );
  NAND2_X2 _f_permutation__U1708  ( .A1(SYNOPSYS_UNCONNECTED_905), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2579 ) );
  NAND2_X2 _f_permutation__U1707  ( .A1(_f_permutation__n2578 ), .A2(
        _f_permutation__n2579 ), .ZN(_f_permutation__n5204 ) );
  NAND2_X2 _f_permutation__U1706  ( .A1(_f_permutation__round_out[182]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2576 ) );
  NAND2_X2 _f_permutation__U1705  ( .A1(SYNOPSYS_UNCONNECTED_906), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2577 ) );
  NAND2_X2 _f_permutation__U1704  ( .A1(_f_permutation__n2576 ), .A2(
        _f_permutation__n2577 ), .ZN(_f_permutation__n5205 ) );
  NAND2_X2 _f_permutation__U1703  ( .A1(_f_permutation__round_out[181]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2574 ) );
  NAND2_X2 _f_permutation__U1702  ( .A1(SYNOPSYS_UNCONNECTED_907), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2575 ) );
  NAND2_X2 _f_permutation__U1701  ( .A1(_f_permutation__n2574 ), .A2(
        _f_permutation__n2575 ), .ZN(_f_permutation__n5206 ) );
  NAND2_X2 _f_permutation__U1700  ( .A1(_f_permutation__round_out[180]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2572 ) );
  NAND2_X2 _f_permutation__U1699  ( .A1(SYNOPSYS_UNCONNECTED_908), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2573 ) );
  NAND2_X2 _f_permutation__U1698  ( .A1(_f_permutation__n2572 ), .A2(
        _f_permutation__n2573 ), .ZN(_f_permutation__n5207 ) );
  NAND2_X2 _f_permutation__U1697  ( .A1(_f_permutation__round_out[179]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2570 ) );
  NAND2_X2 _f_permutation__U1696  ( .A1(SYNOPSYS_UNCONNECTED_909), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2571 ) );
  NAND2_X2 _f_permutation__U1695  ( .A1(_f_permutation__n2570 ), .A2(
        _f_permutation__n2571 ), .ZN(_f_permutation__n5208 ) );
  NAND2_X2 _f_permutation__U1694  ( .A1(_f_permutation__round_out[178]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2568 ) );
  NAND2_X2 _f_permutation__U1693  ( .A1(SYNOPSYS_UNCONNECTED_910), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2569 ) );
  NAND2_X2 _f_permutation__U1692  ( .A1(_f_permutation__n2568 ), .A2(
        _f_permutation__n2569 ), .ZN(_f_permutation__n5209 ) );
  NAND2_X2 _f_permutation__U1691  ( .A1(_f_permutation__round_out[177]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2566 ) );
  NAND2_X2 _f_permutation__U1690  ( .A1(SYNOPSYS_UNCONNECTED_911), .A2(
        _f_permutation__n7290 ), .ZN(_f_permutation__n2567 ) );
  NAND2_X2 _f_permutation__U1689  ( .A1(_f_permutation__n2566 ), .A2(
        _f_permutation__n2567 ), .ZN(_f_permutation__n5210 ) );
  NAND2_X2 _f_permutation__U1688  ( .A1(_f_permutation__round_out[176]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2564 ) );
  NAND2_X2 _f_permutation__U1687  ( .A1(SYNOPSYS_UNCONNECTED_912), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2565 ) );
  NAND2_X2 _f_permutation__U1686  ( .A1(_f_permutation__n2564 ), .A2(
        _f_permutation__n2565 ), .ZN(_f_permutation__n5211 ) );
  NAND2_X2 _f_permutation__U1685  ( .A1(_f_permutation__round_out[175]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2562 ) );
  NAND2_X2 _f_permutation__U1684  ( .A1(SYNOPSYS_UNCONNECTED_913), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2563 ) );
  NAND2_X2 _f_permutation__U1683  ( .A1(_f_permutation__n2562 ), .A2(
        _f_permutation__n2563 ), .ZN(_f_permutation__n5212 ) );
  NAND2_X2 _f_permutation__U1682  ( .A1(_f_permutation__round_out[174]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2560 ) );
  NAND2_X2 _f_permutation__U1681  ( .A1(SYNOPSYS_UNCONNECTED_914), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2561 ) );
  NAND2_X2 _f_permutation__U1680  ( .A1(_f_permutation__n2560 ), .A2(
        _f_permutation__n2561 ), .ZN(_f_permutation__n5213 ) );
  NAND2_X2 _f_permutation__U1679  ( .A1(_f_permutation__round_out[173]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2558 ) );
  NAND2_X2 _f_permutation__U1678  ( .A1(SYNOPSYS_UNCONNECTED_915), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2559 ) );
  NAND2_X2 _f_permutation__U1677  ( .A1(_f_permutation__n2558 ), .A2(
        _f_permutation__n2559 ), .ZN(_f_permutation__n5214 ) );
  NAND2_X2 _f_permutation__U1676  ( .A1(_f_permutation__round_out[172]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2556 ) );
  NAND2_X2 _f_permutation__U1675  ( .A1(SYNOPSYS_UNCONNECTED_916), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2557 ) );
  NAND2_X2 _f_permutation__U1674  ( .A1(_f_permutation__n2556 ), .A2(
        _f_permutation__n2557 ), .ZN(_f_permutation__n5215 ) );
  NAND2_X2 _f_permutation__U1673  ( .A1(_f_permutation__round_out[171]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2554 ) );
  NAND2_X2 _f_permutation__U1672  ( .A1(SYNOPSYS_UNCONNECTED_917), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2555 ) );
  NAND2_X2 _f_permutation__U1671  ( .A1(_f_permutation__n2554 ), .A2(
        _f_permutation__n2555 ), .ZN(_f_permutation__n5216 ) );
  NAND2_X2 _f_permutation__U1670  ( .A1(_f_permutation__round_out[170]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2552 ) );
  NAND2_X2 _f_permutation__U1669  ( .A1(SYNOPSYS_UNCONNECTED_918), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2553 ) );
  NAND2_X2 _f_permutation__U1668  ( .A1(_f_permutation__n2552 ), .A2(
        _f_permutation__n2553 ), .ZN(_f_permutation__n5217 ) );
  NAND2_X2 _f_permutation__U1667  ( .A1(_f_permutation__round_out[169]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2550 ) );
  NAND2_X2 _f_permutation__U1666  ( .A1(SYNOPSYS_UNCONNECTED_919), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2551 ) );
  NAND2_X2 _f_permutation__U1665  ( .A1(_f_permutation__n2550 ), .A2(
        _f_permutation__n2551 ), .ZN(_f_permutation__n5218 ) );
  NAND2_X2 _f_permutation__U1664  ( .A1(_f_permutation__round_out[168]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2548 ) );
  NAND2_X2 _f_permutation__U1663  ( .A1(SYNOPSYS_UNCONNECTED_920), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2549 ) );
  NAND2_X2 _f_permutation__U1662  ( .A1(_f_permutation__n2548 ), .A2(
        _f_permutation__n2549 ), .ZN(_f_permutation__n5219 ) );
  NAND2_X2 _f_permutation__U1661  ( .A1(_f_permutation__round_out[167]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2546 ) );
  NAND2_X2 _f_permutation__U1660  ( .A1(SYNOPSYS_UNCONNECTED_921), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2547 ) );
  NAND2_X2 _f_permutation__U1659  ( .A1(_f_permutation__n2546 ), .A2(
        _f_permutation__n2547 ), .ZN(_f_permutation__n5220 ) );
  NAND2_X2 _f_permutation__U1658  ( .A1(_f_permutation__round_out[166]), .A2(
        _f_permutation__n7086 ), .ZN(_f_permutation__n2544 ) );
  NAND2_X2 _f_permutation__U1657  ( .A1(SYNOPSYS_UNCONNECTED_922), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2545 ) );
  NAND2_X2 _f_permutation__U1656  ( .A1(_f_permutation__n2544 ), .A2(
        _f_permutation__n2545 ), .ZN(_f_permutation__n5221 ) );
  NAND2_X2 _f_permutation__U1655  ( .A1(_f_permutation__round_out[165]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n2542 ) );
  NAND2_X2 _f_permutation__U1654  ( .A1(SYNOPSYS_UNCONNECTED_923), .A2(
        _f_permutation__n7291 ), .ZN(_f_permutation__n2543 ) );
  NAND2_X2 _f_permutation__U1653  ( .A1(_f_permutation__n2542 ), .A2(
        _f_permutation__n2543 ), .ZN(_f_permutation__n5222 ) );
  NAND2_X2 _f_permutation__U1652  ( .A1(_f_permutation__round_out[164]), .A2(
        _f_permutation__n7151 ), .ZN(_f_permutation__n2540 ) );
  NAND2_X2 _f_permutation__U1651  ( .A1(SYNOPSYS_UNCONNECTED_924), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2541 ) );
  NAND2_X2 _f_permutation__U1650  ( .A1(_f_permutation__n2540 ), .A2(
        _f_permutation__n2541 ), .ZN(_f_permutation__n5223 ) );
  NAND2_X2 _f_permutation__U1649  ( .A1(_f_permutation__round_out[163]), .A2(
        _f_permutation__n7150 ), .ZN(_f_permutation__n2538 ) );
  NAND2_X2 _f_permutation__U1648  ( .A1(SYNOPSYS_UNCONNECTED_925), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2539 ) );
  NAND2_X2 _f_permutation__U1647  ( .A1(_f_permutation__n2538 ), .A2(
        _f_permutation__n2539 ), .ZN(_f_permutation__n5224 ) );
  NAND2_X2 _f_permutation__U1646  ( .A1(_f_permutation__round_out[162]), .A2(
        _f_permutation__n7146 ), .ZN(_f_permutation__n2536 ) );
  NAND2_X2 _f_permutation__U1645  ( .A1(SYNOPSYS_UNCONNECTED_926), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2537 ) );
  NAND2_X2 _f_permutation__U1644  ( .A1(_f_permutation__n2536 ), .A2(
        _f_permutation__n2537 ), .ZN(_f_permutation__n5225 ) );
  NAND2_X2 _f_permutation__U1643  ( .A1(_f_permutation__round_out[161]), .A2(
        _f_permutation__n7145 ), .ZN(_f_permutation__n2534 ) );
  NAND2_X2 _f_permutation__U1642  ( .A1(SYNOPSYS_UNCONNECTED_927), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2535 ) );
  NAND2_X2 _f_permutation__U1641  ( .A1(_f_permutation__n2534 ), .A2(
        _f_permutation__n2535 ), .ZN(_f_permutation__n5226 ) );
  NAND2_X2 _f_permutation__U1640  ( .A1(_f_permutation__round_out[160]), .A2(
        _f_permutation__n7144 ), .ZN(_f_permutation__n2532 ) );
  NAND2_X2 _f_permutation__U1639  ( .A1(SYNOPSYS_UNCONNECTED_928), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2533 ) );
  NAND2_X2 _f_permutation__U1638  ( .A1(_f_permutation__n2532 ), .A2(
        _f_permutation__n2533 ), .ZN(_f_permutation__n5227 ) );
  NAND2_X2 _f_permutation__U1637  ( .A1(_f_permutation__round_out[159]), .A2(
        _f_permutation__n7143 ), .ZN(_f_permutation__n2530 ) );
  NAND2_X2 _f_permutation__U1636  ( .A1(SYNOPSYS_UNCONNECTED_929), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2531 ) );
  NAND2_X2 _f_permutation__U1635  ( .A1(_f_permutation__n2530 ), .A2(
        _f_permutation__n2531 ), .ZN(_f_permutation__n5228 ) );
  NAND2_X2 _f_permutation__U1634  ( .A1(_f_permutation__round_out[158]), .A2(
        _f_permutation__n7163 ), .ZN(_f_permutation__n2528 ) );
  NAND2_X2 _f_permutation__U1633  ( .A1(SYNOPSYS_UNCONNECTED_930), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2529 ) );
  NAND2_X2 _f_permutation__U1632  ( .A1(_f_permutation__n2528 ), .A2(
        _f_permutation__n2529 ), .ZN(_f_permutation__n5229 ) );
  NAND2_X2 _f_permutation__U1631  ( .A1(_f_permutation__round_out[157]), .A2(
        _f_permutation__n7162 ), .ZN(_f_permutation__n2526 ) );
  NAND2_X2 _f_permutation__U1630  ( .A1(SYNOPSYS_UNCONNECTED_931), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2527 ) );
  NAND2_X2 _f_permutation__U1629  ( .A1(_f_permutation__n2526 ), .A2(
        _f_permutation__n2527 ), .ZN(_f_permutation__n5230 ) );
  NAND2_X2 _f_permutation__U1628  ( .A1(_f_permutation__round_out[156]), .A2(
        _f_permutation__n7167 ), .ZN(_f_permutation__n2524 ) );
  NAND2_X2 _f_permutation__U1627  ( .A1(SYNOPSYS_UNCONNECTED_932), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2525 ) );
  NAND2_X2 _f_permutation__U1626  ( .A1(_f_permutation__n2524 ), .A2(
        _f_permutation__n2525 ), .ZN(_f_permutation__n5231 ) );
  NAND2_X2 _f_permutation__U1625  ( .A1(_f_permutation__round_out[155]), .A2(
        _f_permutation__n7166 ), .ZN(_f_permutation__n2522 ) );
  NAND2_X2 _f_permutation__U1624  ( .A1(SYNOPSYS_UNCONNECTED_933), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2523 ) );
  NAND2_X2 _f_permutation__U1623  ( .A1(_f_permutation__n2522 ), .A2(
        _f_permutation__n2523 ), .ZN(_f_permutation__n5232 ) );
  NAND2_X2 _f_permutation__U1622  ( .A1(_f_permutation__round_out[154]), .A2(
        _f_permutation__n7165 ), .ZN(_f_permutation__n2520 ) );
  NAND2_X2 _f_permutation__U1621  ( .A1(SYNOPSYS_UNCONNECTED_934), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2521 ) );
  NAND2_X2 _f_permutation__U1620  ( .A1(_f_permutation__n2520 ), .A2(
        _f_permutation__n2521 ), .ZN(_f_permutation__n5233 ) );
  NAND2_X2 _f_permutation__U1619  ( .A1(_f_permutation__round_out[153]), .A2(
        _f_permutation__n7164 ), .ZN(_f_permutation__n2518 ) );
  NAND2_X2 _f_permutation__U1618  ( .A1(SYNOPSYS_UNCONNECTED_935), .A2(
        _f_permutation__n7292 ), .ZN(_f_permutation__n2519 ) );
  NAND2_X2 _f_permutation__U1617  ( .A1(_f_permutation__n2518 ), .A2(
        _f_permutation__n2519 ), .ZN(_f_permutation__n5234 ) );
  NAND2_X2 _f_permutation__U1616  ( .A1(_f_permutation__round_out[152]), .A2(
        _f_permutation__n7156 ), .ZN(_f_permutation__n2516 ) );
  NAND2_X2 _f_permutation__U1615  ( .A1(SYNOPSYS_UNCONNECTED_936), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2517 ) );
  NAND2_X2 _f_permutation__U1614  ( .A1(_f_permutation__n2516 ), .A2(
        _f_permutation__n2517 ), .ZN(_f_permutation__n5235 ) );
  NAND2_X2 _f_permutation__U1613  ( .A1(_f_permutation__round_out[151]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n2514 ) );
  NAND2_X2 _f_permutation__U1612  ( .A1(SYNOPSYS_UNCONNECTED_937), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2515 ) );
  NAND2_X2 _f_permutation__U1611  ( .A1(_f_permutation__n2514 ), .A2(
        _f_permutation__n2515 ), .ZN(_f_permutation__n5236 ) );
  NAND2_X2 _f_permutation__U1610  ( .A1(_f_permutation__round_out[150]), .A2(
        _f_permutation__n7161 ), .ZN(_f_permutation__n2512 ) );
  NAND2_X2 _f_permutation__U1609  ( .A1(SYNOPSYS_UNCONNECTED_938), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2513 ) );
  NAND2_X2 _f_permutation__U1608  ( .A1(_f_permutation__n2512 ), .A2(
        _f_permutation__n2513 ), .ZN(_f_permutation__n5237 ) );
  NAND2_X2 _f_permutation__U1607  ( .A1(_f_permutation__round_out[149]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n2510 ) );
  NAND2_X2 _f_permutation__U1606  ( .A1(SYNOPSYS_UNCONNECTED_939), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2511 ) );
  NAND2_X2 _f_permutation__U1605  ( .A1(_f_permutation__n2510 ), .A2(
        _f_permutation__n2511 ), .ZN(_f_permutation__n5238 ) );
  NAND2_X2 _f_permutation__U1604  ( .A1(_f_permutation__round_out[148]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2508 ) );
  NAND2_X2 _f_permutation__U1603  ( .A1(SYNOPSYS_UNCONNECTED_940), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2509 ) );
  NAND2_X2 _f_permutation__U1602  ( .A1(_f_permutation__n2508 ), .A2(
        _f_permutation__n2509 ), .ZN(_f_permutation__n5239 ) );
  NAND2_X2 _f_permutation__U1601  ( .A1(_f_permutation__round_out[147]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2506 ) );
  NAND2_X2 _f_permutation__U1600  ( .A1(SYNOPSYS_UNCONNECTED_941), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2507 ) );
  NAND2_X2 _f_permutation__U1599  ( .A1(_f_permutation__n2506 ), .A2(
        _f_permutation__n2507 ), .ZN(_f_permutation__n5240 ) );
  NAND2_X2 _f_permutation__U1598  ( .A1(_f_permutation__round_out[146]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2504 ) );
  NAND2_X2 _f_permutation__U1597  ( .A1(SYNOPSYS_UNCONNECTED_942), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2505 ) );
  NAND2_X2 _f_permutation__U1596  ( .A1(_f_permutation__n2504 ), .A2(
        _f_permutation__n2505 ), .ZN(_f_permutation__n5241 ) );
  NAND2_X2 _f_permutation__U1595  ( .A1(_f_permutation__round_out[145]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2502 ) );
  NAND2_X2 _f_permutation__U1594  ( .A1(SYNOPSYS_UNCONNECTED_943), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2503 ) );
  NAND2_X2 _f_permutation__U1593  ( .A1(_f_permutation__n2502 ), .A2(
        _f_permutation__n2503 ), .ZN(_f_permutation__n5242 ) );
  NAND2_X2 _f_permutation__U1592  ( .A1(_f_permutation__round_out[144]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2500 ) );
  NAND2_X2 _f_permutation__U1591  ( .A1(SYNOPSYS_UNCONNECTED_944), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2501 ) );
  NAND2_X2 _f_permutation__U1590  ( .A1(_f_permutation__n2500 ), .A2(
        _f_permutation__n2501 ), .ZN(_f_permutation__n5243 ) );
  NAND2_X2 _f_permutation__U1589  ( .A1(_f_permutation__round_out[143]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2498 ) );
  NAND2_X2 _f_permutation__U1588  ( .A1(SYNOPSYS_UNCONNECTED_945), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2499 ) );
  NAND2_X2 _f_permutation__U1587  ( .A1(_f_permutation__n2498 ), .A2(
        _f_permutation__n2499 ), .ZN(_f_permutation__n5244 ) );
  NAND2_X2 _f_permutation__U1586  ( .A1(_f_permutation__round_out[142]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2496 ) );
  NAND2_X2 _f_permutation__U1585  ( .A1(SYNOPSYS_UNCONNECTED_946), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2497 ) );
  NAND2_X2 _f_permutation__U1584  ( .A1(_f_permutation__n2496 ), .A2(
        _f_permutation__n2497 ), .ZN(_f_permutation__n5245 ) );
  NAND2_X2 _f_permutation__U1583  ( .A1(_f_permutation__round_out[141]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2494 ) );
  NAND2_X2 _f_permutation__U1582  ( .A1(SYNOPSYS_UNCONNECTED_947), .A2(
        _f_permutation__n7293 ), .ZN(_f_permutation__n2495 ) );
  NAND2_X2 _f_permutation__U1581  ( .A1(_f_permutation__n2494 ), .A2(
        _f_permutation__n2495 ), .ZN(_f_permutation__n5246 ) );
  NAND2_X2 _f_permutation__U1580  ( .A1(_f_permutation__round_out[140]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2492 ) );
  NAND2_X2 _f_permutation__U1579  ( .A1(SYNOPSYS_UNCONNECTED_948), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2493 ) );
  NAND2_X2 _f_permutation__U1578  ( .A1(_f_permutation__n2492 ), .A2(
        _f_permutation__n2493 ), .ZN(_f_permutation__n5247 ) );
  NAND2_X2 _f_permutation__U1577  ( .A1(_f_permutation__round_out[139]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2490 ) );
  NAND2_X2 _f_permutation__U1576  ( .A1(SYNOPSYS_UNCONNECTED_949), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2491 ) );
  NAND2_X2 _f_permutation__U1575  ( .A1(_f_permutation__n2490 ), .A2(
        _f_permutation__n2491 ), .ZN(_f_permutation__n5248 ) );
  NAND2_X2 _f_permutation__U1574  ( .A1(_f_permutation__round_out[138]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2488 ) );
  NAND2_X2 _f_permutation__U1573  ( .A1(SYNOPSYS_UNCONNECTED_950), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2489 ) );
  NAND2_X2 _f_permutation__U1572  ( .A1(_f_permutation__n2488 ), .A2(
        _f_permutation__n2489 ), .ZN(_f_permutation__n5249 ) );
  NAND2_X2 _f_permutation__U1571  ( .A1(_f_permutation__round_out[137]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2486 ) );
  NAND2_X2 _f_permutation__U1570  ( .A1(SYNOPSYS_UNCONNECTED_951), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2487 ) );
  NAND2_X2 _f_permutation__U1569  ( .A1(_f_permutation__n2486 ), .A2(
        _f_permutation__n2487 ), .ZN(_f_permutation__n5250 ) );
  NAND2_X2 _f_permutation__U1568  ( .A1(_f_permutation__round_out[136]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2484 ) );
  NAND2_X2 _f_permutation__U1567  ( .A1(SYNOPSYS_UNCONNECTED_952), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2485 ) );
  NAND2_X2 _f_permutation__U1566  ( .A1(_f_permutation__n2484 ), .A2(
        _f_permutation__n2485 ), .ZN(_f_permutation__n5251 ) );
  NAND2_X2 _f_permutation__U1565  ( .A1(_f_permutation__round_out[135]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2482 ) );
  NAND2_X2 _f_permutation__U1564  ( .A1(SYNOPSYS_UNCONNECTED_953), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2483 ) );
  NAND2_X2 _f_permutation__U1563  ( .A1(_f_permutation__n2482 ), .A2(
        _f_permutation__n2483 ), .ZN(_f_permutation__n5252 ) );
  NAND2_X2 _f_permutation__U1562  ( .A1(_f_permutation__round_out[134]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2480 ) );
  NAND2_X2 _f_permutation__U1561  ( .A1(SYNOPSYS_UNCONNECTED_954), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2481 ) );
  NAND2_X2 _f_permutation__U1560  ( .A1(_f_permutation__n2480 ), .A2(
        _f_permutation__n2481 ), .ZN(_f_permutation__n5253 ) );
  NAND2_X2 _f_permutation__U1559  ( .A1(_f_permutation__round_out[133]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2478 ) );
  NAND2_X2 _f_permutation__U1558  ( .A1(SYNOPSYS_UNCONNECTED_955), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2479 ) );
  NAND2_X2 _f_permutation__U1557  ( .A1(_f_permutation__n2478 ), .A2(
        _f_permutation__n2479 ), .ZN(_f_permutation__n5254 ) );
  NAND2_X2 _f_permutation__U1556  ( .A1(_f_permutation__round_out[132]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2476 ) );
  NAND2_X2 _f_permutation__U1555  ( .A1(SYNOPSYS_UNCONNECTED_956), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2477 ) );
  NAND2_X2 _f_permutation__U1554  ( .A1(_f_permutation__n2476 ), .A2(
        _f_permutation__n2477 ), .ZN(_f_permutation__n5255 ) );
  NAND2_X2 _f_permutation__U1553  ( .A1(_f_permutation__round_out[131]), .A2(
        _f_permutation__n7085 ), .ZN(_f_permutation__n2474 ) );
  NAND2_X2 _f_permutation__U1552  ( .A1(SYNOPSYS_UNCONNECTED_957), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2475 ) );
  NAND2_X2 _f_permutation__U1551  ( .A1(_f_permutation__n2474 ), .A2(
        _f_permutation__n2475 ), .ZN(_f_permutation__n5256 ) );
  NAND2_X2 _f_permutation__U1550  ( .A1(_f_permutation__round_out[130]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n2472 ) );
  NAND2_X2 _f_permutation__U1549  ( .A1(SYNOPSYS_UNCONNECTED_958), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2473 ) );
  NAND2_X2 _f_permutation__U1548  ( .A1(_f_permutation__n2472 ), .A2(
        _f_permutation__n2473 ), .ZN(_f_permutation__n5257 ) );
  NAND2_X2 _f_permutation__U1547  ( .A1(_f_permutation__round_out[129]), .A2(
        _f_permutation__n7146 ), .ZN(_f_permutation__n2470 ) );
  NAND2_X2 _f_permutation__U1546  ( .A1(SYNOPSYS_UNCONNECTED_959), .A2(
        _f_permutation__n7294 ), .ZN(_f_permutation__n2471 ) );
  NAND2_X2 _f_permutation__U1545  ( .A1(_f_permutation__n2470 ), .A2(
        _f_permutation__n2471 ), .ZN(_f_permutation__n5258 ) );
  NAND2_X2 _f_permutation__U1544  ( .A1(_f_permutation__round_out[128]), .A2(
        _f_permutation__n7145 ), .ZN(_f_permutation__n2468 ) );
  NAND2_X2 _f_permutation__U1543  ( .A1(SYNOPSYS_UNCONNECTED_960), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2469 ) );
  NAND2_X2 _f_permutation__U1542  ( .A1(_f_permutation__n2468 ), .A2(
        _f_permutation__n2469 ), .ZN(_f_permutation__n5259 ) );
  NAND2_X2 _f_permutation__U1541  ( .A1(_f_permutation__round_out[127]), .A2(
        _f_permutation__n7144 ), .ZN(_f_permutation__n2466 ) );
  NAND2_X2 _f_permutation__U1540  ( .A1(SYNOPSYS_UNCONNECTED_961), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2467 ) );
  NAND2_X2 _f_permutation__U1539  ( .A1(_f_permutation__n2466 ), .A2(
        _f_permutation__n2467 ), .ZN(_f_permutation__n5260 ) );
  NAND2_X2 _f_permutation__U1538  ( .A1(_f_permutation__round_out[126]), .A2(
        _f_permutation__n7143 ), .ZN(_f_permutation__n2464 ) );
  NAND2_X2 _f_permutation__U1537  ( .A1(SYNOPSYS_UNCONNECTED_962), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2465 ) );
  NAND2_X2 _f_permutation__U1536  ( .A1(_f_permutation__n2464 ), .A2(
        _f_permutation__n2465 ), .ZN(_f_permutation__n5261 ) );
  NAND2_X2 _f_permutation__U1535  ( .A1(_f_permutation__round_out[125]), .A2(
        _f_permutation__n7163 ), .ZN(_f_permutation__n2462 ) );
  NAND2_X2 _f_permutation__U1534  ( .A1(SYNOPSYS_UNCONNECTED_963), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2463 ) );
  NAND2_X2 _f_permutation__U1533  ( .A1(_f_permutation__n2462 ), .A2(
        _f_permutation__n2463 ), .ZN(_f_permutation__n5262 ) );
  NAND2_X2 _f_permutation__U1532  ( .A1(_f_permutation__round_out[124]), .A2(
        _f_permutation__n7162 ), .ZN(_f_permutation__n2460 ) );
  NAND2_X2 _f_permutation__U1531  ( .A1(SYNOPSYS_UNCONNECTED_964), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2461 ) );
  NAND2_X2 _f_permutation__U1530  ( .A1(_f_permutation__n2460 ), .A2(
        _f_permutation__n2461 ), .ZN(_f_permutation__n5263 ) );
  NAND2_X2 _f_permutation__U1529  ( .A1(_f_permutation__round_out[123]), .A2(
        _f_permutation__n7167 ), .ZN(_f_permutation__n2458 ) );
  NAND2_X2 _f_permutation__U1528  ( .A1(SYNOPSYS_UNCONNECTED_965), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2459 ) );
  NAND2_X2 _f_permutation__U1527  ( .A1(_f_permutation__n2458 ), .A2(
        _f_permutation__n2459 ), .ZN(_f_permutation__n5264 ) );
  NAND2_X2 _f_permutation__U1526  ( .A1(_f_permutation__round_out[122]), .A2(
        _f_permutation__n7166 ), .ZN(_f_permutation__n2456 ) );
  NAND2_X2 _f_permutation__U1525  ( .A1(SYNOPSYS_UNCONNECTED_966), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2457 ) );
  NAND2_X2 _f_permutation__U1524  ( .A1(_f_permutation__n2456 ), .A2(
        _f_permutation__n2457 ), .ZN(_f_permutation__n5265 ) );
  NAND2_X2 _f_permutation__U1523  ( .A1(_f_permutation__round_out[121]), .A2(
        _f_permutation__n7156 ), .ZN(_f_permutation__n2454 ) );
  NAND2_X2 _f_permutation__U1522  ( .A1(SYNOPSYS_UNCONNECTED_967), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2455 ) );
  NAND2_X2 _f_permutation__U1521  ( .A1(_f_permutation__n2454 ), .A2(
        _f_permutation__n2455 ), .ZN(_f_permutation__n5266 ) );
  NAND2_X2 _f_permutation__U1520  ( .A1(_f_permutation__round_out[120]), .A2(
        _f_permutation__n7141 ), .ZN(_f_permutation__n2452 ) );
  NAND2_X2 _f_permutation__U1519  ( .A1(SYNOPSYS_UNCONNECTED_968), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2453 ) );
  NAND2_X2 _f_permutation__U1518  ( .A1(_f_permutation__n2452 ), .A2(
        _f_permutation__n2453 ), .ZN(_f_permutation__n5267 ) );
  NAND2_X2 _f_permutation__U1517  ( .A1(_f_permutation__round_out[119]), .A2(
        _f_permutation__n7140 ), .ZN(_f_permutation__n2450 ) );
  NAND2_X2 _f_permutation__U1516  ( .A1(SYNOPSYS_UNCONNECTED_969), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2451 ) );
  NAND2_X2 _f_permutation__U1515  ( .A1(_f_permutation__n2450 ), .A2(
        _f_permutation__n2451 ), .ZN(_f_permutation__n5268 ) );
  NAND2_X2 _f_permutation__U1514  ( .A1(_f_permutation__round_out[118]), .A2(
        _f_permutation__n7139 ), .ZN(_f_permutation__n2448 ) );
  NAND2_X2 _f_permutation__U1513  ( .A1(SYNOPSYS_UNCONNECTED_970), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2449 ) );
  NAND2_X2 _f_permutation__U1512  ( .A1(_f_permutation__n2448 ), .A2(
        _f_permutation__n2449 ), .ZN(_f_permutation__n5269 ) );
  NAND2_X2 _f_permutation__U1511  ( .A1(_f_permutation__round_out[117]), .A2(
        _f_permutation__n7142 ), .ZN(_f_permutation__n2446 ) );
  NAND2_X2 _f_permutation__U1510  ( .A1(SYNOPSYS_UNCONNECTED_971), .A2(
        _f_permutation__n7295 ), .ZN(_f_permutation__n2447 ) );
  NAND2_X2 _f_permutation__U1509  ( .A1(_f_permutation__n2446 ), .A2(
        _f_permutation__n2447 ), .ZN(_f_permutation__n5270 ) );
  NAND2_X2 _f_permutation__U1508  ( .A1(_f_permutation__round_out[116]), .A2(
        _f_permutation__n7164 ), .ZN(_f_permutation__n2444 ) );
  NAND2_X2 _f_permutation__U1507  ( .A1(SYNOPSYS_UNCONNECTED_972), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2445 ) );
  NAND2_X2 _f_permutation__U1506  ( .A1(_f_permutation__n2444 ), .A2(
        _f_permutation__n2445 ), .ZN(_f_permutation__n5271 ) );
  NAND2_X2 _f_permutation__U1505  ( .A1(_f_permutation__round_out[115]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n2442 ) );
  NAND2_X2 _f_permutation__U1504  ( .A1(SYNOPSYS_UNCONNECTED_973), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2443 ) );
  NAND2_X2 _f_permutation__U1503  ( .A1(_f_permutation__n2442 ), .A2(
        _f_permutation__n2443 ), .ZN(_f_permutation__n5272 ) );
  NAND2_X2 _f_permutation__U1502  ( .A1(_f_permutation__round_out[114]), .A2(
        _f_permutation__n7154 ), .ZN(_f_permutation__n2440 ) );
  NAND2_X2 _f_permutation__U1501  ( .A1(SYNOPSYS_UNCONNECTED_974), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2441 ) );
  NAND2_X2 _f_permutation__U1500  ( .A1(_f_permutation__n2440 ), .A2(
        _f_permutation__n2441 ), .ZN(_f_permutation__n5273 ) );
  NAND2_X2 _f_permutation__U1499  ( .A1(_f_permutation__round_out[113]), .A2(
        _f_permutation__n7161 ), .ZN(_f_permutation__n2438 ) );
  NAND2_X2 _f_permutation__U1498  ( .A1(SYNOPSYS_UNCONNECTED_975), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2439 ) );
  NAND2_X2 _f_permutation__U1497  ( .A1(_f_permutation__n2438 ), .A2(
        _f_permutation__n2439 ), .ZN(_f_permutation__n5274 ) );
  NAND2_X2 _f_permutation__U1496  ( .A1(_f_permutation__round_out[112]), .A2(
        _f_permutation__n7161 ), .ZN(_f_permutation__n2436 ) );
  NAND2_X2 _f_permutation__U1495  ( .A1(SYNOPSYS_UNCONNECTED_976), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2437 ) );
  NAND2_X2 _f_permutation__U1494  ( .A1(_f_permutation__n2436 ), .A2(
        _f_permutation__n2437 ), .ZN(_f_permutation__n5275 ) );
  NAND2_X2 _f_permutation__U1493  ( .A1(_f_permutation__round_out[111]), .A2(
        _f_permutation__n7162 ), .ZN(_f_permutation__n2434 ) );
  NAND2_X2 _f_permutation__U1492  ( .A1(SYNOPSYS_UNCONNECTED_977), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2435 ) );
  NAND2_X2 _f_permutation__U1491  ( .A1(_f_permutation__n2434 ), .A2(
        _f_permutation__n2435 ), .ZN(_f_permutation__n5276 ) );
  NAND2_X2 _f_permutation__U1490  ( .A1(_f_permutation__round_out[110]), .A2(
        _f_permutation__n7167 ), .ZN(_f_permutation__n2432 ) );
  NAND2_X2 _f_permutation__U1489  ( .A1(SYNOPSYS_UNCONNECTED_978), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2433 ) );
  NAND2_X2 _f_permutation__U1488  ( .A1(_f_permutation__n2432 ), .A2(
        _f_permutation__n2433 ), .ZN(_f_permutation__n5277 ) );
  NAND2_X2 _f_permutation__U1487  ( .A1(_f_permutation__round_out[109]), .A2(
        _f_permutation__n7166 ), .ZN(_f_permutation__n2430 ) );
  NAND2_X2 _f_permutation__U1486  ( .A1(SYNOPSYS_UNCONNECTED_979), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2431 ) );
  NAND2_X2 _f_permutation__U1485  ( .A1(_f_permutation__n2430 ), .A2(
        _f_permutation__n2431 ), .ZN(_f_permutation__n5278 ) );
  NAND2_X2 _f_permutation__U1484  ( .A1(_f_permutation__round_out[108]), .A2(
        _f_permutation__n7165 ), .ZN(_f_permutation__n2428 ) );
  NAND2_X2 _f_permutation__U1483  ( .A1(SYNOPSYS_UNCONNECTED_980), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2429 ) );
  NAND2_X2 _f_permutation__U1482  ( .A1(_f_permutation__n2428 ), .A2(
        _f_permutation__n2429 ), .ZN(_f_permutation__n5279 ) );
  NAND2_X2 _f_permutation__U1481  ( .A1(_f_permutation__round_out[107]), .A2(
        _f_permutation__n7164 ), .ZN(_f_permutation__n2426 ) );
  NAND2_X2 _f_permutation__U1480  ( .A1(SYNOPSYS_UNCONNECTED_981), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2427 ) );
  NAND2_X2 _f_permutation__U1479  ( .A1(_f_permutation__n2426 ), .A2(
        _f_permutation__n2427 ), .ZN(_f_permutation__n5280 ) );
  NAND2_X2 _f_permutation__U1478  ( .A1(_f_permutation__round_out[106]), .A2(
        _f_permutation__n7156 ), .ZN(_f_permutation__n2424 ) );
  NAND2_X2 _f_permutation__U1477  ( .A1(SYNOPSYS_UNCONNECTED_982), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2425 ) );
  NAND2_X2 _f_permutation__U1476  ( .A1(_f_permutation__n2424 ), .A2(
        _f_permutation__n2425 ), .ZN(_f_permutation__n5281 ) );
  NAND2_X2 _f_permutation__U1475  ( .A1(_f_permutation__round_out[105]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n2422 ) );
  NAND2_X2 _f_permutation__U1474  ( .A1(SYNOPSYS_UNCONNECTED_983), .A2(
        _f_permutation__n7296 ), .ZN(_f_permutation__n2423 ) );
  NAND2_X2 _f_permutation__U1473  ( .A1(_f_permutation__n2422 ), .A2(
        _f_permutation__n2423 ), .ZN(_f_permutation__n5282 ) );
  NAND2_X2 _f_permutation__U1472  ( .A1(_f_permutation__round_out[104]), .A2(
        _f_permutation__n7154 ), .ZN(_f_permutation__n2420 ) );
  NAND2_X2 _f_permutation__U1471  ( .A1(SYNOPSYS_UNCONNECTED_984), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2421 ) );
  NAND2_X2 _f_permutation__U1470  ( .A1(_f_permutation__n2420 ), .A2(
        _f_permutation__n2421 ), .ZN(_f_permutation__n5283 ) );
  NAND2_X2 _f_permutation__U1469  ( .A1(_f_permutation__round_out[103]), .A2(
        _f_permutation__n7141 ), .ZN(_f_permutation__n2418 ) );
  NAND2_X2 _f_permutation__U1468  ( .A1(SYNOPSYS_UNCONNECTED_985), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2419 ) );
  NAND2_X2 _f_permutation__U1467  ( .A1(_f_permutation__n2418 ), .A2(
        _f_permutation__n2419 ), .ZN(_f_permutation__n5284 ) );
  NAND2_X2 _f_permutation__U1466  ( .A1(_f_permutation__round_out[102]), .A2(
        _f_permutation__n7140 ), .ZN(_f_permutation__n2416 ) );
  NAND2_X2 _f_permutation__U1465  ( .A1(SYNOPSYS_UNCONNECTED_986), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2417 ) );
  NAND2_X2 _f_permutation__U1464  ( .A1(_f_permutation__n2416 ), .A2(
        _f_permutation__n2417 ), .ZN(_f_permutation__n5285 ) );
  NAND2_X2 _f_permutation__U1463  ( .A1(_f_permutation__round_out[101]), .A2(
        _f_permutation__n7154 ), .ZN(_f_permutation__n2414 ) );
  NAND2_X2 _f_permutation__U1462  ( .A1(SYNOPSYS_UNCONNECTED_987), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2415 ) );
  NAND2_X2 _f_permutation__U1461  ( .A1(_f_permutation__n2414 ), .A2(
        _f_permutation__n2415 ), .ZN(_f_permutation__n5286 ) );
  NAND2_X2 _f_permutation__U1460  ( .A1(_f_permutation__round_out[100]), .A2(
        _f_permutation__n7139 ), .ZN(_f_permutation__n2412 ) );
  NAND2_X2 _f_permutation__U1459  ( .A1(SYNOPSYS_UNCONNECTED_988), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2413 ) );
  NAND2_X2 _f_permutation__U1458  ( .A1(_f_permutation__n2412 ), .A2(
        _f_permutation__n2413 ), .ZN(_f_permutation__n5287 ) );
  NAND2_X2 _f_permutation__U1457  ( .A1(_f_permutation__round_out[99]), .A2(
        _f_permutation__n7146 ), .ZN(_f_permutation__n2410 ) );
  NAND2_X2 _f_permutation__U1456  ( .A1(SYNOPSYS_UNCONNECTED_989), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2411 ) );
  NAND2_X2 _f_permutation__U1455  ( .A1(_f_permutation__n2410 ), .A2(
        _f_permutation__n2411 ), .ZN(_f_permutation__n5288 ) );
  NAND2_X2 _f_permutation__U1454  ( .A1(_f_permutation__round_out[98]), .A2(
        _f_permutation__n7145 ), .ZN(_f_permutation__n2408 ) );
  NAND2_X2 _f_permutation__U1453  ( .A1(SYNOPSYS_UNCONNECTED_990), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2409 ) );
  NAND2_X2 _f_permutation__U1452  ( .A1(_f_permutation__n2408 ), .A2(
        _f_permutation__n2409 ), .ZN(_f_permutation__n5289 ) );
  NAND2_X2 _f_permutation__U1451  ( .A1(_f_permutation__round_out[97]), .A2(
        _f_permutation__n7144 ), .ZN(_f_permutation__n2406 ) );
  NAND2_X2 _f_permutation__U1450  ( .A1(SYNOPSYS_UNCONNECTED_991), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2407 ) );
  NAND2_X2 _f_permutation__U1449  ( .A1(_f_permutation__n2406 ), .A2(
        _f_permutation__n2407 ), .ZN(_f_permutation__n5290 ) );
  NAND2_X2 _f_permutation__U1448  ( .A1(_f_permutation__round_out[96]), .A2(
        _f_permutation__n7143 ), .ZN(_f_permutation__n2404 ) );
  NAND2_X2 _f_permutation__U1447  ( .A1(SYNOPSYS_UNCONNECTED_992), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2405 ) );
  NAND2_X2 _f_permutation__U1446  ( .A1(_f_permutation__n2404 ), .A2(
        _f_permutation__n2405 ), .ZN(_f_permutation__n5291 ) );
  NAND2_X2 _f_permutation__U1445  ( .A1(_f_permutation__round_out[95]), .A2(
        _f_permutation__n7142 ), .ZN(_f_permutation__n2402 ) );
  NAND2_X2 _f_permutation__U1444  ( .A1(SYNOPSYS_UNCONNECTED_993), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2403 ) );
  NAND2_X2 _f_permutation__U1443  ( .A1(_f_permutation__n2402 ), .A2(
        _f_permutation__n2403 ), .ZN(_f_permutation__n5292 ) );
  NAND2_X2 _f_permutation__U1442  ( .A1(_f_permutation__round_out[94]), .A2(
        _f_permutation__n7163 ), .ZN(_f_permutation__n2400 ) );
  NAND2_X2 _f_permutation__U1441  ( .A1(SYNOPSYS_UNCONNECTED_994), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2401 ) );
  NAND2_X2 _f_permutation__U1440  ( .A1(_f_permutation__n2400 ), .A2(
        _f_permutation__n2401 ), .ZN(_f_permutation__n5293 ) );
  NAND2_X2 _f_permutation__U1439  ( .A1(_f_permutation__round_out[93]), .A2(
        _f_permutation__n7162 ), .ZN(_f_permutation__n2398 ) );
  NAND2_X2 _f_permutation__U1438  ( .A1(SYNOPSYS_UNCONNECTED_995), .A2(
        _f_permutation__n7297 ), .ZN(_f_permutation__n2399 ) );
  NAND2_X2 _f_permutation__U1437  ( .A1(_f_permutation__n2398 ), .A2(
        _f_permutation__n2399 ), .ZN(_f_permutation__n5294 ) );
  NAND2_X2 _f_permutation__U1436  ( .A1(_f_permutation__round_out[92]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n2396 ) );
  NAND2_X2 _f_permutation__U1435  ( .A1(SYNOPSYS_UNCONNECTED_996), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2397 ) );
  NAND2_X2 _f_permutation__U1434  ( .A1(_f_permutation__n2396 ), .A2(
        _f_permutation__n2397 ), .ZN(_f_permutation__n5295 ) );
  NAND2_X2 _f_permutation__U1433  ( .A1(_f_permutation__round_out[91]), .A2(
        _f_permutation__n7165 ), .ZN(_f_permutation__n2394 ) );
  NAND2_X2 _f_permutation__U1432  ( .A1(SYNOPSYS_UNCONNECTED_997), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2395 ) );
  NAND2_X2 _f_permutation__U1431  ( .A1(_f_permutation__n2394 ), .A2(
        _f_permutation__n2395 ), .ZN(_f_permutation__n5296 ) );
  NAND2_X2 _f_permutation__U1430  ( .A1(_f_permutation__round_out[90]), .A2(
        _f_permutation__n7154 ), .ZN(_f_permutation__n2392 ) );
  NAND2_X2 _f_permutation__U1429  ( .A1(SYNOPSYS_UNCONNECTED_998), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2393 ) );
  NAND2_X2 _f_permutation__U1428  ( .A1(_f_permutation__n2392 ), .A2(
        _f_permutation__n2393 ), .ZN(_f_permutation__n5297 ) );
  NAND2_X2 _f_permutation__U1427  ( .A1(_f_permutation__round_out[89]), .A2(
        _f_permutation__n7161 ), .ZN(_f_permutation__n2390 ) );
  NAND2_X2 _f_permutation__U1426  ( .A1(SYNOPSYS_UNCONNECTED_999), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2391 ) );
  NAND2_X2 _f_permutation__U1425  ( .A1(_f_permutation__n2390 ), .A2(
        _f_permutation__n2391 ), .ZN(_f_permutation__n5298 ) );
  NAND2_X2 _f_permutation__U1424  ( .A1(_f_permutation__round_out[88]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n2388 ) );
  NAND2_X2 _f_permutation__U1423  ( .A1(SYNOPSYS_UNCONNECTED_1000), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2389 ) );
  NAND2_X2 _f_permutation__U1422  ( .A1(_f_permutation__n2388 ), .A2(
        _f_permutation__n2389 ), .ZN(_f_permutation__n5299 ) );
  NAND2_X2 _f_permutation__U1421  ( .A1(_f_permutation__round_out[87]), .A2(
        _f_permutation__n7164 ), .ZN(_f_permutation__n2386 ) );
  NAND2_X2 _f_permutation__U1420  ( .A1(SYNOPSYS_UNCONNECTED_1001), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2387 ) );
  NAND2_X2 _f_permutation__U1419  ( .A1(_f_permutation__n2386 ), .A2(
        _f_permutation__n2387 ), .ZN(_f_permutation__n5300 ) );
  NAND2_X2 _f_permutation__U1418  ( .A1(_f_permutation__round_out[86]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n2384 ) );
  NAND2_X2 _f_permutation__U1417  ( .A1(SYNOPSYS_UNCONNECTED_1002), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2385 ) );
  NAND2_X2 _f_permutation__U1416  ( .A1(_f_permutation__n2384 ), .A2(
        _f_permutation__n2385 ), .ZN(_f_permutation__n5301 ) );
  NAND2_X2 _f_permutation__U1415  ( .A1(_f_permutation__round_out[85]), .A2(
        _f_permutation__n7153 ), .ZN(_f_permutation__n2382 ) );
  NAND2_X2 _f_permutation__U1414  ( .A1(SYNOPSYS_UNCONNECTED_1003), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2383 ) );
  NAND2_X2 _f_permutation__U1413  ( .A1(_f_permutation__n2382 ), .A2(
        _f_permutation__n2383 ), .ZN(_f_permutation__n5302 ) );
  NAND2_X2 _f_permutation__U1412  ( .A1(_f_permutation__round_out[84]), .A2(
        _f_permutation__n7165 ), .ZN(_f_permutation__n2380 ) );
  NAND2_X2 _f_permutation__U1411  ( .A1(SYNOPSYS_UNCONNECTED_1004), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2381 ) );
  NAND2_X2 _f_permutation__U1410  ( .A1(_f_permutation__n2380 ), .A2(
        _f_permutation__n2381 ), .ZN(_f_permutation__n5303 ) );
  NAND2_X2 _f_permutation__U1409  ( .A1(_f_permutation__round_out[83]), .A2(
        _f_permutation__n7168 ), .ZN(_f_permutation__n2378 ) );
  NAND2_X2 _f_permutation__U1408  ( .A1(SYNOPSYS_UNCONNECTED_1005), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2379 ) );
  NAND2_X2 _f_permutation__U1407  ( .A1(_f_permutation__n2378 ), .A2(
        _f_permutation__n2379 ), .ZN(_f_permutation__n5304 ) );
  NAND2_X2 _f_permutation__U1406  ( .A1(_f_permutation__round_out[82]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n2376 ) );
  NAND2_X2 _f_permutation__U1405  ( .A1(SYNOPSYS_UNCONNECTED_1006), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2377 ) );
  NAND2_X2 _f_permutation__U1404  ( .A1(_f_permutation__n2376 ), .A2(
        _f_permutation__n2377 ), .ZN(_f_permutation__n5305 ) );
  NAND2_X2 _f_permutation__U1403  ( .A1(_f_permutation__round_out[81]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n2374 ) );
  NAND2_X2 _f_permutation__U1402  ( .A1(SYNOPSYS_UNCONNECTED_1007), .A2(
        _f_permutation__n7298 ), .ZN(_f_permutation__n2375 ) );
  NAND2_X2 _f_permutation__U1401  ( .A1(_f_permutation__n2374 ), .A2(
        _f_permutation__n2375 ), .ZN(_f_permutation__n5306 ) );
  NAND2_X2 _f_permutation__U1400  ( .A1(_f_permutation__round_out[80]), .A2(
        _f_permutation__n7149 ), .ZN(_f_permutation__n2372 ) );
  NAND2_X2 _f_permutation__U1399  ( .A1(SYNOPSYS_UNCONNECTED_1008), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2373 ) );
  NAND2_X2 _f_permutation__U1398  ( .A1(_f_permutation__n2372 ), .A2(
        _f_permutation__n2373 ), .ZN(_f_permutation__n5307 ) );
  NAND2_X2 _f_permutation__U1397  ( .A1(_f_permutation__round_out[79]), .A2(
        _f_permutation__n7148 ), .ZN(_f_permutation__n2370 ) );
  NAND2_X2 _f_permutation__U1396  ( .A1(SYNOPSYS_UNCONNECTED_1009), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2371 ) );
  NAND2_X2 _f_permutation__U1395  ( .A1(_f_permutation__n2370 ), .A2(
        _f_permutation__n2371 ), .ZN(_f_permutation__n5308 ) );
  NAND2_X2 _f_permutation__U1394  ( .A1(_f_permutation__round_out[78]), .A2(
        _f_permutation__n7147 ), .ZN(_f_permutation__n2368 ) );
  NAND2_X2 _f_permutation__U1393  ( .A1(SYNOPSYS_UNCONNECTED_1010), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2369 ) );
  NAND2_X2 _f_permutation__U1392  ( .A1(_f_permutation__n2368 ), .A2(
        _f_permutation__n2369 ), .ZN(_f_permutation__n5309 ) );
  NAND2_X2 _f_permutation__U1391  ( .A1(_f_permutation__round_out[77]), .A2(
        _f_permutation__n7152 ), .ZN(_f_permutation__n2366 ) );
  NAND2_X2 _f_permutation__U1390  ( .A1(SYNOPSYS_UNCONNECTED_1011), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2367 ) );
  NAND2_X2 _f_permutation__U1389  ( .A1(_f_permutation__n2366 ), .A2(
        _f_permutation__n2367 ), .ZN(_f_permutation__n5310 ) );
  NAND2_X2 _f_permutation__U1388  ( .A1(_f_permutation__round_out[76]), .A2(
        _f_permutation__n7151 ), .ZN(_f_permutation__n2364 ) );
  NAND2_X2 _f_permutation__U1387  ( .A1(SYNOPSYS_UNCONNECTED_1012), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2365 ) );
  NAND2_X2 _f_permutation__U1386  ( .A1(_f_permutation__n2364 ), .A2(
        _f_permutation__n2365 ), .ZN(_f_permutation__n5311 ) );
  NAND2_X2 _f_permutation__U1385  ( .A1(_f_permutation__round_out[75]), .A2(
        _f_permutation__n7150 ), .ZN(_f_permutation__n2362 ) );
  NAND2_X2 _f_permutation__U1384  ( .A1(SYNOPSYS_UNCONNECTED_1013), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2363 ) );
  NAND2_X2 _f_permutation__U1383  ( .A1(_f_permutation__n2362 ), .A2(
        _f_permutation__n2363 ), .ZN(_f_permutation__n5312 ) );
  NAND2_X2 _f_permutation__U1382  ( .A1(_f_permutation__round_out[74]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2360 ) );
  NAND2_X2 _f_permutation__U1381  ( .A1(SYNOPSYS_UNCONNECTED_1014), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2361 ) );
  NAND2_X2 _f_permutation__U1380  ( .A1(_f_permutation__n2360 ), .A2(
        _f_permutation__n2361 ), .ZN(_f_permutation__n5313 ) );
  NAND2_X2 _f_permutation__U1379  ( .A1(_f_permutation__round_out[73]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2358 ) );
  NAND2_X2 _f_permutation__U1378  ( .A1(SYNOPSYS_UNCONNECTED_1015), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2359 ) );
  NAND2_X2 _f_permutation__U1377  ( .A1(_f_permutation__n2358 ), .A2(
        _f_permutation__n2359 ), .ZN(_f_permutation__n5314 ) );
  NAND2_X2 _f_permutation__U1376  ( .A1(_f_permutation__round_out[72]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2356 ) );
  NAND2_X2 _f_permutation__U1375  ( .A1(SYNOPSYS_UNCONNECTED_1016), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2357 ) );
  NAND2_X2 _f_permutation__U1374  ( .A1(_f_permutation__n2356 ), .A2(
        _f_permutation__n2357 ), .ZN(_f_permutation__n5315 ) );
  NAND2_X2 _f_permutation__U1373  ( .A1(_f_permutation__round_out[71]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2354 ) );
  NAND2_X2 _f_permutation__U1372  ( .A1(SYNOPSYS_UNCONNECTED_1017), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2355 ) );
  NAND2_X2 _f_permutation__U1371  ( .A1(_f_permutation__n2354 ), .A2(
        _f_permutation__n2355 ), .ZN(_f_permutation__n5316 ) );
  NAND2_X2 _f_permutation__U1370  ( .A1(_f_permutation__round_out[70]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2352 ) );
  NAND2_X2 _f_permutation__U1369  ( .A1(SYNOPSYS_UNCONNECTED_1018), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2353 ) );
  NAND2_X2 _f_permutation__U1368  ( .A1(_f_permutation__n2352 ), .A2(
        _f_permutation__n2353 ), .ZN(_f_permutation__n5317 ) );
  NAND2_X2 _f_permutation__U1367  ( .A1(_f_permutation__round_out[69]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2350 ) );
  NAND2_X2 _f_permutation__U1366  ( .A1(SYNOPSYS_UNCONNECTED_1019), .A2(
        _f_permutation__n7299 ), .ZN(_f_permutation__n2351 ) );
  NAND2_X2 _f_permutation__U1365  ( .A1(_f_permutation__n2350 ), .A2(
        _f_permutation__n2351 ), .ZN(_f_permutation__n5318 ) );
  NAND2_X2 _f_permutation__U1364  ( .A1(_f_permutation__round_out[68]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2348 ) );
  NAND2_X2 _f_permutation__U1363  ( .A1(SYNOPSYS_UNCONNECTED_1020), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2349 ) );
  NAND2_X2 _f_permutation__U1362  ( .A1(_f_permutation__n2348 ), .A2(
        _f_permutation__n2349 ), .ZN(_f_permutation__n5319 ) );
  NAND2_X2 _f_permutation__U1361  ( .A1(_f_permutation__round_out[67]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2346 ) );
  NAND2_X2 _f_permutation__U1360  ( .A1(SYNOPSYS_UNCONNECTED_1021), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2347 ) );
  NAND2_X2 _f_permutation__U1359  ( .A1(_f_permutation__n2346 ), .A2(
        _f_permutation__n2347 ), .ZN(_f_permutation__n5320 ) );
  NAND2_X2 _f_permutation__U1358  ( .A1(_f_permutation__round_out[66]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2344 ) );
  NAND2_X2 _f_permutation__U1357  ( .A1(SYNOPSYS_UNCONNECTED_1022), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2345 ) );
  NAND2_X2 _f_permutation__U1356  ( .A1(_f_permutation__n2344 ), .A2(
        _f_permutation__n2345 ), .ZN(_f_permutation__n5321 ) );
  NAND2_X2 _f_permutation__U1355  ( .A1(_f_permutation__round_out[65]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2342 ) );
  NAND2_X2 _f_permutation__U1354  ( .A1(SYNOPSYS_UNCONNECTED_1023), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2343 ) );
  NAND2_X2 _f_permutation__U1353  ( .A1(_f_permutation__n2342 ), .A2(
        _f_permutation__n2343 ), .ZN(_f_permutation__n5322 ) );
  NAND2_X2 _f_permutation__U1352  ( .A1(_f_permutation__round_out[64]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2340 ) );
  NAND2_X2 _f_permutation__U1351  ( .A1(SYNOPSYS_UNCONNECTED_1024), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2341 ) );
  NAND2_X2 _f_permutation__U1350  ( .A1(_f_permutation__n2340 ), .A2(
        _f_permutation__n2341 ), .ZN(_f_permutation__n5323 ) );
  NAND2_X2 _f_permutation__U1349  ( .A1(_f_permutation__round_out[63]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2338 ) );
  NAND2_X2 _f_permutation__U1348  ( .A1(SYNOPSYS_UNCONNECTED_1025), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2339 ) );
  NAND2_X2 _f_permutation__U1347  ( .A1(_f_permutation__n2338 ), .A2(
        _f_permutation__n2339 ), .ZN(_f_permutation__n5324 ) );
  NAND2_X2 _f_permutation__U1346  ( .A1(_f_permutation__round_out[62]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2336 ) );
  NAND2_X2 _f_permutation__U1345  ( .A1(SYNOPSYS_UNCONNECTED_1026), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2337 ) );
  NAND2_X2 _f_permutation__U1344  ( .A1(_f_permutation__n2336 ), .A2(
        _f_permutation__n2337 ), .ZN(_f_permutation__n5325 ) );
  NAND2_X2 _f_permutation__U1343  ( .A1(_f_permutation__round_out[61]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2334 ) );
  NAND2_X2 _f_permutation__U1342  ( .A1(SYNOPSYS_UNCONNECTED_1027), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2335 ) );
  NAND2_X2 _f_permutation__U1341  ( .A1(_f_permutation__n2334 ), .A2(
        _f_permutation__n2335 ), .ZN(_f_permutation__n5326 ) );
  NAND2_X2 _f_permutation__U1340  ( .A1(_f_permutation__round_out[60]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2332 ) );
  NAND2_X2 _f_permutation__U1339  ( .A1(SYNOPSYS_UNCONNECTED_1028), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2333 ) );
  NAND2_X2 _f_permutation__U1338  ( .A1(_f_permutation__n2332 ), .A2(
        _f_permutation__n2333 ), .ZN(_f_permutation__n5327 ) );
  NAND2_X2 _f_permutation__U1337  ( .A1(_f_permutation__round_out[59]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2330 ) );
  NAND2_X2 _f_permutation__U1336  ( .A1(SYNOPSYS_UNCONNECTED_1029), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2331 ) );
  NAND2_X2 _f_permutation__U1335  ( .A1(_f_permutation__n2330 ), .A2(
        _f_permutation__n2331 ), .ZN(_f_permutation__n5328 ) );
  NAND2_X2 _f_permutation__U1334  ( .A1(_f_permutation__round_out[58]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2328 ) );
  NAND2_X2 _f_permutation__U1333  ( .A1(SYNOPSYS_UNCONNECTED_1030), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2329 ) );
  NAND2_X2 _f_permutation__U1332  ( .A1(_f_permutation__n2328 ), .A2(
        _f_permutation__n2329 ), .ZN(_f_permutation__n5329 ) );
  NAND2_X2 _f_permutation__U1331  ( .A1(_f_permutation__round_out[57]), .A2(
        _f_permutation__n7087 ), .ZN(_f_permutation__n2326 ) );
  NAND2_X2 _f_permutation__U1330  ( .A1(SYNOPSYS_UNCONNECTED_1031), .A2(
        _f_permutation__n7300 ), .ZN(_f_permutation__n2327 ) );
  NAND2_X2 _f_permutation__U1329  ( .A1(_f_permutation__n2326 ), .A2(
        _f_permutation__n2327 ), .ZN(_f_permutation__n5330 ) );
  NAND2_X2 _f_permutation__U1328  ( .A1(_f_permutation__round_out[56]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n2324 ) );
  NAND2_X2 _f_permutation__U1327  ( .A1(SYNOPSYS_UNCONNECTED_1032), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2325 ) );
  NAND2_X2 _f_permutation__U1326  ( .A1(_f_permutation__n2324 ), .A2(
        _f_permutation__n2325 ), .ZN(_f_permutation__n5331 ) );
  NAND2_X2 _f_permutation__U1325  ( .A1(_f_permutation__round_out[55]), .A2(
        _f_permutation__n7167 ), .ZN(_f_permutation__n2322 ) );
  NAND2_X2 _f_permutation__U1324  ( .A1(SYNOPSYS_UNCONNECTED_1033), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2323 ) );
  NAND2_X2 _f_permutation__U1323  ( .A1(_f_permutation__n2322 ), .A2(
        _f_permutation__n2323 ), .ZN(_f_permutation__n5332 ) );
  NAND2_X2 _f_permutation__U1322  ( .A1(_f_permutation__round_out[54]), .A2(
        _f_permutation__n7166 ), .ZN(_f_permutation__n2320 ) );
  NAND2_X2 _f_permutation__U1321  ( .A1(SYNOPSYS_UNCONNECTED_1034), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2321 ) );
  NAND2_X2 _f_permutation__U1320  ( .A1(_f_permutation__n2320 ), .A2(
        _f_permutation__n2321 ), .ZN(_f_permutation__n5333 ) );
  NAND2_X2 _f_permutation__U1319  ( .A1(_f_permutation__round_out[53]), .A2(
        _f_permutation__n7165 ), .ZN(_f_permutation__n2318 ) );
  NAND2_X2 _f_permutation__U1318  ( .A1(SYNOPSYS_UNCONNECTED_1035), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2319 ) );
  NAND2_X2 _f_permutation__U1317  ( .A1(_f_permutation__n2318 ), .A2(
        _f_permutation__n2319 ), .ZN(_f_permutation__n5334 ) );
  NAND2_X2 _f_permutation__U1316  ( .A1(_f_permutation__round_out[52]), .A2(
        _f_permutation__n7164 ), .ZN(_f_permutation__n2316 ) );
  NAND2_X2 _f_permutation__U1315  ( .A1(SYNOPSYS_UNCONNECTED_1036), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2317 ) );
  NAND2_X2 _f_permutation__U1314  ( .A1(_f_permutation__n2316 ), .A2(
        _f_permutation__n2317 ), .ZN(_f_permutation__n5335 ) );
  NAND2_X2 _f_permutation__U1313  ( .A1(_f_permutation__round_out[51]), .A2(
        _f_permutation__n7155 ), .ZN(_f_permutation__n2314 ) );
  NAND2_X2 _f_permutation__U1312  ( .A1(SYNOPSYS_UNCONNECTED_1037), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2315 ) );
  NAND2_X2 _f_permutation__U1311  ( .A1(_f_permutation__n2314 ), .A2(
        _f_permutation__n2315 ), .ZN(_f_permutation__n5336 ) );
  NAND2_X2 _f_permutation__U1310  ( .A1(_f_permutation__round_out[50]), .A2(
        _f_permutation__n7154 ), .ZN(_f_permutation__n2312 ) );
  NAND2_X2 _f_permutation__U1309  ( .A1(SYNOPSYS_UNCONNECTED_1038), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2313 ) );
  NAND2_X2 _f_permutation__U1308  ( .A1(_f_permutation__n2312 ), .A2(
        _f_permutation__n2313 ), .ZN(_f_permutation__n5337 ) );
  NAND2_X2 _f_permutation__U1307  ( .A1(_f_permutation__round_out[49]), .A2(
        _f_permutation__n7161 ), .ZN(_f_permutation__n2310 ) );
  NAND2_X2 _f_permutation__U1306  ( .A1(SYNOPSYS_UNCONNECTED_1039), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2311 ) );
  NAND2_X2 _f_permutation__U1305  ( .A1(_f_permutation__n2310 ), .A2(
        _f_permutation__n2311 ), .ZN(_f_permutation__n5338 ) );
  NAND2_X2 _f_permutation__U1304  ( .A1(_f_permutation__round_out[48]), .A2(
        _f_permutation__n7160 ), .ZN(_f_permutation__n2308 ) );
  NAND2_X2 _f_permutation__U1303  ( .A1(SYNOPSYS_UNCONNECTED_1040), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2309 ) );
  NAND2_X2 _f_permutation__U1302  ( .A1(_f_permutation__n2308 ), .A2(
        _f_permutation__n2309 ), .ZN(_f_permutation__n5339 ) );
  NAND2_X2 _f_permutation__U1301  ( .A1(_f_permutation__round_out[47]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n2306 ) );
  NAND2_X2 _f_permutation__U1300  ( .A1(SYNOPSYS_UNCONNECTED_1041), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2307 ) );
  NAND2_X2 _f_permutation__U1299  ( .A1(_f_permutation__n2306 ), .A2(
        _f_permutation__n2307 ), .ZN(_f_permutation__n5340 ) );
  NAND2_X2 _f_permutation__U1298  ( .A1(_f_permutation__round_out[46]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n2304 ) );
  NAND2_X2 _f_permutation__U1297  ( .A1(SYNOPSYS_UNCONNECTED_1042), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2305 ) );
  NAND2_X2 _f_permutation__U1296  ( .A1(_f_permutation__n2304 ), .A2(
        _f_permutation__n2305 ), .ZN(_f_permutation__n5341 ) );
  NAND2_X2 _f_permutation__U1295  ( .A1(_f_permutation__round_out[45]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n2302 ) );
  NAND2_X2 _f_permutation__U1294  ( .A1(SYNOPSYS_UNCONNECTED_1043), .A2(
        _f_permutation__n7301 ), .ZN(_f_permutation__n2303 ) );
  NAND2_X2 _f_permutation__U1293  ( .A1(_f_permutation__n2302 ), .A2(
        _f_permutation__n2303 ), .ZN(_f_permutation__n5342 ) );
  NAND2_X2 _f_permutation__U1292  ( .A1(_f_permutation__round_out[44]), .A2(
        _f_permutation__n7168 ), .ZN(_f_permutation__n2300 ) );
  NAND2_X2 _f_permutation__U1291  ( .A1(SYNOPSYS_UNCONNECTED_1044), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2301 ) );
  NAND2_X2 _f_permutation__U1290  ( .A1(_f_permutation__n2300 ), .A2(
        _f_permutation__n2301 ), .ZN(_f_permutation__n5343 ) );
  NAND2_X2 _f_permutation__U1289  ( .A1(_f_permutation__round_out[43]), .A2(
        _f_permutation__n7167 ), .ZN(_f_permutation__n2298 ) );
  NAND2_X2 _f_permutation__U1288  ( .A1(SYNOPSYS_UNCONNECTED_1045), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2299 ) );
  NAND2_X2 _f_permutation__U1287  ( .A1(_f_permutation__n2298 ), .A2(
        _f_permutation__n2299 ), .ZN(_f_permutation__n5344 ) );
  NAND2_X2 _f_permutation__U1286  ( .A1(_f_permutation__round_out[42]), .A2(
        _f_permutation__n7166 ), .ZN(_f_permutation__n2296 ) );
  NAND2_X2 _f_permutation__U1285  ( .A1(SYNOPSYS_UNCONNECTED_1046), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2297 ) );
  NAND2_X2 _f_permutation__U1284  ( .A1(_f_permutation__n2296 ), .A2(
        _f_permutation__n2297 ), .ZN(_f_permutation__n5345 ) );
  NAND2_X2 _f_permutation__U1283  ( .A1(_f_permutation__round_out[41]), .A2(
        _f_permutation__n7165 ), .ZN(_f_permutation__n2294 ) );
  NAND2_X2 _f_permutation__U1282  ( .A1(SYNOPSYS_UNCONNECTED_1047), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2295 ) );
  NAND2_X2 _f_permutation__U1281  ( .A1(_f_permutation__n2294 ), .A2(
        _f_permutation__n2295 ), .ZN(_f_permutation__n5346 ) );
  NAND2_X2 _f_permutation__U1280  ( .A1(_f_permutation__round_out[40]), .A2(
        _f_permutation__n7164 ), .ZN(_f_permutation__n2292 ) );
  NAND2_X2 _f_permutation__U1279  ( .A1(SYNOPSYS_UNCONNECTED_1048), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2293 ) );
  NAND2_X2 _f_permutation__U1278  ( .A1(_f_permutation__n2292 ), .A2(
        _f_permutation__n2293 ), .ZN(_f_permutation__n5347 ) );
  NAND2_X2 _f_permutation__U1277  ( .A1(_f_permutation__round_out[39]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n2290 ) );
  NAND2_X2 _f_permutation__U1276  ( .A1(SYNOPSYS_UNCONNECTED_1049), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2291 ) );
  NAND2_X2 _f_permutation__U1275  ( .A1(_f_permutation__n2290 ), .A2(
        _f_permutation__n2291 ), .ZN(_f_permutation__n5348 ) );
  NAND2_X2 _f_permutation__U1274  ( .A1(_f_permutation__round_out[38]), .A2(
        _f_permutation__n7153 ), .ZN(_f_permutation__n2288 ) );
  NAND2_X2 _f_permutation__U1273  ( .A1(SYNOPSYS_UNCONNECTED_1050), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2289 ) );
  NAND2_X2 _f_permutation__U1272  ( .A1(_f_permutation__n2288 ), .A2(
        _f_permutation__n2289 ), .ZN(_f_permutation__n5349 ) );
  NAND2_X2 _f_permutation__U1271  ( .A1(_f_permutation__round_out[37]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n2286 ) );
  NAND2_X2 _f_permutation__U1270  ( .A1(SYNOPSYS_UNCONNECTED_1051), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2287 ) );
  NAND2_X2 _f_permutation__U1269  ( .A1(_f_permutation__n2286 ), .A2(
        _f_permutation__n2287 ), .ZN(_f_permutation__n5350 ) );
  NAND2_X2 _f_permutation__U1268  ( .A1(_f_permutation__round_out[36]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n2284 ) );
  NAND2_X2 _f_permutation__U1267  ( .A1(SYNOPSYS_UNCONNECTED_1052), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2285 ) );
  NAND2_X2 _f_permutation__U1266  ( .A1(_f_permutation__n2284 ), .A2(
        _f_permutation__n2285 ), .ZN(_f_permutation__n5351 ) );
  NAND2_X2 _f_permutation__U1265  ( .A1(_f_permutation__round_out[35]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n2282 ) );
  NAND2_X2 _f_permutation__U1264  ( .A1(SYNOPSYS_UNCONNECTED_1053), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2283 ) );
  NAND2_X2 _f_permutation__U1263  ( .A1(_f_permutation__n2282 ), .A2(
        _f_permutation__n2283 ), .ZN(_f_permutation__n5352 ) );
  NAND2_X2 _f_permutation__U1262  ( .A1(_f_permutation__round_out[34]), .A2(
        _f_permutation__n7168 ), .ZN(_f_permutation__n2280 ) );
  NAND2_X2 _f_permutation__U1261  ( .A1(SYNOPSYS_UNCONNECTED_1054), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2281 ) );
  NAND2_X2 _f_permutation__U1260  ( .A1(_f_permutation__n2280 ), .A2(
        _f_permutation__n2281 ), .ZN(_f_permutation__n5353 ) );
  NAND2_X2 _f_permutation__U1259  ( .A1(_f_permutation__round_out[33]), .A2(
        _f_permutation__n7153 ), .ZN(_f_permutation__n2278 ) );
  NAND2_X2 _f_permutation__U1258  ( .A1(SYNOPSYS_UNCONNECTED_1055), .A2(
        _f_permutation__n7302 ), .ZN(_f_permutation__n2279 ) );
  NAND2_X2 _f_permutation__U1257  ( .A1(_f_permutation__n2278 ), .A2(
        _f_permutation__n2279 ), .ZN(_f_permutation__n5354 ) );
  NAND2_X2 _f_permutation__U1256  ( .A1(_f_permutation__round_out[32]), .A2(
        _f_permutation__n7149 ), .ZN(_f_permutation__n2276 ) );
  NAND2_X2 _f_permutation__U1255  ( .A1(SYNOPSYS_UNCONNECTED_1056), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2277 ) );
  NAND2_X2 _f_permutation__U1254  ( .A1(_f_permutation__n2276 ), .A2(
        _f_permutation__n2277 ), .ZN(_f_permutation__n5355 ) );
  NAND2_X2 _f_permutation__U1253  ( .A1(_f_permutation__round_out[31]), .A2(
        _f_permutation__n7148 ), .ZN(_f_permutation__n2274 ) );
  NAND2_X2 _f_permutation__U1252  ( .A1(SYNOPSYS_UNCONNECTED_1057), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2275 ) );
  NAND2_X2 _f_permutation__U1251  ( .A1(_f_permutation__n2274 ), .A2(
        _f_permutation__n2275 ), .ZN(_f_permutation__n5356 ) );
  NAND2_X2 _f_permutation__U1250  ( .A1(_f_permutation__round_out[30]), .A2(
        _f_permutation__n7147 ), .ZN(_f_permutation__n2272 ) );
  NAND2_X2 _f_permutation__U1249  ( .A1(SYNOPSYS_UNCONNECTED_1058), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2273 ) );
  NAND2_X2 _f_permutation__U1248  ( .A1(_f_permutation__n2272 ), .A2(
        _f_permutation__n2273 ), .ZN(_f_permutation__n5357 ) );
  NAND2_X2 _f_permutation__U1247  ( .A1(_f_permutation__round_out[29]), .A2(
        _f_permutation__n7152 ), .ZN(_f_permutation__n2270 ) );
  NAND2_X2 _f_permutation__U1246  ( .A1(SYNOPSYS_UNCONNECTED_1059), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2271 ) );
  NAND2_X2 _f_permutation__U1245  ( .A1(_f_permutation__n2270 ), .A2(
        _f_permutation__n2271 ), .ZN(_f_permutation__n5358 ) );
  NAND2_X2 _f_permutation__U1244  ( .A1(_f_permutation__round_out[28]), .A2(
        _f_permutation__n7151 ), .ZN(_f_permutation__n2268 ) );
  NAND2_X2 _f_permutation__U1243  ( .A1(SYNOPSYS_UNCONNECTED_1060), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2269 ) );
  NAND2_X2 _f_permutation__U1242  ( .A1(_f_permutation__n2268 ), .A2(
        _f_permutation__n2269 ), .ZN(_f_permutation__n5359 ) );
  NAND2_X2 _f_permutation__U1241  ( .A1(_f_permutation__round_out[27]), .A2(
        _f_permutation__n7150 ), .ZN(_f_permutation__n2266 ) );
  NAND2_X2 _f_permutation__U1240  ( .A1(SYNOPSYS_UNCONNECTED_1061), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2267 ) );
  NAND2_X2 _f_permutation__U1239  ( .A1(_f_permutation__n2266 ), .A2(
        _f_permutation__n2267 ), .ZN(_f_permutation__n5360 ) );
  NAND2_X2 _f_permutation__U1238  ( .A1(_f_permutation__round_out[26]), .A2(
        _f_permutation__n7146 ), .ZN(_f_permutation__n2264 ) );
  NAND2_X2 _f_permutation__U1237  ( .A1(SYNOPSYS_UNCONNECTED_1062), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2265 ) );
  NAND2_X2 _f_permutation__U1236  ( .A1(_f_permutation__n2264 ), .A2(
        _f_permutation__n2265 ), .ZN(_f_permutation__n5361 ) );
  NAND2_X2 _f_permutation__U1235  ( .A1(_f_permutation__round_out[25]), .A2(
        _f_permutation__n7145 ), .ZN(_f_permutation__n2262 ) );
  NAND2_X2 _f_permutation__U1234  ( .A1(SYNOPSYS_UNCONNECTED_1063), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2263 ) );
  NAND2_X2 _f_permutation__U1233  ( .A1(_f_permutation__n2262 ), .A2(
        _f_permutation__n2263 ), .ZN(_f_permutation__n5362 ) );
  NAND2_X2 _f_permutation__U1232  ( .A1(_f_permutation__round_out[24]), .A2(
        _f_permutation__n7144 ), .ZN(_f_permutation__n2260 ) );
  NAND2_X2 _f_permutation__U1231  ( .A1(SYNOPSYS_UNCONNECTED_1064), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2261 ) );
  NAND2_X2 _f_permutation__U1230  ( .A1(_f_permutation__n2260 ), .A2(
        _f_permutation__n2261 ), .ZN(_f_permutation__n5363 ) );
  NAND2_X2 _f_permutation__U1229  ( .A1(_f_permutation__round_out[23]), .A2(
        _f_permutation__n7143 ), .ZN(_f_permutation__n2258 ) );
  NAND2_X2 _f_permutation__U1228  ( .A1(SYNOPSYS_UNCONNECTED_1065), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2259 ) );
  NAND2_X2 _f_permutation__U1227  ( .A1(_f_permutation__n2258 ), .A2(
        _f_permutation__n2259 ), .ZN(_f_permutation__n5364 ) );
  NAND2_X2 _f_permutation__U1226  ( .A1(_f_permutation__round_out[22]), .A2(
        _f_permutation__n7163 ), .ZN(_f_permutation__n2256 ) );
  NAND2_X2 _f_permutation__U1225  ( .A1(SYNOPSYS_UNCONNECTED_1066), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2257 ) );
  NAND2_X2 _f_permutation__U1224  ( .A1(_f_permutation__n2256 ), .A2(
        _f_permutation__n2257 ), .ZN(_f_permutation__n5365 ) );
  NAND2_X2 _f_permutation__U1223  ( .A1(_f_permutation__round_out[21]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n2254 ) );
  NAND2_X2 _f_permutation__U1222  ( .A1(SYNOPSYS_UNCONNECTED_1067), .A2(
        _f_permutation__n7303 ), .ZN(_f_permutation__n2255 ) );
  NAND2_X2 _f_permutation__U1221  ( .A1(_f_permutation__n2254 ), .A2(
        _f_permutation__n2255 ), .ZN(_f_permutation__n5366 ) );
  NAND2_X2 _f_permutation__U1220  ( .A1(_f_permutation__round_out[20]), .A2(
        _f_permutation__n7141 ), .ZN(_f_permutation__n2252 ) );
  NAND2_X2 _f_permutation__U1219  ( .A1(SYNOPSYS_UNCONNECTED_1068), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2253 ) );
  NAND2_X2 _f_permutation__U1218  ( .A1(_f_permutation__n2252 ), .A2(
        _f_permutation__n2253 ), .ZN(_f_permutation__n5367 ) );
  NAND2_X2 _f_permutation__U1217  ( .A1(_f_permutation__round_out[19]), .A2(
        _f_permutation__n7140 ), .ZN(_f_permutation__n2250 ) );
  NAND2_X2 _f_permutation__U1216  ( .A1(SYNOPSYS_UNCONNECTED_1069), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2251 ) );
  NAND2_X2 _f_permutation__U1215  ( .A1(_f_permutation__n2250 ), .A2(
        _f_permutation__n2251 ), .ZN(_f_permutation__n5368 ) );
  NAND2_X2 _f_permutation__U1214  ( .A1(_f_permutation__round_out[18]), .A2(
        _f_permutation__n7139 ), .ZN(_f_permutation__n2248 ) );
  NAND2_X2 _f_permutation__U1213  ( .A1(SYNOPSYS_UNCONNECTED_1070), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2249 ) );
  NAND2_X2 _f_permutation__U1212  ( .A1(_f_permutation__n2248 ), .A2(
        _f_permutation__n2249 ), .ZN(_f_permutation__n5369 ) );
  NAND2_X2 _f_permutation__U1211  ( .A1(_f_permutation__round_out[17]), .A2(
        _f_permutation__n7142 ), .ZN(_f_permutation__n2246 ) );
  NAND2_X2 _f_permutation__U1210  ( .A1(SYNOPSYS_UNCONNECTED_1071), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2247 ) );
  NAND2_X2 _f_permutation__U1209  ( .A1(_f_permutation__n2246 ), .A2(
        _f_permutation__n2247 ), .ZN(_f_permutation__n5370 ) );
  NAND2_X2 _f_permutation__U1208  ( .A1(_f_permutation__round_out[16]), .A2(
        _f_permutation__n7158 ), .ZN(_f_permutation__n2244 ) );
  NAND2_X2 _f_permutation__U1207  ( .A1(SYNOPSYS_UNCONNECTED_1072), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2245 ) );
  NAND2_X2 _f_permutation__U1206  ( .A1(_f_permutation__n2244 ), .A2(
        _f_permutation__n2245 ), .ZN(_f_permutation__n5371 ) );
  NAND2_X2 _f_permutation__U1205  ( .A1(_f_permutation__round_out[15]), .A2(
        _f_permutation__n7157 ), .ZN(_f_permutation__n2242 ) );
  NAND2_X2 _f_permutation__U1204  ( .A1(SYNOPSYS_UNCONNECTED_1073), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2243 ) );
  NAND2_X2 _f_permutation__U1203  ( .A1(_f_permutation__n2242 ), .A2(
        _f_permutation__n2243 ), .ZN(_f_permutation__n5372 ) );
  NAND2_X2 _f_permutation__U1202  ( .A1(_f_permutation__round_out[14]), .A2(
        _f_permutation__n7153 ), .ZN(_f_permutation__n2240 ) );
  NAND2_X2 _f_permutation__U1201  ( .A1(SYNOPSYS_UNCONNECTED_1074), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2241 ) );
  NAND2_X2 _f_permutation__U1200  ( .A1(_f_permutation__n2240 ), .A2(
        _f_permutation__n2241 ), .ZN(_f_permutation__n5373 ) );
  NAND2_X2 _f_permutation__U1199  ( .A1(_f_permutation__round_out[13]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n2238 ) );
  NAND2_X2 _f_permutation__U1198  ( .A1(SYNOPSYS_UNCONNECTED_1075), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2239 ) );
  NAND2_X2 _f_permutation__U1197  ( .A1(_f_permutation__n2238 ), .A2(
        _f_permutation__n2239 ), .ZN(_f_permutation__n5374 ) );
  NAND2_X2 _f_permutation__U1196  ( .A1(_f_permutation__round_out[12]), .A2(
        _f_permutation__n7168 ), .ZN(_f_permutation__n2236 ) );
  NAND2_X2 _f_permutation__U1195  ( .A1(SYNOPSYS_UNCONNECTED_1076), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2237 ) );
  NAND2_X2 _f_permutation__U1194  ( .A1(_f_permutation__n2236 ), .A2(
        _f_permutation__n2237 ), .ZN(_f_permutation__n5375 ) );
  NAND2_X2 _f_permutation__U1193  ( .A1(_f_permutation__round_out[11]), .A2(
        _f_permutation__n7141 ), .ZN(_f_permutation__n2234 ) );
  NAND2_X2 _f_permutation__U1192  ( .A1(SYNOPSYS_UNCONNECTED_1077), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2235 ) );
  NAND2_X2 _f_permutation__U1191  ( .A1(_f_permutation__n2234 ), .A2(
        _f_permutation__n2235 ), .ZN(_f_permutation__n5376 ) );
  NAND2_X2 _f_permutation__U1190  ( .A1(_f_permutation__round_out[10]), .A2(
        _f_permutation__n7140 ), .ZN(_f_permutation__n2232 ) );
  NAND2_X2 _f_permutation__U1189  ( .A1(SYNOPSYS_UNCONNECTED_1078), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2233 ) );
  NAND2_X2 _f_permutation__U1188  ( .A1(_f_permutation__n2232 ), .A2(
        _f_permutation__n2233 ), .ZN(_f_permutation__n5377 ) );
  NAND2_X2 _f_permutation__U1187  ( .A1(_f_permutation__round_out[9]), .A2(
        _f_permutation__n7139 ), .ZN(_f_permutation__n2230 ) );
  NAND2_X2 _f_permutation__U1186  ( .A1(SYNOPSYS_UNCONNECTED_1079), .A2(
        _f_permutation__n7304 ), .ZN(_f_permutation__n2231 ) );
  NAND2_X2 _f_permutation__U1185  ( .A1(_f_permutation__n2230 ), .A2(
        _f_permutation__n2231 ), .ZN(_f_permutation__n5378 ) );
  NAND2_X2 _f_permutation__U1184  ( .A1(_f_permutation__round_out[8]), .A2(
        _f_permutation__n7142 ), .ZN(_f_permutation__n2228 ) );
  NAND2_X2 _f_permutation__U1183  ( .A1(SYNOPSYS_UNCONNECTED_1080), .A2(
        _f_permutation__n7220 ), .ZN(_f_permutation__n2229 ) );
  NAND2_X2 _f_permutation__U1182  ( .A1(_f_permutation__n2228 ), .A2(
        _f_permutation__n2229 ), .ZN(_f_permutation__n5379 ) );
  NAND2_X2 _f_permutation__U1181  ( .A1(_f_permutation__round_out[7]), .A2(
        _f_permutation__n7149 ), .ZN(_f_permutation__n2226 ) );
  NAND2_X2 _f_permutation__U1180  ( .A1(SYNOPSYS_UNCONNECTED_1081), .A2(
        _f_permutation__n7310 ), .ZN(_f_permutation__n2227 ) );
  NAND2_X2 _f_permutation__U1179  ( .A1(_f_permutation__n2226 ), .A2(
        _f_permutation__n2227 ), .ZN(_f_permutation__n5380 ) );
  NAND2_X2 _f_permutation__U1178  ( .A1(_f_permutation__round_out[6]), .A2(
        _f_permutation__n7148 ), .ZN(_f_permutation__n2224 ) );
  NAND2_X2 _f_permutation__U1177  ( .A1(SYNOPSYS_UNCONNECTED_1082), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n2225 ) );
  NAND2_X2 _f_permutation__U1176  ( .A1(_f_permutation__n2224 ), .A2(
        _f_permutation__n2225 ), .ZN(_f_permutation__n5381 ) );
  NAND2_X2 _f_permutation__U1175  ( .A1(_f_permutation__round_out[5]), .A2(
        _f_permutation__n7147 ), .ZN(_f_permutation__n2222 ) );
  NAND2_X2 _f_permutation__U1174  ( .A1(SYNOPSYS_UNCONNECTED_1083), .A2(
        _f_permutation__n7308 ), .ZN(_f_permutation__n2223 ) );
  NAND2_X2 _f_permutation__U1173  ( .A1(_f_permutation__n2222 ), .A2(
        _f_permutation__n2223 ), .ZN(_f_permutation__n5382 ) );
  NAND2_X2 _f_permutation__U1172  ( .A1(_f_permutation__round_out[4]), .A2(
        _f_permutation__n7152 ), .ZN(_f_permutation__n2220 ) );
  NAND2_X2 _f_permutation__U1171  ( .A1(SYNOPSYS_UNCONNECTED_1084), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2221 ) );
  NAND2_X2 _f_permutation__U1170  ( .A1(_f_permutation__n2220 ), .A2(
        _f_permutation__n2221 ), .ZN(_f_permutation__n5383 ) );
  NAND2_X2 _f_permutation__U1169  ( .A1(_f_permutation__round_out[3]), .A2(
        _f_permutation__n7159 ), .ZN(_f_permutation__n2218 ) );
  NAND2_X2 _f_permutation__U1168  ( .A1(SYNOPSYS_UNCONNECTED_1085), .A2(
        _f_permutation__n7257 ), .ZN(_f_permutation__n2219 ) );
  NAND2_X2 _f_permutation__U1167  ( .A1(_f_permutation__n2218 ), .A2(
        _f_permutation__n2219 ), .ZN(_f_permutation__n5384 ) );
  NAND2_X2 _f_permutation__U1166  ( .A1(_f_permutation__round_out[2]), .A2(
        _f_permutation__n7156 ), .ZN(_f_permutation__n2216 ) );
  NAND2_X2 _f_permutation__U1165  ( .A1(SYNOPSYS_UNCONNECTED_1086), .A2(
        _f_permutation__n7310 ), .ZN(_f_permutation__n2217 ) );
  NAND2_X2 _f_permutation__U1164  ( .A1(_f_permutation__n2216 ), .A2(
        _f_permutation__n2217 ), .ZN(_f_permutation__n5385 ) );
  NAND2_X2 _f_permutation__U1163  ( .A1(_f_permutation__round_out[1]), .A2(
        _f_permutation__n7141 ), .ZN(_f_permutation__n2214 ) );
  NAND2_X2 _f_permutation__U1162  ( .A1(SYNOPSYS_UNCONNECTED_1087), .A2(
        _f_permutation__n7310 ), .ZN(_f_permutation__n2215 ) );
  NAND2_X2 _f_permutation__U1161  ( .A1(_f_permutation__n2214 ), .A2(
        _f_permutation__n2215 ), .ZN(_f_permutation__n5386 ) );
  NAND2_X2 _f_permutation__U1160  ( .A1(_f_permutation__round_out[0]), .A2(
        _f_permutation__n7165 ), .ZN(_f_permutation__n2210 ) );
  NAND2_X2 _f_permutation__U1159  ( .A1(SYNOPSYS_UNCONNECTED_1088), .A2(
        _f_permutation__n7289 ), .ZN(_f_permutation__n2211 ) );
  NAND2_X2 _f_permutation__U1158  ( .A1(_f_permutation__n2210 ), .A2(
        _f_permutation__n2211 ), .ZN(_f_permutation__n5387 ) );
  NAND2_X2 _f_permutation__U1155  ( .A1(padder_out[0]), .A2(f_ack), .ZN(
        _f_permutation__n2207 ) );
  XNOR2_X2 _f_permutation__U1154  ( .A(SYNOPSYS_UNCONNECTED_64), .B(
        _f_permutation__n2207 ), .ZN(_f_permutation__round_in[1024]) );
  NAND2_X2 _f_permutation__U1153  ( .A1(padder_out[1]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2206 ) );
  XNOR2_X2 _f_permutation__U1152  ( .A(SYNOPSYS_UNCONNECTED_63), .B(
        _f_permutation__n2206 ), .ZN(_f_permutation__round_in[1025]) );
  NAND2_X2 _f_permutation__U1151  ( .A1(padder_out[2]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2205 ) );
  XNOR2_X2 _f_permutation__U1150  ( .A(SYNOPSYS_UNCONNECTED_62), .B(
        _f_permutation__n2205 ), .ZN(_f_permutation__round_in[1026]) );
  NAND2_X2 _f_permutation__U1149  ( .A1(padder_out[3]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2204 ) );
  XNOR2_X2 _f_permutation__U1148  ( .A(SYNOPSYS_UNCONNECTED_61), .B(
        _f_permutation__n2204 ), .ZN(_f_permutation__round_in[1027]) );
  NAND2_X2 _f_permutation__U1147  ( .A1(padder_out[4]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2203 ) );
  XNOR2_X2 _f_permutation__U1146  ( .A(SYNOPSYS_UNCONNECTED_60), .B(
        _f_permutation__n2203 ), .ZN(_f_permutation__round_in[1028]) );
  NAND2_X2 _f_permutation__U1145  ( .A1(padder_out[5]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2202 ) );
  XNOR2_X2 _f_permutation__U1144  ( .A(SYNOPSYS_UNCONNECTED_59), .B(
        _f_permutation__n2202 ), .ZN(_f_permutation__round_in[1029]) );
  NAND2_X2 _f_permutation__U1143  ( .A1(padder_out[6]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2201 ) );
  XNOR2_X2 _f_permutation__U1142  ( .A(SYNOPSYS_UNCONNECTED_58), .B(
        _f_permutation__n2201 ), .ZN(_f_permutation__round_in[1030]) );
  NAND2_X2 _f_permutation__U1141  ( .A1(padder_out[7]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2200 ) );
  XNOR2_X2 _f_permutation__U1140  ( .A(SYNOPSYS_UNCONNECTED_57), .B(
        _f_permutation__n2200 ), .ZN(_f_permutation__round_in[1031]) );
  NAND2_X2 _f_permutation__U1139  ( .A1(padder_out[8]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2199 ) );
  XNOR2_X2 _f_permutation__U1138  ( .A(SYNOPSYS_UNCONNECTED_56), .B(
        _f_permutation__n2199 ), .ZN(_f_permutation__round_in[1032]) );
  NAND2_X2 _f_permutation__U1137  ( .A1(padder_out[9]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2198 ) );
  XNOR2_X2 _f_permutation__U1136  ( .A(SYNOPSYS_UNCONNECTED_55), .B(
        _f_permutation__n2198 ), .ZN(_f_permutation__round_in[1033]) );
  NAND2_X2 _f_permutation__U1135  ( .A1(padder_out[10]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2197 ) );
  XNOR2_X2 _f_permutation__U1134  ( .A(SYNOPSYS_UNCONNECTED_54), .B(
        _f_permutation__n2197 ), .ZN(_f_permutation__round_in[1034]) );
  NAND2_X2 _f_permutation__U1133  ( .A1(padder_out[11]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2196 ) );
  XNOR2_X2 _f_permutation__U1132  ( .A(SYNOPSYS_UNCONNECTED_53), .B(
        _f_permutation__n2196 ), .ZN(_f_permutation__round_in[1035]) );
  NAND2_X2 _f_permutation__U1131  ( .A1(padder_out[12]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2195 ) );
  XNOR2_X2 _f_permutation__U1130  ( .A(SYNOPSYS_UNCONNECTED_52), .B(
        _f_permutation__n2195 ), .ZN(_f_permutation__round_in[1036]) );
  NAND2_X2 _f_permutation__U1129  ( .A1(padder_out[13]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2194 ) );
  XNOR2_X2 _f_permutation__U1128  ( .A(SYNOPSYS_UNCONNECTED_51), .B(
        _f_permutation__n2194 ), .ZN(_f_permutation__round_in[1037]) );
  NAND2_X2 _f_permutation__U1127  ( .A1(padder_out[14]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2193 ) );
  XNOR2_X2 _f_permutation__U1126  ( .A(SYNOPSYS_UNCONNECTED_50), .B(
        _f_permutation__n2193 ), .ZN(_f_permutation__round_in[1038]) );
  NAND2_X2 _f_permutation__U1125  ( .A1(padder_out[15]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2192 ) );
  XNOR2_X2 _f_permutation__U1124  ( .A(SYNOPSYS_UNCONNECTED_49), .B(
        _f_permutation__n2192 ), .ZN(_f_permutation__round_in[1039]) );
  NAND2_X2 _f_permutation__U1123  ( .A1(padder_out[16]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2191 ) );
  XNOR2_X2 _f_permutation__U1122  ( .A(SYNOPSYS_UNCONNECTED_48), .B(
        _f_permutation__n2191 ), .ZN(_f_permutation__round_in[1040]) );
  NAND2_X2 _f_permutation__U1121  ( .A1(padder_out[17]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2190 ) );
  XNOR2_X2 _f_permutation__U1120  ( .A(SYNOPSYS_UNCONNECTED_47), .B(
        _f_permutation__n2190 ), .ZN(_f_permutation__round_in[1041]) );
  NAND2_X2 _f_permutation__U1119  ( .A1(padder_out[18]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2189 ) );
  XNOR2_X2 _f_permutation__U1118  ( .A(SYNOPSYS_UNCONNECTED_46), .B(
        _f_permutation__n2189 ), .ZN(_f_permutation__round_in[1042]) );
  NAND2_X2 _f_permutation__U1117  ( .A1(padder_out[19]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2188 ) );
  XNOR2_X2 _f_permutation__U1116  ( .A(SYNOPSYS_UNCONNECTED_45), .B(
        _f_permutation__n2188 ), .ZN(_f_permutation__round_in[1043]) );
  NAND2_X2 _f_permutation__U1115  ( .A1(padder_out[20]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2187 ) );
  XNOR2_X2 _f_permutation__U1114  ( .A(SYNOPSYS_UNCONNECTED_44), .B(
        _f_permutation__n2187 ), .ZN(_f_permutation__round_in[1044]) );
  NAND2_X2 _f_permutation__U1113  ( .A1(padder_out[21]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2186 ) );
  XNOR2_X2 _f_permutation__U1112  ( .A(SYNOPSYS_UNCONNECTED_43), .B(
        _f_permutation__n2186 ), .ZN(_f_permutation__round_in[1045]) );
  NAND2_X2 _f_permutation__U1111  ( .A1(padder_out[22]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2185 ) );
  XNOR2_X2 _f_permutation__U1110  ( .A(SYNOPSYS_UNCONNECTED_42), .B(
        _f_permutation__n2185 ), .ZN(_f_permutation__round_in[1046]) );
  NAND2_X2 _f_permutation__U1109  ( .A1(padder_out[23]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2184 ) );
  XNOR2_X2 _f_permutation__U1108  ( .A(SYNOPSYS_UNCONNECTED_41), .B(
        _f_permutation__n2184 ), .ZN(_f_permutation__round_in[1047]) );
  NAND2_X2 _f_permutation__U1107  ( .A1(padder_out[24]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2183 ) );
  XNOR2_X2 _f_permutation__U1106  ( .A(SYNOPSYS_UNCONNECTED_40), .B(
        _f_permutation__n2183 ), .ZN(_f_permutation__round_in[1048]) );
  NAND2_X2 _f_permutation__U1105  ( .A1(padder_out[25]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2182 ) );
  XNOR2_X2 _f_permutation__U1104  ( .A(SYNOPSYS_UNCONNECTED_39), .B(
        _f_permutation__n2182 ), .ZN(_f_permutation__round_in[1049]) );
  NAND2_X2 _f_permutation__U1103  ( .A1(padder_out[26]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2181 ) );
  XNOR2_X2 _f_permutation__U1102  ( .A(SYNOPSYS_UNCONNECTED_38), .B(
        _f_permutation__n2181 ), .ZN(_f_permutation__round_in[1050]) );
  NAND2_X2 _f_permutation__U1101  ( .A1(padder_out[27]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2180 ) );
  XNOR2_X2 _f_permutation__U1100  ( .A(SYNOPSYS_UNCONNECTED_37), .B(
        _f_permutation__n2180 ), .ZN(_f_permutation__round_in[1051]) );
  NAND2_X2 _f_permutation__U1099  ( .A1(padder_out[28]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2179 ) );
  XNOR2_X2 _f_permutation__U1098  ( .A(SYNOPSYS_UNCONNECTED_36), .B(
        _f_permutation__n2179 ), .ZN(_f_permutation__round_in[1052]) );
  NAND2_X2 _f_permutation__U1097  ( .A1(padder_out[29]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2178 ) );
  XNOR2_X2 _f_permutation__U1096  ( .A(SYNOPSYS_UNCONNECTED_35), .B(
        _f_permutation__n2178 ), .ZN(_f_permutation__round_in[1053]) );
  NAND2_X2 _f_permutation__U1095  ( .A1(padder_out[30]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2177 ) );
  XNOR2_X2 _f_permutation__U1094  ( .A(SYNOPSYS_UNCONNECTED_34), .B(
        _f_permutation__n2177 ), .ZN(_f_permutation__round_in[1054]) );
  NAND2_X2 _f_permutation__U1093  ( .A1(padder_out[31]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2176 ) );
  XNOR2_X2 _f_permutation__U1092  ( .A(SYNOPSYS_UNCONNECTED_33), .B(
        _f_permutation__n2176 ), .ZN(_f_permutation__round_in[1055]) );
  NAND2_X2 _f_permutation__U1091  ( .A1(padder_out[32]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2175 ) );
  XNOR2_X2 _f_permutation__U1090  ( .A(SYNOPSYS_UNCONNECTED_32), .B(
        _f_permutation__n2175 ), .ZN(_f_permutation__round_in[1056]) );
  NAND2_X2 _f_permutation__U1089  ( .A1(padder_out[33]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2174 ) );
  XNOR2_X2 _f_permutation__U1088  ( .A(SYNOPSYS_UNCONNECTED_31), .B(
        _f_permutation__n2174 ), .ZN(_f_permutation__round_in[1057]) );
  NAND2_X2 _f_permutation__U1087  ( .A1(padder_out[34]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2173 ) );
  XNOR2_X2 _f_permutation__U1086  ( .A(SYNOPSYS_UNCONNECTED_30), .B(
        _f_permutation__n2173 ), .ZN(_f_permutation__round_in[1058]) );
  NAND2_X2 _f_permutation__U1085  ( .A1(padder_out[35]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2172 ) );
  XNOR2_X2 _f_permutation__U1084  ( .A(SYNOPSYS_UNCONNECTED_29), .B(
        _f_permutation__n2172 ), .ZN(_f_permutation__round_in[1059]) );
  NAND2_X2 _f_permutation__U1083  ( .A1(padder_out[36]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2171 ) );
  XNOR2_X2 _f_permutation__U1082  ( .A(SYNOPSYS_UNCONNECTED_28), .B(
        _f_permutation__n2171 ), .ZN(_f_permutation__round_in[1060]) );
  NAND2_X2 _f_permutation__U1081  ( .A1(padder_out[37]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n2170 ) );
  XNOR2_X2 _f_permutation__U1080  ( .A(SYNOPSYS_UNCONNECTED_27), .B(
        _f_permutation__n2170 ), .ZN(_f_permutation__round_in[1061]) );
  NAND2_X2 _f_permutation__U1079  ( .A1(padder_out[38]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2169 ) );
  XNOR2_X2 _f_permutation__U1078  ( .A(SYNOPSYS_UNCONNECTED_26), .B(
        _f_permutation__n2169 ), .ZN(_f_permutation__round_in[1062]) );
  NAND2_X2 _f_permutation__U1077  ( .A1(padder_out[39]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2168 ) );
  XNOR2_X2 _f_permutation__U1076  ( .A(SYNOPSYS_UNCONNECTED_25), .B(
        _f_permutation__n2168 ), .ZN(_f_permutation__round_in[1063]) );
  NAND2_X2 _f_permutation__U1075  ( .A1(padder_out[40]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2167 ) );
  XNOR2_X2 _f_permutation__U1074  ( .A(SYNOPSYS_UNCONNECTED_24), .B(
        _f_permutation__n2167 ), .ZN(_f_permutation__round_in[1064]) );
  NAND2_X2 _f_permutation__U1073  ( .A1(padder_out[41]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2166 ) );
  XNOR2_X2 _f_permutation__U1072  ( .A(SYNOPSYS_UNCONNECTED_23), .B(
        _f_permutation__n2166 ), .ZN(_f_permutation__round_in[1065]) );
  NAND2_X2 _f_permutation__U1071  ( .A1(padder_out[42]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2165 ) );
  XNOR2_X2 _f_permutation__U1070  ( .A(SYNOPSYS_UNCONNECTED_22), .B(
        _f_permutation__n2165 ), .ZN(_f_permutation__round_in[1066]) );
  NAND2_X2 _f_permutation__U1069  ( .A1(padder_out[43]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2164 ) );
  XNOR2_X2 _f_permutation__U1068  ( .A(SYNOPSYS_UNCONNECTED_21), .B(
        _f_permutation__n2164 ), .ZN(_f_permutation__round_in[1067]) );
  NAND2_X2 _f_permutation__U1067  ( .A1(padder_out[44]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2163 ) );
  XNOR2_X2 _f_permutation__U1066  ( .A(SYNOPSYS_UNCONNECTED_20), .B(
        _f_permutation__n2163 ), .ZN(_f_permutation__round_in[1068]) );
  NAND2_X2 _f_permutation__U1065  ( .A1(padder_out[45]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2162 ) );
  XNOR2_X2 _f_permutation__U1064  ( .A(SYNOPSYS_UNCONNECTED_19), .B(
        _f_permutation__n2162 ), .ZN(_f_permutation__round_in[1069]) );
  NAND2_X2 _f_permutation__U1063  ( .A1(padder_out[46]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2161 ) );
  XNOR2_X2 _f_permutation__U1062  ( .A(SYNOPSYS_UNCONNECTED_18), .B(
        _f_permutation__n2161 ), .ZN(_f_permutation__round_in[1070]) );
  NAND2_X2 _f_permutation__U1061  ( .A1(padder_out[47]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2160 ) );
  XNOR2_X2 _f_permutation__U1060  ( .A(SYNOPSYS_UNCONNECTED_17), .B(
        _f_permutation__n2160 ), .ZN(_f_permutation__round_in[1071]) );
  NAND2_X2 _f_permutation__U1059  ( .A1(padder_out[48]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2159 ) );
  XNOR2_X2 _f_permutation__U1058  ( .A(SYNOPSYS_UNCONNECTED_16), .B(
        _f_permutation__n2159 ), .ZN(_f_permutation__round_in[1072]) );
  NAND2_X2 _f_permutation__U1057  ( .A1(padder_out[49]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2158 ) );
  XNOR2_X2 _f_permutation__U1056  ( .A(SYNOPSYS_UNCONNECTED_15), .B(
        _f_permutation__n2158 ), .ZN(_f_permutation__round_in[1073]) );
  NAND2_X2 _f_permutation__U1055  ( .A1(padder_out[50]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2157 ) );
  XNOR2_X2 _f_permutation__U1054  ( .A(SYNOPSYS_UNCONNECTED_14), .B(
        _f_permutation__n2157 ), .ZN(_f_permutation__round_in[1074]) );
  NAND2_X2 _f_permutation__U1053  ( .A1(padder_out[51]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2156 ) );
  XNOR2_X2 _f_permutation__U1052  ( .A(SYNOPSYS_UNCONNECTED_13), .B(
        _f_permutation__n2156 ), .ZN(_f_permutation__round_in[1075]) );
  NAND2_X2 _f_permutation__U1051  ( .A1(padder_out[52]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2155 ) );
  XNOR2_X2 _f_permutation__U1050  ( .A(SYNOPSYS_UNCONNECTED_12), .B(
        _f_permutation__n2155 ), .ZN(_f_permutation__round_in[1076]) );
  NAND2_X2 _f_permutation__U1049  ( .A1(padder_out[53]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2154 ) );
  XNOR2_X2 _f_permutation__U1048  ( .A(SYNOPSYS_UNCONNECTED_11), .B(
        _f_permutation__n2154 ), .ZN(_f_permutation__round_in[1077]) );
  NAND2_X2 _f_permutation__U1047  ( .A1(padder_out[54]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2153 ) );
  XNOR2_X2 _f_permutation__U1046  ( .A(SYNOPSYS_UNCONNECTED_10), .B(
        _f_permutation__n2153 ), .ZN(_f_permutation__round_in[1078]) );
  NAND2_X2 _f_permutation__U1045  ( .A1(padder_out[55]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2152 ) );
  XNOR2_X2 _f_permutation__U1044  ( .A(SYNOPSYS_UNCONNECTED_9), .B(
        _f_permutation__n2152 ), .ZN(_f_permutation__round_in[1079]) );
  NAND2_X2 _f_permutation__U1043  ( .A1(padder_out[56]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2151 ) );
  XNOR2_X2 _f_permutation__U1042  ( .A(SYNOPSYS_UNCONNECTED_8), .B(
        _f_permutation__n2151 ), .ZN(_f_permutation__round_in[1080]) );
  NAND2_X2 _f_permutation__U1041  ( .A1(padder_out[57]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2150 ) );
  XNOR2_X2 _f_permutation__U1040  ( .A(SYNOPSYS_UNCONNECTED_7), .B(
        _f_permutation__n2150 ), .ZN(_f_permutation__round_in[1081]) );
  NAND2_X2 _f_permutation__U1039  ( .A1(padder_out[58]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2149 ) );
  XNOR2_X2 _f_permutation__U1038  ( .A(SYNOPSYS_UNCONNECTED_6), .B(
        _f_permutation__n2149 ), .ZN(_f_permutation__round_in[1082]) );
  NAND2_X2 _f_permutation__U1037  ( .A1(padder_out[59]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2148 ) );
  XNOR2_X2 _f_permutation__U1036  ( .A(SYNOPSYS_UNCONNECTED_5), .B(
        _f_permutation__n2148 ), .ZN(_f_permutation__round_in[1083]) );
  NAND2_X2 _f_permutation__U1035  ( .A1(padder_out[60]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2147 ) );
  XNOR2_X2 _f_permutation__U1034  ( .A(SYNOPSYS_UNCONNECTED_4), .B(
        _f_permutation__n2147 ), .ZN(_f_permutation__round_in[1084]) );
  NAND2_X2 _f_permutation__U1033  ( .A1(padder_out[61]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2146 ) );
  XNOR2_X2 _f_permutation__U1032  ( .A(SYNOPSYS_UNCONNECTED_3), .B(
        _f_permutation__n2146 ), .ZN(_f_permutation__round_in[1085]) );
  NAND2_X2 _f_permutation__U1031  ( .A1(padder_out[62]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2145 ) );
  XNOR2_X2 _f_permutation__U1030  ( .A(SYNOPSYS_UNCONNECTED_2), .B(
        _f_permutation__n2145 ), .ZN(_f_permutation__round_in[1086]) );
  NAND2_X2 _f_permutation__U1029  ( .A1(padder_out[63]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2144 ) );
  XNOR2_X2 _f_permutation__U1028  ( .A(SYNOPSYS_UNCONNECTED_1), .B(
        _f_permutation__n2144 ), .ZN(_f_permutation__round_in[1087]) );
  NAND2_X2 _f_permutation__U1027  ( .A1(padder_out[64]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2143 ) );
  XNOR2_X2 _f_permutation__U1026  ( .A(out[56]), .B(_f_permutation__n2143 ), 
        .ZN(_f_permutation__round_in[1088]) );
  NAND2_X2 _f_permutation__U1025  ( .A1(padder_out[65]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2142 ) );
  XNOR2_X2 _f_permutation__U1024  ( .A(out[57]), .B(_f_permutation__n2142 ), 
        .ZN(_f_permutation__round_in[1089]) );
  NAND2_X2 _f_permutation__U1023  ( .A1(padder_out[66]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2141 ) );
  XNOR2_X2 _f_permutation__U1022  ( .A(out[58]), .B(_f_permutation__n2141 ), 
        .ZN(_f_permutation__round_in[1090]) );
  NAND2_X2 _f_permutation__U1021  ( .A1(padder_out[67]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2140 ) );
  XNOR2_X2 _f_permutation__U1020  ( .A(out[59]), .B(_f_permutation__n2140 ), 
        .ZN(_f_permutation__round_in[1091]) );
  NAND2_X2 _f_permutation__U1019  ( .A1(padder_out[68]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2139 ) );
  XNOR2_X2 _f_permutation__U1018  ( .A(out[60]), .B(_f_permutation__n2139 ), 
        .ZN(_f_permutation__round_in[1092]) );
  NAND2_X2 _f_permutation__U1017  ( .A1(padder_out[69]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2138 ) );
  XNOR2_X2 _f_permutation__U1016  ( .A(out[61]), .B(_f_permutation__n2138 ), 
        .ZN(_f_permutation__round_in[1093]) );
  NAND2_X2 _f_permutation__U1015  ( .A1(padder_out[70]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2137 ) );
  XNOR2_X2 _f_permutation__U1014  ( .A(out[62]), .B(_f_permutation__n2137 ), 
        .ZN(_f_permutation__round_in[1094]) );
  NAND2_X2 _f_permutation__U1013  ( .A1(padder_out[71]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2136 ) );
  XNOR2_X2 _f_permutation__U1012  ( .A(out[63]), .B(_f_permutation__n2136 ), 
        .ZN(_f_permutation__round_in[1095]) );
  NAND2_X2 _f_permutation__U1011  ( .A1(padder_out[72]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2135 ) );
  XNOR2_X2 _f_permutation__U1010  ( .A(out[48]), .B(_f_permutation__n2135 ), 
        .ZN(_f_permutation__round_in[1096]) );
  NAND2_X2 _f_permutation__U1009  ( .A1(padder_out[73]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2134 ) );
  XNOR2_X2 _f_permutation__U1008  ( .A(out[49]), .B(_f_permutation__n2134 ), 
        .ZN(_f_permutation__round_in[1097]) );
  NAND2_X2 _f_permutation__U1007  ( .A1(padder_out[74]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2133 ) );
  XNOR2_X2 _f_permutation__U1006  ( .A(out[50]), .B(_f_permutation__n2133 ), 
        .ZN(_f_permutation__round_in[1098]) );
  NAND2_X2 _f_permutation__U1005  ( .A1(padder_out[75]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2132 ) );
  XNOR2_X2 _f_permutation__U1004  ( .A(out[51]), .B(_f_permutation__n2132 ), 
        .ZN(_f_permutation__round_in[1099]) );
  NAND2_X2 _f_permutation__U1003  ( .A1(padder_out[76]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2131 ) );
  XNOR2_X2 _f_permutation__U1002  ( .A(out[52]), .B(_f_permutation__n2131 ), 
        .ZN(_f_permutation__round_in[1100]) );
  NAND2_X2 _f_permutation__U1001  ( .A1(padder_out[77]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2130 ) );
  XNOR2_X2 _f_permutation__U1000  ( .A(out[53]), .B(_f_permutation__n2130 ), 
        .ZN(_f_permutation__round_in[1101]) );
  NAND2_X2 _f_permutation__U999  ( .A1(padder_out[78]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2129 ) );
  XNOR2_X2 _f_permutation__U998  ( .A(out[54]), .B(_f_permutation__n2129 ), 
        .ZN(_f_permutation__round_in[1102]) );
  NAND2_X2 _f_permutation__U997  ( .A1(padder_out[79]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2128 ) );
  XNOR2_X2 _f_permutation__U996  ( .A(out[55]), .B(_f_permutation__n2128 ), 
        .ZN(_f_permutation__round_in[1103]) );
  NAND2_X2 _f_permutation__U995  ( .A1(padder_out[80]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2127 ) );
  XNOR2_X2 _f_permutation__U994  ( .A(out[40]), .B(_f_permutation__n2127 ), 
        .ZN(_f_permutation__round_in[1104]) );
  NAND2_X2 _f_permutation__U993  ( .A1(padder_out[81]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2126 ) );
  XNOR2_X2 _f_permutation__U992  ( .A(out[41]), .B(_f_permutation__n2126 ), 
        .ZN(_f_permutation__round_in[1105]) );
  NAND2_X2 _f_permutation__U991  ( .A1(padder_out[82]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2125 ) );
  XNOR2_X2 _f_permutation__U990  ( .A(out[42]), .B(_f_permutation__n2125 ), 
        .ZN(_f_permutation__round_in[1106]) );
  NAND2_X2 _f_permutation__U989  ( .A1(padder_out[83]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2124 ) );
  XNOR2_X2 _f_permutation__U988  ( .A(out[43]), .B(_f_permutation__n2124 ), 
        .ZN(_f_permutation__round_in[1107]) );
  NAND2_X2 _f_permutation__U987  ( .A1(padder_out[84]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2123 ) );
  XNOR2_X2 _f_permutation__U986  ( .A(out[44]), .B(_f_permutation__n2123 ), 
        .ZN(_f_permutation__round_in[1108]) );
  NAND2_X2 _f_permutation__U985  ( .A1(padder_out[85]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2122 ) );
  XNOR2_X2 _f_permutation__U984  ( .A(out[45]), .B(_f_permutation__n2122 ), 
        .ZN(_f_permutation__round_in[1109]) );
  NAND2_X2 _f_permutation__U983  ( .A1(padder_out[86]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2121 ) );
  XNOR2_X2 _f_permutation__U982  ( .A(out[46]), .B(_f_permutation__n2121 ), 
        .ZN(_f_permutation__round_in[1110]) );
  NAND2_X2 _f_permutation__U981  ( .A1(padder_out[87]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2120 ) );
  XNOR2_X2 _f_permutation__U980  ( .A(out[47]), .B(_f_permutation__n2120 ), 
        .ZN(_f_permutation__round_in[1111]) );
  NAND2_X2 _f_permutation__U979  ( .A1(padder_out[88]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2119 ) );
  XNOR2_X2 _f_permutation__U978  ( .A(out[32]), .B(_f_permutation__n2119 ), 
        .ZN(_f_permutation__round_in[1112]) );
  NAND2_X2 _f_permutation__U977  ( .A1(padder_out[89]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2118 ) );
  XNOR2_X2 _f_permutation__U976  ( .A(out[33]), .B(_f_permutation__n2118 ), 
        .ZN(_f_permutation__round_in[1113]) );
  NAND2_X2 _f_permutation__U975  ( .A1(padder_out[90]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2117 ) );
  XNOR2_X2 _f_permutation__U974  ( .A(out[34]), .B(_f_permutation__n2117 ), 
        .ZN(_f_permutation__round_in[1114]) );
  NAND2_X2 _f_permutation__U973  ( .A1(padder_out[91]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2116 ) );
  XNOR2_X2 _f_permutation__U972  ( .A(out[35]), .B(_f_permutation__n2116 ), 
        .ZN(_f_permutation__round_in[1115]) );
  NAND2_X2 _f_permutation__U971  ( .A1(padder_out[92]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2115 ) );
  XNOR2_X2 _f_permutation__U970  ( .A(out[36]), .B(_f_permutation__n2115 ), 
        .ZN(_f_permutation__round_in[1116]) );
  NAND2_X2 _f_permutation__U969  ( .A1(padder_out[93]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2114 ) );
  XNOR2_X2 _f_permutation__U968  ( .A(out[37]), .B(_f_permutation__n2114 ), 
        .ZN(_f_permutation__round_in[1117]) );
  NAND2_X2 _f_permutation__U967  ( .A1(padder_out[94]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2113 ) );
  XNOR2_X2 _f_permutation__U966  ( .A(out[38]), .B(_f_permutation__n2113 ), 
        .ZN(_f_permutation__round_in[1118]) );
  NAND2_X2 _f_permutation__U965  ( .A1(padder_out[95]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2112 ) );
  XNOR2_X2 _f_permutation__U964  ( .A(out[39]), .B(_f_permutation__n2112 ), 
        .ZN(_f_permutation__round_in[1119]) );
  NAND2_X2 _f_permutation__U963  ( .A1(padder_out[96]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2111 ) );
  XNOR2_X2 _f_permutation__U962  ( .A(out[24]), .B(_f_permutation__n2111 ), 
        .ZN(_f_permutation__round_in[1120]) );
  NAND2_X2 _f_permutation__U961  ( .A1(padder_out[97]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2110 ) );
  XNOR2_X2 _f_permutation__U960  ( .A(out[25]), .B(_f_permutation__n2110 ), 
        .ZN(_f_permutation__round_in[1121]) );
  NAND2_X2 _f_permutation__U959  ( .A1(padder_out[98]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2109 ) );
  XNOR2_X2 _f_permutation__U958  ( .A(out[26]), .B(_f_permutation__n2109 ), 
        .ZN(_f_permutation__round_in[1122]) );
  NAND2_X2 _f_permutation__U957  ( .A1(padder_out[99]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2108 ) );
  XNOR2_X2 _f_permutation__U956  ( .A(out[27]), .B(_f_permutation__n2108 ), 
        .ZN(_f_permutation__round_in[1123]) );
  NAND2_X2 _f_permutation__U955  ( .A1(padder_out[100]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2107 ) );
  XNOR2_X2 _f_permutation__U954  ( .A(out[28]), .B(_f_permutation__n2107 ), 
        .ZN(_f_permutation__round_in[1124]) );
  NAND2_X2 _f_permutation__U953  ( .A1(padder_out[101]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2106 ) );
  XNOR2_X2 _f_permutation__U952  ( .A(out[29]), .B(_f_permutation__n2106 ), 
        .ZN(_f_permutation__round_in[1125]) );
  NAND2_X2 _f_permutation__U951  ( .A1(padder_out[102]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2105 ) );
  XNOR2_X2 _f_permutation__U950  ( .A(out[30]), .B(_f_permutation__n2105 ), 
        .ZN(_f_permutation__round_in[1126]) );
  NAND2_X2 _f_permutation__U949  ( .A1(padder_out[103]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2104 ) );
  XNOR2_X2 _f_permutation__U948  ( .A(out[31]), .B(_f_permutation__n2104 ), 
        .ZN(_f_permutation__round_in[1127]) );
  NAND2_X2 _f_permutation__U947  ( .A1(padder_out[104]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2103 ) );
  XNOR2_X2 _f_permutation__U946  ( .A(out[16]), .B(_f_permutation__n2103 ), 
        .ZN(_f_permutation__round_in[1128]) );
  NAND2_X2 _f_permutation__U945  ( .A1(padder_out[105]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2102 ) );
  XNOR2_X2 _f_permutation__U944  ( .A(out[17]), .B(_f_permutation__n2102 ), 
        .ZN(_f_permutation__round_in[1129]) );
  NAND2_X2 _f_permutation__U943  ( .A1(padder_out[106]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2101 ) );
  XNOR2_X2 _f_permutation__U942  ( .A(out[18]), .B(_f_permutation__n2101 ), 
        .ZN(_f_permutation__round_in[1130]) );
  NAND2_X2 _f_permutation__U941  ( .A1(padder_out[107]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2100 ) );
  XNOR2_X2 _f_permutation__U940  ( .A(out[19]), .B(_f_permutation__n2100 ), 
        .ZN(_f_permutation__round_in[1131]) );
  NAND2_X2 _f_permutation__U939  ( .A1(padder_out[108]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2099 ) );
  XNOR2_X2 _f_permutation__U938  ( .A(out[20]), .B(_f_permutation__n2099 ), 
        .ZN(_f_permutation__round_in[1132]) );
  NAND2_X2 _f_permutation__U937  ( .A1(padder_out[109]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2098 ) );
  XNOR2_X2 _f_permutation__U936  ( .A(out[21]), .B(_f_permutation__n2098 ), 
        .ZN(_f_permutation__round_in[1133]) );
  NAND2_X2 _f_permutation__U935  ( .A1(padder_out[110]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2097 ) );
  XNOR2_X2 _f_permutation__U934  ( .A(out[22]), .B(_f_permutation__n2097 ), 
        .ZN(_f_permutation__round_in[1134]) );
  NAND2_X2 _f_permutation__U933  ( .A1(padder_out[111]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2096 ) );
  XNOR2_X2 _f_permutation__U932  ( .A(out[23]), .B(_f_permutation__n2096 ), 
        .ZN(_f_permutation__round_in[1135]) );
  NAND2_X2 _f_permutation__U931  ( .A1(padder_out[112]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2095 ) );
  XNOR2_X2 _f_permutation__U930  ( .A(out[8]), .B(_f_permutation__n2095 ), 
        .ZN(_f_permutation__round_in[1136]) );
  NAND2_X2 _f_permutation__U929  ( .A1(padder_out[113]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2094 ) );
  XNOR2_X2 _f_permutation__U928  ( .A(out[9]), .B(_f_permutation__n2094 ), 
        .ZN(_f_permutation__round_in[1137]) );
  NAND2_X2 _f_permutation__U927  ( .A1(padder_out[114]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2093 ) );
  XNOR2_X2 _f_permutation__U926  ( .A(out[10]), .B(_f_permutation__n2093 ), 
        .ZN(_f_permutation__round_in[1138]) );
  NAND2_X2 _f_permutation__U925  ( .A1(padder_out[115]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2092 ) );
  XNOR2_X2 _f_permutation__U924  ( .A(out[11]), .B(_f_permutation__n2092 ), 
        .ZN(_f_permutation__round_in[1139]) );
  NAND2_X2 _f_permutation__U923  ( .A1(padder_out[116]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2091 ) );
  XNOR2_X2 _f_permutation__U922  ( .A(out[12]), .B(_f_permutation__n2091 ), 
        .ZN(_f_permutation__round_in[1140]) );
  NAND2_X2 _f_permutation__U921  ( .A1(padder_out[117]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2090 ) );
  XNOR2_X2 _f_permutation__U920  ( .A(out[13]), .B(_f_permutation__n2090 ), 
        .ZN(_f_permutation__round_in[1141]) );
  NAND2_X2 _f_permutation__U919  ( .A1(padder_out[118]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2089 ) );
  XNOR2_X2 _f_permutation__U918  ( .A(out[14]), .B(_f_permutation__n2089 ), 
        .ZN(_f_permutation__round_in[1142]) );
  NAND2_X2 _f_permutation__U917  ( .A1(padder_out[119]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2088 ) );
  XNOR2_X2 _f_permutation__U916  ( .A(out[15]), .B(_f_permutation__n2088 ), 
        .ZN(_f_permutation__round_in[1143]) );
  NAND2_X2 _f_permutation__U915  ( .A1(padder_out[120]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2087 ) );
  XNOR2_X2 _f_permutation__U914  ( .A(out[0]), .B(_f_permutation__n2087 ), 
        .ZN(_f_permutation__round_in[1144]) );
  NAND2_X2 _f_permutation__U913  ( .A1(padder_out[121]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2086 ) );
  XNOR2_X2 _f_permutation__U912  ( .A(out[1]), .B(_f_permutation__n2086 ), 
        .ZN(_f_permutation__round_in[1145]) );
  NAND2_X2 _f_permutation__U911  ( .A1(padder_out[122]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2085 ) );
  XNOR2_X2 _f_permutation__U910  ( .A(out[2]), .B(_f_permutation__n2085 ), 
        .ZN(_f_permutation__round_in[1146]) );
  NAND2_X2 _f_permutation__U909  ( .A1(padder_out[123]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2084 ) );
  XNOR2_X2 _f_permutation__U908  ( .A(out[3]), .B(_f_permutation__n2084 ), 
        .ZN(_f_permutation__round_in[1147]) );
  NAND2_X2 _f_permutation__U907  ( .A1(padder_out[124]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2083 ) );
  XNOR2_X2 _f_permutation__U906  ( .A(out[4]), .B(_f_permutation__n2083 ), 
        .ZN(_f_permutation__round_in[1148]) );
  NAND2_X2 _f_permutation__U905  ( .A1(padder_out[125]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2082 ) );
  XNOR2_X2 _f_permutation__U904  ( .A(out[5]), .B(_f_permutation__n2082 ), 
        .ZN(_f_permutation__round_in[1149]) );
  NAND2_X2 _f_permutation__U903  ( .A1(padder_out[126]), .A2(
        _f_permutation__n7318 ), .ZN(_f_permutation__n2081 ) );
  XNOR2_X2 _f_permutation__U902  ( .A(out[6]), .B(_f_permutation__n2081 ), 
        .ZN(_f_permutation__round_in[1150]) );
  NAND2_X2 _f_permutation__U901  ( .A1(padder_out[127]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2080 ) );
  XNOR2_X2 _f_permutation__U900  ( .A(out[7]), .B(_f_permutation__n2080 ), 
        .ZN(_f_permutation__round_in[1151]) );
  NAND2_X2 _f_permutation__U899  ( .A1(padder_out[128]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2079 ) );
  XNOR2_X2 _f_permutation__U898  ( .A(out[120]), .B(_f_permutation__n2079 ), 
        .ZN(_f_permutation__round_in[1152]) );
  NAND2_X2 _f_permutation__U897  ( .A1(padder_out[129]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2078 ) );
  XNOR2_X2 _f_permutation__U896  ( .A(out[121]), .B(_f_permutation__n2078 ), 
        .ZN(_f_permutation__round_in[1153]) );
  NAND2_X2 _f_permutation__U895  ( .A1(padder_out[130]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2077 ) );
  XNOR2_X2 _f_permutation__U894  ( .A(out[122]), .B(_f_permutation__n2077 ), 
        .ZN(_f_permutation__round_in[1154]) );
  NAND2_X2 _f_permutation__U893  ( .A1(padder_out[131]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2076 ) );
  XNOR2_X2 _f_permutation__U892  ( .A(out[123]), .B(_f_permutation__n2076 ), 
        .ZN(_f_permutation__round_in[1155]) );
  NAND2_X2 _f_permutation__U891  ( .A1(padder_out[132]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2075 ) );
  XNOR2_X2 _f_permutation__U890  ( .A(out[124]), .B(_f_permutation__n2075 ), 
        .ZN(_f_permutation__round_in[1156]) );
  NAND2_X2 _f_permutation__U889  ( .A1(padder_out[133]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2074 ) );
  XNOR2_X2 _f_permutation__U888  ( .A(out[125]), .B(_f_permutation__n2074 ), 
        .ZN(_f_permutation__round_in[1157]) );
  NAND2_X2 _f_permutation__U887  ( .A1(padder_out[134]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2073 ) );
  XNOR2_X2 _f_permutation__U886  ( .A(out[126]), .B(_f_permutation__n2073 ), 
        .ZN(_f_permutation__round_in[1158]) );
  NAND2_X2 _f_permutation__U885  ( .A1(padder_out[135]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2072 ) );
  XNOR2_X2 _f_permutation__U884  ( .A(out[127]), .B(_f_permutation__n2072 ), 
        .ZN(_f_permutation__round_in[1159]) );
  NAND2_X2 _f_permutation__U883  ( .A1(padder_out[136]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2071 ) );
  XNOR2_X2 _f_permutation__U882  ( .A(out[112]), .B(_f_permutation__n2071 ), 
        .ZN(_f_permutation__round_in[1160]) );
  NAND2_X2 _f_permutation__U881  ( .A1(padder_out[137]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2070 ) );
  XNOR2_X2 _f_permutation__U880  ( .A(out[113]), .B(_f_permutation__n2070 ), 
        .ZN(_f_permutation__round_in[1161]) );
  NAND2_X2 _f_permutation__U879  ( .A1(padder_out[138]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2069 ) );
  XNOR2_X2 _f_permutation__U878  ( .A(out[114]), .B(_f_permutation__n2069 ), 
        .ZN(_f_permutation__round_in[1162]) );
  NAND2_X2 _f_permutation__U877  ( .A1(padder_out[139]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2068 ) );
  XNOR2_X2 _f_permutation__U876  ( .A(out[115]), .B(_f_permutation__n2068 ), 
        .ZN(_f_permutation__round_in[1163]) );
  NAND2_X2 _f_permutation__U875  ( .A1(padder_out[140]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2067 ) );
  XNOR2_X2 _f_permutation__U874  ( .A(out[116]), .B(_f_permutation__n2067 ), 
        .ZN(_f_permutation__round_in[1164]) );
  NAND2_X2 _f_permutation__U873  ( .A1(padder_out[141]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2066 ) );
  XNOR2_X2 _f_permutation__U872  ( .A(out[117]), .B(_f_permutation__n2066 ), 
        .ZN(_f_permutation__round_in[1165]) );
  NAND2_X2 _f_permutation__U871  ( .A1(padder_out[142]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2065 ) );
  XNOR2_X2 _f_permutation__U870  ( .A(out[118]), .B(_f_permutation__n2065 ), 
        .ZN(_f_permutation__round_in[1166]) );
  NAND2_X2 _f_permutation__U869  ( .A1(padder_out[143]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n2064 ) );
  XNOR2_X2 _f_permutation__U868  ( .A(out[119]), .B(_f_permutation__n2064 ), 
        .ZN(_f_permutation__round_in[1167]) );
  NAND2_X2 _f_permutation__U867  ( .A1(padder_out[144]), .A2(
        _f_permutation__n7319 ), .ZN(_f_permutation__n2063 ) );
  XNOR2_X2 _f_permutation__U866  ( .A(out[104]), .B(_f_permutation__n2063 ), 
        .ZN(_f_permutation__round_in[1168]) );
  NAND2_X2 _f_permutation__U865  ( .A1(padder_out[145]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2062 ) );
  XNOR2_X2 _f_permutation__U864  ( .A(out[105]), .B(_f_permutation__n2062 ), 
        .ZN(_f_permutation__round_in[1169]) );
  NAND2_X2 _f_permutation__U863  ( .A1(padder_out[146]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2061 ) );
  XNOR2_X2 _f_permutation__U862  ( .A(out[106]), .B(_f_permutation__n2061 ), 
        .ZN(_f_permutation__round_in[1170]) );
  NAND2_X2 _f_permutation__U861  ( .A1(padder_out[147]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2060 ) );
  XNOR2_X2 _f_permutation__U860  ( .A(out[107]), .B(_f_permutation__n2060 ), 
        .ZN(_f_permutation__round_in[1171]) );
  NAND2_X2 _f_permutation__U859  ( .A1(padder_out[148]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2059 ) );
  XNOR2_X2 _f_permutation__U858  ( .A(out[108]), .B(_f_permutation__n2059 ), 
        .ZN(_f_permutation__round_in[1172]) );
  NAND2_X2 _f_permutation__U857  ( .A1(padder_out[149]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2058 ) );
  XNOR2_X2 _f_permutation__U856  ( .A(out[109]), .B(_f_permutation__n2058 ), 
        .ZN(_f_permutation__round_in[1173]) );
  NAND2_X2 _f_permutation__U855  ( .A1(padder_out[150]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2057 ) );
  XNOR2_X2 _f_permutation__U854  ( .A(out[110]), .B(_f_permutation__n2057 ), 
        .ZN(_f_permutation__round_in[1174]) );
  NAND2_X2 _f_permutation__U853  ( .A1(padder_out[151]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2056 ) );
  XNOR2_X2 _f_permutation__U852  ( .A(out[111]), .B(_f_permutation__n2056 ), 
        .ZN(_f_permutation__round_in[1175]) );
  NAND2_X2 _f_permutation__U851  ( .A1(padder_out[152]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2055 ) );
  XNOR2_X2 _f_permutation__U850  ( .A(out[96]), .B(_f_permutation__n2055 ), 
        .ZN(_f_permutation__round_in[1176]) );
  NAND2_X2 _f_permutation__U849  ( .A1(padder_out[153]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2054 ) );
  XNOR2_X2 _f_permutation__U848  ( .A(out[97]), .B(_f_permutation__n2054 ), 
        .ZN(_f_permutation__round_in[1177]) );
  NAND2_X2 _f_permutation__U847  ( .A1(padder_out[154]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2053 ) );
  XNOR2_X2 _f_permutation__U846  ( .A(out[98]), .B(_f_permutation__n2053 ), 
        .ZN(_f_permutation__round_in[1178]) );
  NAND2_X2 _f_permutation__U845  ( .A1(padder_out[155]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2052 ) );
  XNOR2_X2 _f_permutation__U844  ( .A(out[99]), .B(_f_permutation__n2052 ), 
        .ZN(_f_permutation__round_in[1179]) );
  NAND2_X2 _f_permutation__U843  ( .A1(padder_out[156]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2051 ) );
  XNOR2_X2 _f_permutation__U842  ( .A(out[100]), .B(_f_permutation__n2051 ), 
        .ZN(_f_permutation__round_in[1180]) );
  NAND2_X2 _f_permutation__U841  ( .A1(padder_out[157]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2050 ) );
  XNOR2_X2 _f_permutation__U840  ( .A(out[101]), .B(_f_permutation__n2050 ), 
        .ZN(_f_permutation__round_in[1181]) );
  NAND2_X2 _f_permutation__U839  ( .A1(padder_out[158]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2049 ) );
  XNOR2_X2 _f_permutation__U838  ( .A(out[102]), .B(_f_permutation__n2049 ), 
        .ZN(_f_permutation__round_in[1182]) );
  NAND2_X2 _f_permutation__U837  ( .A1(padder_out[159]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2048 ) );
  XNOR2_X2 _f_permutation__U836  ( .A(out[103]), .B(_f_permutation__n2048 ), 
        .ZN(_f_permutation__round_in[1183]) );
  NAND2_X2 _f_permutation__U835  ( .A1(padder_out[160]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2047 ) );
  XNOR2_X2 _f_permutation__U834  ( .A(out[88]), .B(_f_permutation__n2047 ), 
        .ZN(_f_permutation__round_in[1184]) );
  NAND2_X2 _f_permutation__U833  ( .A1(padder_out[161]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2046 ) );
  XNOR2_X2 _f_permutation__U832  ( .A(out[89]), .B(_f_permutation__n2046 ), 
        .ZN(_f_permutation__round_in[1185]) );
  NAND2_X2 _f_permutation__U831  ( .A1(padder_out[162]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2045 ) );
  XNOR2_X2 _f_permutation__U830  ( .A(out[90]), .B(_f_permutation__n2045 ), 
        .ZN(_f_permutation__round_in[1186]) );
  NAND2_X2 _f_permutation__U829  ( .A1(padder_out[163]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2044 ) );
  XNOR2_X2 _f_permutation__U828  ( .A(out[91]), .B(_f_permutation__n2044 ), 
        .ZN(_f_permutation__round_in[1187]) );
  NAND2_X2 _f_permutation__U827  ( .A1(padder_out[164]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2043 ) );
  XNOR2_X2 _f_permutation__U826  ( .A(out[92]), .B(_f_permutation__n2043 ), 
        .ZN(_f_permutation__round_in[1188]) );
  NAND2_X2 _f_permutation__U825  ( .A1(padder_out[165]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2042 ) );
  XNOR2_X2 _f_permutation__U824  ( .A(out[93]), .B(_f_permutation__n2042 ), 
        .ZN(_f_permutation__round_in[1189]) );
  NAND2_X2 _f_permutation__U823  ( .A1(padder_out[166]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2041 ) );
  XNOR2_X2 _f_permutation__U822  ( .A(out[94]), .B(_f_permutation__n2041 ), 
        .ZN(_f_permutation__round_in[1190]) );
  NAND2_X2 _f_permutation__U821  ( .A1(padder_out[167]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2040 ) );
  XNOR2_X2 _f_permutation__U820  ( .A(out[95]), .B(_f_permutation__n2040 ), 
        .ZN(_f_permutation__round_in[1191]) );
  NAND2_X2 _f_permutation__U819  ( .A1(padder_out[168]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2039 ) );
  XNOR2_X2 _f_permutation__U818  ( .A(out[80]), .B(_f_permutation__n2039 ), 
        .ZN(_f_permutation__round_in[1192]) );
  NAND2_X2 _f_permutation__U817  ( .A1(padder_out[169]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2038 ) );
  XNOR2_X2 _f_permutation__U816  ( .A(out[81]), .B(_f_permutation__n2038 ), 
        .ZN(_f_permutation__round_in[1193]) );
  NAND2_X2 _f_permutation__U815  ( .A1(padder_out[170]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2037 ) );
  XNOR2_X2 _f_permutation__U814  ( .A(out[82]), .B(_f_permutation__n2037 ), 
        .ZN(_f_permutation__round_in[1194]) );
  NAND2_X2 _f_permutation__U813  ( .A1(padder_out[171]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2036 ) );
  XNOR2_X2 _f_permutation__U812  ( .A(out[83]), .B(_f_permutation__n2036 ), 
        .ZN(_f_permutation__round_in[1195]) );
  NAND2_X2 _f_permutation__U811  ( .A1(padder_out[172]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2035 ) );
  XNOR2_X2 _f_permutation__U810  ( .A(out[84]), .B(_f_permutation__n2035 ), 
        .ZN(_f_permutation__round_in[1196]) );
  NAND2_X2 _f_permutation__U809  ( .A1(padder_out[173]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2034 ) );
  XNOR2_X2 _f_permutation__U808  ( .A(out[85]), .B(_f_permutation__n2034 ), 
        .ZN(_f_permutation__round_in[1197]) );
  NAND2_X2 _f_permutation__U807  ( .A1(padder_out[174]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2033 ) );
  XNOR2_X2 _f_permutation__U806  ( .A(out[86]), .B(_f_permutation__n2033 ), 
        .ZN(_f_permutation__round_in[1198]) );
  NAND2_X2 _f_permutation__U805  ( .A1(padder_out[175]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2032 ) );
  XNOR2_X2 _f_permutation__U804  ( .A(out[87]), .B(_f_permutation__n2032 ), 
        .ZN(_f_permutation__round_in[1199]) );
  NAND2_X2 _f_permutation__U803  ( .A1(padder_out[176]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2031 ) );
  XNOR2_X2 _f_permutation__U802  ( .A(out[72]), .B(_f_permutation__n2031 ), 
        .ZN(_f_permutation__round_in[1200]) );
  NAND2_X2 _f_permutation__U801  ( .A1(padder_out[177]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2030 ) );
  XNOR2_X2 _f_permutation__U800  ( .A(out[73]), .B(_f_permutation__n2030 ), 
        .ZN(_f_permutation__round_in[1201]) );
  NAND2_X2 _f_permutation__U799  ( .A1(padder_out[178]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2029 ) );
  XNOR2_X2 _f_permutation__U798  ( .A(out[74]), .B(_f_permutation__n2029 ), 
        .ZN(_f_permutation__round_in[1202]) );
  NAND2_X2 _f_permutation__U797  ( .A1(padder_out[179]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2028 ) );
  XNOR2_X2 _f_permutation__U796  ( .A(out[75]), .B(_f_permutation__n2028 ), 
        .ZN(_f_permutation__round_in[1203]) );
  NAND2_X2 _f_permutation__U795  ( .A1(padder_out[180]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2027 ) );
  XNOR2_X2 _f_permutation__U794  ( .A(out[76]), .B(_f_permutation__n2027 ), 
        .ZN(_f_permutation__round_in[1204]) );
  NAND2_X2 _f_permutation__U793  ( .A1(padder_out[181]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2026 ) );
  XNOR2_X2 _f_permutation__U792  ( .A(out[77]), .B(_f_permutation__n2026 ), 
        .ZN(_f_permutation__round_in[1205]) );
  NAND2_X2 _f_permutation__U791  ( .A1(padder_out[182]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2025 ) );
  XNOR2_X2 _f_permutation__U790  ( .A(out[78]), .B(_f_permutation__n2025 ), 
        .ZN(_f_permutation__round_in[1206]) );
  NAND2_X2 _f_permutation__U789  ( .A1(padder_out[183]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2024 ) );
  XNOR2_X2 _f_permutation__U788  ( .A(out[79]), .B(_f_permutation__n2024 ), 
        .ZN(_f_permutation__round_in[1207]) );
  NAND2_X2 _f_permutation__U787  ( .A1(padder_out[184]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2023 ) );
  XNOR2_X2 _f_permutation__U786  ( .A(out[64]), .B(_f_permutation__n2023 ), 
        .ZN(_f_permutation__round_in[1208]) );
  NAND2_X2 _f_permutation__U785  ( .A1(padder_out[185]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2022 ) );
  XNOR2_X2 _f_permutation__U784  ( .A(out[65]), .B(_f_permutation__n2022 ), 
        .ZN(_f_permutation__round_in[1209]) );
  NAND2_X2 _f_permutation__U783  ( .A1(padder_out[186]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2021 ) );
  XNOR2_X2 _f_permutation__U782  ( .A(out[66]), .B(_f_permutation__n2021 ), 
        .ZN(_f_permutation__round_in[1210]) );
  NAND2_X2 _f_permutation__U781  ( .A1(padder_out[187]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2020 ) );
  XNOR2_X2 _f_permutation__U780  ( .A(out[67]), .B(_f_permutation__n2020 ), 
        .ZN(_f_permutation__round_in[1211]) );
  NAND2_X2 _f_permutation__U779  ( .A1(padder_out[188]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2019 ) );
  XNOR2_X2 _f_permutation__U778  ( .A(out[68]), .B(_f_permutation__n2019 ), 
        .ZN(_f_permutation__round_in[1212]) );
  NAND2_X2 _f_permutation__U777  ( .A1(padder_out[189]), .A2(
        _f_permutation__n7323 ), .ZN(_f_permutation__n2018 ) );
  XNOR2_X2 _f_permutation__U776  ( .A(out[69]), .B(_f_permutation__n2018 ), 
        .ZN(_f_permutation__round_in[1213]) );
  NAND2_X2 _f_permutation__U775  ( .A1(padder_out[190]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2017 ) );
  XNOR2_X2 _f_permutation__U774  ( .A(out[70]), .B(_f_permutation__n2017 ), 
        .ZN(_f_permutation__round_in[1214]) );
  NAND2_X2 _f_permutation__U773  ( .A1(padder_out[191]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2016 ) );
  XNOR2_X2 _f_permutation__U772  ( .A(out[71]), .B(_f_permutation__n2016 ), 
        .ZN(_f_permutation__round_in[1215]) );
  NAND2_X2 _f_permutation__U771  ( .A1(padder_out[192]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2015 ) );
  XNOR2_X2 _f_permutation__U770  ( .A(out[184]), .B(_f_permutation__n2015 ), 
        .ZN(_f_permutation__round_in[1216]) );
  NAND2_X2 _f_permutation__U769  ( .A1(padder_out[193]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2014 ) );
  XNOR2_X2 _f_permutation__U768  ( .A(out[185]), .B(_f_permutation__n2014 ), 
        .ZN(_f_permutation__round_in[1217]) );
  NAND2_X2 _f_permutation__U767  ( .A1(padder_out[194]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2013 ) );
  XNOR2_X2 _f_permutation__U766  ( .A(out[186]), .B(_f_permutation__n2013 ), 
        .ZN(_f_permutation__round_in[1218]) );
  NAND2_X2 _f_permutation__U765  ( .A1(padder_out[195]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2012 ) );
  XNOR2_X2 _f_permutation__U764  ( .A(out[187]), .B(_f_permutation__n2012 ), 
        .ZN(_f_permutation__round_in[1219]) );
  NAND2_X2 _f_permutation__U763  ( .A1(padder_out[196]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2011 ) );
  XNOR2_X2 _f_permutation__U762  ( .A(out[188]), .B(_f_permutation__n2011 ), 
        .ZN(_f_permutation__round_in[1220]) );
  NAND2_X2 _f_permutation__U761  ( .A1(padder_out[197]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2010 ) );
  XNOR2_X2 _f_permutation__U760  ( .A(out[189]), .B(_f_permutation__n2010 ), 
        .ZN(_f_permutation__round_in[1221]) );
  NAND2_X2 _f_permutation__U759  ( .A1(padder_out[198]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2009 ) );
  XNOR2_X2 _f_permutation__U758  ( .A(out[190]), .B(_f_permutation__n2009 ), 
        .ZN(_f_permutation__round_in[1222]) );
  NAND2_X2 _f_permutation__U757  ( .A1(padder_out[199]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2008 ) );
  XNOR2_X2 _f_permutation__U756  ( .A(out[191]), .B(_f_permutation__n2008 ), 
        .ZN(_f_permutation__round_in[1223]) );
  NAND2_X2 _f_permutation__U755  ( .A1(padder_out[200]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2007 ) );
  XNOR2_X2 _f_permutation__U754  ( .A(out[176]), .B(_f_permutation__n2007 ), 
        .ZN(_f_permutation__round_in[1224]) );
  NAND2_X2 _f_permutation__U753  ( .A1(padder_out[201]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2006 ) );
  XNOR2_X2 _f_permutation__U752  ( .A(out[177]), .B(_f_permutation__n2006 ), 
        .ZN(_f_permutation__round_in[1225]) );
  NAND2_X2 _f_permutation__U751  ( .A1(padder_out[202]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2005 ) );
  XNOR2_X2 _f_permutation__U750  ( .A(out[178]), .B(_f_permutation__n2005 ), 
        .ZN(_f_permutation__round_in[1226]) );
  NAND2_X2 _f_permutation__U749  ( .A1(padder_out[203]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2004 ) );
  XNOR2_X2 _f_permutation__U748  ( .A(out[179]), .B(_f_permutation__n2004 ), 
        .ZN(_f_permutation__round_in[1227]) );
  NAND2_X2 _f_permutation__U747  ( .A1(padder_out[204]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2003 ) );
  XNOR2_X2 _f_permutation__U746  ( .A(out[180]), .B(_f_permutation__n2003 ), 
        .ZN(_f_permutation__round_in[1228]) );
  NAND2_X2 _f_permutation__U745  ( .A1(padder_out[205]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2002 ) );
  XNOR2_X2 _f_permutation__U744  ( .A(out[181]), .B(_f_permutation__n2002 ), 
        .ZN(_f_permutation__round_in[1229]) );
  NAND2_X2 _f_permutation__U743  ( .A1(padder_out[206]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2001 ) );
  XNOR2_X2 _f_permutation__U742  ( .A(out[182]), .B(_f_permutation__n2001 ), 
        .ZN(_f_permutation__round_in[1230]) );
  NAND2_X2 _f_permutation__U741  ( .A1(padder_out[207]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n2000 ) );
  XNOR2_X2 _f_permutation__U740  ( .A(out[183]), .B(_f_permutation__n2000 ), 
        .ZN(_f_permutation__round_in[1231]) );
  NAND2_X2 _f_permutation__U739  ( .A1(padder_out[208]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1999 ) );
  XNOR2_X2 _f_permutation__U738  ( .A(out[168]), .B(_f_permutation__n1999 ), 
        .ZN(_f_permutation__round_in[1232]) );
  NAND2_X2 _f_permutation__U737  ( .A1(padder_out[209]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1998 ) );
  XNOR2_X2 _f_permutation__U736  ( .A(out[169]), .B(_f_permutation__n1998 ), 
        .ZN(_f_permutation__round_in[1233]) );
  NAND2_X2 _f_permutation__U735  ( .A1(padder_out[210]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1997 ) );
  XNOR2_X2 _f_permutation__U734  ( .A(out[170]), .B(_f_permutation__n1997 ), 
        .ZN(_f_permutation__round_in[1234]) );
  NAND2_X2 _f_permutation__U733  ( .A1(padder_out[211]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1996 ) );
  XNOR2_X2 _f_permutation__U732  ( .A(out[171]), .B(_f_permutation__n1996 ), 
        .ZN(_f_permutation__round_in[1235]) );
  NAND2_X2 _f_permutation__U731  ( .A1(padder_out[212]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1995 ) );
  XNOR2_X2 _f_permutation__U730  ( .A(out[172]), .B(_f_permutation__n1995 ), 
        .ZN(_f_permutation__round_in[1236]) );
  NAND2_X2 _f_permutation__U729  ( .A1(padder_out[213]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1994 ) );
  XNOR2_X2 _f_permutation__U728  ( .A(out[173]), .B(_f_permutation__n1994 ), 
        .ZN(_f_permutation__round_in[1237]) );
  NAND2_X2 _f_permutation__U727  ( .A1(padder_out[214]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1993 ) );
  XNOR2_X2 _f_permutation__U726  ( .A(out[174]), .B(_f_permutation__n1993 ), 
        .ZN(_f_permutation__round_in[1238]) );
  NAND2_X2 _f_permutation__U725  ( .A1(padder_out[215]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1992 ) );
  XNOR2_X2 _f_permutation__U724  ( .A(out[175]), .B(_f_permutation__n1992 ), 
        .ZN(_f_permutation__round_in[1239]) );
  NAND2_X2 _f_permutation__U723  ( .A1(padder_out[216]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1991 ) );
  XNOR2_X2 _f_permutation__U722  ( .A(out[160]), .B(_f_permutation__n1991 ), 
        .ZN(_f_permutation__round_in[1240]) );
  NAND2_X2 _f_permutation__U721  ( .A1(padder_out[217]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1990 ) );
  XNOR2_X2 _f_permutation__U720  ( .A(out[161]), .B(_f_permutation__n1990 ), 
        .ZN(_f_permutation__round_in[1241]) );
  NAND2_X2 _f_permutation__U719  ( .A1(padder_out[218]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1989 ) );
  XNOR2_X2 _f_permutation__U718  ( .A(out[162]), .B(_f_permutation__n1989 ), 
        .ZN(_f_permutation__round_in[1242]) );
  NAND2_X2 _f_permutation__U717  ( .A1(padder_out[219]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1988 ) );
  XNOR2_X2 _f_permutation__U716  ( .A(out[163]), .B(_f_permutation__n1988 ), 
        .ZN(_f_permutation__round_in[1243]) );
  NAND2_X2 _f_permutation__U715  ( .A1(padder_out[220]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1987 ) );
  XNOR2_X2 _f_permutation__U714  ( .A(out[164]), .B(_f_permutation__n1987 ), 
        .ZN(_f_permutation__round_in[1244]) );
  NAND2_X2 _f_permutation__U713  ( .A1(padder_out[221]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1986 ) );
  XNOR2_X2 _f_permutation__U712  ( .A(out[165]), .B(_f_permutation__n1986 ), 
        .ZN(_f_permutation__round_in[1245]) );
  NAND2_X2 _f_permutation__U711  ( .A1(padder_out[222]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1985 ) );
  XNOR2_X2 _f_permutation__U710  ( .A(out[166]), .B(_f_permutation__n1985 ), 
        .ZN(_f_permutation__round_in[1246]) );
  NAND2_X2 _f_permutation__U709  ( .A1(padder_out[223]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1984 ) );
  XNOR2_X2 _f_permutation__U708  ( .A(out[167]), .B(_f_permutation__n1984 ), 
        .ZN(_f_permutation__round_in[1247]) );
  NAND2_X2 _f_permutation__U707  ( .A1(padder_out[224]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1983 ) );
  XNOR2_X2 _f_permutation__U706  ( .A(out[152]), .B(_f_permutation__n1983 ), 
        .ZN(_f_permutation__round_in[1248]) );
  NAND2_X2 _f_permutation__U705  ( .A1(padder_out[225]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1982 ) );
  XNOR2_X2 _f_permutation__U704  ( .A(out[153]), .B(_f_permutation__n1982 ), 
        .ZN(_f_permutation__round_in[1249]) );
  NAND2_X2 _f_permutation__U703  ( .A1(padder_out[226]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1981 ) );
  XNOR2_X2 _f_permutation__U702  ( .A(out[154]), .B(_f_permutation__n1981 ), 
        .ZN(_f_permutation__round_in[1250]) );
  NAND2_X2 _f_permutation__U701  ( .A1(padder_out[227]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1980 ) );
  XNOR2_X2 _f_permutation__U700  ( .A(out[155]), .B(_f_permutation__n1980 ), 
        .ZN(_f_permutation__round_in[1251]) );
  NAND2_X2 _f_permutation__U699  ( .A1(padder_out[228]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1979 ) );
  XNOR2_X2 _f_permutation__U698  ( .A(out[156]), .B(_f_permutation__n1979 ), 
        .ZN(_f_permutation__round_in[1252]) );
  NAND2_X2 _f_permutation__U697  ( .A1(padder_out[229]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1978 ) );
  XNOR2_X2 _f_permutation__U696  ( .A(out[157]), .B(_f_permutation__n1978 ), 
        .ZN(_f_permutation__round_in[1253]) );
  NAND2_X2 _f_permutation__U695  ( .A1(padder_out[230]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1977 ) );
  XNOR2_X2 _f_permutation__U694  ( .A(out[158]), .B(_f_permutation__n1977 ), 
        .ZN(_f_permutation__round_in[1254]) );
  NAND2_X2 _f_permutation__U693  ( .A1(padder_out[231]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1976 ) );
  XNOR2_X2 _f_permutation__U692  ( .A(out[159]), .B(_f_permutation__n1976 ), 
        .ZN(_f_permutation__round_in[1255]) );
  NAND2_X2 _f_permutation__U691  ( .A1(padder_out[232]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1975 ) );
  XNOR2_X2 _f_permutation__U690  ( .A(out[144]), .B(_f_permutation__n1975 ), 
        .ZN(_f_permutation__round_in[1256]) );
  NAND2_X2 _f_permutation__U689  ( .A1(padder_out[233]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1974 ) );
  XNOR2_X2 _f_permutation__U688  ( .A(out[145]), .B(_f_permutation__n1974 ), 
        .ZN(_f_permutation__round_in[1257]) );
  NAND2_X2 _f_permutation__U687  ( .A1(padder_out[234]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1973 ) );
  XNOR2_X2 _f_permutation__U686  ( .A(out[146]), .B(_f_permutation__n1973 ), 
        .ZN(_f_permutation__round_in[1258]) );
  NAND2_X2 _f_permutation__U685  ( .A1(padder_out[235]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1972 ) );
  XNOR2_X2 _f_permutation__U684  ( .A(out[147]), .B(_f_permutation__n1972 ), 
        .ZN(_f_permutation__round_in[1259]) );
  NAND2_X2 _f_permutation__U683  ( .A1(padder_out[236]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1971 ) );
  XNOR2_X2 _f_permutation__U682  ( .A(out[148]), .B(_f_permutation__n1971 ), 
        .ZN(_f_permutation__round_in[1260]) );
  NAND2_X2 _f_permutation__U681  ( .A1(padder_out[237]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1970 ) );
  XNOR2_X2 _f_permutation__U680  ( .A(out[149]), .B(_f_permutation__n1970 ), 
        .ZN(_f_permutation__round_in[1261]) );
  NAND2_X2 _f_permutation__U679  ( .A1(padder_out[238]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1969 ) );
  XNOR2_X2 _f_permutation__U678  ( .A(out[150]), .B(_f_permutation__n1969 ), 
        .ZN(_f_permutation__round_in[1262]) );
  NAND2_X2 _f_permutation__U677  ( .A1(padder_out[239]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1968 ) );
  XNOR2_X2 _f_permutation__U676  ( .A(out[151]), .B(_f_permutation__n1968 ), 
        .ZN(_f_permutation__round_in[1263]) );
  NAND2_X2 _f_permutation__U675  ( .A1(padder_out[240]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1967 ) );
  XNOR2_X2 _f_permutation__U674  ( .A(out[136]), .B(_f_permutation__n1967 ), 
        .ZN(_f_permutation__round_in[1264]) );
  NAND2_X2 _f_permutation__U673  ( .A1(padder_out[241]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1966 ) );
  XNOR2_X2 _f_permutation__U672  ( .A(out[137]), .B(_f_permutation__n1966 ), 
        .ZN(_f_permutation__round_in[1265]) );
  NAND2_X2 _f_permutation__U671  ( .A1(padder_out[242]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1965 ) );
  XNOR2_X2 _f_permutation__U670  ( .A(out[138]), .B(_f_permutation__n1965 ), 
        .ZN(_f_permutation__round_in[1266]) );
  NAND2_X2 _f_permutation__U669  ( .A1(padder_out[243]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1964 ) );
  XNOR2_X2 _f_permutation__U668  ( .A(out[139]), .B(_f_permutation__n1964 ), 
        .ZN(_f_permutation__round_in[1267]) );
  NAND2_X2 _f_permutation__U667  ( .A1(padder_out[244]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1963 ) );
  XNOR2_X2 _f_permutation__U666  ( .A(out[140]), .B(_f_permutation__n1963 ), 
        .ZN(_f_permutation__round_in[1268]) );
  NAND2_X2 _f_permutation__U665  ( .A1(padder_out[245]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1962 ) );
  XNOR2_X2 _f_permutation__U664  ( .A(out[141]), .B(_f_permutation__n1962 ), 
        .ZN(_f_permutation__round_in[1269]) );
  NAND2_X2 _f_permutation__U663  ( .A1(padder_out[246]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1961 ) );
  XNOR2_X2 _f_permutation__U662  ( .A(out[142]), .B(_f_permutation__n1961 ), 
        .ZN(_f_permutation__round_in[1270]) );
  NAND2_X2 _f_permutation__U661  ( .A1(padder_out[247]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1960 ) );
  XNOR2_X2 _f_permutation__U660  ( .A(out[143]), .B(_f_permutation__n1960 ), 
        .ZN(_f_permutation__round_in[1271]) );
  NAND2_X2 _f_permutation__U659  ( .A1(padder_out[248]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1959 ) );
  XNOR2_X2 _f_permutation__U658  ( .A(out[128]), .B(_f_permutation__n1959 ), 
        .ZN(_f_permutation__round_in[1272]) );
  NAND2_X2 _f_permutation__U657  ( .A1(padder_out[249]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1958 ) );
  XNOR2_X2 _f_permutation__U656  ( .A(out[129]), .B(_f_permutation__n1958 ), 
        .ZN(_f_permutation__round_in[1273]) );
  NAND2_X2 _f_permutation__U655  ( .A1(padder_out[250]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1957 ) );
  XNOR2_X2 _f_permutation__U654  ( .A(out[130]), .B(_f_permutation__n1957 ), 
        .ZN(_f_permutation__round_in[1274]) );
  NAND2_X2 _f_permutation__U653  ( .A1(padder_out[251]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1956 ) );
  XNOR2_X2 _f_permutation__U652  ( .A(out[131]), .B(_f_permutation__n1956 ), 
        .ZN(_f_permutation__round_in[1275]) );
  NAND2_X2 _f_permutation__U651  ( .A1(padder_out[252]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1955 ) );
  XNOR2_X2 _f_permutation__U650  ( .A(out[132]), .B(_f_permutation__n1955 ), 
        .ZN(_f_permutation__round_in[1276]) );
  NAND2_X2 _f_permutation__U649  ( .A1(padder_out[253]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1954 ) );
  XNOR2_X2 _f_permutation__U648  ( .A(out[133]), .B(_f_permutation__n1954 ), 
        .ZN(_f_permutation__round_in[1277]) );
  NAND2_X2 _f_permutation__U647  ( .A1(padder_out[254]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1953 ) );
  XNOR2_X2 _f_permutation__U646  ( .A(out[134]), .B(_f_permutation__n1953 ), 
        .ZN(_f_permutation__round_in[1278]) );
  NAND2_X2 _f_permutation__U645  ( .A1(padder_out[255]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1952 ) );
  XNOR2_X2 _f_permutation__U644  ( .A(out[135]), .B(_f_permutation__n1952 ), 
        .ZN(_f_permutation__round_in[1279]) );
  NAND2_X2 _f_permutation__U643  ( .A1(padder_out[256]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1951 ) );
  XNOR2_X2 _f_permutation__U642  ( .A(out[248]), .B(_f_permutation__n1951 ), 
        .ZN(_f_permutation__round_in[1280]) );
  NAND2_X2 _f_permutation__U641  ( .A1(padder_out[257]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1950 ) );
  XNOR2_X2 _f_permutation__U640  ( .A(out[249]), .B(_f_permutation__n1950 ), 
        .ZN(_f_permutation__round_in[1281]) );
  NAND2_X2 _f_permutation__U639  ( .A1(padder_out[258]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1949 ) );
  XNOR2_X2 _f_permutation__U638  ( .A(out[250]), .B(_f_permutation__n1949 ), 
        .ZN(_f_permutation__round_in[1282]) );
  NAND2_X2 _f_permutation__U637  ( .A1(padder_out[259]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1948 ) );
  XNOR2_X2 _f_permutation__U636  ( .A(out[251]), .B(_f_permutation__n1948 ), 
        .ZN(_f_permutation__round_in[1283]) );
  NAND2_X2 _f_permutation__U635  ( .A1(padder_out[260]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1947 ) );
  XNOR2_X2 _f_permutation__U634  ( .A(out[252]), .B(_f_permutation__n1947 ), 
        .ZN(_f_permutation__round_in[1284]) );
  NAND2_X2 _f_permutation__U633  ( .A1(padder_out[261]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1946 ) );
  XNOR2_X2 _f_permutation__U632  ( .A(out[253]), .B(_f_permutation__n1946 ), 
        .ZN(_f_permutation__round_in[1285]) );
  NAND2_X2 _f_permutation__U631  ( .A1(padder_out[262]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1945 ) );
  XNOR2_X2 _f_permutation__U630  ( .A(out[254]), .B(_f_permutation__n1945 ), 
        .ZN(_f_permutation__round_in[1286]) );
  NAND2_X2 _f_permutation__U629  ( .A1(padder_out[263]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1944 ) );
  XNOR2_X2 _f_permutation__U628  ( .A(out[255]), .B(_f_permutation__n1944 ), 
        .ZN(_f_permutation__round_in[1287]) );
  NAND2_X2 _f_permutation__U627  ( .A1(padder_out[264]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1943 ) );
  XNOR2_X2 _f_permutation__U626  ( .A(out[240]), .B(_f_permutation__n1943 ), 
        .ZN(_f_permutation__round_in[1288]) );
  NAND2_X2 _f_permutation__U625  ( .A1(padder_out[265]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1942 ) );
  XNOR2_X2 _f_permutation__U624  ( .A(out[241]), .B(_f_permutation__n1942 ), 
        .ZN(_f_permutation__round_in[1289]) );
  NAND2_X2 _f_permutation__U623  ( .A1(padder_out[266]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1941 ) );
  XNOR2_X2 _f_permutation__U622  ( .A(out[242]), .B(_f_permutation__n1941 ), 
        .ZN(_f_permutation__round_in[1290]) );
  NAND2_X2 _f_permutation__U621  ( .A1(padder_out[267]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1940 ) );
  XNOR2_X2 _f_permutation__U620  ( .A(out[243]), .B(_f_permutation__n1940 ), 
        .ZN(_f_permutation__round_in[1291]) );
  NAND2_X2 _f_permutation__U619  ( .A1(padder_out[268]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1939 ) );
  XNOR2_X2 _f_permutation__U618  ( .A(out[244]), .B(_f_permutation__n1939 ), 
        .ZN(_f_permutation__round_in[1292]) );
  NAND2_X2 _f_permutation__U617  ( .A1(padder_out[269]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1938 ) );
  XNOR2_X2 _f_permutation__U616  ( .A(out[245]), .B(_f_permutation__n1938 ), 
        .ZN(_f_permutation__round_in[1293]) );
  NAND2_X2 _f_permutation__U615  ( .A1(padder_out[270]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1937 ) );
  XNOR2_X2 _f_permutation__U614  ( .A(out[246]), .B(_f_permutation__n1937 ), 
        .ZN(_f_permutation__round_in[1294]) );
  NAND2_X2 _f_permutation__U613  ( .A1(padder_out[271]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1936 ) );
  XNOR2_X2 _f_permutation__U612  ( .A(out[247]), .B(_f_permutation__n1936 ), 
        .ZN(_f_permutation__round_in[1295]) );
  NAND2_X2 _f_permutation__U611  ( .A1(padder_out[272]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1935 ) );
  XNOR2_X2 _f_permutation__U610  ( .A(out[232]), .B(_f_permutation__n1935 ), 
        .ZN(_f_permutation__round_in[1296]) );
  NAND2_X2 _f_permutation__U609  ( .A1(padder_out[273]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1934 ) );
  XNOR2_X2 _f_permutation__U608  ( .A(out[233]), .B(_f_permutation__n1934 ), 
        .ZN(_f_permutation__round_in[1297]) );
  NAND2_X2 _f_permutation__U607  ( .A1(padder_out[274]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1933 ) );
  XNOR2_X2 _f_permutation__U606  ( .A(out[234]), .B(_f_permutation__n1933 ), 
        .ZN(_f_permutation__round_in[1298]) );
  NAND2_X2 _f_permutation__U605  ( .A1(padder_out[275]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1932 ) );
  XNOR2_X2 _f_permutation__U604  ( .A(out[235]), .B(_f_permutation__n1932 ), 
        .ZN(_f_permutation__round_in[1299]) );
  NAND2_X2 _f_permutation__U603  ( .A1(padder_out[276]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1931 ) );
  XNOR2_X2 _f_permutation__U602  ( .A(out[236]), .B(_f_permutation__n1931 ), 
        .ZN(_f_permutation__round_in[1300]) );
  NAND2_X2 _f_permutation__U601  ( .A1(padder_out[277]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1930 ) );
  XNOR2_X2 _f_permutation__U600  ( .A(out[237]), .B(_f_permutation__n1930 ), 
        .ZN(_f_permutation__round_in[1301]) );
  NAND2_X2 _f_permutation__U599  ( .A1(padder_out[278]), .A2(
        _f_permutation__n7321 ), .ZN(_f_permutation__n1929 ) );
  XNOR2_X2 _f_permutation__U598  ( .A(out[238]), .B(_f_permutation__n1929 ), 
        .ZN(_f_permutation__round_in[1302]) );
  NAND2_X2 _f_permutation__U597  ( .A1(padder_out[279]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n1928 ) );
  XNOR2_X2 _f_permutation__U596  ( .A(out[239]), .B(_f_permutation__n1928 ), 
        .ZN(_f_permutation__round_in[1303]) );
  NAND2_X2 _f_permutation__U595  ( .A1(padder_out[280]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n1927 ) );
  XNOR2_X2 _f_permutation__U594  ( .A(out[224]), .B(_f_permutation__n1927 ), 
        .ZN(_f_permutation__round_in[1304]) );
  NAND2_X2 _f_permutation__U593  ( .A1(padder_out[281]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n1926 ) );
  XNOR2_X2 _f_permutation__U592  ( .A(out[225]), .B(_f_permutation__n1926 ), 
        .ZN(_f_permutation__round_in[1305]) );
  NAND2_X2 _f_permutation__U591  ( .A1(padder_out[282]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n1925 ) );
  XNOR2_X2 _f_permutation__U590  ( .A(out[226]), .B(_f_permutation__n1925 ), 
        .ZN(_f_permutation__round_in[1306]) );
  NAND2_X2 _f_permutation__U589  ( .A1(padder_out[283]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n1924 ) );
  XNOR2_X2 _f_permutation__U588  ( .A(out[227]), .B(_f_permutation__n1924 ), 
        .ZN(_f_permutation__round_in[1307]) );
  NAND2_X2 _f_permutation__U587  ( .A1(padder_out[284]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n1923 ) );
  XNOR2_X2 _f_permutation__U586  ( .A(out[228]), .B(_f_permutation__n1923 ), 
        .ZN(_f_permutation__round_in[1308]) );
  NAND2_X2 _f_permutation__U585  ( .A1(padder_out[285]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n1922 ) );
  XNOR2_X2 _f_permutation__U584  ( .A(out[229]), .B(_f_permutation__n1922 ), 
        .ZN(_f_permutation__round_in[1309]) );
  NAND2_X2 _f_permutation__U583  ( .A1(padder_out[286]), .A2(
        _f_permutation__n7320 ), .ZN(_f_permutation__n1921 ) );
  XNOR2_X2 _f_permutation__U582  ( .A(out[230]), .B(_f_permutation__n1921 ), 
        .ZN(_f_permutation__round_in[1310]) );
  NAND2_X2 _f_permutation__U581  ( .A1(padder_out[287]), .A2(
        _f_permutation__n7322 ), .ZN(_f_permutation__n1920 ) );
  XNOR2_X2 _f_permutation__U580  ( .A(out[231]), .B(_f_permutation__n1920 ), 
        .ZN(_f_permutation__round_in[1311]) );
  NAND2_X2 _f_permutation__U579  ( .A1(padder_out[288]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1919 ) );
  XNOR2_X2 _f_permutation__U578  ( .A(out[216]), .B(_f_permutation__n1919 ), 
        .ZN(_f_permutation__round_in[1312]) );
  NAND2_X2 _f_permutation__U577  ( .A1(padder_out[289]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1918 ) );
  XNOR2_X2 _f_permutation__U576  ( .A(out[217]), .B(_f_permutation__n1918 ), 
        .ZN(_f_permutation__round_in[1313]) );
  NAND2_X2 _f_permutation__U575  ( .A1(padder_out[290]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1917 ) );
  XNOR2_X2 _f_permutation__U574  ( .A(out[218]), .B(_f_permutation__n1917 ), 
        .ZN(_f_permutation__round_in[1314]) );
  NAND2_X2 _f_permutation__U573  ( .A1(padder_out[291]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1916 ) );
  XNOR2_X2 _f_permutation__U572  ( .A(out[219]), .B(_f_permutation__n1916 ), 
        .ZN(_f_permutation__round_in[1315]) );
  NAND2_X2 _f_permutation__U571  ( .A1(padder_out[292]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1915 ) );
  XNOR2_X2 _f_permutation__U570  ( .A(out[220]), .B(_f_permutation__n1915 ), 
        .ZN(_f_permutation__round_in[1316]) );
  NAND2_X2 _f_permutation__U569  ( .A1(padder_out[293]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1914 ) );
  XNOR2_X2 _f_permutation__U568  ( .A(out[221]), .B(_f_permutation__n1914 ), 
        .ZN(_f_permutation__round_in[1317]) );
  NAND2_X2 _f_permutation__U567  ( .A1(padder_out[294]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1913 ) );
  XNOR2_X2 _f_permutation__U566  ( .A(out[222]), .B(_f_permutation__n1913 ), 
        .ZN(_f_permutation__round_in[1318]) );
  NAND2_X2 _f_permutation__U565  ( .A1(padder_out[295]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1912 ) );
  XNOR2_X2 _f_permutation__U564  ( .A(out[223]), .B(_f_permutation__n1912 ), 
        .ZN(_f_permutation__round_in[1319]) );
  NAND2_X2 _f_permutation__U563  ( .A1(padder_out[296]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1911 ) );
  XNOR2_X2 _f_permutation__U562  ( .A(out[208]), .B(_f_permutation__n1911 ), 
        .ZN(_f_permutation__round_in[1320]) );
  NAND2_X2 _f_permutation__U561  ( .A1(padder_out[297]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1910 ) );
  XNOR2_X2 _f_permutation__U560  ( .A(out[209]), .B(_f_permutation__n1910 ), 
        .ZN(_f_permutation__round_in[1321]) );
  NAND2_X2 _f_permutation__U559  ( .A1(padder_out[298]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1909 ) );
  XNOR2_X2 _f_permutation__U558  ( .A(out[210]), .B(_f_permutation__n1909 ), 
        .ZN(_f_permutation__round_in[1322]) );
  NAND2_X2 _f_permutation__U557  ( .A1(padder_out[299]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1908 ) );
  XNOR2_X2 _f_permutation__U556  ( .A(out[211]), .B(_f_permutation__n1908 ), 
        .ZN(_f_permutation__round_in[1323]) );
  NAND2_X2 _f_permutation__U555  ( .A1(padder_out[300]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1907 ) );
  XNOR2_X2 _f_permutation__U554  ( .A(out[212]), .B(_f_permutation__n1907 ), 
        .ZN(_f_permutation__round_in[1324]) );
  NAND2_X2 _f_permutation__U553  ( .A1(padder_out[301]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1906 ) );
  XNOR2_X2 _f_permutation__U552  ( .A(out[213]), .B(_f_permutation__n1906 ), 
        .ZN(_f_permutation__round_in[1325]) );
  NAND2_X2 _f_permutation__U551  ( .A1(padder_out[302]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1905 ) );
  XNOR2_X2 _f_permutation__U550  ( .A(out[214]), .B(_f_permutation__n1905 ), 
        .ZN(_f_permutation__round_in[1326]) );
  NAND2_X2 _f_permutation__U549  ( .A1(padder_out[303]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1904 ) );
  XNOR2_X2 _f_permutation__U548  ( .A(out[215]), .B(_f_permutation__n1904 ), 
        .ZN(_f_permutation__round_in[1327]) );
  NAND2_X2 _f_permutation__U547  ( .A1(padder_out[304]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1903 ) );
  XNOR2_X2 _f_permutation__U546  ( .A(out[200]), .B(_f_permutation__n1903 ), 
        .ZN(_f_permutation__round_in[1328]) );
  NAND2_X2 _f_permutation__U545  ( .A1(padder_out[305]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1902 ) );
  XNOR2_X2 _f_permutation__U544  ( .A(out[201]), .B(_f_permutation__n1902 ), 
        .ZN(_f_permutation__round_in[1329]) );
  NAND2_X2 _f_permutation__U543  ( .A1(padder_out[306]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1901 ) );
  XNOR2_X2 _f_permutation__U542  ( .A(out[202]), .B(_f_permutation__n1901 ), 
        .ZN(_f_permutation__round_in[1330]) );
  NAND2_X2 _f_permutation__U541  ( .A1(padder_out[307]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1900 ) );
  XNOR2_X2 _f_permutation__U540  ( .A(out[203]), .B(_f_permutation__n1900 ), 
        .ZN(_f_permutation__round_in[1331]) );
  NAND2_X2 _f_permutation__U539  ( .A1(padder_out[308]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1899 ) );
  XNOR2_X2 _f_permutation__U538  ( .A(out[204]), .B(_f_permutation__n1899 ), 
        .ZN(_f_permutation__round_in[1332]) );
  NAND2_X2 _f_permutation__U537  ( .A1(padder_out[309]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1898 ) );
  XNOR2_X2 _f_permutation__U536  ( .A(out[205]), .B(_f_permutation__n1898 ), 
        .ZN(_f_permutation__round_in[1333]) );
  NAND2_X2 _f_permutation__U535  ( .A1(padder_out[310]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1897 ) );
  XNOR2_X2 _f_permutation__U534  ( .A(out[206]), .B(_f_permutation__n1897 ), 
        .ZN(_f_permutation__round_in[1334]) );
  NAND2_X2 _f_permutation__U533  ( .A1(padder_out[311]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1896 ) );
  XNOR2_X2 _f_permutation__U532  ( .A(out[207]), .B(_f_permutation__n1896 ), 
        .ZN(_f_permutation__round_in[1335]) );
  NAND2_X2 _f_permutation__U531  ( .A1(padder_out[312]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1895 ) );
  XNOR2_X2 _f_permutation__U530  ( .A(out[192]), .B(_f_permutation__n1895 ), 
        .ZN(_f_permutation__round_in[1336]) );
  NAND2_X2 _f_permutation__U529  ( .A1(padder_out[313]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1894 ) );
  XNOR2_X2 _f_permutation__U528  ( .A(out[193]), .B(_f_permutation__n1894 ), 
        .ZN(_f_permutation__round_in[1337]) );
  NAND2_X2 _f_permutation__U527  ( .A1(padder_out[314]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1893 ) );
  XNOR2_X2 _f_permutation__U526  ( .A(out[194]), .B(_f_permutation__n1893 ), 
        .ZN(_f_permutation__round_in[1338]) );
  NAND2_X2 _f_permutation__U525  ( .A1(padder_out[315]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1892 ) );
  XNOR2_X2 _f_permutation__U524  ( .A(out[195]), .B(_f_permutation__n1892 ), 
        .ZN(_f_permutation__round_in[1339]) );
  NAND2_X2 _f_permutation__U523  ( .A1(padder_out[316]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1891 ) );
  XNOR2_X2 _f_permutation__U522  ( .A(out[196]), .B(_f_permutation__n1891 ), 
        .ZN(_f_permutation__round_in[1340]) );
  NAND2_X2 _f_permutation__U521  ( .A1(padder_out[317]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1890 ) );
  XNOR2_X2 _f_permutation__U520  ( .A(out[197]), .B(_f_permutation__n1890 ), 
        .ZN(_f_permutation__round_in[1341]) );
  NAND2_X2 _f_permutation__U519  ( .A1(padder_out[318]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1889 ) );
  XNOR2_X2 _f_permutation__U518  ( .A(out[198]), .B(_f_permutation__n1889 ), 
        .ZN(_f_permutation__round_in[1342]) );
  NAND2_X2 _f_permutation__U517  ( .A1(padder_out[319]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1888 ) );
  XNOR2_X2 _f_permutation__U516  ( .A(out[199]), .B(_f_permutation__n1888 ), 
        .ZN(_f_permutation__round_in[1343]) );
  NAND2_X2 _f_permutation__U515  ( .A1(padder_out[320]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1887 ) );
  XNOR2_X2 _f_permutation__U514  ( .A(out[312]), .B(_f_permutation__n1887 ), 
        .ZN(_f_permutation__round_in[1344]) );
  NAND2_X2 _f_permutation__U513  ( .A1(padder_out[321]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1886 ) );
  XNOR2_X2 _f_permutation__U512  ( .A(out[313]), .B(_f_permutation__n1886 ), 
        .ZN(_f_permutation__round_in[1345]) );
  NAND2_X2 _f_permutation__U511  ( .A1(padder_out[322]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1885 ) );
  XNOR2_X2 _f_permutation__U510  ( .A(out[314]), .B(_f_permutation__n1885 ), 
        .ZN(_f_permutation__round_in[1346]) );
  NAND2_X2 _f_permutation__U509  ( .A1(padder_out[323]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1884 ) );
  XNOR2_X2 _f_permutation__U508  ( .A(out[315]), .B(_f_permutation__n1884 ), 
        .ZN(_f_permutation__round_in[1347]) );
  NAND2_X2 _f_permutation__U507  ( .A1(padder_out[324]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1883 ) );
  XNOR2_X2 _f_permutation__U506  ( .A(out[316]), .B(_f_permutation__n1883 ), 
        .ZN(_f_permutation__round_in[1348]) );
  NAND2_X2 _f_permutation__U505  ( .A1(padder_out[325]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1882 ) );
  XNOR2_X2 _f_permutation__U504  ( .A(out[317]), .B(_f_permutation__n1882 ), 
        .ZN(_f_permutation__round_in[1349]) );
  NAND2_X2 _f_permutation__U503  ( .A1(padder_out[326]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1881 ) );
  XNOR2_X2 _f_permutation__U502  ( .A(out[318]), .B(_f_permutation__n1881 ), 
        .ZN(_f_permutation__round_in[1350]) );
  NAND2_X2 _f_permutation__U501  ( .A1(padder_out[327]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1880 ) );
  XNOR2_X2 _f_permutation__U500  ( .A(out[319]), .B(_f_permutation__n1880 ), 
        .ZN(_f_permutation__round_in[1351]) );
  NAND2_X2 _f_permutation__U499  ( .A1(padder_out[328]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1879 ) );
  XNOR2_X2 _f_permutation__U498  ( .A(out[304]), .B(_f_permutation__n1879 ), 
        .ZN(_f_permutation__round_in[1352]) );
  NAND2_X2 _f_permutation__U497  ( .A1(padder_out[329]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1878 ) );
  XNOR2_X2 _f_permutation__U496  ( .A(out[305]), .B(_f_permutation__n1878 ), 
        .ZN(_f_permutation__round_in[1353]) );
  NAND2_X2 _f_permutation__U495  ( .A1(padder_out[330]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1877 ) );
  XNOR2_X2 _f_permutation__U494  ( .A(out[306]), .B(_f_permutation__n1877 ), 
        .ZN(_f_permutation__round_in[1354]) );
  NAND2_X2 _f_permutation__U493  ( .A1(padder_out[331]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1876 ) );
  XNOR2_X2 _f_permutation__U492  ( .A(out[307]), .B(_f_permutation__n1876 ), 
        .ZN(_f_permutation__round_in[1355]) );
  NAND2_X2 _f_permutation__U491  ( .A1(padder_out[332]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1875 ) );
  XNOR2_X2 _f_permutation__U490  ( .A(out[308]), .B(_f_permutation__n1875 ), 
        .ZN(_f_permutation__round_in[1356]) );
  NAND2_X2 _f_permutation__U489  ( .A1(padder_out[333]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1874 ) );
  XNOR2_X2 _f_permutation__U488  ( .A(out[309]), .B(_f_permutation__n1874 ), 
        .ZN(_f_permutation__round_in[1357]) );
  NAND2_X2 _f_permutation__U487  ( .A1(padder_out[334]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1873 ) );
  XNOR2_X2 _f_permutation__U486  ( .A(out[310]), .B(_f_permutation__n1873 ), 
        .ZN(_f_permutation__round_in[1358]) );
  NAND2_X2 _f_permutation__U485  ( .A1(padder_out[335]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1872 ) );
  XNOR2_X2 _f_permutation__U484  ( .A(out[311]), .B(_f_permutation__n1872 ), 
        .ZN(_f_permutation__round_in[1359]) );
  NAND2_X2 _f_permutation__U483  ( .A1(padder_out[336]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1871 ) );
  XNOR2_X2 _f_permutation__U482  ( .A(out[296]), .B(_f_permutation__n1871 ), 
        .ZN(_f_permutation__round_in[1360]) );
  NAND2_X2 _f_permutation__U481  ( .A1(padder_out[337]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1870 ) );
  XNOR2_X2 _f_permutation__U480  ( .A(out[297]), .B(_f_permutation__n1870 ), 
        .ZN(_f_permutation__round_in[1361]) );
  NAND2_X2 _f_permutation__U479  ( .A1(padder_out[338]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1869 ) );
  XNOR2_X2 _f_permutation__U478  ( .A(out[298]), .B(_f_permutation__n1869 ), 
        .ZN(_f_permutation__round_in[1362]) );
  NAND2_X2 _f_permutation__U477  ( .A1(padder_out[339]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1868 ) );
  XNOR2_X2 _f_permutation__U476  ( .A(out[299]), .B(_f_permutation__n1868 ), 
        .ZN(_f_permutation__round_in[1363]) );
  NAND2_X2 _f_permutation__U475  ( .A1(padder_out[340]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1867 ) );
  XNOR2_X2 _f_permutation__U474  ( .A(out[300]), .B(_f_permutation__n1867 ), 
        .ZN(_f_permutation__round_in[1364]) );
  NAND2_X2 _f_permutation__U473  ( .A1(padder_out[341]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1866 ) );
  XNOR2_X2 _f_permutation__U472  ( .A(out[301]), .B(_f_permutation__n1866 ), 
        .ZN(_f_permutation__round_in[1365]) );
  NAND2_X2 _f_permutation__U471  ( .A1(padder_out[342]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1865 ) );
  XNOR2_X2 _f_permutation__U470  ( .A(out[302]), .B(_f_permutation__n1865 ), 
        .ZN(_f_permutation__round_in[1366]) );
  NAND2_X2 _f_permutation__U469  ( .A1(padder_out[343]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1864 ) );
  XNOR2_X2 _f_permutation__U468  ( .A(out[303]), .B(_f_permutation__n1864 ), 
        .ZN(_f_permutation__round_in[1367]) );
  NAND2_X2 _f_permutation__U467  ( .A1(padder_out[344]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1863 ) );
  XNOR2_X2 _f_permutation__U466  ( .A(out[288]), .B(_f_permutation__n1863 ), 
        .ZN(_f_permutation__round_in[1368]) );
  NAND2_X2 _f_permutation__U465  ( .A1(padder_out[345]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1862 ) );
  XNOR2_X2 _f_permutation__U464  ( .A(out[289]), .B(_f_permutation__n1862 ), 
        .ZN(_f_permutation__round_in[1369]) );
  NAND2_X2 _f_permutation__U463  ( .A1(padder_out[346]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1861 ) );
  XNOR2_X2 _f_permutation__U462  ( .A(out[290]), .B(_f_permutation__n1861 ), 
        .ZN(_f_permutation__round_in[1370]) );
  NAND2_X2 _f_permutation__U461  ( .A1(padder_out[347]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1860 ) );
  XNOR2_X2 _f_permutation__U460  ( .A(out[291]), .B(_f_permutation__n1860 ), 
        .ZN(_f_permutation__round_in[1371]) );
  NAND2_X2 _f_permutation__U459  ( .A1(padder_out[348]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1859 ) );
  XNOR2_X2 _f_permutation__U458  ( .A(out[292]), .B(_f_permutation__n1859 ), 
        .ZN(_f_permutation__round_in[1372]) );
  NAND2_X2 _f_permutation__U457  ( .A1(padder_out[349]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1858 ) );
  XNOR2_X2 _f_permutation__U456  ( .A(out[293]), .B(_f_permutation__n1858 ), 
        .ZN(_f_permutation__round_in[1373]) );
  NAND2_X2 _f_permutation__U455  ( .A1(padder_out[350]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1857 ) );
  XNOR2_X2 _f_permutation__U454  ( .A(out[294]), .B(_f_permutation__n1857 ), 
        .ZN(_f_permutation__round_in[1374]) );
  NAND2_X2 _f_permutation__U453  ( .A1(padder_out[351]), .A2(
        _f_permutation__n7313 ), .ZN(_f_permutation__n1856 ) );
  XNOR2_X2 _f_permutation__U452  ( .A(out[295]), .B(_f_permutation__n1856 ), 
        .ZN(_f_permutation__round_in[1375]) );
  NAND2_X2 _f_permutation__U451  ( .A1(padder_out[352]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1855 ) );
  XNOR2_X2 _f_permutation__U450  ( .A(out[280]), .B(_f_permutation__n1855 ), 
        .ZN(_f_permutation__round_in[1376]) );
  NAND2_X2 _f_permutation__U449  ( .A1(padder_out[353]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1854 ) );
  XNOR2_X2 _f_permutation__U448  ( .A(out[281]), .B(_f_permutation__n1854 ), 
        .ZN(_f_permutation__round_in[1377]) );
  NAND2_X2 _f_permutation__U447  ( .A1(padder_out[354]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1853 ) );
  XNOR2_X2 _f_permutation__U446  ( .A(out[282]), .B(_f_permutation__n1853 ), 
        .ZN(_f_permutation__round_in[1378]) );
  NAND2_X2 _f_permutation__U445  ( .A1(padder_out[355]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1852 ) );
  XNOR2_X2 _f_permutation__U444  ( .A(out[283]), .B(_f_permutation__n1852 ), 
        .ZN(_f_permutation__round_in[1379]) );
  NAND2_X2 _f_permutation__U443  ( .A1(padder_out[356]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1851 ) );
  XNOR2_X2 _f_permutation__U442  ( .A(out[284]), .B(_f_permutation__n1851 ), 
        .ZN(_f_permutation__round_in[1380]) );
  NAND2_X2 _f_permutation__U441  ( .A1(padder_out[357]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1850 ) );
  XNOR2_X2 _f_permutation__U440  ( .A(out[285]), .B(_f_permutation__n1850 ), 
        .ZN(_f_permutation__round_in[1381]) );
  NAND2_X2 _f_permutation__U439  ( .A1(padder_out[358]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1849 ) );
  XNOR2_X2 _f_permutation__U438  ( .A(out[286]), .B(_f_permutation__n1849 ), 
        .ZN(_f_permutation__round_in[1382]) );
  NAND2_X2 _f_permutation__U437  ( .A1(padder_out[359]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1848 ) );
  XNOR2_X2 _f_permutation__U436  ( .A(out[287]), .B(_f_permutation__n1848 ), 
        .ZN(_f_permutation__round_in[1383]) );
  NAND2_X2 _f_permutation__U435  ( .A1(padder_out[360]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1847 ) );
  XNOR2_X2 _f_permutation__U434  ( .A(out[272]), .B(_f_permutation__n1847 ), 
        .ZN(_f_permutation__round_in[1384]) );
  NAND2_X2 _f_permutation__U433  ( .A1(padder_out[361]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1846 ) );
  XNOR2_X2 _f_permutation__U432  ( .A(out[273]), .B(_f_permutation__n1846 ), 
        .ZN(_f_permutation__round_in[1385]) );
  NAND2_X2 _f_permutation__U431  ( .A1(padder_out[362]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1845 ) );
  XNOR2_X2 _f_permutation__U430  ( .A(out[274]), .B(_f_permutation__n1845 ), 
        .ZN(_f_permutation__round_in[1386]) );
  NAND2_X2 _f_permutation__U429  ( .A1(padder_out[363]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1844 ) );
  XNOR2_X2 _f_permutation__U428  ( .A(out[275]), .B(_f_permutation__n1844 ), 
        .ZN(_f_permutation__round_in[1387]) );
  NAND2_X2 _f_permutation__U427  ( .A1(padder_out[364]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1843 ) );
  XNOR2_X2 _f_permutation__U426  ( .A(out[276]), .B(_f_permutation__n1843 ), 
        .ZN(_f_permutation__round_in[1388]) );
  NAND2_X2 _f_permutation__U425  ( .A1(padder_out[365]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1842 ) );
  XNOR2_X2 _f_permutation__U424  ( .A(out[277]), .B(_f_permutation__n1842 ), 
        .ZN(_f_permutation__round_in[1389]) );
  NAND2_X2 _f_permutation__U423  ( .A1(padder_out[366]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1841 ) );
  XNOR2_X2 _f_permutation__U422  ( .A(out[278]), .B(_f_permutation__n1841 ), 
        .ZN(_f_permutation__round_in[1390]) );
  NAND2_X2 _f_permutation__U421  ( .A1(padder_out[367]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1840 ) );
  XNOR2_X2 _f_permutation__U420  ( .A(out[279]), .B(_f_permutation__n1840 ), 
        .ZN(_f_permutation__round_in[1391]) );
  NAND2_X2 _f_permutation__U419  ( .A1(padder_out[368]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1839 ) );
  XNOR2_X2 _f_permutation__U418  ( .A(out[264]), .B(_f_permutation__n1839 ), 
        .ZN(_f_permutation__round_in[1392]) );
  NAND2_X2 _f_permutation__U417  ( .A1(padder_out[369]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1838 ) );
  XNOR2_X2 _f_permutation__U416  ( .A(out[265]), .B(_f_permutation__n1838 ), 
        .ZN(_f_permutation__round_in[1393]) );
  NAND2_X2 _f_permutation__U415  ( .A1(padder_out[370]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1837 ) );
  XNOR2_X2 _f_permutation__U414  ( .A(out[266]), .B(_f_permutation__n1837 ), 
        .ZN(_f_permutation__round_in[1394]) );
  NAND2_X2 _f_permutation__U413  ( .A1(padder_out[371]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1836 ) );
  XNOR2_X2 _f_permutation__U412  ( .A(out[267]), .B(_f_permutation__n1836 ), 
        .ZN(_f_permutation__round_in[1395]) );
  NAND2_X2 _f_permutation__U411  ( .A1(padder_out[372]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1835 ) );
  XNOR2_X2 _f_permutation__U410  ( .A(out[268]), .B(_f_permutation__n1835 ), 
        .ZN(_f_permutation__round_in[1396]) );
  NAND2_X2 _f_permutation__U409  ( .A1(padder_out[373]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1834 ) );
  XNOR2_X2 _f_permutation__U408  ( .A(out[269]), .B(_f_permutation__n1834 ), 
        .ZN(_f_permutation__round_in[1397]) );
  NAND2_X2 _f_permutation__U407  ( .A1(padder_out[374]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1833 ) );
  XNOR2_X2 _f_permutation__U406  ( .A(out[270]), .B(_f_permutation__n1833 ), 
        .ZN(_f_permutation__round_in[1398]) );
  NAND2_X2 _f_permutation__U405  ( .A1(padder_out[375]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1832 ) );
  XNOR2_X2 _f_permutation__U404  ( .A(out[271]), .B(_f_permutation__n1832 ), 
        .ZN(_f_permutation__round_in[1399]) );
  NAND2_X2 _f_permutation__U403  ( .A1(padder_out[376]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1831 ) );
  XNOR2_X2 _f_permutation__U402  ( .A(out[256]), .B(_f_permutation__n1831 ), 
        .ZN(_f_permutation__round_in[1400]) );
  NAND2_X2 _f_permutation__U401  ( .A1(padder_out[377]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1830 ) );
  XNOR2_X2 _f_permutation__U400  ( .A(out[257]), .B(_f_permutation__n1830 ), 
        .ZN(_f_permutation__round_in[1401]) );
  NAND2_X2 _f_permutation__U399  ( .A1(padder_out[378]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1829 ) );
  XNOR2_X2 _f_permutation__U398  ( .A(out[258]), .B(_f_permutation__n1829 ), 
        .ZN(_f_permutation__round_in[1402]) );
  NAND2_X2 _f_permutation__U397  ( .A1(padder_out[379]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1828 ) );
  XNOR2_X2 _f_permutation__U395  ( .A(out[259]), .B(_f_permutation__n1828 ), 
        .ZN(_f_permutation__round_in[1403]) );
  NAND2_X2 _f_permutation__U394  ( .A1(padder_out[380]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1827 ) );
  XNOR2_X2 _f_permutation__U393  ( .A(out[260]), .B(_f_permutation__n1827 ), 
        .ZN(_f_permutation__round_in[1404]) );
  NAND2_X2 _f_permutation__U392  ( .A1(padder_out[381]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1826 ) );
  XNOR2_X2 _f_permutation__U391  ( .A(out[261]), .B(_f_permutation__n1826 ), 
        .ZN(_f_permutation__round_in[1405]) );
  NAND2_X2 _f_permutation__U390  ( .A1(padder_out[382]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1825 ) );
  XNOR2_X2 _f_permutation__U389  ( .A(out[262]), .B(_f_permutation__n1825 ), 
        .ZN(_f_permutation__round_in[1406]) );
  NAND2_X2 _f_permutation__U388  ( .A1(padder_out[383]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1824 ) );
  XNOR2_X2 _f_permutation__U387  ( .A(out[263]), .B(_f_permutation__n1824 ), 
        .ZN(_f_permutation__round_in[1407]) );
  NAND2_X2 _f_permutation__U386  ( .A1(padder_out[384]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1823 ) );
  XNOR2_X2 _f_permutation__U385  ( .A(out[376]), .B(_f_permutation__n1823 ), 
        .ZN(_f_permutation__round_in[1408]) );
  NAND2_X2 _f_permutation__U384  ( .A1(padder_out[385]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1822 ) );
  XNOR2_X2 _f_permutation__U383  ( .A(out[377]), .B(_f_permutation__n1822 ), 
        .ZN(_f_permutation__round_in[1409]) );
  NAND2_X2 _f_permutation__U382  ( .A1(padder_out[386]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1821 ) );
  XNOR2_X2 _f_permutation__U381  ( .A(out[378]), .B(_f_permutation__n1821 ), 
        .ZN(_f_permutation__round_in[1410]) );
  NAND2_X2 _f_permutation__U380  ( .A1(padder_out[387]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1820 ) );
  XNOR2_X2 _f_permutation__U379  ( .A(out[379]), .B(_f_permutation__n1820 ), 
        .ZN(_f_permutation__round_in[1411]) );
  NAND2_X2 _f_permutation__U378  ( .A1(padder_out[388]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1819 ) );
  XNOR2_X2 _f_permutation__U377  ( .A(out[380]), .B(_f_permutation__n1819 ), 
        .ZN(_f_permutation__round_in[1412]) );
  NAND2_X2 _f_permutation__U376  ( .A1(padder_out[389]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1818 ) );
  XNOR2_X2 _f_permutation__U375  ( .A(out[381]), .B(_f_permutation__n1818 ), 
        .ZN(_f_permutation__round_in[1413]) );
  NAND2_X2 _f_permutation__U374  ( .A1(padder_out[390]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1817 ) );
  XNOR2_X2 _f_permutation__U373  ( .A(out[382]), .B(_f_permutation__n1817 ), 
        .ZN(_f_permutation__round_in[1414]) );
  NAND2_X2 _f_permutation__U372  ( .A1(padder_out[391]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1816 ) );
  XNOR2_X2 _f_permutation__U371  ( .A(out[383]), .B(_f_permutation__n1816 ), 
        .ZN(_f_permutation__round_in[1415]) );
  NAND2_X2 _f_permutation__U370  ( .A1(padder_out[392]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1815 ) );
  XNOR2_X2 _f_permutation__U369  ( .A(out[368]), .B(_f_permutation__n1815 ), 
        .ZN(_f_permutation__round_in[1416]) );
  NAND2_X2 _f_permutation__U368  ( .A1(padder_out[393]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1814 ) );
  XNOR2_X2 _f_permutation__U367  ( .A(out[369]), .B(_f_permutation__n1814 ), 
        .ZN(_f_permutation__round_in[1417]) );
  NAND2_X2 _f_permutation__U366  ( .A1(padder_out[394]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1813 ) );
  XNOR2_X2 _f_permutation__U365  ( .A(out[370]), .B(_f_permutation__n1813 ), 
        .ZN(_f_permutation__round_in[1418]) );
  NAND2_X2 _f_permutation__U364  ( .A1(padder_out[395]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1812 ) );
  XNOR2_X2 _f_permutation__U363  ( .A(out[371]), .B(_f_permutation__n1812 ), 
        .ZN(_f_permutation__round_in[1419]) );
  NAND2_X2 _f_permutation__U362  ( .A1(padder_out[396]), .A2(f_ack), .ZN(
        _f_permutation__n1811 ) );
  XNOR2_X2 _f_permutation__U361  ( .A(out[372]), .B(_f_permutation__n1811 ), 
        .ZN(_f_permutation__round_in[1420]) );
  NAND2_X2 _f_permutation__U360  ( .A1(padder_out[397]), .A2(f_ack), .ZN(
        _f_permutation__n1810 ) );
  XNOR2_X2 _f_permutation__U359  ( .A(out[373]), .B(_f_permutation__n1810 ), 
        .ZN(_f_permutation__round_in[1421]) );
  NAND2_X2 _f_permutation__U358  ( .A1(padder_out[398]), .A2(f_ack), .ZN(
        _f_permutation__n1809 ) );
  XNOR2_X2 _f_permutation__U357  ( .A(out[374]), .B(_f_permutation__n1809 ), 
        .ZN(_f_permutation__round_in[1422]) );
  NAND2_X2 _f_permutation__U356  ( .A1(padder_out[399]), .A2(f_ack), .ZN(
        _f_permutation__n1808 ) );
  XNOR2_X2 _f_permutation__U355  ( .A(out[375]), .B(_f_permutation__n1808 ), 
        .ZN(_f_permutation__round_in[1423]) );
  NAND2_X2 _f_permutation__U354  ( .A1(padder_out[400]), .A2(f_ack), .ZN(
        _f_permutation__n1807 ) );
  XNOR2_X2 _f_permutation__U353  ( .A(out[360]), .B(_f_permutation__n1807 ), 
        .ZN(_f_permutation__round_in[1424]) );
  NAND2_X2 _f_permutation__U352  ( .A1(padder_out[401]), .A2(f_ack), .ZN(
        _f_permutation__n1806 ) );
  XNOR2_X2 _f_permutation__U351  ( .A(out[361]), .B(_f_permutation__n1806 ), 
        .ZN(_f_permutation__round_in[1425]) );
  NAND2_X2 _f_permutation__U350  ( .A1(padder_out[402]), .A2(f_ack), .ZN(
        _f_permutation__n1805 ) );
  XNOR2_X2 _f_permutation__U349  ( .A(out[362]), .B(_f_permutation__n1805 ), 
        .ZN(_f_permutation__round_in[1426]) );
  NAND2_X2 _f_permutation__U348  ( .A1(padder_out[403]), .A2(f_ack), .ZN(
        _f_permutation__n1804 ) );
  XNOR2_X2 _f_permutation__U347  ( .A(out[363]), .B(_f_permutation__n1804 ), 
        .ZN(_f_permutation__round_in[1427]) );
  NAND2_X2 _f_permutation__U346  ( .A1(padder_out[404]), .A2(f_ack), .ZN(
        _f_permutation__n1803 ) );
  XNOR2_X2 _f_permutation__U345  ( .A(out[364]), .B(_f_permutation__n1803 ), 
        .ZN(_f_permutation__round_in[1428]) );
  NAND2_X2 _f_permutation__U344  ( .A1(padder_out[405]), .A2(f_ack), .ZN(
        _f_permutation__n1802 ) );
  XNOR2_X2 _f_permutation__U343  ( .A(out[365]), .B(_f_permutation__n1802 ), 
        .ZN(_f_permutation__round_in[1429]) );
  NAND2_X2 _f_permutation__U342  ( .A1(padder_out[406]), .A2(f_ack), .ZN(
        _f_permutation__n1801 ) );
  XNOR2_X2 _f_permutation__U341  ( .A(out[366]), .B(_f_permutation__n1801 ), 
        .ZN(_f_permutation__round_in[1430]) );
  NAND2_X2 _f_permutation__U340  ( .A1(padder_out[407]), .A2(f_ack), .ZN(
        _f_permutation__n1800 ) );
  XNOR2_X2 _f_permutation__U339  ( .A(out[367]), .B(_f_permutation__n1800 ), 
        .ZN(_f_permutation__round_in[1431]) );
  NAND2_X2 _f_permutation__U338  ( .A1(padder_out[408]), .A2(f_ack), .ZN(
        _f_permutation__n1799 ) );
  XNOR2_X2 _f_permutation__U337  ( .A(out[352]), .B(_f_permutation__n1799 ), 
        .ZN(_f_permutation__round_in[1432]) );
  NAND2_X2 _f_permutation__U336  ( .A1(padder_out[409]), .A2(f_ack), .ZN(
        _f_permutation__n1798 ) );
  XNOR2_X2 _f_permutation__U335  ( .A(out[353]), .B(_f_permutation__n1798 ), 
        .ZN(_f_permutation__round_in[1433]) );
  NAND2_X2 _f_permutation__U334  ( .A1(padder_out[410]), .A2(f_ack), .ZN(
        _f_permutation__n1797 ) );
  XNOR2_X2 _f_permutation__U333  ( .A(out[354]), .B(_f_permutation__n1797 ), 
        .ZN(_f_permutation__round_in[1434]) );
  NAND2_X2 _f_permutation__U332  ( .A1(padder_out[411]), .A2(f_ack), .ZN(
        _f_permutation__n1796 ) );
  XNOR2_X2 _f_permutation__U331  ( .A(out[355]), .B(_f_permutation__n1796 ), 
        .ZN(_f_permutation__round_in[1435]) );
  NAND2_X2 _f_permutation__U330  ( .A1(padder_out[412]), .A2(f_ack), .ZN(
        _f_permutation__n1795 ) );
  XNOR2_X2 _f_permutation__U329  ( .A(out[356]), .B(_f_permutation__n1795 ), 
        .ZN(_f_permutation__round_in[1436]) );
  NAND2_X2 _f_permutation__U328  ( .A1(padder_out[413]), .A2(f_ack), .ZN(
        _f_permutation__n1794 ) );
  XNOR2_X2 _f_permutation__U327  ( .A(out[357]), .B(_f_permutation__n1794 ), 
        .ZN(_f_permutation__round_in[1437]) );
  NAND2_X2 _f_permutation__U326  ( .A1(padder_out[414]), .A2(f_ack), .ZN(
        _f_permutation__n1793 ) );
  XNOR2_X2 _f_permutation__U325  ( .A(out[358]), .B(_f_permutation__n1793 ), 
        .ZN(_f_permutation__round_in[1438]) );
  NAND2_X2 _f_permutation__U324  ( .A1(padder_out[415]), .A2(f_ack), .ZN(
        _f_permutation__n1792 ) );
  XNOR2_X2 _f_permutation__U323  ( .A(out[359]), .B(_f_permutation__n1792 ), 
        .ZN(_f_permutation__round_in[1439]) );
  NAND2_X2 _f_permutation__U322  ( .A1(padder_out[416]), .A2(f_ack), .ZN(
        _f_permutation__n1791 ) );
  XNOR2_X2 _f_permutation__U321  ( .A(out[344]), .B(_f_permutation__n1791 ), 
        .ZN(_f_permutation__round_in[1440]) );
  NAND2_X2 _f_permutation__U320  ( .A1(padder_out[417]), .A2(f_ack), .ZN(
        _f_permutation__n1790 ) );
  XNOR2_X2 _f_permutation__U319  ( .A(out[345]), .B(_f_permutation__n1790 ), 
        .ZN(_f_permutation__round_in[1441]) );
  NAND2_X2 _f_permutation__U318  ( .A1(padder_out[418]), .A2(f_ack), .ZN(
        _f_permutation__n1789 ) );
  XNOR2_X2 _f_permutation__U317  ( .A(out[346]), .B(_f_permutation__n1789 ), 
        .ZN(_f_permutation__round_in[1442]) );
  NAND2_X2 _f_permutation__U316  ( .A1(padder_out[419]), .A2(f_ack), .ZN(
        _f_permutation__n1788 ) );
  XNOR2_X2 _f_permutation__U315  ( .A(out[347]), .B(_f_permutation__n1788 ), 
        .ZN(_f_permutation__round_in[1443]) );
  NAND2_X2 _f_permutation__U314  ( .A1(padder_out[420]), .A2(f_ack), .ZN(
        _f_permutation__n1787 ) );
  XNOR2_X2 _f_permutation__U313  ( .A(out[348]), .B(_f_permutation__n1787 ), 
        .ZN(_f_permutation__round_in[1444]) );
  NAND2_X2 _f_permutation__U312  ( .A1(padder_out[421]), .A2(f_ack), .ZN(
        _f_permutation__n1786 ) );
  XNOR2_X2 _f_permutation__U311  ( .A(out[349]), .B(_f_permutation__n1786 ), 
        .ZN(_f_permutation__round_in[1445]) );
  NAND2_X2 _f_permutation__U310  ( .A1(padder_out[422]), .A2(f_ack), .ZN(
        _f_permutation__n1785 ) );
  XNOR2_X2 _f_permutation__U309  ( .A(out[350]), .B(_f_permutation__n1785 ), 
        .ZN(_f_permutation__round_in[1446]) );
  NAND2_X2 _f_permutation__U308  ( .A1(padder_out[423]), .A2(f_ack), .ZN(
        _f_permutation__n1784 ) );
  XNOR2_X2 _f_permutation__U307  ( .A(out[351]), .B(_f_permutation__n1784 ), 
        .ZN(_f_permutation__round_in[1447]) );
  NAND2_X2 _f_permutation__U306  ( .A1(padder_out[424]), .A2(f_ack), .ZN(
        _f_permutation__n1783 ) );
  XNOR2_X2 _f_permutation__U305  ( .A(out[336]), .B(_f_permutation__n1783 ), 
        .ZN(_f_permutation__round_in[1448]) );
  NAND2_X2 _f_permutation__U304  ( .A1(padder_out[425]), .A2(f_ack), .ZN(
        _f_permutation__n1782 ) );
  XNOR2_X2 _f_permutation__U303  ( .A(out[337]), .B(_f_permutation__n1782 ), 
        .ZN(_f_permutation__round_in[1449]) );
  NAND2_X2 _f_permutation__U302  ( .A1(padder_out[426]), .A2(f_ack), .ZN(
        _f_permutation__n1781 ) );
  XNOR2_X2 _f_permutation__U301  ( .A(out[338]), .B(_f_permutation__n1781 ), 
        .ZN(_f_permutation__round_in[1450]) );
  NAND2_X2 _f_permutation__U300  ( .A1(padder_out[427]), .A2(f_ack), .ZN(
        _f_permutation__n1780 ) );
  XNOR2_X2 _f_permutation__U299  ( .A(out[339]), .B(_f_permutation__n1780 ), 
        .ZN(_f_permutation__round_in[1451]) );
  NAND2_X2 _f_permutation__U298  ( .A1(padder_out[428]), .A2(f_ack), .ZN(
        _f_permutation__n1779 ) );
  XNOR2_X2 _f_permutation__U297  ( .A(out[340]), .B(_f_permutation__n1779 ), 
        .ZN(_f_permutation__round_in[1452]) );
  NAND2_X2 _f_permutation__U296  ( .A1(padder_out[429]), .A2(f_ack), .ZN(
        _f_permutation__n1778 ) );
  XNOR2_X2 _f_permutation__U295  ( .A(out[341]), .B(_f_permutation__n1778 ), 
        .ZN(_f_permutation__round_in[1453]) );
  NAND2_X2 _f_permutation__U294  ( .A1(padder_out[430]), .A2(f_ack), .ZN(
        _f_permutation__n1777 ) );
  XNOR2_X2 _f_permutation__U293  ( .A(out[342]), .B(_f_permutation__n1777 ), 
        .ZN(_f_permutation__round_in[1454]) );
  NAND2_X2 _f_permutation__U292  ( .A1(padder_out[431]), .A2(
        _f_permutation__n7312 ), .ZN(_f_permutation__n1776 ) );
  XNOR2_X2 _f_permutation__U291  ( .A(out[343]), .B(_f_permutation__n1776 ), 
        .ZN(_f_permutation__round_in[1455]) );
  NAND2_X2 _f_permutation__U290  ( .A1(padder_out[432]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1775 ) );
  XNOR2_X2 _f_permutation__U289  ( .A(out[328]), .B(_f_permutation__n1775 ), 
        .ZN(_f_permutation__round_in[1456]) );
  NAND2_X2 _f_permutation__U288  ( .A1(padder_out[433]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1774 ) );
  XNOR2_X2 _f_permutation__U287  ( .A(out[329]), .B(_f_permutation__n1774 ), 
        .ZN(_f_permutation__round_in[1457]) );
  NAND2_X2 _f_permutation__U286  ( .A1(padder_out[434]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1773 ) );
  XNOR2_X2 _f_permutation__U285  ( .A(out[330]), .B(_f_permutation__n1773 ), 
        .ZN(_f_permutation__round_in[1458]) );
  NAND2_X2 _f_permutation__U284  ( .A1(padder_out[435]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1772 ) );
  XNOR2_X2 _f_permutation__U283  ( .A(out[331]), .B(_f_permutation__n1772 ), 
        .ZN(_f_permutation__round_in[1459]) );
  NAND2_X2 _f_permutation__U282  ( .A1(padder_out[436]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1771 ) );
  XNOR2_X2 _f_permutation__U281  ( .A(out[332]), .B(_f_permutation__n1771 ), 
        .ZN(_f_permutation__round_in[1460]) );
  NAND2_X2 _f_permutation__U280  ( .A1(padder_out[437]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1770 ) );
  XNOR2_X2 _f_permutation__U279  ( .A(out[333]), .B(_f_permutation__n1770 ), 
        .ZN(_f_permutation__round_in[1461]) );
  NAND2_X2 _f_permutation__U278  ( .A1(padder_out[438]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1769 ) );
  XNOR2_X2 _f_permutation__U277  ( .A(out[334]), .B(_f_permutation__n1769 ), 
        .ZN(_f_permutation__round_in[1462]) );
  NAND2_X2 _f_permutation__U276  ( .A1(padder_out[439]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1768 ) );
  XNOR2_X2 _f_permutation__U275  ( .A(out[335]), .B(_f_permutation__n1768 ), 
        .ZN(_f_permutation__round_in[1463]) );
  NAND2_X2 _f_permutation__U274  ( .A1(padder_out[440]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1767 ) );
  XNOR2_X2 _f_permutation__U273  ( .A(out[320]), .B(_f_permutation__n1767 ), 
        .ZN(_f_permutation__round_in[1464]) );
  NAND2_X2 _f_permutation__U272  ( .A1(padder_out[441]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1766 ) );
  XNOR2_X2 _f_permutation__U271  ( .A(out[321]), .B(_f_permutation__n1766 ), 
        .ZN(_f_permutation__round_in[1465]) );
  NAND2_X2 _f_permutation__U270  ( .A1(padder_out[442]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1765 ) );
  XNOR2_X2 _f_permutation__U269  ( .A(out[322]), .B(_f_permutation__n1765 ), 
        .ZN(_f_permutation__round_in[1466]) );
  NAND2_X2 _f_permutation__U268  ( .A1(padder_out[443]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1764 ) );
  XNOR2_X2 _f_permutation__U267  ( .A(out[323]), .B(_f_permutation__n1764 ), 
        .ZN(_f_permutation__round_in[1467]) );
  NAND2_X2 _f_permutation__U266  ( .A1(padder_out[444]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1763 ) );
  XNOR2_X2 _f_permutation__U265  ( .A(out[324]), .B(_f_permutation__n1763 ), 
        .ZN(_f_permutation__round_in[1468]) );
  NAND2_X2 _f_permutation__U264  ( .A1(padder_out[445]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1762 ) );
  XNOR2_X2 _f_permutation__U263  ( .A(out[325]), .B(_f_permutation__n1762 ), 
        .ZN(_f_permutation__round_in[1469]) );
  NAND2_X2 _f_permutation__U262  ( .A1(padder_out[446]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1761 ) );
  XNOR2_X2 _f_permutation__U261  ( .A(out[326]), .B(_f_permutation__n1761 ), 
        .ZN(_f_permutation__round_in[1470]) );
  NAND2_X2 _f_permutation__U260  ( .A1(padder_out[447]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1760 ) );
  XNOR2_X2 _f_permutation__U259  ( .A(out[327]), .B(_f_permutation__n1760 ), 
        .ZN(_f_permutation__round_in[1471]) );
  NAND2_X2 _f_permutation__U258  ( .A1(padder_out[448]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1759 ) );
  XNOR2_X2 _f_permutation__U257  ( .A(out[440]), .B(_f_permutation__n1759 ), 
        .ZN(_f_permutation__round_in[1472]) );
  NAND2_X2 _f_permutation__U256  ( .A1(padder_out[449]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1758 ) );
  XNOR2_X2 _f_permutation__U255  ( .A(out[441]), .B(_f_permutation__n1758 ), 
        .ZN(_f_permutation__round_in[1473]) );
  NAND2_X2 _f_permutation__U254  ( .A1(padder_out[450]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1757 ) );
  XNOR2_X2 _f_permutation__U253  ( .A(out[442]), .B(_f_permutation__n1757 ), 
        .ZN(_f_permutation__round_in[1474]) );
  NAND2_X2 _f_permutation__U252  ( .A1(padder_out[451]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1756 ) );
  XNOR2_X2 _f_permutation__U251  ( .A(out[443]), .B(_f_permutation__n1756 ), 
        .ZN(_f_permutation__round_in[1475]) );
  NAND2_X2 _f_permutation__U250  ( .A1(padder_out[452]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1755 ) );
  XNOR2_X2 _f_permutation__U249  ( .A(out[444]), .B(_f_permutation__n1755 ), 
        .ZN(_f_permutation__round_in[1476]) );
  NAND2_X2 _f_permutation__U248  ( .A1(padder_out[453]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1754 ) );
  XNOR2_X2 _f_permutation__U247  ( .A(out[445]), .B(_f_permutation__n1754 ), 
        .ZN(_f_permutation__round_in[1477]) );
  NAND2_X2 _f_permutation__U246  ( .A1(padder_out[454]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1753 ) );
  XNOR2_X2 _f_permutation__U245  ( .A(out[446]), .B(_f_permutation__n1753 ), 
        .ZN(_f_permutation__round_in[1478]) );
  NAND2_X2 _f_permutation__U244  ( .A1(padder_out[455]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1752 ) );
  XNOR2_X2 _f_permutation__U243  ( .A(out[447]), .B(_f_permutation__n1752 ), 
        .ZN(_f_permutation__round_in[1479]) );
  NAND2_X2 _f_permutation__U242  ( .A1(padder_out[456]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1751 ) );
  XNOR2_X2 _f_permutation__U241  ( .A(out[432]), .B(_f_permutation__n1751 ), 
        .ZN(_f_permutation__round_in[1480]) );
  NAND2_X2 _f_permutation__U240  ( .A1(padder_out[457]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1750 ) );
  XNOR2_X2 _f_permutation__U239  ( .A(out[433]), .B(_f_permutation__n1750 ), 
        .ZN(_f_permutation__round_in[1481]) );
  NAND2_X2 _f_permutation__U238  ( .A1(padder_out[458]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1749 ) );
  XNOR2_X2 _f_permutation__U237  ( .A(out[434]), .B(_f_permutation__n1749 ), 
        .ZN(_f_permutation__round_in[1482]) );
  NAND2_X2 _f_permutation__U236  ( .A1(padder_out[459]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1748 ) );
  XNOR2_X2 _f_permutation__U235  ( .A(out[435]), .B(_f_permutation__n1748 ), 
        .ZN(_f_permutation__round_in[1483]) );
  NAND2_X2 _f_permutation__U234  ( .A1(padder_out[460]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1747 ) );
  XNOR2_X2 _f_permutation__U233  ( .A(out[436]), .B(_f_permutation__n1747 ), 
        .ZN(_f_permutation__round_in[1484]) );
  NAND2_X2 _f_permutation__U232  ( .A1(padder_out[461]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1746 ) );
  XNOR2_X2 _f_permutation__U231  ( .A(out[437]), .B(_f_permutation__n1746 ), 
        .ZN(_f_permutation__round_in[1485]) );
  NAND2_X2 _f_permutation__U230  ( .A1(padder_out[462]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1745 ) );
  XNOR2_X2 _f_permutation__U229  ( .A(out[438]), .B(_f_permutation__n1745 ), 
        .ZN(_f_permutation__round_in[1486]) );
  NAND2_X2 _f_permutation__U228  ( .A1(padder_out[463]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1744 ) );
  XNOR2_X2 _f_permutation__U227  ( .A(out[439]), .B(_f_permutation__n1744 ), 
        .ZN(_f_permutation__round_in[1487]) );
  NAND2_X2 _f_permutation__U226  ( .A1(padder_out[464]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1743 ) );
  XNOR2_X2 _f_permutation__U225  ( .A(out[424]), .B(_f_permutation__n1743 ), 
        .ZN(_f_permutation__round_in[1488]) );
  NAND2_X2 _f_permutation__U224  ( .A1(padder_out[465]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1742 ) );
  XNOR2_X2 _f_permutation__U223  ( .A(out[425]), .B(_f_permutation__n1742 ), 
        .ZN(_f_permutation__round_in[1489]) );
  NAND2_X2 _f_permutation__U222  ( .A1(padder_out[466]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1741 ) );
  XNOR2_X2 _f_permutation__U221  ( .A(out[426]), .B(_f_permutation__n1741 ), 
        .ZN(_f_permutation__round_in[1490]) );
  NAND2_X2 _f_permutation__U220  ( .A1(padder_out[467]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1740 ) );
  XNOR2_X2 _f_permutation__U219  ( .A(out[427]), .B(_f_permutation__n1740 ), 
        .ZN(_f_permutation__round_in[1491]) );
  NAND2_X2 _f_permutation__U218  ( .A1(padder_out[468]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1739 ) );
  XNOR2_X2 _f_permutation__U217  ( .A(out[428]), .B(_f_permutation__n1739 ), 
        .ZN(_f_permutation__round_in[1492]) );
  NAND2_X2 _f_permutation__U216  ( .A1(padder_out[469]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1738 ) );
  XNOR2_X2 _f_permutation__U215  ( .A(out[429]), .B(_f_permutation__n1738 ), 
        .ZN(_f_permutation__round_in[1493]) );
  NAND2_X2 _f_permutation__U214  ( .A1(padder_out[470]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1737 ) );
  XNOR2_X2 _f_permutation__U213  ( .A(out[430]), .B(_f_permutation__n1737 ), 
        .ZN(_f_permutation__round_in[1494]) );
  NAND2_X2 _f_permutation__U212  ( .A1(padder_out[471]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1736 ) );
  XNOR2_X2 _f_permutation__U211  ( .A(out[431]), .B(_f_permutation__n1736 ), 
        .ZN(_f_permutation__round_in[1495]) );
  NAND2_X2 _f_permutation__U210  ( .A1(padder_out[472]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1735 ) );
  XNOR2_X2 _f_permutation__U209  ( .A(out[416]), .B(_f_permutation__n1735 ), 
        .ZN(_f_permutation__round_in[1496]) );
  NAND2_X2 _f_permutation__U208  ( .A1(padder_out[473]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1734 ) );
  XNOR2_X2 _f_permutation__U207  ( .A(out[417]), .B(_f_permutation__n1734 ), 
        .ZN(_f_permutation__round_in[1497]) );
  NAND2_X2 _f_permutation__U206  ( .A1(padder_out[474]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1733 ) );
  XNOR2_X2 _f_permutation__U205  ( .A(out[418]), .B(_f_permutation__n1733 ), 
        .ZN(_f_permutation__round_in[1498]) );
  NAND2_X2 _f_permutation__U204  ( .A1(padder_out[475]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1732 ) );
  XNOR2_X2 _f_permutation__U203  ( .A(out[419]), .B(_f_permutation__n1732 ), 
        .ZN(_f_permutation__round_in[1499]) );
  NAND2_X2 _f_permutation__U202  ( .A1(padder_out[476]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1731 ) );
  XNOR2_X2 _f_permutation__U201  ( .A(out[420]), .B(_f_permutation__n1731 ), 
        .ZN(_f_permutation__round_in[1500]) );
  NAND2_X2 _f_permutation__U200  ( .A1(padder_out[477]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1730 ) );
  XNOR2_X2 _f_permutation__U199  ( .A(out[421]), .B(_f_permutation__n1730 ), 
        .ZN(_f_permutation__round_in[1501]) );
  NAND2_X2 _f_permutation__U198  ( .A1(padder_out[478]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1729 ) );
  XNOR2_X2 _f_permutation__U197  ( .A(out[422]), .B(_f_permutation__n1729 ), 
        .ZN(_f_permutation__round_in[1502]) );
  NAND2_X2 _f_permutation__U196  ( .A1(padder_out[479]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1728 ) );
  XNOR2_X2 _f_permutation__U195  ( .A(out[423]), .B(_f_permutation__n1728 ), 
        .ZN(_f_permutation__round_in[1503]) );
  NAND2_X2 _f_permutation__U194  ( .A1(padder_out[480]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1727 ) );
  XNOR2_X2 _f_permutation__U193  ( .A(out[408]), .B(_f_permutation__n1727 ), 
        .ZN(_f_permutation__round_in[1504]) );
  NAND2_X2 _f_permutation__U192  ( .A1(padder_out[481]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1726 ) );
  XNOR2_X2 _f_permutation__U191  ( .A(out[409]), .B(_f_permutation__n1726 ), 
        .ZN(_f_permutation__round_in[1505]) );
  NAND2_X2 _f_permutation__U190  ( .A1(padder_out[482]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1725 ) );
  XNOR2_X2 _f_permutation__U189  ( .A(out[410]), .B(_f_permutation__n1725 ), 
        .ZN(_f_permutation__round_in[1506]) );
  NAND2_X2 _f_permutation__U188  ( .A1(padder_out[483]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1724 ) );
  XNOR2_X2 _f_permutation__U187  ( .A(out[411]), .B(_f_permutation__n1724 ), 
        .ZN(_f_permutation__round_in[1507]) );
  NAND2_X2 _f_permutation__U186  ( .A1(padder_out[484]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1723 ) );
  XNOR2_X2 _f_permutation__U185  ( .A(out[412]), .B(_f_permutation__n1723 ), 
        .ZN(_f_permutation__round_in[1508]) );
  NAND2_X2 _f_permutation__U184  ( .A1(padder_out[485]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1722 ) );
  XNOR2_X2 _f_permutation__U183  ( .A(out[413]), .B(_f_permutation__n1722 ), 
        .ZN(_f_permutation__round_in[1509]) );
  NAND2_X2 _f_permutation__U182  ( .A1(padder_out[486]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1721 ) );
  XNOR2_X2 _f_permutation__U181  ( .A(out[414]), .B(_f_permutation__n1721 ), 
        .ZN(_f_permutation__round_in[1510]) );
  NAND2_X2 _f_permutation__U180  ( .A1(padder_out[487]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1720 ) );
  XNOR2_X2 _f_permutation__U179  ( .A(out[415]), .B(_f_permutation__n1720 ), 
        .ZN(_f_permutation__round_in[1511]) );
  NAND2_X2 _f_permutation__U178  ( .A1(padder_out[488]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1719 ) );
  XNOR2_X2 _f_permutation__U177  ( .A(out[400]), .B(_f_permutation__n1719 ), 
        .ZN(_f_permutation__round_in[1512]) );
  NAND2_X2 _f_permutation__U176  ( .A1(padder_out[489]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1718 ) );
  XNOR2_X2 _f_permutation__U175  ( .A(out[401]), .B(_f_permutation__n1718 ), 
        .ZN(_f_permutation__round_in[1513]) );
  NAND2_X2 _f_permutation__U174  ( .A1(padder_out[490]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1717 ) );
  XNOR2_X2 _f_permutation__U173  ( .A(out[402]), .B(_f_permutation__n1717 ), 
        .ZN(_f_permutation__round_in[1514]) );
  NAND2_X2 _f_permutation__U172  ( .A1(padder_out[491]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1716 ) );
  XNOR2_X2 _f_permutation__U171  ( .A(out[403]), .B(_f_permutation__n1716 ), 
        .ZN(_f_permutation__round_in[1515]) );
  NAND2_X2 _f_permutation__U170  ( .A1(padder_out[492]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1715 ) );
  XNOR2_X2 _f_permutation__U169  ( .A(out[404]), .B(_f_permutation__n1715 ), 
        .ZN(_f_permutation__round_in[1516]) );
  NAND2_X2 _f_permutation__U168  ( .A1(padder_out[493]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1714 ) );
  XNOR2_X2 _f_permutation__U167  ( .A(out[405]), .B(_f_permutation__n1714 ), 
        .ZN(_f_permutation__round_in[1517]) );
  NAND2_X2 _f_permutation__U166  ( .A1(padder_out[494]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1713 ) );
  XNOR2_X2 _f_permutation__U165  ( .A(out[406]), .B(_f_permutation__n1713 ), 
        .ZN(_f_permutation__round_in[1518]) );
  NAND2_X2 _f_permutation__U164  ( .A1(padder_out[495]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1712 ) );
  XNOR2_X2 _f_permutation__U163  ( .A(out[407]), .B(_f_permutation__n1712 ), 
        .ZN(_f_permutation__round_in[1519]) );
  NAND2_X2 _f_permutation__U162  ( .A1(padder_out[496]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1711 ) );
  XNOR2_X2 _f_permutation__U161  ( .A(out[392]), .B(_f_permutation__n1711 ), 
        .ZN(_f_permutation__round_in[1520]) );
  NAND2_X2 _f_permutation__U160  ( .A1(padder_out[497]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1710 ) );
  XNOR2_X2 _f_permutation__U159  ( .A(out[393]), .B(_f_permutation__n1710 ), 
        .ZN(_f_permutation__round_in[1521]) );
  NAND2_X2 _f_permutation__U158  ( .A1(padder_out[498]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1709 ) );
  XNOR2_X2 _f_permutation__U157  ( .A(out[394]), .B(_f_permutation__n1709 ), 
        .ZN(_f_permutation__round_in[1522]) );
  NAND2_X2 _f_permutation__U156  ( .A1(padder_out[499]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1708 ) );
  XNOR2_X2 _f_permutation__U155  ( .A(out[395]), .B(_f_permutation__n1708 ), 
        .ZN(_f_permutation__round_in[1523]) );
  NAND2_X2 _f_permutation__U154  ( .A1(padder_out[500]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1707 ) );
  XNOR2_X2 _f_permutation__U153  ( .A(out[396]), .B(_f_permutation__n1707 ), 
        .ZN(_f_permutation__round_in[1524]) );
  NAND2_X2 _f_permutation__U152  ( .A1(padder_out[501]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1706 ) );
  XNOR2_X2 _f_permutation__U151  ( .A(out[397]), .B(_f_permutation__n1706 ), 
        .ZN(_f_permutation__round_in[1525]) );
  NAND2_X2 _f_permutation__U150  ( .A1(padder_out[502]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1705 ) );
  XNOR2_X2 _f_permutation__U149  ( .A(out[398]), .B(_f_permutation__n1705 ), 
        .ZN(_f_permutation__round_in[1526]) );
  NAND2_X2 _f_permutation__U148  ( .A1(padder_out[503]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1704 ) );
  XNOR2_X2 _f_permutation__U147  ( .A(out[399]), .B(_f_permutation__n1704 ), 
        .ZN(_f_permutation__round_in[1527]) );
  NAND2_X2 _f_permutation__U146  ( .A1(padder_out[504]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1703 ) );
  XNOR2_X2 _f_permutation__U145  ( .A(out[384]), .B(_f_permutation__n1703 ), 
        .ZN(_f_permutation__round_in[1528]) );
  NAND2_X2 _f_permutation__U144  ( .A1(padder_out[505]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1702 ) );
  XNOR2_X2 _f_permutation__U143  ( .A(out[385]), .B(_f_permutation__n1702 ), 
        .ZN(_f_permutation__round_in[1529]) );
  NAND2_X2 _f_permutation__U142  ( .A1(padder_out[506]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1701 ) );
  XNOR2_X2 _f_permutation__U141  ( .A(out[386]), .B(_f_permutation__n1701 ), 
        .ZN(_f_permutation__round_in[1530]) );
  NAND2_X2 _f_permutation__U140  ( .A1(padder_out[507]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1700 ) );
  XNOR2_X2 _f_permutation__U139  ( .A(out[387]), .B(_f_permutation__n1700 ), 
        .ZN(_f_permutation__round_in[1531]) );
  NAND2_X2 _f_permutation__U138  ( .A1(padder_out[508]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1699 ) );
  XNOR2_X2 _f_permutation__U137  ( .A(out[388]), .B(_f_permutation__n1699 ), 
        .ZN(_f_permutation__round_in[1532]) );
  NAND2_X2 _f_permutation__U136  ( .A1(padder_out[509]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1698 ) );
  XNOR2_X2 _f_permutation__U135  ( .A(out[389]), .B(_f_permutation__n1698 ), 
        .ZN(_f_permutation__round_in[1533]) );
  NAND2_X2 _f_permutation__U134  ( .A1(padder_out[510]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1697 ) );
  XNOR2_X2 _f_permutation__U133  ( .A(out[390]), .B(_f_permutation__n1697 ), 
        .ZN(_f_permutation__round_in[1534]) );
  NAND2_X2 _f_permutation__U132  ( .A1(padder_out[511]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1696 ) );
  XNOR2_X2 _f_permutation__U131  ( .A(out[391]), .B(_f_permutation__n1696 ), 
        .ZN(_f_permutation__round_in[1535]) );
  NAND2_X2 _f_permutation__U130  ( .A1(padder_out[512]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1695 ) );
  XNOR2_X2 _f_permutation__U129  ( .A(out[504]), .B(_f_permutation__n1695 ), 
        .ZN(_f_permutation__round_in[1536]) );
  NAND2_X2 _f_permutation__U128  ( .A1(padder_out[513]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1694 ) );
  XNOR2_X2 _f_permutation__U127  ( .A(out[505]), .B(_f_permutation__n1694 ), 
        .ZN(_f_permutation__round_in[1537]) );
  NAND2_X2 _f_permutation__U126  ( .A1(padder_out[514]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1693 ) );
  XNOR2_X2 _f_permutation__U125  ( .A(out[506]), .B(_f_permutation__n1693 ), 
        .ZN(_f_permutation__round_in[1538]) );
  NAND2_X2 _f_permutation__U124  ( .A1(padder_out[515]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1692 ) );
  XNOR2_X2 _f_permutation__U123  ( .A(out[507]), .B(_f_permutation__n1692 ), 
        .ZN(_f_permutation__round_in[1539]) );
  NAND2_X2 _f_permutation__U122  ( .A1(padder_out[516]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1691 ) );
  XNOR2_X2 _f_permutation__U121  ( .A(out[508]), .B(_f_permutation__n1691 ), 
        .ZN(_f_permutation__round_in[1540]) );
  NAND2_X2 _f_permutation__U120  ( .A1(padder_out[517]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1690 ) );
  XNOR2_X2 _f_permutation__U119  ( .A(out[509]), .B(_f_permutation__n1690 ), 
        .ZN(_f_permutation__round_in[1541]) );
  NAND2_X2 _f_permutation__U118  ( .A1(padder_out[518]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1689 ) );
  XNOR2_X2 _f_permutation__U117  ( .A(out[510]), .B(_f_permutation__n1689 ), 
        .ZN(_f_permutation__round_in[1542]) );
  NAND2_X2 _f_permutation__U116  ( .A1(padder_out[519]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1688 ) );
  XNOR2_X2 _f_permutation__U115  ( .A(out[511]), .B(_f_permutation__n1688 ), 
        .ZN(_f_permutation__round_in[1543]) );
  NAND2_X2 _f_permutation__U114  ( .A1(padder_out[520]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1687 ) );
  XNOR2_X2 _f_permutation__U113  ( .A(out[496]), .B(_f_permutation__n1687 ), 
        .ZN(_f_permutation__round_in[1544]) );
  NAND2_X2 _f_permutation__U112  ( .A1(padder_out[521]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1686 ) );
  XNOR2_X2 _f_permutation__U111  ( .A(out[497]), .B(_f_permutation__n1686 ), 
        .ZN(_f_permutation__round_in[1545]) );
  NAND2_X2 _f_permutation__U110  ( .A1(padder_out[522]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1685 ) );
  XNOR2_X2 _f_permutation__U109  ( .A(out[498]), .B(_f_permutation__n1685 ), 
        .ZN(_f_permutation__round_in[1546]) );
  NAND2_X2 _f_permutation__U108  ( .A1(padder_out[523]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1684 ) );
  XNOR2_X2 _f_permutation__U107  ( .A(out[499]), .B(_f_permutation__n1684 ), 
        .ZN(_f_permutation__round_in[1547]) );
  NAND2_X2 _f_permutation__U106  ( .A1(padder_out[524]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1683 ) );
  XNOR2_X2 _f_permutation__U105  ( .A(out[500]), .B(_f_permutation__n1683 ), 
        .ZN(_f_permutation__round_in[1548]) );
  NAND2_X2 _f_permutation__U104  ( .A1(padder_out[525]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1682 ) );
  XNOR2_X2 _f_permutation__U103  ( .A(out[501]), .B(_f_permutation__n1682 ), 
        .ZN(_f_permutation__round_in[1549]) );
  NAND2_X2 _f_permutation__U102  ( .A1(padder_out[526]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1681 ) );
  XNOR2_X2 _f_permutation__U101  ( .A(out[502]), .B(_f_permutation__n1681 ), 
        .ZN(_f_permutation__round_in[1550]) );
  NAND2_X2 _f_permutation__U100  ( .A1(padder_out[527]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1680 ) );
  XNOR2_X2 _f_permutation__U99  ( .A(out[503]), .B(_f_permutation__n1680 ), 
        .ZN(_f_permutation__round_in[1551]) );
  NAND2_X2 _f_permutation__U98  ( .A1(padder_out[528]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1679 ) );
  XNOR2_X2 _f_permutation__U97  ( .A(out[488]), .B(_f_permutation__n1679 ), 
        .ZN(_f_permutation__round_in[1552]) );
  NAND2_X2 _f_permutation__U96  ( .A1(padder_out[529]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1678 ) );
  XNOR2_X2 _f_permutation__U95  ( .A(out[489]), .B(_f_permutation__n1678 ), 
        .ZN(_f_permutation__round_in[1553]) );
  NAND2_X2 _f_permutation__U94  ( .A1(padder_out[530]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1677 ) );
  XNOR2_X2 _f_permutation__U93  ( .A(out[490]), .B(_f_permutation__n1677 ), 
        .ZN(_f_permutation__round_in[1554]) );
  NAND2_X2 _f_permutation__U92  ( .A1(padder_out[531]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1676 ) );
  XNOR2_X2 _f_permutation__U91  ( .A(out[491]), .B(_f_permutation__n1676 ), 
        .ZN(_f_permutation__round_in[1555]) );
  NAND2_X2 _f_permutation__U90  ( .A1(padder_out[532]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1675 ) );
  XNOR2_X2 _f_permutation__U89  ( .A(out[492]), .B(_f_permutation__n1675 ), 
        .ZN(_f_permutation__round_in[1556]) );
  NAND2_X2 _f_permutation__U88  ( .A1(padder_out[533]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1674 ) );
  XNOR2_X2 _f_permutation__U87  ( .A(out[493]), .B(_f_permutation__n1674 ), 
        .ZN(_f_permutation__round_in[1557]) );
  NAND2_X2 _f_permutation__U86  ( .A1(padder_out[534]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1673 ) );
  XNOR2_X2 _f_permutation__U85  ( .A(out[494]), .B(_f_permutation__n1673 ), 
        .ZN(_f_permutation__round_in[1558]) );
  NAND2_X2 _f_permutation__U84  ( .A1(padder_out[535]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1672 ) );
  XNOR2_X2 _f_permutation__U83  ( .A(out[495]), .B(_f_permutation__n1672 ), 
        .ZN(_f_permutation__round_in[1559]) );
  NAND2_X2 _f_permutation__U82  ( .A1(padder_out[536]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1671 ) );
  XNOR2_X2 _f_permutation__U81  ( .A(out[480]), .B(_f_permutation__n1671 ), 
        .ZN(_f_permutation__round_in[1560]) );
  NAND2_X2 _f_permutation__U80  ( .A1(padder_out[537]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1670 ) );
  XNOR2_X2 _f_permutation__U79  ( .A(out[481]), .B(_f_permutation__n1670 ), 
        .ZN(_f_permutation__round_in[1561]) );
  NAND2_X2 _f_permutation__U78  ( .A1(padder_out[538]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1669 ) );
  XNOR2_X2 _f_permutation__U77  ( .A(out[482]), .B(_f_permutation__n1669 ), 
        .ZN(_f_permutation__round_in[1562]) );
  NAND2_X2 _f_permutation__U76  ( .A1(padder_out[539]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1668 ) );
  XNOR2_X2 _f_permutation__U75  ( .A(out[483]), .B(_f_permutation__n1668 ), 
        .ZN(_f_permutation__round_in[1563]) );
  NAND2_X2 _f_permutation__U74  ( .A1(padder_out[540]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1667 ) );
  XNOR2_X2 _f_permutation__U73  ( .A(out[484]), .B(_f_permutation__n1667 ), 
        .ZN(_f_permutation__round_in[1564]) );
  NAND2_X2 _f_permutation__U72  ( .A1(padder_out[541]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1666 ) );
  XNOR2_X2 _f_permutation__U71  ( .A(out[485]), .B(_f_permutation__n1666 ), 
        .ZN(_f_permutation__round_in[1565]) );
  NAND2_X2 _f_permutation__U70  ( .A1(padder_out[542]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1665 ) );
  XNOR2_X2 _f_permutation__U69  ( .A(out[486]), .B(_f_permutation__n1665 ), 
        .ZN(_f_permutation__round_in[1566]) );
  NAND2_X2 _f_permutation__U68  ( .A1(padder_out[543]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1664 ) );
  XNOR2_X2 _f_permutation__U67  ( .A(out[487]), .B(_f_permutation__n1664 ), 
        .ZN(_f_permutation__round_in[1567]) );
  NAND2_X2 _f_permutation__U66  ( .A1(padder_out[544]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1663 ) );
  XNOR2_X2 _f_permutation__U65  ( .A(out[472]), .B(_f_permutation__n1663 ), 
        .ZN(_f_permutation__round_in[1568]) );
  NAND2_X2 _f_permutation__U64  ( .A1(padder_out[545]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1662 ) );
  XNOR2_X2 _f_permutation__U63  ( .A(out[473]), .B(_f_permutation__n1662 ), 
        .ZN(_f_permutation__round_in[1569]) );
  NAND2_X2 _f_permutation__U62  ( .A1(padder_out[546]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1661 ) );
  XNOR2_X2 _f_permutation__U61  ( .A(out[474]), .B(_f_permutation__n1661 ), 
        .ZN(_f_permutation__round_in[1570]) );
  NAND2_X2 _f_permutation__U60  ( .A1(padder_out[547]), .A2(
        _f_permutation__n7315 ), .ZN(_f_permutation__n1660 ) );
  XNOR2_X2 _f_permutation__U59  ( .A(out[475]), .B(_f_permutation__n1660 ), 
        .ZN(_f_permutation__round_in[1571]) );
  NAND2_X2 _f_permutation__U58  ( .A1(padder_out[548]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1659 ) );
  XNOR2_X2 _f_permutation__U57  ( .A(out[476]), .B(_f_permutation__n1659 ), 
        .ZN(_f_permutation__round_in[1572]) );
  NAND2_X2 _f_permutation__U56  ( .A1(padder_out[549]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1658 ) );
  XNOR2_X2 _f_permutation__U55  ( .A(out[477]), .B(_f_permutation__n1658 ), 
        .ZN(_f_permutation__round_in[1573]) );
  NAND2_X2 _f_permutation__U54  ( .A1(padder_out[550]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1657 ) );
  XNOR2_X2 _f_permutation__U53  ( .A(out[478]), .B(_f_permutation__n1657 ), 
        .ZN(_f_permutation__round_in[1574]) );
  NAND2_X2 _f_permutation__U52  ( .A1(padder_out[551]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1656 ) );
  XNOR2_X2 _f_permutation__U51  ( .A(out[479]), .B(_f_permutation__n1656 ), 
        .ZN(_f_permutation__round_in[1575]) );
  NAND2_X2 _f_permutation__U50  ( .A1(padder_out[552]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1655 ) );
  XNOR2_X2 _f_permutation__U49  ( .A(out[464]), .B(_f_permutation__n1655 ), 
        .ZN(_f_permutation__round_in[1576]) );
  NAND2_X2 _f_permutation__U48  ( .A1(padder_out[553]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1654 ) );
  XNOR2_X2 _f_permutation__U47  ( .A(out[465]), .B(_f_permutation__n1654 ), 
        .ZN(_f_permutation__round_in[1577]) );
  NAND2_X2 _f_permutation__U46  ( .A1(padder_out[554]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1653 ) );
  XNOR2_X2 _f_permutation__U45  ( .A(out[466]), .B(_f_permutation__n1653 ), 
        .ZN(_f_permutation__round_in[1578]) );
  NAND2_X2 _f_permutation__U44  ( .A1(padder_out[555]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1652 ) );
  XNOR2_X2 _f_permutation__U43  ( .A(out[467]), .B(_f_permutation__n1652 ), 
        .ZN(_f_permutation__round_in[1579]) );
  NAND2_X2 _f_permutation__U42  ( .A1(padder_out[556]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1651 ) );
  XNOR2_X2 _f_permutation__U41  ( .A(out[468]), .B(_f_permutation__n1651 ), 
        .ZN(_f_permutation__round_in[1580]) );
  NAND2_X2 _f_permutation__U40  ( .A1(padder_out[557]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1650 ) );
  XNOR2_X2 _f_permutation__U39  ( .A(out[469]), .B(_f_permutation__n1650 ), 
        .ZN(_f_permutation__round_in[1581]) );
  NAND2_X2 _f_permutation__U38  ( .A1(padder_out[558]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1649 ) );
  XNOR2_X2 _f_permutation__U37  ( .A(out[470]), .B(_f_permutation__n1649 ), 
        .ZN(_f_permutation__round_in[1582]) );
  NAND2_X2 _f_permutation__U36  ( .A1(padder_out[559]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1648 ) );
  XNOR2_X2 _f_permutation__U35  ( .A(out[471]), .B(_f_permutation__n1648 ), 
        .ZN(_f_permutation__round_in[1583]) );
  NAND2_X2 _f_permutation__U34  ( .A1(padder_out[560]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1647 ) );
  XNOR2_X2 _f_permutation__U33  ( .A(out[456]), .B(_f_permutation__n1647 ), 
        .ZN(_f_permutation__round_in[1584]) );
  NAND2_X2 _f_permutation__U32  ( .A1(padder_out[561]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1646 ) );
  XNOR2_X2 _f_permutation__U31  ( .A(out[457]), .B(_f_permutation__n1646 ), 
        .ZN(_f_permutation__round_in[1585]) );
  NAND2_X2 _f_permutation__U30  ( .A1(padder_out[562]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1645 ) );
  XNOR2_X2 _f_permutation__U29  ( .A(out[458]), .B(_f_permutation__n1645 ), 
        .ZN(_f_permutation__round_in[1586]) );
  NAND2_X2 _f_permutation__U28  ( .A1(padder_out[563]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1644 ) );
  XNOR2_X2 _f_permutation__U27  ( .A(out[459]), .B(_f_permutation__n1644 ), 
        .ZN(_f_permutation__round_in[1587]) );
  NAND2_X2 _f_permutation__U26  ( .A1(padder_out[564]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1643 ) );
  XNOR2_X2 _f_permutation__U25  ( .A(out[460]), .B(_f_permutation__n1643 ), 
        .ZN(_f_permutation__round_in[1588]) );
  NAND2_X2 _f_permutation__U24  ( .A1(padder_out[565]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1642 ) );
  XNOR2_X2 _f_permutation__U23  ( .A(out[461]), .B(_f_permutation__n1642 ), 
        .ZN(_f_permutation__round_in[1589]) );
  NAND2_X2 _f_permutation__U22  ( .A1(padder_out[566]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1641 ) );
  XNOR2_X2 _f_permutation__U21  ( .A(out[462]), .B(_f_permutation__n1641 ), 
        .ZN(_f_permutation__round_in[1590]) );
  NAND2_X2 _f_permutation__U20  ( .A1(padder_out[567]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1640 ) );
  XNOR2_X2 _f_permutation__U19  ( .A(out[463]), .B(_f_permutation__n1640 ), 
        .ZN(_f_permutation__round_in[1591]) );
  NAND2_X2 _f_permutation__U18  ( .A1(padder_out[568]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1639 ) );
  XNOR2_X2 _f_permutation__U17  ( .A(out[448]), .B(_f_permutation__n1639 ), 
        .ZN(_f_permutation__round_in[1592]) );
  NAND2_X2 _f_permutation__U16  ( .A1(padder_out[569]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1638 ) );
  XNOR2_X2 _f_permutation__U15  ( .A(out[449]), .B(_f_permutation__n1638 ), 
        .ZN(_f_permutation__round_in[1593]) );
  NAND2_X2 _f_permutation__U14  ( .A1(padder_out[570]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1637 ) );
  XNOR2_X2 _f_permutation__U13  ( .A(out[450]), .B(_f_permutation__n1637 ), 
        .ZN(_f_permutation__round_in[1594]) );
  NAND2_X2 _f_permutation__U12  ( .A1(padder_out[571]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1636 ) );
  XNOR2_X2 _f_permutation__U11  ( .A(out[451]), .B(_f_permutation__n1636 ), 
        .ZN(_f_permutation__round_in[1595]) );
  NAND2_X2 _f_permutation__U10  ( .A1(padder_out[572]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1635 ) );
  XNOR2_X2 _f_permutation__U9  ( .A(out[452]), .B(_f_permutation__n1635 ), 
        .ZN(_f_permutation__round_in[1596]) );
  NAND2_X2 _f_permutation__U8  ( .A1(padder_out[573]), .A2(
        _f_permutation__n7314 ), .ZN(_f_permutation__n1634 ) );
  XNOR2_X2 _f_permutation__U7  ( .A(out[453]), .B(_f_permutation__n1634 ), 
        .ZN(_f_permutation__round_in[1597]) );
  NAND2_X2 _f_permutation__U6  ( .A1(padder_out[574]), .A2(
        _f_permutation__n7316 ), .ZN(_f_permutation__n1633 ) );
  XNOR2_X2 _f_permutation__U5  ( .A(out[454]), .B(_f_permutation__n1633 ), 
        .ZN(_f_permutation__round_in[1598]) );
  NAND2_X2 _f_permutation__U4  ( .A1(padder_out[575]), .A2(
        _f_permutation__n7317 ), .ZN(_f_permutation__n1632 ) );
  XNOR2_X2 _f_permutation__U3  ( .A(out[455]), .B(_f_permutation__n1632 ), 
        .ZN(_f_permutation__round_in[1599]) );
  DFF_X2 _f_permutation__out_reg_1599_  ( .D(_f_permutation__n3788 ), .CK(clk), 
        .Q(out[455]), .QN() );
  DFF_X2 _f_permutation__out_reg_1598_  ( .D(_f_permutation__n3789 ), .CK(clk), 
        .Q(out[454]), .QN() );
  DFF_X2 _f_permutation__out_reg_1597_  ( .D(_f_permutation__n3790 ), .CK(clk), 
        .Q(out[453]), .QN() );
  DFF_X2 _f_permutation__out_reg_1596_  ( .D(_f_permutation__n3791 ), .CK(clk), 
        .Q(out[452]), .QN() );
  DFF_X2 _f_permutation__out_reg_1595_  ( .D(_f_permutation__n3792 ), .CK(clk), 
        .Q(out[451]), .QN() );
  DFF_X2 _f_permutation__out_reg_1594_  ( .D(_f_permutation__n3793 ), .CK(clk), 
        .Q(out[450]), .QN() );
  DFF_X2 _f_permutation__out_reg_1593_  ( .D(_f_permutation__n3794 ), .CK(clk), 
        .Q(out[449]), .QN() );
  DFF_X2 _f_permutation__out_reg_1592_  ( .D(_f_permutation__n3795 ), .CK(clk), 
        .Q(out[448]), .QN() );
  DFF_X2 _f_permutation__out_reg_1591_  ( .D(_f_permutation__n3796 ), .CK(clk), 
        .Q(out[463]), .QN() );
  DFF_X2 _f_permutation__out_reg_1590_  ( .D(_f_permutation__n3797 ), .CK(clk), 
        .Q(out[462]), .QN() );
  DFF_X2 _f_permutation__out_reg_1589_  ( .D(_f_permutation__n3798 ), .CK(clk), 
        .Q(out[461]), .QN() );
  DFF_X2 _f_permutation__out_reg_1588_  ( .D(_f_permutation__n3799 ), .CK(clk), 
        .Q(out[460]), .QN() );
  DFF_X2 _f_permutation__out_reg_1587_  ( .D(_f_permutation__n3800 ), .CK(clk), 
        .Q(out[459]), .QN() );
  DFF_X2 _f_permutation__out_reg_1586_  ( .D(_f_permutation__n3801 ), .CK(clk), 
        .Q(out[458]), .QN() );
  DFF_X2 _f_permutation__out_reg_1585_  ( .D(_f_permutation__n3802 ), .CK(clk), 
        .Q(out[457]), .QN() );
  DFF_X2 _f_permutation__out_reg_1584_  ( .D(_f_permutation__n3803 ), .CK(clk), 
        .Q(out[456]), .QN() );
  DFF_X2 _f_permutation__out_reg_1583_  ( .D(_f_permutation__n3804 ), .CK(clk), 
        .Q(out[471]), .QN() );
  DFF_X2 _f_permutation__out_reg_1582_  ( .D(_f_permutation__n3805 ), .CK(clk), 
        .Q(out[470]), .QN() );
  DFF_X2 _f_permutation__out_reg_1581_  ( .D(_f_permutation__n3806 ), .CK(clk), 
        .Q(out[469]), .QN() );
  DFF_X2 _f_permutation__out_reg_1580_  ( .D(_f_permutation__n3807 ), .CK(clk), 
        .Q(out[468]), .QN() );
  DFF_X2 _f_permutation__out_reg_1579_  ( .D(_f_permutation__n3808 ), .CK(clk), 
        .Q(out[467]), .QN() );
  DFF_X2 _f_permutation__out_reg_1578_  ( .D(_f_permutation__n3809 ), .CK(clk), 
        .Q(out[466]), .QN() );
  DFF_X2 _f_permutation__out_reg_1577_  ( .D(_f_permutation__n3810 ), .CK(clk), 
        .Q(out[465]), .QN() );
  DFF_X2 _f_permutation__out_reg_1576_  ( .D(_f_permutation__n3811 ), .CK(clk), 
        .Q(out[464]), .QN() );
  DFF_X2 _f_permutation__out_reg_1575_  ( .D(_f_permutation__n3812 ), .CK(clk), 
        .Q(out[479]), .QN() );
  DFF_X2 _f_permutation__out_reg_1574_  ( .D(_f_permutation__n3813 ), .CK(clk), 
        .Q(out[478]), .QN() );
  DFF_X2 _f_permutation__out_reg_1573_  ( .D(_f_permutation__n3814 ), .CK(clk), 
        .Q(out[477]), .QN() );
  DFF_X2 _f_permutation__out_reg_1572_  ( .D(_f_permutation__n3815 ), .CK(clk), 
        .Q(out[476]), .QN() );
  DFF_X2 _f_permutation__out_reg_1571_  ( .D(_f_permutation__n3816 ), .CK(clk), 
        .Q(out[475]), .QN() );
  DFF_X2 _f_permutation__out_reg_1570_  ( .D(_f_permutation__n3817 ), .CK(clk), 
        .Q(out[474]), .QN() );
  DFF_X2 _f_permutation__out_reg_1569_  ( .D(_f_permutation__n3818 ), .CK(clk), 
        .Q(out[473]), .QN() );
  DFF_X2 _f_permutation__out_reg_1568_  ( .D(_f_permutation__n3819 ), .CK(clk), 
        .Q(out[472]), .QN() );
  DFF_X2 _f_permutation__out_reg_1567_  ( .D(_f_permutation__n3820 ), .CK(clk), 
        .Q(out[487]), .QN() );
  DFF_X2 _f_permutation__out_reg_1566_  ( .D(_f_permutation__n3821 ), .CK(clk), 
        .Q(out[486]), .QN() );
  DFF_X2 _f_permutation__out_reg_1565_  ( .D(_f_permutation__n3822 ), .CK(clk), 
        .Q(out[485]), .QN() );
  DFF_X2 _f_permutation__out_reg_1564_  ( .D(_f_permutation__n3823 ), .CK(clk), 
        .Q(out[484]), .QN() );
  DFF_X2 _f_permutation__out_reg_1563_  ( .D(_f_permutation__n3824 ), .CK(clk), 
        .Q(out[483]), .QN() );
  DFF_X2 _f_permutation__out_reg_1562_  ( .D(_f_permutation__n3825 ), .CK(clk), 
        .Q(out[482]), .QN() );
  DFF_X2 _f_permutation__out_reg_1561_  ( .D(_f_permutation__n3826 ), .CK(clk), 
        .Q(out[481]), .QN() );
  DFF_X2 _f_permutation__out_reg_1560_  ( .D(_f_permutation__n3827 ), .CK(clk), 
        .Q(out[480]), .QN() );
  DFF_X2 _f_permutation__out_reg_1559_  ( .D(_f_permutation__n3828 ), .CK(clk), 
        .Q(out[495]), .QN() );
  DFF_X2 _f_permutation__out_reg_1558_  ( .D(_f_permutation__n3829 ), .CK(clk), 
        .Q(out[494]), .QN() );
  DFF_X2 _f_permutation__out_reg_1557_  ( .D(_f_permutation__n3830 ), .CK(clk), 
        .Q(out[493]), .QN() );
  DFF_X2 _f_permutation__out_reg_1556_  ( .D(_f_permutation__n3831 ), .CK(clk), 
        .Q(out[492]), .QN() );
  DFF_X2 _f_permutation__out_reg_1555_  ( .D(_f_permutation__n3832 ), .CK(clk), 
        .Q(out[491]), .QN() );
  DFF_X2 _f_permutation__out_reg_1554_  ( .D(_f_permutation__n3833 ), .CK(clk), 
        .Q(out[490]), .QN() );
  DFF_X2 _f_permutation__out_reg_1553_  ( .D(_f_permutation__n3834 ), .CK(clk), 
        .Q(out[489]), .QN() );
  DFF_X2 _f_permutation__out_reg_1552_  ( .D(_f_permutation__n3835 ), .CK(clk), 
        .Q(out[488]), .QN() );
  DFF_X2 _f_permutation__out_reg_1551_  ( .D(_f_permutation__n3836 ), .CK(clk), 
        .Q(out[503]), .QN() );
  DFF_X2 _f_permutation__out_reg_1550_  ( .D(_f_permutation__n3837 ), .CK(clk), 
        .Q(out[502]), .QN() );
  DFF_X2 _f_permutation__out_reg_1549_  ( .D(_f_permutation__n3838 ), .CK(clk), 
        .Q(out[501]), .QN() );
  DFF_X2 _f_permutation__out_reg_1548_  ( .D(_f_permutation__n3839 ), .CK(clk), 
        .Q(out[500]), .QN() );
  DFF_X2 _f_permutation__out_reg_1547_  ( .D(_f_permutation__n3840 ), .CK(clk), 
        .Q(out[499]), .QN() );
  DFF_X2 _f_permutation__out_reg_1546_  ( .D(_f_permutation__n3841 ), .CK(clk), 
        .Q(out[498]), .QN() );
  DFF_X2 _f_permutation__out_reg_1545_  ( .D(_f_permutation__n3842 ), .CK(clk), 
        .Q(out[497]), .QN() );
  DFF_X2 _f_permutation__out_reg_1544_  ( .D(_f_permutation__n3843 ), .CK(clk), 
        .Q(out[496]), .QN() );
  DFF_X2 _f_permutation__out_reg_1543_  ( .D(_f_permutation__n3844 ), .CK(clk), 
        .Q(out[511]), .QN() );
  DFF_X2 _f_permutation__out_reg_1542_  ( .D(_f_permutation__n3845 ), .CK(clk), 
        .Q(out[510]), .QN() );
  DFF_X2 _f_permutation__out_reg_1541_  ( .D(_f_permutation__n3846 ), .CK(clk), 
        .Q(out[509]), .QN() );
  DFF_X2 _f_permutation__out_reg_1540_  ( .D(_f_permutation__n3847 ), .CK(clk), 
        .Q(out[508]), .QN() );
  DFF_X2 _f_permutation__out_reg_1539_  ( .D(_f_permutation__n3848 ), .CK(clk), 
        .Q(out[507]), .QN() );
  DFF_X2 _f_permutation__out_reg_1538_  ( .D(_f_permutation__n3849 ), .CK(clk), 
        .Q(out[506]), .QN() );
  DFF_X2 _f_permutation__out_reg_1537_  ( .D(_f_permutation__n3850 ), .CK(clk), 
        .Q(out[505]), .QN() );
  DFF_X2 _f_permutation__out_reg_1536_  ( .D(_f_permutation__n3851 ), .CK(clk), 
        .Q(out[504]), .QN() );
  DFF_X2 _f_permutation__out_reg_1535_  ( .D(_f_permutation__n3852 ), .CK(clk), 
        .Q(out[391]), .QN() );
  DFF_X2 _f_permutation__out_reg_1534_  ( .D(_f_permutation__n3853 ), .CK(clk), 
        .Q(out[390]), .QN() );
  DFF_X2 _f_permutation__out_reg_1533_  ( .D(_f_permutation__n3854 ), .CK(clk), 
        .Q(out[389]), .QN() );
  DFF_X2 _f_permutation__out_reg_1532_  ( .D(_f_permutation__n3855 ), .CK(clk), 
        .Q(out[388]), .QN() );
  DFF_X2 _f_permutation__out_reg_1531_  ( .D(_f_permutation__n3856 ), .CK(clk), 
        .Q(out[387]), .QN() );
  DFF_X2 _f_permutation__out_reg_1530_  ( .D(_f_permutation__n3857 ), .CK(clk), 
        .Q(out[386]), .QN() );
  DFF_X2 _f_permutation__out_reg_1529_  ( .D(_f_permutation__n3858 ), .CK(clk), 
        .Q(out[385]), .QN() );
  DFF_X2 _f_permutation__out_reg_1528_  ( .D(_f_permutation__n3859 ), .CK(clk), 
        .Q(out[384]), .QN() );
  DFF_X2 _f_permutation__out_reg_1527_  ( .D(_f_permutation__n3860 ), .CK(clk), 
        .Q(out[399]), .QN() );
  DFF_X2 _f_permutation__out_reg_1526_  ( .D(_f_permutation__n3861 ), .CK(clk), 
        .Q(out[398]), .QN() );
  DFF_X2 _f_permutation__out_reg_1525_  ( .D(_f_permutation__n3862 ), .CK(clk), 
        .Q(out[397]), .QN() );
  DFF_X2 _f_permutation__out_reg_1524_  ( .D(_f_permutation__n3863 ), .CK(clk), 
        .Q(out[396]), .QN() );
  DFF_X2 _f_permutation__out_reg_1523_  ( .D(_f_permutation__n3864 ), .CK(clk), 
        .Q(out[395]), .QN() );
  DFF_X2 _f_permutation__out_reg_1522_  ( .D(_f_permutation__n3865 ), .CK(clk), 
        .Q(out[394]), .QN() );
  DFF_X2 _f_permutation__out_reg_1521_  ( .D(_f_permutation__n3866 ), .CK(clk), 
        .Q(out[393]), .QN() );
  DFF_X2 _f_permutation__out_reg_1520_  ( .D(_f_permutation__n3867 ), .CK(clk), 
        .Q(out[392]), .QN() );
  DFF_X2 _f_permutation__out_reg_1519_  ( .D(_f_permutation__n3868 ), .CK(clk), 
        .Q(out[407]), .QN() );
  DFF_X2 _f_permutation__out_reg_1518_  ( .D(_f_permutation__n3869 ), .CK(clk), 
        .Q(out[406]), .QN() );
  DFF_X2 _f_permutation__out_reg_1517_  ( .D(_f_permutation__n3870 ), .CK(clk), 
        .Q(out[405]), .QN() );
  DFF_X2 _f_permutation__out_reg_1516_  ( .D(_f_permutation__n3871 ), .CK(clk), 
        .Q(out[404]), .QN() );
  DFF_X2 _f_permutation__out_reg_1515_  ( .D(_f_permutation__n3872 ), .CK(clk), 
        .Q(out[403]), .QN() );
  DFF_X2 _f_permutation__out_reg_1514_  ( .D(_f_permutation__n3873 ), .CK(clk), 
        .Q(out[402]), .QN() );
  DFF_X2 _f_permutation__out_reg_1513_  ( .D(_f_permutation__n3874 ), .CK(clk), 
        .Q(out[401]), .QN() );
  DFF_X2 _f_permutation__out_reg_1512_  ( .D(_f_permutation__n3875 ), .CK(clk), 
        .Q(out[400]), .QN() );
  DFF_X2 _f_permutation__out_reg_1511_  ( .D(_f_permutation__n3876 ), .CK(clk), 
        .Q(out[415]), .QN() );
  DFF_X2 _f_permutation__out_reg_1510_  ( .D(_f_permutation__n3877 ), .CK(clk), 
        .Q(out[414]), .QN() );
  DFF_X2 _f_permutation__out_reg_1509_  ( .D(_f_permutation__n3878 ), .CK(clk), 
        .Q(out[413]), .QN() );
  DFF_X2 _f_permutation__out_reg_1508_  ( .D(_f_permutation__n3879 ), .CK(clk), 
        .Q(out[412]), .QN() );
  DFF_X2 _f_permutation__out_reg_1507_  ( .D(_f_permutation__n3880 ), .CK(clk), 
        .Q(out[411]), .QN() );
  DFF_X2 _f_permutation__out_reg_1506_  ( .D(_f_permutation__n3881 ), .CK(clk), 
        .Q(out[410]), .QN() );
  DFF_X2 _f_permutation__out_reg_1505_  ( .D(_f_permutation__n3882 ), .CK(clk), 
        .Q(out[409]), .QN() );
  DFF_X2 _f_permutation__out_reg_1504_  ( .D(_f_permutation__n3883 ), .CK(clk), 
        .Q(out[408]), .QN() );
  DFF_X2 _f_permutation__out_reg_1503_  ( .D(_f_permutation__n3884 ), .CK(clk), 
        .Q(out[423]), .QN() );
  DFF_X2 _f_permutation__out_reg_1502_  ( .D(_f_permutation__n3885 ), .CK(clk), 
        .Q(out[422]), .QN() );
  DFF_X2 _f_permutation__out_reg_1501_  ( .D(_f_permutation__n3886 ), .CK(clk), 
        .Q(out[421]), .QN() );
  DFF_X2 _f_permutation__out_reg_1500_  ( .D(_f_permutation__n3887 ), .CK(clk), 
        .Q(out[420]), .QN() );
  DFF_X2 _f_permutation__out_reg_1499_  ( .D(_f_permutation__n3888 ), .CK(clk), 
        .Q(out[419]), .QN() );
  DFF_X2 _f_permutation__out_reg_1498_  ( .D(_f_permutation__n3889 ), .CK(clk), 
        .Q(out[418]), .QN() );
  DFF_X2 _f_permutation__out_reg_1497_  ( .D(_f_permutation__n3890 ), .CK(clk), 
        .Q(out[417]), .QN() );
  DFF_X2 _f_permutation__out_reg_1496_  ( .D(_f_permutation__n3891 ), .CK(clk), 
        .Q(out[416]), .QN() );
  DFF_X2 _f_permutation__out_reg_1495_  ( .D(_f_permutation__n3892 ), .CK(clk), 
        .Q(out[431]), .QN() );
  DFF_X2 _f_permutation__out_reg_1494_  ( .D(_f_permutation__n3893 ), .CK(clk), 
        .Q(out[430]), .QN() );
  DFF_X2 _f_permutation__out_reg_1493_  ( .D(_f_permutation__n3894 ), .CK(clk), 
        .Q(out[429]), .QN() );
  DFF_X2 _f_permutation__out_reg_1492_  ( .D(_f_permutation__n3895 ), .CK(clk), 
        .Q(out[428]), .QN() );
  DFF_X2 _f_permutation__out_reg_1491_  ( .D(_f_permutation__n3896 ), .CK(clk), 
        .Q(out[427]), .QN() );
  DFF_X2 _f_permutation__out_reg_1490_  ( .D(_f_permutation__n3897 ), .CK(clk), 
        .Q(out[426]), .QN() );
  DFF_X2 _f_permutation__out_reg_1489_  ( .D(_f_permutation__n3898 ), .CK(clk), 
        .Q(out[425]), .QN() );
  DFF_X2 _f_permutation__out_reg_1488_  ( .D(_f_permutation__n3899 ), .CK(clk), 
        .Q(out[424]), .QN() );
  DFF_X2 _f_permutation__out_reg_1487_  ( .D(_f_permutation__n3900 ), .CK(clk), 
        .Q(out[439]), .QN() );
  DFF_X2 _f_permutation__out_reg_1486_  ( .D(_f_permutation__n3901 ), .CK(clk), 
        .Q(out[438]), .QN() );
  DFF_X2 _f_permutation__out_reg_1485_  ( .D(_f_permutation__n3902 ), .CK(clk), 
        .Q(out[437]), .QN() );
  DFF_X2 _f_permutation__out_reg_1484_  ( .D(_f_permutation__n3903 ), .CK(clk), 
        .Q(out[436]), .QN() );
  DFF_X2 _f_permutation__out_reg_1483_  ( .D(_f_permutation__n3904 ), .CK(clk), 
        .Q(out[435]), .QN() );
  DFF_X2 _f_permutation__out_reg_1482_  ( .D(_f_permutation__n3905 ), .CK(clk), 
        .Q(out[434]), .QN() );
  DFF_X2 _f_permutation__out_reg_1481_  ( .D(_f_permutation__n3906 ), .CK(clk), 
        .Q(out[433]), .QN() );
  DFF_X2 _f_permutation__out_reg_1480_  ( .D(_f_permutation__n3907 ), .CK(clk), 
        .Q(out[432]), .QN() );
  DFF_X2 _f_permutation__out_reg_1479_  ( .D(_f_permutation__n3908 ), .CK(clk), 
        .Q(out[447]), .QN() );
  DFF_X2 _f_permutation__out_reg_1478_  ( .D(_f_permutation__n3909 ), .CK(clk), 
        .Q(out[446]), .QN() );
  DFF_X2 _f_permutation__out_reg_1477_  ( .D(_f_permutation__n3910 ), .CK(clk), 
        .Q(out[445]), .QN() );
  DFF_X2 _f_permutation__out_reg_1476_  ( .D(_f_permutation__n3911 ), .CK(clk), 
        .Q(out[444]), .QN() );
  DFF_X2 _f_permutation__out_reg_1475_  ( .D(_f_permutation__n3912 ), .CK(clk), 
        .Q(out[443]), .QN() );
  DFF_X2 _f_permutation__out_reg_1474_  ( .D(_f_permutation__n3913 ), .CK(clk), 
        .Q(out[442]), .QN() );
  DFF_X2 _f_permutation__out_reg_1473_  ( .D(_f_permutation__n3914 ), .CK(clk), 
        .Q(out[441]), .QN() );
  DFF_X2 _f_permutation__out_reg_1472_  ( .D(_f_permutation__n3915 ), .CK(clk), 
        .Q(out[440]), .QN() );
  DFF_X2 _f_permutation__out_reg_1471_  ( .D(_f_permutation__n3916 ), .CK(clk), 
        .Q(out[327]), .QN() );
  DFF_X2 _f_permutation__out_reg_1470_  ( .D(_f_permutation__n3917 ), .CK(clk), 
        .Q(out[326]), .QN() );
  DFF_X2 _f_permutation__out_reg_1469_  ( .D(_f_permutation__n3918 ), .CK(clk), 
        .Q(out[325]), .QN() );
  DFF_X2 _f_permutation__out_reg_1468_  ( .D(_f_permutation__n3919 ), .CK(clk), 
        .Q(out[324]), .QN() );
  DFF_X2 _f_permutation__out_reg_1467_  ( .D(_f_permutation__n3920 ), .CK(clk), 
        .Q(out[323]), .QN() );
  DFF_X2 _f_permutation__out_reg_1466_  ( .D(_f_permutation__n3921 ), .CK(clk), 
        .Q(out[322]), .QN() );
  DFF_X2 _f_permutation__out_reg_1465_  ( .D(_f_permutation__n3922 ), .CK(clk), 
        .Q(out[321]), .QN() );
  DFF_X2 _f_permutation__out_reg_1464_  ( .D(_f_permutation__n3923 ), .CK(clk), 
        .Q(out[320]), .QN() );
  DFF_X2 _f_permutation__out_reg_1463_  ( .D(_f_permutation__n3924 ), .CK(clk), 
        .Q(out[335]), .QN() );
  DFF_X2 _f_permutation__out_reg_1462_  ( .D(_f_permutation__n3925 ), .CK(clk), 
        .Q(out[334]), .QN() );
  DFF_X2 _f_permutation__out_reg_1461_  ( .D(_f_permutation__n3926 ), .CK(clk), 
        .Q(out[333]), .QN() );
  DFF_X2 _f_permutation__out_reg_1460_  ( .D(_f_permutation__n3927 ), .CK(clk), 
        .Q(out[332]), .QN() );
  DFF_X2 _f_permutation__out_reg_1459_  ( .D(_f_permutation__n3928 ), .CK(clk), 
        .Q(out[331]), .QN() );
  DFF_X2 _f_permutation__out_reg_1458_  ( .D(_f_permutation__n3929 ), .CK(clk), 
        .Q(out[330]), .QN() );
  DFF_X2 _f_permutation__out_reg_1457_  ( .D(_f_permutation__n3930 ), .CK(clk), 
        .Q(out[329]), .QN() );
  DFF_X2 _f_permutation__out_reg_1456_  ( .D(_f_permutation__n3931 ), .CK(clk), 
        .Q(out[328]), .QN() );
  DFF_X2 _f_permutation__out_reg_1455_  ( .D(_f_permutation__n3932 ), .CK(clk), 
        .Q(out[343]), .QN() );
  DFF_X2 _f_permutation__out_reg_1454_  ( .D(_f_permutation__n3933 ), .CK(clk), 
        .Q(out[342]), .QN() );
  DFF_X2 _f_permutation__out_reg_1453_  ( .D(_f_permutation__n3934 ), .CK(clk), 
        .Q(out[341]), .QN() );
  DFF_X2 _f_permutation__out_reg_1452_  ( .D(_f_permutation__n3935 ), .CK(clk), 
        .Q(out[340]), .QN() );
  DFF_X2 _f_permutation__out_reg_1451_  ( .D(_f_permutation__n3936 ), .CK(clk), 
        .Q(out[339]), .QN() );
  DFF_X2 _f_permutation__out_reg_1450_  ( .D(_f_permutation__n3937 ), .CK(clk), 
        .Q(out[338]), .QN() );
  DFF_X2 _f_permutation__out_reg_1449_  ( .D(_f_permutation__n3938 ), .CK(clk), 
        .Q(out[337]), .QN() );
  DFF_X2 _f_permutation__out_reg_1448_  ( .D(_f_permutation__n3939 ), .CK(clk), 
        .Q(out[336]), .QN() );
  DFF_X2 _f_permutation__out_reg_1447_  ( .D(_f_permutation__n3940 ), .CK(clk), 
        .Q(out[351]), .QN() );
  DFF_X2 _f_permutation__out_reg_1446_  ( .D(_f_permutation__n3941 ), .CK(clk), 
        .Q(out[350]), .QN() );
  DFF_X2 _f_permutation__out_reg_1445_  ( .D(_f_permutation__n3942 ), .CK(clk), 
        .Q(out[349]), .QN() );
  DFF_X2 _f_permutation__out_reg_1444_  ( .D(_f_permutation__n3943 ), .CK(clk), 
        .Q(out[348]), .QN() );
  DFF_X2 _f_permutation__out_reg_1443_  ( .D(_f_permutation__n3944 ), .CK(clk), 
        .Q(out[347]), .QN() );
  DFF_X2 _f_permutation__out_reg_1442_  ( .D(_f_permutation__n3945 ), .CK(clk), 
        .Q(out[346]), .QN() );
  DFF_X2 _f_permutation__out_reg_1441_  ( .D(_f_permutation__n3946 ), .CK(clk), 
        .Q(out[345]), .QN() );
  DFF_X2 _f_permutation__out_reg_1440_  ( .D(_f_permutation__n3947 ), .CK(clk), 
        .Q(out[344]), .QN() );
  DFF_X2 _f_permutation__out_reg_1439_  ( .D(_f_permutation__n3948 ), .CK(clk), 
        .Q(out[359]), .QN() );
  DFF_X2 _f_permutation__out_reg_1438_  ( .D(_f_permutation__n3949 ), .CK(clk), 
        .Q(out[358]), .QN() );
  DFF_X2 _f_permutation__out_reg_1437_  ( .D(_f_permutation__n3950 ), .CK(clk), 
        .Q(out[357]), .QN() );
  DFF_X2 _f_permutation__out_reg_1436_  ( .D(_f_permutation__n3951 ), .CK(clk), 
        .Q(out[356]), .QN() );
  DFF_X2 _f_permutation__out_reg_1435_  ( .D(_f_permutation__n3952 ), .CK(clk), 
        .Q(out[355]), .QN() );
  DFF_X2 _f_permutation__out_reg_1434_  ( .D(_f_permutation__n3953 ), .CK(clk), 
        .Q(out[354]), .QN() );
  DFF_X2 _f_permutation__out_reg_1433_  ( .D(_f_permutation__n3954 ), .CK(clk), 
        .Q(out[353]), .QN() );
  DFF_X2 _f_permutation__out_reg_1432_  ( .D(_f_permutation__n3955 ), .CK(clk), 
        .Q(out[352]), .QN() );
  DFF_X2 _f_permutation__out_reg_1431_  ( .D(_f_permutation__n3956 ), .CK(clk), 
        .Q(out[367]), .QN() );
  DFF_X2 _f_permutation__out_reg_1430_  ( .D(_f_permutation__n3957 ), .CK(clk), 
        .Q(out[366]), .QN() );
  DFF_X2 _f_permutation__out_reg_1429_  ( .D(_f_permutation__n3958 ), .CK(clk), 
        .Q(out[365]), .QN() );
  DFF_X2 _f_permutation__out_reg_1428_  ( .D(_f_permutation__n3959 ), .CK(clk), 
        .Q(out[364]), .QN() );
  DFF_X2 _f_permutation__out_reg_1427_  ( .D(_f_permutation__n3960 ), .CK(clk), 
        .Q(out[363]), .QN() );
  DFF_X2 _f_permutation__out_reg_1426_  ( .D(_f_permutation__n3961 ), .CK(clk), 
        .Q(out[362]), .QN() );
  DFF_X2 _f_permutation__out_reg_1425_  ( .D(_f_permutation__n3962 ), .CK(clk), 
        .Q(out[361]), .QN() );
  DFF_X2 _f_permutation__out_reg_1424_  ( .D(_f_permutation__n3963 ), .CK(clk), 
        .Q(out[360]), .QN() );
  DFF_X2 _f_permutation__out_reg_1423_  ( .D(_f_permutation__n3964 ), .CK(clk), 
        .Q(out[375]), .QN() );
  DFF_X2 _f_permutation__out_reg_1422_  ( .D(_f_permutation__n3965 ), .CK(clk), 
        .Q(out[374]), .QN() );
  DFF_X2 _f_permutation__out_reg_1421_  ( .D(_f_permutation__n3966 ), .CK(clk), 
        .Q(out[373]), .QN() );
  DFF_X2 _f_permutation__out_reg_1420_  ( .D(_f_permutation__n3967 ), .CK(clk), 
        .Q(out[372]), .QN() );
  DFF_X2 _f_permutation__out_reg_1419_  ( .D(_f_permutation__n3968 ), .CK(clk), 
        .Q(out[371]), .QN() );
  DFF_X2 _f_permutation__out_reg_1418_  ( .D(_f_permutation__n3969 ), .CK(clk), 
        .Q(out[370]), .QN() );
  DFF_X2 _f_permutation__out_reg_1417_  ( .D(_f_permutation__n3970 ), .CK(clk), 
        .Q(out[369]), .QN() );
  DFF_X2 _f_permutation__out_reg_1416_  ( .D(_f_permutation__n3971 ), .CK(clk), 
        .Q(out[368]), .QN() );
  DFF_X2 _f_permutation__out_reg_1415_  ( .D(_f_permutation__n3972 ), .CK(clk), 
        .Q(out[383]), .QN() );
  DFF_X2 _f_permutation__out_reg_1414_  ( .D(_f_permutation__n3973 ), .CK(clk), 
        .Q(out[382]), .QN() );
  DFF_X2 _f_permutation__out_reg_1413_  ( .D(_f_permutation__n3974 ), .CK(clk), 
        .Q(out[381]), .QN() );
  DFF_X2 _f_permutation__out_reg_1412_  ( .D(_f_permutation__n3975 ), .CK(clk), 
        .Q(out[380]), .QN() );
  DFF_X2 _f_permutation__out_reg_1411_  ( .D(_f_permutation__n3976 ), .CK(clk), 
        .Q(out[379]), .QN() );
  DFF_X2 _f_permutation__out_reg_1410_  ( .D(_f_permutation__n3977 ), .CK(clk), 
        .Q(out[378]), .QN() );
  DFF_X2 _f_permutation__out_reg_1409_  ( .D(_f_permutation__n3978 ), .CK(clk), 
        .Q(out[377]), .QN() );
  DFF_X2 _f_permutation__out_reg_1408_  ( .D(_f_permutation__n3979 ), .CK(clk), 
        .Q(out[376]), .QN() );
  DFF_X2 _f_permutation__out_reg_1407_  ( .D(_f_permutation__n3980 ), .CK(clk), 
        .Q(out[263]), .QN() );
  DFF_X2 _f_permutation__out_reg_1406_  ( .D(_f_permutation__n3981 ), .CK(clk), 
        .Q(out[262]), .QN() );
  DFF_X2 _f_permutation__out_reg_1405_  ( .D(_f_permutation__n3982 ), .CK(clk), 
        .Q(out[261]), .QN() );
  DFF_X2 _f_permutation__out_reg_1404_  ( .D(_f_permutation__n3983 ), .CK(clk), 
        .Q(out[260]), .QN() );
  DFF_X2 _f_permutation__out_reg_1403_  ( .D(_f_permutation__n3984 ), .CK(clk), 
        .Q(out[259]), .QN() );
  DFF_X2 _f_permutation__out_reg_1402_  ( .D(_f_permutation__n3985 ), .CK(clk), 
        .Q(out[258]), .QN() );
  DFF_X2 _f_permutation__out_reg_1401_  ( .D(_f_permutation__n3986 ), .CK(clk), 
        .Q(out[257]), .QN() );
  DFF_X2 _f_permutation__out_reg_1400_  ( .D(_f_permutation__n3987 ), .CK(clk), 
        .Q(out[256]), .QN() );
  DFF_X2 _f_permutation__out_reg_1399_  ( .D(_f_permutation__n3988 ), .CK(clk), 
        .Q(out[271]), .QN() );
  DFF_X2 _f_permutation__out_reg_1398_  ( .D(_f_permutation__n3989 ), .CK(clk), 
        .Q(out[270]), .QN() );
  DFF_X2 _f_permutation__out_reg_1397_  ( .D(_f_permutation__n3990 ), .CK(clk), 
        .Q(out[269]), .QN() );
  DFF_X2 _f_permutation__out_reg_1396_  ( .D(_f_permutation__n3991 ), .CK(clk), 
        .Q(out[268]), .QN() );
  DFF_X2 _f_permutation__out_reg_1395_  ( .D(_f_permutation__n3992 ), .CK(clk), 
        .Q(out[267]), .QN() );
  DFF_X2 _f_permutation__out_reg_1394_  ( .D(_f_permutation__n3993 ), .CK(clk), 
        .Q(out[266]), .QN() );
  DFF_X2 _f_permutation__out_reg_1393_  ( .D(_f_permutation__n3994 ), .CK(clk), 
        .Q(out[265]), .QN() );
  DFF_X2 _f_permutation__out_reg_1392_  ( .D(_f_permutation__n3995 ), .CK(clk), 
        .Q(out[264]), .QN() );
  DFF_X2 _f_permutation__out_reg_1391_  ( .D(_f_permutation__n3996 ), .CK(clk), 
        .Q(out[279]), .QN() );
  DFF_X2 _f_permutation__out_reg_1390_  ( .D(_f_permutation__n3997 ), .CK(clk), 
        .Q(out[278]), .QN() );
  DFF_X2 _f_permutation__out_reg_1389_  ( .D(_f_permutation__n3998 ), .CK(clk), 
        .Q(out[277]), .QN() );
  DFF_X2 _f_permutation__out_reg_1388_  ( .D(_f_permutation__n3999 ), .CK(clk), 
        .Q(out[276]), .QN() );
  DFF_X2 _f_permutation__out_reg_1387_  ( .D(_f_permutation__n4000 ), .CK(clk), 
        .Q(out[275]), .QN() );
  DFF_X2 _f_permutation__out_reg_1386_  ( .D(_f_permutation__n4001 ), .CK(clk), 
        .Q(out[274]), .QN() );
  DFF_X2 _f_permutation__out_reg_1385_  ( .D(_f_permutation__n4002 ), .CK(clk), 
        .Q(out[273]), .QN() );
  DFF_X2 _f_permutation__out_reg_1384_  ( .D(_f_permutation__n4003 ), .CK(clk), 
        .Q(out[272]), .QN() );
  DFF_X2 _f_permutation__out_reg_1383_  ( .D(_f_permutation__n4004 ), .CK(clk), 
        .Q(out[287]), .QN() );
  DFF_X2 _f_permutation__out_reg_1382_  ( .D(_f_permutation__n4005 ), .CK(clk), 
        .Q(out[286]), .QN() );
  DFF_X2 _f_permutation__out_reg_1381_  ( .D(_f_permutation__n4006 ), .CK(clk), 
        .Q(out[285]), .QN() );
  DFF_X2 _f_permutation__out_reg_1380_  ( .D(_f_permutation__n4007 ), .CK(clk), 
        .Q(out[284]), .QN() );
  DFF_X2 _f_permutation__out_reg_1379_  ( .D(_f_permutation__n4008 ), .CK(clk), 
        .Q(out[283]), .QN() );
  DFF_X2 _f_permutation__out_reg_1378_  ( .D(_f_permutation__n4009 ), .CK(clk), 
        .Q(out[282]), .QN() );
  DFF_X2 _f_permutation__out_reg_1377_  ( .D(_f_permutation__n4010 ), .CK(clk), 
        .Q(out[281]), .QN() );
  DFF_X2 _f_permutation__out_reg_1376_  ( .D(_f_permutation__n4011 ), .CK(clk), 
        .Q(out[280]), .QN() );
  DFF_X2 _f_permutation__out_reg_1375_  ( .D(_f_permutation__n4012 ), .CK(clk), 
        .Q(out[295]), .QN() );
  DFF_X2 _f_permutation__out_reg_1374_  ( .D(_f_permutation__n4013 ), .CK(clk), 
        .Q(out[294]), .QN() );
  DFF_X2 _f_permutation__out_reg_1373_  ( .D(_f_permutation__n4014 ), .CK(clk), 
        .Q(out[293]), .QN() );
  DFF_X2 _f_permutation__out_reg_1372_  ( .D(_f_permutation__n4015 ), .CK(clk), 
        .Q(out[292]), .QN() );
  DFF_X2 _f_permutation__out_reg_1371_  ( .D(_f_permutation__n4016 ), .CK(clk), 
        .Q(out[291]), .QN() );
  DFF_X2 _f_permutation__out_reg_1370_  ( .D(_f_permutation__n4017 ), .CK(clk), 
        .Q(out[290]), .QN() );
  DFF_X2 _f_permutation__out_reg_1369_  ( .D(_f_permutation__n4018 ), .CK(clk), 
        .Q(out[289]), .QN() );
  DFF_X2 _f_permutation__out_reg_1368_  ( .D(_f_permutation__n4019 ), .CK(clk), 
        .Q(out[288]), .QN() );
  DFF_X2 _f_permutation__out_reg_1367_  ( .D(_f_permutation__n4020 ), .CK(clk), 
        .Q(out[303]), .QN() );
  DFF_X2 _f_permutation__out_reg_1366_  ( .D(_f_permutation__n4021 ), .CK(clk), 
        .Q(out[302]), .QN() );
  DFF_X2 _f_permutation__out_reg_1365_  ( .D(_f_permutation__n4022 ), .CK(clk), 
        .Q(out[301]), .QN() );
  DFF_X2 _f_permutation__out_reg_1364_  ( .D(_f_permutation__n4023 ), .CK(clk), 
        .Q(out[300]), .QN() );
  DFF_X2 _f_permutation__out_reg_1363_  ( .D(_f_permutation__n4024 ), .CK(clk), 
        .Q(out[299]), .QN() );
  DFF_X2 _f_permutation__out_reg_1362_  ( .D(_f_permutation__n4025 ), .CK(clk), 
        .Q(out[298]), .QN() );
  DFF_X2 _f_permutation__out_reg_1361_  ( .D(_f_permutation__n4026 ), .CK(clk), 
        .Q(out[297]), .QN() );
  DFF_X2 _f_permutation__out_reg_1360_  ( .D(_f_permutation__n4027 ), .CK(clk), 
        .Q(out[296]), .QN() );
  DFF_X2 _f_permutation__out_reg_1359_  ( .D(_f_permutation__n4028 ), .CK(clk), 
        .Q(out[311]), .QN() );
  DFF_X2 _f_permutation__out_reg_1358_  ( .D(_f_permutation__n4029 ), .CK(clk), 
        .Q(out[310]), .QN() );
  DFF_X2 _f_permutation__out_reg_1357_  ( .D(_f_permutation__n4030 ), .CK(clk), 
        .Q(out[309]), .QN() );
  DFF_X2 _f_permutation__out_reg_1356_  ( .D(_f_permutation__n4031 ), .CK(clk), 
        .Q(out[308]), .QN() );
  DFF_X2 _f_permutation__out_reg_1355_  ( .D(_f_permutation__n4032 ), .CK(clk), 
        .Q(out[307]), .QN() );
  DFF_X2 _f_permutation__out_reg_1354_  ( .D(_f_permutation__n4033 ), .CK(clk), 
        .Q(out[306]), .QN() );
  DFF_X2 _f_permutation__out_reg_1353_  ( .D(_f_permutation__n4034 ), .CK(clk), 
        .Q(out[305]), .QN() );
  DFF_X2 _f_permutation__out_reg_1352_  ( .D(_f_permutation__n4035 ), .CK(clk), 
        .Q(out[304]), .QN() );
  DFF_X2 _f_permutation__out_reg_1351_  ( .D(_f_permutation__n4036 ), .CK(clk), 
        .Q(out[319]), .QN() );
  DFF_X2 _f_permutation__out_reg_1350_  ( .D(_f_permutation__n4037 ), .CK(clk), 
        .Q(out[318]), .QN() );
  DFF_X2 _f_permutation__out_reg_1349_  ( .D(_f_permutation__n4038 ), .CK(clk), 
        .Q(out[317]), .QN() );
  DFF_X2 _f_permutation__out_reg_1348_  ( .D(_f_permutation__n4039 ), .CK(clk), 
        .Q(out[316]), .QN() );
  DFF_X2 _f_permutation__out_reg_1347_  ( .D(_f_permutation__n4040 ), .CK(clk), 
        .Q(out[315]), .QN() );
  DFF_X2 _f_permutation__out_reg_1346_  ( .D(_f_permutation__n4041 ), .CK(clk), 
        .Q(out[314]), .QN() );
  DFF_X2 _f_permutation__out_reg_1345_  ( .D(_f_permutation__n4042 ), .CK(clk), 
        .Q(out[313]), .QN() );
  DFF_X2 _f_permutation__out_reg_1344_  ( .D(_f_permutation__n4043 ), .CK(clk), 
        .Q(out[312]), .QN() );
  DFF_X2 _f_permutation__out_reg_1343_  ( .D(_f_permutation__n4044 ), .CK(clk), 
        .Q(out[199]), .QN() );
  DFF_X2 _f_permutation__out_reg_1342_  ( .D(_f_permutation__n4045 ), .CK(clk), 
        .Q(out[198]), .QN() );
  DFF_X2 _f_permutation__out_reg_1341_  ( .D(_f_permutation__n4046 ), .CK(clk), 
        .Q(out[197]), .QN() );
  DFF_X2 _f_permutation__out_reg_1340_  ( .D(_f_permutation__n4047 ), .CK(clk), 
        .Q(out[196]), .QN() );
  DFF_X2 _f_permutation__out_reg_1339_  ( .D(_f_permutation__n4048 ), .CK(clk), 
        .Q(out[195]), .QN() );
  DFF_X2 _f_permutation__out_reg_1338_  ( .D(_f_permutation__n4049 ), .CK(clk), 
        .Q(out[194]), .QN() );
  DFF_X2 _f_permutation__out_reg_1337_  ( .D(_f_permutation__n4050 ), .CK(clk), 
        .Q(out[193]), .QN() );
  DFF_X2 _f_permutation__out_reg_1336_  ( .D(_f_permutation__n4051 ), .CK(clk), 
        .Q(out[192]), .QN() );
  DFF_X2 _f_permutation__out_reg_1335_  ( .D(_f_permutation__n4052 ), .CK(clk), 
        .Q(out[207]), .QN() );
  DFF_X2 _f_permutation__out_reg_1334_  ( .D(_f_permutation__n4053 ), .CK(clk), 
        .Q(out[206]), .QN() );
  DFF_X2 _f_permutation__out_reg_1333_  ( .D(_f_permutation__n4054 ), .CK(clk), 
        .Q(out[205]), .QN() );
  DFF_X2 _f_permutation__out_reg_1332_  ( .D(_f_permutation__n4055 ), .CK(clk), 
        .Q(out[204]), .QN() );
  DFF_X2 _f_permutation__out_reg_1331_  ( .D(_f_permutation__n4056 ), .CK(clk), 
        .Q(out[203]), .QN() );
  DFF_X2 _f_permutation__out_reg_1330_  ( .D(_f_permutation__n4057 ), .CK(clk), 
        .Q(out[202]), .QN() );
  DFF_X2 _f_permutation__out_reg_1329_  ( .D(_f_permutation__n4058 ), .CK(clk), 
        .Q(out[201]), .QN() );
  DFF_X2 _f_permutation__out_reg_1328_  ( .D(_f_permutation__n4059 ), .CK(clk), 
        .Q(out[200]), .QN() );
  DFF_X2 _f_permutation__out_reg_1327_  ( .D(_f_permutation__n4060 ), .CK(clk), 
        .Q(out[215]), .QN() );
  DFF_X2 _f_permutation__out_reg_1326_  ( .D(_f_permutation__n4061 ), .CK(clk), 
        .Q(out[214]), .QN() );
  DFF_X2 _f_permutation__out_reg_1325_  ( .D(_f_permutation__n4062 ), .CK(clk), 
        .Q(out[213]), .QN() );
  DFF_X2 _f_permutation__out_reg_1324_  ( .D(_f_permutation__n4063 ), .CK(clk), 
        .Q(out[212]), .QN() );
  DFF_X2 _f_permutation__out_reg_1323_  ( .D(_f_permutation__n4064 ), .CK(clk), 
        .Q(out[211]), .QN() );
  DFF_X2 _f_permutation__out_reg_1322_  ( .D(_f_permutation__n4065 ), .CK(clk), 
        .Q(out[210]), .QN() );
  DFF_X2 _f_permutation__out_reg_1321_  ( .D(_f_permutation__n4066 ), .CK(clk), 
        .Q(out[209]), .QN() );
  DFF_X2 _f_permutation__out_reg_1320_  ( .D(_f_permutation__n4067 ), .CK(clk), 
        .Q(out[208]), .QN() );
  DFF_X2 _f_permutation__out_reg_1319_  ( .D(_f_permutation__n4068 ), .CK(clk), 
        .Q(out[223]), .QN() );
  DFF_X2 _f_permutation__out_reg_1318_  ( .D(_f_permutation__n4069 ), .CK(clk), 
        .Q(out[222]), .QN() );
  DFF_X2 _f_permutation__out_reg_1317_  ( .D(_f_permutation__n4070 ), .CK(clk), 
        .Q(out[221]), .QN() );
  DFF_X2 _f_permutation__out_reg_1316_  ( .D(_f_permutation__n4071 ), .CK(clk), 
        .Q(out[220]), .QN() );
  DFF_X2 _f_permutation__out_reg_1315_  ( .D(_f_permutation__n4072 ), .CK(clk), 
        .Q(out[219]), .QN() );
  DFF_X2 _f_permutation__out_reg_1314_  ( .D(_f_permutation__n4073 ), .CK(clk), 
        .Q(out[218]), .QN() );
  DFF_X2 _f_permutation__out_reg_1313_  ( .D(_f_permutation__n4074 ), .CK(clk), 
        .Q(out[217]), .QN() );
  DFF_X2 _f_permutation__out_reg_1312_  ( .D(_f_permutation__n4075 ), .CK(clk), 
        .Q(out[216]), .QN() );
  DFF_X2 _f_permutation__out_reg_1311_  ( .D(_f_permutation__n4076 ), .CK(clk), 
        .Q(out[231]), .QN() );
  DFF_X2 _f_permutation__out_reg_1310_  ( .D(_f_permutation__n4077 ), .CK(clk), 
        .Q(out[230]), .QN() );
  DFF_X2 _f_permutation__out_reg_1309_  ( .D(_f_permutation__n4078 ), .CK(clk), 
        .Q(out[229]), .QN() );
  DFF_X2 _f_permutation__out_reg_1308_  ( .D(_f_permutation__n4079 ), .CK(clk), 
        .Q(out[228]), .QN() );
  DFF_X2 _f_permutation__out_reg_1307_  ( .D(_f_permutation__n4080 ), .CK(clk), 
        .Q(out[227]), .QN() );
  DFF_X2 _f_permutation__out_reg_1306_  ( .D(_f_permutation__n4081 ), .CK(clk), 
        .Q(out[226]), .QN() );
  DFF_X2 _f_permutation__out_reg_1305_  ( .D(_f_permutation__n4082 ), .CK(clk), 
        .Q(out[225]), .QN() );
  DFF_X2 _f_permutation__out_reg_1304_  ( .D(_f_permutation__n4083 ), .CK(clk), 
        .Q(out[224]), .QN() );
  DFF_X2 _f_permutation__out_reg_1303_  ( .D(_f_permutation__n4084 ), .CK(clk), 
        .Q(out[239]), .QN() );
  DFF_X2 _f_permutation__out_reg_1302_  ( .D(_f_permutation__n4085 ), .CK(clk), 
        .Q(out[238]), .QN() );
  DFF_X2 _f_permutation__out_reg_1301_  ( .D(_f_permutation__n4086 ), .CK(clk), 
        .Q(out[237]), .QN() );
  DFF_X2 _f_permutation__out_reg_1300_  ( .D(_f_permutation__n4087 ), .CK(clk), 
        .Q(out[236]), .QN() );
  DFF_X2 _f_permutation__out_reg_1299_  ( .D(_f_permutation__n4088 ), .CK(clk), 
        .Q(out[235]), .QN() );
  DFF_X2 _f_permutation__out_reg_1298_  ( .D(_f_permutation__n4089 ), .CK(clk), 
        .Q(out[234]), .QN() );
  DFF_X2 _f_permutation__out_reg_1297_  ( .D(_f_permutation__n4090 ), .CK(clk), 
        .Q(out[233]), .QN() );
  DFF_X2 _f_permutation__out_reg_1296_  ( .D(_f_permutation__n4091 ), .CK(clk), 
        .Q(out[232]), .QN() );
  DFF_X2 _f_permutation__out_reg_1295_  ( .D(_f_permutation__n4092 ), .CK(clk), 
        .Q(out[247]), .QN() );
  DFF_X2 _f_permutation__out_reg_1294_  ( .D(_f_permutation__n4093 ), .CK(clk), 
        .Q(out[246]), .QN() );
  DFF_X2 _f_permutation__out_reg_1293_  ( .D(_f_permutation__n4094 ), .CK(clk), 
        .Q(out[245]), .QN() );
  DFF_X2 _f_permutation__out_reg_1292_  ( .D(_f_permutation__n4095 ), .CK(clk), 
        .Q(out[244]), .QN() );
  DFF_X2 _f_permutation__out_reg_1291_  ( .D(_f_permutation__n4096 ), .CK(clk), 
        .Q(out[243]), .QN() );
  DFF_X2 _f_permutation__out_reg_1290_  ( .D(_f_permutation__n4097 ), .CK(clk), 
        .Q(out[242]), .QN() );
  DFF_X2 _f_permutation__out_reg_1289_  ( .D(_f_permutation__n4098 ), .CK(clk), 
        .Q(out[241]), .QN() );
  DFF_X2 _f_permutation__out_reg_1288_  ( .D(_f_permutation__n4099 ), .CK(clk), 
        .Q(out[240]), .QN() );
  DFF_X2 _f_permutation__out_reg_1287_  ( .D(_f_permutation__n4100 ), .CK(clk), 
        .Q(out[255]), .QN() );
  DFF_X2 _f_permutation__out_reg_1286_  ( .D(_f_permutation__n4101 ), .CK(clk), 
        .Q(out[254]), .QN() );
  DFF_X2 _f_permutation__out_reg_1285_  ( .D(_f_permutation__n4102 ), .CK(clk), 
        .Q(out[253]), .QN() );
  DFF_X2 _f_permutation__out_reg_1284_  ( .D(_f_permutation__n4103 ), .CK(clk), 
        .Q(out[252]), .QN() );
  DFF_X2 _f_permutation__out_reg_1283_  ( .D(_f_permutation__n4104 ), .CK(clk), 
        .Q(out[251]), .QN() );
  DFF_X2 _f_permutation__out_reg_1282_  ( .D(_f_permutation__n4105 ), .CK(clk), 
        .Q(out[250]), .QN() );
  DFF_X2 _f_permutation__out_reg_1281_  ( .D(_f_permutation__n4106 ), .CK(clk), 
        .Q(out[249]), .QN() );
  DFF_X2 _f_permutation__out_reg_1280_  ( .D(_f_permutation__n4107 ), .CK(clk), 
        .Q(out[248]), .QN() );
  DFF_X2 _f_permutation__out_reg_1279_  ( .D(_f_permutation__n4108 ), .CK(clk), 
        .Q(out[135]), .QN() );
  DFF_X2 _f_permutation__out_reg_1278_  ( .D(_f_permutation__n4109 ), .CK(clk), 
        .Q(out[134]), .QN() );
  DFF_X2 _f_permutation__out_reg_1277_  ( .D(_f_permutation__n4110 ), .CK(clk), 
        .Q(out[133]), .QN() );
  DFF_X2 _f_permutation__out_reg_1276_  ( .D(_f_permutation__n4111 ), .CK(clk), 
        .Q(out[132]), .QN() );
  DFF_X2 _f_permutation__out_reg_1275_  ( .D(_f_permutation__n4112 ), .CK(clk), 
        .Q(out[131]), .QN() );
  DFF_X2 _f_permutation__out_reg_1274_  ( .D(_f_permutation__n4113 ), .CK(clk), 
        .Q(out[130]), .QN() );
  DFF_X2 _f_permutation__out_reg_1273_  ( .D(_f_permutation__n4114 ), .CK(clk), 
        .Q(out[129]), .QN() );
  DFF_X2 _f_permutation__out_reg_1272_  ( .D(_f_permutation__n4115 ), .CK(clk), 
        .Q(out[128]), .QN() );
  DFF_X2 _f_permutation__out_reg_1271_  ( .D(_f_permutation__n4116 ), .CK(clk), 
        .Q(out[143]), .QN() );
  DFF_X2 _f_permutation__out_reg_1270_  ( .D(_f_permutation__n4117 ), .CK(clk), 
        .Q(out[142]), .QN() );
  DFF_X2 _f_permutation__out_reg_1269_  ( .D(_f_permutation__n4118 ), .CK(clk), 
        .Q(out[141]), .QN() );
  DFF_X2 _f_permutation__out_reg_1268_  ( .D(_f_permutation__n4119 ), .CK(clk), 
        .Q(out[140]), .QN() );
  DFF_X2 _f_permutation__out_reg_1267_  ( .D(_f_permutation__n4120 ), .CK(clk), 
        .Q(out[139]), .QN() );
  DFF_X2 _f_permutation__out_reg_1266_  ( .D(_f_permutation__n4121 ), .CK(clk), 
        .Q(out[138]), .QN() );
  DFF_X2 _f_permutation__out_reg_1265_  ( .D(_f_permutation__n4122 ), .CK(clk), 
        .Q(out[137]), .QN() );
  DFF_X2 _f_permutation__out_reg_1264_  ( .D(_f_permutation__n4123 ), .CK(clk), 
        .Q(out[136]), .QN() );
  DFF_X2 _f_permutation__out_reg_1263_  ( .D(_f_permutation__n4124 ), .CK(clk), 
        .Q(out[151]), .QN() );
  DFF_X2 _f_permutation__out_reg_1262_  ( .D(_f_permutation__n4125 ), .CK(clk), 
        .Q(out[150]), .QN() );
  DFF_X2 _f_permutation__out_reg_1261_  ( .D(_f_permutation__n4126 ), .CK(clk), 
        .Q(out[149]), .QN() );
  DFF_X2 _f_permutation__out_reg_1260_  ( .D(_f_permutation__n4127 ), .CK(clk), 
        .Q(out[148]), .QN() );
  DFF_X2 _f_permutation__out_reg_1259_  ( .D(_f_permutation__n4128 ), .CK(clk), 
        .Q(out[147]), .QN() );
  DFF_X2 _f_permutation__out_reg_1258_  ( .D(_f_permutation__n4129 ), .CK(clk), 
        .Q(out[146]), .QN() );
  DFF_X2 _f_permutation__out_reg_1257_  ( .D(_f_permutation__n4130 ), .CK(clk), 
        .Q(out[145]), .QN() );
  DFF_X2 _f_permutation__out_reg_1256_  ( .D(_f_permutation__n4131 ), .CK(clk), 
        .Q(out[144]), .QN() );
  DFF_X2 _f_permutation__out_reg_1255_  ( .D(_f_permutation__n4132 ), .CK(clk), 
        .Q(out[159]), .QN() );
  DFF_X2 _f_permutation__out_reg_1254_  ( .D(_f_permutation__n4133 ), .CK(clk), 
        .Q(out[158]), .QN() );
  DFF_X2 _f_permutation__out_reg_1253_  ( .D(_f_permutation__n4134 ), .CK(clk), 
        .Q(out[157]), .QN() );
  DFF_X2 _f_permutation__out_reg_1252_  ( .D(_f_permutation__n4135 ), .CK(clk), 
        .Q(out[156]), .QN() );
  DFF_X2 _f_permutation__out_reg_1251_  ( .D(_f_permutation__n4136 ), .CK(clk), 
        .Q(out[155]), .QN() );
  DFF_X2 _f_permutation__out_reg_1250_  ( .D(_f_permutation__n4137 ), .CK(clk), 
        .Q(out[154]), .QN() );
  DFF_X2 _f_permutation__out_reg_1249_  ( .D(_f_permutation__n4138 ), .CK(clk), 
        .Q(out[153]), .QN() );
  DFF_X2 _f_permutation__out_reg_1248_  ( .D(_f_permutation__n4139 ), .CK(clk), 
        .Q(out[152]), .QN() );
  DFF_X2 _f_permutation__out_reg_1247_  ( .D(_f_permutation__n4140 ), .CK(clk), 
        .Q(out[167]), .QN() );
  DFF_X2 _f_permutation__out_reg_1246_  ( .D(_f_permutation__n4141 ), .CK(clk), 
        .Q(out[166]), .QN() );
  DFF_X2 _f_permutation__out_reg_1245_  ( .D(_f_permutation__n4142 ), .CK(clk), 
        .Q(out[165]), .QN() );
  DFF_X2 _f_permutation__out_reg_1244_  ( .D(_f_permutation__n4143 ), .CK(clk), 
        .Q(out[164]), .QN() );
  DFF_X2 _f_permutation__out_reg_1243_  ( .D(_f_permutation__n4144 ), .CK(clk), 
        .Q(out[163]), .QN() );
  DFF_X2 _f_permutation__out_reg_1242_  ( .D(_f_permutation__n4145 ), .CK(clk), 
        .Q(out[162]), .QN() );
  DFF_X2 _f_permutation__out_reg_1241_  ( .D(_f_permutation__n4146 ), .CK(clk), 
        .Q(out[161]), .QN() );
  DFF_X2 _f_permutation__out_reg_1240_  ( .D(_f_permutation__n4147 ), .CK(clk), 
        .Q(out[160]), .QN() );
  DFF_X2 _f_permutation__out_reg_1239_  ( .D(_f_permutation__n4148 ), .CK(clk), 
        .Q(out[175]), .QN() );
  DFF_X2 _f_permutation__out_reg_1238_  ( .D(_f_permutation__n4149 ), .CK(clk), 
        .Q(out[174]), .QN() );
  DFF_X2 _f_permutation__out_reg_1237_  ( .D(_f_permutation__n4150 ), .CK(clk), 
        .Q(out[173]), .QN() );
  DFF_X2 _f_permutation__out_reg_1236_  ( .D(_f_permutation__n4151 ), .CK(clk), 
        .Q(out[172]), .QN() );
  DFF_X2 _f_permutation__out_reg_1235_  ( .D(_f_permutation__n4152 ), .CK(clk), 
        .Q(out[171]), .QN() );
  DFF_X2 _f_permutation__out_reg_1234_  ( .D(_f_permutation__n4153 ), .CK(clk), 
        .Q(out[170]), .QN() );
  DFF_X2 _f_permutation__out_reg_1233_  ( .D(_f_permutation__n4154 ), .CK(clk), 
        .Q(out[169]), .QN() );
  DFF_X2 _f_permutation__out_reg_1232_  ( .D(_f_permutation__n4155 ), .CK(clk), 
        .Q(out[168]), .QN() );
  DFF_X2 _f_permutation__out_reg_1231_  ( .D(_f_permutation__n4156 ), .CK(clk), 
        .Q(out[183]), .QN() );
  DFF_X2 _f_permutation__out_reg_1230_  ( .D(_f_permutation__n4157 ), .CK(clk), 
        .Q(out[182]), .QN() );
  DFF_X2 _f_permutation__out_reg_1229_  ( .D(_f_permutation__n4158 ), .CK(clk), 
        .Q(out[181]), .QN() );
  DFF_X2 _f_permutation__out_reg_1228_  ( .D(_f_permutation__n4159 ), .CK(clk), 
        .Q(out[180]), .QN() );
  DFF_X2 _f_permutation__out_reg_1227_  ( .D(_f_permutation__n4160 ), .CK(clk), 
        .Q(out[179]), .QN() );
  DFF_X2 _f_permutation__out_reg_1226_  ( .D(_f_permutation__n4161 ), .CK(clk), 
        .Q(out[178]), .QN() );
  DFF_X2 _f_permutation__out_reg_1225_  ( .D(_f_permutation__n4162 ), .CK(clk), 
        .Q(out[177]), .QN() );
  DFF_X2 _f_permutation__out_reg_1224_  ( .D(_f_permutation__n4163 ), .CK(clk), 
        .Q(out[176]), .QN() );
  DFF_X2 _f_permutation__out_reg_1223_  ( .D(_f_permutation__n4164 ), .CK(clk), 
        .Q(out[191]), .QN() );
  DFF_X2 _f_permutation__out_reg_1222_  ( .D(_f_permutation__n4165 ), .CK(clk), 
        .Q(out[190]), .QN() );
  DFF_X2 _f_permutation__out_reg_1221_  ( .D(_f_permutation__n4166 ), .CK(clk), 
        .Q(out[189]), .QN() );
  DFF_X2 _f_permutation__out_reg_1220_  ( .D(_f_permutation__n4167 ), .CK(clk), 
        .Q(out[188]), .QN() );
  DFF_X2 _f_permutation__out_reg_1219_  ( .D(_f_permutation__n4168 ), .CK(clk), 
        .Q(out[187]), .QN() );
  DFF_X2 _f_permutation__out_reg_1218_  ( .D(_f_permutation__n4169 ), .CK(clk), 
        .Q(out[186]), .QN() );
  DFF_X2 _f_permutation__out_reg_1217_  ( .D(_f_permutation__n4170 ), .CK(clk), 
        .Q(out[185]), .QN() );
  DFF_X2 _f_permutation__out_reg_1216_  ( .D(_f_permutation__n4171 ), .CK(clk), 
        .Q(out[184]), .QN() );
  DFF_X2 _f_permutation__out_reg_1215_  ( .D(_f_permutation__n4172 ), .CK(clk), 
        .Q(out[71]), .QN() );
  DFF_X2 _f_permutation__out_reg_1214_  ( .D(_f_permutation__n4173 ), .CK(clk), 
        .Q(out[70]), .QN() );
  DFF_X2 _f_permutation__out_reg_1213_  ( .D(_f_permutation__n4174 ), .CK(clk), 
        .Q(out[69]), .QN() );
  DFF_X2 _f_permutation__out_reg_1212_  ( .D(_f_permutation__n4175 ), .CK(clk), 
        .Q(out[68]), .QN() );
  DFF_X2 _f_permutation__out_reg_1211_  ( .D(_f_permutation__n4176 ), .CK(clk), 
        .Q(out[67]), .QN() );
  DFF_X2 _f_permutation__out_reg_1210_  ( .D(_f_permutation__n4177 ), .CK(clk), 
        .Q(out[66]), .QN() );
  DFF_X2 _f_permutation__out_reg_1209_  ( .D(_f_permutation__n4178 ), .CK(clk), 
        .Q(out[65]), .QN() );
  DFF_X2 _f_permutation__out_reg_1208_  ( .D(_f_permutation__n4179 ), .CK(clk), 
        .Q(out[64]), .QN() );
  DFF_X2 _f_permutation__out_reg_1207_  ( .D(_f_permutation__n4180 ), .CK(clk), 
        .Q(out[79]), .QN() );
  DFF_X2 _f_permutation__out_reg_1206_  ( .D(_f_permutation__n4181 ), .CK(clk), 
        .Q(out[78]), .QN() );
  DFF_X2 _f_permutation__out_reg_1205_  ( .D(_f_permutation__n4182 ), .CK(clk), 
        .Q(out[77]), .QN() );
  DFF_X2 _f_permutation__out_reg_1204_  ( .D(_f_permutation__n4183 ), .CK(clk), 
        .Q(out[76]), .QN() );
  DFF_X2 _f_permutation__out_reg_1203_  ( .D(_f_permutation__n4184 ), .CK(clk), 
        .Q(out[75]), .QN() );
  DFF_X2 _f_permutation__out_reg_1202_  ( .D(_f_permutation__n4185 ), .CK(clk), 
        .Q(out[74]), .QN() );
  DFF_X2 _f_permutation__out_reg_1201_  ( .D(_f_permutation__n4186 ), .CK(clk), 
        .Q(out[73]), .QN() );
  DFF_X2 _f_permutation__out_reg_1200_  ( .D(_f_permutation__n4187 ), .CK(clk), 
        .Q(out[72]), .QN() );
  DFF_X2 _f_permutation__out_reg_1199_  ( .D(_f_permutation__n4188 ), .CK(clk), 
        .Q(out[87]), .QN() );
  DFF_X2 _f_permutation__out_reg_1198_  ( .D(_f_permutation__n4189 ), .CK(clk), 
        .Q(out[86]), .QN() );
  DFF_X2 _f_permutation__out_reg_1197_  ( .D(_f_permutation__n4190 ), .CK(clk), 
        .Q(out[85]), .QN() );
  DFF_X2 _f_permutation__out_reg_1196_  ( .D(_f_permutation__n4191 ), .CK(clk), 
        .Q(out[84]), .QN() );
  DFF_X2 _f_permutation__out_reg_1195_  ( .D(_f_permutation__n4192 ), .CK(clk), 
        .Q(out[83]), .QN() );
  DFF_X2 _f_permutation__out_reg_1194_  ( .D(_f_permutation__n4193 ), .CK(clk), 
        .Q(out[82]), .QN() );
  DFF_X2 _f_permutation__out_reg_1193_  ( .D(_f_permutation__n4194 ), .CK(clk), 
        .Q(out[81]), .QN() );
  DFF_X2 _f_permutation__out_reg_1192_  ( .D(_f_permutation__n4195 ), .CK(clk), 
        .Q(out[80]), .QN() );
  DFF_X2 _f_permutation__out_reg_1191_  ( .D(_f_permutation__n4196 ), .CK(clk), 
        .Q(out[95]), .QN() );
  DFF_X2 _f_permutation__out_reg_1190_  ( .D(_f_permutation__n4197 ), .CK(clk), 
        .Q(out[94]), .QN() );
  DFF_X2 _f_permutation__out_reg_1189_  ( .D(_f_permutation__n4198 ), .CK(clk), 
        .Q(out[93]), .QN() );
  DFF_X2 _f_permutation__out_reg_1188_  ( .D(_f_permutation__n4199 ), .CK(clk), 
        .Q(out[92]), .QN() );
  DFF_X2 _f_permutation__out_reg_1187_  ( .D(_f_permutation__n4200 ), .CK(clk), 
        .Q(out[91]), .QN() );
  DFF_X2 _f_permutation__out_reg_1186_  ( .D(_f_permutation__n4201 ), .CK(clk), 
        .Q(out[90]), .QN() );
  DFF_X2 _f_permutation__out_reg_1185_  ( .D(_f_permutation__n4202 ), .CK(clk), 
        .Q(out[89]), .QN() );
  DFF_X2 _f_permutation__out_reg_1184_  ( .D(_f_permutation__n4203 ), .CK(clk), 
        .Q(out[88]), .QN() );
  DFF_X2 _f_permutation__out_reg_1183_  ( .D(_f_permutation__n4204 ), .CK(clk), 
        .Q(out[103]), .QN() );
  DFF_X2 _f_permutation__out_reg_1182_  ( .D(_f_permutation__n4205 ), .CK(clk), 
        .Q(out[102]), .QN() );
  DFF_X2 _f_permutation__out_reg_1181_  ( .D(_f_permutation__n4206 ), .CK(clk), 
        .Q(out[101]), .QN() );
  DFF_X2 _f_permutation__out_reg_1180_  ( .D(_f_permutation__n4207 ), .CK(clk), 
        .Q(out[100]), .QN() );
  DFF_X2 _f_permutation__out_reg_1179_  ( .D(_f_permutation__n4208 ), .CK(clk), 
        .Q(out[99]), .QN() );
  DFF_X2 _f_permutation__out_reg_1178_  ( .D(_f_permutation__n4209 ), .CK(clk), 
        .Q(out[98]), .QN() );
  DFF_X2 _f_permutation__out_reg_1177_  ( .D(_f_permutation__n4210 ), .CK(clk), 
        .Q(out[97]), .QN() );
  DFF_X2 _f_permutation__out_reg_1176_  ( .D(_f_permutation__n4211 ), .CK(clk), 
        .Q(out[96]), .QN() );
  DFF_X2 _f_permutation__out_reg_1175_  ( .D(_f_permutation__n4212 ), .CK(clk), 
        .Q(out[111]), .QN() );
  DFF_X2 _f_permutation__out_reg_1174_  ( .D(_f_permutation__n4213 ), .CK(clk), 
        .Q(out[110]), .QN() );
  DFF_X2 _f_permutation__out_reg_1173_  ( .D(_f_permutation__n4214 ), .CK(clk), 
        .Q(out[109]), .QN() );
  DFF_X2 _f_permutation__out_reg_1172_  ( .D(_f_permutation__n4215 ), .CK(clk), 
        .Q(out[108]), .QN() );
  DFF_X2 _f_permutation__out_reg_1171_  ( .D(_f_permutation__n4216 ), .CK(clk), 
        .Q(out[107]), .QN() );
  DFF_X2 _f_permutation__out_reg_1170_  ( .D(_f_permutation__n4217 ), .CK(clk), 
        .Q(out[106]), .QN() );
  DFF_X2 _f_permutation__out_reg_1169_  ( .D(_f_permutation__n4218 ), .CK(clk), 
        .Q(out[105]), .QN() );
  DFF_X2 _f_permutation__out_reg_1168_  ( .D(_f_permutation__n4219 ), .CK(clk), 
        .Q(out[104]), .QN() );
  DFF_X2 _f_permutation__out_reg_1167_  ( .D(_f_permutation__n4220 ), .CK(clk), 
        .Q(out[119]), .QN() );
  DFF_X2 _f_permutation__out_reg_1166_  ( .D(_f_permutation__n4221 ), .CK(clk), 
        .Q(out[118]), .QN() );
  DFF_X2 _f_permutation__out_reg_1165_  ( .D(_f_permutation__n4222 ), .CK(clk), 
        .Q(out[117]), .QN() );
  DFF_X2 _f_permutation__out_reg_1164_  ( .D(_f_permutation__n4223 ), .CK(clk), 
        .Q(out[116]), .QN() );
  DFF_X2 _f_permutation__out_reg_1163_  ( .D(_f_permutation__n4224 ), .CK(clk), 
        .Q(out[115]), .QN() );
  DFF_X2 _f_permutation__out_reg_1162_  ( .D(_f_permutation__n4225 ), .CK(clk), 
        .Q(out[114]), .QN() );
  DFF_X2 _f_permutation__out_reg_1161_  ( .D(_f_permutation__n4226 ), .CK(clk), 
        .Q(out[113]), .QN() );
  DFF_X2 _f_permutation__out_reg_1160_  ( .D(_f_permutation__n4227 ), .CK(clk), 
        .Q(out[112]), .QN() );
  DFF_X2 _f_permutation__out_reg_1159_  ( .D(_f_permutation__n4228 ), .CK(clk), 
        .Q(out[127]), .QN() );
  DFF_X2 _f_permutation__out_reg_1158_  ( .D(_f_permutation__n4229 ), .CK(clk), 
        .Q(out[126]), .QN() );
  DFF_X2 _f_permutation__out_reg_1157_  ( .D(_f_permutation__n4230 ), .CK(clk), 
        .Q(out[125]), .QN() );
  DFF_X2 _f_permutation__out_reg_1156_  ( .D(_f_permutation__n4231 ), .CK(clk), 
        .Q(out[124]), .QN() );
  DFF_X2 _f_permutation__out_reg_1155_  ( .D(_f_permutation__n4232 ), .CK(clk), 
        .Q(out[123]), .QN() );
  DFF_X2 _f_permutation__out_reg_1154_  ( .D(_f_permutation__n4233 ), .CK(clk), 
        .Q(out[122]), .QN() );
  DFF_X2 _f_permutation__out_reg_1153_  ( .D(_f_permutation__n4234 ), .CK(clk), 
        .Q(out[121]), .QN() );
  DFF_X2 _f_permutation__out_reg_1152_  ( .D(_f_permutation__n4235 ), .CK(clk), 
        .Q(out[120]), .QN() );
  DFF_X2 _f_permutation__out_reg_1151_  ( .D(_f_permutation__n4236 ), .CK(clk), 
        .Q(out[7]), .QN() );
  DFF_X2 _f_permutation__out_reg_1150_  ( .D(_f_permutation__n4237 ), .CK(clk), 
        .Q(out[6]), .QN() );
  DFF_X2 _f_permutation__out_reg_1149_  ( .D(_f_permutation__n4238 ), .CK(clk), 
        .Q(out[5]), .QN() );
  DFF_X2 _f_permutation__out_reg_1148_  ( .D(_f_permutation__n4239 ), .CK(clk), 
        .Q(out[4]), .QN() );
  DFF_X2 _f_permutation__out_reg_1147_  ( .D(_f_permutation__n4240 ), .CK(clk), 
        .Q(out[3]), .QN() );
  DFF_X2 _f_permutation__out_reg_1146_  ( .D(_f_permutation__n4241 ), .CK(clk), 
        .Q(out[2]), .QN() );
  DFF_X2 _f_permutation__out_reg_1145_  ( .D(_f_permutation__n4242 ), .CK(clk), 
        .Q(out[1]), .QN() );
  DFF_X2 _f_permutation__out_reg_1144_  ( .D(_f_permutation__n4243 ), .CK(clk), 
        .Q(out[0]), .QN() );
  DFF_X2 _f_permutation__out_reg_1143_  ( .D(_f_permutation__n4244 ), .CK(clk), 
        .Q(out[15]), .QN() );
  DFF_X2 _f_permutation__out_reg_1142_  ( .D(_f_permutation__n4245 ), .CK(clk), 
        .Q(out[14]), .QN() );
  DFF_X2 _f_permutation__out_reg_1141_  ( .D(_f_permutation__n4246 ), .CK(clk), 
        .Q(out[13]), .QN() );
  DFF_X2 _f_permutation__out_reg_1140_  ( .D(_f_permutation__n4247 ), .CK(clk), 
        .Q(out[12]), .QN() );
  DFF_X2 _f_permutation__out_reg_1139_  ( .D(_f_permutation__n4248 ), .CK(clk), 
        .Q(out[11]), .QN() );
  DFF_X2 _f_permutation__out_reg_1138_  ( .D(_f_permutation__n4249 ), .CK(clk), 
        .Q(out[10]), .QN() );
  DFF_X2 _f_permutation__out_reg_1137_  ( .D(_f_permutation__n4250 ), .CK(clk), 
        .Q(out[9]), .QN() );
  DFF_X2 _f_permutation__out_reg_1136_  ( .D(_f_permutation__n4251 ), .CK(clk), 
        .Q(out[8]), .QN() );
  DFF_X2 _f_permutation__out_reg_1135_  ( .D(_f_permutation__n4252 ), .CK(clk), 
        .Q(out[23]), .QN() );
  DFF_X2 _f_permutation__out_reg_1134_  ( .D(_f_permutation__n4253 ), .CK(clk), 
        .Q(out[22]), .QN() );
  DFF_X2 _f_permutation__out_reg_1133_  ( .D(_f_permutation__n4254 ), .CK(clk), 
        .Q(out[21]), .QN() );
  DFF_X2 _f_permutation__out_reg_1132_  ( .D(_f_permutation__n4255 ), .CK(clk), 
        .Q(out[20]), .QN() );
  DFF_X2 _f_permutation__out_reg_1131_  ( .D(_f_permutation__n4256 ), .CK(clk), 
        .Q(out[19]), .QN() );
  DFF_X2 _f_permutation__out_reg_1130_  ( .D(_f_permutation__n4257 ), .CK(clk), 
        .Q(out[18]), .QN() );
  DFF_X2 _f_permutation__out_reg_1129_  ( .D(_f_permutation__n4258 ), .CK(clk), 
        .Q(out[17]), .QN() );
  DFF_X2 _f_permutation__out_reg_1128_  ( .D(_f_permutation__n4259 ), .CK(clk), 
        .Q(out[16]), .QN() );
  DFF_X2 _f_permutation__out_reg_1127_  ( .D(_f_permutation__n4260 ), .CK(clk), 
        .Q(out[31]), .QN() );
  DFF_X2 _f_permutation__out_reg_1126_  ( .D(_f_permutation__n4261 ), .CK(clk), 
        .Q(out[30]), .QN() );
  DFF_X2 _f_permutation__out_reg_1125_  ( .D(_f_permutation__n4262 ), .CK(clk), 
        .Q(out[29]), .QN() );
  DFF_X2 _f_permutation__out_reg_1124_  ( .D(_f_permutation__n4263 ), .CK(clk), 
        .Q(out[28]), .QN() );
  DFF_X2 _f_permutation__out_reg_1123_  ( .D(_f_permutation__n4264 ), .CK(clk), 
        .Q(out[27]), .QN() );
  DFF_X2 _f_permutation__out_reg_1122_  ( .D(_f_permutation__n4265 ), .CK(clk), 
        .Q(out[26]), .QN() );
  DFF_X2 _f_permutation__out_reg_1121_  ( .D(_f_permutation__n4266 ), .CK(clk), 
        .Q(out[25]), .QN() );
  DFF_X2 _f_permutation__out_reg_1120_  ( .D(_f_permutation__n4267 ), .CK(clk), 
        .Q(out[24]), .QN() );
  DFF_X2 _f_permutation__out_reg_1119_  ( .D(_f_permutation__n4268 ), .CK(clk), 
        .Q(out[39]), .QN() );
  DFF_X2 _f_permutation__out_reg_1118_  ( .D(_f_permutation__n4269 ), .CK(clk), 
        .Q(out[38]), .QN() );
  DFF_X2 _f_permutation__out_reg_1117_  ( .D(_f_permutation__n4270 ), .CK(clk), 
        .Q(out[37]), .QN() );
  DFF_X2 _f_permutation__out_reg_1116_  ( .D(_f_permutation__n4271 ), .CK(clk), 
        .Q(out[36]), .QN() );
  DFF_X2 _f_permutation__out_reg_1115_  ( .D(_f_permutation__n4272 ), .CK(clk), 
        .Q(out[35]), .QN() );
  DFF_X2 _f_permutation__out_reg_1114_  ( .D(_f_permutation__n4273 ), .CK(clk), 
        .Q(out[34]), .QN() );
  DFF_X2 _f_permutation__out_reg_1113_  ( .D(_f_permutation__n4274 ), .CK(clk), 
        .Q(out[33]), .QN() );
  DFF_X2 _f_permutation__out_reg_1112_  ( .D(_f_permutation__n4275 ), .CK(clk), 
        .Q(out[32]), .QN() );
  DFF_X2 _f_permutation__out_reg_1111_  ( .D(_f_permutation__n4276 ), .CK(clk), 
        .Q(out[47]), .QN() );
  DFF_X2 _f_permutation__out_reg_1110_  ( .D(_f_permutation__n4277 ), .CK(clk), 
        .Q(out[46]), .QN() );
  DFF_X2 _f_permutation__out_reg_1109_  ( .D(_f_permutation__n4278 ), .CK(clk), 
        .Q(out[45]), .QN() );
  DFF_X2 _f_permutation__out_reg_1108_  ( .D(_f_permutation__n4279 ), .CK(clk), 
        .Q(out[44]), .QN() );
  DFF_X2 _f_permutation__out_reg_1107_  ( .D(_f_permutation__n4280 ), .CK(clk), 
        .Q(out[43]), .QN() );
  DFF_X2 _f_permutation__out_reg_1106_  ( .D(_f_permutation__n4281 ), .CK(clk), 
        .Q(out[42]), .QN() );
  DFF_X2 _f_permutation__out_reg_1105_  ( .D(_f_permutation__n4282 ), .CK(clk), 
        .Q(out[41]), .QN() );
  DFF_X2 _f_permutation__out_reg_1104_  ( .D(_f_permutation__n4283 ), .CK(clk), 
        .Q(out[40]), .QN() );
  DFF_X2 _f_permutation__out_reg_1103_  ( .D(_f_permutation__n4284 ), .CK(clk), 
        .Q(out[55]), .QN() );
  DFF_X2 _f_permutation__out_reg_1102_  ( .D(_f_permutation__n4285 ), .CK(clk), 
        .Q(out[54]), .QN() );
  DFF_X2 _f_permutation__out_reg_1101_  ( .D(_f_permutation__n4286 ), .CK(clk), 
        .Q(out[53]), .QN() );
  DFF_X2 _f_permutation__out_reg_1100_  ( .D(_f_permutation__n4287 ), .CK(clk), 
        .Q(out[52]), .QN() );
  DFF_X2 _f_permutation__out_reg_1099_  ( .D(_f_permutation__n4288 ), .CK(clk), 
        .Q(out[51]), .QN() );
  DFF_X2 _f_permutation__out_reg_1098_  ( .D(_f_permutation__n4289 ), .CK(clk), 
        .Q(out[50]), .QN() );
  DFF_X2 _f_permutation__out_reg_1097_  ( .D(_f_permutation__n4290 ), .CK(clk), 
        .Q(out[49]), .QN() );
  DFF_X2 _f_permutation__out_reg_1096_  ( .D(_f_permutation__n4291 ), .CK(clk), 
        .Q(out[48]), .QN() );
  DFF_X2 _f_permutation__out_reg_1095_  ( .D(_f_permutation__n4292 ), .CK(clk), 
        .Q(out[63]), .QN() );
  DFF_X2 _f_permutation__out_reg_1094_  ( .D(_f_permutation__n4293 ), .CK(clk), 
        .Q(out[62]), .QN() );
  DFF_X2 _f_permutation__out_reg_1093_  ( .D(_f_permutation__n4294 ), .CK(clk), 
        .Q(out[61]), .QN() );
  DFF_X2 _f_permutation__out_reg_1092_  ( .D(_f_permutation__n4295 ), .CK(clk), 
        .Q(out[60]), .QN() );
  DFF_X2 _f_permutation__out_reg_1091_  ( .D(_f_permutation__n4296 ), .CK(clk), 
        .Q(out[59]), .QN() );
  DFF_X2 _f_permutation__out_reg_1090_  ( .D(_f_permutation__n4297 ), .CK(clk), 
        .Q(out[58]), .QN() );
  DFF_X2 _f_permutation__out_reg_1089_  ( .D(_f_permutation__n4298 ), .CK(clk), 
        .Q(out[57]), .QN() );
  DFF_X2 _f_permutation__out_reg_1088_  ( .D(_f_permutation__n4299 ), .CK(clk), 
        .Q(out[56]), .QN() );
  DFF_X2 _f_permutation__out_reg_1087_  ( .D(_f_permutation__n4300 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1), .QN() );
  DFF_X2 _f_permutation__out_reg_1086_  ( .D(_f_permutation__n4301 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_2), .QN() );
  DFF_X2 _f_permutation__out_reg_1085_  ( .D(_f_permutation__n4302 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_3), .QN() );
  DFF_X2 _f_permutation__out_reg_1084_  ( .D(_f_permutation__n4303 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_4), .QN() );
  DFF_X2 _f_permutation__out_reg_1083_  ( .D(_f_permutation__n4304 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_5), .QN() );
  DFF_X2 _f_permutation__out_reg_1082_  ( .D(_f_permutation__n4305 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_6), .QN() );
  DFF_X2 _f_permutation__out_reg_1081_  ( .D(_f_permutation__n4306 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_7), .QN() );
  DFF_X2 _f_permutation__out_reg_1080_  ( .D(_f_permutation__n4307 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_8), .QN() );
  DFF_X2 _f_permutation__out_reg_1079_  ( .D(_f_permutation__n4308 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_9), .QN() );
  DFF_X2 _f_permutation__out_reg_1078_  ( .D(_f_permutation__n4309 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_10), .QN() );
  DFF_X2 _f_permutation__out_reg_1077_  ( .D(_f_permutation__n4310 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_11), .QN() );
  DFF_X2 _f_permutation__out_reg_1076_  ( .D(_f_permutation__n4311 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_12), .QN() );
  DFF_X2 _f_permutation__out_reg_1075_  ( .D(_f_permutation__n4312 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_13), .QN() );
  DFF_X2 _f_permutation__out_reg_1074_  ( .D(_f_permutation__n4313 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_14), .QN() );
  DFF_X2 _f_permutation__out_reg_1073_  ( .D(_f_permutation__n4314 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_15), .QN() );
  DFF_X2 _f_permutation__out_reg_1072_  ( .D(_f_permutation__n4315 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_16), .QN() );
  DFF_X2 _f_permutation__out_reg_1071_  ( .D(_f_permutation__n4316 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_17), .QN() );
  DFF_X2 _f_permutation__out_reg_1070_  ( .D(_f_permutation__n4317 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_18), .QN() );
  DFF_X2 _f_permutation__out_reg_1069_  ( .D(_f_permutation__n4318 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_19), .QN() );
  DFF_X2 _f_permutation__out_reg_1068_  ( .D(_f_permutation__n4319 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_20), .QN() );
  DFF_X2 _f_permutation__out_reg_1067_  ( .D(_f_permutation__n4320 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_21), .QN() );
  DFF_X2 _f_permutation__out_reg_1066_  ( .D(_f_permutation__n4321 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_22), .QN() );
  DFF_X2 _f_permutation__out_reg_1065_  ( .D(_f_permutation__n4322 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_23), .QN() );
  DFF_X2 _f_permutation__out_reg_1064_  ( .D(_f_permutation__n4323 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_24), .QN() );
  DFF_X2 _f_permutation__out_reg_1063_  ( .D(_f_permutation__n4324 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_25), .QN() );
  DFF_X2 _f_permutation__out_reg_1062_  ( .D(_f_permutation__n4325 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_26), .QN() );
  DFF_X2 _f_permutation__out_reg_1061_  ( .D(_f_permutation__n4326 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_27), .QN() );
  DFF_X2 _f_permutation__out_reg_1060_  ( .D(_f_permutation__n4327 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_28), .QN() );
  DFF_X2 _f_permutation__out_reg_1059_  ( .D(_f_permutation__n4328 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_29), .QN() );
  DFF_X2 _f_permutation__out_reg_1058_  ( .D(_f_permutation__n4329 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_30), .QN() );
  DFF_X2 _f_permutation__out_reg_1057_  ( .D(_f_permutation__n4330 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_31), .QN() );
  DFF_X2 _f_permutation__out_reg_1056_  ( .D(_f_permutation__n4331 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_32), .QN() );
  DFF_X2 _f_permutation__out_reg_1055_  ( .D(_f_permutation__n4332 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_33), .QN() );
  DFF_X2 _f_permutation__out_reg_1054_  ( .D(_f_permutation__n4333 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_34), .QN() );
  DFF_X2 _f_permutation__out_reg_1053_  ( .D(_f_permutation__n4334 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_35), .QN() );
  DFF_X2 _f_permutation__out_reg_1052_  ( .D(_f_permutation__n4335 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_36), .QN() );
  DFF_X2 _f_permutation__out_reg_1051_  ( .D(_f_permutation__n4336 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_37), .QN() );
  DFF_X2 _f_permutation__out_reg_1050_  ( .D(_f_permutation__n4337 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_38), .QN() );
  DFF_X2 _f_permutation__out_reg_1049_  ( .D(_f_permutation__n4338 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_39), .QN() );
  DFF_X2 _f_permutation__out_reg_1048_  ( .D(_f_permutation__n4339 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_40), .QN() );
  DFF_X2 _f_permutation__out_reg_1047_  ( .D(_f_permutation__n4340 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_41), .QN() );
  DFF_X2 _f_permutation__out_reg_1046_  ( .D(_f_permutation__n4341 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_42), .QN() );
  DFF_X2 _f_permutation__out_reg_1045_  ( .D(_f_permutation__n4342 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_43), .QN() );
  DFF_X2 _f_permutation__out_reg_1044_  ( .D(_f_permutation__n4343 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_44), .QN() );
  DFF_X2 _f_permutation__out_reg_1043_  ( .D(_f_permutation__n4344 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_45), .QN() );
  DFF_X2 _f_permutation__out_reg_1042_  ( .D(_f_permutation__n4345 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_46), .QN() );
  DFF_X2 _f_permutation__out_reg_1041_  ( .D(_f_permutation__n4346 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_47), .QN() );
  DFF_X2 _f_permutation__out_reg_1040_  ( .D(_f_permutation__n4347 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_48), .QN() );
  DFF_X2 _f_permutation__out_reg_1039_  ( .D(_f_permutation__n4348 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_49), .QN() );
  DFF_X2 _f_permutation__out_reg_1038_  ( .D(_f_permutation__n4349 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_50), .QN() );
  DFF_X2 _f_permutation__out_reg_1037_  ( .D(_f_permutation__n4350 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_51), .QN() );
  DFF_X2 _f_permutation__out_reg_1036_  ( .D(_f_permutation__n4351 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_52), .QN() );
  DFF_X2 _f_permutation__out_reg_1035_  ( .D(_f_permutation__n4352 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_53), .QN() );
  DFF_X2 _f_permutation__out_reg_1034_  ( .D(_f_permutation__n4353 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_54), .QN() );
  DFF_X2 _f_permutation__out_reg_1033_  ( .D(_f_permutation__n4354 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_55), .QN() );
  DFF_X2 _f_permutation__out_reg_1032_  ( .D(_f_permutation__n4355 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_56), .QN() );
  DFF_X2 _f_permutation__out_reg_1031_  ( .D(_f_permutation__n4356 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_57), .QN() );
  DFF_X2 _f_permutation__out_reg_1030_  ( .D(_f_permutation__n4357 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_58), .QN() );
  DFF_X2 _f_permutation__out_reg_1029_  ( .D(_f_permutation__n4358 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_59), .QN() );
  DFF_X2 _f_permutation__out_reg_1028_  ( .D(_f_permutation__n4359 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_60), .QN() );
  DFF_X2 _f_permutation__out_reg_1027_  ( .D(_f_permutation__n4360 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_61), .QN() );
  DFF_X2 _f_permutation__out_reg_1026_  ( .D(_f_permutation__n4361 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_62), .QN() );
  DFF_X2 _f_permutation__out_reg_1025_  ( .D(_f_permutation__n4362 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_63), .QN() );
  DFF_X2 _f_permutation__out_reg_1024_  ( .D(_f_permutation__n4363 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_64), .QN() );
  DFF_X2 _f_permutation__out_reg_1023_  ( .D(_f_permutation__n4364 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_65), .QN() );
  DFF_X2 _f_permutation__out_reg_1022_  ( .D(_f_permutation__n4365 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_66), .QN() );
  DFF_X2 _f_permutation__out_reg_1021_  ( .D(_f_permutation__n4366 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_67), .QN() );
  DFF_X2 _f_permutation__out_reg_1020_  ( .D(_f_permutation__n4367 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_68), .QN() );
  DFF_X2 _f_permutation__out_reg_1019_  ( .D(_f_permutation__n4368 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_69), .QN() );
  DFF_X2 _f_permutation__out_reg_1018_  ( .D(_f_permutation__n4369 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_70), .QN() );
  DFF_X2 _f_permutation__out_reg_1017_  ( .D(_f_permutation__n4370 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_71), .QN() );
  DFF_X2 _f_permutation__out_reg_1016_  ( .D(_f_permutation__n4371 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_72), .QN() );
  DFF_X2 _f_permutation__out_reg_1015_  ( .D(_f_permutation__n4372 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_73), .QN() );
  DFF_X2 _f_permutation__out_reg_1014_  ( .D(_f_permutation__n4373 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_74), .QN() );
  DFF_X2 _f_permutation__out_reg_1013_  ( .D(_f_permutation__n4374 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_75), .QN() );
  DFF_X2 _f_permutation__out_reg_1012_  ( .D(_f_permutation__n4375 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_76), .QN() );
  DFF_X2 _f_permutation__out_reg_1011_  ( .D(_f_permutation__n4376 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_77), .QN() );
  DFF_X2 _f_permutation__out_reg_1010_  ( .D(_f_permutation__n4377 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_78), .QN() );
  DFF_X2 _f_permutation__out_reg_1009_  ( .D(_f_permutation__n4378 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_79), .QN() );
  DFF_X2 _f_permutation__out_reg_1008_  ( .D(_f_permutation__n4379 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_80), .QN() );
  DFF_X2 _f_permutation__out_reg_1007_  ( .D(_f_permutation__n4380 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_81), .QN() );
  DFF_X2 _f_permutation__out_reg_1006_  ( .D(_f_permutation__n4381 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_82), .QN() );
  DFF_X2 _f_permutation__out_reg_1005_  ( .D(_f_permutation__n4382 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_83), .QN() );
  DFF_X2 _f_permutation__out_reg_1004_  ( .D(_f_permutation__n4383 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_84), .QN() );
  DFF_X2 _f_permutation__out_reg_1003_  ( .D(_f_permutation__n4384 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_85), .QN() );
  DFF_X2 _f_permutation__out_reg_1002_  ( .D(_f_permutation__n4385 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_86), .QN() );
  DFF_X2 _f_permutation__out_reg_1001_  ( .D(_f_permutation__n4386 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_87), .QN() );
  DFF_X2 _f_permutation__out_reg_1000_  ( .D(_f_permutation__n4387 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_88), .QN() );
  DFF_X2 _f_permutation__out_reg_999_  ( .D(_f_permutation__n4388 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_89), .QN() );
  DFF_X2 _f_permutation__out_reg_998_  ( .D(_f_permutation__n4389 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_90), .QN() );
  DFF_X2 _f_permutation__out_reg_997_  ( .D(_f_permutation__n4390 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_91), .QN() );
  DFF_X2 _f_permutation__out_reg_996_  ( .D(_f_permutation__n4391 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_92), .QN() );
  DFF_X2 _f_permutation__out_reg_995_  ( .D(_f_permutation__n4392 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_93), .QN() );
  DFF_X2 _f_permutation__out_reg_994_  ( .D(_f_permutation__n4393 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_94), .QN() );
  DFF_X2 _f_permutation__out_reg_993_  ( .D(_f_permutation__n4394 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_95), .QN() );
  DFF_X2 _f_permutation__out_reg_992_  ( .D(_f_permutation__n4395 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_96), .QN() );
  DFF_X2 _f_permutation__out_reg_991_  ( .D(_f_permutation__n4396 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_97), .QN() );
  DFF_X2 _f_permutation__out_reg_990_  ( .D(_f_permutation__n4397 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_98), .QN() );
  DFF_X2 _f_permutation__out_reg_989_  ( .D(_f_permutation__n4398 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_99), .QN() );
  DFF_X2 _f_permutation__out_reg_988_  ( .D(_f_permutation__n4399 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_100), .QN() );
  DFF_X2 _f_permutation__out_reg_987_  ( .D(_f_permutation__n4400 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_101), .QN() );
  DFF_X2 _f_permutation__out_reg_986_  ( .D(_f_permutation__n4401 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_102), .QN() );
  DFF_X2 _f_permutation__out_reg_985_  ( .D(_f_permutation__n4402 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_103), .QN() );
  DFF_X2 _f_permutation__out_reg_984_  ( .D(_f_permutation__n4403 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_104), .QN() );
  DFF_X2 _f_permutation__out_reg_983_  ( .D(_f_permutation__n4404 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_105), .QN() );
  DFF_X2 _f_permutation__out_reg_982_  ( .D(_f_permutation__n4405 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_106), .QN() );
  DFF_X2 _f_permutation__out_reg_981_  ( .D(_f_permutation__n4406 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_107), .QN() );
  DFF_X2 _f_permutation__out_reg_980_  ( .D(_f_permutation__n4407 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_108), .QN() );
  DFF_X2 _f_permutation__out_reg_979_  ( .D(_f_permutation__n4408 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_109), .QN() );
  DFF_X2 _f_permutation__out_reg_978_  ( .D(_f_permutation__n4409 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_110), .QN() );
  DFF_X2 _f_permutation__out_reg_977_  ( .D(_f_permutation__n4410 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_111), .QN() );
  DFF_X2 _f_permutation__out_reg_976_  ( .D(_f_permutation__n4411 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_112), .QN() );
  DFF_X2 _f_permutation__out_reg_975_  ( .D(_f_permutation__n4412 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_113), .QN() );
  DFF_X2 _f_permutation__out_reg_974_  ( .D(_f_permutation__n4413 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_114), .QN() );
  DFF_X2 _f_permutation__out_reg_973_  ( .D(_f_permutation__n4414 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_115), .QN() );
  DFF_X2 _f_permutation__out_reg_972_  ( .D(_f_permutation__n4415 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_116), .QN() );
  DFF_X2 _f_permutation__out_reg_971_  ( .D(_f_permutation__n4416 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_117), .QN() );
  DFF_X2 _f_permutation__out_reg_970_  ( .D(_f_permutation__n4417 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_118), .QN() );
  DFF_X2 _f_permutation__out_reg_969_  ( .D(_f_permutation__n4418 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_119), .QN() );
  DFF_X2 _f_permutation__out_reg_968_  ( .D(_f_permutation__n4419 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_120), .QN() );
  DFF_X2 _f_permutation__out_reg_967_  ( .D(_f_permutation__n4420 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_121), .QN() );
  DFF_X2 _f_permutation__out_reg_966_  ( .D(_f_permutation__n4421 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_122), .QN() );
  DFF_X2 _f_permutation__out_reg_965_  ( .D(_f_permutation__n4422 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_123), .QN() );
  DFF_X2 _f_permutation__out_reg_964_  ( .D(_f_permutation__n4423 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_124), .QN() );
  DFF_X2 _f_permutation__out_reg_963_  ( .D(_f_permutation__n4424 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_125), .QN() );
  DFF_X2 _f_permutation__out_reg_962_  ( .D(_f_permutation__n4425 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_126), .QN() );
  DFF_X2 _f_permutation__out_reg_961_  ( .D(_f_permutation__n4426 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_127), .QN() );
  DFF_X2 _f_permutation__out_reg_960_  ( .D(_f_permutation__n4427 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_128), .QN() );
  DFF_X2 _f_permutation__out_reg_959_  ( .D(_f_permutation__n4428 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_129), .QN() );
  DFF_X2 _f_permutation__out_reg_958_  ( .D(_f_permutation__n4429 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_130), .QN() );
  DFF_X2 _f_permutation__out_reg_957_  ( .D(_f_permutation__n4430 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_131), .QN() );
  DFF_X2 _f_permutation__out_reg_956_  ( .D(_f_permutation__n4431 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_132), .QN() );
  DFF_X2 _f_permutation__out_reg_955_  ( .D(_f_permutation__n4432 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_133), .QN() );
  DFF_X2 _f_permutation__out_reg_954_  ( .D(_f_permutation__n4433 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_134), .QN() );
  DFF_X2 _f_permutation__out_reg_953_  ( .D(_f_permutation__n4434 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_135), .QN() );
  DFF_X2 _f_permutation__out_reg_952_  ( .D(_f_permutation__n4435 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_136), .QN() );
  DFF_X2 _f_permutation__out_reg_951_  ( .D(_f_permutation__n4436 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_137), .QN() );
  DFF_X2 _f_permutation__out_reg_950_  ( .D(_f_permutation__n4437 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_138), .QN() );
  DFF_X2 _f_permutation__out_reg_949_  ( .D(_f_permutation__n4438 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_139), .QN() );
  DFF_X2 _f_permutation__out_reg_948_  ( .D(_f_permutation__n4439 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_140), .QN() );
  DFF_X2 _f_permutation__out_reg_947_  ( .D(_f_permutation__n4440 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_141), .QN() );
  DFF_X2 _f_permutation__out_reg_946_  ( .D(_f_permutation__n4441 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_142), .QN() );
  DFF_X2 _f_permutation__out_reg_945_  ( .D(_f_permutation__n4442 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_143), .QN() );
  DFF_X2 _f_permutation__out_reg_944_  ( .D(_f_permutation__n4443 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_144), .QN() );
  DFF_X2 _f_permutation__out_reg_943_  ( .D(_f_permutation__n4444 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_145), .QN() );
  DFF_X2 _f_permutation__out_reg_942_  ( .D(_f_permutation__n4445 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_146), .QN() );
  DFF_X2 _f_permutation__out_reg_941_  ( .D(_f_permutation__n4446 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_147), .QN() );
  DFF_X2 _f_permutation__out_reg_940_  ( .D(_f_permutation__n4447 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_148), .QN() );
  DFF_X2 _f_permutation__out_reg_939_  ( .D(_f_permutation__n4448 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_149), .QN() );
  DFF_X2 _f_permutation__out_reg_938_  ( .D(_f_permutation__n4449 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_150), .QN() );
  DFF_X2 _f_permutation__out_reg_937_  ( .D(_f_permutation__n4450 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_151), .QN() );
  DFF_X2 _f_permutation__out_reg_936_  ( .D(_f_permutation__n4451 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_152), .QN() );
  DFF_X2 _f_permutation__out_reg_935_  ( .D(_f_permutation__n4452 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_153), .QN() );
  DFF_X2 _f_permutation__out_reg_934_  ( .D(_f_permutation__n4453 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_154), .QN() );
  DFF_X2 _f_permutation__out_reg_933_  ( .D(_f_permutation__n4454 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_155), .QN() );
  DFF_X2 _f_permutation__out_reg_932_  ( .D(_f_permutation__n4455 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_156), .QN() );
  DFF_X2 _f_permutation__out_reg_931_  ( .D(_f_permutation__n4456 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_157), .QN() );
  DFF_X2 _f_permutation__out_reg_930_  ( .D(_f_permutation__n4457 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_158), .QN() );
  DFF_X2 _f_permutation__out_reg_929_  ( .D(_f_permutation__n4458 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_159), .QN() );
  DFF_X2 _f_permutation__out_reg_928_  ( .D(_f_permutation__n4459 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_160), .QN() );
  DFF_X2 _f_permutation__out_reg_927_  ( .D(_f_permutation__n4460 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_161), .QN() );
  DFF_X2 _f_permutation__out_reg_926_  ( .D(_f_permutation__n4461 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_162), .QN() );
  DFF_X2 _f_permutation__out_reg_925_  ( .D(_f_permutation__n4462 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_163), .QN() );
  DFF_X2 _f_permutation__out_reg_924_  ( .D(_f_permutation__n4463 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_164), .QN() );
  DFF_X2 _f_permutation__out_reg_923_  ( .D(_f_permutation__n4464 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_165), .QN() );
  DFF_X2 _f_permutation__out_reg_922_  ( .D(_f_permutation__n4465 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_166), .QN() );
  DFF_X2 _f_permutation__out_reg_921_  ( .D(_f_permutation__n4466 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_167), .QN() );
  DFF_X2 _f_permutation__out_reg_920_  ( .D(_f_permutation__n4467 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_168), .QN() );
  DFF_X2 _f_permutation__out_reg_919_  ( .D(_f_permutation__n4468 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_169), .QN() );
  DFF_X2 _f_permutation__out_reg_918_  ( .D(_f_permutation__n4469 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_170), .QN() );
  DFF_X2 _f_permutation__out_reg_917_  ( .D(_f_permutation__n4470 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_171), .QN() );
  DFF_X2 _f_permutation__out_reg_916_  ( .D(_f_permutation__n4471 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_172), .QN() );
  DFF_X2 _f_permutation__out_reg_915_  ( .D(_f_permutation__n4472 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_173), .QN() );
  DFF_X2 _f_permutation__out_reg_914_  ( .D(_f_permutation__n4473 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_174), .QN() );
  DFF_X2 _f_permutation__out_reg_913_  ( .D(_f_permutation__n4474 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_175), .QN() );
  DFF_X2 _f_permutation__out_reg_912_  ( .D(_f_permutation__n4475 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_176), .QN() );
  DFF_X2 _f_permutation__out_reg_911_  ( .D(_f_permutation__n4476 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_177), .QN() );
  DFF_X2 _f_permutation__out_reg_910_  ( .D(_f_permutation__n4477 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_178), .QN() );
  DFF_X2 _f_permutation__out_reg_909_  ( .D(_f_permutation__n4478 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_179), .QN() );
  DFF_X2 _f_permutation__out_reg_908_  ( .D(_f_permutation__n4479 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_180), .QN() );
  DFF_X2 _f_permutation__out_reg_907_  ( .D(_f_permutation__n4480 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_181), .QN() );
  DFF_X2 _f_permutation__out_reg_906_  ( .D(_f_permutation__n4481 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_182), .QN() );
  DFF_X2 _f_permutation__out_reg_905_  ( .D(_f_permutation__n4482 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_183), .QN() );
  DFF_X2 _f_permutation__out_reg_904_  ( .D(_f_permutation__n4483 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_184), .QN() );
  DFF_X2 _f_permutation__out_reg_903_  ( .D(_f_permutation__n4484 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_185), .QN() );
  DFF_X2 _f_permutation__out_reg_902_  ( .D(_f_permutation__n4485 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_186), .QN() );
  DFF_X2 _f_permutation__out_reg_901_  ( .D(_f_permutation__n4486 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_187), .QN() );
  DFF_X2 _f_permutation__out_reg_900_  ( .D(_f_permutation__n4487 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_188), .QN() );
  DFF_X2 _f_permutation__out_reg_899_  ( .D(_f_permutation__n4488 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_189), .QN() );
  DFF_X2 _f_permutation__out_reg_898_  ( .D(_f_permutation__n4489 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_190), .QN() );
  DFF_X2 _f_permutation__out_reg_897_  ( .D(_f_permutation__n4490 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_191), .QN() );
  DFF_X2 _f_permutation__out_reg_896_  ( .D(_f_permutation__n4491 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_192), .QN() );
  DFF_X2 _f_permutation__out_reg_895_  ( .D(_f_permutation__n4492 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_193), .QN() );
  DFF_X2 _f_permutation__out_reg_894_  ( .D(_f_permutation__n4493 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_194), .QN() );
  DFF_X2 _f_permutation__out_reg_893_  ( .D(_f_permutation__n4494 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_195), .QN() );
  DFF_X2 _f_permutation__out_reg_892_  ( .D(_f_permutation__n4495 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_196), .QN() );
  DFF_X2 _f_permutation__out_reg_891_  ( .D(_f_permutation__n4496 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_197), .QN() );
  DFF_X2 _f_permutation__out_reg_890_  ( .D(_f_permutation__n4497 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_198), .QN() );
  DFF_X2 _f_permutation__out_reg_889_  ( .D(_f_permutation__n4498 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_199), .QN() );
  DFF_X2 _f_permutation__out_reg_888_  ( .D(_f_permutation__n4499 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_200), .QN() );
  DFF_X2 _f_permutation__out_reg_887_  ( .D(_f_permutation__n4500 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_201), .QN() );
  DFF_X2 _f_permutation__out_reg_886_  ( .D(_f_permutation__n4501 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_202), .QN() );
  DFF_X2 _f_permutation__out_reg_885_  ( .D(_f_permutation__n4502 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_203), .QN() );
  DFF_X2 _f_permutation__out_reg_884_  ( .D(_f_permutation__n4503 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_204), .QN() );
  DFF_X2 _f_permutation__out_reg_883_  ( .D(_f_permutation__n4504 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_205), .QN() );
  DFF_X2 _f_permutation__out_reg_882_  ( .D(_f_permutation__n4505 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_206), .QN() );
  DFF_X2 _f_permutation__out_reg_881_  ( .D(_f_permutation__n4506 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_207), .QN() );
  DFF_X2 _f_permutation__out_reg_880_  ( .D(_f_permutation__n4507 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_208), .QN() );
  DFF_X2 _f_permutation__out_reg_879_  ( .D(_f_permutation__n4508 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_209), .QN() );
  DFF_X2 _f_permutation__out_reg_878_  ( .D(_f_permutation__n4509 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_210), .QN() );
  DFF_X2 _f_permutation__out_reg_877_  ( .D(_f_permutation__n4510 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_211), .QN() );
  DFF_X2 _f_permutation__out_reg_876_  ( .D(_f_permutation__n4511 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_212), .QN() );
  DFF_X2 _f_permutation__out_reg_875_  ( .D(_f_permutation__n4512 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_213), .QN() );
  DFF_X2 _f_permutation__out_reg_874_  ( .D(_f_permutation__n4513 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_214), .QN() );
  DFF_X2 _f_permutation__out_reg_873_  ( .D(_f_permutation__n4514 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_215), .QN() );
  DFF_X2 _f_permutation__out_reg_872_  ( .D(_f_permutation__n4515 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_216), .QN() );
  DFF_X2 _f_permutation__out_reg_871_  ( .D(_f_permutation__n4516 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_217), .QN() );
  DFF_X2 _f_permutation__out_reg_870_  ( .D(_f_permutation__n4517 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_218), .QN() );
  DFF_X2 _f_permutation__out_reg_869_  ( .D(_f_permutation__n4518 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_219), .QN() );
  DFF_X2 _f_permutation__out_reg_868_  ( .D(_f_permutation__n4519 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_220), .QN() );
  DFF_X2 _f_permutation__out_reg_867_  ( .D(_f_permutation__n4520 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_221), .QN() );
  DFF_X2 _f_permutation__out_reg_866_  ( .D(_f_permutation__n4521 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_222), .QN() );
  DFF_X2 _f_permutation__out_reg_865_  ( .D(_f_permutation__n4522 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_223), .QN() );
  DFF_X2 _f_permutation__out_reg_864_  ( .D(_f_permutation__n4523 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_224), .QN() );
  DFF_X2 _f_permutation__out_reg_863_  ( .D(_f_permutation__n4524 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_225), .QN() );
  DFF_X2 _f_permutation__out_reg_862_  ( .D(_f_permutation__n4525 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_226), .QN() );
  DFF_X2 _f_permutation__out_reg_861_  ( .D(_f_permutation__n4526 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_227), .QN() );
  DFF_X2 _f_permutation__out_reg_860_  ( .D(_f_permutation__n4527 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_228), .QN() );
  DFF_X2 _f_permutation__out_reg_859_  ( .D(_f_permutation__n4528 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_229), .QN() );
  DFF_X2 _f_permutation__out_reg_858_  ( .D(_f_permutation__n4529 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_230), .QN() );
  DFF_X2 _f_permutation__out_reg_857_  ( .D(_f_permutation__n4530 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_231), .QN() );
  DFF_X2 _f_permutation__out_reg_856_  ( .D(_f_permutation__n4531 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_232), .QN() );
  DFF_X2 _f_permutation__out_reg_855_  ( .D(_f_permutation__n4532 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_233), .QN() );
  DFF_X2 _f_permutation__out_reg_854_  ( .D(_f_permutation__n4533 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_234), .QN() );
  DFF_X2 _f_permutation__out_reg_853_  ( .D(_f_permutation__n4534 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_235), .QN() );
  DFF_X2 _f_permutation__out_reg_852_  ( .D(_f_permutation__n4535 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_236), .QN() );
  DFF_X2 _f_permutation__out_reg_851_  ( .D(_f_permutation__n4536 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_237), .QN() );
  DFF_X2 _f_permutation__out_reg_850_  ( .D(_f_permutation__n4537 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_238), .QN() );
  DFF_X2 _f_permutation__out_reg_849_  ( .D(_f_permutation__n4538 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_239), .QN() );
  DFF_X2 _f_permutation__out_reg_848_  ( .D(_f_permutation__n4539 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_240), .QN() );
  DFF_X2 _f_permutation__out_reg_847_  ( .D(_f_permutation__n4540 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_241), .QN() );
  DFF_X2 _f_permutation__out_reg_846_  ( .D(_f_permutation__n4541 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_242), .QN() );
  DFF_X2 _f_permutation__out_reg_845_  ( .D(_f_permutation__n4542 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_243), .QN() );
  DFF_X2 _f_permutation__out_reg_844_  ( .D(_f_permutation__n4543 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_244), .QN() );
  DFF_X2 _f_permutation__out_reg_843_  ( .D(_f_permutation__n4544 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_245), .QN() );
  DFF_X2 _f_permutation__out_reg_842_  ( .D(_f_permutation__n4545 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_246), .QN() );
  DFF_X2 _f_permutation__out_reg_841_  ( .D(_f_permutation__n4546 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_247), .QN() );
  DFF_X2 _f_permutation__out_reg_840_  ( .D(_f_permutation__n4547 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_248), .QN() );
  DFF_X2 _f_permutation__out_reg_839_  ( .D(_f_permutation__n4548 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_249), .QN() );
  DFF_X2 _f_permutation__out_reg_838_  ( .D(_f_permutation__n4549 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_250), .QN() );
  DFF_X2 _f_permutation__out_reg_837_  ( .D(_f_permutation__n4550 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_251), .QN() );
  DFF_X2 _f_permutation__out_reg_836_  ( .D(_f_permutation__n4551 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_252), .QN() );
  DFF_X2 _f_permutation__out_reg_835_  ( .D(_f_permutation__n4552 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_253), .QN() );
  DFF_X2 _f_permutation__out_reg_834_  ( .D(_f_permutation__n4553 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_254), .QN() );
  DFF_X2 _f_permutation__out_reg_833_  ( .D(_f_permutation__n4554 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_255), .QN() );
  DFF_X2 _f_permutation__out_reg_832_  ( .D(_f_permutation__n4555 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_256), .QN() );
  DFF_X2 _f_permutation__out_reg_831_  ( .D(_f_permutation__n4556 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_257), .QN() );
  DFF_X2 _f_permutation__out_reg_830_  ( .D(_f_permutation__n4557 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_258), .QN() );
  DFF_X2 _f_permutation__out_reg_829_  ( .D(_f_permutation__n4558 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_259), .QN() );
  DFF_X2 _f_permutation__out_reg_828_  ( .D(_f_permutation__n4559 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_260), .QN() );
  DFF_X2 _f_permutation__out_reg_827_  ( .D(_f_permutation__n4560 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_261), .QN() );
  DFF_X2 _f_permutation__out_reg_826_  ( .D(_f_permutation__n4561 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_262), .QN() );
  DFF_X2 _f_permutation__out_reg_825_  ( .D(_f_permutation__n4562 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_263), .QN() );
  DFF_X2 _f_permutation__out_reg_824_  ( .D(_f_permutation__n4563 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_264), .QN() );
  DFF_X2 _f_permutation__out_reg_823_  ( .D(_f_permutation__n4564 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_265), .QN() );
  DFF_X2 _f_permutation__out_reg_822_  ( .D(_f_permutation__n4565 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_266), .QN() );
  DFF_X2 _f_permutation__out_reg_821_  ( .D(_f_permutation__n4566 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_267), .QN() );
  DFF_X2 _f_permutation__out_reg_820_  ( .D(_f_permutation__n4567 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_268), .QN() );
  DFF_X2 _f_permutation__out_reg_819_  ( .D(_f_permutation__n4568 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_269), .QN() );
  DFF_X2 _f_permutation__out_reg_818_  ( .D(_f_permutation__n4569 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_270), .QN() );
  DFF_X2 _f_permutation__out_reg_817_  ( .D(_f_permutation__n4570 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_271), .QN() );
  DFF_X2 _f_permutation__out_reg_816_  ( .D(_f_permutation__n4571 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_272), .QN() );
  DFF_X2 _f_permutation__out_reg_815_  ( .D(_f_permutation__n4572 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_273), .QN() );
  DFF_X2 _f_permutation__out_reg_814_  ( .D(_f_permutation__n4573 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_274), .QN() );
  DFF_X2 _f_permutation__out_reg_813_  ( .D(_f_permutation__n4574 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_275), .QN() );
  DFF_X2 _f_permutation__out_reg_812_  ( .D(_f_permutation__n4575 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_276), .QN() );
  DFF_X2 _f_permutation__out_reg_811_  ( .D(_f_permutation__n4576 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_277), .QN() );
  DFF_X2 _f_permutation__out_reg_810_  ( .D(_f_permutation__n4577 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_278), .QN() );
  DFF_X2 _f_permutation__out_reg_809_  ( .D(_f_permutation__n4578 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_279), .QN() );
  DFF_X2 _f_permutation__out_reg_808_  ( .D(_f_permutation__n4579 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_280), .QN() );
  DFF_X2 _f_permutation__out_reg_807_  ( .D(_f_permutation__n4580 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_281), .QN() );
  DFF_X2 _f_permutation__out_reg_806_  ( .D(_f_permutation__n4581 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_282), .QN() );
  DFF_X2 _f_permutation__out_reg_805_  ( .D(_f_permutation__n4582 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_283), .QN() );
  DFF_X2 _f_permutation__out_reg_804_  ( .D(_f_permutation__n4583 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_284), .QN() );
  DFF_X2 _f_permutation__out_reg_803_  ( .D(_f_permutation__n4584 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_285), .QN() );
  DFF_X2 _f_permutation__out_reg_802_  ( .D(_f_permutation__n4585 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_286), .QN() );
  DFF_X2 _f_permutation__out_reg_801_  ( .D(_f_permutation__n4586 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_287), .QN() );
  DFF_X2 _f_permutation__out_reg_800_  ( .D(_f_permutation__n4587 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_288), .QN() );
  DFF_X2 _f_permutation__out_reg_799_  ( .D(_f_permutation__n4588 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_289), .QN() );
  DFF_X2 _f_permutation__out_reg_798_  ( .D(_f_permutation__n4589 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_290), .QN() );
  DFF_X2 _f_permutation__out_reg_797_  ( .D(_f_permutation__n4590 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_291), .QN() );
  DFF_X2 _f_permutation__out_reg_796_  ( .D(_f_permutation__n4591 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_292), .QN() );
  DFF_X2 _f_permutation__out_reg_795_  ( .D(_f_permutation__n4592 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_293), .QN() );
  DFF_X2 _f_permutation__out_reg_794_  ( .D(_f_permutation__n4593 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_294), .QN() );
  DFF_X2 _f_permutation__out_reg_793_  ( .D(_f_permutation__n4594 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_295), .QN() );
  DFF_X2 _f_permutation__out_reg_792_  ( .D(_f_permutation__n4595 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_296), .QN() );
  DFF_X2 _f_permutation__out_reg_791_  ( .D(_f_permutation__n4596 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_297), .QN() );
  DFF_X2 _f_permutation__out_reg_790_  ( .D(_f_permutation__n4597 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_298), .QN() );
  DFF_X2 _f_permutation__out_reg_789_  ( .D(_f_permutation__n4598 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_299), .QN() );
  DFF_X2 _f_permutation__out_reg_788_  ( .D(_f_permutation__n4599 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_300), .QN() );
  DFF_X2 _f_permutation__out_reg_787_  ( .D(_f_permutation__n4600 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_301), .QN() );
  DFF_X2 _f_permutation__out_reg_786_  ( .D(_f_permutation__n4601 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_302), .QN() );
  DFF_X2 _f_permutation__out_reg_785_  ( .D(_f_permutation__n4602 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_303), .QN() );
  DFF_X2 _f_permutation__out_reg_784_  ( .D(_f_permutation__n4603 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_304), .QN() );
  DFF_X2 _f_permutation__out_reg_783_  ( .D(_f_permutation__n4604 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_305), .QN() );
  DFF_X2 _f_permutation__out_reg_782_  ( .D(_f_permutation__n4605 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_306), .QN() );
  DFF_X2 _f_permutation__out_reg_781_  ( .D(_f_permutation__n4606 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_307), .QN() );
  DFF_X2 _f_permutation__out_reg_780_  ( .D(_f_permutation__n4607 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_308), .QN() );
  DFF_X2 _f_permutation__out_reg_779_  ( .D(_f_permutation__n4608 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_309), .QN() );
  DFF_X2 _f_permutation__out_reg_778_  ( .D(_f_permutation__n4609 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_310), .QN() );
  DFF_X2 _f_permutation__out_reg_777_  ( .D(_f_permutation__n4610 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_311), .QN() );
  DFF_X2 _f_permutation__out_reg_776_  ( .D(_f_permutation__n4611 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_312), .QN() );
  DFF_X2 _f_permutation__out_reg_775_  ( .D(_f_permutation__n4612 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_313), .QN() );
  DFF_X2 _f_permutation__out_reg_774_  ( .D(_f_permutation__n4613 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_314), .QN() );
  DFF_X2 _f_permutation__out_reg_773_  ( .D(_f_permutation__n4614 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_315), .QN() );
  DFF_X2 _f_permutation__out_reg_772_  ( .D(_f_permutation__n4615 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_316), .QN() );
  DFF_X2 _f_permutation__out_reg_771_  ( .D(_f_permutation__n4616 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_317), .QN() );
  DFF_X2 _f_permutation__out_reg_770_  ( .D(_f_permutation__n4617 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_318), .QN() );
  DFF_X2 _f_permutation__out_reg_769_  ( .D(_f_permutation__n4618 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_319), .QN() );
  DFF_X2 _f_permutation__out_reg_768_  ( .D(_f_permutation__n4619 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_320), .QN() );
  DFF_X2 _f_permutation__out_reg_767_  ( .D(_f_permutation__n4620 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_321), .QN() );
  DFF_X2 _f_permutation__out_reg_766_  ( .D(_f_permutation__n4621 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_322), .QN() );
  DFF_X2 _f_permutation__out_reg_765_  ( .D(_f_permutation__n4622 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_323), .QN() );
  DFF_X2 _f_permutation__out_reg_764_  ( .D(_f_permutation__n4623 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_324), .QN() );
  DFF_X2 _f_permutation__out_reg_763_  ( .D(_f_permutation__n4624 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_325), .QN() );
  DFF_X2 _f_permutation__out_reg_762_  ( .D(_f_permutation__n4625 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_326), .QN() );
  DFF_X2 _f_permutation__out_reg_761_  ( .D(_f_permutation__n4626 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_327), .QN() );
  DFF_X2 _f_permutation__out_reg_760_  ( .D(_f_permutation__n4627 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_328), .QN() );
  DFF_X2 _f_permutation__out_reg_759_  ( .D(_f_permutation__n4628 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_329), .QN() );
  DFF_X2 _f_permutation__out_reg_758_  ( .D(_f_permutation__n4629 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_330), .QN() );
  DFF_X2 _f_permutation__out_reg_757_  ( .D(_f_permutation__n4630 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_331), .QN() );
  DFF_X2 _f_permutation__out_reg_756_  ( .D(_f_permutation__n4631 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_332), .QN() );
  DFF_X2 _f_permutation__out_reg_755_  ( .D(_f_permutation__n4632 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_333), .QN() );
  DFF_X2 _f_permutation__out_reg_754_  ( .D(_f_permutation__n4633 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_334), .QN() );
  DFF_X2 _f_permutation__out_reg_753_  ( .D(_f_permutation__n4634 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_335), .QN() );
  DFF_X2 _f_permutation__out_reg_752_  ( .D(_f_permutation__n4635 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_336), .QN() );
  DFF_X2 _f_permutation__out_reg_751_  ( .D(_f_permutation__n4636 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_337), .QN() );
  DFF_X2 _f_permutation__out_reg_750_  ( .D(_f_permutation__n4637 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_338), .QN() );
  DFF_X2 _f_permutation__out_reg_749_  ( .D(_f_permutation__n4638 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_339), .QN() );
  DFF_X2 _f_permutation__out_reg_748_  ( .D(_f_permutation__n4639 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_340), .QN() );
  DFF_X2 _f_permutation__out_reg_747_  ( .D(_f_permutation__n4640 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_341), .QN() );
  DFF_X2 _f_permutation__out_reg_746_  ( .D(_f_permutation__n4641 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_342), .QN() );
  DFF_X2 _f_permutation__out_reg_745_  ( .D(_f_permutation__n4642 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_343), .QN() );
  DFF_X2 _f_permutation__out_reg_744_  ( .D(_f_permutation__n4643 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_344), .QN() );
  DFF_X2 _f_permutation__out_reg_743_  ( .D(_f_permutation__n4644 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_345), .QN() );
  DFF_X2 _f_permutation__out_reg_742_  ( .D(_f_permutation__n4645 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_346), .QN() );
  DFF_X2 _f_permutation__out_reg_741_  ( .D(_f_permutation__n4646 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_347), .QN() );
  DFF_X2 _f_permutation__out_reg_740_  ( .D(_f_permutation__n4647 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_348), .QN() );
  DFF_X2 _f_permutation__out_reg_739_  ( .D(_f_permutation__n4648 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_349), .QN() );
  DFF_X2 _f_permutation__out_reg_738_  ( .D(_f_permutation__n4649 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_350), .QN() );
  DFF_X2 _f_permutation__out_reg_737_  ( .D(_f_permutation__n4650 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_351), .QN() );
  DFF_X2 _f_permutation__out_reg_736_  ( .D(_f_permutation__n4651 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_352), .QN() );
  DFF_X2 _f_permutation__out_reg_735_  ( .D(_f_permutation__n4652 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_353), .QN() );
  DFF_X2 _f_permutation__out_reg_734_  ( .D(_f_permutation__n4653 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_354), .QN() );
  DFF_X2 _f_permutation__out_reg_733_  ( .D(_f_permutation__n4654 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_355), .QN() );
  DFF_X2 _f_permutation__out_reg_732_  ( .D(_f_permutation__n4655 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_356), .QN() );
  DFF_X2 _f_permutation__out_reg_731_  ( .D(_f_permutation__n4656 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_357), .QN() );
  DFF_X2 _f_permutation__out_reg_730_  ( .D(_f_permutation__n4657 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_358), .QN() );
  DFF_X2 _f_permutation__out_reg_729_  ( .D(_f_permutation__n4658 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_359), .QN() );
  DFF_X2 _f_permutation__out_reg_728_  ( .D(_f_permutation__n4659 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_360), .QN() );
  DFF_X2 _f_permutation__out_reg_727_  ( .D(_f_permutation__n4660 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_361), .QN() );
  DFF_X2 _f_permutation__out_reg_726_  ( .D(_f_permutation__n4661 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_362), .QN() );
  DFF_X2 _f_permutation__out_reg_725_  ( .D(_f_permutation__n4662 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_363), .QN() );
  DFF_X2 _f_permutation__out_reg_724_  ( .D(_f_permutation__n4663 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_364), .QN() );
  DFF_X2 _f_permutation__out_reg_723_  ( .D(_f_permutation__n4664 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_365), .QN() );
  DFF_X2 _f_permutation__out_reg_722_  ( .D(_f_permutation__n4665 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_366), .QN() );
  DFF_X2 _f_permutation__out_reg_721_  ( .D(_f_permutation__n4666 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_367), .QN() );
  DFF_X2 _f_permutation__out_reg_720_  ( .D(_f_permutation__n4667 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_368), .QN() );
  DFF_X2 _f_permutation__out_reg_719_  ( .D(_f_permutation__n4668 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_369), .QN() );
  DFF_X2 _f_permutation__out_reg_718_  ( .D(_f_permutation__n4669 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_370), .QN() );
  DFF_X2 _f_permutation__out_reg_717_  ( .D(_f_permutation__n4670 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_371), .QN() );
  DFF_X2 _f_permutation__out_reg_716_  ( .D(_f_permutation__n4671 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_372), .QN() );
  DFF_X2 _f_permutation__out_reg_715_  ( .D(_f_permutation__n4672 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_373), .QN() );
  DFF_X2 _f_permutation__out_reg_714_  ( .D(_f_permutation__n4673 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_374), .QN() );
  DFF_X2 _f_permutation__out_reg_713_  ( .D(_f_permutation__n4674 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_375), .QN() );
  DFF_X2 _f_permutation__out_reg_712_  ( .D(_f_permutation__n4675 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_376), .QN() );
  DFF_X2 _f_permutation__out_reg_711_  ( .D(_f_permutation__n4676 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_377), .QN() );
  DFF_X2 _f_permutation__out_reg_710_  ( .D(_f_permutation__n4677 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_378), .QN() );
  DFF_X2 _f_permutation__out_reg_709_  ( .D(_f_permutation__n4678 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_379), .QN() );
  DFF_X2 _f_permutation__out_reg_708_  ( .D(_f_permutation__n4679 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_380), .QN() );
  DFF_X2 _f_permutation__out_reg_707_  ( .D(_f_permutation__n4680 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_381), .QN() );
  DFF_X2 _f_permutation__out_reg_706_  ( .D(_f_permutation__n4681 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_382), .QN() );
  DFF_X2 _f_permutation__out_reg_705_  ( .D(_f_permutation__n4682 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_383), .QN() );
  DFF_X2 _f_permutation__out_reg_704_  ( .D(_f_permutation__n4683 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_384), .QN() );
  DFF_X2 _f_permutation__out_reg_703_  ( .D(_f_permutation__n4684 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_385), .QN() );
  DFF_X2 _f_permutation__out_reg_702_  ( .D(_f_permutation__n4685 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_386), .QN() );
  DFF_X2 _f_permutation__out_reg_701_  ( .D(_f_permutation__n4686 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_387), .QN() );
  DFF_X2 _f_permutation__out_reg_700_  ( .D(_f_permutation__n4687 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_388), .QN() );
  DFF_X2 _f_permutation__out_reg_699_  ( .D(_f_permutation__n4688 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_389), .QN() );
  DFF_X2 _f_permutation__out_reg_698_  ( .D(_f_permutation__n4689 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_390), .QN() );
  DFF_X2 _f_permutation__out_reg_697_  ( .D(_f_permutation__n4690 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_391), .QN() );
  DFF_X2 _f_permutation__out_reg_696_  ( .D(_f_permutation__n4691 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_392), .QN() );
  DFF_X2 _f_permutation__out_reg_695_  ( .D(_f_permutation__n4692 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_393), .QN() );
  DFF_X2 _f_permutation__out_reg_694_  ( .D(_f_permutation__n4693 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_394), .QN() );
  DFF_X2 _f_permutation__out_reg_693_  ( .D(_f_permutation__n4694 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_395), .QN() );
  DFF_X2 _f_permutation__out_reg_692_  ( .D(_f_permutation__n4695 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_396), .QN() );
  DFF_X2 _f_permutation__out_reg_691_  ( .D(_f_permutation__n4696 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_397), .QN() );
  DFF_X2 _f_permutation__out_reg_690_  ( .D(_f_permutation__n4697 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_398), .QN() );
  DFF_X2 _f_permutation__out_reg_689_  ( .D(_f_permutation__n4698 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_399), .QN() );
  DFF_X2 _f_permutation__out_reg_688_  ( .D(_f_permutation__n4699 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_400), .QN() );
  DFF_X2 _f_permutation__out_reg_687_  ( .D(_f_permutation__n4700 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_401), .QN() );
  DFF_X2 _f_permutation__out_reg_686_  ( .D(_f_permutation__n4701 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_402), .QN() );
  DFF_X2 _f_permutation__out_reg_685_  ( .D(_f_permutation__n4702 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_403), .QN() );
  DFF_X2 _f_permutation__out_reg_684_  ( .D(_f_permutation__n4703 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_404), .QN() );
  DFF_X2 _f_permutation__out_reg_683_  ( .D(_f_permutation__n4704 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_405), .QN() );
  DFF_X2 _f_permutation__out_reg_682_  ( .D(_f_permutation__n4705 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_406), .QN() );
  DFF_X2 _f_permutation__out_reg_681_  ( .D(_f_permutation__n4706 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_407), .QN() );
  DFF_X2 _f_permutation__out_reg_680_  ( .D(_f_permutation__n4707 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_408), .QN() );
  DFF_X2 _f_permutation__out_reg_679_  ( .D(_f_permutation__n4708 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_409), .QN() );
  DFF_X2 _f_permutation__out_reg_678_  ( .D(_f_permutation__n4709 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_410), .QN() );
  DFF_X2 _f_permutation__out_reg_677_  ( .D(_f_permutation__n4710 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_411), .QN() );
  DFF_X2 _f_permutation__out_reg_676_  ( .D(_f_permutation__n4711 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_412), .QN() );
  DFF_X2 _f_permutation__out_reg_675_  ( .D(_f_permutation__n4712 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_413), .QN() );
  DFF_X2 _f_permutation__out_reg_674_  ( .D(_f_permutation__n4713 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_414), .QN() );
  DFF_X2 _f_permutation__out_reg_673_  ( .D(_f_permutation__n4714 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_415), .QN() );
  DFF_X2 _f_permutation__out_reg_672_  ( .D(_f_permutation__n4715 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_416), .QN() );
  DFF_X2 _f_permutation__out_reg_671_  ( .D(_f_permutation__n4716 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_417), .QN() );
  DFF_X2 _f_permutation__out_reg_670_  ( .D(_f_permutation__n4717 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_418), .QN() );
  DFF_X2 _f_permutation__out_reg_669_  ( .D(_f_permutation__n4718 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_419), .QN() );
  DFF_X2 _f_permutation__out_reg_668_  ( .D(_f_permutation__n4719 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_420), .QN() );
  DFF_X2 _f_permutation__out_reg_667_  ( .D(_f_permutation__n4720 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_421), .QN() );
  DFF_X2 _f_permutation__out_reg_666_  ( .D(_f_permutation__n4721 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_422), .QN() );
  DFF_X2 _f_permutation__out_reg_665_  ( .D(_f_permutation__n4722 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_423), .QN() );
  DFF_X2 _f_permutation__out_reg_664_  ( .D(_f_permutation__n4723 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_424), .QN() );
  DFF_X2 _f_permutation__out_reg_663_  ( .D(_f_permutation__n4724 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_425), .QN() );
  DFF_X2 _f_permutation__out_reg_662_  ( .D(_f_permutation__n4725 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_426), .QN() );
  DFF_X2 _f_permutation__out_reg_661_  ( .D(_f_permutation__n4726 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_427), .QN() );
  DFF_X2 _f_permutation__out_reg_660_  ( .D(_f_permutation__n4727 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_428), .QN() );
  DFF_X2 _f_permutation__out_reg_659_  ( .D(_f_permutation__n4728 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_429), .QN() );
  DFF_X2 _f_permutation__out_reg_658_  ( .D(_f_permutation__n4729 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_430), .QN() );
  DFF_X2 _f_permutation__out_reg_657_  ( .D(_f_permutation__n4730 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_431), .QN() );
  DFF_X2 _f_permutation__out_reg_656_  ( .D(_f_permutation__n4731 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_432), .QN() );
  DFF_X2 _f_permutation__out_reg_655_  ( .D(_f_permutation__n4732 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_433), .QN() );
  DFF_X2 _f_permutation__out_reg_654_  ( .D(_f_permutation__n4733 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_434), .QN() );
  DFF_X2 _f_permutation__out_reg_653_  ( .D(_f_permutation__n4734 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_435), .QN() );
  DFF_X2 _f_permutation__out_reg_652_  ( .D(_f_permutation__n4735 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_436), .QN() );
  DFF_X2 _f_permutation__out_reg_651_  ( .D(_f_permutation__n4736 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_437), .QN() );
  DFF_X2 _f_permutation__out_reg_650_  ( .D(_f_permutation__n4737 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_438), .QN() );
  DFF_X2 _f_permutation__out_reg_649_  ( .D(_f_permutation__n4738 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_439), .QN() );
  DFF_X2 _f_permutation__out_reg_648_  ( .D(_f_permutation__n4739 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_440), .QN() );
  DFF_X2 _f_permutation__out_reg_647_  ( .D(_f_permutation__n4740 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_441), .QN() );
  DFF_X2 _f_permutation__out_reg_646_  ( .D(_f_permutation__n4741 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_442), .QN() );
  DFF_X2 _f_permutation__out_reg_645_  ( .D(_f_permutation__n4742 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_443), .QN() );
  DFF_X2 _f_permutation__out_reg_644_  ( .D(_f_permutation__n4743 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_444), .QN() );
  DFF_X2 _f_permutation__out_reg_643_  ( .D(_f_permutation__n4744 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_445), .QN() );
  DFF_X2 _f_permutation__out_reg_642_  ( .D(_f_permutation__n4745 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_446), .QN() );
  DFF_X2 _f_permutation__out_reg_641_  ( .D(_f_permutation__n4746 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_447), .QN() );
  DFF_X2 _f_permutation__out_reg_640_  ( .D(_f_permutation__n4747 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_448), .QN() );
  DFF_X2 _f_permutation__out_reg_639_  ( .D(_f_permutation__n4748 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_449), .QN() );
  DFF_X2 _f_permutation__out_reg_638_  ( .D(_f_permutation__n4749 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_450), .QN() );
  DFF_X2 _f_permutation__out_reg_637_  ( .D(_f_permutation__n4750 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_451), .QN() );
  DFF_X2 _f_permutation__out_reg_636_  ( .D(_f_permutation__n4751 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_452), .QN() );
  DFF_X2 _f_permutation__out_reg_635_  ( .D(_f_permutation__n4752 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_453), .QN() );
  DFF_X2 _f_permutation__out_reg_634_  ( .D(_f_permutation__n4753 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_454), .QN() );
  DFF_X2 _f_permutation__out_reg_633_  ( .D(_f_permutation__n4754 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_455), .QN() );
  DFF_X2 _f_permutation__out_reg_632_  ( .D(_f_permutation__n4755 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_456), .QN() );
  DFF_X2 _f_permutation__out_reg_631_  ( .D(_f_permutation__n4756 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_457), .QN() );
  DFF_X2 _f_permutation__out_reg_630_  ( .D(_f_permutation__n4757 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_458), .QN() );
  DFF_X2 _f_permutation__out_reg_629_  ( .D(_f_permutation__n4758 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_459), .QN() );
  DFF_X2 _f_permutation__out_reg_628_  ( .D(_f_permutation__n4759 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_460), .QN() );
  DFF_X2 _f_permutation__out_reg_627_  ( .D(_f_permutation__n4760 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_461), .QN() );
  DFF_X2 _f_permutation__out_reg_626_  ( .D(_f_permutation__n4761 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_462), .QN() );
  DFF_X2 _f_permutation__out_reg_625_  ( .D(_f_permutation__n4762 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_463), .QN() );
  DFF_X2 _f_permutation__out_reg_624_  ( .D(_f_permutation__n4763 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_464), .QN() );
  DFF_X2 _f_permutation__out_reg_623_  ( .D(_f_permutation__n4764 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_465), .QN() );
  DFF_X2 _f_permutation__out_reg_622_  ( .D(_f_permutation__n4765 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_466), .QN() );
  DFF_X2 _f_permutation__out_reg_621_  ( .D(_f_permutation__n4766 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_467), .QN() );
  DFF_X2 _f_permutation__out_reg_620_  ( .D(_f_permutation__n4767 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_468), .QN() );
  DFF_X2 _f_permutation__out_reg_619_  ( .D(_f_permutation__n4768 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_469), .QN() );
  DFF_X2 _f_permutation__out_reg_618_  ( .D(_f_permutation__n4769 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_470), .QN() );
  DFF_X2 _f_permutation__out_reg_617_  ( .D(_f_permutation__n4770 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_471), .QN() );
  DFF_X2 _f_permutation__out_reg_616_  ( .D(_f_permutation__n4771 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_472), .QN() );
  DFF_X2 _f_permutation__out_reg_615_  ( .D(_f_permutation__n4772 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_473), .QN() );
  DFF_X2 _f_permutation__out_reg_614_  ( .D(_f_permutation__n4773 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_474), .QN() );
  DFF_X2 _f_permutation__out_reg_613_  ( .D(_f_permutation__n4774 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_475), .QN() );
  DFF_X2 _f_permutation__out_reg_612_  ( .D(_f_permutation__n4775 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_476), .QN() );
  DFF_X2 _f_permutation__out_reg_611_  ( .D(_f_permutation__n4776 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_477), .QN() );
  DFF_X2 _f_permutation__out_reg_610_  ( .D(_f_permutation__n4777 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_478), .QN() );
  DFF_X2 _f_permutation__out_reg_609_  ( .D(_f_permutation__n4778 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_479), .QN() );
  DFF_X2 _f_permutation__out_reg_608_  ( .D(_f_permutation__n4779 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_480), .QN() );
  DFF_X2 _f_permutation__out_reg_607_  ( .D(_f_permutation__n4780 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_481), .QN() );
  DFF_X2 _f_permutation__out_reg_606_  ( .D(_f_permutation__n4781 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_482), .QN() );
  DFF_X2 _f_permutation__out_reg_605_  ( .D(_f_permutation__n4782 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_483), .QN() );
  DFF_X2 _f_permutation__out_reg_604_  ( .D(_f_permutation__n4783 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_484), .QN() );
  DFF_X2 _f_permutation__out_reg_603_  ( .D(_f_permutation__n4784 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_485), .QN() );
  DFF_X2 _f_permutation__out_reg_602_  ( .D(_f_permutation__n4785 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_486), .QN() );
  DFF_X2 _f_permutation__out_reg_601_  ( .D(_f_permutation__n4786 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_487), .QN() );
  DFF_X2 _f_permutation__out_reg_600_  ( .D(_f_permutation__n4787 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_488), .QN() );
  DFF_X2 _f_permutation__out_reg_599_  ( .D(_f_permutation__n4788 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_489), .QN() );
  DFF_X2 _f_permutation__out_reg_598_  ( .D(_f_permutation__n4789 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_490), .QN() );
  DFF_X2 _f_permutation__out_reg_597_  ( .D(_f_permutation__n4790 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_491), .QN() );
  DFF_X2 _f_permutation__out_reg_596_  ( .D(_f_permutation__n4791 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_492), .QN() );
  DFF_X2 _f_permutation__out_reg_595_  ( .D(_f_permutation__n4792 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_493), .QN() );
  DFF_X2 _f_permutation__out_reg_594_  ( .D(_f_permutation__n4793 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_494), .QN() );
  DFF_X2 _f_permutation__out_reg_593_  ( .D(_f_permutation__n4794 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_495), .QN() );
  DFF_X2 _f_permutation__out_reg_592_  ( .D(_f_permutation__n4795 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_496), .QN() );
  DFF_X2 _f_permutation__out_reg_591_  ( .D(_f_permutation__n4796 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_497), .QN() );
  DFF_X2 _f_permutation__out_reg_590_  ( .D(_f_permutation__n4797 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_498), .QN() );
  DFF_X2 _f_permutation__out_reg_589_  ( .D(_f_permutation__n4798 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_499), .QN() );
  DFF_X2 _f_permutation__out_reg_588_  ( .D(_f_permutation__n4799 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_500), .QN() );
  DFF_X2 _f_permutation__out_reg_587_  ( .D(_f_permutation__n4800 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_501), .QN() );
  DFF_X2 _f_permutation__out_reg_586_  ( .D(_f_permutation__n4801 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_502), .QN() );
  DFF_X2 _f_permutation__out_reg_585_  ( .D(_f_permutation__n4802 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_503), .QN() );
  DFF_X2 _f_permutation__out_reg_584_  ( .D(_f_permutation__n4803 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_504), .QN() );
  DFF_X2 _f_permutation__out_reg_583_  ( .D(_f_permutation__n4804 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_505), .QN() );
  DFF_X2 _f_permutation__out_reg_582_  ( .D(_f_permutation__n4805 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_506), .QN() );
  DFF_X2 _f_permutation__out_reg_581_  ( .D(_f_permutation__n4806 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_507), .QN() );
  DFF_X2 _f_permutation__out_reg_580_  ( .D(_f_permutation__n4807 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_508), .QN() );
  DFF_X2 _f_permutation__out_reg_579_  ( .D(_f_permutation__n4808 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_509), .QN() );
  DFF_X2 _f_permutation__out_reg_578_  ( .D(_f_permutation__n4809 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_510), .QN() );
  DFF_X2 _f_permutation__out_reg_577_  ( .D(_f_permutation__n4810 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_511), .QN() );
  DFF_X2 _f_permutation__out_reg_576_  ( .D(_f_permutation__n4811 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_512), .QN() );
  DFF_X2 _f_permutation__out_reg_575_  ( .D(_f_permutation__n4812 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_513), .QN() );
  DFF_X2 _f_permutation__out_reg_574_  ( .D(_f_permutation__n4813 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_514), .QN() );
  DFF_X2 _f_permutation__out_reg_573_  ( .D(_f_permutation__n4814 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_515), .QN() );
  DFF_X2 _f_permutation__out_reg_572_  ( .D(_f_permutation__n4815 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_516), .QN() );
  DFF_X2 _f_permutation__out_reg_571_  ( .D(_f_permutation__n4816 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_517), .QN() );
  DFF_X2 _f_permutation__out_reg_570_  ( .D(_f_permutation__n4817 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_518), .QN() );
  DFF_X2 _f_permutation__out_reg_569_  ( .D(_f_permutation__n4818 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_519), .QN() );
  DFF_X2 _f_permutation__out_reg_568_  ( .D(_f_permutation__n4819 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_520), .QN() );
  DFF_X2 _f_permutation__out_reg_567_  ( .D(_f_permutation__n4820 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_521), .QN() );
  DFF_X2 _f_permutation__out_reg_566_  ( .D(_f_permutation__n4821 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_522), .QN() );
  DFF_X2 _f_permutation__out_reg_565_  ( .D(_f_permutation__n4822 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_523), .QN() );
  DFF_X2 _f_permutation__out_reg_564_  ( .D(_f_permutation__n4823 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_524), .QN() );
  DFF_X2 _f_permutation__out_reg_563_  ( .D(_f_permutation__n4824 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_525), .QN() );
  DFF_X2 _f_permutation__out_reg_562_  ( .D(_f_permutation__n4825 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_526), .QN() );
  DFF_X2 _f_permutation__out_reg_561_  ( .D(_f_permutation__n4826 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_527), .QN() );
  DFF_X2 _f_permutation__out_reg_560_  ( .D(_f_permutation__n4827 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_528), .QN() );
  DFF_X2 _f_permutation__out_reg_559_  ( .D(_f_permutation__n4828 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_529), .QN() );
  DFF_X2 _f_permutation__out_reg_558_  ( .D(_f_permutation__n4829 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_530), .QN() );
  DFF_X2 _f_permutation__out_reg_557_  ( .D(_f_permutation__n4830 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_531), .QN() );
  DFF_X2 _f_permutation__out_reg_556_  ( .D(_f_permutation__n4831 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_532), .QN() );
  DFF_X2 _f_permutation__out_reg_555_  ( .D(_f_permutation__n4832 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_533), .QN() );
  DFF_X2 _f_permutation__out_reg_554_  ( .D(_f_permutation__n4833 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_534), .QN() );
  DFF_X2 _f_permutation__out_reg_553_  ( .D(_f_permutation__n4834 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_535), .QN() );
  DFF_X2 _f_permutation__out_reg_552_  ( .D(_f_permutation__n4835 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_536), .QN() );
  DFF_X2 _f_permutation__out_reg_551_  ( .D(_f_permutation__n4836 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_537), .QN() );
  DFF_X2 _f_permutation__out_reg_550_  ( .D(_f_permutation__n4837 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_538), .QN() );
  DFF_X2 _f_permutation__out_reg_549_  ( .D(_f_permutation__n4838 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_539), .QN() );
  DFF_X2 _f_permutation__out_reg_548_  ( .D(_f_permutation__n4839 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_540), .QN() );
  DFF_X2 _f_permutation__out_reg_547_  ( .D(_f_permutation__n4840 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_541), .QN() );
  DFF_X2 _f_permutation__out_reg_546_  ( .D(_f_permutation__n4841 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_542), .QN() );
  DFF_X2 _f_permutation__out_reg_545_  ( .D(_f_permutation__n4842 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_543), .QN() );
  DFF_X2 _f_permutation__out_reg_544_  ( .D(_f_permutation__n4843 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_544), .QN() );
  DFF_X2 _f_permutation__out_reg_543_  ( .D(_f_permutation__n4844 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_545), .QN() );
  DFF_X2 _f_permutation__out_reg_542_  ( .D(_f_permutation__n4845 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_546), .QN() );
  DFF_X2 _f_permutation__out_reg_541_  ( .D(_f_permutation__n4846 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_547), .QN() );
  DFF_X2 _f_permutation__out_reg_540_  ( .D(_f_permutation__n4847 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_548), .QN() );
  DFF_X2 _f_permutation__out_reg_539_  ( .D(_f_permutation__n4848 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_549), .QN() );
  DFF_X2 _f_permutation__out_reg_538_  ( .D(_f_permutation__n4849 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_550), .QN() );
  DFF_X2 _f_permutation__out_reg_537_  ( .D(_f_permutation__n4850 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_551), .QN() );
  DFF_X2 _f_permutation__out_reg_536_  ( .D(_f_permutation__n4851 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_552), .QN() );
  DFF_X2 _f_permutation__out_reg_535_  ( .D(_f_permutation__n4852 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_553), .QN() );
  DFF_X2 _f_permutation__out_reg_534_  ( .D(_f_permutation__n4853 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_554), .QN() );
  DFF_X2 _f_permutation__out_reg_533_  ( .D(_f_permutation__n4854 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_555), .QN() );
  DFF_X2 _f_permutation__out_reg_532_  ( .D(_f_permutation__n4855 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_556), .QN() );
  DFF_X2 _f_permutation__out_reg_531_  ( .D(_f_permutation__n4856 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_557), .QN() );
  DFF_X2 _f_permutation__out_reg_530_  ( .D(_f_permutation__n4857 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_558), .QN() );
  DFF_X2 _f_permutation__out_reg_529_  ( .D(_f_permutation__n4858 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_559), .QN() );
  DFF_X2 _f_permutation__out_reg_528_  ( .D(_f_permutation__n4859 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_560), .QN() );
  DFF_X2 _f_permutation__out_reg_527_  ( .D(_f_permutation__n4860 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_561), .QN() );
  DFF_X2 _f_permutation__out_reg_526_  ( .D(_f_permutation__n4861 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_562), .QN() );
  DFF_X2 _f_permutation__out_reg_525_  ( .D(_f_permutation__n4862 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_563), .QN() );
  DFF_X2 _f_permutation__out_reg_524_  ( .D(_f_permutation__n4863 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_564), .QN() );
  DFF_X2 _f_permutation__out_reg_523_  ( .D(_f_permutation__n4864 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_565), .QN() );
  DFF_X2 _f_permutation__out_reg_522_  ( .D(_f_permutation__n4865 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_566), .QN() );
  DFF_X2 _f_permutation__out_reg_521_  ( .D(_f_permutation__n4866 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_567), .QN() );
  DFF_X2 _f_permutation__out_reg_520_  ( .D(_f_permutation__n4867 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_568), .QN() );
  DFF_X2 _f_permutation__out_reg_519_  ( .D(_f_permutation__n4868 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_569), .QN() );
  DFF_X2 _f_permutation__out_reg_518_  ( .D(_f_permutation__n4869 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_570), .QN() );
  DFF_X2 _f_permutation__out_reg_517_  ( .D(_f_permutation__n4870 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_571), .QN() );
  DFF_X2 _f_permutation__out_reg_516_  ( .D(_f_permutation__n4871 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_572), .QN() );
  DFF_X2 _f_permutation__out_reg_515_  ( .D(_f_permutation__n4872 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_573), .QN() );
  DFF_X2 _f_permutation__out_reg_514_  ( .D(_f_permutation__n4873 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_574), .QN() );
  DFF_X2 _f_permutation__out_reg_513_  ( .D(_f_permutation__n4874 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_575), .QN() );
  DFF_X2 _f_permutation__out_reg_512_  ( .D(_f_permutation__n4875 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_576), .QN() );
  DFF_X2 _f_permutation__out_reg_511_  ( .D(_f_permutation__n4876 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_577), .QN() );
  DFF_X2 _f_permutation__out_reg_510_  ( .D(_f_permutation__n4877 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_578), .QN() );
  DFF_X2 _f_permutation__out_reg_509_  ( .D(_f_permutation__n4878 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_579), .QN() );
  DFF_X2 _f_permutation__out_reg_508_  ( .D(_f_permutation__n4879 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_580), .QN() );
  DFF_X2 _f_permutation__out_reg_507_  ( .D(_f_permutation__n4880 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_581), .QN() );
  DFF_X2 _f_permutation__out_reg_506_  ( .D(_f_permutation__n4881 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_582), .QN() );
  DFF_X2 _f_permutation__out_reg_505_  ( .D(_f_permutation__n4882 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_583), .QN() );
  DFF_X2 _f_permutation__out_reg_504_  ( .D(_f_permutation__n4883 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_584), .QN() );
  DFF_X2 _f_permutation__out_reg_503_  ( .D(_f_permutation__n4884 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_585), .QN() );
  DFF_X2 _f_permutation__out_reg_502_  ( .D(_f_permutation__n4885 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_586), .QN() );
  DFF_X2 _f_permutation__out_reg_501_  ( .D(_f_permutation__n4886 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_587), .QN() );
  DFF_X2 _f_permutation__out_reg_500_  ( .D(_f_permutation__n4887 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_588), .QN() );
  DFF_X2 _f_permutation__out_reg_499_  ( .D(_f_permutation__n4888 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_589), .QN() );
  DFF_X2 _f_permutation__out_reg_498_  ( .D(_f_permutation__n4889 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_590), .QN() );
  DFF_X2 _f_permutation__out_reg_497_  ( .D(_f_permutation__n4890 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_591), .QN() );
  DFF_X2 _f_permutation__out_reg_496_  ( .D(_f_permutation__n4891 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_592), .QN() );
  DFF_X2 _f_permutation__out_reg_495_  ( .D(_f_permutation__n4892 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_593), .QN() );
  DFF_X2 _f_permutation__out_reg_494_  ( .D(_f_permutation__n4893 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_594), .QN() );
  DFF_X2 _f_permutation__out_reg_493_  ( .D(_f_permutation__n4894 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_595), .QN() );
  DFF_X2 _f_permutation__out_reg_492_  ( .D(_f_permutation__n4895 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_596), .QN() );
  DFF_X2 _f_permutation__out_reg_491_  ( .D(_f_permutation__n4896 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_597), .QN() );
  DFF_X2 _f_permutation__out_reg_490_  ( .D(_f_permutation__n4897 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_598), .QN() );
  DFF_X2 _f_permutation__out_reg_489_  ( .D(_f_permutation__n4898 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_599), .QN() );
  DFF_X2 _f_permutation__out_reg_488_  ( .D(_f_permutation__n4899 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_600), .QN() );
  DFF_X2 _f_permutation__out_reg_487_  ( .D(_f_permutation__n4900 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_601), .QN() );
  DFF_X2 _f_permutation__out_reg_486_  ( .D(_f_permutation__n4901 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_602), .QN() );
  DFF_X2 _f_permutation__out_reg_485_  ( .D(_f_permutation__n4902 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_603), .QN() );
  DFF_X2 _f_permutation__out_reg_484_  ( .D(_f_permutation__n4903 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_604), .QN() );
  DFF_X2 _f_permutation__out_reg_483_  ( .D(_f_permutation__n4904 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_605), .QN() );
  DFF_X2 _f_permutation__out_reg_482_  ( .D(_f_permutation__n4905 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_606), .QN() );
  DFF_X2 _f_permutation__out_reg_481_  ( .D(_f_permutation__n4906 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_607), .QN() );
  DFF_X2 _f_permutation__out_reg_480_  ( .D(_f_permutation__n4907 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_608), .QN() );
  DFF_X2 _f_permutation__out_reg_479_  ( .D(_f_permutation__n4908 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_609), .QN() );
  DFF_X2 _f_permutation__out_reg_478_  ( .D(_f_permutation__n4909 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_610), .QN() );
  DFF_X2 _f_permutation__out_reg_477_  ( .D(_f_permutation__n4910 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_611), .QN() );
  DFF_X2 _f_permutation__out_reg_476_  ( .D(_f_permutation__n4911 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_612), .QN() );
  DFF_X2 _f_permutation__out_reg_475_  ( .D(_f_permutation__n4912 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_613), .QN() );
  DFF_X2 _f_permutation__out_reg_474_  ( .D(_f_permutation__n4913 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_614), .QN() );
  DFF_X2 _f_permutation__out_reg_473_  ( .D(_f_permutation__n4914 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_615), .QN() );
  DFF_X2 _f_permutation__out_reg_472_  ( .D(_f_permutation__n4915 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_616), .QN() );
  DFF_X2 _f_permutation__out_reg_471_  ( .D(_f_permutation__n4916 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_617), .QN() );
  DFF_X2 _f_permutation__out_reg_470_  ( .D(_f_permutation__n4917 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_618), .QN() );
  DFF_X2 _f_permutation__out_reg_469_  ( .D(_f_permutation__n4918 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_619), .QN() );
  DFF_X2 _f_permutation__out_reg_468_  ( .D(_f_permutation__n4919 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_620), .QN() );
  DFF_X2 _f_permutation__out_reg_467_  ( .D(_f_permutation__n4920 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_621), .QN() );
  DFF_X2 _f_permutation__out_reg_466_  ( .D(_f_permutation__n4921 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_622), .QN() );
  DFF_X2 _f_permutation__out_reg_465_  ( .D(_f_permutation__n4922 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_623), .QN() );
  DFF_X2 _f_permutation__out_reg_464_  ( .D(_f_permutation__n4923 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_624), .QN() );
  DFF_X2 _f_permutation__out_reg_463_  ( .D(_f_permutation__n4924 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_625), .QN() );
  DFF_X2 _f_permutation__out_reg_462_  ( .D(_f_permutation__n4925 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_626), .QN() );
  DFF_X2 _f_permutation__out_reg_461_  ( .D(_f_permutation__n4926 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_627), .QN() );
  DFF_X2 _f_permutation__out_reg_460_  ( .D(_f_permutation__n4927 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_628), .QN() );
  DFF_X2 _f_permutation__out_reg_459_  ( .D(_f_permutation__n4928 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_629), .QN() );
  DFF_X2 _f_permutation__out_reg_458_  ( .D(_f_permutation__n4929 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_630), .QN() );
  DFF_X2 _f_permutation__out_reg_457_  ( .D(_f_permutation__n4930 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_631), .QN() );
  DFF_X2 _f_permutation__out_reg_456_  ( .D(_f_permutation__n4931 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_632), .QN() );
  DFF_X2 _f_permutation__out_reg_455_  ( .D(_f_permutation__n4932 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_633), .QN() );
  DFF_X2 _f_permutation__out_reg_454_  ( .D(_f_permutation__n4933 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_634), .QN() );
  DFF_X2 _f_permutation__out_reg_453_  ( .D(_f_permutation__n4934 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_635), .QN() );
  DFF_X2 _f_permutation__out_reg_452_  ( .D(_f_permutation__n4935 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_636), .QN() );
  DFF_X2 _f_permutation__out_reg_451_  ( .D(_f_permutation__n4936 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_637), .QN() );
  DFF_X2 _f_permutation__out_reg_450_  ( .D(_f_permutation__n4937 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_638), .QN() );
  DFF_X2 _f_permutation__out_reg_449_  ( .D(_f_permutation__n4938 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_639), .QN() );
  DFF_X2 _f_permutation__out_reg_448_  ( .D(_f_permutation__n4939 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_640), .QN() );
  DFF_X2 _f_permutation__out_reg_447_  ( .D(_f_permutation__n4940 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_641), .QN() );
  DFF_X2 _f_permutation__out_reg_446_  ( .D(_f_permutation__n4941 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_642), .QN() );
  DFF_X2 _f_permutation__out_reg_445_  ( .D(_f_permutation__n4942 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_643), .QN() );
  DFF_X2 _f_permutation__out_reg_444_  ( .D(_f_permutation__n4943 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_644), .QN() );
  DFF_X2 _f_permutation__out_reg_443_  ( .D(_f_permutation__n4944 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_645), .QN() );
  DFF_X2 _f_permutation__out_reg_442_  ( .D(_f_permutation__n4945 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_646), .QN() );
  DFF_X2 _f_permutation__out_reg_441_  ( .D(_f_permutation__n4946 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_647), .QN() );
  DFF_X2 _f_permutation__out_reg_440_  ( .D(_f_permutation__n4947 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_648), .QN() );
  DFF_X2 _f_permutation__out_reg_439_  ( .D(_f_permutation__n4948 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_649), .QN() );
  DFF_X2 _f_permutation__out_reg_438_  ( .D(_f_permutation__n4949 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_650), .QN() );
  DFF_X2 _f_permutation__out_reg_437_  ( .D(_f_permutation__n4950 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_651), .QN() );
  DFF_X2 _f_permutation__out_reg_436_  ( .D(_f_permutation__n4951 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_652), .QN() );
  DFF_X2 _f_permutation__out_reg_435_  ( .D(_f_permutation__n4952 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_653), .QN() );
  DFF_X2 _f_permutation__out_reg_434_  ( .D(_f_permutation__n4953 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_654), .QN() );
  DFF_X2 _f_permutation__out_reg_433_  ( .D(_f_permutation__n4954 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_655), .QN() );
  DFF_X2 _f_permutation__out_reg_432_  ( .D(_f_permutation__n4955 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_656), .QN() );
  DFF_X2 _f_permutation__out_reg_431_  ( .D(_f_permutation__n4956 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_657), .QN() );
  DFF_X2 _f_permutation__out_reg_430_  ( .D(_f_permutation__n4957 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_658), .QN() );
  DFF_X2 _f_permutation__out_reg_429_  ( .D(_f_permutation__n4958 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_659), .QN() );
  DFF_X2 _f_permutation__out_reg_428_  ( .D(_f_permutation__n4959 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_660), .QN() );
  DFF_X2 _f_permutation__out_reg_427_  ( .D(_f_permutation__n4960 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_661), .QN() );
  DFF_X2 _f_permutation__out_reg_426_  ( .D(_f_permutation__n4961 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_662), .QN() );
  DFF_X2 _f_permutation__out_reg_425_  ( .D(_f_permutation__n4962 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_663), .QN() );
  DFF_X2 _f_permutation__out_reg_424_  ( .D(_f_permutation__n4963 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_664), .QN() );
  DFF_X2 _f_permutation__out_reg_423_  ( .D(_f_permutation__n4964 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_665), .QN() );
  DFF_X2 _f_permutation__out_reg_422_  ( .D(_f_permutation__n4965 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_666), .QN() );
  DFF_X2 _f_permutation__out_reg_421_  ( .D(_f_permutation__n4966 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_667), .QN() );
  DFF_X2 _f_permutation__out_reg_420_  ( .D(_f_permutation__n4967 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_668), .QN() );
  DFF_X2 _f_permutation__out_reg_419_  ( .D(_f_permutation__n4968 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_669), .QN() );
  DFF_X2 _f_permutation__out_reg_418_  ( .D(_f_permutation__n4969 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_670), .QN() );
  DFF_X2 _f_permutation__out_reg_417_  ( .D(_f_permutation__n4970 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_671), .QN() );
  DFF_X2 _f_permutation__out_reg_416_  ( .D(_f_permutation__n4971 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_672), .QN() );
  DFF_X2 _f_permutation__out_reg_415_  ( .D(_f_permutation__n4972 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_673), .QN() );
  DFF_X2 _f_permutation__out_reg_414_  ( .D(_f_permutation__n4973 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_674), .QN() );
  DFF_X2 _f_permutation__out_reg_413_  ( .D(_f_permutation__n4974 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_675), .QN() );
  DFF_X2 _f_permutation__out_reg_412_  ( .D(_f_permutation__n4975 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_676), .QN() );
  DFF_X2 _f_permutation__out_reg_411_  ( .D(_f_permutation__n4976 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_677), .QN() );
  DFF_X2 _f_permutation__out_reg_410_  ( .D(_f_permutation__n4977 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_678), .QN() );
  DFF_X2 _f_permutation__out_reg_409_  ( .D(_f_permutation__n4978 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_679), .QN() );
  DFF_X2 _f_permutation__out_reg_408_  ( .D(_f_permutation__n4979 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_680), .QN() );
  DFF_X2 _f_permutation__out_reg_407_  ( .D(_f_permutation__n4980 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_681), .QN() );
  DFF_X2 _f_permutation__out_reg_406_  ( .D(_f_permutation__n4981 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_682), .QN() );
  DFF_X2 _f_permutation__out_reg_405_  ( .D(_f_permutation__n4982 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_683), .QN() );
  DFF_X2 _f_permutation__out_reg_404_  ( .D(_f_permutation__n4983 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_684), .QN() );
  DFF_X2 _f_permutation__out_reg_403_  ( .D(_f_permutation__n4984 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_685), .QN() );
  DFF_X2 _f_permutation__out_reg_402_  ( .D(_f_permutation__n4985 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_686), .QN() );
  DFF_X2 _f_permutation__out_reg_401_  ( .D(_f_permutation__n4986 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_687), .QN() );
  DFF_X2 _f_permutation__out_reg_400_  ( .D(_f_permutation__n4987 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_688), .QN() );
  DFF_X2 _f_permutation__out_reg_399_  ( .D(_f_permutation__n4988 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_689), .QN() );
  DFF_X2 _f_permutation__out_reg_398_  ( .D(_f_permutation__n4989 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_690), .QN() );
  DFF_X2 _f_permutation__out_reg_397_  ( .D(_f_permutation__n4990 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_691), .QN() );
  DFF_X2 _f_permutation__out_reg_396_  ( .D(_f_permutation__n4991 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_692), .QN() );
  DFF_X2 _f_permutation__out_reg_395_  ( .D(_f_permutation__n4992 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_693), .QN() );
  DFF_X2 _f_permutation__out_reg_394_  ( .D(_f_permutation__n4993 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_694), .QN() );
  DFF_X2 _f_permutation__out_reg_393_  ( .D(_f_permutation__n4994 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_695), .QN() );
  DFF_X2 _f_permutation__out_reg_392_  ( .D(_f_permutation__n4995 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_696), .QN() );
  DFF_X2 _f_permutation__out_reg_391_  ( .D(_f_permutation__n4996 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_697), .QN() );
  DFF_X2 _f_permutation__out_reg_390_  ( .D(_f_permutation__n4997 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_698), .QN() );
  DFF_X2 _f_permutation__out_reg_389_  ( .D(_f_permutation__n4998 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_699), .QN() );
  DFF_X2 _f_permutation__out_reg_388_  ( .D(_f_permutation__n4999 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_700), .QN() );
  DFF_X2 _f_permutation__out_reg_387_  ( .D(_f_permutation__n5000 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_701), .QN() );
  DFF_X2 _f_permutation__out_reg_386_  ( .D(_f_permutation__n5001 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_702), .QN() );
  DFF_X2 _f_permutation__out_reg_385_  ( .D(_f_permutation__n5002 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_703), .QN() );
  DFF_X2 _f_permutation__out_reg_384_  ( .D(_f_permutation__n5003 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_704), .QN() );
  DFF_X2 _f_permutation__out_reg_383_  ( .D(_f_permutation__n5004 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_705), .QN() );
  DFF_X2 _f_permutation__out_reg_382_  ( .D(_f_permutation__n5005 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_706), .QN() );
  DFF_X2 _f_permutation__out_reg_381_  ( .D(_f_permutation__n5006 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_707), .QN() );
  DFF_X2 _f_permutation__out_reg_380_  ( .D(_f_permutation__n5007 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_708), .QN() );
  DFF_X2 _f_permutation__out_reg_379_  ( .D(_f_permutation__n5008 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_709), .QN() );
  DFF_X2 _f_permutation__out_reg_378_  ( .D(_f_permutation__n5009 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_710), .QN() );
  DFF_X2 _f_permutation__out_reg_377_  ( .D(_f_permutation__n5010 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_711), .QN() );
  DFF_X2 _f_permutation__out_reg_376_  ( .D(_f_permutation__n5011 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_712), .QN() );
  DFF_X2 _f_permutation__out_reg_375_  ( .D(_f_permutation__n5012 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_713), .QN() );
  DFF_X2 _f_permutation__out_reg_374_  ( .D(_f_permutation__n5013 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_714), .QN() );
  DFF_X2 _f_permutation__out_reg_373_  ( .D(_f_permutation__n5014 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_715), .QN() );
  DFF_X2 _f_permutation__out_reg_372_  ( .D(_f_permutation__n5015 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_716), .QN() );
  DFF_X2 _f_permutation__out_reg_371_  ( .D(_f_permutation__n5016 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_717), .QN() );
  DFF_X2 _f_permutation__out_reg_370_  ( .D(_f_permutation__n5017 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_718), .QN() );
  DFF_X2 _f_permutation__out_reg_369_  ( .D(_f_permutation__n5018 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_719), .QN() );
  DFF_X2 _f_permutation__out_reg_368_  ( .D(_f_permutation__n5019 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_720), .QN() );
  DFF_X2 _f_permutation__out_reg_367_  ( .D(_f_permutation__n5020 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_721), .QN() );
  DFF_X2 _f_permutation__out_reg_366_  ( .D(_f_permutation__n5021 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_722), .QN() );
  DFF_X2 _f_permutation__out_reg_365_  ( .D(_f_permutation__n5022 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_723), .QN() );
  DFF_X2 _f_permutation__out_reg_364_  ( .D(_f_permutation__n5023 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_724), .QN() );
  DFF_X2 _f_permutation__out_reg_363_  ( .D(_f_permutation__n5024 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_725), .QN() );
  DFF_X2 _f_permutation__out_reg_362_  ( .D(_f_permutation__n5025 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_726), .QN() );
  DFF_X2 _f_permutation__out_reg_361_  ( .D(_f_permutation__n5026 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_727), .QN() );
  DFF_X2 _f_permutation__out_reg_360_  ( .D(_f_permutation__n5027 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_728), .QN() );
  DFF_X2 _f_permutation__out_reg_359_  ( .D(_f_permutation__n5028 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_729), .QN() );
  DFF_X2 _f_permutation__out_reg_358_  ( .D(_f_permutation__n5029 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_730), .QN() );
  DFF_X2 _f_permutation__out_reg_357_  ( .D(_f_permutation__n5030 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_731), .QN() );
  DFF_X2 _f_permutation__out_reg_356_  ( .D(_f_permutation__n5031 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_732), .QN() );
  DFF_X2 _f_permutation__out_reg_355_  ( .D(_f_permutation__n5032 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_733), .QN() );
  DFF_X2 _f_permutation__out_reg_354_  ( .D(_f_permutation__n5033 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_734), .QN() );
  DFF_X2 _f_permutation__out_reg_353_  ( .D(_f_permutation__n5034 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_735), .QN() );
  DFF_X2 _f_permutation__out_reg_352_  ( .D(_f_permutation__n5035 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_736), .QN() );
  DFF_X2 _f_permutation__out_reg_351_  ( .D(_f_permutation__n5036 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_737), .QN() );
  DFF_X2 _f_permutation__out_reg_350_  ( .D(_f_permutation__n5037 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_738), .QN() );
  DFF_X2 _f_permutation__out_reg_349_  ( .D(_f_permutation__n5038 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_739), .QN() );
  DFF_X2 _f_permutation__out_reg_348_  ( .D(_f_permutation__n5039 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_740), .QN() );
  DFF_X2 _f_permutation__out_reg_347_  ( .D(_f_permutation__n5040 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_741), .QN() );
  DFF_X2 _f_permutation__out_reg_346_  ( .D(_f_permutation__n5041 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_742), .QN() );
  DFF_X2 _f_permutation__out_reg_345_  ( .D(_f_permutation__n5042 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_743), .QN() );
  DFF_X2 _f_permutation__out_reg_344_  ( .D(_f_permutation__n5043 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_744), .QN() );
  DFF_X2 _f_permutation__out_reg_343_  ( .D(_f_permutation__n5044 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_745), .QN() );
  DFF_X2 _f_permutation__out_reg_342_  ( .D(_f_permutation__n5045 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_746), .QN() );
  DFF_X2 _f_permutation__out_reg_341_  ( .D(_f_permutation__n5046 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_747), .QN() );
  DFF_X2 _f_permutation__out_reg_340_  ( .D(_f_permutation__n5047 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_748), .QN() );
  DFF_X2 _f_permutation__out_reg_339_  ( .D(_f_permutation__n5048 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_749), .QN() );
  DFF_X2 _f_permutation__out_reg_338_  ( .D(_f_permutation__n5049 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_750), .QN() );
  DFF_X2 _f_permutation__out_reg_337_  ( .D(_f_permutation__n5050 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_751), .QN() );
  DFF_X2 _f_permutation__out_reg_336_  ( .D(_f_permutation__n5051 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_752), .QN() );
  DFF_X2 _f_permutation__out_reg_335_  ( .D(_f_permutation__n5052 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_753), .QN() );
  DFF_X2 _f_permutation__out_reg_334_  ( .D(_f_permutation__n5053 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_754), .QN() );
  DFF_X2 _f_permutation__out_reg_333_  ( .D(_f_permutation__n5054 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_755), .QN() );
  DFF_X2 _f_permutation__out_reg_332_  ( .D(_f_permutation__n5055 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_756), .QN() );
  DFF_X2 _f_permutation__out_reg_331_  ( .D(_f_permutation__n5056 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_757), .QN() );
  DFF_X2 _f_permutation__out_reg_330_  ( .D(_f_permutation__n5057 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_758), .QN() );
  DFF_X2 _f_permutation__out_reg_329_  ( .D(_f_permutation__n5058 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_759), .QN() );
  DFF_X2 _f_permutation__out_reg_328_  ( .D(_f_permutation__n5059 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_760), .QN() );
  DFF_X2 _f_permutation__out_reg_327_  ( .D(_f_permutation__n5060 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_761), .QN() );
  DFF_X2 _f_permutation__out_reg_326_  ( .D(_f_permutation__n5061 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_762), .QN() );
  DFF_X2 _f_permutation__out_reg_325_  ( .D(_f_permutation__n5062 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_763), .QN() );
  DFF_X2 _f_permutation__out_reg_324_  ( .D(_f_permutation__n5063 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_764), .QN() );
  DFF_X2 _f_permutation__out_reg_323_  ( .D(_f_permutation__n5064 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_765), .QN() );
  DFF_X2 _f_permutation__out_reg_322_  ( .D(_f_permutation__n5065 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_766), .QN() );
  DFF_X2 _f_permutation__out_reg_321_  ( .D(_f_permutation__n5066 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_767), .QN() );
  DFF_X2 _f_permutation__out_reg_320_  ( .D(_f_permutation__n5067 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_768), .QN() );
  DFF_X2 _f_permutation__out_reg_319_  ( .D(_f_permutation__n5068 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_769), .QN() );
  DFF_X2 _f_permutation__out_reg_318_  ( .D(_f_permutation__n5069 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_770), .QN() );
  DFF_X2 _f_permutation__out_reg_317_  ( .D(_f_permutation__n5070 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_771), .QN() );
  DFF_X2 _f_permutation__out_reg_316_  ( .D(_f_permutation__n5071 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_772), .QN() );
  DFF_X2 _f_permutation__out_reg_315_  ( .D(_f_permutation__n5072 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_773), .QN() );
  DFF_X2 _f_permutation__out_reg_314_  ( .D(_f_permutation__n5073 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_774), .QN() );
  DFF_X2 _f_permutation__out_reg_313_  ( .D(_f_permutation__n5074 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_775), .QN() );
  DFF_X2 _f_permutation__out_reg_312_  ( .D(_f_permutation__n5075 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_776), .QN() );
  DFF_X2 _f_permutation__out_reg_311_  ( .D(_f_permutation__n5076 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_777), .QN() );
  DFF_X2 _f_permutation__out_reg_310_  ( .D(_f_permutation__n5077 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_778), .QN() );
  DFF_X2 _f_permutation__out_reg_309_  ( .D(_f_permutation__n5078 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_779), .QN() );
  DFF_X2 _f_permutation__out_reg_308_  ( .D(_f_permutation__n5079 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_780), .QN() );
  DFF_X2 _f_permutation__out_reg_307_  ( .D(_f_permutation__n5080 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_781), .QN() );
  DFF_X2 _f_permutation__out_reg_306_  ( .D(_f_permutation__n5081 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_782), .QN() );
  DFF_X2 _f_permutation__out_reg_305_  ( .D(_f_permutation__n5082 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_783), .QN() );
  DFF_X2 _f_permutation__out_reg_304_  ( .D(_f_permutation__n5083 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_784), .QN() );
  DFF_X2 _f_permutation__out_reg_303_  ( .D(_f_permutation__n5084 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_785), .QN() );
  DFF_X2 _f_permutation__out_reg_302_  ( .D(_f_permutation__n5085 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_786), .QN() );
  DFF_X2 _f_permutation__out_reg_301_  ( .D(_f_permutation__n5086 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_787), .QN() );
  DFF_X2 _f_permutation__out_reg_300_  ( .D(_f_permutation__n5087 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_788), .QN() );
  DFF_X2 _f_permutation__out_reg_299_  ( .D(_f_permutation__n5088 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_789), .QN() );
  DFF_X2 _f_permutation__out_reg_298_  ( .D(_f_permutation__n5089 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_790), .QN() );
  DFF_X2 _f_permutation__out_reg_297_  ( .D(_f_permutation__n5090 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_791), .QN() );
  DFF_X2 _f_permutation__out_reg_296_  ( .D(_f_permutation__n5091 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_792), .QN() );
  DFF_X2 _f_permutation__out_reg_295_  ( .D(_f_permutation__n5092 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_793), .QN() );
  DFF_X2 _f_permutation__out_reg_294_  ( .D(_f_permutation__n5093 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_794), .QN() );
  DFF_X2 _f_permutation__out_reg_293_  ( .D(_f_permutation__n5094 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_795), .QN() );
  DFF_X2 _f_permutation__out_reg_292_  ( .D(_f_permutation__n5095 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_796), .QN() );
  DFF_X2 _f_permutation__out_reg_291_  ( .D(_f_permutation__n5096 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_797), .QN() );
  DFF_X2 _f_permutation__out_reg_290_  ( .D(_f_permutation__n5097 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_798), .QN() );
  DFF_X2 _f_permutation__out_reg_289_  ( .D(_f_permutation__n5098 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_799), .QN() );
  DFF_X2 _f_permutation__out_reg_288_  ( .D(_f_permutation__n5099 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_800), .QN() );
  DFF_X2 _f_permutation__out_reg_287_  ( .D(_f_permutation__n5100 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_801), .QN() );
  DFF_X2 _f_permutation__out_reg_286_  ( .D(_f_permutation__n5101 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_802), .QN() );
  DFF_X2 _f_permutation__out_reg_285_  ( .D(_f_permutation__n5102 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_803), .QN() );
  DFF_X2 _f_permutation__out_reg_284_  ( .D(_f_permutation__n5103 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_804), .QN() );
  DFF_X2 _f_permutation__out_reg_283_  ( .D(_f_permutation__n5104 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_805), .QN() );
  DFF_X2 _f_permutation__out_reg_282_  ( .D(_f_permutation__n5105 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_806), .QN() );
  DFF_X2 _f_permutation__out_reg_281_  ( .D(_f_permutation__n5106 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_807), .QN() );
  DFF_X2 _f_permutation__out_reg_280_  ( .D(_f_permutation__n5107 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_808), .QN() );
  DFF_X2 _f_permutation__out_reg_279_  ( .D(_f_permutation__n5108 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_809), .QN() );
  DFF_X2 _f_permutation__out_reg_278_  ( .D(_f_permutation__n5109 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_810), .QN() );
  DFF_X2 _f_permutation__out_reg_277_  ( .D(_f_permutation__n5110 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_811), .QN() );
  DFF_X2 _f_permutation__out_reg_276_  ( .D(_f_permutation__n5111 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_812), .QN() );
  DFF_X2 _f_permutation__out_reg_275_  ( .D(_f_permutation__n5112 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_813), .QN() );
  DFF_X2 _f_permutation__out_reg_274_  ( .D(_f_permutation__n5113 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_814), .QN() );
  DFF_X2 _f_permutation__out_reg_273_  ( .D(_f_permutation__n5114 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_815), .QN() );
  DFF_X2 _f_permutation__out_reg_272_  ( .D(_f_permutation__n5115 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_816), .QN() );
  DFF_X2 _f_permutation__out_reg_271_  ( .D(_f_permutation__n5116 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_817), .QN() );
  DFF_X2 _f_permutation__out_reg_270_  ( .D(_f_permutation__n5117 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_818), .QN() );
  DFF_X2 _f_permutation__out_reg_269_  ( .D(_f_permutation__n5118 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_819), .QN() );
  DFF_X2 _f_permutation__out_reg_268_  ( .D(_f_permutation__n5119 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_820), .QN() );
  DFF_X2 _f_permutation__out_reg_267_  ( .D(_f_permutation__n5120 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_821), .QN() );
  DFF_X2 _f_permutation__out_reg_266_  ( .D(_f_permutation__n5121 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_822), .QN() );
  DFF_X2 _f_permutation__out_reg_265_  ( .D(_f_permutation__n5122 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_823), .QN() );
  DFF_X2 _f_permutation__out_reg_264_  ( .D(_f_permutation__n5123 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_824), .QN() );
  DFF_X2 _f_permutation__out_reg_263_  ( .D(_f_permutation__n5124 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_825), .QN() );
  DFF_X2 _f_permutation__out_reg_262_  ( .D(_f_permutation__n5125 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_826), .QN() );
  DFF_X2 _f_permutation__out_reg_261_  ( .D(_f_permutation__n5126 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_827), .QN() );
  DFF_X2 _f_permutation__out_reg_260_  ( .D(_f_permutation__n5127 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_828), .QN() );
  DFF_X2 _f_permutation__out_reg_259_  ( .D(_f_permutation__n5128 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_829), .QN() );
  DFF_X2 _f_permutation__out_reg_258_  ( .D(_f_permutation__n5129 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_830), .QN() );
  DFF_X2 _f_permutation__out_reg_257_  ( .D(_f_permutation__n5130 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_831), .QN() );
  DFF_X2 _f_permutation__out_reg_256_  ( .D(_f_permutation__n5131 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_832), .QN() );
  DFF_X2 _f_permutation__out_reg_255_  ( .D(_f_permutation__n5132 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_833), .QN() );
  DFF_X2 _f_permutation__out_reg_254_  ( .D(_f_permutation__n5133 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_834), .QN() );
  DFF_X2 _f_permutation__out_reg_253_  ( .D(_f_permutation__n5134 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_835), .QN() );
  DFF_X2 _f_permutation__out_reg_252_  ( .D(_f_permutation__n5135 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_836), .QN() );
  DFF_X2 _f_permutation__out_reg_251_  ( .D(_f_permutation__n5136 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_837), .QN() );
  DFF_X2 _f_permutation__out_reg_250_  ( .D(_f_permutation__n5137 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_838), .QN() );
  DFF_X2 _f_permutation__out_reg_249_  ( .D(_f_permutation__n5138 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_839), .QN() );
  DFF_X2 _f_permutation__out_reg_248_  ( .D(_f_permutation__n5139 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_840), .QN() );
  DFF_X2 _f_permutation__out_reg_247_  ( .D(_f_permutation__n5140 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_841), .QN() );
  DFF_X2 _f_permutation__out_reg_246_  ( .D(_f_permutation__n5141 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_842), .QN() );
  DFF_X2 _f_permutation__out_reg_245_  ( .D(_f_permutation__n5142 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_843), .QN() );
  DFF_X2 _f_permutation__out_reg_244_  ( .D(_f_permutation__n5143 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_844), .QN() );
  DFF_X2 _f_permutation__out_reg_243_  ( .D(_f_permutation__n5144 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_845), .QN() );
  DFF_X2 _f_permutation__out_reg_242_  ( .D(_f_permutation__n5145 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_846), .QN() );
  DFF_X2 _f_permutation__out_reg_241_  ( .D(_f_permutation__n5146 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_847), .QN() );
  DFF_X2 _f_permutation__out_reg_240_  ( .D(_f_permutation__n5147 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_848), .QN() );
  DFF_X2 _f_permutation__out_reg_239_  ( .D(_f_permutation__n5148 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_849), .QN() );
  DFF_X2 _f_permutation__out_reg_238_  ( .D(_f_permutation__n5149 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_850), .QN() );
  DFF_X2 _f_permutation__out_reg_237_  ( .D(_f_permutation__n5150 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_851), .QN() );
  DFF_X2 _f_permutation__out_reg_236_  ( .D(_f_permutation__n5151 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_852), .QN() );
  DFF_X2 _f_permutation__out_reg_235_  ( .D(_f_permutation__n5152 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_853), .QN() );
  DFF_X2 _f_permutation__out_reg_234_  ( .D(_f_permutation__n5153 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_854), .QN() );
  DFF_X2 _f_permutation__out_reg_233_  ( .D(_f_permutation__n5154 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_855), .QN() );
  DFF_X2 _f_permutation__out_reg_232_  ( .D(_f_permutation__n5155 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_856), .QN() );
  DFF_X2 _f_permutation__out_reg_231_  ( .D(_f_permutation__n5156 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_857), .QN() );
  DFF_X2 _f_permutation__out_reg_230_  ( .D(_f_permutation__n5157 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_858), .QN() );
  DFF_X2 _f_permutation__out_reg_229_  ( .D(_f_permutation__n5158 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_859), .QN() );
  DFF_X2 _f_permutation__out_reg_228_  ( .D(_f_permutation__n5159 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_860), .QN() );
  DFF_X2 _f_permutation__out_reg_227_  ( .D(_f_permutation__n5160 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_861), .QN() );
  DFF_X2 _f_permutation__out_reg_226_  ( .D(_f_permutation__n5161 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_862), .QN() );
  DFF_X2 _f_permutation__out_reg_225_  ( .D(_f_permutation__n5162 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_863), .QN() );
  DFF_X2 _f_permutation__out_reg_224_  ( .D(_f_permutation__n5163 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_864), .QN() );
  DFF_X2 _f_permutation__out_reg_223_  ( .D(_f_permutation__n5164 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_865), .QN() );
  DFF_X2 _f_permutation__out_reg_222_  ( .D(_f_permutation__n5165 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_866), .QN() );
  DFF_X2 _f_permutation__out_reg_221_  ( .D(_f_permutation__n5166 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_867), .QN() );
  DFF_X2 _f_permutation__out_reg_220_  ( .D(_f_permutation__n5167 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_868), .QN() );
  DFF_X2 _f_permutation__out_reg_219_  ( .D(_f_permutation__n5168 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_869), .QN() );
  DFF_X2 _f_permutation__out_reg_218_  ( .D(_f_permutation__n5169 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_870), .QN() );
  DFF_X2 _f_permutation__out_reg_217_  ( .D(_f_permutation__n5170 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_871), .QN() );
  DFF_X2 _f_permutation__out_reg_216_  ( .D(_f_permutation__n5171 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_872), .QN() );
  DFF_X2 _f_permutation__out_reg_215_  ( .D(_f_permutation__n5172 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_873), .QN() );
  DFF_X2 _f_permutation__out_reg_214_  ( .D(_f_permutation__n5173 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_874), .QN() );
  DFF_X2 _f_permutation__out_reg_213_  ( .D(_f_permutation__n5174 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_875), .QN() );
  DFF_X2 _f_permutation__out_reg_212_  ( .D(_f_permutation__n5175 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_876), .QN() );
  DFF_X2 _f_permutation__out_reg_211_  ( .D(_f_permutation__n5176 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_877), .QN() );
  DFF_X2 _f_permutation__out_reg_210_  ( .D(_f_permutation__n5177 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_878), .QN() );
  DFF_X2 _f_permutation__out_reg_209_  ( .D(_f_permutation__n5178 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_879), .QN() );
  DFF_X2 _f_permutation__out_reg_208_  ( .D(_f_permutation__n5179 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_880), .QN() );
  DFF_X2 _f_permutation__out_reg_207_  ( .D(_f_permutation__n5180 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_881), .QN() );
  DFF_X2 _f_permutation__out_reg_206_  ( .D(_f_permutation__n5181 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_882), .QN() );
  DFF_X2 _f_permutation__out_reg_205_  ( .D(_f_permutation__n5182 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_883), .QN() );
  DFF_X2 _f_permutation__out_reg_204_  ( .D(_f_permutation__n5183 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_884), .QN() );
  DFF_X2 _f_permutation__out_reg_203_  ( .D(_f_permutation__n5184 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_885), .QN() );
  DFF_X2 _f_permutation__out_reg_202_  ( .D(_f_permutation__n5185 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_886), .QN() );
  DFF_X2 _f_permutation__out_reg_201_  ( .D(_f_permutation__n5186 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_887), .QN() );
  DFF_X2 _f_permutation__out_reg_200_  ( .D(_f_permutation__n5187 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_888), .QN() );
  DFF_X2 _f_permutation__out_reg_199_  ( .D(_f_permutation__n5188 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_889), .QN() );
  DFF_X2 _f_permutation__out_reg_198_  ( .D(_f_permutation__n5189 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_890), .QN() );
  DFF_X2 _f_permutation__out_reg_197_  ( .D(_f_permutation__n5190 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_891), .QN() );
  DFF_X2 _f_permutation__out_reg_196_  ( .D(_f_permutation__n5191 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_892), .QN() );
  DFF_X2 _f_permutation__out_reg_195_  ( .D(_f_permutation__n5192 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_893), .QN() );
  DFF_X2 _f_permutation__out_reg_194_  ( .D(_f_permutation__n5193 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_894), .QN() );
  DFF_X2 _f_permutation__out_reg_193_  ( .D(_f_permutation__n5194 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_895), .QN() );
  DFF_X2 _f_permutation__out_reg_192_  ( .D(_f_permutation__n5195 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_896), .QN() );
  DFF_X2 _f_permutation__out_reg_191_  ( .D(_f_permutation__n5196 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_897), .QN() );
  DFF_X2 _f_permutation__out_reg_190_  ( .D(_f_permutation__n5197 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_898), .QN() );
  DFF_X2 _f_permutation__out_reg_189_  ( .D(_f_permutation__n5198 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_899), .QN() );
  DFF_X2 _f_permutation__out_reg_188_  ( .D(_f_permutation__n5199 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_900), .QN() );
  DFF_X2 _f_permutation__out_reg_187_  ( .D(_f_permutation__n5200 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_901), .QN() );
  DFF_X2 _f_permutation__out_reg_186_  ( .D(_f_permutation__n5201 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_902), .QN() );
  DFF_X2 _f_permutation__out_reg_185_  ( .D(_f_permutation__n5202 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_903), .QN() );
  DFF_X2 _f_permutation__out_reg_184_  ( .D(_f_permutation__n5203 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_904), .QN() );
  DFF_X2 _f_permutation__out_reg_183_  ( .D(_f_permutation__n5204 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_905), .QN() );
  DFF_X2 _f_permutation__out_reg_182_  ( .D(_f_permutation__n5205 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_906), .QN() );
  DFF_X2 _f_permutation__out_reg_181_  ( .D(_f_permutation__n5206 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_907), .QN() );
  DFF_X2 _f_permutation__out_reg_180_  ( .D(_f_permutation__n5207 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_908), .QN() );
  DFF_X2 _f_permutation__out_reg_179_  ( .D(_f_permutation__n5208 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_909), .QN() );
  DFF_X2 _f_permutation__out_reg_178_  ( .D(_f_permutation__n5209 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_910), .QN() );
  DFF_X2 _f_permutation__out_reg_177_  ( .D(_f_permutation__n5210 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_911), .QN() );
  DFF_X2 _f_permutation__out_reg_176_  ( .D(_f_permutation__n5211 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_912), .QN() );
  DFF_X2 _f_permutation__out_reg_175_  ( .D(_f_permutation__n5212 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_913), .QN() );
  DFF_X2 _f_permutation__out_reg_174_  ( .D(_f_permutation__n5213 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_914), .QN() );
  DFF_X2 _f_permutation__out_reg_173_  ( .D(_f_permutation__n5214 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_915), .QN() );
  DFF_X2 _f_permutation__out_reg_172_  ( .D(_f_permutation__n5215 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_916), .QN() );
  DFF_X2 _f_permutation__out_reg_171_  ( .D(_f_permutation__n5216 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_917), .QN() );
  DFF_X2 _f_permutation__out_reg_170_  ( .D(_f_permutation__n5217 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_918), .QN() );
  DFF_X2 _f_permutation__out_reg_169_  ( .D(_f_permutation__n5218 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_919), .QN() );
  DFF_X2 _f_permutation__out_reg_168_  ( .D(_f_permutation__n5219 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_920), .QN() );
  DFF_X2 _f_permutation__out_reg_167_  ( .D(_f_permutation__n5220 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_921), .QN() );
  DFF_X2 _f_permutation__out_reg_166_  ( .D(_f_permutation__n5221 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_922), .QN() );
  DFF_X2 _f_permutation__out_reg_165_  ( .D(_f_permutation__n5222 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_923), .QN() );
  DFF_X2 _f_permutation__out_reg_164_  ( .D(_f_permutation__n5223 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_924), .QN() );
  DFF_X2 _f_permutation__out_reg_163_  ( .D(_f_permutation__n5224 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_925), .QN() );
  DFF_X2 _f_permutation__out_reg_162_  ( .D(_f_permutation__n5225 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_926), .QN() );
  DFF_X2 _f_permutation__out_reg_161_  ( .D(_f_permutation__n5226 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_927), .QN() );
  DFF_X2 _f_permutation__out_reg_160_  ( .D(_f_permutation__n5227 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_928), .QN() );
  DFF_X2 _f_permutation__out_reg_159_  ( .D(_f_permutation__n5228 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_929), .QN() );
  DFF_X2 _f_permutation__out_reg_158_  ( .D(_f_permutation__n5229 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_930), .QN() );
  DFF_X2 _f_permutation__out_reg_157_  ( .D(_f_permutation__n5230 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_931), .QN() );
  DFF_X2 _f_permutation__out_reg_156_  ( .D(_f_permutation__n5231 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_932), .QN() );
  DFF_X2 _f_permutation__out_reg_155_  ( .D(_f_permutation__n5232 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_933), .QN() );
  DFF_X2 _f_permutation__out_reg_154_  ( .D(_f_permutation__n5233 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_934), .QN() );
  DFF_X2 _f_permutation__out_reg_153_  ( .D(_f_permutation__n5234 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_935), .QN() );
  DFF_X2 _f_permutation__out_reg_152_  ( .D(_f_permutation__n5235 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_936), .QN() );
  DFF_X2 _f_permutation__out_reg_151_  ( .D(_f_permutation__n5236 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_937), .QN() );
  DFF_X2 _f_permutation__out_reg_150_  ( .D(_f_permutation__n5237 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_938), .QN() );
  DFF_X2 _f_permutation__out_reg_149_  ( .D(_f_permutation__n5238 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_939), .QN() );
  DFF_X2 _f_permutation__out_reg_148_  ( .D(_f_permutation__n5239 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_940), .QN() );
  DFF_X2 _f_permutation__out_reg_147_  ( .D(_f_permutation__n5240 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_941), .QN() );
  DFF_X2 _f_permutation__out_reg_146_  ( .D(_f_permutation__n5241 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_942), .QN() );
  DFF_X2 _f_permutation__out_reg_145_  ( .D(_f_permutation__n5242 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_943), .QN() );
  DFF_X2 _f_permutation__out_reg_144_  ( .D(_f_permutation__n5243 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_944), .QN() );
  DFF_X2 _f_permutation__out_reg_143_  ( .D(_f_permutation__n5244 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_945), .QN() );
  DFF_X2 _f_permutation__out_reg_142_  ( .D(_f_permutation__n5245 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_946), .QN() );
  DFF_X2 _f_permutation__out_reg_141_  ( .D(_f_permutation__n5246 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_947), .QN() );
  DFF_X2 _f_permutation__out_reg_140_  ( .D(_f_permutation__n5247 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_948), .QN() );
  DFF_X2 _f_permutation__out_reg_139_  ( .D(_f_permutation__n5248 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_949), .QN() );
  DFF_X2 _f_permutation__out_reg_138_  ( .D(_f_permutation__n5249 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_950), .QN() );
  DFF_X2 _f_permutation__out_reg_137_  ( .D(_f_permutation__n5250 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_951), .QN() );
  DFF_X2 _f_permutation__out_reg_136_  ( .D(_f_permutation__n5251 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_952), .QN() );
  DFF_X2 _f_permutation__out_reg_135_  ( .D(_f_permutation__n5252 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_953), .QN() );
  DFF_X2 _f_permutation__out_reg_134_  ( .D(_f_permutation__n5253 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_954), .QN() );
  DFF_X2 _f_permutation__out_reg_133_  ( .D(_f_permutation__n5254 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_955), .QN() );
  DFF_X2 _f_permutation__out_reg_132_  ( .D(_f_permutation__n5255 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_956), .QN() );
  DFF_X2 _f_permutation__out_reg_131_  ( .D(_f_permutation__n5256 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_957), .QN() );
  DFF_X2 _f_permutation__out_reg_130_  ( .D(_f_permutation__n5257 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_958), .QN() );
  DFF_X2 _f_permutation__out_reg_129_  ( .D(_f_permutation__n5258 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_959), .QN() );
  DFF_X2 _f_permutation__out_reg_128_  ( .D(_f_permutation__n5259 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_960), .QN() );
  DFF_X2 _f_permutation__out_reg_127_  ( .D(_f_permutation__n5260 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_961), .QN() );
  DFF_X2 _f_permutation__out_reg_126_  ( .D(_f_permutation__n5261 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_962), .QN() );
  DFF_X2 _f_permutation__out_reg_125_  ( .D(_f_permutation__n5262 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_963), .QN() );
  DFF_X2 _f_permutation__out_reg_124_  ( .D(_f_permutation__n5263 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_964), .QN() );
  DFF_X2 _f_permutation__out_reg_123_  ( .D(_f_permutation__n5264 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_965), .QN() );
  DFF_X2 _f_permutation__out_reg_122_  ( .D(_f_permutation__n5265 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_966), .QN() );
  DFF_X2 _f_permutation__out_reg_121_  ( .D(_f_permutation__n5266 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_967), .QN() );
  DFF_X2 _f_permutation__out_reg_120_  ( .D(_f_permutation__n5267 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_968), .QN() );
  DFF_X2 _f_permutation__out_reg_119_  ( .D(_f_permutation__n5268 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_969), .QN() );
  DFF_X2 _f_permutation__out_reg_118_  ( .D(_f_permutation__n5269 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_970), .QN() );
  DFF_X2 _f_permutation__out_reg_117_  ( .D(_f_permutation__n5270 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_971), .QN() );
  DFF_X2 _f_permutation__out_reg_116_  ( .D(_f_permutation__n5271 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_972), .QN() );
  DFF_X2 _f_permutation__out_reg_115_  ( .D(_f_permutation__n5272 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_973), .QN() );
  DFF_X2 _f_permutation__out_reg_114_  ( .D(_f_permutation__n5273 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_974), .QN() );
  DFF_X2 _f_permutation__out_reg_113_  ( .D(_f_permutation__n5274 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_975), .QN() );
  DFF_X2 _f_permutation__out_reg_112_  ( .D(_f_permutation__n5275 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_976), .QN() );
  DFF_X2 _f_permutation__out_reg_111_  ( .D(_f_permutation__n5276 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_977), .QN() );
  DFF_X2 _f_permutation__out_reg_110_  ( .D(_f_permutation__n5277 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_978), .QN() );
  DFF_X2 _f_permutation__out_reg_109_  ( .D(_f_permutation__n5278 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_979), .QN() );
  DFF_X2 _f_permutation__out_reg_108_  ( .D(_f_permutation__n5279 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_980), .QN() );
  DFF_X2 _f_permutation__out_reg_107_  ( .D(_f_permutation__n5280 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_981), .QN() );
  DFF_X2 _f_permutation__out_reg_106_  ( .D(_f_permutation__n5281 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_982), .QN() );
  DFF_X2 _f_permutation__out_reg_105_  ( .D(_f_permutation__n5282 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_983), .QN() );
  DFF_X2 _f_permutation__out_reg_104_  ( .D(_f_permutation__n5283 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_984), .QN() );
  DFF_X2 _f_permutation__out_reg_103_  ( .D(_f_permutation__n5284 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_985), .QN() );
  DFF_X2 _f_permutation__out_reg_102_  ( .D(_f_permutation__n5285 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_986), .QN() );
  DFF_X2 _f_permutation__out_reg_101_  ( .D(_f_permutation__n5286 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_987), .QN() );
  DFF_X2 _f_permutation__out_reg_100_  ( .D(_f_permutation__n5287 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_988), .QN() );
  DFF_X2 _f_permutation__out_reg_99_  ( .D(_f_permutation__n5288 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_989), .QN() );
  DFF_X2 _f_permutation__out_reg_98_  ( .D(_f_permutation__n5289 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_990), .QN() );
  DFF_X2 _f_permutation__out_reg_97_  ( .D(_f_permutation__n5290 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_991), .QN() );
  DFF_X2 _f_permutation__out_reg_96_  ( .D(_f_permutation__n5291 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_992), .QN() );
  DFF_X2 _f_permutation__out_reg_95_  ( .D(_f_permutation__n5292 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_993), .QN() );
  DFF_X2 _f_permutation__out_reg_94_  ( .D(_f_permutation__n5293 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_994), .QN() );
  DFF_X2 _f_permutation__out_reg_93_  ( .D(_f_permutation__n5294 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_995), .QN() );
  DFF_X2 _f_permutation__out_reg_92_  ( .D(_f_permutation__n5295 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_996), .QN() );
  DFF_X2 _f_permutation__out_reg_91_  ( .D(_f_permutation__n5296 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_997), .QN() );
  DFF_X2 _f_permutation__out_reg_90_  ( .D(_f_permutation__n5297 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_998), .QN() );
  DFF_X2 _f_permutation__out_reg_89_  ( .D(_f_permutation__n5298 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_999), .QN() );
  DFF_X2 _f_permutation__out_reg_88_  ( .D(_f_permutation__n5299 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1000), .QN() );
  DFF_X2 _f_permutation__out_reg_87_  ( .D(_f_permutation__n5300 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1001), .QN() );
  DFF_X2 _f_permutation__out_reg_86_  ( .D(_f_permutation__n5301 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1002), .QN() );
  DFF_X2 _f_permutation__out_reg_85_  ( .D(_f_permutation__n5302 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1003), .QN() );
  DFF_X2 _f_permutation__out_reg_84_  ( .D(_f_permutation__n5303 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1004), .QN() );
  DFF_X2 _f_permutation__out_reg_83_  ( .D(_f_permutation__n5304 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1005), .QN() );
  DFF_X2 _f_permutation__out_reg_82_  ( .D(_f_permutation__n5305 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1006), .QN() );
  DFF_X2 _f_permutation__out_reg_81_  ( .D(_f_permutation__n5306 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1007), .QN() );
  DFF_X2 _f_permutation__out_reg_80_  ( .D(_f_permutation__n5307 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1008), .QN() );
  DFF_X2 _f_permutation__out_reg_79_  ( .D(_f_permutation__n5308 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1009), .QN() );
  DFF_X2 _f_permutation__out_reg_78_  ( .D(_f_permutation__n5309 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1010), .QN() );
  DFF_X2 _f_permutation__out_reg_77_  ( .D(_f_permutation__n5310 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1011), .QN() );
  DFF_X2 _f_permutation__out_reg_76_  ( .D(_f_permutation__n5311 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1012), .QN() );
  DFF_X2 _f_permutation__out_reg_75_  ( .D(_f_permutation__n5312 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1013), .QN() );
  DFF_X2 _f_permutation__out_reg_74_  ( .D(_f_permutation__n5313 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1014), .QN() );
  DFF_X2 _f_permutation__out_reg_73_  ( .D(_f_permutation__n5314 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1015), .QN() );
  DFF_X2 _f_permutation__out_reg_72_  ( .D(_f_permutation__n5315 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1016), .QN() );
  DFF_X2 _f_permutation__out_reg_71_  ( .D(_f_permutation__n5316 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1017), .QN() );
  DFF_X2 _f_permutation__out_reg_70_  ( .D(_f_permutation__n5317 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1018), .QN() );
  DFF_X2 _f_permutation__out_reg_69_  ( .D(_f_permutation__n5318 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1019), .QN() );
  DFF_X2 _f_permutation__out_reg_68_  ( .D(_f_permutation__n5319 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1020), .QN() );
  DFF_X2 _f_permutation__out_reg_67_  ( .D(_f_permutation__n5320 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1021), .QN() );
  DFF_X2 _f_permutation__out_reg_66_  ( .D(_f_permutation__n5321 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1022), .QN() );
  DFF_X2 _f_permutation__out_reg_65_  ( .D(_f_permutation__n5322 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1023), .QN() );
  DFF_X2 _f_permutation__out_reg_64_  ( .D(_f_permutation__n5323 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1024), .QN() );
  DFF_X2 _f_permutation__out_reg_63_  ( .D(_f_permutation__n5324 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1025), .QN() );
  DFF_X2 _f_permutation__out_reg_62_  ( .D(_f_permutation__n5325 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1026), .QN() );
  DFF_X2 _f_permutation__out_reg_61_  ( .D(_f_permutation__n5326 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1027), .QN() );
  DFF_X2 _f_permutation__out_reg_60_  ( .D(_f_permutation__n5327 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1028), .QN() );
  DFF_X2 _f_permutation__out_reg_59_  ( .D(_f_permutation__n5328 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1029), .QN() );
  DFF_X2 _f_permutation__out_reg_58_  ( .D(_f_permutation__n5329 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1030), .QN() );
  DFF_X2 _f_permutation__out_reg_57_  ( .D(_f_permutation__n5330 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1031), .QN() );
  DFF_X2 _f_permutation__out_reg_56_  ( .D(_f_permutation__n5331 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1032), .QN() );
  DFF_X2 _f_permutation__out_reg_55_  ( .D(_f_permutation__n5332 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1033), .QN() );
  DFF_X2 _f_permutation__out_reg_54_  ( .D(_f_permutation__n5333 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1034), .QN() );
  DFF_X2 _f_permutation__out_reg_53_  ( .D(_f_permutation__n5334 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1035), .QN() );
  DFF_X2 _f_permutation__out_reg_52_  ( .D(_f_permutation__n5335 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1036), .QN() );
  DFF_X2 _f_permutation__out_reg_51_  ( .D(_f_permutation__n5336 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1037), .QN() );
  DFF_X2 _f_permutation__out_reg_50_  ( .D(_f_permutation__n5337 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1038), .QN() );
  DFF_X2 _f_permutation__out_reg_49_  ( .D(_f_permutation__n5338 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1039), .QN() );
  DFF_X2 _f_permutation__out_reg_48_  ( .D(_f_permutation__n5339 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1040), .QN() );
  DFF_X2 _f_permutation__out_reg_47_  ( .D(_f_permutation__n5340 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1041), .QN() );
  DFF_X2 _f_permutation__out_reg_46_  ( .D(_f_permutation__n5341 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1042), .QN() );
  DFF_X2 _f_permutation__out_reg_45_  ( .D(_f_permutation__n5342 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1043), .QN() );
  DFF_X2 _f_permutation__out_reg_44_  ( .D(_f_permutation__n5343 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1044), .QN() );
  DFF_X2 _f_permutation__out_reg_43_  ( .D(_f_permutation__n5344 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1045), .QN() );
  DFF_X2 _f_permutation__out_reg_42_  ( .D(_f_permutation__n5345 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1046), .QN() );
  DFF_X2 _f_permutation__out_reg_41_  ( .D(_f_permutation__n5346 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1047), .QN() );
  DFF_X2 _f_permutation__out_reg_40_  ( .D(_f_permutation__n5347 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1048), .QN() );
  DFF_X2 _f_permutation__out_reg_39_  ( .D(_f_permutation__n5348 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1049), .QN() );
  DFF_X2 _f_permutation__out_reg_38_  ( .D(_f_permutation__n5349 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1050), .QN() );
  DFF_X2 _f_permutation__out_reg_37_  ( .D(_f_permutation__n5350 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1051), .QN() );
  DFF_X2 _f_permutation__out_reg_36_  ( .D(_f_permutation__n5351 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1052), .QN() );
  DFF_X2 _f_permutation__out_reg_35_  ( .D(_f_permutation__n5352 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1053), .QN() );
  DFF_X2 _f_permutation__out_reg_34_  ( .D(_f_permutation__n5353 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1054), .QN() );
  DFF_X2 _f_permutation__out_reg_33_  ( .D(_f_permutation__n5354 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1055), .QN() );
  DFF_X2 _f_permutation__out_reg_32_  ( .D(_f_permutation__n5355 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1056), .QN() );
  DFF_X2 _f_permutation__out_reg_31_  ( .D(_f_permutation__n5356 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1057), .QN() );
  DFF_X2 _f_permutation__out_reg_30_  ( .D(_f_permutation__n5357 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1058), .QN() );
  DFF_X2 _f_permutation__out_reg_29_  ( .D(_f_permutation__n5358 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1059), .QN() );
  DFF_X2 _f_permutation__out_reg_28_  ( .D(_f_permutation__n5359 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1060), .QN() );
  DFF_X2 _f_permutation__out_reg_27_  ( .D(_f_permutation__n5360 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1061), .QN() );
  DFF_X2 _f_permutation__out_reg_26_  ( .D(_f_permutation__n5361 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1062), .QN() );
  DFF_X2 _f_permutation__out_reg_25_  ( .D(_f_permutation__n5362 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1063), .QN() );
  DFF_X2 _f_permutation__out_reg_24_  ( .D(_f_permutation__n5363 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1064), .QN() );
  DFF_X2 _f_permutation__out_reg_23_  ( .D(_f_permutation__n5364 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1065), .QN() );
  DFF_X2 _f_permutation__out_reg_22_  ( .D(_f_permutation__n5365 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1066), .QN() );
  DFF_X2 _f_permutation__out_reg_21_  ( .D(_f_permutation__n5366 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1067), .QN() );
  DFF_X2 _f_permutation__out_reg_20_  ( .D(_f_permutation__n5367 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1068), .QN() );
  DFF_X2 _f_permutation__out_reg_19_  ( .D(_f_permutation__n5368 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1069), .QN() );
  DFF_X2 _f_permutation__out_reg_18_  ( .D(_f_permutation__n5369 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1070), .QN() );
  DFF_X2 _f_permutation__out_reg_17_  ( .D(_f_permutation__n5370 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1071), .QN() );
  DFF_X2 _f_permutation__out_reg_16_  ( .D(_f_permutation__n5371 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1072), .QN() );
  DFF_X2 _f_permutation__out_reg_15_  ( .D(_f_permutation__n5372 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1073), .QN() );
  DFF_X2 _f_permutation__out_reg_14_  ( .D(_f_permutation__n5373 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1074), .QN() );
  DFF_X2 _f_permutation__out_reg_13_  ( .D(_f_permutation__n5374 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1075), .QN() );
  DFF_X2 _f_permutation__out_reg_12_  ( .D(_f_permutation__n5375 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1076), .QN() );
  DFF_X2 _f_permutation__out_reg_11_  ( .D(_f_permutation__n5376 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1077), .QN() );
  DFF_X2 _f_permutation__out_reg_10_  ( .D(_f_permutation__n5377 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1078), .QN() );
  DFF_X2 _f_permutation__out_reg_9_  ( .D(_f_permutation__n5378 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1079), .QN() );
  DFF_X2 _f_permutation__out_reg_8_  ( .D(_f_permutation__n5379 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1080), .QN() );
  DFF_X2 _f_permutation__out_reg_7_  ( .D(_f_permutation__n5380 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1081), .QN() );
  DFF_X2 _f_permutation__out_reg_6_  ( .D(_f_permutation__n5381 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1082), .QN() );
  DFF_X2 _f_permutation__out_reg_5_  ( .D(_f_permutation__n5382 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1083), .QN() );
  DFF_X2 _f_permutation__out_reg_4_  ( .D(_f_permutation__n5383 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1084), .QN() );
  DFF_X2 _f_permutation__out_reg_3_  ( .D(_f_permutation__n5384 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1085), .QN() );
  DFF_X2 _f_permutation__out_reg_2_  ( .D(_f_permutation__n5385 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1086), .QN() );
  DFF_X2 _f_permutation__out_reg_1_  ( .D(_f_permutation__n5386 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1087), .QN() );
  DFF_X2 _f_permutation__out_reg_0_  ( .D(_f_permutation__n5387 ), .CK(clk), 
        .Q(SYNOPSYS_UNCONNECTED_1088), .QN() );
  NOR4_X2 _f_permutation__rconst__U145  ( .A1(_f_permutation__i[7] ), .A2(
        _f_permutation__i[3] ), .A3(_f_permutation__i[1] ), .A4(
        _f_permutation__i[18] ), .ZN(_f_permutation__rconst__n21 ) );
  NOR4_X2 _f_permutation__rconst__U144  ( .A1(_f_permutation__i[17] ), .A2(
        _f_permutation__i[12] ), .A3(_f_permutation__i[11] ), .A4(
        _f_permutation__i[10] ), .ZN(_f_permutation__rconst__n20 ) );
  NOR4_X2 _f_permutation__rconst__U143  ( .A1(_f_permutation__i[6] ), .A2(
        _f_permutation__i[1] ), .A3(_f_permutation__i[20] ), .A4(
        _f_permutation__i[15] ), .ZN(_f_permutation__rconst__n19 ) );
  NOR3_X2 _f_permutation__rconst__U142  ( .A1(_f_permutation__i[19] ), .A2(
        _f_permutation__i[5] ), .A3(_f_permutation__i[3] ), .ZN(
        _f_permutation__rconst__n23 ) );
  NOR3_X2 _f_permutation__rconst__U141  ( .A1(_f_permutation__i[4] ), .A2(
        _f_permutation__i[21] ), .A3(_f_permutation__i[9] ), .ZN(
        _f_permutation__rconst__n13 ) );
  NOR4_X2 _f_permutation__rconst__U140  ( .A1(_f_permutation__i[22] ), .A2(
        _f_permutation__i[19] ), .A3(_f_permutation__i[5] ), .A4(
        _f_permutation__i[2] ), .ZN(_f_permutation__rconst__n14 ) );
  NOR3_X2 _f_permutation__rconst__U139  ( .A1(f_ack), .A2(
        _f_permutation__i[6] ), .A3(_f_permutation__i[14] ), .ZN(
        _f_permutation__rconst__n22 ) );
  NAND3_X2 _f_permutation__rconst__U138  ( .A1(_f_permutation__rconst__n13 ), 
        .A2(_f_permutation__rconst__n10 ), .A3(_f_permutation__rconst__n22 ), 
        .ZN(_f_permutation__rc[0]) );
  NOR3_X2 _f_permutation__rconst__U137  ( .A1(_f_permutation__i[22] ), .A2(
        _f_permutation__i[8] ), .A3(_f_permutation__i[6] ), .ZN(
        _f_permutation__rconst__n17 ) );
  NOR4_X2 _f_permutation__rconst__U136  ( .A1(_f_permutation__i[8] ), .A2(
        _f_permutation__i[7] ), .A3(_f_permutation__i[1] ), .A4(
        _f_permutation__i[20] ), .ZN(_f_permutation__rconst__n11 ) );
  NOR3_X2 _f_permutation__rconst__U135  ( .A1(_f_permutation__i[17] ), .A2(
        _f_permutation__i[3] ), .A3(_f_permutation__i[0] ), .ZN(
        _f_permutation__rconst__n18 ) );
  NOR3_X2 _f_permutation__rconst__U134  ( .A1(_f_permutation__i[10] ), .A2(
        _f_permutation__i[18] ), .A3(_f_permutation__i[11] ), .ZN(
        _f_permutation__rconst__n15 ) );
  NAND3_X2 _f_permutation__rconst__U133  ( .A1(_f_permutation__rconst__n13 ), 
        .A2(_f_permutation__rconst__n14 ), .A3(_f_permutation__rconst__n15 ), 
        .ZN(_f_permutation__rc[31]) );
  INV_X4 _f_permutation__rconst__U131  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[62] ) );
  INV_X4 _f_permutation__rconst__U129  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[61] ) );
  INV_X4 _f_permutation__rconst__U127  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[60] ) );
  INV_X4 _f_permutation__rconst__U125  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[59] ) );
  INV_X4 _f_permutation__rconst__U123  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[58] ) );
  INV_X4 _f_permutation__rconst__U121  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[57] ) );
  INV_X4 _f_permutation__rconst__U119  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[56] ) );
  INV_X4 _f_permutation__rconst__U117  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[55] ) );
  INV_X4 _f_permutation__rconst__U115  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[54] ) );
  INV_X4 _f_permutation__rconst__U113  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[53] ) );
  INV_X4 _f_permutation__rconst__U111  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[52] ) );
  INV_X4 _f_permutation__rconst__U109  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[51] ) );
  INV_X4 _f_permutation__rconst__U107  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[50] ) );
  INV_X4 _f_permutation__rconst__U105  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[49] ) );
  INV_X4 _f_permutation__rconst__U103  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[48] ) );
  INV_X4 _f_permutation__rconst__U101  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[47] ) );
  INV_X4 _f_permutation__rconst__U99  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[46] ) );
  INV_X4 _f_permutation__rconst__U97  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[45] ) );
  INV_X4 _f_permutation__rconst__U95  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[44] ) );
  INV_X4 _f_permutation__rconst__U93  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[43] ) );
  INV_X4 _f_permutation__rconst__U91  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[42] ) );
  INV_X4 _f_permutation__rconst__U89  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[41] ) );
  INV_X4 _f_permutation__rconst__U87  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[40] ) );
  INV_X4 _f_permutation__rconst__U85  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[39] ) );
  INV_X4 _f_permutation__rconst__U83  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[38] ) );
  INV_X4 _f_permutation__rconst__U81  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[37] ) );
  INV_X4 _f_permutation__rconst__U79  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[36] ) );
  INV_X4 _f_permutation__rconst__U77  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[35] ) );
  INV_X4 _f_permutation__rconst__U75  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[34] ) );
  INV_X4 _f_permutation__rconst__U73  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[33] ) );
  INV_X4 _f_permutation__rconst__U71  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[32] ) );
  INV_X4 _f_permutation__rconst__U69  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[30] ) );
  INV_X4 _f_permutation__rconst__U67  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[29] ) );
  INV_X4 _f_permutation__rconst__U65  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[28] ) );
  INV_X4 _f_permutation__rconst__U63  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[27] ) );
  INV_X4 _f_permutation__rconst__U61  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[26] ) );
  INV_X4 _f_permutation__rconst__U59  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[25] ) );
  INV_X4 _f_permutation__rconst__U57  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[24] ) );
  INV_X4 _f_permutation__rconst__U55  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[23] ) );
  INV_X4 _f_permutation__rconst__U53  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[22] ) );
  INV_X4 _f_permutation__rconst__U51  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[21] ) );
  INV_X4 _f_permutation__rconst__U49  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[20] ) );
  INV_X4 _f_permutation__rconst__U47  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[19] ) );
  INV_X4 _f_permutation__rconst__U45  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[18] ) );
  INV_X4 _f_permutation__rconst__U43  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[17] ) );
  INV_X4 _f_permutation__rconst__U41  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[16] ) );
  INV_X4 _f_permutation__rconst__U39  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[14] ) );
  INV_X4 _f_permutation__rconst__U37  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[13] ) );
  INV_X4 _f_permutation__rconst__U35  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[12] ) );
  INV_X4 _f_permutation__rconst__U33  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[11] ) );
  INV_X4 _f_permutation__rconst__U22  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[10] ) );
  INV_X4 _f_permutation__rconst__U19  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[9] ) );
  INV_X4 _f_permutation__rconst__U17  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[8] ) );
  INV_X4 _f_permutation__rconst__U13  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[6] ) );
  INV_X4 _f_permutation__rconst__U10  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[5] ) );
  INV_X4 _f_permutation__rconst__U6  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[4] ) );
  INV_X4 _f_permutation__rconst__U3  ( .A(1'b1), .ZN(
        _f_permutation__rconst__rc[2] ) );
  INV_X4 _f_permutation__rconst__U31  ( .A(_f_permutation__i[0] ), .ZN(
        _f_permutation__rconst__n9 ) );
  INV_X4 _f_permutation__rconst__U30  ( .A(_f_permutation__i[9] ), .ZN(
        _f_permutation__rconst__n8 ) );
  INV_X4 _f_permutation__rconst__U29  ( .A(_f_permutation__i[11] ), .ZN(
        _f_permutation__rconst__n7 ) );
  INV_X4 _f_permutation__rconst__U28  ( .A(_f_permutation__i[12] ), .ZN(
        _f_permutation__rconst__n6 ) );
  INV_X4 _f_permutation__rconst__U27  ( .A(_f_permutation__i[13] ), .ZN(
        _f_permutation__rconst__n5 ) );
  INV_X4 _f_permutation__rconst__U26  ( .A(_f_permutation__i[14] ), .ZN(
        _f_permutation__rconst__n4 ) );
  INV_X4 _f_permutation__rconst__U25  ( .A(_f_permutation__i[15] ), .ZN(
        _f_permutation__rconst__n3 ) );
  INV_X4 _f_permutation__rconst__U24  ( .A(_f_permutation__i[16] ), .ZN(
        _f_permutation__rconst__n2 ) );
  INV_X4 _f_permutation__rconst__U23  ( .A(_f_permutation__i[18] ), .ZN(
        _f_permutation__rconst__n1 ) );
  AND4_X2 _f_permutation__rconst__U20  ( .A1(_f_permutation__rconst__n6 ), 
        .A2(_f_permutation__rconst__n5 ), .A3(_f_permutation__rconst__n7 ), 
        .A4(_f_permutation__rconst__n23 ), .ZN(_f_permutation__rconst__n10 )
         );
  AND2_X2 _f_permutation__rconst__U15  ( .A1(_f_permutation__rconst__n20 ), 
        .A2(_f_permutation__rconst__n21 ), .ZN(_f_permutation__rconst__n16 )
         );
  NAND4_X2 _f_permutation__rconst__U14  ( .A1(_f_permutation__rconst__n16 ), 
        .A2(_f_permutation__rconst__n4 ), .A3(_f_permutation__rconst__n3 ), 
        .A4(_f_permutation__rconst__n9 ), .ZN(_f_permutation__rc[1]) );
  AND4_X2 _f_permutation__rconst__U11  ( .A1(_f_permutation__rconst__n5 ), 
        .A2(_f_permutation__rconst__n4 ), .A3(_f_permutation__rconst__n14 ), 
        .A4(_f_permutation__rconst__n19 ), .ZN(_f_permutation__rconst__n12 )
         );
  NAND4_X2 _f_permutation__rconst__U9  ( .A1(_f_permutation__rconst__n8 ), 
        .A2(_f_permutation__rconst__n7 ), .A3(_f_permutation__rconst__n12 ), 
        .A4(_f_permutation__rconst__n18 ), .ZN(_f_permutation__rc[15]) );
  NAND4_X2 _f_permutation__rconst__U7  ( .A1(_f_permutation__rconst__n8 ), 
        .A2(_f_permutation__rconst__n5 ), .A3(_f_permutation__rconst__n16 ), 
        .A4(_f_permutation__rconst__n17 ), .ZN(_f_permutation__rc[3]) );
  NAND4_X2 _f_permutation__rconst__U4  ( .A1(_f_permutation__rconst__n12 ), 
        .A2(_f_permutation__rconst__n6 ), .A3(_f_permutation__rconst__n2 ), 
        .A4(_f_permutation__rconst__n1 ), .ZN(_f_permutation__rc[63]) );
  NAND4_X2 _f_permutation__rconst__U2  ( .A1(_f_permutation__rconst__n2 ), 
        .A2(_f_permutation__rconst__n9 ), .A3(_f_permutation__rconst__n10 ), 
        .A4(_f_permutation__rconst__n11 ), .ZN(_f_permutation__rc[7]) );
  NOR2_X2 _f_permutation__round__U1600  ( .A1(_f_permutation__round__c[404] ), 
        .A2(_f_permutation__round__n660 ), .ZN(_f_permutation__round__N2687 )
         );
  NOR2_X2 _f_permutation__round__U1599  ( .A1(_f_permutation__round__c[405] ), 
        .A2(_f_permutation__round__n655 ), .ZN(_f_permutation__round__N2685 )
         );
  NOR2_X2 _f_permutation__round__U1598  ( .A1(_f_permutation__round__c[407] ), 
        .A2(_f_permutation__round__n645 ), .ZN(_f_permutation__round__N2681 )
         );
  NOR2_X2 _f_permutation__round__U1597  ( .A1(_f_permutation__round__c[411] ), 
        .A2(_f_permutation__round__n625 ), .ZN(_f_permutation__round__N2673 )
         );
  NOR2_X2 _f_permutation__round__U1596  ( .A1(_f_permutation__round__c[419] ), 
        .A2(_f_permutation__round__n585 ), .ZN(_f_permutation__round__N2657 )
         );
  NOR2_X2 _f_permutation__round__U1595  ( .A1(_f_permutation__round__c[435] ), 
        .A2(_f_permutation__round__n505 ), .ZN(_f_permutation__round__N2625 )
         );
  NOR2_X2 _f_permutation__round__U1594  ( .A1(_f_permutation__round__c[403] ), 
        .A2(_f_permutation__round__n665 ), .ZN(_f_permutation__round__N2561 )
         );
  NOR2_X2 _f_permutation__round__U1593  ( .A1(_f_permutation__round__c[638] ), 
        .A2(_f_permutation__round__n754 ), .ZN(_f_permutation__round__N5631 )
         );
  NOR2_X2 _f_permutation__round__U1592  ( .A1(_f_permutation__round__c[639] ), 
        .A2(_f_permutation__round__n749 ), .ZN(_f_permutation__round__N5629 )
         );
  NOR2_X2 _f_permutation__round__U1591  ( .A1(_f_permutation__round__c[576] ), 
        .A2(_f_permutation__round__n744 ), .ZN(_f_permutation__round__N5627 )
         );
  NOR2_X2 _f_permutation__round__U1590  ( .A1(_f_permutation__round__c[577] ), 
        .A2(_f_permutation__round__n739 ), .ZN(_f_permutation__round__N5625 )
         );
  NOR2_X2 _f_permutation__round__U1589  ( .A1(_f_permutation__round__c[578] ), 
        .A2(_f_permutation__round__n734 ), .ZN(_f_permutation__round__N5623 )
         );
  NOR2_X2 _f_permutation__round__U1588  ( .A1(_f_permutation__round__c[579] ), 
        .A2(_f_permutation__round__n729 ), .ZN(_f_permutation__round__N5621 )
         );
  NOR2_X2 _f_permutation__round__U1587  ( .A1(_f_permutation__round__c[580] ), 
        .A2(_f_permutation__round__n724 ), .ZN(_f_permutation__round__N5619 )
         );
  NOR2_X2 _f_permutation__round__U1586  ( .A1(_f_permutation__round__c[581] ), 
        .A2(_f_permutation__round__n719 ), .ZN(_f_permutation__round__N5617 )
         );
  NOR2_X2 _f_permutation__round__U1585  ( .A1(_f_permutation__round__c[582] ), 
        .A2(_f_permutation__round__n714 ), .ZN(_f_permutation__round__N5615 )
         );
  NOR2_X2 _f_permutation__round__U1584  ( .A1(_f_permutation__round__c[583] ), 
        .A2(_f_permutation__round__n709 ), .ZN(_f_permutation__round__N5613 )
         );
  NOR2_X2 _f_permutation__round__U1583  ( .A1(_f_permutation__round__c[584] ), 
        .A2(_f_permutation__round__n704 ), .ZN(_f_permutation__round__N5611 )
         );
  NOR2_X2 _f_permutation__round__U1582  ( .A1(_f_permutation__round__c[585] ), 
        .A2(_f_permutation__round__n699 ), .ZN(_f_permutation__round__N5609 )
         );
  NOR2_X2 _f_permutation__round__U1581  ( .A1(_f_permutation__round__c[586] ), 
        .A2(_f_permutation__round__n694 ), .ZN(_f_permutation__round__N5607 )
         );
  NOR2_X2 _f_permutation__round__U1580  ( .A1(_f_permutation__round__c[587] ), 
        .A2(_f_permutation__round__n689 ), .ZN(_f_permutation__round__N5605 )
         );
  NOR2_X2 _f_permutation__round__U1579  ( .A1(_f_permutation__round__c[588] ), 
        .A2(_f_permutation__round__n684 ), .ZN(_f_permutation__round__N5603 )
         );
  NOR2_X2 _f_permutation__round__U1578  ( .A1(_f_permutation__round__c[589] ), 
        .A2(_f_permutation__round__n679 ), .ZN(_f_permutation__round__N5601 )
         );
  NOR2_X2 _f_permutation__round__U1577  ( .A1(_f_permutation__round__c[590] ), 
        .A2(_f_permutation__round__n674 ), .ZN(_f_permutation__round__N5599 )
         );
  NOR2_X2 _f_permutation__round__U1576  ( .A1(_f_permutation__round__c[591] ), 
        .A2(_f_permutation__round__n669 ), .ZN(_f_permutation__round__N5597 )
         );
  NOR2_X2 _f_permutation__round__U1575  ( .A1(_f_permutation__round__c[592] ), 
        .A2(_f_permutation__round__n664 ), .ZN(_f_permutation__round__N5595 )
         );
  NOR2_X2 _f_permutation__round__U1574  ( .A1(_f_permutation__round__c[593] ), 
        .A2(_f_permutation__round__n659 ), .ZN(_f_permutation__round__N5593 )
         );
  NOR2_X2 _f_permutation__round__U1573  ( .A1(_f_permutation__round__c[594] ), 
        .A2(_f_permutation__round__n654 ), .ZN(_f_permutation__round__N5591 )
         );
  NOR2_X2 _f_permutation__round__U1572  ( .A1(_f_permutation__round__c[595] ), 
        .A2(_f_permutation__round__n649 ), .ZN(_f_permutation__round__N5589 )
         );
  NOR2_X2 _f_permutation__round__U1571  ( .A1(_f_permutation__round__c[596] ), 
        .A2(_f_permutation__round__n644 ), .ZN(_f_permutation__round__N5587 )
         );
  NOR2_X2 _f_permutation__round__U1570  ( .A1(_f_permutation__round__c[597] ), 
        .A2(_f_permutation__round__n639 ), .ZN(_f_permutation__round__N5585 )
         );
  NOR2_X2 _f_permutation__round__U1569  ( .A1(_f_permutation__round__c[598] ), 
        .A2(_f_permutation__round__n634 ), .ZN(_f_permutation__round__N5583 )
         );
  NOR2_X2 _f_permutation__round__U1568  ( .A1(_f_permutation__round__c[599] ), 
        .A2(_f_permutation__round__n629 ), .ZN(_f_permutation__round__N5581 )
         );
  NOR2_X2 _f_permutation__round__U1567  ( .A1(_f_permutation__round__c[600] ), 
        .A2(_f_permutation__round__n624 ), .ZN(_f_permutation__round__N5579 )
         );
  NOR2_X2 _f_permutation__round__U1566  ( .A1(_f_permutation__round__c[601] ), 
        .A2(_f_permutation__round__n619 ), .ZN(_f_permutation__round__N5577 )
         );
  NOR2_X2 _f_permutation__round__U1565  ( .A1(_f_permutation__round__c[602] ), 
        .A2(_f_permutation__round__n614 ), .ZN(_f_permutation__round__N5575 )
         );
  NOR2_X2 _f_permutation__round__U1564  ( .A1(_f_permutation__round__c[603] ), 
        .A2(_f_permutation__round__n609 ), .ZN(_f_permutation__round__N5573 )
         );
  NOR2_X2 _f_permutation__round__U1563  ( .A1(_f_permutation__round__c[604] ), 
        .A2(_f_permutation__round__n604 ), .ZN(_f_permutation__round__N5571 )
         );
  NOR2_X2 _f_permutation__round__U1562  ( .A1(_f_permutation__round__c[605] ), 
        .A2(_f_permutation__round__n599 ), .ZN(_f_permutation__round__N5569 )
         );
  NOR2_X2 _f_permutation__round__U1561  ( .A1(_f_permutation__round__c[606] ), 
        .A2(_f_permutation__round__n594 ), .ZN(_f_permutation__round__N5567 )
         );
  NOR2_X2 _f_permutation__round__U1560  ( .A1(_f_permutation__round__c[607] ), 
        .A2(_f_permutation__round__n589 ), .ZN(_f_permutation__round__N5565 )
         );
  NOR2_X2 _f_permutation__round__U1559  ( .A1(_f_permutation__round__c[608] ), 
        .A2(_f_permutation__round__n584 ), .ZN(_f_permutation__round__N5563 )
         );
  NOR2_X2 _f_permutation__round__U1558  ( .A1(_f_permutation__round__c[609] ), 
        .A2(_f_permutation__round__n579 ), .ZN(_f_permutation__round__N5561 )
         );
  NOR2_X2 _f_permutation__round__U1557  ( .A1(_f_permutation__round__c[610] ), 
        .A2(_f_permutation__round__n574 ), .ZN(_f_permutation__round__N5559 )
         );
  NOR2_X2 _f_permutation__round__U1556  ( .A1(_f_permutation__round__c[611] ), 
        .A2(_f_permutation__round__n569 ), .ZN(_f_permutation__round__N5557 )
         );
  NOR2_X2 _f_permutation__round__U1555  ( .A1(_f_permutation__round__c[612] ), 
        .A2(_f_permutation__round__n564 ), .ZN(_f_permutation__round__N5555 )
         );
  NOR2_X2 _f_permutation__round__U1554  ( .A1(_f_permutation__round__c[613] ), 
        .A2(_f_permutation__round__n559 ), .ZN(_f_permutation__round__N5553 )
         );
  NOR2_X2 _f_permutation__round__U1553  ( .A1(_f_permutation__round__c[614] ), 
        .A2(_f_permutation__round__n554 ), .ZN(_f_permutation__round__N5551 )
         );
  NOR2_X2 _f_permutation__round__U1552  ( .A1(_f_permutation__round__c[615] ), 
        .A2(_f_permutation__round__n549 ), .ZN(_f_permutation__round__N5549 )
         );
  NOR2_X2 _f_permutation__round__U1551  ( .A1(_f_permutation__round__c[616] ), 
        .A2(_f_permutation__round__n544 ), .ZN(_f_permutation__round__N5547 )
         );
  NOR2_X2 _f_permutation__round__U1550  ( .A1(_f_permutation__round__c[617] ), 
        .A2(_f_permutation__round__n539 ), .ZN(_f_permutation__round__N5545 )
         );
  NOR2_X2 _f_permutation__round__U1549  ( .A1(_f_permutation__round__c[618] ), 
        .A2(_f_permutation__round__n534 ), .ZN(_f_permutation__round__N5543 )
         );
  NOR2_X2 _f_permutation__round__U1548  ( .A1(_f_permutation__round__c[619] ), 
        .A2(_f_permutation__round__n529 ), .ZN(_f_permutation__round__N5541 )
         );
  NOR2_X2 _f_permutation__round__U1547  ( .A1(_f_permutation__round__c[620] ), 
        .A2(_f_permutation__round__n524 ), .ZN(_f_permutation__round__N5539 )
         );
  NOR2_X2 _f_permutation__round__U1546  ( .A1(_f_permutation__round__c[621] ), 
        .A2(_f_permutation__round__n519 ), .ZN(_f_permutation__round__N5537 )
         );
  NOR2_X2 _f_permutation__round__U1545  ( .A1(_f_permutation__round__c[622] ), 
        .A2(_f_permutation__round__n514 ), .ZN(_f_permutation__round__N5535 )
         );
  NOR2_X2 _f_permutation__round__U1544  ( .A1(_f_permutation__round__c[623] ), 
        .A2(_f_permutation__round__n509 ), .ZN(_f_permutation__round__N5533 )
         );
  NOR2_X2 _f_permutation__round__U1543  ( .A1(_f_permutation__round__c[624] ), 
        .A2(_f_permutation__round__n504 ), .ZN(_f_permutation__round__N5531 )
         );
  NOR2_X2 _f_permutation__round__U1542  ( .A1(_f_permutation__round__c[625] ), 
        .A2(_f_permutation__round__n499 ), .ZN(_f_permutation__round__N5529 )
         );
  NOR2_X2 _f_permutation__round__U1541  ( .A1(_f_permutation__round__c[626] ), 
        .A2(_f_permutation__round__n494 ), .ZN(_f_permutation__round__N5527 )
         );
  NOR2_X2 _f_permutation__round__U1540  ( .A1(_f_permutation__round__c[627] ), 
        .A2(_f_permutation__round__n489 ), .ZN(_f_permutation__round__N5525 )
         );
  NOR2_X2 _f_permutation__round__U1539  ( .A1(_f_permutation__round__c[628] ), 
        .A2(_f_permutation__round__n484 ), .ZN(_f_permutation__round__N5523 )
         );
  NOR2_X2 _f_permutation__round__U1538  ( .A1(_f_permutation__round__c[629] ), 
        .A2(_f_permutation__round__n479 ), .ZN(_f_permutation__round__N5521 )
         );
  NOR2_X2 _f_permutation__round__U1537  ( .A1(_f_permutation__round__c[630] ), 
        .A2(_f_permutation__round__n474 ), .ZN(_f_permutation__round__N5519 )
         );
  NOR2_X2 _f_permutation__round__U1536  ( .A1(_f_permutation__round__c[631] ), 
        .A2(_f_permutation__round__n469 ), .ZN(_f_permutation__round__N5517 )
         );
  NOR2_X2 _f_permutation__round__U1535  ( .A1(_f_permutation__round__c[632] ), 
        .A2(_f_permutation__round__n464 ), .ZN(_f_permutation__round__N5515 )
         );
  NOR2_X2 _f_permutation__round__U1534  ( .A1(_f_permutation__round__c[633] ), 
        .A2(_f_permutation__round__n459 ), .ZN(_f_permutation__round__N5513 )
         );
  NOR2_X2 _f_permutation__round__U1533  ( .A1(_f_permutation__round__c[634] ), 
        .A2(_f_permutation__round__n454 ), .ZN(_f_permutation__round__N5511 )
         );
  NOR2_X2 _f_permutation__round__U1532  ( .A1(_f_permutation__round__c[635] ), 
        .A2(_f_permutation__round__n449 ), .ZN(_f_permutation__round__N5509 )
         );
  NOR2_X2 _f_permutation__round__U1531  ( .A1(_f_permutation__round__c[636] ), 
        .A2(_f_permutation__round__n764 ), .ZN(_f_permutation__round__N5507 )
         );
  NOR2_X2 _f_permutation__round__U1530  ( .A1(_f_permutation__round__c[637] ), 
        .A2(_f_permutation__round__n759 ), .ZN(_f_permutation__round__N5505 )
         );
  NOR2_X2 _f_permutation__round__U1529  ( .A1(_f_permutation__round__c[1033] ), 
        .A2(_f_permutation__round__n278 ), .ZN(_f_permutation__round__N5247 )
         );
  NOR2_X2 _f_permutation__round__U1528  ( .A1(_f_permutation__round__c[1034] ), 
        .A2(_f_permutation__round__n271 ), .ZN(_f_permutation__round__N5245 )
         );
  NOR2_X2 _f_permutation__round__U1527  ( .A1(_f_permutation__round__c[1035] ), 
        .A2(_f_permutation__round__n264 ), .ZN(_f_permutation__round__N5243 )
         );
  NOR2_X2 _f_permutation__round__U1526  ( .A1(_f_permutation__round__c[1036] ), 
        .A2(_f_permutation__round__n257 ), .ZN(_f_permutation__round__N5241 )
         );
  NOR2_X2 _f_permutation__round__U1525  ( .A1(_f_permutation__round__c[1037] ), 
        .A2(_f_permutation__round__n250 ), .ZN(_f_permutation__round__N5239 )
         );
  NOR2_X2 _f_permutation__round__U1524  ( .A1(_f_permutation__round__c[1038] ), 
        .A2(_f_permutation__round__n243 ), .ZN(_f_permutation__round__N5237 )
         );
  NOR2_X2 _f_permutation__round__U1523  ( .A1(_f_permutation__round__c[1039] ), 
        .A2(_f_permutation__round__n236 ), .ZN(_f_permutation__round__N5235 )
         );
  NOR2_X2 _f_permutation__round__U1522  ( .A1(_f_permutation__round__c[1040] ), 
        .A2(_f_permutation__round__n229 ), .ZN(_f_permutation__round__N5233 )
         );
  NOR2_X2 _f_permutation__round__U1521  ( .A1(_f_permutation__round__c[1041] ), 
        .A2(_f_permutation__round__n222 ), .ZN(_f_permutation__round__N5231 )
         );
  NOR2_X2 _f_permutation__round__U1520  ( .A1(_f_permutation__round__c[1042] ), 
        .A2(_f_permutation__round__n215 ), .ZN(_f_permutation__round__N5229 )
         );
  NOR2_X2 _f_permutation__round__U1519  ( .A1(_f_permutation__round__c[1043] ), 
        .A2(_f_permutation__round__n208 ), .ZN(_f_permutation__round__N5227 )
         );
  NOR2_X2 _f_permutation__round__U1518  ( .A1(_f_permutation__round__c[1044] ), 
        .A2(_f_permutation__round__n201 ), .ZN(_f_permutation__round__N5225 )
         );
  NOR2_X2 _f_permutation__round__U1517  ( .A1(_f_permutation__round__c[1045] ), 
        .A2(_f_permutation__round__n194 ), .ZN(_f_permutation__round__N5223 )
         );
  NOR2_X2 _f_permutation__round__U1516  ( .A1(_f_permutation__round__c[1046] ), 
        .A2(_f_permutation__round__n187 ), .ZN(_f_permutation__round__N5221 )
         );
  NOR2_X2 _f_permutation__round__U1515  ( .A1(_f_permutation__round__c[1047] ), 
        .A2(_f_permutation__round__n180 ), .ZN(_f_permutation__round__N5219 )
         );
  NOR2_X2 _f_permutation__round__U1514  ( .A1(_f_permutation__round__c[1048] ), 
        .A2(_f_permutation__round__n173 ), .ZN(_f_permutation__round__N5217 )
         );
  NOR2_X2 _f_permutation__round__U1513  ( .A1(_f_permutation__round__c[1049] ), 
        .A2(_f_permutation__round__n166 ), .ZN(_f_permutation__round__N5215 )
         );
  NOR2_X2 _f_permutation__round__U1512  ( .A1(_f_permutation__round__c[1050] ), 
        .A2(_f_permutation__round__n159 ), .ZN(_f_permutation__round__N5213 )
         );
  NOR2_X2 _f_permutation__round__U1511  ( .A1(_f_permutation__round__c[1051] ), 
        .A2(_f_permutation__round__n152 ), .ZN(_f_permutation__round__N5211 )
         );
  NOR2_X2 _f_permutation__round__U1510  ( .A1(_f_permutation__round__c[1052] ), 
        .A2(_f_permutation__round__n145 ), .ZN(_f_permutation__round__N5209 )
         );
  NOR2_X2 _f_permutation__round__U1509  ( .A1(_f_permutation__round__c[1053] ), 
        .A2(_f_permutation__round__n138 ), .ZN(_f_permutation__round__N5207 )
         );
  NOR2_X2 _f_permutation__round__U1508  ( .A1(_f_permutation__round__c[1054] ), 
        .A2(_f_permutation__round__n131 ), .ZN(_f_permutation__round__N5205 )
         );
  NOR2_X2 _f_permutation__round__U1507  ( .A1(_f_permutation__round__c[1055] ), 
        .A2(_f_permutation__round__n124 ), .ZN(_f_permutation__round__N5203 )
         );
  NOR2_X2 _f_permutation__round__U1506  ( .A1(_f_permutation__round__c[1056] ), 
        .A2(_f_permutation__round__n117 ), .ZN(_f_permutation__round__N5201 )
         );
  NOR2_X2 _f_permutation__round__U1505  ( .A1(_f_permutation__round__c[1057] ), 
        .A2(_f_permutation__round__n110 ), .ZN(_f_permutation__round__N5199 )
         );
  NOR2_X2 _f_permutation__round__U1504  ( .A1(_f_permutation__round__c[1058] ), 
        .A2(_f_permutation__round__n103 ), .ZN(_f_permutation__round__N5197 )
         );
  NOR2_X2 _f_permutation__round__U1503  ( .A1(_f_permutation__round__c[1059] ), 
        .A2(_f_permutation__round__n96 ), .ZN(_f_permutation__round__N5195 )
         );
  NOR2_X2 _f_permutation__round__U1502  ( .A1(_f_permutation__round__c[1060] ), 
        .A2(_f_permutation__round__n89 ), .ZN(_f_permutation__round__N5193 )
         );
  NOR2_X2 _f_permutation__round__U1501  ( .A1(_f_permutation__round__c[1061] ), 
        .A2(_f_permutation__round__n82 ), .ZN(_f_permutation__round__N5191 )
         );
  NOR2_X2 _f_permutation__round__U1500  ( .A1(_f_permutation__round__c[1062] ), 
        .A2(_f_permutation__round__n75 ), .ZN(_f_permutation__round__N5189 )
         );
  NOR2_X2 _f_permutation__round__U1499  ( .A1(_f_permutation__round__c[1063] ), 
        .A2(_f_permutation__round__n68 ), .ZN(_f_permutation__round__N5187 )
         );
  NOR2_X2 _f_permutation__round__U1498  ( .A1(_f_permutation__round__c[1064] ), 
        .A2(_f_permutation__round__n61 ), .ZN(_f_permutation__round__N5185 )
         );
  NOR2_X2 _f_permutation__round__U1497  ( .A1(_f_permutation__round__c[1065] ), 
        .A2(_f_permutation__round__n54 ), .ZN(_f_permutation__round__N5183 )
         );
  NOR2_X2 _f_permutation__round__U1496  ( .A1(_f_permutation__round__c[1066] ), 
        .A2(_f_permutation__round__n47 ), .ZN(_f_permutation__round__N5181 )
         );
  NOR2_X2 _f_permutation__round__U1495  ( .A1(_f_permutation__round__c[1067] ), 
        .A2(_f_permutation__round__n40 ), .ZN(_f_permutation__round__N5179 )
         );
  NOR2_X2 _f_permutation__round__U1494  ( .A1(_f_permutation__round__c[1068] ), 
        .A2(_f_permutation__round__n33 ), .ZN(_f_permutation__round__N5177 )
         );
  NOR2_X2 _f_permutation__round__U1493  ( .A1(_f_permutation__round__c[1069] ), 
        .A2(_f_permutation__round__n26 ), .ZN(_f_permutation__round__N5175 )
         );
  NOR2_X2 _f_permutation__round__U1492  ( .A1(_f_permutation__round__c[1070] ), 
        .A2(_f_permutation__round__n19 ), .ZN(_f_permutation__round__N5173 )
         );
  NOR2_X2 _f_permutation__round__U1491  ( .A1(_f_permutation__round__c[1071] ), 
        .A2(_f_permutation__round__n12 ), .ZN(_f_permutation__round__N5171 )
         );
  NOR2_X2 _f_permutation__round__U1490  ( .A1(_f_permutation__round__c[1072] ), 
        .A2(_f_permutation__round__n5 ), .ZN(_f_permutation__round__N5169 ) );
  NOR2_X2 _f_permutation__round__U1489  ( .A1(_f_permutation__round__c[1073] ), 
        .A2(_f_permutation__round__n446 ), .ZN(_f_permutation__round__N5167 )
         );
  NOR2_X2 _f_permutation__round__U1488  ( .A1(_f_permutation__round__c[1074] ), 
        .A2(_f_permutation__round__n439 ), .ZN(_f_permutation__round__N5165 )
         );
  NOR2_X2 _f_permutation__round__U1487  ( .A1(_f_permutation__round__c[1075] ), 
        .A2(_f_permutation__round__n432 ), .ZN(_f_permutation__round__N5163 )
         );
  NOR2_X2 _f_permutation__round__U1486  ( .A1(_f_permutation__round__c[1076] ), 
        .A2(_f_permutation__round__n425 ), .ZN(_f_permutation__round__N5161 )
         );
  NOR2_X2 _f_permutation__round__U1485  ( .A1(_f_permutation__round__c[1077] ), 
        .A2(_f_permutation__round__n418 ), .ZN(_f_permutation__round__N5159 )
         );
  NOR2_X2 _f_permutation__round__U1484  ( .A1(_f_permutation__round__c[1078] ), 
        .A2(_f_permutation__round__n411 ), .ZN(_f_permutation__round__N5157 )
         );
  NOR2_X2 _f_permutation__round__U1483  ( .A1(_f_permutation__round__c[1079] ), 
        .A2(_f_permutation__round__n404 ), .ZN(_f_permutation__round__N5155 )
         );
  NOR2_X2 _f_permutation__round__U1482  ( .A1(_f_permutation__round__c[1080] ), 
        .A2(_f_permutation__round__n397 ), .ZN(_f_permutation__round__N5153 )
         );
  NOR2_X2 _f_permutation__round__U1481  ( .A1(_f_permutation__round__c[1081] ), 
        .A2(_f_permutation__round__n390 ), .ZN(_f_permutation__round__N5151 )
         );
  NOR2_X2 _f_permutation__round__U1480  ( .A1(_f_permutation__round__c[1082] ), 
        .A2(_f_permutation__round__n383 ), .ZN(_f_permutation__round__N5149 )
         );
  NOR2_X2 _f_permutation__round__U1479  ( .A1(_f_permutation__round__c[1083] ), 
        .A2(_f_permutation__round__n376 ), .ZN(_f_permutation__round__N5147 )
         );
  NOR2_X2 _f_permutation__round__U1478  ( .A1(_f_permutation__round__c[1084] ), 
        .A2(_f_permutation__round__n369 ), .ZN(_f_permutation__round__N5145 )
         );
  NOR2_X2 _f_permutation__round__U1477  ( .A1(_f_permutation__round__c[1085] ), 
        .A2(_f_permutation__round__n362 ), .ZN(_f_permutation__round__N5143 )
         );
  NOR2_X2 _f_permutation__round__U1476  ( .A1(_f_permutation__round__c[1086] ), 
        .A2(_f_permutation__round__n355 ), .ZN(_f_permutation__round__N5141 )
         );
  NOR2_X2 _f_permutation__round__U1475  ( .A1(_f_permutation__round__c[1087] ), 
        .A2(_f_permutation__round__n348 ), .ZN(_f_permutation__round__N5139 )
         );
  NOR2_X2 _f_permutation__round__U1474  ( .A1(_f_permutation__round__c[1024] ), 
        .A2(_f_permutation__round__n341 ), .ZN(_f_permutation__round__N5137 )
         );
  NOR2_X2 _f_permutation__round__U1473  ( .A1(_f_permutation__round__c[1025] ), 
        .A2(_f_permutation__round__n334 ), .ZN(_f_permutation__round__N5135 )
         );
  NOR2_X2 _f_permutation__round__U1408  ( .A1(_f_permutation__round__c[1026] ), 
        .A2(_f_permutation__round__n327 ), .ZN(_f_permutation__round__N5133 )
         );
  NOR2_X2 _f_permutation__round__U1407  ( .A1(_f_permutation__round__c[1027] ), 
        .A2(_f_permutation__round__n320 ), .ZN(_f_permutation__round__N5131 )
         );
  NOR2_X2 _f_permutation__round__U1406  ( .A1(_f_permutation__round__c[1028] ), 
        .A2(_f_permutation__round__n313 ), .ZN(_f_permutation__round__N5129 )
         );
  NOR2_X2 _f_permutation__round__U1405  ( .A1(_f_permutation__round__c[1029] ), 
        .A2(_f_permutation__round__n306 ), .ZN(_f_permutation__round__N5127 )
         );
  NOR2_X2 _f_permutation__round__U1404  ( .A1(_f_permutation__round__c[1030] ), 
        .A2(_f_permutation__round__n299 ), .ZN(_f_permutation__round__N5125 )
         );
  NOR2_X2 _f_permutation__round__U1403  ( .A1(_f_permutation__round__c[1031] ), 
        .A2(_f_permutation__round__n292 ), .ZN(_f_permutation__round__N5123 )
         );
  NOR2_X2 _f_permutation__round__U1402  ( .A1(_f_permutation__round__c[1032] ), 
        .A2(_f_permutation__round__n285 ), .ZN(_f_permutation__round__N5121 )
         );
  NOR2_X2 _f_permutation__round__U1401  ( .A1(_f_permutation__round__c[1224] ), 
        .A2(_f_permutation__round__n193 ), .ZN(_f_permutation__round__N4991 )
         );
  NOR2_X2 _f_permutation__round__U1400  ( .A1(_f_permutation__round__c[1225] ), 
        .A2(_f_permutation__round__n186 ), .ZN(_f_permutation__round__N4989 )
         );
  NOR2_X2 _f_permutation__round__U1399  ( .A1(_f_permutation__round__c[1226] ), 
        .A2(_f_permutation__round__n179 ), .ZN(_f_permutation__round__N4987 )
         );
  NOR2_X2 _f_permutation__round__U1398  ( .A1(_f_permutation__round__c[1227] ), 
        .A2(_f_permutation__round__n172 ), .ZN(_f_permutation__round__N4985 )
         );
  NOR2_X2 _f_permutation__round__U1397  ( .A1(_f_permutation__round__c[1228] ), 
        .A2(_f_permutation__round__n165 ), .ZN(_f_permutation__round__N4983 )
         );
  NOR2_X2 _f_permutation__round__U1396  ( .A1(_f_permutation__round__c[1229] ), 
        .A2(_f_permutation__round__n158 ), .ZN(_f_permutation__round__N4981 )
         );
  NOR2_X2 _f_permutation__round__U1395  ( .A1(_f_permutation__round__c[1230] ), 
        .A2(_f_permutation__round__n151 ), .ZN(_f_permutation__round__N4979 )
         );
  NOR2_X2 _f_permutation__round__U1394  ( .A1(_f_permutation__round__c[1231] ), 
        .A2(_f_permutation__round__n144 ), .ZN(_f_permutation__round__N4977 )
         );
  NOR2_X2 _f_permutation__round__U1393  ( .A1(_f_permutation__round__c[1232] ), 
        .A2(_f_permutation__round__n137 ), .ZN(_f_permutation__round__N4975 )
         );
  NOR2_X2 _f_permutation__round__U1392  ( .A1(_f_permutation__round__c[1233] ), 
        .A2(_f_permutation__round__n130 ), .ZN(_f_permutation__round__N4973 )
         );
  NOR2_X2 _f_permutation__round__U1391  ( .A1(_f_permutation__round__c[1234] ), 
        .A2(_f_permutation__round__n123 ), .ZN(_f_permutation__round__N4971 )
         );
  NOR2_X2 _f_permutation__round__U1390  ( .A1(_f_permutation__round__c[1235] ), 
        .A2(_f_permutation__round__n116 ), .ZN(_f_permutation__round__N4969 )
         );
  NOR2_X2 _f_permutation__round__U1389  ( .A1(_f_permutation__round__c[1236] ), 
        .A2(_f_permutation__round__n109 ), .ZN(_f_permutation__round__N4967 )
         );
  NOR2_X2 _f_permutation__round__U1388  ( .A1(_f_permutation__round__c[1237] ), 
        .A2(_f_permutation__round__n102 ), .ZN(_f_permutation__round__N4965 )
         );
  NOR2_X2 _f_permutation__round__U1387  ( .A1(_f_permutation__round__c[1238] ), 
        .A2(_f_permutation__round__n95 ), .ZN(_f_permutation__round__N4963 )
         );
  NOR2_X2 _f_permutation__round__U1386  ( .A1(_f_permutation__round__c[1239] ), 
        .A2(_f_permutation__round__n88 ), .ZN(_f_permutation__round__N4961 )
         );
  NOR2_X2 _f_permutation__round__U1385  ( .A1(_f_permutation__round__c[1240] ), 
        .A2(_f_permutation__round__n81 ), .ZN(_f_permutation__round__N4959 )
         );
  NOR2_X2 _f_permutation__round__U1384  ( .A1(_f_permutation__round__c[1241] ), 
        .A2(_f_permutation__round__n74 ), .ZN(_f_permutation__round__N4957 )
         );
  NOR2_X2 _f_permutation__round__U1383  ( .A1(_f_permutation__round__c[1242] ), 
        .A2(_f_permutation__round__n67 ), .ZN(_f_permutation__round__N4955 )
         );
  NOR2_X2 _f_permutation__round__U1382  ( .A1(_f_permutation__round__c[1243] ), 
        .A2(_f_permutation__round__n60 ), .ZN(_f_permutation__round__N4953 )
         );
  NOR2_X2 _f_permutation__round__U1381  ( .A1(_f_permutation__round__c[1244] ), 
        .A2(_f_permutation__round__n53 ), .ZN(_f_permutation__round__N4951 )
         );
  NOR2_X2 _f_permutation__round__U1380  ( .A1(_f_permutation__round__c[1245] ), 
        .A2(_f_permutation__round__n46 ), .ZN(_f_permutation__round__N4949 )
         );
  NOR2_X2 _f_permutation__round__U1379  ( .A1(_f_permutation__round__c[1246] ), 
        .A2(_f_permutation__round__n39 ), .ZN(_f_permutation__round__N4947 )
         );
  NOR2_X2 _f_permutation__round__U1378  ( .A1(_f_permutation__round__c[1247] ), 
        .A2(_f_permutation__round__n32 ), .ZN(_f_permutation__round__N4945 )
         );
  NOR2_X2 _f_permutation__round__U1377  ( .A1(_f_permutation__round__c[1248] ), 
        .A2(_f_permutation__round__n25 ), .ZN(_f_permutation__round__N4943 )
         );
  NOR2_X2 _f_permutation__round__U1376  ( .A1(_f_permutation__round__c[1249] ), 
        .A2(_f_permutation__round__n18 ), .ZN(_f_permutation__round__N4941 )
         );
  NOR2_X2 _f_permutation__round__U1375  ( .A1(_f_permutation__round__c[1250] ), 
        .A2(_f_permutation__round__n11 ), .ZN(_f_permutation__round__N4939 )
         );
  NOR2_X2 _f_permutation__round__U1374  ( .A1(_f_permutation__round__c[1251] ), 
        .A2(_f_permutation__round__n4 ), .ZN(_f_permutation__round__N4937 ) );
  NOR2_X2 _f_permutation__round__U1373  ( .A1(_f_permutation__round__c[1252] ), 
        .A2(_f_permutation__round__n445 ), .ZN(_f_permutation__round__N4935 )
         );
  NOR2_X2 _f_permutation__round__U1372  ( .A1(_f_permutation__round__c[1253] ), 
        .A2(_f_permutation__round__n438 ), .ZN(_f_permutation__round__N4933 )
         );
  NOR2_X2 _f_permutation__round__U1371  ( .A1(_f_permutation__round__c[1254] ), 
        .A2(_f_permutation__round__n431 ), .ZN(_f_permutation__round__N4931 )
         );
  NOR2_X2 _f_permutation__round__U1370  ( .A1(_f_permutation__round__c[1255] ), 
        .A2(_f_permutation__round__n424 ), .ZN(_f_permutation__round__N4929 )
         );
  NOR2_X2 _f_permutation__round__U1369  ( .A1(_f_permutation__round__c[1256] ), 
        .A2(_f_permutation__round__n417 ), .ZN(_f_permutation__round__N4927 )
         );
  NOR2_X2 _f_permutation__round__U1368  ( .A1(_f_permutation__round__c[1257] ), 
        .A2(_f_permutation__round__n410 ), .ZN(_f_permutation__round__N4925 )
         );
  NOR2_X2 _f_permutation__round__U1367  ( .A1(_f_permutation__round__c[1258] ), 
        .A2(_f_permutation__round__n403 ), .ZN(_f_permutation__round__N4923 )
         );
  NOR2_X2 _f_permutation__round__U1366  ( .A1(_f_permutation__round__c[1259] ), 
        .A2(_f_permutation__round__n396 ), .ZN(_f_permutation__round__N4921 )
         );
  NOR2_X2 _f_permutation__round__U1365  ( .A1(_f_permutation__round__c[1260] ), 
        .A2(_f_permutation__round__n389 ), .ZN(_f_permutation__round__N4919 )
         );
  NOR2_X2 _f_permutation__round__U1364  ( .A1(_f_permutation__round__c[1261] ), 
        .A2(_f_permutation__round__n382 ), .ZN(_f_permutation__round__N4917 )
         );
  NOR2_X2 _f_permutation__round__U1363  ( .A1(_f_permutation__round__c[1262] ), 
        .A2(_f_permutation__round__n375 ), .ZN(_f_permutation__round__N4915 )
         );
  NOR2_X2 _f_permutation__round__U1362  ( .A1(_f_permutation__round__c[1263] ), 
        .A2(_f_permutation__round__n368 ), .ZN(_f_permutation__round__N4913 )
         );
  NOR2_X2 _f_permutation__round__U1361  ( .A1(_f_permutation__round__c[1264] ), 
        .A2(_f_permutation__round__n361 ), .ZN(_f_permutation__round__N4911 )
         );
  NOR2_X2 _f_permutation__round__U1360  ( .A1(_f_permutation__round__c[1265] ), 
        .A2(_f_permutation__round__n354 ), .ZN(_f_permutation__round__N4909 )
         );
  NOR2_X2 _f_permutation__round__U1359  ( .A1(_f_permutation__round__c[1266] ), 
        .A2(_f_permutation__round__n347 ), .ZN(_f_permutation__round__N4907 )
         );
  NOR2_X2 _f_permutation__round__U1358  ( .A1(_f_permutation__round__c[1267] ), 
        .A2(_f_permutation__round__n340 ), .ZN(_f_permutation__round__N4905 )
         );
  NOR2_X2 _f_permutation__round__U1357  ( .A1(_f_permutation__round__c[1268] ), 
        .A2(_f_permutation__round__n333 ), .ZN(_f_permutation__round__N4903 )
         );
  NOR2_X2 _f_permutation__round__U1356  ( .A1(_f_permutation__round__c[1269] ), 
        .A2(_f_permutation__round__n326 ), .ZN(_f_permutation__round__N4901 )
         );
  NOR2_X2 _f_permutation__round__U1355  ( .A1(_f_permutation__round__c[1270] ), 
        .A2(_f_permutation__round__n319 ), .ZN(_f_permutation__round__N4899 )
         );
  NOR2_X2 _f_permutation__round__U1354  ( .A1(_f_permutation__round__c[1271] ), 
        .A2(_f_permutation__round__n312 ), .ZN(_f_permutation__round__N4897 )
         );
  NOR2_X2 _f_permutation__round__U1353  ( .A1(_f_permutation__round__c[1272] ), 
        .A2(_f_permutation__round__n305 ), .ZN(_f_permutation__round__N4895 )
         );
  NOR2_X2 _f_permutation__round__U1352  ( .A1(_f_permutation__round__c[1273] ), 
        .A2(_f_permutation__round__n298 ), .ZN(_f_permutation__round__N4893 )
         );
  NOR2_X2 _f_permutation__round__U1351  ( .A1(_f_permutation__round__c[1274] ), 
        .A2(_f_permutation__round__n291 ), .ZN(_f_permutation__round__N4891 )
         );
  NOR2_X2 _f_permutation__round__U1350  ( .A1(_f_permutation__round__c[1275] ), 
        .A2(_f_permutation__round__n284 ), .ZN(_f_permutation__round__N4889 )
         );
  NOR2_X2 _f_permutation__round__U1349  ( .A1(_f_permutation__round__c[1276] ), 
        .A2(_f_permutation__round__n277 ), .ZN(_f_permutation__round__N4887 )
         );
  NOR2_X2 _f_permutation__round__U1348  ( .A1(_f_permutation__round__c[1277] ), 
        .A2(_f_permutation__round__n270 ), .ZN(_f_permutation__round__N4885 )
         );
  NOR2_X2 _f_permutation__round__U1347  ( .A1(_f_permutation__round__c[1278] ), 
        .A2(_f_permutation__round__n263 ), .ZN(_f_permutation__round__N4883 )
         );
  NOR2_X2 _f_permutation__round__U1346  ( .A1(_f_permutation__round__c[1279] ), 
        .A2(_f_permutation__round__n256 ), .ZN(_f_permutation__round__N4881 )
         );
  NOR2_X2 _f_permutation__round__U1345  ( .A1(_f_permutation__round__c[1216] ), 
        .A2(_f_permutation__round__n249 ), .ZN(_f_permutation__round__N4879 )
         );
  NOR2_X2 _f_permutation__round__U1280  ( .A1(_f_permutation__round__c[1217] ), 
        .A2(_f_permutation__round__n242 ), .ZN(_f_permutation__round__N4877 )
         );
  NOR2_X2 _f_permutation__round__U1279  ( .A1(_f_permutation__round__c[1218] ), 
        .A2(_f_permutation__round__n235 ), .ZN(_f_permutation__round__N4875 )
         );
  NOR2_X2 _f_permutation__round__U1278  ( .A1(_f_permutation__round__c[1219] ), 
        .A2(_f_permutation__round__n228 ), .ZN(_f_permutation__round__N4873 )
         );
  NOR2_X2 _f_permutation__round__U1277  ( .A1(_f_permutation__round__c[1220] ), 
        .A2(_f_permutation__round__n221 ), .ZN(_f_permutation__round__N4871 )
         );
  NOR2_X2 _f_permutation__round__U1276  ( .A1(_f_permutation__round__c[1221] ), 
        .A2(_f_permutation__round__n214 ), .ZN(_f_permutation__round__N4869 )
         );
  NOR2_X2 _f_permutation__round__U1275  ( .A1(_f_permutation__round__c[1222] ), 
        .A2(_f_permutation__round__n207 ), .ZN(_f_permutation__round__N4867 )
         );
  NOR2_X2 _f_permutation__round__U1274  ( .A1(_f_permutation__round__c[1223] ), 
        .A2(_f_permutation__round__n200 ), .ZN(_f_permutation__round__N4865 )
         );
  NOR2_X2 _f_permutation__round__U1273  ( .A1(_f_permutation__round__c[92] ), 
        .A2(_f_permutation__round__n65 ), .ZN(_f_permutation__round__N4607 )
         );
  NOR2_X2 _f_permutation__round__U1272  ( .A1(_f_permutation__round__c[93] ), 
        .A2(_f_permutation__round__n58 ), .ZN(_f_permutation__round__N4605 )
         );
  NOR2_X2 _f_permutation__round__U1271  ( .A1(_f_permutation__round__c[94] ), 
        .A2(_f_permutation__round__n51 ), .ZN(_f_permutation__round__N4603 )
         );
  NOR2_X2 _f_permutation__round__U1270  ( .A1(_f_permutation__round__c[95] ), 
        .A2(_f_permutation__round__n44 ), .ZN(_f_permutation__round__N4601 )
         );
  NOR2_X2 _f_permutation__round__U1269  ( .A1(_f_permutation__round__c[96] ), 
        .A2(_f_permutation__round__n37 ), .ZN(_f_permutation__round__N4599 )
         );
  NOR2_X2 _f_permutation__round__U1268  ( .A1(_f_permutation__round__c[97] ), 
        .A2(_f_permutation__round__n30 ), .ZN(_f_permutation__round__N4597 )
         );
  NOR2_X2 _f_permutation__round__U1267  ( .A1(_f_permutation__round__c[98] ), 
        .A2(_f_permutation__round__n23 ), .ZN(_f_permutation__round__N4595 )
         );
  NOR2_X2 _f_permutation__round__U1266  ( .A1(_f_permutation__round__c[99] ), 
        .A2(_f_permutation__round__n16 ), .ZN(_f_permutation__round__N4593 )
         );
  NOR2_X2 _f_permutation__round__U1265  ( .A1(_f_permutation__round__c[100] ), 
        .A2(_f_permutation__round__n9 ), .ZN(_f_permutation__round__N4591 ) );
  NOR2_X2 _f_permutation__round__U1264  ( .A1(_f_permutation__round__c[101] ), 
        .A2(_f_permutation__round__n2 ), .ZN(_f_permutation__round__N4589 ) );
  NOR2_X2 _f_permutation__round__U1263  ( .A1(_f_permutation__round__c[102] ), 
        .A2(_f_permutation__round__n443 ), .ZN(_f_permutation__round__N4587 )
         );
  NOR2_X2 _f_permutation__round__U1262  ( .A1(_f_permutation__round__c[103] ), 
        .A2(_f_permutation__round__n436 ), .ZN(_f_permutation__round__N4585 )
         );
  NOR2_X2 _f_permutation__round__U1261  ( .A1(_f_permutation__round__c[104] ), 
        .A2(_f_permutation__round__n429 ), .ZN(_f_permutation__round__N4583 )
         );
  NOR2_X2 _f_permutation__round__U1260  ( .A1(_f_permutation__round__c[105] ), 
        .A2(_f_permutation__round__n422 ), .ZN(_f_permutation__round__N4581 )
         );
  NOR2_X2 _f_permutation__round__U1259  ( .A1(_f_permutation__round__c[106] ), 
        .A2(_f_permutation__round__n415 ), .ZN(_f_permutation__round__N4579 )
         );
  NOR2_X2 _f_permutation__round__U1258  ( .A1(_f_permutation__round__c[107] ), 
        .A2(_f_permutation__round__n408 ), .ZN(_f_permutation__round__N4577 )
         );
  NOR2_X2 _f_permutation__round__U1257  ( .A1(_f_permutation__round__c[108] ), 
        .A2(_f_permutation__round__n401 ), .ZN(_f_permutation__round__N4575 )
         );
  NOR2_X2 _f_permutation__round__U1256  ( .A1(_f_permutation__round__c[109] ), 
        .A2(_f_permutation__round__n394 ), .ZN(_f_permutation__round__N4573 )
         );
  NOR2_X2 _f_permutation__round__U1255  ( .A1(_f_permutation__round__c[110] ), 
        .A2(_f_permutation__round__n387 ), .ZN(_f_permutation__round__N4571 )
         );
  NOR2_X2 _f_permutation__round__U1254  ( .A1(_f_permutation__round__c[111] ), 
        .A2(_f_permutation__round__n380 ), .ZN(_f_permutation__round__N4569 )
         );
  NOR2_X2 _f_permutation__round__U1253  ( .A1(_f_permutation__round__c[112] ), 
        .A2(_f_permutation__round__n373 ), .ZN(_f_permutation__round__N4567 )
         );
  NOR2_X2 _f_permutation__round__U1252  ( .A1(_f_permutation__round__c[113] ), 
        .A2(_f_permutation__round__n366 ), .ZN(_f_permutation__round__N4565 )
         );
  NOR2_X2 _f_permutation__round__U1251  ( .A1(_f_permutation__round__c[114] ), 
        .A2(_f_permutation__round__n359 ), .ZN(_f_permutation__round__N4563 )
         );
  NOR2_X2 _f_permutation__round__U1250  ( .A1(_f_permutation__round__c[115] ), 
        .A2(_f_permutation__round__n352 ), .ZN(_f_permutation__round__N4561 )
         );
  NOR2_X2 _f_permutation__round__U1249  ( .A1(_f_permutation__round__c[116] ), 
        .A2(_f_permutation__round__n345 ), .ZN(_f_permutation__round__N4559 )
         );
  NOR2_X2 _f_permutation__round__U1248  ( .A1(_f_permutation__round__c[117] ), 
        .A2(_f_permutation__round__n338 ), .ZN(_f_permutation__round__N4557 )
         );
  NOR2_X2 _f_permutation__round__U1247  ( .A1(_f_permutation__round__c[118] ), 
        .A2(_f_permutation__round__n331 ), .ZN(_f_permutation__round__N4555 )
         );
  NOR2_X2 _f_permutation__round__U1246  ( .A1(_f_permutation__round__c[119] ), 
        .A2(_f_permutation__round__n324 ), .ZN(_f_permutation__round__N4553 )
         );
  NOR2_X2 _f_permutation__round__U1245  ( .A1(_f_permutation__round__c[120] ), 
        .A2(_f_permutation__round__n317 ), .ZN(_f_permutation__round__N4551 )
         );
  NOR2_X2 _f_permutation__round__U1244  ( .A1(_f_permutation__round__c[121] ), 
        .A2(_f_permutation__round__n310 ), .ZN(_f_permutation__round__N4549 )
         );
  NOR2_X2 _f_permutation__round__U1243  ( .A1(_f_permutation__round__c[122] ), 
        .A2(_f_permutation__round__n303 ), .ZN(_f_permutation__round__N4547 )
         );
  NOR2_X2 _f_permutation__round__U1242  ( .A1(_f_permutation__round__c[123] ), 
        .A2(_f_permutation__round__n296 ), .ZN(_f_permutation__round__N4545 )
         );
  NOR2_X2 _f_permutation__round__U1241  ( .A1(_f_permutation__round__c[124] ), 
        .A2(_f_permutation__round__n289 ), .ZN(_f_permutation__round__N4543 )
         );
  NOR2_X2 _f_permutation__round__U1240  ( .A1(_f_permutation__round__c[125] ), 
        .A2(_f_permutation__round__n282 ), .ZN(_f_permutation__round__N4541 )
         );
  NOR2_X2 _f_permutation__round__U1239  ( .A1(_f_permutation__round__c[126] ), 
        .A2(_f_permutation__round__n275 ), .ZN(_f_permutation__round__N4539 )
         );
  NOR2_X2 _f_permutation__round__U1238  ( .A1(_f_permutation__round__c[127] ), 
        .A2(_f_permutation__round__n268 ), .ZN(_f_permutation__round__N4537 )
         );
  NOR2_X2 _f_permutation__round__U1237  ( .A1(_f_permutation__round__c[64] ), 
        .A2(_f_permutation__round__n261 ), .ZN(_f_permutation__round__N4535 )
         );
  NOR2_X2 _f_permutation__round__U1236  ( .A1(_f_permutation__round__c[65] ), 
        .A2(_f_permutation__round__n254 ), .ZN(_f_permutation__round__N4533 )
         );
  NOR2_X2 _f_permutation__round__U1235  ( .A1(_f_permutation__round__c[66] ), 
        .A2(_f_permutation__round__n247 ), .ZN(_f_permutation__round__N4531 )
         );
  NOR2_X2 _f_permutation__round__U1234  ( .A1(_f_permutation__round__c[67] ), 
        .A2(_f_permutation__round__n240 ), .ZN(_f_permutation__round__N4529 )
         );
  NOR2_X2 _f_permutation__round__U1233  ( .A1(_f_permutation__round__c[68] ), 
        .A2(_f_permutation__round__n233 ), .ZN(_f_permutation__round__N4527 )
         );
  NOR2_X2 _f_permutation__round__U1232  ( .A1(_f_permutation__round__c[69] ), 
        .A2(_f_permutation__round__n226 ), .ZN(_f_permutation__round__N4525 )
         );
  NOR2_X2 _f_permutation__round__U1231  ( .A1(_f_permutation__round__c[70] ), 
        .A2(_f_permutation__round__n219 ), .ZN(_f_permutation__round__N4523 )
         );
  NOR2_X2 _f_permutation__round__U1230  ( .A1(_f_permutation__round__c[71] ), 
        .A2(_f_permutation__round__n212 ), .ZN(_f_permutation__round__N4521 )
         );
  NOR2_X2 _f_permutation__round__U1229  ( .A1(_f_permutation__round__c[72] ), 
        .A2(_f_permutation__round__n205 ), .ZN(_f_permutation__round__N4519 )
         );
  NOR2_X2 _f_permutation__round__U1228  ( .A1(_f_permutation__round__c[73] ), 
        .A2(_f_permutation__round__n198 ), .ZN(_f_permutation__round__N4517 )
         );
  NOR2_X2 _f_permutation__round__U1227  ( .A1(_f_permutation__round__c[74] ), 
        .A2(_f_permutation__round__n191 ), .ZN(_f_permutation__round__N4515 )
         );
  NOR2_X2 _f_permutation__round__U1226  ( .A1(_f_permutation__round__c[75] ), 
        .A2(_f_permutation__round__n184 ), .ZN(_f_permutation__round__N4513 )
         );
  NOR2_X2 _f_permutation__round__U1225  ( .A1(_f_permutation__round__c[76] ), 
        .A2(_f_permutation__round__n177 ), .ZN(_f_permutation__round__N4511 )
         );
  NOR2_X2 _f_permutation__round__U1224  ( .A1(_f_permutation__round__c[77] ), 
        .A2(_f_permutation__round__n170 ), .ZN(_f_permutation__round__N4509 )
         );
  NOR2_X2 _f_permutation__round__U1223  ( .A1(_f_permutation__round__c[78] ), 
        .A2(_f_permutation__round__n163 ), .ZN(_f_permutation__round__N4507 )
         );
  NOR2_X2 _f_permutation__round__U1222  ( .A1(_f_permutation__round__c[79] ), 
        .A2(_f_permutation__round__n156 ), .ZN(_f_permutation__round__N4505 )
         );
  NOR2_X2 _f_permutation__round__U1221  ( .A1(_f_permutation__round__c[80] ), 
        .A2(_f_permutation__round__n149 ), .ZN(_f_permutation__round__N4503 )
         );
  NOR2_X2 _f_permutation__round__U1220  ( .A1(_f_permutation__round__c[81] ), 
        .A2(_f_permutation__round__n142 ), .ZN(_f_permutation__round__N4501 )
         );
  NOR2_X2 _f_permutation__round__U1219  ( .A1(_f_permutation__round__c[82] ), 
        .A2(_f_permutation__round__n135 ), .ZN(_f_permutation__round__N4499 )
         );
  NOR2_X2 _f_permutation__round__U1218  ( .A1(_f_permutation__round__c[83] ), 
        .A2(_f_permutation__round__n128 ), .ZN(_f_permutation__round__N4497 )
         );
  NOR2_X2 _f_permutation__round__U1217  ( .A1(_f_permutation__round__c[84] ), 
        .A2(_f_permutation__round__n121 ), .ZN(_f_permutation__round__N4495 )
         );
  NOR2_X2 _f_permutation__round__U1216  ( .A1(_f_permutation__round__c[85] ), 
        .A2(_f_permutation__round__n114 ), .ZN(_f_permutation__round__N4493 )
         );
  NOR2_X2 _f_permutation__round__U1215  ( .A1(_f_permutation__round__c[86] ), 
        .A2(_f_permutation__round__n107 ), .ZN(_f_permutation__round__N4491 )
         );
  NOR2_X2 _f_permutation__round__U1214  ( .A1(_f_permutation__round__c[87] ), 
        .A2(_f_permutation__round__n100 ), .ZN(_f_permutation__round__N4489 )
         );
  NOR2_X2 _f_permutation__round__U1213  ( .A1(_f_permutation__round__c[88] ), 
        .A2(_f_permutation__round__n93 ), .ZN(_f_permutation__round__N4487 )
         );
  NOR2_X2 _f_permutation__round__U1212  ( .A1(_f_permutation__round__c[89] ), 
        .A2(_f_permutation__round__n86 ), .ZN(_f_permutation__round__N4485 )
         );
  NOR2_X2 _f_permutation__round__U1211  ( .A1(_f_permutation__round__c[90] ), 
        .A2(_f_permutation__round__n79 ), .ZN(_f_permutation__round__N4483 )
         );
  NOR2_X2 _f_permutation__round__U1210  ( .A1(_f_permutation__round__c[91] ), 
        .A2(_f_permutation__round__n72 ), .ZN(_f_permutation__round__N4481 )
         );
  NOR2_X2 _f_permutation__round__U1209  ( .A1(_f_permutation__round__c[302] ), 
        .A2(_f_permutation__round__n1 ), .ZN(_f_permutation__round__N4351 ) );
  NOR2_X2 _f_permutation__round__U1208  ( .A1(_f_permutation__round__c[303] ), 
        .A2(_f_permutation__round__n442 ), .ZN(_f_permutation__round__N4349 )
         );
  NOR2_X2 _f_permutation__round__U1207  ( .A1(_f_permutation__round__c[304] ), 
        .A2(_f_permutation__round__n435 ), .ZN(_f_permutation__round__N4347 )
         );
  NOR2_X2 _f_permutation__round__U1206  ( .A1(_f_permutation__round__c[305] ), 
        .A2(_f_permutation__round__n428 ), .ZN(_f_permutation__round__N4345 )
         );
  NOR2_X2 _f_permutation__round__U1205  ( .A1(_f_permutation__round__c[306] ), 
        .A2(_f_permutation__round__n421 ), .ZN(_f_permutation__round__N4343 )
         );
  NOR2_X2 _f_permutation__round__U1204  ( .A1(_f_permutation__round__c[307] ), 
        .A2(_f_permutation__round__n414 ), .ZN(_f_permutation__round__N4341 )
         );
  NOR2_X2 _f_permutation__round__U1203  ( .A1(_f_permutation__round__c[308] ), 
        .A2(_f_permutation__round__n407 ), .ZN(_f_permutation__round__N4339 )
         );
  NOR2_X2 _f_permutation__round__U1202  ( .A1(_f_permutation__round__c[309] ), 
        .A2(_f_permutation__round__n400 ), .ZN(_f_permutation__round__N4337 )
         );
  NOR2_X2 _f_permutation__round__U1201  ( .A1(_f_permutation__round__c[310] ), 
        .A2(_f_permutation__round__n393 ), .ZN(_f_permutation__round__N4335 )
         );
  NOR2_X2 _f_permutation__round__U1200  ( .A1(_f_permutation__round__c[311] ), 
        .A2(_f_permutation__round__n386 ), .ZN(_f_permutation__round__N4333 )
         );
  NOR2_X2 _f_permutation__round__U1199  ( .A1(_f_permutation__round__c[312] ), 
        .A2(_f_permutation__round__n379 ), .ZN(_f_permutation__round__N4331 )
         );
  NOR2_X2 _f_permutation__round__U1198  ( .A1(_f_permutation__round__c[313] ), 
        .A2(_f_permutation__round__n372 ), .ZN(_f_permutation__round__N4329 )
         );
  NOR2_X2 _f_permutation__round__U1197  ( .A1(_f_permutation__round__c[314] ), 
        .A2(_f_permutation__round__n365 ), .ZN(_f_permutation__round__N4327 )
         );
  NOR2_X2 _f_permutation__round__U1196  ( .A1(_f_permutation__round__c[315] ), 
        .A2(_f_permutation__round__n358 ), .ZN(_f_permutation__round__N4325 )
         );
  NOR2_X2 _f_permutation__round__U1195  ( .A1(_f_permutation__round__c[316] ), 
        .A2(_f_permutation__round__n351 ), .ZN(_f_permutation__round__N4323 )
         );
  NOR2_X2 _f_permutation__round__U1194  ( .A1(_f_permutation__round__c[317] ), 
        .A2(_f_permutation__round__n344 ), .ZN(_f_permutation__round__N4321 )
         );
  NOR2_X2 _f_permutation__round__U1193  ( .A1(_f_permutation__round__c[318] ), 
        .A2(_f_permutation__round__n337 ), .ZN(_f_permutation__round__N4319 )
         );
  NOR2_X2 _f_permutation__round__U1192  ( .A1(_f_permutation__round__c[319] ), 
        .A2(_f_permutation__round__n330 ), .ZN(_f_permutation__round__N4317 )
         );
  NOR2_X2 _f_permutation__round__U1191  ( .A1(_f_permutation__round__c[256] ), 
        .A2(_f_permutation__round__n323 ), .ZN(_f_permutation__round__N4315 )
         );
  NOR2_X2 _f_permutation__round__U1190  ( .A1(_f_permutation__round__c[257] ), 
        .A2(_f_permutation__round__n316 ), .ZN(_f_permutation__round__N4313 )
         );
  NOR2_X2 _f_permutation__round__U1189  ( .A1(_f_permutation__round__c[258] ), 
        .A2(_f_permutation__round__n309 ), .ZN(_f_permutation__round__N4311 )
         );
  NOR2_X2 _f_permutation__round__U1188  ( .A1(_f_permutation__round__c[259] ), 
        .A2(_f_permutation__round__n302 ), .ZN(_f_permutation__round__N4309 )
         );
  NOR2_X2 _f_permutation__round__U1187  ( .A1(_f_permutation__round__c[260] ), 
        .A2(_f_permutation__round__n295 ), .ZN(_f_permutation__round__N4307 )
         );
  NOR2_X2 _f_permutation__round__U1186  ( .A1(_f_permutation__round__c[261] ), 
        .A2(_f_permutation__round__n288 ), .ZN(_f_permutation__round__N4305 )
         );
  NOR2_X2 _f_permutation__round__U1185  ( .A1(_f_permutation__round__c[262] ), 
        .A2(_f_permutation__round__n281 ), .ZN(_f_permutation__round__N4303 )
         );
  NOR2_X2 _f_permutation__round__U1184  ( .A1(_f_permutation__round__c[263] ), 
        .A2(_f_permutation__round__n274 ), .ZN(_f_permutation__round__N4301 )
         );
  NOR2_X2 _f_permutation__round__U1183  ( .A1(_f_permutation__round__c[264] ), 
        .A2(_f_permutation__round__n267 ), .ZN(_f_permutation__round__N4299 )
         );
  NOR2_X2 _f_permutation__round__U1182  ( .A1(_f_permutation__round__c[265] ), 
        .A2(_f_permutation__round__n260 ), .ZN(_f_permutation__round__N4297 )
         );
  NOR2_X2 _f_permutation__round__U1181  ( .A1(_f_permutation__round__c[266] ), 
        .A2(_f_permutation__round__n253 ), .ZN(_f_permutation__round__N4295 )
         );
  NOR2_X2 _f_permutation__round__U1180  ( .A1(_f_permutation__round__c[267] ), 
        .A2(_f_permutation__round__n246 ), .ZN(_f_permutation__round__N4293 )
         );
  NOR2_X2 _f_permutation__round__U1179  ( .A1(_f_permutation__round__c[268] ), 
        .A2(_f_permutation__round__n239 ), .ZN(_f_permutation__round__N4291 )
         );
  NOR2_X2 _f_permutation__round__U1178  ( .A1(_f_permutation__round__c[269] ), 
        .A2(_f_permutation__round__n232 ), .ZN(_f_permutation__round__N4289 )
         );
  NOR2_X2 _f_permutation__round__U1177  ( .A1(_f_permutation__round__c[270] ), 
        .A2(_f_permutation__round__n225 ), .ZN(_f_permutation__round__N4287 )
         );
  NOR2_X2 _f_permutation__round__U1176  ( .A1(_f_permutation__round__c[271] ), 
        .A2(_f_permutation__round__n218 ), .ZN(_f_permutation__round__N4285 )
         );
  NOR2_X2 _f_permutation__round__U1175  ( .A1(_f_permutation__round__c[272] ), 
        .A2(_f_permutation__round__n211 ), .ZN(_f_permutation__round__N4283 )
         );
  NOR2_X2 _f_permutation__round__U1174  ( .A1(_f_permutation__round__c[273] ), 
        .A2(_f_permutation__round__n204 ), .ZN(_f_permutation__round__N4281 )
         );
  NOR2_X2 _f_permutation__round__U1173  ( .A1(_f_permutation__round__c[274] ), 
        .A2(_f_permutation__round__n197 ), .ZN(_f_permutation__round__N4279 )
         );
  NOR2_X2 _f_permutation__round__U1172  ( .A1(_f_permutation__round__c[275] ), 
        .A2(_f_permutation__round__n190 ), .ZN(_f_permutation__round__N4277 )
         );
  NOR2_X2 _f_permutation__round__U1171  ( .A1(_f_permutation__round__c[276] ), 
        .A2(_f_permutation__round__n183 ), .ZN(_f_permutation__round__N4275 )
         );
  NOR2_X2 _f_permutation__round__U1170  ( .A1(_f_permutation__round__c[277] ), 
        .A2(_f_permutation__round__n176 ), .ZN(_f_permutation__round__N4273 )
         );
  NOR2_X2 _f_permutation__round__U1169  ( .A1(_f_permutation__round__c[278] ), 
        .A2(_f_permutation__round__n169 ), .ZN(_f_permutation__round__N4271 )
         );
  NOR2_X2 _f_permutation__round__U1168  ( .A1(_f_permutation__round__c[279] ), 
        .A2(_f_permutation__round__n162 ), .ZN(_f_permutation__round__N4269 )
         );
  NOR2_X2 _f_permutation__round__U1167  ( .A1(_f_permutation__round__c[280] ), 
        .A2(_f_permutation__round__n155 ), .ZN(_f_permutation__round__N4267 )
         );
  NOR2_X2 _f_permutation__round__U1166  ( .A1(_f_permutation__round__c[281] ), 
        .A2(_f_permutation__round__n148 ), .ZN(_f_permutation__round__N4265 )
         );
  NOR2_X2 _f_permutation__round__U1165  ( .A1(_f_permutation__round__c[282] ), 
        .A2(_f_permutation__round__n141 ), .ZN(_f_permutation__round__N4263 )
         );
  NOR2_X2 _f_permutation__round__U1164  ( .A1(_f_permutation__round__c[283] ), 
        .A2(_f_permutation__round__n134 ), .ZN(_f_permutation__round__N4261 )
         );
  NOR2_X2 _f_permutation__round__U1163  ( .A1(_f_permutation__round__c[284] ), 
        .A2(_f_permutation__round__n127 ), .ZN(_f_permutation__round__N4259 )
         );
  NOR2_X2 _f_permutation__round__U1162  ( .A1(_f_permutation__round__c[285] ), 
        .A2(_f_permutation__round__n120 ), .ZN(_f_permutation__round__N4257 )
         );
  NOR2_X2 _f_permutation__round__U1161  ( .A1(_f_permutation__round__c[286] ), 
        .A2(_f_permutation__round__n113 ), .ZN(_f_permutation__round__N4255 )
         );
  NOR2_X2 _f_permutation__round__U1160  ( .A1(_f_permutation__round__c[287] ), 
        .A2(_f_permutation__round__n106 ), .ZN(_f_permutation__round__N4253 )
         );
  NOR2_X2 _f_permutation__round__U1159  ( .A1(_f_permutation__round__c[288] ), 
        .A2(_f_permutation__round__n99 ), .ZN(_f_permutation__round__N4251 )
         );
  NOR2_X2 _f_permutation__round__U1158  ( .A1(_f_permutation__round__c[289] ), 
        .A2(_f_permutation__round__n92 ), .ZN(_f_permutation__round__N4249 )
         );
  NOR2_X2 _f_permutation__round__U1157  ( .A1(_f_permutation__round__c[290] ), 
        .A2(_f_permutation__round__n85 ), .ZN(_f_permutation__round__N4247 )
         );
  NOR2_X2 _f_permutation__round__U1156  ( .A1(_f_permutation__round__c[291] ), 
        .A2(_f_permutation__round__n78 ), .ZN(_f_permutation__round__N4245 )
         );
  NOR2_X2 _f_permutation__round__U1155  ( .A1(_f_permutation__round__c[292] ), 
        .A2(_f_permutation__round__n71 ), .ZN(_f_permutation__round__N4243 )
         );
  NOR2_X2 _f_permutation__round__U1154  ( .A1(_f_permutation__round__c[293] ), 
        .A2(_f_permutation__round__n64 ), .ZN(_f_permutation__round__N4241 )
         );
  NOR2_X2 _f_permutation__round__U1153  ( .A1(_f_permutation__round__c[294] ), 
        .A2(_f_permutation__round__n57 ), .ZN(_f_permutation__round__N4239 )
         );
  NOR2_X2 _f_permutation__round__U1088  ( .A1(_f_permutation__round__c[295] ), 
        .A2(_f_permutation__round__n50 ), .ZN(_f_permutation__round__N4237 )
         );
  NOR2_X2 _f_permutation__round__U1087  ( .A1(_f_permutation__round__c[296] ), 
        .A2(_f_permutation__round__n43 ), .ZN(_f_permutation__round__N4235 )
         );
  NOR2_X2 _f_permutation__round__U1086  ( .A1(_f_permutation__round__c[297] ), 
        .A2(_f_permutation__round__n36 ), .ZN(_f_permutation__round__N4233 )
         );
  NOR2_X2 _f_permutation__round__U1085  ( .A1(_f_permutation__round__c[298] ), 
        .A2(_f_permutation__round__n29 ), .ZN(_f_permutation__round__N4231 )
         );
  NOR2_X2 _f_permutation__round__U1084  ( .A1(_f_permutation__round__c[299] ), 
        .A2(_f_permutation__round__n22 ), .ZN(_f_permutation__round__N4229 )
         );
  NOR2_X2 _f_permutation__round__U1083  ( .A1(_f_permutation__round__c[300] ), 
        .A2(_f_permutation__round__n15 ), .ZN(_f_permutation__round__N4227 )
         );
  NOR2_X2 _f_permutation__round__U1082  ( .A1(_f_permutation__round__c[301] ), 
        .A2(_f_permutation__round__n8 ), .ZN(_f_permutation__round__N4225 ) );
  NOR2_X2 _f_permutation__round__U1081  ( .A1(_f_permutation__round__c[762] ), 
        .A2(_f_permutation__round__n842 ), .ZN(_f_permutation__round__N3967 )
         );
  NOR2_X2 _f_permutation__round__U1080  ( .A1(_f_permutation__round__c[763] ), 
        .A2(_f_permutation__round__n839 ), .ZN(_f_permutation__round__N3965 )
         );
  NOR2_X2 _f_permutation__round__U1079  ( .A1(_f_permutation__round__c[764] ), 
        .A2(_f_permutation__round__n836 ), .ZN(_f_permutation__round__N3963 )
         );
  NOR2_X2 _f_permutation__round__U1078  ( .A1(_f_permutation__round__c[765] ), 
        .A2(_f_permutation__round__n833 ), .ZN(_f_permutation__round__N3961 )
         );
  NOR2_X2 _f_permutation__round__U1077  ( .A1(_f_permutation__round__c[766] ), 
        .A2(_f_permutation__round__n830 ), .ZN(_f_permutation__round__N3959 )
         );
  NOR2_X2 _f_permutation__round__U1076  ( .A1(_f_permutation__round__c[767] ), 
        .A2(_f_permutation__round__n827 ), .ZN(_f_permutation__round__N3957 )
         );
  NOR2_X2 _f_permutation__round__U1075  ( .A1(_f_permutation__round__c[704] ), 
        .A2(_f_permutation__round__n824 ), .ZN(_f_permutation__round__N3955 )
         );
  NOR2_X2 _f_permutation__round__U1074  ( .A1(_f_permutation__round__c[705] ), 
        .A2(_f_permutation__round__n821 ), .ZN(_f_permutation__round__N3953 )
         );
  NOR2_X2 _f_permutation__round__U1073  ( .A1(_f_permutation__round__c[706] ), 
        .A2(_f_permutation__round__n818 ), .ZN(_f_permutation__round__N3951 )
         );
  NOR2_X2 _f_permutation__round__U1072  ( .A1(_f_permutation__round__c[707] ), 
        .A2(_f_permutation__round__n815 ), .ZN(_f_permutation__round__N3949 )
         );
  NOR2_X2 _f_permutation__round__U1071  ( .A1(_f_permutation__round__c[708] ), 
        .A2(_f_permutation__round__n812 ), .ZN(_f_permutation__round__N3947 )
         );
  NOR2_X2 _f_permutation__round__U1070  ( .A1(_f_permutation__round__c[709] ), 
        .A2(_f_permutation__round__n809 ), .ZN(_f_permutation__round__N3945 )
         );
  NOR2_X2 _f_permutation__round__U1069  ( .A1(_f_permutation__round__c[710] ), 
        .A2(_f_permutation__round__n806 ), .ZN(_f_permutation__round__N3943 )
         );
  NOR2_X2 _f_permutation__round__U1068  ( .A1(_f_permutation__round__c[711] ), 
        .A2(_f_permutation__round__n803 ), .ZN(_f_permutation__round__N3941 )
         );
  NOR2_X2 _f_permutation__round__U1067  ( .A1(_f_permutation__round__c[712] ), 
        .A2(_f_permutation__round__n800 ), .ZN(_f_permutation__round__N3939 )
         );
  NOR2_X2 _f_permutation__round__U1066  ( .A1(_f_permutation__round__c[713] ), 
        .A2(_f_permutation__round__n797 ), .ZN(_f_permutation__round__N3937 )
         );
  NOR2_X2 _f_permutation__round__U1065  ( .A1(_f_permutation__round__c[714] ), 
        .A2(_f_permutation__round__n794 ), .ZN(_f_permutation__round__N3935 )
         );
  NOR2_X2 _f_permutation__round__U1064  ( .A1(_f_permutation__round__c[715] ), 
        .A2(_f_permutation__round__n791 ), .ZN(_f_permutation__round__N3933 )
         );
  NOR2_X2 _f_permutation__round__U1063  ( .A1(_f_permutation__round__c[716] ), 
        .A2(_f_permutation__round__n788 ), .ZN(_f_permutation__round__N3931 )
         );
  NOR2_X2 _f_permutation__round__U1062  ( .A1(_f_permutation__round__c[717] ), 
        .A2(_f_permutation__round__n785 ), .ZN(_f_permutation__round__N3929 )
         );
  NOR2_X2 _f_permutation__round__U1061  ( .A1(_f_permutation__round__c[718] ), 
        .A2(_f_permutation__round__n782 ), .ZN(_f_permutation__round__N3927 )
         );
  NOR2_X2 _f_permutation__round__U1060  ( .A1(_f_permutation__round__c[719] ), 
        .A2(_f_permutation__round__n779 ), .ZN(_f_permutation__round__N3925 )
         );
  NOR2_X2 _f_permutation__round__U1059  ( .A1(_f_permutation__round__c[720] ), 
        .A2(_f_permutation__round__n776 ), .ZN(_f_permutation__round__N3923 )
         );
  NOR2_X2 _f_permutation__round__U1058  ( .A1(_f_permutation__round__c[721] ), 
        .A2(_f_permutation__round__n773 ), .ZN(_f_permutation__round__N3921 )
         );
  NOR2_X2 _f_permutation__round__U1057  ( .A1(_f_permutation__round__c[722] ), 
        .A2(_f_permutation__round__n770 ), .ZN(_f_permutation__round__N3919 )
         );
  NOR2_X2 _f_permutation__round__U1056  ( .A1(_f_permutation__round__c[723] ), 
        .A2(_f_permutation__round__n959 ), .ZN(_f_permutation__round__N3917 )
         );
  NOR2_X2 _f_permutation__round__U1055  ( .A1(_f_permutation__round__c[724] ), 
        .A2(_f_permutation__round__n956 ), .ZN(_f_permutation__round__N3915 )
         );
  NOR2_X2 _f_permutation__round__U1054  ( .A1(_f_permutation__round__c[725] ), 
        .A2(_f_permutation__round__n953 ), .ZN(_f_permutation__round__N3913 )
         );
  NOR2_X2 _f_permutation__round__U1053  ( .A1(_f_permutation__round__c[726] ), 
        .A2(_f_permutation__round__n950 ), .ZN(_f_permutation__round__N3911 )
         );
  NOR2_X2 _f_permutation__round__U1052  ( .A1(_f_permutation__round__c[727] ), 
        .A2(_f_permutation__round__n947 ), .ZN(_f_permutation__round__N3909 )
         );
  NOR2_X2 _f_permutation__round__U1051  ( .A1(_f_permutation__round__c[728] ), 
        .A2(_f_permutation__round__n944 ), .ZN(_f_permutation__round__N3907 )
         );
  NOR2_X2 _f_permutation__round__U1050  ( .A1(_f_permutation__round__c[729] ), 
        .A2(_f_permutation__round__n941 ), .ZN(_f_permutation__round__N3905 )
         );
  NOR2_X2 _f_permutation__round__U1049  ( .A1(_f_permutation__round__c[730] ), 
        .A2(_f_permutation__round__n938 ), .ZN(_f_permutation__round__N3903 )
         );
  NOR2_X2 _f_permutation__round__U1048  ( .A1(_f_permutation__round__c[731] ), 
        .A2(_f_permutation__round__n935 ), .ZN(_f_permutation__round__N3901 )
         );
  NOR2_X2 _f_permutation__round__U1047  ( .A1(_f_permutation__round__c[732] ), 
        .A2(_f_permutation__round__n932 ), .ZN(_f_permutation__round__N3899 )
         );
  NOR2_X2 _f_permutation__round__U1046  ( .A1(_f_permutation__round__c[733] ), 
        .A2(_f_permutation__round__n929 ), .ZN(_f_permutation__round__N3897 )
         );
  NOR2_X2 _f_permutation__round__U1045  ( .A1(_f_permutation__round__c[734] ), 
        .A2(_f_permutation__round__n926 ), .ZN(_f_permutation__round__N3895 )
         );
  NOR2_X2 _f_permutation__round__U1044  ( .A1(_f_permutation__round__c[735] ), 
        .A2(_f_permutation__round__n923 ), .ZN(_f_permutation__round__N3893 )
         );
  NOR2_X2 _f_permutation__round__U1043  ( .A1(_f_permutation__round__c[736] ), 
        .A2(_f_permutation__round__n920 ), .ZN(_f_permutation__round__N3891 )
         );
  NOR2_X2 _f_permutation__round__U1042  ( .A1(_f_permutation__round__c[737] ), 
        .A2(_f_permutation__round__n917 ), .ZN(_f_permutation__round__N3889 )
         );
  NOR2_X2 _f_permutation__round__U1041  ( .A1(_f_permutation__round__c[738] ), 
        .A2(_f_permutation__round__n914 ), .ZN(_f_permutation__round__N3887 )
         );
  NOR2_X2 _f_permutation__round__U1040  ( .A1(_f_permutation__round__c[739] ), 
        .A2(_f_permutation__round__n911 ), .ZN(_f_permutation__round__N3885 )
         );
  NOR2_X2 _f_permutation__round__U1039  ( .A1(_f_permutation__round__c[740] ), 
        .A2(_f_permutation__round__n908 ), .ZN(_f_permutation__round__N3883 )
         );
  NOR2_X2 _f_permutation__round__U1038  ( .A1(_f_permutation__round__c[741] ), 
        .A2(_f_permutation__round__n905 ), .ZN(_f_permutation__round__N3881 )
         );
  NOR2_X2 _f_permutation__round__U1037  ( .A1(_f_permutation__round__c[742] ), 
        .A2(_f_permutation__round__n902 ), .ZN(_f_permutation__round__N3879 )
         );
  NOR2_X2 _f_permutation__round__U1036  ( .A1(_f_permutation__round__c[743] ), 
        .A2(_f_permutation__round__n899 ), .ZN(_f_permutation__round__N3877 )
         );
  NOR2_X2 _f_permutation__round__U1035  ( .A1(_f_permutation__round__c[744] ), 
        .A2(_f_permutation__round__n896 ), .ZN(_f_permutation__round__N3875 )
         );
  NOR2_X2 _f_permutation__round__U1034  ( .A1(_f_permutation__round__c[745] ), 
        .A2(_f_permutation__round__n893 ), .ZN(_f_permutation__round__N3873 )
         );
  NOR2_X2 _f_permutation__round__U1033  ( .A1(_f_permutation__round__c[746] ), 
        .A2(_f_permutation__round__n890 ), .ZN(_f_permutation__round__N3871 )
         );
  NOR2_X2 _f_permutation__round__U1032  ( .A1(_f_permutation__round__c[747] ), 
        .A2(_f_permutation__round__n887 ), .ZN(_f_permutation__round__N3869 )
         );
  NOR2_X2 _f_permutation__round__U1031  ( .A1(_f_permutation__round__c[748] ), 
        .A2(_f_permutation__round__n884 ), .ZN(_f_permutation__round__N3867 )
         );
  NOR2_X2 _f_permutation__round__U1030  ( .A1(_f_permutation__round__c[749] ), 
        .A2(_f_permutation__round__n881 ), .ZN(_f_permutation__round__N3865 )
         );
  NOR2_X2 _f_permutation__round__U1029  ( .A1(_f_permutation__round__c[750] ), 
        .A2(_f_permutation__round__n878 ), .ZN(_f_permutation__round__N3863 )
         );
  NOR2_X2 _f_permutation__round__U1028  ( .A1(_f_permutation__round__c[751] ), 
        .A2(_f_permutation__round__n875 ), .ZN(_f_permutation__round__N3861 )
         );
  NOR2_X2 _f_permutation__round__U1027  ( .A1(_f_permutation__round__c[752] ), 
        .A2(_f_permutation__round__n872 ), .ZN(_f_permutation__round__N3859 )
         );
  NOR2_X2 _f_permutation__round__U1026  ( .A1(_f_permutation__round__c[753] ), 
        .A2(_f_permutation__round__n869 ), .ZN(_f_permutation__round__N3857 )
         );
  NOR2_X2 _f_permutation__round__U1025  ( .A1(_f_permutation__round__c[754] ), 
        .A2(_f_permutation__round__n866 ), .ZN(_f_permutation__round__N3855 )
         );
  NOR2_X2 _f_permutation__round__U960  ( .A1(_f_permutation__round__c[755] ), 
        .A2(_f_permutation__round__n863 ), .ZN(_f_permutation__round__N3853 )
         );
  NOR2_X2 _f_permutation__round__U959  ( .A1(_f_permutation__round__c[756] ), 
        .A2(_f_permutation__round__n860 ), .ZN(_f_permutation__round__N3851 )
         );
  NOR2_X2 _f_permutation__round__U958  ( .A1(_f_permutation__round__c[757] ), 
        .A2(_f_permutation__round__n857 ), .ZN(_f_permutation__round__N3849 )
         );
  NOR2_X2 _f_permutation__round__U957  ( .A1(_f_permutation__round__c[758] ), 
        .A2(_f_permutation__round__n854 ), .ZN(_f_permutation__round__N3847 )
         );
  NOR2_X2 _f_permutation__round__U956  ( .A1(_f_permutation__round__c[759] ), 
        .A2(_f_permutation__round__n851 ), .ZN(_f_permutation__round__N3845 )
         );
  NOR2_X2 _f_permutation__round__U955  ( .A1(_f_permutation__round__c[760] ), 
        .A2(_f_permutation__round__n848 ), .ZN(_f_permutation__round__N3843 )
         );
  NOR2_X2 _f_permutation__round__U954  ( .A1(_f_permutation__round__c[761] ), 
        .A2(_f_permutation__round__n845 ), .ZN(_f_permutation__round__N3841 )
         );
  NOR2_X2 _f_permutation__round__U953  ( .A1(_f_permutation__round__c[899] ), 
        .A2(_f_permutation__round__n850 ), .ZN(_f_permutation__round__N3711 )
         );
  NOR2_X2 _f_permutation__round__U952  ( .A1(_f_permutation__round__c[900] ), 
        .A2(_f_permutation__round__n847 ), .ZN(_f_permutation__round__N3709 )
         );
  NOR2_X2 _f_permutation__round__U951  ( .A1(_f_permutation__round__c[901] ), 
        .A2(_f_permutation__round__n844 ), .ZN(_f_permutation__round__N3707 )
         );
  NOR2_X2 _f_permutation__round__U950  ( .A1(_f_permutation__round__c[902] ), 
        .A2(_f_permutation__round__n841 ), .ZN(_f_permutation__round__N3705 )
         );
  NOR2_X2 _f_permutation__round__U949  ( .A1(_f_permutation__round__c[903] ), 
        .A2(_f_permutation__round__n838 ), .ZN(_f_permutation__round__N3703 )
         );
  NOR2_X2 _f_permutation__round__U948  ( .A1(_f_permutation__round__c[904] ), 
        .A2(_f_permutation__round__n835 ), .ZN(_f_permutation__round__N3701 )
         );
  NOR2_X2 _f_permutation__round__U947  ( .A1(_f_permutation__round__c[905] ), 
        .A2(_f_permutation__round__n832 ), .ZN(_f_permutation__round__N3699 )
         );
  NOR2_X2 _f_permutation__round__U946  ( .A1(_f_permutation__round__c[906] ), 
        .A2(_f_permutation__round__n829 ), .ZN(_f_permutation__round__N3697 )
         );
  NOR2_X2 _f_permutation__round__U945  ( .A1(_f_permutation__round__c[907] ), 
        .A2(_f_permutation__round__n826 ), .ZN(_f_permutation__round__N3695 )
         );
  NOR2_X2 _f_permutation__round__U944  ( .A1(_f_permutation__round__c[908] ), 
        .A2(_f_permutation__round__n823 ), .ZN(_f_permutation__round__N3693 )
         );
  NOR2_X2 _f_permutation__round__U943  ( .A1(_f_permutation__round__c[909] ), 
        .A2(_f_permutation__round__n820 ), .ZN(_f_permutation__round__N3691 )
         );
  NOR2_X2 _f_permutation__round__U942  ( .A1(_f_permutation__round__c[910] ), 
        .A2(_f_permutation__round__n817 ), .ZN(_f_permutation__round__N3689 )
         );
  NOR2_X2 _f_permutation__round__U941  ( .A1(_f_permutation__round__c[911] ), 
        .A2(_f_permutation__round__n814 ), .ZN(_f_permutation__round__N3687 )
         );
  NOR2_X2 _f_permutation__round__U940  ( .A1(_f_permutation__round__c[912] ), 
        .A2(_f_permutation__round__n811 ), .ZN(_f_permutation__round__N3685 )
         );
  NOR2_X2 _f_permutation__round__U939  ( .A1(_f_permutation__round__c[913] ), 
        .A2(_f_permutation__round__n808 ), .ZN(_f_permutation__round__N3683 )
         );
  NOR2_X2 _f_permutation__round__U938  ( .A1(_f_permutation__round__c[914] ), 
        .A2(_f_permutation__round__n805 ), .ZN(_f_permutation__round__N3681 )
         );
  NOR2_X2 _f_permutation__round__U937  ( .A1(_f_permutation__round__c[915] ), 
        .A2(_f_permutation__round__n802 ), .ZN(_f_permutation__round__N3679 )
         );
  NOR2_X2 _f_permutation__round__U936  ( .A1(_f_permutation__round__c[916] ), 
        .A2(_f_permutation__round__n799 ), .ZN(_f_permutation__round__N3677 )
         );
  NOR2_X2 _f_permutation__round__U935  ( .A1(_f_permutation__round__c[917] ), 
        .A2(_f_permutation__round__n796 ), .ZN(_f_permutation__round__N3675 )
         );
  NOR2_X2 _f_permutation__round__U934  ( .A1(_f_permutation__round__c[918] ), 
        .A2(_f_permutation__round__n793 ), .ZN(_f_permutation__round__N3673 )
         );
  NOR2_X2 _f_permutation__round__U933  ( .A1(_f_permutation__round__c[919] ), 
        .A2(_f_permutation__round__n790 ), .ZN(_f_permutation__round__N3671 )
         );
  NOR2_X2 _f_permutation__round__U932  ( .A1(_f_permutation__round__c[920] ), 
        .A2(_f_permutation__round__n787 ), .ZN(_f_permutation__round__N3669 )
         );
  NOR2_X2 _f_permutation__round__U931  ( .A1(_f_permutation__round__c[921] ), 
        .A2(_f_permutation__round__n784 ), .ZN(_f_permutation__round__N3667 )
         );
  NOR2_X2 _f_permutation__round__U930  ( .A1(_f_permutation__round__c[922] ), 
        .A2(_f_permutation__round__n781 ), .ZN(_f_permutation__round__N3665 )
         );
  NOR2_X2 _f_permutation__round__U929  ( .A1(_f_permutation__round__c[923] ), 
        .A2(_f_permutation__round__n778 ), .ZN(_f_permutation__round__N3663 )
         );
  NOR2_X2 _f_permutation__round__U928  ( .A1(_f_permutation__round__c[924] ), 
        .A2(_f_permutation__round__n775 ), .ZN(_f_permutation__round__N3661 )
         );
  NOR2_X2 _f_permutation__round__U927  ( .A1(_f_permutation__round__c[925] ), 
        .A2(_f_permutation__round__n772 ), .ZN(_f_permutation__round__N3659 )
         );
  NOR2_X2 _f_permutation__round__U926  ( .A1(_f_permutation__round__c[926] ), 
        .A2(_f_permutation__round__n769 ), .ZN(_f_permutation__round__N3657 )
         );
  NOR2_X2 _f_permutation__round__U925  ( .A1(_f_permutation__round__c[927] ), 
        .A2(_f_permutation__round__n958 ), .ZN(_f_permutation__round__N3655 )
         );
  NOR2_X2 _f_permutation__round__U924  ( .A1(_f_permutation__round__c[928] ), 
        .A2(_f_permutation__round__n955 ), .ZN(_f_permutation__round__N3653 )
         );
  NOR2_X2 _f_permutation__round__U923  ( .A1(_f_permutation__round__c[929] ), 
        .A2(_f_permutation__round__n952 ), .ZN(_f_permutation__round__N3651 )
         );
  NOR2_X2 _f_permutation__round__U922  ( .A1(_f_permutation__round__c[930] ), 
        .A2(_f_permutation__round__n949 ), .ZN(_f_permutation__round__N3649 )
         );
  NOR2_X2 _f_permutation__round__U921  ( .A1(_f_permutation__round__c[931] ), 
        .A2(_f_permutation__round__n946 ), .ZN(_f_permutation__round__N3647 )
         );
  NOR2_X2 _f_permutation__round__U920  ( .A1(_f_permutation__round__c[932] ), 
        .A2(_f_permutation__round__n943 ), .ZN(_f_permutation__round__N3645 )
         );
  NOR2_X2 _f_permutation__round__U919  ( .A1(_f_permutation__round__c[933] ), 
        .A2(_f_permutation__round__n940 ), .ZN(_f_permutation__round__N3643 )
         );
  NOR2_X2 _f_permutation__round__U918  ( .A1(_f_permutation__round__c[934] ), 
        .A2(_f_permutation__round__n937 ), .ZN(_f_permutation__round__N3641 )
         );
  NOR2_X2 _f_permutation__round__U917  ( .A1(_f_permutation__round__c[935] ), 
        .A2(_f_permutation__round__n934 ), .ZN(_f_permutation__round__N3639 )
         );
  NOR2_X2 _f_permutation__round__U916  ( .A1(_f_permutation__round__c[936] ), 
        .A2(_f_permutation__round__n931 ), .ZN(_f_permutation__round__N3637 )
         );
  NOR2_X2 _f_permutation__round__U915  ( .A1(_f_permutation__round__c[937] ), 
        .A2(_f_permutation__round__n928 ), .ZN(_f_permutation__round__N3635 )
         );
  NOR2_X2 _f_permutation__round__U914  ( .A1(_f_permutation__round__c[938] ), 
        .A2(_f_permutation__round__n925 ), .ZN(_f_permutation__round__N3633 )
         );
  NOR2_X2 _f_permutation__round__U913  ( .A1(_f_permutation__round__c[939] ), 
        .A2(_f_permutation__round__n922 ), .ZN(_f_permutation__round__N3631 )
         );
  NOR2_X2 _f_permutation__round__U912  ( .A1(_f_permutation__round__c[940] ), 
        .A2(_f_permutation__round__n919 ), .ZN(_f_permutation__round__N3629 )
         );
  NOR2_X2 _f_permutation__round__U911  ( .A1(_f_permutation__round__c[941] ), 
        .A2(_f_permutation__round__n916 ), .ZN(_f_permutation__round__N3627 )
         );
  NOR2_X2 _f_permutation__round__U910  ( .A1(_f_permutation__round__c[942] ), 
        .A2(_f_permutation__round__n913 ), .ZN(_f_permutation__round__N3625 )
         );
  NOR2_X2 _f_permutation__round__U909  ( .A1(_f_permutation__round__c[943] ), 
        .A2(_f_permutation__round__n910 ), .ZN(_f_permutation__round__N3623 )
         );
  NOR2_X2 _f_permutation__round__U908  ( .A1(_f_permutation__round__c[944] ), 
        .A2(_f_permutation__round__n907 ), .ZN(_f_permutation__round__N3621 )
         );
  NOR2_X2 _f_permutation__round__U907  ( .A1(_f_permutation__round__c[945] ), 
        .A2(_f_permutation__round__n904 ), .ZN(_f_permutation__round__N3619 )
         );
  NOR2_X2 _f_permutation__round__U906  ( .A1(_f_permutation__round__c[946] ), 
        .A2(_f_permutation__round__n901 ), .ZN(_f_permutation__round__N3617 )
         );
  NOR2_X2 _f_permutation__round__U905  ( .A1(_f_permutation__round__c[947] ), 
        .A2(_f_permutation__round__n898 ), .ZN(_f_permutation__round__N3615 )
         );
  NOR2_X2 _f_permutation__round__U904  ( .A1(_f_permutation__round__c[948] ), 
        .A2(_f_permutation__round__n895 ), .ZN(_f_permutation__round__N3613 )
         );
  NOR2_X2 _f_permutation__round__U903  ( .A1(_f_permutation__round__c[949] ), 
        .A2(_f_permutation__round__n892 ), .ZN(_f_permutation__round__N3611 )
         );
  NOR2_X2 _f_permutation__round__U902  ( .A1(_f_permutation__round__c[950] ), 
        .A2(_f_permutation__round__n889 ), .ZN(_f_permutation__round__N3609 )
         );
  NOR2_X2 _f_permutation__round__U901  ( .A1(_f_permutation__round__c[951] ), 
        .A2(_f_permutation__round__n886 ), .ZN(_f_permutation__round__N3607 )
         );
  NOR2_X2 _f_permutation__round__U900  ( .A1(_f_permutation__round__c[952] ), 
        .A2(_f_permutation__round__n883 ), .ZN(_f_permutation__round__N3605 )
         );
  NOR2_X2 _f_permutation__round__U899  ( .A1(_f_permutation__round__c[953] ), 
        .A2(_f_permutation__round__n880 ), .ZN(_f_permutation__round__N3603 )
         );
  NOR2_X2 _f_permutation__round__U898  ( .A1(_f_permutation__round__c[954] ), 
        .A2(_f_permutation__round__n877 ), .ZN(_f_permutation__round__N3601 )
         );
  NOR2_X2 _f_permutation__round__U897  ( .A1(_f_permutation__round__c[955] ), 
        .A2(_f_permutation__round__n874 ), .ZN(_f_permutation__round__N3599 )
         );
  NOR2_X2 _f_permutation__round__U896  ( .A1(_f_permutation__round__c[956] ), 
        .A2(_f_permutation__round__n871 ), .ZN(_f_permutation__round__N3597 )
         );
  NOR2_X2 _f_permutation__round__U895  ( .A1(_f_permutation__round__c[957] ), 
        .A2(_f_permutation__round__n868 ), .ZN(_f_permutation__round__N3595 )
         );
  NOR2_X2 _f_permutation__round__U894  ( .A1(_f_permutation__round__c[958] ), 
        .A2(_f_permutation__round__n865 ), .ZN(_f_permutation__round__N3593 )
         );
  NOR2_X2 _f_permutation__round__U893  ( .A1(_f_permutation__round__c[959] ), 
        .A2(_f_permutation__round__n862 ), .ZN(_f_permutation__round__N3591 )
         );
  NOR2_X2 _f_permutation__round__U892  ( .A1(_f_permutation__round__c[896] ), 
        .A2(_f_permutation__round__n859 ), .ZN(_f_permutation__round__N3589 )
         );
  NOR2_X2 _f_permutation__round__U891  ( .A1(_f_permutation__round__c[897] ), 
        .A2(_f_permutation__round__n856 ), .ZN(_f_permutation__round__N3587 )
         );
  NOR2_X2 _f_permutation__round__U890  ( .A1(_f_permutation__round__c[898] ), 
        .A2(_f_permutation__round__n853 ), .ZN(_f_permutation__round__N3585 )
         );
  NOR2_X2 _f_permutation__round__U889  ( .A1(_f_permutation__round__c[1388] ), 
        .A2(_f_permutation__round__n467 ), .ZN(_f_permutation__round__N3327 )
         );
  NOR2_X2 _f_permutation__round__U888  ( .A1(_f_permutation__round__c[1389] ), 
        .A2(_f_permutation__round__n462 ), .ZN(_f_permutation__round__N3325 )
         );
  NOR2_X2 _f_permutation__round__U887  ( .A1(_f_permutation__round__c[1390] ), 
        .A2(_f_permutation__round__n457 ), .ZN(_f_permutation__round__N3323 )
         );
  NOR2_X2 _f_permutation__round__U886  ( .A1(_f_permutation__round__c[1391] ), 
        .A2(_f_permutation__round__n452 ), .ZN(_f_permutation__round__N3321 )
         );
  NOR2_X2 _f_permutation__round__U885  ( .A1(_f_permutation__round__c[1392] ), 
        .A2(_f_permutation__round__n767 ), .ZN(_f_permutation__round__N3319 )
         );
  NOR2_X2 _f_permutation__round__U884  ( .A1(_f_permutation__round__c[1393] ), 
        .A2(_f_permutation__round__n762 ), .ZN(_f_permutation__round__N3317 )
         );
  NOR2_X2 _f_permutation__round__U883  ( .A1(_f_permutation__round__c[1394] ), 
        .A2(_f_permutation__round__n757 ), .ZN(_f_permutation__round__N3315 )
         );
  NOR2_X2 _f_permutation__round__U882  ( .A1(_f_permutation__round__c[1395] ), 
        .A2(_f_permutation__round__n752 ), .ZN(_f_permutation__round__N3313 )
         );
  NOR2_X2 _f_permutation__round__U881  ( .A1(_f_permutation__round__c[1396] ), 
        .A2(_f_permutation__round__n747 ), .ZN(_f_permutation__round__N3311 )
         );
  NOR2_X2 _f_permutation__round__U880  ( .A1(_f_permutation__round__c[1397] ), 
        .A2(_f_permutation__round__n742 ), .ZN(_f_permutation__round__N3309 )
         );
  NOR2_X2 _f_permutation__round__U879  ( .A1(_f_permutation__round__c[1398] ), 
        .A2(_f_permutation__round__n737 ), .ZN(_f_permutation__round__N3307 )
         );
  NOR2_X2 _f_permutation__round__U878  ( .A1(_f_permutation__round__c[1399] ), 
        .A2(_f_permutation__round__n732 ), .ZN(_f_permutation__round__N3305 )
         );
  NOR2_X2 _f_permutation__round__U877  ( .A1(_f_permutation__round__c[1400] ), 
        .A2(_f_permutation__round__n727 ), .ZN(_f_permutation__round__N3303 )
         );
  NOR2_X2 _f_permutation__round__U876  ( .A1(_f_permutation__round__c[1401] ), 
        .A2(_f_permutation__round__n722 ), .ZN(_f_permutation__round__N3301 )
         );
  NOR2_X2 _f_permutation__round__U875  ( .A1(_f_permutation__round__c[1402] ), 
        .A2(_f_permutation__round__n717 ), .ZN(_f_permutation__round__N3299 )
         );
  NOR2_X2 _f_permutation__round__U874  ( .A1(_f_permutation__round__c[1403] ), 
        .A2(_f_permutation__round__n712 ), .ZN(_f_permutation__round__N3297 )
         );
  NOR2_X2 _f_permutation__round__U873  ( .A1(_f_permutation__round__c[1404] ), 
        .A2(_f_permutation__round__n707 ), .ZN(_f_permutation__round__N3295 )
         );
  NOR2_X2 _f_permutation__round__U872  ( .A1(_f_permutation__round__c[1405] ), 
        .A2(_f_permutation__round__n702 ), .ZN(_f_permutation__round__N3293 )
         );
  NOR2_X2 _f_permutation__round__U871  ( .A1(_f_permutation__round__c[1406] ), 
        .A2(_f_permutation__round__n697 ), .ZN(_f_permutation__round__N3291 )
         );
  NOR2_X2 _f_permutation__round__U870  ( .A1(_f_permutation__round__c[1407] ), 
        .A2(_f_permutation__round__n692 ), .ZN(_f_permutation__round__N3289 )
         );
  NOR2_X2 _f_permutation__round__U869  ( .A1(_f_permutation__round__c[1344] ), 
        .A2(_f_permutation__round__n687 ), .ZN(_f_permutation__round__N3287 )
         );
  NOR2_X2 _f_permutation__round__U868  ( .A1(_f_permutation__round__c[1345] ), 
        .A2(_f_permutation__round__n682 ), .ZN(_f_permutation__round__N3285 )
         );
  NOR2_X2 _f_permutation__round__U867  ( .A1(_f_permutation__round__c[1346] ), 
        .A2(_f_permutation__round__n677 ), .ZN(_f_permutation__round__N3283 )
         );
  NOR2_X2 _f_permutation__round__U866  ( .A1(_f_permutation__round__c[1347] ), 
        .A2(_f_permutation__round__n672 ), .ZN(_f_permutation__round__N3281 )
         );
  NOR2_X2 _f_permutation__round__U865  ( .A1(_f_permutation__round__c[1348] ), 
        .A2(_f_permutation__round__n667 ), .ZN(_f_permutation__round__N3279 )
         );
  NOR2_X2 _f_permutation__round__U864  ( .A1(_f_permutation__round__c[1349] ), 
        .A2(_f_permutation__round__n662 ), .ZN(_f_permutation__round__N3277 )
         );
  NOR2_X2 _f_permutation__round__U863  ( .A1(_f_permutation__round__c[1350] ), 
        .A2(_f_permutation__round__n657 ), .ZN(_f_permutation__round__N3275 )
         );
  NOR2_X2 _f_permutation__round__U862  ( .A1(_f_permutation__round__c[1351] ), 
        .A2(_f_permutation__round__n652 ), .ZN(_f_permutation__round__N3273 )
         );
  NOR2_X2 _f_permutation__round__U861  ( .A1(_f_permutation__round__c[1352] ), 
        .A2(_f_permutation__round__n647 ), .ZN(_f_permutation__round__N3271 )
         );
  NOR2_X2 _f_permutation__round__U860  ( .A1(_f_permutation__round__c[1353] ), 
        .A2(_f_permutation__round__n642 ), .ZN(_f_permutation__round__N3269 )
         );
  NOR2_X2 _f_permutation__round__U859  ( .A1(_f_permutation__round__c[1354] ), 
        .A2(_f_permutation__round__n637 ), .ZN(_f_permutation__round__N3267 )
         );
  NOR2_X2 _f_permutation__round__U858  ( .A1(_f_permutation__round__c[1355] ), 
        .A2(_f_permutation__round__n632 ), .ZN(_f_permutation__round__N3265 )
         );
  NOR2_X2 _f_permutation__round__U857  ( .A1(_f_permutation__round__c[1356] ), 
        .A2(_f_permutation__round__n627 ), .ZN(_f_permutation__round__N3263 )
         );
  NOR2_X2 _f_permutation__round__U856  ( .A1(_f_permutation__round__c[1357] ), 
        .A2(_f_permutation__round__n622 ), .ZN(_f_permutation__round__N3261 )
         );
  NOR2_X2 _f_permutation__round__U855  ( .A1(_f_permutation__round__c[1358] ), 
        .A2(_f_permutation__round__n617 ), .ZN(_f_permutation__round__N3259 )
         );
  NOR2_X2 _f_permutation__round__U854  ( .A1(_f_permutation__round__c[1359] ), 
        .A2(_f_permutation__round__n612 ), .ZN(_f_permutation__round__N3257 )
         );
  NOR2_X2 _f_permutation__round__U853  ( .A1(_f_permutation__round__c[1360] ), 
        .A2(_f_permutation__round__n607 ), .ZN(_f_permutation__round__N3255 )
         );
  NOR2_X2 _f_permutation__round__U852  ( .A1(_f_permutation__round__c[1361] ), 
        .A2(_f_permutation__round__n602 ), .ZN(_f_permutation__round__N3253 )
         );
  NOR2_X2 _f_permutation__round__U851  ( .A1(_f_permutation__round__c[1362] ), 
        .A2(_f_permutation__round__n597 ), .ZN(_f_permutation__round__N3251 )
         );
  NOR2_X2 _f_permutation__round__U850  ( .A1(_f_permutation__round__c[1363] ), 
        .A2(_f_permutation__round__n592 ), .ZN(_f_permutation__round__N3249 )
         );
  NOR2_X2 _f_permutation__round__U849  ( .A1(_f_permutation__round__c[1364] ), 
        .A2(_f_permutation__round__n587 ), .ZN(_f_permutation__round__N3247 )
         );
  NOR2_X2 _f_permutation__round__U848  ( .A1(_f_permutation__round__c[1365] ), 
        .A2(_f_permutation__round__n582 ), .ZN(_f_permutation__round__N3245 )
         );
  NOR2_X2 _f_permutation__round__U847  ( .A1(_f_permutation__round__c[1366] ), 
        .A2(_f_permutation__round__n577 ), .ZN(_f_permutation__round__N3243 )
         );
  NOR2_X2 _f_permutation__round__U846  ( .A1(_f_permutation__round__c[1367] ), 
        .A2(_f_permutation__round__n572 ), .ZN(_f_permutation__round__N3241 )
         );
  NOR2_X2 _f_permutation__round__U845  ( .A1(_f_permutation__round__c[1368] ), 
        .A2(_f_permutation__round__n567 ), .ZN(_f_permutation__round__N3239 )
         );
  NOR2_X2 _f_permutation__round__U844  ( .A1(_f_permutation__round__c[1369] ), 
        .A2(_f_permutation__round__n562 ), .ZN(_f_permutation__round__N3237 )
         );
  NOR2_X2 _f_permutation__round__U843  ( .A1(_f_permutation__round__c[1370] ), 
        .A2(_f_permutation__round__n557 ), .ZN(_f_permutation__round__N3235 )
         );
  NOR2_X2 _f_permutation__round__U842  ( .A1(_f_permutation__round__c[1371] ), 
        .A2(_f_permutation__round__n552 ), .ZN(_f_permutation__round__N3233 )
         );
  NOR2_X2 _f_permutation__round__U841  ( .A1(_f_permutation__round__c[1372] ), 
        .A2(_f_permutation__round__n547 ), .ZN(_f_permutation__round__N3231 )
         );
  NOR2_X2 _f_permutation__round__U840  ( .A1(_f_permutation__round__c[1373] ), 
        .A2(_f_permutation__round__n542 ), .ZN(_f_permutation__round__N3229 )
         );
  NOR2_X2 _f_permutation__round__U839  ( .A1(_f_permutation__round__c[1374] ), 
        .A2(_f_permutation__round__n537 ), .ZN(_f_permutation__round__N3227 )
         );
  NOR2_X2 _f_permutation__round__U838  ( .A1(_f_permutation__round__c[1375] ), 
        .A2(_f_permutation__round__n532 ), .ZN(_f_permutation__round__N3225 )
         );
  NOR2_X2 _f_permutation__round__U837  ( .A1(_f_permutation__round__c[1376] ), 
        .A2(_f_permutation__round__n527 ), .ZN(_f_permutation__round__N3223 )
         );
  NOR2_X2 _f_permutation__round__U836  ( .A1(_f_permutation__round__c[1377] ), 
        .A2(_f_permutation__round__n522 ), .ZN(_f_permutation__round__N3221 )
         );
  NOR2_X2 _f_permutation__round__U835  ( .A1(_f_permutation__round__c[1378] ), 
        .A2(_f_permutation__round__n517 ), .ZN(_f_permutation__round__N3219 )
         );
  NOR2_X2 _f_permutation__round__U834  ( .A1(_f_permutation__round__c[1379] ), 
        .A2(_f_permutation__round__n512 ), .ZN(_f_permutation__round__N3217 )
         );
  NOR2_X2 _f_permutation__round__U833  ( .A1(_f_permutation__round__c[1380] ), 
        .A2(_f_permutation__round__n507 ), .ZN(_f_permutation__round__N3215 )
         );
  NOR2_X2 _f_permutation__round__U768  ( .A1(_f_permutation__round__c[1381] ), 
        .A2(_f_permutation__round__n502 ), .ZN(_f_permutation__round__N3213 )
         );
  NOR2_X2 _f_permutation__round__U767  ( .A1(_f_permutation__round__c[1382] ), 
        .A2(_f_permutation__round__n497 ), .ZN(_f_permutation__round__N3211 )
         );
  NOR2_X2 _f_permutation__round__U766  ( .A1(_f_permutation__round__c[1383] ), 
        .A2(_f_permutation__round__n492 ), .ZN(_f_permutation__round__N3209 )
         );
  NOR2_X2 _f_permutation__round__U765  ( .A1(_f_permutation__round__c[1384] ), 
        .A2(_f_permutation__round__n487 ), .ZN(_f_permutation__round__N3207 )
         );
  NOR2_X2 _f_permutation__round__U764  ( .A1(_f_permutation__round__c[1385] ), 
        .A2(_f_permutation__round__n482 ), .ZN(_f_permutation__round__N3205 )
         );
  NOR2_X2 _f_permutation__round__U763  ( .A1(_f_permutation__round__c[1386] ), 
        .A2(_f_permutation__round__n477 ), .ZN(_f_permutation__round__N3203 )
         );
  NOR2_X2 _f_permutation__round__U762  ( .A1(_f_permutation__round__c[1387] ), 
        .A2(_f_permutation__round__n472 ), .ZN(_f_permutation__round__N3201 )
         );
  NOR2_X2 _f_permutation__round__U761  ( .A1(_f_permutation__round__c[1586] ), 
        .A2(_f_permutation__round__n448 ), .ZN(_f_permutation__round__N3071 )
         );
  NOR2_X2 _f_permutation__round__U760  ( .A1(_f_permutation__round__c[1587] ), 
        .A2(_f_permutation__round__n441 ), .ZN(_f_permutation__round__N3069 )
         );
  NOR2_X2 _f_permutation__round__U759  ( .A1(_f_permutation__round__c[1588] ), 
        .A2(_f_permutation__round__n434 ), .ZN(_f_permutation__round__N3067 )
         );
  NOR2_X2 _f_permutation__round__U758  ( .A1(_f_permutation__round__c[1589] ), 
        .A2(_f_permutation__round__n427 ), .ZN(_f_permutation__round__N3065 )
         );
  NOR2_X2 _f_permutation__round__U757  ( .A1(_f_permutation__round__c[1590] ), 
        .A2(_f_permutation__round__n420 ), .ZN(_f_permutation__round__N3063 )
         );
  NOR2_X2 _f_permutation__round__U756  ( .A1(_f_permutation__round__c[1591] ), 
        .A2(_f_permutation__round__n413 ), .ZN(_f_permutation__round__N3061 )
         );
  NOR2_X2 _f_permutation__round__U755  ( .A1(_f_permutation__round__c[1592] ), 
        .A2(_f_permutation__round__n406 ), .ZN(_f_permutation__round__N3059 )
         );
  NOR2_X2 _f_permutation__round__U754  ( .A1(_f_permutation__round__c[1593] ), 
        .A2(_f_permutation__round__n399 ), .ZN(_f_permutation__round__N3057 )
         );
  NOR2_X2 _f_permutation__round__U753  ( .A1(_f_permutation__round__c[1594] ), 
        .A2(_f_permutation__round__n392 ), .ZN(_f_permutation__round__N3055 )
         );
  NOR2_X2 _f_permutation__round__U752  ( .A1(_f_permutation__round__c[1595] ), 
        .A2(_f_permutation__round__n385 ), .ZN(_f_permutation__round__N3053 )
         );
  NOR2_X2 _f_permutation__round__U751  ( .A1(_f_permutation__round__c[1596] ), 
        .A2(_f_permutation__round__n378 ), .ZN(_f_permutation__round__N3051 )
         );
  NOR2_X2 _f_permutation__round__U750  ( .A1(_f_permutation__round__c[1597] ), 
        .A2(_f_permutation__round__n371 ), .ZN(_f_permutation__round__N3049 )
         );
  NOR2_X2 _f_permutation__round__U749  ( .A1(_f_permutation__round__c[1598] ), 
        .A2(_f_permutation__round__n364 ), .ZN(_f_permutation__round__N3047 )
         );
  NOR2_X2 _f_permutation__round__U748  ( .A1(_f_permutation__round__c[1599] ), 
        .A2(_f_permutation__round__n357 ), .ZN(_f_permutation__round__N3045 )
         );
  NOR2_X2 _f_permutation__round__U747  ( .A1(_f_permutation__round__c[1536] ), 
        .A2(_f_permutation__round__n350 ), .ZN(_f_permutation__round__N3043 )
         );
  NOR2_X2 _f_permutation__round__U746  ( .A1(_f_permutation__round__c[1537] ), 
        .A2(_f_permutation__round__n343 ), .ZN(_f_permutation__round__N3041 )
         );
  NOR2_X2 _f_permutation__round__U745  ( .A1(_f_permutation__round__c[1538] ), 
        .A2(_f_permutation__round__n336 ), .ZN(_f_permutation__round__N3039 )
         );
  NOR2_X2 _f_permutation__round__U744  ( .A1(_f_permutation__round__c[1539] ), 
        .A2(_f_permutation__round__n329 ), .ZN(_f_permutation__round__N3037 )
         );
  NOR2_X2 _f_permutation__round__U743  ( .A1(_f_permutation__round__c[1540] ), 
        .A2(_f_permutation__round__n322 ), .ZN(_f_permutation__round__N3035 )
         );
  NOR2_X2 _f_permutation__round__U742  ( .A1(_f_permutation__round__c[1541] ), 
        .A2(_f_permutation__round__n315 ), .ZN(_f_permutation__round__N3033 )
         );
  NOR2_X2 _f_permutation__round__U741  ( .A1(_f_permutation__round__c[1542] ), 
        .A2(_f_permutation__round__n308 ), .ZN(_f_permutation__round__N3031 )
         );
  NOR2_X2 _f_permutation__round__U740  ( .A1(_f_permutation__round__c[1543] ), 
        .A2(_f_permutation__round__n301 ), .ZN(_f_permutation__round__N3029 )
         );
  NOR2_X2 _f_permutation__round__U739  ( .A1(_f_permutation__round__c[1544] ), 
        .A2(_f_permutation__round__n294 ), .ZN(_f_permutation__round__N3027 )
         );
  NOR2_X2 _f_permutation__round__U738  ( .A1(_f_permutation__round__c[1545] ), 
        .A2(_f_permutation__round__n287 ), .ZN(_f_permutation__round__N3025 )
         );
  NOR2_X2 _f_permutation__round__U737  ( .A1(_f_permutation__round__c[1546] ), 
        .A2(_f_permutation__round__n280 ), .ZN(_f_permutation__round__N3023 )
         );
  NOR2_X2 _f_permutation__round__U736  ( .A1(_f_permutation__round__c[1547] ), 
        .A2(_f_permutation__round__n273 ), .ZN(_f_permutation__round__N3021 )
         );
  NOR2_X2 _f_permutation__round__U735  ( .A1(_f_permutation__round__c[1548] ), 
        .A2(_f_permutation__round__n266 ), .ZN(_f_permutation__round__N3019 )
         );
  NOR2_X2 _f_permutation__round__U734  ( .A1(_f_permutation__round__c[1549] ), 
        .A2(_f_permutation__round__n259 ), .ZN(_f_permutation__round__N3017 )
         );
  NOR2_X2 _f_permutation__round__U733  ( .A1(_f_permutation__round__c[1550] ), 
        .A2(_f_permutation__round__n252 ), .ZN(_f_permutation__round__N3015 )
         );
  NOR2_X2 _f_permutation__round__U732  ( .A1(_f_permutation__round__c[1551] ), 
        .A2(_f_permutation__round__n245 ), .ZN(_f_permutation__round__N3013 )
         );
  NOR2_X2 _f_permutation__round__U731  ( .A1(_f_permutation__round__c[1552] ), 
        .A2(_f_permutation__round__n238 ), .ZN(_f_permutation__round__N3011 )
         );
  NOR2_X2 _f_permutation__round__U730  ( .A1(_f_permutation__round__c[1553] ), 
        .A2(_f_permutation__round__n231 ), .ZN(_f_permutation__round__N3009 )
         );
  NOR2_X2 _f_permutation__round__U729  ( .A1(_f_permutation__round__c[1554] ), 
        .A2(_f_permutation__round__n224 ), .ZN(_f_permutation__round__N3007 )
         );
  NOR2_X2 _f_permutation__round__U728  ( .A1(_f_permutation__round__c[1555] ), 
        .A2(_f_permutation__round__n217 ), .ZN(_f_permutation__round__N3005 )
         );
  NOR2_X2 _f_permutation__round__U727  ( .A1(_f_permutation__round__c[1556] ), 
        .A2(_f_permutation__round__n210 ), .ZN(_f_permutation__round__N3003 )
         );
  NOR2_X2 _f_permutation__round__U726  ( .A1(_f_permutation__round__c[1557] ), 
        .A2(_f_permutation__round__n203 ), .ZN(_f_permutation__round__N3001 )
         );
  NOR2_X2 _f_permutation__round__U725  ( .A1(_f_permutation__round__c[1558] ), 
        .A2(_f_permutation__round__n196 ), .ZN(_f_permutation__round__N2999 )
         );
  NOR2_X2 _f_permutation__round__U724  ( .A1(_f_permutation__round__c[1559] ), 
        .A2(_f_permutation__round__n189 ), .ZN(_f_permutation__round__N2997 )
         );
  NOR2_X2 _f_permutation__round__U723  ( .A1(_f_permutation__round__c[1560] ), 
        .A2(_f_permutation__round__n182 ), .ZN(_f_permutation__round__N2995 )
         );
  NOR2_X2 _f_permutation__round__U722  ( .A1(_f_permutation__round__c[1561] ), 
        .A2(_f_permutation__round__n175 ), .ZN(_f_permutation__round__N2993 )
         );
  NOR2_X2 _f_permutation__round__U721  ( .A1(_f_permutation__round__c[1562] ), 
        .A2(_f_permutation__round__n168 ), .ZN(_f_permutation__round__N2991 )
         );
  NOR2_X2 _f_permutation__round__U720  ( .A1(_f_permutation__round__c[1563] ), 
        .A2(_f_permutation__round__n161 ), .ZN(_f_permutation__round__N2989 )
         );
  NOR2_X2 _f_permutation__round__U719  ( .A1(_f_permutation__round__c[1564] ), 
        .A2(_f_permutation__round__n154 ), .ZN(_f_permutation__round__N2987 )
         );
  NOR2_X2 _f_permutation__round__U718  ( .A1(_f_permutation__round__c[1565] ), 
        .A2(_f_permutation__round__n147 ), .ZN(_f_permutation__round__N2985 )
         );
  NOR2_X2 _f_permutation__round__U717  ( .A1(_f_permutation__round__c[1566] ), 
        .A2(_f_permutation__round__n140 ), .ZN(_f_permutation__round__N2983 )
         );
  NOR2_X2 _f_permutation__round__U716  ( .A1(_f_permutation__round__c[1567] ), 
        .A2(_f_permutation__round__n133 ), .ZN(_f_permutation__round__N2981 )
         );
  NOR2_X2 _f_permutation__round__U715  ( .A1(_f_permutation__round__c[1568] ), 
        .A2(_f_permutation__round__n126 ), .ZN(_f_permutation__round__N2979 )
         );
  NOR2_X2 _f_permutation__round__U714  ( .A1(_f_permutation__round__c[1569] ), 
        .A2(_f_permutation__round__n119 ), .ZN(_f_permutation__round__N2977 )
         );
  NOR2_X2 _f_permutation__round__U713  ( .A1(_f_permutation__round__c[1570] ), 
        .A2(_f_permutation__round__n112 ), .ZN(_f_permutation__round__N2975 )
         );
  NOR2_X2 _f_permutation__round__U712  ( .A1(_f_permutation__round__c[1571] ), 
        .A2(_f_permutation__round__n105 ), .ZN(_f_permutation__round__N2973 )
         );
  NOR2_X2 _f_permutation__round__U711  ( .A1(_f_permutation__round__c[1572] ), 
        .A2(_f_permutation__round__n98 ), .ZN(_f_permutation__round__N2971 )
         );
  NOR2_X2 _f_permutation__round__U710  ( .A1(_f_permutation__round__c[1573] ), 
        .A2(_f_permutation__round__n91 ), .ZN(_f_permutation__round__N2969 )
         );
  NOR2_X2 _f_permutation__round__U709  ( .A1(_f_permutation__round__c[1574] ), 
        .A2(_f_permutation__round__n84 ), .ZN(_f_permutation__round__N2967 )
         );
  NOR2_X2 _f_permutation__round__U708  ( .A1(_f_permutation__round__c[1575] ), 
        .A2(_f_permutation__round__n77 ), .ZN(_f_permutation__round__N2965 )
         );
  NOR2_X2 _f_permutation__round__U707  ( .A1(_f_permutation__round__c[1576] ), 
        .A2(_f_permutation__round__n70 ), .ZN(_f_permutation__round__N2963 )
         );
  NOR2_X2 _f_permutation__round__U706  ( .A1(_f_permutation__round__c[1577] ), 
        .A2(_f_permutation__round__n63 ), .ZN(_f_permutation__round__N2961 )
         );
  NOR2_X2 _f_permutation__round__U705  ( .A1(_f_permutation__round__c[1578] ), 
        .A2(_f_permutation__round__n56 ), .ZN(_f_permutation__round__N2959 )
         );
  NOR2_X2 _f_permutation__round__U640  ( .A1(_f_permutation__round__c[1579] ), 
        .A2(_f_permutation__round__n49 ), .ZN(_f_permutation__round__N2957 )
         );
  NOR2_X2 _f_permutation__round__U639  ( .A1(_f_permutation__round__c[1580] ), 
        .A2(_f_permutation__round__n42 ), .ZN(_f_permutation__round__N2955 )
         );
  NOR2_X2 _f_permutation__round__U638  ( .A1(_f_permutation__round__c[1581] ), 
        .A2(_f_permutation__round__n35 ), .ZN(_f_permutation__round__N2953 )
         );
  NOR2_X2 _f_permutation__round__U637  ( .A1(_f_permutation__round__c[1582] ), 
        .A2(_f_permutation__round__n28 ), .ZN(_f_permutation__round__N2951 )
         );
  NOR2_X2 _f_permutation__round__U636  ( .A1(_f_permutation__round__c[1583] ), 
        .A2(_f_permutation__round__n21 ), .ZN(_f_permutation__round__N2949 )
         );
  NOR2_X2 _f_permutation__round__U635  ( .A1(_f_permutation__round__c[1584] ), 
        .A2(_f_permutation__round__n14 ), .ZN(_f_permutation__round__N2947 )
         );
  NOR2_X2 _f_permutation__round__U634  ( .A1(_f_permutation__round__c[1585] ), 
        .A2(_f_permutation__round__n7 ), .ZN(_f_permutation__round__N2945 ) );
  NOR2_X2 _f_permutation__round__U633  ( .A1(_f_permutation__round__c[406] ), 
        .A2(_f_permutation__round__n650 ), .ZN(_f_permutation__round__N2683 )
         );
  NOR2_X2 _f_permutation__round__U632  ( .A1(_f_permutation__round__c[408] ), 
        .A2(_f_permutation__round__n640 ), .ZN(_f_permutation__round__N2679 )
         );
  NOR2_X2 _f_permutation__round__U631  ( .A1(_f_permutation__round__c[409] ), 
        .A2(_f_permutation__round__n635 ), .ZN(_f_permutation__round__N2677 )
         );
  NOR2_X2 _f_permutation__round__U630  ( .A1(_f_permutation__round__c[410] ), 
        .A2(_f_permutation__round__n630 ), .ZN(_f_permutation__round__N2675 )
         );
  NOR2_X2 _f_permutation__round__U629  ( .A1(_f_permutation__round__c[412] ), 
        .A2(_f_permutation__round__n620 ), .ZN(_f_permutation__round__N2671 )
         );
  NOR2_X2 _f_permutation__round__U628  ( .A1(_f_permutation__round__c[413] ), 
        .A2(_f_permutation__round__n615 ), .ZN(_f_permutation__round__N2669 )
         );
  NOR2_X2 _f_permutation__round__U627  ( .A1(_f_permutation__round__c[414] ), 
        .A2(_f_permutation__round__n610 ), .ZN(_f_permutation__round__N2667 )
         );
  NOR2_X2 _f_permutation__round__U626  ( .A1(_f_permutation__round__c[415] ), 
        .A2(_f_permutation__round__n605 ), .ZN(_f_permutation__round__N2665 )
         );
  NOR2_X2 _f_permutation__round__U625  ( .A1(_f_permutation__round__c[416] ), 
        .A2(_f_permutation__round__n600 ), .ZN(_f_permutation__round__N2663 )
         );
  NOR2_X2 _f_permutation__round__U624  ( .A1(_f_permutation__round__c[417] ), 
        .A2(_f_permutation__round__n595 ), .ZN(_f_permutation__round__N2661 )
         );
  NOR2_X2 _f_permutation__round__U623  ( .A1(_f_permutation__round__c[418] ), 
        .A2(_f_permutation__round__n590 ), .ZN(_f_permutation__round__N2659 )
         );
  NOR2_X2 _f_permutation__round__U622  ( .A1(_f_permutation__round__c[420] ), 
        .A2(_f_permutation__round__n580 ), .ZN(_f_permutation__round__N2655 )
         );
  NOR2_X2 _f_permutation__round__U621  ( .A1(_f_permutation__round__c[421] ), 
        .A2(_f_permutation__round__n575 ), .ZN(_f_permutation__round__N2653 )
         );
  NOR2_X2 _f_permutation__round__U620  ( .A1(_f_permutation__round__c[422] ), 
        .A2(_f_permutation__round__n570 ), .ZN(_f_permutation__round__N2651 )
         );
  NOR2_X2 _f_permutation__round__U619  ( .A1(_f_permutation__round__c[423] ), 
        .A2(_f_permutation__round__n565 ), .ZN(_f_permutation__round__N2649 )
         );
  NOR2_X2 _f_permutation__round__U618  ( .A1(_f_permutation__round__c[424] ), 
        .A2(_f_permutation__round__n560 ), .ZN(_f_permutation__round__N2647 )
         );
  NOR2_X2 _f_permutation__round__U617  ( .A1(_f_permutation__round__c[425] ), 
        .A2(_f_permutation__round__n555 ), .ZN(_f_permutation__round__N2645 )
         );
  NOR2_X2 _f_permutation__round__U616  ( .A1(_f_permutation__round__c[426] ), 
        .A2(_f_permutation__round__n550 ), .ZN(_f_permutation__round__N2643 )
         );
  NOR2_X2 _f_permutation__round__U615  ( .A1(_f_permutation__round__c[427] ), 
        .A2(_f_permutation__round__n545 ), .ZN(_f_permutation__round__N2641 )
         );
  NOR2_X2 _f_permutation__round__U614  ( .A1(_f_permutation__round__c[428] ), 
        .A2(_f_permutation__round__n540 ), .ZN(_f_permutation__round__N2639 )
         );
  NOR2_X2 _f_permutation__round__U613  ( .A1(_f_permutation__round__c[429] ), 
        .A2(_f_permutation__round__n535 ), .ZN(_f_permutation__round__N2637 )
         );
  NOR2_X2 _f_permutation__round__U612  ( .A1(_f_permutation__round__c[430] ), 
        .A2(_f_permutation__round__n530 ), .ZN(_f_permutation__round__N2635 )
         );
  NOR2_X2 _f_permutation__round__U611  ( .A1(_f_permutation__round__c[431] ), 
        .A2(_f_permutation__round__n525 ), .ZN(_f_permutation__round__N2633 )
         );
  NOR2_X2 _f_permutation__round__U610  ( .A1(_f_permutation__round__c[432] ), 
        .A2(_f_permutation__round__n520 ), .ZN(_f_permutation__round__N2631 )
         );
  NOR2_X2 _f_permutation__round__U609  ( .A1(_f_permutation__round__c[433] ), 
        .A2(_f_permutation__round__n515 ), .ZN(_f_permutation__round__N2629 )
         );
  NOR2_X2 _f_permutation__round__U608  ( .A1(_f_permutation__round__c[434] ), 
        .A2(_f_permutation__round__n510 ), .ZN(_f_permutation__round__N2627 )
         );
  NOR2_X2 _f_permutation__round__U607  ( .A1(_f_permutation__round__c[436] ), 
        .A2(_f_permutation__round__n500 ), .ZN(_f_permutation__round__N2623 )
         );
  NOR2_X2 _f_permutation__round__U606  ( .A1(_f_permutation__round__c[437] ), 
        .A2(_f_permutation__round__n495 ), .ZN(_f_permutation__round__N2621 )
         );
  NOR2_X2 _f_permutation__round__U605  ( .A1(_f_permutation__round__c[438] ), 
        .A2(_f_permutation__round__n490 ), .ZN(_f_permutation__round__N2619 )
         );
  NOR2_X2 _f_permutation__round__U604  ( .A1(_f_permutation__round__c[439] ), 
        .A2(_f_permutation__round__n485 ), .ZN(_f_permutation__round__N2617 )
         );
  NOR2_X2 _f_permutation__round__U603  ( .A1(_f_permutation__round__c[440] ), 
        .A2(_f_permutation__round__n480 ), .ZN(_f_permutation__round__N2615 )
         );
  NOR2_X2 _f_permutation__round__U602  ( .A1(_f_permutation__round__c[441] ), 
        .A2(_f_permutation__round__n475 ), .ZN(_f_permutation__round__N2613 )
         );
  NOR2_X2 _f_permutation__round__U601  ( .A1(_f_permutation__round__c[442] ), 
        .A2(_f_permutation__round__n470 ), .ZN(_f_permutation__round__N2611 )
         );
  NOR2_X2 _f_permutation__round__U600  ( .A1(_f_permutation__round__c[443] ), 
        .A2(_f_permutation__round__n465 ), .ZN(_f_permutation__round__N2609 )
         );
  NOR2_X2 _f_permutation__round__U599  ( .A1(_f_permutation__round__c[444] ), 
        .A2(_f_permutation__round__n460 ), .ZN(_f_permutation__round__N2607 )
         );
  NOR2_X2 _f_permutation__round__U598  ( .A1(_f_permutation__round__c[445] ), 
        .A2(_f_permutation__round__n455 ), .ZN(_f_permutation__round__N2605 )
         );
  NOR2_X2 _f_permutation__round__U597  ( .A1(_f_permutation__round__c[446] ), 
        .A2(_f_permutation__round__n450 ), .ZN(_f_permutation__round__N2603 )
         );
  NOR2_X2 _f_permutation__round__U596  ( .A1(_f_permutation__round__c[447] ), 
        .A2(_f_permutation__round__n765 ), .ZN(_f_permutation__round__N2601 )
         );
  NOR2_X2 _f_permutation__round__U595  ( .A1(_f_permutation__round__c[384] ), 
        .A2(_f_permutation__round__n760 ), .ZN(_f_permutation__round__N2599 )
         );
  NOR2_X2 _f_permutation__round__U594  ( .A1(_f_permutation__round__c[385] ), 
        .A2(_f_permutation__round__n755 ), .ZN(_f_permutation__round__N2597 )
         );
  NOR2_X2 _f_permutation__round__U593  ( .A1(_f_permutation__round__c[386] ), 
        .A2(_f_permutation__round__n750 ), .ZN(_f_permutation__round__N2595 )
         );
  NOR2_X2 _f_permutation__round__U592  ( .A1(_f_permutation__round__c[387] ), 
        .A2(_f_permutation__round__n745 ), .ZN(_f_permutation__round__N2593 )
         );
  NOR2_X2 _f_permutation__round__U591  ( .A1(_f_permutation__round__c[388] ), 
        .A2(_f_permutation__round__n740 ), .ZN(_f_permutation__round__N2591 )
         );
  NOR2_X2 _f_permutation__round__U590  ( .A1(_f_permutation__round__c[389] ), 
        .A2(_f_permutation__round__n735 ), .ZN(_f_permutation__round__N2589 )
         );
  NOR2_X2 _f_permutation__round__U589  ( .A1(_f_permutation__round__c[390] ), 
        .A2(_f_permutation__round__n730 ), .ZN(_f_permutation__round__N2587 )
         );
  NOR2_X2 _f_permutation__round__U588  ( .A1(_f_permutation__round__c[391] ), 
        .A2(_f_permutation__round__n725 ), .ZN(_f_permutation__round__N2585 )
         );
  NOR2_X2 _f_permutation__round__U587  ( .A1(_f_permutation__round__c[392] ), 
        .A2(_f_permutation__round__n720 ), .ZN(_f_permutation__round__N2583 )
         );
  NOR2_X2 _f_permutation__round__U586  ( .A1(_f_permutation__round__c[393] ), 
        .A2(_f_permutation__round__n715 ), .ZN(_f_permutation__round__N2581 )
         );
  NOR2_X2 _f_permutation__round__U585  ( .A1(_f_permutation__round__c[394] ), 
        .A2(_f_permutation__round__n710 ), .ZN(_f_permutation__round__N2579 )
         );
  NOR2_X2 _f_permutation__round__U584  ( .A1(_f_permutation__round__c[395] ), 
        .A2(_f_permutation__round__n705 ), .ZN(_f_permutation__round__N2577 )
         );
  NOR2_X2 _f_permutation__round__U583  ( .A1(_f_permutation__round__c[396] ), 
        .A2(_f_permutation__round__n700 ), .ZN(_f_permutation__round__N2575 )
         );
  NOR2_X2 _f_permutation__round__U582  ( .A1(_f_permutation__round__c[397] ), 
        .A2(_f_permutation__round__n695 ), .ZN(_f_permutation__round__N2573 )
         );
  NOR2_X2 _f_permutation__round__U581  ( .A1(_f_permutation__round__c[398] ), 
        .A2(_f_permutation__round__n690 ), .ZN(_f_permutation__round__N2571 )
         );
  NOR2_X2 _f_permutation__round__U580  ( .A1(_f_permutation__round__c[399] ), 
        .A2(_f_permutation__round__n685 ), .ZN(_f_permutation__round__N2569 )
         );
  NOR2_X2 _f_permutation__round__U579  ( .A1(_f_permutation__round__c[400] ), 
        .A2(_f_permutation__round__n680 ), .ZN(_f_permutation__round__N2567 )
         );
  NOR2_X2 _f_permutation__round__U578  ( .A1(_f_permutation__round__c[401] ), 
        .A2(_f_permutation__round__n675 ), .ZN(_f_permutation__round__N2565 )
         );
  NOR2_X2 _f_permutation__round__U577  ( .A1(_f_permutation__round__c[402] ), 
        .A2(_f_permutation__round__n670 ), .ZN(_f_permutation__round__N2563 )
         );
  NOR2_X2 _f_permutation__round__U576  ( .A1(_f_permutation__round__c[1433] ), 
        .A2(_f_permutation__round__n658 ), .ZN(_f_permutation__round__N5375 )
         );
  NOR2_X2 _f_permutation__round__U575  ( .A1(_f_permutation__round__c[1434] ), 
        .A2(_f_permutation__round__n653 ), .ZN(_f_permutation__round__N5373 )
         );
  NOR2_X2 _f_permutation__round__U574  ( .A1(_f_permutation__round__c[1435] ), 
        .A2(_f_permutation__round__n648 ), .ZN(_f_permutation__round__N5371 )
         );
  NOR2_X2 _f_permutation__round__U573  ( .A1(_f_permutation__round__c[1436] ), 
        .A2(_f_permutation__round__n643 ), .ZN(_f_permutation__round__N5369 )
         );
  NOR2_X2 _f_permutation__round__U572  ( .A1(_f_permutation__round__c[1437] ), 
        .A2(_f_permutation__round__n638 ), .ZN(_f_permutation__round__N5367 )
         );
  NOR2_X2 _f_permutation__round__U571  ( .A1(_f_permutation__round__c[1438] ), 
        .A2(_f_permutation__round__n633 ), .ZN(_f_permutation__round__N5365 )
         );
  NOR2_X2 _f_permutation__round__U570  ( .A1(_f_permutation__round__c[1439] ), 
        .A2(_f_permutation__round__n628 ), .ZN(_f_permutation__round__N5363 )
         );
  NOR2_X2 _f_permutation__round__U569  ( .A1(_f_permutation__round__c[1440] ), 
        .A2(_f_permutation__round__n623 ), .ZN(_f_permutation__round__N5361 )
         );
  NOR2_X2 _f_permutation__round__U568  ( .A1(_f_permutation__round__c[1441] ), 
        .A2(_f_permutation__round__n618 ), .ZN(_f_permutation__round__N5359 )
         );
  NOR2_X2 _f_permutation__round__U567  ( .A1(_f_permutation__round__c[1442] ), 
        .A2(_f_permutation__round__n613 ), .ZN(_f_permutation__round__N5357 )
         );
  NOR2_X2 _f_permutation__round__U566  ( .A1(_f_permutation__round__c[1443] ), 
        .A2(_f_permutation__round__n608 ), .ZN(_f_permutation__round__N5355 )
         );
  NOR2_X2 _f_permutation__round__U565  ( .A1(_f_permutation__round__c[1444] ), 
        .A2(_f_permutation__round__n603 ), .ZN(_f_permutation__round__N5353 )
         );
  NOR2_X2 _f_permutation__round__U564  ( .A1(_f_permutation__round__c[1445] ), 
        .A2(_f_permutation__round__n598 ), .ZN(_f_permutation__round__N5351 )
         );
  NOR2_X2 _f_permutation__round__U563  ( .A1(_f_permutation__round__c[1446] ), 
        .A2(_f_permutation__round__n593 ), .ZN(_f_permutation__round__N5349 )
         );
  NOR2_X2 _f_permutation__round__U562  ( .A1(_f_permutation__round__c[1447] ), 
        .A2(_f_permutation__round__n588 ), .ZN(_f_permutation__round__N5347 )
         );
  NOR2_X2 _f_permutation__round__U561  ( .A1(_f_permutation__round__c[1448] ), 
        .A2(_f_permutation__round__n583 ), .ZN(_f_permutation__round__N5345 )
         );
  NOR2_X2 _f_permutation__round__U560  ( .A1(_f_permutation__round__c[1449] ), 
        .A2(_f_permutation__round__n578 ), .ZN(_f_permutation__round__N5343 )
         );
  NOR2_X2 _f_permutation__round__U559  ( .A1(_f_permutation__round__c[1450] ), 
        .A2(_f_permutation__round__n573 ), .ZN(_f_permutation__round__N5341 )
         );
  NOR2_X2 _f_permutation__round__U558  ( .A1(_f_permutation__round__c[1451] ), 
        .A2(_f_permutation__round__n568 ), .ZN(_f_permutation__round__N5339 )
         );
  NOR2_X2 _f_permutation__round__U557  ( .A1(_f_permutation__round__c[1452] ), 
        .A2(_f_permutation__round__n563 ), .ZN(_f_permutation__round__N5337 )
         );
  NOR2_X2 _f_permutation__round__U556  ( .A1(_f_permutation__round__c[1453] ), 
        .A2(_f_permutation__round__n558 ), .ZN(_f_permutation__round__N5335 )
         );
  NOR2_X2 _f_permutation__round__U555  ( .A1(_f_permutation__round__c[1454] ), 
        .A2(_f_permutation__round__n553 ), .ZN(_f_permutation__round__N5333 )
         );
  NOR2_X2 _f_permutation__round__U554  ( .A1(_f_permutation__round__c[1455] ), 
        .A2(_f_permutation__round__n548 ), .ZN(_f_permutation__round__N5331 )
         );
  NOR2_X2 _f_permutation__round__U553  ( .A1(_f_permutation__round__c[1456] ), 
        .A2(_f_permutation__round__n543 ), .ZN(_f_permutation__round__N5329 )
         );
  NOR2_X2 _f_permutation__round__U552  ( .A1(_f_permutation__round__c[1457] ), 
        .A2(_f_permutation__round__n538 ), .ZN(_f_permutation__round__N5327 )
         );
  NOR2_X2 _f_permutation__round__U551  ( .A1(_f_permutation__round__c[1458] ), 
        .A2(_f_permutation__round__n533 ), .ZN(_f_permutation__round__N5325 )
         );
  NOR2_X2 _f_permutation__round__U550  ( .A1(_f_permutation__round__c[1459] ), 
        .A2(_f_permutation__round__n528 ), .ZN(_f_permutation__round__N5323 )
         );
  NOR2_X2 _f_permutation__round__U549  ( .A1(_f_permutation__round__c[1460] ), 
        .A2(_f_permutation__round__n523 ), .ZN(_f_permutation__round__N5321 )
         );
  NOR2_X2 _f_permutation__round__U548  ( .A1(_f_permutation__round__c[1461] ), 
        .A2(_f_permutation__round__n518 ), .ZN(_f_permutation__round__N5319 )
         );
  NOR2_X2 _f_permutation__round__U547  ( .A1(_f_permutation__round__c[1462] ), 
        .A2(_f_permutation__round__n513 ), .ZN(_f_permutation__round__N5317 )
         );
  NOR2_X2 _f_permutation__round__U546  ( .A1(_f_permutation__round__c[1463] ), 
        .A2(_f_permutation__round__n508 ), .ZN(_f_permutation__round__N5315 )
         );
  NOR2_X2 _f_permutation__round__U545  ( .A1(_f_permutation__round__c[1464] ), 
        .A2(_f_permutation__round__n503 ), .ZN(_f_permutation__round__N5313 )
         );
  NOR2_X2 _f_permutation__round__U544  ( .A1(_f_permutation__round__c[1465] ), 
        .A2(_f_permutation__round__n498 ), .ZN(_f_permutation__round__N5311 )
         );
  NOR2_X2 _f_permutation__round__U543  ( .A1(_f_permutation__round__c[1466] ), 
        .A2(_f_permutation__round__n493 ), .ZN(_f_permutation__round__N5309 )
         );
  NOR2_X2 _f_permutation__round__U542  ( .A1(_f_permutation__round__c[1467] ), 
        .A2(_f_permutation__round__n488 ), .ZN(_f_permutation__round__N5307 )
         );
  NOR2_X2 _f_permutation__round__U541  ( .A1(_f_permutation__round__c[1468] ), 
        .A2(_f_permutation__round__n483 ), .ZN(_f_permutation__round__N5305 )
         );
  NOR2_X2 _f_permutation__round__U540  ( .A1(_f_permutation__round__c[1469] ), 
        .A2(_f_permutation__round__n478 ), .ZN(_f_permutation__round__N5303 )
         );
  NOR2_X2 _f_permutation__round__U539  ( .A1(_f_permutation__round__c[1470] ), 
        .A2(_f_permutation__round__n473 ), .ZN(_f_permutation__round__N5301 )
         );
  NOR2_X2 _f_permutation__round__U538  ( .A1(_f_permutation__round__c[1471] ), 
        .A2(_f_permutation__round__n468 ), .ZN(_f_permutation__round__N5299 )
         );
  NOR2_X2 _f_permutation__round__U537  ( .A1(_f_permutation__round__c[1408] ), 
        .A2(_f_permutation__round__n463 ), .ZN(_f_permutation__round__N5297 )
         );
  NOR2_X2 _f_permutation__round__U536  ( .A1(_f_permutation__round__c[1409] ), 
        .A2(_f_permutation__round__n458 ), .ZN(_f_permutation__round__N5295 )
         );
  NOR2_X2 _f_permutation__round__U535  ( .A1(_f_permutation__round__c[1410] ), 
        .A2(_f_permutation__round__n453 ), .ZN(_f_permutation__round__N5293 )
         );
  NOR2_X2 _f_permutation__round__U534  ( .A1(_f_permutation__round__c[1411] ), 
        .A2(_f_permutation__round__n768 ), .ZN(_f_permutation__round__N5291 )
         );
  NOR2_X2 _f_permutation__round__U533  ( .A1(_f_permutation__round__c[1412] ), 
        .A2(_f_permutation__round__n763 ), .ZN(_f_permutation__round__N5289 )
         );
  NOR2_X2 _f_permutation__round__U532  ( .A1(_f_permutation__round__c[1413] ), 
        .A2(_f_permutation__round__n758 ), .ZN(_f_permutation__round__N5287 )
         );
  NOR2_X2 _f_permutation__round__U531  ( .A1(_f_permutation__round__c[1414] ), 
        .A2(_f_permutation__round__n753 ), .ZN(_f_permutation__round__N5285 )
         );
  NOR2_X2 _f_permutation__round__U530  ( .A1(_f_permutation__round__c[1415] ), 
        .A2(_f_permutation__round__n748 ), .ZN(_f_permutation__round__N5283 )
         );
  NOR2_X2 _f_permutation__round__U529  ( .A1(_f_permutation__round__c[1416] ), 
        .A2(_f_permutation__round__n743 ), .ZN(_f_permutation__round__N5281 )
         );
  NOR2_X2 _f_permutation__round__U528  ( .A1(_f_permutation__round__c[1417] ), 
        .A2(_f_permutation__round__n738 ), .ZN(_f_permutation__round__N5279 )
         );
  NOR2_X2 _f_permutation__round__U527  ( .A1(_f_permutation__round__c[1418] ), 
        .A2(_f_permutation__round__n733 ), .ZN(_f_permutation__round__N5277 )
         );
  NOR2_X2 _f_permutation__round__U526  ( .A1(_f_permutation__round__c[1419] ), 
        .A2(_f_permutation__round__n728 ), .ZN(_f_permutation__round__N5275 )
         );
  NOR2_X2 _f_permutation__round__U525  ( .A1(_f_permutation__round__c[1420] ), 
        .A2(_f_permutation__round__n723 ), .ZN(_f_permutation__round__N5273 )
         );
  NOR2_X2 _f_permutation__round__U524  ( .A1(_f_permutation__round__c[1421] ), 
        .A2(_f_permutation__round__n718 ), .ZN(_f_permutation__round__N5271 )
         );
  NOR2_X2 _f_permutation__round__U523  ( .A1(_f_permutation__round__c[1422] ), 
        .A2(_f_permutation__round__n713 ), .ZN(_f_permutation__round__N5269 )
         );
  NOR2_X2 _f_permutation__round__U522  ( .A1(_f_permutation__round__c[1423] ), 
        .A2(_f_permutation__round__n708 ), .ZN(_f_permutation__round__N5267 )
         );
  NOR2_X2 _f_permutation__round__U521  ( .A1(_f_permutation__round__c[1424] ), 
        .A2(_f_permutation__round__n703 ), .ZN(_f_permutation__round__N5265 )
         );
  NOR2_X2 _f_permutation__round__U520  ( .A1(_f_permutation__round__c[1425] ), 
        .A2(_f_permutation__round__n698 ), .ZN(_f_permutation__round__N5263 )
         );
  NOR2_X2 _f_permutation__round__U519  ( .A1(_f_permutation__round__c[1426] ), 
        .A2(_f_permutation__round__n693 ), .ZN(_f_permutation__round__N5261 )
         );
  NOR2_X2 _f_permutation__round__U518  ( .A1(_f_permutation__round__c[1427] ), 
        .A2(_f_permutation__round__n688 ), .ZN(_f_permutation__round__N5259 )
         );
  NOR2_X2 _f_permutation__round__U517  ( .A1(_f_permutation__round__c[1428] ), 
        .A2(_f_permutation__round__n683 ), .ZN(_f_permutation__round__N5257 )
         );
  NOR2_X2 _f_permutation__round__U516  ( .A1(_f_permutation__round__c[1429] ), 
        .A2(_f_permutation__round__n678 ), .ZN(_f_permutation__round__N5255 )
         );
  NOR2_X2 _f_permutation__round__U515  ( .A1(_f_permutation__round__c[1430] ), 
        .A2(_f_permutation__round__n673 ), .ZN(_f_permutation__round__N5253 )
         );
  NOR2_X2 _f_permutation__round__U514  ( .A1(_f_permutation__round__c[1431] ), 
        .A2(_f_permutation__round__n668 ), .ZN(_f_permutation__round__N5251 )
         );
  NOR2_X2 _f_permutation__round__U513  ( .A1(_f_permutation__round__c[1432] ), 
        .A2(_f_permutation__round__n663 ), .ZN(_f_permutation__round__N5249 )
         );
  NOR2_X2 _f_permutation__round__U448  ( .A1(_f_permutation__round__c[502] ), 
        .A2(_f_permutation__round__n521 ), .ZN(_f_permutation__round__N4735 )
         );
  NOR2_X2 _f_permutation__round__U447  ( .A1(_f_permutation__round__c[503] ), 
        .A2(_f_permutation__round__n516 ), .ZN(_f_permutation__round__N4733 )
         );
  NOR2_X2 _f_permutation__round__U446  ( .A1(_f_permutation__round__c[504] ), 
        .A2(_f_permutation__round__n511 ), .ZN(_f_permutation__round__N4731 )
         );
  NOR2_X2 _f_permutation__round__U445  ( .A1(_f_permutation__round__c[505] ), 
        .A2(_f_permutation__round__n506 ), .ZN(_f_permutation__round__N4729 )
         );
  NOR2_X2 _f_permutation__round__U444  ( .A1(_f_permutation__round__c[506] ), 
        .A2(_f_permutation__round__n501 ), .ZN(_f_permutation__round__N4727 )
         );
  NOR2_X2 _f_permutation__round__U443  ( .A1(_f_permutation__round__c[507] ), 
        .A2(_f_permutation__round__n496 ), .ZN(_f_permutation__round__N4725 )
         );
  NOR2_X2 _f_permutation__round__U442  ( .A1(_f_permutation__round__c[508] ), 
        .A2(_f_permutation__round__n491 ), .ZN(_f_permutation__round__N4723 )
         );
  NOR2_X2 _f_permutation__round__U441  ( .A1(_f_permutation__round__c[509] ), 
        .A2(_f_permutation__round__n486 ), .ZN(_f_permutation__round__N4721 )
         );
  NOR2_X2 _f_permutation__round__U440  ( .A1(_f_permutation__round__c[510] ), 
        .A2(_f_permutation__round__n481 ), .ZN(_f_permutation__round__N4719 )
         );
  NOR2_X2 _f_permutation__round__U439  ( .A1(_f_permutation__round__c[511] ), 
        .A2(_f_permutation__round__n476 ), .ZN(_f_permutation__round__N4717 )
         );
  NOR2_X2 _f_permutation__round__U438  ( .A1(_f_permutation__round__c[448] ), 
        .A2(_f_permutation__round__n471 ), .ZN(_f_permutation__round__N4715 )
         );
  NOR2_X2 _f_permutation__round__U437  ( .A1(_f_permutation__round__c[449] ), 
        .A2(_f_permutation__round__n466 ), .ZN(_f_permutation__round__N4713 )
         );
  NOR2_X2 _f_permutation__round__U436  ( .A1(_f_permutation__round__c[450] ), 
        .A2(_f_permutation__round__n461 ), .ZN(_f_permutation__round__N4711 )
         );
  NOR2_X2 _f_permutation__round__U435  ( .A1(_f_permutation__round__c[451] ), 
        .A2(_f_permutation__round__n456 ), .ZN(_f_permutation__round__N4709 )
         );
  NOR2_X2 _f_permutation__round__U434  ( .A1(_f_permutation__round__c[452] ), 
        .A2(_f_permutation__round__n451 ), .ZN(_f_permutation__round__N4707 )
         );
  NOR2_X2 _f_permutation__round__U433  ( .A1(_f_permutation__round__c[453] ), 
        .A2(_f_permutation__round__n766 ), .ZN(_f_permutation__round__N4705 )
         );
  NOR2_X2 _f_permutation__round__U432  ( .A1(_f_permutation__round__c[454] ), 
        .A2(_f_permutation__round__n761 ), .ZN(_f_permutation__round__N4703 )
         );
  NOR2_X2 _f_permutation__round__U431  ( .A1(_f_permutation__round__c[455] ), 
        .A2(_f_permutation__round__n756 ), .ZN(_f_permutation__round__N4701 )
         );
  NOR2_X2 _f_permutation__round__U430  ( .A1(_f_permutation__round__c[456] ), 
        .A2(_f_permutation__round__n751 ), .ZN(_f_permutation__round__N4699 )
         );
  NOR2_X2 _f_permutation__round__U429  ( .A1(_f_permutation__round__c[457] ), 
        .A2(_f_permutation__round__n746 ), .ZN(_f_permutation__round__N4697 )
         );
  NOR2_X2 _f_permutation__round__U428  ( .A1(_f_permutation__round__c[458] ), 
        .A2(_f_permutation__round__n741 ), .ZN(_f_permutation__round__N4695 )
         );
  NOR2_X2 _f_permutation__round__U427  ( .A1(_f_permutation__round__c[459] ), 
        .A2(_f_permutation__round__n736 ), .ZN(_f_permutation__round__N4693 )
         );
  NOR2_X2 _f_permutation__round__U426  ( .A1(_f_permutation__round__c[460] ), 
        .A2(_f_permutation__round__n731 ), .ZN(_f_permutation__round__N4691 )
         );
  NOR2_X2 _f_permutation__round__U425  ( .A1(_f_permutation__round__c[461] ), 
        .A2(_f_permutation__round__n726 ), .ZN(_f_permutation__round__N4689 )
         );
  NOR2_X2 _f_permutation__round__U424  ( .A1(_f_permutation__round__c[462] ), 
        .A2(_f_permutation__round__n721 ), .ZN(_f_permutation__round__N4687 )
         );
  NOR2_X2 _f_permutation__round__U423  ( .A1(_f_permutation__round__c[463] ), 
        .A2(_f_permutation__round__n716 ), .ZN(_f_permutation__round__N4685 )
         );
  NOR2_X2 _f_permutation__round__U422  ( .A1(_f_permutation__round__c[464] ), 
        .A2(_f_permutation__round__n711 ), .ZN(_f_permutation__round__N4683 )
         );
  NOR2_X2 _f_permutation__round__U421  ( .A1(_f_permutation__round__c[465] ), 
        .A2(_f_permutation__round__n706 ), .ZN(_f_permutation__round__N4681 )
         );
  NOR2_X2 _f_permutation__round__U420  ( .A1(_f_permutation__round__c[466] ), 
        .A2(_f_permutation__round__n701 ), .ZN(_f_permutation__round__N4679 )
         );
  NOR2_X2 _f_permutation__round__U419  ( .A1(_f_permutation__round__c[467] ), 
        .A2(_f_permutation__round__n696 ), .ZN(_f_permutation__round__N4677 )
         );
  NOR2_X2 _f_permutation__round__U418  ( .A1(_f_permutation__round__c[468] ), 
        .A2(_f_permutation__round__n691 ), .ZN(_f_permutation__round__N4675 )
         );
  NOR2_X2 _f_permutation__round__U417  ( .A1(_f_permutation__round__c[469] ), 
        .A2(_f_permutation__round__n686 ), .ZN(_f_permutation__round__N4673 )
         );
  NOR2_X2 _f_permutation__round__U416  ( .A1(_f_permutation__round__c[470] ), 
        .A2(_f_permutation__round__n681 ), .ZN(_f_permutation__round__N4671 )
         );
  NOR2_X2 _f_permutation__round__U415  ( .A1(_f_permutation__round__c[471] ), 
        .A2(_f_permutation__round__n676 ), .ZN(_f_permutation__round__N4669 )
         );
  NOR2_X2 _f_permutation__round__U414  ( .A1(_f_permutation__round__c[472] ), 
        .A2(_f_permutation__round__n671 ), .ZN(_f_permutation__round__N4667 )
         );
  NOR2_X2 _f_permutation__round__U413  ( .A1(_f_permutation__round__c[473] ), 
        .A2(_f_permutation__round__n666 ), .ZN(_f_permutation__round__N4665 )
         );
  NOR2_X2 _f_permutation__round__U412  ( .A1(_f_permutation__round__c[474] ), 
        .A2(_f_permutation__round__n661 ), .ZN(_f_permutation__round__N4663 )
         );
  NOR2_X2 _f_permutation__round__U411  ( .A1(_f_permutation__round__c[475] ), 
        .A2(_f_permutation__round__n656 ), .ZN(_f_permutation__round__N4661 )
         );
  NOR2_X2 _f_permutation__round__U410  ( .A1(_f_permutation__round__c[476] ), 
        .A2(_f_permutation__round__n651 ), .ZN(_f_permutation__round__N4659 )
         );
  NOR2_X2 _f_permutation__round__U409  ( .A1(_f_permutation__round__c[477] ), 
        .A2(_f_permutation__round__n646 ), .ZN(_f_permutation__round__N4657 )
         );
  NOR2_X2 _f_permutation__round__U408  ( .A1(_f_permutation__round__c[478] ), 
        .A2(_f_permutation__round__n641 ), .ZN(_f_permutation__round__N4655 )
         );
  NOR2_X2 _f_permutation__round__U407  ( .A1(_f_permutation__round__c[479] ), 
        .A2(_f_permutation__round__n636 ), .ZN(_f_permutation__round__N4653 )
         );
  NOR2_X2 _f_permutation__round__U406  ( .A1(_f_permutation__round__c[480] ), 
        .A2(_f_permutation__round__n631 ), .ZN(_f_permutation__round__N4651 )
         );
  NOR2_X2 _f_permutation__round__U405  ( .A1(_f_permutation__round__c[481] ), 
        .A2(_f_permutation__round__n626 ), .ZN(_f_permutation__round__N4649 )
         );
  NOR2_X2 _f_permutation__round__U404  ( .A1(_f_permutation__round__c[482] ), 
        .A2(_f_permutation__round__n621 ), .ZN(_f_permutation__round__N4647 )
         );
  NOR2_X2 _f_permutation__round__U403  ( .A1(_f_permutation__round__c[483] ), 
        .A2(_f_permutation__round__n616 ), .ZN(_f_permutation__round__N4645 )
         );
  NOR2_X2 _f_permutation__round__U402  ( .A1(_f_permutation__round__c[484] ), 
        .A2(_f_permutation__round__n611 ), .ZN(_f_permutation__round__N4643 )
         );
  NOR2_X2 _f_permutation__round__U401  ( .A1(_f_permutation__round__c[485] ), 
        .A2(_f_permutation__round__n606 ), .ZN(_f_permutation__round__N4641 )
         );
  NOR2_X2 _f_permutation__round__U400  ( .A1(_f_permutation__round__c[486] ), 
        .A2(_f_permutation__round__n601 ), .ZN(_f_permutation__round__N4639 )
         );
  NOR2_X2 _f_permutation__round__U399  ( .A1(_f_permutation__round__c[487] ), 
        .A2(_f_permutation__round__n596 ), .ZN(_f_permutation__round__N4637 )
         );
  NOR2_X2 _f_permutation__round__U398  ( .A1(_f_permutation__round__c[488] ), 
        .A2(_f_permutation__round__n591 ), .ZN(_f_permutation__round__N4635 )
         );
  NOR2_X2 _f_permutation__round__U397  ( .A1(_f_permutation__round__c[489] ), 
        .A2(_f_permutation__round__n586 ), .ZN(_f_permutation__round__N4633 )
         );
  NOR2_X2 _f_permutation__round__U396  ( .A1(_f_permutation__round__c[490] ), 
        .A2(_f_permutation__round__n581 ), .ZN(_f_permutation__round__N4631 )
         );
  NOR2_X2 _f_permutation__round__U395  ( .A1(_f_permutation__round__c[491] ), 
        .A2(_f_permutation__round__n576 ), .ZN(_f_permutation__round__N4629 )
         );
  NOR2_X2 _f_permutation__round__U394  ( .A1(_f_permutation__round__c[492] ), 
        .A2(_f_permutation__round__n571 ), .ZN(_f_permutation__round__N4627 )
         );
  NOR2_X2 _f_permutation__round__U393  ( .A1(_f_permutation__round__c[493] ), 
        .A2(_f_permutation__round__n566 ), .ZN(_f_permutation__round__N4625 )
         );
  NOR2_X2 _f_permutation__round__U392  ( .A1(_f_permutation__round__c[494] ), 
        .A2(_f_permutation__round__n561 ), .ZN(_f_permutation__round__N4623 )
         );
  NOR2_X2 _f_permutation__round__U391  ( .A1(_f_permutation__round__c[495] ), 
        .A2(_f_permutation__round__n556 ), .ZN(_f_permutation__round__N4621 )
         );
  NOR2_X2 _f_permutation__round__U390  ( .A1(_f_permutation__round__c[496] ), 
        .A2(_f_permutation__round__n551 ), .ZN(_f_permutation__round__N4619 )
         );
  NOR2_X2 _f_permutation__round__U389  ( .A1(_f_permutation__round__c[497] ), 
        .A2(_f_permutation__round__n546 ), .ZN(_f_permutation__round__N4617 )
         );
  NOR2_X2 _f_permutation__round__U388  ( .A1(_f_permutation__round__c[498] ), 
        .A2(_f_permutation__round__n541 ), .ZN(_f_permutation__round__N4615 )
         );
  NOR2_X2 _f_permutation__round__U387  ( .A1(_f_permutation__round__c[499] ), 
        .A2(_f_permutation__round__n536 ), .ZN(_f_permutation__round__N4613 )
         );
  NOR2_X2 _f_permutation__round__U386  ( .A1(_f_permutation__round__c[500] ), 
        .A2(_f_permutation__round__n531 ), .ZN(_f_permutation__round__N4611 )
         );
  NOR2_X2 _f_permutation__round__U385  ( .A1(_f_permutation__round__c[501] ), 
        .A2(_f_permutation__round__n526 ), .ZN(_f_permutation__round__N4609 )
         );
  NOR2_X2 _f_permutation__round__U320  ( .A1(_f_permutation__round__c[1127] ), 
        .A2(_f_permutation__round__n62 ), .ZN(_f_permutation__round__N4095 )
         );
  NOR2_X2 _f_permutation__round__U319  ( .A1(_f_permutation__round__c[1128] ), 
        .A2(_f_permutation__round__n55 ), .ZN(_f_permutation__round__N4093 )
         );
  NOR2_X2 _f_permutation__round__U318  ( .A1(_f_permutation__round__c[1129] ), 
        .A2(_f_permutation__round__n48 ), .ZN(_f_permutation__round__N4091 )
         );
  NOR2_X2 _f_permutation__round__U317  ( .A1(_f_permutation__round__c[1130] ), 
        .A2(_f_permutation__round__n41 ), .ZN(_f_permutation__round__N4089 )
         );
  NOR2_X2 _f_permutation__round__U316  ( .A1(_f_permutation__round__c[1131] ), 
        .A2(_f_permutation__round__n34 ), .ZN(_f_permutation__round__N4087 )
         );
  NOR2_X2 _f_permutation__round__U315  ( .A1(_f_permutation__round__c[1132] ), 
        .A2(_f_permutation__round__n27 ), .ZN(_f_permutation__round__N4085 )
         );
  NOR2_X2 _f_permutation__round__U314  ( .A1(_f_permutation__round__c[1133] ), 
        .A2(_f_permutation__round__n20 ), .ZN(_f_permutation__round__N4083 )
         );
  NOR2_X2 _f_permutation__round__U313  ( .A1(_f_permutation__round__c[1134] ), 
        .A2(_f_permutation__round__n13 ), .ZN(_f_permutation__round__N4081 )
         );
  NOR2_X2 _f_permutation__round__U312  ( .A1(_f_permutation__round__c[1135] ), 
        .A2(_f_permutation__round__n6 ), .ZN(_f_permutation__round__N4079 ) );
  NOR2_X2 _f_permutation__round__U311  ( .A1(_f_permutation__round__c[1136] ), 
        .A2(_f_permutation__round__n447 ), .ZN(_f_permutation__round__N4077 )
         );
  NOR2_X2 _f_permutation__round__U310  ( .A1(_f_permutation__round__c[1137] ), 
        .A2(_f_permutation__round__n440 ), .ZN(_f_permutation__round__N4075 )
         );
  NOR2_X2 _f_permutation__round__U309  ( .A1(_f_permutation__round__c[1138] ), 
        .A2(_f_permutation__round__n433 ), .ZN(_f_permutation__round__N4073 )
         );
  NOR2_X2 _f_permutation__round__U308  ( .A1(_f_permutation__round__c[1139] ), 
        .A2(_f_permutation__round__n426 ), .ZN(_f_permutation__round__N4071 )
         );
  NOR2_X2 _f_permutation__round__U307  ( .A1(_f_permutation__round__c[1140] ), 
        .A2(_f_permutation__round__n419 ), .ZN(_f_permutation__round__N4069 )
         );
  NOR2_X2 _f_permutation__round__U306  ( .A1(_f_permutation__round__c[1141] ), 
        .A2(_f_permutation__round__n412 ), .ZN(_f_permutation__round__N4067 )
         );
  NOR2_X2 _f_permutation__round__U305  ( .A1(_f_permutation__round__c[1142] ), 
        .A2(_f_permutation__round__n405 ), .ZN(_f_permutation__round__N4065 )
         );
  NOR2_X2 _f_permutation__round__U304  ( .A1(_f_permutation__round__c[1143] ), 
        .A2(_f_permutation__round__n398 ), .ZN(_f_permutation__round__N4063 )
         );
  NOR2_X2 _f_permutation__round__U303  ( .A1(_f_permutation__round__c[1144] ), 
        .A2(_f_permutation__round__n391 ), .ZN(_f_permutation__round__N4061 )
         );
  NOR2_X2 _f_permutation__round__U302  ( .A1(_f_permutation__round__c[1145] ), 
        .A2(_f_permutation__round__n384 ), .ZN(_f_permutation__round__N4059 )
         );
  NOR2_X2 _f_permutation__round__U301  ( .A1(_f_permutation__round__c[1146] ), 
        .A2(_f_permutation__round__n377 ), .ZN(_f_permutation__round__N4057 )
         );
  NOR2_X2 _f_permutation__round__U300  ( .A1(_f_permutation__round__c[1147] ), 
        .A2(_f_permutation__round__n370 ), .ZN(_f_permutation__round__N4055 )
         );
  NOR2_X2 _f_permutation__round__U299  ( .A1(_f_permutation__round__c[1148] ), 
        .A2(_f_permutation__round__n363 ), .ZN(_f_permutation__round__N4053 )
         );
  NOR2_X2 _f_permutation__round__U298  ( .A1(_f_permutation__round__c[1149] ), 
        .A2(_f_permutation__round__n356 ), .ZN(_f_permutation__round__N4051 )
         );
  NOR2_X2 _f_permutation__round__U297  ( .A1(_f_permutation__round__c[1150] ), 
        .A2(_f_permutation__round__n349 ), .ZN(_f_permutation__round__N4049 )
         );
  NOR2_X2 _f_permutation__round__U296  ( .A1(_f_permutation__round__c[1151] ), 
        .A2(_f_permutation__round__n342 ), .ZN(_f_permutation__round__N4047 )
         );
  NOR2_X2 _f_permutation__round__U295  ( .A1(_f_permutation__round__c[1088] ), 
        .A2(_f_permutation__round__n335 ), .ZN(_f_permutation__round__N4045 )
         );
  NOR2_X2 _f_permutation__round__U294  ( .A1(_f_permutation__round__c[1089] ), 
        .A2(_f_permutation__round__n328 ), .ZN(_f_permutation__round__N4043 )
         );
  NOR2_X2 _f_permutation__round__U293  ( .A1(_f_permutation__round__c[1090] ), 
        .A2(_f_permutation__round__n321 ), .ZN(_f_permutation__round__N4041 )
         );
  NOR2_X2 _f_permutation__round__U292  ( .A1(_f_permutation__round__c[1091] ), 
        .A2(_f_permutation__round__n314 ), .ZN(_f_permutation__round__N4039 )
         );
  NOR2_X2 _f_permutation__round__U291  ( .A1(_f_permutation__round__c[1092] ), 
        .A2(_f_permutation__round__n307 ), .ZN(_f_permutation__round__N4037 )
         );
  NOR2_X2 _f_permutation__round__U290  ( .A1(_f_permutation__round__c[1093] ), 
        .A2(_f_permutation__round__n300 ), .ZN(_f_permutation__round__N4035 )
         );
  NOR2_X2 _f_permutation__round__U289  ( .A1(_f_permutation__round__c[1094] ), 
        .A2(_f_permutation__round__n293 ), .ZN(_f_permutation__round__N4033 )
         );
  NOR2_X2 _f_permutation__round__U288  ( .A1(_f_permutation__round__c[1095] ), 
        .A2(_f_permutation__round__n286 ), .ZN(_f_permutation__round__N4031 )
         );
  NOR2_X2 _f_permutation__round__U287  ( .A1(_f_permutation__round__c[1096] ), 
        .A2(_f_permutation__round__n279 ), .ZN(_f_permutation__round__N4029 )
         );
  NOR2_X2 _f_permutation__round__U286  ( .A1(_f_permutation__round__c[1097] ), 
        .A2(_f_permutation__round__n272 ), .ZN(_f_permutation__round__N4027 )
         );
  NOR2_X2 _f_permutation__round__U285  ( .A1(_f_permutation__round__c[1098] ), 
        .A2(_f_permutation__round__n265 ), .ZN(_f_permutation__round__N4025 )
         );
  NOR2_X2 _f_permutation__round__U284  ( .A1(_f_permutation__round__c[1099] ), 
        .A2(_f_permutation__round__n258 ), .ZN(_f_permutation__round__N4023 )
         );
  NOR2_X2 _f_permutation__round__U283  ( .A1(_f_permutation__round__c[1100] ), 
        .A2(_f_permutation__round__n251 ), .ZN(_f_permutation__round__N4021 )
         );
  NOR2_X2 _f_permutation__round__U282  ( .A1(_f_permutation__round__c[1101] ), 
        .A2(_f_permutation__round__n244 ), .ZN(_f_permutation__round__N4019 )
         );
  NOR2_X2 _f_permutation__round__U281  ( .A1(_f_permutation__round__c[1102] ), 
        .A2(_f_permutation__round__n237 ), .ZN(_f_permutation__round__N4017 )
         );
  NOR2_X2 _f_permutation__round__U280  ( .A1(_f_permutation__round__c[1103] ), 
        .A2(_f_permutation__round__n230 ), .ZN(_f_permutation__round__N4015 )
         );
  NOR2_X2 _f_permutation__round__U279  ( .A1(_f_permutation__round__c[1104] ), 
        .A2(_f_permutation__round__n223 ), .ZN(_f_permutation__round__N4013 )
         );
  NOR2_X2 _f_permutation__round__U278  ( .A1(_f_permutation__round__c[1105] ), 
        .A2(_f_permutation__round__n216 ), .ZN(_f_permutation__round__N4011 )
         );
  NOR2_X2 _f_permutation__round__U277  ( .A1(_f_permutation__round__c[1106] ), 
        .A2(_f_permutation__round__n209 ), .ZN(_f_permutation__round__N4009 )
         );
  NOR2_X2 _f_permutation__round__U276  ( .A1(_f_permutation__round__c[1107] ), 
        .A2(_f_permutation__round__n202 ), .ZN(_f_permutation__round__N4007 )
         );
  NOR2_X2 _f_permutation__round__U275  ( .A1(_f_permutation__round__c[1108] ), 
        .A2(_f_permutation__round__n195 ), .ZN(_f_permutation__round__N4005 )
         );
  NOR2_X2 _f_permutation__round__U274  ( .A1(_f_permutation__round__c[1109] ), 
        .A2(_f_permutation__round__n188 ), .ZN(_f_permutation__round__N4003 )
         );
  NOR2_X2 _f_permutation__round__U273  ( .A1(_f_permutation__round__c[1110] ), 
        .A2(_f_permutation__round__n181 ), .ZN(_f_permutation__round__N4001 )
         );
  NOR2_X2 _f_permutation__round__U272  ( .A1(_f_permutation__round__c[1111] ), 
        .A2(_f_permutation__round__n174 ), .ZN(_f_permutation__round__N3999 )
         );
  NOR2_X2 _f_permutation__round__U271  ( .A1(_f_permutation__round__c[1112] ), 
        .A2(_f_permutation__round__n167 ), .ZN(_f_permutation__round__N3997 )
         );
  NOR2_X2 _f_permutation__round__U270  ( .A1(_f_permutation__round__c[1113] ), 
        .A2(_f_permutation__round__n160 ), .ZN(_f_permutation__round__N3995 )
         );
  NOR2_X2 _f_permutation__round__U269  ( .A1(_f_permutation__round__c[1114] ), 
        .A2(_f_permutation__round__n153 ), .ZN(_f_permutation__round__N3993 )
         );
  NOR2_X2 _f_permutation__round__U268  ( .A1(_f_permutation__round__c[1115] ), 
        .A2(_f_permutation__round__n146 ), .ZN(_f_permutation__round__N3991 )
         );
  NOR2_X2 _f_permutation__round__U267  ( .A1(_f_permutation__round__c[1116] ), 
        .A2(_f_permutation__round__n139 ), .ZN(_f_permutation__round__N3989 )
         );
  NOR2_X2 _f_permutation__round__U266  ( .A1(_f_permutation__round__c[1117] ), 
        .A2(_f_permutation__round__n132 ), .ZN(_f_permutation__round__N3987 )
         );
  NOR2_X2 _f_permutation__round__U265  ( .A1(_f_permutation__round__c[1118] ), 
        .A2(_f_permutation__round__n125 ), .ZN(_f_permutation__round__N3985 )
         );
  NOR2_X2 _f_permutation__round__U264  ( .A1(_f_permutation__round__c[1119] ), 
        .A2(_f_permutation__round__n118 ), .ZN(_f_permutation__round__N3983 )
         );
  NOR2_X2 _f_permutation__round__U263  ( .A1(_f_permutation__round__c[1120] ), 
        .A2(_f_permutation__round__n111 ), .ZN(_f_permutation__round__N3981 )
         );
  NOR2_X2 _f_permutation__round__U262  ( .A1(_f_permutation__round__c[1121] ), 
        .A2(_f_permutation__round__n104 ), .ZN(_f_permutation__round__N3979 )
         );
  NOR2_X2 _f_permutation__round__U261  ( .A1(_f_permutation__round__c[1122] ), 
        .A2(_f_permutation__round__n97 ), .ZN(_f_permutation__round__N3977 )
         );
  NOR2_X2 _f_permutation__round__U260  ( .A1(_f_permutation__round__c[1123] ), 
        .A2(_f_permutation__round__n90 ), .ZN(_f_permutation__round__N3975 )
         );
  NOR2_X2 _f_permutation__round__U259  ( .A1(_f_permutation__round__c[1124] ), 
        .A2(_f_permutation__round__n83 ), .ZN(_f_permutation__round__N3973 )
         );
  NOR2_X2 _f_permutation__round__U258  ( .A1(_f_permutation__round__c[1125] ), 
        .A2(_f_permutation__round__n76 ), .ZN(_f_permutation__round__N3971 )
         );
  NOR2_X2 _f_permutation__round__U257  ( .A1(_f_permutation__round__c[1126] ), 
        .A2(_f_permutation__round__n69 ), .ZN(_f_permutation__round__N3969 )
         );
  NOR2_X2 _f_permutation__round__U256  ( .A1(_f_permutation__round__c[189] ), 
        .A2(_f_permutation__round__n311 ), .ZN(_f_permutation__round__N3455 )
         );
  NOR2_X2 _f_permutation__round__U255  ( .A1(_f_permutation__round__c[190] ), 
        .A2(_f_permutation__round__n304 ), .ZN(_f_permutation__round__N3453 )
         );
  NOR2_X2 _f_permutation__round__U254  ( .A1(_f_permutation__round__c[191] ), 
        .A2(_f_permutation__round__n297 ), .ZN(_f_permutation__round__N3451 )
         );
  NOR2_X2 _f_permutation__round__U253  ( .A1(_f_permutation__round__c[128] ), 
        .A2(_f_permutation__round__n290 ), .ZN(_f_permutation__round__N3449 )
         );
  NOR2_X2 _f_permutation__round__U252  ( .A1(_f_permutation__round__c[129] ), 
        .A2(_f_permutation__round__n283 ), .ZN(_f_permutation__round__N3447 )
         );
  NOR2_X2 _f_permutation__round__U251  ( .A1(_f_permutation__round__c[130] ), 
        .A2(_f_permutation__round__n276 ), .ZN(_f_permutation__round__N3445 )
         );
  NOR2_X2 _f_permutation__round__U250  ( .A1(_f_permutation__round__c[131] ), 
        .A2(_f_permutation__round__n269 ), .ZN(_f_permutation__round__N3443 )
         );
  NOR2_X2 _f_permutation__round__U249  ( .A1(_f_permutation__round__c[132] ), 
        .A2(_f_permutation__round__n262 ), .ZN(_f_permutation__round__N3441 )
         );
  NOR2_X2 _f_permutation__round__U248  ( .A1(_f_permutation__round__c[133] ), 
        .A2(_f_permutation__round__n255 ), .ZN(_f_permutation__round__N3439 )
         );
  NOR2_X2 _f_permutation__round__U247  ( .A1(_f_permutation__round__c[134] ), 
        .A2(_f_permutation__round__n248 ), .ZN(_f_permutation__round__N3437 )
         );
  NOR2_X2 _f_permutation__round__U246  ( .A1(_f_permutation__round__c[135] ), 
        .A2(_f_permutation__round__n241 ), .ZN(_f_permutation__round__N3435 )
         );
  NOR2_X2 _f_permutation__round__U245  ( .A1(_f_permutation__round__c[136] ), 
        .A2(_f_permutation__round__n234 ), .ZN(_f_permutation__round__N3433 )
         );
  NOR2_X2 _f_permutation__round__U244  ( .A1(_f_permutation__round__c[137] ), 
        .A2(_f_permutation__round__n227 ), .ZN(_f_permutation__round__N3431 )
         );
  NOR2_X2 _f_permutation__round__U243  ( .A1(_f_permutation__round__c[138] ), 
        .A2(_f_permutation__round__n220 ), .ZN(_f_permutation__round__N3429 )
         );
  NOR2_X2 _f_permutation__round__U242  ( .A1(_f_permutation__round__c[139] ), 
        .A2(_f_permutation__round__n213 ), .ZN(_f_permutation__round__N3427 )
         );
  NOR2_X2 _f_permutation__round__U241  ( .A1(_f_permutation__round__c[140] ), 
        .A2(_f_permutation__round__n206 ), .ZN(_f_permutation__round__N3425 )
         );
  NOR2_X2 _f_permutation__round__U240  ( .A1(_f_permutation__round__c[141] ), 
        .A2(_f_permutation__round__n199 ), .ZN(_f_permutation__round__N3423 )
         );
  NOR2_X2 _f_permutation__round__U239  ( .A1(_f_permutation__round__c[142] ), 
        .A2(_f_permutation__round__n192 ), .ZN(_f_permutation__round__N3421 )
         );
  NOR2_X2 _f_permutation__round__U238  ( .A1(_f_permutation__round__c[143] ), 
        .A2(_f_permutation__round__n185 ), .ZN(_f_permutation__round__N3419 )
         );
  NOR2_X2 _f_permutation__round__U237  ( .A1(_f_permutation__round__c[144] ), 
        .A2(_f_permutation__round__n178 ), .ZN(_f_permutation__round__N3417 )
         );
  NOR2_X2 _f_permutation__round__U236  ( .A1(_f_permutation__round__c[145] ), 
        .A2(_f_permutation__round__n171 ), .ZN(_f_permutation__round__N3415 )
         );
  NOR2_X2 _f_permutation__round__U235  ( .A1(_f_permutation__round__c[146] ), 
        .A2(_f_permutation__round__n164 ), .ZN(_f_permutation__round__N3413 )
         );
  NOR2_X2 _f_permutation__round__U234  ( .A1(_f_permutation__round__c[147] ), 
        .A2(_f_permutation__round__n157 ), .ZN(_f_permutation__round__N3411 )
         );
  NOR2_X2 _f_permutation__round__U233  ( .A1(_f_permutation__round__c[148] ), 
        .A2(_f_permutation__round__n150 ), .ZN(_f_permutation__round__N3409 )
         );
  NOR2_X2 _f_permutation__round__U232  ( .A1(_f_permutation__round__c[149] ), 
        .A2(_f_permutation__round__n143 ), .ZN(_f_permutation__round__N3407 )
         );
  NOR2_X2 _f_permutation__round__U231  ( .A1(_f_permutation__round__c[150] ), 
        .A2(_f_permutation__round__n136 ), .ZN(_f_permutation__round__N3405 )
         );
  NOR2_X2 _f_permutation__round__U230  ( .A1(_f_permutation__round__c[151] ), 
        .A2(_f_permutation__round__n129 ), .ZN(_f_permutation__round__N3403 )
         );
  NOR2_X2 _f_permutation__round__U229  ( .A1(_f_permutation__round__c[152] ), 
        .A2(_f_permutation__round__n122 ), .ZN(_f_permutation__round__N3401 )
         );
  NOR2_X2 _f_permutation__round__U228  ( .A1(_f_permutation__round__c[153] ), 
        .A2(_f_permutation__round__n115 ), .ZN(_f_permutation__round__N3399 )
         );
  NOR2_X2 _f_permutation__round__U227  ( .A1(_f_permutation__round__c[154] ), 
        .A2(_f_permutation__round__n108 ), .ZN(_f_permutation__round__N3397 )
         );
  NOR2_X2 _f_permutation__round__U226  ( .A1(_f_permutation__round__c[155] ), 
        .A2(_f_permutation__round__n101 ), .ZN(_f_permutation__round__N3395 )
         );
  NOR2_X2 _f_permutation__round__U225  ( .A1(_f_permutation__round__c[156] ), 
        .A2(_f_permutation__round__n94 ), .ZN(_f_permutation__round__N3393 )
         );
  NOR2_X2 _f_permutation__round__U224  ( .A1(_f_permutation__round__c[157] ), 
        .A2(_f_permutation__round__n87 ), .ZN(_f_permutation__round__N3391 )
         );
  NOR2_X2 _f_permutation__round__U223  ( .A1(_f_permutation__round__c[158] ), 
        .A2(_f_permutation__round__n80 ), .ZN(_f_permutation__round__N3389 )
         );
  NOR2_X2 _f_permutation__round__U222  ( .A1(_f_permutation__round__c[159] ), 
        .A2(_f_permutation__round__n73 ), .ZN(_f_permutation__round__N3387 )
         );
  NOR2_X2 _f_permutation__round__U221  ( .A1(_f_permutation__round__c[160] ), 
        .A2(_f_permutation__round__n66 ), .ZN(_f_permutation__round__N3385 )
         );
  NOR2_X2 _f_permutation__round__U220  ( .A1(_f_permutation__round__c[161] ), 
        .A2(_f_permutation__round__n59 ), .ZN(_f_permutation__round__N3383 )
         );
  NOR2_X2 _f_permutation__round__U219  ( .A1(_f_permutation__round__c[162] ), 
        .A2(_f_permutation__round__n52 ), .ZN(_f_permutation__round__N3381 )
         );
  NOR2_X2 _f_permutation__round__U218  ( .A1(_f_permutation__round__c[163] ), 
        .A2(_f_permutation__round__n45 ), .ZN(_f_permutation__round__N3379 )
         );
  NOR2_X2 _f_permutation__round__U217  ( .A1(_f_permutation__round__c[164] ), 
        .A2(_f_permutation__round__n38 ), .ZN(_f_permutation__round__N3377 )
         );
  NOR2_X2 _f_permutation__round__U216  ( .A1(_f_permutation__round__c[165] ), 
        .A2(_f_permutation__round__n31 ), .ZN(_f_permutation__round__N3375 )
         );
  NOR2_X2 _f_permutation__round__U215  ( .A1(_f_permutation__round__c[166] ), 
        .A2(_f_permutation__round__n24 ), .ZN(_f_permutation__round__N3373 )
         );
  NOR2_X2 _f_permutation__round__U214  ( .A1(_f_permutation__round__c[167] ), 
        .A2(_f_permutation__round__n17 ), .ZN(_f_permutation__round__N3371 )
         );
  NOR2_X2 _f_permutation__round__U213  ( .A1(_f_permutation__round__c[168] ), 
        .A2(_f_permutation__round__n10 ), .ZN(_f_permutation__round__N3369 )
         );
  NOR2_X2 _f_permutation__round__U212  ( .A1(_f_permutation__round__c[169] ), 
        .A2(_f_permutation__round__n3 ), .ZN(_f_permutation__round__N3367 ) );
  NOR2_X2 _f_permutation__round__U211  ( .A1(_f_permutation__round__c[170] ), 
        .A2(_f_permutation__round__n444 ), .ZN(_f_permutation__round__N3365 )
         );
  NOR2_X2 _f_permutation__round__U210  ( .A1(_f_permutation__round__c[171] ), 
        .A2(_f_permutation__round__n437 ), .ZN(_f_permutation__round__N3363 )
         );
  NOR2_X2 _f_permutation__round__U209  ( .A1(_f_permutation__round__c[172] ), 
        .A2(_f_permutation__round__n430 ), .ZN(_f_permutation__round__N3361 )
         );
  NOR2_X2 _f_permutation__round__U208  ( .A1(_f_permutation__round__c[173] ), 
        .A2(_f_permutation__round__n423 ), .ZN(_f_permutation__round__N3359 )
         );
  NOR2_X2 _f_permutation__round__U207  ( .A1(_f_permutation__round__c[174] ), 
        .A2(_f_permutation__round__n416 ), .ZN(_f_permutation__round__N3357 )
         );
  NOR2_X2 _f_permutation__round__U206  ( .A1(_f_permutation__round__c[175] ), 
        .A2(_f_permutation__round__n409 ), .ZN(_f_permutation__round__N3355 )
         );
  NOR2_X2 _f_permutation__round__U205  ( .A1(_f_permutation__round__c[176] ), 
        .A2(_f_permutation__round__n402 ), .ZN(_f_permutation__round__N3353 )
         );
  NOR2_X2 _f_permutation__round__U204  ( .A1(_f_permutation__round__c[177] ), 
        .A2(_f_permutation__round__n395 ), .ZN(_f_permutation__round__N3351 )
         );
  NOR2_X2 _f_permutation__round__U203  ( .A1(_f_permutation__round__c[178] ), 
        .A2(_f_permutation__round__n388 ), .ZN(_f_permutation__round__N3349 )
         );
  NOR2_X2 _f_permutation__round__U202  ( .A1(_f_permutation__round__c[179] ), 
        .A2(_f_permutation__round__n381 ), .ZN(_f_permutation__round__N3347 )
         );
  NOR2_X2 _f_permutation__round__U201  ( .A1(_f_permutation__round__c[180] ), 
        .A2(_f_permutation__round__n374 ), .ZN(_f_permutation__round__N3345 )
         );
  NOR2_X2 _f_permutation__round__U200  ( .A1(_f_permutation__round__c[181] ), 
        .A2(_f_permutation__round__n367 ), .ZN(_f_permutation__round__N3343 )
         );
  NOR2_X2 _f_permutation__round__U199  ( .A1(_f_permutation__round__c[182] ), 
        .A2(_f_permutation__round__n360 ), .ZN(_f_permutation__round__N3341 )
         );
  NOR2_X2 _f_permutation__round__U198  ( .A1(_f_permutation__round__c[183] ), 
        .A2(_f_permutation__round__n353 ), .ZN(_f_permutation__round__N3339 )
         );
  NOR2_X2 _f_permutation__round__U197  ( .A1(_f_permutation__round__c[184] ), 
        .A2(_f_permutation__round__n346 ), .ZN(_f_permutation__round__N3337 )
         );
  NOR2_X2 _f_permutation__round__U196  ( .A1(_f_permutation__round__c[185] ), 
        .A2(_f_permutation__round__n339 ), .ZN(_f_permutation__round__N3335 )
         );
  NOR2_X2 _f_permutation__round__U195  ( .A1(_f_permutation__round__c[186] ), 
        .A2(_f_permutation__round__n332 ), .ZN(_f_permutation__round__N3333 )
         );
  NOR2_X2 _f_permutation__round__U194  ( .A1(_f_permutation__round__c[187] ), 
        .A2(_f_permutation__round__n325 ), .ZN(_f_permutation__round__N3331 )
         );
  NOR2_X2 _f_permutation__round__U193  ( .A1(_f_permutation__round__c[188] ), 
        .A2(_f_permutation__round__n318 ), .ZN(_f_permutation__round__N3329 )
         );
  NOR2_X2 _f_permutation__round__U128  ( .A1(_f_permutation__round__c[789] ), 
        .A2(_f_permutation__round__n831 ), .ZN(_f_permutation__round__N2815 )
         );
  NOR2_X2 _f_permutation__round__U127  ( .A1(_f_permutation__round__c[790] ), 
        .A2(_f_permutation__round__n828 ), .ZN(_f_permutation__round__N2813 )
         );
  NOR2_X2 _f_permutation__round__U126  ( .A1(_f_permutation__round__c[791] ), 
        .A2(_f_permutation__round__n825 ), .ZN(_f_permutation__round__N2811 )
         );
  NOR2_X2 _f_permutation__round__U125  ( .A1(_f_permutation__round__c[792] ), 
        .A2(_f_permutation__round__n822 ), .ZN(_f_permutation__round__N2809 )
         );
  NOR2_X2 _f_permutation__round__U124  ( .A1(_f_permutation__round__c[793] ), 
        .A2(_f_permutation__round__n819 ), .ZN(_f_permutation__round__N2807 )
         );
  NOR2_X2 _f_permutation__round__U123  ( .A1(_f_permutation__round__c[794] ), 
        .A2(_f_permutation__round__n816 ), .ZN(_f_permutation__round__N2805 )
         );
  NOR2_X2 _f_permutation__round__U122  ( .A1(_f_permutation__round__c[795] ), 
        .A2(_f_permutation__round__n813 ), .ZN(_f_permutation__round__N2803 )
         );
  NOR2_X2 _f_permutation__round__U121  ( .A1(_f_permutation__round__c[796] ), 
        .A2(_f_permutation__round__n810 ), .ZN(_f_permutation__round__N2801 )
         );
  NOR2_X2 _f_permutation__round__U120  ( .A1(_f_permutation__round__c[797] ), 
        .A2(_f_permutation__round__n807 ), .ZN(_f_permutation__round__N2799 )
         );
  NOR2_X2 _f_permutation__round__U119  ( .A1(_f_permutation__round__c[798] ), 
        .A2(_f_permutation__round__n804 ), .ZN(_f_permutation__round__N2797 )
         );
  NOR2_X2 _f_permutation__round__U118  ( .A1(_f_permutation__round__c[799] ), 
        .A2(_f_permutation__round__n801 ), .ZN(_f_permutation__round__N2795 )
         );
  NOR2_X2 _f_permutation__round__U117  ( .A1(_f_permutation__round__c[800] ), 
        .A2(_f_permutation__round__n798 ), .ZN(_f_permutation__round__N2793 )
         );
  NOR2_X2 _f_permutation__round__U116  ( .A1(_f_permutation__round__c[801] ), 
        .A2(_f_permutation__round__n795 ), .ZN(_f_permutation__round__N2791 )
         );
  NOR2_X2 _f_permutation__round__U115  ( .A1(_f_permutation__round__c[802] ), 
        .A2(_f_permutation__round__n792 ), .ZN(_f_permutation__round__N2789 )
         );
  NOR2_X2 _f_permutation__round__U114  ( .A1(_f_permutation__round__c[803] ), 
        .A2(_f_permutation__round__n789 ), .ZN(_f_permutation__round__N2787 )
         );
  NOR2_X2 _f_permutation__round__U113  ( .A1(_f_permutation__round__c[804] ), 
        .A2(_f_permutation__round__n786 ), .ZN(_f_permutation__round__N2785 )
         );
  NOR2_X2 _f_permutation__round__U112  ( .A1(_f_permutation__round__c[805] ), 
        .A2(_f_permutation__round__n783 ), .ZN(_f_permutation__round__N2783 )
         );
  NOR2_X2 _f_permutation__round__U111  ( .A1(_f_permutation__round__c[806] ), 
        .A2(_f_permutation__round__n780 ), .ZN(_f_permutation__round__N2781 )
         );
  NOR2_X2 _f_permutation__round__U110  ( .A1(_f_permutation__round__c[807] ), 
        .A2(_f_permutation__round__n777 ), .ZN(_f_permutation__round__N2779 )
         );
  NOR2_X2 _f_permutation__round__U109  ( .A1(_f_permutation__round__c[808] ), 
        .A2(_f_permutation__round__n774 ), .ZN(_f_permutation__round__N2777 )
         );
  NOR2_X2 _f_permutation__round__U108  ( .A1(_f_permutation__round__c[809] ), 
        .A2(_f_permutation__round__n771 ), .ZN(_f_permutation__round__N2775 )
         );
  NOR2_X2 _f_permutation__round__U107  ( .A1(_f_permutation__round__c[810] ), 
        .A2(_f_permutation__round__n960 ), .ZN(_f_permutation__round__N2773 )
         );
  NOR2_X2 _f_permutation__round__U106  ( .A1(_f_permutation__round__c[811] ), 
        .A2(_f_permutation__round__n957 ), .ZN(_f_permutation__round__N2771 )
         );
  NOR2_X2 _f_permutation__round__U105  ( .A1(_f_permutation__round__c[812] ), 
        .A2(_f_permutation__round__n954 ), .ZN(_f_permutation__round__N2769 )
         );
  NOR2_X2 _f_permutation__round__U104  ( .A1(_f_permutation__round__c[813] ), 
        .A2(_f_permutation__round__n951 ), .ZN(_f_permutation__round__N2767 )
         );
  NOR2_X2 _f_permutation__round__U103  ( .A1(_f_permutation__round__c[814] ), 
        .A2(_f_permutation__round__n948 ), .ZN(_f_permutation__round__N2765 )
         );
  NOR2_X2 _f_permutation__round__U102  ( .A1(_f_permutation__round__c[815] ), 
        .A2(_f_permutation__round__n945 ), .ZN(_f_permutation__round__N2763 )
         );
  NOR2_X2 _f_permutation__round__U101  ( .A1(_f_permutation__round__c[816] ), 
        .A2(_f_permutation__round__n942 ), .ZN(_f_permutation__round__N2761 )
         );
  NOR2_X2 _f_permutation__round__U100  ( .A1(_f_permutation__round__c[817] ), 
        .A2(_f_permutation__round__n939 ), .ZN(_f_permutation__round__N2759 )
         );
  NOR2_X2 _f_permutation__round__U99  ( .A1(_f_permutation__round__c[818] ), 
        .A2(_f_permutation__round__n936 ), .ZN(_f_permutation__round__N2757 )
         );
  NOR2_X2 _f_permutation__round__U98  ( .A1(_f_permutation__round__c[819] ), 
        .A2(_f_permutation__round__n933 ), .ZN(_f_permutation__round__N2755 )
         );
  NOR2_X2 _f_permutation__round__U97  ( .A1(_f_permutation__round__c[820] ), 
        .A2(_f_permutation__round__n930 ), .ZN(_f_permutation__round__N2753 )
         );
  NOR2_X2 _f_permutation__round__U96  ( .A1(_f_permutation__round__c[821] ), 
        .A2(_f_permutation__round__n927 ), .ZN(_f_permutation__round__N2751 )
         );
  NOR2_X2 _f_permutation__round__U95  ( .A1(_f_permutation__round__c[822] ), 
        .A2(_f_permutation__round__n924 ), .ZN(_f_permutation__round__N2749 )
         );
  NOR2_X2 _f_permutation__round__U94  ( .A1(_f_permutation__round__c[823] ), 
        .A2(_f_permutation__round__n921 ), .ZN(_f_permutation__round__N2747 )
         );
  NOR2_X2 _f_permutation__round__U93  ( .A1(_f_permutation__round__c[824] ), 
        .A2(_f_permutation__round__n918 ), .ZN(_f_permutation__round__N2745 )
         );
  NOR2_X2 _f_permutation__round__U92  ( .A1(_f_permutation__round__c[825] ), 
        .A2(_f_permutation__round__n915 ), .ZN(_f_permutation__round__N2743 )
         );
  NOR2_X2 _f_permutation__round__U91  ( .A1(_f_permutation__round__c[826] ), 
        .A2(_f_permutation__round__n912 ), .ZN(_f_permutation__round__N2741 )
         );
  NOR2_X2 _f_permutation__round__U90  ( .A1(_f_permutation__round__c[827] ), 
        .A2(_f_permutation__round__n909 ), .ZN(_f_permutation__round__N2739 )
         );
  NOR2_X2 _f_permutation__round__U89  ( .A1(_f_permutation__round__c[828] ), 
        .A2(_f_permutation__round__n906 ), .ZN(_f_permutation__round__N2737 )
         );
  NOR2_X2 _f_permutation__round__U88  ( .A1(_f_permutation__round__c[829] ), 
        .A2(_f_permutation__round__n903 ), .ZN(_f_permutation__round__N2735 )
         );
  NOR2_X2 _f_permutation__round__U87  ( .A1(_f_permutation__round__c[830] ), 
        .A2(_f_permutation__round__n900 ), .ZN(_f_permutation__round__N2733 )
         );
  NOR2_X2 _f_permutation__round__U86  ( .A1(_f_permutation__round__c[831] ), 
        .A2(_f_permutation__round__n897 ), .ZN(_f_permutation__round__N2731 )
         );
  NOR2_X2 _f_permutation__round__U85  ( .A1(_f_permutation__round__c[768] ), 
        .A2(_f_permutation__round__n894 ), .ZN(_f_permutation__round__N2729 )
         );
  NOR2_X2 _f_permutation__round__U84  ( .A1(_f_permutation__round__c[769] ), 
        .A2(_f_permutation__round__n891 ), .ZN(_f_permutation__round__N2727 )
         );
  NOR2_X2 _f_permutation__round__U83  ( .A1(_f_permutation__round__c[770] ), 
        .A2(_f_permutation__round__n888 ), .ZN(_f_permutation__round__N2725 )
         );
  NOR2_X2 _f_permutation__round__U82  ( .A1(_f_permutation__round__c[771] ), 
        .A2(_f_permutation__round__n885 ), .ZN(_f_permutation__round__N2723 )
         );
  NOR2_X2 _f_permutation__round__U81  ( .A1(_f_permutation__round__c[772] ), 
        .A2(_f_permutation__round__n882 ), .ZN(_f_permutation__round__N2721 )
         );
  NOR2_X2 _f_permutation__round__U80  ( .A1(_f_permutation__round__c[773] ), 
        .A2(_f_permutation__round__n879 ), .ZN(_f_permutation__round__N2719 )
         );
  NOR2_X2 _f_permutation__round__U79  ( .A1(_f_permutation__round__c[774] ), 
        .A2(_f_permutation__round__n876 ), .ZN(_f_permutation__round__N2717 )
         );
  NOR2_X2 _f_permutation__round__U78  ( .A1(_f_permutation__round__c[775] ), 
        .A2(_f_permutation__round__n873 ), .ZN(_f_permutation__round__N2715 )
         );
  NOR2_X2 _f_permutation__round__U77  ( .A1(_f_permutation__round__c[776] ), 
        .A2(_f_permutation__round__n870 ), .ZN(_f_permutation__round__N2713 )
         );
  NOR2_X2 _f_permutation__round__U76  ( .A1(_f_permutation__round__c[777] ), 
        .A2(_f_permutation__round__n867 ), .ZN(_f_permutation__round__N2711 )
         );
  NOR2_X2 _f_permutation__round__U75  ( .A1(_f_permutation__round__c[778] ), 
        .A2(_f_permutation__round__n864 ), .ZN(_f_permutation__round__N2709 )
         );
  NOR2_X2 _f_permutation__round__U74  ( .A1(_f_permutation__round__c[779] ), 
        .A2(_f_permutation__round__n861 ), .ZN(_f_permutation__round__N2707 )
         );
  NOR2_X2 _f_permutation__round__U73  ( .A1(_f_permutation__round__c[780] ), 
        .A2(_f_permutation__round__n858 ), .ZN(_f_permutation__round__N2705 )
         );
  NOR2_X2 _f_permutation__round__U72  ( .A1(_f_permutation__round__c[781] ), 
        .A2(_f_permutation__round__n855 ), .ZN(_f_permutation__round__N2703 )
         );
  NOR2_X2 _f_permutation__round__U71  ( .A1(_f_permutation__round__c[782] ), 
        .A2(_f_permutation__round__n852 ), .ZN(_f_permutation__round__N2701 )
         );
  NOR2_X2 _f_permutation__round__U70  ( .A1(_f_permutation__round__c[783] ), 
        .A2(_f_permutation__round__n849 ), .ZN(_f_permutation__round__N2699 )
         );
  NOR2_X2 _f_permutation__round__U69  ( .A1(_f_permutation__round__c[784] ), 
        .A2(_f_permutation__round__n846 ), .ZN(_f_permutation__round__N2697 )
         );
  NOR2_X2 _f_permutation__round__U68  ( .A1(_f_permutation__round__c[785] ), 
        .A2(_f_permutation__round__n843 ), .ZN(_f_permutation__round__N2695 )
         );
  NOR2_X2 _f_permutation__round__U67  ( .A1(_f_permutation__round__c[786] ), 
        .A2(_f_permutation__round__n840 ), .ZN(_f_permutation__round__N2693 )
         );
  NOR2_X2 _f_permutation__round__U66  ( .A1(_f_permutation__round__c[787] ), 
        .A2(_f_permutation__round__n837 ), .ZN(_f_permutation__round__N2691 )
         );
  NOR2_X2 _f_permutation__round__U65  ( .A1(_f_permutation__round__c[788] ), 
        .A2(_f_permutation__round__n834 ), .ZN(_f_permutation__round__N2689 )
         );
  INV_X4 _f_permutation__round__U2560  ( .A(_f_permutation__round__c[1152] ), 
        .ZN(_f_permutation__round__n960 ) );
  INV_X4 _f_permutation__round__U2559  ( .A(_f_permutation__round__c[1088] ), 
        .ZN(_f_permutation__round__n959 ) );
  INV_X4 _f_permutation__round__U2558  ( .A(_f_permutation__round__c[960] ), 
        .ZN(_f_permutation__round__n958 ) );
  INV_X4 _f_permutation__round__U2557  ( .A(_f_permutation__round__c[1153] ), 
        .ZN(_f_permutation__round__n957 ) );
  INV_X4 _f_permutation__round__U2556  ( .A(_f_permutation__round__c[1089] ), 
        .ZN(_f_permutation__round__n956 ) );
  INV_X4 _f_permutation__round__U2555  ( .A(_f_permutation__round__c[961] ), 
        .ZN(_f_permutation__round__n955 ) );
  INV_X4 _f_permutation__round__U2554  ( .A(_f_permutation__round__c[1154] ), 
        .ZN(_f_permutation__round__n954 ) );
  INV_X4 _f_permutation__round__U2553  ( .A(_f_permutation__round__c[1090] ), 
        .ZN(_f_permutation__round__n953 ) );
  INV_X4 _f_permutation__round__U2552  ( .A(_f_permutation__round__c[962] ), 
        .ZN(_f_permutation__round__n952 ) );
  INV_X4 _f_permutation__round__U2551  ( .A(_f_permutation__round__c[1155] ), 
        .ZN(_f_permutation__round__n951 ) );
  INV_X4 _f_permutation__round__U2550  ( .A(_f_permutation__round__c[1091] ), 
        .ZN(_f_permutation__round__n950 ) );
  INV_X4 _f_permutation__round__U2549  ( .A(_f_permutation__round__c[963] ), 
        .ZN(_f_permutation__round__n949 ) );
  INV_X4 _f_permutation__round__U2548  ( .A(_f_permutation__round__c[1156] ), 
        .ZN(_f_permutation__round__n948 ) );
  INV_X4 _f_permutation__round__U2547  ( .A(_f_permutation__round__c[1092] ), 
        .ZN(_f_permutation__round__n947 ) );
  INV_X4 _f_permutation__round__U2546  ( .A(_f_permutation__round__c[964] ), 
        .ZN(_f_permutation__round__n946 ) );
  INV_X4 _f_permutation__round__U2545  ( .A(_f_permutation__round__c[1157] ), 
        .ZN(_f_permutation__round__n945 ) );
  INV_X4 _f_permutation__round__U2544  ( .A(_f_permutation__round__c[1093] ), 
        .ZN(_f_permutation__round__n944 ) );
  INV_X4 _f_permutation__round__U2543  ( .A(_f_permutation__round__c[965] ), 
        .ZN(_f_permutation__round__n943 ) );
  INV_X4 _f_permutation__round__U2542  ( .A(_f_permutation__round__c[1158] ), 
        .ZN(_f_permutation__round__n942 ) );
  INV_X4 _f_permutation__round__U2541  ( .A(_f_permutation__round__c[1094] ), 
        .ZN(_f_permutation__round__n941 ) );
  INV_X4 _f_permutation__round__U2540  ( .A(_f_permutation__round__c[966] ), 
        .ZN(_f_permutation__round__n940 ) );
  INV_X4 _f_permutation__round__U2539  ( .A(_f_permutation__round__c[1159] ), 
        .ZN(_f_permutation__round__n939 ) );
  INV_X4 _f_permutation__round__U2538  ( .A(_f_permutation__round__c[1095] ), 
        .ZN(_f_permutation__round__n938 ) );
  INV_X4 _f_permutation__round__U2537  ( .A(_f_permutation__round__c[967] ), 
        .ZN(_f_permutation__round__n937 ) );
  INV_X4 _f_permutation__round__U2536  ( .A(_f_permutation__round__c[1160] ), 
        .ZN(_f_permutation__round__n936 ) );
  INV_X4 _f_permutation__round__U2535  ( .A(_f_permutation__round__c[1096] ), 
        .ZN(_f_permutation__round__n935 ) );
  INV_X4 _f_permutation__round__U2534  ( .A(_f_permutation__round__c[968] ), 
        .ZN(_f_permutation__round__n934 ) );
  INV_X4 _f_permutation__round__U2533  ( .A(_f_permutation__round__c[1161] ), 
        .ZN(_f_permutation__round__n933 ) );
  INV_X4 _f_permutation__round__U2532  ( .A(_f_permutation__round__c[1097] ), 
        .ZN(_f_permutation__round__n932 ) );
  INV_X4 _f_permutation__round__U2531  ( .A(_f_permutation__round__c[969] ), 
        .ZN(_f_permutation__round__n931 ) );
  INV_X4 _f_permutation__round__U2530  ( .A(_f_permutation__round__c[1162] ), 
        .ZN(_f_permutation__round__n930 ) );
  INV_X4 _f_permutation__round__U2529  ( .A(_f_permutation__round__c[1098] ), 
        .ZN(_f_permutation__round__n929 ) );
  INV_X4 _f_permutation__round__U2528  ( .A(_f_permutation__round__c[970] ), 
        .ZN(_f_permutation__round__n928 ) );
  INV_X4 _f_permutation__round__U2527  ( .A(_f_permutation__round__c[1163] ), 
        .ZN(_f_permutation__round__n927 ) );
  INV_X4 _f_permutation__round__U2526  ( .A(_f_permutation__round__c[1099] ), 
        .ZN(_f_permutation__round__n926 ) );
  INV_X4 _f_permutation__round__U2525  ( .A(_f_permutation__round__c[971] ), 
        .ZN(_f_permutation__round__n925 ) );
  INV_X4 _f_permutation__round__U2524  ( .A(_f_permutation__round__c[1164] ), 
        .ZN(_f_permutation__round__n924 ) );
  INV_X4 _f_permutation__round__U2523  ( .A(_f_permutation__round__c[1100] ), 
        .ZN(_f_permutation__round__n923 ) );
  INV_X4 _f_permutation__round__U2522  ( .A(_f_permutation__round__c[972] ), 
        .ZN(_f_permutation__round__n922 ) );
  INV_X4 _f_permutation__round__U2521  ( .A(_f_permutation__round__c[1165] ), 
        .ZN(_f_permutation__round__n921 ) );
  INV_X4 _f_permutation__round__U2520  ( .A(_f_permutation__round__c[1101] ), 
        .ZN(_f_permutation__round__n920 ) );
  INV_X4 _f_permutation__round__U2519  ( .A(_f_permutation__round__c[973] ), 
        .ZN(_f_permutation__round__n919 ) );
  INV_X4 _f_permutation__round__U2518  ( .A(_f_permutation__round__c[1166] ), 
        .ZN(_f_permutation__round__n918 ) );
  INV_X4 _f_permutation__round__U2517  ( .A(_f_permutation__round__c[1102] ), 
        .ZN(_f_permutation__round__n917 ) );
  INV_X4 _f_permutation__round__U2516  ( .A(_f_permutation__round__c[974] ), 
        .ZN(_f_permutation__round__n916 ) );
  INV_X4 _f_permutation__round__U2515  ( .A(_f_permutation__round__c[1167] ), 
        .ZN(_f_permutation__round__n915 ) );
  INV_X4 _f_permutation__round__U2514  ( .A(_f_permutation__round__c[1103] ), 
        .ZN(_f_permutation__round__n914 ) );
  INV_X4 _f_permutation__round__U2513  ( .A(_f_permutation__round__c[975] ), 
        .ZN(_f_permutation__round__n913 ) );
  INV_X4 _f_permutation__round__U2512  ( .A(_f_permutation__round__c[1168] ), 
        .ZN(_f_permutation__round__n912 ) );
  INV_X4 _f_permutation__round__U2511  ( .A(_f_permutation__round__c[1104] ), 
        .ZN(_f_permutation__round__n911 ) );
  INV_X4 _f_permutation__round__U2510  ( .A(_f_permutation__round__c[976] ), 
        .ZN(_f_permutation__round__n910 ) );
  INV_X4 _f_permutation__round__U2509  ( .A(_f_permutation__round__c[1169] ), 
        .ZN(_f_permutation__round__n909 ) );
  INV_X4 _f_permutation__round__U2508  ( .A(_f_permutation__round__c[1105] ), 
        .ZN(_f_permutation__round__n908 ) );
  INV_X4 _f_permutation__round__U2507  ( .A(_f_permutation__round__c[977] ), 
        .ZN(_f_permutation__round__n907 ) );
  INV_X4 _f_permutation__round__U2506  ( .A(_f_permutation__round__c[1170] ), 
        .ZN(_f_permutation__round__n906 ) );
  INV_X4 _f_permutation__round__U2505  ( .A(_f_permutation__round__c[1106] ), 
        .ZN(_f_permutation__round__n905 ) );
  INV_X4 _f_permutation__round__U2504  ( .A(_f_permutation__round__c[978] ), 
        .ZN(_f_permutation__round__n904 ) );
  INV_X4 _f_permutation__round__U2503  ( .A(_f_permutation__round__c[1171] ), 
        .ZN(_f_permutation__round__n903 ) );
  INV_X4 _f_permutation__round__U2502  ( .A(_f_permutation__round__c[1107] ), 
        .ZN(_f_permutation__round__n902 ) );
  INV_X4 _f_permutation__round__U2501  ( .A(_f_permutation__round__c[979] ), 
        .ZN(_f_permutation__round__n901 ) );
  INV_X4 _f_permutation__round__U2500  ( .A(_f_permutation__round__c[1172] ), 
        .ZN(_f_permutation__round__n900 ) );
  INV_X4 _f_permutation__round__U2499  ( .A(_f_permutation__round__c[1108] ), 
        .ZN(_f_permutation__round__n899 ) );
  INV_X4 _f_permutation__round__U2498  ( .A(_f_permutation__round__c[980] ), 
        .ZN(_f_permutation__round__n898 ) );
  INV_X4 _f_permutation__round__U2497  ( .A(_f_permutation__round__c[1173] ), 
        .ZN(_f_permutation__round__n897 ) );
  INV_X4 _f_permutation__round__U2496  ( .A(_f_permutation__round__c[1109] ), 
        .ZN(_f_permutation__round__n896 ) );
  INV_X4 _f_permutation__round__U2495  ( .A(_f_permutation__round__c[981] ), 
        .ZN(_f_permutation__round__n895 ) );
  INV_X4 _f_permutation__round__U2494  ( .A(_f_permutation__round__c[1174] ), 
        .ZN(_f_permutation__round__n894 ) );
  INV_X4 _f_permutation__round__U2493  ( .A(_f_permutation__round__c[1110] ), 
        .ZN(_f_permutation__round__n893 ) );
  INV_X4 _f_permutation__round__U2492  ( .A(_f_permutation__round__c[982] ), 
        .ZN(_f_permutation__round__n892 ) );
  INV_X4 _f_permutation__round__U2491  ( .A(_f_permutation__round__c[1175] ), 
        .ZN(_f_permutation__round__n891 ) );
  INV_X4 _f_permutation__round__U2490  ( .A(_f_permutation__round__c[1111] ), 
        .ZN(_f_permutation__round__n890 ) );
  INV_X4 _f_permutation__round__U2489  ( .A(_f_permutation__round__c[983] ), 
        .ZN(_f_permutation__round__n889 ) );
  INV_X4 _f_permutation__round__U2488  ( .A(_f_permutation__round__c[1176] ), 
        .ZN(_f_permutation__round__n888 ) );
  INV_X4 _f_permutation__round__U2487  ( .A(_f_permutation__round__c[1112] ), 
        .ZN(_f_permutation__round__n887 ) );
  INV_X4 _f_permutation__round__U2486  ( .A(_f_permutation__round__c[984] ), 
        .ZN(_f_permutation__round__n886 ) );
  INV_X4 _f_permutation__round__U2485  ( .A(_f_permutation__round__c[1177] ), 
        .ZN(_f_permutation__round__n885 ) );
  INV_X4 _f_permutation__round__U2484  ( .A(_f_permutation__round__c[1113] ), 
        .ZN(_f_permutation__round__n884 ) );
  INV_X4 _f_permutation__round__U2483  ( .A(_f_permutation__round__c[985] ), 
        .ZN(_f_permutation__round__n883 ) );
  INV_X4 _f_permutation__round__U2482  ( .A(_f_permutation__round__c[1178] ), 
        .ZN(_f_permutation__round__n882 ) );
  INV_X4 _f_permutation__round__U2481  ( .A(_f_permutation__round__c[1114] ), 
        .ZN(_f_permutation__round__n881 ) );
  INV_X4 _f_permutation__round__U2480  ( .A(_f_permutation__round__c[986] ), 
        .ZN(_f_permutation__round__n880 ) );
  INV_X4 _f_permutation__round__U2479  ( .A(_f_permutation__round__c[1179] ), 
        .ZN(_f_permutation__round__n879 ) );
  INV_X4 _f_permutation__round__U2478  ( .A(_f_permutation__round__c[1115] ), 
        .ZN(_f_permutation__round__n878 ) );
  INV_X4 _f_permutation__round__U2477  ( .A(_f_permutation__round__c[987] ), 
        .ZN(_f_permutation__round__n877 ) );
  INV_X4 _f_permutation__round__U2476  ( .A(_f_permutation__round__c[1180] ), 
        .ZN(_f_permutation__round__n876 ) );
  INV_X4 _f_permutation__round__U2475  ( .A(_f_permutation__round__c[1116] ), 
        .ZN(_f_permutation__round__n875 ) );
  INV_X4 _f_permutation__round__U2474  ( .A(_f_permutation__round__c[988] ), 
        .ZN(_f_permutation__round__n874 ) );
  INV_X4 _f_permutation__round__U2473  ( .A(_f_permutation__round__c[1181] ), 
        .ZN(_f_permutation__round__n873 ) );
  INV_X4 _f_permutation__round__U2472  ( .A(_f_permutation__round__c[1117] ), 
        .ZN(_f_permutation__round__n872 ) );
  INV_X4 _f_permutation__round__U2471  ( .A(_f_permutation__round__c[989] ), 
        .ZN(_f_permutation__round__n871 ) );
  INV_X4 _f_permutation__round__U2470  ( .A(_f_permutation__round__c[1182] ), 
        .ZN(_f_permutation__round__n870 ) );
  INV_X4 _f_permutation__round__U2469  ( .A(_f_permutation__round__c[1118] ), 
        .ZN(_f_permutation__round__n869 ) );
  INV_X4 _f_permutation__round__U2468  ( .A(_f_permutation__round__c[990] ), 
        .ZN(_f_permutation__round__n868 ) );
  INV_X4 _f_permutation__round__U2467  ( .A(_f_permutation__round__c[1183] ), 
        .ZN(_f_permutation__round__n867 ) );
  INV_X4 _f_permutation__round__U2466  ( .A(_f_permutation__round__c[1119] ), 
        .ZN(_f_permutation__round__n866 ) );
  INV_X4 _f_permutation__round__U2465  ( .A(_f_permutation__round__c[991] ), 
        .ZN(_f_permutation__round__n865 ) );
  INV_X4 _f_permutation__round__U2464  ( .A(_f_permutation__round__c[1184] ), 
        .ZN(_f_permutation__round__n864 ) );
  INV_X4 _f_permutation__round__U2463  ( .A(_f_permutation__round__c[1120] ), 
        .ZN(_f_permutation__round__n863 ) );
  INV_X4 _f_permutation__round__U2462  ( .A(_f_permutation__round__c[992] ), 
        .ZN(_f_permutation__round__n862 ) );
  INV_X4 _f_permutation__round__U2461  ( .A(_f_permutation__round__c[1185] ), 
        .ZN(_f_permutation__round__n861 ) );
  INV_X4 _f_permutation__round__U2460  ( .A(_f_permutation__round__c[1121] ), 
        .ZN(_f_permutation__round__n860 ) );
  INV_X4 _f_permutation__round__U2459  ( .A(_f_permutation__round__c[993] ), 
        .ZN(_f_permutation__round__n859 ) );
  INV_X4 _f_permutation__round__U2458  ( .A(_f_permutation__round__c[1186] ), 
        .ZN(_f_permutation__round__n858 ) );
  INV_X4 _f_permutation__round__U2457  ( .A(_f_permutation__round__c[1122] ), 
        .ZN(_f_permutation__round__n857 ) );
  INV_X4 _f_permutation__round__U2456  ( .A(_f_permutation__round__c[994] ), 
        .ZN(_f_permutation__round__n856 ) );
  INV_X4 _f_permutation__round__U2455  ( .A(_f_permutation__round__c[1187] ), 
        .ZN(_f_permutation__round__n855 ) );
  INV_X4 _f_permutation__round__U2454  ( .A(_f_permutation__round__c[1123] ), 
        .ZN(_f_permutation__round__n854 ) );
  INV_X4 _f_permutation__round__U2453  ( .A(_f_permutation__round__c[995] ), 
        .ZN(_f_permutation__round__n853 ) );
  INV_X4 _f_permutation__round__U2452  ( .A(_f_permutation__round__c[1188] ), 
        .ZN(_f_permutation__round__n852 ) );
  INV_X4 _f_permutation__round__U2451  ( .A(_f_permutation__round__c[1124] ), 
        .ZN(_f_permutation__round__n851 ) );
  INV_X4 _f_permutation__round__U2450  ( .A(_f_permutation__round__c[996] ), 
        .ZN(_f_permutation__round__n850 ) );
  INV_X4 _f_permutation__round__U2449  ( .A(_f_permutation__round__c[1189] ), 
        .ZN(_f_permutation__round__n849 ) );
  INV_X4 _f_permutation__round__U2448  ( .A(_f_permutation__round__c[1125] ), 
        .ZN(_f_permutation__round__n848 ) );
  INV_X4 _f_permutation__round__U2447  ( .A(_f_permutation__round__c[997] ), 
        .ZN(_f_permutation__round__n847 ) );
  INV_X4 _f_permutation__round__U2446  ( .A(_f_permutation__round__c[1190] ), 
        .ZN(_f_permutation__round__n846 ) );
  INV_X4 _f_permutation__round__U2445  ( .A(_f_permutation__round__c[1126] ), 
        .ZN(_f_permutation__round__n845 ) );
  INV_X4 _f_permutation__round__U2444  ( .A(_f_permutation__round__c[998] ), 
        .ZN(_f_permutation__round__n844 ) );
  INV_X4 _f_permutation__round__U2443  ( .A(_f_permutation__round__c[1191] ), 
        .ZN(_f_permutation__round__n843 ) );
  INV_X4 _f_permutation__round__U2442  ( .A(_f_permutation__round__c[1127] ), 
        .ZN(_f_permutation__round__n842 ) );
  INV_X4 _f_permutation__round__U2441  ( .A(_f_permutation__round__c[999] ), 
        .ZN(_f_permutation__round__n841 ) );
  INV_X4 _f_permutation__round__U2440  ( .A(_f_permutation__round__c[1192] ), 
        .ZN(_f_permutation__round__n840 ) );
  INV_X4 _f_permutation__round__U2439  ( .A(_f_permutation__round__c[1128] ), 
        .ZN(_f_permutation__round__n839 ) );
  INV_X4 _f_permutation__round__U2438  ( .A(_f_permutation__round__c[1000] ), 
        .ZN(_f_permutation__round__n838 ) );
  INV_X4 _f_permutation__round__U2437  ( .A(_f_permutation__round__c[1193] ), 
        .ZN(_f_permutation__round__n837 ) );
  INV_X4 _f_permutation__round__U2436  ( .A(_f_permutation__round__c[1129] ), 
        .ZN(_f_permutation__round__n836 ) );
  INV_X4 _f_permutation__round__U2435  ( .A(_f_permutation__round__c[1001] ), 
        .ZN(_f_permutation__round__n835 ) );
  INV_X4 _f_permutation__round__U2434  ( .A(_f_permutation__round__c[1194] ), 
        .ZN(_f_permutation__round__n834 ) );
  INV_X4 _f_permutation__round__U2433  ( .A(_f_permutation__round__c[1130] ), 
        .ZN(_f_permutation__round__n833 ) );
  INV_X4 _f_permutation__round__U2432  ( .A(_f_permutation__round__c[1002] ), 
        .ZN(_f_permutation__round__n832 ) );
  INV_X4 _f_permutation__round__U2431  ( .A(_f_permutation__round__c[1195] ), 
        .ZN(_f_permutation__round__n831 ) );
  INV_X4 _f_permutation__round__U2430  ( .A(_f_permutation__round__c[1131] ), 
        .ZN(_f_permutation__round__n830 ) );
  INV_X4 _f_permutation__round__U2429  ( .A(_f_permutation__round__c[1003] ), 
        .ZN(_f_permutation__round__n829 ) );
  INV_X4 _f_permutation__round__U2428  ( .A(_f_permutation__round__c[1196] ), 
        .ZN(_f_permutation__round__n828 ) );
  INV_X4 _f_permutation__round__U2427  ( .A(_f_permutation__round__c[1132] ), 
        .ZN(_f_permutation__round__n827 ) );
  INV_X4 _f_permutation__round__U2426  ( .A(_f_permutation__round__c[1004] ), 
        .ZN(_f_permutation__round__n826 ) );
  INV_X4 _f_permutation__round__U2425  ( .A(_f_permutation__round__c[1197] ), 
        .ZN(_f_permutation__round__n825 ) );
  INV_X4 _f_permutation__round__U2424  ( .A(_f_permutation__round__c[1133] ), 
        .ZN(_f_permutation__round__n824 ) );
  INV_X4 _f_permutation__round__U2423  ( .A(_f_permutation__round__c[1005] ), 
        .ZN(_f_permutation__round__n823 ) );
  INV_X4 _f_permutation__round__U2422  ( .A(_f_permutation__round__c[1198] ), 
        .ZN(_f_permutation__round__n822 ) );
  INV_X4 _f_permutation__round__U2421  ( .A(_f_permutation__round__c[1134] ), 
        .ZN(_f_permutation__round__n821 ) );
  INV_X4 _f_permutation__round__U2420  ( .A(_f_permutation__round__c[1006] ), 
        .ZN(_f_permutation__round__n820 ) );
  INV_X4 _f_permutation__round__U2419  ( .A(_f_permutation__round__c[1199] ), 
        .ZN(_f_permutation__round__n819 ) );
  INV_X4 _f_permutation__round__U2418  ( .A(_f_permutation__round__c[1135] ), 
        .ZN(_f_permutation__round__n818 ) );
  INV_X4 _f_permutation__round__U2417  ( .A(_f_permutation__round__c[1007] ), 
        .ZN(_f_permutation__round__n817 ) );
  INV_X4 _f_permutation__round__U2416  ( .A(_f_permutation__round__c[1200] ), 
        .ZN(_f_permutation__round__n816 ) );
  INV_X4 _f_permutation__round__U2415  ( .A(_f_permutation__round__c[1136] ), 
        .ZN(_f_permutation__round__n815 ) );
  INV_X4 _f_permutation__round__U2414  ( .A(_f_permutation__round__c[1008] ), 
        .ZN(_f_permutation__round__n814 ) );
  INV_X4 _f_permutation__round__U2413  ( .A(_f_permutation__round__c[1201] ), 
        .ZN(_f_permutation__round__n813 ) );
  INV_X4 _f_permutation__round__U2412  ( .A(_f_permutation__round__c[1137] ), 
        .ZN(_f_permutation__round__n812 ) );
  INV_X4 _f_permutation__round__U2411  ( .A(_f_permutation__round__c[1009] ), 
        .ZN(_f_permutation__round__n811 ) );
  INV_X4 _f_permutation__round__U2410  ( .A(_f_permutation__round__c[1202] ), 
        .ZN(_f_permutation__round__n810 ) );
  INV_X4 _f_permutation__round__U2409  ( .A(_f_permutation__round__c[1138] ), 
        .ZN(_f_permutation__round__n809 ) );
  INV_X4 _f_permutation__round__U2408  ( .A(_f_permutation__round__c[1010] ), 
        .ZN(_f_permutation__round__n808 ) );
  INV_X4 _f_permutation__round__U2407  ( .A(_f_permutation__round__c[1203] ), 
        .ZN(_f_permutation__round__n807 ) );
  INV_X4 _f_permutation__round__U2406  ( .A(_f_permutation__round__c[1139] ), 
        .ZN(_f_permutation__round__n806 ) );
  INV_X4 _f_permutation__round__U2405  ( .A(_f_permutation__round__c[1011] ), 
        .ZN(_f_permutation__round__n805 ) );
  INV_X4 _f_permutation__round__U2404  ( .A(_f_permutation__round__c[1204] ), 
        .ZN(_f_permutation__round__n804 ) );
  INV_X4 _f_permutation__round__U2403  ( .A(_f_permutation__round__c[1140] ), 
        .ZN(_f_permutation__round__n803 ) );
  INV_X4 _f_permutation__round__U2402  ( .A(_f_permutation__round__c[1012] ), 
        .ZN(_f_permutation__round__n802 ) );
  INV_X4 _f_permutation__round__U2401  ( .A(_f_permutation__round__c[1205] ), 
        .ZN(_f_permutation__round__n801 ) );
  INV_X4 _f_permutation__round__U2400  ( .A(_f_permutation__round__c[1141] ), 
        .ZN(_f_permutation__round__n800 ) );
  INV_X4 _f_permutation__round__U2399  ( .A(_f_permutation__round__c[1013] ), 
        .ZN(_f_permutation__round__n799 ) );
  INV_X4 _f_permutation__round__U2398  ( .A(_f_permutation__round__c[1206] ), 
        .ZN(_f_permutation__round__n798 ) );
  INV_X4 _f_permutation__round__U2397  ( .A(_f_permutation__round__c[1142] ), 
        .ZN(_f_permutation__round__n797 ) );
  INV_X4 _f_permutation__round__U2396  ( .A(_f_permutation__round__c[1014] ), 
        .ZN(_f_permutation__round__n796 ) );
  INV_X4 _f_permutation__round__U2395  ( .A(_f_permutation__round__c[1207] ), 
        .ZN(_f_permutation__round__n795 ) );
  INV_X4 _f_permutation__round__U2394  ( .A(_f_permutation__round__c[1143] ), 
        .ZN(_f_permutation__round__n794 ) );
  INV_X4 _f_permutation__round__U2393  ( .A(_f_permutation__round__c[1015] ), 
        .ZN(_f_permutation__round__n793 ) );
  INV_X4 _f_permutation__round__U2392  ( .A(_f_permutation__round__c[1208] ), 
        .ZN(_f_permutation__round__n792 ) );
  INV_X4 _f_permutation__round__U2391  ( .A(_f_permutation__round__c[1144] ), 
        .ZN(_f_permutation__round__n791 ) );
  INV_X4 _f_permutation__round__U2390  ( .A(_f_permutation__round__c[1016] ), 
        .ZN(_f_permutation__round__n790 ) );
  INV_X4 _f_permutation__round__U2389  ( .A(_f_permutation__round__c[1209] ), 
        .ZN(_f_permutation__round__n789 ) );
  INV_X4 _f_permutation__round__U2388  ( .A(_f_permutation__round__c[1145] ), 
        .ZN(_f_permutation__round__n788 ) );
  INV_X4 _f_permutation__round__U2387  ( .A(_f_permutation__round__c[1017] ), 
        .ZN(_f_permutation__round__n787 ) );
  INV_X4 _f_permutation__round__U2386  ( .A(_f_permutation__round__c[1210] ), 
        .ZN(_f_permutation__round__n786 ) );
  INV_X4 _f_permutation__round__U2385  ( .A(_f_permutation__round__c[1146] ), 
        .ZN(_f_permutation__round__n785 ) );
  INV_X4 _f_permutation__round__U2384  ( .A(_f_permutation__round__c[1018] ), 
        .ZN(_f_permutation__round__n784 ) );
  INV_X4 _f_permutation__round__U2383  ( .A(_f_permutation__round__c[1211] ), 
        .ZN(_f_permutation__round__n783 ) );
  INV_X4 _f_permutation__round__U2382  ( .A(_f_permutation__round__c[1147] ), 
        .ZN(_f_permutation__round__n782 ) );
  INV_X4 _f_permutation__round__U2381  ( .A(_f_permutation__round__c[1019] ), 
        .ZN(_f_permutation__round__n781 ) );
  INV_X4 _f_permutation__round__U2380  ( .A(_f_permutation__round__c[1212] ), 
        .ZN(_f_permutation__round__n780 ) );
  INV_X4 _f_permutation__round__U2379  ( .A(_f_permutation__round__c[1148] ), 
        .ZN(_f_permutation__round__n779 ) );
  INV_X4 _f_permutation__round__U2378  ( .A(_f_permutation__round__c[1020] ), 
        .ZN(_f_permutation__round__n778 ) );
  INV_X4 _f_permutation__round__U2377  ( .A(_f_permutation__round__c[1213] ), 
        .ZN(_f_permutation__round__n777 ) );
  INV_X4 _f_permutation__round__U2376  ( .A(_f_permutation__round__c[1149] ), 
        .ZN(_f_permutation__round__n776 ) );
  INV_X4 _f_permutation__round__U2375  ( .A(_f_permutation__round__c[1021] ), 
        .ZN(_f_permutation__round__n775 ) );
  INV_X4 _f_permutation__round__U2374  ( .A(_f_permutation__round__c[1214] ), 
        .ZN(_f_permutation__round__n774 ) );
  INV_X4 _f_permutation__round__U2373  ( .A(_f_permutation__round__c[1150] ), 
        .ZN(_f_permutation__round__n773 ) );
  INV_X4 _f_permutation__round__U2372  ( .A(_f_permutation__round__c[1022] ), 
        .ZN(_f_permutation__round__n772 ) );
  INV_X4 _f_permutation__round__U2371  ( .A(_f_permutation__round__c[1215] ), 
        .ZN(_f_permutation__round__n771 ) );
  INV_X4 _f_permutation__round__U2370  ( .A(_f_permutation__round__c[1151] ), 
        .ZN(_f_permutation__round__n770 ) );
  INV_X4 _f_permutation__round__U2369  ( .A(_f_permutation__round__c[1023] ), 
        .ZN(_f_permutation__round__n769 ) );
  INV_X4 _f_permutation__round__U2368  ( .A(_f_permutation__round__c[193] ), 
        .ZN(_f_permutation__round__n768 ) );
  INV_X4 _f_permutation__round__U2367  ( .A(_f_permutation__round__c[129] ), 
        .ZN(_f_permutation__round__n767 ) );
  INV_X4 _f_permutation__round__U2366  ( .A(_f_permutation__round__c[832] ), 
        .ZN(_f_permutation__round__n766 ) );
  INV_X4 _f_permutation__round__U2365  ( .A(_f_permutation__round__c[768] ), 
        .ZN(_f_permutation__round__n765 ) );
  INV_X4 _f_permutation__round__U2364  ( .A(_f_permutation__round__c[640] ), 
        .ZN(_f_permutation__round__n764 ) );
  INV_X4 _f_permutation__round__U2363  ( .A(_f_permutation__round__c[194] ), 
        .ZN(_f_permutation__round__n763 ) );
  INV_X4 _f_permutation__round__U2362  ( .A(_f_permutation__round__c[130] ), 
        .ZN(_f_permutation__round__n762 ) );
  INV_X4 _f_permutation__round__U2361  ( .A(_f_permutation__round__c[833] ), 
        .ZN(_f_permutation__round__n761 ) );
  INV_X4 _f_permutation__round__U2360  ( .A(_f_permutation__round__c[769] ), 
        .ZN(_f_permutation__round__n760 ) );
  INV_X4 _f_permutation__round__U2359  ( .A(_f_permutation__round__c[641] ), 
        .ZN(_f_permutation__round__n759 ) );
  INV_X4 _f_permutation__round__U2358  ( .A(_f_permutation__round__c[195] ), 
        .ZN(_f_permutation__round__n758 ) );
  INV_X4 _f_permutation__round__U2357  ( .A(_f_permutation__round__c[131] ), 
        .ZN(_f_permutation__round__n757 ) );
  INV_X4 _f_permutation__round__U2356  ( .A(_f_permutation__round__c[834] ), 
        .ZN(_f_permutation__round__n756 ) );
  INV_X4 _f_permutation__round__U2355  ( .A(_f_permutation__round__c[770] ), 
        .ZN(_f_permutation__round__n755 ) );
  INV_X4 _f_permutation__round__U2354  ( .A(_f_permutation__round__c[642] ), 
        .ZN(_f_permutation__round__n754 ) );
  INV_X4 _f_permutation__round__U2353  ( .A(_f_permutation__round__c[196] ), 
        .ZN(_f_permutation__round__n753 ) );
  INV_X4 _f_permutation__round__U2352  ( .A(_f_permutation__round__c[132] ), 
        .ZN(_f_permutation__round__n752 ) );
  INV_X4 _f_permutation__round__U2351  ( .A(_f_permutation__round__c[835] ), 
        .ZN(_f_permutation__round__n751 ) );
  INV_X4 _f_permutation__round__U2350  ( .A(_f_permutation__round__c[771] ), 
        .ZN(_f_permutation__round__n750 ) );
  INV_X4 _f_permutation__round__U2349  ( .A(_f_permutation__round__c[643] ), 
        .ZN(_f_permutation__round__n749 ) );
  INV_X4 _f_permutation__round__U2348  ( .A(_f_permutation__round__c[197] ), 
        .ZN(_f_permutation__round__n748 ) );
  INV_X4 _f_permutation__round__U2347  ( .A(_f_permutation__round__c[133] ), 
        .ZN(_f_permutation__round__n747 ) );
  INV_X4 _f_permutation__round__U2346  ( .A(_f_permutation__round__c[836] ), 
        .ZN(_f_permutation__round__n746 ) );
  INV_X4 _f_permutation__round__U2345  ( .A(_f_permutation__round__c[772] ), 
        .ZN(_f_permutation__round__n745 ) );
  INV_X4 _f_permutation__round__U2344  ( .A(_f_permutation__round__c[644] ), 
        .ZN(_f_permutation__round__n744 ) );
  INV_X4 _f_permutation__round__U2343  ( .A(_f_permutation__round__c[198] ), 
        .ZN(_f_permutation__round__n743 ) );
  INV_X4 _f_permutation__round__U2342  ( .A(_f_permutation__round__c[134] ), 
        .ZN(_f_permutation__round__n742 ) );
  INV_X4 _f_permutation__round__U2341  ( .A(_f_permutation__round__c[837] ), 
        .ZN(_f_permutation__round__n741 ) );
  INV_X4 _f_permutation__round__U2340  ( .A(_f_permutation__round__c[773] ), 
        .ZN(_f_permutation__round__n740 ) );
  INV_X4 _f_permutation__round__U2339  ( .A(_f_permutation__round__c[645] ), 
        .ZN(_f_permutation__round__n739 ) );
  INV_X4 _f_permutation__round__U2338  ( .A(_f_permutation__round__c[199] ), 
        .ZN(_f_permutation__round__n738 ) );
  INV_X4 _f_permutation__round__U2337  ( .A(_f_permutation__round__c[135] ), 
        .ZN(_f_permutation__round__n737 ) );
  INV_X4 _f_permutation__round__U2336  ( .A(_f_permutation__round__c[838] ), 
        .ZN(_f_permutation__round__n736 ) );
  INV_X4 _f_permutation__round__U2335  ( .A(_f_permutation__round__c[774] ), 
        .ZN(_f_permutation__round__n735 ) );
  INV_X4 _f_permutation__round__U2334  ( .A(_f_permutation__round__c[646] ), 
        .ZN(_f_permutation__round__n734 ) );
  INV_X4 _f_permutation__round__U2333  ( .A(_f_permutation__round__c[200] ), 
        .ZN(_f_permutation__round__n733 ) );
  INV_X4 _f_permutation__round__U2332  ( .A(_f_permutation__round__c[136] ), 
        .ZN(_f_permutation__round__n732 ) );
  INV_X4 _f_permutation__round__U2331  ( .A(_f_permutation__round__c[839] ), 
        .ZN(_f_permutation__round__n731 ) );
  INV_X4 _f_permutation__round__U2330  ( .A(_f_permutation__round__c[775] ), 
        .ZN(_f_permutation__round__n730 ) );
  INV_X4 _f_permutation__round__U2329  ( .A(_f_permutation__round__c[647] ), 
        .ZN(_f_permutation__round__n729 ) );
  INV_X4 _f_permutation__round__U2328  ( .A(_f_permutation__round__c[201] ), 
        .ZN(_f_permutation__round__n728 ) );
  INV_X4 _f_permutation__round__U2327  ( .A(_f_permutation__round__c[137] ), 
        .ZN(_f_permutation__round__n727 ) );
  INV_X4 _f_permutation__round__U2326  ( .A(_f_permutation__round__c[840] ), 
        .ZN(_f_permutation__round__n726 ) );
  INV_X4 _f_permutation__round__U2325  ( .A(_f_permutation__round__c[776] ), 
        .ZN(_f_permutation__round__n725 ) );
  INV_X4 _f_permutation__round__U2324  ( .A(_f_permutation__round__c[648] ), 
        .ZN(_f_permutation__round__n724 ) );
  INV_X4 _f_permutation__round__U2323  ( .A(_f_permutation__round__c[202] ), 
        .ZN(_f_permutation__round__n723 ) );
  INV_X4 _f_permutation__round__U2322  ( .A(_f_permutation__round__c[138] ), 
        .ZN(_f_permutation__round__n722 ) );
  INV_X4 _f_permutation__round__U2321  ( .A(_f_permutation__round__c[841] ), 
        .ZN(_f_permutation__round__n721 ) );
  INV_X4 _f_permutation__round__U2320  ( .A(_f_permutation__round__c[777] ), 
        .ZN(_f_permutation__round__n720 ) );
  INV_X4 _f_permutation__round__U2319  ( .A(_f_permutation__round__c[649] ), 
        .ZN(_f_permutation__round__n719 ) );
  INV_X4 _f_permutation__round__U2318  ( .A(_f_permutation__round__c[203] ), 
        .ZN(_f_permutation__round__n718 ) );
  INV_X4 _f_permutation__round__U2317  ( .A(_f_permutation__round__c[139] ), 
        .ZN(_f_permutation__round__n717 ) );
  INV_X4 _f_permutation__round__U2316  ( .A(_f_permutation__round__c[842] ), 
        .ZN(_f_permutation__round__n716 ) );
  INV_X4 _f_permutation__round__U2315  ( .A(_f_permutation__round__c[778] ), 
        .ZN(_f_permutation__round__n715 ) );
  INV_X4 _f_permutation__round__U2314  ( .A(_f_permutation__round__c[650] ), 
        .ZN(_f_permutation__round__n714 ) );
  INV_X4 _f_permutation__round__U2313  ( .A(_f_permutation__round__c[204] ), 
        .ZN(_f_permutation__round__n713 ) );
  INV_X4 _f_permutation__round__U2312  ( .A(_f_permutation__round__c[140] ), 
        .ZN(_f_permutation__round__n712 ) );
  INV_X4 _f_permutation__round__U2311  ( .A(_f_permutation__round__c[843] ), 
        .ZN(_f_permutation__round__n711 ) );
  INV_X4 _f_permutation__round__U2310  ( .A(_f_permutation__round__c[779] ), 
        .ZN(_f_permutation__round__n710 ) );
  INV_X4 _f_permutation__round__U2309  ( .A(_f_permutation__round__c[651] ), 
        .ZN(_f_permutation__round__n709 ) );
  INV_X4 _f_permutation__round__U2308  ( .A(_f_permutation__round__c[205] ), 
        .ZN(_f_permutation__round__n708 ) );
  INV_X4 _f_permutation__round__U2307  ( .A(_f_permutation__round__c[141] ), 
        .ZN(_f_permutation__round__n707 ) );
  INV_X4 _f_permutation__round__U2306  ( .A(_f_permutation__round__c[844] ), 
        .ZN(_f_permutation__round__n706 ) );
  INV_X4 _f_permutation__round__U2305  ( .A(_f_permutation__round__c[780] ), 
        .ZN(_f_permutation__round__n705 ) );
  INV_X4 _f_permutation__round__U2304  ( .A(_f_permutation__round__c[652] ), 
        .ZN(_f_permutation__round__n704 ) );
  INV_X4 _f_permutation__round__U2303  ( .A(_f_permutation__round__c[206] ), 
        .ZN(_f_permutation__round__n703 ) );
  INV_X4 _f_permutation__round__U2302  ( .A(_f_permutation__round__c[142] ), 
        .ZN(_f_permutation__round__n702 ) );
  INV_X4 _f_permutation__round__U2301  ( .A(_f_permutation__round__c[845] ), 
        .ZN(_f_permutation__round__n701 ) );
  INV_X4 _f_permutation__round__U2300  ( .A(_f_permutation__round__c[781] ), 
        .ZN(_f_permutation__round__n700 ) );
  INV_X4 _f_permutation__round__U2299  ( .A(_f_permutation__round__c[653] ), 
        .ZN(_f_permutation__round__n699 ) );
  INV_X4 _f_permutation__round__U2298  ( .A(_f_permutation__round__c[207] ), 
        .ZN(_f_permutation__round__n698 ) );
  INV_X4 _f_permutation__round__U2297  ( .A(_f_permutation__round__c[143] ), 
        .ZN(_f_permutation__round__n697 ) );
  INV_X4 _f_permutation__round__U2296  ( .A(_f_permutation__round__c[846] ), 
        .ZN(_f_permutation__round__n696 ) );
  INV_X4 _f_permutation__round__U2295  ( .A(_f_permutation__round__c[782] ), 
        .ZN(_f_permutation__round__n695 ) );
  INV_X4 _f_permutation__round__U2294  ( .A(_f_permutation__round__c[654] ), 
        .ZN(_f_permutation__round__n694 ) );
  INV_X4 _f_permutation__round__U2293  ( .A(_f_permutation__round__c[208] ), 
        .ZN(_f_permutation__round__n693 ) );
  INV_X4 _f_permutation__round__U2292  ( .A(_f_permutation__round__c[144] ), 
        .ZN(_f_permutation__round__n692 ) );
  INV_X4 _f_permutation__round__U2291  ( .A(_f_permutation__round__c[847] ), 
        .ZN(_f_permutation__round__n691 ) );
  INV_X4 _f_permutation__round__U2290  ( .A(_f_permutation__round__c[783] ), 
        .ZN(_f_permutation__round__n690 ) );
  INV_X4 _f_permutation__round__U2289  ( .A(_f_permutation__round__c[655] ), 
        .ZN(_f_permutation__round__n689 ) );
  INV_X4 _f_permutation__round__U2288  ( .A(_f_permutation__round__c[209] ), 
        .ZN(_f_permutation__round__n688 ) );
  INV_X4 _f_permutation__round__U2287  ( .A(_f_permutation__round__c[145] ), 
        .ZN(_f_permutation__round__n687 ) );
  INV_X4 _f_permutation__round__U2286  ( .A(_f_permutation__round__c[848] ), 
        .ZN(_f_permutation__round__n686 ) );
  INV_X4 _f_permutation__round__U2285  ( .A(_f_permutation__round__c[784] ), 
        .ZN(_f_permutation__round__n685 ) );
  INV_X4 _f_permutation__round__U2284  ( .A(_f_permutation__round__c[656] ), 
        .ZN(_f_permutation__round__n684 ) );
  INV_X4 _f_permutation__round__U2283  ( .A(_f_permutation__round__c[210] ), 
        .ZN(_f_permutation__round__n683 ) );
  INV_X4 _f_permutation__round__U2282  ( .A(_f_permutation__round__c[146] ), 
        .ZN(_f_permutation__round__n682 ) );
  INV_X4 _f_permutation__round__U2281  ( .A(_f_permutation__round__c[849] ), 
        .ZN(_f_permutation__round__n681 ) );
  INV_X4 _f_permutation__round__U2280  ( .A(_f_permutation__round__c[785] ), 
        .ZN(_f_permutation__round__n680 ) );
  INV_X4 _f_permutation__round__U2279  ( .A(_f_permutation__round__c[657] ), 
        .ZN(_f_permutation__round__n679 ) );
  INV_X4 _f_permutation__round__U2278  ( .A(_f_permutation__round__c[211] ), 
        .ZN(_f_permutation__round__n678 ) );
  INV_X4 _f_permutation__round__U2277  ( .A(_f_permutation__round__c[147] ), 
        .ZN(_f_permutation__round__n677 ) );
  INV_X4 _f_permutation__round__U2276  ( .A(_f_permutation__round__c[850] ), 
        .ZN(_f_permutation__round__n676 ) );
  INV_X4 _f_permutation__round__U2275  ( .A(_f_permutation__round__c[786] ), 
        .ZN(_f_permutation__round__n675 ) );
  INV_X4 _f_permutation__round__U2274  ( .A(_f_permutation__round__c[658] ), 
        .ZN(_f_permutation__round__n674 ) );
  INV_X4 _f_permutation__round__U2273  ( .A(_f_permutation__round__c[212] ), 
        .ZN(_f_permutation__round__n673 ) );
  INV_X4 _f_permutation__round__U2272  ( .A(_f_permutation__round__c[148] ), 
        .ZN(_f_permutation__round__n672 ) );
  INV_X4 _f_permutation__round__U2271  ( .A(_f_permutation__round__c[851] ), 
        .ZN(_f_permutation__round__n671 ) );
  INV_X4 _f_permutation__round__U2270  ( .A(_f_permutation__round__c[787] ), 
        .ZN(_f_permutation__round__n670 ) );
  INV_X4 _f_permutation__round__U2269  ( .A(_f_permutation__round__c[659] ), 
        .ZN(_f_permutation__round__n669 ) );
  INV_X4 _f_permutation__round__U2268  ( .A(_f_permutation__round__c[213] ), 
        .ZN(_f_permutation__round__n668 ) );
  INV_X4 _f_permutation__round__U2267  ( .A(_f_permutation__round__c[149] ), 
        .ZN(_f_permutation__round__n667 ) );
  INV_X4 _f_permutation__round__U2266  ( .A(_f_permutation__round__c[852] ), 
        .ZN(_f_permutation__round__n666 ) );
  INV_X4 _f_permutation__round__U2265  ( .A(_f_permutation__round__c[788] ), 
        .ZN(_f_permutation__round__n665 ) );
  INV_X4 _f_permutation__round__U2264  ( .A(_f_permutation__round__c[660] ), 
        .ZN(_f_permutation__round__n664 ) );
  INV_X4 _f_permutation__round__U2263  ( .A(_f_permutation__round__c[214] ), 
        .ZN(_f_permutation__round__n663 ) );
  INV_X4 _f_permutation__round__U2262  ( .A(_f_permutation__round__c[150] ), 
        .ZN(_f_permutation__round__n662 ) );
  INV_X4 _f_permutation__round__U2261  ( .A(_f_permutation__round__c[853] ), 
        .ZN(_f_permutation__round__n661 ) );
  INV_X4 _f_permutation__round__U2260  ( .A(_f_permutation__round__c[789] ), 
        .ZN(_f_permutation__round__n660 ) );
  INV_X4 _f_permutation__round__U2259  ( .A(_f_permutation__round__c[661] ), 
        .ZN(_f_permutation__round__n659 ) );
  INV_X4 _f_permutation__round__U2258  ( .A(_f_permutation__round__c[215] ), 
        .ZN(_f_permutation__round__n658 ) );
  INV_X4 _f_permutation__round__U2257  ( .A(_f_permutation__round__c[151] ), 
        .ZN(_f_permutation__round__n657 ) );
  INV_X4 _f_permutation__round__U2256  ( .A(_f_permutation__round__c[854] ), 
        .ZN(_f_permutation__round__n656 ) );
  INV_X4 _f_permutation__round__U2255  ( .A(_f_permutation__round__c[790] ), 
        .ZN(_f_permutation__round__n655 ) );
  INV_X4 _f_permutation__round__U2254  ( .A(_f_permutation__round__c[662] ), 
        .ZN(_f_permutation__round__n654 ) );
  INV_X4 _f_permutation__round__U2253  ( .A(_f_permutation__round__c[216] ), 
        .ZN(_f_permutation__round__n653 ) );
  INV_X4 _f_permutation__round__U2252  ( .A(_f_permutation__round__c[152] ), 
        .ZN(_f_permutation__round__n652 ) );
  INV_X4 _f_permutation__round__U2251  ( .A(_f_permutation__round__c[855] ), 
        .ZN(_f_permutation__round__n651 ) );
  INV_X4 _f_permutation__round__U2250  ( .A(_f_permutation__round__c[791] ), 
        .ZN(_f_permutation__round__n650 ) );
  INV_X4 _f_permutation__round__U2249  ( .A(_f_permutation__round__c[663] ), 
        .ZN(_f_permutation__round__n649 ) );
  INV_X4 _f_permutation__round__U2248  ( .A(_f_permutation__round__c[217] ), 
        .ZN(_f_permutation__round__n648 ) );
  INV_X4 _f_permutation__round__U2247  ( .A(_f_permutation__round__c[153] ), 
        .ZN(_f_permutation__round__n647 ) );
  INV_X4 _f_permutation__round__U2246  ( .A(_f_permutation__round__c[856] ), 
        .ZN(_f_permutation__round__n646 ) );
  INV_X4 _f_permutation__round__U2245  ( .A(_f_permutation__round__c[792] ), 
        .ZN(_f_permutation__round__n645 ) );
  INV_X4 _f_permutation__round__U2244  ( .A(_f_permutation__round__c[664] ), 
        .ZN(_f_permutation__round__n644 ) );
  INV_X4 _f_permutation__round__U2243  ( .A(_f_permutation__round__c[218] ), 
        .ZN(_f_permutation__round__n643 ) );
  INV_X4 _f_permutation__round__U2242  ( .A(_f_permutation__round__c[154] ), 
        .ZN(_f_permutation__round__n642 ) );
  INV_X4 _f_permutation__round__U2241  ( .A(_f_permutation__round__c[857] ), 
        .ZN(_f_permutation__round__n641 ) );
  INV_X4 _f_permutation__round__U2240  ( .A(_f_permutation__round__c[793] ), 
        .ZN(_f_permutation__round__n640 ) );
  INV_X4 _f_permutation__round__U2239  ( .A(_f_permutation__round__c[665] ), 
        .ZN(_f_permutation__round__n639 ) );
  INV_X4 _f_permutation__round__U2238  ( .A(_f_permutation__round__c[219] ), 
        .ZN(_f_permutation__round__n638 ) );
  INV_X4 _f_permutation__round__U2237  ( .A(_f_permutation__round__c[155] ), 
        .ZN(_f_permutation__round__n637 ) );
  INV_X4 _f_permutation__round__U2236  ( .A(_f_permutation__round__c[858] ), 
        .ZN(_f_permutation__round__n636 ) );
  INV_X4 _f_permutation__round__U2235  ( .A(_f_permutation__round__c[794] ), 
        .ZN(_f_permutation__round__n635 ) );
  INV_X4 _f_permutation__round__U2234  ( .A(_f_permutation__round__c[666] ), 
        .ZN(_f_permutation__round__n634 ) );
  INV_X4 _f_permutation__round__U2233  ( .A(_f_permutation__round__c[220] ), 
        .ZN(_f_permutation__round__n633 ) );
  INV_X4 _f_permutation__round__U2232  ( .A(_f_permutation__round__c[156] ), 
        .ZN(_f_permutation__round__n632 ) );
  INV_X4 _f_permutation__round__U2231  ( .A(_f_permutation__round__c[859] ), 
        .ZN(_f_permutation__round__n631 ) );
  INV_X4 _f_permutation__round__U2230  ( .A(_f_permutation__round__c[795] ), 
        .ZN(_f_permutation__round__n630 ) );
  INV_X4 _f_permutation__round__U2229  ( .A(_f_permutation__round__c[667] ), 
        .ZN(_f_permutation__round__n629 ) );
  INV_X4 _f_permutation__round__U2228  ( .A(_f_permutation__round__c[221] ), 
        .ZN(_f_permutation__round__n628 ) );
  INV_X4 _f_permutation__round__U2227  ( .A(_f_permutation__round__c[157] ), 
        .ZN(_f_permutation__round__n627 ) );
  INV_X4 _f_permutation__round__U2226  ( .A(_f_permutation__round__c[860] ), 
        .ZN(_f_permutation__round__n626 ) );
  INV_X4 _f_permutation__round__U2225  ( .A(_f_permutation__round__c[796] ), 
        .ZN(_f_permutation__round__n625 ) );
  INV_X4 _f_permutation__round__U2224  ( .A(_f_permutation__round__c[668] ), 
        .ZN(_f_permutation__round__n624 ) );
  INV_X4 _f_permutation__round__U2223  ( .A(_f_permutation__round__c[222] ), 
        .ZN(_f_permutation__round__n623 ) );
  INV_X4 _f_permutation__round__U2222  ( .A(_f_permutation__round__c[158] ), 
        .ZN(_f_permutation__round__n622 ) );
  INV_X4 _f_permutation__round__U2221  ( .A(_f_permutation__round__c[861] ), 
        .ZN(_f_permutation__round__n621 ) );
  INV_X4 _f_permutation__round__U2220  ( .A(_f_permutation__round__c[797] ), 
        .ZN(_f_permutation__round__n620 ) );
  INV_X4 _f_permutation__round__U2219  ( .A(_f_permutation__round__c[669] ), 
        .ZN(_f_permutation__round__n619 ) );
  INV_X4 _f_permutation__round__U2218  ( .A(_f_permutation__round__c[223] ), 
        .ZN(_f_permutation__round__n618 ) );
  INV_X4 _f_permutation__round__U2217  ( .A(_f_permutation__round__c[159] ), 
        .ZN(_f_permutation__round__n617 ) );
  INV_X4 _f_permutation__round__U2216  ( .A(_f_permutation__round__c[862] ), 
        .ZN(_f_permutation__round__n616 ) );
  INV_X4 _f_permutation__round__U2215  ( .A(_f_permutation__round__c[798] ), 
        .ZN(_f_permutation__round__n615 ) );
  INV_X4 _f_permutation__round__U2214  ( .A(_f_permutation__round__c[670] ), 
        .ZN(_f_permutation__round__n614 ) );
  INV_X4 _f_permutation__round__U2213  ( .A(_f_permutation__round__c[224] ), 
        .ZN(_f_permutation__round__n613 ) );
  INV_X4 _f_permutation__round__U2212  ( .A(_f_permutation__round__c[160] ), 
        .ZN(_f_permutation__round__n612 ) );
  INV_X4 _f_permutation__round__U2211  ( .A(_f_permutation__round__c[863] ), 
        .ZN(_f_permutation__round__n611 ) );
  INV_X4 _f_permutation__round__U2210  ( .A(_f_permutation__round__c[799] ), 
        .ZN(_f_permutation__round__n610 ) );
  INV_X4 _f_permutation__round__U2209  ( .A(_f_permutation__round__c[671] ), 
        .ZN(_f_permutation__round__n609 ) );
  INV_X4 _f_permutation__round__U2208  ( .A(_f_permutation__round__c[225] ), 
        .ZN(_f_permutation__round__n608 ) );
  INV_X4 _f_permutation__round__U2207  ( .A(_f_permutation__round__c[161] ), 
        .ZN(_f_permutation__round__n607 ) );
  INV_X4 _f_permutation__round__U2206  ( .A(_f_permutation__round__c[864] ), 
        .ZN(_f_permutation__round__n606 ) );
  INV_X4 _f_permutation__round__U2205  ( .A(_f_permutation__round__c[800] ), 
        .ZN(_f_permutation__round__n605 ) );
  INV_X4 _f_permutation__round__U2204  ( .A(_f_permutation__round__c[672] ), 
        .ZN(_f_permutation__round__n604 ) );
  INV_X4 _f_permutation__round__U2203  ( .A(_f_permutation__round__c[226] ), 
        .ZN(_f_permutation__round__n603 ) );
  INV_X4 _f_permutation__round__U2202  ( .A(_f_permutation__round__c[162] ), 
        .ZN(_f_permutation__round__n602 ) );
  INV_X4 _f_permutation__round__U2201  ( .A(_f_permutation__round__c[865] ), 
        .ZN(_f_permutation__round__n601 ) );
  INV_X4 _f_permutation__round__U2200  ( .A(_f_permutation__round__c[801] ), 
        .ZN(_f_permutation__round__n600 ) );
  INV_X4 _f_permutation__round__U2199  ( .A(_f_permutation__round__c[673] ), 
        .ZN(_f_permutation__round__n599 ) );
  INV_X4 _f_permutation__round__U2198  ( .A(_f_permutation__round__c[227] ), 
        .ZN(_f_permutation__round__n598 ) );
  INV_X4 _f_permutation__round__U2197  ( .A(_f_permutation__round__c[163] ), 
        .ZN(_f_permutation__round__n597 ) );
  INV_X4 _f_permutation__round__U2196  ( .A(_f_permutation__round__c[866] ), 
        .ZN(_f_permutation__round__n596 ) );
  INV_X4 _f_permutation__round__U2195  ( .A(_f_permutation__round__c[802] ), 
        .ZN(_f_permutation__round__n595 ) );
  INV_X4 _f_permutation__round__U2194  ( .A(_f_permutation__round__c[674] ), 
        .ZN(_f_permutation__round__n594 ) );
  INV_X4 _f_permutation__round__U2193  ( .A(_f_permutation__round__c[228] ), 
        .ZN(_f_permutation__round__n593 ) );
  INV_X4 _f_permutation__round__U2192  ( .A(_f_permutation__round__c[164] ), 
        .ZN(_f_permutation__round__n592 ) );
  INV_X4 _f_permutation__round__U2191  ( .A(_f_permutation__round__c[867] ), 
        .ZN(_f_permutation__round__n591 ) );
  INV_X4 _f_permutation__round__U2190  ( .A(_f_permutation__round__c[803] ), 
        .ZN(_f_permutation__round__n590 ) );
  INV_X4 _f_permutation__round__U2189  ( .A(_f_permutation__round__c[675] ), 
        .ZN(_f_permutation__round__n589 ) );
  INV_X4 _f_permutation__round__U2188  ( .A(_f_permutation__round__c[229] ), 
        .ZN(_f_permutation__round__n588 ) );
  INV_X4 _f_permutation__round__U2187  ( .A(_f_permutation__round__c[165] ), 
        .ZN(_f_permutation__round__n587 ) );
  INV_X4 _f_permutation__round__U2186  ( .A(_f_permutation__round__c[868] ), 
        .ZN(_f_permutation__round__n586 ) );
  INV_X4 _f_permutation__round__U2185  ( .A(_f_permutation__round__c[804] ), 
        .ZN(_f_permutation__round__n585 ) );
  INV_X4 _f_permutation__round__U2184  ( .A(_f_permutation__round__c[676] ), 
        .ZN(_f_permutation__round__n584 ) );
  INV_X4 _f_permutation__round__U2183  ( .A(_f_permutation__round__c[230] ), 
        .ZN(_f_permutation__round__n583 ) );
  INV_X4 _f_permutation__round__U2182  ( .A(_f_permutation__round__c[166] ), 
        .ZN(_f_permutation__round__n582 ) );
  INV_X4 _f_permutation__round__U2181  ( .A(_f_permutation__round__c[869] ), 
        .ZN(_f_permutation__round__n581 ) );
  INV_X4 _f_permutation__round__U2180  ( .A(_f_permutation__round__c[805] ), 
        .ZN(_f_permutation__round__n580 ) );
  INV_X4 _f_permutation__round__U2179  ( .A(_f_permutation__round__c[677] ), 
        .ZN(_f_permutation__round__n579 ) );
  INV_X4 _f_permutation__round__U2178  ( .A(_f_permutation__round__c[231] ), 
        .ZN(_f_permutation__round__n578 ) );
  INV_X4 _f_permutation__round__U2177  ( .A(_f_permutation__round__c[167] ), 
        .ZN(_f_permutation__round__n577 ) );
  INV_X4 _f_permutation__round__U2176  ( .A(_f_permutation__round__c[870] ), 
        .ZN(_f_permutation__round__n576 ) );
  INV_X4 _f_permutation__round__U2175  ( .A(_f_permutation__round__c[806] ), 
        .ZN(_f_permutation__round__n575 ) );
  INV_X4 _f_permutation__round__U2174  ( .A(_f_permutation__round__c[678] ), 
        .ZN(_f_permutation__round__n574 ) );
  INV_X4 _f_permutation__round__U2173  ( .A(_f_permutation__round__c[232] ), 
        .ZN(_f_permutation__round__n573 ) );
  INV_X4 _f_permutation__round__U2172  ( .A(_f_permutation__round__c[168] ), 
        .ZN(_f_permutation__round__n572 ) );
  INV_X4 _f_permutation__round__U2171  ( .A(_f_permutation__round__c[871] ), 
        .ZN(_f_permutation__round__n571 ) );
  INV_X4 _f_permutation__round__U2170  ( .A(_f_permutation__round__c[807] ), 
        .ZN(_f_permutation__round__n570 ) );
  INV_X4 _f_permutation__round__U2169  ( .A(_f_permutation__round__c[679] ), 
        .ZN(_f_permutation__round__n569 ) );
  INV_X4 _f_permutation__round__U2168  ( .A(_f_permutation__round__c[233] ), 
        .ZN(_f_permutation__round__n568 ) );
  INV_X4 _f_permutation__round__U2167  ( .A(_f_permutation__round__c[169] ), 
        .ZN(_f_permutation__round__n567 ) );
  INV_X4 _f_permutation__round__U2166  ( .A(_f_permutation__round__c[872] ), 
        .ZN(_f_permutation__round__n566 ) );
  INV_X4 _f_permutation__round__U2165  ( .A(_f_permutation__round__c[808] ), 
        .ZN(_f_permutation__round__n565 ) );
  INV_X4 _f_permutation__round__U2164  ( .A(_f_permutation__round__c[680] ), 
        .ZN(_f_permutation__round__n564 ) );
  INV_X4 _f_permutation__round__U2163  ( .A(_f_permutation__round__c[234] ), 
        .ZN(_f_permutation__round__n563 ) );
  INV_X4 _f_permutation__round__U2162  ( .A(_f_permutation__round__c[170] ), 
        .ZN(_f_permutation__round__n562 ) );
  INV_X4 _f_permutation__round__U2161  ( .A(_f_permutation__round__c[873] ), 
        .ZN(_f_permutation__round__n561 ) );
  INV_X4 _f_permutation__round__U2160  ( .A(_f_permutation__round__c[809] ), 
        .ZN(_f_permutation__round__n560 ) );
  INV_X4 _f_permutation__round__U2159  ( .A(_f_permutation__round__c[681] ), 
        .ZN(_f_permutation__round__n559 ) );
  INV_X4 _f_permutation__round__U2158  ( .A(_f_permutation__round__c[235] ), 
        .ZN(_f_permutation__round__n558 ) );
  INV_X4 _f_permutation__round__U2157  ( .A(_f_permutation__round__c[171] ), 
        .ZN(_f_permutation__round__n557 ) );
  INV_X4 _f_permutation__round__U2156  ( .A(_f_permutation__round__c[874] ), 
        .ZN(_f_permutation__round__n556 ) );
  INV_X4 _f_permutation__round__U2155  ( .A(_f_permutation__round__c[810] ), 
        .ZN(_f_permutation__round__n555 ) );
  INV_X4 _f_permutation__round__U2154  ( .A(_f_permutation__round__c[682] ), 
        .ZN(_f_permutation__round__n554 ) );
  INV_X4 _f_permutation__round__U2153  ( .A(_f_permutation__round__c[236] ), 
        .ZN(_f_permutation__round__n553 ) );
  INV_X4 _f_permutation__round__U2152  ( .A(_f_permutation__round__c[172] ), 
        .ZN(_f_permutation__round__n552 ) );
  INV_X4 _f_permutation__round__U2151  ( .A(_f_permutation__round__c[875] ), 
        .ZN(_f_permutation__round__n551 ) );
  INV_X4 _f_permutation__round__U2150  ( .A(_f_permutation__round__c[811] ), 
        .ZN(_f_permutation__round__n550 ) );
  INV_X4 _f_permutation__round__U2149  ( .A(_f_permutation__round__c[683] ), 
        .ZN(_f_permutation__round__n549 ) );
  INV_X4 _f_permutation__round__U2148  ( .A(_f_permutation__round__c[237] ), 
        .ZN(_f_permutation__round__n548 ) );
  INV_X4 _f_permutation__round__U2147  ( .A(_f_permutation__round__c[173] ), 
        .ZN(_f_permutation__round__n547 ) );
  INV_X4 _f_permutation__round__U2146  ( .A(_f_permutation__round__c[876] ), 
        .ZN(_f_permutation__round__n546 ) );
  INV_X4 _f_permutation__round__U2145  ( .A(_f_permutation__round__c[812] ), 
        .ZN(_f_permutation__round__n545 ) );
  INV_X4 _f_permutation__round__U2144  ( .A(_f_permutation__round__c[684] ), 
        .ZN(_f_permutation__round__n544 ) );
  INV_X4 _f_permutation__round__U2143  ( .A(_f_permutation__round__c[238] ), 
        .ZN(_f_permutation__round__n543 ) );
  INV_X4 _f_permutation__round__U2142  ( .A(_f_permutation__round__c[174] ), 
        .ZN(_f_permutation__round__n542 ) );
  INV_X4 _f_permutation__round__U2141  ( .A(_f_permutation__round__c[877] ), 
        .ZN(_f_permutation__round__n541 ) );
  INV_X4 _f_permutation__round__U2140  ( .A(_f_permutation__round__c[813] ), 
        .ZN(_f_permutation__round__n540 ) );
  INV_X4 _f_permutation__round__U2139  ( .A(_f_permutation__round__c[685] ), 
        .ZN(_f_permutation__round__n539 ) );
  INV_X4 _f_permutation__round__U2138  ( .A(_f_permutation__round__c[239] ), 
        .ZN(_f_permutation__round__n538 ) );
  INV_X4 _f_permutation__round__U2137  ( .A(_f_permutation__round__c[175] ), 
        .ZN(_f_permutation__round__n537 ) );
  INV_X4 _f_permutation__round__U2136  ( .A(_f_permutation__round__c[878] ), 
        .ZN(_f_permutation__round__n536 ) );
  INV_X4 _f_permutation__round__U2135  ( .A(_f_permutation__round__c[814] ), 
        .ZN(_f_permutation__round__n535 ) );
  INV_X4 _f_permutation__round__U2134  ( .A(_f_permutation__round__c[686] ), 
        .ZN(_f_permutation__round__n534 ) );
  INV_X4 _f_permutation__round__U2133  ( .A(_f_permutation__round__c[240] ), 
        .ZN(_f_permutation__round__n533 ) );
  INV_X4 _f_permutation__round__U2132  ( .A(_f_permutation__round__c[176] ), 
        .ZN(_f_permutation__round__n532 ) );
  INV_X4 _f_permutation__round__U2131  ( .A(_f_permutation__round__c[879] ), 
        .ZN(_f_permutation__round__n531 ) );
  INV_X4 _f_permutation__round__U2130  ( .A(_f_permutation__round__c[815] ), 
        .ZN(_f_permutation__round__n530 ) );
  INV_X4 _f_permutation__round__U2129  ( .A(_f_permutation__round__c[687] ), 
        .ZN(_f_permutation__round__n529 ) );
  INV_X4 _f_permutation__round__U2128  ( .A(_f_permutation__round__c[241] ), 
        .ZN(_f_permutation__round__n528 ) );
  INV_X4 _f_permutation__round__U2127  ( .A(_f_permutation__round__c[177] ), 
        .ZN(_f_permutation__round__n527 ) );
  INV_X4 _f_permutation__round__U2126  ( .A(_f_permutation__round__c[880] ), 
        .ZN(_f_permutation__round__n526 ) );
  INV_X4 _f_permutation__round__U2125  ( .A(_f_permutation__round__c[816] ), 
        .ZN(_f_permutation__round__n525 ) );
  INV_X4 _f_permutation__round__U2124  ( .A(_f_permutation__round__c[688] ), 
        .ZN(_f_permutation__round__n524 ) );
  INV_X4 _f_permutation__round__U2123  ( .A(_f_permutation__round__c[242] ), 
        .ZN(_f_permutation__round__n523 ) );
  INV_X4 _f_permutation__round__U2122  ( .A(_f_permutation__round__c[178] ), 
        .ZN(_f_permutation__round__n522 ) );
  INV_X4 _f_permutation__round__U2121  ( .A(_f_permutation__round__c[881] ), 
        .ZN(_f_permutation__round__n521 ) );
  INV_X4 _f_permutation__round__U2120  ( .A(_f_permutation__round__c[817] ), 
        .ZN(_f_permutation__round__n520 ) );
  INV_X4 _f_permutation__round__U2119  ( .A(_f_permutation__round__c[689] ), 
        .ZN(_f_permutation__round__n519 ) );
  INV_X4 _f_permutation__round__U2118  ( .A(_f_permutation__round__c[243] ), 
        .ZN(_f_permutation__round__n518 ) );
  INV_X4 _f_permutation__round__U2117  ( .A(_f_permutation__round__c[179] ), 
        .ZN(_f_permutation__round__n517 ) );
  INV_X4 _f_permutation__round__U2116  ( .A(_f_permutation__round__c[882] ), 
        .ZN(_f_permutation__round__n516 ) );
  INV_X4 _f_permutation__round__U2115  ( .A(_f_permutation__round__c[818] ), 
        .ZN(_f_permutation__round__n515 ) );
  INV_X4 _f_permutation__round__U2114  ( .A(_f_permutation__round__c[690] ), 
        .ZN(_f_permutation__round__n514 ) );
  INV_X4 _f_permutation__round__U2113  ( .A(_f_permutation__round__c[244] ), 
        .ZN(_f_permutation__round__n513 ) );
  INV_X4 _f_permutation__round__U2112  ( .A(_f_permutation__round__c[180] ), 
        .ZN(_f_permutation__round__n512 ) );
  INV_X4 _f_permutation__round__U2111  ( .A(_f_permutation__round__c[883] ), 
        .ZN(_f_permutation__round__n511 ) );
  INV_X4 _f_permutation__round__U2110  ( .A(_f_permutation__round__c[819] ), 
        .ZN(_f_permutation__round__n510 ) );
  INV_X4 _f_permutation__round__U2109  ( .A(_f_permutation__round__c[691] ), 
        .ZN(_f_permutation__round__n509 ) );
  INV_X4 _f_permutation__round__U2108  ( .A(_f_permutation__round__c[245] ), 
        .ZN(_f_permutation__round__n508 ) );
  INV_X4 _f_permutation__round__U2107  ( .A(_f_permutation__round__c[181] ), 
        .ZN(_f_permutation__round__n507 ) );
  INV_X4 _f_permutation__round__U2106  ( .A(_f_permutation__round__c[884] ), 
        .ZN(_f_permutation__round__n506 ) );
  INV_X4 _f_permutation__round__U2105  ( .A(_f_permutation__round__c[820] ), 
        .ZN(_f_permutation__round__n505 ) );
  INV_X4 _f_permutation__round__U2104  ( .A(_f_permutation__round__c[692] ), 
        .ZN(_f_permutation__round__n504 ) );
  INV_X4 _f_permutation__round__U2103  ( .A(_f_permutation__round__c[246] ), 
        .ZN(_f_permutation__round__n503 ) );
  INV_X4 _f_permutation__round__U2102  ( .A(_f_permutation__round__c[182] ), 
        .ZN(_f_permutation__round__n502 ) );
  INV_X4 _f_permutation__round__U2101  ( .A(_f_permutation__round__c[885] ), 
        .ZN(_f_permutation__round__n501 ) );
  INV_X4 _f_permutation__round__U2100  ( .A(_f_permutation__round__c[821] ), 
        .ZN(_f_permutation__round__n500 ) );
  INV_X4 _f_permutation__round__U2099  ( .A(_f_permutation__round__c[693] ), 
        .ZN(_f_permutation__round__n499 ) );
  INV_X4 _f_permutation__round__U2098  ( .A(_f_permutation__round__c[247] ), 
        .ZN(_f_permutation__round__n498 ) );
  INV_X4 _f_permutation__round__U2097  ( .A(_f_permutation__round__c[183] ), 
        .ZN(_f_permutation__round__n497 ) );
  INV_X4 _f_permutation__round__U2096  ( .A(_f_permutation__round__c[886] ), 
        .ZN(_f_permutation__round__n496 ) );
  INV_X4 _f_permutation__round__U2095  ( .A(_f_permutation__round__c[822] ), 
        .ZN(_f_permutation__round__n495 ) );
  INV_X4 _f_permutation__round__U2094  ( .A(_f_permutation__round__c[694] ), 
        .ZN(_f_permutation__round__n494 ) );
  INV_X4 _f_permutation__round__U2093  ( .A(_f_permutation__round__c[248] ), 
        .ZN(_f_permutation__round__n493 ) );
  INV_X4 _f_permutation__round__U2092  ( .A(_f_permutation__round__c[184] ), 
        .ZN(_f_permutation__round__n492 ) );
  INV_X4 _f_permutation__round__U2091  ( .A(_f_permutation__round__c[887] ), 
        .ZN(_f_permutation__round__n491 ) );
  INV_X4 _f_permutation__round__U2090  ( .A(_f_permutation__round__c[823] ), 
        .ZN(_f_permutation__round__n490 ) );
  INV_X4 _f_permutation__round__U2089  ( .A(_f_permutation__round__c[695] ), 
        .ZN(_f_permutation__round__n489 ) );
  INV_X4 _f_permutation__round__U2088  ( .A(_f_permutation__round__c[249] ), 
        .ZN(_f_permutation__round__n488 ) );
  INV_X4 _f_permutation__round__U2087  ( .A(_f_permutation__round__c[185] ), 
        .ZN(_f_permutation__round__n487 ) );
  INV_X4 _f_permutation__round__U2086  ( .A(_f_permutation__round__c[888] ), 
        .ZN(_f_permutation__round__n486 ) );
  INV_X4 _f_permutation__round__U2085  ( .A(_f_permutation__round__c[824] ), 
        .ZN(_f_permutation__round__n485 ) );
  INV_X4 _f_permutation__round__U2084  ( .A(_f_permutation__round__c[696] ), 
        .ZN(_f_permutation__round__n484 ) );
  INV_X4 _f_permutation__round__U2083  ( .A(_f_permutation__round__c[250] ), 
        .ZN(_f_permutation__round__n483 ) );
  INV_X4 _f_permutation__round__U2082  ( .A(_f_permutation__round__c[186] ), 
        .ZN(_f_permutation__round__n482 ) );
  INV_X4 _f_permutation__round__U2081  ( .A(_f_permutation__round__c[889] ), 
        .ZN(_f_permutation__round__n481 ) );
  INV_X4 _f_permutation__round__U2080  ( .A(_f_permutation__round__c[825] ), 
        .ZN(_f_permutation__round__n480 ) );
  INV_X4 _f_permutation__round__U2079  ( .A(_f_permutation__round__c[697] ), 
        .ZN(_f_permutation__round__n479 ) );
  INV_X4 _f_permutation__round__U2078  ( .A(_f_permutation__round__c[251] ), 
        .ZN(_f_permutation__round__n478 ) );
  INV_X4 _f_permutation__round__U2077  ( .A(_f_permutation__round__c[187] ), 
        .ZN(_f_permutation__round__n477 ) );
  INV_X4 _f_permutation__round__U2076  ( .A(_f_permutation__round__c[890] ), 
        .ZN(_f_permutation__round__n476 ) );
  INV_X4 _f_permutation__round__U2075  ( .A(_f_permutation__round__c[826] ), 
        .ZN(_f_permutation__round__n475 ) );
  INV_X4 _f_permutation__round__U2074  ( .A(_f_permutation__round__c[698] ), 
        .ZN(_f_permutation__round__n474 ) );
  INV_X4 _f_permutation__round__U2073  ( .A(_f_permutation__round__c[252] ), 
        .ZN(_f_permutation__round__n473 ) );
  INV_X4 _f_permutation__round__U2072  ( .A(_f_permutation__round__c[188] ), 
        .ZN(_f_permutation__round__n472 ) );
  INV_X4 _f_permutation__round__U2071  ( .A(_f_permutation__round__c[891] ), 
        .ZN(_f_permutation__round__n471 ) );
  INV_X4 _f_permutation__round__U2070  ( .A(_f_permutation__round__c[827] ), 
        .ZN(_f_permutation__round__n470 ) );
  INV_X4 _f_permutation__round__U2069  ( .A(_f_permutation__round__c[699] ), 
        .ZN(_f_permutation__round__n469 ) );
  INV_X4 _f_permutation__round__U2068  ( .A(_f_permutation__round__c[253] ), 
        .ZN(_f_permutation__round__n468 ) );
  INV_X4 _f_permutation__round__U2067  ( .A(_f_permutation__round__c[189] ), 
        .ZN(_f_permutation__round__n467 ) );
  INV_X4 _f_permutation__round__U2066  ( .A(_f_permutation__round__c[892] ), 
        .ZN(_f_permutation__round__n466 ) );
  INV_X4 _f_permutation__round__U2065  ( .A(_f_permutation__round__c[828] ), 
        .ZN(_f_permutation__round__n465 ) );
  INV_X4 _f_permutation__round__U2064  ( .A(_f_permutation__round__c[700] ), 
        .ZN(_f_permutation__round__n464 ) );
  INV_X4 _f_permutation__round__U2063  ( .A(_f_permutation__round__c[254] ), 
        .ZN(_f_permutation__round__n463 ) );
  INV_X4 _f_permutation__round__U2062  ( .A(_f_permutation__round__c[190] ), 
        .ZN(_f_permutation__round__n462 ) );
  INV_X4 _f_permutation__round__U2061  ( .A(_f_permutation__round__c[893] ), 
        .ZN(_f_permutation__round__n461 ) );
  INV_X4 _f_permutation__round__U2060  ( .A(_f_permutation__round__c[829] ), 
        .ZN(_f_permutation__round__n460 ) );
  INV_X4 _f_permutation__round__U2059  ( .A(_f_permutation__round__c[701] ), 
        .ZN(_f_permutation__round__n459 ) );
  INV_X4 _f_permutation__round__U2058  ( .A(_f_permutation__round__c[255] ), 
        .ZN(_f_permutation__round__n458 ) );
  INV_X4 _f_permutation__round__U2057  ( .A(_f_permutation__round__c[191] ), 
        .ZN(_f_permutation__round__n457 ) );
  INV_X4 _f_permutation__round__U2056  ( .A(_f_permutation__round__c[894] ), 
        .ZN(_f_permutation__round__n456 ) );
  INV_X4 _f_permutation__round__U2055  ( .A(_f_permutation__round__c[830] ), 
        .ZN(_f_permutation__round__n455 ) );
  INV_X4 _f_permutation__round__U2054  ( .A(_f_permutation__round__c[702] ), 
        .ZN(_f_permutation__round__n454 ) );
  INV_X4 _f_permutation__round__U2053  ( .A(_f_permutation__round__c[192] ), 
        .ZN(_f_permutation__round__n453 ) );
  INV_X4 _f_permutation__round__U2052  ( .A(_f_permutation__round__c[128] ), 
        .ZN(_f_permutation__round__n452 ) );
  INV_X4 _f_permutation__round__U2051  ( .A(_f_permutation__round__c[895] ), 
        .ZN(_f_permutation__round__n451 ) );
  INV_X4 _f_permutation__round__U2050  ( .A(_f_permutation__round__c[831] ), 
        .ZN(_f_permutation__round__n450 ) );
  INV_X4 _f_permutation__round__U2049  ( .A(_f_permutation__round__c[703] ), 
        .ZN(_f_permutation__round__n449 ) );
  INV_X4 _f_permutation__round__U2048  ( .A(_f_permutation__round__c[0] ), 
        .ZN(_f_permutation__round__n448 ) );
  INV_X4 _f_permutation__round__U2047  ( .A(_f_permutation__round__c[1473] ), 
        .ZN(_f_permutation__round__n447 ) );
  INV_X4 _f_permutation__round__U2046  ( .A(_f_permutation__round__c[1409] ), 
        .ZN(_f_permutation__round__n446 ) );
  INV_X4 _f_permutation__round__U2045  ( .A(_f_permutation__round__c[1281] ), 
        .ZN(_f_permutation__round__n445 ) );
  INV_X4 _f_permutation__round__U2044  ( .A(_f_permutation__round__c[512] ), 
        .ZN(_f_permutation__round__n444 ) );
  INV_X4 _f_permutation__round__U2043  ( .A(_f_permutation__round__c[448] ), 
        .ZN(_f_permutation__round__n443 ) );
  INV_X4 _f_permutation__round__U2042  ( .A(_f_permutation__round__c[320] ), 
        .ZN(_f_permutation__round__n442 ) );
  INV_X4 _f_permutation__round__U2041  ( .A(_f_permutation__round__c[1] ), 
        .ZN(_f_permutation__round__n441 ) );
  INV_X4 _f_permutation__round__U2040  ( .A(_f_permutation__round__c[1474] ), 
        .ZN(_f_permutation__round__n440 ) );
  INV_X4 _f_permutation__round__U2039  ( .A(_f_permutation__round__c[1410] ), 
        .ZN(_f_permutation__round__n439 ) );
  INV_X4 _f_permutation__round__U2038  ( .A(_f_permutation__round__c[1282] ), 
        .ZN(_f_permutation__round__n438 ) );
  INV_X4 _f_permutation__round__U2037  ( .A(_f_permutation__round__c[513] ), 
        .ZN(_f_permutation__round__n437 ) );
  INV_X4 _f_permutation__round__U2036  ( .A(_f_permutation__round__c[449] ), 
        .ZN(_f_permutation__round__n436 ) );
  INV_X4 _f_permutation__round__U2035  ( .A(_f_permutation__round__c[321] ), 
        .ZN(_f_permutation__round__n435 ) );
  INV_X4 _f_permutation__round__U2034  ( .A(_f_permutation__round__c[2] ), 
        .ZN(_f_permutation__round__n434 ) );
  INV_X4 _f_permutation__round__U2033  ( .A(_f_permutation__round__c[1475] ), 
        .ZN(_f_permutation__round__n433 ) );
  INV_X4 _f_permutation__round__U2032  ( .A(_f_permutation__round__c[1411] ), 
        .ZN(_f_permutation__round__n432 ) );
  INV_X4 _f_permutation__round__U2031  ( .A(_f_permutation__round__c[1283] ), 
        .ZN(_f_permutation__round__n431 ) );
  INV_X4 _f_permutation__round__U2030  ( .A(_f_permutation__round__c[514] ), 
        .ZN(_f_permutation__round__n430 ) );
  INV_X4 _f_permutation__round__U2029  ( .A(_f_permutation__round__c[450] ), 
        .ZN(_f_permutation__round__n429 ) );
  INV_X4 _f_permutation__round__U2028  ( .A(_f_permutation__round__c[322] ), 
        .ZN(_f_permutation__round__n428 ) );
  INV_X4 _f_permutation__round__U2027  ( .A(_f_permutation__round__c[3] ), 
        .ZN(_f_permutation__round__n427 ) );
  INV_X4 _f_permutation__round__U2026  ( .A(_f_permutation__round__c[1476] ), 
        .ZN(_f_permutation__round__n426 ) );
  INV_X4 _f_permutation__round__U2025  ( .A(_f_permutation__round__c[1412] ), 
        .ZN(_f_permutation__round__n425 ) );
  INV_X4 _f_permutation__round__U2024  ( .A(_f_permutation__round__c[1284] ), 
        .ZN(_f_permutation__round__n424 ) );
  INV_X4 _f_permutation__round__U2023  ( .A(_f_permutation__round__c[515] ), 
        .ZN(_f_permutation__round__n423 ) );
  INV_X4 _f_permutation__round__U2022  ( .A(_f_permutation__round__c[451] ), 
        .ZN(_f_permutation__round__n422 ) );
  INV_X4 _f_permutation__round__U2021  ( .A(_f_permutation__round__c[323] ), 
        .ZN(_f_permutation__round__n421 ) );
  INV_X4 _f_permutation__round__U2020  ( .A(_f_permutation__round__c[4] ), 
        .ZN(_f_permutation__round__n420 ) );
  INV_X4 _f_permutation__round__U2019  ( .A(_f_permutation__round__c[1477] ), 
        .ZN(_f_permutation__round__n419 ) );
  INV_X4 _f_permutation__round__U2018  ( .A(_f_permutation__round__c[1413] ), 
        .ZN(_f_permutation__round__n418 ) );
  INV_X4 _f_permutation__round__U2017  ( .A(_f_permutation__round__c[1285] ), 
        .ZN(_f_permutation__round__n417 ) );
  INV_X4 _f_permutation__round__U2016  ( .A(_f_permutation__round__c[516] ), 
        .ZN(_f_permutation__round__n416 ) );
  INV_X4 _f_permutation__round__U2015  ( .A(_f_permutation__round__c[452] ), 
        .ZN(_f_permutation__round__n415 ) );
  INV_X4 _f_permutation__round__U2014  ( .A(_f_permutation__round__c[324] ), 
        .ZN(_f_permutation__round__n414 ) );
  INV_X4 _f_permutation__round__U2013  ( .A(_f_permutation__round__c[5] ), 
        .ZN(_f_permutation__round__n413 ) );
  INV_X4 _f_permutation__round__U2012  ( .A(_f_permutation__round__c[1478] ), 
        .ZN(_f_permutation__round__n412 ) );
  INV_X4 _f_permutation__round__U2011  ( .A(_f_permutation__round__c[1414] ), 
        .ZN(_f_permutation__round__n411 ) );
  INV_X4 _f_permutation__round__U2010  ( .A(_f_permutation__round__c[1286] ), 
        .ZN(_f_permutation__round__n410 ) );
  INV_X4 _f_permutation__round__U2009  ( .A(_f_permutation__round__c[517] ), 
        .ZN(_f_permutation__round__n409 ) );
  INV_X4 _f_permutation__round__U2008  ( .A(_f_permutation__round__c[453] ), 
        .ZN(_f_permutation__round__n408 ) );
  INV_X4 _f_permutation__round__U2007  ( .A(_f_permutation__round__c[325] ), 
        .ZN(_f_permutation__round__n407 ) );
  INV_X4 _f_permutation__round__U2006  ( .A(_f_permutation__round__c[6] ), 
        .ZN(_f_permutation__round__n406 ) );
  INV_X4 _f_permutation__round__U2005  ( .A(_f_permutation__round__c[1479] ), 
        .ZN(_f_permutation__round__n405 ) );
  INV_X4 _f_permutation__round__U2004  ( .A(_f_permutation__round__c[1415] ), 
        .ZN(_f_permutation__round__n404 ) );
  INV_X4 _f_permutation__round__U2003  ( .A(_f_permutation__round__c[1287] ), 
        .ZN(_f_permutation__round__n403 ) );
  INV_X4 _f_permutation__round__U2002  ( .A(_f_permutation__round__c[518] ), 
        .ZN(_f_permutation__round__n402 ) );
  INV_X4 _f_permutation__round__U2001  ( .A(_f_permutation__round__c[454] ), 
        .ZN(_f_permutation__round__n401 ) );
  INV_X4 _f_permutation__round__U2000  ( .A(_f_permutation__round__c[326] ), 
        .ZN(_f_permutation__round__n400 ) );
  INV_X4 _f_permutation__round__U1999  ( .A(_f_permutation__round__c[7] ), 
        .ZN(_f_permutation__round__n399 ) );
  INV_X4 _f_permutation__round__U1998  ( .A(_f_permutation__round__c[1480] ), 
        .ZN(_f_permutation__round__n398 ) );
  INV_X4 _f_permutation__round__U1997  ( .A(_f_permutation__round__c[1416] ), 
        .ZN(_f_permutation__round__n397 ) );
  INV_X4 _f_permutation__round__U1996  ( .A(_f_permutation__round__c[1288] ), 
        .ZN(_f_permutation__round__n396 ) );
  INV_X4 _f_permutation__round__U1995  ( .A(_f_permutation__round__c[519] ), 
        .ZN(_f_permutation__round__n395 ) );
  INV_X4 _f_permutation__round__U1994  ( .A(_f_permutation__round__c[455] ), 
        .ZN(_f_permutation__round__n394 ) );
  INV_X4 _f_permutation__round__U1993  ( .A(_f_permutation__round__c[327] ), 
        .ZN(_f_permutation__round__n393 ) );
  INV_X4 _f_permutation__round__U1992  ( .A(_f_permutation__round__c[8] ), 
        .ZN(_f_permutation__round__n392 ) );
  INV_X4 _f_permutation__round__U1991  ( .A(_f_permutation__round__c[1481] ), 
        .ZN(_f_permutation__round__n391 ) );
  INV_X4 _f_permutation__round__U1990  ( .A(_f_permutation__round__c[1417] ), 
        .ZN(_f_permutation__round__n390 ) );
  INV_X4 _f_permutation__round__U1989  ( .A(_f_permutation__round__c[1289] ), 
        .ZN(_f_permutation__round__n389 ) );
  INV_X4 _f_permutation__round__U1988  ( .A(_f_permutation__round__c[520] ), 
        .ZN(_f_permutation__round__n388 ) );
  INV_X4 _f_permutation__round__U1987  ( .A(_f_permutation__round__c[456] ), 
        .ZN(_f_permutation__round__n387 ) );
  INV_X4 _f_permutation__round__U1986  ( .A(_f_permutation__round__c[328] ), 
        .ZN(_f_permutation__round__n386 ) );
  INV_X4 _f_permutation__round__U1985  ( .A(_f_permutation__round__c[9] ), 
        .ZN(_f_permutation__round__n385 ) );
  INV_X4 _f_permutation__round__U1984  ( .A(_f_permutation__round__c[1482] ), 
        .ZN(_f_permutation__round__n384 ) );
  INV_X4 _f_permutation__round__U1983  ( .A(_f_permutation__round__c[1418] ), 
        .ZN(_f_permutation__round__n383 ) );
  INV_X4 _f_permutation__round__U1982  ( .A(_f_permutation__round__c[1290] ), 
        .ZN(_f_permutation__round__n382 ) );
  INV_X4 _f_permutation__round__U1981  ( .A(_f_permutation__round__c[521] ), 
        .ZN(_f_permutation__round__n381 ) );
  INV_X4 _f_permutation__round__U1980  ( .A(_f_permutation__round__c[457] ), 
        .ZN(_f_permutation__round__n380 ) );
  INV_X4 _f_permutation__round__U1979  ( .A(_f_permutation__round__c[329] ), 
        .ZN(_f_permutation__round__n379 ) );
  INV_X4 _f_permutation__round__U1978  ( .A(_f_permutation__round__c[10] ), 
        .ZN(_f_permutation__round__n378 ) );
  INV_X4 _f_permutation__round__U1977  ( .A(_f_permutation__round__c[1483] ), 
        .ZN(_f_permutation__round__n377 ) );
  INV_X4 _f_permutation__round__U1976  ( .A(_f_permutation__round__c[1419] ), 
        .ZN(_f_permutation__round__n376 ) );
  INV_X4 _f_permutation__round__U1975  ( .A(_f_permutation__round__c[1291] ), 
        .ZN(_f_permutation__round__n375 ) );
  INV_X4 _f_permutation__round__U1974  ( .A(_f_permutation__round__c[522] ), 
        .ZN(_f_permutation__round__n374 ) );
  INV_X4 _f_permutation__round__U1973  ( .A(_f_permutation__round__c[458] ), 
        .ZN(_f_permutation__round__n373 ) );
  INV_X4 _f_permutation__round__U1972  ( .A(_f_permutation__round__c[330] ), 
        .ZN(_f_permutation__round__n372 ) );
  INV_X4 _f_permutation__round__U1971  ( .A(_f_permutation__round__c[11] ), 
        .ZN(_f_permutation__round__n371 ) );
  INV_X4 _f_permutation__round__U1970  ( .A(_f_permutation__round__c[1484] ), 
        .ZN(_f_permutation__round__n370 ) );
  INV_X4 _f_permutation__round__U1969  ( .A(_f_permutation__round__c[1420] ), 
        .ZN(_f_permutation__round__n369 ) );
  INV_X4 _f_permutation__round__U1968  ( .A(_f_permutation__round__c[1292] ), 
        .ZN(_f_permutation__round__n368 ) );
  INV_X4 _f_permutation__round__U1967  ( .A(_f_permutation__round__c[523] ), 
        .ZN(_f_permutation__round__n367 ) );
  INV_X4 _f_permutation__round__U1966  ( .A(_f_permutation__round__c[459] ), 
        .ZN(_f_permutation__round__n366 ) );
  INV_X4 _f_permutation__round__U1965  ( .A(_f_permutation__round__c[331] ), 
        .ZN(_f_permutation__round__n365 ) );
  INV_X4 _f_permutation__round__U1964  ( .A(_f_permutation__round__c[12] ), 
        .ZN(_f_permutation__round__n364 ) );
  INV_X4 _f_permutation__round__U1963  ( .A(_f_permutation__round__c[1485] ), 
        .ZN(_f_permutation__round__n363 ) );
  INV_X4 _f_permutation__round__U1962  ( .A(_f_permutation__round__c[1421] ), 
        .ZN(_f_permutation__round__n362 ) );
  INV_X4 _f_permutation__round__U1961  ( .A(_f_permutation__round__c[1293] ), 
        .ZN(_f_permutation__round__n361 ) );
  INV_X4 _f_permutation__round__U1960  ( .A(_f_permutation__round__c[524] ), 
        .ZN(_f_permutation__round__n360 ) );
  INV_X4 _f_permutation__round__U1959  ( .A(_f_permutation__round__c[460] ), 
        .ZN(_f_permutation__round__n359 ) );
  INV_X4 _f_permutation__round__U1958  ( .A(_f_permutation__round__c[332] ), 
        .ZN(_f_permutation__round__n358 ) );
  INV_X4 _f_permutation__round__U1957  ( .A(_f_permutation__round__c[13] ), 
        .ZN(_f_permutation__round__n357 ) );
  INV_X4 _f_permutation__round__U1956  ( .A(_f_permutation__round__c[1486] ), 
        .ZN(_f_permutation__round__n356 ) );
  INV_X4 _f_permutation__round__U1955  ( .A(_f_permutation__round__c[1422] ), 
        .ZN(_f_permutation__round__n355 ) );
  INV_X4 _f_permutation__round__U1954  ( .A(_f_permutation__round__c[1294] ), 
        .ZN(_f_permutation__round__n354 ) );
  INV_X4 _f_permutation__round__U1953  ( .A(_f_permutation__round__c[525] ), 
        .ZN(_f_permutation__round__n353 ) );
  INV_X4 _f_permutation__round__U1952  ( .A(_f_permutation__round__c[461] ), 
        .ZN(_f_permutation__round__n352 ) );
  INV_X4 _f_permutation__round__U1951  ( .A(_f_permutation__round__c[333] ), 
        .ZN(_f_permutation__round__n351 ) );
  INV_X4 _f_permutation__round__U1950  ( .A(_f_permutation__round__c[14] ), 
        .ZN(_f_permutation__round__n350 ) );
  INV_X4 _f_permutation__round__U1949  ( .A(_f_permutation__round__c[1487] ), 
        .ZN(_f_permutation__round__n349 ) );
  INV_X4 _f_permutation__round__U1948  ( .A(_f_permutation__round__c[1423] ), 
        .ZN(_f_permutation__round__n348 ) );
  INV_X4 _f_permutation__round__U1947  ( .A(_f_permutation__round__c[1295] ), 
        .ZN(_f_permutation__round__n347 ) );
  INV_X4 _f_permutation__round__U1946  ( .A(_f_permutation__round__c[526] ), 
        .ZN(_f_permutation__round__n346 ) );
  INV_X4 _f_permutation__round__U1945  ( .A(_f_permutation__round__c[462] ), 
        .ZN(_f_permutation__round__n345 ) );
  INV_X4 _f_permutation__round__U1944  ( .A(_f_permutation__round__c[334] ), 
        .ZN(_f_permutation__round__n344 ) );
  INV_X4 _f_permutation__round__U1943  ( .A(_f_permutation__round__c[15] ), 
        .ZN(_f_permutation__round__n343 ) );
  INV_X4 _f_permutation__round__U1942  ( .A(_f_permutation__round__c[1488] ), 
        .ZN(_f_permutation__round__n342 ) );
  INV_X4 _f_permutation__round__U1941  ( .A(_f_permutation__round__c[1424] ), 
        .ZN(_f_permutation__round__n341 ) );
  INV_X4 _f_permutation__round__U1940  ( .A(_f_permutation__round__c[1296] ), 
        .ZN(_f_permutation__round__n340 ) );
  INV_X4 _f_permutation__round__U1939  ( .A(_f_permutation__round__c[527] ), 
        .ZN(_f_permutation__round__n339 ) );
  INV_X4 _f_permutation__round__U1938  ( .A(_f_permutation__round__c[463] ), 
        .ZN(_f_permutation__round__n338 ) );
  INV_X4 _f_permutation__round__U1937  ( .A(_f_permutation__round__c[335] ), 
        .ZN(_f_permutation__round__n337 ) );
  INV_X4 _f_permutation__round__U1936  ( .A(_f_permutation__round__c[16] ), 
        .ZN(_f_permutation__round__n336 ) );
  INV_X4 _f_permutation__round__U1935  ( .A(_f_permutation__round__c[1489] ), 
        .ZN(_f_permutation__round__n335 ) );
  INV_X4 _f_permutation__round__U1934  ( .A(_f_permutation__round__c[1425] ), 
        .ZN(_f_permutation__round__n334 ) );
  INV_X4 _f_permutation__round__U1933  ( .A(_f_permutation__round__c[1297] ), 
        .ZN(_f_permutation__round__n333 ) );
  INV_X4 _f_permutation__round__U1932  ( .A(_f_permutation__round__c[528] ), 
        .ZN(_f_permutation__round__n332 ) );
  INV_X4 _f_permutation__round__U1931  ( .A(_f_permutation__round__c[464] ), 
        .ZN(_f_permutation__round__n331 ) );
  INV_X4 _f_permutation__round__U1930  ( .A(_f_permutation__round__c[336] ), 
        .ZN(_f_permutation__round__n330 ) );
  INV_X4 _f_permutation__round__U1929  ( .A(_f_permutation__round__c[17] ), 
        .ZN(_f_permutation__round__n329 ) );
  INV_X4 _f_permutation__round__U1928  ( .A(_f_permutation__round__c[1490] ), 
        .ZN(_f_permutation__round__n328 ) );
  INV_X4 _f_permutation__round__U1927  ( .A(_f_permutation__round__c[1426] ), 
        .ZN(_f_permutation__round__n327 ) );
  INV_X4 _f_permutation__round__U1926  ( .A(_f_permutation__round__c[1298] ), 
        .ZN(_f_permutation__round__n326 ) );
  INV_X4 _f_permutation__round__U1925  ( .A(_f_permutation__round__c[529] ), 
        .ZN(_f_permutation__round__n325 ) );
  INV_X4 _f_permutation__round__U1924  ( .A(_f_permutation__round__c[465] ), 
        .ZN(_f_permutation__round__n324 ) );
  INV_X4 _f_permutation__round__U1923  ( .A(_f_permutation__round__c[337] ), 
        .ZN(_f_permutation__round__n323 ) );
  INV_X4 _f_permutation__round__U1922  ( .A(_f_permutation__round__c[18] ), 
        .ZN(_f_permutation__round__n322 ) );
  INV_X4 _f_permutation__round__U1921  ( .A(_f_permutation__round__c[1491] ), 
        .ZN(_f_permutation__round__n321 ) );
  INV_X4 _f_permutation__round__U1920  ( .A(_f_permutation__round__c[1427] ), 
        .ZN(_f_permutation__round__n320 ) );
  INV_X4 _f_permutation__round__U1919  ( .A(_f_permutation__round__c[1299] ), 
        .ZN(_f_permutation__round__n319 ) );
  INV_X4 _f_permutation__round__U1918  ( .A(_f_permutation__round__c[530] ), 
        .ZN(_f_permutation__round__n318 ) );
  INV_X4 _f_permutation__round__U1917  ( .A(_f_permutation__round__c[466] ), 
        .ZN(_f_permutation__round__n317 ) );
  INV_X4 _f_permutation__round__U1916  ( .A(_f_permutation__round__c[338] ), 
        .ZN(_f_permutation__round__n316 ) );
  INV_X4 _f_permutation__round__U1915  ( .A(_f_permutation__round__c[19] ), 
        .ZN(_f_permutation__round__n315 ) );
  INV_X4 _f_permutation__round__U1914  ( .A(_f_permutation__round__c[1492] ), 
        .ZN(_f_permutation__round__n314 ) );
  INV_X4 _f_permutation__round__U1913  ( .A(_f_permutation__round__c[1428] ), 
        .ZN(_f_permutation__round__n313 ) );
  INV_X4 _f_permutation__round__U1912  ( .A(_f_permutation__round__c[1300] ), 
        .ZN(_f_permutation__round__n312 ) );
  INV_X4 _f_permutation__round__U1911  ( .A(_f_permutation__round__c[531] ), 
        .ZN(_f_permutation__round__n311 ) );
  INV_X4 _f_permutation__round__U1910  ( .A(_f_permutation__round__c[467] ), 
        .ZN(_f_permutation__round__n310 ) );
  INV_X4 _f_permutation__round__U1909  ( .A(_f_permutation__round__c[339] ), 
        .ZN(_f_permutation__round__n309 ) );
  INV_X4 _f_permutation__round__U1908  ( .A(_f_permutation__round__c[20] ), 
        .ZN(_f_permutation__round__n308 ) );
  INV_X4 _f_permutation__round__U1907  ( .A(_f_permutation__round__c[1493] ), 
        .ZN(_f_permutation__round__n307 ) );
  INV_X4 _f_permutation__round__U1906  ( .A(_f_permutation__round__c[1429] ), 
        .ZN(_f_permutation__round__n306 ) );
  INV_X4 _f_permutation__round__U1905  ( .A(_f_permutation__round__c[1301] ), 
        .ZN(_f_permutation__round__n305 ) );
  INV_X4 _f_permutation__round__U1904  ( .A(_f_permutation__round__c[532] ), 
        .ZN(_f_permutation__round__n304 ) );
  INV_X4 _f_permutation__round__U1903  ( .A(_f_permutation__round__c[468] ), 
        .ZN(_f_permutation__round__n303 ) );
  INV_X4 _f_permutation__round__U1902  ( .A(_f_permutation__round__c[340] ), 
        .ZN(_f_permutation__round__n302 ) );
  INV_X4 _f_permutation__round__U1901  ( .A(_f_permutation__round__c[21] ), 
        .ZN(_f_permutation__round__n301 ) );
  INV_X4 _f_permutation__round__U1900  ( .A(_f_permutation__round__c[1494] ), 
        .ZN(_f_permutation__round__n300 ) );
  INV_X4 _f_permutation__round__U1899  ( .A(_f_permutation__round__c[1430] ), 
        .ZN(_f_permutation__round__n299 ) );
  INV_X4 _f_permutation__round__U1898  ( .A(_f_permutation__round__c[1302] ), 
        .ZN(_f_permutation__round__n298 ) );
  INV_X4 _f_permutation__round__U1897  ( .A(_f_permutation__round__c[533] ), 
        .ZN(_f_permutation__round__n297 ) );
  INV_X4 _f_permutation__round__U1896  ( .A(_f_permutation__round__c[469] ), 
        .ZN(_f_permutation__round__n296 ) );
  INV_X4 _f_permutation__round__U1895  ( .A(_f_permutation__round__c[341] ), 
        .ZN(_f_permutation__round__n295 ) );
  INV_X4 _f_permutation__round__U1894  ( .A(_f_permutation__round__c[22] ), 
        .ZN(_f_permutation__round__n294 ) );
  INV_X4 _f_permutation__round__U1893  ( .A(_f_permutation__round__c[1495] ), 
        .ZN(_f_permutation__round__n293 ) );
  INV_X4 _f_permutation__round__U1892  ( .A(_f_permutation__round__c[1431] ), 
        .ZN(_f_permutation__round__n292 ) );
  INV_X4 _f_permutation__round__U1891  ( .A(_f_permutation__round__c[1303] ), 
        .ZN(_f_permutation__round__n291 ) );
  INV_X4 _f_permutation__round__U1890  ( .A(_f_permutation__round__c[534] ), 
        .ZN(_f_permutation__round__n290 ) );
  INV_X4 _f_permutation__round__U1889  ( .A(_f_permutation__round__c[470] ), 
        .ZN(_f_permutation__round__n289 ) );
  INV_X4 _f_permutation__round__U1888  ( .A(_f_permutation__round__c[342] ), 
        .ZN(_f_permutation__round__n288 ) );
  INV_X4 _f_permutation__round__U1887  ( .A(_f_permutation__round__c[23] ), 
        .ZN(_f_permutation__round__n287 ) );
  INV_X4 _f_permutation__round__U1886  ( .A(_f_permutation__round__c[1496] ), 
        .ZN(_f_permutation__round__n286 ) );
  INV_X4 _f_permutation__round__U1885  ( .A(_f_permutation__round__c[1432] ), 
        .ZN(_f_permutation__round__n285 ) );
  INV_X4 _f_permutation__round__U1884  ( .A(_f_permutation__round__c[1304] ), 
        .ZN(_f_permutation__round__n284 ) );
  INV_X4 _f_permutation__round__U1883  ( .A(_f_permutation__round__c[535] ), 
        .ZN(_f_permutation__round__n283 ) );
  INV_X4 _f_permutation__round__U1882  ( .A(_f_permutation__round__c[471] ), 
        .ZN(_f_permutation__round__n282 ) );
  INV_X4 _f_permutation__round__U1881  ( .A(_f_permutation__round__c[343] ), 
        .ZN(_f_permutation__round__n281 ) );
  INV_X4 _f_permutation__round__U1880  ( .A(_f_permutation__round__c[24] ), 
        .ZN(_f_permutation__round__n280 ) );
  INV_X4 _f_permutation__round__U1879  ( .A(_f_permutation__round__c[1497] ), 
        .ZN(_f_permutation__round__n279 ) );
  INV_X4 _f_permutation__round__U1878  ( .A(_f_permutation__round__c[1433] ), 
        .ZN(_f_permutation__round__n278 ) );
  INV_X4 _f_permutation__round__U1877  ( .A(_f_permutation__round__c[1305] ), 
        .ZN(_f_permutation__round__n277 ) );
  INV_X4 _f_permutation__round__U1876  ( .A(_f_permutation__round__c[536] ), 
        .ZN(_f_permutation__round__n276 ) );
  INV_X4 _f_permutation__round__U1875  ( .A(_f_permutation__round__c[472] ), 
        .ZN(_f_permutation__round__n275 ) );
  INV_X4 _f_permutation__round__U1874  ( .A(_f_permutation__round__c[344] ), 
        .ZN(_f_permutation__round__n274 ) );
  INV_X4 _f_permutation__round__U1873  ( .A(_f_permutation__round__c[25] ), 
        .ZN(_f_permutation__round__n273 ) );
  INV_X4 _f_permutation__round__U1872  ( .A(_f_permutation__round__c[1498] ), 
        .ZN(_f_permutation__round__n272 ) );
  INV_X4 _f_permutation__round__U1871  ( .A(_f_permutation__round__c[1434] ), 
        .ZN(_f_permutation__round__n271 ) );
  INV_X4 _f_permutation__round__U1870  ( .A(_f_permutation__round__c[1306] ), 
        .ZN(_f_permutation__round__n270 ) );
  INV_X4 _f_permutation__round__U1869  ( .A(_f_permutation__round__c[537] ), 
        .ZN(_f_permutation__round__n269 ) );
  INV_X4 _f_permutation__round__U1868  ( .A(_f_permutation__round__c[473] ), 
        .ZN(_f_permutation__round__n268 ) );
  INV_X4 _f_permutation__round__U1867  ( .A(_f_permutation__round__c[345] ), 
        .ZN(_f_permutation__round__n267 ) );
  INV_X4 _f_permutation__round__U1866  ( .A(_f_permutation__round__c[26] ), 
        .ZN(_f_permutation__round__n266 ) );
  INV_X4 _f_permutation__round__U1865  ( .A(_f_permutation__round__c[1499] ), 
        .ZN(_f_permutation__round__n265 ) );
  INV_X4 _f_permutation__round__U1864  ( .A(_f_permutation__round__c[1435] ), 
        .ZN(_f_permutation__round__n264 ) );
  INV_X4 _f_permutation__round__U1863  ( .A(_f_permutation__round__c[1307] ), 
        .ZN(_f_permutation__round__n263 ) );
  INV_X4 _f_permutation__round__U1862  ( .A(_f_permutation__round__c[538] ), 
        .ZN(_f_permutation__round__n262 ) );
  INV_X4 _f_permutation__round__U1861  ( .A(_f_permutation__round__c[474] ), 
        .ZN(_f_permutation__round__n261 ) );
  INV_X4 _f_permutation__round__U1860  ( .A(_f_permutation__round__c[346] ), 
        .ZN(_f_permutation__round__n260 ) );
  INV_X4 _f_permutation__round__U1859  ( .A(_f_permutation__round__c[27] ), 
        .ZN(_f_permutation__round__n259 ) );
  INV_X4 _f_permutation__round__U1858  ( .A(_f_permutation__round__c[1500] ), 
        .ZN(_f_permutation__round__n258 ) );
  INV_X4 _f_permutation__round__U1857  ( .A(_f_permutation__round__c[1436] ), 
        .ZN(_f_permutation__round__n257 ) );
  INV_X4 _f_permutation__round__U1856  ( .A(_f_permutation__round__c[1308] ), 
        .ZN(_f_permutation__round__n256 ) );
  INV_X4 _f_permutation__round__U1855  ( .A(_f_permutation__round__c[539] ), 
        .ZN(_f_permutation__round__n255 ) );
  INV_X4 _f_permutation__round__U1854  ( .A(_f_permutation__round__c[475] ), 
        .ZN(_f_permutation__round__n254 ) );
  INV_X4 _f_permutation__round__U1853  ( .A(_f_permutation__round__c[347] ), 
        .ZN(_f_permutation__round__n253 ) );
  INV_X4 _f_permutation__round__U1852  ( .A(_f_permutation__round__c[28] ), 
        .ZN(_f_permutation__round__n252 ) );
  INV_X4 _f_permutation__round__U1851  ( .A(_f_permutation__round__c[1501] ), 
        .ZN(_f_permutation__round__n251 ) );
  INV_X4 _f_permutation__round__U1850  ( .A(_f_permutation__round__c[1437] ), 
        .ZN(_f_permutation__round__n250 ) );
  INV_X4 _f_permutation__round__U1849  ( .A(_f_permutation__round__c[1309] ), 
        .ZN(_f_permutation__round__n249 ) );
  INV_X4 _f_permutation__round__U1848  ( .A(_f_permutation__round__c[540] ), 
        .ZN(_f_permutation__round__n248 ) );
  INV_X4 _f_permutation__round__U1847  ( .A(_f_permutation__round__c[476] ), 
        .ZN(_f_permutation__round__n247 ) );
  INV_X4 _f_permutation__round__U1846  ( .A(_f_permutation__round__c[348] ), 
        .ZN(_f_permutation__round__n246 ) );
  INV_X4 _f_permutation__round__U1845  ( .A(_f_permutation__round__c[29] ), 
        .ZN(_f_permutation__round__n245 ) );
  INV_X4 _f_permutation__round__U1844  ( .A(_f_permutation__round__c[1502] ), 
        .ZN(_f_permutation__round__n244 ) );
  INV_X4 _f_permutation__round__U1843  ( .A(_f_permutation__round__c[1438] ), 
        .ZN(_f_permutation__round__n243 ) );
  INV_X4 _f_permutation__round__U1842  ( .A(_f_permutation__round__c[1310] ), 
        .ZN(_f_permutation__round__n242 ) );
  INV_X4 _f_permutation__round__U1841  ( .A(_f_permutation__round__c[541] ), 
        .ZN(_f_permutation__round__n241 ) );
  INV_X4 _f_permutation__round__U1840  ( .A(_f_permutation__round__c[477] ), 
        .ZN(_f_permutation__round__n240 ) );
  INV_X4 _f_permutation__round__U1839  ( .A(_f_permutation__round__c[349] ), 
        .ZN(_f_permutation__round__n239 ) );
  INV_X4 _f_permutation__round__U1838  ( .A(_f_permutation__round__c[30] ), 
        .ZN(_f_permutation__round__n238 ) );
  INV_X4 _f_permutation__round__U1837  ( .A(_f_permutation__round__c[1503] ), 
        .ZN(_f_permutation__round__n237 ) );
  INV_X4 _f_permutation__round__U1836  ( .A(_f_permutation__round__c[1439] ), 
        .ZN(_f_permutation__round__n236 ) );
  INV_X4 _f_permutation__round__U1835  ( .A(_f_permutation__round__c[1311] ), 
        .ZN(_f_permutation__round__n235 ) );
  INV_X4 _f_permutation__round__U1834  ( .A(_f_permutation__round__c[542] ), 
        .ZN(_f_permutation__round__n234 ) );
  INV_X4 _f_permutation__round__U1833  ( .A(_f_permutation__round__c[478] ), 
        .ZN(_f_permutation__round__n233 ) );
  INV_X4 _f_permutation__round__U1832  ( .A(_f_permutation__round__c[350] ), 
        .ZN(_f_permutation__round__n232 ) );
  INV_X4 _f_permutation__round__U1831  ( .A(_f_permutation__round__c[31] ), 
        .ZN(_f_permutation__round__n231 ) );
  INV_X4 _f_permutation__round__U1830  ( .A(_f_permutation__round__c[1504] ), 
        .ZN(_f_permutation__round__n230 ) );
  INV_X4 _f_permutation__round__U1829  ( .A(_f_permutation__round__c[1440] ), 
        .ZN(_f_permutation__round__n229 ) );
  INV_X4 _f_permutation__round__U1828  ( .A(_f_permutation__round__c[1312] ), 
        .ZN(_f_permutation__round__n228 ) );
  INV_X4 _f_permutation__round__U1827  ( .A(_f_permutation__round__c[543] ), 
        .ZN(_f_permutation__round__n227 ) );
  INV_X4 _f_permutation__round__U1826  ( .A(_f_permutation__round__c[479] ), 
        .ZN(_f_permutation__round__n226 ) );
  INV_X4 _f_permutation__round__U1825  ( .A(_f_permutation__round__c[351] ), 
        .ZN(_f_permutation__round__n225 ) );
  INV_X4 _f_permutation__round__U1824  ( .A(_f_permutation__round__c[32] ), 
        .ZN(_f_permutation__round__n224 ) );
  INV_X4 _f_permutation__round__U1823  ( .A(_f_permutation__round__c[1505] ), 
        .ZN(_f_permutation__round__n223 ) );
  INV_X4 _f_permutation__round__U1822  ( .A(_f_permutation__round__c[1441] ), 
        .ZN(_f_permutation__round__n222 ) );
  INV_X4 _f_permutation__round__U1821  ( .A(_f_permutation__round__c[1313] ), 
        .ZN(_f_permutation__round__n221 ) );
  INV_X4 _f_permutation__round__U1820  ( .A(_f_permutation__round__c[544] ), 
        .ZN(_f_permutation__round__n220 ) );
  INV_X4 _f_permutation__round__U1819  ( .A(_f_permutation__round__c[480] ), 
        .ZN(_f_permutation__round__n219 ) );
  INV_X4 _f_permutation__round__U1818  ( .A(_f_permutation__round__c[352] ), 
        .ZN(_f_permutation__round__n218 ) );
  INV_X4 _f_permutation__round__U1817  ( .A(_f_permutation__round__c[33] ), 
        .ZN(_f_permutation__round__n217 ) );
  INV_X4 _f_permutation__round__U1816  ( .A(_f_permutation__round__c[1506] ), 
        .ZN(_f_permutation__round__n216 ) );
  INV_X4 _f_permutation__round__U1815  ( .A(_f_permutation__round__c[1442] ), 
        .ZN(_f_permutation__round__n215 ) );
  INV_X4 _f_permutation__round__U1814  ( .A(_f_permutation__round__c[1314] ), 
        .ZN(_f_permutation__round__n214 ) );
  INV_X4 _f_permutation__round__U1813  ( .A(_f_permutation__round__c[545] ), 
        .ZN(_f_permutation__round__n213 ) );
  INV_X4 _f_permutation__round__U1812  ( .A(_f_permutation__round__c[481] ), 
        .ZN(_f_permutation__round__n212 ) );
  INV_X4 _f_permutation__round__U1811  ( .A(_f_permutation__round__c[353] ), 
        .ZN(_f_permutation__round__n211 ) );
  INV_X4 _f_permutation__round__U1810  ( .A(_f_permutation__round__c[34] ), 
        .ZN(_f_permutation__round__n210 ) );
  INV_X4 _f_permutation__round__U1809  ( .A(_f_permutation__round__c[1507] ), 
        .ZN(_f_permutation__round__n209 ) );
  INV_X4 _f_permutation__round__U1808  ( .A(_f_permutation__round__c[1443] ), 
        .ZN(_f_permutation__round__n208 ) );
  INV_X4 _f_permutation__round__U1807  ( .A(_f_permutation__round__c[1315] ), 
        .ZN(_f_permutation__round__n207 ) );
  INV_X4 _f_permutation__round__U1806  ( .A(_f_permutation__round__c[546] ), 
        .ZN(_f_permutation__round__n206 ) );
  INV_X4 _f_permutation__round__U1805  ( .A(_f_permutation__round__c[482] ), 
        .ZN(_f_permutation__round__n205 ) );
  INV_X4 _f_permutation__round__U1804  ( .A(_f_permutation__round__c[354] ), 
        .ZN(_f_permutation__round__n204 ) );
  INV_X4 _f_permutation__round__U1803  ( .A(_f_permutation__round__c[35] ), 
        .ZN(_f_permutation__round__n203 ) );
  INV_X4 _f_permutation__round__U1802  ( .A(_f_permutation__round__c[1508] ), 
        .ZN(_f_permutation__round__n202 ) );
  INV_X4 _f_permutation__round__U1801  ( .A(_f_permutation__round__c[1444] ), 
        .ZN(_f_permutation__round__n201 ) );
  INV_X4 _f_permutation__round__U1800  ( .A(_f_permutation__round__c[1316] ), 
        .ZN(_f_permutation__round__n200 ) );
  INV_X4 _f_permutation__round__U1799  ( .A(_f_permutation__round__c[547] ), 
        .ZN(_f_permutation__round__n199 ) );
  INV_X4 _f_permutation__round__U1798  ( .A(_f_permutation__round__c[483] ), 
        .ZN(_f_permutation__round__n198 ) );
  INV_X4 _f_permutation__round__U1797  ( .A(_f_permutation__round__c[355] ), 
        .ZN(_f_permutation__round__n197 ) );
  INV_X4 _f_permutation__round__U1796  ( .A(_f_permutation__round__c[36] ), 
        .ZN(_f_permutation__round__n196 ) );
  INV_X4 _f_permutation__round__U1795  ( .A(_f_permutation__round__c[1509] ), 
        .ZN(_f_permutation__round__n195 ) );
  INV_X4 _f_permutation__round__U1794  ( .A(_f_permutation__round__c[1445] ), 
        .ZN(_f_permutation__round__n194 ) );
  INV_X4 _f_permutation__round__U1793  ( .A(_f_permutation__round__c[1317] ), 
        .ZN(_f_permutation__round__n193 ) );
  INV_X4 _f_permutation__round__U1792  ( .A(_f_permutation__round__c[548] ), 
        .ZN(_f_permutation__round__n192 ) );
  INV_X4 _f_permutation__round__U1791  ( .A(_f_permutation__round__c[484] ), 
        .ZN(_f_permutation__round__n191 ) );
  INV_X4 _f_permutation__round__U1790  ( .A(_f_permutation__round__c[356] ), 
        .ZN(_f_permutation__round__n190 ) );
  INV_X4 _f_permutation__round__U1789  ( .A(_f_permutation__round__c[37] ), 
        .ZN(_f_permutation__round__n189 ) );
  INV_X4 _f_permutation__round__U1788  ( .A(_f_permutation__round__c[1510] ), 
        .ZN(_f_permutation__round__n188 ) );
  INV_X4 _f_permutation__round__U1787  ( .A(_f_permutation__round__c[1446] ), 
        .ZN(_f_permutation__round__n187 ) );
  INV_X4 _f_permutation__round__U1786  ( .A(_f_permutation__round__c[1318] ), 
        .ZN(_f_permutation__round__n186 ) );
  INV_X4 _f_permutation__round__U1785  ( .A(_f_permutation__round__c[549] ), 
        .ZN(_f_permutation__round__n185 ) );
  INV_X4 _f_permutation__round__U1784  ( .A(_f_permutation__round__c[485] ), 
        .ZN(_f_permutation__round__n184 ) );
  INV_X4 _f_permutation__round__U1783  ( .A(_f_permutation__round__c[357] ), 
        .ZN(_f_permutation__round__n183 ) );
  INV_X4 _f_permutation__round__U1782  ( .A(_f_permutation__round__c[38] ), 
        .ZN(_f_permutation__round__n182 ) );
  INV_X4 _f_permutation__round__U1781  ( .A(_f_permutation__round__c[1511] ), 
        .ZN(_f_permutation__round__n181 ) );
  INV_X4 _f_permutation__round__U1780  ( .A(_f_permutation__round__c[1447] ), 
        .ZN(_f_permutation__round__n180 ) );
  INV_X4 _f_permutation__round__U1779  ( .A(_f_permutation__round__c[1319] ), 
        .ZN(_f_permutation__round__n179 ) );
  INV_X4 _f_permutation__round__U1778  ( .A(_f_permutation__round__c[550] ), 
        .ZN(_f_permutation__round__n178 ) );
  INV_X4 _f_permutation__round__U1777  ( .A(_f_permutation__round__c[486] ), 
        .ZN(_f_permutation__round__n177 ) );
  INV_X4 _f_permutation__round__U1776  ( .A(_f_permutation__round__c[358] ), 
        .ZN(_f_permutation__round__n176 ) );
  INV_X4 _f_permutation__round__U1775  ( .A(_f_permutation__round__c[39] ), 
        .ZN(_f_permutation__round__n175 ) );
  INV_X4 _f_permutation__round__U1774  ( .A(_f_permutation__round__c[1512] ), 
        .ZN(_f_permutation__round__n174 ) );
  INV_X4 _f_permutation__round__U1773  ( .A(_f_permutation__round__c[1448] ), 
        .ZN(_f_permutation__round__n173 ) );
  INV_X4 _f_permutation__round__U1772  ( .A(_f_permutation__round__c[1320] ), 
        .ZN(_f_permutation__round__n172 ) );
  INV_X4 _f_permutation__round__U1771  ( .A(_f_permutation__round__c[551] ), 
        .ZN(_f_permutation__round__n171 ) );
  INV_X4 _f_permutation__round__U1770  ( .A(_f_permutation__round__c[487] ), 
        .ZN(_f_permutation__round__n170 ) );
  INV_X4 _f_permutation__round__U1769  ( .A(_f_permutation__round__c[359] ), 
        .ZN(_f_permutation__round__n169 ) );
  INV_X4 _f_permutation__round__U1768  ( .A(_f_permutation__round__c[40] ), 
        .ZN(_f_permutation__round__n168 ) );
  INV_X4 _f_permutation__round__U1767  ( .A(_f_permutation__round__c[1513] ), 
        .ZN(_f_permutation__round__n167 ) );
  INV_X4 _f_permutation__round__U1766  ( .A(_f_permutation__round__c[1449] ), 
        .ZN(_f_permutation__round__n166 ) );
  INV_X4 _f_permutation__round__U1765  ( .A(_f_permutation__round__c[1321] ), 
        .ZN(_f_permutation__round__n165 ) );
  INV_X4 _f_permutation__round__U1764  ( .A(_f_permutation__round__c[552] ), 
        .ZN(_f_permutation__round__n164 ) );
  INV_X4 _f_permutation__round__U1763  ( .A(_f_permutation__round__c[488] ), 
        .ZN(_f_permutation__round__n163 ) );
  INV_X4 _f_permutation__round__U1762  ( .A(_f_permutation__round__c[360] ), 
        .ZN(_f_permutation__round__n162 ) );
  INV_X4 _f_permutation__round__U1761  ( .A(_f_permutation__round__c[41] ), 
        .ZN(_f_permutation__round__n161 ) );
  INV_X4 _f_permutation__round__U1760  ( .A(_f_permutation__round__c[1514] ), 
        .ZN(_f_permutation__round__n160 ) );
  INV_X4 _f_permutation__round__U1759  ( .A(_f_permutation__round__c[1450] ), 
        .ZN(_f_permutation__round__n159 ) );
  INV_X4 _f_permutation__round__U1758  ( .A(_f_permutation__round__c[1322] ), 
        .ZN(_f_permutation__round__n158 ) );
  INV_X4 _f_permutation__round__U1757  ( .A(_f_permutation__round__c[553] ), 
        .ZN(_f_permutation__round__n157 ) );
  INV_X4 _f_permutation__round__U1756  ( .A(_f_permutation__round__c[489] ), 
        .ZN(_f_permutation__round__n156 ) );
  INV_X4 _f_permutation__round__U1755  ( .A(_f_permutation__round__c[361] ), 
        .ZN(_f_permutation__round__n155 ) );
  INV_X4 _f_permutation__round__U1754  ( .A(_f_permutation__round__c[42] ), 
        .ZN(_f_permutation__round__n154 ) );
  INV_X4 _f_permutation__round__U1753  ( .A(_f_permutation__round__c[1515] ), 
        .ZN(_f_permutation__round__n153 ) );
  INV_X4 _f_permutation__round__U1752  ( .A(_f_permutation__round__c[1451] ), 
        .ZN(_f_permutation__round__n152 ) );
  INV_X4 _f_permutation__round__U1751  ( .A(_f_permutation__round__c[1323] ), 
        .ZN(_f_permutation__round__n151 ) );
  INV_X4 _f_permutation__round__U1750  ( .A(_f_permutation__round__c[554] ), 
        .ZN(_f_permutation__round__n150 ) );
  INV_X4 _f_permutation__round__U1749  ( .A(_f_permutation__round__c[490] ), 
        .ZN(_f_permutation__round__n149 ) );
  INV_X4 _f_permutation__round__U1748  ( .A(_f_permutation__round__c[362] ), 
        .ZN(_f_permutation__round__n148 ) );
  INV_X4 _f_permutation__round__U1747  ( .A(_f_permutation__round__c[43] ), 
        .ZN(_f_permutation__round__n147 ) );
  INV_X4 _f_permutation__round__U1746  ( .A(_f_permutation__round__c[1516] ), 
        .ZN(_f_permutation__round__n146 ) );
  INV_X4 _f_permutation__round__U1745  ( .A(_f_permutation__round__c[1452] ), 
        .ZN(_f_permutation__round__n145 ) );
  INV_X4 _f_permutation__round__U1744  ( .A(_f_permutation__round__c[1324] ), 
        .ZN(_f_permutation__round__n144 ) );
  INV_X4 _f_permutation__round__U1743  ( .A(_f_permutation__round__c[555] ), 
        .ZN(_f_permutation__round__n143 ) );
  INV_X4 _f_permutation__round__U1742  ( .A(_f_permutation__round__c[491] ), 
        .ZN(_f_permutation__round__n142 ) );
  INV_X4 _f_permutation__round__U1741  ( .A(_f_permutation__round__c[363] ), 
        .ZN(_f_permutation__round__n141 ) );
  INV_X4 _f_permutation__round__U1740  ( .A(_f_permutation__round__c[44] ), 
        .ZN(_f_permutation__round__n140 ) );
  INV_X4 _f_permutation__round__U1739  ( .A(_f_permutation__round__c[1517] ), 
        .ZN(_f_permutation__round__n139 ) );
  INV_X4 _f_permutation__round__U1738  ( .A(_f_permutation__round__c[1453] ), 
        .ZN(_f_permutation__round__n138 ) );
  INV_X4 _f_permutation__round__U1737  ( .A(_f_permutation__round__c[1325] ), 
        .ZN(_f_permutation__round__n137 ) );
  INV_X4 _f_permutation__round__U1736  ( .A(_f_permutation__round__c[556] ), 
        .ZN(_f_permutation__round__n136 ) );
  INV_X4 _f_permutation__round__U1735  ( .A(_f_permutation__round__c[492] ), 
        .ZN(_f_permutation__round__n135 ) );
  INV_X4 _f_permutation__round__U1734  ( .A(_f_permutation__round__c[364] ), 
        .ZN(_f_permutation__round__n134 ) );
  INV_X4 _f_permutation__round__U1733  ( .A(_f_permutation__round__c[45] ), 
        .ZN(_f_permutation__round__n133 ) );
  INV_X4 _f_permutation__round__U1732  ( .A(_f_permutation__round__c[1518] ), 
        .ZN(_f_permutation__round__n132 ) );
  INV_X4 _f_permutation__round__U1731  ( .A(_f_permutation__round__c[1454] ), 
        .ZN(_f_permutation__round__n131 ) );
  INV_X4 _f_permutation__round__U1730  ( .A(_f_permutation__round__c[1326] ), 
        .ZN(_f_permutation__round__n130 ) );
  INV_X4 _f_permutation__round__U1729  ( .A(_f_permutation__round__c[557] ), 
        .ZN(_f_permutation__round__n129 ) );
  INV_X4 _f_permutation__round__U1728  ( .A(_f_permutation__round__c[493] ), 
        .ZN(_f_permutation__round__n128 ) );
  INV_X4 _f_permutation__round__U1727  ( .A(_f_permutation__round__c[365] ), 
        .ZN(_f_permutation__round__n127 ) );
  INV_X4 _f_permutation__round__U1726  ( .A(_f_permutation__round__c[46] ), 
        .ZN(_f_permutation__round__n126 ) );
  INV_X4 _f_permutation__round__U1725  ( .A(_f_permutation__round__c[1519] ), 
        .ZN(_f_permutation__round__n125 ) );
  INV_X4 _f_permutation__round__U1724  ( .A(_f_permutation__round__c[1455] ), 
        .ZN(_f_permutation__round__n124 ) );
  INV_X4 _f_permutation__round__U1723  ( .A(_f_permutation__round__c[1327] ), 
        .ZN(_f_permutation__round__n123 ) );
  INV_X4 _f_permutation__round__U1722  ( .A(_f_permutation__round__c[558] ), 
        .ZN(_f_permutation__round__n122 ) );
  INV_X4 _f_permutation__round__U1721  ( .A(_f_permutation__round__c[494] ), 
        .ZN(_f_permutation__round__n121 ) );
  INV_X4 _f_permutation__round__U1720  ( .A(_f_permutation__round__c[366] ), 
        .ZN(_f_permutation__round__n120 ) );
  INV_X4 _f_permutation__round__U1719  ( .A(_f_permutation__round__c[47] ), 
        .ZN(_f_permutation__round__n119 ) );
  INV_X4 _f_permutation__round__U1718  ( .A(_f_permutation__round__c[1520] ), 
        .ZN(_f_permutation__round__n118 ) );
  INV_X4 _f_permutation__round__U1717  ( .A(_f_permutation__round__c[1456] ), 
        .ZN(_f_permutation__round__n117 ) );
  INV_X4 _f_permutation__round__U1716  ( .A(_f_permutation__round__c[1328] ), 
        .ZN(_f_permutation__round__n116 ) );
  INV_X4 _f_permutation__round__U1715  ( .A(_f_permutation__round__c[559] ), 
        .ZN(_f_permutation__round__n115 ) );
  INV_X4 _f_permutation__round__U1714  ( .A(_f_permutation__round__c[495] ), 
        .ZN(_f_permutation__round__n114 ) );
  INV_X4 _f_permutation__round__U1713  ( .A(_f_permutation__round__c[367] ), 
        .ZN(_f_permutation__round__n113 ) );
  INV_X4 _f_permutation__round__U1712  ( .A(_f_permutation__round__c[48] ), 
        .ZN(_f_permutation__round__n112 ) );
  INV_X4 _f_permutation__round__U1711  ( .A(_f_permutation__round__c[1521] ), 
        .ZN(_f_permutation__round__n111 ) );
  INV_X4 _f_permutation__round__U1710  ( .A(_f_permutation__round__c[1457] ), 
        .ZN(_f_permutation__round__n110 ) );
  INV_X4 _f_permutation__round__U1709  ( .A(_f_permutation__round__c[1329] ), 
        .ZN(_f_permutation__round__n109 ) );
  INV_X4 _f_permutation__round__U1708  ( .A(_f_permutation__round__c[560] ), 
        .ZN(_f_permutation__round__n108 ) );
  INV_X4 _f_permutation__round__U1707  ( .A(_f_permutation__round__c[496] ), 
        .ZN(_f_permutation__round__n107 ) );
  INV_X4 _f_permutation__round__U1706  ( .A(_f_permutation__round__c[368] ), 
        .ZN(_f_permutation__round__n106 ) );
  INV_X4 _f_permutation__round__U1705  ( .A(_f_permutation__round__c[49] ), 
        .ZN(_f_permutation__round__n105 ) );
  INV_X4 _f_permutation__round__U1704  ( .A(_f_permutation__round__c[1522] ), 
        .ZN(_f_permutation__round__n104 ) );
  INV_X4 _f_permutation__round__U1703  ( .A(_f_permutation__round__c[1458] ), 
        .ZN(_f_permutation__round__n103 ) );
  INV_X4 _f_permutation__round__U1702  ( .A(_f_permutation__round__c[1330] ), 
        .ZN(_f_permutation__round__n102 ) );
  INV_X4 _f_permutation__round__U1701  ( .A(_f_permutation__round__c[561] ), 
        .ZN(_f_permutation__round__n101 ) );
  INV_X4 _f_permutation__round__U1700  ( .A(_f_permutation__round__c[497] ), 
        .ZN(_f_permutation__round__n100 ) );
  INV_X4 _f_permutation__round__U1699  ( .A(_f_permutation__round__c[369] ), 
        .ZN(_f_permutation__round__n99 ) );
  INV_X4 _f_permutation__round__U1698  ( .A(_f_permutation__round__c[50] ), 
        .ZN(_f_permutation__round__n98 ) );
  INV_X4 _f_permutation__round__U1697  ( .A(_f_permutation__round__c[1523] ), 
        .ZN(_f_permutation__round__n97 ) );
  INV_X4 _f_permutation__round__U1696  ( .A(_f_permutation__round__c[1459] ), 
        .ZN(_f_permutation__round__n96 ) );
  INV_X4 _f_permutation__round__U1695  ( .A(_f_permutation__round__c[1331] ), 
        .ZN(_f_permutation__round__n95 ) );
  INV_X4 _f_permutation__round__U1694  ( .A(_f_permutation__round__c[562] ), 
        .ZN(_f_permutation__round__n94 ) );
  INV_X4 _f_permutation__round__U1693  ( .A(_f_permutation__round__c[498] ), 
        .ZN(_f_permutation__round__n93 ) );
  INV_X4 _f_permutation__round__U1692  ( .A(_f_permutation__round__c[370] ), 
        .ZN(_f_permutation__round__n92 ) );
  INV_X4 _f_permutation__round__U1691  ( .A(_f_permutation__round__c[51] ), 
        .ZN(_f_permutation__round__n91 ) );
  INV_X4 _f_permutation__round__U1690  ( .A(_f_permutation__round__c[1524] ), 
        .ZN(_f_permutation__round__n90 ) );
  INV_X4 _f_permutation__round__U1689  ( .A(_f_permutation__round__c[1460] ), 
        .ZN(_f_permutation__round__n89 ) );
  INV_X4 _f_permutation__round__U1688  ( .A(_f_permutation__round__c[1332] ), 
        .ZN(_f_permutation__round__n88 ) );
  INV_X4 _f_permutation__round__U1687  ( .A(_f_permutation__round__c[563] ), 
        .ZN(_f_permutation__round__n87 ) );
  INV_X4 _f_permutation__round__U1686  ( .A(_f_permutation__round__c[499] ), 
        .ZN(_f_permutation__round__n86 ) );
  INV_X4 _f_permutation__round__U1685  ( .A(_f_permutation__round__c[371] ), 
        .ZN(_f_permutation__round__n85 ) );
  INV_X4 _f_permutation__round__U1684  ( .A(_f_permutation__round__c[52] ), 
        .ZN(_f_permutation__round__n84 ) );
  INV_X4 _f_permutation__round__U1683  ( .A(_f_permutation__round__c[1525] ), 
        .ZN(_f_permutation__round__n83 ) );
  INV_X4 _f_permutation__round__U1682  ( .A(_f_permutation__round__c[1461] ), 
        .ZN(_f_permutation__round__n82 ) );
  INV_X4 _f_permutation__round__U1681  ( .A(_f_permutation__round__c[1333] ), 
        .ZN(_f_permutation__round__n81 ) );
  INV_X4 _f_permutation__round__U1680  ( .A(_f_permutation__round__c[564] ), 
        .ZN(_f_permutation__round__n80 ) );
  INV_X4 _f_permutation__round__U1679  ( .A(_f_permutation__round__c[500] ), 
        .ZN(_f_permutation__round__n79 ) );
  INV_X4 _f_permutation__round__U1678  ( .A(_f_permutation__round__c[372] ), 
        .ZN(_f_permutation__round__n78 ) );
  INV_X4 _f_permutation__round__U1677  ( .A(_f_permutation__round__c[53] ), 
        .ZN(_f_permutation__round__n77 ) );
  INV_X4 _f_permutation__round__U1676  ( .A(_f_permutation__round__c[1526] ), 
        .ZN(_f_permutation__round__n76 ) );
  INV_X4 _f_permutation__round__U1675  ( .A(_f_permutation__round__c[1462] ), 
        .ZN(_f_permutation__round__n75 ) );
  INV_X4 _f_permutation__round__U1674  ( .A(_f_permutation__round__c[1334] ), 
        .ZN(_f_permutation__round__n74 ) );
  INV_X4 _f_permutation__round__U1673  ( .A(_f_permutation__round__c[565] ), 
        .ZN(_f_permutation__round__n73 ) );
  INV_X4 _f_permutation__round__U1672  ( .A(_f_permutation__round__c[501] ), 
        .ZN(_f_permutation__round__n72 ) );
  INV_X4 _f_permutation__round__U1671  ( .A(_f_permutation__round__c[373] ), 
        .ZN(_f_permutation__round__n71 ) );
  INV_X4 _f_permutation__round__U1670  ( .A(_f_permutation__round__c[54] ), 
        .ZN(_f_permutation__round__n70 ) );
  INV_X4 _f_permutation__round__U1669  ( .A(_f_permutation__round__c[1527] ), 
        .ZN(_f_permutation__round__n69 ) );
  INV_X4 _f_permutation__round__U1668  ( .A(_f_permutation__round__c[1463] ), 
        .ZN(_f_permutation__round__n68 ) );
  INV_X4 _f_permutation__round__U1667  ( .A(_f_permutation__round__c[1335] ), 
        .ZN(_f_permutation__round__n67 ) );
  INV_X4 _f_permutation__round__U1666  ( .A(_f_permutation__round__c[566] ), 
        .ZN(_f_permutation__round__n66 ) );
  INV_X4 _f_permutation__round__U1665  ( .A(_f_permutation__round__c[502] ), 
        .ZN(_f_permutation__round__n65 ) );
  INV_X4 _f_permutation__round__U1664  ( .A(_f_permutation__round__c[374] ), 
        .ZN(_f_permutation__round__n64 ) );
  INV_X4 _f_permutation__round__U1663  ( .A(_f_permutation__round__c[55] ), 
        .ZN(_f_permutation__round__n63 ) );
  INV_X4 _f_permutation__round__U1662  ( .A(_f_permutation__round__c[1528] ), 
        .ZN(_f_permutation__round__n62 ) );
  INV_X4 _f_permutation__round__U1661  ( .A(_f_permutation__round__c[1464] ), 
        .ZN(_f_permutation__round__n61 ) );
  INV_X4 _f_permutation__round__U1660  ( .A(_f_permutation__round__c[1336] ), 
        .ZN(_f_permutation__round__n60 ) );
  INV_X4 _f_permutation__round__U1659  ( .A(_f_permutation__round__c[567] ), 
        .ZN(_f_permutation__round__n59 ) );
  INV_X4 _f_permutation__round__U1658  ( .A(_f_permutation__round__c[503] ), 
        .ZN(_f_permutation__round__n58 ) );
  INV_X4 _f_permutation__round__U1657  ( .A(_f_permutation__round__c[375] ), 
        .ZN(_f_permutation__round__n57 ) );
  INV_X4 _f_permutation__round__U1656  ( .A(_f_permutation__round__c[56] ), 
        .ZN(_f_permutation__round__n56 ) );
  INV_X4 _f_permutation__round__U1655  ( .A(_f_permutation__round__c[1529] ), 
        .ZN(_f_permutation__round__n55 ) );
  INV_X4 _f_permutation__round__U1654  ( .A(_f_permutation__round__c[1465] ), 
        .ZN(_f_permutation__round__n54 ) );
  INV_X4 _f_permutation__round__U1653  ( .A(_f_permutation__round__c[1337] ), 
        .ZN(_f_permutation__round__n53 ) );
  INV_X4 _f_permutation__round__U1652  ( .A(_f_permutation__round__c[568] ), 
        .ZN(_f_permutation__round__n52 ) );
  INV_X4 _f_permutation__round__U1651  ( .A(_f_permutation__round__c[504] ), 
        .ZN(_f_permutation__round__n51 ) );
  INV_X4 _f_permutation__round__U1650  ( .A(_f_permutation__round__c[376] ), 
        .ZN(_f_permutation__round__n50 ) );
  INV_X4 _f_permutation__round__U1649  ( .A(_f_permutation__round__c[57] ), 
        .ZN(_f_permutation__round__n49 ) );
  INV_X4 _f_permutation__round__U1648  ( .A(_f_permutation__round__c[1530] ), 
        .ZN(_f_permutation__round__n48 ) );
  INV_X4 _f_permutation__round__U1647  ( .A(_f_permutation__round__c[1466] ), 
        .ZN(_f_permutation__round__n47 ) );
  INV_X4 _f_permutation__round__U1646  ( .A(_f_permutation__round__c[1338] ), 
        .ZN(_f_permutation__round__n46 ) );
  INV_X4 _f_permutation__round__U1645  ( .A(_f_permutation__round__c[569] ), 
        .ZN(_f_permutation__round__n45 ) );
  INV_X4 _f_permutation__round__U1644  ( .A(_f_permutation__round__c[505] ), 
        .ZN(_f_permutation__round__n44 ) );
  INV_X4 _f_permutation__round__U1643  ( .A(_f_permutation__round__c[377] ), 
        .ZN(_f_permutation__round__n43 ) );
  INV_X4 _f_permutation__round__U1642  ( .A(_f_permutation__round__c[58] ), 
        .ZN(_f_permutation__round__n42 ) );
  INV_X4 _f_permutation__round__U1641  ( .A(_f_permutation__round__c[1531] ), 
        .ZN(_f_permutation__round__n41 ) );
  INV_X4 _f_permutation__round__U1640  ( .A(_f_permutation__round__c[1467] ), 
        .ZN(_f_permutation__round__n40 ) );
  INV_X4 _f_permutation__round__U1639  ( .A(_f_permutation__round__c[1339] ), 
        .ZN(_f_permutation__round__n39 ) );
  INV_X4 _f_permutation__round__U1638  ( .A(_f_permutation__round__c[570] ), 
        .ZN(_f_permutation__round__n38 ) );
  INV_X4 _f_permutation__round__U1637  ( .A(_f_permutation__round__c[506] ), 
        .ZN(_f_permutation__round__n37 ) );
  INV_X4 _f_permutation__round__U1636  ( .A(_f_permutation__round__c[378] ), 
        .ZN(_f_permutation__round__n36 ) );
  INV_X4 _f_permutation__round__U1635  ( .A(_f_permutation__round__c[59] ), 
        .ZN(_f_permutation__round__n35 ) );
  INV_X4 _f_permutation__round__U1634  ( .A(_f_permutation__round__c[1532] ), 
        .ZN(_f_permutation__round__n34 ) );
  INV_X4 _f_permutation__round__U1633  ( .A(_f_permutation__round__c[1468] ), 
        .ZN(_f_permutation__round__n33 ) );
  INV_X4 _f_permutation__round__U1632  ( .A(_f_permutation__round__c[1340] ), 
        .ZN(_f_permutation__round__n32 ) );
  INV_X4 _f_permutation__round__U1631  ( .A(_f_permutation__round__c[571] ), 
        .ZN(_f_permutation__round__n31 ) );
  INV_X4 _f_permutation__round__U1630  ( .A(_f_permutation__round__c[507] ), 
        .ZN(_f_permutation__round__n30 ) );
  INV_X4 _f_permutation__round__U1629  ( .A(_f_permutation__round__c[379] ), 
        .ZN(_f_permutation__round__n29 ) );
  INV_X4 _f_permutation__round__U1628  ( .A(_f_permutation__round__c[60] ), 
        .ZN(_f_permutation__round__n28 ) );
  INV_X4 _f_permutation__round__U1627  ( .A(_f_permutation__round__c[1533] ), 
        .ZN(_f_permutation__round__n27 ) );
  INV_X4 _f_permutation__round__U1626  ( .A(_f_permutation__round__c[1469] ), 
        .ZN(_f_permutation__round__n26 ) );
  INV_X4 _f_permutation__round__U1625  ( .A(_f_permutation__round__c[1341] ), 
        .ZN(_f_permutation__round__n25 ) );
  INV_X4 _f_permutation__round__U1624  ( .A(_f_permutation__round__c[572] ), 
        .ZN(_f_permutation__round__n24 ) );
  INV_X4 _f_permutation__round__U1623  ( .A(_f_permutation__round__c[508] ), 
        .ZN(_f_permutation__round__n23 ) );
  INV_X4 _f_permutation__round__U1622  ( .A(_f_permutation__round__c[380] ), 
        .ZN(_f_permutation__round__n22 ) );
  INV_X4 _f_permutation__round__U1621  ( .A(_f_permutation__round__c[61] ), 
        .ZN(_f_permutation__round__n21 ) );
  INV_X4 _f_permutation__round__U1620  ( .A(_f_permutation__round__c[1534] ), 
        .ZN(_f_permutation__round__n20 ) );
  INV_X4 _f_permutation__round__U1619  ( .A(_f_permutation__round__c[1470] ), 
        .ZN(_f_permutation__round__n19 ) );
  INV_X4 _f_permutation__round__U1618  ( .A(_f_permutation__round__c[1342] ), 
        .ZN(_f_permutation__round__n18 ) );
  INV_X4 _f_permutation__round__U1617  ( .A(_f_permutation__round__c[573] ), 
        .ZN(_f_permutation__round__n17 ) );
  INV_X4 _f_permutation__round__U1616  ( .A(_f_permutation__round__c[509] ), 
        .ZN(_f_permutation__round__n16 ) );
  INV_X4 _f_permutation__round__U1615  ( .A(_f_permutation__round__c[381] ), 
        .ZN(_f_permutation__round__n15 ) );
  INV_X4 _f_permutation__round__U1614  ( .A(_f_permutation__round__c[62] ), 
        .ZN(_f_permutation__round__n14 ) );
  INV_X4 _f_permutation__round__U1613  ( .A(_f_permutation__round__c[1535] ), 
        .ZN(_f_permutation__round__n13 ) );
  INV_X4 _f_permutation__round__U1612  ( .A(_f_permutation__round__c[1471] ), 
        .ZN(_f_permutation__round__n12 ) );
  INV_X4 _f_permutation__round__U1611  ( .A(_f_permutation__round__c[1343] ), 
        .ZN(_f_permutation__round__n11 ) );
  INV_X4 _f_permutation__round__U1610  ( .A(_f_permutation__round__c[574] ), 
        .ZN(_f_permutation__round__n10 ) );
  INV_X4 _f_permutation__round__U1609  ( .A(_f_permutation__round__c[510] ), 
        .ZN(_f_permutation__round__n9 ) );
  INV_X4 _f_permutation__round__U1608  ( .A(_f_permutation__round__c[382] ), 
        .ZN(_f_permutation__round__n8 ) );
  INV_X4 _f_permutation__round__U1607  ( .A(_f_permutation__round__c[63] ), 
        .ZN(_f_permutation__round__n7 ) );
  INV_X4 _f_permutation__round__U1606  ( .A(_f_permutation__round__c[1472] ), 
        .ZN(_f_permutation__round__n6 ) );
  INV_X4 _f_permutation__round__U1605  ( .A(_f_permutation__round__c[1408] ), 
        .ZN(_f_permutation__round__n5 ) );
  INV_X4 _f_permutation__round__U1604  ( .A(_f_permutation__round__c[1280] ), 
        .ZN(_f_permutation__round__n4 ) );
  INV_X4 _f_permutation__round__U1603  ( .A(_f_permutation__round__c[575] ), 
        .ZN(_f_permutation__round__n3 ) );
  INV_X4 _f_permutation__round__U1602  ( .A(_f_permutation__round__c[511] ), 
        .ZN(_f_permutation__round__n2 ) );
  INV_X4 _f_permutation__round__U1601  ( .A(_f_permutation__round__c[383] ), 
        .ZN(_f_permutation__round__n1 ) );
  AND2_X2 _f_permutation__round__U1472  ( .A1(_f_permutation__round__n834 ), 
        .A2(_f_permutation__round__c[1585] ), .ZN(
        _f_permutation__round__N2817 ) );
  AND2_X2 _f_permutation__round__U1471  ( .A1(_f_permutation__round__n837 ), 
        .A2(_f_permutation__round__c[1584] ), .ZN(
        _f_permutation__round__N2819 ) );
  AND2_X2 _f_permutation__round__U1470  ( .A1(_f_permutation__round__n840 ), 
        .A2(_f_permutation__round__c[1583] ), .ZN(
        _f_permutation__round__N2821 ) );
  AND2_X2 _f_permutation__round__U1469  ( .A1(_f_permutation__round__n843 ), 
        .A2(_f_permutation__round__c[1582] ), .ZN(
        _f_permutation__round__N2823 ) );
  AND2_X2 _f_permutation__round__U1468  ( .A1(_f_permutation__round__n846 ), 
        .A2(_f_permutation__round__c[1581] ), .ZN(
        _f_permutation__round__N2825 ) );
  AND2_X2 _f_permutation__round__U1467  ( .A1(_f_permutation__round__n849 ), 
        .A2(_f_permutation__round__c[1580] ), .ZN(
        _f_permutation__round__N2827 ) );
  AND2_X2 _f_permutation__round__U1466  ( .A1(_f_permutation__round__n852 ), 
        .A2(_f_permutation__round__c[1579] ), .ZN(
        _f_permutation__round__N2829 ) );
  AND2_X2 _f_permutation__round__U1465  ( .A1(_f_permutation__round__n855 ), 
        .A2(_f_permutation__round__c[1578] ), .ZN(
        _f_permutation__round__N2831 ) );
  AND2_X2 _f_permutation__round__U1464  ( .A1(_f_permutation__round__n858 ), 
        .A2(_f_permutation__round__c[1577] ), .ZN(
        _f_permutation__round__N2833 ) );
  AND2_X2 _f_permutation__round__U1463  ( .A1(_f_permutation__round__n861 ), 
        .A2(_f_permutation__round__c[1576] ), .ZN(
        _f_permutation__round__N2835 ) );
  AND2_X2 _f_permutation__round__U1462  ( .A1(_f_permutation__round__n864 ), 
        .A2(_f_permutation__round__c[1575] ), .ZN(
        _f_permutation__round__N2837 ) );
  AND2_X2 _f_permutation__round__U1461  ( .A1(_f_permutation__round__n867 ), 
        .A2(_f_permutation__round__c[1574] ), .ZN(
        _f_permutation__round__N2839 ) );
  AND2_X2 _f_permutation__round__U1460  ( .A1(_f_permutation__round__n870 ), 
        .A2(_f_permutation__round__c[1573] ), .ZN(
        _f_permutation__round__N2841 ) );
  AND2_X2 _f_permutation__round__U1459  ( .A1(_f_permutation__round__n873 ), 
        .A2(_f_permutation__round__c[1572] ), .ZN(
        _f_permutation__round__N2843 ) );
  AND2_X2 _f_permutation__round__U1458  ( .A1(_f_permutation__round__n876 ), 
        .A2(_f_permutation__round__c[1571] ), .ZN(
        _f_permutation__round__N2845 ) );
  AND2_X2 _f_permutation__round__U1457  ( .A1(_f_permutation__round__n879 ), 
        .A2(_f_permutation__round__c[1570] ), .ZN(
        _f_permutation__round__N2847 ) );
  AND2_X2 _f_permutation__round__U1456  ( .A1(_f_permutation__round__n882 ), 
        .A2(_f_permutation__round__c[1569] ), .ZN(
        _f_permutation__round__N2849 ) );
  AND2_X2 _f_permutation__round__U1455  ( .A1(_f_permutation__round__n885 ), 
        .A2(_f_permutation__round__c[1568] ), .ZN(
        _f_permutation__round__N2851 ) );
  AND2_X2 _f_permutation__round__U1454  ( .A1(_f_permutation__round__n888 ), 
        .A2(_f_permutation__round__c[1567] ), .ZN(
        _f_permutation__round__N2853 ) );
  AND2_X2 _f_permutation__round__U1453  ( .A1(_f_permutation__round__n891 ), 
        .A2(_f_permutation__round__c[1566] ), .ZN(
        _f_permutation__round__N2855 ) );
  AND2_X2 _f_permutation__round__U1452  ( .A1(_f_permutation__round__n894 ), 
        .A2(_f_permutation__round__c[1565] ), .ZN(
        _f_permutation__round__N2857 ) );
  AND2_X2 _f_permutation__round__U1451  ( .A1(_f_permutation__round__n897 ), 
        .A2(_f_permutation__round__c[1564] ), .ZN(
        _f_permutation__round__N2859 ) );
  AND2_X2 _f_permutation__round__U1450  ( .A1(_f_permutation__round__n900 ), 
        .A2(_f_permutation__round__c[1563] ), .ZN(
        _f_permutation__round__N2861 ) );
  AND2_X2 _f_permutation__round__U1449  ( .A1(_f_permutation__round__n903 ), 
        .A2(_f_permutation__round__c[1562] ), .ZN(
        _f_permutation__round__N2863 ) );
  AND2_X2 _f_permutation__round__U1448  ( .A1(_f_permutation__round__n906 ), 
        .A2(_f_permutation__round__c[1561] ), .ZN(
        _f_permutation__round__N2865 ) );
  AND2_X2 _f_permutation__round__U1447  ( .A1(_f_permutation__round__n909 ), 
        .A2(_f_permutation__round__c[1560] ), .ZN(
        _f_permutation__round__N2867 ) );
  AND2_X2 _f_permutation__round__U1446  ( .A1(_f_permutation__round__n912 ), 
        .A2(_f_permutation__round__c[1559] ), .ZN(
        _f_permutation__round__N2869 ) );
  AND2_X2 _f_permutation__round__U1445  ( .A1(_f_permutation__round__n915 ), 
        .A2(_f_permutation__round__c[1558] ), .ZN(
        _f_permutation__round__N2871 ) );
  AND2_X2 _f_permutation__round__U1444  ( .A1(_f_permutation__round__n918 ), 
        .A2(_f_permutation__round__c[1557] ), .ZN(
        _f_permutation__round__N2873 ) );
  AND2_X2 _f_permutation__round__U1443  ( .A1(_f_permutation__round__n921 ), 
        .A2(_f_permutation__round__c[1556] ), .ZN(
        _f_permutation__round__N2875 ) );
  AND2_X2 _f_permutation__round__U1442  ( .A1(_f_permutation__round__n924 ), 
        .A2(_f_permutation__round__c[1555] ), .ZN(
        _f_permutation__round__N2877 ) );
  AND2_X2 _f_permutation__round__U1441  ( .A1(_f_permutation__round__n927 ), 
        .A2(_f_permutation__round__c[1554] ), .ZN(
        _f_permutation__round__N2879 ) );
  AND2_X2 _f_permutation__round__U1440  ( .A1(_f_permutation__round__n930 ), 
        .A2(_f_permutation__round__c[1553] ), .ZN(
        _f_permutation__round__N2881 ) );
  AND2_X2 _f_permutation__round__U1439  ( .A1(_f_permutation__round__n933 ), 
        .A2(_f_permutation__round__c[1552] ), .ZN(
        _f_permutation__round__N2883 ) );
  AND2_X2 _f_permutation__round__U1438  ( .A1(_f_permutation__round__n936 ), 
        .A2(_f_permutation__round__c[1551] ), .ZN(
        _f_permutation__round__N2885 ) );
  AND2_X2 _f_permutation__round__U1437  ( .A1(_f_permutation__round__n939 ), 
        .A2(_f_permutation__round__c[1550] ), .ZN(
        _f_permutation__round__N2887 ) );
  AND2_X2 _f_permutation__round__U1436  ( .A1(_f_permutation__round__n942 ), 
        .A2(_f_permutation__round__c[1549] ), .ZN(
        _f_permutation__round__N2889 ) );
  AND2_X2 _f_permutation__round__U1435  ( .A1(_f_permutation__round__n945 ), 
        .A2(_f_permutation__round__c[1548] ), .ZN(
        _f_permutation__round__N2891 ) );
  AND2_X2 _f_permutation__round__U1434  ( .A1(_f_permutation__round__n948 ), 
        .A2(_f_permutation__round__c[1547] ), .ZN(
        _f_permutation__round__N2893 ) );
  AND2_X2 _f_permutation__round__U1433  ( .A1(_f_permutation__round__n951 ), 
        .A2(_f_permutation__round__c[1546] ), .ZN(
        _f_permutation__round__N2895 ) );
  AND2_X2 _f_permutation__round__U1432  ( .A1(_f_permutation__round__n954 ), 
        .A2(_f_permutation__round__c[1545] ), .ZN(
        _f_permutation__round__N2897 ) );
  AND2_X2 _f_permutation__round__U1431  ( .A1(_f_permutation__round__n957 ), 
        .A2(_f_permutation__round__c[1544] ), .ZN(
        _f_permutation__round__N2899 ) );
  AND2_X2 _f_permutation__round__U1430  ( .A1(_f_permutation__round__n960 ), 
        .A2(_f_permutation__round__c[1543] ), .ZN(
        _f_permutation__round__N2901 ) );
  AND2_X2 _f_permutation__round__U1429  ( .A1(_f_permutation__round__n771 ), 
        .A2(_f_permutation__round__c[1542] ), .ZN(
        _f_permutation__round__N2903 ) );
  AND2_X2 _f_permutation__round__U1428  ( .A1(_f_permutation__round__n774 ), 
        .A2(_f_permutation__round__c[1541] ), .ZN(
        _f_permutation__round__N2905 ) );
  AND2_X2 _f_permutation__round__U1427  ( .A1(_f_permutation__round__n777 ), 
        .A2(_f_permutation__round__c[1540] ), .ZN(
        _f_permutation__round__N2907 ) );
  AND2_X2 _f_permutation__round__U1426  ( .A1(_f_permutation__round__n780 ), 
        .A2(_f_permutation__round__c[1539] ), .ZN(
        _f_permutation__round__N2909 ) );
  AND2_X2 _f_permutation__round__U1425  ( .A1(_f_permutation__round__n783 ), 
        .A2(_f_permutation__round__c[1538] ), .ZN(
        _f_permutation__round__N2911 ) );
  AND2_X2 _f_permutation__round__U1424  ( .A1(_f_permutation__round__n786 ), 
        .A2(_f_permutation__round__c[1537] ), .ZN(
        _f_permutation__round__N2913 ) );
  AND2_X2 _f_permutation__round__U1423  ( .A1(_f_permutation__round__n789 ), 
        .A2(_f_permutation__round__c[1536] ), .ZN(
        _f_permutation__round__N2915 ) );
  AND2_X2 _f_permutation__round__U1422  ( .A1(_f_permutation__round__n792 ), 
        .A2(_f_permutation__round__c[1599] ), .ZN(
        _f_permutation__round__N2917 ) );
  AND2_X2 _f_permutation__round__U1421  ( .A1(_f_permutation__round__n795 ), 
        .A2(_f_permutation__round__c[1598] ), .ZN(
        _f_permutation__round__N2919 ) );
  AND2_X2 _f_permutation__round__U1420  ( .A1(_f_permutation__round__n798 ), 
        .A2(_f_permutation__round__c[1597] ), .ZN(
        _f_permutation__round__N2921 ) );
  AND2_X2 _f_permutation__round__U1419  ( .A1(_f_permutation__round__n801 ), 
        .A2(_f_permutation__round__c[1596] ), .ZN(
        _f_permutation__round__N2923 ) );
  AND2_X2 _f_permutation__round__U1418  ( .A1(_f_permutation__round__n804 ), 
        .A2(_f_permutation__round__c[1595] ), .ZN(
        _f_permutation__round__N2925 ) );
  AND2_X2 _f_permutation__round__U1417  ( .A1(_f_permutation__round__n807 ), 
        .A2(_f_permutation__round__c[1594] ), .ZN(
        _f_permutation__round__N2927 ) );
  AND2_X2 _f_permutation__round__U1416  ( .A1(_f_permutation__round__n810 ), 
        .A2(_f_permutation__round__c[1593] ), .ZN(
        _f_permutation__round__N2929 ) );
  AND2_X2 _f_permutation__round__U1415  ( .A1(_f_permutation__round__n813 ), 
        .A2(_f_permutation__round__c[1592] ), .ZN(
        _f_permutation__round__N2931 ) );
  AND2_X2 _f_permutation__round__U1414  ( .A1(_f_permutation__round__n816 ), 
        .A2(_f_permutation__round__c[1591] ), .ZN(
        _f_permutation__round__N2933 ) );
  AND2_X2 _f_permutation__round__U1413  ( .A1(_f_permutation__round__n819 ), 
        .A2(_f_permutation__round__c[1590] ), .ZN(
        _f_permutation__round__N2935 ) );
  AND2_X2 _f_permutation__round__U1412  ( .A1(_f_permutation__round__n822 ), 
        .A2(_f_permutation__round__c[1589] ), .ZN(
        _f_permutation__round__N2937 ) );
  AND2_X2 _f_permutation__round__U1411  ( .A1(_f_permutation__round__n825 ), 
        .A2(_f_permutation__round__c[1588] ), .ZN(
        _f_permutation__round__N2939 ) );
  AND2_X2 _f_permutation__round__U1410  ( .A1(_f_permutation__round__n828 ), 
        .A2(_f_permutation__round__c[1587] ), .ZN(
        _f_permutation__round__N2941 ) );
  AND2_X2 _f_permutation__round__U1409  ( .A1(_f_permutation__round__n831 ), 
        .A2(_f_permutation__round__c[1586] ), .ZN(
        _f_permutation__round__N2943 ) );
  AND2_X2 _f_permutation__round__U1344  ( .A1(_f_permutation__round__n7 ), 
        .A2(_f_permutation__round__c[403] ), .ZN(_f_permutation__round__N3073 ) );
  AND2_X2 _f_permutation__round__U1343  ( .A1(_f_permutation__round__n14 ), 
        .A2(_f_permutation__round__c[402] ), .ZN(_f_permutation__round__N3075 ) );
  AND2_X2 _f_permutation__round__U1342  ( .A1(_f_permutation__round__n21 ), 
        .A2(_f_permutation__round__c[401] ), .ZN(_f_permutation__round__N3077 ) );
  AND2_X2 _f_permutation__round__U1341  ( .A1(_f_permutation__round__n28 ), 
        .A2(_f_permutation__round__c[400] ), .ZN(_f_permutation__round__N3079 ) );
  AND2_X2 _f_permutation__round__U1340  ( .A1(_f_permutation__round__n35 ), 
        .A2(_f_permutation__round__c[399] ), .ZN(_f_permutation__round__N3081 ) );
  AND2_X2 _f_permutation__round__U1339  ( .A1(_f_permutation__round__n42 ), 
        .A2(_f_permutation__round__c[398] ), .ZN(_f_permutation__round__N3083 ) );
  AND2_X2 _f_permutation__round__U1338  ( .A1(_f_permutation__round__n49 ), 
        .A2(_f_permutation__round__c[397] ), .ZN(_f_permutation__round__N3085 ) );
  AND2_X2 _f_permutation__round__U1337  ( .A1(_f_permutation__round__n56 ), 
        .A2(_f_permutation__round__c[396] ), .ZN(_f_permutation__round__N3087 ) );
  AND2_X2 _f_permutation__round__U1336  ( .A1(_f_permutation__round__n63 ), 
        .A2(_f_permutation__round__c[395] ), .ZN(_f_permutation__round__N3089 ) );
  AND2_X2 _f_permutation__round__U1335  ( .A1(_f_permutation__round__n70 ), 
        .A2(_f_permutation__round__c[394] ), .ZN(_f_permutation__round__N3091 ) );
  AND2_X2 _f_permutation__round__U1334  ( .A1(_f_permutation__round__n77 ), 
        .A2(_f_permutation__round__c[393] ), .ZN(_f_permutation__round__N3093 ) );
  AND2_X2 _f_permutation__round__U1333  ( .A1(_f_permutation__round__n84 ), 
        .A2(_f_permutation__round__c[392] ), .ZN(_f_permutation__round__N3095 ) );
  AND2_X2 _f_permutation__round__U1332  ( .A1(_f_permutation__round__n91 ), 
        .A2(_f_permutation__round__c[391] ), .ZN(_f_permutation__round__N3097 ) );
  AND2_X2 _f_permutation__round__U1331  ( .A1(_f_permutation__round__n98 ), 
        .A2(_f_permutation__round__c[390] ), .ZN(_f_permutation__round__N3099 ) );
  AND2_X2 _f_permutation__round__U1330  ( .A1(_f_permutation__round__n105 ), 
        .A2(_f_permutation__round__c[389] ), .ZN(_f_permutation__round__N3101 ) );
  AND2_X2 _f_permutation__round__U1329  ( .A1(_f_permutation__round__n112 ), 
        .A2(_f_permutation__round__c[388] ), .ZN(_f_permutation__round__N3103 ) );
  AND2_X2 _f_permutation__round__U1328  ( .A1(_f_permutation__round__n119 ), 
        .A2(_f_permutation__round__c[387] ), .ZN(_f_permutation__round__N3105 ) );
  AND2_X2 _f_permutation__round__U1327  ( .A1(_f_permutation__round__n126 ), 
        .A2(_f_permutation__round__c[386] ), .ZN(_f_permutation__round__N3107 ) );
  AND2_X2 _f_permutation__round__U1326  ( .A1(_f_permutation__round__n133 ), 
        .A2(_f_permutation__round__c[385] ), .ZN(_f_permutation__round__N3109 ) );
  AND2_X2 _f_permutation__round__U1325  ( .A1(_f_permutation__round__n140 ), 
        .A2(_f_permutation__round__c[384] ), .ZN(_f_permutation__round__N3111 ) );
  AND2_X2 _f_permutation__round__U1324  ( .A1(_f_permutation__round__n147 ), 
        .A2(_f_permutation__round__c[447] ), .ZN(_f_permutation__round__N3113 ) );
  AND2_X2 _f_permutation__round__U1323  ( .A1(_f_permutation__round__n154 ), 
        .A2(_f_permutation__round__c[446] ), .ZN(_f_permutation__round__N3115 ) );
  AND2_X2 _f_permutation__round__U1322  ( .A1(_f_permutation__round__n161 ), 
        .A2(_f_permutation__round__c[445] ), .ZN(_f_permutation__round__N3117 ) );
  AND2_X2 _f_permutation__round__U1321  ( .A1(_f_permutation__round__n168 ), 
        .A2(_f_permutation__round__c[444] ), .ZN(_f_permutation__round__N3119 ) );
  AND2_X2 _f_permutation__round__U1320  ( .A1(_f_permutation__round__n175 ), 
        .A2(_f_permutation__round__c[443] ), .ZN(_f_permutation__round__N3121 ) );
  AND2_X2 _f_permutation__round__U1319  ( .A1(_f_permutation__round__n182 ), 
        .A2(_f_permutation__round__c[442] ), .ZN(_f_permutation__round__N3123 ) );
  AND2_X2 _f_permutation__round__U1318  ( .A1(_f_permutation__round__n189 ), 
        .A2(_f_permutation__round__c[441] ), .ZN(_f_permutation__round__N3125 ) );
  AND2_X2 _f_permutation__round__U1317  ( .A1(_f_permutation__round__n196 ), 
        .A2(_f_permutation__round__c[440] ), .ZN(_f_permutation__round__N3127 ) );
  AND2_X2 _f_permutation__round__U1316  ( .A1(_f_permutation__round__n203 ), 
        .A2(_f_permutation__round__c[439] ), .ZN(_f_permutation__round__N3129 ) );
  AND2_X2 _f_permutation__round__U1315  ( .A1(_f_permutation__round__n210 ), 
        .A2(_f_permutation__round__c[438] ), .ZN(_f_permutation__round__N3131 ) );
  AND2_X2 _f_permutation__round__U1314  ( .A1(_f_permutation__round__n217 ), 
        .A2(_f_permutation__round__c[437] ), .ZN(_f_permutation__round__N3133 ) );
  AND2_X2 _f_permutation__round__U1313  ( .A1(_f_permutation__round__n224 ), 
        .A2(_f_permutation__round__c[436] ), .ZN(_f_permutation__round__N3135 ) );
  AND2_X2 _f_permutation__round__U1312  ( .A1(_f_permutation__round__n231 ), 
        .A2(_f_permutation__round__c[435] ), .ZN(_f_permutation__round__N3137 ) );
  AND2_X2 _f_permutation__round__U1311  ( .A1(_f_permutation__round__n238 ), 
        .A2(_f_permutation__round__c[434] ), .ZN(_f_permutation__round__N3139 ) );
  AND2_X2 _f_permutation__round__U1310  ( .A1(_f_permutation__round__n245 ), 
        .A2(_f_permutation__round__c[433] ), .ZN(_f_permutation__round__N3141 ) );
  AND2_X2 _f_permutation__round__U1309  ( .A1(_f_permutation__round__n252 ), 
        .A2(_f_permutation__round__c[432] ), .ZN(_f_permutation__round__N3143 ) );
  AND2_X2 _f_permutation__round__U1308  ( .A1(_f_permutation__round__n259 ), 
        .A2(_f_permutation__round__c[431] ), .ZN(_f_permutation__round__N3145 ) );
  AND2_X2 _f_permutation__round__U1307  ( .A1(_f_permutation__round__n266 ), 
        .A2(_f_permutation__round__c[430] ), .ZN(_f_permutation__round__N3147 ) );
  AND2_X2 _f_permutation__round__U1306  ( .A1(_f_permutation__round__n273 ), 
        .A2(_f_permutation__round__c[429] ), .ZN(_f_permutation__round__N3149 ) );
  AND2_X2 _f_permutation__round__U1305  ( .A1(_f_permutation__round__n280 ), 
        .A2(_f_permutation__round__c[428] ), .ZN(_f_permutation__round__N3151 ) );
  AND2_X2 _f_permutation__round__U1304  ( .A1(_f_permutation__round__n287 ), 
        .A2(_f_permutation__round__c[427] ), .ZN(_f_permutation__round__N3153 ) );
  AND2_X2 _f_permutation__round__U1303  ( .A1(_f_permutation__round__n294 ), 
        .A2(_f_permutation__round__c[426] ), .ZN(_f_permutation__round__N3155 ) );
  AND2_X2 _f_permutation__round__U1302  ( .A1(_f_permutation__round__n301 ), 
        .A2(_f_permutation__round__c[425] ), .ZN(_f_permutation__round__N3157 ) );
  AND2_X2 _f_permutation__round__U1301  ( .A1(_f_permutation__round__n308 ), 
        .A2(_f_permutation__round__c[424] ), .ZN(_f_permutation__round__N3159 ) );
  AND2_X2 _f_permutation__round__U1300  ( .A1(_f_permutation__round__n315 ), 
        .A2(_f_permutation__round__c[423] ), .ZN(_f_permutation__round__N3161 ) );
  AND2_X2 _f_permutation__round__U1299  ( .A1(_f_permutation__round__n322 ), 
        .A2(_f_permutation__round__c[422] ), .ZN(_f_permutation__round__N3163 ) );
  AND2_X2 _f_permutation__round__U1298  ( .A1(_f_permutation__round__n329 ), 
        .A2(_f_permutation__round__c[421] ), .ZN(_f_permutation__round__N3165 ) );
  AND2_X2 _f_permutation__round__U1297  ( .A1(_f_permutation__round__n336 ), 
        .A2(_f_permutation__round__c[420] ), .ZN(_f_permutation__round__N3167 ) );
  AND2_X2 _f_permutation__round__U1296  ( .A1(_f_permutation__round__n343 ), 
        .A2(_f_permutation__round__c[419] ), .ZN(_f_permutation__round__N3169 ) );
  AND2_X2 _f_permutation__round__U1295  ( .A1(_f_permutation__round__n350 ), 
        .A2(_f_permutation__round__c[418] ), .ZN(_f_permutation__round__N3171 ) );
  AND2_X2 _f_permutation__round__U1294  ( .A1(_f_permutation__round__n357 ), 
        .A2(_f_permutation__round__c[417] ), .ZN(_f_permutation__round__N3173 ) );
  AND2_X2 _f_permutation__round__U1293  ( .A1(_f_permutation__round__n364 ), 
        .A2(_f_permutation__round__c[416] ), .ZN(_f_permutation__round__N3175 ) );
  AND2_X2 _f_permutation__round__U1292  ( .A1(_f_permutation__round__n371 ), 
        .A2(_f_permutation__round__c[415] ), .ZN(_f_permutation__round__N3177 ) );
  AND2_X2 _f_permutation__round__U1291  ( .A1(_f_permutation__round__n378 ), 
        .A2(_f_permutation__round__c[414] ), .ZN(_f_permutation__round__N3179 ) );
  AND2_X2 _f_permutation__round__U1290  ( .A1(_f_permutation__round__n385 ), 
        .A2(_f_permutation__round__c[413] ), .ZN(_f_permutation__round__N3181 ) );
  AND2_X2 _f_permutation__round__U1289  ( .A1(_f_permutation__round__n392 ), 
        .A2(_f_permutation__round__c[412] ), .ZN(_f_permutation__round__N3183 ) );
  AND2_X2 _f_permutation__round__U1288  ( .A1(_f_permutation__round__n399 ), 
        .A2(_f_permutation__round__c[411] ), .ZN(_f_permutation__round__N3185 ) );
  AND2_X2 _f_permutation__round__U1287  ( .A1(_f_permutation__round__n406 ), 
        .A2(_f_permutation__round__c[410] ), .ZN(_f_permutation__round__N3187 ) );
  AND2_X2 _f_permutation__round__U1286  ( .A1(_f_permutation__round__n413 ), 
        .A2(_f_permutation__round__c[409] ), .ZN(_f_permutation__round__N3189 ) );
  AND2_X2 _f_permutation__round__U1285  ( .A1(_f_permutation__round__n420 ), 
        .A2(_f_permutation__round__c[408] ), .ZN(_f_permutation__round__N3191 ) );
  AND2_X2 _f_permutation__round__U1284  ( .A1(_f_permutation__round__n427 ), 
        .A2(_f_permutation__round__c[407] ), .ZN(_f_permutation__round__N3193 ) );
  AND2_X2 _f_permutation__round__U1283  ( .A1(_f_permutation__round__n434 ), 
        .A2(_f_permutation__round__c[406] ), .ZN(_f_permutation__round__N3195 ) );
  AND2_X2 _f_permutation__round__U1282  ( .A1(_f_permutation__round__n441 ), 
        .A2(_f_permutation__round__c[405] ), .ZN(_f_permutation__round__N3197 ) );
  AND2_X2 _f_permutation__round__U1281  ( .A1(_f_permutation__round__n448 ), 
        .A2(_f_permutation__round__c[404] ), .ZN(_f_permutation__round__N3199 ) );
  AND2_X2 _f_permutation__round__U1152  ( .A1(_f_permutation__round__n318 ), 
        .A2(_f_permutation__round__c[898] ), .ZN(_f_permutation__round__N3457 ) );
  AND2_X2 _f_permutation__round__U1151  ( .A1(_f_permutation__round__n325 ), 
        .A2(_f_permutation__round__c[897] ), .ZN(_f_permutation__round__N3459 ) );
  AND2_X2 _f_permutation__round__U1150  ( .A1(_f_permutation__round__n332 ), 
        .A2(_f_permutation__round__c[896] ), .ZN(_f_permutation__round__N3461 ) );
  AND2_X2 _f_permutation__round__U1149  ( .A1(_f_permutation__round__n339 ), 
        .A2(_f_permutation__round__c[959] ), .ZN(_f_permutation__round__N3463 ) );
  AND2_X2 _f_permutation__round__U1148  ( .A1(_f_permutation__round__n346 ), 
        .A2(_f_permutation__round__c[958] ), .ZN(_f_permutation__round__N3465 ) );
  AND2_X2 _f_permutation__round__U1147  ( .A1(_f_permutation__round__n353 ), 
        .A2(_f_permutation__round__c[957] ), .ZN(_f_permutation__round__N3467 ) );
  AND2_X2 _f_permutation__round__U1146  ( .A1(_f_permutation__round__n360 ), 
        .A2(_f_permutation__round__c[956] ), .ZN(_f_permutation__round__N3469 ) );
  AND2_X2 _f_permutation__round__U1145  ( .A1(_f_permutation__round__n367 ), 
        .A2(_f_permutation__round__c[955] ), .ZN(_f_permutation__round__N3471 ) );
  AND2_X2 _f_permutation__round__U1144  ( .A1(_f_permutation__round__n374 ), 
        .A2(_f_permutation__round__c[954] ), .ZN(_f_permutation__round__N3473 ) );
  AND2_X2 _f_permutation__round__U1143  ( .A1(_f_permutation__round__n381 ), 
        .A2(_f_permutation__round__c[953] ), .ZN(_f_permutation__round__N3475 ) );
  AND2_X2 _f_permutation__round__U1142  ( .A1(_f_permutation__round__n388 ), 
        .A2(_f_permutation__round__c[952] ), .ZN(_f_permutation__round__N3477 ) );
  AND2_X2 _f_permutation__round__U1141  ( .A1(_f_permutation__round__n395 ), 
        .A2(_f_permutation__round__c[951] ), .ZN(_f_permutation__round__N3479 ) );
  AND2_X2 _f_permutation__round__U1140  ( .A1(_f_permutation__round__n402 ), 
        .A2(_f_permutation__round__c[950] ), .ZN(_f_permutation__round__N3481 ) );
  AND2_X2 _f_permutation__round__U1139  ( .A1(_f_permutation__round__n409 ), 
        .A2(_f_permutation__round__c[949] ), .ZN(_f_permutation__round__N3483 ) );
  AND2_X2 _f_permutation__round__U1138  ( .A1(_f_permutation__round__n416 ), 
        .A2(_f_permutation__round__c[948] ), .ZN(_f_permutation__round__N3485 ) );
  AND2_X2 _f_permutation__round__U1137  ( .A1(_f_permutation__round__n423 ), 
        .A2(_f_permutation__round__c[947] ), .ZN(_f_permutation__round__N3487 ) );
  AND2_X2 _f_permutation__round__U1136  ( .A1(_f_permutation__round__n430 ), 
        .A2(_f_permutation__round__c[946] ), .ZN(_f_permutation__round__N3489 ) );
  AND2_X2 _f_permutation__round__U1135  ( .A1(_f_permutation__round__n437 ), 
        .A2(_f_permutation__round__c[945] ), .ZN(_f_permutation__round__N3491 ) );
  AND2_X2 _f_permutation__round__U1134  ( .A1(_f_permutation__round__n444 ), 
        .A2(_f_permutation__round__c[944] ), .ZN(_f_permutation__round__N3493 ) );
  AND2_X2 _f_permutation__round__U1133  ( .A1(_f_permutation__round__n3 ), 
        .A2(_f_permutation__round__c[943] ), .ZN(_f_permutation__round__N3495 ) );
  AND2_X2 _f_permutation__round__U1132  ( .A1(_f_permutation__round__n10 ), 
        .A2(_f_permutation__round__c[942] ), .ZN(_f_permutation__round__N3497 ) );
  AND2_X2 _f_permutation__round__U1131  ( .A1(_f_permutation__round__n17 ), 
        .A2(_f_permutation__round__c[941] ), .ZN(_f_permutation__round__N3499 ) );
  AND2_X2 _f_permutation__round__U1130  ( .A1(_f_permutation__round__n24 ), 
        .A2(_f_permutation__round__c[940] ), .ZN(_f_permutation__round__N3501 ) );
  AND2_X2 _f_permutation__round__U1129  ( .A1(_f_permutation__round__n31 ), 
        .A2(_f_permutation__round__c[939] ), .ZN(_f_permutation__round__N3503 ) );
  AND2_X2 _f_permutation__round__U1128  ( .A1(_f_permutation__round__n38 ), 
        .A2(_f_permutation__round__c[938] ), .ZN(_f_permutation__round__N3505 ) );
  AND2_X2 _f_permutation__round__U1127  ( .A1(_f_permutation__round__n45 ), 
        .A2(_f_permutation__round__c[937] ), .ZN(_f_permutation__round__N3507 ) );
  AND2_X2 _f_permutation__round__U1126  ( .A1(_f_permutation__round__n52 ), 
        .A2(_f_permutation__round__c[936] ), .ZN(_f_permutation__round__N3509 ) );
  AND2_X2 _f_permutation__round__U1125  ( .A1(_f_permutation__round__n59 ), 
        .A2(_f_permutation__round__c[935] ), .ZN(_f_permutation__round__N3511 ) );
  AND2_X2 _f_permutation__round__U1124  ( .A1(_f_permutation__round__n66 ), 
        .A2(_f_permutation__round__c[934] ), .ZN(_f_permutation__round__N3513 ) );
  AND2_X2 _f_permutation__round__U1123  ( .A1(_f_permutation__round__n73 ), 
        .A2(_f_permutation__round__c[933] ), .ZN(_f_permutation__round__N3515 ) );
  AND2_X2 _f_permutation__round__U1122  ( .A1(_f_permutation__round__n80 ), 
        .A2(_f_permutation__round__c[932] ), .ZN(_f_permutation__round__N3517 ) );
  AND2_X2 _f_permutation__round__U1121  ( .A1(_f_permutation__round__n87 ), 
        .A2(_f_permutation__round__c[931] ), .ZN(_f_permutation__round__N3519 ) );
  AND2_X2 _f_permutation__round__U1120  ( .A1(_f_permutation__round__n94 ), 
        .A2(_f_permutation__round__c[930] ), .ZN(_f_permutation__round__N3521 ) );
  AND2_X2 _f_permutation__round__U1119  ( .A1(_f_permutation__round__n101 ), 
        .A2(_f_permutation__round__c[929] ), .ZN(_f_permutation__round__N3523 ) );
  AND2_X2 _f_permutation__round__U1118  ( .A1(_f_permutation__round__n108 ), 
        .A2(_f_permutation__round__c[928] ), .ZN(_f_permutation__round__N3525 ) );
  AND2_X2 _f_permutation__round__U1117  ( .A1(_f_permutation__round__n115 ), 
        .A2(_f_permutation__round__c[927] ), .ZN(_f_permutation__round__N3527 ) );
  AND2_X2 _f_permutation__round__U1116  ( .A1(_f_permutation__round__n122 ), 
        .A2(_f_permutation__round__c[926] ), .ZN(_f_permutation__round__N3529 ) );
  AND2_X2 _f_permutation__round__U1115  ( .A1(_f_permutation__round__n129 ), 
        .A2(_f_permutation__round__c[925] ), .ZN(_f_permutation__round__N3531 ) );
  AND2_X2 _f_permutation__round__U1114  ( .A1(_f_permutation__round__n136 ), 
        .A2(_f_permutation__round__c[924] ), .ZN(_f_permutation__round__N3533 ) );
  AND2_X2 _f_permutation__round__U1113  ( .A1(_f_permutation__round__n143 ), 
        .A2(_f_permutation__round__c[923] ), .ZN(_f_permutation__round__N3535 ) );
  AND2_X2 _f_permutation__round__U1112  ( .A1(_f_permutation__round__n150 ), 
        .A2(_f_permutation__round__c[922] ), .ZN(_f_permutation__round__N3537 ) );
  AND2_X2 _f_permutation__round__U1111  ( .A1(_f_permutation__round__n157 ), 
        .A2(_f_permutation__round__c[921] ), .ZN(_f_permutation__round__N3539 ) );
  AND2_X2 _f_permutation__round__U1110  ( .A1(_f_permutation__round__n164 ), 
        .A2(_f_permutation__round__c[920] ), .ZN(_f_permutation__round__N3541 ) );
  AND2_X2 _f_permutation__round__U1109  ( .A1(_f_permutation__round__n171 ), 
        .A2(_f_permutation__round__c[919] ), .ZN(_f_permutation__round__N3543 ) );
  AND2_X2 _f_permutation__round__U1108  ( .A1(_f_permutation__round__n178 ), 
        .A2(_f_permutation__round__c[918] ), .ZN(_f_permutation__round__N3545 ) );
  AND2_X2 _f_permutation__round__U1107  ( .A1(_f_permutation__round__n185 ), 
        .A2(_f_permutation__round__c[917] ), .ZN(_f_permutation__round__N3547 ) );
  AND2_X2 _f_permutation__round__U1106  ( .A1(_f_permutation__round__n192 ), 
        .A2(_f_permutation__round__c[916] ), .ZN(_f_permutation__round__N3549 ) );
  AND2_X2 _f_permutation__round__U1105  ( .A1(_f_permutation__round__n199 ), 
        .A2(_f_permutation__round__c[915] ), .ZN(_f_permutation__round__N3551 ) );
  AND2_X2 _f_permutation__round__U1104  ( .A1(_f_permutation__round__n206 ), 
        .A2(_f_permutation__round__c[914] ), .ZN(_f_permutation__round__N3553 ) );
  AND2_X2 _f_permutation__round__U1103  ( .A1(_f_permutation__round__n213 ), 
        .A2(_f_permutation__round__c[913] ), .ZN(_f_permutation__round__N3555 ) );
  AND2_X2 _f_permutation__round__U1102  ( .A1(_f_permutation__round__n220 ), 
        .A2(_f_permutation__round__c[912] ), .ZN(_f_permutation__round__N3557 ) );
  AND2_X2 _f_permutation__round__U1101  ( .A1(_f_permutation__round__n227 ), 
        .A2(_f_permutation__round__c[911] ), .ZN(_f_permutation__round__N3559 ) );
  AND2_X2 _f_permutation__round__U1100  ( .A1(_f_permutation__round__n234 ), 
        .A2(_f_permutation__round__c[910] ), .ZN(_f_permutation__round__N3561 ) );
  AND2_X2 _f_permutation__round__U1099  ( .A1(_f_permutation__round__n241 ), 
        .A2(_f_permutation__round__c[909] ), .ZN(_f_permutation__round__N3563 ) );
  AND2_X2 _f_permutation__round__U1098  ( .A1(_f_permutation__round__n248 ), 
        .A2(_f_permutation__round__c[908] ), .ZN(_f_permutation__round__N3565 ) );
  AND2_X2 _f_permutation__round__U1097  ( .A1(_f_permutation__round__n255 ), 
        .A2(_f_permutation__round__c[907] ), .ZN(_f_permutation__round__N3567 ) );
  AND2_X2 _f_permutation__round__U1096  ( .A1(_f_permutation__round__n262 ), 
        .A2(_f_permutation__round__c[906] ), .ZN(_f_permutation__round__N3569 ) );
  AND2_X2 _f_permutation__round__U1095  ( .A1(_f_permutation__round__n269 ), 
        .A2(_f_permutation__round__c[905] ), .ZN(_f_permutation__round__N3571 ) );
  AND2_X2 _f_permutation__round__U1094  ( .A1(_f_permutation__round__n276 ), 
        .A2(_f_permutation__round__c[904] ), .ZN(_f_permutation__round__N3573 ) );
  AND2_X2 _f_permutation__round__U1093  ( .A1(_f_permutation__round__n283 ), 
        .A2(_f_permutation__round__c[903] ), .ZN(_f_permutation__round__N3575 ) );
  AND2_X2 _f_permutation__round__U1092  ( .A1(_f_permutation__round__n290 ), 
        .A2(_f_permutation__round__c[902] ), .ZN(_f_permutation__round__N3577 ) );
  AND2_X2 _f_permutation__round__U1091  ( .A1(_f_permutation__round__n297 ), 
        .A2(_f_permutation__round__c[901] ), .ZN(_f_permutation__round__N3579 ) );
  AND2_X2 _f_permutation__round__U1090  ( .A1(_f_permutation__round__n304 ), 
        .A2(_f_permutation__round__c[900] ), .ZN(_f_permutation__round__N3581 ) );
  AND2_X2 _f_permutation__round__U1089  ( .A1(_f_permutation__round__n311 ), 
        .A2(_f_permutation__round__c[899] ), .ZN(_f_permutation__round__N3583 ) );
  AND2_X2 _f_permutation__round__U1024  ( .A1(_f_permutation__round__n853 ), 
        .A2(_f_permutation__round__c[1387] ), .ZN(
        _f_permutation__round__N3713 ) );
  AND2_X2 _f_permutation__round__U1023  ( .A1(_f_permutation__round__n856 ), 
        .A2(_f_permutation__round__c[1386] ), .ZN(
        _f_permutation__round__N3715 ) );
  AND2_X2 _f_permutation__round__U1022  ( .A1(_f_permutation__round__n859 ), 
        .A2(_f_permutation__round__c[1385] ), .ZN(
        _f_permutation__round__N3717 ) );
  AND2_X2 _f_permutation__round__U1021  ( .A1(_f_permutation__round__n862 ), 
        .A2(_f_permutation__round__c[1384] ), .ZN(
        _f_permutation__round__N3719 ) );
  AND2_X2 _f_permutation__round__U1020  ( .A1(_f_permutation__round__n865 ), 
        .A2(_f_permutation__round__c[1383] ), .ZN(
        _f_permutation__round__N3721 ) );
  AND2_X2 _f_permutation__round__U1019  ( .A1(_f_permutation__round__n868 ), 
        .A2(_f_permutation__round__c[1382] ), .ZN(
        _f_permutation__round__N3723 ) );
  AND2_X2 _f_permutation__round__U1018  ( .A1(_f_permutation__round__n871 ), 
        .A2(_f_permutation__round__c[1381] ), .ZN(
        _f_permutation__round__N3725 ) );
  AND2_X2 _f_permutation__round__U1017  ( .A1(_f_permutation__round__n874 ), 
        .A2(_f_permutation__round__c[1380] ), .ZN(
        _f_permutation__round__N3727 ) );
  AND2_X2 _f_permutation__round__U1016  ( .A1(_f_permutation__round__n877 ), 
        .A2(_f_permutation__round__c[1379] ), .ZN(
        _f_permutation__round__N3729 ) );
  AND2_X2 _f_permutation__round__U1015  ( .A1(_f_permutation__round__n880 ), 
        .A2(_f_permutation__round__c[1378] ), .ZN(
        _f_permutation__round__N3731 ) );
  AND2_X2 _f_permutation__round__U1014  ( .A1(_f_permutation__round__n883 ), 
        .A2(_f_permutation__round__c[1377] ), .ZN(
        _f_permutation__round__N3733 ) );
  AND2_X2 _f_permutation__round__U1013  ( .A1(_f_permutation__round__n886 ), 
        .A2(_f_permutation__round__c[1376] ), .ZN(
        _f_permutation__round__N3735 ) );
  AND2_X2 _f_permutation__round__U1012  ( .A1(_f_permutation__round__n889 ), 
        .A2(_f_permutation__round__c[1375] ), .ZN(
        _f_permutation__round__N3737 ) );
  AND2_X2 _f_permutation__round__U1011  ( .A1(_f_permutation__round__n892 ), 
        .A2(_f_permutation__round__c[1374] ), .ZN(
        _f_permutation__round__N3739 ) );
  AND2_X2 _f_permutation__round__U1010  ( .A1(_f_permutation__round__n895 ), 
        .A2(_f_permutation__round__c[1373] ), .ZN(
        _f_permutation__round__N3741 ) );
  AND2_X2 _f_permutation__round__U1009  ( .A1(_f_permutation__round__n898 ), 
        .A2(_f_permutation__round__c[1372] ), .ZN(
        _f_permutation__round__N3743 ) );
  AND2_X2 _f_permutation__round__U1008  ( .A1(_f_permutation__round__n901 ), 
        .A2(_f_permutation__round__c[1371] ), .ZN(
        _f_permutation__round__N3745 ) );
  AND2_X2 _f_permutation__round__U1007  ( .A1(_f_permutation__round__n904 ), 
        .A2(_f_permutation__round__c[1370] ), .ZN(
        _f_permutation__round__N3747 ) );
  AND2_X2 _f_permutation__round__U1006  ( .A1(_f_permutation__round__n907 ), 
        .A2(_f_permutation__round__c[1369] ), .ZN(
        _f_permutation__round__N3749 ) );
  AND2_X2 _f_permutation__round__U1005  ( .A1(_f_permutation__round__n910 ), 
        .A2(_f_permutation__round__c[1368] ), .ZN(
        _f_permutation__round__N3751 ) );
  AND2_X2 _f_permutation__round__U1004  ( .A1(_f_permutation__round__n913 ), 
        .A2(_f_permutation__round__c[1367] ), .ZN(
        _f_permutation__round__N3753 ) );
  AND2_X2 _f_permutation__round__U1003  ( .A1(_f_permutation__round__n916 ), 
        .A2(_f_permutation__round__c[1366] ), .ZN(
        _f_permutation__round__N3755 ) );
  AND2_X2 _f_permutation__round__U1002  ( .A1(_f_permutation__round__n919 ), 
        .A2(_f_permutation__round__c[1365] ), .ZN(
        _f_permutation__round__N3757 ) );
  AND2_X2 _f_permutation__round__U1001  ( .A1(_f_permutation__round__n922 ), 
        .A2(_f_permutation__round__c[1364] ), .ZN(
        _f_permutation__round__N3759 ) );
  AND2_X2 _f_permutation__round__U1000  ( .A1(_f_permutation__round__n925 ), 
        .A2(_f_permutation__round__c[1363] ), .ZN(
        _f_permutation__round__N3761 ) );
  AND2_X2 _f_permutation__round__U999  ( .A1(_f_permutation__round__n928 ), 
        .A2(_f_permutation__round__c[1362] ), .ZN(
        _f_permutation__round__N3763 ) );
  AND2_X2 _f_permutation__round__U998  ( .A1(_f_permutation__round__n931 ), 
        .A2(_f_permutation__round__c[1361] ), .ZN(
        _f_permutation__round__N3765 ) );
  AND2_X2 _f_permutation__round__U997  ( .A1(_f_permutation__round__n934 ), 
        .A2(_f_permutation__round__c[1360] ), .ZN(
        _f_permutation__round__N3767 ) );
  AND2_X2 _f_permutation__round__U996  ( .A1(_f_permutation__round__n937 ), 
        .A2(_f_permutation__round__c[1359] ), .ZN(
        _f_permutation__round__N3769 ) );
  AND2_X2 _f_permutation__round__U995  ( .A1(_f_permutation__round__n940 ), 
        .A2(_f_permutation__round__c[1358] ), .ZN(
        _f_permutation__round__N3771 ) );
  AND2_X2 _f_permutation__round__U994  ( .A1(_f_permutation__round__n943 ), 
        .A2(_f_permutation__round__c[1357] ), .ZN(
        _f_permutation__round__N3773 ) );
  AND2_X2 _f_permutation__round__U993  ( .A1(_f_permutation__round__n946 ), 
        .A2(_f_permutation__round__c[1356] ), .ZN(
        _f_permutation__round__N3775 ) );
  AND2_X2 _f_permutation__round__U992  ( .A1(_f_permutation__round__n949 ), 
        .A2(_f_permutation__round__c[1355] ), .ZN(
        _f_permutation__round__N3777 ) );
  AND2_X2 _f_permutation__round__U991  ( .A1(_f_permutation__round__n952 ), 
        .A2(_f_permutation__round__c[1354] ), .ZN(
        _f_permutation__round__N3779 ) );
  AND2_X2 _f_permutation__round__U990  ( .A1(_f_permutation__round__n955 ), 
        .A2(_f_permutation__round__c[1353] ), .ZN(
        _f_permutation__round__N3781 ) );
  AND2_X2 _f_permutation__round__U989  ( .A1(_f_permutation__round__n958 ), 
        .A2(_f_permutation__round__c[1352] ), .ZN(
        _f_permutation__round__N3783 ) );
  AND2_X2 _f_permutation__round__U988  ( .A1(_f_permutation__round__n769 ), 
        .A2(_f_permutation__round__c[1351] ), .ZN(
        _f_permutation__round__N3785 ) );
  AND2_X2 _f_permutation__round__U987  ( .A1(_f_permutation__round__n772 ), 
        .A2(_f_permutation__round__c[1350] ), .ZN(
        _f_permutation__round__N3787 ) );
  AND2_X2 _f_permutation__round__U986  ( .A1(_f_permutation__round__n775 ), 
        .A2(_f_permutation__round__c[1349] ), .ZN(
        _f_permutation__round__N3789 ) );
  AND2_X2 _f_permutation__round__U985  ( .A1(_f_permutation__round__n778 ), 
        .A2(_f_permutation__round__c[1348] ), .ZN(
        _f_permutation__round__N3791 ) );
  AND2_X2 _f_permutation__round__U984  ( .A1(_f_permutation__round__n781 ), 
        .A2(_f_permutation__round__c[1347] ), .ZN(
        _f_permutation__round__N3793 ) );
  AND2_X2 _f_permutation__round__U983  ( .A1(_f_permutation__round__n784 ), 
        .A2(_f_permutation__round__c[1346] ), .ZN(
        _f_permutation__round__N3795 ) );
  AND2_X2 _f_permutation__round__U982  ( .A1(_f_permutation__round__n787 ), 
        .A2(_f_permutation__round__c[1345] ), .ZN(
        _f_permutation__round__N3797 ) );
  AND2_X2 _f_permutation__round__U981  ( .A1(_f_permutation__round__n790 ), 
        .A2(_f_permutation__round__c[1344] ), .ZN(
        _f_permutation__round__N3799 ) );
  AND2_X2 _f_permutation__round__U980  ( .A1(_f_permutation__round__n793 ), 
        .A2(_f_permutation__round__c[1407] ), .ZN(
        _f_permutation__round__N3801 ) );
  AND2_X2 _f_permutation__round__U979  ( .A1(_f_permutation__round__n796 ), 
        .A2(_f_permutation__round__c[1406] ), .ZN(
        _f_permutation__round__N3803 ) );
  AND2_X2 _f_permutation__round__U978  ( .A1(_f_permutation__round__n799 ), 
        .A2(_f_permutation__round__c[1405] ), .ZN(
        _f_permutation__round__N3805 ) );
  AND2_X2 _f_permutation__round__U977  ( .A1(_f_permutation__round__n802 ), 
        .A2(_f_permutation__round__c[1404] ), .ZN(
        _f_permutation__round__N3807 ) );
  AND2_X2 _f_permutation__round__U976  ( .A1(_f_permutation__round__n805 ), 
        .A2(_f_permutation__round__c[1403] ), .ZN(
        _f_permutation__round__N3809 ) );
  AND2_X2 _f_permutation__round__U975  ( .A1(_f_permutation__round__n808 ), 
        .A2(_f_permutation__round__c[1402] ), .ZN(
        _f_permutation__round__N3811 ) );
  AND2_X2 _f_permutation__round__U974  ( .A1(_f_permutation__round__n811 ), 
        .A2(_f_permutation__round__c[1401] ), .ZN(
        _f_permutation__round__N3813 ) );
  AND2_X2 _f_permutation__round__U973  ( .A1(_f_permutation__round__n814 ), 
        .A2(_f_permutation__round__c[1400] ), .ZN(
        _f_permutation__round__N3815 ) );
  AND2_X2 _f_permutation__round__U972  ( .A1(_f_permutation__round__n817 ), 
        .A2(_f_permutation__round__c[1399] ), .ZN(
        _f_permutation__round__N3817 ) );
  AND2_X2 _f_permutation__round__U971  ( .A1(_f_permutation__round__n820 ), 
        .A2(_f_permutation__round__c[1398] ), .ZN(
        _f_permutation__round__N3819 ) );
  AND2_X2 _f_permutation__round__U970  ( .A1(_f_permutation__round__n823 ), 
        .A2(_f_permutation__round__c[1397] ), .ZN(
        _f_permutation__round__N3821 ) );
  AND2_X2 _f_permutation__round__U969  ( .A1(_f_permutation__round__n826 ), 
        .A2(_f_permutation__round__c[1396] ), .ZN(
        _f_permutation__round__N3823 ) );
  AND2_X2 _f_permutation__round__U968  ( .A1(_f_permutation__round__n829 ), 
        .A2(_f_permutation__round__c[1395] ), .ZN(
        _f_permutation__round__N3825 ) );
  AND2_X2 _f_permutation__round__U967  ( .A1(_f_permutation__round__n832 ), 
        .A2(_f_permutation__round__c[1394] ), .ZN(
        _f_permutation__round__N3827 ) );
  AND2_X2 _f_permutation__round__U966  ( .A1(_f_permutation__round__n835 ), 
        .A2(_f_permutation__round__c[1393] ), .ZN(
        _f_permutation__round__N3829 ) );
  AND2_X2 _f_permutation__round__U965  ( .A1(_f_permutation__round__n838 ), 
        .A2(_f_permutation__round__c[1392] ), .ZN(
        _f_permutation__round__N3831 ) );
  AND2_X2 _f_permutation__round__U964  ( .A1(_f_permutation__round__n841 ), 
        .A2(_f_permutation__round__c[1391] ), .ZN(
        _f_permutation__round__N3833 ) );
  AND2_X2 _f_permutation__round__U963  ( .A1(_f_permutation__round__n844 ), 
        .A2(_f_permutation__round__c[1390] ), .ZN(
        _f_permutation__round__N3835 ) );
  AND2_X2 _f_permutation__round__U962  ( .A1(_f_permutation__round__n847 ), 
        .A2(_f_permutation__round__c[1389] ), .ZN(
        _f_permutation__round__N3837 ) );
  AND2_X2 _f_permutation__round__U961  ( .A1(_f_permutation__round__n850 ), 
        .A2(_f_permutation__round__c[1388] ), .ZN(
        _f_permutation__round__N3839 ) );
  AND2_X2 _f_permutation__round__U832  ( .A1(_f_permutation__round__n69 ), 
        .A2(_f_permutation__round__c[301] ), .ZN(_f_permutation__round__N4097 ) );
  AND2_X2 _f_permutation__round__U831  ( .A1(_f_permutation__round__n76 ), 
        .A2(_f_permutation__round__c[300] ), .ZN(_f_permutation__round__N4099 ) );
  AND2_X2 _f_permutation__round__U830  ( .A1(_f_permutation__round__n83 ), 
        .A2(_f_permutation__round__c[299] ), .ZN(_f_permutation__round__N4101 ) );
  AND2_X2 _f_permutation__round__U829  ( .A1(_f_permutation__round__n90 ), 
        .A2(_f_permutation__round__c[298] ), .ZN(_f_permutation__round__N4103 ) );
  AND2_X2 _f_permutation__round__U828  ( .A1(_f_permutation__round__n97 ), 
        .A2(_f_permutation__round__c[297] ), .ZN(_f_permutation__round__N4105 ) );
  AND2_X2 _f_permutation__round__U827  ( .A1(_f_permutation__round__n104 ), 
        .A2(_f_permutation__round__c[296] ), .ZN(_f_permutation__round__N4107 ) );
  AND2_X2 _f_permutation__round__U826  ( .A1(_f_permutation__round__n111 ), 
        .A2(_f_permutation__round__c[295] ), .ZN(_f_permutation__round__N4109 ) );
  AND2_X2 _f_permutation__round__U825  ( .A1(_f_permutation__round__n118 ), 
        .A2(_f_permutation__round__c[294] ), .ZN(_f_permutation__round__N4111 ) );
  AND2_X2 _f_permutation__round__U824  ( .A1(_f_permutation__round__n125 ), 
        .A2(_f_permutation__round__c[293] ), .ZN(_f_permutation__round__N4113 ) );
  AND2_X2 _f_permutation__round__U823  ( .A1(_f_permutation__round__n132 ), 
        .A2(_f_permutation__round__c[292] ), .ZN(_f_permutation__round__N4115 ) );
  AND2_X2 _f_permutation__round__U822  ( .A1(_f_permutation__round__n139 ), 
        .A2(_f_permutation__round__c[291] ), .ZN(_f_permutation__round__N4117 ) );
  AND2_X2 _f_permutation__round__U821  ( .A1(_f_permutation__round__n146 ), 
        .A2(_f_permutation__round__c[290] ), .ZN(_f_permutation__round__N4119 ) );
  AND2_X2 _f_permutation__round__U820  ( .A1(_f_permutation__round__n153 ), 
        .A2(_f_permutation__round__c[289] ), .ZN(_f_permutation__round__N4121 ) );
  AND2_X2 _f_permutation__round__U819  ( .A1(_f_permutation__round__n160 ), 
        .A2(_f_permutation__round__c[288] ), .ZN(_f_permutation__round__N4123 ) );
  AND2_X2 _f_permutation__round__U818  ( .A1(_f_permutation__round__n167 ), 
        .A2(_f_permutation__round__c[287] ), .ZN(_f_permutation__round__N4125 ) );
  AND2_X2 _f_permutation__round__U817  ( .A1(_f_permutation__round__n174 ), 
        .A2(_f_permutation__round__c[286] ), .ZN(_f_permutation__round__N4127 ) );
  AND2_X2 _f_permutation__round__U816  ( .A1(_f_permutation__round__n181 ), 
        .A2(_f_permutation__round__c[285] ), .ZN(_f_permutation__round__N4129 ) );
  AND2_X2 _f_permutation__round__U815  ( .A1(_f_permutation__round__n188 ), 
        .A2(_f_permutation__round__c[284] ), .ZN(_f_permutation__round__N4131 ) );
  AND2_X2 _f_permutation__round__U814  ( .A1(_f_permutation__round__n195 ), 
        .A2(_f_permutation__round__c[283] ), .ZN(_f_permutation__round__N4133 ) );
  AND2_X2 _f_permutation__round__U813  ( .A1(_f_permutation__round__n202 ), 
        .A2(_f_permutation__round__c[282] ), .ZN(_f_permutation__round__N4135 ) );
  AND2_X2 _f_permutation__round__U812  ( .A1(_f_permutation__round__n209 ), 
        .A2(_f_permutation__round__c[281] ), .ZN(_f_permutation__round__N4137 ) );
  AND2_X2 _f_permutation__round__U811  ( .A1(_f_permutation__round__n216 ), 
        .A2(_f_permutation__round__c[280] ), .ZN(_f_permutation__round__N4139 ) );
  AND2_X2 _f_permutation__round__U810  ( .A1(_f_permutation__round__n223 ), 
        .A2(_f_permutation__round__c[279] ), .ZN(_f_permutation__round__N4141 ) );
  AND2_X2 _f_permutation__round__U809  ( .A1(_f_permutation__round__n230 ), 
        .A2(_f_permutation__round__c[278] ), .ZN(_f_permutation__round__N4143 ) );
  AND2_X2 _f_permutation__round__U808  ( .A1(_f_permutation__round__n237 ), 
        .A2(_f_permutation__round__c[277] ), .ZN(_f_permutation__round__N4145 ) );
  AND2_X2 _f_permutation__round__U807  ( .A1(_f_permutation__round__n244 ), 
        .A2(_f_permutation__round__c[276] ), .ZN(_f_permutation__round__N4147 ) );
  AND2_X2 _f_permutation__round__U806  ( .A1(_f_permutation__round__n251 ), 
        .A2(_f_permutation__round__c[275] ), .ZN(_f_permutation__round__N4149 ) );
  AND2_X2 _f_permutation__round__U805  ( .A1(_f_permutation__round__n258 ), 
        .A2(_f_permutation__round__c[274] ), .ZN(_f_permutation__round__N4151 ) );
  AND2_X2 _f_permutation__round__U804  ( .A1(_f_permutation__round__n265 ), 
        .A2(_f_permutation__round__c[273] ), .ZN(_f_permutation__round__N4153 ) );
  AND2_X2 _f_permutation__round__U803  ( .A1(_f_permutation__round__n272 ), 
        .A2(_f_permutation__round__c[272] ), .ZN(_f_permutation__round__N4155 ) );
  AND2_X2 _f_permutation__round__U802  ( .A1(_f_permutation__round__n279 ), 
        .A2(_f_permutation__round__c[271] ), .ZN(_f_permutation__round__N4157 ) );
  AND2_X2 _f_permutation__round__U801  ( .A1(_f_permutation__round__n286 ), 
        .A2(_f_permutation__round__c[270] ), .ZN(_f_permutation__round__N4159 ) );
  AND2_X2 _f_permutation__round__U800  ( .A1(_f_permutation__round__n293 ), 
        .A2(_f_permutation__round__c[269] ), .ZN(_f_permutation__round__N4161 ) );
  AND2_X2 _f_permutation__round__U799  ( .A1(_f_permutation__round__n300 ), 
        .A2(_f_permutation__round__c[268] ), .ZN(_f_permutation__round__N4163 ) );
  AND2_X2 _f_permutation__round__U798  ( .A1(_f_permutation__round__n307 ), 
        .A2(_f_permutation__round__c[267] ), .ZN(_f_permutation__round__N4165 ) );
  AND2_X2 _f_permutation__round__U797  ( .A1(_f_permutation__round__n314 ), 
        .A2(_f_permutation__round__c[266] ), .ZN(_f_permutation__round__N4167 ) );
  AND2_X2 _f_permutation__round__U796  ( .A1(_f_permutation__round__n321 ), 
        .A2(_f_permutation__round__c[265] ), .ZN(_f_permutation__round__N4169 ) );
  AND2_X2 _f_permutation__round__U795  ( .A1(_f_permutation__round__n328 ), 
        .A2(_f_permutation__round__c[264] ), .ZN(_f_permutation__round__N4171 ) );
  AND2_X2 _f_permutation__round__U794  ( .A1(_f_permutation__round__n335 ), 
        .A2(_f_permutation__round__c[263] ), .ZN(_f_permutation__round__N4173 ) );
  AND2_X2 _f_permutation__round__U793  ( .A1(_f_permutation__round__n342 ), 
        .A2(_f_permutation__round__c[262] ), .ZN(_f_permutation__round__N4175 ) );
  AND2_X2 _f_permutation__round__U792  ( .A1(_f_permutation__round__n349 ), 
        .A2(_f_permutation__round__c[261] ), .ZN(_f_permutation__round__N4177 ) );
  AND2_X2 _f_permutation__round__U791  ( .A1(_f_permutation__round__n356 ), 
        .A2(_f_permutation__round__c[260] ), .ZN(_f_permutation__round__N4179 ) );
  AND2_X2 _f_permutation__round__U790  ( .A1(_f_permutation__round__n363 ), 
        .A2(_f_permutation__round__c[259] ), .ZN(_f_permutation__round__N4181 ) );
  AND2_X2 _f_permutation__round__U789  ( .A1(_f_permutation__round__n370 ), 
        .A2(_f_permutation__round__c[258] ), .ZN(_f_permutation__round__N4183 ) );
  AND2_X2 _f_permutation__round__U788  ( .A1(_f_permutation__round__n377 ), 
        .A2(_f_permutation__round__c[257] ), .ZN(_f_permutation__round__N4185 ) );
  AND2_X2 _f_permutation__round__U787  ( .A1(_f_permutation__round__n384 ), 
        .A2(_f_permutation__round__c[256] ), .ZN(_f_permutation__round__N4187 ) );
  AND2_X2 _f_permutation__round__U786  ( .A1(_f_permutation__round__n391 ), 
        .A2(_f_permutation__round__c[319] ), .ZN(_f_permutation__round__N4189 ) );
  AND2_X2 _f_permutation__round__U785  ( .A1(_f_permutation__round__n398 ), 
        .A2(_f_permutation__round__c[318] ), .ZN(_f_permutation__round__N4191 ) );
  AND2_X2 _f_permutation__round__U784  ( .A1(_f_permutation__round__n405 ), 
        .A2(_f_permutation__round__c[317] ), .ZN(_f_permutation__round__N4193 ) );
  AND2_X2 _f_permutation__round__U783  ( .A1(_f_permutation__round__n412 ), 
        .A2(_f_permutation__round__c[316] ), .ZN(_f_permutation__round__N4195 ) );
  AND2_X2 _f_permutation__round__U782  ( .A1(_f_permutation__round__n419 ), 
        .A2(_f_permutation__round__c[315] ), .ZN(_f_permutation__round__N4197 ) );
  AND2_X2 _f_permutation__round__U781  ( .A1(_f_permutation__round__n426 ), 
        .A2(_f_permutation__round__c[314] ), .ZN(_f_permutation__round__N4199 ) );
  AND2_X2 _f_permutation__round__U780  ( .A1(_f_permutation__round__n433 ), 
        .A2(_f_permutation__round__c[313] ), .ZN(_f_permutation__round__N4201 ) );
  AND2_X2 _f_permutation__round__U779  ( .A1(_f_permutation__round__n440 ), 
        .A2(_f_permutation__round__c[312] ), .ZN(_f_permutation__round__N4203 ) );
  AND2_X2 _f_permutation__round__U778  ( .A1(_f_permutation__round__n447 ), 
        .A2(_f_permutation__round__c[311] ), .ZN(_f_permutation__round__N4205 ) );
  AND2_X2 _f_permutation__round__U777  ( .A1(_f_permutation__round__n6 ), .A2(
        _f_permutation__round__c[310] ), .ZN(_f_permutation__round__N4207 ) );
  AND2_X2 _f_permutation__round__U776  ( .A1(_f_permutation__round__n13 ), 
        .A2(_f_permutation__round__c[309] ), .ZN(_f_permutation__round__N4209 ) );
  AND2_X2 _f_permutation__round__U775  ( .A1(_f_permutation__round__n20 ), 
        .A2(_f_permutation__round__c[308] ), .ZN(_f_permutation__round__N4211 ) );
  AND2_X2 _f_permutation__round__U774  ( .A1(_f_permutation__round__n27 ), 
        .A2(_f_permutation__round__c[307] ), .ZN(_f_permutation__round__N4213 ) );
  AND2_X2 _f_permutation__round__U773  ( .A1(_f_permutation__round__n34 ), 
        .A2(_f_permutation__round__c[306] ), .ZN(_f_permutation__round__N4215 ) );
  AND2_X2 _f_permutation__round__U772  ( .A1(_f_permutation__round__n41 ), 
        .A2(_f_permutation__round__c[305] ), .ZN(_f_permutation__round__N4217 ) );
  AND2_X2 _f_permutation__round__U771  ( .A1(_f_permutation__round__n48 ), 
        .A2(_f_permutation__round__c[304] ), .ZN(_f_permutation__round__N4219 ) );
  AND2_X2 _f_permutation__round__U770  ( .A1(_f_permutation__round__n55 ), 
        .A2(_f_permutation__round__c[303] ), .ZN(_f_permutation__round__N4221 ) );
  AND2_X2 _f_permutation__round__U769  ( .A1(_f_permutation__round__n62 ), 
        .A2(_f_permutation__round__c[302] ), .ZN(_f_permutation__round__N4223 ) );
  AND2_X2 _f_permutation__round__U704  ( .A1(_f_permutation__round__n8 ), .A2(
        _f_permutation__round__c[761] ), .ZN(_f_permutation__round__N4353 ) );
  AND2_X2 _f_permutation__round__U703  ( .A1(_f_permutation__round__n15 ), 
        .A2(_f_permutation__round__c[760] ), .ZN(_f_permutation__round__N4355 ) );
  AND2_X2 _f_permutation__round__U702  ( .A1(_f_permutation__round__n22 ), 
        .A2(_f_permutation__round__c[759] ), .ZN(_f_permutation__round__N4357 ) );
  AND2_X2 _f_permutation__round__U701  ( .A1(_f_permutation__round__n29 ), 
        .A2(_f_permutation__round__c[758] ), .ZN(_f_permutation__round__N4359 ) );
  AND2_X2 _f_permutation__round__U700  ( .A1(_f_permutation__round__n36 ), 
        .A2(_f_permutation__round__c[757] ), .ZN(_f_permutation__round__N4361 ) );
  AND2_X2 _f_permutation__round__U699  ( .A1(_f_permutation__round__n43 ), 
        .A2(_f_permutation__round__c[756] ), .ZN(_f_permutation__round__N4363 ) );
  AND2_X2 _f_permutation__round__U698  ( .A1(_f_permutation__round__n50 ), 
        .A2(_f_permutation__round__c[755] ), .ZN(_f_permutation__round__N4365 ) );
  AND2_X2 _f_permutation__round__U697  ( .A1(_f_permutation__round__n57 ), 
        .A2(_f_permutation__round__c[754] ), .ZN(_f_permutation__round__N4367 ) );
  AND2_X2 _f_permutation__round__U696  ( .A1(_f_permutation__round__n64 ), 
        .A2(_f_permutation__round__c[753] ), .ZN(_f_permutation__round__N4369 ) );
  AND2_X2 _f_permutation__round__U695  ( .A1(_f_permutation__round__n71 ), 
        .A2(_f_permutation__round__c[752] ), .ZN(_f_permutation__round__N4371 ) );
  AND2_X2 _f_permutation__round__U694  ( .A1(_f_permutation__round__n78 ), 
        .A2(_f_permutation__round__c[751] ), .ZN(_f_permutation__round__N4373 ) );
  AND2_X2 _f_permutation__round__U693  ( .A1(_f_permutation__round__n85 ), 
        .A2(_f_permutation__round__c[750] ), .ZN(_f_permutation__round__N4375 ) );
  AND2_X2 _f_permutation__round__U692  ( .A1(_f_permutation__round__n92 ), 
        .A2(_f_permutation__round__c[749] ), .ZN(_f_permutation__round__N4377 ) );
  AND2_X2 _f_permutation__round__U691  ( .A1(_f_permutation__round__n99 ), 
        .A2(_f_permutation__round__c[748] ), .ZN(_f_permutation__round__N4379 ) );
  AND2_X2 _f_permutation__round__U690  ( .A1(_f_permutation__round__n106 ), 
        .A2(_f_permutation__round__c[747] ), .ZN(_f_permutation__round__N4381 ) );
  AND2_X2 _f_permutation__round__U689  ( .A1(_f_permutation__round__n113 ), 
        .A2(_f_permutation__round__c[746] ), .ZN(_f_permutation__round__N4383 ) );
  AND2_X2 _f_permutation__round__U688  ( .A1(_f_permutation__round__n120 ), 
        .A2(_f_permutation__round__c[745] ), .ZN(_f_permutation__round__N4385 ) );
  AND2_X2 _f_permutation__round__U687  ( .A1(_f_permutation__round__n127 ), 
        .A2(_f_permutation__round__c[744] ), .ZN(_f_permutation__round__N4387 ) );
  AND2_X2 _f_permutation__round__U686  ( .A1(_f_permutation__round__n134 ), 
        .A2(_f_permutation__round__c[743] ), .ZN(_f_permutation__round__N4389 ) );
  AND2_X2 _f_permutation__round__U685  ( .A1(_f_permutation__round__n141 ), 
        .A2(_f_permutation__round__c[742] ), .ZN(_f_permutation__round__N4391 ) );
  AND2_X2 _f_permutation__round__U684  ( .A1(_f_permutation__round__n148 ), 
        .A2(_f_permutation__round__c[741] ), .ZN(_f_permutation__round__N4393 ) );
  AND2_X2 _f_permutation__round__U683  ( .A1(_f_permutation__round__n155 ), 
        .A2(_f_permutation__round__c[740] ), .ZN(_f_permutation__round__N4395 ) );
  AND2_X2 _f_permutation__round__U682  ( .A1(_f_permutation__round__n162 ), 
        .A2(_f_permutation__round__c[739] ), .ZN(_f_permutation__round__N4397 ) );
  AND2_X2 _f_permutation__round__U681  ( .A1(_f_permutation__round__n169 ), 
        .A2(_f_permutation__round__c[738] ), .ZN(_f_permutation__round__N4399 ) );
  AND2_X2 _f_permutation__round__U680  ( .A1(_f_permutation__round__n176 ), 
        .A2(_f_permutation__round__c[737] ), .ZN(_f_permutation__round__N4401 ) );
  AND2_X2 _f_permutation__round__U679  ( .A1(_f_permutation__round__n183 ), 
        .A2(_f_permutation__round__c[736] ), .ZN(_f_permutation__round__N4403 ) );
  AND2_X2 _f_permutation__round__U678  ( .A1(_f_permutation__round__n190 ), 
        .A2(_f_permutation__round__c[735] ), .ZN(_f_permutation__round__N4405 ) );
  AND2_X2 _f_permutation__round__U677  ( .A1(_f_permutation__round__n197 ), 
        .A2(_f_permutation__round__c[734] ), .ZN(_f_permutation__round__N4407 ) );
  AND2_X2 _f_permutation__round__U676  ( .A1(_f_permutation__round__n204 ), 
        .A2(_f_permutation__round__c[733] ), .ZN(_f_permutation__round__N4409 ) );
  AND2_X2 _f_permutation__round__U675  ( .A1(_f_permutation__round__n211 ), 
        .A2(_f_permutation__round__c[732] ), .ZN(_f_permutation__round__N4411 ) );
  AND2_X2 _f_permutation__round__U674  ( .A1(_f_permutation__round__n218 ), 
        .A2(_f_permutation__round__c[731] ), .ZN(_f_permutation__round__N4413 ) );
  AND2_X2 _f_permutation__round__U673  ( .A1(_f_permutation__round__n225 ), 
        .A2(_f_permutation__round__c[730] ), .ZN(_f_permutation__round__N4415 ) );
  AND2_X2 _f_permutation__round__U672  ( .A1(_f_permutation__round__n232 ), 
        .A2(_f_permutation__round__c[729] ), .ZN(_f_permutation__round__N4417 ) );
  AND2_X2 _f_permutation__round__U671  ( .A1(_f_permutation__round__n239 ), 
        .A2(_f_permutation__round__c[728] ), .ZN(_f_permutation__round__N4419 ) );
  AND2_X2 _f_permutation__round__U670  ( .A1(_f_permutation__round__n246 ), 
        .A2(_f_permutation__round__c[727] ), .ZN(_f_permutation__round__N4421 ) );
  AND2_X2 _f_permutation__round__U669  ( .A1(_f_permutation__round__n253 ), 
        .A2(_f_permutation__round__c[726] ), .ZN(_f_permutation__round__N4423 ) );
  AND2_X2 _f_permutation__round__U668  ( .A1(_f_permutation__round__n260 ), 
        .A2(_f_permutation__round__c[725] ), .ZN(_f_permutation__round__N4425 ) );
  AND2_X2 _f_permutation__round__U667  ( .A1(_f_permutation__round__n267 ), 
        .A2(_f_permutation__round__c[724] ), .ZN(_f_permutation__round__N4427 ) );
  AND2_X2 _f_permutation__round__U666  ( .A1(_f_permutation__round__n274 ), 
        .A2(_f_permutation__round__c[723] ), .ZN(_f_permutation__round__N4429 ) );
  AND2_X2 _f_permutation__round__U665  ( .A1(_f_permutation__round__n281 ), 
        .A2(_f_permutation__round__c[722] ), .ZN(_f_permutation__round__N4431 ) );
  AND2_X2 _f_permutation__round__U664  ( .A1(_f_permutation__round__n288 ), 
        .A2(_f_permutation__round__c[721] ), .ZN(_f_permutation__round__N4433 ) );
  AND2_X2 _f_permutation__round__U663  ( .A1(_f_permutation__round__n295 ), 
        .A2(_f_permutation__round__c[720] ), .ZN(_f_permutation__round__N4435 ) );
  AND2_X2 _f_permutation__round__U662  ( .A1(_f_permutation__round__n302 ), 
        .A2(_f_permutation__round__c[719] ), .ZN(_f_permutation__round__N4437 ) );
  AND2_X2 _f_permutation__round__U661  ( .A1(_f_permutation__round__n309 ), 
        .A2(_f_permutation__round__c[718] ), .ZN(_f_permutation__round__N4439 ) );
  AND2_X2 _f_permutation__round__U660  ( .A1(_f_permutation__round__n316 ), 
        .A2(_f_permutation__round__c[717] ), .ZN(_f_permutation__round__N4441 ) );
  AND2_X2 _f_permutation__round__U659  ( .A1(_f_permutation__round__n323 ), 
        .A2(_f_permutation__round__c[716] ), .ZN(_f_permutation__round__N4443 ) );
  AND2_X2 _f_permutation__round__U658  ( .A1(_f_permutation__round__n330 ), 
        .A2(_f_permutation__round__c[715] ), .ZN(_f_permutation__round__N4445 ) );
  AND2_X2 _f_permutation__round__U657  ( .A1(_f_permutation__round__n337 ), 
        .A2(_f_permutation__round__c[714] ), .ZN(_f_permutation__round__N4447 ) );
  AND2_X2 _f_permutation__round__U656  ( .A1(_f_permutation__round__n344 ), 
        .A2(_f_permutation__round__c[713] ), .ZN(_f_permutation__round__N4449 ) );
  AND2_X2 _f_permutation__round__U655  ( .A1(_f_permutation__round__n351 ), 
        .A2(_f_permutation__round__c[712] ), .ZN(_f_permutation__round__N4451 ) );
  AND2_X2 _f_permutation__round__U654  ( .A1(_f_permutation__round__n358 ), 
        .A2(_f_permutation__round__c[711] ), .ZN(_f_permutation__round__N4453 ) );
  AND2_X2 _f_permutation__round__U653  ( .A1(_f_permutation__round__n365 ), 
        .A2(_f_permutation__round__c[710] ), .ZN(_f_permutation__round__N4455 ) );
  AND2_X2 _f_permutation__round__U652  ( .A1(_f_permutation__round__n372 ), 
        .A2(_f_permutation__round__c[709] ), .ZN(_f_permutation__round__N4457 ) );
  AND2_X2 _f_permutation__round__U651  ( .A1(_f_permutation__round__n379 ), 
        .A2(_f_permutation__round__c[708] ), .ZN(_f_permutation__round__N4459 ) );
  AND2_X2 _f_permutation__round__U650  ( .A1(_f_permutation__round__n386 ), 
        .A2(_f_permutation__round__c[707] ), .ZN(_f_permutation__round__N4461 ) );
  AND2_X2 _f_permutation__round__U649  ( .A1(_f_permutation__round__n393 ), 
        .A2(_f_permutation__round__c[706] ), .ZN(_f_permutation__round__N4463 ) );
  AND2_X2 _f_permutation__round__U648  ( .A1(_f_permutation__round__n400 ), 
        .A2(_f_permutation__round__c[705] ), .ZN(_f_permutation__round__N4465 ) );
  AND2_X2 _f_permutation__round__U647  ( .A1(_f_permutation__round__n407 ), 
        .A2(_f_permutation__round__c[704] ), .ZN(_f_permutation__round__N4467 ) );
  AND2_X2 _f_permutation__round__U646  ( .A1(_f_permutation__round__n414 ), 
        .A2(_f_permutation__round__c[767] ), .ZN(_f_permutation__round__N4469 ) );
  AND2_X2 _f_permutation__round__U645  ( .A1(_f_permutation__round__n421 ), 
        .A2(_f_permutation__round__c[766] ), .ZN(_f_permutation__round__N4471 ) );
  AND2_X2 _f_permutation__round__U644  ( .A1(_f_permutation__round__n428 ), 
        .A2(_f_permutation__round__c[765] ), .ZN(_f_permutation__round__N4473 ) );
  AND2_X2 _f_permutation__round__U643  ( .A1(_f_permutation__round__n435 ), 
        .A2(_f_permutation__round__c[764] ), .ZN(_f_permutation__round__N4475 ) );
  AND2_X2 _f_permutation__round__U642  ( .A1(_f_permutation__round__n442 ), 
        .A2(_f_permutation__round__c[763] ), .ZN(_f_permutation__round__N4477 ) );
  AND2_X2 _f_permutation__round__U641  ( .A1(_f_permutation__round__n1 ), .A2(
        _f_permutation__round__c[762] ), .ZN(_f_permutation__round__N4479 ) );
  AND2_X2 _f_permutation__round__U512  ( .A1(_f_permutation__round__n526 ), 
        .A2(_f_permutation__round__c[1223] ), .ZN(
        _f_permutation__round__N4737 ) );
  AND2_X2 _f_permutation__round__U511  ( .A1(_f_permutation__round__n531 ), 
        .A2(_f_permutation__round__c[1222] ), .ZN(
        _f_permutation__round__N4739 ) );
  AND2_X2 _f_permutation__round__U510  ( .A1(_f_permutation__round__n536 ), 
        .A2(_f_permutation__round__c[1221] ), .ZN(
        _f_permutation__round__N4741 ) );
  AND2_X2 _f_permutation__round__U509  ( .A1(_f_permutation__round__n541 ), 
        .A2(_f_permutation__round__c[1220] ), .ZN(
        _f_permutation__round__N4743 ) );
  AND2_X2 _f_permutation__round__U508  ( .A1(_f_permutation__round__n546 ), 
        .A2(_f_permutation__round__c[1219] ), .ZN(
        _f_permutation__round__N4745 ) );
  AND2_X2 _f_permutation__round__U507  ( .A1(_f_permutation__round__n551 ), 
        .A2(_f_permutation__round__c[1218] ), .ZN(
        _f_permutation__round__N4747 ) );
  AND2_X2 _f_permutation__round__U506  ( .A1(_f_permutation__round__n556 ), 
        .A2(_f_permutation__round__c[1217] ), .ZN(
        _f_permutation__round__N4749 ) );
  AND2_X2 _f_permutation__round__U505  ( .A1(_f_permutation__round__n561 ), 
        .A2(_f_permutation__round__c[1216] ), .ZN(
        _f_permutation__round__N4751 ) );
  AND2_X2 _f_permutation__round__U504  ( .A1(_f_permutation__round__n566 ), 
        .A2(_f_permutation__round__c[1279] ), .ZN(
        _f_permutation__round__N4753 ) );
  AND2_X2 _f_permutation__round__U503  ( .A1(_f_permutation__round__n571 ), 
        .A2(_f_permutation__round__c[1278] ), .ZN(
        _f_permutation__round__N4755 ) );
  AND2_X2 _f_permutation__round__U502  ( .A1(_f_permutation__round__n576 ), 
        .A2(_f_permutation__round__c[1277] ), .ZN(
        _f_permutation__round__N4757 ) );
  AND2_X2 _f_permutation__round__U501  ( .A1(_f_permutation__round__n581 ), 
        .A2(_f_permutation__round__c[1276] ), .ZN(
        _f_permutation__round__N4759 ) );
  AND2_X2 _f_permutation__round__U500  ( .A1(_f_permutation__round__n586 ), 
        .A2(_f_permutation__round__c[1275] ), .ZN(
        _f_permutation__round__N4761 ) );
  AND2_X2 _f_permutation__round__U499  ( .A1(_f_permutation__round__n591 ), 
        .A2(_f_permutation__round__c[1274] ), .ZN(
        _f_permutation__round__N4763 ) );
  AND2_X2 _f_permutation__round__U498  ( .A1(_f_permutation__round__n596 ), 
        .A2(_f_permutation__round__c[1273] ), .ZN(
        _f_permutation__round__N4765 ) );
  AND2_X2 _f_permutation__round__U497  ( .A1(_f_permutation__round__n601 ), 
        .A2(_f_permutation__round__c[1272] ), .ZN(
        _f_permutation__round__N4767 ) );
  AND2_X2 _f_permutation__round__U496  ( .A1(_f_permutation__round__n606 ), 
        .A2(_f_permutation__round__c[1271] ), .ZN(
        _f_permutation__round__N4769 ) );
  AND2_X2 _f_permutation__round__U495  ( .A1(_f_permutation__round__n611 ), 
        .A2(_f_permutation__round__c[1270] ), .ZN(
        _f_permutation__round__N4771 ) );
  AND2_X2 _f_permutation__round__U494  ( .A1(_f_permutation__round__n616 ), 
        .A2(_f_permutation__round__c[1269] ), .ZN(
        _f_permutation__round__N4773 ) );
  AND2_X2 _f_permutation__round__U493  ( .A1(_f_permutation__round__n621 ), 
        .A2(_f_permutation__round__c[1268] ), .ZN(
        _f_permutation__round__N4775 ) );
  AND2_X2 _f_permutation__round__U492  ( .A1(_f_permutation__round__n626 ), 
        .A2(_f_permutation__round__c[1267] ), .ZN(
        _f_permutation__round__N4777 ) );
  AND2_X2 _f_permutation__round__U491  ( .A1(_f_permutation__round__n631 ), 
        .A2(_f_permutation__round__c[1266] ), .ZN(
        _f_permutation__round__N4779 ) );
  AND2_X2 _f_permutation__round__U490  ( .A1(_f_permutation__round__n636 ), 
        .A2(_f_permutation__round__c[1265] ), .ZN(
        _f_permutation__round__N4781 ) );
  AND2_X2 _f_permutation__round__U489  ( .A1(_f_permutation__round__n641 ), 
        .A2(_f_permutation__round__c[1264] ), .ZN(
        _f_permutation__round__N4783 ) );
  AND2_X2 _f_permutation__round__U488  ( .A1(_f_permutation__round__n646 ), 
        .A2(_f_permutation__round__c[1263] ), .ZN(
        _f_permutation__round__N4785 ) );
  AND2_X2 _f_permutation__round__U487  ( .A1(_f_permutation__round__n651 ), 
        .A2(_f_permutation__round__c[1262] ), .ZN(
        _f_permutation__round__N4787 ) );
  AND2_X2 _f_permutation__round__U486  ( .A1(_f_permutation__round__n656 ), 
        .A2(_f_permutation__round__c[1261] ), .ZN(
        _f_permutation__round__N4789 ) );
  AND2_X2 _f_permutation__round__U485  ( .A1(_f_permutation__round__n661 ), 
        .A2(_f_permutation__round__c[1260] ), .ZN(
        _f_permutation__round__N4791 ) );
  AND2_X2 _f_permutation__round__U484  ( .A1(_f_permutation__round__n666 ), 
        .A2(_f_permutation__round__c[1259] ), .ZN(
        _f_permutation__round__N4793 ) );
  AND2_X2 _f_permutation__round__U483  ( .A1(_f_permutation__round__n671 ), 
        .A2(_f_permutation__round__c[1258] ), .ZN(
        _f_permutation__round__N4795 ) );
  AND2_X2 _f_permutation__round__U482  ( .A1(_f_permutation__round__n676 ), 
        .A2(_f_permutation__round__c[1257] ), .ZN(
        _f_permutation__round__N4797 ) );
  AND2_X2 _f_permutation__round__U481  ( .A1(_f_permutation__round__n681 ), 
        .A2(_f_permutation__round__c[1256] ), .ZN(
        _f_permutation__round__N4799 ) );
  AND2_X2 _f_permutation__round__U480  ( .A1(_f_permutation__round__n686 ), 
        .A2(_f_permutation__round__c[1255] ), .ZN(
        _f_permutation__round__N4801 ) );
  AND2_X2 _f_permutation__round__U479  ( .A1(_f_permutation__round__n691 ), 
        .A2(_f_permutation__round__c[1254] ), .ZN(
        _f_permutation__round__N4803 ) );
  AND2_X2 _f_permutation__round__U478  ( .A1(_f_permutation__round__n696 ), 
        .A2(_f_permutation__round__c[1253] ), .ZN(
        _f_permutation__round__N4805 ) );
  AND2_X2 _f_permutation__round__U477  ( .A1(_f_permutation__round__n701 ), 
        .A2(_f_permutation__round__c[1252] ), .ZN(
        _f_permutation__round__N4807 ) );
  AND2_X2 _f_permutation__round__U476  ( .A1(_f_permutation__round__n706 ), 
        .A2(_f_permutation__round__c[1251] ), .ZN(
        _f_permutation__round__N4809 ) );
  AND2_X2 _f_permutation__round__U475  ( .A1(_f_permutation__round__n711 ), 
        .A2(_f_permutation__round__c[1250] ), .ZN(
        _f_permutation__round__N4811 ) );
  AND2_X2 _f_permutation__round__U474  ( .A1(_f_permutation__round__n716 ), 
        .A2(_f_permutation__round__c[1249] ), .ZN(
        _f_permutation__round__N4813 ) );
  AND2_X2 _f_permutation__round__U473  ( .A1(_f_permutation__round__n721 ), 
        .A2(_f_permutation__round__c[1248] ), .ZN(
        _f_permutation__round__N4815 ) );
  AND2_X2 _f_permutation__round__U472  ( .A1(_f_permutation__round__n726 ), 
        .A2(_f_permutation__round__c[1247] ), .ZN(
        _f_permutation__round__N4817 ) );
  AND2_X2 _f_permutation__round__U471  ( .A1(_f_permutation__round__n731 ), 
        .A2(_f_permutation__round__c[1246] ), .ZN(
        _f_permutation__round__N4819 ) );
  AND2_X2 _f_permutation__round__U470  ( .A1(_f_permutation__round__n736 ), 
        .A2(_f_permutation__round__c[1245] ), .ZN(
        _f_permutation__round__N4821 ) );
  AND2_X2 _f_permutation__round__U469  ( .A1(_f_permutation__round__n741 ), 
        .A2(_f_permutation__round__c[1244] ), .ZN(
        _f_permutation__round__N4823 ) );
  AND2_X2 _f_permutation__round__U468  ( .A1(_f_permutation__round__n746 ), 
        .A2(_f_permutation__round__c[1243] ), .ZN(
        _f_permutation__round__N4825 ) );
  AND2_X2 _f_permutation__round__U467  ( .A1(_f_permutation__round__n751 ), 
        .A2(_f_permutation__round__c[1242] ), .ZN(
        _f_permutation__round__N4827 ) );
  AND2_X2 _f_permutation__round__U466  ( .A1(_f_permutation__round__n756 ), 
        .A2(_f_permutation__round__c[1241] ), .ZN(
        _f_permutation__round__N4829 ) );
  AND2_X2 _f_permutation__round__U465  ( .A1(_f_permutation__round__n761 ), 
        .A2(_f_permutation__round__c[1240] ), .ZN(
        _f_permutation__round__N4831 ) );
  AND2_X2 _f_permutation__round__U464  ( .A1(_f_permutation__round__n766 ), 
        .A2(_f_permutation__round__c[1239] ), .ZN(
        _f_permutation__round__N4833 ) );
  AND2_X2 _f_permutation__round__U463  ( .A1(_f_permutation__round__n451 ), 
        .A2(_f_permutation__round__c[1238] ), .ZN(
        _f_permutation__round__N4835 ) );
  AND2_X2 _f_permutation__round__U462  ( .A1(_f_permutation__round__n456 ), 
        .A2(_f_permutation__round__c[1237] ), .ZN(
        _f_permutation__round__N4837 ) );
  AND2_X2 _f_permutation__round__U461  ( .A1(_f_permutation__round__n461 ), 
        .A2(_f_permutation__round__c[1236] ), .ZN(
        _f_permutation__round__N4839 ) );
  AND2_X2 _f_permutation__round__U460  ( .A1(_f_permutation__round__n466 ), 
        .A2(_f_permutation__round__c[1235] ), .ZN(
        _f_permutation__round__N4841 ) );
  AND2_X2 _f_permutation__round__U459  ( .A1(_f_permutation__round__n471 ), 
        .A2(_f_permutation__round__c[1234] ), .ZN(
        _f_permutation__round__N4843 ) );
  AND2_X2 _f_permutation__round__U458  ( .A1(_f_permutation__round__n476 ), 
        .A2(_f_permutation__round__c[1233] ), .ZN(
        _f_permutation__round__N4845 ) );
  AND2_X2 _f_permutation__round__U457  ( .A1(_f_permutation__round__n481 ), 
        .A2(_f_permutation__round__c[1232] ), .ZN(
        _f_permutation__round__N4847 ) );
  AND2_X2 _f_permutation__round__U456  ( .A1(_f_permutation__round__n486 ), 
        .A2(_f_permutation__round__c[1231] ), .ZN(
        _f_permutation__round__N4849 ) );
  AND2_X2 _f_permutation__round__U455  ( .A1(_f_permutation__round__n491 ), 
        .A2(_f_permutation__round__c[1230] ), .ZN(
        _f_permutation__round__N4851 ) );
  AND2_X2 _f_permutation__round__U454  ( .A1(_f_permutation__round__n496 ), 
        .A2(_f_permutation__round__c[1229] ), .ZN(
        _f_permutation__round__N4853 ) );
  AND2_X2 _f_permutation__round__U453  ( .A1(_f_permutation__round__n501 ), 
        .A2(_f_permutation__round__c[1228] ), .ZN(
        _f_permutation__round__N4855 ) );
  AND2_X2 _f_permutation__round__U452  ( .A1(_f_permutation__round__n506 ), 
        .A2(_f_permutation__round__c[1227] ), .ZN(
        _f_permutation__round__N4857 ) );
  AND2_X2 _f_permutation__round__U451  ( .A1(_f_permutation__round__n511 ), 
        .A2(_f_permutation__round__c[1226] ), .ZN(
        _f_permutation__round__N4859 ) );
  AND2_X2 _f_permutation__round__U450  ( .A1(_f_permutation__round__n516 ), 
        .A2(_f_permutation__round__c[1225] ), .ZN(
        _f_permutation__round__N4861 ) );
  AND2_X2 _f_permutation__round__U449  ( .A1(_f_permutation__round__n521 ), 
        .A2(_f_permutation__round__c[1224] ), .ZN(
        _f_permutation__round__N4863 ) );
  AND2_X2 _f_permutation__round__U384  ( .A1(_f_permutation__round__n200 ), 
        .A2(_f_permutation__round__c[91] ), .ZN(_f_permutation__round__N4993 )
         );
  AND2_X2 _f_permutation__round__U383  ( .A1(_f_permutation__round__n207 ), 
        .A2(_f_permutation__round__c[90] ), .ZN(_f_permutation__round__N4995 )
         );
  AND2_X2 _f_permutation__round__U382  ( .A1(_f_permutation__round__n214 ), 
        .A2(_f_permutation__round__c[89] ), .ZN(_f_permutation__round__N4997 )
         );
  AND2_X2 _f_permutation__round__U381  ( .A1(_f_permutation__round__n221 ), 
        .A2(_f_permutation__round__c[88] ), .ZN(_f_permutation__round__N4999 )
         );
  AND2_X2 _f_permutation__round__U380  ( .A1(_f_permutation__round__n228 ), 
        .A2(_f_permutation__round__c[87] ), .ZN(_f_permutation__round__N5001 )
         );
  AND2_X2 _f_permutation__round__U379  ( .A1(_f_permutation__round__n235 ), 
        .A2(_f_permutation__round__c[86] ), .ZN(_f_permutation__round__N5003 )
         );
  AND2_X2 _f_permutation__round__U378  ( .A1(_f_permutation__round__n242 ), 
        .A2(_f_permutation__round__c[85] ), .ZN(_f_permutation__round__N5005 )
         );
  AND2_X2 _f_permutation__round__U377  ( .A1(_f_permutation__round__n249 ), 
        .A2(_f_permutation__round__c[84] ), .ZN(_f_permutation__round__N5007 )
         );
  AND2_X2 _f_permutation__round__U376  ( .A1(_f_permutation__round__n256 ), 
        .A2(_f_permutation__round__c[83] ), .ZN(_f_permutation__round__N5009 )
         );
  AND2_X2 _f_permutation__round__U375  ( .A1(_f_permutation__round__n263 ), 
        .A2(_f_permutation__round__c[82] ), .ZN(_f_permutation__round__N5011 )
         );
  AND2_X2 _f_permutation__round__U374  ( .A1(_f_permutation__round__n270 ), 
        .A2(_f_permutation__round__c[81] ), .ZN(_f_permutation__round__N5013 )
         );
  AND2_X2 _f_permutation__round__U373  ( .A1(_f_permutation__round__n277 ), 
        .A2(_f_permutation__round__c[80] ), .ZN(_f_permutation__round__N5015 )
         );
  AND2_X2 _f_permutation__round__U372  ( .A1(_f_permutation__round__n284 ), 
        .A2(_f_permutation__round__c[79] ), .ZN(_f_permutation__round__N5017 )
         );
  AND2_X2 _f_permutation__round__U371  ( .A1(_f_permutation__round__n291 ), 
        .A2(_f_permutation__round__c[78] ), .ZN(_f_permutation__round__N5019 )
         );
  AND2_X2 _f_permutation__round__U370  ( .A1(_f_permutation__round__n298 ), 
        .A2(_f_permutation__round__c[77] ), .ZN(_f_permutation__round__N5021 )
         );
  AND2_X2 _f_permutation__round__U369  ( .A1(_f_permutation__round__n305 ), 
        .A2(_f_permutation__round__c[76] ), .ZN(_f_permutation__round__N5023 )
         );
  AND2_X2 _f_permutation__round__U368  ( .A1(_f_permutation__round__n312 ), 
        .A2(_f_permutation__round__c[75] ), .ZN(_f_permutation__round__N5025 )
         );
  AND2_X2 _f_permutation__round__U367  ( .A1(_f_permutation__round__n319 ), 
        .A2(_f_permutation__round__c[74] ), .ZN(_f_permutation__round__N5027 )
         );
  AND2_X2 _f_permutation__round__U366  ( .A1(_f_permutation__round__n326 ), 
        .A2(_f_permutation__round__c[73] ), .ZN(_f_permutation__round__N5029 )
         );
  AND2_X2 _f_permutation__round__U365  ( .A1(_f_permutation__round__n333 ), 
        .A2(_f_permutation__round__c[72] ), .ZN(_f_permutation__round__N5031 )
         );
  AND2_X2 _f_permutation__round__U364  ( .A1(_f_permutation__round__n340 ), 
        .A2(_f_permutation__round__c[71] ), .ZN(_f_permutation__round__N5033 )
         );
  AND2_X2 _f_permutation__round__U363  ( .A1(_f_permutation__round__n347 ), 
        .A2(_f_permutation__round__c[70] ), .ZN(_f_permutation__round__N5035 )
         );
  AND2_X2 _f_permutation__round__U362  ( .A1(_f_permutation__round__n354 ), 
        .A2(_f_permutation__round__c[69] ), .ZN(_f_permutation__round__N5037 )
         );
  AND2_X2 _f_permutation__round__U361  ( .A1(_f_permutation__round__n361 ), 
        .A2(_f_permutation__round__c[68] ), .ZN(_f_permutation__round__N5039 )
         );
  AND2_X2 _f_permutation__round__U360  ( .A1(_f_permutation__round__n368 ), 
        .A2(_f_permutation__round__c[67] ), .ZN(_f_permutation__round__N5041 )
         );
  AND2_X2 _f_permutation__round__U359  ( .A1(_f_permutation__round__n375 ), 
        .A2(_f_permutation__round__c[66] ), .ZN(_f_permutation__round__N5043 )
         );
  AND2_X2 _f_permutation__round__U358  ( .A1(_f_permutation__round__n382 ), 
        .A2(_f_permutation__round__c[65] ), .ZN(_f_permutation__round__N5045 )
         );
  AND2_X2 _f_permutation__round__U357  ( .A1(_f_permutation__round__n389 ), 
        .A2(_f_permutation__round__c[64] ), .ZN(_f_permutation__round__N5047 )
         );
  AND2_X2 _f_permutation__round__U356  ( .A1(_f_permutation__round__n396 ), 
        .A2(_f_permutation__round__c[127] ), .ZN(_f_permutation__round__N5049 ) );
  AND2_X2 _f_permutation__round__U355  ( .A1(_f_permutation__round__n403 ), 
        .A2(_f_permutation__round__c[126] ), .ZN(_f_permutation__round__N5051 ) );
  AND2_X2 _f_permutation__round__U354  ( .A1(_f_permutation__round__n410 ), 
        .A2(_f_permutation__round__c[125] ), .ZN(_f_permutation__round__N5053 ) );
  AND2_X2 _f_permutation__round__U353  ( .A1(_f_permutation__round__n417 ), 
        .A2(_f_permutation__round__c[124] ), .ZN(_f_permutation__round__N5055 ) );
  AND2_X2 _f_permutation__round__U352  ( .A1(_f_permutation__round__n424 ), 
        .A2(_f_permutation__round__c[123] ), .ZN(_f_permutation__round__N5057 ) );
  AND2_X2 _f_permutation__round__U351  ( .A1(_f_permutation__round__n431 ), 
        .A2(_f_permutation__round__c[122] ), .ZN(_f_permutation__round__N5059 ) );
  AND2_X2 _f_permutation__round__U350  ( .A1(_f_permutation__round__n438 ), 
        .A2(_f_permutation__round__c[121] ), .ZN(_f_permutation__round__N5061 ) );
  AND2_X2 _f_permutation__round__U349  ( .A1(_f_permutation__round__n445 ), 
        .A2(_f_permutation__round__c[120] ), .ZN(_f_permutation__round__N5063 ) );
  AND2_X2 _f_permutation__round__U348  ( .A1(_f_permutation__round__n4 ), .A2(
        _f_permutation__round__c[119] ), .ZN(_f_permutation__round__N5065 ) );
  AND2_X2 _f_permutation__round__U347  ( .A1(_f_permutation__round__n11 ), 
        .A2(_f_permutation__round__c[118] ), .ZN(_f_permutation__round__N5067 ) );
  AND2_X2 _f_permutation__round__U346  ( .A1(_f_permutation__round__n18 ), 
        .A2(_f_permutation__round__c[117] ), .ZN(_f_permutation__round__N5069 ) );
  AND2_X2 _f_permutation__round__U345  ( .A1(_f_permutation__round__n25 ), 
        .A2(_f_permutation__round__c[116] ), .ZN(_f_permutation__round__N5071 ) );
  AND2_X2 _f_permutation__round__U344  ( .A1(_f_permutation__round__n32 ), 
        .A2(_f_permutation__round__c[115] ), .ZN(_f_permutation__round__N5073 ) );
  AND2_X2 _f_permutation__round__U343  ( .A1(_f_permutation__round__n39 ), 
        .A2(_f_permutation__round__c[114] ), .ZN(_f_permutation__round__N5075 ) );
  AND2_X2 _f_permutation__round__U342  ( .A1(_f_permutation__round__n46 ), 
        .A2(_f_permutation__round__c[113] ), .ZN(_f_permutation__round__N5077 ) );
  AND2_X2 _f_permutation__round__U341  ( .A1(_f_permutation__round__n53 ), 
        .A2(_f_permutation__round__c[112] ), .ZN(_f_permutation__round__N5079 ) );
  AND2_X2 _f_permutation__round__U340  ( .A1(_f_permutation__round__n60 ), 
        .A2(_f_permutation__round__c[111] ), .ZN(_f_permutation__round__N5081 ) );
  AND2_X2 _f_permutation__round__U339  ( .A1(_f_permutation__round__n67 ), 
        .A2(_f_permutation__round__c[110] ), .ZN(_f_permutation__round__N5083 ) );
  AND2_X2 _f_permutation__round__U338  ( .A1(_f_permutation__round__n74 ), 
        .A2(_f_permutation__round__c[109] ), .ZN(_f_permutation__round__N5085 ) );
  AND2_X2 _f_permutation__round__U337  ( .A1(_f_permutation__round__n81 ), 
        .A2(_f_permutation__round__c[108] ), .ZN(_f_permutation__round__N5087 ) );
  AND2_X2 _f_permutation__round__U336  ( .A1(_f_permutation__round__n88 ), 
        .A2(_f_permutation__round__c[107] ), .ZN(_f_permutation__round__N5089 ) );
  AND2_X2 _f_permutation__round__U335  ( .A1(_f_permutation__round__n95 ), 
        .A2(_f_permutation__round__c[106] ), .ZN(_f_permutation__round__N5091 ) );
  AND2_X2 _f_permutation__round__U334  ( .A1(_f_permutation__round__n102 ), 
        .A2(_f_permutation__round__c[105] ), .ZN(_f_permutation__round__N5093 ) );
  AND2_X2 _f_permutation__round__U333  ( .A1(_f_permutation__round__n109 ), 
        .A2(_f_permutation__round__c[104] ), .ZN(_f_permutation__round__N5095 ) );
  AND2_X2 _f_permutation__round__U332  ( .A1(_f_permutation__round__n116 ), 
        .A2(_f_permutation__round__c[103] ), .ZN(_f_permutation__round__N5097 ) );
  AND2_X2 _f_permutation__round__U331  ( .A1(_f_permutation__round__n123 ), 
        .A2(_f_permutation__round__c[102] ), .ZN(_f_permutation__round__N5099 ) );
  AND2_X2 _f_permutation__round__U330  ( .A1(_f_permutation__round__n130 ), 
        .A2(_f_permutation__round__c[101] ), .ZN(_f_permutation__round__N5101 ) );
  AND2_X2 _f_permutation__round__U329  ( .A1(_f_permutation__round__n137 ), 
        .A2(_f_permutation__round__c[100] ), .ZN(_f_permutation__round__N5103 ) );
  AND2_X2 _f_permutation__round__U328  ( .A1(_f_permutation__round__n144 ), 
        .A2(_f_permutation__round__c[99] ), .ZN(_f_permutation__round__N5105 )
         );
  AND2_X2 _f_permutation__round__U327  ( .A1(_f_permutation__round__n151 ), 
        .A2(_f_permutation__round__c[98] ), .ZN(_f_permutation__round__N5107 )
         );
  AND2_X2 _f_permutation__round__U326  ( .A1(_f_permutation__round__n158 ), 
        .A2(_f_permutation__round__c[97] ), .ZN(_f_permutation__round__N5109 )
         );
  AND2_X2 _f_permutation__round__U325  ( .A1(_f_permutation__round__n165 ), 
        .A2(_f_permutation__round__c[96] ), .ZN(_f_permutation__round__N5111 )
         );
  AND2_X2 _f_permutation__round__U324  ( .A1(_f_permutation__round__n172 ), 
        .A2(_f_permutation__round__c[95] ), .ZN(_f_permutation__round__N5113 )
         );
  AND2_X2 _f_permutation__round__U323  ( .A1(_f_permutation__round__n179 ), 
        .A2(_f_permutation__round__c[94] ), .ZN(_f_permutation__round__N5115 )
         );
  AND2_X2 _f_permutation__round__U322  ( .A1(_f_permutation__round__n186 ), 
        .A2(_f_permutation__round__c[93] ), .ZN(_f_permutation__round__N5117 )
         );
  AND2_X2 _f_permutation__round__U321  ( .A1(_f_permutation__round__n193 ), 
        .A2(_f_permutation__round__c[92] ), .ZN(_f_permutation__round__N5119 )
         );
  AND2_X2 _f_permutation__round__U192  ( .A1(_f_permutation__round__n663 ), 
        .A2(_f_permutation__round__c[637] ), .ZN(_f_permutation__round__N5377 ) );
  AND2_X2 _f_permutation__round__U191  ( .A1(_f_permutation__round__n668 ), 
        .A2(_f_permutation__round__c[636] ), .ZN(_f_permutation__round__N5379 ) );
  AND2_X2 _f_permutation__round__U190  ( .A1(_f_permutation__round__n673 ), 
        .A2(_f_permutation__round__c[635] ), .ZN(_f_permutation__round__N5381 ) );
  AND2_X2 _f_permutation__round__U189  ( .A1(_f_permutation__round__n678 ), 
        .A2(_f_permutation__round__c[634] ), .ZN(_f_permutation__round__N5383 ) );
  AND2_X2 _f_permutation__round__U188  ( .A1(_f_permutation__round__n683 ), 
        .A2(_f_permutation__round__c[633] ), .ZN(_f_permutation__round__N5385 ) );
  AND2_X2 _f_permutation__round__U187  ( .A1(_f_permutation__round__n688 ), 
        .A2(_f_permutation__round__c[632] ), .ZN(_f_permutation__round__N5387 ) );
  AND2_X2 _f_permutation__round__U186  ( .A1(_f_permutation__round__n693 ), 
        .A2(_f_permutation__round__c[631] ), .ZN(_f_permutation__round__N5389 ) );
  AND2_X2 _f_permutation__round__U185  ( .A1(_f_permutation__round__n698 ), 
        .A2(_f_permutation__round__c[630] ), .ZN(_f_permutation__round__N5391 ) );
  AND2_X2 _f_permutation__round__U184  ( .A1(_f_permutation__round__n703 ), 
        .A2(_f_permutation__round__c[629] ), .ZN(_f_permutation__round__N5393 ) );
  AND2_X2 _f_permutation__round__U183  ( .A1(_f_permutation__round__n708 ), 
        .A2(_f_permutation__round__c[628] ), .ZN(_f_permutation__round__N5395 ) );
  AND2_X2 _f_permutation__round__U182  ( .A1(_f_permutation__round__n713 ), 
        .A2(_f_permutation__round__c[627] ), .ZN(_f_permutation__round__N5397 ) );
  AND2_X2 _f_permutation__round__U181  ( .A1(_f_permutation__round__n718 ), 
        .A2(_f_permutation__round__c[626] ), .ZN(_f_permutation__round__N5399 ) );
  AND2_X2 _f_permutation__round__U180  ( .A1(_f_permutation__round__n723 ), 
        .A2(_f_permutation__round__c[625] ), .ZN(_f_permutation__round__N5401 ) );
  AND2_X2 _f_permutation__round__U179  ( .A1(_f_permutation__round__n728 ), 
        .A2(_f_permutation__round__c[624] ), .ZN(_f_permutation__round__N5403 ) );
  AND2_X2 _f_permutation__round__U178  ( .A1(_f_permutation__round__n733 ), 
        .A2(_f_permutation__round__c[623] ), .ZN(_f_permutation__round__N5405 ) );
  AND2_X2 _f_permutation__round__U177  ( .A1(_f_permutation__round__n738 ), 
        .A2(_f_permutation__round__c[622] ), .ZN(_f_permutation__round__N5407 ) );
  AND2_X2 _f_permutation__round__U176  ( .A1(_f_permutation__round__n743 ), 
        .A2(_f_permutation__round__c[621] ), .ZN(_f_permutation__round__N5409 ) );
  AND2_X2 _f_permutation__round__U175  ( .A1(_f_permutation__round__n748 ), 
        .A2(_f_permutation__round__c[620] ), .ZN(_f_permutation__round__N5411 ) );
  AND2_X2 _f_permutation__round__U174  ( .A1(_f_permutation__round__n753 ), 
        .A2(_f_permutation__round__c[619] ), .ZN(_f_permutation__round__N5413 ) );
  AND2_X2 _f_permutation__round__U173  ( .A1(_f_permutation__round__n758 ), 
        .A2(_f_permutation__round__c[618] ), .ZN(_f_permutation__round__N5415 ) );
  AND2_X2 _f_permutation__round__U172  ( .A1(_f_permutation__round__n763 ), 
        .A2(_f_permutation__round__c[617] ), .ZN(_f_permutation__round__N5417 ) );
  AND2_X2 _f_permutation__round__U171  ( .A1(_f_permutation__round__n768 ), 
        .A2(_f_permutation__round__c[616] ), .ZN(_f_permutation__round__N5419 ) );
  AND2_X2 _f_permutation__round__U170  ( .A1(_f_permutation__round__n453 ), 
        .A2(_f_permutation__round__c[615] ), .ZN(_f_permutation__round__N5421 ) );
  AND2_X2 _f_permutation__round__U169  ( .A1(_f_permutation__round__n458 ), 
        .A2(_f_permutation__round__c[614] ), .ZN(_f_permutation__round__N5423 ) );
  AND2_X2 _f_permutation__round__U168  ( .A1(_f_permutation__round__n463 ), 
        .A2(_f_permutation__round__c[613] ), .ZN(_f_permutation__round__N5425 ) );
  AND2_X2 _f_permutation__round__U167  ( .A1(_f_permutation__round__n468 ), 
        .A2(_f_permutation__round__c[612] ), .ZN(_f_permutation__round__N5427 ) );
  AND2_X2 _f_permutation__round__U166  ( .A1(_f_permutation__round__n473 ), 
        .A2(_f_permutation__round__c[611] ), .ZN(_f_permutation__round__N5429 ) );
  AND2_X2 _f_permutation__round__U165  ( .A1(_f_permutation__round__n478 ), 
        .A2(_f_permutation__round__c[610] ), .ZN(_f_permutation__round__N5431 ) );
  AND2_X2 _f_permutation__round__U164  ( .A1(_f_permutation__round__n483 ), 
        .A2(_f_permutation__round__c[609] ), .ZN(_f_permutation__round__N5433 ) );
  AND2_X2 _f_permutation__round__U163  ( .A1(_f_permutation__round__n488 ), 
        .A2(_f_permutation__round__c[608] ), .ZN(_f_permutation__round__N5435 ) );
  AND2_X2 _f_permutation__round__U162  ( .A1(_f_permutation__round__n493 ), 
        .A2(_f_permutation__round__c[607] ), .ZN(_f_permutation__round__N5437 ) );
  AND2_X2 _f_permutation__round__U161  ( .A1(_f_permutation__round__n498 ), 
        .A2(_f_permutation__round__c[606] ), .ZN(_f_permutation__round__N5439 ) );
  AND2_X2 _f_permutation__round__U160  ( .A1(_f_permutation__round__n503 ), 
        .A2(_f_permutation__round__c[605] ), .ZN(_f_permutation__round__N5441 ) );
  AND2_X2 _f_permutation__round__U159  ( .A1(_f_permutation__round__n508 ), 
        .A2(_f_permutation__round__c[604] ), .ZN(_f_permutation__round__N5443 ) );
  AND2_X2 _f_permutation__round__U158  ( .A1(_f_permutation__round__n513 ), 
        .A2(_f_permutation__round__c[603] ), .ZN(_f_permutation__round__N5445 ) );
  AND2_X2 _f_permutation__round__U157  ( .A1(_f_permutation__round__n518 ), 
        .A2(_f_permutation__round__c[602] ), .ZN(_f_permutation__round__N5447 ) );
  AND2_X2 _f_permutation__round__U156  ( .A1(_f_permutation__round__n523 ), 
        .A2(_f_permutation__round__c[601] ), .ZN(_f_permutation__round__N5449 ) );
  AND2_X2 _f_permutation__round__U155  ( .A1(_f_permutation__round__n528 ), 
        .A2(_f_permutation__round__c[600] ), .ZN(_f_permutation__round__N5451 ) );
  AND2_X2 _f_permutation__round__U154  ( .A1(_f_permutation__round__n533 ), 
        .A2(_f_permutation__round__c[599] ), .ZN(_f_permutation__round__N5453 ) );
  AND2_X2 _f_permutation__round__U153  ( .A1(_f_permutation__round__n538 ), 
        .A2(_f_permutation__round__c[598] ), .ZN(_f_permutation__round__N5455 ) );
  AND2_X2 _f_permutation__round__U152  ( .A1(_f_permutation__round__n543 ), 
        .A2(_f_permutation__round__c[597] ), .ZN(_f_permutation__round__N5457 ) );
  AND2_X2 _f_permutation__round__U151  ( .A1(_f_permutation__round__n548 ), 
        .A2(_f_permutation__round__c[596] ), .ZN(_f_permutation__round__N5459 ) );
  AND2_X2 _f_permutation__round__U150  ( .A1(_f_permutation__round__n553 ), 
        .A2(_f_permutation__round__c[595] ), .ZN(_f_permutation__round__N5461 ) );
  AND2_X2 _f_permutation__round__U149  ( .A1(_f_permutation__round__n558 ), 
        .A2(_f_permutation__round__c[594] ), .ZN(_f_permutation__round__N5463 ) );
  AND2_X2 _f_permutation__round__U148  ( .A1(_f_permutation__round__n563 ), 
        .A2(_f_permutation__round__c[593] ), .ZN(_f_permutation__round__N5465 ) );
  AND2_X2 _f_permutation__round__U147  ( .A1(_f_permutation__round__n568 ), 
        .A2(_f_permutation__round__c[592] ), .ZN(_f_permutation__round__N5467 ) );
  AND2_X2 _f_permutation__round__U146  ( .A1(_f_permutation__round__n573 ), 
        .A2(_f_permutation__round__c[591] ), .ZN(_f_permutation__round__N5469 ) );
  AND2_X2 _f_permutation__round__U145  ( .A1(_f_permutation__round__n578 ), 
        .A2(_f_permutation__round__c[590] ), .ZN(_f_permutation__round__N5471 ) );
  AND2_X2 _f_permutation__round__U144  ( .A1(_f_permutation__round__n583 ), 
        .A2(_f_permutation__round__c[589] ), .ZN(_f_permutation__round__N5473 ) );
  AND2_X2 _f_permutation__round__U143  ( .A1(_f_permutation__round__n588 ), 
        .A2(_f_permutation__round__c[588] ), .ZN(_f_permutation__round__N5475 ) );
  AND2_X2 _f_permutation__round__U142  ( .A1(_f_permutation__round__n593 ), 
        .A2(_f_permutation__round__c[587] ), .ZN(_f_permutation__round__N5477 ) );
  AND2_X2 _f_permutation__round__U141  ( .A1(_f_permutation__round__n598 ), 
        .A2(_f_permutation__round__c[586] ), .ZN(_f_permutation__round__N5479 ) );
  AND2_X2 _f_permutation__round__U140  ( .A1(_f_permutation__round__n603 ), 
        .A2(_f_permutation__round__c[585] ), .ZN(_f_permutation__round__N5481 ) );
  AND2_X2 _f_permutation__round__U139  ( .A1(_f_permutation__round__n608 ), 
        .A2(_f_permutation__round__c[584] ), .ZN(_f_permutation__round__N5483 ) );
  AND2_X2 _f_permutation__round__U138  ( .A1(_f_permutation__round__n613 ), 
        .A2(_f_permutation__round__c[583] ), .ZN(_f_permutation__round__N5485 ) );
  AND2_X2 _f_permutation__round__U137  ( .A1(_f_permutation__round__n618 ), 
        .A2(_f_permutation__round__c[582] ), .ZN(_f_permutation__round__N5487 ) );
  AND2_X2 _f_permutation__round__U136  ( .A1(_f_permutation__round__n623 ), 
        .A2(_f_permutation__round__c[581] ), .ZN(_f_permutation__round__N5489 ) );
  AND2_X2 _f_permutation__round__U135  ( .A1(_f_permutation__round__n628 ), 
        .A2(_f_permutation__round__c[580] ), .ZN(_f_permutation__round__N5491 ) );
  AND2_X2 _f_permutation__round__U134  ( .A1(_f_permutation__round__n633 ), 
        .A2(_f_permutation__round__c[579] ), .ZN(_f_permutation__round__N5493 ) );
  AND2_X2 _f_permutation__round__U133  ( .A1(_f_permutation__round__n638 ), 
        .A2(_f_permutation__round__c[578] ), .ZN(_f_permutation__round__N5495 ) );
  AND2_X2 _f_permutation__round__U132  ( .A1(_f_permutation__round__n643 ), 
        .A2(_f_permutation__round__c[577] ), .ZN(_f_permutation__round__N5497 ) );
  AND2_X2 _f_permutation__round__U131  ( .A1(_f_permutation__round__n648 ), 
        .A2(_f_permutation__round__c[576] ), .ZN(_f_permutation__round__N5499 ) );
  AND2_X2 _f_permutation__round__U130  ( .A1(_f_permutation__round__n653 ), 
        .A2(_f_permutation__round__c[639] ), .ZN(_f_permutation__round__N5501 ) );
  AND2_X2 _f_permutation__round__U129  ( .A1(_f_permutation__round__n658 ), 
        .A2(_f_permutation__round__c[638] ), .ZN(_f_permutation__round__N5503 ) );
  AND2_X2 _f_permutation__round__U64  ( .A1(_f_permutation__round__n759 ), 
        .A2(_f_permutation__round__c[1032] ), .ZN(
        _f_permutation__round__N5633 ) );
  AND2_X2 _f_permutation__round__U63  ( .A1(_f_permutation__round__n764 ), 
        .A2(_f_permutation__round__c[1031] ), .ZN(
        _f_permutation__round__N5635 ) );
  AND2_X2 _f_permutation__round__U62  ( .A1(_f_permutation__round__n449 ), 
        .A2(_f_permutation__round__c[1030] ), .ZN(
        _f_permutation__round__N5637 ) );
  AND2_X2 _f_permutation__round__U61  ( .A1(_f_permutation__round__n454 ), 
        .A2(_f_permutation__round__c[1029] ), .ZN(
        _f_permutation__round__N5639 ) );
  AND2_X2 _f_permutation__round__U60  ( .A1(_f_permutation__round__n459 ), 
        .A2(_f_permutation__round__c[1028] ), .ZN(
        _f_permutation__round__N5641 ) );
  AND2_X2 _f_permutation__round__U59  ( .A1(_f_permutation__round__n464 ), 
        .A2(_f_permutation__round__c[1027] ), .ZN(
        _f_permutation__round__N5643 ) );
  AND2_X2 _f_permutation__round__U58  ( .A1(_f_permutation__round__n469 ), 
        .A2(_f_permutation__round__c[1026] ), .ZN(
        _f_permutation__round__N5645 ) );
  AND2_X2 _f_permutation__round__U57  ( .A1(_f_permutation__round__n474 ), 
        .A2(_f_permutation__round__c[1025] ), .ZN(
        _f_permutation__round__N5647 ) );
  AND2_X2 _f_permutation__round__U56  ( .A1(_f_permutation__round__n479 ), 
        .A2(_f_permutation__round__c[1024] ), .ZN(
        _f_permutation__round__N5649 ) );
  AND2_X2 _f_permutation__round__U55  ( .A1(_f_permutation__round__n484 ), 
        .A2(_f_permutation__round__c[1087] ), .ZN(
        _f_permutation__round__N5651 ) );
  AND2_X2 _f_permutation__round__U54  ( .A1(_f_permutation__round__n489 ), 
        .A2(_f_permutation__round__c[1086] ), .ZN(
        _f_permutation__round__N5653 ) );
  AND2_X2 _f_permutation__round__U53  ( .A1(_f_permutation__round__n494 ), 
        .A2(_f_permutation__round__c[1085] ), .ZN(
        _f_permutation__round__N5655 ) );
  AND2_X2 _f_permutation__round__U52  ( .A1(_f_permutation__round__n499 ), 
        .A2(_f_permutation__round__c[1084] ), .ZN(
        _f_permutation__round__N5657 ) );
  AND2_X2 _f_permutation__round__U51  ( .A1(_f_permutation__round__n504 ), 
        .A2(_f_permutation__round__c[1083] ), .ZN(
        _f_permutation__round__N5659 ) );
  AND2_X2 _f_permutation__round__U50  ( .A1(_f_permutation__round__n509 ), 
        .A2(_f_permutation__round__c[1082] ), .ZN(
        _f_permutation__round__N5661 ) );
  AND2_X2 _f_permutation__round__U49  ( .A1(_f_permutation__round__n514 ), 
        .A2(_f_permutation__round__c[1081] ), .ZN(
        _f_permutation__round__N5663 ) );
  AND2_X2 _f_permutation__round__U48  ( .A1(_f_permutation__round__n519 ), 
        .A2(_f_permutation__round__c[1080] ), .ZN(
        _f_permutation__round__N5665 ) );
  AND2_X2 _f_permutation__round__U47  ( .A1(_f_permutation__round__n524 ), 
        .A2(_f_permutation__round__c[1079] ), .ZN(
        _f_permutation__round__N5667 ) );
  AND2_X2 _f_permutation__round__U46  ( .A1(_f_permutation__round__n529 ), 
        .A2(_f_permutation__round__c[1078] ), .ZN(
        _f_permutation__round__N5669 ) );
  AND2_X2 _f_permutation__round__U45  ( .A1(_f_permutation__round__n534 ), 
        .A2(_f_permutation__round__c[1077] ), .ZN(
        _f_permutation__round__N5671 ) );
  AND2_X2 _f_permutation__round__U44  ( .A1(_f_permutation__round__n539 ), 
        .A2(_f_permutation__round__c[1076] ), .ZN(
        _f_permutation__round__N5673 ) );
  AND2_X2 _f_permutation__round__U43  ( .A1(_f_permutation__round__n544 ), 
        .A2(_f_permutation__round__c[1075] ), .ZN(
        _f_permutation__round__N5675 ) );
  AND2_X2 _f_permutation__round__U42  ( .A1(_f_permutation__round__n549 ), 
        .A2(_f_permutation__round__c[1074] ), .ZN(
        _f_permutation__round__N5677 ) );
  AND2_X2 _f_permutation__round__U41  ( .A1(_f_permutation__round__n554 ), 
        .A2(_f_permutation__round__c[1073] ), .ZN(
        _f_permutation__round__N5679 ) );
  AND2_X2 _f_permutation__round__U40  ( .A1(_f_permutation__round__n559 ), 
        .A2(_f_permutation__round__c[1072] ), .ZN(
        _f_permutation__round__N5681 ) );
  AND2_X2 _f_permutation__round__U39  ( .A1(_f_permutation__round__n564 ), 
        .A2(_f_permutation__round__c[1071] ), .ZN(
        _f_permutation__round__N5683 ) );
  AND2_X2 _f_permutation__round__U38  ( .A1(_f_permutation__round__n569 ), 
        .A2(_f_permutation__round__c[1070] ), .ZN(
        _f_permutation__round__N5685 ) );
  AND2_X2 _f_permutation__round__U37  ( .A1(_f_permutation__round__n574 ), 
        .A2(_f_permutation__round__c[1069] ), .ZN(
        _f_permutation__round__N5687 ) );
  AND2_X2 _f_permutation__round__U36  ( .A1(_f_permutation__round__n579 ), 
        .A2(_f_permutation__round__c[1068] ), .ZN(
        _f_permutation__round__N5689 ) );
  AND2_X2 _f_permutation__round__U35  ( .A1(_f_permutation__round__n584 ), 
        .A2(_f_permutation__round__c[1067] ), .ZN(
        _f_permutation__round__N5691 ) );
  AND2_X2 _f_permutation__round__U34  ( .A1(_f_permutation__round__n589 ), 
        .A2(_f_permutation__round__c[1066] ), .ZN(
        _f_permutation__round__N5693 ) );
  AND2_X2 _f_permutation__round__U33  ( .A1(_f_permutation__round__n594 ), 
        .A2(_f_permutation__round__c[1065] ), .ZN(
        _f_permutation__round__N5695 ) );
  AND2_X2 _f_permutation__round__U32  ( .A1(_f_permutation__round__n599 ), 
        .A2(_f_permutation__round__c[1064] ), .ZN(
        _f_permutation__round__N5697 ) );
  AND2_X2 _f_permutation__round__U31  ( .A1(_f_permutation__round__n604 ), 
        .A2(_f_permutation__round__c[1063] ), .ZN(
        _f_permutation__round__N5699 ) );
  AND2_X2 _f_permutation__round__U30  ( .A1(_f_permutation__round__n609 ), 
        .A2(_f_permutation__round__c[1062] ), .ZN(
        _f_permutation__round__N5701 ) );
  AND2_X2 _f_permutation__round__U29  ( .A1(_f_permutation__round__n614 ), 
        .A2(_f_permutation__round__c[1061] ), .ZN(
        _f_permutation__round__N5703 ) );
  AND2_X2 _f_permutation__round__U28  ( .A1(_f_permutation__round__n619 ), 
        .A2(_f_permutation__round__c[1060] ), .ZN(
        _f_permutation__round__N5705 ) );
  AND2_X2 _f_permutation__round__U27  ( .A1(_f_permutation__round__n624 ), 
        .A2(_f_permutation__round__c[1059] ), .ZN(
        _f_permutation__round__N5707 ) );
  AND2_X2 _f_permutation__round__U26  ( .A1(_f_permutation__round__n629 ), 
        .A2(_f_permutation__round__c[1058] ), .ZN(
        _f_permutation__round__N5709 ) );
  AND2_X2 _f_permutation__round__U25  ( .A1(_f_permutation__round__n634 ), 
        .A2(_f_permutation__round__c[1057] ), .ZN(
        _f_permutation__round__N5711 ) );
  AND2_X2 _f_permutation__round__U24  ( .A1(_f_permutation__round__n639 ), 
        .A2(_f_permutation__round__c[1056] ), .ZN(
        _f_permutation__round__N5713 ) );
  AND2_X2 _f_permutation__round__U23  ( .A1(_f_permutation__round__n644 ), 
        .A2(_f_permutation__round__c[1055] ), .ZN(
        _f_permutation__round__N5715 ) );
  AND2_X2 _f_permutation__round__U22  ( .A1(_f_permutation__round__n649 ), 
        .A2(_f_permutation__round__c[1054] ), .ZN(
        _f_permutation__round__N5717 ) );
  AND2_X2 _f_permutation__round__U21  ( .A1(_f_permutation__round__n654 ), 
        .A2(_f_permutation__round__c[1053] ), .ZN(
        _f_permutation__round__N5719 ) );
  AND2_X2 _f_permutation__round__U20  ( .A1(_f_permutation__round__n659 ), 
        .A2(_f_permutation__round__c[1052] ), .ZN(
        _f_permutation__round__N5721 ) );
  AND2_X2 _f_permutation__round__U19  ( .A1(_f_permutation__round__n664 ), 
        .A2(_f_permutation__round__c[1051] ), .ZN(
        _f_permutation__round__N5723 ) );
  AND2_X2 _f_permutation__round__U18  ( .A1(_f_permutation__round__n669 ), 
        .A2(_f_permutation__round__c[1050] ), .ZN(
        _f_permutation__round__N5725 ) );
  AND2_X2 _f_permutation__round__U17  ( .A1(_f_permutation__round__n674 ), 
        .A2(_f_permutation__round__c[1049] ), .ZN(
        _f_permutation__round__N5727 ) );
  AND2_X2 _f_permutation__round__U16  ( .A1(_f_permutation__round__n679 ), 
        .A2(_f_permutation__round__c[1048] ), .ZN(
        _f_permutation__round__N5729 ) );
  AND2_X2 _f_permutation__round__U15  ( .A1(_f_permutation__round__n684 ), 
        .A2(_f_permutation__round__c[1047] ), .ZN(
        _f_permutation__round__N5731 ) );
  AND2_X2 _f_permutation__round__U14  ( .A1(_f_permutation__round__n689 ), 
        .A2(_f_permutation__round__c[1046] ), .ZN(
        _f_permutation__round__N5733 ) );
  AND2_X2 _f_permutation__round__U13  ( .A1(_f_permutation__round__n694 ), 
        .A2(_f_permutation__round__c[1045] ), .ZN(
        _f_permutation__round__N5735 ) );
  AND2_X2 _f_permutation__round__U12  ( .A1(_f_permutation__round__n699 ), 
        .A2(_f_permutation__round__c[1044] ), .ZN(
        _f_permutation__round__N5737 ) );
  AND2_X2 _f_permutation__round__U11  ( .A1(_f_permutation__round__n704 ), 
        .A2(_f_permutation__round__c[1043] ), .ZN(
        _f_permutation__round__N5739 ) );
  AND2_X2 _f_permutation__round__U10  ( .A1(_f_permutation__round__n709 ), 
        .A2(_f_permutation__round__c[1042] ), .ZN(
        _f_permutation__round__N5741 ) );
  AND2_X2 _f_permutation__round__U9  ( .A1(_f_permutation__round__n714 ), .A2(
        _f_permutation__round__c[1041] ), .ZN(_f_permutation__round__N5743 )
         );
  AND2_X2 _f_permutation__round__U8  ( .A1(_f_permutation__round__n719 ), .A2(
        _f_permutation__round__c[1040] ), .ZN(_f_permutation__round__N5745 )
         );
  AND2_X2 _f_permutation__round__U7  ( .A1(_f_permutation__round__n724 ), .A2(
        _f_permutation__round__c[1039] ), .ZN(_f_permutation__round__N5747 )
         );
  AND2_X2 _f_permutation__round__U6  ( .A1(_f_permutation__round__n729 ), .A2(
        _f_permutation__round__c[1038] ), .ZN(_f_permutation__round__N5749 )
         );
  AND2_X2 _f_permutation__round__U5  ( .A1(_f_permutation__round__n734 ), .A2(
        _f_permutation__round__c[1037] ), .ZN(_f_permutation__round__N5751 )
         );
  AND2_X2 _f_permutation__round__U4  ( .A1(_f_permutation__round__n739 ), .A2(
        _f_permutation__round__c[1036] ), .ZN(_f_permutation__round__N5753 )
         );
  AND2_X2 _f_permutation__round__U3  ( .A1(_f_permutation__round__n744 ), .A2(
        _f_permutation__round__c[1035] ), .ZN(_f_permutation__round__N5755 )
         );
  AND2_X2 _f_permutation__round__U2  ( .A1(_f_permutation__round__n749 ), .A2(
        _f_permutation__round__c[1034] ), .ZN(_f_permutation__round__N5757 )
         );
  AND2_X2 _f_permutation__round__U1  ( .A1(_f_permutation__round__n754 ), .A2(
        _f_permutation__round__c[1033] ), .ZN(_f_permutation__round__N5759 )
         );
  XOR2_X2 _f_permutation__round__U7367  ( .A(_f_permutation__round__n962 ), 
        .B(_f_permutation__round__n961 ), .Z(_f_permutation__round__n2125 ) );
  XOR2_X2 _f_permutation__round__U7366  ( .A(SYNOPSYS_UNCONNECTED_834), .B(
        _f_permutation__round__n963 ), .Z(_f_permutation__round__n961 ) );
  XOR2_X2 _f_permutation__round__U7365  ( .A(SYNOPSYS_UNCONNECTED_194), .B(
        SYNOPSYS_UNCONNECTED_514), .Z(_f_permutation__round__n962 ) );
  XOR2_X2 _f_permutation__round__U7364  ( .A(_f_permutation__round_in[1534]), 
        .B(_f_permutation__round_in[1214]), .Z(_f_permutation__round__n963 )
         );
  XOR2_X2 _f_permutation__round__U7363  ( .A(_f_permutation__round__n965 ), 
        .B(_f_permutation__round__n964 ), .Z(_f_permutation__round__n25650 )
         );
  XOR2_X2 _f_permutation__round__U7362  ( .A(SYNOPSYS_UNCONNECTED_1025), .B(
        _f_permutation__round__n966 ), .Z(_f_permutation__round__n964 ) );
  XOR2_X2 _f_permutation__round__U7361  ( .A(SYNOPSYS_UNCONNECTED_385), .B(
        SYNOPSYS_UNCONNECTED_705), .Z(_f_permutation__round__n965 ) );
  XOR2_X2 _f_permutation__round__U7360  ( .A(_f_permutation__round_in[1343]), 
        .B(SYNOPSYS_UNCONNECTED_65), .Z(_f_permutation__round__n966 ) );
  XOR2_X2 _f_permutation__round__U7359  ( .A(_f_permutation__round__n2125 ), 
        .B(_f_permutation__round__n25650 ), .Z(_f_permutation__round__n2126 )
         );
  XOR2_X2 _f_permutation__round__U7358  ( .A(_f_permutation__round_in[1599]), 
        .B(_f_permutation__round__n2126 ), .Z(_f_permutation__round__c[63] )
         );
  XOR2_X2 _f_permutation__round__U7357  ( .A(_f_permutation__round__n968 ), 
        .B(_f_permutation__round__n967 ), .Z(_f_permutation__round__n1928 ) );
  XOR2_X2 _f_permutation__round__U7356  ( .A(SYNOPSYS_UNCONNECTED_769), .B(
        _f_permutation__round__n969 ), .Z(_f_permutation__round__n967 ) );
  XOR2_X2 _f_permutation__round__U7355  ( .A(SYNOPSYS_UNCONNECTED_129), .B(
        SYNOPSYS_UNCONNECTED_449), .Z(_f_permutation__round__n968 ) );
  XOR2_X2 _f_permutation__round__U7354  ( .A(_f_permutation__round_in[1599]), 
        .B(_f_permutation__round_in[1279]), .Z(_f_permutation__round__n969 )
         );
  XOR2_X2 _f_permutation__round__U7353  ( .A(_f_permutation__round__n971 ), 
        .B(_f_permutation__round__n970 ), .Z(_f_permutation__round__n2368 ) );
  XOR2_X2 _f_permutation__round__U7352  ( .A(SYNOPSYS_UNCONNECTED_1024), .B(
        _f_permutation__round__n972 ), .Z(_f_permutation__round__n970 ) );
  XOR2_X2 _f_permutation__round__U7351  ( .A(SYNOPSYS_UNCONNECTED_384), .B(
        SYNOPSYS_UNCONNECTED_704), .Z(_f_permutation__round__n971 ) );
  XOR2_X2 _f_permutation__round__U7350  ( .A(_f_permutation__round_in[1344]), 
        .B(_f_permutation__round_in[1024]), .Z(_f_permutation__round__n972 )
         );
  XOR2_X2 _f_permutation__round__U7349  ( .A(_f_permutation__round__n1928 ), 
        .B(_f_permutation__round__n2368 ), .Z(_f_permutation__round__n1929 )
         );
  XOR2_X2 _f_permutation__round__U7348  ( .A(SYNOPSYS_UNCONNECTED_1088), .B(
        _f_permutation__round__n1929 ), .Z(_f_permutation__round__c[1536] ) );
  XOR2_X2 _f_permutation__round__U7347  ( .A(_f_permutation__round__n974 ), 
        .B(_f_permutation__round__n973 ), .Z(_f_permutation__round__n2380 ) );
  XOR2_X2 _f_permutation__round__U7346  ( .A(SYNOPSYS_UNCONNECTED_898), .B(
        _f_permutation__round__n975 ), .Z(_f_permutation__round__n973 ) );
  XOR2_X2 _f_permutation__round__U7345  ( .A(SYNOPSYS_UNCONNECTED_258), .B(
        SYNOPSYS_UNCONNECTED_578), .Z(_f_permutation__round__n974 ) );
  XOR2_X2 _f_permutation__round__U7344  ( .A(_f_permutation__round_in[1470]), 
        .B(_f_permutation__round_in[1150]), .Z(_f_permutation__round__n975 )
         );
  XOR2_X2 _f_permutation__round__U7343  ( .A(_f_permutation__round__n1928 ), 
        .B(_f_permutation__round__n2380 ), .Z(_f_permutation__round__n1930 )
         );
  XOR2_X2 _f_permutation__round__U7342  ( .A(SYNOPSYS_UNCONNECTED_833), .B(
        _f_permutation__round__n1930 ), .Z(_f_permutation__round__c[639] ) );
  XOR2_X2 _f_permutation__round__U7341  ( .A(SYNOPSYS_UNCONNECTED_768), .B(
        _f_permutation__round__n1929 ), .Z(_f_permutation__round__c[1472] ) );
  XOR2_X2 _f_permutation__round__U7340  ( .A(SYNOPSYS_UNCONNECTED_513), .B(
        _f_permutation__round__n1930 ), .Z(_f_permutation__round__c[575] ) );
  XOR2_X2 _f_permutation__round__U7339  ( .A(SYNOPSYS_UNCONNECTED_448), .B(
        _f_permutation__round__n1929 ), .Z(_f_permutation__round__c[1408] ) );
  XOR2_X2 _f_permutation__round__U7338  ( .A(SYNOPSYS_UNCONNECTED_193), .B(
        _f_permutation__round__n1930 ), .Z(_f_permutation__round__c[511] ) );
  XOR2_X2 _f_permutation__round__U7337  ( .A(SYNOPSYS_UNCONNECTED_128), .B(
        _f_permutation__round__n1929 ), .Z(_f_permutation__round__c[1344] ) );
  XOR2_X2 _f_permutation__round__U7336  ( .A(_f_permutation__round_in[1215]), 
        .B(_f_permutation__round__n1930 ), .Z(_f_permutation__round__c[447] )
         );
  XOR2_X2 _f_permutation__round__U7335  ( .A(_f_permutation__round_in[1280]), 
        .B(_f_permutation__round__n1929 ), .Z(_f_permutation__round__c[1280] )
         );
  XOR2_X2 _f_permutation__round__U7334  ( .A(_f_permutation__round_in[1535]), 
        .B(_f_permutation__round__n1930 ), .Z(_f_permutation__round__c[383] )
         );
  XOR2_X2 _f_permutation__round__U7333  ( .A(_f_permutation__round__n977 ), 
        .B(_f_permutation__round__n976 ), .Z(_f_permutation__round__n2129 ) );
  XOR2_X2 _f_permutation__round__U7332  ( .A(SYNOPSYS_UNCONNECTED_835), .B(
        _f_permutation__round__n978 ), .Z(_f_permutation__round__n976 ) );
  XOR2_X2 _f_permutation__round__U7331  ( .A(SYNOPSYS_UNCONNECTED_195), .B(
        SYNOPSYS_UNCONNECTED_515), .Z(_f_permutation__round__n977 ) );
  XOR2_X2 _f_permutation__round__U7330  ( .A(_f_permutation__round_in[1533]), 
        .B(_f_permutation__round_in[1213]), .Z(_f_permutation__round__n978 )
         );
  XOR2_X2 _f_permutation__round__U7329  ( .A(_f_permutation__round__n980 ), 
        .B(_f_permutation__round__n979 ), .Z(_f_permutation__round__n2376 ) );
  XOR2_X2 _f_permutation__round__U7328  ( .A(SYNOPSYS_UNCONNECTED_1026), .B(
        _f_permutation__round__n981 ), .Z(_f_permutation__round__n979 ) );
  XOR2_X2 _f_permutation__round__U7327  ( .A(SYNOPSYS_UNCONNECTED_386), .B(
        SYNOPSYS_UNCONNECTED_706), .Z(_f_permutation__round__n980 ) );
  XOR2_X2 _f_permutation__round__U7326  ( .A(_f_permutation__round_in[1342]), 
        .B(SYNOPSYS_UNCONNECTED_66), .Z(_f_permutation__round__n981 ) );
  XOR2_X2 _f_permutation__round__U7325  ( .A(_f_permutation__round__n2129 ), 
        .B(_f_permutation__round__n2376 ), .Z(_f_permutation__round__n2130 )
         );
  XOR2_X2 _f_permutation__round__U7324  ( .A(_f_permutation__round_in[1598]), 
        .B(_f_permutation__round__n2130 ), .Z(_f_permutation__round__c[62] )
         );
  XOR2_X2 _f_permutation__round__U7323  ( .A(_f_permutation__round__n983 ), 
        .B(_f_permutation__round__n982 ), .Z(_f_permutation__round__n1931 ) );
  XOR2_X2 _f_permutation__round__U7322  ( .A(SYNOPSYS_UNCONNECTED_770), .B(
        _f_permutation__round__n984 ), .Z(_f_permutation__round__n982 ) );
  XOR2_X2 _f_permutation__round__U7321  ( .A(SYNOPSYS_UNCONNECTED_130), .B(
        SYNOPSYS_UNCONNECTED_450), .Z(_f_permutation__round__n983 ) );
  XOR2_X2 _f_permutation__round__U7320  ( .A(_f_permutation__round_in[1598]), 
        .B(_f_permutation__round_in[1278]), .Z(_f_permutation__round__n984 )
         );
  XOR2_X2 _f_permutation__round__U7319  ( .A(_f_permutation__round__n986 ), 
        .B(_f_permutation__round__n985 ), .Z(_f_permutation__round__n2372 ) );
  XOR2_X2 _f_permutation__round__U7318  ( .A(SYNOPSYS_UNCONNECTED_961), .B(
        _f_permutation__round__n987 ), .Z(_f_permutation__round__n985 ) );
  XOR2_X2 _f_permutation__round__U7317  ( .A(SYNOPSYS_UNCONNECTED_321), .B(
        SYNOPSYS_UNCONNECTED_641), .Z(_f_permutation__round__n986 ) );
  XOR2_X2 _f_permutation__round__U7316  ( .A(_f_permutation__round_in[1407]), 
        .B(_f_permutation__round_in[1087]), .Z(_f_permutation__round__n987 )
         );
  XOR2_X2 _f_permutation__round__U7315  ( .A(_f_permutation__round__n1931 ), 
        .B(_f_permutation__round__n2372 ), .Z(_f_permutation__round__n1932 )
         );
  XOR2_X2 _f_permutation__round__U7314  ( .A(SYNOPSYS_UNCONNECTED_1025), .B(
        _f_permutation__round__n1932 ), .Z(_f_permutation__round__c[1599] ) );
  XOR2_X2 _f_permutation__round__U7313  ( .A(_f_permutation__round__n989 ), 
        .B(_f_permutation__round__n988 ), .Z(_f_permutation__round__n2383 ) );
  XOR2_X2 _f_permutation__round__U7312  ( .A(SYNOPSYS_UNCONNECTED_899), .B(
        _f_permutation__round__n990 ), .Z(_f_permutation__round__n988 ) );
  XOR2_X2 _f_permutation__round__U7311  ( .A(SYNOPSYS_UNCONNECTED_259), .B(
        SYNOPSYS_UNCONNECTED_579), .Z(_f_permutation__round__n989 ) );
  XOR2_X2 _f_permutation__round__U7310  ( .A(_f_permutation__round_in[1469]), 
        .B(_f_permutation__round_in[1149]), .Z(_f_permutation__round__n990 )
         );
  XOR2_X2 _f_permutation__round__U7309  ( .A(_f_permutation__round__n1931 ), 
        .B(_f_permutation__round__n2383 ), .Z(_f_permutation__round__n1933 )
         );
  XOR2_X2 _f_permutation__round__U7308  ( .A(SYNOPSYS_UNCONNECTED_834), .B(
        _f_permutation__round__n1933 ), .Z(_f_permutation__round__c[638] ) );
  XOR2_X2 _f_permutation__round__U7307  ( .A(SYNOPSYS_UNCONNECTED_705), .B(
        _f_permutation__round__n1932 ), .Z(_f_permutation__round__c[1535] ) );
  XOR2_X2 _f_permutation__round__U7306  ( .A(SYNOPSYS_UNCONNECTED_514), .B(
        _f_permutation__round__n1933 ), .Z(_f_permutation__round__c[574] ) );
  XOR2_X2 _f_permutation__round__U7305  ( .A(SYNOPSYS_UNCONNECTED_385), .B(
        _f_permutation__round__n1932 ), .Z(_f_permutation__round__c[1471] ) );
  XOR2_X2 _f_permutation__round__U7304  ( .A(SYNOPSYS_UNCONNECTED_194), .B(
        _f_permutation__round__n1933 ), .Z(_f_permutation__round__c[510] ) );
  XOR2_X2 _f_permutation__round__U7303  ( .A(SYNOPSYS_UNCONNECTED_65), .B(
        _f_permutation__round__n1932 ), .Z(_f_permutation__round__c[1407] ) );
  XOR2_X2 _f_permutation__round__U7302  ( .A(_f_permutation__round_in[1214]), 
        .B(_f_permutation__round__n1933 ), .Z(_f_permutation__round__c[446] )
         );
  XOR2_X2 _f_permutation__round__U7301  ( .A(_f_permutation__round_in[1343]), 
        .B(_f_permutation__round__n1932 ), .Z(_f_permutation__round__c[1343] )
         );
  XOR2_X2 _f_permutation__round__U7300  ( .A(_f_permutation__round_in[1534]), 
        .B(_f_permutation__round__n1933 ), .Z(_f_permutation__round__c[382] )
         );
  XOR2_X2 _f_permutation__round__U7299  ( .A(_f_permutation__round__n992 ), 
        .B(_f_permutation__round__n991 ), .Z(_f_permutation__round__n2133 ) );
  XOR2_X2 _f_permutation__round__U7298  ( .A(SYNOPSYS_UNCONNECTED_836), .B(
        _f_permutation__round__n993 ), .Z(_f_permutation__round__n991 ) );
  XOR2_X2 _f_permutation__round__U7297  ( .A(SYNOPSYS_UNCONNECTED_196), .B(
        SYNOPSYS_UNCONNECTED_516), .Z(_f_permutation__round__n992 ) );
  XOR2_X2 _f_permutation__round__U7296  ( .A(_f_permutation__round_in[1532]), 
        .B(_f_permutation__round_in[1212]), .Z(_f_permutation__round__n993 )
         );
  XOR2_X2 _f_permutation__round__U7295  ( .A(_f_permutation__round__n995 ), 
        .B(_f_permutation__round__n994 ), .Z(_f_permutation__round__n2379 ) );
  XOR2_X2 _f_permutation__round__U7294  ( .A(SYNOPSYS_UNCONNECTED_1027), .B(
        _f_permutation__round__n996 ), .Z(_f_permutation__round__n994 ) );
  XOR2_X2 _f_permutation__round__U7293  ( .A(SYNOPSYS_UNCONNECTED_387), .B(
        SYNOPSYS_UNCONNECTED_707), .Z(_f_permutation__round__n995 ) );
  XOR2_X2 _f_permutation__round__U7292  ( .A(_f_permutation__round_in[1341]), 
        .B(SYNOPSYS_UNCONNECTED_67), .Z(_f_permutation__round__n996 ) );
  XOR2_X2 _f_permutation__round__U7291  ( .A(_f_permutation__round__n2133 ), 
        .B(_f_permutation__round__n2379 ), .Z(_f_permutation__round__n2134 )
         );
  XOR2_X2 _f_permutation__round__U7290  ( .A(_f_permutation__round_in[1597]), 
        .B(_f_permutation__round__n2134 ), .Z(_f_permutation__round__c[61] )
         );
  XOR2_X2 _f_permutation__round__U7289  ( .A(_f_permutation__round__n998 ), 
        .B(_f_permutation__round__n997 ), .Z(_f_permutation__round__n1934 ) );
  XOR2_X2 _f_permutation__round__U7288  ( .A(SYNOPSYS_UNCONNECTED_771), .B(
        _f_permutation__round__n999 ), .Z(_f_permutation__round__n997 ) );
  XOR2_X2 _f_permutation__round__U7287  ( .A(SYNOPSYS_UNCONNECTED_131), .B(
        SYNOPSYS_UNCONNECTED_451), .Z(_f_permutation__round__n998 ) );
  XOR2_X2 _f_permutation__round__U7286  ( .A(_f_permutation__round_in[1597]), 
        .B(_f_permutation__round_in[1277]), .Z(_f_permutation__round__n999 )
         );
  XOR2_X2 _f_permutation__round__U7285  ( .A(_f_permutation__round__n1001 ), 
        .B(_f_permutation__round__n1000 ), .Z(_f_permutation__round__n2120 )
         );
  XOR2_X2 _f_permutation__round__U7284  ( .A(SYNOPSYS_UNCONNECTED_962), .B(
        _f_permutation__round__n1002 ), .Z(_f_permutation__round__n1000 ) );
  XOR2_X2 _f_permutation__round__U7283  ( .A(SYNOPSYS_UNCONNECTED_322), .B(
        SYNOPSYS_UNCONNECTED_642), .Z(_f_permutation__round__n1001 ) );
  XOR2_X2 _f_permutation__round__U7282  ( .A(_f_permutation__round_in[1406]), 
        .B(_f_permutation__round_in[1086]), .Z(_f_permutation__round__n1002 )
         );
  XOR2_X2 _f_permutation__round__U7281  ( .A(_f_permutation__round__n1934 ), 
        .B(_f_permutation__round__n2120 ), .Z(_f_permutation__round__n1935 )
         );
  XOR2_X2 _f_permutation__round__U7280  ( .A(SYNOPSYS_UNCONNECTED_1026), .B(
        _f_permutation__round__n1935 ), .Z(_f_permutation__round__c[1598] ) );
  XOR2_X2 _f_permutation__round__U7279  ( .A(_f_permutation__round__n1004 ), 
        .B(_f_permutation__round__n1003 ), .Z(_f_permutation__round__n2386 )
         );
  XOR2_X2 _f_permutation__round__U7278  ( .A(SYNOPSYS_UNCONNECTED_900), .B(
        _f_permutation__round__n1005 ), .Z(_f_permutation__round__n1003 ) );
  XOR2_X2 _f_permutation__round__U7277  ( .A(SYNOPSYS_UNCONNECTED_260), .B(
        SYNOPSYS_UNCONNECTED_580), .Z(_f_permutation__round__n1004 ) );
  XOR2_X2 _f_permutation__round__U7276  ( .A(_f_permutation__round_in[1468]), 
        .B(_f_permutation__round_in[1148]), .Z(_f_permutation__round__n1005 )
         );
  XOR2_X2 _f_permutation__round__U7275  ( .A(_f_permutation__round__n1934 ), 
        .B(_f_permutation__round__n2386 ), .Z(_f_permutation__round__n1936 )
         );
  XOR2_X2 _f_permutation__round__U7274  ( .A(SYNOPSYS_UNCONNECTED_835), .B(
        _f_permutation__round__n1936 ), .Z(_f_permutation__round__c[637] ) );
  XOR2_X2 _f_permutation__round__U7273  ( .A(SYNOPSYS_UNCONNECTED_706), .B(
        _f_permutation__round__n1935 ), .Z(_f_permutation__round__c[1534] ) );
  XOR2_X2 _f_permutation__round__U7272  ( .A(SYNOPSYS_UNCONNECTED_515), .B(
        _f_permutation__round__n1936 ), .Z(_f_permutation__round__c[573] ) );
  XOR2_X2 _f_permutation__round__U7271  ( .A(SYNOPSYS_UNCONNECTED_386), .B(
        _f_permutation__round__n1935 ), .Z(_f_permutation__round__c[1470] ) );
  XOR2_X2 _f_permutation__round__U7270  ( .A(SYNOPSYS_UNCONNECTED_195), .B(
        _f_permutation__round__n1936 ), .Z(_f_permutation__round__c[509] ) );
  XOR2_X2 _f_permutation__round__U7269  ( .A(SYNOPSYS_UNCONNECTED_66), .B(
        _f_permutation__round__n1935 ), .Z(_f_permutation__round__c[1406] ) );
  XOR2_X2 _f_permutation__round__U7268  ( .A(_f_permutation__round_in[1213]), 
        .B(_f_permutation__round__n1936 ), .Z(_f_permutation__round__c[445] )
         );
  XOR2_X2 _f_permutation__round__U7267  ( .A(_f_permutation__round_in[1342]), 
        .B(_f_permutation__round__n1935 ), .Z(_f_permutation__round__c[1342] )
         );
  XOR2_X2 _f_permutation__round__U7266  ( .A(_f_permutation__round_in[1533]), 
        .B(_f_permutation__round__n1936 ), .Z(_f_permutation__round__c[381] )
         );
  XOR2_X2 _f_permutation__round__U7265  ( .A(_f_permutation__round__n1007 ), 
        .B(_f_permutation__round__n1006 ), .Z(_f_permutation__round__n2137 )
         );
  XOR2_X2 _f_permutation__round__U7264  ( .A(SYNOPSYS_UNCONNECTED_837), .B(
        _f_permutation__round__n1008 ), .Z(_f_permutation__round__n1006 ) );
  XOR2_X2 _f_permutation__round__U7263  ( .A(SYNOPSYS_UNCONNECTED_197), .B(
        SYNOPSYS_UNCONNECTED_517), .Z(_f_permutation__round__n1007 ) );
  XOR2_X2 _f_permutation__round__U7262  ( .A(_f_permutation__round_in[1531]), 
        .B(_f_permutation__round_in[1211]), .Z(_f_permutation__round__n1008 )
         );
  XOR2_X2 _f_permutation__round__U7261  ( .A(_f_permutation__round__n1010 ), 
        .B(_f_permutation__round__n1009 ), .Z(_f_permutation__round__n2382 )
         );
  XOR2_X2 _f_permutation__round__U7260  ( .A(SYNOPSYS_UNCONNECTED_1028), .B(
        _f_permutation__round__n1011 ), .Z(_f_permutation__round__n1009 ) );
  XOR2_X2 _f_permutation__round__U7259  ( .A(SYNOPSYS_UNCONNECTED_388), .B(
        SYNOPSYS_UNCONNECTED_708), .Z(_f_permutation__round__n1010 ) );
  XOR2_X2 _f_permutation__round__U7258  ( .A(_f_permutation__round_in[1340]), 
        .B(SYNOPSYS_UNCONNECTED_68), .Z(_f_permutation__round__n1011 ) );
  XOR2_X2 _f_permutation__round__U7257  ( .A(_f_permutation__round__n2137 ), 
        .B(_f_permutation__round__n2382 ), .Z(_f_permutation__round__n2138 )
         );
  XOR2_X2 _f_permutation__round__U7256  ( .A(_f_permutation__round_in[1596]), 
        .B(_f_permutation__round__n2138 ), .Z(_f_permutation__round__c[60] )
         );
  XOR2_X2 _f_permutation__round__U7255  ( .A(_f_permutation__round__n1013 ), 
        .B(_f_permutation__round__n1012 ), .Z(_f_permutation__round__n1937 )
         );
  XOR2_X2 _f_permutation__round__U7254  ( .A(SYNOPSYS_UNCONNECTED_772), .B(
        _f_permutation__round__n1014 ), .Z(_f_permutation__round__n1012 ) );
  XOR2_X2 _f_permutation__round__U7253  ( .A(SYNOPSYS_UNCONNECTED_132), .B(
        SYNOPSYS_UNCONNECTED_452), .Z(_f_permutation__round__n1013 ) );
  XOR2_X2 _f_permutation__round__U7252  ( .A(_f_permutation__round_in[1596]), 
        .B(_f_permutation__round_in[1276]), .Z(_f_permutation__round__n1014 )
         );
  XOR2_X2 _f_permutation__round__U7251  ( .A(_f_permutation__round__n1016 ), 
        .B(_f_permutation__round__n1015 ), .Z(_f_permutation__round__n2124 )
         );
  XOR2_X2 _f_permutation__round__U7250  ( .A(SYNOPSYS_UNCONNECTED_963), .B(
        _f_permutation__round__n1017 ), .Z(_f_permutation__round__n1015 ) );
  XOR2_X2 _f_permutation__round__U7249  ( .A(SYNOPSYS_UNCONNECTED_323), .B(
        SYNOPSYS_UNCONNECTED_643), .Z(_f_permutation__round__n1016 ) );
  XOR2_X2 _f_permutation__round__U7248  ( .A(_f_permutation__round_in[1405]), 
        .B(_f_permutation__round_in[1085]), .Z(_f_permutation__round__n1017 )
         );
  XOR2_X2 _f_permutation__round__U7247  ( .A(_f_permutation__round__n1937 ), 
        .B(_f_permutation__round__n2124 ), .Z(_f_permutation__round__n1938 )
         );
  XOR2_X2 _f_permutation__round__U7246  ( .A(SYNOPSYS_UNCONNECTED_1027), .B(
        _f_permutation__round__n1938 ), .Z(_f_permutation__round__c[1597] ) );
  XOR2_X2 _f_permutation__round__U7245  ( .A(_f_permutation__round__n1019 ), 
        .B(_f_permutation__round__n1018 ), .Z(_f_permutation__round__n2389 )
         );
  XOR2_X2 _f_permutation__round__U7244  ( .A(SYNOPSYS_UNCONNECTED_901), .B(
        _f_permutation__round__n1020 ), .Z(_f_permutation__round__n1018 ) );
  XOR2_X2 _f_permutation__round__U7243  ( .A(SYNOPSYS_UNCONNECTED_261), .B(
        SYNOPSYS_UNCONNECTED_581), .Z(_f_permutation__round__n1019 ) );
  XOR2_X2 _f_permutation__round__U7242  ( .A(_f_permutation__round_in[1467]), 
        .B(_f_permutation__round_in[1147]), .Z(_f_permutation__round__n1020 )
         );
  XOR2_X2 _f_permutation__round__U7241  ( .A(_f_permutation__round__n1937 ), 
        .B(_f_permutation__round__n2389 ), .Z(_f_permutation__round__n1939 )
         );
  XOR2_X2 _f_permutation__round__U7240  ( .A(SYNOPSYS_UNCONNECTED_836), .B(
        _f_permutation__round__n1939 ), .Z(_f_permutation__round__c[636] ) );
  XOR2_X2 _f_permutation__round__U7239  ( .A(SYNOPSYS_UNCONNECTED_707), .B(
        _f_permutation__round__n1938 ), .Z(_f_permutation__round__c[1533] ) );
  XOR2_X2 _f_permutation__round__U7238  ( .A(SYNOPSYS_UNCONNECTED_516), .B(
        _f_permutation__round__n1939 ), .Z(_f_permutation__round__c[572] ) );
  XOR2_X2 _f_permutation__round__U7237  ( .A(SYNOPSYS_UNCONNECTED_387), .B(
        _f_permutation__round__n1938 ), .Z(_f_permutation__round__c[1469] ) );
  XOR2_X2 _f_permutation__round__U7236  ( .A(SYNOPSYS_UNCONNECTED_196), .B(
        _f_permutation__round__n1939 ), .Z(_f_permutation__round__c[508] ) );
  XOR2_X2 _f_permutation__round__U7235  ( .A(SYNOPSYS_UNCONNECTED_67), .B(
        _f_permutation__round__n1938 ), .Z(_f_permutation__round__c[1405] ) );
  XOR2_X2 _f_permutation__round__U7234  ( .A(_f_permutation__round_in[1212]), 
        .B(_f_permutation__round__n1939 ), .Z(_f_permutation__round__c[444] )
         );
  XOR2_X2 _f_permutation__round__U7233  ( .A(_f_permutation__round_in[1341]), 
        .B(_f_permutation__round__n1938 ), .Z(_f_permutation__round__c[1341] )
         );
  XOR2_X2 _f_permutation__round__U7232  ( .A(_f_permutation__round_in[1532]), 
        .B(_f_permutation__round__n1939 ), .Z(_f_permutation__round__c[380] )
         );
  XOR2_X2 _f_permutation__round__U7231  ( .A(_f_permutation__round__n1022 ), 
        .B(_f_permutation__round__n1021 ), .Z(_f_permutation__round__n2141 )
         );
  XOR2_X2 _f_permutation__round__U7230  ( .A(SYNOPSYS_UNCONNECTED_838), .B(
        _f_permutation__round__n1023 ), .Z(_f_permutation__round__n1021 ) );
  XOR2_X2 _f_permutation__round__U7229  ( .A(SYNOPSYS_UNCONNECTED_198), .B(
        SYNOPSYS_UNCONNECTED_518), .Z(_f_permutation__round__n1022 ) );
  XOR2_X2 _f_permutation__round__U7228  ( .A(_f_permutation__round_in[1530]), 
        .B(_f_permutation__round_in[1210]), .Z(_f_permutation__round__n1023 )
         );
  XOR2_X2 _f_permutation__round__U7227  ( .A(_f_permutation__round__n1025 ), 
        .B(_f_permutation__round__n1024 ), .Z(_f_permutation__round__n2385 )
         );
  XOR2_X2 _f_permutation__round__U7226  ( .A(SYNOPSYS_UNCONNECTED_1029), .B(
        _f_permutation__round__n1026 ), .Z(_f_permutation__round__n1024 ) );
  XOR2_X2 _f_permutation__round__U7225  ( .A(SYNOPSYS_UNCONNECTED_389), .B(
        SYNOPSYS_UNCONNECTED_709), .Z(_f_permutation__round__n1025 ) );
  XOR2_X2 _f_permutation__round__U7224  ( .A(_f_permutation__round_in[1339]), 
        .B(SYNOPSYS_UNCONNECTED_69), .Z(_f_permutation__round__n1026 ) );
  XOR2_X2 _f_permutation__round__U7223  ( .A(_f_permutation__round__n2141 ), 
        .B(_f_permutation__round__n2385 ), .Z(_f_permutation__round__n2142 )
         );
  XOR2_X2 _f_permutation__round__U7222  ( .A(_f_permutation__round_in[1595]), 
        .B(_f_permutation__round__n2142 ), .Z(_f_permutation__round__c[59] )
         );
  XOR2_X2 _f_permutation__round__U7221  ( .A(_f_permutation__round__n1028 ), 
        .B(_f_permutation__round__n1027 ), .Z(_f_permutation__round__n1940 )
         );
  XOR2_X2 _f_permutation__round__U7220  ( .A(SYNOPSYS_UNCONNECTED_773), .B(
        _f_permutation__round__n1029 ), .Z(_f_permutation__round__n1027 ) );
  XOR2_X2 _f_permutation__round__U7219  ( .A(SYNOPSYS_UNCONNECTED_133), .B(
        SYNOPSYS_UNCONNECTED_453), .Z(_f_permutation__round__n1028 ) );
  XOR2_X2 _f_permutation__round__U7218  ( .A(_f_permutation__round_in[1595]), 
        .B(_f_permutation__round_in[1275]), .Z(_f_permutation__round__n1029 )
         );
  XOR2_X2 _f_permutation__round__U7217  ( .A(_f_permutation__round__n1031 ), 
        .B(_f_permutation__round__n1030 ), .Z(_f_permutation__round__n2128 )
         );
  XOR2_X2 _f_permutation__round__U7216  ( .A(SYNOPSYS_UNCONNECTED_964), .B(
        _f_permutation__round__n1032 ), .Z(_f_permutation__round__n1030 ) );
  XOR2_X2 _f_permutation__round__U7215  ( .A(SYNOPSYS_UNCONNECTED_324), .B(
        SYNOPSYS_UNCONNECTED_644), .Z(_f_permutation__round__n1031 ) );
  XOR2_X2 _f_permutation__round__U7214  ( .A(_f_permutation__round_in[1404]), 
        .B(_f_permutation__round_in[1084]), .Z(_f_permutation__round__n1032 )
         );
  XOR2_X2 _f_permutation__round__U7213  ( .A(_f_permutation__round__n1940 ), 
        .B(_f_permutation__round__n2128 ), .Z(_f_permutation__round__n1941 )
         );
  XOR2_X2 _f_permutation__round__U7212  ( .A(SYNOPSYS_UNCONNECTED_1028), .B(
        _f_permutation__round__n1941 ), .Z(_f_permutation__round__c[1596] ) );
  XOR2_X2 _f_permutation__round__U7211  ( .A(_f_permutation__round__n1034 ), 
        .B(_f_permutation__round__n1033 ), .Z(_f_permutation__round__n2392 )
         );
  XOR2_X2 _f_permutation__round__U7210  ( .A(SYNOPSYS_UNCONNECTED_902), .B(
        _f_permutation__round__n1035 ), .Z(_f_permutation__round__n1033 ) );
  XOR2_X2 _f_permutation__round__U7209  ( .A(SYNOPSYS_UNCONNECTED_262), .B(
        SYNOPSYS_UNCONNECTED_582), .Z(_f_permutation__round__n1034 ) );
  XOR2_X2 _f_permutation__round__U7208  ( .A(_f_permutation__round_in[1466]), 
        .B(_f_permutation__round_in[1146]), .Z(_f_permutation__round__n1035 )
         );
  XOR2_X2 _f_permutation__round__U7207  ( .A(_f_permutation__round__n1940 ), 
        .B(_f_permutation__round__n2392 ), .Z(_f_permutation__round__n1942 )
         );
  XOR2_X2 _f_permutation__round__U7206  ( .A(SYNOPSYS_UNCONNECTED_837), .B(
        _f_permutation__round__n1942 ), .Z(_f_permutation__round__c[635] ) );
  XOR2_X2 _f_permutation__round__U7205  ( .A(SYNOPSYS_UNCONNECTED_708), .B(
        _f_permutation__round__n1941 ), .Z(_f_permutation__round__c[1532] ) );
  XOR2_X2 _f_permutation__round__U7204  ( .A(SYNOPSYS_UNCONNECTED_517), .B(
        _f_permutation__round__n1942 ), .Z(_f_permutation__round__c[571] ) );
  XOR2_X2 _f_permutation__round__U7203  ( .A(SYNOPSYS_UNCONNECTED_388), .B(
        _f_permutation__round__n1941 ), .Z(_f_permutation__round__c[1468] ) );
  XOR2_X2 _f_permutation__round__U7202  ( .A(SYNOPSYS_UNCONNECTED_197), .B(
        _f_permutation__round__n1942 ), .Z(_f_permutation__round__c[507] ) );
  XOR2_X2 _f_permutation__round__U7201  ( .A(SYNOPSYS_UNCONNECTED_68), .B(
        _f_permutation__round__n1941 ), .Z(_f_permutation__round__c[1404] ) );
  XOR2_X2 _f_permutation__round__U7200  ( .A(_f_permutation__round_in[1211]), 
        .B(_f_permutation__round__n1942 ), .Z(_f_permutation__round__c[443] )
         );
  XOR2_X2 _f_permutation__round__U7199  ( .A(_f_permutation__round_in[1340]), 
        .B(_f_permutation__round__n1941 ), .Z(_f_permutation__round__c[1340] )
         );
  XOR2_X2 _f_permutation__round__U7198  ( .A(_f_permutation__round_in[1531]), 
        .B(_f_permutation__round__n1942 ), .Z(_f_permutation__round__c[379] )
         );
  XOR2_X2 _f_permutation__round__U7197  ( .A(_f_permutation__round__n1037 ), 
        .B(_f_permutation__round__n1036 ), .Z(_f_permutation__round__n2145 )
         );
  XOR2_X2 _f_permutation__round__U7196  ( .A(SYNOPSYS_UNCONNECTED_839), .B(
        _f_permutation__round__n1038 ), .Z(_f_permutation__round__n1036 ) );
  XOR2_X2 _f_permutation__round__U7195  ( .A(SYNOPSYS_UNCONNECTED_199), .B(
        SYNOPSYS_UNCONNECTED_519), .Z(_f_permutation__round__n1037 ) );
  XOR2_X2 _f_permutation__round__U7194  ( .A(_f_permutation__round_in[1529]), 
        .B(_f_permutation__round_in[1209]), .Z(_f_permutation__round__n1038 )
         );
  XOR2_X2 _f_permutation__round__U7193  ( .A(_f_permutation__round__n1040 ), 
        .B(_f_permutation__round__n1039 ), .Z(_f_permutation__round__n2388 )
         );
  XOR2_X2 _f_permutation__round__U7192  ( .A(SYNOPSYS_UNCONNECTED_1030), .B(
        _f_permutation__round__n1041 ), .Z(_f_permutation__round__n1039 ) );
  XOR2_X2 _f_permutation__round__U7191  ( .A(SYNOPSYS_UNCONNECTED_390), .B(
        SYNOPSYS_UNCONNECTED_710), .Z(_f_permutation__round__n1040 ) );
  XOR2_X2 _f_permutation__round__U7190  ( .A(_f_permutation__round_in[1338]), 
        .B(SYNOPSYS_UNCONNECTED_70), .Z(_f_permutation__round__n1041 ) );
  XOR2_X2 _f_permutation__round__U7189  ( .A(_f_permutation__round__n2145 ), 
        .B(_f_permutation__round__n2388 ), .Z(_f_permutation__round__n2146 )
         );
  XOR2_X2 _f_permutation__round__U7188  ( .A(_f_permutation__round_in[1594]), 
        .B(_f_permutation__round__n2146 ), .Z(_f_permutation__round__c[58] )
         );
  XOR2_X2 _f_permutation__round__U7187  ( .A(_f_permutation__round__n1043 ), 
        .B(_f_permutation__round__n1042 ), .Z(_f_permutation__round__n1943 )
         );
  XOR2_X2 _f_permutation__round__U7186  ( .A(SYNOPSYS_UNCONNECTED_774), .B(
        _f_permutation__round__n1044 ), .Z(_f_permutation__round__n1042 ) );
  XOR2_X2 _f_permutation__round__U7185  ( .A(SYNOPSYS_UNCONNECTED_134), .B(
        SYNOPSYS_UNCONNECTED_454), .Z(_f_permutation__round__n1043 ) );
  XOR2_X2 _f_permutation__round__U7184  ( .A(_f_permutation__round_in[1594]), 
        .B(_f_permutation__round_in[1274]), .Z(_f_permutation__round__n1044 )
         );
  XOR2_X2 _f_permutation__round__U7183  ( .A(_f_permutation__round__n1046 ), 
        .B(_f_permutation__round__n1045 ), .Z(_f_permutation__round__n2132 )
         );
  XOR2_X2 _f_permutation__round__U7182  ( .A(SYNOPSYS_UNCONNECTED_965), .B(
        _f_permutation__round__n1047 ), .Z(_f_permutation__round__n1045 ) );
  XOR2_X2 _f_permutation__round__U7181  ( .A(SYNOPSYS_UNCONNECTED_325), .B(
        SYNOPSYS_UNCONNECTED_645), .Z(_f_permutation__round__n1046 ) );
  XOR2_X2 _f_permutation__round__U7180  ( .A(_f_permutation__round_in[1403]), 
        .B(_f_permutation__round_in[1083]), .Z(_f_permutation__round__n1047 )
         );
  XOR2_X2 _f_permutation__round__U7179  ( .A(_f_permutation__round__n1943 ), 
        .B(_f_permutation__round__n2132 ), .Z(_f_permutation__round__n1944 )
         );
  XOR2_X2 _f_permutation__round__U7178  ( .A(SYNOPSYS_UNCONNECTED_1029), .B(
        _f_permutation__round__n1944 ), .Z(_f_permutation__round__c[1595] ) );
  XOR2_X2 _f_permutation__round__U7177  ( .A(_f_permutation__round__n1049 ), 
        .B(_f_permutation__round__n1048 ), .Z(_f_permutation__round__n2395 )
         );
  XOR2_X2 _f_permutation__round__U7176  ( .A(SYNOPSYS_UNCONNECTED_903), .B(
        _f_permutation__round__n1050 ), .Z(_f_permutation__round__n1048 ) );
  XOR2_X2 _f_permutation__round__U7175  ( .A(SYNOPSYS_UNCONNECTED_263), .B(
        SYNOPSYS_UNCONNECTED_583), .Z(_f_permutation__round__n1049 ) );
  XOR2_X2 _f_permutation__round__U7174  ( .A(_f_permutation__round_in[1465]), 
        .B(_f_permutation__round_in[1145]), .Z(_f_permutation__round__n1050 )
         );
  XOR2_X2 _f_permutation__round__U7173  ( .A(_f_permutation__round__n1943 ), 
        .B(_f_permutation__round__n2395 ), .Z(_f_permutation__round__n1945 )
         );
  XOR2_X2 _f_permutation__round__U7172  ( .A(SYNOPSYS_UNCONNECTED_838), .B(
        _f_permutation__round__n1945 ), .Z(_f_permutation__round__c[634] ) );
  XOR2_X2 _f_permutation__round__U7171  ( .A(SYNOPSYS_UNCONNECTED_709), .B(
        _f_permutation__round__n1944 ), .Z(_f_permutation__round__c[1531] ) );
  XOR2_X2 _f_permutation__round__U7170  ( .A(SYNOPSYS_UNCONNECTED_518), .B(
        _f_permutation__round__n1945 ), .Z(_f_permutation__round__c[570] ) );
  XOR2_X2 _f_permutation__round__U7169  ( .A(SYNOPSYS_UNCONNECTED_389), .B(
        _f_permutation__round__n1944 ), .Z(_f_permutation__round__c[1467] ) );
  XOR2_X2 _f_permutation__round__U7168  ( .A(SYNOPSYS_UNCONNECTED_198), .B(
        _f_permutation__round__n1945 ), .Z(_f_permutation__round__c[506] ) );
  XOR2_X2 _f_permutation__round__U7167  ( .A(SYNOPSYS_UNCONNECTED_69), .B(
        _f_permutation__round__n1944 ), .Z(_f_permutation__round__c[1403] ) );
  XOR2_X2 _f_permutation__round__U7166  ( .A(_f_permutation__round_in[1210]), 
        .B(_f_permutation__round__n1945 ), .Z(_f_permutation__round__c[442] )
         );
  XOR2_X2 _f_permutation__round__U7165  ( .A(_f_permutation__round_in[1339]), 
        .B(_f_permutation__round__n1944 ), .Z(_f_permutation__round__c[1339] )
         );
  XOR2_X2 _f_permutation__round__U7164  ( .A(_f_permutation__round_in[1530]), 
        .B(_f_permutation__round__n1945 ), .Z(_f_permutation__round__c[378] )
         );
  XOR2_X2 _f_permutation__round__U7163  ( .A(_f_permutation__round__n1052 ), 
        .B(_f_permutation__round__n1051 ), .Z(_f_permutation__round__n2149 )
         );
  XOR2_X2 _f_permutation__round__U7162  ( .A(SYNOPSYS_UNCONNECTED_840), .B(
        _f_permutation__round__n1053 ), .Z(_f_permutation__round__n1051 ) );
  XOR2_X2 _f_permutation__round__U7161  ( .A(SYNOPSYS_UNCONNECTED_200), .B(
        SYNOPSYS_UNCONNECTED_520), .Z(_f_permutation__round__n1052 ) );
  XOR2_X2 _f_permutation__round__U7160  ( .A(_f_permutation__round_in[1528]), 
        .B(_f_permutation__round_in[1208]), .Z(_f_permutation__round__n1053 )
         );
  XOR2_X2 _f_permutation__round__U7159  ( .A(_f_permutation__round__n1055 ), 
        .B(_f_permutation__round__n1054 ), .Z(_f_permutation__round__n2391 )
         );
  XOR2_X2 _f_permutation__round__U7158  ( .A(SYNOPSYS_UNCONNECTED_1031), .B(
        _f_permutation__round__n1056 ), .Z(_f_permutation__round__n1054 ) );
  XOR2_X2 _f_permutation__round__U7157  ( .A(SYNOPSYS_UNCONNECTED_391), .B(
        SYNOPSYS_UNCONNECTED_711), .Z(_f_permutation__round__n1055 ) );
  XOR2_X2 _f_permutation__round__U7156  ( .A(_f_permutation__round_in[1337]), 
        .B(SYNOPSYS_UNCONNECTED_71), .Z(_f_permutation__round__n1056 ) );
  XOR2_X2 _f_permutation__round__U7155  ( .A(_f_permutation__round__n2149 ), 
        .B(_f_permutation__round__n2391 ), .Z(_f_permutation__round__n2150 )
         );
  XOR2_X2 _f_permutation__round__U7154  ( .A(_f_permutation__round_in[1593]), 
        .B(_f_permutation__round__n2150 ), .Z(_f_permutation__round__c[57] )
         );
  XOR2_X2 _f_permutation__round__U7153  ( .A(_f_permutation__round__n1058 ), 
        .B(_f_permutation__round__n1057 ), .Z(_f_permutation__round__n1946 )
         );
  XOR2_X2 _f_permutation__round__U7152  ( .A(SYNOPSYS_UNCONNECTED_775), .B(
        _f_permutation__round__n1059 ), .Z(_f_permutation__round__n1057 ) );
  XOR2_X2 _f_permutation__round__U7151  ( .A(SYNOPSYS_UNCONNECTED_135), .B(
        SYNOPSYS_UNCONNECTED_455), .Z(_f_permutation__round__n1058 ) );
  XOR2_X2 _f_permutation__round__U7150  ( .A(_f_permutation__round_in[1593]), 
        .B(_f_permutation__round_in[1273]), .Z(_f_permutation__round__n1059 )
         );
  XOR2_X2 _f_permutation__round__U7149  ( .A(_f_permutation__round__n1061 ), 
        .B(_f_permutation__round__n1060 ), .Z(_f_permutation__round__n2136 )
         );
  XOR2_X2 _f_permutation__round__U7148  ( .A(SYNOPSYS_UNCONNECTED_966), .B(
        _f_permutation__round__n1062 ), .Z(_f_permutation__round__n1060 ) );
  XOR2_X2 _f_permutation__round__U7147  ( .A(SYNOPSYS_UNCONNECTED_326), .B(
        SYNOPSYS_UNCONNECTED_646), .Z(_f_permutation__round__n1061 ) );
  XOR2_X2 _f_permutation__round__U7146  ( .A(_f_permutation__round_in[1402]), 
        .B(_f_permutation__round_in[1082]), .Z(_f_permutation__round__n1062 )
         );
  XOR2_X2 _f_permutation__round__U7145  ( .A(_f_permutation__round__n1946 ), 
        .B(_f_permutation__round__n2136 ), .Z(_f_permutation__round__n1947 )
         );
  XOR2_X2 _f_permutation__round__U7144  ( .A(SYNOPSYS_UNCONNECTED_1030), .B(
        _f_permutation__round__n1947 ), .Z(_f_permutation__round__c[1594] ) );
  XOR2_X2 _f_permutation__round__U7143  ( .A(_f_permutation__round__n1064 ), 
        .B(_f_permutation__round__n1063 ), .Z(_f_permutation__round__n2398 )
         );
  XOR2_X2 _f_permutation__round__U7142  ( .A(SYNOPSYS_UNCONNECTED_904), .B(
        _f_permutation__round__n1065 ), .Z(_f_permutation__round__n1063 ) );
  XOR2_X2 _f_permutation__round__U7141  ( .A(SYNOPSYS_UNCONNECTED_264), .B(
        SYNOPSYS_UNCONNECTED_584), .Z(_f_permutation__round__n1064 ) );
  XOR2_X2 _f_permutation__round__U7140  ( .A(_f_permutation__round_in[1464]), 
        .B(_f_permutation__round_in[1144]), .Z(_f_permutation__round__n1065 )
         );
  XOR2_X2 _f_permutation__round__U7139  ( .A(_f_permutation__round__n1946 ), 
        .B(_f_permutation__round__n2398 ), .Z(_f_permutation__round__n1948 )
         );
  XOR2_X2 _f_permutation__round__U7138  ( .A(SYNOPSYS_UNCONNECTED_839), .B(
        _f_permutation__round__n1948 ), .Z(_f_permutation__round__c[633] ) );
  XOR2_X2 _f_permutation__round__U7137  ( .A(SYNOPSYS_UNCONNECTED_710), .B(
        _f_permutation__round__n1947 ), .Z(_f_permutation__round__c[1530] ) );
  XOR2_X2 _f_permutation__round__U7136  ( .A(SYNOPSYS_UNCONNECTED_519), .B(
        _f_permutation__round__n1948 ), .Z(_f_permutation__round__c[569] ) );
  XOR2_X2 _f_permutation__round__U7135  ( .A(SYNOPSYS_UNCONNECTED_390), .B(
        _f_permutation__round__n1947 ), .Z(_f_permutation__round__c[1466] ) );
  XOR2_X2 _f_permutation__round__U7134  ( .A(SYNOPSYS_UNCONNECTED_199), .B(
        _f_permutation__round__n1948 ), .Z(_f_permutation__round__c[505] ) );
  XOR2_X2 _f_permutation__round__U7133  ( .A(SYNOPSYS_UNCONNECTED_70), .B(
        _f_permutation__round__n1947 ), .Z(_f_permutation__round__c[1402] ) );
  XOR2_X2 _f_permutation__round__U7132  ( .A(_f_permutation__round_in[1209]), 
        .B(_f_permutation__round__n1948 ), .Z(_f_permutation__round__c[441] )
         );
  XOR2_X2 _f_permutation__round__U7131  ( .A(_f_permutation__round_in[1338]), 
        .B(_f_permutation__round__n1947 ), .Z(_f_permutation__round__c[1338] )
         );
  XOR2_X2 _f_permutation__round__U7130  ( .A(_f_permutation__round_in[1529]), 
        .B(_f_permutation__round__n1948 ), .Z(_f_permutation__round__c[377] )
         );
  XOR2_X2 _f_permutation__round__U7129  ( .A(_f_permutation__round__n1067 ), 
        .B(_f_permutation__round__n1066 ), .Z(_f_permutation__round__n2153 )
         );
  XOR2_X2 _f_permutation__round__U7128  ( .A(SYNOPSYS_UNCONNECTED_841), .B(
        _f_permutation__round__n1068 ), .Z(_f_permutation__round__n1066 ) );
  XOR2_X2 _f_permutation__round__U7127  ( .A(SYNOPSYS_UNCONNECTED_201), .B(
        SYNOPSYS_UNCONNECTED_521), .Z(_f_permutation__round__n1067 ) );
  XOR2_X2 _f_permutation__round__U7126  ( .A(_f_permutation__round_in[1527]), 
        .B(_f_permutation__round_in[1207]), .Z(_f_permutation__round__n1068 )
         );
  XOR2_X2 _f_permutation__round__U7125  ( .A(_f_permutation__round__n1070 ), 
        .B(_f_permutation__round__n1069 ), .Z(_f_permutation__round__n2394 )
         );
  XOR2_X2 _f_permutation__round__U7124  ( .A(SYNOPSYS_UNCONNECTED_1032), .B(
        _f_permutation__round__n1071 ), .Z(_f_permutation__round__n1069 ) );
  XOR2_X2 _f_permutation__round__U7123  ( .A(SYNOPSYS_UNCONNECTED_392), .B(
        SYNOPSYS_UNCONNECTED_712), .Z(_f_permutation__round__n1070 ) );
  XOR2_X2 _f_permutation__round__U7122  ( .A(_f_permutation__round_in[1336]), 
        .B(SYNOPSYS_UNCONNECTED_72), .Z(_f_permutation__round__n1071 ) );
  XOR2_X2 _f_permutation__round__U7121  ( .A(_f_permutation__round__n2153 ), 
        .B(_f_permutation__round__n2394 ), .Z(_f_permutation__round__n2154 )
         );
  XOR2_X2 _f_permutation__round__U7120  ( .A(_f_permutation__round_in[1592]), 
        .B(_f_permutation__round__n2154 ), .Z(_f_permutation__round__c[56] )
         );
  XOR2_X2 _f_permutation__round__U7119  ( .A(_f_permutation__round__n1073 ), 
        .B(_f_permutation__round__n1072 ), .Z(_f_permutation__round__n1949 )
         );
  XOR2_X2 _f_permutation__round__U7118  ( .A(SYNOPSYS_UNCONNECTED_776), .B(
        _f_permutation__round__n1074 ), .Z(_f_permutation__round__n1072 ) );
  XOR2_X2 _f_permutation__round__U7117  ( .A(SYNOPSYS_UNCONNECTED_136), .B(
        SYNOPSYS_UNCONNECTED_456), .Z(_f_permutation__round__n1073 ) );
  XOR2_X2 _f_permutation__round__U7116  ( .A(_f_permutation__round_in[1592]), 
        .B(_f_permutation__round_in[1272]), .Z(_f_permutation__round__n1074 )
         );
  XOR2_X2 _f_permutation__round__U7115  ( .A(_f_permutation__round__n1076 ), 
        .B(_f_permutation__round__n1075 ), .Z(_f_permutation__round__n2140 )
         );
  XOR2_X2 _f_permutation__round__U7114  ( .A(SYNOPSYS_UNCONNECTED_967), .B(
        _f_permutation__round__n1077 ), .Z(_f_permutation__round__n1075 ) );
  XOR2_X2 _f_permutation__round__U7113  ( .A(SYNOPSYS_UNCONNECTED_327), .B(
        SYNOPSYS_UNCONNECTED_647), .Z(_f_permutation__round__n1076 ) );
  XOR2_X2 _f_permutation__round__U7112  ( .A(_f_permutation__round_in[1401]), 
        .B(_f_permutation__round_in[1081]), .Z(_f_permutation__round__n1077 )
         );
  XOR2_X2 _f_permutation__round__U7111  ( .A(_f_permutation__round__n1949 ), 
        .B(_f_permutation__round__n2140 ), .Z(_f_permutation__round__n1950 )
         );
  XOR2_X2 _f_permutation__round__U7110  ( .A(SYNOPSYS_UNCONNECTED_1031), .B(
        _f_permutation__round__n1950 ), .Z(_f_permutation__round__c[1593] ) );
  XOR2_X2 _f_permutation__round__U7109  ( .A(_f_permutation__round__n1079 ), 
        .B(_f_permutation__round__n1078 ), .Z(_f_permutation__round__n2401 )
         );
  XOR2_X2 _f_permutation__round__U7108  ( .A(SYNOPSYS_UNCONNECTED_905), .B(
        _f_permutation__round__n1080 ), .Z(_f_permutation__round__n1078 ) );
  XOR2_X2 _f_permutation__round__U7107  ( .A(SYNOPSYS_UNCONNECTED_265), .B(
        SYNOPSYS_UNCONNECTED_585), .Z(_f_permutation__round__n1079 ) );
  XOR2_X2 _f_permutation__round__U7106  ( .A(_f_permutation__round_in[1463]), 
        .B(_f_permutation__round_in[1143]), .Z(_f_permutation__round__n1080 )
         );
  XOR2_X2 _f_permutation__round__U7105  ( .A(_f_permutation__round__n1949 ), 
        .B(_f_permutation__round__n2401 ), .Z(_f_permutation__round__n1951 )
         );
  XOR2_X2 _f_permutation__round__U7104  ( .A(SYNOPSYS_UNCONNECTED_840), .B(
        _f_permutation__round__n1951 ), .Z(_f_permutation__round__c[632] ) );
  XOR2_X2 _f_permutation__round__U7103  ( .A(SYNOPSYS_UNCONNECTED_711), .B(
        _f_permutation__round__n1950 ), .Z(_f_permutation__round__c[1529] ) );
  XOR2_X2 _f_permutation__round__U7102  ( .A(SYNOPSYS_UNCONNECTED_520), .B(
        _f_permutation__round__n1951 ), .Z(_f_permutation__round__c[568] ) );
  XOR2_X2 _f_permutation__round__U7101  ( .A(SYNOPSYS_UNCONNECTED_391), .B(
        _f_permutation__round__n1950 ), .Z(_f_permutation__round__c[1465] ) );
  XOR2_X2 _f_permutation__round__U7100  ( .A(SYNOPSYS_UNCONNECTED_200), .B(
        _f_permutation__round__n1951 ), .Z(_f_permutation__round__c[504] ) );
  XOR2_X2 _f_permutation__round__U7099  ( .A(SYNOPSYS_UNCONNECTED_71), .B(
        _f_permutation__round__n1950 ), .Z(_f_permutation__round__c[1401] ) );
  XOR2_X2 _f_permutation__round__U7098  ( .A(_f_permutation__round_in[1208]), 
        .B(_f_permutation__round__n1951 ), .Z(_f_permutation__round__c[440] )
         );
  XOR2_X2 _f_permutation__round__U7097  ( .A(_f_permutation__round_in[1337]), 
        .B(_f_permutation__round__n1950 ), .Z(_f_permutation__round__c[1337] )
         );
  XOR2_X2 _f_permutation__round__U7096  ( .A(_f_permutation__round_in[1528]), 
        .B(_f_permutation__round__n1951 ), .Z(_f_permutation__round__c[376] )
         );
  XOR2_X2 _f_permutation__round__U7095  ( .A(_f_permutation__round__n1082 ), 
        .B(_f_permutation__round__n1081 ), .Z(_f_permutation__round__n2157 )
         );
  XOR2_X2 _f_permutation__round__U7094  ( .A(SYNOPSYS_UNCONNECTED_842), .B(
        _f_permutation__round__n1083 ), .Z(_f_permutation__round__n1081 ) );
  XOR2_X2 _f_permutation__round__U7093  ( .A(SYNOPSYS_UNCONNECTED_202), .B(
        SYNOPSYS_UNCONNECTED_522), .Z(_f_permutation__round__n1082 ) );
  XOR2_X2 _f_permutation__round__U7092  ( .A(_f_permutation__round_in[1526]), 
        .B(_f_permutation__round_in[1206]), .Z(_f_permutation__round__n1083 )
         );
  XOR2_X2 _f_permutation__round__U7091  ( .A(_f_permutation__round__n1085 ), 
        .B(_f_permutation__round__n1084 ), .Z(_f_permutation__round__n2397 )
         );
  XOR2_X2 _f_permutation__round__U7090  ( .A(SYNOPSYS_UNCONNECTED_1033), .B(
        _f_permutation__round__n1086 ), .Z(_f_permutation__round__n1084 ) );
  XOR2_X2 _f_permutation__round__U7089  ( .A(SYNOPSYS_UNCONNECTED_393), .B(
        SYNOPSYS_UNCONNECTED_713), .Z(_f_permutation__round__n1085 ) );
  XOR2_X2 _f_permutation__round__U7088  ( .A(_f_permutation__round_in[1335]), 
        .B(SYNOPSYS_UNCONNECTED_73), .Z(_f_permutation__round__n1086 ) );
  XOR2_X2 _f_permutation__round__U7087  ( .A(_f_permutation__round__n2157 ), 
        .B(_f_permutation__round__n2397 ), .Z(_f_permutation__round__n2158 )
         );
  XOR2_X2 _f_permutation__round__U7086  ( .A(_f_permutation__round_in[1591]), 
        .B(_f_permutation__round__n2158 ), .Z(_f_permutation__round__c[55] )
         );
  XOR2_X2 _f_permutation__round__U7085  ( .A(_f_permutation__round__n1088 ), 
        .B(_f_permutation__round__n1087 ), .Z(_f_permutation__round__n1952 )
         );
  XOR2_X2 _f_permutation__round__U7084  ( .A(SYNOPSYS_UNCONNECTED_777), .B(
        _f_permutation__round__n1089 ), .Z(_f_permutation__round__n1087 ) );
  XOR2_X2 _f_permutation__round__U7083  ( .A(SYNOPSYS_UNCONNECTED_137), .B(
        SYNOPSYS_UNCONNECTED_457), .Z(_f_permutation__round__n1088 ) );
  XOR2_X2 _f_permutation__round__U7082  ( .A(_f_permutation__round_in[1591]), 
        .B(_f_permutation__round_in[1271]), .Z(_f_permutation__round__n1089 )
         );
  XOR2_X2 _f_permutation__round__U7081  ( .A(_f_permutation__round__n1091 ), 
        .B(_f_permutation__round__n1090 ), .Z(_f_permutation__round__n2144 )
         );
  XOR2_X2 _f_permutation__round__U7080  ( .A(SYNOPSYS_UNCONNECTED_968), .B(
        _f_permutation__round__n1092 ), .Z(_f_permutation__round__n1090 ) );
  XOR2_X2 _f_permutation__round__U7079  ( .A(SYNOPSYS_UNCONNECTED_328), .B(
        SYNOPSYS_UNCONNECTED_648), .Z(_f_permutation__round__n1091 ) );
  XOR2_X2 _f_permutation__round__U7078  ( .A(_f_permutation__round_in[1400]), 
        .B(_f_permutation__round_in[1080]), .Z(_f_permutation__round__n1092 )
         );
  XOR2_X2 _f_permutation__round__U7077  ( .A(_f_permutation__round__n1952 ), 
        .B(_f_permutation__round__n2144 ), .Z(_f_permutation__round__n1953 )
         );
  XOR2_X2 _f_permutation__round__U7076  ( .A(SYNOPSYS_UNCONNECTED_1032), .B(
        _f_permutation__round__n1953 ), .Z(_f_permutation__round__c[1592] ) );
  XOR2_X2 _f_permutation__round__U7075  ( .A(_f_permutation__round__n1094 ), 
        .B(_f_permutation__round__n1093 ), .Z(_f_permutation__round__n2404 )
         );
  XOR2_X2 _f_permutation__round__U7074  ( .A(SYNOPSYS_UNCONNECTED_906), .B(
        _f_permutation__round__n1095 ), .Z(_f_permutation__round__n1093 ) );
  XOR2_X2 _f_permutation__round__U7073  ( .A(SYNOPSYS_UNCONNECTED_266), .B(
        SYNOPSYS_UNCONNECTED_586), .Z(_f_permutation__round__n1094 ) );
  XOR2_X2 _f_permutation__round__U7072  ( .A(_f_permutation__round_in[1462]), 
        .B(_f_permutation__round_in[1142]), .Z(_f_permutation__round__n1095 )
         );
  XOR2_X2 _f_permutation__round__U7071  ( .A(_f_permutation__round__n1952 ), 
        .B(_f_permutation__round__n2404 ), .Z(_f_permutation__round__n1954 )
         );
  XOR2_X2 _f_permutation__round__U7070  ( .A(SYNOPSYS_UNCONNECTED_841), .B(
        _f_permutation__round__n1954 ), .Z(_f_permutation__round__c[631] ) );
  XOR2_X2 _f_permutation__round__U7069  ( .A(SYNOPSYS_UNCONNECTED_712), .B(
        _f_permutation__round__n1953 ), .Z(_f_permutation__round__c[1528] ) );
  XOR2_X2 _f_permutation__round__U7068  ( .A(SYNOPSYS_UNCONNECTED_521), .B(
        _f_permutation__round__n1954 ), .Z(_f_permutation__round__c[567] ) );
  XOR2_X2 _f_permutation__round__U7067  ( .A(SYNOPSYS_UNCONNECTED_392), .B(
        _f_permutation__round__n1953 ), .Z(_f_permutation__round__c[1464] ) );
  XOR2_X2 _f_permutation__round__U7066  ( .A(SYNOPSYS_UNCONNECTED_201), .B(
        _f_permutation__round__n1954 ), .Z(_f_permutation__round__c[503] ) );
  XOR2_X2 _f_permutation__round__U7065  ( .A(SYNOPSYS_UNCONNECTED_72), .B(
        _f_permutation__round__n1953 ), .Z(_f_permutation__round__c[1400] ) );
  XOR2_X2 _f_permutation__round__U7064  ( .A(_f_permutation__round_in[1207]), 
        .B(_f_permutation__round__n1954 ), .Z(_f_permutation__round__c[439] )
         );
  XOR2_X2 _f_permutation__round__U7063  ( .A(_f_permutation__round_in[1336]), 
        .B(_f_permutation__round__n1953 ), .Z(_f_permutation__round__c[1336] )
         );
  XOR2_X2 _f_permutation__round__U7062  ( .A(_f_permutation__round_in[1527]), 
        .B(_f_permutation__round__n1954 ), .Z(_f_permutation__round__c[375] )
         );
  XOR2_X2 _f_permutation__round__U7061  ( .A(_f_permutation__round__n1097 ), 
        .B(_f_permutation__round__n1096 ), .Z(_f_permutation__round__n2161 )
         );
  XOR2_X2 _f_permutation__round__U7060  ( .A(SYNOPSYS_UNCONNECTED_843), .B(
        _f_permutation__round__n1098 ), .Z(_f_permutation__round__n1096 ) );
  XOR2_X2 _f_permutation__round__U7059  ( .A(SYNOPSYS_UNCONNECTED_203), .B(
        SYNOPSYS_UNCONNECTED_523), .Z(_f_permutation__round__n1097 ) );
  XOR2_X2 _f_permutation__round__U7058  ( .A(_f_permutation__round_in[1525]), 
        .B(_f_permutation__round_in[1205]), .Z(_f_permutation__round__n1098 )
         );
  XOR2_X2 _f_permutation__round__U7057  ( .A(_f_permutation__round__n1100 ), 
        .B(_f_permutation__round__n1099 ), .Z(_f_permutation__round__n2400 )
         );
  XOR2_X2 _f_permutation__round__U7056  ( .A(SYNOPSYS_UNCONNECTED_1034), .B(
        _f_permutation__round__n1101 ), .Z(_f_permutation__round__n1099 ) );
  XOR2_X2 _f_permutation__round__U7055  ( .A(SYNOPSYS_UNCONNECTED_394), .B(
        SYNOPSYS_UNCONNECTED_714), .Z(_f_permutation__round__n1100 ) );
  XOR2_X2 _f_permutation__round__U7054  ( .A(_f_permutation__round_in[1334]), 
        .B(SYNOPSYS_UNCONNECTED_74), .Z(_f_permutation__round__n1101 ) );
  XOR2_X2 _f_permutation__round__U7053  ( .A(_f_permutation__round__n2161 ), 
        .B(_f_permutation__round__n2400 ), .Z(_f_permutation__round__n2162 )
         );
  XOR2_X2 _f_permutation__round__U7052  ( .A(_f_permutation__round_in[1590]), 
        .B(_f_permutation__round__n2162 ), .Z(_f_permutation__round__c[54] )
         );
  XOR2_X2 _f_permutation__round__U7051  ( .A(_f_permutation__round__n1103 ), 
        .B(_f_permutation__round__n1102 ), .Z(_f_permutation__round__n1955 )
         );
  XOR2_X2 _f_permutation__round__U7050  ( .A(SYNOPSYS_UNCONNECTED_778), .B(
        _f_permutation__round__n1104 ), .Z(_f_permutation__round__n1102 ) );
  XOR2_X2 _f_permutation__round__U7049  ( .A(SYNOPSYS_UNCONNECTED_138), .B(
        SYNOPSYS_UNCONNECTED_458), .Z(_f_permutation__round__n1103 ) );
  XOR2_X2 _f_permutation__round__U7048  ( .A(_f_permutation__round_in[1590]), 
        .B(_f_permutation__round_in[1270]), .Z(_f_permutation__round__n1104 )
         );
  XOR2_X2 _f_permutation__round__U7047  ( .A(_f_permutation__round__n1106 ), 
        .B(_f_permutation__round__n1105 ), .Z(_f_permutation__round__n2148 )
         );
  XOR2_X2 _f_permutation__round__U7046  ( .A(SYNOPSYS_UNCONNECTED_969), .B(
        _f_permutation__round__n1107 ), .Z(_f_permutation__round__n1105 ) );
  XOR2_X2 _f_permutation__round__U7045  ( .A(SYNOPSYS_UNCONNECTED_329), .B(
        SYNOPSYS_UNCONNECTED_649), .Z(_f_permutation__round__n1106 ) );
  XOR2_X2 _f_permutation__round__U7044  ( .A(_f_permutation__round_in[1399]), 
        .B(_f_permutation__round_in[1079]), .Z(_f_permutation__round__n1107 )
         );
  XOR2_X2 _f_permutation__round__U7043  ( .A(_f_permutation__round__n1955 ), 
        .B(_f_permutation__round__n2148 ), .Z(_f_permutation__round__n1956 )
         );
  XOR2_X2 _f_permutation__round__U7042  ( .A(SYNOPSYS_UNCONNECTED_1033), .B(
        _f_permutation__round__n1956 ), .Z(_f_permutation__round__c[1591] ) );
  XOR2_X2 _f_permutation__round__U7041  ( .A(_f_permutation__round__n1109 ), 
        .B(_f_permutation__round__n1108 ), .Z(_f_permutation__round__n2407 )
         );
  XOR2_X2 _f_permutation__round__U7040  ( .A(SYNOPSYS_UNCONNECTED_907), .B(
        _f_permutation__round__n1110 ), .Z(_f_permutation__round__n1108 ) );
  XOR2_X2 _f_permutation__round__U7039  ( .A(SYNOPSYS_UNCONNECTED_267), .B(
        SYNOPSYS_UNCONNECTED_587), .Z(_f_permutation__round__n1109 ) );
  XOR2_X2 _f_permutation__round__U7038  ( .A(_f_permutation__round_in[1461]), 
        .B(_f_permutation__round_in[1141]), .Z(_f_permutation__round__n1110 )
         );
  XOR2_X2 _f_permutation__round__U7037  ( .A(_f_permutation__round__n1955 ), 
        .B(_f_permutation__round__n2407 ), .Z(_f_permutation__round__n1957 )
         );
  XOR2_X2 _f_permutation__round__U7036  ( .A(SYNOPSYS_UNCONNECTED_842), .B(
        _f_permutation__round__n1957 ), .Z(_f_permutation__round__c[630] ) );
  XOR2_X2 _f_permutation__round__U7035  ( .A(SYNOPSYS_UNCONNECTED_713), .B(
        _f_permutation__round__n1956 ), .Z(_f_permutation__round__c[1527] ) );
  XOR2_X2 _f_permutation__round__U7034  ( .A(SYNOPSYS_UNCONNECTED_522), .B(
        _f_permutation__round__n1957 ), .Z(_f_permutation__round__c[566] ) );
  XOR2_X2 _f_permutation__round__U7033  ( .A(SYNOPSYS_UNCONNECTED_393), .B(
        _f_permutation__round__n1956 ), .Z(_f_permutation__round__c[1463] ) );
  XOR2_X2 _f_permutation__round__U7032  ( .A(SYNOPSYS_UNCONNECTED_202), .B(
        _f_permutation__round__n1957 ), .Z(_f_permutation__round__c[502] ) );
  XOR2_X2 _f_permutation__round__U7031  ( .A(SYNOPSYS_UNCONNECTED_73), .B(
        _f_permutation__round__n1956 ), .Z(_f_permutation__round__c[1399] ) );
  XOR2_X2 _f_permutation__round__U7030  ( .A(_f_permutation__round_in[1206]), 
        .B(_f_permutation__round__n1957 ), .Z(_f_permutation__round__c[438] )
         );
  XOR2_X2 _f_permutation__round__U7029  ( .A(_f_permutation__round_in[1335]), 
        .B(_f_permutation__round__n1956 ), .Z(_f_permutation__round__c[1335] )
         );
  XOR2_X2 _f_permutation__round__U7028  ( .A(_f_permutation__round_in[1526]), 
        .B(_f_permutation__round__n1957 ), .Z(_f_permutation__round__c[374] )
         );
  XOR2_X2 _f_permutation__round__U7027  ( .A(_f_permutation__round__n1112 ), 
        .B(_f_permutation__round__n1111 ), .Z(_f_permutation__round__n2165 )
         );
  XOR2_X2 _f_permutation__round__U7026  ( .A(SYNOPSYS_UNCONNECTED_844), .B(
        _f_permutation__round__n1113 ), .Z(_f_permutation__round__n1111 ) );
  XOR2_X2 _f_permutation__round__U7025  ( .A(SYNOPSYS_UNCONNECTED_204), .B(
        SYNOPSYS_UNCONNECTED_524), .Z(_f_permutation__round__n1112 ) );
  XOR2_X2 _f_permutation__round__U7024  ( .A(_f_permutation__round_in[1524]), 
        .B(_f_permutation__round_in[1204]), .Z(_f_permutation__round__n1113 )
         );
  XOR2_X2 _f_permutation__round__U7023  ( .A(_f_permutation__round__n1115 ), 
        .B(_f_permutation__round__n1114 ), .Z(_f_permutation__round__n2403 )
         );
  XOR2_X2 _f_permutation__round__U7022  ( .A(SYNOPSYS_UNCONNECTED_1035), .B(
        _f_permutation__round__n1116 ), .Z(_f_permutation__round__n1114 ) );
  XOR2_X2 _f_permutation__round__U7021  ( .A(SYNOPSYS_UNCONNECTED_395), .B(
        SYNOPSYS_UNCONNECTED_715), .Z(_f_permutation__round__n1115 ) );
  XOR2_X2 _f_permutation__round__U7020  ( .A(_f_permutation__round_in[1333]), 
        .B(SYNOPSYS_UNCONNECTED_75), .Z(_f_permutation__round__n1116 ) );
  XOR2_X2 _f_permutation__round__U7019  ( .A(_f_permutation__round__n2165 ), 
        .B(_f_permutation__round__n2403 ), .Z(_f_permutation__round__n2166 )
         );
  XOR2_X2 _f_permutation__round__U7018  ( .A(_f_permutation__round_in[1589]), 
        .B(_f_permutation__round__n2166 ), .Z(_f_permutation__round__c[53] )
         );
  XOR2_X2 _f_permutation__round__U7017  ( .A(_f_permutation__round__n1118 ), 
        .B(_f_permutation__round__n1117 ), .Z(_f_permutation__round__n1958 )
         );
  XOR2_X2 _f_permutation__round__U7016  ( .A(SYNOPSYS_UNCONNECTED_779), .B(
        _f_permutation__round__n1119 ), .Z(_f_permutation__round__n1117 ) );
  XOR2_X2 _f_permutation__round__U7015  ( .A(SYNOPSYS_UNCONNECTED_139), .B(
        SYNOPSYS_UNCONNECTED_459), .Z(_f_permutation__round__n1118 ) );
  XOR2_X2 _f_permutation__round__U7014  ( .A(_f_permutation__round_in[1589]), 
        .B(_f_permutation__round_in[1269]), .Z(_f_permutation__round__n1119 )
         );
  XOR2_X2 _f_permutation__round__U7013  ( .A(_f_permutation__round__n1121 ), 
        .B(_f_permutation__round__n1120 ), .Z(_f_permutation__round__n2152 )
         );
  XOR2_X2 _f_permutation__round__U7012  ( .A(SYNOPSYS_UNCONNECTED_970), .B(
        _f_permutation__round__n1122 ), .Z(_f_permutation__round__n1120 ) );
  XOR2_X2 _f_permutation__round__U7011  ( .A(SYNOPSYS_UNCONNECTED_330), .B(
        SYNOPSYS_UNCONNECTED_650), .Z(_f_permutation__round__n1121 ) );
  XOR2_X2 _f_permutation__round__U7010  ( .A(_f_permutation__round_in[1398]), 
        .B(_f_permutation__round_in[1078]), .Z(_f_permutation__round__n1122 )
         );
  XOR2_X2 _f_permutation__round__U7009  ( .A(_f_permutation__round__n1958 ), 
        .B(_f_permutation__round__n2152 ), .Z(_f_permutation__round__n1959 )
         );
  XOR2_X2 _f_permutation__round__U7008  ( .A(SYNOPSYS_UNCONNECTED_1034), .B(
        _f_permutation__round__n1959 ), .Z(_f_permutation__round__c[1590] ) );
  XOR2_X2 _f_permutation__round__U7007  ( .A(_f_permutation__round__n1124 ), 
        .B(_f_permutation__round__n1123 ), .Z(_f_permutation__round__n2410 )
         );
  XOR2_X2 _f_permutation__round__U7006  ( .A(SYNOPSYS_UNCONNECTED_908), .B(
        _f_permutation__round__n1125 ), .Z(_f_permutation__round__n1123 ) );
  XOR2_X2 _f_permutation__round__U7005  ( .A(SYNOPSYS_UNCONNECTED_268), .B(
        SYNOPSYS_UNCONNECTED_588), .Z(_f_permutation__round__n1124 ) );
  XOR2_X2 _f_permutation__round__U7004  ( .A(_f_permutation__round_in[1460]), 
        .B(_f_permutation__round_in[1140]), .Z(_f_permutation__round__n1125 )
         );
  XOR2_X2 _f_permutation__round__U7003  ( .A(_f_permutation__round__n1958 ), 
        .B(_f_permutation__round__n2410 ), .Z(_f_permutation__round__n1960 )
         );
  XOR2_X2 _f_permutation__round__U7002  ( .A(SYNOPSYS_UNCONNECTED_843), .B(
        _f_permutation__round__n1960 ), .Z(_f_permutation__round__c[629] ) );
  XOR2_X2 _f_permutation__round__U7001  ( .A(SYNOPSYS_UNCONNECTED_714), .B(
        _f_permutation__round__n1959 ), .Z(_f_permutation__round__c[1526] ) );
  XOR2_X2 _f_permutation__round__U7000  ( .A(SYNOPSYS_UNCONNECTED_523), .B(
        _f_permutation__round__n1960 ), .Z(_f_permutation__round__c[565] ) );
  XOR2_X2 _f_permutation__round__U6999  ( .A(SYNOPSYS_UNCONNECTED_394), .B(
        _f_permutation__round__n1959 ), .Z(_f_permutation__round__c[1462] ) );
  XOR2_X2 _f_permutation__round__U6998  ( .A(SYNOPSYS_UNCONNECTED_203), .B(
        _f_permutation__round__n1960 ), .Z(_f_permutation__round__c[501] ) );
  XOR2_X2 _f_permutation__round__U6997  ( .A(SYNOPSYS_UNCONNECTED_74), .B(
        _f_permutation__round__n1959 ), .Z(_f_permutation__round__c[1398] ) );
  XOR2_X2 _f_permutation__round__U6996  ( .A(_f_permutation__round_in[1205]), 
        .B(_f_permutation__round__n1960 ), .Z(_f_permutation__round__c[437] )
         );
  XOR2_X2 _f_permutation__round__U6995  ( .A(_f_permutation__round_in[1334]), 
        .B(_f_permutation__round__n1959 ), .Z(_f_permutation__round__c[1334] )
         );
  XOR2_X2 _f_permutation__round__U6994  ( .A(_f_permutation__round_in[1525]), 
        .B(_f_permutation__round__n1960 ), .Z(_f_permutation__round__c[373] )
         );
  XOR2_X2 _f_permutation__round__U6993  ( .A(_f_permutation__round__n1127 ), 
        .B(_f_permutation__round__n1126 ), .Z(_f_permutation__round__n2169 )
         );
  XOR2_X2 _f_permutation__round__U6992  ( .A(SYNOPSYS_UNCONNECTED_845), .B(
        _f_permutation__round__n1128 ), .Z(_f_permutation__round__n1126 ) );
  XOR2_X2 _f_permutation__round__U6991  ( .A(SYNOPSYS_UNCONNECTED_205), .B(
        SYNOPSYS_UNCONNECTED_525), .Z(_f_permutation__round__n1127 ) );
  XOR2_X2 _f_permutation__round__U6990  ( .A(_f_permutation__round_in[1523]), 
        .B(_f_permutation__round_in[1203]), .Z(_f_permutation__round__n1128 )
         );
  XOR2_X2 _f_permutation__round__U6989  ( .A(_f_permutation__round__n1130 ), 
        .B(_f_permutation__round__n1129 ), .Z(_f_permutation__round__n2406 )
         );
  XOR2_X2 _f_permutation__round__U6988  ( .A(SYNOPSYS_UNCONNECTED_1036), .B(
        _f_permutation__round__n1131 ), .Z(_f_permutation__round__n1129 ) );
  XOR2_X2 _f_permutation__round__U6987  ( .A(SYNOPSYS_UNCONNECTED_396), .B(
        SYNOPSYS_UNCONNECTED_716), .Z(_f_permutation__round__n1130 ) );
  XOR2_X2 _f_permutation__round__U6986  ( .A(_f_permutation__round_in[1332]), 
        .B(SYNOPSYS_UNCONNECTED_76), .Z(_f_permutation__round__n1131 ) );
  XOR2_X2 _f_permutation__round__U6985  ( .A(_f_permutation__round__n2169 ), 
        .B(_f_permutation__round__n2406 ), .Z(_f_permutation__round__n2170 )
         );
  XOR2_X2 _f_permutation__round__U6984  ( .A(_f_permutation__round_in[1588]), 
        .B(_f_permutation__round__n2170 ), .Z(_f_permutation__round__c[52] )
         );
  XOR2_X2 _f_permutation__round__U6983  ( .A(_f_permutation__round__n1133 ), 
        .B(_f_permutation__round__n1132 ), .Z(_f_permutation__round__n1961 )
         );
  XOR2_X2 _f_permutation__round__U6982  ( .A(SYNOPSYS_UNCONNECTED_780), .B(
        _f_permutation__round__n1134 ), .Z(_f_permutation__round__n1132 ) );
  XOR2_X2 _f_permutation__round__U6981  ( .A(SYNOPSYS_UNCONNECTED_140), .B(
        SYNOPSYS_UNCONNECTED_460), .Z(_f_permutation__round__n1133 ) );
  XOR2_X2 _f_permutation__round__U6980  ( .A(_f_permutation__round_in[1588]), 
        .B(_f_permutation__round_in[1268]), .Z(_f_permutation__round__n1134 )
         );
  XOR2_X2 _f_permutation__round__U6979  ( .A(_f_permutation__round__n1136 ), 
        .B(_f_permutation__round__n1135 ), .Z(_f_permutation__round__n2156 )
         );
  XOR2_X2 _f_permutation__round__U6978  ( .A(SYNOPSYS_UNCONNECTED_971), .B(
        _f_permutation__round__n1137 ), .Z(_f_permutation__round__n1135 ) );
  XOR2_X2 _f_permutation__round__U6977  ( .A(SYNOPSYS_UNCONNECTED_331), .B(
        SYNOPSYS_UNCONNECTED_651), .Z(_f_permutation__round__n1136 ) );
  XOR2_X2 _f_permutation__round__U6976  ( .A(_f_permutation__round_in[1397]), 
        .B(_f_permutation__round_in[1077]), .Z(_f_permutation__round__n1137 )
         );
  XOR2_X2 _f_permutation__round__U6975  ( .A(_f_permutation__round__n1961 ), 
        .B(_f_permutation__round__n2156 ), .Z(_f_permutation__round__n1962 )
         );
  XOR2_X2 _f_permutation__round__U6974  ( .A(SYNOPSYS_UNCONNECTED_1035), .B(
        _f_permutation__round__n1962 ), .Z(_f_permutation__round__c[1589] ) );
  XOR2_X2 _f_permutation__round__U6973  ( .A(_f_permutation__round__n1139 ), 
        .B(_f_permutation__round__n1138 ), .Z(_f_permutation__round__n2413 )
         );
  XOR2_X2 _f_permutation__round__U6972  ( .A(SYNOPSYS_UNCONNECTED_909), .B(
        _f_permutation__round__n1140 ), .Z(_f_permutation__round__n1138 ) );
  XOR2_X2 _f_permutation__round__U6971  ( .A(SYNOPSYS_UNCONNECTED_269), .B(
        SYNOPSYS_UNCONNECTED_589), .Z(_f_permutation__round__n1139 ) );
  XOR2_X2 _f_permutation__round__U6970  ( .A(_f_permutation__round_in[1459]), 
        .B(_f_permutation__round_in[1139]), .Z(_f_permutation__round__n1140 )
         );
  XOR2_X2 _f_permutation__round__U6969  ( .A(_f_permutation__round__n1961 ), 
        .B(_f_permutation__round__n2413 ), .Z(_f_permutation__round__n1963 )
         );
  XOR2_X2 _f_permutation__round__U6968  ( .A(SYNOPSYS_UNCONNECTED_844), .B(
        _f_permutation__round__n1963 ), .Z(_f_permutation__round__c[628] ) );
  XOR2_X2 _f_permutation__round__U6967  ( .A(SYNOPSYS_UNCONNECTED_715), .B(
        _f_permutation__round__n1962 ), .Z(_f_permutation__round__c[1525] ) );
  XOR2_X2 _f_permutation__round__U6966  ( .A(SYNOPSYS_UNCONNECTED_524), .B(
        _f_permutation__round__n1963 ), .Z(_f_permutation__round__c[564] ) );
  XOR2_X2 _f_permutation__round__U6965  ( .A(SYNOPSYS_UNCONNECTED_395), .B(
        _f_permutation__round__n1962 ), .Z(_f_permutation__round__c[1461] ) );
  XOR2_X2 _f_permutation__round__U6964  ( .A(SYNOPSYS_UNCONNECTED_204), .B(
        _f_permutation__round__n1963 ), .Z(_f_permutation__round__c[500] ) );
  XOR2_X2 _f_permutation__round__U6963  ( .A(SYNOPSYS_UNCONNECTED_75), .B(
        _f_permutation__round__n1962 ), .Z(_f_permutation__round__c[1397] ) );
  XOR2_X2 _f_permutation__round__U6962  ( .A(_f_permutation__round_in[1204]), 
        .B(_f_permutation__round__n1963 ), .Z(_f_permutation__round__c[436] )
         );
  XOR2_X2 _f_permutation__round__U6961  ( .A(_f_permutation__round_in[1333]), 
        .B(_f_permutation__round__n1962 ), .Z(_f_permutation__round__c[1333] )
         );
  XOR2_X2 _f_permutation__round__U6960  ( .A(_f_permutation__round_in[1524]), 
        .B(_f_permutation__round__n1963 ), .Z(_f_permutation__round__c[372] )
         );
  XOR2_X2 _f_permutation__round__U6959  ( .A(_f_permutation__round__n1142 ), 
        .B(_f_permutation__round__n1141 ), .Z(_f_permutation__round__n2173 )
         );
  XOR2_X2 _f_permutation__round__U6958  ( .A(SYNOPSYS_UNCONNECTED_846), .B(
        _f_permutation__round__n1143 ), .Z(_f_permutation__round__n1141 ) );
  XOR2_X2 _f_permutation__round__U6957  ( .A(SYNOPSYS_UNCONNECTED_206), .B(
        SYNOPSYS_UNCONNECTED_526), .Z(_f_permutation__round__n1142 ) );
  XOR2_X2 _f_permutation__round__U6956  ( .A(_f_permutation__round_in[1522]), 
        .B(_f_permutation__round_in[1202]), .Z(_f_permutation__round__n1143 )
         );
  XOR2_X2 _f_permutation__round__U6955  ( .A(_f_permutation__round__n1145 ), 
        .B(_f_permutation__round__n1144 ), .Z(_f_permutation__round__n2409 )
         );
  XOR2_X2 _f_permutation__round__U6954  ( .A(SYNOPSYS_UNCONNECTED_1037), .B(
        _f_permutation__round__n1146 ), .Z(_f_permutation__round__n1144 ) );
  XOR2_X2 _f_permutation__round__U6953  ( .A(SYNOPSYS_UNCONNECTED_397), .B(
        SYNOPSYS_UNCONNECTED_717), .Z(_f_permutation__round__n1145 ) );
  XOR2_X2 _f_permutation__round__U6952  ( .A(_f_permutation__round_in[1331]), 
        .B(SYNOPSYS_UNCONNECTED_77), .Z(_f_permutation__round__n1146 ) );
  XOR2_X2 _f_permutation__round__U6951  ( .A(_f_permutation__round__n2173 ), 
        .B(_f_permutation__round__n2409 ), .Z(_f_permutation__round__n2174 )
         );
  XOR2_X2 _f_permutation__round__U6950  ( .A(_f_permutation__round_in[1587]), 
        .B(_f_permutation__round__n2174 ), .Z(_f_permutation__round__c[51] )
         );
  XOR2_X2 _f_permutation__round__U6949  ( .A(_f_permutation__round__n1148 ), 
        .B(_f_permutation__round__n1147 ), .Z(_f_permutation__round__n1964 )
         );
  XOR2_X2 _f_permutation__round__U6948  ( .A(SYNOPSYS_UNCONNECTED_781), .B(
        _f_permutation__round__n1149 ), .Z(_f_permutation__round__n1147 ) );
  XOR2_X2 _f_permutation__round__U6947  ( .A(SYNOPSYS_UNCONNECTED_141), .B(
        SYNOPSYS_UNCONNECTED_461), .Z(_f_permutation__round__n1148 ) );
  XOR2_X2 _f_permutation__round__U6946  ( .A(_f_permutation__round_in[1587]), 
        .B(_f_permutation__round_in[1267]), .Z(_f_permutation__round__n1149 )
         );
  XOR2_X2 _f_permutation__round__U6945  ( .A(_f_permutation__round__n1151 ), 
        .B(_f_permutation__round__n1150 ), .Z(_f_permutation__round__n2160 )
         );
  XOR2_X2 _f_permutation__round__U6944  ( .A(SYNOPSYS_UNCONNECTED_972), .B(
        _f_permutation__round__n1152 ), .Z(_f_permutation__round__n1150 ) );
  XOR2_X2 _f_permutation__round__U6943  ( .A(SYNOPSYS_UNCONNECTED_332), .B(
        SYNOPSYS_UNCONNECTED_652), .Z(_f_permutation__round__n1151 ) );
  XOR2_X2 _f_permutation__round__U6942  ( .A(_f_permutation__round_in[1396]), 
        .B(_f_permutation__round_in[1076]), .Z(_f_permutation__round__n1152 )
         );
  XOR2_X2 _f_permutation__round__U6941  ( .A(_f_permutation__round__n1964 ), 
        .B(_f_permutation__round__n2160 ), .Z(_f_permutation__round__n1965 )
         );
  XOR2_X2 _f_permutation__round__U6940  ( .A(SYNOPSYS_UNCONNECTED_1036), .B(
        _f_permutation__round__n1965 ), .Z(_f_permutation__round__c[1588] ) );
  XOR2_X2 _f_permutation__round__U6939  ( .A(_f_permutation__round__n1154 ), 
        .B(_f_permutation__round__n1153 ), .Z(_f_permutation__round__n2416 )
         );
  XOR2_X2 _f_permutation__round__U6938  ( .A(SYNOPSYS_UNCONNECTED_910), .B(
        _f_permutation__round__n1155 ), .Z(_f_permutation__round__n1153 ) );
  XOR2_X2 _f_permutation__round__U6937  ( .A(SYNOPSYS_UNCONNECTED_270), .B(
        SYNOPSYS_UNCONNECTED_590), .Z(_f_permutation__round__n1154 ) );
  XOR2_X2 _f_permutation__round__U6936  ( .A(_f_permutation__round_in[1458]), 
        .B(_f_permutation__round_in[1138]), .Z(_f_permutation__round__n1155 )
         );
  XOR2_X2 _f_permutation__round__U6935  ( .A(_f_permutation__round__n1964 ), 
        .B(_f_permutation__round__n2416 ), .Z(_f_permutation__round__n1966 )
         );
  XOR2_X2 _f_permutation__round__U6934  ( .A(SYNOPSYS_UNCONNECTED_845), .B(
        _f_permutation__round__n1966 ), .Z(_f_permutation__round__c[627] ) );
  XOR2_X2 _f_permutation__round__U6933  ( .A(SYNOPSYS_UNCONNECTED_716), .B(
        _f_permutation__round__n1965 ), .Z(_f_permutation__round__c[1524] ) );
  XOR2_X2 _f_permutation__round__U6932  ( .A(SYNOPSYS_UNCONNECTED_525), .B(
        _f_permutation__round__n1966 ), .Z(_f_permutation__round__c[563] ) );
  XOR2_X2 _f_permutation__round__U6931  ( .A(SYNOPSYS_UNCONNECTED_396), .B(
        _f_permutation__round__n1965 ), .Z(_f_permutation__round__c[1460] ) );
  XOR2_X2 _f_permutation__round__U6930  ( .A(SYNOPSYS_UNCONNECTED_205), .B(
        _f_permutation__round__n1966 ), .Z(_f_permutation__round__c[499] ) );
  XOR2_X2 _f_permutation__round__U6929  ( .A(SYNOPSYS_UNCONNECTED_76), .B(
        _f_permutation__round__n1965 ), .Z(_f_permutation__round__c[1396] ) );
  XOR2_X2 _f_permutation__round__U6928  ( .A(_f_permutation__round_in[1203]), 
        .B(_f_permutation__round__n1966 ), .Z(_f_permutation__round__c[435] )
         );
  XOR2_X2 _f_permutation__round__U6927  ( .A(_f_permutation__round_in[1332]), 
        .B(_f_permutation__round__n1965 ), .Z(_f_permutation__round__c[1332] )
         );
  XOR2_X2 _f_permutation__round__U6926  ( .A(_f_permutation__round_in[1523]), 
        .B(_f_permutation__round__n1966 ), .Z(_f_permutation__round__c[371] )
         );
  XOR2_X2 _f_permutation__round__U6925  ( .A(_f_permutation__round__n1157 ), 
        .B(_f_permutation__round__n1156 ), .Z(_f_permutation__round__n2177 )
         );
  XOR2_X2 _f_permutation__round__U6924  ( .A(SYNOPSYS_UNCONNECTED_847), .B(
        _f_permutation__round__n1158 ), .Z(_f_permutation__round__n1156 ) );
  XOR2_X2 _f_permutation__round__U6923  ( .A(SYNOPSYS_UNCONNECTED_207), .B(
        SYNOPSYS_UNCONNECTED_527), .Z(_f_permutation__round__n1157 ) );
  XOR2_X2 _f_permutation__round__U6922  ( .A(_f_permutation__round_in[1521]), 
        .B(_f_permutation__round_in[1201]), .Z(_f_permutation__round__n1158 )
         );
  XOR2_X2 _f_permutation__round__U6921  ( .A(_f_permutation__round__n1160 ), 
        .B(_f_permutation__round__n1159 ), .Z(_f_permutation__round__n2412 )
         );
  XOR2_X2 _f_permutation__round__U6920  ( .A(SYNOPSYS_UNCONNECTED_1038), .B(
        _f_permutation__round__n1161 ), .Z(_f_permutation__round__n1159 ) );
  XOR2_X2 _f_permutation__round__U6919  ( .A(SYNOPSYS_UNCONNECTED_398), .B(
        SYNOPSYS_UNCONNECTED_718), .Z(_f_permutation__round__n1160 ) );
  XOR2_X2 _f_permutation__round__U6918  ( .A(_f_permutation__round_in[1330]), 
        .B(SYNOPSYS_UNCONNECTED_78), .Z(_f_permutation__round__n1161 ) );
  XOR2_X2 _f_permutation__round__U6917  ( .A(_f_permutation__round__n2177 ), 
        .B(_f_permutation__round__n2412 ), .Z(_f_permutation__round__n2178 )
         );
  XOR2_X2 _f_permutation__round__U6916  ( .A(_f_permutation__round_in[1586]), 
        .B(_f_permutation__round__n2178 ), .Z(_f_permutation__round__c[50] )
         );
  XOR2_X2 _f_permutation__round__U6915  ( .A(_f_permutation__round__n1163 ), 
        .B(_f_permutation__round__n1162 ), .Z(_f_permutation__round__n1967 )
         );
  XOR2_X2 _f_permutation__round__U6914  ( .A(SYNOPSYS_UNCONNECTED_782), .B(
        _f_permutation__round__n1164 ), .Z(_f_permutation__round__n1162 ) );
  XOR2_X2 _f_permutation__round__U6913  ( .A(SYNOPSYS_UNCONNECTED_142), .B(
        SYNOPSYS_UNCONNECTED_462), .Z(_f_permutation__round__n1163 ) );
  XOR2_X2 _f_permutation__round__U6912  ( .A(_f_permutation__round_in[1586]), 
        .B(_f_permutation__round_in[1266]), .Z(_f_permutation__round__n1164 )
         );
  XOR2_X2 _f_permutation__round__U6911  ( .A(_f_permutation__round__n1166 ), 
        .B(_f_permutation__round__n1165 ), .Z(_f_permutation__round__n2164 )
         );
  XOR2_X2 _f_permutation__round__U6910  ( .A(SYNOPSYS_UNCONNECTED_973), .B(
        _f_permutation__round__n1167 ), .Z(_f_permutation__round__n1165 ) );
  XOR2_X2 _f_permutation__round__U6909  ( .A(SYNOPSYS_UNCONNECTED_333), .B(
        SYNOPSYS_UNCONNECTED_653), .Z(_f_permutation__round__n1166 ) );
  XOR2_X2 _f_permutation__round__U6908  ( .A(_f_permutation__round_in[1395]), 
        .B(_f_permutation__round_in[1075]), .Z(_f_permutation__round__n1167 )
         );
  XOR2_X2 _f_permutation__round__U6907  ( .A(_f_permutation__round__n1967 ), 
        .B(_f_permutation__round__n2164 ), .Z(_f_permutation__round__n1968 )
         );
  XOR2_X2 _f_permutation__round__U6906  ( .A(SYNOPSYS_UNCONNECTED_1037), .B(
        _f_permutation__round__n1968 ), .Z(_f_permutation__round__c[1587] ) );
  XOR2_X2 _f_permutation__round__U6905  ( .A(_f_permutation__round__n1169 ), 
        .B(_f_permutation__round__n1168 ), .Z(_f_permutation__round__n2419 )
         );
  XOR2_X2 _f_permutation__round__U6904  ( .A(SYNOPSYS_UNCONNECTED_911), .B(
        _f_permutation__round__n1170 ), .Z(_f_permutation__round__n1168 ) );
  XOR2_X2 _f_permutation__round__U6903  ( .A(SYNOPSYS_UNCONNECTED_271), .B(
        SYNOPSYS_UNCONNECTED_591), .Z(_f_permutation__round__n1169 ) );
  XOR2_X2 _f_permutation__round__U6902  ( .A(_f_permutation__round_in[1457]), 
        .B(_f_permutation__round_in[1137]), .Z(_f_permutation__round__n1170 )
         );
  XOR2_X2 _f_permutation__round__U6901  ( .A(_f_permutation__round__n1967 ), 
        .B(_f_permutation__round__n2419 ), .Z(_f_permutation__round__n1969 )
         );
  XOR2_X2 _f_permutation__round__U6900  ( .A(SYNOPSYS_UNCONNECTED_846), .B(
        _f_permutation__round__n1969 ), .Z(_f_permutation__round__c[626] ) );
  XOR2_X2 _f_permutation__round__U6899  ( .A(SYNOPSYS_UNCONNECTED_717), .B(
        _f_permutation__round__n1968 ), .Z(_f_permutation__round__c[1523] ) );
  XOR2_X2 _f_permutation__round__U6898  ( .A(SYNOPSYS_UNCONNECTED_526), .B(
        _f_permutation__round__n1969 ), .Z(_f_permutation__round__c[562] ) );
  XOR2_X2 _f_permutation__round__U6897  ( .A(SYNOPSYS_UNCONNECTED_397), .B(
        _f_permutation__round__n1968 ), .Z(_f_permutation__round__c[1459] ) );
  XOR2_X2 _f_permutation__round__U6896  ( .A(SYNOPSYS_UNCONNECTED_206), .B(
        _f_permutation__round__n1969 ), .Z(_f_permutation__round__c[498] ) );
  XOR2_X2 _f_permutation__round__U6895  ( .A(SYNOPSYS_UNCONNECTED_77), .B(
        _f_permutation__round__n1968 ), .Z(_f_permutation__round__c[1395] ) );
  XOR2_X2 _f_permutation__round__U6894  ( .A(_f_permutation__round_in[1202]), 
        .B(_f_permutation__round__n1969 ), .Z(_f_permutation__round__c[434] )
         );
  XOR2_X2 _f_permutation__round__U6893  ( .A(_f_permutation__round_in[1331]), 
        .B(_f_permutation__round__n1968 ), .Z(_f_permutation__round__c[1331] )
         );
  XOR2_X2 _f_permutation__round__U6892  ( .A(_f_permutation__round_in[1522]), 
        .B(_f_permutation__round__n1969 ), .Z(_f_permutation__round__c[370] )
         );
  XOR2_X2 _f_permutation__round__U6891  ( .A(_f_permutation__round__n1172 ), 
        .B(_f_permutation__round__n1171 ), .Z(_f_permutation__round__n2181 )
         );
  XOR2_X2 _f_permutation__round__U6890  ( .A(SYNOPSYS_UNCONNECTED_848), .B(
        _f_permutation__round__n1173 ), .Z(_f_permutation__round__n1171 ) );
  XOR2_X2 _f_permutation__round__U6889  ( .A(SYNOPSYS_UNCONNECTED_208), .B(
        SYNOPSYS_UNCONNECTED_528), .Z(_f_permutation__round__n1172 ) );
  XOR2_X2 _f_permutation__round__U6888  ( .A(_f_permutation__round_in[1520]), 
        .B(_f_permutation__round_in[1200]), .Z(_f_permutation__round__n1173 )
         );
  XOR2_X2 _f_permutation__round__U6887  ( .A(_f_permutation__round__n1175 ), 
        .B(_f_permutation__round__n1174 ), .Z(_f_permutation__round__n2415 )
         );
  XOR2_X2 _f_permutation__round__U6886  ( .A(SYNOPSYS_UNCONNECTED_1039), .B(
        _f_permutation__round__n1176 ), .Z(_f_permutation__round__n1174 ) );
  XOR2_X2 _f_permutation__round__U6885  ( .A(SYNOPSYS_UNCONNECTED_399), .B(
        SYNOPSYS_UNCONNECTED_719), .Z(_f_permutation__round__n1175 ) );
  XOR2_X2 _f_permutation__round__U6884  ( .A(_f_permutation__round_in[1329]), 
        .B(SYNOPSYS_UNCONNECTED_79), .Z(_f_permutation__round__n1176 ) );
  XOR2_X2 _f_permutation__round__U6883  ( .A(_f_permutation__round__n2181 ), 
        .B(_f_permutation__round__n2415 ), .Z(_f_permutation__round__n2182 )
         );
  XOR2_X2 _f_permutation__round__U6882  ( .A(_f_permutation__round_in[1585]), 
        .B(_f_permutation__round__n2182 ), .Z(_f_permutation__round__c[49] )
         );
  XOR2_X2 _f_permutation__round__U6881  ( .A(_f_permutation__round__n1178 ), 
        .B(_f_permutation__round__n1177 ), .Z(_f_permutation__round__n1970 )
         );
  XOR2_X2 _f_permutation__round__U6880  ( .A(SYNOPSYS_UNCONNECTED_783), .B(
        _f_permutation__round__n1179 ), .Z(_f_permutation__round__n1177 ) );
  XOR2_X2 _f_permutation__round__U6879  ( .A(SYNOPSYS_UNCONNECTED_143), .B(
        SYNOPSYS_UNCONNECTED_463), .Z(_f_permutation__round__n1178 ) );
  XOR2_X2 _f_permutation__round__U6878  ( .A(_f_permutation__round_in[1585]), 
        .B(_f_permutation__round_in[1265]), .Z(_f_permutation__round__n1179 )
         );
  XOR2_X2 _f_permutation__round__U6877  ( .A(_f_permutation__round__n1181 ), 
        .B(_f_permutation__round__n1180 ), .Z(_f_permutation__round__n2168 )
         );
  XOR2_X2 _f_permutation__round__U6876  ( .A(SYNOPSYS_UNCONNECTED_974), .B(
        _f_permutation__round__n1182 ), .Z(_f_permutation__round__n1180 ) );
  XOR2_X2 _f_permutation__round__U6875  ( .A(SYNOPSYS_UNCONNECTED_334), .B(
        SYNOPSYS_UNCONNECTED_654), .Z(_f_permutation__round__n1181 ) );
  XOR2_X2 _f_permutation__round__U6874  ( .A(_f_permutation__round_in[1394]), 
        .B(_f_permutation__round_in[1074]), .Z(_f_permutation__round__n1182 )
         );
  XOR2_X2 _f_permutation__round__U6873  ( .A(_f_permutation__round__n1970 ), 
        .B(_f_permutation__round__n2168 ), .Z(_f_permutation__round__n1971 )
         );
  XOR2_X2 _f_permutation__round__U6872  ( .A(SYNOPSYS_UNCONNECTED_1038), .B(
        _f_permutation__round__n1971 ), .Z(_f_permutation__round__c[1586] ) );
  XOR2_X2 _f_permutation__round__U6871  ( .A(_f_permutation__round__n1184 ), 
        .B(_f_permutation__round__n1183 ), .Z(_f_permutation__round__n2422 )
         );
  XOR2_X2 _f_permutation__round__U6870  ( .A(SYNOPSYS_UNCONNECTED_912), .B(
        _f_permutation__round__n1185 ), .Z(_f_permutation__round__n1183 ) );
  XOR2_X2 _f_permutation__round__U6869  ( .A(SYNOPSYS_UNCONNECTED_272), .B(
        SYNOPSYS_UNCONNECTED_592), .Z(_f_permutation__round__n1184 ) );
  XOR2_X2 _f_permutation__round__U6868  ( .A(_f_permutation__round_in[1456]), 
        .B(_f_permutation__round_in[1136]), .Z(_f_permutation__round__n1185 )
         );
  XOR2_X2 _f_permutation__round__U6867  ( .A(_f_permutation__round__n1970 ), 
        .B(_f_permutation__round__n2422 ), .Z(_f_permutation__round__n1972 )
         );
  XOR2_X2 _f_permutation__round__U6866  ( .A(SYNOPSYS_UNCONNECTED_847), .B(
        _f_permutation__round__n1972 ), .Z(_f_permutation__round__c[625] ) );
  XOR2_X2 _f_permutation__round__U6865  ( .A(SYNOPSYS_UNCONNECTED_718), .B(
        _f_permutation__round__n1971 ), .Z(_f_permutation__round__c[1522] ) );
  XOR2_X2 _f_permutation__round__U6864  ( .A(SYNOPSYS_UNCONNECTED_527), .B(
        _f_permutation__round__n1972 ), .Z(_f_permutation__round__c[561] ) );
  XOR2_X2 _f_permutation__round__U6863  ( .A(SYNOPSYS_UNCONNECTED_398), .B(
        _f_permutation__round__n1971 ), .Z(_f_permutation__round__c[1458] ) );
  XOR2_X2 _f_permutation__round__U6862  ( .A(SYNOPSYS_UNCONNECTED_207), .B(
        _f_permutation__round__n1972 ), .Z(_f_permutation__round__c[497] ) );
  XOR2_X2 _f_permutation__round__U6861  ( .A(SYNOPSYS_UNCONNECTED_78), .B(
        _f_permutation__round__n1971 ), .Z(_f_permutation__round__c[1394] ) );
  XOR2_X2 _f_permutation__round__U6860  ( .A(_f_permutation__round_in[1201]), 
        .B(_f_permutation__round__n1972 ), .Z(_f_permutation__round__c[433] )
         );
  XOR2_X2 _f_permutation__round__U6859  ( .A(_f_permutation__round_in[1330]), 
        .B(_f_permutation__round__n1971 ), .Z(_f_permutation__round__c[1330] )
         );
  XOR2_X2 _f_permutation__round__U6858  ( .A(_f_permutation__round_in[1521]), 
        .B(_f_permutation__round__n1972 ), .Z(_f_permutation__round__c[369] )
         );
  XOR2_X2 _f_permutation__round__U6857  ( .A(_f_permutation__round__n1187 ), 
        .B(_f_permutation__round__n1186 ), .Z(_f_permutation__round__n2185 )
         );
  XOR2_X2 _f_permutation__round__U6856  ( .A(SYNOPSYS_UNCONNECTED_849), .B(
        _f_permutation__round__n1188 ), .Z(_f_permutation__round__n1186 ) );
  XOR2_X2 _f_permutation__round__U6855  ( .A(SYNOPSYS_UNCONNECTED_209), .B(
        SYNOPSYS_UNCONNECTED_529), .Z(_f_permutation__round__n1187 ) );
  XOR2_X2 _f_permutation__round__U6854  ( .A(_f_permutation__round_in[1519]), 
        .B(_f_permutation__round_in[1199]), .Z(_f_permutation__round__n1188 )
         );
  XOR2_X2 _f_permutation__round__U6853  ( .A(_f_permutation__round__n1190 ), 
        .B(_f_permutation__round__n1189 ), .Z(_f_permutation__round__n2418 )
         );
  XOR2_X2 _f_permutation__round__U6852  ( .A(SYNOPSYS_UNCONNECTED_1040), .B(
        _f_permutation__round__n1191 ), .Z(_f_permutation__round__n1189 ) );
  XOR2_X2 _f_permutation__round__U6851  ( .A(SYNOPSYS_UNCONNECTED_400), .B(
        SYNOPSYS_UNCONNECTED_720), .Z(_f_permutation__round__n1190 ) );
  XOR2_X2 _f_permutation__round__U6850  ( .A(_f_permutation__round_in[1328]), 
        .B(SYNOPSYS_UNCONNECTED_80), .Z(_f_permutation__round__n1191 ) );
  XOR2_X2 _f_permutation__round__U6849  ( .A(_f_permutation__round__n2185 ), 
        .B(_f_permutation__round__n2418 ), .Z(_f_permutation__round__n2186 )
         );
  XOR2_X2 _f_permutation__round__U6848  ( .A(_f_permutation__round_in[1584]), 
        .B(_f_permutation__round__n2186 ), .Z(_f_permutation__round__c[48] )
         );
  XOR2_X2 _f_permutation__round__U6847  ( .A(_f_permutation__round__n1193 ), 
        .B(_f_permutation__round__n1192 ), .Z(_f_permutation__round__n1973 )
         );
  XOR2_X2 _f_permutation__round__U6846  ( .A(SYNOPSYS_UNCONNECTED_784), .B(
        _f_permutation__round__n1194 ), .Z(_f_permutation__round__n1192 ) );
  XOR2_X2 _f_permutation__round__U6845  ( .A(SYNOPSYS_UNCONNECTED_144), .B(
        SYNOPSYS_UNCONNECTED_464), .Z(_f_permutation__round__n1193 ) );
  XOR2_X2 _f_permutation__round__U6844  ( .A(_f_permutation__round_in[1584]), 
        .B(_f_permutation__round_in[1264]), .Z(_f_permutation__round__n1194 )
         );
  XOR2_X2 _f_permutation__round__U6843  ( .A(_f_permutation__round__n1196 ), 
        .B(_f_permutation__round__n1195 ), .Z(_f_permutation__round__n2172 )
         );
  XOR2_X2 _f_permutation__round__U6842  ( .A(SYNOPSYS_UNCONNECTED_975), .B(
        _f_permutation__round__n1197 ), .Z(_f_permutation__round__n1195 ) );
  XOR2_X2 _f_permutation__round__U6841  ( .A(SYNOPSYS_UNCONNECTED_335), .B(
        SYNOPSYS_UNCONNECTED_655), .Z(_f_permutation__round__n1196 ) );
  XOR2_X2 _f_permutation__round__U6840  ( .A(_f_permutation__round_in[1393]), 
        .B(_f_permutation__round_in[1073]), .Z(_f_permutation__round__n1197 )
         );
  XOR2_X2 _f_permutation__round__U6839  ( .A(_f_permutation__round__n1973 ), 
        .B(_f_permutation__round__n2172 ), .Z(_f_permutation__round__n1974 )
         );
  XOR2_X2 _f_permutation__round__U6838  ( .A(SYNOPSYS_UNCONNECTED_1039), .B(
        _f_permutation__round__n1974 ), .Z(_f_permutation__round__c[1585] ) );
  XOR2_X2 _f_permutation__round__U6837  ( .A(_f_permutation__round__n1199 ), 
        .B(_f_permutation__round__n1198 ), .Z(_f_permutation__round__n2425 )
         );
  XOR2_X2 _f_permutation__round__U6836  ( .A(SYNOPSYS_UNCONNECTED_913), .B(
        _f_permutation__round__n1200 ), .Z(_f_permutation__round__n1198 ) );
  XOR2_X2 _f_permutation__round__U6835  ( .A(SYNOPSYS_UNCONNECTED_273), .B(
        SYNOPSYS_UNCONNECTED_593), .Z(_f_permutation__round__n1199 ) );
  XOR2_X2 _f_permutation__round__U6834  ( .A(_f_permutation__round_in[1455]), 
        .B(_f_permutation__round_in[1135]), .Z(_f_permutation__round__n1200 )
         );
  XOR2_X2 _f_permutation__round__U6833  ( .A(_f_permutation__round__n1973 ), 
        .B(_f_permutation__round__n2425 ), .Z(_f_permutation__round__n1975 )
         );
  XOR2_X2 _f_permutation__round__U6832  ( .A(SYNOPSYS_UNCONNECTED_848), .B(
        _f_permutation__round__n1975 ), .Z(_f_permutation__round__c[624] ) );
  XOR2_X2 _f_permutation__round__U6831  ( .A(SYNOPSYS_UNCONNECTED_719), .B(
        _f_permutation__round__n1974 ), .Z(_f_permutation__round__c[1521] ) );
  XOR2_X2 _f_permutation__round__U6830  ( .A(SYNOPSYS_UNCONNECTED_528), .B(
        _f_permutation__round__n1975 ), .Z(_f_permutation__round__c[560] ) );
  XOR2_X2 _f_permutation__round__U6829  ( .A(SYNOPSYS_UNCONNECTED_399), .B(
        _f_permutation__round__n1974 ), .Z(_f_permutation__round__c[1457] ) );
  XOR2_X2 _f_permutation__round__U6828  ( .A(SYNOPSYS_UNCONNECTED_208), .B(
        _f_permutation__round__n1975 ), .Z(_f_permutation__round__c[496] ) );
  XOR2_X2 _f_permutation__round__U6827  ( .A(SYNOPSYS_UNCONNECTED_79), .B(
        _f_permutation__round__n1974 ), .Z(_f_permutation__round__c[1393] ) );
  XOR2_X2 _f_permutation__round__U6826  ( .A(_f_permutation__round_in[1200]), 
        .B(_f_permutation__round__n1975 ), .Z(_f_permutation__round__c[432] )
         );
  XOR2_X2 _f_permutation__round__U6825  ( .A(_f_permutation__round_in[1329]), 
        .B(_f_permutation__round__n1974 ), .Z(_f_permutation__round__c[1329] )
         );
  XOR2_X2 _f_permutation__round__U6824  ( .A(_f_permutation__round_in[1520]), 
        .B(_f_permutation__round__n1975 ), .Z(_f_permutation__round__c[368] )
         );
  XOR2_X2 _f_permutation__round__U6823  ( .A(_f_permutation__round__n1202 ), 
        .B(_f_permutation__round__n1201 ), .Z(_f_permutation__round__n2189 )
         );
  XOR2_X2 _f_permutation__round__U6822  ( .A(SYNOPSYS_UNCONNECTED_850), .B(
        _f_permutation__round__n1203 ), .Z(_f_permutation__round__n1201 ) );
  XOR2_X2 _f_permutation__round__U6821  ( .A(SYNOPSYS_UNCONNECTED_210), .B(
        SYNOPSYS_UNCONNECTED_530), .Z(_f_permutation__round__n1202 ) );
  XOR2_X2 _f_permutation__round__U6820  ( .A(_f_permutation__round_in[1518]), 
        .B(_f_permutation__round_in[1198]), .Z(_f_permutation__round__n1203 )
         );
  XOR2_X2 _f_permutation__round__U6819  ( .A(_f_permutation__round__n1205 ), 
        .B(_f_permutation__round__n1204 ), .Z(_f_permutation__round__n2421 )
         );
  XOR2_X2 _f_permutation__round__U6818  ( .A(SYNOPSYS_UNCONNECTED_1041), .B(
        _f_permutation__round__n1206 ), .Z(_f_permutation__round__n1204 ) );
  XOR2_X2 _f_permutation__round__U6817  ( .A(SYNOPSYS_UNCONNECTED_401), .B(
        SYNOPSYS_UNCONNECTED_721), .Z(_f_permutation__round__n1205 ) );
  XOR2_X2 _f_permutation__round__U6816  ( .A(_f_permutation__round_in[1327]), 
        .B(SYNOPSYS_UNCONNECTED_81), .Z(_f_permutation__round__n1206 ) );
  XOR2_X2 _f_permutation__round__U6815  ( .A(_f_permutation__round__n2189 ), 
        .B(_f_permutation__round__n2421 ), .Z(_f_permutation__round__n2190 )
         );
  XOR2_X2 _f_permutation__round__U6814  ( .A(_f_permutation__round_in[1583]), 
        .B(_f_permutation__round__n2190 ), .Z(_f_permutation__round__c[47] )
         );
  XOR2_X2 _f_permutation__round__U6813  ( .A(_f_permutation__round__n1208 ), 
        .B(_f_permutation__round__n1207 ), .Z(_f_permutation__round__n1976 )
         );
  XOR2_X2 _f_permutation__round__U6812  ( .A(SYNOPSYS_UNCONNECTED_785), .B(
        _f_permutation__round__n1209 ), .Z(_f_permutation__round__n1207 ) );
  XOR2_X2 _f_permutation__round__U6811  ( .A(SYNOPSYS_UNCONNECTED_145), .B(
        SYNOPSYS_UNCONNECTED_465), .Z(_f_permutation__round__n1208 ) );
  XOR2_X2 _f_permutation__round__U6810  ( .A(_f_permutation__round_in[1583]), 
        .B(_f_permutation__round_in[1263]), .Z(_f_permutation__round__n1209 )
         );
  XOR2_X2 _f_permutation__round__U6809  ( .A(_f_permutation__round__n1211 ), 
        .B(_f_permutation__round__n1210 ), .Z(_f_permutation__round__n2176 )
         );
  XOR2_X2 _f_permutation__round__U6808  ( .A(SYNOPSYS_UNCONNECTED_976), .B(
        _f_permutation__round__n1212 ), .Z(_f_permutation__round__n1210 ) );
  XOR2_X2 _f_permutation__round__U6807  ( .A(SYNOPSYS_UNCONNECTED_336), .B(
        SYNOPSYS_UNCONNECTED_656), .Z(_f_permutation__round__n1211 ) );
  XOR2_X2 _f_permutation__round__U6806  ( .A(_f_permutation__round_in[1392]), 
        .B(_f_permutation__round_in[1072]), .Z(_f_permutation__round__n1212 )
         );
  XOR2_X2 _f_permutation__round__U6805  ( .A(_f_permutation__round__n1976 ), 
        .B(_f_permutation__round__n2176 ), .Z(_f_permutation__round__n1977 )
         );
  XOR2_X2 _f_permutation__round__U6804  ( .A(SYNOPSYS_UNCONNECTED_1040), .B(
        _f_permutation__round__n1977 ), .Z(_f_permutation__round__c[1584] ) );
  XOR2_X2 _f_permutation__round__U6803  ( .A(_f_permutation__round__n1214 ), 
        .B(_f_permutation__round__n1213 ), .Z(_f_permutation__round__n2428 )
         );
  XOR2_X2 _f_permutation__round__U6802  ( .A(SYNOPSYS_UNCONNECTED_914), .B(
        _f_permutation__round__n1215 ), .Z(_f_permutation__round__n1213 ) );
  XOR2_X2 _f_permutation__round__U6801  ( .A(SYNOPSYS_UNCONNECTED_274), .B(
        SYNOPSYS_UNCONNECTED_594), .Z(_f_permutation__round__n1214 ) );
  XOR2_X2 _f_permutation__round__U6800  ( .A(_f_permutation__round_in[1454]), 
        .B(_f_permutation__round_in[1134]), .Z(_f_permutation__round__n1215 )
         );
  XOR2_X2 _f_permutation__round__U6799  ( .A(_f_permutation__round__n1976 ), 
        .B(_f_permutation__round__n2428 ), .Z(_f_permutation__round__n1978 )
         );
  XOR2_X2 _f_permutation__round__U6798  ( .A(SYNOPSYS_UNCONNECTED_849), .B(
        _f_permutation__round__n1978 ), .Z(_f_permutation__round__c[623] ) );
  XOR2_X2 _f_permutation__round__U6797  ( .A(SYNOPSYS_UNCONNECTED_720), .B(
        _f_permutation__round__n1977 ), .Z(_f_permutation__round__c[1520] ) );
  XOR2_X2 _f_permutation__round__U6796  ( .A(SYNOPSYS_UNCONNECTED_529), .B(
        _f_permutation__round__n1978 ), .Z(_f_permutation__round__c[559] ) );
  XOR2_X2 _f_permutation__round__U6795  ( .A(SYNOPSYS_UNCONNECTED_400), .B(
        _f_permutation__round__n1977 ), .Z(_f_permutation__round__c[1456] ) );
  XOR2_X2 _f_permutation__round__U6794  ( .A(SYNOPSYS_UNCONNECTED_209), .B(
        _f_permutation__round__n1978 ), .Z(_f_permutation__round__c[495] ) );
  XOR2_X2 _f_permutation__round__U6793  ( .A(SYNOPSYS_UNCONNECTED_80), .B(
        _f_permutation__round__n1977 ), .Z(_f_permutation__round__c[1392] ) );
  XOR2_X2 _f_permutation__round__U6792  ( .A(_f_permutation__round_in[1199]), 
        .B(_f_permutation__round__n1978 ), .Z(_f_permutation__round__c[431] )
         );
  XOR2_X2 _f_permutation__round__U6791  ( .A(_f_permutation__round_in[1328]), 
        .B(_f_permutation__round__n1977 ), .Z(_f_permutation__round__c[1328] )
         );
  XOR2_X2 _f_permutation__round__U6790  ( .A(_f_permutation__round_in[1519]), 
        .B(_f_permutation__round__n1978 ), .Z(_f_permutation__round__c[367] )
         );
  XOR2_X2 _f_permutation__round__U6789  ( .A(_f_permutation__round__n1217 ), 
        .B(_f_permutation__round__n1216 ), .Z(_f_permutation__round__n2193 )
         );
  XOR2_X2 _f_permutation__round__U6788  ( .A(SYNOPSYS_UNCONNECTED_851), .B(
        _f_permutation__round__n1218 ), .Z(_f_permutation__round__n1216 ) );
  XOR2_X2 _f_permutation__round__U6787  ( .A(SYNOPSYS_UNCONNECTED_211), .B(
        SYNOPSYS_UNCONNECTED_531), .Z(_f_permutation__round__n1217 ) );
  XOR2_X2 _f_permutation__round__U6786  ( .A(_f_permutation__round_in[1517]), 
        .B(_f_permutation__round_in[1197]), .Z(_f_permutation__round__n1218 )
         );
  XOR2_X2 _f_permutation__round__U6785  ( .A(_f_permutation__round__n1220 ), 
        .B(_f_permutation__round__n1219 ), .Z(_f_permutation__round__n2424 )
         );
  XOR2_X2 _f_permutation__round__U6784  ( .A(SYNOPSYS_UNCONNECTED_1042), .B(
        _f_permutation__round__n1221 ), .Z(_f_permutation__round__n1219 ) );
  XOR2_X2 _f_permutation__round__U6783  ( .A(SYNOPSYS_UNCONNECTED_402), .B(
        SYNOPSYS_UNCONNECTED_722), .Z(_f_permutation__round__n1220 ) );
  XOR2_X2 _f_permutation__round__U6782  ( .A(_f_permutation__round_in[1326]), 
        .B(SYNOPSYS_UNCONNECTED_82), .Z(_f_permutation__round__n1221 ) );
  XOR2_X2 _f_permutation__round__U6781  ( .A(_f_permutation__round__n2193 ), 
        .B(_f_permutation__round__n2424 ), .Z(_f_permutation__round__n2194 )
         );
  XOR2_X2 _f_permutation__round__U6780  ( .A(_f_permutation__round_in[1582]), 
        .B(_f_permutation__round__n2194 ), .Z(_f_permutation__round__c[46] )
         );
  XOR2_X2 _f_permutation__round__U6779  ( .A(_f_permutation__round__n1223 ), 
        .B(_f_permutation__round__n1222 ), .Z(_f_permutation__round__n1979 )
         );
  XOR2_X2 _f_permutation__round__U6778  ( .A(SYNOPSYS_UNCONNECTED_786), .B(
        _f_permutation__round__n1224 ), .Z(_f_permutation__round__n1222 ) );
  XOR2_X2 _f_permutation__round__U6777  ( .A(SYNOPSYS_UNCONNECTED_146), .B(
        SYNOPSYS_UNCONNECTED_466), .Z(_f_permutation__round__n1223 ) );
  XOR2_X2 _f_permutation__round__U6776  ( .A(_f_permutation__round_in[1582]), 
        .B(_f_permutation__round_in[1262]), .Z(_f_permutation__round__n1224 )
         );
  XOR2_X2 _f_permutation__round__U6775  ( .A(_f_permutation__round__n1226 ), 
        .B(_f_permutation__round__n1225 ), .Z(_f_permutation__round__n2180 )
         );
  XOR2_X2 _f_permutation__round__U6774  ( .A(SYNOPSYS_UNCONNECTED_977), .B(
        _f_permutation__round__n1227 ), .Z(_f_permutation__round__n1225 ) );
  XOR2_X2 _f_permutation__round__U6773  ( .A(SYNOPSYS_UNCONNECTED_337), .B(
        SYNOPSYS_UNCONNECTED_657), .Z(_f_permutation__round__n1226 ) );
  XOR2_X2 _f_permutation__round__U6772  ( .A(_f_permutation__round_in[1391]), 
        .B(_f_permutation__round_in[1071]), .Z(_f_permutation__round__n1227 )
         );
  XOR2_X2 _f_permutation__round__U6771  ( .A(_f_permutation__round__n1979 ), 
        .B(_f_permutation__round__n2180 ), .Z(_f_permutation__round__n1980 )
         );
  XOR2_X2 _f_permutation__round__U6770  ( .A(SYNOPSYS_UNCONNECTED_1041), .B(
        _f_permutation__round__n1980 ), .Z(_f_permutation__round__c[1583] ) );
  XOR2_X2 _f_permutation__round__U6769  ( .A(_f_permutation__round__n1229 ), 
        .B(_f_permutation__round__n1228 ), .Z(_f_permutation__round__n2431 )
         );
  XOR2_X2 _f_permutation__round__U6768  ( .A(SYNOPSYS_UNCONNECTED_915), .B(
        _f_permutation__round__n1230 ), .Z(_f_permutation__round__n1228 ) );
  XOR2_X2 _f_permutation__round__U6767  ( .A(SYNOPSYS_UNCONNECTED_275), .B(
        SYNOPSYS_UNCONNECTED_595), .Z(_f_permutation__round__n1229 ) );
  XOR2_X2 _f_permutation__round__U6766  ( .A(_f_permutation__round_in[1453]), 
        .B(_f_permutation__round_in[1133]), .Z(_f_permutation__round__n1230 )
         );
  XOR2_X2 _f_permutation__round__U6765  ( .A(_f_permutation__round__n1979 ), 
        .B(_f_permutation__round__n2431 ), .Z(_f_permutation__round__n1981 )
         );
  XOR2_X2 _f_permutation__round__U6764  ( .A(SYNOPSYS_UNCONNECTED_850), .B(
        _f_permutation__round__n1981 ), .Z(_f_permutation__round__c[622] ) );
  XOR2_X2 _f_permutation__round__U6763  ( .A(SYNOPSYS_UNCONNECTED_721), .B(
        _f_permutation__round__n1980 ), .Z(_f_permutation__round__c[1519] ) );
  XOR2_X2 _f_permutation__round__U6762  ( .A(SYNOPSYS_UNCONNECTED_530), .B(
        _f_permutation__round__n1981 ), .Z(_f_permutation__round__c[558] ) );
  XOR2_X2 _f_permutation__round__U6761  ( .A(SYNOPSYS_UNCONNECTED_401), .B(
        _f_permutation__round__n1980 ), .Z(_f_permutation__round__c[1455] ) );
  XOR2_X2 _f_permutation__round__U6760  ( .A(SYNOPSYS_UNCONNECTED_210), .B(
        _f_permutation__round__n1981 ), .Z(_f_permutation__round__c[494] ) );
  XOR2_X2 _f_permutation__round__U6759  ( .A(SYNOPSYS_UNCONNECTED_81), .B(
        _f_permutation__round__n1980 ), .Z(_f_permutation__round__c[1391] ) );
  XOR2_X2 _f_permutation__round__U6758  ( .A(_f_permutation__round_in[1198]), 
        .B(_f_permutation__round__n1981 ), .Z(_f_permutation__round__c[430] )
         );
  XOR2_X2 _f_permutation__round__U6757  ( .A(_f_permutation__round_in[1327]), 
        .B(_f_permutation__round__n1980 ), .Z(_f_permutation__round__c[1327] )
         );
  XOR2_X2 _f_permutation__round__U6756  ( .A(_f_permutation__round_in[1518]), 
        .B(_f_permutation__round__n1981 ), .Z(_f_permutation__round__c[366] )
         );
  XOR2_X2 _f_permutation__round__U6755  ( .A(_f_permutation__round__n1232 ), 
        .B(_f_permutation__round__n1231 ), .Z(_f_permutation__round__n2197 )
         );
  XOR2_X2 _f_permutation__round__U6754  ( .A(SYNOPSYS_UNCONNECTED_852), .B(
        _f_permutation__round__n1233 ), .Z(_f_permutation__round__n1231 ) );
  XOR2_X2 _f_permutation__round__U6753  ( .A(SYNOPSYS_UNCONNECTED_212), .B(
        SYNOPSYS_UNCONNECTED_532), .Z(_f_permutation__round__n1232 ) );
  XOR2_X2 _f_permutation__round__U6752  ( .A(_f_permutation__round_in[1516]), 
        .B(_f_permutation__round_in[1196]), .Z(_f_permutation__round__n1233 )
         );
  XOR2_X2 _f_permutation__round__U6751  ( .A(_f_permutation__round__n1235 ), 
        .B(_f_permutation__round__n1234 ), .Z(_f_permutation__round__n2427 )
         );
  XOR2_X2 _f_permutation__round__U6750  ( .A(SYNOPSYS_UNCONNECTED_1043), .B(
        _f_permutation__round__n1236 ), .Z(_f_permutation__round__n1234 ) );
  XOR2_X2 _f_permutation__round__U6749  ( .A(SYNOPSYS_UNCONNECTED_403), .B(
        SYNOPSYS_UNCONNECTED_723), .Z(_f_permutation__round__n1235 ) );
  XOR2_X2 _f_permutation__round__U6748  ( .A(_f_permutation__round_in[1325]), 
        .B(SYNOPSYS_UNCONNECTED_83), .Z(_f_permutation__round__n1236 ) );
  XOR2_X2 _f_permutation__round__U6747  ( .A(_f_permutation__round__n2197 ), 
        .B(_f_permutation__round__n2427 ), .Z(_f_permutation__round__n2198 )
         );
  XOR2_X2 _f_permutation__round__U6746  ( .A(_f_permutation__round_in[1581]), 
        .B(_f_permutation__round__n2198 ), .Z(_f_permutation__round__c[45] )
         );
  XOR2_X2 _f_permutation__round__U6745  ( .A(_f_permutation__round__n1238 ), 
        .B(_f_permutation__round__n1237 ), .Z(_f_permutation__round__n1982 )
         );
  XOR2_X2 _f_permutation__round__U6744  ( .A(SYNOPSYS_UNCONNECTED_787), .B(
        _f_permutation__round__n1239 ), .Z(_f_permutation__round__n1237 ) );
  XOR2_X2 _f_permutation__round__U6743  ( .A(SYNOPSYS_UNCONNECTED_147), .B(
        SYNOPSYS_UNCONNECTED_467), .Z(_f_permutation__round__n1238 ) );
  XOR2_X2 _f_permutation__round__U6742  ( .A(_f_permutation__round_in[1581]), 
        .B(_f_permutation__round_in[1261]), .Z(_f_permutation__round__n1239 )
         );
  XOR2_X2 _f_permutation__round__U6741  ( .A(_f_permutation__round__n1241 ), 
        .B(_f_permutation__round__n1240 ), .Z(_f_permutation__round__n2184 )
         );
  XOR2_X2 _f_permutation__round__U6740  ( .A(SYNOPSYS_UNCONNECTED_978), .B(
        _f_permutation__round__n1242 ), .Z(_f_permutation__round__n1240 ) );
  XOR2_X2 _f_permutation__round__U6739  ( .A(SYNOPSYS_UNCONNECTED_338), .B(
        SYNOPSYS_UNCONNECTED_658), .Z(_f_permutation__round__n1241 ) );
  XOR2_X2 _f_permutation__round__U6738  ( .A(_f_permutation__round_in[1390]), 
        .B(_f_permutation__round_in[1070]), .Z(_f_permutation__round__n1242 )
         );
  XOR2_X2 _f_permutation__round__U6737  ( .A(_f_permutation__round__n1982 ), 
        .B(_f_permutation__round__n2184 ), .Z(_f_permutation__round__n1983 )
         );
  XOR2_X2 _f_permutation__round__U6736  ( .A(SYNOPSYS_UNCONNECTED_1042), .B(
        _f_permutation__round__n1983 ), .Z(_f_permutation__round__c[1582] ) );
  XOR2_X2 _f_permutation__round__U6735  ( .A(_f_permutation__round__n1244 ), 
        .B(_f_permutation__round__n1243 ), .Z(_f_permutation__round__n2434 )
         );
  XOR2_X2 _f_permutation__round__U6734  ( .A(SYNOPSYS_UNCONNECTED_916), .B(
        _f_permutation__round__n1245 ), .Z(_f_permutation__round__n1243 ) );
  XOR2_X2 _f_permutation__round__U6733  ( .A(SYNOPSYS_UNCONNECTED_276), .B(
        SYNOPSYS_UNCONNECTED_596), .Z(_f_permutation__round__n1244 ) );
  XOR2_X2 _f_permutation__round__U6732  ( .A(_f_permutation__round_in[1452]), 
        .B(_f_permutation__round_in[1132]), .Z(_f_permutation__round__n1245 )
         );
  XOR2_X2 _f_permutation__round__U6731  ( .A(_f_permutation__round__n1982 ), 
        .B(_f_permutation__round__n2434 ), .Z(_f_permutation__round__n1984 )
         );
  XOR2_X2 _f_permutation__round__U6730  ( .A(SYNOPSYS_UNCONNECTED_851), .B(
        _f_permutation__round__n1984 ), .Z(_f_permutation__round__c[621] ) );
  XOR2_X2 _f_permutation__round__U6729  ( .A(SYNOPSYS_UNCONNECTED_722), .B(
        _f_permutation__round__n1983 ), .Z(_f_permutation__round__c[1518] ) );
  XOR2_X2 _f_permutation__round__U6728  ( .A(SYNOPSYS_UNCONNECTED_531), .B(
        _f_permutation__round__n1984 ), .Z(_f_permutation__round__c[557] ) );
  XOR2_X2 _f_permutation__round__U6727  ( .A(SYNOPSYS_UNCONNECTED_402), .B(
        _f_permutation__round__n1983 ), .Z(_f_permutation__round__c[1454] ) );
  XOR2_X2 _f_permutation__round__U6726  ( .A(SYNOPSYS_UNCONNECTED_211), .B(
        _f_permutation__round__n1984 ), .Z(_f_permutation__round__c[493] ) );
  XOR2_X2 _f_permutation__round__U6725  ( .A(SYNOPSYS_UNCONNECTED_82), .B(
        _f_permutation__round__n1983 ), .Z(_f_permutation__round__c[1390] ) );
  XOR2_X2 _f_permutation__round__U6724  ( .A(_f_permutation__round_in[1197]), 
        .B(_f_permutation__round__n1984 ), .Z(_f_permutation__round__c[429] )
         );
  XOR2_X2 _f_permutation__round__U6723  ( .A(_f_permutation__round_in[1326]), 
        .B(_f_permutation__round__n1983 ), .Z(_f_permutation__round__c[1326] )
         );
  XOR2_X2 _f_permutation__round__U6722  ( .A(_f_permutation__round_in[1517]), 
        .B(_f_permutation__round__n1984 ), .Z(_f_permutation__round__c[365] )
         );
  XOR2_X2 _f_permutation__round__U6721  ( .A(_f_permutation__round__n1247 ), 
        .B(_f_permutation__round__n1246 ), .Z(_f_permutation__round__n2201 )
         );
  XOR2_X2 _f_permutation__round__U6720  ( .A(SYNOPSYS_UNCONNECTED_853), .B(
        _f_permutation__round__n1248 ), .Z(_f_permutation__round__n1246 ) );
  XOR2_X2 _f_permutation__round__U6719  ( .A(SYNOPSYS_UNCONNECTED_213), .B(
        SYNOPSYS_UNCONNECTED_533), .Z(_f_permutation__round__n1247 ) );
  XOR2_X2 _f_permutation__round__U6718  ( .A(_f_permutation__round_in[1515]), 
        .B(_f_permutation__round_in[1195]), .Z(_f_permutation__round__n1248 )
         );
  XOR2_X2 _f_permutation__round__U6717  ( .A(_f_permutation__round__n1250 ), 
        .B(_f_permutation__round__n1249 ), .Z(_f_permutation__round__n2430 )
         );
  XOR2_X2 _f_permutation__round__U6716  ( .A(SYNOPSYS_UNCONNECTED_1044), .B(
        _f_permutation__round__n1251 ), .Z(_f_permutation__round__n1249 ) );
  XOR2_X2 _f_permutation__round__U6715  ( .A(SYNOPSYS_UNCONNECTED_404), .B(
        SYNOPSYS_UNCONNECTED_724), .Z(_f_permutation__round__n1250 ) );
  XOR2_X2 _f_permutation__round__U6714  ( .A(_f_permutation__round_in[1324]), 
        .B(SYNOPSYS_UNCONNECTED_84), .Z(_f_permutation__round__n1251 ) );
  XOR2_X2 _f_permutation__round__U6713  ( .A(_f_permutation__round__n2201 ), 
        .B(_f_permutation__round__n2430 ), .Z(_f_permutation__round__n2202 )
         );
  XOR2_X2 _f_permutation__round__U6712  ( .A(_f_permutation__round_in[1580]), 
        .B(_f_permutation__round__n2202 ), .Z(_f_permutation__round__c[44] )
         );
  XOR2_X2 _f_permutation__round__U6711  ( .A(_f_permutation__round__n1253 ), 
        .B(_f_permutation__round__n1252 ), .Z(_f_permutation__round__n1985 )
         );
  XOR2_X2 _f_permutation__round__U6710  ( .A(SYNOPSYS_UNCONNECTED_788), .B(
        _f_permutation__round__n1254 ), .Z(_f_permutation__round__n1252 ) );
  XOR2_X2 _f_permutation__round__U6709  ( .A(SYNOPSYS_UNCONNECTED_148), .B(
        SYNOPSYS_UNCONNECTED_468), .Z(_f_permutation__round__n1253 ) );
  XOR2_X2 _f_permutation__round__U6708  ( .A(_f_permutation__round_in[1580]), 
        .B(_f_permutation__round_in[1260]), .Z(_f_permutation__round__n1254 )
         );
  XOR2_X2 _f_permutation__round__U6707  ( .A(_f_permutation__round__n1256 ), 
        .B(_f_permutation__round__n1255 ), .Z(_f_permutation__round__n2188 )
         );
  XOR2_X2 _f_permutation__round__U6706  ( .A(SYNOPSYS_UNCONNECTED_979), .B(
        _f_permutation__round__n1257 ), .Z(_f_permutation__round__n1255 ) );
  XOR2_X2 _f_permutation__round__U6705  ( .A(SYNOPSYS_UNCONNECTED_339), .B(
        SYNOPSYS_UNCONNECTED_659), .Z(_f_permutation__round__n1256 ) );
  XOR2_X2 _f_permutation__round__U6704  ( .A(_f_permutation__round_in[1389]), 
        .B(_f_permutation__round_in[1069]), .Z(_f_permutation__round__n1257 )
         );
  XOR2_X2 _f_permutation__round__U6703  ( .A(_f_permutation__round__n1985 ), 
        .B(_f_permutation__round__n2188 ), .Z(_f_permutation__round__n1986 )
         );
  XOR2_X2 _f_permutation__round__U6702  ( .A(SYNOPSYS_UNCONNECTED_1043), .B(
        _f_permutation__round__n1986 ), .Z(_f_permutation__round__c[1581] ) );
  XOR2_X2 _f_permutation__round__U6701  ( .A(_f_permutation__round__n1259 ), 
        .B(_f_permutation__round__n1258 ), .Z(_f_permutation__round__n2437 )
         );
  XOR2_X2 _f_permutation__round__U6700  ( .A(SYNOPSYS_UNCONNECTED_917), .B(
        _f_permutation__round__n1260 ), .Z(_f_permutation__round__n1258 ) );
  XOR2_X2 _f_permutation__round__U6699  ( .A(SYNOPSYS_UNCONNECTED_277), .B(
        SYNOPSYS_UNCONNECTED_597), .Z(_f_permutation__round__n1259 ) );
  XOR2_X2 _f_permutation__round__U6698  ( .A(_f_permutation__round_in[1451]), 
        .B(_f_permutation__round_in[1131]), .Z(_f_permutation__round__n1260 )
         );
  XOR2_X2 _f_permutation__round__U6697  ( .A(_f_permutation__round__n1985 ), 
        .B(_f_permutation__round__n2437 ), .Z(_f_permutation__round__n1987 )
         );
  XOR2_X2 _f_permutation__round__U6696  ( .A(SYNOPSYS_UNCONNECTED_852), .B(
        _f_permutation__round__n1987 ), .Z(_f_permutation__round__c[620] ) );
  XOR2_X2 _f_permutation__round__U6695  ( .A(SYNOPSYS_UNCONNECTED_723), .B(
        _f_permutation__round__n1986 ), .Z(_f_permutation__round__c[1517] ) );
  XOR2_X2 _f_permutation__round__U6694  ( .A(SYNOPSYS_UNCONNECTED_532), .B(
        _f_permutation__round__n1987 ), .Z(_f_permutation__round__c[556] ) );
  XOR2_X2 _f_permutation__round__U6693  ( .A(SYNOPSYS_UNCONNECTED_403), .B(
        _f_permutation__round__n1986 ), .Z(_f_permutation__round__c[1453] ) );
  XOR2_X2 _f_permutation__round__U6692  ( .A(SYNOPSYS_UNCONNECTED_212), .B(
        _f_permutation__round__n1987 ), .Z(_f_permutation__round__c[492] ) );
  XOR2_X2 _f_permutation__round__U6691  ( .A(SYNOPSYS_UNCONNECTED_83), .B(
        _f_permutation__round__n1986 ), .Z(_f_permutation__round__c[1389] ) );
  XOR2_X2 _f_permutation__round__U6690  ( .A(_f_permutation__round_in[1196]), 
        .B(_f_permutation__round__n1987 ), .Z(_f_permutation__round__c[428] )
         );
  XOR2_X2 _f_permutation__round__U6689  ( .A(_f_permutation__round_in[1325]), 
        .B(_f_permutation__round__n1986 ), .Z(_f_permutation__round__c[1325] )
         );
  XOR2_X2 _f_permutation__round__U6688  ( .A(_f_permutation__round_in[1516]), 
        .B(_f_permutation__round__n1987 ), .Z(_f_permutation__round__c[364] )
         );
  XOR2_X2 _f_permutation__round__U6687  ( .A(_f_permutation__round__n1262 ), 
        .B(_f_permutation__round__n1261 ), .Z(_f_permutation__round__n2205 )
         );
  XOR2_X2 _f_permutation__round__U6686  ( .A(SYNOPSYS_UNCONNECTED_854), .B(
        _f_permutation__round__n1263 ), .Z(_f_permutation__round__n1261 ) );
  XOR2_X2 _f_permutation__round__U6685  ( .A(SYNOPSYS_UNCONNECTED_214), .B(
        SYNOPSYS_UNCONNECTED_534), .Z(_f_permutation__round__n1262 ) );
  XOR2_X2 _f_permutation__round__U6684  ( .A(_f_permutation__round_in[1514]), 
        .B(_f_permutation__round_in[1194]), .Z(_f_permutation__round__n1263 )
         );
  XOR2_X2 _f_permutation__round__U6683  ( .A(_f_permutation__round__n1265 ), 
        .B(_f_permutation__round__n1264 ), .Z(_f_permutation__round__n2433 )
         );
  XOR2_X2 _f_permutation__round__U6682  ( .A(SYNOPSYS_UNCONNECTED_1045), .B(
        _f_permutation__round__n1266 ), .Z(_f_permutation__round__n1264 ) );
  XOR2_X2 _f_permutation__round__U6681  ( .A(SYNOPSYS_UNCONNECTED_405), .B(
        SYNOPSYS_UNCONNECTED_725), .Z(_f_permutation__round__n1265 ) );
  XOR2_X2 _f_permutation__round__U6680  ( .A(_f_permutation__round_in[1323]), 
        .B(SYNOPSYS_UNCONNECTED_85), .Z(_f_permutation__round__n1266 ) );
  XOR2_X2 _f_permutation__round__U6679  ( .A(_f_permutation__round__n2205 ), 
        .B(_f_permutation__round__n2433 ), .Z(_f_permutation__round__n2206 )
         );
  XOR2_X2 _f_permutation__round__U6678  ( .A(_f_permutation__round_in[1579]), 
        .B(_f_permutation__round__n2206 ), .Z(_f_permutation__round__c[43] )
         );
  XOR2_X2 _f_permutation__round__U6677  ( .A(_f_permutation__round__n1268 ), 
        .B(_f_permutation__round__n1267 ), .Z(_f_permutation__round__n1988 )
         );
  XOR2_X2 _f_permutation__round__U6676  ( .A(SYNOPSYS_UNCONNECTED_789), .B(
        _f_permutation__round__n1269 ), .Z(_f_permutation__round__n1267 ) );
  XOR2_X2 _f_permutation__round__U6675  ( .A(SYNOPSYS_UNCONNECTED_149), .B(
        SYNOPSYS_UNCONNECTED_469), .Z(_f_permutation__round__n1268 ) );
  XOR2_X2 _f_permutation__round__U6674  ( .A(_f_permutation__round_in[1579]), 
        .B(_f_permutation__round_in[1259]), .Z(_f_permutation__round__n1269 )
         );
  XOR2_X2 _f_permutation__round__U6673  ( .A(_f_permutation__round__n1271 ), 
        .B(_f_permutation__round__n1270 ), .Z(_f_permutation__round__n2192 )
         );
  XOR2_X2 _f_permutation__round__U6672  ( .A(SYNOPSYS_UNCONNECTED_980), .B(
        _f_permutation__round__n1272 ), .Z(_f_permutation__round__n1270 ) );
  XOR2_X2 _f_permutation__round__U6671  ( .A(SYNOPSYS_UNCONNECTED_340), .B(
        SYNOPSYS_UNCONNECTED_660), .Z(_f_permutation__round__n1271 ) );
  XOR2_X2 _f_permutation__round__U6670  ( .A(_f_permutation__round_in[1388]), 
        .B(_f_permutation__round_in[1068]), .Z(_f_permutation__round__n1272 )
         );
  XOR2_X2 _f_permutation__round__U6669  ( .A(_f_permutation__round__n1988 ), 
        .B(_f_permutation__round__n2192 ), .Z(_f_permutation__round__n1989 )
         );
  XOR2_X2 _f_permutation__round__U6668  ( .A(SYNOPSYS_UNCONNECTED_1044), .B(
        _f_permutation__round__n1989 ), .Z(_f_permutation__round__c[1580] ) );
  XOR2_X2 _f_permutation__round__U6667  ( .A(_f_permutation__round__n1274 ), 
        .B(_f_permutation__round__n1273 ), .Z(_f_permutation__round__n2440 )
         );
  XOR2_X2 _f_permutation__round__U6666  ( .A(SYNOPSYS_UNCONNECTED_918), .B(
        _f_permutation__round__n1275 ), .Z(_f_permutation__round__n1273 ) );
  XOR2_X2 _f_permutation__round__U6665  ( .A(SYNOPSYS_UNCONNECTED_278), .B(
        SYNOPSYS_UNCONNECTED_598), .Z(_f_permutation__round__n1274 ) );
  XOR2_X2 _f_permutation__round__U6664  ( .A(_f_permutation__round_in[1450]), 
        .B(_f_permutation__round_in[1130]), .Z(_f_permutation__round__n1275 )
         );
  XOR2_X2 _f_permutation__round__U6663  ( .A(_f_permutation__round__n1988 ), 
        .B(_f_permutation__round__n2440 ), .Z(_f_permutation__round__n1990 )
         );
  XOR2_X2 _f_permutation__round__U6662  ( .A(SYNOPSYS_UNCONNECTED_853), .B(
        _f_permutation__round__n1990 ), .Z(_f_permutation__round__c[619] ) );
  XOR2_X2 _f_permutation__round__U6661  ( .A(SYNOPSYS_UNCONNECTED_724), .B(
        _f_permutation__round__n1989 ), .Z(_f_permutation__round__c[1516] ) );
  XOR2_X2 _f_permutation__round__U6660  ( .A(SYNOPSYS_UNCONNECTED_533), .B(
        _f_permutation__round__n1990 ), .Z(_f_permutation__round__c[555] ) );
  XOR2_X2 _f_permutation__round__U6659  ( .A(SYNOPSYS_UNCONNECTED_404), .B(
        _f_permutation__round__n1989 ), .Z(_f_permutation__round__c[1452] ) );
  XOR2_X2 _f_permutation__round__U6658  ( .A(SYNOPSYS_UNCONNECTED_213), .B(
        _f_permutation__round__n1990 ), .Z(_f_permutation__round__c[491] ) );
  XOR2_X2 _f_permutation__round__U6657  ( .A(SYNOPSYS_UNCONNECTED_84), .B(
        _f_permutation__round__n1989 ), .Z(_f_permutation__round__c[1388] ) );
  XOR2_X2 _f_permutation__round__U6656  ( .A(_f_permutation__round_in[1195]), 
        .B(_f_permutation__round__n1990 ), .Z(_f_permutation__round__c[427] )
         );
  XOR2_X2 _f_permutation__round__U6655  ( .A(_f_permutation__round_in[1324]), 
        .B(_f_permutation__round__n1989 ), .Z(_f_permutation__round__c[1324] )
         );
  XOR2_X2 _f_permutation__round__U6654  ( .A(_f_permutation__round_in[1515]), 
        .B(_f_permutation__round__n1990 ), .Z(_f_permutation__round__c[363] )
         );
  XOR2_X2 _f_permutation__round__U6653  ( .A(_f_permutation__round__n1277 ), 
        .B(_f_permutation__round__n1276 ), .Z(_f_permutation__round__n2209 )
         );
  XOR2_X2 _f_permutation__round__U6652  ( .A(SYNOPSYS_UNCONNECTED_855), .B(
        _f_permutation__round__n1278 ), .Z(_f_permutation__round__n1276 ) );
  XOR2_X2 _f_permutation__round__U6651  ( .A(SYNOPSYS_UNCONNECTED_215), .B(
        SYNOPSYS_UNCONNECTED_535), .Z(_f_permutation__round__n1277 ) );
  XOR2_X2 _f_permutation__round__U6650  ( .A(_f_permutation__round_in[1513]), 
        .B(_f_permutation__round_in[1193]), .Z(_f_permutation__round__n1278 )
         );
  XOR2_X2 _f_permutation__round__U6649  ( .A(_f_permutation__round__n1280 ), 
        .B(_f_permutation__round__n1279 ), .Z(_f_permutation__round__n2436 )
         );
  XOR2_X2 _f_permutation__round__U6648  ( .A(SYNOPSYS_UNCONNECTED_1046), .B(
        _f_permutation__round__n1281 ), .Z(_f_permutation__round__n1279 ) );
  XOR2_X2 _f_permutation__round__U6647  ( .A(SYNOPSYS_UNCONNECTED_406), .B(
        SYNOPSYS_UNCONNECTED_726), .Z(_f_permutation__round__n1280 ) );
  XOR2_X2 _f_permutation__round__U6646  ( .A(_f_permutation__round_in[1322]), 
        .B(SYNOPSYS_UNCONNECTED_86), .Z(_f_permutation__round__n1281 ) );
  XOR2_X2 _f_permutation__round__U6645  ( .A(_f_permutation__round__n2209 ), 
        .B(_f_permutation__round__n2436 ), .Z(_f_permutation__round__n2210 )
         );
  XOR2_X2 _f_permutation__round__U6644  ( .A(_f_permutation__round_in[1578]), 
        .B(_f_permutation__round__n2210 ), .Z(_f_permutation__round__c[42] )
         );
  XOR2_X2 _f_permutation__round__U6643  ( .A(_f_permutation__round__n1283 ), 
        .B(_f_permutation__round__n1282 ), .Z(_f_permutation__round__n1991 )
         );
  XOR2_X2 _f_permutation__round__U6642  ( .A(SYNOPSYS_UNCONNECTED_790), .B(
        _f_permutation__round__n1284 ), .Z(_f_permutation__round__n1282 ) );
  XOR2_X2 _f_permutation__round__U6641  ( .A(SYNOPSYS_UNCONNECTED_150), .B(
        SYNOPSYS_UNCONNECTED_470), .Z(_f_permutation__round__n1283 ) );
  XOR2_X2 _f_permutation__round__U6640  ( .A(_f_permutation__round_in[1578]), 
        .B(_f_permutation__round_in[1258]), .Z(_f_permutation__round__n1284 )
         );
  XOR2_X2 _f_permutation__round__U6639  ( .A(_f_permutation__round__n1286 ), 
        .B(_f_permutation__round__n1285 ), .Z(_f_permutation__round__n2196 )
         );
  XOR2_X2 _f_permutation__round__U6638  ( .A(SYNOPSYS_UNCONNECTED_981), .B(
        _f_permutation__round__n1287 ), .Z(_f_permutation__round__n1285 ) );
  XOR2_X2 _f_permutation__round__U6637  ( .A(SYNOPSYS_UNCONNECTED_341), .B(
        SYNOPSYS_UNCONNECTED_661), .Z(_f_permutation__round__n1286 ) );
  XOR2_X2 _f_permutation__round__U6636  ( .A(_f_permutation__round_in[1387]), 
        .B(_f_permutation__round_in[1067]), .Z(_f_permutation__round__n1287 )
         );
  XOR2_X2 _f_permutation__round__U6635  ( .A(_f_permutation__round__n1991 ), 
        .B(_f_permutation__round__n2196 ), .Z(_f_permutation__round__n1992 )
         );
  XOR2_X2 _f_permutation__round__U6634  ( .A(SYNOPSYS_UNCONNECTED_1045), .B(
        _f_permutation__round__n1992 ), .Z(_f_permutation__round__c[1579] ) );
  XOR2_X2 _f_permutation__round__U6633  ( .A(_f_permutation__round__n1289 ), 
        .B(_f_permutation__round__n1288 ), .Z(_f_permutation__round__n2443 )
         );
  XOR2_X2 _f_permutation__round__U6632  ( .A(SYNOPSYS_UNCONNECTED_919), .B(
        _f_permutation__round__n1290 ), .Z(_f_permutation__round__n1288 ) );
  XOR2_X2 _f_permutation__round__U6631  ( .A(SYNOPSYS_UNCONNECTED_279), .B(
        SYNOPSYS_UNCONNECTED_599), .Z(_f_permutation__round__n1289 ) );
  XOR2_X2 _f_permutation__round__U6630  ( .A(_f_permutation__round_in[1449]), 
        .B(_f_permutation__round_in[1129]), .Z(_f_permutation__round__n1290 )
         );
  XOR2_X2 _f_permutation__round__U6629  ( .A(_f_permutation__round__n1991 ), 
        .B(_f_permutation__round__n2443 ), .Z(_f_permutation__round__n1993 )
         );
  XOR2_X2 _f_permutation__round__U6628  ( .A(SYNOPSYS_UNCONNECTED_854), .B(
        _f_permutation__round__n1993 ), .Z(_f_permutation__round__c[618] ) );
  XOR2_X2 _f_permutation__round__U6627  ( .A(SYNOPSYS_UNCONNECTED_725), .B(
        _f_permutation__round__n1992 ), .Z(_f_permutation__round__c[1515] ) );
  XOR2_X2 _f_permutation__round__U6626  ( .A(SYNOPSYS_UNCONNECTED_534), .B(
        _f_permutation__round__n1993 ), .Z(_f_permutation__round__c[554] ) );
  XOR2_X2 _f_permutation__round__U6625  ( .A(SYNOPSYS_UNCONNECTED_405), .B(
        _f_permutation__round__n1992 ), .Z(_f_permutation__round__c[1451] ) );
  XOR2_X2 _f_permutation__round__U6624  ( .A(SYNOPSYS_UNCONNECTED_214), .B(
        _f_permutation__round__n1993 ), .Z(_f_permutation__round__c[490] ) );
  XOR2_X2 _f_permutation__round__U6623  ( .A(SYNOPSYS_UNCONNECTED_85), .B(
        _f_permutation__round__n1992 ), .Z(_f_permutation__round__c[1387] ) );
  XOR2_X2 _f_permutation__round__U6622  ( .A(_f_permutation__round_in[1194]), 
        .B(_f_permutation__round__n1993 ), .Z(_f_permutation__round__c[426] )
         );
  XOR2_X2 _f_permutation__round__U6621  ( .A(_f_permutation__round_in[1323]), 
        .B(_f_permutation__round__n1992 ), .Z(_f_permutation__round__c[1323] )
         );
  XOR2_X2 _f_permutation__round__U6620  ( .A(_f_permutation__round_in[1514]), 
        .B(_f_permutation__round__n1993 ), .Z(_f_permutation__round__c[362] )
         );
  XOR2_X2 _f_permutation__round__U6619  ( .A(_f_permutation__round__n1292 ), 
        .B(_f_permutation__round__n1291 ), .Z(_f_permutation__round__n2213 )
         );
  XOR2_X2 _f_permutation__round__U6618  ( .A(SYNOPSYS_UNCONNECTED_856), .B(
        _f_permutation__round__n1293 ), .Z(_f_permutation__round__n1291 ) );
  XOR2_X2 _f_permutation__round__U6617  ( .A(SYNOPSYS_UNCONNECTED_216), .B(
        SYNOPSYS_UNCONNECTED_536), .Z(_f_permutation__round__n1292 ) );
  XOR2_X2 _f_permutation__round__U6616  ( .A(_f_permutation__round_in[1512]), 
        .B(_f_permutation__round_in[1192]), .Z(_f_permutation__round__n1293 )
         );
  XOR2_X2 _f_permutation__round__U6615  ( .A(_f_permutation__round__n1295 ), 
        .B(_f_permutation__round__n1294 ), .Z(_f_permutation__round__n2439 )
         );
  XOR2_X2 _f_permutation__round__U6614  ( .A(SYNOPSYS_UNCONNECTED_1047), .B(
        _f_permutation__round__n1296 ), .Z(_f_permutation__round__n1294 ) );
  XOR2_X2 _f_permutation__round__U6613  ( .A(SYNOPSYS_UNCONNECTED_407), .B(
        SYNOPSYS_UNCONNECTED_727), .Z(_f_permutation__round__n1295 ) );
  XOR2_X2 _f_permutation__round__U6612  ( .A(_f_permutation__round_in[1321]), 
        .B(SYNOPSYS_UNCONNECTED_87), .Z(_f_permutation__round__n1296 ) );
  XOR2_X2 _f_permutation__round__U6611  ( .A(_f_permutation__round__n2213 ), 
        .B(_f_permutation__round__n2439 ), .Z(_f_permutation__round__n2214 )
         );
  XOR2_X2 _f_permutation__round__U6610  ( .A(_f_permutation__round_in[1577]), 
        .B(_f_permutation__round__n2214 ), .Z(_f_permutation__round__c[41] )
         );
  XOR2_X2 _f_permutation__round__U6609  ( .A(_f_permutation__round__n1298 ), 
        .B(_f_permutation__round__n1297 ), .Z(_f_permutation__round__n1994 )
         );
  XOR2_X2 _f_permutation__round__U6608  ( .A(SYNOPSYS_UNCONNECTED_791), .B(
        _f_permutation__round__n1299 ), .Z(_f_permutation__round__n1297 ) );
  XOR2_X2 _f_permutation__round__U6607  ( .A(SYNOPSYS_UNCONNECTED_151), .B(
        SYNOPSYS_UNCONNECTED_471), .Z(_f_permutation__round__n1298 ) );
  XOR2_X2 _f_permutation__round__U6606  ( .A(_f_permutation__round_in[1577]), 
        .B(_f_permutation__round_in[1257]), .Z(_f_permutation__round__n1299 )
         );
  XOR2_X2 _f_permutation__round__U6605  ( .A(_f_permutation__round__n1301 ), 
        .B(_f_permutation__round__n1300 ), .Z(_f_permutation__round__n2200 )
         );
  XOR2_X2 _f_permutation__round__U6604  ( .A(SYNOPSYS_UNCONNECTED_982), .B(
        _f_permutation__round__n1302 ), .Z(_f_permutation__round__n1300 ) );
  XOR2_X2 _f_permutation__round__U6603  ( .A(SYNOPSYS_UNCONNECTED_342), .B(
        SYNOPSYS_UNCONNECTED_662), .Z(_f_permutation__round__n1301 ) );
  XOR2_X2 _f_permutation__round__U6602  ( .A(_f_permutation__round_in[1386]), 
        .B(_f_permutation__round_in[1066]), .Z(_f_permutation__round__n1302 )
         );
  XOR2_X2 _f_permutation__round__U6601  ( .A(_f_permutation__round__n1994 ), 
        .B(_f_permutation__round__n2200 ), .Z(_f_permutation__round__n1995 )
         );
  XOR2_X2 _f_permutation__round__U6600  ( .A(SYNOPSYS_UNCONNECTED_1046), .B(
        _f_permutation__round__n1995 ), .Z(_f_permutation__round__c[1578] ) );
  XOR2_X2 _f_permutation__round__U6599  ( .A(_f_permutation__round__n1304 ), 
        .B(_f_permutation__round__n1303 ), .Z(_f_permutation__round__n2446 )
         );
  XOR2_X2 _f_permutation__round__U6598  ( .A(SYNOPSYS_UNCONNECTED_920), .B(
        _f_permutation__round__n1305 ), .Z(_f_permutation__round__n1303 ) );
  XOR2_X2 _f_permutation__round__U6597  ( .A(SYNOPSYS_UNCONNECTED_280), .B(
        SYNOPSYS_UNCONNECTED_600), .Z(_f_permutation__round__n1304 ) );
  XOR2_X2 _f_permutation__round__U6596  ( .A(_f_permutation__round_in[1448]), 
        .B(_f_permutation__round_in[1128]), .Z(_f_permutation__round__n1305 )
         );
  XOR2_X2 _f_permutation__round__U6595  ( .A(_f_permutation__round__n1994 ), 
        .B(_f_permutation__round__n2446 ), .Z(_f_permutation__round__n1996 )
         );
  XOR2_X2 _f_permutation__round__U6594  ( .A(SYNOPSYS_UNCONNECTED_855), .B(
        _f_permutation__round__n1996 ), .Z(_f_permutation__round__c[617] ) );
  XOR2_X2 _f_permutation__round__U6593  ( .A(SYNOPSYS_UNCONNECTED_726), .B(
        _f_permutation__round__n1995 ), .Z(_f_permutation__round__c[1514] ) );
  XOR2_X2 _f_permutation__round__U6592  ( .A(SYNOPSYS_UNCONNECTED_535), .B(
        _f_permutation__round__n1996 ), .Z(_f_permutation__round__c[553] ) );
  XOR2_X2 _f_permutation__round__U6591  ( .A(SYNOPSYS_UNCONNECTED_406), .B(
        _f_permutation__round__n1995 ), .Z(_f_permutation__round__c[1450] ) );
  XOR2_X2 _f_permutation__round__U6590  ( .A(SYNOPSYS_UNCONNECTED_215), .B(
        _f_permutation__round__n1996 ), .Z(_f_permutation__round__c[489] ) );
  XOR2_X2 _f_permutation__round__U6589  ( .A(SYNOPSYS_UNCONNECTED_86), .B(
        _f_permutation__round__n1995 ), .Z(_f_permutation__round__c[1386] ) );
  XOR2_X2 _f_permutation__round__U6588  ( .A(_f_permutation__round_in[1193]), 
        .B(_f_permutation__round__n1996 ), .Z(_f_permutation__round__c[425] )
         );
  XOR2_X2 _f_permutation__round__U6587  ( .A(_f_permutation__round_in[1322]), 
        .B(_f_permutation__round__n1995 ), .Z(_f_permutation__round__c[1322] )
         );
  XOR2_X2 _f_permutation__round__U6586  ( .A(_f_permutation__round_in[1513]), 
        .B(_f_permutation__round__n1996 ), .Z(_f_permutation__round__c[361] )
         );
  XOR2_X2 _f_permutation__round__U6585  ( .A(_f_permutation__round__n1307 ), 
        .B(_f_permutation__round__n1306 ), .Z(_f_permutation__round__n2217 )
         );
  XOR2_X2 _f_permutation__round__U6584  ( .A(SYNOPSYS_UNCONNECTED_857), .B(
        _f_permutation__round__n1308 ), .Z(_f_permutation__round__n1306 ) );
  XOR2_X2 _f_permutation__round__U6583  ( .A(SYNOPSYS_UNCONNECTED_217), .B(
        SYNOPSYS_UNCONNECTED_537), .Z(_f_permutation__round__n1307 ) );
  XOR2_X2 _f_permutation__round__U6582  ( .A(_f_permutation__round_in[1511]), 
        .B(_f_permutation__round_in[1191]), .Z(_f_permutation__round__n1308 )
         );
  XOR2_X2 _f_permutation__round__U6581  ( .A(_f_permutation__round__n1310 ), 
        .B(_f_permutation__round__n1309 ), .Z(_f_permutation__round__n2442 )
         );
  XOR2_X2 _f_permutation__round__U6580  ( .A(SYNOPSYS_UNCONNECTED_1048), .B(
        _f_permutation__round__n1311 ), .Z(_f_permutation__round__n1309 ) );
  XOR2_X2 _f_permutation__round__U6579  ( .A(SYNOPSYS_UNCONNECTED_408), .B(
        SYNOPSYS_UNCONNECTED_728), .Z(_f_permutation__round__n1310 ) );
  XOR2_X2 _f_permutation__round__U6578  ( .A(_f_permutation__round_in[1320]), 
        .B(SYNOPSYS_UNCONNECTED_88), .Z(_f_permutation__round__n1311 ) );
  XOR2_X2 _f_permutation__round__U6577  ( .A(_f_permutation__round__n2217 ), 
        .B(_f_permutation__round__n2442 ), .Z(_f_permutation__round__n2218 )
         );
  XOR2_X2 _f_permutation__round__U6576  ( .A(_f_permutation__round_in[1576]), 
        .B(_f_permutation__round__n2218 ), .Z(_f_permutation__round__c[40] )
         );
  XOR2_X2 _f_permutation__round__U6575  ( .A(_f_permutation__round__n1313 ), 
        .B(_f_permutation__round__n1312 ), .Z(_f_permutation__round__n1997 )
         );
  XOR2_X2 _f_permutation__round__U6574  ( .A(SYNOPSYS_UNCONNECTED_792), .B(
        _f_permutation__round__n1314 ), .Z(_f_permutation__round__n1312 ) );
  XOR2_X2 _f_permutation__round__U6573  ( .A(SYNOPSYS_UNCONNECTED_152), .B(
        SYNOPSYS_UNCONNECTED_472), .Z(_f_permutation__round__n1313 ) );
  XOR2_X2 _f_permutation__round__U6572  ( .A(_f_permutation__round_in[1576]), 
        .B(_f_permutation__round_in[1256]), .Z(_f_permutation__round__n1314 )
         );
  XOR2_X2 _f_permutation__round__U6571  ( .A(_f_permutation__round__n1316 ), 
        .B(_f_permutation__round__n1315 ), .Z(_f_permutation__round__n2204 )
         );
  XOR2_X2 _f_permutation__round__U6570  ( .A(SYNOPSYS_UNCONNECTED_983), .B(
        _f_permutation__round__n1317 ), .Z(_f_permutation__round__n1315 ) );
  XOR2_X2 _f_permutation__round__U6569  ( .A(SYNOPSYS_UNCONNECTED_343), .B(
        SYNOPSYS_UNCONNECTED_663), .Z(_f_permutation__round__n1316 ) );
  XOR2_X2 _f_permutation__round__U6568  ( .A(_f_permutation__round_in[1385]), 
        .B(_f_permutation__round_in[1065]), .Z(_f_permutation__round__n1317 )
         );
  XOR2_X2 _f_permutation__round__U6567  ( .A(_f_permutation__round__n1997 ), 
        .B(_f_permutation__round__n2204 ), .Z(_f_permutation__round__n1998 )
         );
  XOR2_X2 _f_permutation__round__U6566  ( .A(SYNOPSYS_UNCONNECTED_1047), .B(
        _f_permutation__round__n1998 ), .Z(_f_permutation__round__c[1577] ) );
  XOR2_X2 _f_permutation__round__U6565  ( .A(_f_permutation__round__n1319 ), 
        .B(_f_permutation__round__n1318 ), .Z(_f_permutation__round__n2449 )
         );
  XOR2_X2 _f_permutation__round__U6564  ( .A(SYNOPSYS_UNCONNECTED_921), .B(
        _f_permutation__round__n1320 ), .Z(_f_permutation__round__n1318 ) );
  XOR2_X2 _f_permutation__round__U6563  ( .A(SYNOPSYS_UNCONNECTED_281), .B(
        SYNOPSYS_UNCONNECTED_601), .Z(_f_permutation__round__n1319 ) );
  XOR2_X2 _f_permutation__round__U6562  ( .A(_f_permutation__round_in[1447]), 
        .B(_f_permutation__round_in[1127]), .Z(_f_permutation__round__n1320 )
         );
  XOR2_X2 _f_permutation__round__U6561  ( .A(_f_permutation__round__n1997 ), 
        .B(_f_permutation__round__n2449 ), .Z(_f_permutation__round__n1999 )
         );
  XOR2_X2 _f_permutation__round__U6560  ( .A(SYNOPSYS_UNCONNECTED_856), .B(
        _f_permutation__round__n1999 ), .Z(_f_permutation__round__c[616] ) );
  XOR2_X2 _f_permutation__round__U6559  ( .A(SYNOPSYS_UNCONNECTED_727), .B(
        _f_permutation__round__n1998 ), .Z(_f_permutation__round__c[1513] ) );
  XOR2_X2 _f_permutation__round__U6558  ( .A(SYNOPSYS_UNCONNECTED_536), .B(
        _f_permutation__round__n1999 ), .Z(_f_permutation__round__c[552] ) );
  XOR2_X2 _f_permutation__round__U6557  ( .A(SYNOPSYS_UNCONNECTED_407), .B(
        _f_permutation__round__n1998 ), .Z(_f_permutation__round__c[1449] ) );
  XOR2_X2 _f_permutation__round__U6556  ( .A(SYNOPSYS_UNCONNECTED_216), .B(
        _f_permutation__round__n1999 ), .Z(_f_permutation__round__c[488] ) );
  XOR2_X2 _f_permutation__round__U6555  ( .A(SYNOPSYS_UNCONNECTED_87), .B(
        _f_permutation__round__n1998 ), .Z(_f_permutation__round__c[1385] ) );
  XOR2_X2 _f_permutation__round__U6554  ( .A(_f_permutation__round_in[1192]), 
        .B(_f_permutation__round__n1999 ), .Z(_f_permutation__round__c[424] )
         );
  XOR2_X2 _f_permutation__round__U6553  ( .A(_f_permutation__round_in[1321]), 
        .B(_f_permutation__round__n1998 ), .Z(_f_permutation__round__c[1321] )
         );
  XOR2_X2 _f_permutation__round__U6552  ( .A(_f_permutation__round_in[1512]), 
        .B(_f_permutation__round__n1999 ), .Z(_f_permutation__round__c[360] )
         );
  XOR2_X2 _f_permutation__round__U6551  ( .A(_f_permutation__round__n1322 ), 
        .B(_f_permutation__round__n1321 ), .Z(_f_permutation__round__n2221 )
         );
  XOR2_X2 _f_permutation__round__U6550  ( .A(SYNOPSYS_UNCONNECTED_858), .B(
        _f_permutation__round__n1323 ), .Z(_f_permutation__round__n1321 ) );
  XOR2_X2 _f_permutation__round__U6549  ( .A(SYNOPSYS_UNCONNECTED_218), .B(
        SYNOPSYS_UNCONNECTED_538), .Z(_f_permutation__round__n1322 ) );
  XOR2_X2 _f_permutation__round__U6548  ( .A(_f_permutation__round_in[1510]), 
        .B(_f_permutation__round_in[1190]), .Z(_f_permutation__round__n1323 )
         );
  XOR2_X2 _f_permutation__round__U6547  ( .A(_f_permutation__round__n1325 ), 
        .B(_f_permutation__round__n1324 ), .Z(_f_permutation__round__n2445 )
         );
  XOR2_X2 _f_permutation__round__U6546  ( .A(SYNOPSYS_UNCONNECTED_1049), .B(
        _f_permutation__round__n1326 ), .Z(_f_permutation__round__n1324 ) );
  XOR2_X2 _f_permutation__round__U6545  ( .A(SYNOPSYS_UNCONNECTED_409), .B(
        SYNOPSYS_UNCONNECTED_729), .Z(_f_permutation__round__n1325 ) );
  XOR2_X2 _f_permutation__round__U6544  ( .A(_f_permutation__round_in[1319]), 
        .B(SYNOPSYS_UNCONNECTED_89), .Z(_f_permutation__round__n1326 ) );
  XOR2_X2 _f_permutation__round__U6543  ( .A(_f_permutation__round__n2221 ), 
        .B(_f_permutation__round__n2445 ), .Z(_f_permutation__round__n2222 )
         );
  XOR2_X2 _f_permutation__round__U6542  ( .A(_f_permutation__round_in[1575]), 
        .B(_f_permutation__round__n2222 ), .Z(_f_permutation__round__c[39] )
         );
  XOR2_X2 _f_permutation__round__U6541  ( .A(_f_permutation__round__n1328 ), 
        .B(_f_permutation__round__n1327 ), .Z(_f_permutation__round__n2000 )
         );
  XOR2_X2 _f_permutation__round__U6540  ( .A(SYNOPSYS_UNCONNECTED_793), .B(
        _f_permutation__round__n1329 ), .Z(_f_permutation__round__n1327 ) );
  XOR2_X2 _f_permutation__round__U6539  ( .A(SYNOPSYS_UNCONNECTED_153), .B(
        SYNOPSYS_UNCONNECTED_473), .Z(_f_permutation__round__n1328 ) );
  XOR2_X2 _f_permutation__round__U6538  ( .A(_f_permutation__round_in[1575]), 
        .B(_f_permutation__round_in[1255]), .Z(_f_permutation__round__n1329 )
         );
  XOR2_X2 _f_permutation__round__U6537  ( .A(_f_permutation__round__n1331 ), 
        .B(_f_permutation__round__n1330 ), .Z(_f_permutation__round__n2208 )
         );
  XOR2_X2 _f_permutation__round__U6536  ( .A(SYNOPSYS_UNCONNECTED_984), .B(
        _f_permutation__round__n1332 ), .Z(_f_permutation__round__n1330 ) );
  XOR2_X2 _f_permutation__round__U6535  ( .A(SYNOPSYS_UNCONNECTED_344), .B(
        SYNOPSYS_UNCONNECTED_664), .Z(_f_permutation__round__n1331 ) );
  XOR2_X2 _f_permutation__round__U6534  ( .A(_f_permutation__round_in[1384]), 
        .B(_f_permutation__round_in[1064]), .Z(_f_permutation__round__n1332 )
         );
  XOR2_X2 _f_permutation__round__U6533  ( .A(_f_permutation__round__n2000 ), 
        .B(_f_permutation__round__n2208 ), .Z(_f_permutation__round__n2001 )
         );
  XOR2_X2 _f_permutation__round__U6532  ( .A(SYNOPSYS_UNCONNECTED_1048), .B(
        _f_permutation__round__n2001 ), .Z(_f_permutation__round__c[1576] ) );
  XOR2_X2 _f_permutation__round__U6531  ( .A(_f_permutation__round__n1334 ), 
        .B(_f_permutation__round__n1333 ), .Z(_f_permutation__round__n2452 )
         );
  XOR2_X2 _f_permutation__round__U6530  ( .A(SYNOPSYS_UNCONNECTED_922), .B(
        _f_permutation__round__n1335 ), .Z(_f_permutation__round__n1333 ) );
  XOR2_X2 _f_permutation__round__U6529  ( .A(SYNOPSYS_UNCONNECTED_282), .B(
        SYNOPSYS_UNCONNECTED_602), .Z(_f_permutation__round__n1334 ) );
  XOR2_X2 _f_permutation__round__U6528  ( .A(_f_permutation__round_in[1446]), 
        .B(_f_permutation__round_in[1126]), .Z(_f_permutation__round__n1335 )
         );
  XOR2_X2 _f_permutation__round__U6527  ( .A(_f_permutation__round__n2000 ), 
        .B(_f_permutation__round__n2452 ), .Z(_f_permutation__round__n2002 )
         );
  XOR2_X2 _f_permutation__round__U6526  ( .A(SYNOPSYS_UNCONNECTED_857), .B(
        _f_permutation__round__n2002 ), .Z(_f_permutation__round__c[615] ) );
  XOR2_X2 _f_permutation__round__U6525  ( .A(SYNOPSYS_UNCONNECTED_728), .B(
        _f_permutation__round__n2001 ), .Z(_f_permutation__round__c[1512] ) );
  XOR2_X2 _f_permutation__round__U6524  ( .A(SYNOPSYS_UNCONNECTED_537), .B(
        _f_permutation__round__n2002 ), .Z(_f_permutation__round__c[551] ) );
  XOR2_X2 _f_permutation__round__U6523  ( .A(SYNOPSYS_UNCONNECTED_408), .B(
        _f_permutation__round__n2001 ), .Z(_f_permutation__round__c[1448] ) );
  XOR2_X2 _f_permutation__round__U6522  ( .A(SYNOPSYS_UNCONNECTED_217), .B(
        _f_permutation__round__n2002 ), .Z(_f_permutation__round__c[487] ) );
  XOR2_X2 _f_permutation__round__U6521  ( .A(SYNOPSYS_UNCONNECTED_88), .B(
        _f_permutation__round__n2001 ), .Z(_f_permutation__round__c[1384] ) );
  XOR2_X2 _f_permutation__round__U6520  ( .A(_f_permutation__round_in[1191]), 
        .B(_f_permutation__round__n2002 ), .Z(_f_permutation__round__c[423] )
         );
  XOR2_X2 _f_permutation__round__U6519  ( .A(_f_permutation__round_in[1320]), 
        .B(_f_permutation__round__n2001 ), .Z(_f_permutation__round__c[1320] )
         );
  XOR2_X2 _f_permutation__round__U6518  ( .A(_f_permutation__round_in[1511]), 
        .B(_f_permutation__round__n2002 ), .Z(_f_permutation__round__c[359] )
         );
  XOR2_X2 _f_permutation__round__U6517  ( .A(_f_permutation__round__n1337 ), 
        .B(_f_permutation__round__n1336 ), .Z(_f_permutation__round__n2225 )
         );
  XOR2_X2 _f_permutation__round__U6516  ( .A(SYNOPSYS_UNCONNECTED_859), .B(
        _f_permutation__round__n1338 ), .Z(_f_permutation__round__n1336 ) );
  XOR2_X2 _f_permutation__round__U6515  ( .A(SYNOPSYS_UNCONNECTED_219), .B(
        SYNOPSYS_UNCONNECTED_539), .Z(_f_permutation__round__n1337 ) );
  XOR2_X2 _f_permutation__round__U6514  ( .A(_f_permutation__round_in[1509]), 
        .B(_f_permutation__round_in[1189]), .Z(_f_permutation__round__n1338 )
         );
  XOR2_X2 _f_permutation__round__U6513  ( .A(_f_permutation__round__n1340 ), 
        .B(_f_permutation__round__n1339 ), .Z(_f_permutation__round__n2448 )
         );
  XOR2_X2 _f_permutation__round__U6512  ( .A(SYNOPSYS_UNCONNECTED_1050), .B(
        _f_permutation__round__n1341 ), .Z(_f_permutation__round__n1339 ) );
  XOR2_X2 _f_permutation__round__U6511  ( .A(SYNOPSYS_UNCONNECTED_410), .B(
        SYNOPSYS_UNCONNECTED_730), .Z(_f_permutation__round__n1340 ) );
  XOR2_X2 _f_permutation__round__U6510  ( .A(_f_permutation__round_in[1318]), 
        .B(SYNOPSYS_UNCONNECTED_90), .Z(_f_permutation__round__n1341 ) );
  XOR2_X2 _f_permutation__round__U6509  ( .A(_f_permutation__round__n2225 ), 
        .B(_f_permutation__round__n2448 ), .Z(_f_permutation__round__n2226 )
         );
  XOR2_X2 _f_permutation__round__U6508  ( .A(_f_permutation__round_in[1574]), 
        .B(_f_permutation__round__n2226 ), .Z(_f_permutation__round__c[38] )
         );
  XOR2_X2 _f_permutation__round__U6507  ( .A(_f_permutation__round__n1343 ), 
        .B(_f_permutation__round__n1342 ), .Z(_f_permutation__round__n2003 )
         );
  XOR2_X2 _f_permutation__round__U6506  ( .A(SYNOPSYS_UNCONNECTED_794), .B(
        _f_permutation__round__n1344 ), .Z(_f_permutation__round__n1342 ) );
  XOR2_X2 _f_permutation__round__U6505  ( .A(SYNOPSYS_UNCONNECTED_154), .B(
        SYNOPSYS_UNCONNECTED_474), .Z(_f_permutation__round__n1343 ) );
  XOR2_X2 _f_permutation__round__U6504  ( .A(_f_permutation__round_in[1574]), 
        .B(_f_permutation__round_in[1254]), .Z(_f_permutation__round__n1344 )
         );
  XOR2_X2 _f_permutation__round__U6503  ( .A(_f_permutation__round__n1346 ), 
        .B(_f_permutation__round__n1345 ), .Z(_f_permutation__round__n2212 )
         );
  XOR2_X2 _f_permutation__round__U6502  ( .A(SYNOPSYS_UNCONNECTED_985), .B(
        _f_permutation__round__n1347 ), .Z(_f_permutation__round__n1345 ) );
  XOR2_X2 _f_permutation__round__U6501  ( .A(SYNOPSYS_UNCONNECTED_345), .B(
        SYNOPSYS_UNCONNECTED_665), .Z(_f_permutation__round__n1346 ) );
  XOR2_X2 _f_permutation__round__U6500  ( .A(_f_permutation__round_in[1383]), 
        .B(_f_permutation__round_in[1063]), .Z(_f_permutation__round__n1347 )
         );
  XOR2_X2 _f_permutation__round__U6499  ( .A(_f_permutation__round__n2003 ), 
        .B(_f_permutation__round__n2212 ), .Z(_f_permutation__round__n2004 )
         );
  XOR2_X2 _f_permutation__round__U6498  ( .A(SYNOPSYS_UNCONNECTED_1049), .B(
        _f_permutation__round__n2004 ), .Z(_f_permutation__round__c[1575] ) );
  XOR2_X2 _f_permutation__round__U6497  ( .A(_f_permutation__round__n1349 ), 
        .B(_f_permutation__round__n1348 ), .Z(_f_permutation__round__n2455 )
         );
  XOR2_X2 _f_permutation__round__U6496  ( .A(SYNOPSYS_UNCONNECTED_923), .B(
        _f_permutation__round__n1350 ), .Z(_f_permutation__round__n1348 ) );
  XOR2_X2 _f_permutation__round__U6495  ( .A(SYNOPSYS_UNCONNECTED_283), .B(
        SYNOPSYS_UNCONNECTED_603), .Z(_f_permutation__round__n1349 ) );
  XOR2_X2 _f_permutation__round__U6494  ( .A(_f_permutation__round_in[1445]), 
        .B(_f_permutation__round_in[1125]), .Z(_f_permutation__round__n1350 )
         );
  XOR2_X2 _f_permutation__round__U6493  ( .A(_f_permutation__round__n2003 ), 
        .B(_f_permutation__round__n2455 ), .Z(_f_permutation__round__n2005 )
         );
  XOR2_X2 _f_permutation__round__U6492  ( .A(SYNOPSYS_UNCONNECTED_858), .B(
        _f_permutation__round__n2005 ), .Z(_f_permutation__round__c[614] ) );
  XOR2_X2 _f_permutation__round__U6491  ( .A(SYNOPSYS_UNCONNECTED_729), .B(
        _f_permutation__round__n2004 ), .Z(_f_permutation__round__c[1511] ) );
  XOR2_X2 _f_permutation__round__U6490  ( .A(SYNOPSYS_UNCONNECTED_538), .B(
        _f_permutation__round__n2005 ), .Z(_f_permutation__round__c[550] ) );
  XOR2_X2 _f_permutation__round__U6489  ( .A(SYNOPSYS_UNCONNECTED_409), .B(
        _f_permutation__round__n2004 ), .Z(_f_permutation__round__c[1447] ) );
  XOR2_X2 _f_permutation__round__U6488  ( .A(SYNOPSYS_UNCONNECTED_218), .B(
        _f_permutation__round__n2005 ), .Z(_f_permutation__round__c[486] ) );
  XOR2_X2 _f_permutation__round__U6487  ( .A(SYNOPSYS_UNCONNECTED_89), .B(
        _f_permutation__round__n2004 ), .Z(_f_permutation__round__c[1383] ) );
  XOR2_X2 _f_permutation__round__U6486  ( .A(_f_permutation__round_in[1190]), 
        .B(_f_permutation__round__n2005 ), .Z(_f_permutation__round__c[422] )
         );
  XOR2_X2 _f_permutation__round__U6485  ( .A(_f_permutation__round_in[1319]), 
        .B(_f_permutation__round__n2004 ), .Z(_f_permutation__round__c[1319] )
         );
  XOR2_X2 _f_permutation__round__U6484  ( .A(_f_permutation__round_in[1510]), 
        .B(_f_permutation__round__n2005 ), .Z(_f_permutation__round__c[358] )
         );
  XOR2_X2 _f_permutation__round__U6483  ( .A(_f_permutation__round__n1352 ), 
        .B(_f_permutation__round__n1351 ), .Z(_f_permutation__round__n2229 )
         );
  XOR2_X2 _f_permutation__round__U6482  ( .A(SYNOPSYS_UNCONNECTED_860), .B(
        _f_permutation__round__n1353 ), .Z(_f_permutation__round__n1351 ) );
  XOR2_X2 _f_permutation__round__U6481  ( .A(SYNOPSYS_UNCONNECTED_220), .B(
        SYNOPSYS_UNCONNECTED_540), .Z(_f_permutation__round__n1352 ) );
  XOR2_X2 _f_permutation__round__U6480  ( .A(_f_permutation__round_in[1508]), 
        .B(_f_permutation__round_in[1188]), .Z(_f_permutation__round__n1353 )
         );
  XOR2_X2 _f_permutation__round__U6479  ( .A(_f_permutation__round__n1355 ), 
        .B(_f_permutation__round__n1354 ), .Z(_f_permutation__round__n2451 )
         );
  XOR2_X2 _f_permutation__round__U6478  ( .A(SYNOPSYS_UNCONNECTED_1051), .B(
        _f_permutation__round__n1356 ), .Z(_f_permutation__round__n1354 ) );
  XOR2_X2 _f_permutation__round__U6477  ( .A(SYNOPSYS_UNCONNECTED_411), .B(
        SYNOPSYS_UNCONNECTED_731), .Z(_f_permutation__round__n1355 ) );
  XOR2_X2 _f_permutation__round__U6476  ( .A(_f_permutation__round_in[1317]), 
        .B(SYNOPSYS_UNCONNECTED_91), .Z(_f_permutation__round__n1356 ) );
  XOR2_X2 _f_permutation__round__U6475  ( .A(_f_permutation__round__n2229 ), 
        .B(_f_permutation__round__n2451 ), .Z(_f_permutation__round__n2230 )
         );
  XOR2_X2 _f_permutation__round__U6474  ( .A(_f_permutation__round_in[1573]), 
        .B(_f_permutation__round__n2230 ), .Z(_f_permutation__round__c[37] )
         );
  XOR2_X2 _f_permutation__round__U6473  ( .A(_f_permutation__round__n1358 ), 
        .B(_f_permutation__round__n1357 ), .Z(_f_permutation__round__n2006 )
         );
  XOR2_X2 _f_permutation__round__U6472  ( .A(SYNOPSYS_UNCONNECTED_795), .B(
        _f_permutation__round__n1359 ), .Z(_f_permutation__round__n1357 ) );
  XOR2_X2 _f_permutation__round__U6471  ( .A(SYNOPSYS_UNCONNECTED_155), .B(
        SYNOPSYS_UNCONNECTED_475), .Z(_f_permutation__round__n1358 ) );
  XOR2_X2 _f_permutation__round__U6470  ( .A(_f_permutation__round_in[1573]), 
        .B(_f_permutation__round_in[1253]), .Z(_f_permutation__round__n1359 )
         );
  XOR2_X2 _f_permutation__round__U6469  ( .A(_f_permutation__round__n1361 ), 
        .B(_f_permutation__round__n1360 ), .Z(_f_permutation__round__n2216 )
         );
  XOR2_X2 _f_permutation__round__U6468  ( .A(SYNOPSYS_UNCONNECTED_986), .B(
        _f_permutation__round__n1362 ), .Z(_f_permutation__round__n1360 ) );
  XOR2_X2 _f_permutation__round__U6467  ( .A(SYNOPSYS_UNCONNECTED_346), .B(
        SYNOPSYS_UNCONNECTED_666), .Z(_f_permutation__round__n1361 ) );
  XOR2_X2 _f_permutation__round__U6466  ( .A(_f_permutation__round_in[1382]), 
        .B(_f_permutation__round_in[1062]), .Z(_f_permutation__round__n1362 )
         );
  XOR2_X2 _f_permutation__round__U6465  ( .A(_f_permutation__round__n2006 ), 
        .B(_f_permutation__round__n2216 ), .Z(_f_permutation__round__n2007 )
         );
  XOR2_X2 _f_permutation__round__U6464  ( .A(SYNOPSYS_UNCONNECTED_1050), .B(
        _f_permutation__round__n2007 ), .Z(_f_permutation__round__c[1574] ) );
  XOR2_X2 _f_permutation__round__U6463  ( .A(_f_permutation__round__n1364 ), 
        .B(_f_permutation__round__n1363 ), .Z(_f_permutation__round__n2458 )
         );
  XOR2_X2 _f_permutation__round__U6462  ( .A(SYNOPSYS_UNCONNECTED_924), .B(
        _f_permutation__round__n1365 ), .Z(_f_permutation__round__n1363 ) );
  XOR2_X2 _f_permutation__round__U6461  ( .A(SYNOPSYS_UNCONNECTED_284), .B(
        SYNOPSYS_UNCONNECTED_604), .Z(_f_permutation__round__n1364 ) );
  XOR2_X2 _f_permutation__round__U6460  ( .A(_f_permutation__round_in[1444]), 
        .B(_f_permutation__round_in[1124]), .Z(_f_permutation__round__n1365 )
         );
  XOR2_X2 _f_permutation__round__U6459  ( .A(_f_permutation__round__n2006 ), 
        .B(_f_permutation__round__n2458 ), .Z(_f_permutation__round__n2008 )
         );
  XOR2_X2 _f_permutation__round__U6458  ( .A(SYNOPSYS_UNCONNECTED_859), .B(
        _f_permutation__round__n2008 ), .Z(_f_permutation__round__c[613] ) );
  XOR2_X2 _f_permutation__round__U6457  ( .A(SYNOPSYS_UNCONNECTED_730), .B(
        _f_permutation__round__n2007 ), .Z(_f_permutation__round__c[1510] ) );
  XOR2_X2 _f_permutation__round__U6456  ( .A(SYNOPSYS_UNCONNECTED_539), .B(
        _f_permutation__round__n2008 ), .Z(_f_permutation__round__c[549] ) );
  XOR2_X2 _f_permutation__round__U6455  ( .A(SYNOPSYS_UNCONNECTED_410), .B(
        _f_permutation__round__n2007 ), .Z(_f_permutation__round__c[1446] ) );
  XOR2_X2 _f_permutation__round__U6454  ( .A(SYNOPSYS_UNCONNECTED_219), .B(
        _f_permutation__round__n2008 ), .Z(_f_permutation__round__c[485] ) );
  XOR2_X2 _f_permutation__round__U6453  ( .A(SYNOPSYS_UNCONNECTED_90), .B(
        _f_permutation__round__n2007 ), .Z(_f_permutation__round__c[1382] ) );
  XOR2_X2 _f_permutation__round__U6452  ( .A(_f_permutation__round_in[1189]), 
        .B(_f_permutation__round__n2008 ), .Z(_f_permutation__round__c[421] )
         );
  XOR2_X2 _f_permutation__round__U6451  ( .A(_f_permutation__round_in[1318]), 
        .B(_f_permutation__round__n2007 ), .Z(_f_permutation__round__c[1318] )
         );
  XOR2_X2 _f_permutation__round__U6450  ( .A(_f_permutation__round_in[1509]), 
        .B(_f_permutation__round__n2008 ), .Z(_f_permutation__round__c[357] )
         );
  XOR2_X2 _f_permutation__round__U6449  ( .A(_f_permutation__round__n1367 ), 
        .B(_f_permutation__round__n1366 ), .Z(_f_permutation__round__n2233 )
         );
  XOR2_X2 _f_permutation__round__U6448  ( .A(SYNOPSYS_UNCONNECTED_861), .B(
        _f_permutation__round__n1368 ), .Z(_f_permutation__round__n1366 ) );
  XOR2_X2 _f_permutation__round__U6447  ( .A(SYNOPSYS_UNCONNECTED_221), .B(
        SYNOPSYS_UNCONNECTED_541), .Z(_f_permutation__round__n1367 ) );
  XOR2_X2 _f_permutation__round__U6446  ( .A(_f_permutation__round_in[1507]), 
        .B(_f_permutation__round_in[1187]), .Z(_f_permutation__round__n1368 )
         );
  XOR2_X2 _f_permutation__round__U6445  ( .A(_f_permutation__round__n1370 ), 
        .B(_f_permutation__round__n1369 ), .Z(_f_permutation__round__n2454 )
         );
  XOR2_X2 _f_permutation__round__U6444  ( .A(SYNOPSYS_UNCONNECTED_1052), .B(
        _f_permutation__round__n1371 ), .Z(_f_permutation__round__n1369 ) );
  XOR2_X2 _f_permutation__round__U6443  ( .A(SYNOPSYS_UNCONNECTED_412), .B(
        SYNOPSYS_UNCONNECTED_732), .Z(_f_permutation__round__n1370 ) );
  XOR2_X2 _f_permutation__round__U6442  ( .A(_f_permutation__round_in[1316]), 
        .B(SYNOPSYS_UNCONNECTED_92), .Z(_f_permutation__round__n1371 ) );
  XOR2_X2 _f_permutation__round__U6441  ( .A(_f_permutation__round__n2233 ), 
        .B(_f_permutation__round__n2454 ), .Z(_f_permutation__round__n2234 )
         );
  XOR2_X2 _f_permutation__round__U6440  ( .A(_f_permutation__round_in[1572]), 
        .B(_f_permutation__round__n2234 ), .Z(_f_permutation__round__c[36] )
         );
  XOR2_X2 _f_permutation__round__U6439  ( .A(_f_permutation__round__n1373 ), 
        .B(_f_permutation__round__n1372 ), .Z(_f_permutation__round__n2009 )
         );
  XOR2_X2 _f_permutation__round__U6438  ( .A(SYNOPSYS_UNCONNECTED_796), .B(
        _f_permutation__round__n1374 ), .Z(_f_permutation__round__n1372 ) );
  XOR2_X2 _f_permutation__round__U6437  ( .A(SYNOPSYS_UNCONNECTED_156), .B(
        SYNOPSYS_UNCONNECTED_476), .Z(_f_permutation__round__n1373 ) );
  XOR2_X2 _f_permutation__round__U6436  ( .A(_f_permutation__round_in[1572]), 
        .B(_f_permutation__round_in[1252]), .Z(_f_permutation__round__n1374 )
         );
  XOR2_X2 _f_permutation__round__U6435  ( .A(_f_permutation__round__n1376 ), 
        .B(_f_permutation__round__n1375 ), .Z(_f_permutation__round__n2220 )
         );
  XOR2_X2 _f_permutation__round__U6434  ( .A(SYNOPSYS_UNCONNECTED_987), .B(
        _f_permutation__round__n1377 ), .Z(_f_permutation__round__n1375 ) );
  XOR2_X2 _f_permutation__round__U6433  ( .A(SYNOPSYS_UNCONNECTED_347), .B(
        SYNOPSYS_UNCONNECTED_667), .Z(_f_permutation__round__n1376 ) );
  XOR2_X2 _f_permutation__round__U6432  ( .A(_f_permutation__round_in[1381]), 
        .B(_f_permutation__round_in[1061]), .Z(_f_permutation__round__n1377 )
         );
  XOR2_X2 _f_permutation__round__U6431  ( .A(_f_permutation__round__n2009 ), 
        .B(_f_permutation__round__n2220 ), .Z(_f_permutation__round__n2010 )
         );
  XOR2_X2 _f_permutation__round__U6430  ( .A(SYNOPSYS_UNCONNECTED_1051), .B(
        _f_permutation__round__n2010 ), .Z(_f_permutation__round__c[1573] ) );
  XOR2_X2 _f_permutation__round__U6429  ( .A(_f_permutation__round__n1379 ), 
        .B(_f_permutation__round__n1378 ), .Z(_f_permutation__round__n2461 )
         );
  XOR2_X2 _f_permutation__round__U6428  ( .A(SYNOPSYS_UNCONNECTED_925), .B(
        _f_permutation__round__n1380 ), .Z(_f_permutation__round__n1378 ) );
  XOR2_X2 _f_permutation__round__U6427  ( .A(SYNOPSYS_UNCONNECTED_285), .B(
        SYNOPSYS_UNCONNECTED_605), .Z(_f_permutation__round__n1379 ) );
  XOR2_X2 _f_permutation__round__U6426  ( .A(_f_permutation__round_in[1443]), 
        .B(_f_permutation__round_in[1123]), .Z(_f_permutation__round__n1380 )
         );
  XOR2_X2 _f_permutation__round__U6425  ( .A(_f_permutation__round__n2009 ), 
        .B(_f_permutation__round__n2461 ), .Z(_f_permutation__round__n2011 )
         );
  XOR2_X2 _f_permutation__round__U6424  ( .A(SYNOPSYS_UNCONNECTED_860), .B(
        _f_permutation__round__n2011 ), .Z(_f_permutation__round__c[612] ) );
  XOR2_X2 _f_permutation__round__U6423  ( .A(SYNOPSYS_UNCONNECTED_731), .B(
        _f_permutation__round__n2010 ), .Z(_f_permutation__round__c[1509] ) );
  XOR2_X2 _f_permutation__round__U6422  ( .A(SYNOPSYS_UNCONNECTED_540), .B(
        _f_permutation__round__n2011 ), .Z(_f_permutation__round__c[548] ) );
  XOR2_X2 _f_permutation__round__U6421  ( .A(SYNOPSYS_UNCONNECTED_411), .B(
        _f_permutation__round__n2010 ), .Z(_f_permutation__round__c[1445] ) );
  XOR2_X2 _f_permutation__round__U6420  ( .A(SYNOPSYS_UNCONNECTED_220), .B(
        _f_permutation__round__n2011 ), .Z(_f_permutation__round__c[484] ) );
  XOR2_X2 _f_permutation__round__U6419  ( .A(SYNOPSYS_UNCONNECTED_91), .B(
        _f_permutation__round__n2010 ), .Z(_f_permutation__round__c[1381] ) );
  XOR2_X2 _f_permutation__round__U6418  ( .A(_f_permutation__round_in[1188]), 
        .B(_f_permutation__round__n2011 ), .Z(_f_permutation__round__c[420] )
         );
  XOR2_X2 _f_permutation__round__U6417  ( .A(_f_permutation__round_in[1317]), 
        .B(_f_permutation__round__n2010 ), .Z(_f_permutation__round__c[1317] )
         );
  XOR2_X2 _f_permutation__round__U6416  ( .A(_f_permutation__round_in[1508]), 
        .B(_f_permutation__round__n2011 ), .Z(_f_permutation__round__c[356] )
         );
  XOR2_X2 _f_permutation__round__U6415  ( .A(_f_permutation__round__n1382 ), 
        .B(_f_permutation__round__n1381 ), .Z(_f_permutation__round__n2237 )
         );
  XOR2_X2 _f_permutation__round__U6414  ( .A(SYNOPSYS_UNCONNECTED_862), .B(
        _f_permutation__round__n1383 ), .Z(_f_permutation__round__n1381 ) );
  XOR2_X2 _f_permutation__round__U6413  ( .A(SYNOPSYS_UNCONNECTED_222), .B(
        SYNOPSYS_UNCONNECTED_542), .Z(_f_permutation__round__n1382 ) );
  XOR2_X2 _f_permutation__round__U6412  ( .A(_f_permutation__round_in[1506]), 
        .B(_f_permutation__round_in[1186]), .Z(_f_permutation__round__n1383 )
         );
  XOR2_X2 _f_permutation__round__U6411  ( .A(_f_permutation__round__n1385 ), 
        .B(_f_permutation__round__n1384 ), .Z(_f_permutation__round__n2457 )
         );
  XOR2_X2 _f_permutation__round__U6410  ( .A(SYNOPSYS_UNCONNECTED_1053), .B(
        _f_permutation__round__n1386 ), .Z(_f_permutation__round__n1384 ) );
  XOR2_X2 _f_permutation__round__U6409  ( .A(SYNOPSYS_UNCONNECTED_413), .B(
        SYNOPSYS_UNCONNECTED_733), .Z(_f_permutation__round__n1385 ) );
  XOR2_X2 _f_permutation__round__U6408  ( .A(_f_permutation__round_in[1315]), 
        .B(SYNOPSYS_UNCONNECTED_93), .Z(_f_permutation__round__n1386 ) );
  XOR2_X2 _f_permutation__round__U6407  ( .A(_f_permutation__round__n2237 ), 
        .B(_f_permutation__round__n2457 ), .Z(_f_permutation__round__n2238 )
         );
  XOR2_X2 _f_permutation__round__U6406  ( .A(_f_permutation__round_in[1571]), 
        .B(_f_permutation__round__n2238 ), .Z(_f_permutation__round__c[35] )
         );
  XOR2_X2 _f_permutation__round__U6405  ( .A(_f_permutation__round__n1388 ), 
        .B(_f_permutation__round__n1387 ), .Z(_f_permutation__round__n2012 )
         );
  XOR2_X2 _f_permutation__round__U6404  ( .A(SYNOPSYS_UNCONNECTED_797), .B(
        _f_permutation__round__n1389 ), .Z(_f_permutation__round__n1387 ) );
  XOR2_X2 _f_permutation__round__U6403  ( .A(SYNOPSYS_UNCONNECTED_157), .B(
        SYNOPSYS_UNCONNECTED_477), .Z(_f_permutation__round__n1388 ) );
  XOR2_X2 _f_permutation__round__U6402  ( .A(_f_permutation__round_in[1571]), 
        .B(_f_permutation__round_in[1251]), .Z(_f_permutation__round__n1389 )
         );
  XOR2_X2 _f_permutation__round__U6401  ( .A(_f_permutation__round__n1391 ), 
        .B(_f_permutation__round__n1390 ), .Z(_f_permutation__round__n2224 )
         );
  XOR2_X2 _f_permutation__round__U6400  ( .A(SYNOPSYS_UNCONNECTED_988), .B(
        _f_permutation__round__n1392 ), .Z(_f_permutation__round__n1390 ) );
  XOR2_X2 _f_permutation__round__U6399  ( .A(SYNOPSYS_UNCONNECTED_348), .B(
        SYNOPSYS_UNCONNECTED_668), .Z(_f_permutation__round__n1391 ) );
  XOR2_X2 _f_permutation__round__U6398  ( .A(_f_permutation__round_in[1380]), 
        .B(_f_permutation__round_in[1060]), .Z(_f_permutation__round__n1392 )
         );
  XOR2_X2 _f_permutation__round__U6397  ( .A(_f_permutation__round__n2012 ), 
        .B(_f_permutation__round__n2224 ), .Z(_f_permutation__round__n2013 )
         );
  XOR2_X2 _f_permutation__round__U6396  ( .A(SYNOPSYS_UNCONNECTED_1052), .B(
        _f_permutation__round__n2013 ), .Z(_f_permutation__round__c[1572] ) );
  XOR2_X2 _f_permutation__round__U6395  ( .A(_f_permutation__round__n1394 ), 
        .B(_f_permutation__round__n1393 ), .Z(_f_permutation__round__n2464 )
         );
  XOR2_X2 _f_permutation__round__U6394  ( .A(SYNOPSYS_UNCONNECTED_926), .B(
        _f_permutation__round__n1395 ), .Z(_f_permutation__round__n1393 ) );
  XOR2_X2 _f_permutation__round__U6393  ( .A(SYNOPSYS_UNCONNECTED_286), .B(
        SYNOPSYS_UNCONNECTED_606), .Z(_f_permutation__round__n1394 ) );
  XOR2_X2 _f_permutation__round__U6392  ( .A(_f_permutation__round_in[1442]), 
        .B(_f_permutation__round_in[1122]), .Z(_f_permutation__round__n1395 )
         );
  XOR2_X2 _f_permutation__round__U6391  ( .A(_f_permutation__round__n2012 ), 
        .B(_f_permutation__round__n2464 ), .Z(_f_permutation__round__n2014 )
         );
  XOR2_X2 _f_permutation__round__U6390  ( .A(SYNOPSYS_UNCONNECTED_861), .B(
        _f_permutation__round__n2014 ), .Z(_f_permutation__round__c[611] ) );
  XOR2_X2 _f_permutation__round__U6389  ( .A(SYNOPSYS_UNCONNECTED_732), .B(
        _f_permutation__round__n2013 ), .Z(_f_permutation__round__c[1508] ) );
  XOR2_X2 _f_permutation__round__U6388  ( .A(SYNOPSYS_UNCONNECTED_541), .B(
        _f_permutation__round__n2014 ), .Z(_f_permutation__round__c[547] ) );
  XOR2_X2 _f_permutation__round__U6387  ( .A(SYNOPSYS_UNCONNECTED_412), .B(
        _f_permutation__round__n2013 ), .Z(_f_permutation__round__c[1444] ) );
  XOR2_X2 _f_permutation__round__U6386  ( .A(SYNOPSYS_UNCONNECTED_221), .B(
        _f_permutation__round__n2014 ), .Z(_f_permutation__round__c[483] ) );
  XOR2_X2 _f_permutation__round__U6385  ( .A(SYNOPSYS_UNCONNECTED_92), .B(
        _f_permutation__round__n2013 ), .Z(_f_permutation__round__c[1380] ) );
  XOR2_X2 _f_permutation__round__U6384  ( .A(_f_permutation__round_in[1187]), 
        .B(_f_permutation__round__n2014 ), .Z(_f_permutation__round__c[419] )
         );
  XOR2_X2 _f_permutation__round__U6383  ( .A(_f_permutation__round_in[1316]), 
        .B(_f_permutation__round__n2013 ), .Z(_f_permutation__round__c[1316] )
         );
  XOR2_X2 _f_permutation__round__U6382  ( .A(_f_permutation__round_in[1507]), 
        .B(_f_permutation__round__n2014 ), .Z(_f_permutation__round__c[355] )
         );
  XOR2_X2 _f_permutation__round__U6381  ( .A(_f_permutation__round__n1397 ), 
        .B(_f_permutation__round__n1396 ), .Z(_f_permutation__round__n2241 )
         );
  XOR2_X2 _f_permutation__round__U6380  ( .A(SYNOPSYS_UNCONNECTED_863), .B(
        _f_permutation__round__n1398 ), .Z(_f_permutation__round__n1396 ) );
  XOR2_X2 _f_permutation__round__U6379  ( .A(SYNOPSYS_UNCONNECTED_223), .B(
        SYNOPSYS_UNCONNECTED_543), .Z(_f_permutation__round__n1397 ) );
  XOR2_X2 _f_permutation__round__U6378  ( .A(_f_permutation__round_in[1505]), 
        .B(_f_permutation__round_in[1185]), .Z(_f_permutation__round__n1398 )
         );
  XOR2_X2 _f_permutation__round__U6377  ( .A(_f_permutation__round__n1400 ), 
        .B(_f_permutation__round__n1399 ), .Z(_f_permutation__round__n2460 )
         );
  XOR2_X2 _f_permutation__round__U6376  ( .A(SYNOPSYS_UNCONNECTED_1054), .B(
        _f_permutation__round__n1401 ), .Z(_f_permutation__round__n1399 ) );
  XOR2_X2 _f_permutation__round__U6375  ( .A(SYNOPSYS_UNCONNECTED_414), .B(
        SYNOPSYS_UNCONNECTED_734), .Z(_f_permutation__round__n1400 ) );
  XOR2_X2 _f_permutation__round__U6374  ( .A(_f_permutation__round_in[1314]), 
        .B(SYNOPSYS_UNCONNECTED_94), .Z(_f_permutation__round__n1401 ) );
  XOR2_X2 _f_permutation__round__U6373  ( .A(_f_permutation__round__n2241 ), 
        .B(_f_permutation__round__n2460 ), .Z(_f_permutation__round__n2242 )
         );
  XOR2_X2 _f_permutation__round__U6372  ( .A(_f_permutation__round_in[1570]), 
        .B(_f_permutation__round__n2242 ), .Z(_f_permutation__round__c[34] )
         );
  XOR2_X2 _f_permutation__round__U6371  ( .A(_f_permutation__round__n1403 ), 
        .B(_f_permutation__round__n1402 ), .Z(_f_permutation__round__n2015 )
         );
  XOR2_X2 _f_permutation__round__U6370  ( .A(SYNOPSYS_UNCONNECTED_798), .B(
        _f_permutation__round__n1404 ), .Z(_f_permutation__round__n1402 ) );
  XOR2_X2 _f_permutation__round__U6369  ( .A(SYNOPSYS_UNCONNECTED_158), .B(
        SYNOPSYS_UNCONNECTED_478), .Z(_f_permutation__round__n1403 ) );
  XOR2_X2 _f_permutation__round__U6368  ( .A(_f_permutation__round_in[1570]), 
        .B(_f_permutation__round_in[1250]), .Z(_f_permutation__round__n1404 )
         );
  XOR2_X2 _f_permutation__round__U6367  ( .A(_f_permutation__round__n1406 ), 
        .B(_f_permutation__round__n1405 ), .Z(_f_permutation__round__n2228 )
         );
  XOR2_X2 _f_permutation__round__U6366  ( .A(SYNOPSYS_UNCONNECTED_989), .B(
        _f_permutation__round__n1407 ), .Z(_f_permutation__round__n1405 ) );
  XOR2_X2 _f_permutation__round__U6365  ( .A(SYNOPSYS_UNCONNECTED_349), .B(
        SYNOPSYS_UNCONNECTED_669), .Z(_f_permutation__round__n1406 ) );
  XOR2_X2 _f_permutation__round__U6364  ( .A(_f_permutation__round_in[1379]), 
        .B(_f_permutation__round_in[1059]), .Z(_f_permutation__round__n1407 )
         );
  XOR2_X2 _f_permutation__round__U6363  ( .A(_f_permutation__round__n2015 ), 
        .B(_f_permutation__round__n2228 ), .Z(_f_permutation__round__n2016 )
         );
  XOR2_X2 _f_permutation__round__U6362  ( .A(SYNOPSYS_UNCONNECTED_1053), .B(
        _f_permutation__round__n2016 ), .Z(_f_permutation__round__c[1571] ) );
  XOR2_X2 _f_permutation__round__U6361  ( .A(_f_permutation__round__n1409 ), 
        .B(_f_permutation__round__n1408 ), .Z(_f_permutation__round__n2467 )
         );
  XOR2_X2 _f_permutation__round__U6360  ( .A(SYNOPSYS_UNCONNECTED_927), .B(
        _f_permutation__round__n1410 ), .Z(_f_permutation__round__n1408 ) );
  XOR2_X2 _f_permutation__round__U6359  ( .A(SYNOPSYS_UNCONNECTED_287), .B(
        SYNOPSYS_UNCONNECTED_607), .Z(_f_permutation__round__n1409 ) );
  XOR2_X2 _f_permutation__round__U6358  ( .A(_f_permutation__round_in[1441]), 
        .B(_f_permutation__round_in[1121]), .Z(_f_permutation__round__n1410 )
         );
  XOR2_X2 _f_permutation__round__U6357  ( .A(_f_permutation__round__n2015 ), 
        .B(_f_permutation__round__n2467 ), .Z(_f_permutation__round__n2017 )
         );
  XOR2_X2 _f_permutation__round__U6356  ( .A(SYNOPSYS_UNCONNECTED_862), .B(
        _f_permutation__round__n2017 ), .Z(_f_permutation__round__c[610] ) );
  XOR2_X2 _f_permutation__round__U6355  ( .A(SYNOPSYS_UNCONNECTED_733), .B(
        _f_permutation__round__n2016 ), .Z(_f_permutation__round__c[1507] ) );
  XOR2_X2 _f_permutation__round__U6354  ( .A(SYNOPSYS_UNCONNECTED_542), .B(
        _f_permutation__round__n2017 ), .Z(_f_permutation__round__c[546] ) );
  XOR2_X2 _f_permutation__round__U6353  ( .A(SYNOPSYS_UNCONNECTED_413), .B(
        _f_permutation__round__n2016 ), .Z(_f_permutation__round__c[1443] ) );
  XOR2_X2 _f_permutation__round__U6352  ( .A(SYNOPSYS_UNCONNECTED_222), .B(
        _f_permutation__round__n2017 ), .Z(_f_permutation__round__c[482] ) );
  XOR2_X2 _f_permutation__round__U6351  ( .A(SYNOPSYS_UNCONNECTED_93), .B(
        _f_permutation__round__n2016 ), .Z(_f_permutation__round__c[1379] ) );
  XOR2_X2 _f_permutation__round__U6350  ( .A(_f_permutation__round_in[1186]), 
        .B(_f_permutation__round__n2017 ), .Z(_f_permutation__round__c[418] )
         );
  XOR2_X2 _f_permutation__round__U6349  ( .A(_f_permutation__round_in[1315]), 
        .B(_f_permutation__round__n2016 ), .Z(_f_permutation__round__c[1315] )
         );
  XOR2_X2 _f_permutation__round__U6348  ( .A(_f_permutation__round_in[1506]), 
        .B(_f_permutation__round__n2017 ), .Z(_f_permutation__round__c[354] )
         );
  XOR2_X2 _f_permutation__round__U6347  ( .A(_f_permutation__round__n1412 ), 
        .B(_f_permutation__round__n1411 ), .Z(_f_permutation__round__n2245 )
         );
  XOR2_X2 _f_permutation__round__U6346  ( .A(SYNOPSYS_UNCONNECTED_864), .B(
        _f_permutation__round__n1413 ), .Z(_f_permutation__round__n1411 ) );
  XOR2_X2 _f_permutation__round__U6345  ( .A(SYNOPSYS_UNCONNECTED_224), .B(
        SYNOPSYS_UNCONNECTED_544), .Z(_f_permutation__round__n1412 ) );
  XOR2_X2 _f_permutation__round__U6344  ( .A(_f_permutation__round_in[1504]), 
        .B(_f_permutation__round_in[1184]), .Z(_f_permutation__round__n1413 )
         );
  XOR2_X2 _f_permutation__round__U6343  ( .A(_f_permutation__round__n1415 ), 
        .B(_f_permutation__round__n1414 ), .Z(_f_permutation__round__n2463 )
         );
  XOR2_X2 _f_permutation__round__U6342  ( .A(SYNOPSYS_UNCONNECTED_1055), .B(
        _f_permutation__round__n1416 ), .Z(_f_permutation__round__n1414 ) );
  XOR2_X2 _f_permutation__round__U6341  ( .A(SYNOPSYS_UNCONNECTED_415), .B(
        SYNOPSYS_UNCONNECTED_735), .Z(_f_permutation__round__n1415 ) );
  XOR2_X2 _f_permutation__round__U6340  ( .A(_f_permutation__round_in[1313]), 
        .B(SYNOPSYS_UNCONNECTED_95), .Z(_f_permutation__round__n1416 ) );
  XOR2_X2 _f_permutation__round__U6339  ( .A(_f_permutation__round__n2245 ), 
        .B(_f_permutation__round__n2463 ), .Z(_f_permutation__round__n2246 )
         );
  XOR2_X2 _f_permutation__round__U6338  ( .A(_f_permutation__round_in[1569]), 
        .B(_f_permutation__round__n2246 ), .Z(_f_permutation__round__c[33] )
         );
  XOR2_X2 _f_permutation__round__U6337  ( .A(_f_permutation__round__n1418 ), 
        .B(_f_permutation__round__n1417 ), .Z(_f_permutation__round__n2018 )
         );
  XOR2_X2 _f_permutation__round__U6336  ( .A(SYNOPSYS_UNCONNECTED_799), .B(
        _f_permutation__round__n1419 ), .Z(_f_permutation__round__n1417 ) );
  XOR2_X2 _f_permutation__round__U6335  ( .A(SYNOPSYS_UNCONNECTED_159), .B(
        SYNOPSYS_UNCONNECTED_479), .Z(_f_permutation__round__n1418 ) );
  XOR2_X2 _f_permutation__round__U6334  ( .A(_f_permutation__round_in[1569]), 
        .B(_f_permutation__round_in[1249]), .Z(_f_permutation__round__n1419 )
         );
  XOR2_X2 _f_permutation__round__U6333  ( .A(_f_permutation__round__n1421 ), 
        .B(_f_permutation__round__n1420 ), .Z(_f_permutation__round__n2232 )
         );
  XOR2_X2 _f_permutation__round__U6332  ( .A(SYNOPSYS_UNCONNECTED_990), .B(
        _f_permutation__round__n1422 ), .Z(_f_permutation__round__n1420 ) );
  XOR2_X2 _f_permutation__round__U6331  ( .A(SYNOPSYS_UNCONNECTED_350), .B(
        SYNOPSYS_UNCONNECTED_670), .Z(_f_permutation__round__n1421 ) );
  XOR2_X2 _f_permutation__round__U6330  ( .A(_f_permutation__round_in[1378]), 
        .B(_f_permutation__round_in[1058]), .Z(_f_permutation__round__n1422 )
         );
  XOR2_X2 _f_permutation__round__U6329  ( .A(_f_permutation__round__n2018 ), 
        .B(_f_permutation__round__n2232 ), .Z(_f_permutation__round__n2019 )
         );
  XOR2_X2 _f_permutation__round__U6328  ( .A(SYNOPSYS_UNCONNECTED_1054), .B(
        _f_permutation__round__n2019 ), .Z(_f_permutation__round__c[1570] ) );
  XOR2_X2 _f_permutation__round__U6327  ( .A(_f_permutation__round__n1424 ), 
        .B(_f_permutation__round__n1423 ), .Z(_f_permutation__round__n2470 )
         );
  XOR2_X2 _f_permutation__round__U6326  ( .A(SYNOPSYS_UNCONNECTED_928), .B(
        _f_permutation__round__n1425 ), .Z(_f_permutation__round__n1423 ) );
  XOR2_X2 _f_permutation__round__U6325  ( .A(SYNOPSYS_UNCONNECTED_288), .B(
        SYNOPSYS_UNCONNECTED_608), .Z(_f_permutation__round__n1424 ) );
  XOR2_X2 _f_permutation__round__U6324  ( .A(_f_permutation__round_in[1440]), 
        .B(_f_permutation__round_in[1120]), .Z(_f_permutation__round__n1425 )
         );
  XOR2_X2 _f_permutation__round__U6323  ( .A(_f_permutation__round__n2018 ), 
        .B(_f_permutation__round__n2470 ), .Z(_f_permutation__round__n2020 )
         );
  XOR2_X2 _f_permutation__round__U6322  ( .A(SYNOPSYS_UNCONNECTED_863), .B(
        _f_permutation__round__n2020 ), .Z(_f_permutation__round__c[609] ) );
  XOR2_X2 _f_permutation__round__U6321  ( .A(SYNOPSYS_UNCONNECTED_734), .B(
        _f_permutation__round__n2019 ), .Z(_f_permutation__round__c[1506] ) );
  XOR2_X2 _f_permutation__round__U6320  ( .A(SYNOPSYS_UNCONNECTED_543), .B(
        _f_permutation__round__n2020 ), .Z(_f_permutation__round__c[545] ) );
  XOR2_X2 _f_permutation__round__U6319  ( .A(SYNOPSYS_UNCONNECTED_414), .B(
        _f_permutation__round__n2019 ), .Z(_f_permutation__round__c[1442] ) );
  XOR2_X2 _f_permutation__round__U6318  ( .A(SYNOPSYS_UNCONNECTED_223), .B(
        _f_permutation__round__n2020 ), .Z(_f_permutation__round__c[481] ) );
  XOR2_X2 _f_permutation__round__U6317  ( .A(SYNOPSYS_UNCONNECTED_94), .B(
        _f_permutation__round__n2019 ), .Z(_f_permutation__round__c[1378] ) );
  XOR2_X2 _f_permutation__round__U6316  ( .A(_f_permutation__round_in[1185]), 
        .B(_f_permutation__round__n2020 ), .Z(_f_permutation__round__c[417] )
         );
  XOR2_X2 _f_permutation__round__U6315  ( .A(_f_permutation__round_in[1314]), 
        .B(_f_permutation__round__n2019 ), .Z(_f_permutation__round__c[1314] )
         );
  XOR2_X2 _f_permutation__round__U6314  ( .A(_f_permutation__round_in[1505]), 
        .B(_f_permutation__round__n2020 ), .Z(_f_permutation__round__c[353] )
         );
  XOR2_X2 _f_permutation__round__U6313  ( .A(_f_permutation__round__n1427 ), 
        .B(_f_permutation__round__n1426 ), .Z(_f_permutation__round__n2249 )
         );
  XOR2_X2 _f_permutation__round__U6312  ( .A(SYNOPSYS_UNCONNECTED_865), .B(
        _f_permutation__round__n1428 ), .Z(_f_permutation__round__n1426 ) );
  XOR2_X2 _f_permutation__round__U6311  ( .A(SYNOPSYS_UNCONNECTED_225), .B(
        SYNOPSYS_UNCONNECTED_545), .Z(_f_permutation__round__n1427 ) );
  XOR2_X2 _f_permutation__round__U6310  ( .A(_f_permutation__round_in[1503]), 
        .B(_f_permutation__round_in[1183]), .Z(_f_permutation__round__n1428 )
         );
  XOR2_X2 _f_permutation__round__U6309  ( .A(_f_permutation__round__n1430 ), 
        .B(_f_permutation__round__n1429 ), .Z(_f_permutation__round__n2466 )
         );
  XOR2_X2 _f_permutation__round__U6308  ( .A(SYNOPSYS_UNCONNECTED_1056), .B(
        _f_permutation__round__n1431 ), .Z(_f_permutation__round__n1429 ) );
  XOR2_X2 _f_permutation__round__U6307  ( .A(SYNOPSYS_UNCONNECTED_416), .B(
        SYNOPSYS_UNCONNECTED_736), .Z(_f_permutation__round__n1430 ) );
  XOR2_X2 _f_permutation__round__U6306  ( .A(_f_permutation__round_in[1312]), 
        .B(SYNOPSYS_UNCONNECTED_96), .Z(_f_permutation__round__n1431 ) );
  XOR2_X2 _f_permutation__round__U6305  ( .A(_f_permutation__round__n2249 ), 
        .B(_f_permutation__round__n2466 ), .Z(_f_permutation__round__n2250 )
         );
  XOR2_X2 _f_permutation__round__U6304  ( .A(_f_permutation__round_in[1568]), 
        .B(_f_permutation__round__n2250 ), .Z(_f_permutation__round__c[32] )
         );
  XOR2_X2 _f_permutation__round__U6303  ( .A(_f_permutation__round__n1433 ), 
        .B(_f_permutation__round__n1432 ), .Z(_f_permutation__round__n2021 )
         );
  XOR2_X2 _f_permutation__round__U6302  ( .A(SYNOPSYS_UNCONNECTED_800), .B(
        _f_permutation__round__n1434 ), .Z(_f_permutation__round__n1432 ) );
  XOR2_X2 _f_permutation__round__U6301  ( .A(SYNOPSYS_UNCONNECTED_160), .B(
        SYNOPSYS_UNCONNECTED_480), .Z(_f_permutation__round__n1433 ) );
  XOR2_X2 _f_permutation__round__U6300  ( .A(_f_permutation__round_in[1568]), 
        .B(_f_permutation__round_in[1248]), .Z(_f_permutation__round__n1434 )
         );
  XOR2_X2 _f_permutation__round__U6299  ( .A(_f_permutation__round__n1436 ), 
        .B(_f_permutation__round__n1435 ), .Z(_f_permutation__round__n2236 )
         );
  XOR2_X2 _f_permutation__round__U6298  ( .A(SYNOPSYS_UNCONNECTED_991), .B(
        _f_permutation__round__n1437 ), .Z(_f_permutation__round__n1435 ) );
  XOR2_X2 _f_permutation__round__U6297  ( .A(SYNOPSYS_UNCONNECTED_351), .B(
        SYNOPSYS_UNCONNECTED_671), .Z(_f_permutation__round__n1436 ) );
  XOR2_X2 _f_permutation__round__U6296  ( .A(_f_permutation__round_in[1377]), 
        .B(_f_permutation__round_in[1057]), .Z(_f_permutation__round__n1437 )
         );
  XOR2_X2 _f_permutation__round__U6295  ( .A(_f_permutation__round__n2021 ), 
        .B(_f_permutation__round__n2236 ), .Z(_f_permutation__round__n2022 )
         );
  XOR2_X2 _f_permutation__round__U6294  ( .A(SYNOPSYS_UNCONNECTED_1055), .B(
        _f_permutation__round__n2022 ), .Z(_f_permutation__round__c[1569] ) );
  XOR2_X2 _f_permutation__round__U6293  ( .A(_f_permutation__round__n1439 ), 
        .B(_f_permutation__round__n1438 ), .Z(_f_permutation__round__n2473 )
         );
  XOR2_X2 _f_permutation__round__U6292  ( .A(SYNOPSYS_UNCONNECTED_929), .B(
        _f_permutation__round__n1440 ), .Z(_f_permutation__round__n1438 ) );
  XOR2_X2 _f_permutation__round__U6291  ( .A(SYNOPSYS_UNCONNECTED_289), .B(
        SYNOPSYS_UNCONNECTED_609), .Z(_f_permutation__round__n1439 ) );
  XOR2_X2 _f_permutation__round__U6290  ( .A(_f_permutation__round_in[1439]), 
        .B(_f_permutation__round_in[1119]), .Z(_f_permutation__round__n1440 )
         );
  XOR2_X2 _f_permutation__round__U6289  ( .A(_f_permutation__round__n2021 ), 
        .B(_f_permutation__round__n2473 ), .Z(_f_permutation__round__n2023 )
         );
  XOR2_X2 _f_permutation__round__U6288  ( .A(SYNOPSYS_UNCONNECTED_864), .B(
        _f_permutation__round__n2023 ), .Z(_f_permutation__round__c[608] ) );
  XOR2_X2 _f_permutation__round__U6287  ( .A(SYNOPSYS_UNCONNECTED_735), .B(
        _f_permutation__round__n2022 ), .Z(_f_permutation__round__c[1505] ) );
  XOR2_X2 _f_permutation__round__U6286  ( .A(SYNOPSYS_UNCONNECTED_544), .B(
        _f_permutation__round__n2023 ), .Z(_f_permutation__round__c[544] ) );
  XOR2_X2 _f_permutation__round__U6285  ( .A(SYNOPSYS_UNCONNECTED_415), .B(
        _f_permutation__round__n2022 ), .Z(_f_permutation__round__c[1441] ) );
  XOR2_X2 _f_permutation__round__U6284  ( .A(SYNOPSYS_UNCONNECTED_224), .B(
        _f_permutation__round__n2023 ), .Z(_f_permutation__round__c[480] ) );
  XOR2_X2 _f_permutation__round__U6283  ( .A(SYNOPSYS_UNCONNECTED_95), .B(
        _f_permutation__round__n2022 ), .Z(_f_permutation__round__c[1377] ) );
  XOR2_X2 _f_permutation__round__U6282  ( .A(_f_permutation__round_in[1184]), 
        .B(_f_permutation__round__n2023 ), .Z(_f_permutation__round__c[416] )
         );
  XOR2_X2 _f_permutation__round__U6281  ( .A(_f_permutation__round_in[1313]), 
        .B(_f_permutation__round__n2022 ), .Z(_f_permutation__round__c[1313] )
         );
  XOR2_X2 _f_permutation__round__U6280  ( .A(_f_permutation__round_in[1504]), 
        .B(_f_permutation__round__n2023 ), .Z(_f_permutation__round__c[352] )
         );
  XOR2_X2 _f_permutation__round__U6279  ( .A(_f_permutation__round__n1442 ), 
        .B(_f_permutation__round__n1441 ), .Z(_f_permutation__round__n2253 )
         );
  XOR2_X2 _f_permutation__round__U6278  ( .A(SYNOPSYS_UNCONNECTED_866), .B(
        _f_permutation__round__n1443 ), .Z(_f_permutation__round__n1441 ) );
  XOR2_X2 _f_permutation__round__U6277  ( .A(SYNOPSYS_UNCONNECTED_226), .B(
        SYNOPSYS_UNCONNECTED_546), .Z(_f_permutation__round__n1442 ) );
  XOR2_X2 _f_permutation__round__U6276  ( .A(_f_permutation__round_in[1502]), 
        .B(_f_permutation__round_in[1182]), .Z(_f_permutation__round__n1443 )
         );
  XOR2_X2 _f_permutation__round__U6275  ( .A(_f_permutation__round__n1445 ), 
        .B(_f_permutation__round__n1444 ), .Z(_f_permutation__round__n2469 )
         );
  XOR2_X2 _f_permutation__round__U6274  ( .A(SYNOPSYS_UNCONNECTED_1057), .B(
        _f_permutation__round__n1446 ), .Z(_f_permutation__round__n1444 ) );
  XOR2_X2 _f_permutation__round__U6273  ( .A(SYNOPSYS_UNCONNECTED_417), .B(
        SYNOPSYS_UNCONNECTED_737), .Z(_f_permutation__round__n1445 ) );
  XOR2_X2 _f_permutation__round__U6272  ( .A(_f_permutation__round_in[1311]), 
        .B(SYNOPSYS_UNCONNECTED_97), .Z(_f_permutation__round__n1446 ) );
  XOR2_X2 _f_permutation__round__U6271  ( .A(_f_permutation__round__n2253 ), 
        .B(_f_permutation__round__n2469 ), .Z(_f_permutation__round__n2254 )
         );
  XOR2_X2 _f_permutation__round__U6270  ( .A(_f_permutation__round_in[1567]), 
        .B(_f_permutation__round__n2254 ), .Z(_f_permutation__round__c[31] )
         );
  XOR2_X2 _f_permutation__round__U6269  ( .A(_f_permutation__round__n1448 ), 
        .B(_f_permutation__round__n1447 ), .Z(_f_permutation__round__n2024 )
         );
  XOR2_X2 _f_permutation__round__U6268  ( .A(SYNOPSYS_UNCONNECTED_801), .B(
        _f_permutation__round__n1449 ), .Z(_f_permutation__round__n1447 ) );
  XOR2_X2 _f_permutation__round__U6267  ( .A(SYNOPSYS_UNCONNECTED_161), .B(
        SYNOPSYS_UNCONNECTED_481), .Z(_f_permutation__round__n1448 ) );
  XOR2_X2 _f_permutation__round__U6266  ( .A(_f_permutation__round_in[1567]), 
        .B(_f_permutation__round_in[1247]), .Z(_f_permutation__round__n1449 )
         );
  XOR2_X2 _f_permutation__round__U6265  ( .A(_f_permutation__round__n1451 ), 
        .B(_f_permutation__round__n1450 ), .Z(_f_permutation__round__n2240 )
         );
  XOR2_X2 _f_permutation__round__U6264  ( .A(SYNOPSYS_UNCONNECTED_992), .B(
        _f_permutation__round__n1452 ), .Z(_f_permutation__round__n1450 ) );
  XOR2_X2 _f_permutation__round__U6263  ( .A(SYNOPSYS_UNCONNECTED_352), .B(
        SYNOPSYS_UNCONNECTED_672), .Z(_f_permutation__round__n1451 ) );
  XOR2_X2 _f_permutation__round__U6262  ( .A(_f_permutation__round_in[1376]), 
        .B(_f_permutation__round_in[1056]), .Z(_f_permutation__round__n1452 )
         );
  XOR2_X2 _f_permutation__round__U6261  ( .A(_f_permutation__round__n2024 ), 
        .B(_f_permutation__round__n2240 ), .Z(_f_permutation__round__n2025 )
         );
  XOR2_X2 _f_permutation__round__U6260  ( .A(SYNOPSYS_UNCONNECTED_1056), .B(
        _f_permutation__round__n2025 ), .Z(_f_permutation__round__c[1568] ) );
  XOR2_X2 _f_permutation__round__U6259  ( .A(_f_permutation__round__n1454 ), 
        .B(_f_permutation__round__n1453 ), .Z(_f_permutation__round__n2476 )
         );
  XOR2_X2 _f_permutation__round__U6258  ( .A(SYNOPSYS_UNCONNECTED_930), .B(
        _f_permutation__round__n1455 ), .Z(_f_permutation__round__n1453 ) );
  XOR2_X2 _f_permutation__round__U6257  ( .A(SYNOPSYS_UNCONNECTED_290), .B(
        SYNOPSYS_UNCONNECTED_610), .Z(_f_permutation__round__n1454 ) );
  XOR2_X2 _f_permutation__round__U6256  ( .A(_f_permutation__round_in[1438]), 
        .B(_f_permutation__round_in[1118]), .Z(_f_permutation__round__n1455 )
         );
  XOR2_X2 _f_permutation__round__U6255  ( .A(_f_permutation__round__n2024 ), 
        .B(_f_permutation__round__n2476 ), .Z(_f_permutation__round__n2026 )
         );
  XOR2_X2 _f_permutation__round__U6254  ( .A(SYNOPSYS_UNCONNECTED_865), .B(
        _f_permutation__round__n2026 ), .Z(_f_permutation__round__c[607] ) );
  XOR2_X2 _f_permutation__round__U6253  ( .A(SYNOPSYS_UNCONNECTED_736), .B(
        _f_permutation__round__n2025 ), .Z(_f_permutation__round__c[1504] ) );
  XOR2_X2 _f_permutation__round__U6252  ( .A(SYNOPSYS_UNCONNECTED_545), .B(
        _f_permutation__round__n2026 ), .Z(_f_permutation__round__c[543] ) );
  XOR2_X2 _f_permutation__round__U6251  ( .A(SYNOPSYS_UNCONNECTED_416), .B(
        _f_permutation__round__n2025 ), .Z(_f_permutation__round__c[1440] ) );
  XOR2_X2 _f_permutation__round__U6250  ( .A(SYNOPSYS_UNCONNECTED_225), .B(
        _f_permutation__round__n2026 ), .Z(_f_permutation__round__c[479] ) );
  XOR2_X2 _f_permutation__round__U6249  ( .A(SYNOPSYS_UNCONNECTED_96), .B(
        _f_permutation__round__n2025 ), .Z(_f_permutation__round__c[1376] ) );
  XOR2_X2 _f_permutation__round__U6248  ( .A(_f_permutation__round_in[1183]), 
        .B(_f_permutation__round__n2026 ), .Z(_f_permutation__round__c[415] )
         );
  XOR2_X2 _f_permutation__round__U6247  ( .A(_f_permutation__round_in[1312]), 
        .B(_f_permutation__round__n2025 ), .Z(_f_permutation__round__c[1312] )
         );
  XOR2_X2 _f_permutation__round__U6246  ( .A(_f_permutation__round_in[1503]), 
        .B(_f_permutation__round__n2026 ), .Z(_f_permutation__round__c[351] )
         );
  XOR2_X2 _f_permutation__round__U6245  ( .A(_f_permutation__round__n1457 ), 
        .B(_f_permutation__round__n1456 ), .Z(_f_permutation__round__n2257 )
         );
  XOR2_X2 _f_permutation__round__U6244  ( .A(SYNOPSYS_UNCONNECTED_867), .B(
        _f_permutation__round__n1458 ), .Z(_f_permutation__round__n1456 ) );
  XOR2_X2 _f_permutation__round__U6243  ( .A(SYNOPSYS_UNCONNECTED_227), .B(
        SYNOPSYS_UNCONNECTED_547), .Z(_f_permutation__round__n1457 ) );
  XOR2_X2 _f_permutation__round__U6242  ( .A(_f_permutation__round_in[1501]), 
        .B(_f_permutation__round_in[1181]), .Z(_f_permutation__round__n1458 )
         );
  XOR2_X2 _f_permutation__round__U6241  ( .A(_f_permutation__round__n1460 ), 
        .B(_f_permutation__round__n1459 ), .Z(_f_permutation__round__n2472 )
         );
  XOR2_X2 _f_permutation__round__U6240  ( .A(SYNOPSYS_UNCONNECTED_1058), .B(
        _f_permutation__round__n1461 ), .Z(_f_permutation__round__n1459 ) );
  XOR2_X2 _f_permutation__round__U6239  ( .A(SYNOPSYS_UNCONNECTED_418), .B(
        SYNOPSYS_UNCONNECTED_738), .Z(_f_permutation__round__n1460 ) );
  XOR2_X2 _f_permutation__round__U6238  ( .A(_f_permutation__round_in[1310]), 
        .B(SYNOPSYS_UNCONNECTED_98), .Z(_f_permutation__round__n1461 ) );
  XOR2_X2 _f_permutation__round__U6237  ( .A(_f_permutation__round__n2257 ), 
        .B(_f_permutation__round__n2472 ), .Z(_f_permutation__round__n2258 )
         );
  XOR2_X2 _f_permutation__round__U6236  ( .A(_f_permutation__round_in[1566]), 
        .B(_f_permutation__round__n2258 ), .Z(_f_permutation__round__c[30] )
         );
  XOR2_X2 _f_permutation__round__U6235  ( .A(_f_permutation__round__n1463 ), 
        .B(_f_permutation__round__n1462 ), .Z(_f_permutation__round__n2027 )
         );
  XOR2_X2 _f_permutation__round__U6234  ( .A(SYNOPSYS_UNCONNECTED_802), .B(
        _f_permutation__round__n1464 ), .Z(_f_permutation__round__n1462 ) );
  XOR2_X2 _f_permutation__round__U6233  ( .A(SYNOPSYS_UNCONNECTED_162), .B(
        SYNOPSYS_UNCONNECTED_482), .Z(_f_permutation__round__n1463 ) );
  XOR2_X2 _f_permutation__round__U6232  ( .A(_f_permutation__round_in[1566]), 
        .B(_f_permutation__round_in[1246]), .Z(_f_permutation__round__n1464 )
         );
  XOR2_X2 _f_permutation__round__U6231  ( .A(_f_permutation__round__n1466 ), 
        .B(_f_permutation__round__n1465 ), .Z(_f_permutation__round__n2244 )
         );
  XOR2_X2 _f_permutation__round__U6230  ( .A(SYNOPSYS_UNCONNECTED_993), .B(
        _f_permutation__round__n1467 ), .Z(_f_permutation__round__n1465 ) );
  XOR2_X2 _f_permutation__round__U6229  ( .A(SYNOPSYS_UNCONNECTED_353), .B(
        SYNOPSYS_UNCONNECTED_673), .Z(_f_permutation__round__n1466 ) );
  XOR2_X2 _f_permutation__round__U6228  ( .A(_f_permutation__round_in[1375]), 
        .B(_f_permutation__round_in[1055]), .Z(_f_permutation__round__n1467 )
         );
  XOR2_X2 _f_permutation__round__U6227  ( .A(_f_permutation__round__n2027 ), 
        .B(_f_permutation__round__n2244 ), .Z(_f_permutation__round__n2028 )
         );
  XOR2_X2 _f_permutation__round__U6226  ( .A(SYNOPSYS_UNCONNECTED_1057), .B(
        _f_permutation__round__n2028 ), .Z(_f_permutation__round__c[1567] ) );
  XOR2_X2 _f_permutation__round__U6225  ( .A(_f_permutation__round__n1469 ), 
        .B(_f_permutation__round__n1468 ), .Z(_f_permutation__round__n2479 )
         );
  XOR2_X2 _f_permutation__round__U6224  ( .A(SYNOPSYS_UNCONNECTED_931), .B(
        _f_permutation__round__n1470 ), .Z(_f_permutation__round__n1468 ) );
  XOR2_X2 _f_permutation__round__U6223  ( .A(SYNOPSYS_UNCONNECTED_291), .B(
        SYNOPSYS_UNCONNECTED_611), .Z(_f_permutation__round__n1469 ) );
  XOR2_X2 _f_permutation__round__U6222  ( .A(_f_permutation__round_in[1437]), 
        .B(_f_permutation__round_in[1117]), .Z(_f_permutation__round__n1470 )
         );
  XOR2_X2 _f_permutation__round__U6221  ( .A(_f_permutation__round__n2027 ), 
        .B(_f_permutation__round__n2479 ), .Z(_f_permutation__round__n2029 )
         );
  XOR2_X2 _f_permutation__round__U6220  ( .A(SYNOPSYS_UNCONNECTED_866), .B(
        _f_permutation__round__n2029 ), .Z(_f_permutation__round__c[606] ) );
  XOR2_X2 _f_permutation__round__U6219  ( .A(SYNOPSYS_UNCONNECTED_737), .B(
        _f_permutation__round__n2028 ), .Z(_f_permutation__round__c[1503] ) );
  XOR2_X2 _f_permutation__round__U6218  ( .A(SYNOPSYS_UNCONNECTED_546), .B(
        _f_permutation__round__n2029 ), .Z(_f_permutation__round__c[542] ) );
  XOR2_X2 _f_permutation__round__U6217  ( .A(SYNOPSYS_UNCONNECTED_417), .B(
        _f_permutation__round__n2028 ), .Z(_f_permutation__round__c[1439] ) );
  XOR2_X2 _f_permutation__round__U6216  ( .A(SYNOPSYS_UNCONNECTED_226), .B(
        _f_permutation__round__n2029 ), .Z(_f_permutation__round__c[478] ) );
  XOR2_X2 _f_permutation__round__U6215  ( .A(SYNOPSYS_UNCONNECTED_97), .B(
        _f_permutation__round__n2028 ), .Z(_f_permutation__round__c[1375] ) );
  XOR2_X2 _f_permutation__round__U6214  ( .A(_f_permutation__round_in[1182]), 
        .B(_f_permutation__round__n2029 ), .Z(_f_permutation__round__c[414] )
         );
  XOR2_X2 _f_permutation__round__U6213  ( .A(_f_permutation__round_in[1311]), 
        .B(_f_permutation__round__n2028 ), .Z(_f_permutation__round__c[1311] )
         );
  XOR2_X2 _f_permutation__round__U6212  ( .A(_f_permutation__round_in[1502]), 
        .B(_f_permutation__round__n2029 ), .Z(_f_permutation__round__c[350] )
         );
  XOR2_X2 _f_permutation__round__U6211  ( .A(_f_permutation__round__n1472 ), 
        .B(_f_permutation__round__n1471 ), .Z(_f_permutation__round__n2261 )
         );
  XOR2_X2 _f_permutation__round__U6210  ( .A(SYNOPSYS_UNCONNECTED_868), .B(
        _f_permutation__round__n1473 ), .Z(_f_permutation__round__n1471 ) );
  XOR2_X2 _f_permutation__round__U6209  ( .A(SYNOPSYS_UNCONNECTED_228), .B(
        SYNOPSYS_UNCONNECTED_548), .Z(_f_permutation__round__n1472 ) );
  XOR2_X2 _f_permutation__round__U6208  ( .A(_f_permutation__round_in[1500]), 
        .B(_f_permutation__round_in[1180]), .Z(_f_permutation__round__n1473 )
         );
  XOR2_X2 _f_permutation__round__U6207  ( .A(_f_permutation__round__n1475 ), 
        .B(_f_permutation__round__n1474 ), .Z(_f_permutation__round__n2475 )
         );
  XOR2_X2 _f_permutation__round__U6206  ( .A(SYNOPSYS_UNCONNECTED_1059), .B(
        _f_permutation__round__n1476 ), .Z(_f_permutation__round__n1474 ) );
  XOR2_X2 _f_permutation__round__U6205  ( .A(SYNOPSYS_UNCONNECTED_419), .B(
        SYNOPSYS_UNCONNECTED_739), .Z(_f_permutation__round__n1475 ) );
  XOR2_X2 _f_permutation__round__U6204  ( .A(_f_permutation__round_in[1309]), 
        .B(SYNOPSYS_UNCONNECTED_99), .Z(_f_permutation__round__n1476 ) );
  XOR2_X2 _f_permutation__round__U6203  ( .A(_f_permutation__round__n2261 ), 
        .B(_f_permutation__round__n2475 ), .Z(_f_permutation__round__n2262 )
         );
  XOR2_X2 _f_permutation__round__U6202  ( .A(_f_permutation__round_in[1565]), 
        .B(_f_permutation__round__n2262 ), .Z(_f_permutation__round__c[29] )
         );
  XOR2_X2 _f_permutation__round__U6201  ( .A(_f_permutation__round__n1478 ), 
        .B(_f_permutation__round__n1477 ), .Z(_f_permutation__round__n2030 )
         );
  XOR2_X2 _f_permutation__round__U6200  ( .A(SYNOPSYS_UNCONNECTED_803), .B(
        _f_permutation__round__n1479 ), .Z(_f_permutation__round__n1477 ) );
  XOR2_X2 _f_permutation__round__U6199  ( .A(SYNOPSYS_UNCONNECTED_163), .B(
        SYNOPSYS_UNCONNECTED_483), .Z(_f_permutation__round__n1478 ) );
  XOR2_X2 _f_permutation__round__U6198  ( .A(_f_permutation__round_in[1565]), 
        .B(_f_permutation__round_in[1245]), .Z(_f_permutation__round__n1479 )
         );
  XOR2_X2 _f_permutation__round__U6197  ( .A(_f_permutation__round__n1481 ), 
        .B(_f_permutation__round__n1480 ), .Z(_f_permutation__round__n2248 )
         );
  XOR2_X2 _f_permutation__round__U6196  ( .A(SYNOPSYS_UNCONNECTED_994), .B(
        _f_permutation__round__n1482 ), .Z(_f_permutation__round__n1480 ) );
  XOR2_X2 _f_permutation__round__U6195  ( .A(SYNOPSYS_UNCONNECTED_354), .B(
        SYNOPSYS_UNCONNECTED_674), .Z(_f_permutation__round__n1481 ) );
  XOR2_X2 _f_permutation__round__U6194  ( .A(_f_permutation__round_in[1374]), 
        .B(_f_permutation__round_in[1054]), .Z(_f_permutation__round__n1482 )
         );
  XOR2_X2 _f_permutation__round__U6193  ( .A(_f_permutation__round__n2030 ), 
        .B(_f_permutation__round__n2248 ), .Z(_f_permutation__round__n2031 )
         );
  XOR2_X2 _f_permutation__round__U6192  ( .A(SYNOPSYS_UNCONNECTED_1058), .B(
        _f_permutation__round__n2031 ), .Z(_f_permutation__round__c[1566] ) );
  XOR2_X2 _f_permutation__round__U6191  ( .A(_f_permutation__round__n1484 ), 
        .B(_f_permutation__round__n1483 ), .Z(_f_permutation__round__n2482 )
         );
  XOR2_X2 _f_permutation__round__U6190  ( .A(SYNOPSYS_UNCONNECTED_932), .B(
        _f_permutation__round__n1485 ), .Z(_f_permutation__round__n1483 ) );
  XOR2_X2 _f_permutation__round__U6189  ( .A(SYNOPSYS_UNCONNECTED_292), .B(
        SYNOPSYS_UNCONNECTED_612), .Z(_f_permutation__round__n1484 ) );
  XOR2_X2 _f_permutation__round__U6188  ( .A(_f_permutation__round_in[1436]), 
        .B(_f_permutation__round_in[1116]), .Z(_f_permutation__round__n1485 )
         );
  XOR2_X2 _f_permutation__round__U6187  ( .A(_f_permutation__round__n2030 ), 
        .B(_f_permutation__round__n2482 ), .Z(_f_permutation__round__n2032 )
         );
  XOR2_X2 _f_permutation__round__U6186  ( .A(SYNOPSYS_UNCONNECTED_867), .B(
        _f_permutation__round__n2032 ), .Z(_f_permutation__round__c[605] ) );
  XOR2_X2 _f_permutation__round__U6185  ( .A(SYNOPSYS_UNCONNECTED_738), .B(
        _f_permutation__round__n2031 ), .Z(_f_permutation__round__c[1502] ) );
  XOR2_X2 _f_permutation__round__U6184  ( .A(SYNOPSYS_UNCONNECTED_547), .B(
        _f_permutation__round__n2032 ), .Z(_f_permutation__round__c[541] ) );
  XOR2_X2 _f_permutation__round__U6183  ( .A(SYNOPSYS_UNCONNECTED_418), .B(
        _f_permutation__round__n2031 ), .Z(_f_permutation__round__c[1438] ) );
  XOR2_X2 _f_permutation__round__U6182  ( .A(SYNOPSYS_UNCONNECTED_227), .B(
        _f_permutation__round__n2032 ), .Z(_f_permutation__round__c[477] ) );
  XOR2_X2 _f_permutation__round__U6181  ( .A(SYNOPSYS_UNCONNECTED_98), .B(
        _f_permutation__round__n2031 ), .Z(_f_permutation__round__c[1374] ) );
  XOR2_X2 _f_permutation__round__U6180  ( .A(_f_permutation__round_in[1181]), 
        .B(_f_permutation__round__n2032 ), .Z(_f_permutation__round__c[413] )
         );
  XOR2_X2 _f_permutation__round__U6179  ( .A(_f_permutation__round_in[1310]), 
        .B(_f_permutation__round__n2031 ), .Z(_f_permutation__round__c[1310] )
         );
  XOR2_X2 _f_permutation__round__U6178  ( .A(_f_permutation__round_in[1501]), 
        .B(_f_permutation__round__n2032 ), .Z(_f_permutation__round__c[349] )
         );
  XOR2_X2 _f_permutation__round__U6177  ( .A(_f_permutation__round__n1487 ), 
        .B(_f_permutation__round__n1486 ), .Z(_f_permutation__round__n2265 )
         );
  XOR2_X2 _f_permutation__round__U6176  ( .A(SYNOPSYS_UNCONNECTED_869), .B(
        _f_permutation__round__n1488 ), .Z(_f_permutation__round__n1486 ) );
  XOR2_X2 _f_permutation__round__U6175  ( .A(SYNOPSYS_UNCONNECTED_229), .B(
        SYNOPSYS_UNCONNECTED_549), .Z(_f_permutation__round__n1487 ) );
  XOR2_X2 _f_permutation__round__U6174  ( .A(_f_permutation__round_in[1499]), 
        .B(_f_permutation__round_in[1179]), .Z(_f_permutation__round__n1488 )
         );
  XOR2_X2 _f_permutation__round__U6173  ( .A(_f_permutation__round__n1490 ), 
        .B(_f_permutation__round__n1489 ), .Z(_f_permutation__round__n2478 )
         );
  XOR2_X2 _f_permutation__round__U6172  ( .A(SYNOPSYS_UNCONNECTED_1060), .B(
        _f_permutation__round__n1491 ), .Z(_f_permutation__round__n1489 ) );
  XOR2_X2 _f_permutation__round__U6171  ( .A(SYNOPSYS_UNCONNECTED_420), .B(
        SYNOPSYS_UNCONNECTED_740), .Z(_f_permutation__round__n1490 ) );
  XOR2_X2 _f_permutation__round__U6170  ( .A(_f_permutation__round_in[1308]), 
        .B(SYNOPSYS_UNCONNECTED_100), .Z(_f_permutation__round__n1491 ) );
  XOR2_X2 _f_permutation__round__U6169  ( .A(_f_permutation__round__n2265 ), 
        .B(_f_permutation__round__n2478 ), .Z(_f_permutation__round__n2266 )
         );
  XOR2_X2 _f_permutation__round__U6168  ( .A(_f_permutation__round_in[1564]), 
        .B(_f_permutation__round__n2266 ), .Z(_f_permutation__round__c[28] )
         );
  XOR2_X2 _f_permutation__round__U6167  ( .A(_f_permutation__round__n1493 ), 
        .B(_f_permutation__round__n1492 ), .Z(_f_permutation__round__n2033 )
         );
  XOR2_X2 _f_permutation__round__U6166  ( .A(SYNOPSYS_UNCONNECTED_804), .B(
        _f_permutation__round__n1494 ), .Z(_f_permutation__round__n1492 ) );
  XOR2_X2 _f_permutation__round__U6165  ( .A(SYNOPSYS_UNCONNECTED_164), .B(
        SYNOPSYS_UNCONNECTED_484), .Z(_f_permutation__round__n1493 ) );
  XOR2_X2 _f_permutation__round__U6164  ( .A(_f_permutation__round_in[1564]), 
        .B(_f_permutation__round_in[1244]), .Z(_f_permutation__round__n1494 )
         );
  XOR2_X2 _f_permutation__round__U6163  ( .A(_f_permutation__round__n1496 ), 
        .B(_f_permutation__round__n1495 ), .Z(_f_permutation__round__n2252 )
         );
  XOR2_X2 _f_permutation__round__U6162  ( .A(SYNOPSYS_UNCONNECTED_995), .B(
        _f_permutation__round__n1497 ), .Z(_f_permutation__round__n1495 ) );
  XOR2_X2 _f_permutation__round__U6161  ( .A(SYNOPSYS_UNCONNECTED_355), .B(
        SYNOPSYS_UNCONNECTED_675), .Z(_f_permutation__round__n1496 ) );
  XOR2_X2 _f_permutation__round__U6160  ( .A(_f_permutation__round_in[1373]), 
        .B(_f_permutation__round_in[1053]), .Z(_f_permutation__round__n1497 )
         );
  XOR2_X2 _f_permutation__round__U6159  ( .A(_f_permutation__round__n2033 ), 
        .B(_f_permutation__round__n2252 ), .Z(_f_permutation__round__n2034 )
         );
  XOR2_X2 _f_permutation__round__U6158  ( .A(SYNOPSYS_UNCONNECTED_1059), .B(
        _f_permutation__round__n2034 ), .Z(_f_permutation__round__c[1565] ) );
  XOR2_X2 _f_permutation__round__U6157  ( .A(_f_permutation__round__n1499 ), 
        .B(_f_permutation__round__n1498 ), .Z(_f_permutation__round__n2485 )
         );
  XOR2_X2 _f_permutation__round__U6156  ( .A(SYNOPSYS_UNCONNECTED_933), .B(
        _f_permutation__round__n1500 ), .Z(_f_permutation__round__n1498 ) );
  XOR2_X2 _f_permutation__round__U6155  ( .A(SYNOPSYS_UNCONNECTED_293), .B(
        SYNOPSYS_UNCONNECTED_613), .Z(_f_permutation__round__n1499 ) );
  XOR2_X2 _f_permutation__round__U6154  ( .A(_f_permutation__round_in[1435]), 
        .B(_f_permutation__round_in[1115]), .Z(_f_permutation__round__n1500 )
         );
  XOR2_X2 _f_permutation__round__U6153  ( .A(_f_permutation__round__n2033 ), 
        .B(_f_permutation__round__n2485 ), .Z(_f_permutation__round__n2035 )
         );
  XOR2_X2 _f_permutation__round__U6152  ( .A(SYNOPSYS_UNCONNECTED_868), .B(
        _f_permutation__round__n2035 ), .Z(_f_permutation__round__c[604] ) );
  XOR2_X2 _f_permutation__round__U6151  ( .A(SYNOPSYS_UNCONNECTED_739), .B(
        _f_permutation__round__n2034 ), .Z(_f_permutation__round__c[1501] ) );
  XOR2_X2 _f_permutation__round__U6150  ( .A(SYNOPSYS_UNCONNECTED_548), .B(
        _f_permutation__round__n2035 ), .Z(_f_permutation__round__c[540] ) );
  XOR2_X2 _f_permutation__round__U6149  ( .A(SYNOPSYS_UNCONNECTED_419), .B(
        _f_permutation__round__n2034 ), .Z(_f_permutation__round__c[1437] ) );
  XOR2_X2 _f_permutation__round__U6148  ( .A(SYNOPSYS_UNCONNECTED_228), .B(
        _f_permutation__round__n2035 ), .Z(_f_permutation__round__c[476] ) );
  XOR2_X2 _f_permutation__round__U6147  ( .A(SYNOPSYS_UNCONNECTED_99), .B(
        _f_permutation__round__n2034 ), .Z(_f_permutation__round__c[1373] ) );
  XOR2_X2 _f_permutation__round__U6146  ( .A(_f_permutation__round_in[1180]), 
        .B(_f_permutation__round__n2035 ), .Z(_f_permutation__round__c[412] )
         );
  XOR2_X2 _f_permutation__round__U6145  ( .A(_f_permutation__round_in[1309]), 
        .B(_f_permutation__round__n2034 ), .Z(_f_permutation__round__c[1309] )
         );
  XOR2_X2 _f_permutation__round__U6144  ( .A(_f_permutation__round_in[1500]), 
        .B(_f_permutation__round__n2035 ), .Z(_f_permutation__round__c[348] )
         );
  XOR2_X2 _f_permutation__round__U6143  ( .A(_f_permutation__round__n1502 ), 
        .B(_f_permutation__round__n1501 ), .Z(_f_permutation__round__n2269 )
         );
  XOR2_X2 _f_permutation__round__U6142  ( .A(SYNOPSYS_UNCONNECTED_870), .B(
        _f_permutation__round__n1503 ), .Z(_f_permutation__round__n1501 ) );
  XOR2_X2 _f_permutation__round__U6141  ( .A(SYNOPSYS_UNCONNECTED_230), .B(
        SYNOPSYS_UNCONNECTED_550), .Z(_f_permutation__round__n1502 ) );
  XOR2_X2 _f_permutation__round__U6140  ( .A(_f_permutation__round_in[1498]), 
        .B(_f_permutation__round_in[1178]), .Z(_f_permutation__round__n1503 )
         );
  XOR2_X2 _f_permutation__round__U6139  ( .A(_f_permutation__round__n1505 ), 
        .B(_f_permutation__round__n1504 ), .Z(_f_permutation__round__n2481 )
         );
  XOR2_X2 _f_permutation__round__U6138  ( .A(SYNOPSYS_UNCONNECTED_1061), .B(
        _f_permutation__round__n1506 ), .Z(_f_permutation__round__n1504 ) );
  XOR2_X2 _f_permutation__round__U6137  ( .A(SYNOPSYS_UNCONNECTED_421), .B(
        SYNOPSYS_UNCONNECTED_741), .Z(_f_permutation__round__n1505 ) );
  XOR2_X2 _f_permutation__round__U6136  ( .A(_f_permutation__round_in[1307]), 
        .B(SYNOPSYS_UNCONNECTED_101), .Z(_f_permutation__round__n1506 ) );
  XOR2_X2 _f_permutation__round__U6135  ( .A(_f_permutation__round__n2269 ), 
        .B(_f_permutation__round__n2481 ), .Z(_f_permutation__round__n2270 )
         );
  XOR2_X2 _f_permutation__round__U6134  ( .A(_f_permutation__round_in[1563]), 
        .B(_f_permutation__round__n2270 ), .Z(_f_permutation__round__c[27] )
         );
  XOR2_X2 _f_permutation__round__U6133  ( .A(_f_permutation__round__n1508 ), 
        .B(_f_permutation__round__n1507 ), .Z(_f_permutation__round__n2036 )
         );
  XOR2_X2 _f_permutation__round__U6132  ( .A(SYNOPSYS_UNCONNECTED_805), .B(
        _f_permutation__round__n1509 ), .Z(_f_permutation__round__n1507 ) );
  XOR2_X2 _f_permutation__round__U6131  ( .A(SYNOPSYS_UNCONNECTED_165), .B(
        SYNOPSYS_UNCONNECTED_485), .Z(_f_permutation__round__n1508 ) );
  XOR2_X2 _f_permutation__round__U6130  ( .A(_f_permutation__round_in[1563]), 
        .B(_f_permutation__round_in[1243]), .Z(_f_permutation__round__n1509 )
         );
  XOR2_X2 _f_permutation__round__U6129  ( .A(_f_permutation__round__n1511 ), 
        .B(_f_permutation__round__n1510 ), .Z(_f_permutation__round__n2256 )
         );
  XOR2_X2 _f_permutation__round__U6128  ( .A(SYNOPSYS_UNCONNECTED_996), .B(
        _f_permutation__round__n1512 ), .Z(_f_permutation__round__n1510 ) );
  XOR2_X2 _f_permutation__round__U6127  ( .A(SYNOPSYS_UNCONNECTED_356), .B(
        SYNOPSYS_UNCONNECTED_676), .Z(_f_permutation__round__n1511 ) );
  XOR2_X2 _f_permutation__round__U6126  ( .A(_f_permutation__round_in[1372]), 
        .B(_f_permutation__round_in[1052]), .Z(_f_permutation__round__n1512 )
         );
  XOR2_X2 _f_permutation__round__U6125  ( .A(_f_permutation__round__n2036 ), 
        .B(_f_permutation__round__n2256 ), .Z(_f_permutation__round__n2037 )
         );
  XOR2_X2 _f_permutation__round__U6124  ( .A(SYNOPSYS_UNCONNECTED_1060), .B(
        _f_permutation__round__n2037 ), .Z(_f_permutation__round__c[1564] ) );
  XOR2_X2 _f_permutation__round__U6123  ( .A(_f_permutation__round__n1514 ), 
        .B(_f_permutation__round__n1513 ), .Z(_f_permutation__round__n2488 )
         );
  XOR2_X2 _f_permutation__round__U6122  ( .A(SYNOPSYS_UNCONNECTED_934), .B(
        _f_permutation__round__n1515 ), .Z(_f_permutation__round__n1513 ) );
  XOR2_X2 _f_permutation__round__U6121  ( .A(SYNOPSYS_UNCONNECTED_294), .B(
        SYNOPSYS_UNCONNECTED_614), .Z(_f_permutation__round__n1514 ) );
  XOR2_X2 _f_permutation__round__U6120  ( .A(_f_permutation__round_in[1434]), 
        .B(_f_permutation__round_in[1114]), .Z(_f_permutation__round__n1515 )
         );
  XOR2_X2 _f_permutation__round__U6119  ( .A(_f_permutation__round__n2036 ), 
        .B(_f_permutation__round__n2488 ), .Z(_f_permutation__round__n2038 )
         );
  XOR2_X2 _f_permutation__round__U6118  ( .A(SYNOPSYS_UNCONNECTED_869), .B(
        _f_permutation__round__n2038 ), .Z(_f_permutation__round__c[603] ) );
  XOR2_X2 _f_permutation__round__U6117  ( .A(SYNOPSYS_UNCONNECTED_740), .B(
        _f_permutation__round__n2037 ), .Z(_f_permutation__round__c[1500] ) );
  XOR2_X2 _f_permutation__round__U6116  ( .A(SYNOPSYS_UNCONNECTED_549), .B(
        _f_permutation__round__n2038 ), .Z(_f_permutation__round__c[539] ) );
  XOR2_X2 _f_permutation__round__U6115  ( .A(SYNOPSYS_UNCONNECTED_420), .B(
        _f_permutation__round__n2037 ), .Z(_f_permutation__round__c[1436] ) );
  XOR2_X2 _f_permutation__round__U6114  ( .A(SYNOPSYS_UNCONNECTED_229), .B(
        _f_permutation__round__n2038 ), .Z(_f_permutation__round__c[475] ) );
  XOR2_X2 _f_permutation__round__U6113  ( .A(SYNOPSYS_UNCONNECTED_100), .B(
        _f_permutation__round__n2037 ), .Z(_f_permutation__round__c[1372] ) );
  XOR2_X2 _f_permutation__round__U6112  ( .A(_f_permutation__round_in[1179]), 
        .B(_f_permutation__round__n2038 ), .Z(_f_permutation__round__c[411] )
         );
  XOR2_X2 _f_permutation__round__U6111  ( .A(_f_permutation__round_in[1308]), 
        .B(_f_permutation__round__n2037 ), .Z(_f_permutation__round__c[1308] )
         );
  XOR2_X2 _f_permutation__round__U6110  ( .A(_f_permutation__round_in[1499]), 
        .B(_f_permutation__round__n2038 ), .Z(_f_permutation__round__c[347] )
         );
  XOR2_X2 _f_permutation__round__U6109  ( .A(_f_permutation__round__n1517 ), 
        .B(_f_permutation__round__n1516 ), .Z(_f_permutation__round__n2273 )
         );
  XOR2_X2 _f_permutation__round__U6108  ( .A(SYNOPSYS_UNCONNECTED_871), .B(
        _f_permutation__round__n1518 ), .Z(_f_permutation__round__n1516 ) );
  XOR2_X2 _f_permutation__round__U6107  ( .A(SYNOPSYS_UNCONNECTED_231), .B(
        SYNOPSYS_UNCONNECTED_551), .Z(_f_permutation__round__n1517 ) );
  XOR2_X2 _f_permutation__round__U6106  ( .A(_f_permutation__round_in[1497]), 
        .B(_f_permutation__round_in[1177]), .Z(_f_permutation__round__n1518 )
         );
  XOR2_X2 _f_permutation__round__U6105  ( .A(_f_permutation__round__n1520 ), 
        .B(_f_permutation__round__n1519 ), .Z(_f_permutation__round__n2484 )
         );
  XOR2_X2 _f_permutation__round__U6104  ( .A(SYNOPSYS_UNCONNECTED_1062), .B(
        _f_permutation__round__n1521 ), .Z(_f_permutation__round__n1519 ) );
  XOR2_X2 _f_permutation__round__U6103  ( .A(SYNOPSYS_UNCONNECTED_422), .B(
        SYNOPSYS_UNCONNECTED_742), .Z(_f_permutation__round__n1520 ) );
  XOR2_X2 _f_permutation__round__U6102  ( .A(_f_permutation__round_in[1306]), 
        .B(SYNOPSYS_UNCONNECTED_102), .Z(_f_permutation__round__n1521 ) );
  XOR2_X2 _f_permutation__round__U6101  ( .A(_f_permutation__round__n2273 ), 
        .B(_f_permutation__round__n2484 ), .Z(_f_permutation__round__n2274 )
         );
  XOR2_X2 _f_permutation__round__U6100  ( .A(_f_permutation__round_in[1562]), 
        .B(_f_permutation__round__n2274 ), .Z(_f_permutation__round__c[26] )
         );
  XOR2_X2 _f_permutation__round__U6099  ( .A(_f_permutation__round__n1523 ), 
        .B(_f_permutation__round__n1522 ), .Z(_f_permutation__round__n2039 )
         );
  XOR2_X2 _f_permutation__round__U6098  ( .A(SYNOPSYS_UNCONNECTED_806), .B(
        _f_permutation__round__n1524 ), .Z(_f_permutation__round__n1522 ) );
  XOR2_X2 _f_permutation__round__U6097  ( .A(SYNOPSYS_UNCONNECTED_166), .B(
        SYNOPSYS_UNCONNECTED_486), .Z(_f_permutation__round__n1523 ) );
  XOR2_X2 _f_permutation__round__U6096  ( .A(_f_permutation__round_in[1562]), 
        .B(_f_permutation__round_in[1242]), .Z(_f_permutation__round__n1524 )
         );
  XOR2_X2 _f_permutation__round__U6095  ( .A(_f_permutation__round__n1526 ), 
        .B(_f_permutation__round__n1525 ), .Z(_f_permutation__round__n2260 )
         );
  XOR2_X2 _f_permutation__round__U6094  ( .A(SYNOPSYS_UNCONNECTED_997), .B(
        _f_permutation__round__n1527 ), .Z(_f_permutation__round__n1525 ) );
  XOR2_X2 _f_permutation__round__U6093  ( .A(SYNOPSYS_UNCONNECTED_357), .B(
        SYNOPSYS_UNCONNECTED_677), .Z(_f_permutation__round__n1526 ) );
  XOR2_X2 _f_permutation__round__U6092  ( .A(_f_permutation__round_in[1371]), 
        .B(_f_permutation__round_in[1051]), .Z(_f_permutation__round__n1527 )
         );
  XOR2_X2 _f_permutation__round__U6091  ( .A(_f_permutation__round__n2039 ), 
        .B(_f_permutation__round__n2260 ), .Z(_f_permutation__round__n2040 )
         );
  XOR2_X2 _f_permutation__round__U6090  ( .A(SYNOPSYS_UNCONNECTED_1061), .B(
        _f_permutation__round__n2040 ), .Z(_f_permutation__round__c[1563] ) );
  XOR2_X2 _f_permutation__round__U6089  ( .A(_f_permutation__round__n1529 ), 
        .B(_f_permutation__round__n1528 ), .Z(_f_permutation__round__n2491 )
         );
  XOR2_X2 _f_permutation__round__U6088  ( .A(SYNOPSYS_UNCONNECTED_935), .B(
        _f_permutation__round__n1530 ), .Z(_f_permutation__round__n1528 ) );
  XOR2_X2 _f_permutation__round__U6087  ( .A(SYNOPSYS_UNCONNECTED_295), .B(
        SYNOPSYS_UNCONNECTED_615), .Z(_f_permutation__round__n1529 ) );
  XOR2_X2 _f_permutation__round__U6086  ( .A(_f_permutation__round_in[1433]), 
        .B(_f_permutation__round_in[1113]), .Z(_f_permutation__round__n1530 )
         );
  XOR2_X2 _f_permutation__round__U6085  ( .A(_f_permutation__round__n2039 ), 
        .B(_f_permutation__round__n2491 ), .Z(_f_permutation__round__n2041 )
         );
  XOR2_X2 _f_permutation__round__U6084  ( .A(SYNOPSYS_UNCONNECTED_870), .B(
        _f_permutation__round__n2041 ), .Z(_f_permutation__round__c[602] ) );
  XOR2_X2 _f_permutation__round__U6083  ( .A(SYNOPSYS_UNCONNECTED_741), .B(
        _f_permutation__round__n2040 ), .Z(_f_permutation__round__c[1499] ) );
  XOR2_X2 _f_permutation__round__U6082  ( .A(SYNOPSYS_UNCONNECTED_550), .B(
        _f_permutation__round__n2041 ), .Z(_f_permutation__round__c[538] ) );
  XOR2_X2 _f_permutation__round__U6081  ( .A(SYNOPSYS_UNCONNECTED_421), .B(
        _f_permutation__round__n2040 ), .Z(_f_permutation__round__c[1435] ) );
  XOR2_X2 _f_permutation__round__U6080  ( .A(SYNOPSYS_UNCONNECTED_230), .B(
        _f_permutation__round__n2041 ), .Z(_f_permutation__round__c[474] ) );
  XOR2_X2 _f_permutation__round__U6079  ( .A(SYNOPSYS_UNCONNECTED_101), .B(
        _f_permutation__round__n2040 ), .Z(_f_permutation__round__c[1371] ) );
  XOR2_X2 _f_permutation__round__U6078  ( .A(_f_permutation__round_in[1178]), 
        .B(_f_permutation__round__n2041 ), .Z(_f_permutation__round__c[410] )
         );
  XOR2_X2 _f_permutation__round__U6077  ( .A(_f_permutation__round_in[1307]), 
        .B(_f_permutation__round__n2040 ), .Z(_f_permutation__round__c[1307] )
         );
  XOR2_X2 _f_permutation__round__U6076  ( .A(_f_permutation__round_in[1498]), 
        .B(_f_permutation__round__n2041 ), .Z(_f_permutation__round__c[346] )
         );
  XOR2_X2 _f_permutation__round__U6075  ( .A(_f_permutation__round__n1532 ), 
        .B(_f_permutation__round__n1531 ), .Z(_f_permutation__round__n2277 )
         );
  XOR2_X2 _f_permutation__round__U6074  ( .A(SYNOPSYS_UNCONNECTED_872), .B(
        _f_permutation__round__n1533 ), .Z(_f_permutation__round__n1531 ) );
  XOR2_X2 _f_permutation__round__U6073  ( .A(SYNOPSYS_UNCONNECTED_232), .B(
        SYNOPSYS_UNCONNECTED_552), .Z(_f_permutation__round__n1532 ) );
  XOR2_X2 _f_permutation__round__U6072  ( .A(_f_permutation__round_in[1496]), 
        .B(_f_permutation__round_in[1176]), .Z(_f_permutation__round__n1533 )
         );
  XOR2_X2 _f_permutation__round__U6071  ( .A(_f_permutation__round__n1535 ), 
        .B(_f_permutation__round__n1534 ), .Z(_f_permutation__round__n2487 )
         );
  XOR2_X2 _f_permutation__round__U6070  ( .A(SYNOPSYS_UNCONNECTED_1063), .B(
        _f_permutation__round__n1536 ), .Z(_f_permutation__round__n1534 ) );
  XOR2_X2 _f_permutation__round__U6069  ( .A(SYNOPSYS_UNCONNECTED_423), .B(
        SYNOPSYS_UNCONNECTED_743), .Z(_f_permutation__round__n1535 ) );
  XOR2_X2 _f_permutation__round__U6068  ( .A(_f_permutation__round_in[1305]), 
        .B(SYNOPSYS_UNCONNECTED_103), .Z(_f_permutation__round__n1536 ) );
  XOR2_X2 _f_permutation__round__U6067  ( .A(_f_permutation__round__n2277 ), 
        .B(_f_permutation__round__n2487 ), .Z(_f_permutation__round__n2278 )
         );
  XOR2_X2 _f_permutation__round__U6066  ( .A(_f_permutation__round_in[1561]), 
        .B(_f_permutation__round__n2278 ), .Z(_f_permutation__round__c[25] )
         );
  XOR2_X2 _f_permutation__round__U6065  ( .A(_f_permutation__round__n1538 ), 
        .B(_f_permutation__round__n1537 ), .Z(_f_permutation__round__n2042 )
         );
  XOR2_X2 _f_permutation__round__U6064  ( .A(SYNOPSYS_UNCONNECTED_807), .B(
        _f_permutation__round__n1539 ), .Z(_f_permutation__round__n1537 ) );
  XOR2_X2 _f_permutation__round__U6063  ( .A(SYNOPSYS_UNCONNECTED_167), .B(
        SYNOPSYS_UNCONNECTED_487), .Z(_f_permutation__round__n1538 ) );
  XOR2_X2 _f_permutation__round__U6062  ( .A(_f_permutation__round_in[1561]), 
        .B(_f_permutation__round_in[1241]), .Z(_f_permutation__round__n1539 )
         );
  XOR2_X2 _f_permutation__round__U6061  ( .A(_f_permutation__round__n1541 ), 
        .B(_f_permutation__round__n1540 ), .Z(_f_permutation__round__n2264 )
         );
  XOR2_X2 _f_permutation__round__U6060  ( .A(SYNOPSYS_UNCONNECTED_998), .B(
        _f_permutation__round__n1542 ), .Z(_f_permutation__round__n1540 ) );
  XOR2_X2 _f_permutation__round__U6059  ( .A(SYNOPSYS_UNCONNECTED_358), .B(
        SYNOPSYS_UNCONNECTED_678), .Z(_f_permutation__round__n1541 ) );
  XOR2_X2 _f_permutation__round__U6058  ( .A(_f_permutation__round_in[1370]), 
        .B(_f_permutation__round_in[1050]), .Z(_f_permutation__round__n1542 )
         );
  XOR2_X2 _f_permutation__round__U6057  ( .A(_f_permutation__round__n2042 ), 
        .B(_f_permutation__round__n2264 ), .Z(_f_permutation__round__n2043 )
         );
  XOR2_X2 _f_permutation__round__U6056  ( .A(SYNOPSYS_UNCONNECTED_1062), .B(
        _f_permutation__round__n2043 ), .Z(_f_permutation__round__c[1562] ) );
  XOR2_X2 _f_permutation__round__U6055  ( .A(_f_permutation__round__n1544 ), 
        .B(_f_permutation__round__n1543 ), .Z(_f_permutation__round__n2494 )
         );
  XOR2_X2 _f_permutation__round__U6054  ( .A(SYNOPSYS_UNCONNECTED_936), .B(
        _f_permutation__round__n1545 ), .Z(_f_permutation__round__n1543 ) );
  XOR2_X2 _f_permutation__round__U6053  ( .A(SYNOPSYS_UNCONNECTED_296), .B(
        SYNOPSYS_UNCONNECTED_616), .Z(_f_permutation__round__n1544 ) );
  XOR2_X2 _f_permutation__round__U6052  ( .A(_f_permutation__round_in[1432]), 
        .B(_f_permutation__round_in[1112]), .Z(_f_permutation__round__n1545 )
         );
  XOR2_X2 _f_permutation__round__U6051  ( .A(_f_permutation__round__n2042 ), 
        .B(_f_permutation__round__n2494 ), .Z(_f_permutation__round__n2044 )
         );
  XOR2_X2 _f_permutation__round__U6050  ( .A(SYNOPSYS_UNCONNECTED_871), .B(
        _f_permutation__round__n2044 ), .Z(_f_permutation__round__c[601] ) );
  XOR2_X2 _f_permutation__round__U6049  ( .A(SYNOPSYS_UNCONNECTED_742), .B(
        _f_permutation__round__n2043 ), .Z(_f_permutation__round__c[1498] ) );
  XOR2_X2 _f_permutation__round__U6048  ( .A(SYNOPSYS_UNCONNECTED_551), .B(
        _f_permutation__round__n2044 ), .Z(_f_permutation__round__c[537] ) );
  XOR2_X2 _f_permutation__round__U6047  ( .A(SYNOPSYS_UNCONNECTED_422), .B(
        _f_permutation__round__n2043 ), .Z(_f_permutation__round__c[1434] ) );
  XOR2_X2 _f_permutation__round__U6046  ( .A(SYNOPSYS_UNCONNECTED_231), .B(
        _f_permutation__round__n2044 ), .Z(_f_permutation__round__c[473] ) );
  XOR2_X2 _f_permutation__round__U6045  ( .A(SYNOPSYS_UNCONNECTED_102), .B(
        _f_permutation__round__n2043 ), .Z(_f_permutation__round__c[1370] ) );
  XOR2_X2 _f_permutation__round__U6044  ( .A(_f_permutation__round_in[1177]), 
        .B(_f_permutation__round__n2044 ), .Z(_f_permutation__round__c[409] )
         );
  XOR2_X2 _f_permutation__round__U6043  ( .A(_f_permutation__round_in[1306]), 
        .B(_f_permutation__round__n2043 ), .Z(_f_permutation__round__c[1306] )
         );
  XOR2_X2 _f_permutation__round__U6042  ( .A(_f_permutation__round_in[1497]), 
        .B(_f_permutation__round__n2044 ), .Z(_f_permutation__round__c[345] )
         );
  XOR2_X2 _f_permutation__round__U6041  ( .A(_f_permutation__round__n1547 ), 
        .B(_f_permutation__round__n1546 ), .Z(_f_permutation__round__n2281 )
         );
  XOR2_X2 _f_permutation__round__U6040  ( .A(SYNOPSYS_UNCONNECTED_873), .B(
        _f_permutation__round__n1548 ), .Z(_f_permutation__round__n1546 ) );
  XOR2_X2 _f_permutation__round__U6039  ( .A(SYNOPSYS_UNCONNECTED_233), .B(
        SYNOPSYS_UNCONNECTED_553), .Z(_f_permutation__round__n1547 ) );
  XOR2_X2 _f_permutation__round__U6038  ( .A(_f_permutation__round_in[1495]), 
        .B(_f_permutation__round_in[1175]), .Z(_f_permutation__round__n1548 )
         );
  XOR2_X2 _f_permutation__round__U6037  ( .A(_f_permutation__round__n1550 ), 
        .B(_f_permutation__round__n1549 ), .Z(_f_permutation__round__n2490 )
         );
  XOR2_X2 _f_permutation__round__U6036  ( .A(SYNOPSYS_UNCONNECTED_1064), .B(
        _f_permutation__round__n1551 ), .Z(_f_permutation__round__n1549 ) );
  XOR2_X2 _f_permutation__round__U6035  ( .A(SYNOPSYS_UNCONNECTED_424), .B(
        SYNOPSYS_UNCONNECTED_744), .Z(_f_permutation__round__n1550 ) );
  XOR2_X2 _f_permutation__round__U6034  ( .A(_f_permutation__round_in[1304]), 
        .B(SYNOPSYS_UNCONNECTED_104), .Z(_f_permutation__round__n1551 ) );
  XOR2_X2 _f_permutation__round__U6033  ( .A(_f_permutation__round__n2281 ), 
        .B(_f_permutation__round__n2490 ), .Z(_f_permutation__round__n2282 )
         );
  XOR2_X2 _f_permutation__round__U6032  ( .A(_f_permutation__round_in[1560]), 
        .B(_f_permutation__round__n2282 ), .Z(_f_permutation__round__c[24] )
         );
  XOR2_X2 _f_permutation__round__U6031  ( .A(_f_permutation__round__n1553 ), 
        .B(_f_permutation__round__n1552 ), .Z(_f_permutation__round__n2045 )
         );
  XOR2_X2 _f_permutation__round__U6030  ( .A(SYNOPSYS_UNCONNECTED_808), .B(
        _f_permutation__round__n1554 ), .Z(_f_permutation__round__n1552 ) );
  XOR2_X2 _f_permutation__round__U6029  ( .A(SYNOPSYS_UNCONNECTED_168), .B(
        SYNOPSYS_UNCONNECTED_488), .Z(_f_permutation__round__n1553 ) );
  XOR2_X2 _f_permutation__round__U6028  ( .A(_f_permutation__round_in[1560]), 
        .B(_f_permutation__round_in[1240]), .Z(_f_permutation__round__n1554 )
         );
  XOR2_X2 _f_permutation__round__U6027  ( .A(_f_permutation__round__n1556 ), 
        .B(_f_permutation__round__n1555 ), .Z(_f_permutation__round__n2268 )
         );
  XOR2_X2 _f_permutation__round__U6026  ( .A(SYNOPSYS_UNCONNECTED_999), .B(
        _f_permutation__round__n1557 ), .Z(_f_permutation__round__n1555 ) );
  XOR2_X2 _f_permutation__round__U6025  ( .A(SYNOPSYS_UNCONNECTED_359), .B(
        SYNOPSYS_UNCONNECTED_679), .Z(_f_permutation__round__n1556 ) );
  XOR2_X2 _f_permutation__round__U6024  ( .A(_f_permutation__round_in[1369]), 
        .B(_f_permutation__round_in[1049]), .Z(_f_permutation__round__n1557 )
         );
  XOR2_X2 _f_permutation__round__U6023  ( .A(_f_permutation__round__n2045 ), 
        .B(_f_permutation__round__n2268 ), .Z(_f_permutation__round__n2046 )
         );
  XOR2_X2 _f_permutation__round__U6022  ( .A(SYNOPSYS_UNCONNECTED_1063), .B(
        _f_permutation__round__n2046 ), .Z(_f_permutation__round__c[1561] ) );
  XOR2_X2 _f_permutation__round__U6021  ( .A(_f_permutation__round__n1559 ), 
        .B(_f_permutation__round__n1558 ), .Z(_f_permutation__round__n2497 )
         );
  XOR2_X2 _f_permutation__round__U6020  ( .A(SYNOPSYS_UNCONNECTED_937), .B(
        _f_permutation__round__n1560 ), .Z(_f_permutation__round__n1558 ) );
  XOR2_X2 _f_permutation__round__U6019  ( .A(SYNOPSYS_UNCONNECTED_297), .B(
        SYNOPSYS_UNCONNECTED_617), .Z(_f_permutation__round__n1559 ) );
  XOR2_X2 _f_permutation__round__U6018  ( .A(_f_permutation__round_in[1431]), 
        .B(_f_permutation__round_in[1111]), .Z(_f_permutation__round__n1560 )
         );
  XOR2_X2 _f_permutation__round__U6017  ( .A(_f_permutation__round__n2045 ), 
        .B(_f_permutation__round__n2497 ), .Z(_f_permutation__round__n2047 )
         );
  XOR2_X2 _f_permutation__round__U6016  ( .A(SYNOPSYS_UNCONNECTED_872), .B(
        _f_permutation__round__n2047 ), .Z(_f_permutation__round__c[600] ) );
  XOR2_X2 _f_permutation__round__U6015  ( .A(SYNOPSYS_UNCONNECTED_743), .B(
        _f_permutation__round__n2046 ), .Z(_f_permutation__round__c[1497] ) );
  XOR2_X2 _f_permutation__round__U6014  ( .A(SYNOPSYS_UNCONNECTED_552), .B(
        _f_permutation__round__n2047 ), .Z(_f_permutation__round__c[536] ) );
  XOR2_X2 _f_permutation__round__U6013  ( .A(SYNOPSYS_UNCONNECTED_423), .B(
        _f_permutation__round__n2046 ), .Z(_f_permutation__round__c[1433] ) );
  XOR2_X2 _f_permutation__round__U6012  ( .A(SYNOPSYS_UNCONNECTED_232), .B(
        _f_permutation__round__n2047 ), .Z(_f_permutation__round__c[472] ) );
  XOR2_X2 _f_permutation__round__U6011  ( .A(SYNOPSYS_UNCONNECTED_103), .B(
        _f_permutation__round__n2046 ), .Z(_f_permutation__round__c[1369] ) );
  XOR2_X2 _f_permutation__round__U6010  ( .A(_f_permutation__round_in[1176]), 
        .B(_f_permutation__round__n2047 ), .Z(_f_permutation__round__c[408] )
         );
  XOR2_X2 _f_permutation__round__U6009  ( .A(_f_permutation__round_in[1305]), 
        .B(_f_permutation__round__n2046 ), .Z(_f_permutation__round__c[1305] )
         );
  XOR2_X2 _f_permutation__round__U6008  ( .A(_f_permutation__round_in[1496]), 
        .B(_f_permutation__round__n2047 ), .Z(_f_permutation__round__c[344] )
         );
  XOR2_X2 _f_permutation__round__U6007  ( .A(_f_permutation__round__n1562 ), 
        .B(_f_permutation__round__n1561 ), .Z(_f_permutation__round__n2285 )
         );
  XOR2_X2 _f_permutation__round__U6006  ( .A(SYNOPSYS_UNCONNECTED_874), .B(
        _f_permutation__round__n1563 ), .Z(_f_permutation__round__n1561 ) );
  XOR2_X2 _f_permutation__round__U6005  ( .A(SYNOPSYS_UNCONNECTED_234), .B(
        SYNOPSYS_UNCONNECTED_554), .Z(_f_permutation__round__n1562 ) );
  XOR2_X2 _f_permutation__round__U6004  ( .A(_f_permutation__round_in[1494]), 
        .B(_f_permutation__round_in[1174]), .Z(_f_permutation__round__n1563 )
         );
  XOR2_X2 _f_permutation__round__U6003  ( .A(_f_permutation__round__n1565 ), 
        .B(_f_permutation__round__n1564 ), .Z(_f_permutation__round__n2493 )
         );
  XOR2_X2 _f_permutation__round__U6002  ( .A(SYNOPSYS_UNCONNECTED_1065), .B(
        _f_permutation__round__n1566 ), .Z(_f_permutation__round__n1564 ) );
  XOR2_X2 _f_permutation__round__U6001  ( .A(SYNOPSYS_UNCONNECTED_425), .B(
        SYNOPSYS_UNCONNECTED_745), .Z(_f_permutation__round__n1565 ) );
  XOR2_X2 _f_permutation__round__U6000  ( .A(_f_permutation__round_in[1303]), 
        .B(SYNOPSYS_UNCONNECTED_105), .Z(_f_permutation__round__n1566 ) );
  XOR2_X2 _f_permutation__round__U5999  ( .A(_f_permutation__round__n2285 ), 
        .B(_f_permutation__round__n2493 ), .Z(_f_permutation__round__n2286 )
         );
  XOR2_X2 _f_permutation__round__U5998  ( .A(_f_permutation__round_in[1559]), 
        .B(_f_permutation__round__n2286 ), .Z(_f_permutation__round__c[23] )
         );
  XOR2_X2 _f_permutation__round__U5997  ( .A(_f_permutation__round__n1568 ), 
        .B(_f_permutation__round__n1567 ), .Z(_f_permutation__round__n2048 )
         );
  XOR2_X2 _f_permutation__round__U5996  ( .A(SYNOPSYS_UNCONNECTED_809), .B(
        _f_permutation__round__n1569 ), .Z(_f_permutation__round__n1567 ) );
  XOR2_X2 _f_permutation__round__U5995  ( .A(SYNOPSYS_UNCONNECTED_169), .B(
        SYNOPSYS_UNCONNECTED_489), .Z(_f_permutation__round__n1568 ) );
  XOR2_X2 _f_permutation__round__U5994  ( .A(_f_permutation__round_in[1559]), 
        .B(_f_permutation__round_in[1239]), .Z(_f_permutation__round__n1569 )
         );
  XOR2_X2 _f_permutation__round__U5993  ( .A(_f_permutation__round__n1571 ), 
        .B(_f_permutation__round__n1570 ), .Z(_f_permutation__round__n2272 )
         );
  XOR2_X2 _f_permutation__round__U5992  ( .A(SYNOPSYS_UNCONNECTED_1000), .B(
        _f_permutation__round__n1572 ), .Z(_f_permutation__round__n1570 ) );
  XOR2_X2 _f_permutation__round__U5991  ( .A(SYNOPSYS_UNCONNECTED_360), .B(
        SYNOPSYS_UNCONNECTED_680), .Z(_f_permutation__round__n1571 ) );
  XOR2_X2 _f_permutation__round__U5990  ( .A(_f_permutation__round_in[1368]), 
        .B(_f_permutation__round_in[1048]), .Z(_f_permutation__round__n1572 )
         );
  XOR2_X2 _f_permutation__round__U5989  ( .A(_f_permutation__round__n2048 ), 
        .B(_f_permutation__round__n2272 ), .Z(_f_permutation__round__n2049 )
         );
  XOR2_X2 _f_permutation__round__U5988  ( .A(SYNOPSYS_UNCONNECTED_1064), .B(
        _f_permutation__round__n2049 ), .Z(_f_permutation__round__c[1560] ) );
  XOR2_X2 _f_permutation__round__U5987  ( .A(_f_permutation__round__n1574 ), 
        .B(_f_permutation__round__n1573 ), .Z(_f_permutation__round__n2500 )
         );
  XOR2_X2 _f_permutation__round__U5986  ( .A(SYNOPSYS_UNCONNECTED_938), .B(
        _f_permutation__round__n1575 ), .Z(_f_permutation__round__n1573 ) );
  XOR2_X2 _f_permutation__round__U5985  ( .A(SYNOPSYS_UNCONNECTED_298), .B(
        SYNOPSYS_UNCONNECTED_618), .Z(_f_permutation__round__n1574 ) );
  XOR2_X2 _f_permutation__round__U5984  ( .A(_f_permutation__round_in[1430]), 
        .B(_f_permutation__round_in[1110]), .Z(_f_permutation__round__n1575 )
         );
  XOR2_X2 _f_permutation__round__U5983  ( .A(_f_permutation__round__n2048 ), 
        .B(_f_permutation__round__n2500 ), .Z(_f_permutation__round__n2050 )
         );
  XOR2_X2 _f_permutation__round__U5982  ( .A(SYNOPSYS_UNCONNECTED_873), .B(
        _f_permutation__round__n2050 ), .Z(_f_permutation__round__c[599] ) );
  XOR2_X2 _f_permutation__round__U5981  ( .A(SYNOPSYS_UNCONNECTED_744), .B(
        _f_permutation__round__n2049 ), .Z(_f_permutation__round__c[1496] ) );
  XOR2_X2 _f_permutation__round__U5980  ( .A(SYNOPSYS_UNCONNECTED_553), .B(
        _f_permutation__round__n2050 ), .Z(_f_permutation__round__c[535] ) );
  XOR2_X2 _f_permutation__round__U5979  ( .A(SYNOPSYS_UNCONNECTED_424), .B(
        _f_permutation__round__n2049 ), .Z(_f_permutation__round__c[1432] ) );
  XOR2_X2 _f_permutation__round__U5978  ( .A(SYNOPSYS_UNCONNECTED_233), .B(
        _f_permutation__round__n2050 ), .Z(_f_permutation__round__c[471] ) );
  XOR2_X2 _f_permutation__round__U5977  ( .A(SYNOPSYS_UNCONNECTED_104), .B(
        _f_permutation__round__n2049 ), .Z(_f_permutation__round__c[1368] ) );
  XOR2_X2 _f_permutation__round__U5976  ( .A(_f_permutation__round_in[1175]), 
        .B(_f_permutation__round__n2050 ), .Z(_f_permutation__round__c[407] )
         );
  XOR2_X2 _f_permutation__round__U5975  ( .A(_f_permutation__round_in[1304]), 
        .B(_f_permutation__round__n2049 ), .Z(_f_permutation__round__c[1304] )
         );
  XOR2_X2 _f_permutation__round__U5974  ( .A(_f_permutation__round_in[1495]), 
        .B(_f_permutation__round__n2050 ), .Z(_f_permutation__round__c[343] )
         );
  XOR2_X2 _f_permutation__round__U5973  ( .A(_f_permutation__round__n1577 ), 
        .B(_f_permutation__round__n1576 ), .Z(_f_permutation__round__n2289 )
         );
  XOR2_X2 _f_permutation__round__U5972  ( .A(SYNOPSYS_UNCONNECTED_875), .B(
        _f_permutation__round__n1578 ), .Z(_f_permutation__round__n1576 ) );
  XOR2_X2 _f_permutation__round__U5971  ( .A(SYNOPSYS_UNCONNECTED_235), .B(
        SYNOPSYS_UNCONNECTED_555), .Z(_f_permutation__round__n1577 ) );
  XOR2_X2 _f_permutation__round__U5970  ( .A(_f_permutation__round_in[1493]), 
        .B(_f_permutation__round_in[1173]), .Z(_f_permutation__round__n1578 )
         );
  XOR2_X2 _f_permutation__round__U5969  ( .A(_f_permutation__round__n1580 ), 
        .B(_f_permutation__round__n1579 ), .Z(_f_permutation__round__n2496 )
         );
  XOR2_X2 _f_permutation__round__U5968  ( .A(SYNOPSYS_UNCONNECTED_1066), .B(
        _f_permutation__round__n1581 ), .Z(_f_permutation__round__n1579 ) );
  XOR2_X2 _f_permutation__round__U5967  ( .A(SYNOPSYS_UNCONNECTED_426), .B(
        SYNOPSYS_UNCONNECTED_746), .Z(_f_permutation__round__n1580 ) );
  XOR2_X2 _f_permutation__round__U5966  ( .A(_f_permutation__round_in[1302]), 
        .B(SYNOPSYS_UNCONNECTED_106), .Z(_f_permutation__round__n1581 ) );
  XOR2_X2 _f_permutation__round__U5965  ( .A(_f_permutation__round__n2289 ), 
        .B(_f_permutation__round__n2496 ), .Z(_f_permutation__round__n2290 )
         );
  XOR2_X2 _f_permutation__round__U5964  ( .A(_f_permutation__round_in[1558]), 
        .B(_f_permutation__round__n2290 ), .Z(_f_permutation__round__c[22] )
         );
  XOR2_X2 _f_permutation__round__U5963  ( .A(_f_permutation__round__n1583 ), 
        .B(_f_permutation__round__n1582 ), .Z(_f_permutation__round__n2051 )
         );
  XOR2_X2 _f_permutation__round__U5962  ( .A(SYNOPSYS_UNCONNECTED_810), .B(
        _f_permutation__round__n1584 ), .Z(_f_permutation__round__n1582 ) );
  XOR2_X2 _f_permutation__round__U5961  ( .A(SYNOPSYS_UNCONNECTED_170), .B(
        SYNOPSYS_UNCONNECTED_490), .Z(_f_permutation__round__n1583 ) );
  XOR2_X2 _f_permutation__round__U5960  ( .A(_f_permutation__round_in[1558]), 
        .B(_f_permutation__round_in[1238]), .Z(_f_permutation__round__n1584 )
         );
  XOR2_X2 _f_permutation__round__U5959  ( .A(_f_permutation__round__n1586 ), 
        .B(_f_permutation__round__n1585 ), .Z(_f_permutation__round__n2276 )
         );
  XOR2_X2 _f_permutation__round__U5958  ( .A(SYNOPSYS_UNCONNECTED_1001), .B(
        _f_permutation__round__n1587 ), .Z(_f_permutation__round__n1585 ) );
  XOR2_X2 _f_permutation__round__U5957  ( .A(SYNOPSYS_UNCONNECTED_361), .B(
        SYNOPSYS_UNCONNECTED_681), .Z(_f_permutation__round__n1586 ) );
  XOR2_X2 _f_permutation__round__U5956  ( .A(_f_permutation__round_in[1367]), 
        .B(_f_permutation__round_in[1047]), .Z(_f_permutation__round__n1587 )
         );
  XOR2_X2 _f_permutation__round__U5955  ( .A(_f_permutation__round__n2051 ), 
        .B(_f_permutation__round__n2276 ), .Z(_f_permutation__round__n2052 )
         );
  XOR2_X2 _f_permutation__round__U5954  ( .A(SYNOPSYS_UNCONNECTED_1065), .B(
        _f_permutation__round__n2052 ), .Z(_f_permutation__round__c[1559] ) );
  XOR2_X2 _f_permutation__round__U5953  ( .A(_f_permutation__round__n1589 ), 
        .B(_f_permutation__round__n1588 ), .Z(_f_permutation__round__n2503 )
         );
  XOR2_X2 _f_permutation__round__U5952  ( .A(SYNOPSYS_UNCONNECTED_939), .B(
        _f_permutation__round__n1590 ), .Z(_f_permutation__round__n1588 ) );
  XOR2_X2 _f_permutation__round__U5951  ( .A(SYNOPSYS_UNCONNECTED_299), .B(
        SYNOPSYS_UNCONNECTED_619), .Z(_f_permutation__round__n1589 ) );
  XOR2_X2 _f_permutation__round__U5950  ( .A(_f_permutation__round_in[1429]), 
        .B(_f_permutation__round_in[1109]), .Z(_f_permutation__round__n1590 )
         );
  XOR2_X2 _f_permutation__round__U5949  ( .A(_f_permutation__round__n2051 ), 
        .B(_f_permutation__round__n2503 ), .Z(_f_permutation__round__n2053 )
         );
  XOR2_X2 _f_permutation__round__U5948  ( .A(SYNOPSYS_UNCONNECTED_874), .B(
        _f_permutation__round__n2053 ), .Z(_f_permutation__round__c[598] ) );
  XOR2_X2 _f_permutation__round__U5947  ( .A(SYNOPSYS_UNCONNECTED_745), .B(
        _f_permutation__round__n2052 ), .Z(_f_permutation__round__c[1495] ) );
  XOR2_X2 _f_permutation__round__U5946  ( .A(SYNOPSYS_UNCONNECTED_554), .B(
        _f_permutation__round__n2053 ), .Z(_f_permutation__round__c[534] ) );
  XOR2_X2 _f_permutation__round__U5945  ( .A(SYNOPSYS_UNCONNECTED_425), .B(
        _f_permutation__round__n2052 ), .Z(_f_permutation__round__c[1431] ) );
  XOR2_X2 _f_permutation__round__U5944  ( .A(SYNOPSYS_UNCONNECTED_234), .B(
        _f_permutation__round__n2053 ), .Z(_f_permutation__round__c[470] ) );
  XOR2_X2 _f_permutation__round__U5943  ( .A(SYNOPSYS_UNCONNECTED_105), .B(
        _f_permutation__round__n2052 ), .Z(_f_permutation__round__c[1367] ) );
  XOR2_X2 _f_permutation__round__U5942  ( .A(_f_permutation__round_in[1174]), 
        .B(_f_permutation__round__n2053 ), .Z(_f_permutation__round__c[406] )
         );
  XOR2_X2 _f_permutation__round__U5941  ( .A(_f_permutation__round_in[1303]), 
        .B(_f_permutation__round__n2052 ), .Z(_f_permutation__round__c[1303] )
         );
  XOR2_X2 _f_permutation__round__U5940  ( .A(_f_permutation__round_in[1494]), 
        .B(_f_permutation__round__n2053 ), .Z(_f_permutation__round__c[342] )
         );
  XOR2_X2 _f_permutation__round__U5939  ( .A(_f_permutation__round__n1592 ), 
        .B(_f_permutation__round__n1591 ), .Z(_f_permutation__round__n2293 )
         );
  XOR2_X2 _f_permutation__round__U5938  ( .A(SYNOPSYS_UNCONNECTED_876), .B(
        _f_permutation__round__n1593 ), .Z(_f_permutation__round__n1591 ) );
  XOR2_X2 _f_permutation__round__U5937  ( .A(SYNOPSYS_UNCONNECTED_236), .B(
        SYNOPSYS_UNCONNECTED_556), .Z(_f_permutation__round__n1592 ) );
  XOR2_X2 _f_permutation__round__U5936  ( .A(_f_permutation__round_in[1492]), 
        .B(_f_permutation__round_in[1172]), .Z(_f_permutation__round__n1593 )
         );
  XOR2_X2 _f_permutation__round__U5935  ( .A(_f_permutation__round__n1595 ), 
        .B(_f_permutation__round__n1594 ), .Z(_f_permutation__round__n2499 )
         );
  XOR2_X2 _f_permutation__round__U5934  ( .A(SYNOPSYS_UNCONNECTED_1067), .B(
        _f_permutation__round__n1596 ), .Z(_f_permutation__round__n1594 ) );
  XOR2_X2 _f_permutation__round__U5933  ( .A(SYNOPSYS_UNCONNECTED_427), .B(
        SYNOPSYS_UNCONNECTED_747), .Z(_f_permutation__round__n1595 ) );
  XOR2_X2 _f_permutation__round__U5932  ( .A(_f_permutation__round_in[1301]), 
        .B(SYNOPSYS_UNCONNECTED_107), .Z(_f_permutation__round__n1596 ) );
  XOR2_X2 _f_permutation__round__U5931  ( .A(_f_permutation__round__n2293 ), 
        .B(_f_permutation__round__n2499 ), .Z(_f_permutation__round__n2294 )
         );
  XOR2_X2 _f_permutation__round__U5930  ( .A(_f_permutation__round_in[1557]), 
        .B(_f_permutation__round__n2294 ), .Z(_f_permutation__round__c[21] )
         );
  XOR2_X2 _f_permutation__round__U5929  ( .A(_f_permutation__round__n1598 ), 
        .B(_f_permutation__round__n1597 ), .Z(_f_permutation__round__n2054 )
         );
  XOR2_X2 _f_permutation__round__U5928  ( .A(SYNOPSYS_UNCONNECTED_811), .B(
        _f_permutation__round__n1599 ), .Z(_f_permutation__round__n1597 ) );
  XOR2_X2 _f_permutation__round__U5927  ( .A(SYNOPSYS_UNCONNECTED_171), .B(
        SYNOPSYS_UNCONNECTED_491), .Z(_f_permutation__round__n1598 ) );
  XOR2_X2 _f_permutation__round__U5926  ( .A(_f_permutation__round_in[1557]), 
        .B(_f_permutation__round_in[1237]), .Z(_f_permutation__round__n1599 )
         );
  XOR2_X2 _f_permutation__round__U5925  ( .A(_f_permutation__round__n1601 ), 
        .B(_f_permutation__round__n1600 ), .Z(_f_permutation__round__n2280 )
         );
  XOR2_X2 _f_permutation__round__U5924  ( .A(SYNOPSYS_UNCONNECTED_1002), .B(
        _f_permutation__round__n1602 ), .Z(_f_permutation__round__n1600 ) );
  XOR2_X2 _f_permutation__round__U5923  ( .A(SYNOPSYS_UNCONNECTED_362), .B(
        SYNOPSYS_UNCONNECTED_682), .Z(_f_permutation__round__n1601 ) );
  XOR2_X2 _f_permutation__round__U5922  ( .A(_f_permutation__round_in[1366]), 
        .B(_f_permutation__round_in[1046]), .Z(_f_permutation__round__n1602 )
         );
  XOR2_X2 _f_permutation__round__U5921  ( .A(_f_permutation__round__n2054 ), 
        .B(_f_permutation__round__n2280 ), .Z(_f_permutation__round__n2055 )
         );
  XOR2_X2 _f_permutation__round__U5920  ( .A(SYNOPSYS_UNCONNECTED_1066), .B(
        _f_permutation__round__n2055 ), .Z(_f_permutation__round__c[1558] ) );
  XOR2_X2 _f_permutation__round__U5919  ( .A(_f_permutation__round__n1604 ), 
        .B(_f_permutation__round__n1603 ), .Z(_f_permutation__round__n2506 )
         );
  XOR2_X2 _f_permutation__round__U5918  ( .A(SYNOPSYS_UNCONNECTED_940), .B(
        _f_permutation__round__n1605 ), .Z(_f_permutation__round__n1603 ) );
  XOR2_X2 _f_permutation__round__U5917  ( .A(SYNOPSYS_UNCONNECTED_300), .B(
        SYNOPSYS_UNCONNECTED_620), .Z(_f_permutation__round__n1604 ) );
  XOR2_X2 _f_permutation__round__U5916  ( .A(_f_permutation__round_in[1428]), 
        .B(_f_permutation__round_in[1108]), .Z(_f_permutation__round__n1605 )
         );
  XOR2_X2 _f_permutation__round__U5915  ( .A(_f_permutation__round__n2054 ), 
        .B(_f_permutation__round__n2506 ), .Z(_f_permutation__round__n2056 )
         );
  XOR2_X2 _f_permutation__round__U5914  ( .A(SYNOPSYS_UNCONNECTED_875), .B(
        _f_permutation__round__n2056 ), .Z(_f_permutation__round__c[597] ) );
  XOR2_X2 _f_permutation__round__U5913  ( .A(SYNOPSYS_UNCONNECTED_746), .B(
        _f_permutation__round__n2055 ), .Z(_f_permutation__round__c[1494] ) );
  XOR2_X2 _f_permutation__round__U5912  ( .A(SYNOPSYS_UNCONNECTED_555), .B(
        _f_permutation__round__n2056 ), .Z(_f_permutation__round__c[533] ) );
  XOR2_X2 _f_permutation__round__U5911  ( .A(SYNOPSYS_UNCONNECTED_426), .B(
        _f_permutation__round__n2055 ), .Z(_f_permutation__round__c[1430] ) );
  XOR2_X2 _f_permutation__round__U5910  ( .A(SYNOPSYS_UNCONNECTED_235), .B(
        _f_permutation__round__n2056 ), .Z(_f_permutation__round__c[469] ) );
  XOR2_X2 _f_permutation__round__U5909  ( .A(SYNOPSYS_UNCONNECTED_106), .B(
        _f_permutation__round__n2055 ), .Z(_f_permutation__round__c[1366] ) );
  XOR2_X2 _f_permutation__round__U5908  ( .A(_f_permutation__round_in[1173]), 
        .B(_f_permutation__round__n2056 ), .Z(_f_permutation__round__c[405] )
         );
  XOR2_X2 _f_permutation__round__U5907  ( .A(_f_permutation__round_in[1302]), 
        .B(_f_permutation__round__n2055 ), .Z(_f_permutation__round__c[1302] )
         );
  XOR2_X2 _f_permutation__round__U5906  ( .A(_f_permutation__round_in[1493]), 
        .B(_f_permutation__round__n2056 ), .Z(_f_permutation__round__c[341] )
         );
  XOR2_X2 _f_permutation__round__U5905  ( .A(_f_permutation__round__n1607 ), 
        .B(_f_permutation__round__n1606 ), .Z(_f_permutation__round__n2297 )
         );
  XOR2_X2 _f_permutation__round__U5904  ( .A(SYNOPSYS_UNCONNECTED_877), .B(
        _f_permutation__round__n1608 ), .Z(_f_permutation__round__n1606 ) );
  XOR2_X2 _f_permutation__round__U5903  ( .A(SYNOPSYS_UNCONNECTED_237), .B(
        SYNOPSYS_UNCONNECTED_557), .Z(_f_permutation__round__n1607 ) );
  XOR2_X2 _f_permutation__round__U5902  ( .A(_f_permutation__round_in[1491]), 
        .B(_f_permutation__round_in[1171]), .Z(_f_permutation__round__n1608 )
         );
  XOR2_X2 _f_permutation__round__U5901  ( .A(_f_permutation__round__n1610 ), 
        .B(_f_permutation__round__n1609 ), .Z(_f_permutation__round__n2502 )
         );
  XOR2_X2 _f_permutation__round__U5900  ( .A(SYNOPSYS_UNCONNECTED_1068), .B(
        _f_permutation__round__n1611 ), .Z(_f_permutation__round__n1609 ) );
  XOR2_X2 _f_permutation__round__U5899  ( .A(SYNOPSYS_UNCONNECTED_428), .B(
        SYNOPSYS_UNCONNECTED_748), .Z(_f_permutation__round__n1610 ) );
  XOR2_X2 _f_permutation__round__U5898  ( .A(_f_permutation__round_in[1300]), 
        .B(SYNOPSYS_UNCONNECTED_108), .Z(_f_permutation__round__n1611 ) );
  XOR2_X2 _f_permutation__round__U5897  ( .A(_f_permutation__round__n2297 ), 
        .B(_f_permutation__round__n2502 ), .Z(_f_permutation__round__n2298 )
         );
  XOR2_X2 _f_permutation__round__U5896  ( .A(_f_permutation__round_in[1556]), 
        .B(_f_permutation__round__n2298 ), .Z(_f_permutation__round__c[20] )
         );
  XOR2_X2 _f_permutation__round__U5895  ( .A(_f_permutation__round__n1613 ), 
        .B(_f_permutation__round__n1612 ), .Z(_f_permutation__round__n2057 )
         );
  XOR2_X2 _f_permutation__round__U5894  ( .A(SYNOPSYS_UNCONNECTED_812), .B(
        _f_permutation__round__n1614 ), .Z(_f_permutation__round__n1612 ) );
  XOR2_X2 _f_permutation__round__U5893  ( .A(SYNOPSYS_UNCONNECTED_172), .B(
        SYNOPSYS_UNCONNECTED_492), .Z(_f_permutation__round__n1613 ) );
  XOR2_X2 _f_permutation__round__U5892  ( .A(_f_permutation__round_in[1556]), 
        .B(_f_permutation__round_in[1236]), .Z(_f_permutation__round__n1614 )
         );
  XOR2_X2 _f_permutation__round__U5891  ( .A(_f_permutation__round__n1616 ), 
        .B(_f_permutation__round__n1615 ), .Z(_f_permutation__round__n2284 )
         );
  XOR2_X2 _f_permutation__round__U5890  ( .A(SYNOPSYS_UNCONNECTED_1003), .B(
        _f_permutation__round__n1617 ), .Z(_f_permutation__round__n1615 ) );
  XOR2_X2 _f_permutation__round__U5889  ( .A(SYNOPSYS_UNCONNECTED_363), .B(
        SYNOPSYS_UNCONNECTED_683), .Z(_f_permutation__round__n1616 ) );
  XOR2_X2 _f_permutation__round__U5888  ( .A(_f_permutation__round_in[1365]), 
        .B(_f_permutation__round_in[1045]), .Z(_f_permutation__round__n1617 )
         );
  XOR2_X2 _f_permutation__round__U5887  ( .A(_f_permutation__round__n2057 ), 
        .B(_f_permutation__round__n2284 ), .Z(_f_permutation__round__n2058 )
         );
  XOR2_X2 _f_permutation__round__U5886  ( .A(SYNOPSYS_UNCONNECTED_1067), .B(
        _f_permutation__round__n2058 ), .Z(_f_permutation__round__c[1557] ) );
  XOR2_X2 _f_permutation__round__U5885  ( .A(_f_permutation__round__n1619 ), 
        .B(_f_permutation__round__n1618 ), .Z(_f_permutation__round__n2509 )
         );
  XOR2_X2 _f_permutation__round__U5884  ( .A(SYNOPSYS_UNCONNECTED_941), .B(
        _f_permutation__round__n1620 ), .Z(_f_permutation__round__n1618 ) );
  XOR2_X2 _f_permutation__round__U5883  ( .A(SYNOPSYS_UNCONNECTED_301), .B(
        SYNOPSYS_UNCONNECTED_621), .Z(_f_permutation__round__n1619 ) );
  XOR2_X2 _f_permutation__round__U5882  ( .A(_f_permutation__round_in[1427]), 
        .B(_f_permutation__round_in[1107]), .Z(_f_permutation__round__n1620 )
         );
  XOR2_X2 _f_permutation__round__U5881  ( .A(_f_permutation__round__n2057 ), 
        .B(_f_permutation__round__n2509 ), .Z(_f_permutation__round__n2059 )
         );
  XOR2_X2 _f_permutation__round__U5880  ( .A(SYNOPSYS_UNCONNECTED_876), .B(
        _f_permutation__round__n2059 ), .Z(_f_permutation__round__c[596] ) );
  XOR2_X2 _f_permutation__round__U5879  ( .A(SYNOPSYS_UNCONNECTED_747), .B(
        _f_permutation__round__n2058 ), .Z(_f_permutation__round__c[1493] ) );
  XOR2_X2 _f_permutation__round__U5878  ( .A(SYNOPSYS_UNCONNECTED_556), .B(
        _f_permutation__round__n2059 ), .Z(_f_permutation__round__c[532] ) );
  XOR2_X2 _f_permutation__round__U5877  ( .A(SYNOPSYS_UNCONNECTED_427), .B(
        _f_permutation__round__n2058 ), .Z(_f_permutation__round__c[1429] ) );
  XOR2_X2 _f_permutation__round__U5876  ( .A(SYNOPSYS_UNCONNECTED_236), .B(
        _f_permutation__round__n2059 ), .Z(_f_permutation__round__c[468] ) );
  XOR2_X2 _f_permutation__round__U5875  ( .A(SYNOPSYS_UNCONNECTED_107), .B(
        _f_permutation__round__n2058 ), .Z(_f_permutation__round__c[1365] ) );
  XOR2_X2 _f_permutation__round__U5874  ( .A(_f_permutation__round_in[1172]), 
        .B(_f_permutation__round__n2059 ), .Z(_f_permutation__round__c[404] )
         );
  XOR2_X2 _f_permutation__round__U5873  ( .A(_f_permutation__round_in[1301]), 
        .B(_f_permutation__round__n2058 ), .Z(_f_permutation__round__c[1301] )
         );
  XOR2_X2 _f_permutation__round__U5872  ( .A(_f_permutation__round_in[1492]), 
        .B(_f_permutation__round__n2059 ), .Z(_f_permutation__round__c[340] )
         );
  XOR2_X2 _f_permutation__round__U5871  ( .A(_f_permutation__round__n1622 ), 
        .B(_f_permutation__round__n1621 ), .Z(_f_permutation__round__n2301 )
         );
  XOR2_X2 _f_permutation__round__U5870  ( .A(SYNOPSYS_UNCONNECTED_878), .B(
        _f_permutation__round__n1623 ), .Z(_f_permutation__round__n1621 ) );
  XOR2_X2 _f_permutation__round__U5869  ( .A(SYNOPSYS_UNCONNECTED_238), .B(
        SYNOPSYS_UNCONNECTED_558), .Z(_f_permutation__round__n1622 ) );
  XOR2_X2 _f_permutation__round__U5868  ( .A(_f_permutation__round_in[1490]), 
        .B(_f_permutation__round_in[1170]), .Z(_f_permutation__round__n1623 )
         );
  XOR2_X2 _f_permutation__round__U5867  ( .A(_f_permutation__round__n1625 ), 
        .B(_f_permutation__round__n1624 ), .Z(_f_permutation__round__n2505 )
         );
  XOR2_X2 _f_permutation__round__U5866  ( .A(SYNOPSYS_UNCONNECTED_1069), .B(
        _f_permutation__round__n1626 ), .Z(_f_permutation__round__n1624 ) );
  XOR2_X2 _f_permutation__round__U5865  ( .A(SYNOPSYS_UNCONNECTED_429), .B(
        SYNOPSYS_UNCONNECTED_749), .Z(_f_permutation__round__n1625 ) );
  XOR2_X2 _f_permutation__round__U5864  ( .A(_f_permutation__round_in[1299]), 
        .B(SYNOPSYS_UNCONNECTED_109), .Z(_f_permutation__round__n1626 ) );
  XOR2_X2 _f_permutation__round__U5863  ( .A(_f_permutation__round__n2301 ), 
        .B(_f_permutation__round__n2505 ), .Z(_f_permutation__round__n2302 )
         );
  XOR2_X2 _f_permutation__round__U5862  ( .A(_f_permutation__round_in[1555]), 
        .B(_f_permutation__round__n2302 ), .Z(_f_permutation__round__c[19] )
         );
  XOR2_X2 _f_permutation__round__U5861  ( .A(_f_permutation__round__n1628 ), 
        .B(_f_permutation__round__n1627 ), .Z(_f_permutation__round__n2060 )
         );
  XOR2_X2 _f_permutation__round__U5860  ( .A(SYNOPSYS_UNCONNECTED_813), .B(
        _f_permutation__round__n1629 ), .Z(_f_permutation__round__n1627 ) );
  XOR2_X2 _f_permutation__round__U5859  ( .A(SYNOPSYS_UNCONNECTED_173), .B(
        SYNOPSYS_UNCONNECTED_493), .Z(_f_permutation__round__n1628 ) );
  XOR2_X2 _f_permutation__round__U5858  ( .A(_f_permutation__round_in[1555]), 
        .B(_f_permutation__round_in[1235]), .Z(_f_permutation__round__n1629 )
         );
  XOR2_X2 _f_permutation__round__U5857  ( .A(_f_permutation__round__n1631 ), 
        .B(_f_permutation__round__n1630 ), .Z(_f_permutation__round__n2288 )
         );
  XOR2_X2 _f_permutation__round__U5856  ( .A(SYNOPSYS_UNCONNECTED_1004), .B(
        _f_permutation__round__n1632 ), .Z(_f_permutation__round__n1630 ) );
  XOR2_X2 _f_permutation__round__U5855  ( .A(SYNOPSYS_UNCONNECTED_364), .B(
        SYNOPSYS_UNCONNECTED_684), .Z(_f_permutation__round__n1631 ) );
  XOR2_X2 _f_permutation__round__U5854  ( .A(_f_permutation__round_in[1364]), 
        .B(_f_permutation__round_in[1044]), .Z(_f_permutation__round__n1632 )
         );
  XOR2_X2 _f_permutation__round__U5853  ( .A(_f_permutation__round__n2060 ), 
        .B(_f_permutation__round__n2288 ), .Z(_f_permutation__round__n2061 )
         );
  XOR2_X2 _f_permutation__round__U5852  ( .A(SYNOPSYS_UNCONNECTED_1068), .B(
        _f_permutation__round__n2061 ), .Z(_f_permutation__round__c[1556] ) );
  XOR2_X2 _f_permutation__round__U5851  ( .A(_f_permutation__round__n1634 ), 
        .B(_f_permutation__round__n1633 ), .Z(_f_permutation__round__n2512 )
         );
  XOR2_X2 _f_permutation__round__U5850  ( .A(SYNOPSYS_UNCONNECTED_942), .B(
        _f_permutation__round__n1635 ), .Z(_f_permutation__round__n1633 ) );
  XOR2_X2 _f_permutation__round__U5849  ( .A(SYNOPSYS_UNCONNECTED_302), .B(
        SYNOPSYS_UNCONNECTED_622), .Z(_f_permutation__round__n1634 ) );
  XOR2_X2 _f_permutation__round__U5848  ( .A(_f_permutation__round_in[1426]), 
        .B(_f_permutation__round_in[1106]), .Z(_f_permutation__round__n1635 )
         );
  XOR2_X2 _f_permutation__round__U5847  ( .A(_f_permutation__round__n2060 ), 
        .B(_f_permutation__round__n2512 ), .Z(_f_permutation__round__n2062 )
         );
  XOR2_X2 _f_permutation__round__U5846  ( .A(SYNOPSYS_UNCONNECTED_877), .B(
        _f_permutation__round__n2062 ), .Z(_f_permutation__round__c[595] ) );
  XOR2_X2 _f_permutation__round__U5845  ( .A(SYNOPSYS_UNCONNECTED_748), .B(
        _f_permutation__round__n2061 ), .Z(_f_permutation__round__c[1492] ) );
  XOR2_X2 _f_permutation__round__U5844  ( .A(SYNOPSYS_UNCONNECTED_557), .B(
        _f_permutation__round__n2062 ), .Z(_f_permutation__round__c[531] ) );
  XOR2_X2 _f_permutation__round__U5843  ( .A(SYNOPSYS_UNCONNECTED_428), .B(
        _f_permutation__round__n2061 ), .Z(_f_permutation__round__c[1428] ) );
  XOR2_X2 _f_permutation__round__U5842  ( .A(SYNOPSYS_UNCONNECTED_237), .B(
        _f_permutation__round__n2062 ), .Z(_f_permutation__round__c[467] ) );
  XOR2_X2 _f_permutation__round__U5841  ( .A(SYNOPSYS_UNCONNECTED_108), .B(
        _f_permutation__round__n2061 ), .Z(_f_permutation__round__c[1364] ) );
  XOR2_X2 _f_permutation__round__U5840  ( .A(_f_permutation__round_in[1171]), 
        .B(_f_permutation__round__n2062 ), .Z(_f_permutation__round__c[403] )
         );
  XOR2_X2 _f_permutation__round__U5839  ( .A(_f_permutation__round_in[1300]), 
        .B(_f_permutation__round__n2061 ), .Z(_f_permutation__round__c[1300] )
         );
  XOR2_X2 _f_permutation__round__U5838  ( .A(_f_permutation__round_in[1491]), 
        .B(_f_permutation__round__n2062 ), .Z(_f_permutation__round__c[339] )
         );
  XOR2_X2 _f_permutation__round__U5837  ( .A(_f_permutation__round__n1637 ), 
        .B(_f_permutation__round__n1636 ), .Z(_f_permutation__round__n2305 )
         );
  XOR2_X2 _f_permutation__round__U5836  ( .A(SYNOPSYS_UNCONNECTED_879), .B(
        _f_permutation__round__n1638 ), .Z(_f_permutation__round__n1636 ) );
  XOR2_X2 _f_permutation__round__U5835  ( .A(SYNOPSYS_UNCONNECTED_239), .B(
        SYNOPSYS_UNCONNECTED_559), .Z(_f_permutation__round__n1637 ) );
  XOR2_X2 _f_permutation__round__U5834  ( .A(_f_permutation__round_in[1489]), 
        .B(_f_permutation__round_in[1169]), .Z(_f_permutation__round__n1638 )
         );
  XOR2_X2 _f_permutation__round__U5833  ( .A(_f_permutation__round__n1640 ), 
        .B(_f_permutation__round__n1639 ), .Z(_f_permutation__round__n2508 )
         );
  XOR2_X2 _f_permutation__round__U5832  ( .A(SYNOPSYS_UNCONNECTED_1070), .B(
        _f_permutation__round__n1641 ), .Z(_f_permutation__round__n1639 ) );
  XOR2_X2 _f_permutation__round__U5831  ( .A(SYNOPSYS_UNCONNECTED_430), .B(
        SYNOPSYS_UNCONNECTED_750), .Z(_f_permutation__round__n1640 ) );
  XOR2_X2 _f_permutation__round__U5830  ( .A(_f_permutation__round_in[1298]), 
        .B(SYNOPSYS_UNCONNECTED_110), .Z(_f_permutation__round__n1641 ) );
  XOR2_X2 _f_permutation__round__U5829  ( .A(_f_permutation__round__n2305 ), 
        .B(_f_permutation__round__n2508 ), .Z(_f_permutation__round__n2306 )
         );
  XOR2_X2 _f_permutation__round__U5828  ( .A(_f_permutation__round_in[1554]), 
        .B(_f_permutation__round__n2306 ), .Z(_f_permutation__round__c[18] )
         );
  XOR2_X2 _f_permutation__round__U5827  ( .A(_f_permutation__round__n1643 ), 
        .B(_f_permutation__round__n1642 ), .Z(_f_permutation__round__n2063 )
         );
  XOR2_X2 _f_permutation__round__U5826  ( .A(SYNOPSYS_UNCONNECTED_814), .B(
        _f_permutation__round__n1644 ), .Z(_f_permutation__round__n1642 ) );
  XOR2_X2 _f_permutation__round__U5825  ( .A(SYNOPSYS_UNCONNECTED_174), .B(
        SYNOPSYS_UNCONNECTED_494), .Z(_f_permutation__round__n1643 ) );
  XOR2_X2 _f_permutation__round__U5824  ( .A(_f_permutation__round_in[1554]), 
        .B(_f_permutation__round_in[1234]), .Z(_f_permutation__round__n1644 )
         );
  XOR2_X2 _f_permutation__round__U5823  ( .A(_f_permutation__round__n1646 ), 
        .B(_f_permutation__round__n1645 ), .Z(_f_permutation__round__n2292 )
         );
  XOR2_X2 _f_permutation__round__U5822  ( .A(SYNOPSYS_UNCONNECTED_1005), .B(
        _f_permutation__round__n1647 ), .Z(_f_permutation__round__n1645 ) );
  XOR2_X2 _f_permutation__round__U5821  ( .A(SYNOPSYS_UNCONNECTED_365), .B(
        SYNOPSYS_UNCONNECTED_685), .Z(_f_permutation__round__n1646 ) );
  XOR2_X2 _f_permutation__round__U5820  ( .A(_f_permutation__round_in[1363]), 
        .B(_f_permutation__round_in[1043]), .Z(_f_permutation__round__n1647 )
         );
  XOR2_X2 _f_permutation__round__U5819  ( .A(_f_permutation__round__n2063 ), 
        .B(_f_permutation__round__n2292 ), .Z(_f_permutation__round__n2064 )
         );
  XOR2_X2 _f_permutation__round__U5818  ( .A(SYNOPSYS_UNCONNECTED_1069), .B(
        _f_permutation__round__n2064 ), .Z(_f_permutation__round__c[1555] ) );
  XOR2_X2 _f_permutation__round__U5817  ( .A(_f_permutation__round__n1649 ), 
        .B(_f_permutation__round__n1648 ), .Z(_f_permutation__round__n2515 )
         );
  XOR2_X2 _f_permutation__round__U5816  ( .A(SYNOPSYS_UNCONNECTED_943), .B(
        _f_permutation__round__n1650 ), .Z(_f_permutation__round__n1648 ) );
  XOR2_X2 _f_permutation__round__U5815  ( .A(SYNOPSYS_UNCONNECTED_303), .B(
        SYNOPSYS_UNCONNECTED_623), .Z(_f_permutation__round__n1649 ) );
  XOR2_X2 _f_permutation__round__U5814  ( .A(_f_permutation__round_in[1425]), 
        .B(_f_permutation__round_in[1105]), .Z(_f_permutation__round__n1650 )
         );
  XOR2_X2 _f_permutation__round__U5813  ( .A(_f_permutation__round__n2063 ), 
        .B(_f_permutation__round__n2515 ), .Z(_f_permutation__round__n2065 )
         );
  XOR2_X2 _f_permutation__round__U5812  ( .A(SYNOPSYS_UNCONNECTED_878), .B(
        _f_permutation__round__n2065 ), .Z(_f_permutation__round__c[594] ) );
  XOR2_X2 _f_permutation__round__U5811  ( .A(SYNOPSYS_UNCONNECTED_749), .B(
        _f_permutation__round__n2064 ), .Z(_f_permutation__round__c[1491] ) );
  XOR2_X2 _f_permutation__round__U5810  ( .A(SYNOPSYS_UNCONNECTED_558), .B(
        _f_permutation__round__n2065 ), .Z(_f_permutation__round__c[530] ) );
  XOR2_X2 _f_permutation__round__U5809  ( .A(SYNOPSYS_UNCONNECTED_429), .B(
        _f_permutation__round__n2064 ), .Z(_f_permutation__round__c[1427] ) );
  XOR2_X2 _f_permutation__round__U5808  ( .A(SYNOPSYS_UNCONNECTED_238), .B(
        _f_permutation__round__n2065 ), .Z(_f_permutation__round__c[466] ) );
  XOR2_X2 _f_permutation__round__U5807  ( .A(SYNOPSYS_UNCONNECTED_109), .B(
        _f_permutation__round__n2064 ), .Z(_f_permutation__round__c[1363] ) );
  XOR2_X2 _f_permutation__round__U5806  ( .A(_f_permutation__round_in[1170]), 
        .B(_f_permutation__round__n2065 ), .Z(_f_permutation__round__c[402] )
         );
  XOR2_X2 _f_permutation__round__U5805  ( .A(_f_permutation__round_in[1299]), 
        .B(_f_permutation__round__n2064 ), .Z(_f_permutation__round__c[1299] )
         );
  XOR2_X2 _f_permutation__round__U5804  ( .A(_f_permutation__round_in[1490]), 
        .B(_f_permutation__round__n2065 ), .Z(_f_permutation__round__c[338] )
         );
  XOR2_X2 _f_permutation__round__U5803  ( .A(_f_permutation__round__n1652 ), 
        .B(_f_permutation__round__n1651 ), .Z(_f_permutation__round__n2309 )
         );
  XOR2_X2 _f_permutation__round__U5802  ( .A(SYNOPSYS_UNCONNECTED_880), .B(
        _f_permutation__round__n1653 ), .Z(_f_permutation__round__n1651 ) );
  XOR2_X2 _f_permutation__round__U5801  ( .A(SYNOPSYS_UNCONNECTED_240), .B(
        SYNOPSYS_UNCONNECTED_560), .Z(_f_permutation__round__n1652 ) );
  XOR2_X2 _f_permutation__round__U5800  ( .A(_f_permutation__round_in[1488]), 
        .B(_f_permutation__round_in[1168]), .Z(_f_permutation__round__n1653 )
         );
  XOR2_X2 _f_permutation__round__U5799  ( .A(_f_permutation__round__n1655 ), 
        .B(_f_permutation__round__n1654 ), .Z(_f_permutation__round__n2511 )
         );
  XOR2_X2 _f_permutation__round__U5798  ( .A(SYNOPSYS_UNCONNECTED_1071), .B(
        _f_permutation__round__n1656 ), .Z(_f_permutation__round__n1654 ) );
  XOR2_X2 _f_permutation__round__U5797  ( .A(SYNOPSYS_UNCONNECTED_431), .B(
        SYNOPSYS_UNCONNECTED_751), .Z(_f_permutation__round__n1655 ) );
  XOR2_X2 _f_permutation__round__U5796  ( .A(_f_permutation__round_in[1297]), 
        .B(SYNOPSYS_UNCONNECTED_111), .Z(_f_permutation__round__n1656 ) );
  XOR2_X2 _f_permutation__round__U5795  ( .A(_f_permutation__round__n2309 ), 
        .B(_f_permutation__round__n2511 ), .Z(_f_permutation__round__n2310 )
         );
  XOR2_X2 _f_permutation__round__U5794  ( .A(_f_permutation__round_in[1553]), 
        .B(_f_permutation__round__n2310 ), .Z(_f_permutation__round__c[17] )
         );
  XOR2_X2 _f_permutation__round__U5793  ( .A(_f_permutation__round__n1658 ), 
        .B(_f_permutation__round__n1657 ), .Z(_f_permutation__round__n2066 )
         );
  XOR2_X2 _f_permutation__round__U5792  ( .A(SYNOPSYS_UNCONNECTED_815), .B(
        _f_permutation__round__n1659 ), .Z(_f_permutation__round__n1657 ) );
  XOR2_X2 _f_permutation__round__U5791  ( .A(SYNOPSYS_UNCONNECTED_175), .B(
        SYNOPSYS_UNCONNECTED_495), .Z(_f_permutation__round__n1658 ) );
  XOR2_X2 _f_permutation__round__U5790  ( .A(_f_permutation__round_in[1553]), 
        .B(_f_permutation__round_in[1233]), .Z(_f_permutation__round__n1659 )
         );
  XOR2_X2 _f_permutation__round__U5789  ( .A(_f_permutation__round__n1661 ), 
        .B(_f_permutation__round__n1660 ), .Z(_f_permutation__round__n2296 )
         );
  XOR2_X2 _f_permutation__round__U5788  ( .A(SYNOPSYS_UNCONNECTED_1006), .B(
        _f_permutation__round__n1662 ), .Z(_f_permutation__round__n1660 ) );
  XOR2_X2 _f_permutation__round__U5787  ( .A(SYNOPSYS_UNCONNECTED_366), .B(
        SYNOPSYS_UNCONNECTED_686), .Z(_f_permutation__round__n1661 ) );
  XOR2_X2 _f_permutation__round__U5786  ( .A(_f_permutation__round_in[1362]), 
        .B(_f_permutation__round_in[1042]), .Z(_f_permutation__round__n1662 )
         );
  XOR2_X2 _f_permutation__round__U5785  ( .A(_f_permutation__round__n2066 ), 
        .B(_f_permutation__round__n2296 ), .Z(_f_permutation__round__n2067 )
         );
  XOR2_X2 _f_permutation__round__U5784  ( .A(SYNOPSYS_UNCONNECTED_1070), .B(
        _f_permutation__round__n2067 ), .Z(_f_permutation__round__c[1554] ) );
  XOR2_X2 _f_permutation__round__U5783  ( .A(_f_permutation__round__n1664 ), 
        .B(_f_permutation__round__n1663 ), .Z(_f_permutation__round__n2518 )
         );
  XOR2_X2 _f_permutation__round__U5782  ( .A(SYNOPSYS_UNCONNECTED_944), .B(
        _f_permutation__round__n1665 ), .Z(_f_permutation__round__n1663 ) );
  XOR2_X2 _f_permutation__round__U5781  ( .A(SYNOPSYS_UNCONNECTED_304), .B(
        SYNOPSYS_UNCONNECTED_624), .Z(_f_permutation__round__n1664 ) );
  XOR2_X2 _f_permutation__round__U5780  ( .A(_f_permutation__round_in[1424]), 
        .B(_f_permutation__round_in[1104]), .Z(_f_permutation__round__n1665 )
         );
  XOR2_X2 _f_permutation__round__U5779  ( .A(_f_permutation__round__n2066 ), 
        .B(_f_permutation__round__n2518 ), .Z(_f_permutation__round__n2068 )
         );
  XOR2_X2 _f_permutation__round__U5778  ( .A(SYNOPSYS_UNCONNECTED_879), .B(
        _f_permutation__round__n2068 ), .Z(_f_permutation__round__c[593] ) );
  XOR2_X2 _f_permutation__round__U5777  ( .A(SYNOPSYS_UNCONNECTED_750), .B(
        _f_permutation__round__n2067 ), .Z(_f_permutation__round__c[1490] ) );
  XOR2_X2 _f_permutation__round__U5776  ( .A(SYNOPSYS_UNCONNECTED_559), .B(
        _f_permutation__round__n2068 ), .Z(_f_permutation__round__c[529] ) );
  XOR2_X2 _f_permutation__round__U5775  ( .A(SYNOPSYS_UNCONNECTED_430), .B(
        _f_permutation__round__n2067 ), .Z(_f_permutation__round__c[1426] ) );
  XOR2_X2 _f_permutation__round__U5774  ( .A(SYNOPSYS_UNCONNECTED_239), .B(
        _f_permutation__round__n2068 ), .Z(_f_permutation__round__c[465] ) );
  XOR2_X2 _f_permutation__round__U5773  ( .A(SYNOPSYS_UNCONNECTED_110), .B(
        _f_permutation__round__n2067 ), .Z(_f_permutation__round__c[1362] ) );
  XOR2_X2 _f_permutation__round__U5772  ( .A(_f_permutation__round_in[1169]), 
        .B(_f_permutation__round__n2068 ), .Z(_f_permutation__round__c[401] )
         );
  XOR2_X2 _f_permutation__round__U5771  ( .A(_f_permutation__round_in[1298]), 
        .B(_f_permutation__round__n2067 ), .Z(_f_permutation__round__c[1298] )
         );
  XOR2_X2 _f_permutation__round__U5770  ( .A(_f_permutation__round_in[1489]), 
        .B(_f_permutation__round__n2068 ), .Z(_f_permutation__round__c[337] )
         );
  XOR2_X2 _f_permutation__round__U5769  ( .A(_f_permutation__round__n1667 ), 
        .B(_f_permutation__round__n1666 ), .Z(_f_permutation__round__n2313 )
         );
  XOR2_X2 _f_permutation__round__U5768  ( .A(SYNOPSYS_UNCONNECTED_881), .B(
        _f_permutation__round__n1668 ), .Z(_f_permutation__round__n1666 ) );
  XOR2_X2 _f_permutation__round__U5767  ( .A(SYNOPSYS_UNCONNECTED_241), .B(
        SYNOPSYS_UNCONNECTED_561), .Z(_f_permutation__round__n1667 ) );
  XOR2_X2 _f_permutation__round__U5766  ( .A(_f_permutation__round_in[1487]), 
        .B(_f_permutation__round_in[1167]), .Z(_f_permutation__round__n1668 )
         );
  XOR2_X2 _f_permutation__round__U5765  ( .A(_f_permutation__round__n1670 ), 
        .B(_f_permutation__round__n1669 ), .Z(_f_permutation__round__n2514 )
         );
  XOR2_X2 _f_permutation__round__U5764  ( .A(SYNOPSYS_UNCONNECTED_1072), .B(
        _f_permutation__round__n1671 ), .Z(_f_permutation__round__n1669 ) );
  XOR2_X2 _f_permutation__round__U5763  ( .A(SYNOPSYS_UNCONNECTED_432), .B(
        SYNOPSYS_UNCONNECTED_752), .Z(_f_permutation__round__n1670 ) );
  XOR2_X2 _f_permutation__round__U5762  ( .A(_f_permutation__round_in[1296]), 
        .B(SYNOPSYS_UNCONNECTED_112), .Z(_f_permutation__round__n1671 ) );
  XOR2_X2 _f_permutation__round__U5761  ( .A(_f_permutation__round__n2313 ), 
        .B(_f_permutation__round__n2514 ), .Z(_f_permutation__round__n2314 )
         );
  XOR2_X2 _f_permutation__round__U5760  ( .A(_f_permutation__round_in[1552]), 
        .B(_f_permutation__round__n2314 ), .Z(_f_permutation__round__c[16] )
         );
  XOR2_X2 _f_permutation__round__U5759  ( .A(_f_permutation__round__n1673 ), 
        .B(_f_permutation__round__n1672 ), .Z(_f_permutation__round__n2069 )
         );
  XOR2_X2 _f_permutation__round__U5758  ( .A(SYNOPSYS_UNCONNECTED_816), .B(
        _f_permutation__round__n1674 ), .Z(_f_permutation__round__n1672 ) );
  XOR2_X2 _f_permutation__round__U5757  ( .A(SYNOPSYS_UNCONNECTED_176), .B(
        SYNOPSYS_UNCONNECTED_496), .Z(_f_permutation__round__n1673 ) );
  XOR2_X2 _f_permutation__round__U5756  ( .A(_f_permutation__round_in[1552]), 
        .B(_f_permutation__round_in[1232]), .Z(_f_permutation__round__n1674 )
         );
  XOR2_X2 _f_permutation__round__U5755  ( .A(_f_permutation__round__n1676 ), 
        .B(_f_permutation__round__n1675 ), .Z(_f_permutation__round__n2300 )
         );
  XOR2_X2 _f_permutation__round__U5754  ( .A(SYNOPSYS_UNCONNECTED_1007), .B(
        _f_permutation__round__n1677 ), .Z(_f_permutation__round__n1675 ) );
  XOR2_X2 _f_permutation__round__U5753  ( .A(SYNOPSYS_UNCONNECTED_367), .B(
        SYNOPSYS_UNCONNECTED_687), .Z(_f_permutation__round__n1676 ) );
  XOR2_X2 _f_permutation__round__U5752  ( .A(_f_permutation__round_in[1361]), 
        .B(_f_permutation__round_in[1041]), .Z(_f_permutation__round__n1677 )
         );
  XOR2_X2 _f_permutation__round__U5751  ( .A(_f_permutation__round__n2069 ), 
        .B(_f_permutation__round__n2300 ), .Z(_f_permutation__round__n2070 )
         );
  XOR2_X2 _f_permutation__round__U5750  ( .A(SYNOPSYS_UNCONNECTED_1071), .B(
        _f_permutation__round__n2070 ), .Z(_f_permutation__round__c[1553] ) );
  XOR2_X2 _f_permutation__round__U5749  ( .A(_f_permutation__round__n1679 ), 
        .B(_f_permutation__round__n1678 ), .Z(_f_permutation__round__n2521 )
         );
  XOR2_X2 _f_permutation__round__U5748  ( .A(SYNOPSYS_UNCONNECTED_945), .B(
        _f_permutation__round__n1680 ), .Z(_f_permutation__round__n1678 ) );
  XOR2_X2 _f_permutation__round__U5747  ( .A(SYNOPSYS_UNCONNECTED_305), .B(
        SYNOPSYS_UNCONNECTED_625), .Z(_f_permutation__round__n1679 ) );
  XOR2_X2 _f_permutation__round__U5746  ( .A(_f_permutation__round_in[1423]), 
        .B(_f_permutation__round_in[1103]), .Z(_f_permutation__round__n1680 )
         );
  XOR2_X2 _f_permutation__round__U5745  ( .A(_f_permutation__round__n2069 ), 
        .B(_f_permutation__round__n2521 ), .Z(_f_permutation__round__n2071 )
         );
  XOR2_X2 _f_permutation__round__U5744  ( .A(SYNOPSYS_UNCONNECTED_880), .B(
        _f_permutation__round__n2071 ), .Z(_f_permutation__round__c[592] ) );
  XOR2_X2 _f_permutation__round__U5743  ( .A(SYNOPSYS_UNCONNECTED_751), .B(
        _f_permutation__round__n2070 ), .Z(_f_permutation__round__c[1489] ) );
  XOR2_X2 _f_permutation__round__U5742  ( .A(SYNOPSYS_UNCONNECTED_560), .B(
        _f_permutation__round__n2071 ), .Z(_f_permutation__round__c[528] ) );
  XOR2_X2 _f_permutation__round__U5741  ( .A(SYNOPSYS_UNCONNECTED_431), .B(
        _f_permutation__round__n2070 ), .Z(_f_permutation__round__c[1425] ) );
  XOR2_X2 _f_permutation__round__U5740  ( .A(SYNOPSYS_UNCONNECTED_240), .B(
        _f_permutation__round__n2071 ), .Z(_f_permutation__round__c[464] ) );
  XOR2_X2 _f_permutation__round__U5739  ( .A(SYNOPSYS_UNCONNECTED_111), .B(
        _f_permutation__round__n2070 ), .Z(_f_permutation__round__c[1361] ) );
  XOR2_X2 _f_permutation__round__U5738  ( .A(_f_permutation__round_in[1168]), 
        .B(_f_permutation__round__n2071 ), .Z(_f_permutation__round__c[400] )
         );
  XOR2_X2 _f_permutation__round__U5737  ( .A(_f_permutation__round_in[1297]), 
        .B(_f_permutation__round__n2070 ), .Z(_f_permutation__round__c[1297] )
         );
  XOR2_X2 _f_permutation__round__U5736  ( .A(_f_permutation__round_in[1488]), 
        .B(_f_permutation__round__n2071 ), .Z(_f_permutation__round__c[336] )
         );
  XOR2_X2 _f_permutation__round__U5735  ( .A(_f_permutation__round__n1682 ), 
        .B(_f_permutation__round__n1681 ), .Z(_f_permutation__round__n2317 )
         );
  XOR2_X2 _f_permutation__round__U5734  ( .A(SYNOPSYS_UNCONNECTED_882), .B(
        _f_permutation__round__n1683 ), .Z(_f_permutation__round__n1681 ) );
  XOR2_X2 _f_permutation__round__U5733  ( .A(SYNOPSYS_UNCONNECTED_242), .B(
        SYNOPSYS_UNCONNECTED_562), .Z(_f_permutation__round__n1682 ) );
  XOR2_X2 _f_permutation__round__U5732  ( .A(_f_permutation__round_in[1486]), 
        .B(_f_permutation__round_in[1166]), .Z(_f_permutation__round__n1683 )
         );
  XOR2_X2 _f_permutation__round__U5731  ( .A(_f_permutation__round__n1685 ), 
        .B(_f_permutation__round__n1684 ), .Z(_f_permutation__round__n2517 )
         );
  XOR2_X2 _f_permutation__round__U5730  ( .A(SYNOPSYS_UNCONNECTED_1073), .B(
        _f_permutation__round__n1686 ), .Z(_f_permutation__round__n1684 ) );
  XOR2_X2 _f_permutation__round__U5729  ( .A(SYNOPSYS_UNCONNECTED_433), .B(
        SYNOPSYS_UNCONNECTED_753), .Z(_f_permutation__round__n1685 ) );
  XOR2_X2 _f_permutation__round__U5728  ( .A(_f_permutation__round_in[1295]), 
        .B(SYNOPSYS_UNCONNECTED_113), .Z(_f_permutation__round__n1686 ) );
  XOR2_X2 _f_permutation__round__U5727  ( .A(_f_permutation__round__n2317 ), 
        .B(_f_permutation__round__n2517 ), .Z(_f_permutation__round__n2318 )
         );
  XOR2_X2 _f_permutation__round__U5726  ( .A(_f_permutation__round_in[1551]), 
        .B(_f_permutation__round__n2318 ), .Z(_f_permutation__round__c[15] )
         );
  XOR2_X2 _f_permutation__round__U5725  ( .A(_f_permutation__round__n1688 ), 
        .B(_f_permutation__round__n1687 ), .Z(_f_permutation__round__n2072 )
         );
  XOR2_X2 _f_permutation__round__U5724  ( .A(SYNOPSYS_UNCONNECTED_817), .B(
        _f_permutation__round__n1689 ), .Z(_f_permutation__round__n1687 ) );
  XOR2_X2 _f_permutation__round__U5723  ( .A(SYNOPSYS_UNCONNECTED_177), .B(
        SYNOPSYS_UNCONNECTED_497), .Z(_f_permutation__round__n1688 ) );
  XOR2_X2 _f_permutation__round__U5722  ( .A(_f_permutation__round_in[1551]), 
        .B(_f_permutation__round_in[1231]), .Z(_f_permutation__round__n1689 )
         );
  XOR2_X2 _f_permutation__round__U5721  ( .A(_f_permutation__round__n1691 ), 
        .B(_f_permutation__round__n1690 ), .Z(_f_permutation__round__n2304 )
         );
  XOR2_X2 _f_permutation__round__U5720  ( .A(SYNOPSYS_UNCONNECTED_1008), .B(
        _f_permutation__round__n1692 ), .Z(_f_permutation__round__n1690 ) );
  XOR2_X2 _f_permutation__round__U5719  ( .A(SYNOPSYS_UNCONNECTED_368), .B(
        SYNOPSYS_UNCONNECTED_688), .Z(_f_permutation__round__n1691 ) );
  XOR2_X2 _f_permutation__round__U5718  ( .A(_f_permutation__round_in[1360]), 
        .B(_f_permutation__round_in[1040]), .Z(_f_permutation__round__n1692 )
         );
  XOR2_X2 _f_permutation__round__U5717  ( .A(_f_permutation__round__n2072 ), 
        .B(_f_permutation__round__n2304 ), .Z(_f_permutation__round__n2073 )
         );
  XOR2_X2 _f_permutation__round__U5716  ( .A(SYNOPSYS_UNCONNECTED_1072), .B(
        _f_permutation__round__n2073 ), .Z(_f_permutation__round__c[1552] ) );
  XOR2_X2 _f_permutation__round__U5715  ( .A(_f_permutation__round__n1694 ), 
        .B(_f_permutation__round__n1693 ), .Z(_f_permutation__round__n2524 )
         );
  XOR2_X2 _f_permutation__round__U5714  ( .A(SYNOPSYS_UNCONNECTED_946), .B(
        _f_permutation__round__n1695 ), .Z(_f_permutation__round__n1693 ) );
  XOR2_X2 _f_permutation__round__U5713  ( .A(SYNOPSYS_UNCONNECTED_306), .B(
        SYNOPSYS_UNCONNECTED_626), .Z(_f_permutation__round__n1694 ) );
  XOR2_X2 _f_permutation__round__U5712  ( .A(_f_permutation__round_in[1422]), 
        .B(_f_permutation__round_in[1102]), .Z(_f_permutation__round__n1695 )
         );
  XOR2_X2 _f_permutation__round__U5711  ( .A(_f_permutation__round__n2072 ), 
        .B(_f_permutation__round__n2524 ), .Z(_f_permutation__round__n2074 )
         );
  XOR2_X2 _f_permutation__round__U5710  ( .A(SYNOPSYS_UNCONNECTED_881), .B(
        _f_permutation__round__n2074 ), .Z(_f_permutation__round__c[591] ) );
  XOR2_X2 _f_permutation__round__U5709  ( .A(SYNOPSYS_UNCONNECTED_752), .B(
        _f_permutation__round__n2073 ), .Z(_f_permutation__round__c[1488] ) );
  XOR2_X2 _f_permutation__round__U5708  ( .A(SYNOPSYS_UNCONNECTED_561), .B(
        _f_permutation__round__n2074 ), .Z(_f_permutation__round__c[527] ) );
  XOR2_X2 _f_permutation__round__U5707  ( .A(SYNOPSYS_UNCONNECTED_432), .B(
        _f_permutation__round__n2073 ), .Z(_f_permutation__round__c[1424] ) );
  XOR2_X2 _f_permutation__round__U5706  ( .A(SYNOPSYS_UNCONNECTED_241), .B(
        _f_permutation__round__n2074 ), .Z(_f_permutation__round__c[463] ) );
  XOR2_X2 _f_permutation__round__U5705  ( .A(SYNOPSYS_UNCONNECTED_112), .B(
        _f_permutation__round__n2073 ), .Z(_f_permutation__round__c[1360] ) );
  XOR2_X2 _f_permutation__round__U5704  ( .A(_f_permutation__round_in[1167]), 
        .B(_f_permutation__round__n2074 ), .Z(_f_permutation__round__c[399] )
         );
  XOR2_X2 _f_permutation__round__U5703  ( .A(_f_permutation__round_in[1296]), 
        .B(_f_permutation__round__n2073 ), .Z(_f_permutation__round__c[1296] )
         );
  XOR2_X2 _f_permutation__round__U5702  ( .A(_f_permutation__round_in[1487]), 
        .B(_f_permutation__round__n2074 ), .Z(_f_permutation__round__c[335] )
         );
  XOR2_X2 _f_permutation__round__U5701  ( .A(_f_permutation__round__n1697 ), 
        .B(_f_permutation__round__n1696 ), .Z(_f_permutation__round__n2321 )
         );
  XOR2_X2 _f_permutation__round__U5700  ( .A(SYNOPSYS_UNCONNECTED_883), .B(
        _f_permutation__round__n1698 ), .Z(_f_permutation__round__n1696 ) );
  XOR2_X2 _f_permutation__round__U5699  ( .A(SYNOPSYS_UNCONNECTED_243), .B(
        SYNOPSYS_UNCONNECTED_563), .Z(_f_permutation__round__n1697 ) );
  XOR2_X2 _f_permutation__round__U5698  ( .A(_f_permutation__round_in[1485]), 
        .B(_f_permutation__round_in[1165]), .Z(_f_permutation__round__n1698 )
         );
  XOR2_X2 _f_permutation__round__U5697  ( .A(_f_permutation__round__n1700 ), 
        .B(_f_permutation__round__n1699 ), .Z(_f_permutation__round__n2520 )
         );
  XOR2_X2 _f_permutation__round__U5696  ( .A(SYNOPSYS_UNCONNECTED_1074), .B(
        _f_permutation__round__n1701 ), .Z(_f_permutation__round__n1699 ) );
  XOR2_X2 _f_permutation__round__U5695  ( .A(SYNOPSYS_UNCONNECTED_434), .B(
        SYNOPSYS_UNCONNECTED_754), .Z(_f_permutation__round__n1700 ) );
  XOR2_X2 _f_permutation__round__U5694  ( .A(_f_permutation__round_in[1294]), 
        .B(SYNOPSYS_UNCONNECTED_114), .Z(_f_permutation__round__n1701 ) );
  XOR2_X2 _f_permutation__round__U5693  ( .A(_f_permutation__round__n2321 ), 
        .B(_f_permutation__round__n2520 ), .Z(_f_permutation__round__n2322 )
         );
  XOR2_X2 _f_permutation__round__U5692  ( .A(_f_permutation__round_in[1550]), 
        .B(_f_permutation__round__n2322 ), .Z(_f_permutation__round__c[14] )
         );
  XOR2_X2 _f_permutation__round__U5691  ( .A(_f_permutation__round__n1703 ), 
        .B(_f_permutation__round__n1702 ), .Z(_f_permutation__round__n2075 )
         );
  XOR2_X2 _f_permutation__round__U5690  ( .A(SYNOPSYS_UNCONNECTED_818), .B(
        _f_permutation__round__n1704 ), .Z(_f_permutation__round__n1702 ) );
  XOR2_X2 _f_permutation__round__U5689  ( .A(SYNOPSYS_UNCONNECTED_178), .B(
        SYNOPSYS_UNCONNECTED_498), .Z(_f_permutation__round__n1703 ) );
  XOR2_X2 _f_permutation__round__U5688  ( .A(_f_permutation__round_in[1550]), 
        .B(_f_permutation__round_in[1230]), .Z(_f_permutation__round__n1704 )
         );
  XOR2_X2 _f_permutation__round__U5687  ( .A(_f_permutation__round__n1706 ), 
        .B(_f_permutation__round__n1705 ), .Z(_f_permutation__round__n2308 )
         );
  XOR2_X2 _f_permutation__round__U5686  ( .A(SYNOPSYS_UNCONNECTED_1009), .B(
        _f_permutation__round__n1707 ), .Z(_f_permutation__round__n1705 ) );
  XOR2_X2 _f_permutation__round__U5685  ( .A(SYNOPSYS_UNCONNECTED_369), .B(
        SYNOPSYS_UNCONNECTED_689), .Z(_f_permutation__round__n1706 ) );
  XOR2_X2 _f_permutation__round__U5684  ( .A(_f_permutation__round_in[1359]), 
        .B(_f_permutation__round_in[1039]), .Z(_f_permutation__round__n1707 )
         );
  XOR2_X2 _f_permutation__round__U5683  ( .A(_f_permutation__round__n2075 ), 
        .B(_f_permutation__round__n2308 ), .Z(_f_permutation__round__n2076 )
         );
  XOR2_X2 _f_permutation__round__U5682  ( .A(SYNOPSYS_UNCONNECTED_1073), .B(
        _f_permutation__round__n2076 ), .Z(_f_permutation__round__c[1551] ) );
  XOR2_X2 _f_permutation__round__U5681  ( .A(_f_permutation__round__n1709 ), 
        .B(_f_permutation__round__n1708 ), .Z(_f_permutation__round__n2527 )
         );
  XOR2_X2 _f_permutation__round__U5680  ( .A(SYNOPSYS_UNCONNECTED_947), .B(
        _f_permutation__round__n1710 ), .Z(_f_permutation__round__n1708 ) );
  XOR2_X2 _f_permutation__round__U5679  ( .A(SYNOPSYS_UNCONNECTED_307), .B(
        SYNOPSYS_UNCONNECTED_627), .Z(_f_permutation__round__n1709 ) );
  XOR2_X2 _f_permutation__round__U5678  ( .A(_f_permutation__round_in[1421]), 
        .B(_f_permutation__round_in[1101]), .Z(_f_permutation__round__n1710 )
         );
  XOR2_X2 _f_permutation__round__U5677  ( .A(_f_permutation__round__n2075 ), 
        .B(_f_permutation__round__n2527 ), .Z(_f_permutation__round__n2077 )
         );
  XOR2_X2 _f_permutation__round__U5676  ( .A(SYNOPSYS_UNCONNECTED_882), .B(
        _f_permutation__round__n2077 ), .Z(_f_permutation__round__c[590] ) );
  XOR2_X2 _f_permutation__round__U5675  ( .A(SYNOPSYS_UNCONNECTED_753), .B(
        _f_permutation__round__n2076 ), .Z(_f_permutation__round__c[1487] ) );
  XOR2_X2 _f_permutation__round__U5674  ( .A(SYNOPSYS_UNCONNECTED_562), .B(
        _f_permutation__round__n2077 ), .Z(_f_permutation__round__c[526] ) );
  XOR2_X2 _f_permutation__round__U5673  ( .A(SYNOPSYS_UNCONNECTED_433), .B(
        _f_permutation__round__n2076 ), .Z(_f_permutation__round__c[1423] ) );
  XOR2_X2 _f_permutation__round__U5672  ( .A(SYNOPSYS_UNCONNECTED_242), .B(
        _f_permutation__round__n2077 ), .Z(_f_permutation__round__c[462] ) );
  XOR2_X2 _f_permutation__round__U5671  ( .A(SYNOPSYS_UNCONNECTED_113), .B(
        _f_permutation__round__n2076 ), .Z(_f_permutation__round__c[1359] ) );
  XOR2_X2 _f_permutation__round__U5670  ( .A(_f_permutation__round_in[1166]), 
        .B(_f_permutation__round__n2077 ), .Z(_f_permutation__round__c[398] )
         );
  XOR2_X2 _f_permutation__round__U5669  ( .A(_f_permutation__round_in[1295]), 
        .B(_f_permutation__round__n2076 ), .Z(_f_permutation__round__c[1295] )
         );
  XOR2_X2 _f_permutation__round__U5668  ( .A(_f_permutation__round_in[1486]), 
        .B(_f_permutation__round__n2077 ), .Z(_f_permutation__round__c[334] )
         );
  XOR2_X2 _f_permutation__round__U5667  ( .A(_f_permutation__round__n1712 ), 
        .B(_f_permutation__round__n1711 ), .Z(_f_permutation__round__n2325 )
         );
  XOR2_X2 _f_permutation__round__U5666  ( .A(SYNOPSYS_UNCONNECTED_884), .B(
        _f_permutation__round__n1713 ), .Z(_f_permutation__round__n1711 ) );
  XOR2_X2 _f_permutation__round__U5665  ( .A(SYNOPSYS_UNCONNECTED_244), .B(
        SYNOPSYS_UNCONNECTED_564), .Z(_f_permutation__round__n1712 ) );
  XOR2_X2 _f_permutation__round__U5664  ( .A(_f_permutation__round_in[1484]), 
        .B(_f_permutation__round_in[1164]), .Z(_f_permutation__round__n1713 )
         );
  XOR2_X2 _f_permutation__round__U5663  ( .A(_f_permutation__round__n1715 ), 
        .B(_f_permutation__round__n1714 ), .Z(_f_permutation__round__n2523 )
         );
  XOR2_X2 _f_permutation__round__U5662  ( .A(SYNOPSYS_UNCONNECTED_1075), .B(
        _f_permutation__round__n1716 ), .Z(_f_permutation__round__n1714 ) );
  XOR2_X2 _f_permutation__round__U5661  ( .A(SYNOPSYS_UNCONNECTED_435), .B(
        SYNOPSYS_UNCONNECTED_755), .Z(_f_permutation__round__n1715 ) );
  XOR2_X2 _f_permutation__round__U5660  ( .A(_f_permutation__round_in[1293]), 
        .B(SYNOPSYS_UNCONNECTED_115), .Z(_f_permutation__round__n1716 ) );
  XOR2_X2 _f_permutation__round__U5659  ( .A(_f_permutation__round__n2325 ), 
        .B(_f_permutation__round__n2523 ), .Z(_f_permutation__round__n2326 )
         );
  XOR2_X2 _f_permutation__round__U5658  ( .A(_f_permutation__round_in[1549]), 
        .B(_f_permutation__round__n2326 ), .Z(_f_permutation__round__c[13] )
         );
  XOR2_X2 _f_permutation__round__U5657  ( .A(_f_permutation__round__n1718 ), 
        .B(_f_permutation__round__n1717 ), .Z(_f_permutation__round__n2078 )
         );
  XOR2_X2 _f_permutation__round__U5656  ( .A(SYNOPSYS_UNCONNECTED_819), .B(
        _f_permutation__round__n1719 ), .Z(_f_permutation__round__n1717 ) );
  XOR2_X2 _f_permutation__round__U5655  ( .A(SYNOPSYS_UNCONNECTED_179), .B(
        SYNOPSYS_UNCONNECTED_499), .Z(_f_permutation__round__n1718 ) );
  XOR2_X2 _f_permutation__round__U5654  ( .A(_f_permutation__round_in[1549]), 
        .B(_f_permutation__round_in[1229]), .Z(_f_permutation__round__n1719 )
         );
  XOR2_X2 _f_permutation__round__U5653  ( .A(_f_permutation__round__n1721 ), 
        .B(_f_permutation__round__n1720 ), .Z(_f_permutation__round__n2312 )
         );
  XOR2_X2 _f_permutation__round__U5652  ( .A(SYNOPSYS_UNCONNECTED_1010), .B(
        _f_permutation__round__n1722 ), .Z(_f_permutation__round__n1720 ) );
  XOR2_X2 _f_permutation__round__U5651  ( .A(SYNOPSYS_UNCONNECTED_370), .B(
        SYNOPSYS_UNCONNECTED_690), .Z(_f_permutation__round__n1721 ) );
  XOR2_X2 _f_permutation__round__U5650  ( .A(_f_permutation__round_in[1358]), 
        .B(_f_permutation__round_in[1038]), .Z(_f_permutation__round__n1722 )
         );
  XOR2_X2 _f_permutation__round__U5649  ( .A(_f_permutation__round__n2078 ), 
        .B(_f_permutation__round__n2312 ), .Z(_f_permutation__round__n2079 )
         );
  XOR2_X2 _f_permutation__round__U5648  ( .A(SYNOPSYS_UNCONNECTED_1074), .B(
        _f_permutation__round__n2079 ), .Z(_f_permutation__round__c[1550] ) );
  XOR2_X2 _f_permutation__round__U5647  ( .A(_f_permutation__round__n1724 ), 
        .B(_f_permutation__round__n1723 ), .Z(_f_permutation__round__n2530 )
         );
  XOR2_X2 _f_permutation__round__U5646  ( .A(SYNOPSYS_UNCONNECTED_948), .B(
        _f_permutation__round__n1725 ), .Z(_f_permutation__round__n1723 ) );
  XOR2_X2 _f_permutation__round__U5645  ( .A(SYNOPSYS_UNCONNECTED_308), .B(
        SYNOPSYS_UNCONNECTED_628), .Z(_f_permutation__round__n1724 ) );
  XOR2_X2 _f_permutation__round__U5644  ( .A(_f_permutation__round_in[1420]), 
        .B(_f_permutation__round_in[1100]), .Z(_f_permutation__round__n1725 )
         );
  XOR2_X2 _f_permutation__round__U5643  ( .A(_f_permutation__round__n2078 ), 
        .B(_f_permutation__round__n2530 ), .Z(_f_permutation__round__n2080 )
         );
  XOR2_X2 _f_permutation__round__U5642  ( .A(SYNOPSYS_UNCONNECTED_883), .B(
        _f_permutation__round__n2080 ), .Z(_f_permutation__round__c[589] ) );
  XOR2_X2 _f_permutation__round__U5641  ( .A(SYNOPSYS_UNCONNECTED_754), .B(
        _f_permutation__round__n2079 ), .Z(_f_permutation__round__c[1486] ) );
  XOR2_X2 _f_permutation__round__U5640  ( .A(SYNOPSYS_UNCONNECTED_563), .B(
        _f_permutation__round__n2080 ), .Z(_f_permutation__round__c[525] ) );
  XOR2_X2 _f_permutation__round__U5639  ( .A(SYNOPSYS_UNCONNECTED_434), .B(
        _f_permutation__round__n2079 ), .Z(_f_permutation__round__c[1422] ) );
  XOR2_X2 _f_permutation__round__U5638  ( .A(SYNOPSYS_UNCONNECTED_243), .B(
        _f_permutation__round__n2080 ), .Z(_f_permutation__round__c[461] ) );
  XOR2_X2 _f_permutation__round__U5637  ( .A(SYNOPSYS_UNCONNECTED_114), .B(
        _f_permutation__round__n2079 ), .Z(_f_permutation__round__c[1358] ) );
  XOR2_X2 _f_permutation__round__U5636  ( .A(_f_permutation__round_in[1165]), 
        .B(_f_permutation__round__n2080 ), .Z(_f_permutation__round__c[397] )
         );
  XOR2_X2 _f_permutation__round__U5635  ( .A(_f_permutation__round_in[1294]), 
        .B(_f_permutation__round__n2079 ), .Z(_f_permutation__round__c[1294] )
         );
  XOR2_X2 _f_permutation__round__U5634  ( .A(_f_permutation__round_in[1485]), 
        .B(_f_permutation__round__n2080 ), .Z(_f_permutation__round__c[333] )
         );
  XOR2_X2 _f_permutation__round__U5633  ( .A(_f_permutation__round__n1727 ), 
        .B(_f_permutation__round__n1726 ), .Z(_f_permutation__round__n2329 )
         );
  XOR2_X2 _f_permutation__round__U5632  ( .A(SYNOPSYS_UNCONNECTED_885), .B(
        _f_permutation__round__n1728 ), .Z(_f_permutation__round__n1726 ) );
  XOR2_X2 _f_permutation__round__U5631  ( .A(SYNOPSYS_UNCONNECTED_245), .B(
        SYNOPSYS_UNCONNECTED_565), .Z(_f_permutation__round__n1727 ) );
  XOR2_X2 _f_permutation__round__U5630  ( .A(_f_permutation__round_in[1483]), 
        .B(_f_permutation__round_in[1163]), .Z(_f_permutation__round__n1728 )
         );
  XOR2_X2 _f_permutation__round__U5629  ( .A(_f_permutation__round__n1730 ), 
        .B(_f_permutation__round__n1729 ), .Z(_f_permutation__round__n2526 )
         );
  XOR2_X2 _f_permutation__round__U5628  ( .A(SYNOPSYS_UNCONNECTED_1076), .B(
        _f_permutation__round__n1731 ), .Z(_f_permutation__round__n1729 ) );
  XOR2_X2 _f_permutation__round__U5627  ( .A(SYNOPSYS_UNCONNECTED_436), .B(
        SYNOPSYS_UNCONNECTED_756), .Z(_f_permutation__round__n1730 ) );
  XOR2_X2 _f_permutation__round__U5626  ( .A(_f_permutation__round_in[1292]), 
        .B(SYNOPSYS_UNCONNECTED_116), .Z(_f_permutation__round__n1731 ) );
  XOR2_X2 _f_permutation__round__U5625  ( .A(_f_permutation__round__n2329 ), 
        .B(_f_permutation__round__n2526 ), .Z(_f_permutation__round__n2330 )
         );
  XOR2_X2 _f_permutation__round__U5624  ( .A(_f_permutation__round_in[1548]), 
        .B(_f_permutation__round__n2330 ), .Z(_f_permutation__round__c[12] )
         );
  XOR2_X2 _f_permutation__round__U5623  ( .A(_f_permutation__round__n1733 ), 
        .B(_f_permutation__round__n1732 ), .Z(_f_permutation__round__n2081 )
         );
  XOR2_X2 _f_permutation__round__U5622  ( .A(SYNOPSYS_UNCONNECTED_820), .B(
        _f_permutation__round__n1734 ), .Z(_f_permutation__round__n1732 ) );
  XOR2_X2 _f_permutation__round__U5621  ( .A(SYNOPSYS_UNCONNECTED_180), .B(
        SYNOPSYS_UNCONNECTED_500), .Z(_f_permutation__round__n1733 ) );
  XOR2_X2 _f_permutation__round__U5620  ( .A(_f_permutation__round_in[1548]), 
        .B(_f_permutation__round_in[1228]), .Z(_f_permutation__round__n1734 )
         );
  XOR2_X2 _f_permutation__round__U5619  ( .A(_f_permutation__round__n1736 ), 
        .B(_f_permutation__round__n1735 ), .Z(_f_permutation__round__n2316 )
         );
  XOR2_X2 _f_permutation__round__U5618  ( .A(SYNOPSYS_UNCONNECTED_1011), .B(
        _f_permutation__round__n1737 ), .Z(_f_permutation__round__n1735 ) );
  XOR2_X2 _f_permutation__round__U5617  ( .A(SYNOPSYS_UNCONNECTED_371), .B(
        SYNOPSYS_UNCONNECTED_691), .Z(_f_permutation__round__n1736 ) );
  XOR2_X2 _f_permutation__round__U5616  ( .A(_f_permutation__round_in[1357]), 
        .B(_f_permutation__round_in[1037]), .Z(_f_permutation__round__n1737 )
         );
  XOR2_X2 _f_permutation__round__U5615  ( .A(_f_permutation__round__n2081 ), 
        .B(_f_permutation__round__n2316 ), .Z(_f_permutation__round__n2082 )
         );
  XOR2_X2 _f_permutation__round__U5614  ( .A(SYNOPSYS_UNCONNECTED_1075), .B(
        _f_permutation__round__n2082 ), .Z(_f_permutation__round__c[1549] ) );
  XOR2_X2 _f_permutation__round__U5613  ( .A(_f_permutation__round__n1739 ), 
        .B(_f_permutation__round__n1738 ), .Z(_f_permutation__round__n2533 )
         );
  XOR2_X2 _f_permutation__round__U5612  ( .A(SYNOPSYS_UNCONNECTED_949), .B(
        _f_permutation__round__n1740 ), .Z(_f_permutation__round__n1738 ) );
  XOR2_X2 _f_permutation__round__U5611  ( .A(SYNOPSYS_UNCONNECTED_309), .B(
        SYNOPSYS_UNCONNECTED_629), .Z(_f_permutation__round__n1739 ) );
  XOR2_X2 _f_permutation__round__U5610  ( .A(_f_permutation__round_in[1419]), 
        .B(_f_permutation__round_in[1099]), .Z(_f_permutation__round__n1740 )
         );
  XOR2_X2 _f_permutation__round__U5609  ( .A(_f_permutation__round__n2081 ), 
        .B(_f_permutation__round__n2533 ), .Z(_f_permutation__round__n2083 )
         );
  XOR2_X2 _f_permutation__round__U5608  ( .A(SYNOPSYS_UNCONNECTED_884), .B(
        _f_permutation__round__n2083 ), .Z(_f_permutation__round__c[588] ) );
  XOR2_X2 _f_permutation__round__U5607  ( .A(SYNOPSYS_UNCONNECTED_755), .B(
        _f_permutation__round__n2082 ), .Z(_f_permutation__round__c[1485] ) );
  XOR2_X2 _f_permutation__round__U5606  ( .A(SYNOPSYS_UNCONNECTED_564), .B(
        _f_permutation__round__n2083 ), .Z(_f_permutation__round__c[524] ) );
  XOR2_X2 _f_permutation__round__U5605  ( .A(SYNOPSYS_UNCONNECTED_435), .B(
        _f_permutation__round__n2082 ), .Z(_f_permutation__round__c[1421] ) );
  XOR2_X2 _f_permutation__round__U5604  ( .A(SYNOPSYS_UNCONNECTED_244), .B(
        _f_permutation__round__n2083 ), .Z(_f_permutation__round__c[460] ) );
  XOR2_X2 _f_permutation__round__U5603  ( .A(SYNOPSYS_UNCONNECTED_115), .B(
        _f_permutation__round__n2082 ), .Z(_f_permutation__round__c[1357] ) );
  XOR2_X2 _f_permutation__round__U5602  ( .A(_f_permutation__round_in[1164]), 
        .B(_f_permutation__round__n2083 ), .Z(_f_permutation__round__c[396] )
         );
  XOR2_X2 _f_permutation__round__U5601  ( .A(_f_permutation__round_in[1293]), 
        .B(_f_permutation__round__n2082 ), .Z(_f_permutation__round__c[1293] )
         );
  XOR2_X2 _f_permutation__round__U5600  ( .A(_f_permutation__round_in[1484]), 
        .B(_f_permutation__round__n2083 ), .Z(_f_permutation__round__c[332] )
         );
  XOR2_X2 _f_permutation__round__U5599  ( .A(_f_permutation__round__n1742 ), 
        .B(_f_permutation__round__n1741 ), .Z(_f_permutation__round__n2333 )
         );
  XOR2_X2 _f_permutation__round__U5598  ( .A(SYNOPSYS_UNCONNECTED_886), .B(
        _f_permutation__round__n1743 ), .Z(_f_permutation__round__n1741 ) );
  XOR2_X2 _f_permutation__round__U5597  ( .A(SYNOPSYS_UNCONNECTED_246), .B(
        SYNOPSYS_UNCONNECTED_566), .Z(_f_permutation__round__n1742 ) );
  XOR2_X2 _f_permutation__round__U5596  ( .A(_f_permutation__round_in[1482]), 
        .B(_f_permutation__round_in[1162]), .Z(_f_permutation__round__n1743 )
         );
  XOR2_X2 _f_permutation__round__U5595  ( .A(_f_permutation__round__n1745 ), 
        .B(_f_permutation__round__n1744 ), .Z(_f_permutation__round__n2529 )
         );
  XOR2_X2 _f_permutation__round__U5594  ( .A(SYNOPSYS_UNCONNECTED_1077), .B(
        _f_permutation__round__n1746 ), .Z(_f_permutation__round__n1744 ) );
  XOR2_X2 _f_permutation__round__U5593  ( .A(SYNOPSYS_UNCONNECTED_437), .B(
        SYNOPSYS_UNCONNECTED_757), .Z(_f_permutation__round__n1745 ) );
  XOR2_X2 _f_permutation__round__U5592  ( .A(_f_permutation__round_in[1291]), 
        .B(SYNOPSYS_UNCONNECTED_117), .Z(_f_permutation__round__n1746 ) );
  XOR2_X2 _f_permutation__round__U5591  ( .A(_f_permutation__round__n2333 ), 
        .B(_f_permutation__round__n2529 ), .Z(_f_permutation__round__n2334 )
         );
  XOR2_X2 _f_permutation__round__U5590  ( .A(_f_permutation__round_in[1547]), 
        .B(_f_permutation__round__n2334 ), .Z(_f_permutation__round__c[11] )
         );
  XOR2_X2 _f_permutation__round__U5589  ( .A(_f_permutation__round__n1748 ), 
        .B(_f_permutation__round__n1747 ), .Z(_f_permutation__round__n2084 )
         );
  XOR2_X2 _f_permutation__round__U5588  ( .A(SYNOPSYS_UNCONNECTED_821), .B(
        _f_permutation__round__n1749 ), .Z(_f_permutation__round__n1747 ) );
  XOR2_X2 _f_permutation__round__U5587  ( .A(SYNOPSYS_UNCONNECTED_181), .B(
        SYNOPSYS_UNCONNECTED_501), .Z(_f_permutation__round__n1748 ) );
  XOR2_X2 _f_permutation__round__U5586  ( .A(_f_permutation__round_in[1547]), 
        .B(_f_permutation__round_in[1227]), .Z(_f_permutation__round__n1749 )
         );
  XOR2_X2 _f_permutation__round__U5585  ( .A(_f_permutation__round__n1751 ), 
        .B(_f_permutation__round__n1750 ), .Z(_f_permutation__round__n2320 )
         );
  XOR2_X2 _f_permutation__round__U5584  ( .A(SYNOPSYS_UNCONNECTED_1012), .B(
        _f_permutation__round__n1752 ), .Z(_f_permutation__round__n1750 ) );
  XOR2_X2 _f_permutation__round__U5583  ( .A(SYNOPSYS_UNCONNECTED_372), .B(
        SYNOPSYS_UNCONNECTED_692), .Z(_f_permutation__round__n1751 ) );
  XOR2_X2 _f_permutation__round__U5582  ( .A(_f_permutation__round_in[1356]), 
        .B(_f_permutation__round_in[1036]), .Z(_f_permutation__round__n1752 )
         );
  XOR2_X2 _f_permutation__round__U5581  ( .A(_f_permutation__round__n2084 ), 
        .B(_f_permutation__round__n2320 ), .Z(_f_permutation__round__n2085 )
         );
  XOR2_X2 _f_permutation__round__U5580  ( .A(SYNOPSYS_UNCONNECTED_1076), .B(
        _f_permutation__round__n2085 ), .Z(_f_permutation__round__c[1548] ) );
  XOR2_X2 _f_permutation__round__U5579  ( .A(_f_permutation__round__n1754 ), 
        .B(_f_permutation__round__n1753 ), .Z(_f_permutation__round__n2536 )
         );
  XOR2_X2 _f_permutation__round__U5578  ( .A(SYNOPSYS_UNCONNECTED_950), .B(
        _f_permutation__round__n1755 ), .Z(_f_permutation__round__n1753 ) );
  XOR2_X2 _f_permutation__round__U5577  ( .A(SYNOPSYS_UNCONNECTED_310), .B(
        SYNOPSYS_UNCONNECTED_630), .Z(_f_permutation__round__n1754 ) );
  XOR2_X2 _f_permutation__round__U5576  ( .A(_f_permutation__round_in[1418]), 
        .B(_f_permutation__round_in[1098]), .Z(_f_permutation__round__n1755 )
         );
  XOR2_X2 _f_permutation__round__U5575  ( .A(_f_permutation__round__n2084 ), 
        .B(_f_permutation__round__n2536 ), .Z(_f_permutation__round__n2086 )
         );
  XOR2_X2 _f_permutation__round__U5574  ( .A(SYNOPSYS_UNCONNECTED_885), .B(
        _f_permutation__round__n2086 ), .Z(_f_permutation__round__c[587] ) );
  XOR2_X2 _f_permutation__round__U5573  ( .A(SYNOPSYS_UNCONNECTED_756), .B(
        _f_permutation__round__n2085 ), .Z(_f_permutation__round__c[1484] ) );
  XOR2_X2 _f_permutation__round__U5572  ( .A(SYNOPSYS_UNCONNECTED_565), .B(
        _f_permutation__round__n2086 ), .Z(_f_permutation__round__c[523] ) );
  XOR2_X2 _f_permutation__round__U5571  ( .A(SYNOPSYS_UNCONNECTED_436), .B(
        _f_permutation__round__n2085 ), .Z(_f_permutation__round__c[1420] ) );
  XOR2_X2 _f_permutation__round__U5570  ( .A(SYNOPSYS_UNCONNECTED_245), .B(
        _f_permutation__round__n2086 ), .Z(_f_permutation__round__c[459] ) );
  XOR2_X2 _f_permutation__round__U5569  ( .A(SYNOPSYS_UNCONNECTED_116), .B(
        _f_permutation__round__n2085 ), .Z(_f_permutation__round__c[1356] ) );
  XOR2_X2 _f_permutation__round__U5568  ( .A(_f_permutation__round_in[1163]), 
        .B(_f_permutation__round__n2086 ), .Z(_f_permutation__round__c[395] )
         );
  XOR2_X2 _f_permutation__round__U5567  ( .A(_f_permutation__round_in[1292]), 
        .B(_f_permutation__round__n2085 ), .Z(_f_permutation__round__c[1292] )
         );
  XOR2_X2 _f_permutation__round__U5566  ( .A(_f_permutation__round_in[1483]), 
        .B(_f_permutation__round__n2086 ), .Z(_f_permutation__round__c[331] )
         );
  XOR2_X2 _f_permutation__round__U5565  ( .A(_f_permutation__round__n1757 ), 
        .B(_f_permutation__round__n1756 ), .Z(_f_permutation__round__n2337 )
         );
  XOR2_X2 _f_permutation__round__U5564  ( .A(SYNOPSYS_UNCONNECTED_887), .B(
        _f_permutation__round__n1758 ), .Z(_f_permutation__round__n1756 ) );
  XOR2_X2 _f_permutation__round__U5563  ( .A(SYNOPSYS_UNCONNECTED_247), .B(
        SYNOPSYS_UNCONNECTED_567), .Z(_f_permutation__round__n1757 ) );
  XOR2_X2 _f_permutation__round__U5562  ( .A(_f_permutation__round_in[1481]), 
        .B(_f_permutation__round_in[1161]), .Z(_f_permutation__round__n1758 )
         );
  XOR2_X2 _f_permutation__round__U5561  ( .A(_f_permutation__round__n1760 ), 
        .B(_f_permutation__round__n1759 ), .Z(_f_permutation__round__n2532 )
         );
  XOR2_X2 _f_permutation__round__U5560  ( .A(SYNOPSYS_UNCONNECTED_1078), .B(
        _f_permutation__round__n1761 ), .Z(_f_permutation__round__n1759 ) );
  XOR2_X2 _f_permutation__round__U5559  ( .A(SYNOPSYS_UNCONNECTED_438), .B(
        SYNOPSYS_UNCONNECTED_758), .Z(_f_permutation__round__n1760 ) );
  XOR2_X2 _f_permutation__round__U5558  ( .A(_f_permutation__round_in[1290]), 
        .B(SYNOPSYS_UNCONNECTED_118), .Z(_f_permutation__round__n1761 ) );
  XOR2_X2 _f_permutation__round__U5557  ( .A(_f_permutation__round__n2337 ), 
        .B(_f_permutation__round__n2532 ), .Z(_f_permutation__round__n2338 )
         );
  XOR2_X2 _f_permutation__round__U5556  ( .A(_f_permutation__round_in[1546]), 
        .B(_f_permutation__round__n2338 ), .Z(_f_permutation__round__c[10] )
         );
  XOR2_X2 _f_permutation__round__U5555  ( .A(_f_permutation__round__n1763 ), 
        .B(_f_permutation__round__n1762 ), .Z(_f_permutation__round__n2087 )
         );
  XOR2_X2 _f_permutation__round__U5554  ( .A(SYNOPSYS_UNCONNECTED_822), .B(
        _f_permutation__round__n1764 ), .Z(_f_permutation__round__n1762 ) );
  XOR2_X2 _f_permutation__round__U5553  ( .A(SYNOPSYS_UNCONNECTED_182), .B(
        SYNOPSYS_UNCONNECTED_502), .Z(_f_permutation__round__n1763 ) );
  XOR2_X2 _f_permutation__round__U5552  ( .A(_f_permutation__round_in[1546]), 
        .B(_f_permutation__round_in[1226]), .Z(_f_permutation__round__n1764 )
         );
  XOR2_X2 _f_permutation__round__U5551  ( .A(_f_permutation__round__n1766 ), 
        .B(_f_permutation__round__n1765 ), .Z(_f_permutation__round__n2324 )
         );
  XOR2_X2 _f_permutation__round__U5550  ( .A(SYNOPSYS_UNCONNECTED_1013), .B(
        _f_permutation__round__n1767 ), .Z(_f_permutation__round__n1765 ) );
  XOR2_X2 _f_permutation__round__U5549  ( .A(SYNOPSYS_UNCONNECTED_373), .B(
        SYNOPSYS_UNCONNECTED_693), .Z(_f_permutation__round__n1766 ) );
  XOR2_X2 _f_permutation__round__U5548  ( .A(_f_permutation__round_in[1355]), 
        .B(_f_permutation__round_in[1035]), .Z(_f_permutation__round__n1767 )
         );
  XOR2_X2 _f_permutation__round__U5547  ( .A(_f_permutation__round__n2087 ), 
        .B(_f_permutation__round__n2324 ), .Z(_f_permutation__round__n2088 )
         );
  XOR2_X2 _f_permutation__round__U5546  ( .A(SYNOPSYS_UNCONNECTED_1077), .B(
        _f_permutation__round__n2088 ), .Z(_f_permutation__round__c[1547] ) );
  XOR2_X2 _f_permutation__round__U5545  ( .A(_f_permutation__round__n1769 ), 
        .B(_f_permutation__round__n1768 ), .Z(_f_permutation__round__n2539 )
         );
  XOR2_X2 _f_permutation__round__U5544  ( .A(SYNOPSYS_UNCONNECTED_951), .B(
        _f_permutation__round__n1770 ), .Z(_f_permutation__round__n1768 ) );
  XOR2_X2 _f_permutation__round__U5543  ( .A(SYNOPSYS_UNCONNECTED_311), .B(
        SYNOPSYS_UNCONNECTED_631), .Z(_f_permutation__round__n1769 ) );
  XOR2_X2 _f_permutation__round__U5542  ( .A(_f_permutation__round_in[1417]), 
        .B(_f_permutation__round_in[1097]), .Z(_f_permutation__round__n1770 )
         );
  XOR2_X2 _f_permutation__round__U5541  ( .A(_f_permutation__round__n2087 ), 
        .B(_f_permutation__round__n2539 ), .Z(_f_permutation__round__n2089 )
         );
  XOR2_X2 _f_permutation__round__U5540  ( .A(SYNOPSYS_UNCONNECTED_886), .B(
        _f_permutation__round__n2089 ), .Z(_f_permutation__round__c[586] ) );
  XOR2_X2 _f_permutation__round__U5539  ( .A(SYNOPSYS_UNCONNECTED_757), .B(
        _f_permutation__round__n2088 ), .Z(_f_permutation__round__c[1483] ) );
  XOR2_X2 _f_permutation__round__U5538  ( .A(SYNOPSYS_UNCONNECTED_566), .B(
        _f_permutation__round__n2089 ), .Z(_f_permutation__round__c[522] ) );
  XOR2_X2 _f_permutation__round__U5537  ( .A(SYNOPSYS_UNCONNECTED_437), .B(
        _f_permutation__round__n2088 ), .Z(_f_permutation__round__c[1419] ) );
  XOR2_X2 _f_permutation__round__U5536  ( .A(SYNOPSYS_UNCONNECTED_246), .B(
        _f_permutation__round__n2089 ), .Z(_f_permutation__round__c[458] ) );
  XOR2_X2 _f_permutation__round__U5535  ( .A(SYNOPSYS_UNCONNECTED_117), .B(
        _f_permutation__round__n2088 ), .Z(_f_permutation__round__c[1355] ) );
  XOR2_X2 _f_permutation__round__U5534  ( .A(_f_permutation__round_in[1162]), 
        .B(_f_permutation__round__n2089 ), .Z(_f_permutation__round__c[394] )
         );
  XOR2_X2 _f_permutation__round__U5533  ( .A(_f_permutation__round_in[1291]), 
        .B(_f_permutation__round__n2088 ), .Z(_f_permutation__round__c[1291] )
         );
  XOR2_X2 _f_permutation__round__U5532  ( .A(_f_permutation__round_in[1482]), 
        .B(_f_permutation__round__n2089 ), .Z(_f_permutation__round__c[330] )
         );
  XOR2_X2 _f_permutation__round__U5531  ( .A(_f_permutation__round__n1772 ), 
        .B(_f_permutation__round__n1771 ), .Z(_f_permutation__round__n2341 )
         );
  XOR2_X2 _f_permutation__round__U5530  ( .A(SYNOPSYS_UNCONNECTED_888), .B(
        _f_permutation__round__n1773 ), .Z(_f_permutation__round__n1771 ) );
  XOR2_X2 _f_permutation__round__U5529  ( .A(SYNOPSYS_UNCONNECTED_248), .B(
        SYNOPSYS_UNCONNECTED_568), .Z(_f_permutation__round__n1772 ) );
  XOR2_X2 _f_permutation__round__U5528  ( .A(_f_permutation__round_in[1480]), 
        .B(_f_permutation__round_in[1160]), .Z(_f_permutation__round__n1773 )
         );
  XOR2_X2 _f_permutation__round__U5527  ( .A(_f_permutation__round__n1775 ), 
        .B(_f_permutation__round__n1774 ), .Z(_f_permutation__round__n2535 )
         );
  XOR2_X2 _f_permutation__round__U5526  ( .A(SYNOPSYS_UNCONNECTED_1079), .B(
        _f_permutation__round__n1776 ), .Z(_f_permutation__round__n1774 ) );
  XOR2_X2 _f_permutation__round__U5525  ( .A(SYNOPSYS_UNCONNECTED_439), .B(
        SYNOPSYS_UNCONNECTED_759), .Z(_f_permutation__round__n1775 ) );
  XOR2_X2 _f_permutation__round__U5524  ( .A(_f_permutation__round_in[1289]), 
        .B(SYNOPSYS_UNCONNECTED_119), .Z(_f_permutation__round__n1776 ) );
  XOR2_X2 _f_permutation__round__U5523  ( .A(_f_permutation__round__n2341 ), 
        .B(_f_permutation__round__n2535 ), .Z(_f_permutation__round__n2342 )
         );
  XOR2_X2 _f_permutation__round__U5522  ( .A(_f_permutation__round_in[1545]), 
        .B(_f_permutation__round__n2342 ), .Z(_f_permutation__round__c[9] ) );
  XOR2_X2 _f_permutation__round__U5521  ( .A(_f_permutation__round__n1778 ), 
        .B(_f_permutation__round__n1777 ), .Z(_f_permutation__round__n2090 )
         );
  XOR2_X2 _f_permutation__round__U5520  ( .A(SYNOPSYS_UNCONNECTED_823), .B(
        _f_permutation__round__n1779 ), .Z(_f_permutation__round__n1777 ) );
  XOR2_X2 _f_permutation__round__U5519  ( .A(SYNOPSYS_UNCONNECTED_183), .B(
        SYNOPSYS_UNCONNECTED_503), .Z(_f_permutation__round__n1778 ) );
  XOR2_X2 _f_permutation__round__U5518  ( .A(_f_permutation__round_in[1545]), 
        .B(_f_permutation__round_in[1225]), .Z(_f_permutation__round__n1779 )
         );
  XOR2_X2 _f_permutation__round__U5517  ( .A(_f_permutation__round__n1781 ), 
        .B(_f_permutation__round__n1780 ), .Z(_f_permutation__round__n2328 )
         );
  XOR2_X2 _f_permutation__round__U5516  ( .A(SYNOPSYS_UNCONNECTED_1014), .B(
        _f_permutation__round__n1782 ), .Z(_f_permutation__round__n1780 ) );
  XOR2_X2 _f_permutation__round__U5515  ( .A(SYNOPSYS_UNCONNECTED_374), .B(
        SYNOPSYS_UNCONNECTED_694), .Z(_f_permutation__round__n1781 ) );
  XOR2_X2 _f_permutation__round__U5514  ( .A(_f_permutation__round_in[1354]), 
        .B(_f_permutation__round_in[1034]), .Z(_f_permutation__round__n1782 )
         );
  XOR2_X2 _f_permutation__round__U5513  ( .A(_f_permutation__round__n2090 ), 
        .B(_f_permutation__round__n2328 ), .Z(_f_permutation__round__n2091 )
         );
  XOR2_X2 _f_permutation__round__U5512  ( .A(SYNOPSYS_UNCONNECTED_1078), .B(
        _f_permutation__round__n2091 ), .Z(_f_permutation__round__c[1546] ) );
  XOR2_X2 _f_permutation__round__U5511  ( .A(_f_permutation__round__n1784 ), 
        .B(_f_permutation__round__n1783 ), .Z(_f_permutation__round__n2542 )
         );
  XOR2_X2 _f_permutation__round__U5510  ( .A(SYNOPSYS_UNCONNECTED_952), .B(
        _f_permutation__round__n1785 ), .Z(_f_permutation__round__n1783 ) );
  XOR2_X2 _f_permutation__round__U5509  ( .A(SYNOPSYS_UNCONNECTED_312), .B(
        SYNOPSYS_UNCONNECTED_632), .Z(_f_permutation__round__n1784 ) );
  XOR2_X2 _f_permutation__round__U5508  ( .A(_f_permutation__round_in[1416]), 
        .B(_f_permutation__round_in[1096]), .Z(_f_permutation__round__n1785 )
         );
  XOR2_X2 _f_permutation__round__U5507  ( .A(_f_permutation__round__n2090 ), 
        .B(_f_permutation__round__n2542 ), .Z(_f_permutation__round__n2092 )
         );
  XOR2_X2 _f_permutation__round__U5506  ( .A(SYNOPSYS_UNCONNECTED_887), .B(
        _f_permutation__round__n2092 ), .Z(_f_permutation__round__c[585] ) );
  XOR2_X2 _f_permutation__round__U5505  ( .A(SYNOPSYS_UNCONNECTED_758), .B(
        _f_permutation__round__n2091 ), .Z(_f_permutation__round__c[1482] ) );
  XOR2_X2 _f_permutation__round__U5504  ( .A(SYNOPSYS_UNCONNECTED_567), .B(
        _f_permutation__round__n2092 ), .Z(_f_permutation__round__c[521] ) );
  XOR2_X2 _f_permutation__round__U5503  ( .A(SYNOPSYS_UNCONNECTED_438), .B(
        _f_permutation__round__n2091 ), .Z(_f_permutation__round__c[1418] ) );
  XOR2_X2 _f_permutation__round__U5502  ( .A(SYNOPSYS_UNCONNECTED_247), .B(
        _f_permutation__round__n2092 ), .Z(_f_permutation__round__c[457] ) );
  XOR2_X2 _f_permutation__round__U5501  ( .A(SYNOPSYS_UNCONNECTED_118), .B(
        _f_permutation__round__n2091 ), .Z(_f_permutation__round__c[1354] ) );
  XOR2_X2 _f_permutation__round__U5500  ( .A(_f_permutation__round_in[1161]), 
        .B(_f_permutation__round__n2092 ), .Z(_f_permutation__round__c[393] )
         );
  XOR2_X2 _f_permutation__round__U5499  ( .A(_f_permutation__round_in[1290]), 
        .B(_f_permutation__round__n2091 ), .Z(_f_permutation__round__c[1290] )
         );
  XOR2_X2 _f_permutation__round__U5498  ( .A(_f_permutation__round_in[1481]), 
        .B(_f_permutation__round__n2092 ), .Z(_f_permutation__round__c[329] )
         );
  XOR2_X2 _f_permutation__round__U5497  ( .A(_f_permutation__round__n1787 ), 
        .B(_f_permutation__round__n1786 ), .Z(_f_permutation__round__n2345 )
         );
  XOR2_X2 _f_permutation__round__U5496  ( .A(SYNOPSYS_UNCONNECTED_889), .B(
        _f_permutation__round__n1788 ), .Z(_f_permutation__round__n1786 ) );
  XOR2_X2 _f_permutation__round__U5495  ( .A(SYNOPSYS_UNCONNECTED_249), .B(
        SYNOPSYS_UNCONNECTED_569), .Z(_f_permutation__round__n1787 ) );
  XOR2_X2 _f_permutation__round__U5494  ( .A(_f_permutation__round_in[1479]), 
        .B(_f_permutation__round_in[1159]), .Z(_f_permutation__round__n1788 )
         );
  XOR2_X2 _f_permutation__round__U5493  ( .A(_f_permutation__round__n1790 ), 
        .B(_f_permutation__round__n1789 ), .Z(_f_permutation__round__n2538 )
         );
  XOR2_X2 _f_permutation__round__U5492  ( .A(SYNOPSYS_UNCONNECTED_1080), .B(
        _f_permutation__round__n1791 ), .Z(_f_permutation__round__n1789 ) );
  XOR2_X2 _f_permutation__round__U5491  ( .A(SYNOPSYS_UNCONNECTED_440), .B(
        SYNOPSYS_UNCONNECTED_760), .Z(_f_permutation__round__n1790 ) );
  XOR2_X2 _f_permutation__round__U5490  ( .A(_f_permutation__round_in[1288]), 
        .B(SYNOPSYS_UNCONNECTED_120), .Z(_f_permutation__round__n1791 ) );
  XOR2_X2 _f_permutation__round__U5489  ( .A(_f_permutation__round__n2345 ), 
        .B(_f_permutation__round__n2538 ), .Z(_f_permutation__round__n2346 )
         );
  XOR2_X2 _f_permutation__round__U5488  ( .A(_f_permutation__round_in[1544]), 
        .B(_f_permutation__round__n2346 ), .Z(_f_permutation__round__c[8] ) );
  XOR2_X2 _f_permutation__round__U5487  ( .A(_f_permutation__round__n1793 ), 
        .B(_f_permutation__round__n1792 ), .Z(_f_permutation__round__n2093 )
         );
  XOR2_X2 _f_permutation__round__U5486  ( .A(SYNOPSYS_UNCONNECTED_824), .B(
        _f_permutation__round__n1794 ), .Z(_f_permutation__round__n1792 ) );
  XOR2_X2 _f_permutation__round__U5485  ( .A(SYNOPSYS_UNCONNECTED_184), .B(
        SYNOPSYS_UNCONNECTED_504), .Z(_f_permutation__round__n1793 ) );
  XOR2_X2 _f_permutation__round__U5484  ( .A(_f_permutation__round_in[1544]), 
        .B(_f_permutation__round_in[1224]), .Z(_f_permutation__round__n1794 )
         );
  XOR2_X2 _f_permutation__round__U5483  ( .A(_f_permutation__round__n1796 ), 
        .B(_f_permutation__round__n1795 ), .Z(_f_permutation__round__n2332 )
         );
  XOR2_X2 _f_permutation__round__U5482  ( .A(SYNOPSYS_UNCONNECTED_1015), .B(
        _f_permutation__round__n1797 ), .Z(_f_permutation__round__n1795 ) );
  XOR2_X2 _f_permutation__round__U5481  ( .A(SYNOPSYS_UNCONNECTED_375), .B(
        SYNOPSYS_UNCONNECTED_695), .Z(_f_permutation__round__n1796 ) );
  XOR2_X2 _f_permutation__round__U5480  ( .A(_f_permutation__round_in[1353]), 
        .B(_f_permutation__round_in[1033]), .Z(_f_permutation__round__n1797 )
         );
  XOR2_X2 _f_permutation__round__U5479  ( .A(_f_permutation__round__n2093 ), 
        .B(_f_permutation__round__n2332 ), .Z(_f_permutation__round__n2094 )
         );
  XOR2_X2 _f_permutation__round__U5478  ( .A(SYNOPSYS_UNCONNECTED_1079), .B(
        _f_permutation__round__n2094 ), .Z(_f_permutation__round__c[1545] ) );
  XOR2_X2 _f_permutation__round__U5477  ( .A(_f_permutation__round__n1799 ), 
        .B(_f_permutation__round__n1798 ), .Z(_f_permutation__round__n2545 )
         );
  XOR2_X2 _f_permutation__round__U5476  ( .A(SYNOPSYS_UNCONNECTED_953), .B(
        _f_permutation__round__n1800 ), .Z(_f_permutation__round__n1798 ) );
  XOR2_X2 _f_permutation__round__U5475  ( .A(SYNOPSYS_UNCONNECTED_313), .B(
        SYNOPSYS_UNCONNECTED_633), .Z(_f_permutation__round__n1799 ) );
  XOR2_X2 _f_permutation__round__U5474  ( .A(_f_permutation__round_in[1415]), 
        .B(_f_permutation__round_in[1095]), .Z(_f_permutation__round__n1800 )
         );
  XOR2_X2 _f_permutation__round__U5473  ( .A(_f_permutation__round__n2093 ), 
        .B(_f_permutation__round__n2545 ), .Z(_f_permutation__round__n2095 )
         );
  XOR2_X2 _f_permutation__round__U5472  ( .A(SYNOPSYS_UNCONNECTED_888), .B(
        _f_permutation__round__n2095 ), .Z(_f_permutation__round__c[584] ) );
  XOR2_X2 _f_permutation__round__U5471  ( .A(SYNOPSYS_UNCONNECTED_759), .B(
        _f_permutation__round__n2094 ), .Z(_f_permutation__round__c[1481] ) );
  XOR2_X2 _f_permutation__round__U5470  ( .A(SYNOPSYS_UNCONNECTED_568), .B(
        _f_permutation__round__n2095 ), .Z(_f_permutation__round__c[520] ) );
  XOR2_X2 _f_permutation__round__U5469  ( .A(SYNOPSYS_UNCONNECTED_439), .B(
        _f_permutation__round__n2094 ), .Z(_f_permutation__round__c[1417] ) );
  XOR2_X2 _f_permutation__round__U5468  ( .A(SYNOPSYS_UNCONNECTED_248), .B(
        _f_permutation__round__n2095 ), .Z(_f_permutation__round__c[456] ) );
  XOR2_X2 _f_permutation__round__U5467  ( .A(SYNOPSYS_UNCONNECTED_119), .B(
        _f_permutation__round__n2094 ), .Z(_f_permutation__round__c[1353] ) );
  XOR2_X2 _f_permutation__round__U5466  ( .A(_f_permutation__round_in[1160]), 
        .B(_f_permutation__round__n2095 ), .Z(_f_permutation__round__c[392] )
         );
  XOR2_X2 _f_permutation__round__U5465  ( .A(_f_permutation__round_in[1289]), 
        .B(_f_permutation__round__n2094 ), .Z(_f_permutation__round__c[1289] )
         );
  XOR2_X2 _f_permutation__round__U5464  ( .A(_f_permutation__round_in[1480]), 
        .B(_f_permutation__round__n2095 ), .Z(_f_permutation__round__c[328] )
         );
  XOR2_X2 _f_permutation__round__U5463  ( .A(_f_permutation__round__n1802 ), 
        .B(_f_permutation__round__n1801 ), .Z(_f_permutation__round__n2349 )
         );
  XOR2_X2 _f_permutation__round__U5462  ( .A(SYNOPSYS_UNCONNECTED_890), .B(
        _f_permutation__round__n1803 ), .Z(_f_permutation__round__n1801 ) );
  XOR2_X2 _f_permutation__round__U5461  ( .A(SYNOPSYS_UNCONNECTED_250), .B(
        SYNOPSYS_UNCONNECTED_570), .Z(_f_permutation__round__n1802 ) );
  XOR2_X2 _f_permutation__round__U5460  ( .A(_f_permutation__round_in[1478]), 
        .B(_f_permutation__round_in[1158]), .Z(_f_permutation__round__n1803 )
         );
  XOR2_X2 _f_permutation__round__U5459  ( .A(_f_permutation__round__n1805 ), 
        .B(_f_permutation__round__n1804 ), .Z(_f_permutation__round__n2541 )
         );
  XOR2_X2 _f_permutation__round__U5458  ( .A(SYNOPSYS_UNCONNECTED_1081), .B(
        _f_permutation__round__n1806 ), .Z(_f_permutation__round__n1804 ) );
  XOR2_X2 _f_permutation__round__U5457  ( .A(SYNOPSYS_UNCONNECTED_441), .B(
        SYNOPSYS_UNCONNECTED_761), .Z(_f_permutation__round__n1805 ) );
  XOR2_X2 _f_permutation__round__U5456  ( .A(_f_permutation__round_in[1287]), 
        .B(SYNOPSYS_UNCONNECTED_121), .Z(_f_permutation__round__n1806 ) );
  XOR2_X2 _f_permutation__round__U5455  ( .A(_f_permutation__round__n2349 ), 
        .B(_f_permutation__round__n2541 ), .Z(_f_permutation__round__n2350 )
         );
  XOR2_X2 _f_permutation__round__U5454  ( .A(_f_permutation__round_in[1543]), 
        .B(_f_permutation__round__n2350 ), .Z(_f_permutation__round__c[7] ) );
  XOR2_X2 _f_permutation__round__U5453  ( .A(_f_permutation__round__n1808 ), 
        .B(_f_permutation__round__n1807 ), .Z(_f_permutation__round__n2096 )
         );
  XOR2_X2 _f_permutation__round__U5452  ( .A(SYNOPSYS_UNCONNECTED_825), .B(
        _f_permutation__round__n1809 ), .Z(_f_permutation__round__n1807 ) );
  XOR2_X2 _f_permutation__round__U5451  ( .A(SYNOPSYS_UNCONNECTED_185), .B(
        SYNOPSYS_UNCONNECTED_505), .Z(_f_permutation__round__n1808 ) );
  XOR2_X2 _f_permutation__round__U5450  ( .A(_f_permutation__round_in[1543]), 
        .B(_f_permutation__round_in[1223]), .Z(_f_permutation__round__n1809 )
         );
  XOR2_X2 _f_permutation__round__U5449  ( .A(_f_permutation__round__n1811 ), 
        .B(_f_permutation__round__n1810 ), .Z(_f_permutation__round__n2336 )
         );
  XOR2_X2 _f_permutation__round__U5448  ( .A(SYNOPSYS_UNCONNECTED_1016), .B(
        _f_permutation__round__n1812 ), .Z(_f_permutation__round__n1810 ) );
  XOR2_X2 _f_permutation__round__U5447  ( .A(SYNOPSYS_UNCONNECTED_376), .B(
        SYNOPSYS_UNCONNECTED_696), .Z(_f_permutation__round__n1811 ) );
  XOR2_X2 _f_permutation__round__U5446  ( .A(_f_permutation__round_in[1352]), 
        .B(_f_permutation__round_in[1032]), .Z(_f_permutation__round__n1812 )
         );
  XOR2_X2 _f_permutation__round__U5445  ( .A(_f_permutation__round__n2096 ), 
        .B(_f_permutation__round__n2336 ), .Z(_f_permutation__round__n2097 )
         );
  XOR2_X2 _f_permutation__round__U5444  ( .A(SYNOPSYS_UNCONNECTED_1080), .B(
        _f_permutation__round__n2097 ), .Z(_f_permutation__round__c[1544] ) );
  XOR2_X2 _f_permutation__round__U5443  ( .A(_f_permutation__round__n1814 ), 
        .B(_f_permutation__round__n1813 ), .Z(_f_permutation__round__n2548 )
         );
  XOR2_X2 _f_permutation__round__U5442  ( .A(SYNOPSYS_UNCONNECTED_954), .B(
        _f_permutation__round__n1815 ), .Z(_f_permutation__round__n1813 ) );
  XOR2_X2 _f_permutation__round__U5441  ( .A(SYNOPSYS_UNCONNECTED_314), .B(
        SYNOPSYS_UNCONNECTED_634), .Z(_f_permutation__round__n1814 ) );
  XOR2_X2 _f_permutation__round__U5440  ( .A(_f_permutation__round_in[1414]), 
        .B(_f_permutation__round_in[1094]), .Z(_f_permutation__round__n1815 )
         );
  XOR2_X2 _f_permutation__round__U5439  ( .A(_f_permutation__round__n2096 ), 
        .B(_f_permutation__round__n2548 ), .Z(_f_permutation__round__n2098 )
         );
  XOR2_X2 _f_permutation__round__U5438  ( .A(SYNOPSYS_UNCONNECTED_889), .B(
        _f_permutation__round__n2098 ), .Z(_f_permutation__round__c[583] ) );
  XOR2_X2 _f_permutation__round__U5437  ( .A(SYNOPSYS_UNCONNECTED_760), .B(
        _f_permutation__round__n2097 ), .Z(_f_permutation__round__c[1480] ) );
  XOR2_X2 _f_permutation__round__U5436  ( .A(SYNOPSYS_UNCONNECTED_569), .B(
        _f_permutation__round__n2098 ), .Z(_f_permutation__round__c[519] ) );
  XOR2_X2 _f_permutation__round__U5435  ( .A(SYNOPSYS_UNCONNECTED_440), .B(
        _f_permutation__round__n2097 ), .Z(_f_permutation__round__c[1416] ) );
  XOR2_X2 _f_permutation__round__U5434  ( .A(SYNOPSYS_UNCONNECTED_249), .B(
        _f_permutation__round__n2098 ), .Z(_f_permutation__round__c[455] ) );
  XOR2_X2 _f_permutation__round__U5433  ( .A(SYNOPSYS_UNCONNECTED_120), .B(
        _f_permutation__round__n2097 ), .Z(_f_permutation__round__c[1352] ) );
  XOR2_X2 _f_permutation__round__U5432  ( .A(_f_permutation__round_in[1159]), 
        .B(_f_permutation__round__n2098 ), .Z(_f_permutation__round__c[391] )
         );
  XOR2_X2 _f_permutation__round__U5431  ( .A(_f_permutation__round_in[1288]), 
        .B(_f_permutation__round__n2097 ), .Z(_f_permutation__round__c[1288] )
         );
  XOR2_X2 _f_permutation__round__U5430  ( .A(_f_permutation__round_in[1479]), 
        .B(_f_permutation__round__n2098 ), .Z(_f_permutation__round__c[327] )
         );
  XOR2_X2 _f_permutation__round__U5429  ( .A(_f_permutation__round__n1817 ), 
        .B(_f_permutation__round__n1816 ), .Z(_f_permutation__round__n2353 )
         );
  XOR2_X2 _f_permutation__round__U5428  ( .A(SYNOPSYS_UNCONNECTED_891), .B(
        _f_permutation__round__n1818 ), .Z(_f_permutation__round__n1816 ) );
  XOR2_X2 _f_permutation__round__U5427  ( .A(SYNOPSYS_UNCONNECTED_251), .B(
        SYNOPSYS_UNCONNECTED_571), .Z(_f_permutation__round__n1817 ) );
  XOR2_X2 _f_permutation__round__U5426  ( .A(_f_permutation__round_in[1477]), 
        .B(_f_permutation__round_in[1157]), .Z(_f_permutation__round__n1818 )
         );
  XOR2_X2 _f_permutation__round__U5425  ( .A(_f_permutation__round__n1820 ), 
        .B(_f_permutation__round__n1819 ), .Z(_f_permutation__round__n2544 )
         );
  XOR2_X2 _f_permutation__round__U5424  ( .A(SYNOPSYS_UNCONNECTED_1082), .B(
        _f_permutation__round__n1821 ), .Z(_f_permutation__round__n1819 ) );
  XOR2_X2 _f_permutation__round__U5423  ( .A(SYNOPSYS_UNCONNECTED_442), .B(
        SYNOPSYS_UNCONNECTED_762), .Z(_f_permutation__round__n1820 ) );
  XOR2_X2 _f_permutation__round__U5422  ( .A(_f_permutation__round_in[1286]), 
        .B(SYNOPSYS_UNCONNECTED_122), .Z(_f_permutation__round__n1821 ) );
  XOR2_X2 _f_permutation__round__U5421  ( .A(_f_permutation__round__n2353 ), 
        .B(_f_permutation__round__n2544 ), .Z(_f_permutation__round__n2354 )
         );
  XOR2_X2 _f_permutation__round__U5420  ( .A(_f_permutation__round_in[1542]), 
        .B(_f_permutation__round__n2354 ), .Z(_f_permutation__round__c[6] ) );
  XOR2_X2 _f_permutation__round__U5419  ( .A(_f_permutation__round__n1823 ), 
        .B(_f_permutation__round__n1822 ), .Z(_f_permutation__round__n2099 )
         );
  XOR2_X2 _f_permutation__round__U5418  ( .A(SYNOPSYS_UNCONNECTED_826), .B(
        _f_permutation__round__n1824 ), .Z(_f_permutation__round__n1822 ) );
  XOR2_X2 _f_permutation__round__U5417  ( .A(SYNOPSYS_UNCONNECTED_186), .B(
        SYNOPSYS_UNCONNECTED_506), .Z(_f_permutation__round__n1823 ) );
  XOR2_X2 _f_permutation__round__U5416  ( .A(_f_permutation__round_in[1542]), 
        .B(_f_permutation__round_in[1222]), .Z(_f_permutation__round__n1824 )
         );
  XOR2_X2 _f_permutation__round__U5415  ( .A(_f_permutation__round__n1826 ), 
        .B(_f_permutation__round__n1825 ), .Z(_f_permutation__round__n2340 )
         );
  XOR2_X2 _f_permutation__round__U5414  ( .A(SYNOPSYS_UNCONNECTED_1017), .B(
        _f_permutation__round__n1827 ), .Z(_f_permutation__round__n1825 ) );
  XOR2_X2 _f_permutation__round__U5413  ( .A(SYNOPSYS_UNCONNECTED_377), .B(
        SYNOPSYS_UNCONNECTED_697), .Z(_f_permutation__round__n1826 ) );
  XOR2_X2 _f_permutation__round__U5412  ( .A(_f_permutation__round_in[1351]), 
        .B(_f_permutation__round_in[1031]), .Z(_f_permutation__round__n1827 )
         );
  XOR2_X2 _f_permutation__round__U5411  ( .A(_f_permutation__round__n2099 ), 
        .B(_f_permutation__round__n2340 ), .Z(_f_permutation__round__n2100 )
         );
  XOR2_X2 _f_permutation__round__U5410  ( .A(SYNOPSYS_UNCONNECTED_1081), .B(
        _f_permutation__round__n2100 ), .Z(_f_permutation__round__c[1543] ) );
  XOR2_X2 _f_permutation__round__U5409  ( .A(_f_permutation__round__n1829 ), 
        .B(_f_permutation__round__n1828 ), .Z(_f_permutation__round__n2551 )
         );
  XOR2_X2 _f_permutation__round__U5408  ( .A(SYNOPSYS_UNCONNECTED_955), .B(
        _f_permutation__round__n1830 ), .Z(_f_permutation__round__n1828 ) );
  XOR2_X2 _f_permutation__round__U5407  ( .A(SYNOPSYS_UNCONNECTED_315), .B(
        SYNOPSYS_UNCONNECTED_635), .Z(_f_permutation__round__n1829 ) );
  XOR2_X2 _f_permutation__round__U5406  ( .A(_f_permutation__round_in[1413]), 
        .B(_f_permutation__round_in[1093]), .Z(_f_permutation__round__n1830 )
         );
  XOR2_X2 _f_permutation__round__U5405  ( .A(_f_permutation__round__n2099 ), 
        .B(_f_permutation__round__n2551 ), .Z(_f_permutation__round__n2101 )
         );
  XOR2_X2 _f_permutation__round__U5404  ( .A(SYNOPSYS_UNCONNECTED_890), .B(
        _f_permutation__round__n2101 ), .Z(_f_permutation__round__c[582] ) );
  XOR2_X2 _f_permutation__round__U5403  ( .A(SYNOPSYS_UNCONNECTED_761), .B(
        _f_permutation__round__n2100 ), .Z(_f_permutation__round__c[1479] ) );
  XOR2_X2 _f_permutation__round__U5402  ( .A(SYNOPSYS_UNCONNECTED_570), .B(
        _f_permutation__round__n2101 ), .Z(_f_permutation__round__c[518] ) );
  XOR2_X2 _f_permutation__round__U5401  ( .A(SYNOPSYS_UNCONNECTED_441), .B(
        _f_permutation__round__n2100 ), .Z(_f_permutation__round__c[1415] ) );
  XOR2_X2 _f_permutation__round__U5400  ( .A(SYNOPSYS_UNCONNECTED_250), .B(
        _f_permutation__round__n2101 ), .Z(_f_permutation__round__c[454] ) );
  XOR2_X2 _f_permutation__round__U5399  ( .A(SYNOPSYS_UNCONNECTED_121), .B(
        _f_permutation__round__n2100 ), .Z(_f_permutation__round__c[1351] ) );
  XOR2_X2 _f_permutation__round__U5398  ( .A(_f_permutation__round_in[1158]), 
        .B(_f_permutation__round__n2101 ), .Z(_f_permutation__round__c[390] )
         );
  XOR2_X2 _f_permutation__round__U5397  ( .A(_f_permutation__round_in[1287]), 
        .B(_f_permutation__round__n2100 ), .Z(_f_permutation__round__c[1287] )
         );
  XOR2_X2 _f_permutation__round__U5396  ( .A(_f_permutation__round_in[1478]), 
        .B(_f_permutation__round__n2101 ), .Z(_f_permutation__round__c[326] )
         );
  XOR2_X2 _f_permutation__round__U5395  ( .A(_f_permutation__round__n1832 ), 
        .B(_f_permutation__round__n1831 ), .Z(_f_permutation__round__n2357 )
         );
  XOR2_X2 _f_permutation__round__U5394  ( .A(SYNOPSYS_UNCONNECTED_892), .B(
        _f_permutation__round__n1833 ), .Z(_f_permutation__round__n1831 ) );
  XOR2_X2 _f_permutation__round__U5393  ( .A(SYNOPSYS_UNCONNECTED_252), .B(
        SYNOPSYS_UNCONNECTED_572), .Z(_f_permutation__round__n1832 ) );
  XOR2_X2 _f_permutation__round__U5392  ( .A(_f_permutation__round_in[1476]), 
        .B(_f_permutation__round_in[1156]), .Z(_f_permutation__round__n1833 )
         );
  XOR2_X2 _f_permutation__round__U5391  ( .A(_f_permutation__round__n1835 ), 
        .B(_f_permutation__round__n1834 ), .Z(_f_permutation__round__n2547 )
         );
  XOR2_X2 _f_permutation__round__U5390  ( .A(SYNOPSYS_UNCONNECTED_1083), .B(
        _f_permutation__round__n1836 ), .Z(_f_permutation__round__n1834 ) );
  XOR2_X2 _f_permutation__round__U5389  ( .A(SYNOPSYS_UNCONNECTED_443), .B(
        SYNOPSYS_UNCONNECTED_763), .Z(_f_permutation__round__n1835 ) );
  XOR2_X2 _f_permutation__round__U5388  ( .A(_f_permutation__round_in[1285]), 
        .B(SYNOPSYS_UNCONNECTED_123), .Z(_f_permutation__round__n1836 ) );
  XOR2_X2 _f_permutation__round__U5387  ( .A(_f_permutation__round__n2357 ), 
        .B(_f_permutation__round__n2547 ), .Z(_f_permutation__round__n2358 )
         );
  XOR2_X2 _f_permutation__round__U5386  ( .A(_f_permutation__round_in[1541]), 
        .B(_f_permutation__round__n2358 ), .Z(_f_permutation__round__c[5] ) );
  XOR2_X2 _f_permutation__round__U5385  ( .A(_f_permutation__round__n1838 ), 
        .B(_f_permutation__round__n1837 ), .Z(_f_permutation__round__n2102 )
         );
  XOR2_X2 _f_permutation__round__U5384  ( .A(SYNOPSYS_UNCONNECTED_827), .B(
        _f_permutation__round__n1839 ), .Z(_f_permutation__round__n1837 ) );
  XOR2_X2 _f_permutation__round__U5383  ( .A(SYNOPSYS_UNCONNECTED_187), .B(
        SYNOPSYS_UNCONNECTED_507), .Z(_f_permutation__round__n1838 ) );
  XOR2_X2 _f_permutation__round__U5382  ( .A(_f_permutation__round_in[1541]), 
        .B(_f_permutation__round_in[1221]), .Z(_f_permutation__round__n1839 )
         );
  XOR2_X2 _f_permutation__round__U5381  ( .A(_f_permutation__round__n1841 ), 
        .B(_f_permutation__round__n1840 ), .Z(_f_permutation__round__n2344 )
         );
  XOR2_X2 _f_permutation__round__U5380  ( .A(SYNOPSYS_UNCONNECTED_1018), .B(
        _f_permutation__round__n1842 ), .Z(_f_permutation__round__n1840 ) );
  XOR2_X2 _f_permutation__round__U5379  ( .A(SYNOPSYS_UNCONNECTED_378), .B(
        SYNOPSYS_UNCONNECTED_698), .Z(_f_permutation__round__n1841 ) );
  XOR2_X2 _f_permutation__round__U5378  ( .A(_f_permutation__round_in[1350]), 
        .B(_f_permutation__round_in[1030]), .Z(_f_permutation__round__n1842 )
         );
  XOR2_X2 _f_permutation__round__U5377  ( .A(_f_permutation__round__n2102 ), 
        .B(_f_permutation__round__n2344 ), .Z(_f_permutation__round__n2103 )
         );
  XOR2_X2 _f_permutation__round__U5376  ( .A(SYNOPSYS_UNCONNECTED_1082), .B(
        _f_permutation__round__n2103 ), .Z(_f_permutation__round__c[1542] ) );
  XOR2_X2 _f_permutation__round__U5375  ( .A(_f_permutation__round__n1844 ), 
        .B(_f_permutation__round__n1843 ), .Z(_f_permutation__round__n2554 )
         );
  XOR2_X2 _f_permutation__round__U5374  ( .A(SYNOPSYS_UNCONNECTED_956), .B(
        _f_permutation__round__n1845 ), .Z(_f_permutation__round__n1843 ) );
  XOR2_X2 _f_permutation__round__U5373  ( .A(SYNOPSYS_UNCONNECTED_316), .B(
        SYNOPSYS_UNCONNECTED_636), .Z(_f_permutation__round__n1844 ) );
  XOR2_X2 _f_permutation__round__U5372  ( .A(_f_permutation__round_in[1412]), 
        .B(_f_permutation__round_in[1092]), .Z(_f_permutation__round__n1845 )
         );
  XOR2_X2 _f_permutation__round__U5371  ( .A(_f_permutation__round__n2102 ), 
        .B(_f_permutation__round__n2554 ), .Z(_f_permutation__round__n2104 )
         );
  XOR2_X2 _f_permutation__round__U5370  ( .A(SYNOPSYS_UNCONNECTED_891), .B(
        _f_permutation__round__n2104 ), .Z(_f_permutation__round__c[581] ) );
  XOR2_X2 _f_permutation__round__U5369  ( .A(SYNOPSYS_UNCONNECTED_762), .B(
        _f_permutation__round__n2103 ), .Z(_f_permutation__round__c[1478] ) );
  XOR2_X2 _f_permutation__round__U5368  ( .A(SYNOPSYS_UNCONNECTED_571), .B(
        _f_permutation__round__n2104 ), .Z(_f_permutation__round__c[517] ) );
  XOR2_X2 _f_permutation__round__U5367  ( .A(SYNOPSYS_UNCONNECTED_442), .B(
        _f_permutation__round__n2103 ), .Z(_f_permutation__round__c[1414] ) );
  XOR2_X2 _f_permutation__round__U5366  ( .A(SYNOPSYS_UNCONNECTED_251), .B(
        _f_permutation__round__n2104 ), .Z(_f_permutation__round__c[453] ) );
  XOR2_X2 _f_permutation__round__U5365  ( .A(SYNOPSYS_UNCONNECTED_122), .B(
        _f_permutation__round__n2103 ), .Z(_f_permutation__round__c[1350] ) );
  XOR2_X2 _f_permutation__round__U5364  ( .A(_f_permutation__round_in[1157]), 
        .B(_f_permutation__round__n2104 ), .Z(_f_permutation__round__c[389] )
         );
  XOR2_X2 _f_permutation__round__U5363  ( .A(_f_permutation__round_in[1286]), 
        .B(_f_permutation__round__n2103 ), .Z(_f_permutation__round__c[1286] )
         );
  XOR2_X2 _f_permutation__round__U5362  ( .A(_f_permutation__round_in[1477]), 
        .B(_f_permutation__round__n2104 ), .Z(_f_permutation__round__c[325] )
         );
  XOR2_X2 _f_permutation__round__U5361  ( .A(_f_permutation__round__n1847 ), 
        .B(_f_permutation__round__n1846 ), .Z(_f_permutation__round__n2361 )
         );
  XOR2_X2 _f_permutation__round__U5360  ( .A(SYNOPSYS_UNCONNECTED_893), .B(
        _f_permutation__round__n1848 ), .Z(_f_permutation__round__n1846 ) );
  XOR2_X2 _f_permutation__round__U5359  ( .A(SYNOPSYS_UNCONNECTED_253), .B(
        SYNOPSYS_UNCONNECTED_573), .Z(_f_permutation__round__n1847 ) );
  XOR2_X2 _f_permutation__round__U5358  ( .A(_f_permutation__round_in[1475]), 
        .B(_f_permutation__round_in[1155]), .Z(_f_permutation__round__n1848 )
         );
  XOR2_X2 _f_permutation__round__U5357  ( .A(_f_permutation__round__n1850 ), 
        .B(_f_permutation__round__n1849 ), .Z(_f_permutation__round__n2550 )
         );
  XOR2_X2 _f_permutation__round__U5356  ( .A(SYNOPSYS_UNCONNECTED_1084), .B(
        _f_permutation__round__n1851 ), .Z(_f_permutation__round__n1849 ) );
  XOR2_X2 _f_permutation__round__U5355  ( .A(SYNOPSYS_UNCONNECTED_444), .B(
        SYNOPSYS_UNCONNECTED_764), .Z(_f_permutation__round__n1850 ) );
  XOR2_X2 _f_permutation__round__U5354  ( .A(_f_permutation__round_in[1284]), 
        .B(SYNOPSYS_UNCONNECTED_124), .Z(_f_permutation__round__n1851 ) );
  XOR2_X2 _f_permutation__round__U5353  ( .A(_f_permutation__round__n2361 ), 
        .B(_f_permutation__round__n2550 ), .Z(_f_permutation__round__n2362 )
         );
  XOR2_X2 _f_permutation__round__U5352  ( .A(_f_permutation__round_in[1540]), 
        .B(_f_permutation__round__n2362 ), .Z(_f_permutation__round__c[4] ) );
  XOR2_X2 _f_permutation__round__U5351  ( .A(_f_permutation__round__n1853 ), 
        .B(_f_permutation__round__n1852 ), .Z(_f_permutation__round__n2105 )
         );
  XOR2_X2 _f_permutation__round__U5350  ( .A(SYNOPSYS_UNCONNECTED_828), .B(
        _f_permutation__round__n1854 ), .Z(_f_permutation__round__n1852 ) );
  XOR2_X2 _f_permutation__round__U5349  ( .A(SYNOPSYS_UNCONNECTED_188), .B(
        SYNOPSYS_UNCONNECTED_508), .Z(_f_permutation__round__n1853 ) );
  XOR2_X2 _f_permutation__round__U5348  ( .A(_f_permutation__round_in[1540]), 
        .B(_f_permutation__round_in[1220]), .Z(_f_permutation__round__n1854 )
         );
  XOR2_X2 _f_permutation__round__U5347  ( .A(_f_permutation__round__n1856 ), 
        .B(_f_permutation__round__n1855 ), .Z(_f_permutation__round__n2348 )
         );
  XOR2_X2 _f_permutation__round__U5346  ( .A(SYNOPSYS_UNCONNECTED_1019), .B(
        _f_permutation__round__n1857 ), .Z(_f_permutation__round__n1855 ) );
  XOR2_X2 _f_permutation__round__U5345  ( .A(SYNOPSYS_UNCONNECTED_379), .B(
        SYNOPSYS_UNCONNECTED_699), .Z(_f_permutation__round__n1856 ) );
  XOR2_X2 _f_permutation__round__U5344  ( .A(_f_permutation__round_in[1349]), 
        .B(_f_permutation__round_in[1029]), .Z(_f_permutation__round__n1857 )
         );
  XOR2_X2 _f_permutation__round__U5343  ( .A(_f_permutation__round__n2105 ), 
        .B(_f_permutation__round__n2348 ), .Z(_f_permutation__round__n2106 )
         );
  XOR2_X2 _f_permutation__round__U5342  ( .A(SYNOPSYS_UNCONNECTED_1083), .B(
        _f_permutation__round__n2106 ), .Z(_f_permutation__round__c[1541] ) );
  XOR2_X2 _f_permutation__round__U5341  ( .A(_f_permutation__round__n1859 ), 
        .B(_f_permutation__round__n1858 ), .Z(_f_permutation__round__n2557 )
         );
  XOR2_X2 _f_permutation__round__U5340  ( .A(SYNOPSYS_UNCONNECTED_957), .B(
        _f_permutation__round__n1860 ), .Z(_f_permutation__round__n1858 ) );
  XOR2_X2 _f_permutation__round__U5339  ( .A(SYNOPSYS_UNCONNECTED_317), .B(
        SYNOPSYS_UNCONNECTED_637), .Z(_f_permutation__round__n1859 ) );
  XOR2_X2 _f_permutation__round__U5338  ( .A(_f_permutation__round_in[1411]), 
        .B(_f_permutation__round_in[1091]), .Z(_f_permutation__round__n1860 )
         );
  XOR2_X2 _f_permutation__round__U5337  ( .A(_f_permutation__round__n2105 ), 
        .B(_f_permutation__round__n2557 ), .Z(_f_permutation__round__n2107 )
         );
  XOR2_X2 _f_permutation__round__U5336  ( .A(SYNOPSYS_UNCONNECTED_892), .B(
        _f_permutation__round__n2107 ), .Z(_f_permutation__round__c[580] ) );
  XOR2_X2 _f_permutation__round__U5335  ( .A(SYNOPSYS_UNCONNECTED_763), .B(
        _f_permutation__round__n2106 ), .Z(_f_permutation__round__c[1477] ) );
  XOR2_X2 _f_permutation__round__U5334  ( .A(SYNOPSYS_UNCONNECTED_572), .B(
        _f_permutation__round__n2107 ), .Z(_f_permutation__round__c[516] ) );
  XOR2_X2 _f_permutation__round__U5333  ( .A(SYNOPSYS_UNCONNECTED_443), .B(
        _f_permutation__round__n2106 ), .Z(_f_permutation__round__c[1413] ) );
  XOR2_X2 _f_permutation__round__U5332  ( .A(SYNOPSYS_UNCONNECTED_252), .B(
        _f_permutation__round__n2107 ), .Z(_f_permutation__round__c[452] ) );
  XOR2_X2 _f_permutation__round__U5331  ( .A(SYNOPSYS_UNCONNECTED_123), .B(
        _f_permutation__round__n2106 ), .Z(_f_permutation__round__c[1349] ) );
  XOR2_X2 _f_permutation__round__U5330  ( .A(_f_permutation__round_in[1156]), 
        .B(_f_permutation__round__n2107 ), .Z(_f_permutation__round__c[388] )
         );
  XOR2_X2 _f_permutation__round__U5329  ( .A(_f_permutation__round_in[1285]), 
        .B(_f_permutation__round__n2106 ), .Z(_f_permutation__round__c[1285] )
         );
  XOR2_X2 _f_permutation__round__U5328  ( .A(_f_permutation__round_in[1476]), 
        .B(_f_permutation__round__n2107 ), .Z(_f_permutation__round__c[324] )
         );
  XOR2_X2 _f_permutation__round__U5327  ( .A(_f_permutation__round__n1862 ), 
        .B(_f_permutation__round__n1861 ), .Z(_f_permutation__round__n2365 )
         );
  XOR2_X2 _f_permutation__round__U5326  ( .A(SYNOPSYS_UNCONNECTED_894), .B(
        _f_permutation__round__n1863 ), .Z(_f_permutation__round__n1861 ) );
  XOR2_X2 _f_permutation__round__U5325  ( .A(SYNOPSYS_UNCONNECTED_254), .B(
        SYNOPSYS_UNCONNECTED_574), .Z(_f_permutation__round__n1862 ) );
  XOR2_X2 _f_permutation__round__U5324  ( .A(_f_permutation__round_in[1474]), 
        .B(_f_permutation__round_in[1154]), .Z(_f_permutation__round__n1863 )
         );
  XOR2_X2 _f_permutation__round__U5323  ( .A(_f_permutation__round__n1865 ), 
        .B(_f_permutation__round__n1864 ), .Z(_f_permutation__round__n2553 )
         );
  XOR2_X2 _f_permutation__round__U5322  ( .A(SYNOPSYS_UNCONNECTED_1085), .B(
        _f_permutation__round__n1866 ), .Z(_f_permutation__round__n1864 ) );
  XOR2_X2 _f_permutation__round__U5321  ( .A(SYNOPSYS_UNCONNECTED_445), .B(
        SYNOPSYS_UNCONNECTED_765), .Z(_f_permutation__round__n1865 ) );
  XOR2_X2 _f_permutation__round__U5320  ( .A(_f_permutation__round_in[1283]), 
        .B(SYNOPSYS_UNCONNECTED_125), .Z(_f_permutation__round__n1866 ) );
  XOR2_X2 _f_permutation__round__U5319  ( .A(_f_permutation__round__n2365 ), 
        .B(_f_permutation__round__n2553 ), .Z(_f_permutation__round__n2366 )
         );
  XOR2_X2 _f_permutation__round__U5318  ( .A(_f_permutation__round_in[1539]), 
        .B(_f_permutation__round__n2366 ), .Z(_f_permutation__round__c[3] ) );
  XOR2_X2 _f_permutation__round__U5317  ( .A(_f_permutation__round__n1868 ), 
        .B(_f_permutation__round__n1867 ), .Z(_f_permutation__round__n2108 )
         );
  XOR2_X2 _f_permutation__round__U5316  ( .A(SYNOPSYS_UNCONNECTED_829), .B(
        _f_permutation__round__n1869 ), .Z(_f_permutation__round__n1867 ) );
  XOR2_X2 _f_permutation__round__U5315  ( .A(SYNOPSYS_UNCONNECTED_189), .B(
        SYNOPSYS_UNCONNECTED_509), .Z(_f_permutation__round__n1868 ) );
  XOR2_X2 _f_permutation__round__U5314  ( .A(_f_permutation__round_in[1539]), 
        .B(_f_permutation__round_in[1219]), .Z(_f_permutation__round__n1869 )
         );
  XOR2_X2 _f_permutation__round__U5313  ( .A(_f_permutation__round__n1871 ), 
        .B(_f_permutation__round__n1870 ), .Z(_f_permutation__round__n2352 )
         );
  XOR2_X2 _f_permutation__round__U5312  ( .A(SYNOPSYS_UNCONNECTED_1020), .B(
        _f_permutation__round__n1872 ), .Z(_f_permutation__round__n1870 ) );
  XOR2_X2 _f_permutation__round__U5311  ( .A(SYNOPSYS_UNCONNECTED_380), .B(
        SYNOPSYS_UNCONNECTED_700), .Z(_f_permutation__round__n1871 ) );
  XOR2_X2 _f_permutation__round__U5310  ( .A(_f_permutation__round_in[1348]), 
        .B(_f_permutation__round_in[1028]), .Z(_f_permutation__round__n1872 )
         );
  XOR2_X2 _f_permutation__round__U5309  ( .A(_f_permutation__round__n2108 ), 
        .B(_f_permutation__round__n2352 ), .Z(_f_permutation__round__n2109 )
         );
  XOR2_X2 _f_permutation__round__U5308  ( .A(SYNOPSYS_UNCONNECTED_1084), .B(
        _f_permutation__round__n2109 ), .Z(_f_permutation__round__c[1540] ) );
  XOR2_X2 _f_permutation__round__U5307  ( .A(_f_permutation__round__n1874 ), 
        .B(_f_permutation__round__n1873 ), .Z(_f_permutation__round__n2560 )
         );
  XOR2_X2 _f_permutation__round__U5306  ( .A(SYNOPSYS_UNCONNECTED_958), .B(
        _f_permutation__round__n1875 ), .Z(_f_permutation__round__n1873 ) );
  XOR2_X2 _f_permutation__round__U5305  ( .A(SYNOPSYS_UNCONNECTED_318), .B(
        SYNOPSYS_UNCONNECTED_638), .Z(_f_permutation__round__n1874 ) );
  XOR2_X2 _f_permutation__round__U5304  ( .A(_f_permutation__round_in[1410]), 
        .B(_f_permutation__round_in[1090]), .Z(_f_permutation__round__n1875 )
         );
  XOR2_X2 _f_permutation__round__U5303  ( .A(_f_permutation__round__n2108 ), 
        .B(_f_permutation__round__n2560 ), .Z(_f_permutation__round__n2110 )
         );
  XOR2_X2 _f_permutation__round__U5302  ( .A(SYNOPSYS_UNCONNECTED_893), .B(
        _f_permutation__round__n2110 ), .Z(_f_permutation__round__c[579] ) );
  XOR2_X2 _f_permutation__round__U5301  ( .A(SYNOPSYS_UNCONNECTED_764), .B(
        _f_permutation__round__n2109 ), .Z(_f_permutation__round__c[1476] ) );
  XOR2_X2 _f_permutation__round__U5300  ( .A(SYNOPSYS_UNCONNECTED_573), .B(
        _f_permutation__round__n2110 ), .Z(_f_permutation__round__c[515] ) );
  XOR2_X2 _f_permutation__round__U5299  ( .A(SYNOPSYS_UNCONNECTED_444), .B(
        _f_permutation__round__n2109 ), .Z(_f_permutation__round__c[1412] ) );
  XOR2_X2 _f_permutation__round__U5298  ( .A(SYNOPSYS_UNCONNECTED_253), .B(
        _f_permutation__round__n2110 ), .Z(_f_permutation__round__c[451] ) );
  XOR2_X2 _f_permutation__round__U5297  ( .A(SYNOPSYS_UNCONNECTED_124), .B(
        _f_permutation__round__n2109 ), .Z(_f_permutation__round__c[1348] ) );
  XOR2_X2 _f_permutation__round__U5296  ( .A(_f_permutation__round_in[1155]), 
        .B(_f_permutation__round__n2110 ), .Z(_f_permutation__round__c[387] )
         );
  XOR2_X2 _f_permutation__round__U5295  ( .A(_f_permutation__round_in[1284]), 
        .B(_f_permutation__round__n2109 ), .Z(_f_permutation__round__c[1284] )
         );
  XOR2_X2 _f_permutation__round__U5294  ( .A(_f_permutation__round_in[1475]), 
        .B(_f_permutation__round__n2110 ), .Z(_f_permutation__round__c[323] )
         );
  XOR2_X2 _f_permutation__round__U5293  ( .A(_f_permutation__round__n1877 ), 
        .B(_f_permutation__round__n1876 ), .Z(_f_permutation__round__n2369 )
         );
  XOR2_X2 _f_permutation__round__U5292  ( .A(SYNOPSYS_UNCONNECTED_895), .B(
        _f_permutation__round__n1878 ), .Z(_f_permutation__round__n1876 ) );
  XOR2_X2 _f_permutation__round__U5291  ( .A(SYNOPSYS_UNCONNECTED_255), .B(
        SYNOPSYS_UNCONNECTED_575), .Z(_f_permutation__round__n1877 ) );
  XOR2_X2 _f_permutation__round__U5290  ( .A(_f_permutation__round_in[1473]), 
        .B(_f_permutation__round_in[1153]), .Z(_f_permutation__round__n1878 )
         );
  XOR2_X2 _f_permutation__round__U5289  ( .A(_f_permutation__round__n1880 ), 
        .B(_f_permutation__round__n1879 ), .Z(_f_permutation__round__n2556 )
         );
  XOR2_X2 _f_permutation__round__U5288  ( .A(SYNOPSYS_UNCONNECTED_1086), .B(
        _f_permutation__round__n1881 ), .Z(_f_permutation__round__n1879 ) );
  XOR2_X2 _f_permutation__round__U5287  ( .A(SYNOPSYS_UNCONNECTED_446), .B(
        SYNOPSYS_UNCONNECTED_766), .Z(_f_permutation__round__n1880 ) );
  XOR2_X2 _f_permutation__round__U5286  ( .A(_f_permutation__round_in[1282]), 
        .B(SYNOPSYS_UNCONNECTED_126), .Z(_f_permutation__round__n1881 ) );
  XOR2_X2 _f_permutation__round__U5285  ( .A(_f_permutation__round__n2369 ), 
        .B(_f_permutation__round__n2556 ), .Z(_f_permutation__round__n2370 )
         );
  XOR2_X2 _f_permutation__round__U5284  ( .A(_f_permutation__round_in[1538]), 
        .B(_f_permutation__round__n2370 ), .Z(_f_permutation__round__c[2] ) );
  XOR2_X2 _f_permutation__round__U5283  ( .A(_f_permutation__round__n1883 ), 
        .B(_f_permutation__round__n1882 ), .Z(_f_permutation__round__n2111 )
         );
  XOR2_X2 _f_permutation__round__U5282  ( .A(SYNOPSYS_UNCONNECTED_830), .B(
        _f_permutation__round__n1884 ), .Z(_f_permutation__round__n1882 ) );
  XOR2_X2 _f_permutation__round__U5281  ( .A(SYNOPSYS_UNCONNECTED_190), .B(
        SYNOPSYS_UNCONNECTED_510), .Z(_f_permutation__round__n1883 ) );
  XOR2_X2 _f_permutation__round__U5280  ( .A(_f_permutation__round_in[1538]), 
        .B(_f_permutation__round_in[1218]), .Z(_f_permutation__round__n1884 )
         );
  XOR2_X2 _f_permutation__round__U5279  ( .A(_f_permutation__round__n1886 ), 
        .B(_f_permutation__round__n1885 ), .Z(_f_permutation__round__n2356 )
         );
  XOR2_X2 _f_permutation__round__U5278  ( .A(SYNOPSYS_UNCONNECTED_1021), .B(
        _f_permutation__round__n1887 ), .Z(_f_permutation__round__n1885 ) );
  XOR2_X2 _f_permutation__round__U5277  ( .A(SYNOPSYS_UNCONNECTED_381), .B(
        SYNOPSYS_UNCONNECTED_701), .Z(_f_permutation__round__n1886 ) );
  XOR2_X2 _f_permutation__round__U5276  ( .A(_f_permutation__round_in[1347]), 
        .B(_f_permutation__round_in[1027]), .Z(_f_permutation__round__n1887 )
         );
  XOR2_X2 _f_permutation__round__U5275  ( .A(_f_permutation__round__n2111 ), 
        .B(_f_permutation__round__n2356 ), .Z(_f_permutation__round__n2112 )
         );
  XOR2_X2 _f_permutation__round__U5274  ( .A(SYNOPSYS_UNCONNECTED_1085), .B(
        _f_permutation__round__n2112 ), .Z(_f_permutation__round__c[1539] ) );
  XOR2_X2 _f_permutation__round__U5273  ( .A(_f_permutation__round__n1889 ), 
        .B(_f_permutation__round__n1888 ), .Z(_f_permutation__round__n25630 )
         );
  XOR2_X2 _f_permutation__round__U5272  ( .A(SYNOPSYS_UNCONNECTED_959), .B(
        _f_permutation__round__n1890 ), .Z(_f_permutation__round__n1888 ) );
  XOR2_X2 _f_permutation__round__U5271  ( .A(SYNOPSYS_UNCONNECTED_319), .B(
        SYNOPSYS_UNCONNECTED_639), .Z(_f_permutation__round__n1889 ) );
  XOR2_X2 _f_permutation__round__U5270  ( .A(_f_permutation__round_in[1409]), 
        .B(_f_permutation__round_in[1089]), .Z(_f_permutation__round__n1890 )
         );
  XOR2_X2 _f_permutation__round__U5269  ( .A(_f_permutation__round__n2111 ), 
        .B(_f_permutation__round__n25630 ), .Z(_f_permutation__round__n2113 )
         );
  XOR2_X2 _f_permutation__round__U5268  ( .A(SYNOPSYS_UNCONNECTED_894), .B(
        _f_permutation__round__n2113 ), .Z(_f_permutation__round__c[578] ) );
  XOR2_X2 _f_permutation__round__U5267  ( .A(SYNOPSYS_UNCONNECTED_765), .B(
        _f_permutation__round__n2112 ), .Z(_f_permutation__round__c[1475] ) );
  XOR2_X2 _f_permutation__round__U5266  ( .A(SYNOPSYS_UNCONNECTED_574), .B(
        _f_permutation__round__n2113 ), .Z(_f_permutation__round__c[514] ) );
  XOR2_X2 _f_permutation__round__U5265  ( .A(SYNOPSYS_UNCONNECTED_445), .B(
        _f_permutation__round__n2112 ), .Z(_f_permutation__round__c[1411] ) );
  XOR2_X2 _f_permutation__round__U5264  ( .A(SYNOPSYS_UNCONNECTED_254), .B(
        _f_permutation__round__n2113 ), .Z(_f_permutation__round__c[450] ) );
  XOR2_X2 _f_permutation__round__U5263  ( .A(SYNOPSYS_UNCONNECTED_125), .B(
        _f_permutation__round__n2112 ), .Z(_f_permutation__round__c[1347] ) );
  XOR2_X2 _f_permutation__round__U5262  ( .A(_f_permutation__round_in[1154]), 
        .B(_f_permutation__round__n2113 ), .Z(_f_permutation__round__c[386] )
         );
  XOR2_X2 _f_permutation__round__U5261  ( .A(_f_permutation__round_in[1283]), 
        .B(_f_permutation__round__n2112 ), .Z(_f_permutation__round__c[1283] )
         );
  XOR2_X2 _f_permutation__round__U5260  ( .A(_f_permutation__round_in[1474]), 
        .B(_f_permutation__round__n2113 ), .Z(_f_permutation__round__c[322] )
         );
  XOR2_X2 _f_permutation__round__U5259  ( .A(_f_permutation__round__n1892 ), 
        .B(_f_permutation__round__n1891 ), .Z(_f_permutation__round__n2373 )
         );
  XOR2_X2 _f_permutation__round__U5258  ( .A(SYNOPSYS_UNCONNECTED_896), .B(
        _f_permutation__round__n1893 ), .Z(_f_permutation__round__n1891 ) );
  XOR2_X2 _f_permutation__round__U5257  ( .A(SYNOPSYS_UNCONNECTED_256), .B(
        SYNOPSYS_UNCONNECTED_576), .Z(_f_permutation__round__n1892 ) );
  XOR2_X2 _f_permutation__round__U5256  ( .A(_f_permutation__round_in[1472]), 
        .B(_f_permutation__round_in[1152]), .Z(_f_permutation__round__n1893 )
         );
  XOR2_X2 _f_permutation__round__U5255  ( .A(_f_permutation__round__n1895 ), 
        .B(_f_permutation__round__n1894 ), .Z(_f_permutation__round__n2559 )
         );
  XOR2_X2 _f_permutation__round__U5254  ( .A(SYNOPSYS_UNCONNECTED_1087), .B(
        _f_permutation__round__n1896 ), .Z(_f_permutation__round__n1894 ) );
  XOR2_X2 _f_permutation__round__U5253  ( .A(SYNOPSYS_UNCONNECTED_447), .B(
        SYNOPSYS_UNCONNECTED_767), .Z(_f_permutation__round__n1895 ) );
  XOR2_X2 _f_permutation__round__U5252  ( .A(_f_permutation__round_in[1281]), 
        .B(SYNOPSYS_UNCONNECTED_127), .Z(_f_permutation__round__n1896 ) );
  XOR2_X2 _f_permutation__round__U5251  ( .A(_f_permutation__round__n2373 ), 
        .B(_f_permutation__round__n2559 ), .Z(_f_permutation__round__n2374 )
         );
  XOR2_X2 _f_permutation__round__U5250  ( .A(_f_permutation__round_in[1537]), 
        .B(_f_permutation__round__n2374 ), .Z(_f_permutation__round__c[1] ) );
  XOR2_X2 _f_permutation__round__U5249  ( .A(_f_permutation__round__n1898 ), 
        .B(_f_permutation__round__n1897 ), .Z(_f_permutation__round__n2114 )
         );
  XOR2_X2 _f_permutation__round__U5248  ( .A(SYNOPSYS_UNCONNECTED_831), .B(
        _f_permutation__round__n1899 ), .Z(_f_permutation__round__n1897 ) );
  XOR2_X2 _f_permutation__round__U5247  ( .A(SYNOPSYS_UNCONNECTED_191), .B(
        SYNOPSYS_UNCONNECTED_511), .Z(_f_permutation__round__n1898 ) );
  XOR2_X2 _f_permutation__round__U5246  ( .A(_f_permutation__round_in[1537]), 
        .B(_f_permutation__round_in[1217]), .Z(_f_permutation__round__n1899 )
         );
  XOR2_X2 _f_permutation__round__U5245  ( .A(_f_permutation__round__n1901 ), 
        .B(_f_permutation__round__n1900 ), .Z(_f_permutation__round__n2360 )
         );
  XOR2_X2 _f_permutation__round__U5244  ( .A(SYNOPSYS_UNCONNECTED_1022), .B(
        _f_permutation__round__n1902 ), .Z(_f_permutation__round__n1900 ) );
  XOR2_X2 _f_permutation__round__U5243  ( .A(SYNOPSYS_UNCONNECTED_382), .B(
        SYNOPSYS_UNCONNECTED_702), .Z(_f_permutation__round__n1901 ) );
  XOR2_X2 _f_permutation__round__U5242  ( .A(_f_permutation__round_in[1346]), 
        .B(_f_permutation__round_in[1026]), .Z(_f_permutation__round__n1902 )
         );
  XOR2_X2 _f_permutation__round__U5241  ( .A(_f_permutation__round__n2114 ), 
        .B(_f_permutation__round__n2360 ), .Z(_f_permutation__round__n2115 )
         );
  XOR2_X2 _f_permutation__round__U5240  ( .A(SYNOPSYS_UNCONNECTED_1086), .B(
        _f_permutation__round__n2115 ), .Z(_f_permutation__round__c[1538] ) );
  XOR2_X2 _f_permutation__round__U5239  ( .A(_f_permutation__round__n1904 ), 
        .B(_f_permutation__round__n1903 ), .Z(_f_permutation__round__n2566 )
         );
  XOR2_X2 _f_permutation__round__U5238  ( .A(SYNOPSYS_UNCONNECTED_960), .B(
        _f_permutation__round__n1905 ), .Z(_f_permutation__round__n1903 ) );
  XOR2_X2 _f_permutation__round__U5237  ( .A(SYNOPSYS_UNCONNECTED_320), .B(
        SYNOPSYS_UNCONNECTED_640), .Z(_f_permutation__round__n1904 ) );
  XOR2_X2 _f_permutation__round__U5236  ( .A(_f_permutation__round_in[1408]), 
        .B(_f_permutation__round_in[1088]), .Z(_f_permutation__round__n1905 )
         );
  XOR2_X2 _f_permutation__round__U5235  ( .A(_f_permutation__round__n2114 ), 
        .B(_f_permutation__round__n2566 ), .Z(_f_permutation__round__n2116 )
         );
  XOR2_X2 _f_permutation__round__U5234  ( .A(SYNOPSYS_UNCONNECTED_895), .B(
        _f_permutation__round__n2116 ), .Z(_f_permutation__round__c[577] ) );
  XOR2_X2 _f_permutation__round__U5233  ( .A(SYNOPSYS_UNCONNECTED_766), .B(
        _f_permutation__round__n2115 ), .Z(_f_permutation__round__c[1474] ) );
  XOR2_X2 _f_permutation__round__U5232  ( .A(SYNOPSYS_UNCONNECTED_575), .B(
        _f_permutation__round__n2116 ), .Z(_f_permutation__round__c[513] ) );
  XOR2_X2 _f_permutation__round__U5231  ( .A(SYNOPSYS_UNCONNECTED_446), .B(
        _f_permutation__round__n2115 ), .Z(_f_permutation__round__c[1410] ) );
  XOR2_X2 _f_permutation__round__U5230  ( .A(SYNOPSYS_UNCONNECTED_255), .B(
        _f_permutation__round__n2116 ), .Z(_f_permutation__round__c[449] ) );
  XOR2_X2 _f_permutation__round__U5229  ( .A(SYNOPSYS_UNCONNECTED_126), .B(
        _f_permutation__round__n2115 ), .Z(_f_permutation__round__c[1346] ) );
  XOR2_X2 _f_permutation__round__U5228  ( .A(_f_permutation__round_in[1153]), 
        .B(_f_permutation__round__n2116 ), .Z(_f_permutation__round__c[385] )
         );
  XOR2_X2 _f_permutation__round__U5227  ( .A(_f_permutation__round_in[1282]), 
        .B(_f_permutation__round__n2115 ), .Z(_f_permutation__round__c[1282] )
         );
  XOR2_X2 _f_permutation__round__U5226  ( .A(_f_permutation__round_in[1473]), 
        .B(_f_permutation__round__n2116 ), .Z(_f_permutation__round__c[321] )
         );
  XOR2_X2 _f_permutation__round__U5225  ( .A(_f_permutation__round__n1907 ), 
        .B(_f_permutation__round__n1906 ), .Z(_f_permutation__round__n2121 )
         );
  XOR2_X2 _f_permutation__round__U5224  ( .A(SYNOPSYS_UNCONNECTED_833), .B(
        _f_permutation__round__n1908 ), .Z(_f_permutation__round__n1906 ) );
  XOR2_X2 _f_permutation__round__U5223  ( .A(SYNOPSYS_UNCONNECTED_193), .B(
        SYNOPSYS_UNCONNECTED_513), .Z(_f_permutation__round__n1907 ) );
  XOR2_X2 _f_permutation__round__U5222  ( .A(_f_permutation__round_in[1535]), 
        .B(_f_permutation__round_in[1215]), .Z(_f_permutation__round__n1908 )
         );
  XOR2_X2 _f_permutation__round__U5221  ( .A(_f_permutation__round__n1910 ), 
        .B(_f_permutation__round__n1909 ), .Z(_f_permutation__round__n2562 )
         );
  XOR2_X2 _f_permutation__round__U5220  ( .A(SYNOPSYS_UNCONNECTED_1088), .B(
        _f_permutation__round__n1911 ), .Z(_f_permutation__round__n1909 ) );
  XOR2_X2 _f_permutation__round__U5219  ( .A(SYNOPSYS_UNCONNECTED_448), .B(
        SYNOPSYS_UNCONNECTED_768), .Z(_f_permutation__round__n1910 ) );
  XOR2_X2 _f_permutation__round__U5218  ( .A(_f_permutation__round_in[1280]), 
        .B(SYNOPSYS_UNCONNECTED_128), .Z(_f_permutation__round__n1911 ) );
  XOR2_X2 _f_permutation__round__U5217  ( .A(_f_permutation__round__n2121 ), 
        .B(_f_permutation__round__n2562 ), .Z(_f_permutation__round__n2122 )
         );
  XOR2_X2 _f_permutation__round__U5216  ( .A(_f_permutation__round_in[1536]), 
        .B(_f_permutation__round__n2122 ), .Z(_f_permutation__round__c[0] ) );
  XOR2_X2 _f_permutation__round__U5215  ( .A(_f_permutation__round__n1913 ), 
        .B(_f_permutation__round__n1912 ), .Z(_f_permutation__round__n2117 )
         );
  XOR2_X2 _f_permutation__round__U5214  ( .A(SYNOPSYS_UNCONNECTED_832), .B(
        _f_permutation__round__n1914 ), .Z(_f_permutation__round__n1912 ) );
  XOR2_X2 _f_permutation__round__U5213  ( .A(SYNOPSYS_UNCONNECTED_192), .B(
        SYNOPSYS_UNCONNECTED_512), .Z(_f_permutation__round__n1913 ) );
  XOR2_X2 _f_permutation__round__U5212  ( .A(_f_permutation__round_in[1536]), 
        .B(_f_permutation__round_in[1216]), .Z(_f_permutation__round__n1914 )
         );
  XOR2_X2 _f_permutation__round__U5211  ( .A(_f_permutation__round__n1916 ), 
        .B(_f_permutation__round__n1915 ), .Z(_f_permutation__round__n2364 )
         );
  XOR2_X2 _f_permutation__round__U5210  ( .A(SYNOPSYS_UNCONNECTED_1023), .B(
        _f_permutation__round__n1917 ), .Z(_f_permutation__round__n1915 ) );
  XOR2_X2 _f_permutation__round__U5209  ( .A(SYNOPSYS_UNCONNECTED_383), .B(
        SYNOPSYS_UNCONNECTED_703), .Z(_f_permutation__round__n1916 ) );
  XOR2_X2 _f_permutation__round__U5208  ( .A(_f_permutation__round_in[1345]), 
        .B(_f_permutation__round_in[1025]), .Z(_f_permutation__round__n1917 )
         );
  XOR2_X2 _f_permutation__round__U5207  ( .A(_f_permutation__round__n2117 ), 
        .B(_f_permutation__round__n2364 ), .Z(_f_permutation__round__n2118 )
         );
  XOR2_X2 _f_permutation__round__U5206  ( .A(SYNOPSYS_UNCONNECTED_1087), .B(
        _f_permutation__round__n2118 ), .Z(_f_permutation__round__c[1537] ) );
  XOR2_X2 _f_permutation__round__U5205  ( .A(_f_permutation__round__n1919 ), 
        .B(_f_permutation__round__n1918 ), .Z(_f_permutation__round__n2377 )
         );
  XOR2_X2 _f_permutation__round__U5204  ( .A(SYNOPSYS_UNCONNECTED_897), .B(
        _f_permutation__round__n1920 ), .Z(_f_permutation__round__n1918 ) );
  XOR2_X2 _f_permutation__round__U5203  ( .A(SYNOPSYS_UNCONNECTED_257), .B(
        SYNOPSYS_UNCONNECTED_577), .Z(_f_permutation__round__n1919 ) );
  XOR2_X2 _f_permutation__round__U5202  ( .A(_f_permutation__round_in[1471]), 
        .B(_f_permutation__round_in[1151]), .Z(_f_permutation__round__n1920 )
         );
  XOR2_X2 _f_permutation__round__U5201  ( .A(_f_permutation__round__n2117 ), 
        .B(_f_permutation__round__n2377 ), .Z(_f_permutation__round__n2119 )
         );
  XOR2_X2 _f_permutation__round__U5200  ( .A(SYNOPSYS_UNCONNECTED_896), .B(
        _f_permutation__round__n2119 ), .Z(_f_permutation__round__c[576] ) );
  XOR2_X2 _f_permutation__round__U5199  ( .A(SYNOPSYS_UNCONNECTED_767), .B(
        _f_permutation__round__n2118 ), .Z(_f_permutation__round__c[1473] ) );
  XOR2_X2 _f_permutation__round__U5198  ( .A(SYNOPSYS_UNCONNECTED_576), .B(
        _f_permutation__round__n2119 ), .Z(_f_permutation__round__c[512] ) );
  XOR2_X2 _f_permutation__round__U5197  ( .A(SYNOPSYS_UNCONNECTED_447), .B(
        _f_permutation__round__n2118 ), .Z(_f_permutation__round__c[1409] ) );
  XOR2_X2 _f_permutation__round__U5196  ( .A(SYNOPSYS_UNCONNECTED_256), .B(
        _f_permutation__round__n2119 ), .Z(_f_permutation__round__c[448] ) );
  XOR2_X2 _f_permutation__round__U5195  ( .A(SYNOPSYS_UNCONNECTED_127), .B(
        _f_permutation__round__n2118 ), .Z(_f_permutation__round__c[1345] ) );
  XOR2_X2 _f_permutation__round__U5194  ( .A(_f_permutation__round_in[1152]), 
        .B(_f_permutation__round__n2119 ), .Z(_f_permutation__round__c[384] )
         );
  XOR2_X2 _f_permutation__round__U5193  ( .A(_f_permutation__round_in[1281]), 
        .B(_f_permutation__round__n2118 ), .Z(_f_permutation__round__c[1281] )
         );
  XOR2_X2 _f_permutation__round__U5192  ( .A(_f_permutation__round_in[1472]), 
        .B(_f_permutation__round__n2119 ), .Z(_f_permutation__round__c[320] )
         );
  XOR2_X2 _f_permutation__round__U5191  ( .A(_f_permutation__round__n2121 ), 
        .B(_f_permutation__round__n2120 ), .Z(_f_permutation__round__n2123 )
         );
  XOR2_X2 _f_permutation__round__U5190  ( .A(SYNOPSYS_UNCONNECTED_897), .B(
        _f_permutation__round__n2123 ), .Z(_f_permutation__round__c[959] ) );
  XOR2_X2 _f_permutation__round__U5189  ( .A(SYNOPSYS_UNCONNECTED_832), .B(
        _f_permutation__round__n2122 ), .Z(_f_permutation__round__c[256] ) );
  XOR2_X2 _f_permutation__round__U5188  ( .A(SYNOPSYS_UNCONNECTED_577), .B(
        _f_permutation__round__n2123 ), .Z(_f_permutation__round__c[895] ) );
  XOR2_X2 _f_permutation__round__U5187  ( .A(SYNOPSYS_UNCONNECTED_512), .B(
        _f_permutation__round__n2122 ), .Z(_f_permutation__round__c[192] ) );
  XOR2_X2 _f_permutation__round__U5186  ( .A(SYNOPSYS_UNCONNECTED_257), .B(
        _f_permutation__round__n2123 ), .Z(_f_permutation__round__c[831] ) );
  XOR2_X2 _f_permutation__round__U5185  ( .A(SYNOPSYS_UNCONNECTED_192), .B(
        _f_permutation__round__n2122 ), .Z(_f_permutation__round__c[128] ) );
  XOR2_X2 _f_permutation__round__U5184  ( .A(_f_permutation__round_in[1151]), 
        .B(_f_permutation__round__n2123 ), .Z(_f_permutation__round__c[767] )
         );
  XOR2_X2 _f_permutation__round__U5183  ( .A(_f_permutation__round_in[1216]), 
        .B(_f_permutation__round__n2122 ), .Z(_f_permutation__round__c[64] )
         );
  XOR2_X2 _f_permutation__round__U5182  ( .A(_f_permutation__round_in[1471]), 
        .B(_f_permutation__round__n2123 ), .Z(_f_permutation__round__c[703] )
         );
  XOR2_X2 _f_permutation__round__U5181  ( .A(_f_permutation__round__n2125 ), 
        .B(_f_permutation__round__n2124 ), .Z(_f_permutation__round__n2127 )
         );
  XOR2_X2 _f_permutation__round__U5180  ( .A(SYNOPSYS_UNCONNECTED_898), .B(
        _f_permutation__round__n2127 ), .Z(_f_permutation__round__c[958] ) );
  XOR2_X2 _f_permutation__round__U5179  ( .A(SYNOPSYS_UNCONNECTED_769), .B(
        _f_permutation__round__n2126 ), .Z(_f_permutation__round__c[319] ) );
  XOR2_X2 _f_permutation__round__U5178  ( .A(SYNOPSYS_UNCONNECTED_578), .B(
        _f_permutation__round__n2127 ), .Z(_f_permutation__round__c[894] ) );
  XOR2_X2 _f_permutation__round__U5177  ( .A(SYNOPSYS_UNCONNECTED_449), .B(
        _f_permutation__round__n2126 ), .Z(_f_permutation__round__c[255] ) );
  XOR2_X2 _f_permutation__round__U5176  ( .A(SYNOPSYS_UNCONNECTED_258), .B(
        _f_permutation__round__n2127 ), .Z(_f_permutation__round__c[830] ) );
  XOR2_X2 _f_permutation__round__U5175  ( .A(SYNOPSYS_UNCONNECTED_129), .B(
        _f_permutation__round__n2126 ), .Z(_f_permutation__round__c[191] ) );
  XOR2_X2 _f_permutation__round__U5174  ( .A(_f_permutation__round_in[1150]), 
        .B(_f_permutation__round__n2127 ), .Z(_f_permutation__round__c[766] )
         );
  XOR2_X2 _f_permutation__round__U5173  ( .A(_f_permutation__round_in[1279]), 
        .B(_f_permutation__round__n2126 ), .Z(_f_permutation__round__c[127] )
         );
  XOR2_X2 _f_permutation__round__U5172  ( .A(_f_permutation__round_in[1470]), 
        .B(_f_permutation__round__n2127 ), .Z(_f_permutation__round__c[702] )
         );
  XOR2_X2 _f_permutation__round__U5171  ( .A(_f_permutation__round__n2129 ), 
        .B(_f_permutation__round__n2128 ), .Z(_f_permutation__round__n2131 )
         );
  XOR2_X2 _f_permutation__round__U5170  ( .A(SYNOPSYS_UNCONNECTED_899), .B(
        _f_permutation__round__n2131 ), .Z(_f_permutation__round__c[957] ) );
  XOR2_X2 _f_permutation__round__U5169  ( .A(SYNOPSYS_UNCONNECTED_770), .B(
        _f_permutation__round__n2130 ), .Z(_f_permutation__round__c[318] ) );
  XOR2_X2 _f_permutation__round__U5168  ( .A(SYNOPSYS_UNCONNECTED_579), .B(
        _f_permutation__round__n2131 ), .Z(_f_permutation__round__c[893] ) );
  XOR2_X2 _f_permutation__round__U5167  ( .A(SYNOPSYS_UNCONNECTED_450), .B(
        _f_permutation__round__n2130 ), .Z(_f_permutation__round__c[254] ) );
  XOR2_X2 _f_permutation__round__U5166  ( .A(SYNOPSYS_UNCONNECTED_259), .B(
        _f_permutation__round__n2131 ), .Z(_f_permutation__round__c[829] ) );
  XOR2_X2 _f_permutation__round__U5165  ( .A(SYNOPSYS_UNCONNECTED_130), .B(
        _f_permutation__round__n2130 ), .Z(_f_permutation__round__c[190] ) );
  XOR2_X2 _f_permutation__round__U5164  ( .A(_f_permutation__round_in[1149]), 
        .B(_f_permutation__round__n2131 ), .Z(_f_permutation__round__c[765] )
         );
  XOR2_X2 _f_permutation__round__U5163  ( .A(_f_permutation__round_in[1278]), 
        .B(_f_permutation__round__n2130 ), .Z(_f_permutation__round__c[126] )
         );
  XOR2_X2 _f_permutation__round__U5162  ( .A(_f_permutation__round_in[1469]), 
        .B(_f_permutation__round__n2131 ), .Z(_f_permutation__round__c[701] )
         );
  XOR2_X2 _f_permutation__round__U5161  ( .A(_f_permutation__round__n2133 ), 
        .B(_f_permutation__round__n2132 ), .Z(_f_permutation__round__n2135 )
         );
  XOR2_X2 _f_permutation__round__U5160  ( .A(SYNOPSYS_UNCONNECTED_900), .B(
        _f_permutation__round__n2135 ), .Z(_f_permutation__round__c[956] ) );
  XOR2_X2 _f_permutation__round__U5159  ( .A(SYNOPSYS_UNCONNECTED_771), .B(
        _f_permutation__round__n2134 ), .Z(_f_permutation__round__c[317] ) );
  XOR2_X2 _f_permutation__round__U5158  ( .A(SYNOPSYS_UNCONNECTED_580), .B(
        _f_permutation__round__n2135 ), .Z(_f_permutation__round__c[892] ) );
  XOR2_X2 _f_permutation__round__U5157  ( .A(SYNOPSYS_UNCONNECTED_451), .B(
        _f_permutation__round__n2134 ), .Z(_f_permutation__round__c[253] ) );
  XOR2_X2 _f_permutation__round__U5156  ( .A(SYNOPSYS_UNCONNECTED_260), .B(
        _f_permutation__round__n2135 ), .Z(_f_permutation__round__c[828] ) );
  XOR2_X2 _f_permutation__round__U5155  ( .A(SYNOPSYS_UNCONNECTED_131), .B(
        _f_permutation__round__n2134 ), .Z(_f_permutation__round__c[189] ) );
  XOR2_X2 _f_permutation__round__U5154  ( .A(_f_permutation__round_in[1148]), 
        .B(_f_permutation__round__n2135 ), .Z(_f_permutation__round__c[764] )
         );
  XOR2_X2 _f_permutation__round__U5153  ( .A(_f_permutation__round_in[1277]), 
        .B(_f_permutation__round__n2134 ), .Z(_f_permutation__round__c[125] )
         );
  XOR2_X2 _f_permutation__round__U5152  ( .A(_f_permutation__round_in[1468]), 
        .B(_f_permutation__round__n2135 ), .Z(_f_permutation__round__c[700] )
         );
  XOR2_X2 _f_permutation__round__U5151  ( .A(_f_permutation__round__n2137 ), 
        .B(_f_permutation__round__n2136 ), .Z(_f_permutation__round__n2139 )
         );
  XOR2_X2 _f_permutation__round__U5150  ( .A(SYNOPSYS_UNCONNECTED_901), .B(
        _f_permutation__round__n2139 ), .Z(_f_permutation__round__c[955] ) );
  XOR2_X2 _f_permutation__round__U5149  ( .A(SYNOPSYS_UNCONNECTED_772), .B(
        _f_permutation__round__n2138 ), .Z(_f_permutation__round__c[316] ) );
  XOR2_X2 _f_permutation__round__U5148  ( .A(SYNOPSYS_UNCONNECTED_581), .B(
        _f_permutation__round__n2139 ), .Z(_f_permutation__round__c[891] ) );
  XOR2_X2 _f_permutation__round__U5147  ( .A(SYNOPSYS_UNCONNECTED_452), .B(
        _f_permutation__round__n2138 ), .Z(_f_permutation__round__c[252] ) );
  XOR2_X2 _f_permutation__round__U5146  ( .A(SYNOPSYS_UNCONNECTED_261), .B(
        _f_permutation__round__n2139 ), .Z(_f_permutation__round__c[827] ) );
  XOR2_X2 _f_permutation__round__U5145  ( .A(SYNOPSYS_UNCONNECTED_132), .B(
        _f_permutation__round__n2138 ), .Z(_f_permutation__round__c[188] ) );
  XOR2_X2 _f_permutation__round__U5144  ( .A(_f_permutation__round_in[1147]), 
        .B(_f_permutation__round__n2139 ), .Z(_f_permutation__round__c[763] )
         );
  XOR2_X2 _f_permutation__round__U5143  ( .A(_f_permutation__round_in[1276]), 
        .B(_f_permutation__round__n2138 ), .Z(_f_permutation__round__c[124] )
         );
  XOR2_X2 _f_permutation__round__U5142  ( .A(_f_permutation__round_in[1467]), 
        .B(_f_permutation__round__n2139 ), .Z(_f_permutation__round__c[699] )
         );
  XOR2_X2 _f_permutation__round__U5141  ( .A(_f_permutation__round__n2141 ), 
        .B(_f_permutation__round__n2140 ), .Z(_f_permutation__round__n2143 )
         );
  XOR2_X2 _f_permutation__round__U5140  ( .A(SYNOPSYS_UNCONNECTED_902), .B(
        _f_permutation__round__n2143 ), .Z(_f_permutation__round__c[954] ) );
  XOR2_X2 _f_permutation__round__U5139  ( .A(SYNOPSYS_UNCONNECTED_773), .B(
        _f_permutation__round__n2142 ), .Z(_f_permutation__round__c[315] ) );
  XOR2_X2 _f_permutation__round__U5138  ( .A(SYNOPSYS_UNCONNECTED_582), .B(
        _f_permutation__round__n2143 ), .Z(_f_permutation__round__c[890] ) );
  XOR2_X2 _f_permutation__round__U5137  ( .A(SYNOPSYS_UNCONNECTED_453), .B(
        _f_permutation__round__n2142 ), .Z(_f_permutation__round__c[251] ) );
  XOR2_X2 _f_permutation__round__U5136  ( .A(SYNOPSYS_UNCONNECTED_262), .B(
        _f_permutation__round__n2143 ), .Z(_f_permutation__round__c[826] ) );
  XOR2_X2 _f_permutation__round__U5135  ( .A(SYNOPSYS_UNCONNECTED_133), .B(
        _f_permutation__round__n2142 ), .Z(_f_permutation__round__c[187] ) );
  XOR2_X2 _f_permutation__round__U5134  ( .A(_f_permutation__round_in[1146]), 
        .B(_f_permutation__round__n2143 ), .Z(_f_permutation__round__c[762] )
         );
  XOR2_X2 _f_permutation__round__U5133  ( .A(_f_permutation__round_in[1275]), 
        .B(_f_permutation__round__n2142 ), .Z(_f_permutation__round__c[123] )
         );
  XOR2_X2 _f_permutation__round__U5132  ( .A(_f_permutation__round_in[1466]), 
        .B(_f_permutation__round__n2143 ), .Z(_f_permutation__round__c[698] )
         );
  XOR2_X2 _f_permutation__round__U5131  ( .A(_f_permutation__round__n2145 ), 
        .B(_f_permutation__round__n2144 ), .Z(_f_permutation__round__n2147 )
         );
  XOR2_X2 _f_permutation__round__U5130  ( .A(SYNOPSYS_UNCONNECTED_903), .B(
        _f_permutation__round__n2147 ), .Z(_f_permutation__round__c[953] ) );
  XOR2_X2 _f_permutation__round__U5129  ( .A(SYNOPSYS_UNCONNECTED_774), .B(
        _f_permutation__round__n2146 ), .Z(_f_permutation__round__c[314] ) );
  XOR2_X2 _f_permutation__round__U5128  ( .A(SYNOPSYS_UNCONNECTED_583), .B(
        _f_permutation__round__n2147 ), .Z(_f_permutation__round__c[889] ) );
  XOR2_X2 _f_permutation__round__U5127  ( .A(SYNOPSYS_UNCONNECTED_454), .B(
        _f_permutation__round__n2146 ), .Z(_f_permutation__round__c[250] ) );
  XOR2_X2 _f_permutation__round__U5126  ( .A(SYNOPSYS_UNCONNECTED_263), .B(
        _f_permutation__round__n2147 ), .Z(_f_permutation__round__c[825] ) );
  XOR2_X2 _f_permutation__round__U5125  ( .A(SYNOPSYS_UNCONNECTED_134), .B(
        _f_permutation__round__n2146 ), .Z(_f_permutation__round__c[186] ) );
  XOR2_X2 _f_permutation__round__U5124  ( .A(_f_permutation__round_in[1145]), 
        .B(_f_permutation__round__n2147 ), .Z(_f_permutation__round__c[761] )
         );
  XOR2_X2 _f_permutation__round__U5123  ( .A(_f_permutation__round_in[1274]), 
        .B(_f_permutation__round__n2146 ), .Z(_f_permutation__round__c[122] )
         );
  XOR2_X2 _f_permutation__round__U5122  ( .A(_f_permutation__round_in[1465]), 
        .B(_f_permutation__round__n2147 ), .Z(_f_permutation__round__c[697] )
         );
  XOR2_X2 _f_permutation__round__U5121  ( .A(_f_permutation__round__n2149 ), 
        .B(_f_permutation__round__n2148 ), .Z(_f_permutation__round__n2151 )
         );
  XOR2_X2 _f_permutation__round__U5120  ( .A(SYNOPSYS_UNCONNECTED_904), .B(
        _f_permutation__round__n2151 ), .Z(_f_permutation__round__c[952] ) );
  XOR2_X2 _f_permutation__round__U5119  ( .A(SYNOPSYS_UNCONNECTED_775), .B(
        _f_permutation__round__n2150 ), .Z(_f_permutation__round__c[313] ) );
  XOR2_X2 _f_permutation__round__U5118  ( .A(SYNOPSYS_UNCONNECTED_584), .B(
        _f_permutation__round__n2151 ), .Z(_f_permutation__round__c[888] ) );
  XOR2_X2 _f_permutation__round__U5117  ( .A(SYNOPSYS_UNCONNECTED_455), .B(
        _f_permutation__round__n2150 ), .Z(_f_permutation__round__c[249] ) );
  XOR2_X2 _f_permutation__round__U5116  ( .A(SYNOPSYS_UNCONNECTED_264), .B(
        _f_permutation__round__n2151 ), .Z(_f_permutation__round__c[824] ) );
  XOR2_X2 _f_permutation__round__U5115  ( .A(SYNOPSYS_UNCONNECTED_135), .B(
        _f_permutation__round__n2150 ), .Z(_f_permutation__round__c[185] ) );
  XOR2_X2 _f_permutation__round__U5114  ( .A(_f_permutation__round_in[1144]), 
        .B(_f_permutation__round__n2151 ), .Z(_f_permutation__round__c[760] )
         );
  XOR2_X2 _f_permutation__round__U5113  ( .A(_f_permutation__round_in[1273]), 
        .B(_f_permutation__round__n2150 ), .Z(_f_permutation__round__c[121] )
         );
  XOR2_X2 _f_permutation__round__U5112  ( .A(_f_permutation__round_in[1464]), 
        .B(_f_permutation__round__n2151 ), .Z(_f_permutation__round__c[696] )
         );
  XOR2_X2 _f_permutation__round__U5111  ( .A(_f_permutation__round__n2153 ), 
        .B(_f_permutation__round__n2152 ), .Z(_f_permutation__round__n2155 )
         );
  XOR2_X2 _f_permutation__round__U5110  ( .A(SYNOPSYS_UNCONNECTED_905), .B(
        _f_permutation__round__n2155 ), .Z(_f_permutation__round__c[951] ) );
  XOR2_X2 _f_permutation__round__U5109  ( .A(SYNOPSYS_UNCONNECTED_776), .B(
        _f_permutation__round__n2154 ), .Z(_f_permutation__round__c[312] ) );
  XOR2_X2 _f_permutation__round__U5108  ( .A(SYNOPSYS_UNCONNECTED_585), .B(
        _f_permutation__round__n2155 ), .Z(_f_permutation__round__c[887] ) );
  XOR2_X2 _f_permutation__round__U5107  ( .A(SYNOPSYS_UNCONNECTED_456), .B(
        _f_permutation__round__n2154 ), .Z(_f_permutation__round__c[248] ) );
  XOR2_X2 _f_permutation__round__U5106  ( .A(SYNOPSYS_UNCONNECTED_265), .B(
        _f_permutation__round__n2155 ), .Z(_f_permutation__round__c[823] ) );
  XOR2_X2 _f_permutation__round__U5105  ( .A(SYNOPSYS_UNCONNECTED_136), .B(
        _f_permutation__round__n2154 ), .Z(_f_permutation__round__c[184] ) );
  XOR2_X2 _f_permutation__round__U5104  ( .A(_f_permutation__round_in[1143]), 
        .B(_f_permutation__round__n2155 ), .Z(_f_permutation__round__c[759] )
         );
  XOR2_X2 _f_permutation__round__U5103  ( .A(_f_permutation__round_in[1272]), 
        .B(_f_permutation__round__n2154 ), .Z(_f_permutation__round__c[120] )
         );
  XOR2_X2 _f_permutation__round__U5102  ( .A(_f_permutation__round_in[1463]), 
        .B(_f_permutation__round__n2155 ), .Z(_f_permutation__round__c[695] )
         );
  XOR2_X2 _f_permutation__round__U5101  ( .A(_f_permutation__round__n2157 ), 
        .B(_f_permutation__round__n2156 ), .Z(_f_permutation__round__n2159 )
         );
  XOR2_X2 _f_permutation__round__U5100  ( .A(SYNOPSYS_UNCONNECTED_906), .B(
        _f_permutation__round__n2159 ), .Z(_f_permutation__round__c[950] ) );
  XOR2_X2 _f_permutation__round__U5099  ( .A(SYNOPSYS_UNCONNECTED_777), .B(
        _f_permutation__round__n2158 ), .Z(_f_permutation__round__c[311] ) );
  XOR2_X2 _f_permutation__round__U5098  ( .A(SYNOPSYS_UNCONNECTED_586), .B(
        _f_permutation__round__n2159 ), .Z(_f_permutation__round__c[886] ) );
  XOR2_X2 _f_permutation__round__U5097  ( .A(SYNOPSYS_UNCONNECTED_457), .B(
        _f_permutation__round__n2158 ), .Z(_f_permutation__round__c[247] ) );
  XOR2_X2 _f_permutation__round__U5096  ( .A(SYNOPSYS_UNCONNECTED_266), .B(
        _f_permutation__round__n2159 ), .Z(_f_permutation__round__c[822] ) );
  XOR2_X2 _f_permutation__round__U5095  ( .A(SYNOPSYS_UNCONNECTED_137), .B(
        _f_permutation__round__n2158 ), .Z(_f_permutation__round__c[183] ) );
  XOR2_X2 _f_permutation__round__U5094  ( .A(_f_permutation__round_in[1142]), 
        .B(_f_permutation__round__n2159 ), .Z(_f_permutation__round__c[758] )
         );
  XOR2_X2 _f_permutation__round__U5093  ( .A(_f_permutation__round_in[1271]), 
        .B(_f_permutation__round__n2158 ), .Z(_f_permutation__round__c[119] )
         );
  XOR2_X2 _f_permutation__round__U5092  ( .A(_f_permutation__round_in[1462]), 
        .B(_f_permutation__round__n2159 ), .Z(_f_permutation__round__c[694] )
         );
  XOR2_X2 _f_permutation__round__U5091  ( .A(_f_permutation__round__n2161 ), 
        .B(_f_permutation__round__n2160 ), .Z(_f_permutation__round__n2163 )
         );
  XOR2_X2 _f_permutation__round__U5090  ( .A(SYNOPSYS_UNCONNECTED_907), .B(
        _f_permutation__round__n2163 ), .Z(_f_permutation__round__c[949] ) );
  XOR2_X2 _f_permutation__round__U5089  ( .A(SYNOPSYS_UNCONNECTED_778), .B(
        _f_permutation__round__n2162 ), .Z(_f_permutation__round__c[310] ) );
  XOR2_X2 _f_permutation__round__U5088  ( .A(SYNOPSYS_UNCONNECTED_587), .B(
        _f_permutation__round__n2163 ), .Z(_f_permutation__round__c[885] ) );
  XOR2_X2 _f_permutation__round__U5087  ( .A(SYNOPSYS_UNCONNECTED_458), .B(
        _f_permutation__round__n2162 ), .Z(_f_permutation__round__c[246] ) );
  XOR2_X2 _f_permutation__round__U5086  ( .A(SYNOPSYS_UNCONNECTED_267), .B(
        _f_permutation__round__n2163 ), .Z(_f_permutation__round__c[821] ) );
  XOR2_X2 _f_permutation__round__U5085  ( .A(SYNOPSYS_UNCONNECTED_138), .B(
        _f_permutation__round__n2162 ), .Z(_f_permutation__round__c[182] ) );
  XOR2_X2 _f_permutation__round__U5084  ( .A(_f_permutation__round_in[1141]), 
        .B(_f_permutation__round__n2163 ), .Z(_f_permutation__round__c[757] )
         );
  XOR2_X2 _f_permutation__round__U5083  ( .A(_f_permutation__round_in[1270]), 
        .B(_f_permutation__round__n2162 ), .Z(_f_permutation__round__c[118] )
         );
  XOR2_X2 _f_permutation__round__U5082  ( .A(_f_permutation__round_in[1461]), 
        .B(_f_permutation__round__n2163 ), .Z(_f_permutation__round__c[693] )
         );
  XOR2_X2 _f_permutation__round__U5081  ( .A(_f_permutation__round__n2165 ), 
        .B(_f_permutation__round__n2164 ), .Z(_f_permutation__round__n2167 )
         );
  XOR2_X2 _f_permutation__round__U5080  ( .A(SYNOPSYS_UNCONNECTED_908), .B(
        _f_permutation__round__n2167 ), .Z(_f_permutation__round__c[948] ) );
  XOR2_X2 _f_permutation__round__U5079  ( .A(SYNOPSYS_UNCONNECTED_779), .B(
        _f_permutation__round__n2166 ), .Z(_f_permutation__round__c[309] ) );
  XOR2_X2 _f_permutation__round__U5078  ( .A(SYNOPSYS_UNCONNECTED_588), .B(
        _f_permutation__round__n2167 ), .Z(_f_permutation__round__c[884] ) );
  XOR2_X2 _f_permutation__round__U5077  ( .A(SYNOPSYS_UNCONNECTED_459), .B(
        _f_permutation__round__n2166 ), .Z(_f_permutation__round__c[245] ) );
  XOR2_X2 _f_permutation__round__U5076  ( .A(SYNOPSYS_UNCONNECTED_268), .B(
        _f_permutation__round__n2167 ), .Z(_f_permutation__round__c[820] ) );
  XOR2_X2 _f_permutation__round__U5075  ( .A(SYNOPSYS_UNCONNECTED_139), .B(
        _f_permutation__round__n2166 ), .Z(_f_permutation__round__c[181] ) );
  XOR2_X2 _f_permutation__round__U5074  ( .A(_f_permutation__round_in[1140]), 
        .B(_f_permutation__round__n2167 ), .Z(_f_permutation__round__c[756] )
         );
  XOR2_X2 _f_permutation__round__U5073  ( .A(_f_permutation__round_in[1269]), 
        .B(_f_permutation__round__n2166 ), .Z(_f_permutation__round__c[117] )
         );
  XOR2_X2 _f_permutation__round__U5072  ( .A(_f_permutation__round_in[1460]), 
        .B(_f_permutation__round__n2167 ), .Z(_f_permutation__round__c[692] )
         );
  XOR2_X2 _f_permutation__round__U5071  ( .A(_f_permutation__round__n2169 ), 
        .B(_f_permutation__round__n2168 ), .Z(_f_permutation__round__n2171 )
         );
  XOR2_X2 _f_permutation__round__U5070  ( .A(SYNOPSYS_UNCONNECTED_909), .B(
        _f_permutation__round__n2171 ), .Z(_f_permutation__round__c[947] ) );
  XOR2_X2 _f_permutation__round__U5069  ( .A(SYNOPSYS_UNCONNECTED_780), .B(
        _f_permutation__round__n2170 ), .Z(_f_permutation__round__c[308] ) );
  XOR2_X2 _f_permutation__round__U5068  ( .A(SYNOPSYS_UNCONNECTED_589), .B(
        _f_permutation__round__n2171 ), .Z(_f_permutation__round__c[883] ) );
  XOR2_X2 _f_permutation__round__U5067  ( .A(SYNOPSYS_UNCONNECTED_460), .B(
        _f_permutation__round__n2170 ), .Z(_f_permutation__round__c[244] ) );
  XOR2_X2 _f_permutation__round__U5066  ( .A(SYNOPSYS_UNCONNECTED_269), .B(
        _f_permutation__round__n2171 ), .Z(_f_permutation__round__c[819] ) );
  XOR2_X2 _f_permutation__round__U5065  ( .A(SYNOPSYS_UNCONNECTED_140), .B(
        _f_permutation__round__n2170 ), .Z(_f_permutation__round__c[180] ) );
  XOR2_X2 _f_permutation__round__U5064  ( .A(_f_permutation__round_in[1139]), 
        .B(_f_permutation__round__n2171 ), .Z(_f_permutation__round__c[755] )
         );
  XOR2_X2 _f_permutation__round__U5063  ( .A(_f_permutation__round_in[1268]), 
        .B(_f_permutation__round__n2170 ), .Z(_f_permutation__round__c[116] )
         );
  XOR2_X2 _f_permutation__round__U5062  ( .A(_f_permutation__round_in[1459]), 
        .B(_f_permutation__round__n2171 ), .Z(_f_permutation__round__c[691] )
         );
  XOR2_X2 _f_permutation__round__U5061  ( .A(_f_permutation__round__n2173 ), 
        .B(_f_permutation__round__n2172 ), .Z(_f_permutation__round__n2175 )
         );
  XOR2_X2 _f_permutation__round__U5060  ( .A(SYNOPSYS_UNCONNECTED_910), .B(
        _f_permutation__round__n2175 ), .Z(_f_permutation__round__c[946] ) );
  XOR2_X2 _f_permutation__round__U5059  ( .A(SYNOPSYS_UNCONNECTED_781), .B(
        _f_permutation__round__n2174 ), .Z(_f_permutation__round__c[307] ) );
  XOR2_X2 _f_permutation__round__U5058  ( .A(SYNOPSYS_UNCONNECTED_590), .B(
        _f_permutation__round__n2175 ), .Z(_f_permutation__round__c[882] ) );
  XOR2_X2 _f_permutation__round__U5057  ( .A(SYNOPSYS_UNCONNECTED_461), .B(
        _f_permutation__round__n2174 ), .Z(_f_permutation__round__c[243] ) );
  XOR2_X2 _f_permutation__round__U5056  ( .A(SYNOPSYS_UNCONNECTED_270), .B(
        _f_permutation__round__n2175 ), .Z(_f_permutation__round__c[818] ) );
  XOR2_X2 _f_permutation__round__U5055  ( .A(SYNOPSYS_UNCONNECTED_141), .B(
        _f_permutation__round__n2174 ), .Z(_f_permutation__round__c[179] ) );
  XOR2_X2 _f_permutation__round__U5054  ( .A(_f_permutation__round_in[1138]), 
        .B(_f_permutation__round__n2175 ), .Z(_f_permutation__round__c[754] )
         );
  XOR2_X2 _f_permutation__round__U5053  ( .A(_f_permutation__round_in[1267]), 
        .B(_f_permutation__round__n2174 ), .Z(_f_permutation__round__c[115] )
         );
  XOR2_X2 _f_permutation__round__U5052  ( .A(_f_permutation__round_in[1458]), 
        .B(_f_permutation__round__n2175 ), .Z(_f_permutation__round__c[690] )
         );
  XOR2_X2 _f_permutation__round__U5051  ( .A(_f_permutation__round__n2177 ), 
        .B(_f_permutation__round__n2176 ), .Z(_f_permutation__round__n2179 )
         );
  XOR2_X2 _f_permutation__round__U5050  ( .A(SYNOPSYS_UNCONNECTED_911), .B(
        _f_permutation__round__n2179 ), .Z(_f_permutation__round__c[945] ) );
  XOR2_X2 _f_permutation__round__U5049  ( .A(SYNOPSYS_UNCONNECTED_782), .B(
        _f_permutation__round__n2178 ), .Z(_f_permutation__round__c[306] ) );
  XOR2_X2 _f_permutation__round__U5048  ( .A(SYNOPSYS_UNCONNECTED_591), .B(
        _f_permutation__round__n2179 ), .Z(_f_permutation__round__c[881] ) );
  XOR2_X2 _f_permutation__round__U5047  ( .A(SYNOPSYS_UNCONNECTED_462), .B(
        _f_permutation__round__n2178 ), .Z(_f_permutation__round__c[242] ) );
  XOR2_X2 _f_permutation__round__U5046  ( .A(SYNOPSYS_UNCONNECTED_271), .B(
        _f_permutation__round__n2179 ), .Z(_f_permutation__round__c[817] ) );
  XOR2_X2 _f_permutation__round__U5045  ( .A(SYNOPSYS_UNCONNECTED_142), .B(
        _f_permutation__round__n2178 ), .Z(_f_permutation__round__c[178] ) );
  XOR2_X2 _f_permutation__round__U5044  ( .A(_f_permutation__round_in[1137]), 
        .B(_f_permutation__round__n2179 ), .Z(_f_permutation__round__c[753] )
         );
  XOR2_X2 _f_permutation__round__U5043  ( .A(_f_permutation__round_in[1266]), 
        .B(_f_permutation__round__n2178 ), .Z(_f_permutation__round__c[114] )
         );
  XOR2_X2 _f_permutation__round__U5042  ( .A(_f_permutation__round_in[1457]), 
        .B(_f_permutation__round__n2179 ), .Z(_f_permutation__round__c[689] )
         );
  XOR2_X2 _f_permutation__round__U5041  ( .A(_f_permutation__round__n2181 ), 
        .B(_f_permutation__round__n2180 ), .Z(_f_permutation__round__n2183 )
         );
  XOR2_X2 _f_permutation__round__U5040  ( .A(SYNOPSYS_UNCONNECTED_912), .B(
        _f_permutation__round__n2183 ), .Z(_f_permutation__round__c[944] ) );
  XOR2_X2 _f_permutation__round__U5039  ( .A(SYNOPSYS_UNCONNECTED_783), .B(
        _f_permutation__round__n2182 ), .Z(_f_permutation__round__c[305] ) );
  XOR2_X2 _f_permutation__round__U5038  ( .A(SYNOPSYS_UNCONNECTED_592), .B(
        _f_permutation__round__n2183 ), .Z(_f_permutation__round__c[880] ) );
  XOR2_X2 _f_permutation__round__U5037  ( .A(SYNOPSYS_UNCONNECTED_463), .B(
        _f_permutation__round__n2182 ), .Z(_f_permutation__round__c[241] ) );
  XOR2_X2 _f_permutation__round__U5036  ( .A(SYNOPSYS_UNCONNECTED_272), .B(
        _f_permutation__round__n2183 ), .Z(_f_permutation__round__c[816] ) );
  XOR2_X2 _f_permutation__round__U5035  ( .A(SYNOPSYS_UNCONNECTED_143), .B(
        _f_permutation__round__n2182 ), .Z(_f_permutation__round__c[177] ) );
  XOR2_X2 _f_permutation__round__U5034  ( .A(_f_permutation__round_in[1136]), 
        .B(_f_permutation__round__n2183 ), .Z(_f_permutation__round__c[752] )
         );
  XOR2_X2 _f_permutation__round__U5033  ( .A(_f_permutation__round_in[1265]), 
        .B(_f_permutation__round__n2182 ), .Z(_f_permutation__round__c[113] )
         );
  XOR2_X2 _f_permutation__round__U5032  ( .A(_f_permutation__round_in[1456]), 
        .B(_f_permutation__round__n2183 ), .Z(_f_permutation__round__c[688] )
         );
  XOR2_X2 _f_permutation__round__U5031  ( .A(_f_permutation__round__n2185 ), 
        .B(_f_permutation__round__n2184 ), .Z(_f_permutation__round__n2187 )
         );
  XOR2_X2 _f_permutation__round__U5030  ( .A(SYNOPSYS_UNCONNECTED_913), .B(
        _f_permutation__round__n2187 ), .Z(_f_permutation__round__c[943] ) );
  XOR2_X2 _f_permutation__round__U5029  ( .A(SYNOPSYS_UNCONNECTED_784), .B(
        _f_permutation__round__n2186 ), .Z(_f_permutation__round__c[304] ) );
  XOR2_X2 _f_permutation__round__U5028  ( .A(SYNOPSYS_UNCONNECTED_593), .B(
        _f_permutation__round__n2187 ), .Z(_f_permutation__round__c[879] ) );
  XOR2_X2 _f_permutation__round__U5027  ( .A(SYNOPSYS_UNCONNECTED_464), .B(
        _f_permutation__round__n2186 ), .Z(_f_permutation__round__c[240] ) );
  XOR2_X2 _f_permutation__round__U5026  ( .A(SYNOPSYS_UNCONNECTED_273), .B(
        _f_permutation__round__n2187 ), .Z(_f_permutation__round__c[815] ) );
  XOR2_X2 _f_permutation__round__U5025  ( .A(SYNOPSYS_UNCONNECTED_144), .B(
        _f_permutation__round__n2186 ), .Z(_f_permutation__round__c[176] ) );
  XOR2_X2 _f_permutation__round__U5024  ( .A(_f_permutation__round_in[1135]), 
        .B(_f_permutation__round__n2187 ), .Z(_f_permutation__round__c[751] )
         );
  XOR2_X2 _f_permutation__round__U5023  ( .A(_f_permutation__round_in[1264]), 
        .B(_f_permutation__round__n2186 ), .Z(_f_permutation__round__c[112] )
         );
  XOR2_X2 _f_permutation__round__U5022  ( .A(_f_permutation__round_in[1455]), 
        .B(_f_permutation__round__n2187 ), .Z(_f_permutation__round__c[687] )
         );
  XOR2_X2 _f_permutation__round__U5021  ( .A(_f_permutation__round__n2189 ), 
        .B(_f_permutation__round__n2188 ), .Z(_f_permutation__round__n2191 )
         );
  XOR2_X2 _f_permutation__round__U5020  ( .A(SYNOPSYS_UNCONNECTED_914), .B(
        _f_permutation__round__n2191 ), .Z(_f_permutation__round__c[942] ) );
  XOR2_X2 _f_permutation__round__U5019  ( .A(SYNOPSYS_UNCONNECTED_785), .B(
        _f_permutation__round__n2190 ), .Z(_f_permutation__round__c[303] ) );
  XOR2_X2 _f_permutation__round__U5018  ( .A(SYNOPSYS_UNCONNECTED_594), .B(
        _f_permutation__round__n2191 ), .Z(_f_permutation__round__c[878] ) );
  XOR2_X2 _f_permutation__round__U5017  ( .A(SYNOPSYS_UNCONNECTED_465), .B(
        _f_permutation__round__n2190 ), .Z(_f_permutation__round__c[239] ) );
  XOR2_X2 _f_permutation__round__U5016  ( .A(SYNOPSYS_UNCONNECTED_274), .B(
        _f_permutation__round__n2191 ), .Z(_f_permutation__round__c[814] ) );
  XOR2_X2 _f_permutation__round__U5015  ( .A(SYNOPSYS_UNCONNECTED_145), .B(
        _f_permutation__round__n2190 ), .Z(_f_permutation__round__c[175] ) );
  XOR2_X2 _f_permutation__round__U5014  ( .A(_f_permutation__round_in[1134]), 
        .B(_f_permutation__round__n2191 ), .Z(_f_permutation__round__c[750] )
         );
  XOR2_X2 _f_permutation__round__U5013  ( .A(_f_permutation__round_in[1263]), 
        .B(_f_permutation__round__n2190 ), .Z(_f_permutation__round__c[111] )
         );
  XOR2_X2 _f_permutation__round__U5012  ( .A(_f_permutation__round_in[1454]), 
        .B(_f_permutation__round__n2191 ), .Z(_f_permutation__round__c[686] )
         );
  XOR2_X2 _f_permutation__round__U5011  ( .A(_f_permutation__round__n2193 ), 
        .B(_f_permutation__round__n2192 ), .Z(_f_permutation__round__n2195 )
         );
  XOR2_X2 _f_permutation__round__U5010  ( .A(SYNOPSYS_UNCONNECTED_915), .B(
        _f_permutation__round__n2195 ), .Z(_f_permutation__round__c[941] ) );
  XOR2_X2 _f_permutation__round__U5009  ( .A(SYNOPSYS_UNCONNECTED_786), .B(
        _f_permutation__round__n2194 ), .Z(_f_permutation__round__c[302] ) );
  XOR2_X2 _f_permutation__round__U5008  ( .A(SYNOPSYS_UNCONNECTED_595), .B(
        _f_permutation__round__n2195 ), .Z(_f_permutation__round__c[877] ) );
  XOR2_X2 _f_permutation__round__U5007  ( .A(SYNOPSYS_UNCONNECTED_466), .B(
        _f_permutation__round__n2194 ), .Z(_f_permutation__round__c[238] ) );
  XOR2_X2 _f_permutation__round__U5006  ( .A(SYNOPSYS_UNCONNECTED_275), .B(
        _f_permutation__round__n2195 ), .Z(_f_permutation__round__c[813] ) );
  XOR2_X2 _f_permutation__round__U5005  ( .A(SYNOPSYS_UNCONNECTED_146), .B(
        _f_permutation__round__n2194 ), .Z(_f_permutation__round__c[174] ) );
  XOR2_X2 _f_permutation__round__U5004  ( .A(_f_permutation__round_in[1133]), 
        .B(_f_permutation__round__n2195 ), .Z(_f_permutation__round__c[749] )
         );
  XOR2_X2 _f_permutation__round__U5003  ( .A(_f_permutation__round_in[1262]), 
        .B(_f_permutation__round__n2194 ), .Z(_f_permutation__round__c[110] )
         );
  XOR2_X2 _f_permutation__round__U5002  ( .A(_f_permutation__round_in[1453]), 
        .B(_f_permutation__round__n2195 ), .Z(_f_permutation__round__c[685] )
         );
  XOR2_X2 _f_permutation__round__U5001  ( .A(_f_permutation__round__n2197 ), 
        .B(_f_permutation__round__n2196 ), .Z(_f_permutation__round__n2199 )
         );
  XOR2_X2 _f_permutation__round__U5000  ( .A(SYNOPSYS_UNCONNECTED_916), .B(
        _f_permutation__round__n2199 ), .Z(_f_permutation__round__c[940] ) );
  XOR2_X2 _f_permutation__round__U4999  ( .A(SYNOPSYS_UNCONNECTED_787), .B(
        _f_permutation__round__n2198 ), .Z(_f_permutation__round__c[301] ) );
  XOR2_X2 _f_permutation__round__U4998  ( .A(SYNOPSYS_UNCONNECTED_596), .B(
        _f_permutation__round__n2199 ), .Z(_f_permutation__round__c[876] ) );
  XOR2_X2 _f_permutation__round__U4997  ( .A(SYNOPSYS_UNCONNECTED_467), .B(
        _f_permutation__round__n2198 ), .Z(_f_permutation__round__c[237] ) );
  XOR2_X2 _f_permutation__round__U4996  ( .A(SYNOPSYS_UNCONNECTED_276), .B(
        _f_permutation__round__n2199 ), .Z(_f_permutation__round__c[812] ) );
  XOR2_X2 _f_permutation__round__U4995  ( .A(SYNOPSYS_UNCONNECTED_147), .B(
        _f_permutation__round__n2198 ), .Z(_f_permutation__round__c[173] ) );
  XOR2_X2 _f_permutation__round__U4994  ( .A(_f_permutation__round_in[1132]), 
        .B(_f_permutation__round__n2199 ), .Z(_f_permutation__round__c[748] )
         );
  XOR2_X2 _f_permutation__round__U4993  ( .A(_f_permutation__round_in[1261]), 
        .B(_f_permutation__round__n2198 ), .Z(_f_permutation__round__c[109] )
         );
  XOR2_X2 _f_permutation__round__U4992  ( .A(_f_permutation__round_in[1452]), 
        .B(_f_permutation__round__n2199 ), .Z(_f_permutation__round__c[684] )
         );
  XOR2_X2 _f_permutation__round__U4991  ( .A(_f_permutation__round__n2201 ), 
        .B(_f_permutation__round__n2200 ), .Z(_f_permutation__round__n2203 )
         );
  XOR2_X2 _f_permutation__round__U4990  ( .A(SYNOPSYS_UNCONNECTED_917), .B(
        _f_permutation__round__n2203 ), .Z(_f_permutation__round__c[939] ) );
  XOR2_X2 _f_permutation__round__U4989  ( .A(SYNOPSYS_UNCONNECTED_788), .B(
        _f_permutation__round__n2202 ), .Z(_f_permutation__round__c[300] ) );
  XOR2_X2 _f_permutation__round__U4988  ( .A(SYNOPSYS_UNCONNECTED_597), .B(
        _f_permutation__round__n2203 ), .Z(_f_permutation__round__c[875] ) );
  XOR2_X2 _f_permutation__round__U4987  ( .A(SYNOPSYS_UNCONNECTED_468), .B(
        _f_permutation__round__n2202 ), .Z(_f_permutation__round__c[236] ) );
  XOR2_X2 _f_permutation__round__U4986  ( .A(SYNOPSYS_UNCONNECTED_277), .B(
        _f_permutation__round__n2203 ), .Z(_f_permutation__round__c[811] ) );
  XOR2_X2 _f_permutation__round__U4985  ( .A(SYNOPSYS_UNCONNECTED_148), .B(
        _f_permutation__round__n2202 ), .Z(_f_permutation__round__c[172] ) );
  XOR2_X2 _f_permutation__round__U4984  ( .A(_f_permutation__round_in[1131]), 
        .B(_f_permutation__round__n2203 ), .Z(_f_permutation__round__c[747] )
         );
  XOR2_X2 _f_permutation__round__U4983  ( .A(_f_permutation__round_in[1260]), 
        .B(_f_permutation__round__n2202 ), .Z(_f_permutation__round__c[108] )
         );
  XOR2_X2 _f_permutation__round__U4982  ( .A(_f_permutation__round_in[1451]), 
        .B(_f_permutation__round__n2203 ), .Z(_f_permutation__round__c[683] )
         );
  XOR2_X2 _f_permutation__round__U4981  ( .A(_f_permutation__round__n2205 ), 
        .B(_f_permutation__round__n2204 ), .Z(_f_permutation__round__n2207 )
         );
  XOR2_X2 _f_permutation__round__U4980  ( .A(SYNOPSYS_UNCONNECTED_918), .B(
        _f_permutation__round__n2207 ), .Z(_f_permutation__round__c[938] ) );
  XOR2_X2 _f_permutation__round__U4979  ( .A(SYNOPSYS_UNCONNECTED_789), .B(
        _f_permutation__round__n2206 ), .Z(_f_permutation__round__c[299] ) );
  XOR2_X2 _f_permutation__round__U4978  ( .A(SYNOPSYS_UNCONNECTED_598), .B(
        _f_permutation__round__n2207 ), .Z(_f_permutation__round__c[874] ) );
  XOR2_X2 _f_permutation__round__U4977  ( .A(SYNOPSYS_UNCONNECTED_469), .B(
        _f_permutation__round__n2206 ), .Z(_f_permutation__round__c[235] ) );
  XOR2_X2 _f_permutation__round__U4976  ( .A(SYNOPSYS_UNCONNECTED_278), .B(
        _f_permutation__round__n2207 ), .Z(_f_permutation__round__c[810] ) );
  XOR2_X2 _f_permutation__round__U4975  ( .A(SYNOPSYS_UNCONNECTED_149), .B(
        _f_permutation__round__n2206 ), .Z(_f_permutation__round__c[171] ) );
  XOR2_X2 _f_permutation__round__U4974  ( .A(_f_permutation__round_in[1130]), 
        .B(_f_permutation__round__n2207 ), .Z(_f_permutation__round__c[746] )
         );
  XOR2_X2 _f_permutation__round__U4973  ( .A(_f_permutation__round_in[1259]), 
        .B(_f_permutation__round__n2206 ), .Z(_f_permutation__round__c[107] )
         );
  XOR2_X2 _f_permutation__round__U4972  ( .A(_f_permutation__round_in[1450]), 
        .B(_f_permutation__round__n2207 ), .Z(_f_permutation__round__c[682] )
         );
  XOR2_X2 _f_permutation__round__U4971  ( .A(_f_permutation__round__n2209 ), 
        .B(_f_permutation__round__n2208 ), .Z(_f_permutation__round__n2211 )
         );
  XOR2_X2 _f_permutation__round__U4970  ( .A(SYNOPSYS_UNCONNECTED_919), .B(
        _f_permutation__round__n2211 ), .Z(_f_permutation__round__c[937] ) );
  XOR2_X2 _f_permutation__round__U4969  ( .A(SYNOPSYS_UNCONNECTED_790), .B(
        _f_permutation__round__n2210 ), .Z(_f_permutation__round__c[298] ) );
  XOR2_X2 _f_permutation__round__U4968  ( .A(SYNOPSYS_UNCONNECTED_599), .B(
        _f_permutation__round__n2211 ), .Z(_f_permutation__round__c[873] ) );
  XOR2_X2 _f_permutation__round__U4967  ( .A(SYNOPSYS_UNCONNECTED_470), .B(
        _f_permutation__round__n2210 ), .Z(_f_permutation__round__c[234] ) );
  XOR2_X2 _f_permutation__round__U4966  ( .A(SYNOPSYS_UNCONNECTED_279), .B(
        _f_permutation__round__n2211 ), .Z(_f_permutation__round__c[809] ) );
  XOR2_X2 _f_permutation__round__U4965  ( .A(SYNOPSYS_UNCONNECTED_150), .B(
        _f_permutation__round__n2210 ), .Z(_f_permutation__round__c[170] ) );
  XOR2_X2 _f_permutation__round__U4964  ( .A(_f_permutation__round_in[1129]), 
        .B(_f_permutation__round__n2211 ), .Z(_f_permutation__round__c[745] )
         );
  XOR2_X2 _f_permutation__round__U4963  ( .A(_f_permutation__round_in[1258]), 
        .B(_f_permutation__round__n2210 ), .Z(_f_permutation__round__c[106] )
         );
  XOR2_X2 _f_permutation__round__U4962  ( .A(_f_permutation__round_in[1449]), 
        .B(_f_permutation__round__n2211 ), .Z(_f_permutation__round__c[681] )
         );
  XOR2_X2 _f_permutation__round__U4961  ( .A(_f_permutation__round__n2213 ), 
        .B(_f_permutation__round__n2212 ), .Z(_f_permutation__round__n2215 )
         );
  XOR2_X2 _f_permutation__round__U4960  ( .A(SYNOPSYS_UNCONNECTED_920), .B(
        _f_permutation__round__n2215 ), .Z(_f_permutation__round__c[936] ) );
  XOR2_X2 _f_permutation__round__U4959  ( .A(SYNOPSYS_UNCONNECTED_791), .B(
        _f_permutation__round__n2214 ), .Z(_f_permutation__round__c[297] ) );
  XOR2_X2 _f_permutation__round__U4958  ( .A(SYNOPSYS_UNCONNECTED_600), .B(
        _f_permutation__round__n2215 ), .Z(_f_permutation__round__c[872] ) );
  XOR2_X2 _f_permutation__round__U4957  ( .A(SYNOPSYS_UNCONNECTED_471), .B(
        _f_permutation__round__n2214 ), .Z(_f_permutation__round__c[233] ) );
  XOR2_X2 _f_permutation__round__U4956  ( .A(SYNOPSYS_UNCONNECTED_280), .B(
        _f_permutation__round__n2215 ), .Z(_f_permutation__round__c[808] ) );
  XOR2_X2 _f_permutation__round__U4955  ( .A(SYNOPSYS_UNCONNECTED_151), .B(
        _f_permutation__round__n2214 ), .Z(_f_permutation__round__c[169] ) );
  XOR2_X2 _f_permutation__round__U4954  ( .A(_f_permutation__round_in[1128]), 
        .B(_f_permutation__round__n2215 ), .Z(_f_permutation__round__c[744] )
         );
  XOR2_X2 _f_permutation__round__U4953  ( .A(_f_permutation__round_in[1257]), 
        .B(_f_permutation__round__n2214 ), .Z(_f_permutation__round__c[105] )
         );
  XOR2_X2 _f_permutation__round__U4952  ( .A(_f_permutation__round_in[1448]), 
        .B(_f_permutation__round__n2215 ), .Z(_f_permutation__round__c[680] )
         );
  XOR2_X2 _f_permutation__round__U4951  ( .A(_f_permutation__round__n2217 ), 
        .B(_f_permutation__round__n2216 ), .Z(_f_permutation__round__n2219 )
         );
  XOR2_X2 _f_permutation__round__U4950  ( .A(SYNOPSYS_UNCONNECTED_921), .B(
        _f_permutation__round__n2219 ), .Z(_f_permutation__round__c[935] ) );
  XOR2_X2 _f_permutation__round__U4949  ( .A(SYNOPSYS_UNCONNECTED_792), .B(
        _f_permutation__round__n2218 ), .Z(_f_permutation__round__c[296] ) );
  XOR2_X2 _f_permutation__round__U4948  ( .A(SYNOPSYS_UNCONNECTED_601), .B(
        _f_permutation__round__n2219 ), .Z(_f_permutation__round__c[871] ) );
  XOR2_X2 _f_permutation__round__U4947  ( .A(SYNOPSYS_UNCONNECTED_472), .B(
        _f_permutation__round__n2218 ), .Z(_f_permutation__round__c[232] ) );
  XOR2_X2 _f_permutation__round__U4946  ( .A(SYNOPSYS_UNCONNECTED_281), .B(
        _f_permutation__round__n2219 ), .Z(_f_permutation__round__c[807] ) );
  XOR2_X2 _f_permutation__round__U4945  ( .A(SYNOPSYS_UNCONNECTED_152), .B(
        _f_permutation__round__n2218 ), .Z(_f_permutation__round__c[168] ) );
  XOR2_X2 _f_permutation__round__U4944  ( .A(_f_permutation__round_in[1127]), 
        .B(_f_permutation__round__n2219 ), .Z(_f_permutation__round__c[743] )
         );
  XOR2_X2 _f_permutation__round__U4943  ( .A(_f_permutation__round_in[1256]), 
        .B(_f_permutation__round__n2218 ), .Z(_f_permutation__round__c[104] )
         );
  XOR2_X2 _f_permutation__round__U4942  ( .A(_f_permutation__round_in[1447]), 
        .B(_f_permutation__round__n2219 ), .Z(_f_permutation__round__c[679] )
         );
  XOR2_X2 _f_permutation__round__U4941  ( .A(_f_permutation__round__n2221 ), 
        .B(_f_permutation__round__n2220 ), .Z(_f_permutation__round__n2223 )
         );
  XOR2_X2 _f_permutation__round__U4940  ( .A(SYNOPSYS_UNCONNECTED_922), .B(
        _f_permutation__round__n2223 ), .Z(_f_permutation__round__c[934] ) );
  XOR2_X2 _f_permutation__round__U4939  ( .A(SYNOPSYS_UNCONNECTED_793), .B(
        _f_permutation__round__n2222 ), .Z(_f_permutation__round__c[295] ) );
  XOR2_X2 _f_permutation__round__U4938  ( .A(SYNOPSYS_UNCONNECTED_602), .B(
        _f_permutation__round__n2223 ), .Z(_f_permutation__round__c[870] ) );
  XOR2_X2 _f_permutation__round__U4937  ( .A(SYNOPSYS_UNCONNECTED_473), .B(
        _f_permutation__round__n2222 ), .Z(_f_permutation__round__c[231] ) );
  XOR2_X2 _f_permutation__round__U4936  ( .A(SYNOPSYS_UNCONNECTED_282), .B(
        _f_permutation__round__n2223 ), .Z(_f_permutation__round__c[806] ) );
  XOR2_X2 _f_permutation__round__U4935  ( .A(SYNOPSYS_UNCONNECTED_153), .B(
        _f_permutation__round__n2222 ), .Z(_f_permutation__round__c[167] ) );
  XOR2_X2 _f_permutation__round__U4934  ( .A(_f_permutation__round_in[1126]), 
        .B(_f_permutation__round__n2223 ), .Z(_f_permutation__round__c[742] )
         );
  XOR2_X2 _f_permutation__round__U4933  ( .A(_f_permutation__round_in[1255]), 
        .B(_f_permutation__round__n2222 ), .Z(_f_permutation__round__c[103] )
         );
  XOR2_X2 _f_permutation__round__U4932  ( .A(_f_permutation__round_in[1446]), 
        .B(_f_permutation__round__n2223 ), .Z(_f_permutation__round__c[678] )
         );
  XOR2_X2 _f_permutation__round__U4931  ( .A(_f_permutation__round__n2225 ), 
        .B(_f_permutation__round__n2224 ), .Z(_f_permutation__round__n2227 )
         );
  XOR2_X2 _f_permutation__round__U4930  ( .A(SYNOPSYS_UNCONNECTED_923), .B(
        _f_permutation__round__n2227 ), .Z(_f_permutation__round__c[933] ) );
  XOR2_X2 _f_permutation__round__U4929  ( .A(SYNOPSYS_UNCONNECTED_794), .B(
        _f_permutation__round__n2226 ), .Z(_f_permutation__round__c[294] ) );
  XOR2_X2 _f_permutation__round__U4928  ( .A(SYNOPSYS_UNCONNECTED_603), .B(
        _f_permutation__round__n2227 ), .Z(_f_permutation__round__c[869] ) );
  XOR2_X2 _f_permutation__round__U4927  ( .A(SYNOPSYS_UNCONNECTED_474), .B(
        _f_permutation__round__n2226 ), .Z(_f_permutation__round__c[230] ) );
  XOR2_X2 _f_permutation__round__U4926  ( .A(SYNOPSYS_UNCONNECTED_283), .B(
        _f_permutation__round__n2227 ), .Z(_f_permutation__round__c[805] ) );
  XOR2_X2 _f_permutation__round__U4925  ( .A(SYNOPSYS_UNCONNECTED_154), .B(
        _f_permutation__round__n2226 ), .Z(_f_permutation__round__c[166] ) );
  XOR2_X2 _f_permutation__round__U4924  ( .A(_f_permutation__round_in[1125]), 
        .B(_f_permutation__round__n2227 ), .Z(_f_permutation__round__c[741] )
         );
  XOR2_X2 _f_permutation__round__U4923  ( .A(_f_permutation__round_in[1254]), 
        .B(_f_permutation__round__n2226 ), .Z(_f_permutation__round__c[102] )
         );
  XOR2_X2 _f_permutation__round__U4922  ( .A(_f_permutation__round_in[1445]), 
        .B(_f_permutation__round__n2227 ), .Z(_f_permutation__round__c[677] )
         );
  XOR2_X2 _f_permutation__round__U4921  ( .A(_f_permutation__round__n2229 ), 
        .B(_f_permutation__round__n2228 ), .Z(_f_permutation__round__n2231 )
         );
  XOR2_X2 _f_permutation__round__U4920  ( .A(SYNOPSYS_UNCONNECTED_924), .B(
        _f_permutation__round__n2231 ), .Z(_f_permutation__round__c[932] ) );
  XOR2_X2 _f_permutation__round__U4919  ( .A(SYNOPSYS_UNCONNECTED_795), .B(
        _f_permutation__round__n2230 ), .Z(_f_permutation__round__c[293] ) );
  XOR2_X2 _f_permutation__round__U4918  ( .A(SYNOPSYS_UNCONNECTED_604), .B(
        _f_permutation__round__n2231 ), .Z(_f_permutation__round__c[868] ) );
  XOR2_X2 _f_permutation__round__U4917  ( .A(SYNOPSYS_UNCONNECTED_475), .B(
        _f_permutation__round__n2230 ), .Z(_f_permutation__round__c[229] ) );
  XOR2_X2 _f_permutation__round__U4916  ( .A(SYNOPSYS_UNCONNECTED_284), .B(
        _f_permutation__round__n2231 ), .Z(_f_permutation__round__c[804] ) );
  XOR2_X2 _f_permutation__round__U4915  ( .A(SYNOPSYS_UNCONNECTED_155), .B(
        _f_permutation__round__n2230 ), .Z(_f_permutation__round__c[165] ) );
  XOR2_X2 _f_permutation__round__U4914  ( .A(_f_permutation__round_in[1124]), 
        .B(_f_permutation__round__n2231 ), .Z(_f_permutation__round__c[740] )
         );
  XOR2_X2 _f_permutation__round__U4913  ( .A(_f_permutation__round_in[1253]), 
        .B(_f_permutation__round__n2230 ), .Z(_f_permutation__round__c[101] )
         );
  XOR2_X2 _f_permutation__round__U4912  ( .A(_f_permutation__round_in[1444]), 
        .B(_f_permutation__round__n2231 ), .Z(_f_permutation__round__c[676] )
         );
  XOR2_X2 _f_permutation__round__U4911  ( .A(_f_permutation__round__n2233 ), 
        .B(_f_permutation__round__n2232 ), .Z(_f_permutation__round__n2235 )
         );
  XOR2_X2 _f_permutation__round__U4910  ( .A(SYNOPSYS_UNCONNECTED_925), .B(
        _f_permutation__round__n2235 ), .Z(_f_permutation__round__c[931] ) );
  XOR2_X2 _f_permutation__round__U4909  ( .A(SYNOPSYS_UNCONNECTED_796), .B(
        _f_permutation__round__n2234 ), .Z(_f_permutation__round__c[292] ) );
  XOR2_X2 _f_permutation__round__U4908  ( .A(SYNOPSYS_UNCONNECTED_605), .B(
        _f_permutation__round__n2235 ), .Z(_f_permutation__round__c[867] ) );
  XOR2_X2 _f_permutation__round__U4907  ( .A(SYNOPSYS_UNCONNECTED_476), .B(
        _f_permutation__round__n2234 ), .Z(_f_permutation__round__c[228] ) );
  XOR2_X2 _f_permutation__round__U4906  ( .A(SYNOPSYS_UNCONNECTED_285), .B(
        _f_permutation__round__n2235 ), .Z(_f_permutation__round__c[803] ) );
  XOR2_X2 _f_permutation__round__U4905  ( .A(SYNOPSYS_UNCONNECTED_156), .B(
        _f_permutation__round__n2234 ), .Z(_f_permutation__round__c[164] ) );
  XOR2_X2 _f_permutation__round__U4904  ( .A(_f_permutation__round_in[1123]), 
        .B(_f_permutation__round__n2235 ), .Z(_f_permutation__round__c[739] )
         );
  XOR2_X2 _f_permutation__round__U4903  ( .A(_f_permutation__round_in[1252]), 
        .B(_f_permutation__round__n2234 ), .Z(_f_permutation__round__c[100] )
         );
  XOR2_X2 _f_permutation__round__U4902  ( .A(_f_permutation__round_in[1443]), 
        .B(_f_permutation__round__n2235 ), .Z(_f_permutation__round__c[675] )
         );
  XOR2_X2 _f_permutation__round__U4901  ( .A(_f_permutation__round__n2237 ), 
        .B(_f_permutation__round__n2236 ), .Z(_f_permutation__round__n2239 )
         );
  XOR2_X2 _f_permutation__round__U4900  ( .A(SYNOPSYS_UNCONNECTED_926), .B(
        _f_permutation__round__n2239 ), .Z(_f_permutation__round__c[930] ) );
  XOR2_X2 _f_permutation__round__U4899  ( .A(SYNOPSYS_UNCONNECTED_797), .B(
        _f_permutation__round__n2238 ), .Z(_f_permutation__round__c[291] ) );
  XOR2_X2 _f_permutation__round__U4898  ( .A(SYNOPSYS_UNCONNECTED_606), .B(
        _f_permutation__round__n2239 ), .Z(_f_permutation__round__c[866] ) );
  XOR2_X2 _f_permutation__round__U4897  ( .A(SYNOPSYS_UNCONNECTED_477), .B(
        _f_permutation__round__n2238 ), .Z(_f_permutation__round__c[227] ) );
  XOR2_X2 _f_permutation__round__U4896  ( .A(SYNOPSYS_UNCONNECTED_286), .B(
        _f_permutation__round__n2239 ), .Z(_f_permutation__round__c[802] ) );
  XOR2_X2 _f_permutation__round__U4895  ( .A(SYNOPSYS_UNCONNECTED_157), .B(
        _f_permutation__round__n2238 ), .Z(_f_permutation__round__c[163] ) );
  XOR2_X2 _f_permutation__round__U4894  ( .A(_f_permutation__round_in[1122]), 
        .B(_f_permutation__round__n2239 ), .Z(_f_permutation__round__c[738] )
         );
  XOR2_X2 _f_permutation__round__U4893  ( .A(_f_permutation__round_in[1251]), 
        .B(_f_permutation__round__n2238 ), .Z(_f_permutation__round__c[99] )
         );
  XOR2_X2 _f_permutation__round__U4892  ( .A(_f_permutation__round_in[1442]), 
        .B(_f_permutation__round__n2239 ), .Z(_f_permutation__round__c[674] )
         );
  XOR2_X2 _f_permutation__round__U4891  ( .A(_f_permutation__round__n2241 ), 
        .B(_f_permutation__round__n2240 ), .Z(_f_permutation__round__n2243 )
         );
  XOR2_X2 _f_permutation__round__U4890  ( .A(SYNOPSYS_UNCONNECTED_927), .B(
        _f_permutation__round__n2243 ), .Z(_f_permutation__round__c[929] ) );
  XOR2_X2 _f_permutation__round__U4889  ( .A(SYNOPSYS_UNCONNECTED_798), .B(
        _f_permutation__round__n2242 ), .Z(_f_permutation__round__c[290] ) );
  XOR2_X2 _f_permutation__round__U4888  ( .A(SYNOPSYS_UNCONNECTED_607), .B(
        _f_permutation__round__n2243 ), .Z(_f_permutation__round__c[865] ) );
  XOR2_X2 _f_permutation__round__U4887  ( .A(SYNOPSYS_UNCONNECTED_478), .B(
        _f_permutation__round__n2242 ), .Z(_f_permutation__round__c[226] ) );
  XOR2_X2 _f_permutation__round__U4886  ( .A(SYNOPSYS_UNCONNECTED_287), .B(
        _f_permutation__round__n2243 ), .Z(_f_permutation__round__c[801] ) );
  XOR2_X2 _f_permutation__round__U4885  ( .A(SYNOPSYS_UNCONNECTED_158), .B(
        _f_permutation__round__n2242 ), .Z(_f_permutation__round__c[162] ) );
  XOR2_X2 _f_permutation__round__U4884  ( .A(_f_permutation__round_in[1121]), 
        .B(_f_permutation__round__n2243 ), .Z(_f_permutation__round__c[737] )
         );
  XOR2_X2 _f_permutation__round__U4883  ( .A(_f_permutation__round_in[1250]), 
        .B(_f_permutation__round__n2242 ), .Z(_f_permutation__round__c[98] )
         );
  XOR2_X2 _f_permutation__round__U4882  ( .A(_f_permutation__round_in[1441]), 
        .B(_f_permutation__round__n2243 ), .Z(_f_permutation__round__c[673] )
         );
  XOR2_X2 _f_permutation__round__U4881  ( .A(_f_permutation__round__n2245 ), 
        .B(_f_permutation__round__n2244 ), .Z(_f_permutation__round__n2247 )
         );
  XOR2_X2 _f_permutation__round__U4880  ( .A(SYNOPSYS_UNCONNECTED_928), .B(
        _f_permutation__round__n2247 ), .Z(_f_permutation__round__c[928] ) );
  XOR2_X2 _f_permutation__round__U4879  ( .A(SYNOPSYS_UNCONNECTED_799), .B(
        _f_permutation__round__n2246 ), .Z(_f_permutation__round__c[289] ) );
  XOR2_X2 _f_permutation__round__U4878  ( .A(SYNOPSYS_UNCONNECTED_608), .B(
        _f_permutation__round__n2247 ), .Z(_f_permutation__round__c[864] ) );
  XOR2_X2 _f_permutation__round__U4877  ( .A(SYNOPSYS_UNCONNECTED_479), .B(
        _f_permutation__round__n2246 ), .Z(_f_permutation__round__c[225] ) );
  XOR2_X2 _f_permutation__round__U4876  ( .A(SYNOPSYS_UNCONNECTED_288), .B(
        _f_permutation__round__n2247 ), .Z(_f_permutation__round__c[800] ) );
  XOR2_X2 _f_permutation__round__U4875  ( .A(SYNOPSYS_UNCONNECTED_159), .B(
        _f_permutation__round__n2246 ), .Z(_f_permutation__round__c[161] ) );
  XOR2_X2 _f_permutation__round__U4874  ( .A(_f_permutation__round_in[1120]), 
        .B(_f_permutation__round__n2247 ), .Z(_f_permutation__round__c[736] )
         );
  XOR2_X2 _f_permutation__round__U4873  ( .A(_f_permutation__round_in[1249]), 
        .B(_f_permutation__round__n2246 ), .Z(_f_permutation__round__c[97] )
         );
  XOR2_X2 _f_permutation__round__U4872  ( .A(_f_permutation__round_in[1440]), 
        .B(_f_permutation__round__n2247 ), .Z(_f_permutation__round__c[672] )
         );
  XOR2_X2 _f_permutation__round__U4871  ( .A(_f_permutation__round__n2249 ), 
        .B(_f_permutation__round__n2248 ), .Z(_f_permutation__round__n2251 )
         );
  XOR2_X2 _f_permutation__round__U4870  ( .A(SYNOPSYS_UNCONNECTED_929), .B(
        _f_permutation__round__n2251 ), .Z(_f_permutation__round__c[927] ) );
  XOR2_X2 _f_permutation__round__U4869  ( .A(SYNOPSYS_UNCONNECTED_800), .B(
        _f_permutation__round__n2250 ), .Z(_f_permutation__round__c[288] ) );
  XOR2_X2 _f_permutation__round__U4868  ( .A(SYNOPSYS_UNCONNECTED_609), .B(
        _f_permutation__round__n2251 ), .Z(_f_permutation__round__c[863] ) );
  XOR2_X2 _f_permutation__round__U4867  ( .A(SYNOPSYS_UNCONNECTED_480), .B(
        _f_permutation__round__n2250 ), .Z(_f_permutation__round__c[224] ) );
  XOR2_X2 _f_permutation__round__U4866  ( .A(SYNOPSYS_UNCONNECTED_289), .B(
        _f_permutation__round__n2251 ), .Z(_f_permutation__round__c[799] ) );
  XOR2_X2 _f_permutation__round__U4865  ( .A(SYNOPSYS_UNCONNECTED_160), .B(
        _f_permutation__round__n2250 ), .Z(_f_permutation__round__c[160] ) );
  XOR2_X2 _f_permutation__round__U4864  ( .A(_f_permutation__round_in[1119]), 
        .B(_f_permutation__round__n2251 ), .Z(_f_permutation__round__c[735] )
         );
  XOR2_X2 _f_permutation__round__U4863  ( .A(_f_permutation__round_in[1248]), 
        .B(_f_permutation__round__n2250 ), .Z(_f_permutation__round__c[96] )
         );
  XOR2_X2 _f_permutation__round__U4862  ( .A(_f_permutation__round_in[1439]), 
        .B(_f_permutation__round__n2251 ), .Z(_f_permutation__round__c[671] )
         );
  XOR2_X2 _f_permutation__round__U4861  ( .A(_f_permutation__round__n2253 ), 
        .B(_f_permutation__round__n2252 ), .Z(_f_permutation__round__n2255 )
         );
  XOR2_X2 _f_permutation__round__U4860  ( .A(SYNOPSYS_UNCONNECTED_930), .B(
        _f_permutation__round__n2255 ), .Z(_f_permutation__round__c[926] ) );
  XOR2_X2 _f_permutation__round__U4859  ( .A(SYNOPSYS_UNCONNECTED_801), .B(
        _f_permutation__round__n2254 ), .Z(_f_permutation__round__c[287] ) );
  XOR2_X2 _f_permutation__round__U4858  ( .A(SYNOPSYS_UNCONNECTED_610), .B(
        _f_permutation__round__n2255 ), .Z(_f_permutation__round__c[862] ) );
  XOR2_X2 _f_permutation__round__U4857  ( .A(SYNOPSYS_UNCONNECTED_481), .B(
        _f_permutation__round__n2254 ), .Z(_f_permutation__round__c[223] ) );
  XOR2_X2 _f_permutation__round__U4856  ( .A(SYNOPSYS_UNCONNECTED_290), .B(
        _f_permutation__round__n2255 ), .Z(_f_permutation__round__c[798] ) );
  XOR2_X2 _f_permutation__round__U4855  ( .A(SYNOPSYS_UNCONNECTED_161), .B(
        _f_permutation__round__n2254 ), .Z(_f_permutation__round__c[159] ) );
  XOR2_X2 _f_permutation__round__U4854  ( .A(_f_permutation__round_in[1118]), 
        .B(_f_permutation__round__n2255 ), .Z(_f_permutation__round__c[734] )
         );
  XOR2_X2 _f_permutation__round__U4853  ( .A(_f_permutation__round_in[1247]), 
        .B(_f_permutation__round__n2254 ), .Z(_f_permutation__round__c[95] )
         );
  XOR2_X2 _f_permutation__round__U4852  ( .A(_f_permutation__round_in[1438]), 
        .B(_f_permutation__round__n2255 ), .Z(_f_permutation__round__c[670] )
         );
  XOR2_X2 _f_permutation__round__U4851  ( .A(_f_permutation__round__n2257 ), 
        .B(_f_permutation__round__n2256 ), .Z(_f_permutation__round__n2259 )
         );
  XOR2_X2 _f_permutation__round__U4850  ( .A(SYNOPSYS_UNCONNECTED_931), .B(
        _f_permutation__round__n2259 ), .Z(_f_permutation__round__c[925] ) );
  XOR2_X2 _f_permutation__round__U4849  ( .A(SYNOPSYS_UNCONNECTED_802), .B(
        _f_permutation__round__n2258 ), .Z(_f_permutation__round__c[286] ) );
  XOR2_X2 _f_permutation__round__U4848  ( .A(SYNOPSYS_UNCONNECTED_611), .B(
        _f_permutation__round__n2259 ), .Z(_f_permutation__round__c[861] ) );
  XOR2_X2 _f_permutation__round__U4847  ( .A(SYNOPSYS_UNCONNECTED_482), .B(
        _f_permutation__round__n2258 ), .Z(_f_permutation__round__c[222] ) );
  XOR2_X2 _f_permutation__round__U4846  ( .A(SYNOPSYS_UNCONNECTED_291), .B(
        _f_permutation__round__n2259 ), .Z(_f_permutation__round__c[797] ) );
  XOR2_X2 _f_permutation__round__U4845  ( .A(SYNOPSYS_UNCONNECTED_162), .B(
        _f_permutation__round__n2258 ), .Z(_f_permutation__round__c[158] ) );
  XOR2_X2 _f_permutation__round__U4844  ( .A(_f_permutation__round_in[1117]), 
        .B(_f_permutation__round__n2259 ), .Z(_f_permutation__round__c[733] )
         );
  XOR2_X2 _f_permutation__round__U4843  ( .A(_f_permutation__round_in[1246]), 
        .B(_f_permutation__round__n2258 ), .Z(_f_permutation__round__c[94] )
         );
  XOR2_X2 _f_permutation__round__U4842  ( .A(_f_permutation__round_in[1437]), 
        .B(_f_permutation__round__n2259 ), .Z(_f_permutation__round__c[669] )
         );
  XOR2_X2 _f_permutation__round__U4841  ( .A(_f_permutation__round__n2261 ), 
        .B(_f_permutation__round__n2260 ), .Z(_f_permutation__round__n2263 )
         );
  XOR2_X2 _f_permutation__round__U4840  ( .A(SYNOPSYS_UNCONNECTED_932), .B(
        _f_permutation__round__n2263 ), .Z(_f_permutation__round__c[924] ) );
  XOR2_X2 _f_permutation__round__U4839  ( .A(SYNOPSYS_UNCONNECTED_803), .B(
        _f_permutation__round__n2262 ), .Z(_f_permutation__round__c[285] ) );
  XOR2_X2 _f_permutation__round__U4838  ( .A(SYNOPSYS_UNCONNECTED_612), .B(
        _f_permutation__round__n2263 ), .Z(_f_permutation__round__c[860] ) );
  XOR2_X2 _f_permutation__round__U4837  ( .A(SYNOPSYS_UNCONNECTED_483), .B(
        _f_permutation__round__n2262 ), .Z(_f_permutation__round__c[221] ) );
  XOR2_X2 _f_permutation__round__U4836  ( .A(SYNOPSYS_UNCONNECTED_292), .B(
        _f_permutation__round__n2263 ), .Z(_f_permutation__round__c[796] ) );
  XOR2_X2 _f_permutation__round__U4835  ( .A(SYNOPSYS_UNCONNECTED_163), .B(
        _f_permutation__round__n2262 ), .Z(_f_permutation__round__c[157] ) );
  XOR2_X2 _f_permutation__round__U4834  ( .A(_f_permutation__round_in[1116]), 
        .B(_f_permutation__round__n2263 ), .Z(_f_permutation__round__c[732] )
         );
  XOR2_X2 _f_permutation__round__U4833  ( .A(_f_permutation__round_in[1245]), 
        .B(_f_permutation__round__n2262 ), .Z(_f_permutation__round__c[93] )
         );
  XOR2_X2 _f_permutation__round__U4832  ( .A(_f_permutation__round_in[1436]), 
        .B(_f_permutation__round__n2263 ), .Z(_f_permutation__round__c[668] )
         );
  XOR2_X2 _f_permutation__round__U4831  ( .A(_f_permutation__round__n2265 ), 
        .B(_f_permutation__round__n2264 ), .Z(_f_permutation__round__n2267 )
         );
  XOR2_X2 _f_permutation__round__U4830  ( .A(SYNOPSYS_UNCONNECTED_933), .B(
        _f_permutation__round__n2267 ), .Z(_f_permutation__round__c[923] ) );
  XOR2_X2 _f_permutation__round__U4829  ( .A(SYNOPSYS_UNCONNECTED_804), .B(
        _f_permutation__round__n2266 ), .Z(_f_permutation__round__c[284] ) );
  XOR2_X2 _f_permutation__round__U4828  ( .A(SYNOPSYS_UNCONNECTED_613), .B(
        _f_permutation__round__n2267 ), .Z(_f_permutation__round__c[859] ) );
  XOR2_X2 _f_permutation__round__U4827  ( .A(SYNOPSYS_UNCONNECTED_484), .B(
        _f_permutation__round__n2266 ), .Z(_f_permutation__round__c[220] ) );
  XOR2_X2 _f_permutation__round__U4826  ( .A(SYNOPSYS_UNCONNECTED_293), .B(
        _f_permutation__round__n2267 ), .Z(_f_permutation__round__c[795] ) );
  XOR2_X2 _f_permutation__round__U4825  ( .A(SYNOPSYS_UNCONNECTED_164), .B(
        _f_permutation__round__n2266 ), .Z(_f_permutation__round__c[156] ) );
  XOR2_X2 _f_permutation__round__U4824  ( .A(_f_permutation__round_in[1115]), 
        .B(_f_permutation__round__n2267 ), .Z(_f_permutation__round__c[731] )
         );
  XOR2_X2 _f_permutation__round__U4823  ( .A(_f_permutation__round_in[1244]), 
        .B(_f_permutation__round__n2266 ), .Z(_f_permutation__round__c[92] )
         );
  XOR2_X2 _f_permutation__round__U4822  ( .A(_f_permutation__round_in[1435]), 
        .B(_f_permutation__round__n2267 ), .Z(_f_permutation__round__c[667] )
         );
  XOR2_X2 _f_permutation__round__U4821  ( .A(_f_permutation__round__n2269 ), 
        .B(_f_permutation__round__n2268 ), .Z(_f_permutation__round__n2271 )
         );
  XOR2_X2 _f_permutation__round__U4820  ( .A(SYNOPSYS_UNCONNECTED_934), .B(
        _f_permutation__round__n2271 ), .Z(_f_permutation__round__c[922] ) );
  XOR2_X2 _f_permutation__round__U4819  ( .A(SYNOPSYS_UNCONNECTED_805), .B(
        _f_permutation__round__n2270 ), .Z(_f_permutation__round__c[283] ) );
  XOR2_X2 _f_permutation__round__U4818  ( .A(SYNOPSYS_UNCONNECTED_614), .B(
        _f_permutation__round__n2271 ), .Z(_f_permutation__round__c[858] ) );
  XOR2_X2 _f_permutation__round__U4817  ( .A(SYNOPSYS_UNCONNECTED_485), .B(
        _f_permutation__round__n2270 ), .Z(_f_permutation__round__c[219] ) );
  XOR2_X2 _f_permutation__round__U4816  ( .A(SYNOPSYS_UNCONNECTED_294), .B(
        _f_permutation__round__n2271 ), .Z(_f_permutation__round__c[794] ) );
  XOR2_X2 _f_permutation__round__U4815  ( .A(SYNOPSYS_UNCONNECTED_165), .B(
        _f_permutation__round__n2270 ), .Z(_f_permutation__round__c[155] ) );
  XOR2_X2 _f_permutation__round__U4814  ( .A(_f_permutation__round_in[1114]), 
        .B(_f_permutation__round__n2271 ), .Z(_f_permutation__round__c[730] )
         );
  XOR2_X2 _f_permutation__round__U4813  ( .A(_f_permutation__round_in[1243]), 
        .B(_f_permutation__round__n2270 ), .Z(_f_permutation__round__c[91] )
         );
  XOR2_X2 _f_permutation__round__U4812  ( .A(_f_permutation__round_in[1434]), 
        .B(_f_permutation__round__n2271 ), .Z(_f_permutation__round__c[666] )
         );
  XOR2_X2 _f_permutation__round__U4811  ( .A(_f_permutation__round__n2273 ), 
        .B(_f_permutation__round__n2272 ), .Z(_f_permutation__round__n2275 )
         );
  XOR2_X2 _f_permutation__round__U4810  ( .A(SYNOPSYS_UNCONNECTED_935), .B(
        _f_permutation__round__n2275 ), .Z(_f_permutation__round__c[921] ) );
  XOR2_X2 _f_permutation__round__U4809  ( .A(SYNOPSYS_UNCONNECTED_806), .B(
        _f_permutation__round__n2274 ), .Z(_f_permutation__round__c[282] ) );
  XOR2_X2 _f_permutation__round__U4808  ( .A(SYNOPSYS_UNCONNECTED_615), .B(
        _f_permutation__round__n2275 ), .Z(_f_permutation__round__c[857] ) );
  XOR2_X2 _f_permutation__round__U4807  ( .A(SYNOPSYS_UNCONNECTED_486), .B(
        _f_permutation__round__n2274 ), .Z(_f_permutation__round__c[218] ) );
  XOR2_X2 _f_permutation__round__U4806  ( .A(SYNOPSYS_UNCONNECTED_295), .B(
        _f_permutation__round__n2275 ), .Z(_f_permutation__round__c[793] ) );
  XOR2_X2 _f_permutation__round__U4805  ( .A(SYNOPSYS_UNCONNECTED_166), .B(
        _f_permutation__round__n2274 ), .Z(_f_permutation__round__c[154] ) );
  XOR2_X2 _f_permutation__round__U4804  ( .A(_f_permutation__round_in[1113]), 
        .B(_f_permutation__round__n2275 ), .Z(_f_permutation__round__c[729] )
         );
  XOR2_X2 _f_permutation__round__U4803  ( .A(_f_permutation__round_in[1242]), 
        .B(_f_permutation__round__n2274 ), .Z(_f_permutation__round__c[90] )
         );
  XOR2_X2 _f_permutation__round__U4802  ( .A(_f_permutation__round_in[1433]), 
        .B(_f_permutation__round__n2275 ), .Z(_f_permutation__round__c[665] )
         );
  XOR2_X2 _f_permutation__round__U4801  ( .A(_f_permutation__round__n2277 ), 
        .B(_f_permutation__round__n2276 ), .Z(_f_permutation__round__n2279 )
         );
  XOR2_X2 _f_permutation__round__U4800  ( .A(SYNOPSYS_UNCONNECTED_936), .B(
        _f_permutation__round__n2279 ), .Z(_f_permutation__round__c[920] ) );
  XOR2_X2 _f_permutation__round__U4799  ( .A(SYNOPSYS_UNCONNECTED_807), .B(
        _f_permutation__round__n2278 ), .Z(_f_permutation__round__c[281] ) );
  XOR2_X2 _f_permutation__round__U4798  ( .A(SYNOPSYS_UNCONNECTED_616), .B(
        _f_permutation__round__n2279 ), .Z(_f_permutation__round__c[856] ) );
  XOR2_X2 _f_permutation__round__U4797  ( .A(SYNOPSYS_UNCONNECTED_487), .B(
        _f_permutation__round__n2278 ), .Z(_f_permutation__round__c[217] ) );
  XOR2_X2 _f_permutation__round__U4796  ( .A(SYNOPSYS_UNCONNECTED_296), .B(
        _f_permutation__round__n2279 ), .Z(_f_permutation__round__c[792] ) );
  XOR2_X2 _f_permutation__round__U4795  ( .A(SYNOPSYS_UNCONNECTED_167), .B(
        _f_permutation__round__n2278 ), .Z(_f_permutation__round__c[153] ) );
  XOR2_X2 _f_permutation__round__U4794  ( .A(_f_permutation__round_in[1112]), 
        .B(_f_permutation__round__n2279 ), .Z(_f_permutation__round__c[728] )
         );
  XOR2_X2 _f_permutation__round__U4793  ( .A(_f_permutation__round_in[1241]), 
        .B(_f_permutation__round__n2278 ), .Z(_f_permutation__round__c[89] )
         );
  XOR2_X2 _f_permutation__round__U4792  ( .A(_f_permutation__round_in[1432]), 
        .B(_f_permutation__round__n2279 ), .Z(_f_permutation__round__c[664] )
         );
  XOR2_X2 _f_permutation__round__U4791  ( .A(_f_permutation__round__n2281 ), 
        .B(_f_permutation__round__n2280 ), .Z(_f_permutation__round__n2283 )
         );
  XOR2_X2 _f_permutation__round__U4790  ( .A(SYNOPSYS_UNCONNECTED_937), .B(
        _f_permutation__round__n2283 ), .Z(_f_permutation__round__c[919] ) );
  XOR2_X2 _f_permutation__round__U4789  ( .A(SYNOPSYS_UNCONNECTED_808), .B(
        _f_permutation__round__n2282 ), .Z(_f_permutation__round__c[280] ) );
  XOR2_X2 _f_permutation__round__U4788  ( .A(SYNOPSYS_UNCONNECTED_617), .B(
        _f_permutation__round__n2283 ), .Z(_f_permutation__round__c[855] ) );
  XOR2_X2 _f_permutation__round__U4787  ( .A(SYNOPSYS_UNCONNECTED_488), .B(
        _f_permutation__round__n2282 ), .Z(_f_permutation__round__c[216] ) );
  XOR2_X2 _f_permutation__round__U4786  ( .A(SYNOPSYS_UNCONNECTED_297), .B(
        _f_permutation__round__n2283 ), .Z(_f_permutation__round__c[791] ) );
  XOR2_X2 _f_permutation__round__U4785  ( .A(SYNOPSYS_UNCONNECTED_168), .B(
        _f_permutation__round__n2282 ), .Z(_f_permutation__round__c[152] ) );
  XOR2_X2 _f_permutation__round__U4784  ( .A(_f_permutation__round_in[1111]), 
        .B(_f_permutation__round__n2283 ), .Z(_f_permutation__round__c[727] )
         );
  XOR2_X2 _f_permutation__round__U4783  ( .A(_f_permutation__round_in[1240]), 
        .B(_f_permutation__round__n2282 ), .Z(_f_permutation__round__c[88] )
         );
  XOR2_X2 _f_permutation__round__U4782  ( .A(_f_permutation__round_in[1431]), 
        .B(_f_permutation__round__n2283 ), .Z(_f_permutation__round__c[663] )
         );
  XOR2_X2 _f_permutation__round__U4781  ( .A(_f_permutation__round__n2285 ), 
        .B(_f_permutation__round__n2284 ), .Z(_f_permutation__round__n2287 )
         );
  XOR2_X2 _f_permutation__round__U4780  ( .A(SYNOPSYS_UNCONNECTED_938), .B(
        _f_permutation__round__n2287 ), .Z(_f_permutation__round__c[918] ) );
  XOR2_X2 _f_permutation__round__U4779  ( .A(SYNOPSYS_UNCONNECTED_809), .B(
        _f_permutation__round__n2286 ), .Z(_f_permutation__round__c[279] ) );
  XOR2_X2 _f_permutation__round__U4778  ( .A(SYNOPSYS_UNCONNECTED_618), .B(
        _f_permutation__round__n2287 ), .Z(_f_permutation__round__c[854] ) );
  XOR2_X2 _f_permutation__round__U4777  ( .A(SYNOPSYS_UNCONNECTED_489), .B(
        _f_permutation__round__n2286 ), .Z(_f_permutation__round__c[215] ) );
  XOR2_X2 _f_permutation__round__U4776  ( .A(SYNOPSYS_UNCONNECTED_298), .B(
        _f_permutation__round__n2287 ), .Z(_f_permutation__round__c[790] ) );
  XOR2_X2 _f_permutation__round__U4775  ( .A(SYNOPSYS_UNCONNECTED_169), .B(
        _f_permutation__round__n2286 ), .Z(_f_permutation__round__c[151] ) );
  XOR2_X2 _f_permutation__round__U4774  ( .A(_f_permutation__round_in[1110]), 
        .B(_f_permutation__round__n2287 ), .Z(_f_permutation__round__c[726] )
         );
  XOR2_X2 _f_permutation__round__U4773  ( .A(_f_permutation__round_in[1239]), 
        .B(_f_permutation__round__n2286 ), .Z(_f_permutation__round__c[87] )
         );
  XOR2_X2 _f_permutation__round__U4772  ( .A(_f_permutation__round_in[1430]), 
        .B(_f_permutation__round__n2287 ), .Z(_f_permutation__round__c[662] )
         );
  XOR2_X2 _f_permutation__round__U4771  ( .A(_f_permutation__round__n2289 ), 
        .B(_f_permutation__round__n2288 ), .Z(_f_permutation__round__n2291 )
         );
  XOR2_X2 _f_permutation__round__U4770  ( .A(SYNOPSYS_UNCONNECTED_939), .B(
        _f_permutation__round__n2291 ), .Z(_f_permutation__round__c[917] ) );
  XOR2_X2 _f_permutation__round__U4769  ( .A(SYNOPSYS_UNCONNECTED_810), .B(
        _f_permutation__round__n2290 ), .Z(_f_permutation__round__c[278] ) );
  XOR2_X2 _f_permutation__round__U4768  ( .A(SYNOPSYS_UNCONNECTED_619), .B(
        _f_permutation__round__n2291 ), .Z(_f_permutation__round__c[853] ) );
  XOR2_X2 _f_permutation__round__U4767  ( .A(SYNOPSYS_UNCONNECTED_490), .B(
        _f_permutation__round__n2290 ), .Z(_f_permutation__round__c[214] ) );
  XOR2_X2 _f_permutation__round__U4766  ( .A(SYNOPSYS_UNCONNECTED_299), .B(
        _f_permutation__round__n2291 ), .Z(_f_permutation__round__c[789] ) );
  XOR2_X2 _f_permutation__round__U4765  ( .A(SYNOPSYS_UNCONNECTED_170), .B(
        _f_permutation__round__n2290 ), .Z(_f_permutation__round__c[150] ) );
  XOR2_X2 _f_permutation__round__U4764  ( .A(_f_permutation__round_in[1109]), 
        .B(_f_permutation__round__n2291 ), .Z(_f_permutation__round__c[725] )
         );
  XOR2_X2 _f_permutation__round__U4763  ( .A(_f_permutation__round_in[1238]), 
        .B(_f_permutation__round__n2290 ), .Z(_f_permutation__round__c[86] )
         );
  XOR2_X2 _f_permutation__round__U4762  ( .A(_f_permutation__round_in[1429]), 
        .B(_f_permutation__round__n2291 ), .Z(_f_permutation__round__c[661] )
         );
  XOR2_X2 _f_permutation__round__U4761  ( .A(_f_permutation__round__n2293 ), 
        .B(_f_permutation__round__n2292 ), .Z(_f_permutation__round__n2295 )
         );
  XOR2_X2 _f_permutation__round__U4760  ( .A(SYNOPSYS_UNCONNECTED_940), .B(
        _f_permutation__round__n2295 ), .Z(_f_permutation__round__c[916] ) );
  XOR2_X2 _f_permutation__round__U4759  ( .A(SYNOPSYS_UNCONNECTED_811), .B(
        _f_permutation__round__n2294 ), .Z(_f_permutation__round__c[277] ) );
  XOR2_X2 _f_permutation__round__U4758  ( .A(SYNOPSYS_UNCONNECTED_620), .B(
        _f_permutation__round__n2295 ), .Z(_f_permutation__round__c[852] ) );
  XOR2_X2 _f_permutation__round__U4757  ( .A(SYNOPSYS_UNCONNECTED_491), .B(
        _f_permutation__round__n2294 ), .Z(_f_permutation__round__c[213] ) );
  XOR2_X2 _f_permutation__round__U4756  ( .A(SYNOPSYS_UNCONNECTED_300), .B(
        _f_permutation__round__n2295 ), .Z(_f_permutation__round__c[788] ) );
  XOR2_X2 _f_permutation__round__U4755  ( .A(SYNOPSYS_UNCONNECTED_171), .B(
        _f_permutation__round__n2294 ), .Z(_f_permutation__round__c[149] ) );
  XOR2_X2 _f_permutation__round__U4754  ( .A(_f_permutation__round_in[1108]), 
        .B(_f_permutation__round__n2295 ), .Z(_f_permutation__round__c[724] )
         );
  XOR2_X2 _f_permutation__round__U4753  ( .A(_f_permutation__round_in[1237]), 
        .B(_f_permutation__round__n2294 ), .Z(_f_permutation__round__c[85] )
         );
  XOR2_X2 _f_permutation__round__U4752  ( .A(_f_permutation__round_in[1428]), 
        .B(_f_permutation__round__n2295 ), .Z(_f_permutation__round__c[660] )
         );
  XOR2_X2 _f_permutation__round__U4751  ( .A(_f_permutation__round__n2297 ), 
        .B(_f_permutation__round__n2296 ), .Z(_f_permutation__round__n2299 )
         );
  XOR2_X2 _f_permutation__round__U4750  ( .A(SYNOPSYS_UNCONNECTED_941), .B(
        _f_permutation__round__n2299 ), .Z(_f_permutation__round__c[915] ) );
  XOR2_X2 _f_permutation__round__U4749  ( .A(SYNOPSYS_UNCONNECTED_812), .B(
        _f_permutation__round__n2298 ), .Z(_f_permutation__round__c[276] ) );
  XOR2_X2 _f_permutation__round__U4748  ( .A(SYNOPSYS_UNCONNECTED_621), .B(
        _f_permutation__round__n2299 ), .Z(_f_permutation__round__c[851] ) );
  XOR2_X2 _f_permutation__round__U4747  ( .A(SYNOPSYS_UNCONNECTED_492), .B(
        _f_permutation__round__n2298 ), .Z(_f_permutation__round__c[212] ) );
  XOR2_X2 _f_permutation__round__U4746  ( .A(SYNOPSYS_UNCONNECTED_301), .B(
        _f_permutation__round__n2299 ), .Z(_f_permutation__round__c[787] ) );
  XOR2_X2 _f_permutation__round__U4745  ( .A(SYNOPSYS_UNCONNECTED_172), .B(
        _f_permutation__round__n2298 ), .Z(_f_permutation__round__c[148] ) );
  XOR2_X2 _f_permutation__round__U4744  ( .A(_f_permutation__round_in[1107]), 
        .B(_f_permutation__round__n2299 ), .Z(_f_permutation__round__c[723] )
         );
  XOR2_X2 _f_permutation__round__U4743  ( .A(_f_permutation__round_in[1236]), 
        .B(_f_permutation__round__n2298 ), .Z(_f_permutation__round__c[84] )
         );
  XOR2_X2 _f_permutation__round__U4742  ( .A(_f_permutation__round_in[1427]), 
        .B(_f_permutation__round__n2299 ), .Z(_f_permutation__round__c[659] )
         );
  XOR2_X2 _f_permutation__round__U4741  ( .A(_f_permutation__round__n2301 ), 
        .B(_f_permutation__round__n2300 ), .Z(_f_permutation__round__n2303 )
         );
  XOR2_X2 _f_permutation__round__U4740  ( .A(SYNOPSYS_UNCONNECTED_942), .B(
        _f_permutation__round__n2303 ), .Z(_f_permutation__round__c[914] ) );
  XOR2_X2 _f_permutation__round__U4739  ( .A(SYNOPSYS_UNCONNECTED_813), .B(
        _f_permutation__round__n2302 ), .Z(_f_permutation__round__c[275] ) );
  XOR2_X2 _f_permutation__round__U4738  ( .A(SYNOPSYS_UNCONNECTED_622), .B(
        _f_permutation__round__n2303 ), .Z(_f_permutation__round__c[850] ) );
  XOR2_X2 _f_permutation__round__U4737  ( .A(SYNOPSYS_UNCONNECTED_493), .B(
        _f_permutation__round__n2302 ), .Z(_f_permutation__round__c[211] ) );
  XOR2_X2 _f_permutation__round__U4736  ( .A(SYNOPSYS_UNCONNECTED_302), .B(
        _f_permutation__round__n2303 ), .Z(_f_permutation__round__c[786] ) );
  XOR2_X2 _f_permutation__round__U4735  ( .A(SYNOPSYS_UNCONNECTED_173), .B(
        _f_permutation__round__n2302 ), .Z(_f_permutation__round__c[147] ) );
  XOR2_X2 _f_permutation__round__U4734  ( .A(_f_permutation__round_in[1106]), 
        .B(_f_permutation__round__n2303 ), .Z(_f_permutation__round__c[722] )
         );
  XOR2_X2 _f_permutation__round__U4733  ( .A(_f_permutation__round_in[1235]), 
        .B(_f_permutation__round__n2302 ), .Z(_f_permutation__round__c[83] )
         );
  XOR2_X2 _f_permutation__round__U4732  ( .A(_f_permutation__round_in[1426]), 
        .B(_f_permutation__round__n2303 ), .Z(_f_permutation__round__c[658] )
         );
  XOR2_X2 _f_permutation__round__U4731  ( .A(_f_permutation__round__n2305 ), 
        .B(_f_permutation__round__n2304 ), .Z(_f_permutation__round__n2307 )
         );
  XOR2_X2 _f_permutation__round__U4730  ( .A(SYNOPSYS_UNCONNECTED_943), .B(
        _f_permutation__round__n2307 ), .Z(_f_permutation__round__c[913] ) );
  XOR2_X2 _f_permutation__round__U4729  ( .A(SYNOPSYS_UNCONNECTED_814), .B(
        _f_permutation__round__n2306 ), .Z(_f_permutation__round__c[274] ) );
  XOR2_X2 _f_permutation__round__U4728  ( .A(SYNOPSYS_UNCONNECTED_623), .B(
        _f_permutation__round__n2307 ), .Z(_f_permutation__round__c[849] ) );
  XOR2_X2 _f_permutation__round__U4727  ( .A(SYNOPSYS_UNCONNECTED_494), .B(
        _f_permutation__round__n2306 ), .Z(_f_permutation__round__c[210] ) );
  XOR2_X2 _f_permutation__round__U4726  ( .A(SYNOPSYS_UNCONNECTED_303), .B(
        _f_permutation__round__n2307 ), .Z(_f_permutation__round__c[785] ) );
  XOR2_X2 _f_permutation__round__U4725  ( .A(SYNOPSYS_UNCONNECTED_174), .B(
        _f_permutation__round__n2306 ), .Z(_f_permutation__round__c[146] ) );
  XOR2_X2 _f_permutation__round__U4724  ( .A(_f_permutation__round_in[1105]), 
        .B(_f_permutation__round__n2307 ), .Z(_f_permutation__round__c[721] )
         );
  XOR2_X2 _f_permutation__round__U4723  ( .A(_f_permutation__round_in[1234]), 
        .B(_f_permutation__round__n2306 ), .Z(_f_permutation__round__c[82] )
         );
  XOR2_X2 _f_permutation__round__U4722  ( .A(_f_permutation__round_in[1425]), 
        .B(_f_permutation__round__n2307 ), .Z(_f_permutation__round__c[657] )
         );
  XOR2_X2 _f_permutation__round__U4721  ( .A(_f_permutation__round__n2309 ), 
        .B(_f_permutation__round__n2308 ), .Z(_f_permutation__round__n2311 )
         );
  XOR2_X2 _f_permutation__round__U4720  ( .A(SYNOPSYS_UNCONNECTED_944), .B(
        _f_permutation__round__n2311 ), .Z(_f_permutation__round__c[912] ) );
  XOR2_X2 _f_permutation__round__U4719  ( .A(SYNOPSYS_UNCONNECTED_815), .B(
        _f_permutation__round__n2310 ), .Z(_f_permutation__round__c[273] ) );
  XOR2_X2 _f_permutation__round__U4718  ( .A(SYNOPSYS_UNCONNECTED_624), .B(
        _f_permutation__round__n2311 ), .Z(_f_permutation__round__c[848] ) );
  XOR2_X2 _f_permutation__round__U4717  ( .A(SYNOPSYS_UNCONNECTED_495), .B(
        _f_permutation__round__n2310 ), .Z(_f_permutation__round__c[209] ) );
  XOR2_X2 _f_permutation__round__U4716  ( .A(SYNOPSYS_UNCONNECTED_304), .B(
        _f_permutation__round__n2311 ), .Z(_f_permutation__round__c[784] ) );
  XOR2_X2 _f_permutation__round__U4715  ( .A(SYNOPSYS_UNCONNECTED_175), .B(
        _f_permutation__round__n2310 ), .Z(_f_permutation__round__c[145] ) );
  XOR2_X2 _f_permutation__round__U4714  ( .A(_f_permutation__round_in[1104]), 
        .B(_f_permutation__round__n2311 ), .Z(_f_permutation__round__c[720] )
         );
  XOR2_X2 _f_permutation__round__U4713  ( .A(_f_permutation__round_in[1233]), 
        .B(_f_permutation__round__n2310 ), .Z(_f_permutation__round__c[81] )
         );
  XOR2_X2 _f_permutation__round__U4712  ( .A(_f_permutation__round_in[1424]), 
        .B(_f_permutation__round__n2311 ), .Z(_f_permutation__round__c[656] )
         );
  XOR2_X2 _f_permutation__round__U4711  ( .A(_f_permutation__round__n2313 ), 
        .B(_f_permutation__round__n2312 ), .Z(_f_permutation__round__n2315 )
         );
  XOR2_X2 _f_permutation__round__U4710  ( .A(SYNOPSYS_UNCONNECTED_945), .B(
        _f_permutation__round__n2315 ), .Z(_f_permutation__round__c[911] ) );
  XOR2_X2 _f_permutation__round__U4709  ( .A(SYNOPSYS_UNCONNECTED_816), .B(
        _f_permutation__round__n2314 ), .Z(_f_permutation__round__c[272] ) );
  XOR2_X2 _f_permutation__round__U4708  ( .A(SYNOPSYS_UNCONNECTED_625), .B(
        _f_permutation__round__n2315 ), .Z(_f_permutation__round__c[847] ) );
  XOR2_X2 _f_permutation__round__U4707  ( .A(SYNOPSYS_UNCONNECTED_496), .B(
        _f_permutation__round__n2314 ), .Z(_f_permutation__round__c[208] ) );
  XOR2_X2 _f_permutation__round__U4706  ( .A(SYNOPSYS_UNCONNECTED_305), .B(
        _f_permutation__round__n2315 ), .Z(_f_permutation__round__c[783] ) );
  XOR2_X2 _f_permutation__round__U4705  ( .A(SYNOPSYS_UNCONNECTED_176), .B(
        _f_permutation__round__n2314 ), .Z(_f_permutation__round__c[144] ) );
  XOR2_X2 _f_permutation__round__U4704  ( .A(_f_permutation__round_in[1103]), 
        .B(_f_permutation__round__n2315 ), .Z(_f_permutation__round__c[719] )
         );
  XOR2_X2 _f_permutation__round__U4703  ( .A(_f_permutation__round_in[1232]), 
        .B(_f_permutation__round__n2314 ), .Z(_f_permutation__round__c[80] )
         );
  XOR2_X2 _f_permutation__round__U4702  ( .A(_f_permutation__round_in[1423]), 
        .B(_f_permutation__round__n2315 ), .Z(_f_permutation__round__c[655] )
         );
  XOR2_X2 _f_permutation__round__U4701  ( .A(_f_permutation__round__n2317 ), 
        .B(_f_permutation__round__n2316 ), .Z(_f_permutation__round__n2319 )
         );
  XOR2_X2 _f_permutation__round__U4700  ( .A(SYNOPSYS_UNCONNECTED_946), .B(
        _f_permutation__round__n2319 ), .Z(_f_permutation__round__c[910] ) );
  XOR2_X2 _f_permutation__round__U4699  ( .A(SYNOPSYS_UNCONNECTED_817), .B(
        _f_permutation__round__n2318 ), .Z(_f_permutation__round__c[271] ) );
  XOR2_X2 _f_permutation__round__U4698  ( .A(SYNOPSYS_UNCONNECTED_626), .B(
        _f_permutation__round__n2319 ), .Z(_f_permutation__round__c[846] ) );
  XOR2_X2 _f_permutation__round__U4697  ( .A(SYNOPSYS_UNCONNECTED_497), .B(
        _f_permutation__round__n2318 ), .Z(_f_permutation__round__c[207] ) );
  XOR2_X2 _f_permutation__round__U4696  ( .A(SYNOPSYS_UNCONNECTED_306), .B(
        _f_permutation__round__n2319 ), .Z(_f_permutation__round__c[782] ) );
  XOR2_X2 _f_permutation__round__U4695  ( .A(SYNOPSYS_UNCONNECTED_177), .B(
        _f_permutation__round__n2318 ), .Z(_f_permutation__round__c[143] ) );
  XOR2_X2 _f_permutation__round__U4694  ( .A(_f_permutation__round_in[1102]), 
        .B(_f_permutation__round__n2319 ), .Z(_f_permutation__round__c[718] )
         );
  XOR2_X2 _f_permutation__round__U4693  ( .A(_f_permutation__round_in[1231]), 
        .B(_f_permutation__round__n2318 ), .Z(_f_permutation__round__c[79] )
         );
  XOR2_X2 _f_permutation__round__U4692  ( .A(_f_permutation__round_in[1422]), 
        .B(_f_permutation__round__n2319 ), .Z(_f_permutation__round__c[654] )
         );
  XOR2_X2 _f_permutation__round__U4691  ( .A(_f_permutation__round__n2321 ), 
        .B(_f_permutation__round__n2320 ), .Z(_f_permutation__round__n2323 )
         );
  XOR2_X2 _f_permutation__round__U4690  ( .A(SYNOPSYS_UNCONNECTED_947), .B(
        _f_permutation__round__n2323 ), .Z(_f_permutation__round__c[909] ) );
  XOR2_X2 _f_permutation__round__U4689  ( .A(SYNOPSYS_UNCONNECTED_818), .B(
        _f_permutation__round__n2322 ), .Z(_f_permutation__round__c[270] ) );
  XOR2_X2 _f_permutation__round__U4688  ( .A(SYNOPSYS_UNCONNECTED_627), .B(
        _f_permutation__round__n2323 ), .Z(_f_permutation__round__c[845] ) );
  XOR2_X2 _f_permutation__round__U4687  ( .A(SYNOPSYS_UNCONNECTED_498), .B(
        _f_permutation__round__n2322 ), .Z(_f_permutation__round__c[206] ) );
  XOR2_X2 _f_permutation__round__U4686  ( .A(SYNOPSYS_UNCONNECTED_307), .B(
        _f_permutation__round__n2323 ), .Z(_f_permutation__round__c[781] ) );
  XOR2_X2 _f_permutation__round__U4685  ( .A(SYNOPSYS_UNCONNECTED_178), .B(
        _f_permutation__round__n2322 ), .Z(_f_permutation__round__c[142] ) );
  XOR2_X2 _f_permutation__round__U4684  ( .A(_f_permutation__round_in[1101]), 
        .B(_f_permutation__round__n2323 ), .Z(_f_permutation__round__c[717] )
         );
  XOR2_X2 _f_permutation__round__U4683  ( .A(_f_permutation__round_in[1230]), 
        .B(_f_permutation__round__n2322 ), .Z(_f_permutation__round__c[78] )
         );
  XOR2_X2 _f_permutation__round__U4682  ( .A(_f_permutation__round_in[1421]), 
        .B(_f_permutation__round__n2323 ), .Z(_f_permutation__round__c[653] )
         );
  XOR2_X2 _f_permutation__round__U4681  ( .A(_f_permutation__round__n2325 ), 
        .B(_f_permutation__round__n2324 ), .Z(_f_permutation__round__n2327 )
         );
  XOR2_X2 _f_permutation__round__U4680  ( .A(SYNOPSYS_UNCONNECTED_948), .B(
        _f_permutation__round__n2327 ), .Z(_f_permutation__round__c[908] ) );
  XOR2_X2 _f_permutation__round__U4679  ( .A(SYNOPSYS_UNCONNECTED_819), .B(
        _f_permutation__round__n2326 ), .Z(_f_permutation__round__c[269] ) );
  XOR2_X2 _f_permutation__round__U4678  ( .A(SYNOPSYS_UNCONNECTED_628), .B(
        _f_permutation__round__n2327 ), .Z(_f_permutation__round__c[844] ) );
  XOR2_X2 _f_permutation__round__U4677  ( .A(SYNOPSYS_UNCONNECTED_499), .B(
        _f_permutation__round__n2326 ), .Z(_f_permutation__round__c[205] ) );
  XOR2_X2 _f_permutation__round__U4676  ( .A(SYNOPSYS_UNCONNECTED_308), .B(
        _f_permutation__round__n2327 ), .Z(_f_permutation__round__c[780] ) );
  XOR2_X2 _f_permutation__round__U4675  ( .A(SYNOPSYS_UNCONNECTED_179), .B(
        _f_permutation__round__n2326 ), .Z(_f_permutation__round__c[141] ) );
  XOR2_X2 _f_permutation__round__U4674  ( .A(_f_permutation__round_in[1100]), 
        .B(_f_permutation__round__n2327 ), .Z(_f_permutation__round__c[716] )
         );
  XOR2_X2 _f_permutation__round__U4673  ( .A(_f_permutation__round_in[1229]), 
        .B(_f_permutation__round__n2326 ), .Z(_f_permutation__round__c[77] )
         );
  XOR2_X2 _f_permutation__round__U4672  ( .A(_f_permutation__round_in[1420]), 
        .B(_f_permutation__round__n2327 ), .Z(_f_permutation__round__c[652] )
         );
  XOR2_X2 _f_permutation__round__U4671  ( .A(_f_permutation__round__n2329 ), 
        .B(_f_permutation__round__n2328 ), .Z(_f_permutation__round__n2331 )
         );
  XOR2_X2 _f_permutation__round__U4670  ( .A(SYNOPSYS_UNCONNECTED_949), .B(
        _f_permutation__round__n2331 ), .Z(_f_permutation__round__c[907] ) );
  XOR2_X2 _f_permutation__round__U4669  ( .A(SYNOPSYS_UNCONNECTED_820), .B(
        _f_permutation__round__n2330 ), .Z(_f_permutation__round__c[268] ) );
  XOR2_X2 _f_permutation__round__U4668  ( .A(SYNOPSYS_UNCONNECTED_629), .B(
        _f_permutation__round__n2331 ), .Z(_f_permutation__round__c[843] ) );
  XOR2_X2 _f_permutation__round__U4667  ( .A(SYNOPSYS_UNCONNECTED_500), .B(
        _f_permutation__round__n2330 ), .Z(_f_permutation__round__c[204] ) );
  XOR2_X2 _f_permutation__round__U4666  ( .A(SYNOPSYS_UNCONNECTED_309), .B(
        _f_permutation__round__n2331 ), .Z(_f_permutation__round__c[779] ) );
  XOR2_X2 _f_permutation__round__U4665  ( .A(SYNOPSYS_UNCONNECTED_180), .B(
        _f_permutation__round__n2330 ), .Z(_f_permutation__round__c[140] ) );
  XOR2_X2 _f_permutation__round__U4664  ( .A(_f_permutation__round_in[1099]), 
        .B(_f_permutation__round__n2331 ), .Z(_f_permutation__round__c[715] )
         );
  XOR2_X2 _f_permutation__round__U4663  ( .A(_f_permutation__round_in[1228]), 
        .B(_f_permutation__round__n2330 ), .Z(_f_permutation__round__c[76] )
         );
  XOR2_X2 _f_permutation__round__U4662  ( .A(_f_permutation__round_in[1419]), 
        .B(_f_permutation__round__n2331 ), .Z(_f_permutation__round__c[651] )
         );
  XOR2_X2 _f_permutation__round__U4661  ( .A(_f_permutation__round__n2333 ), 
        .B(_f_permutation__round__n2332 ), .Z(_f_permutation__round__n2335 )
         );
  XOR2_X2 _f_permutation__round__U4660  ( .A(SYNOPSYS_UNCONNECTED_950), .B(
        _f_permutation__round__n2335 ), .Z(_f_permutation__round__c[906] ) );
  XOR2_X2 _f_permutation__round__U4659  ( .A(SYNOPSYS_UNCONNECTED_821), .B(
        _f_permutation__round__n2334 ), .Z(_f_permutation__round__c[267] ) );
  XOR2_X2 _f_permutation__round__U4658  ( .A(SYNOPSYS_UNCONNECTED_630), .B(
        _f_permutation__round__n2335 ), .Z(_f_permutation__round__c[842] ) );
  XOR2_X2 _f_permutation__round__U4657  ( .A(SYNOPSYS_UNCONNECTED_501), .B(
        _f_permutation__round__n2334 ), .Z(_f_permutation__round__c[203] ) );
  XOR2_X2 _f_permutation__round__U4656  ( .A(SYNOPSYS_UNCONNECTED_310), .B(
        _f_permutation__round__n2335 ), .Z(_f_permutation__round__c[778] ) );
  XOR2_X2 _f_permutation__round__U4655  ( .A(SYNOPSYS_UNCONNECTED_181), .B(
        _f_permutation__round__n2334 ), .Z(_f_permutation__round__c[139] ) );
  XOR2_X2 _f_permutation__round__U4654  ( .A(_f_permutation__round_in[1098]), 
        .B(_f_permutation__round__n2335 ), .Z(_f_permutation__round__c[714] )
         );
  XOR2_X2 _f_permutation__round__U4653  ( .A(_f_permutation__round_in[1227]), 
        .B(_f_permutation__round__n2334 ), .Z(_f_permutation__round__c[75] )
         );
  XOR2_X2 _f_permutation__round__U4652  ( .A(_f_permutation__round_in[1418]), 
        .B(_f_permutation__round__n2335 ), .Z(_f_permutation__round__c[650] )
         );
  XOR2_X2 _f_permutation__round__U4651  ( .A(_f_permutation__round__n2337 ), 
        .B(_f_permutation__round__n2336 ), .Z(_f_permutation__round__n2339 )
         );
  XOR2_X2 _f_permutation__round__U4650  ( .A(SYNOPSYS_UNCONNECTED_951), .B(
        _f_permutation__round__n2339 ), .Z(_f_permutation__round__c[905] ) );
  XOR2_X2 _f_permutation__round__U4649  ( .A(SYNOPSYS_UNCONNECTED_822), .B(
        _f_permutation__round__n2338 ), .Z(_f_permutation__round__c[266] ) );
  XOR2_X2 _f_permutation__round__U4648  ( .A(SYNOPSYS_UNCONNECTED_631), .B(
        _f_permutation__round__n2339 ), .Z(_f_permutation__round__c[841] ) );
  XOR2_X2 _f_permutation__round__U4647  ( .A(SYNOPSYS_UNCONNECTED_502), .B(
        _f_permutation__round__n2338 ), .Z(_f_permutation__round__c[202] ) );
  XOR2_X2 _f_permutation__round__U4646  ( .A(SYNOPSYS_UNCONNECTED_311), .B(
        _f_permutation__round__n2339 ), .Z(_f_permutation__round__c[777] ) );
  XOR2_X2 _f_permutation__round__U4645  ( .A(SYNOPSYS_UNCONNECTED_182), .B(
        _f_permutation__round__n2338 ), .Z(_f_permutation__round__c[138] ) );
  XOR2_X2 _f_permutation__round__U4644  ( .A(_f_permutation__round_in[1097]), 
        .B(_f_permutation__round__n2339 ), .Z(_f_permutation__round__c[713] )
         );
  XOR2_X2 _f_permutation__round__U4643  ( .A(_f_permutation__round_in[1226]), 
        .B(_f_permutation__round__n2338 ), .Z(_f_permutation__round__c[74] )
         );
  XOR2_X2 _f_permutation__round__U4642  ( .A(_f_permutation__round_in[1417]), 
        .B(_f_permutation__round__n2339 ), .Z(_f_permutation__round__c[649] )
         );
  XOR2_X2 _f_permutation__round__U4641  ( .A(_f_permutation__round__n2341 ), 
        .B(_f_permutation__round__n2340 ), .Z(_f_permutation__round__n2343 )
         );
  XOR2_X2 _f_permutation__round__U4640  ( .A(SYNOPSYS_UNCONNECTED_952), .B(
        _f_permutation__round__n2343 ), .Z(_f_permutation__round__c[904] ) );
  XOR2_X2 _f_permutation__round__U4639  ( .A(SYNOPSYS_UNCONNECTED_823), .B(
        _f_permutation__round__n2342 ), .Z(_f_permutation__round__c[265] ) );
  XOR2_X2 _f_permutation__round__U4638  ( .A(SYNOPSYS_UNCONNECTED_632), .B(
        _f_permutation__round__n2343 ), .Z(_f_permutation__round__c[840] ) );
  XOR2_X2 _f_permutation__round__U4637  ( .A(SYNOPSYS_UNCONNECTED_503), .B(
        _f_permutation__round__n2342 ), .Z(_f_permutation__round__c[201] ) );
  XOR2_X2 _f_permutation__round__U4636  ( .A(SYNOPSYS_UNCONNECTED_312), .B(
        _f_permutation__round__n2343 ), .Z(_f_permutation__round__c[776] ) );
  XOR2_X2 _f_permutation__round__U4635  ( .A(SYNOPSYS_UNCONNECTED_183), .B(
        _f_permutation__round__n2342 ), .Z(_f_permutation__round__c[137] ) );
  XOR2_X2 _f_permutation__round__U4634  ( .A(_f_permutation__round_in[1096]), 
        .B(_f_permutation__round__n2343 ), .Z(_f_permutation__round__c[712] )
         );
  XOR2_X2 _f_permutation__round__U4633  ( .A(_f_permutation__round_in[1225]), 
        .B(_f_permutation__round__n2342 ), .Z(_f_permutation__round__c[73] )
         );
  XOR2_X2 _f_permutation__round__U4632  ( .A(_f_permutation__round_in[1416]), 
        .B(_f_permutation__round__n2343 ), .Z(_f_permutation__round__c[648] )
         );
  XOR2_X2 _f_permutation__round__U4631  ( .A(_f_permutation__round__n2345 ), 
        .B(_f_permutation__round__n2344 ), .Z(_f_permutation__round__n2347 )
         );
  XOR2_X2 _f_permutation__round__U4630  ( .A(SYNOPSYS_UNCONNECTED_953), .B(
        _f_permutation__round__n2347 ), .Z(_f_permutation__round__c[903] ) );
  XOR2_X2 _f_permutation__round__U4629  ( .A(SYNOPSYS_UNCONNECTED_824), .B(
        _f_permutation__round__n2346 ), .Z(_f_permutation__round__c[264] ) );
  XOR2_X2 _f_permutation__round__U4628  ( .A(SYNOPSYS_UNCONNECTED_633), .B(
        _f_permutation__round__n2347 ), .Z(_f_permutation__round__c[839] ) );
  XOR2_X2 _f_permutation__round__U4627  ( .A(SYNOPSYS_UNCONNECTED_504), .B(
        _f_permutation__round__n2346 ), .Z(_f_permutation__round__c[200] ) );
  XOR2_X2 _f_permutation__round__U4626  ( .A(SYNOPSYS_UNCONNECTED_313), .B(
        _f_permutation__round__n2347 ), .Z(_f_permutation__round__c[775] ) );
  XOR2_X2 _f_permutation__round__U4625  ( .A(SYNOPSYS_UNCONNECTED_184), .B(
        _f_permutation__round__n2346 ), .Z(_f_permutation__round__c[136] ) );
  XOR2_X2 _f_permutation__round__U4624  ( .A(_f_permutation__round_in[1095]), 
        .B(_f_permutation__round__n2347 ), .Z(_f_permutation__round__c[711] )
         );
  XOR2_X2 _f_permutation__round__U4623  ( .A(_f_permutation__round_in[1224]), 
        .B(_f_permutation__round__n2346 ), .Z(_f_permutation__round__c[72] )
         );
  XOR2_X2 _f_permutation__round__U4622  ( .A(_f_permutation__round_in[1415]), 
        .B(_f_permutation__round__n2347 ), .Z(_f_permutation__round__c[647] )
         );
  XOR2_X2 _f_permutation__round__U4621  ( .A(_f_permutation__round__n2349 ), 
        .B(_f_permutation__round__n2348 ), .Z(_f_permutation__round__n2351 )
         );
  XOR2_X2 _f_permutation__round__U4620  ( .A(SYNOPSYS_UNCONNECTED_954), .B(
        _f_permutation__round__n2351 ), .Z(_f_permutation__round__c[902] ) );
  XOR2_X2 _f_permutation__round__U4619  ( .A(SYNOPSYS_UNCONNECTED_825), .B(
        _f_permutation__round__n2350 ), .Z(_f_permutation__round__c[263] ) );
  XOR2_X2 _f_permutation__round__U4618  ( .A(SYNOPSYS_UNCONNECTED_634), .B(
        _f_permutation__round__n2351 ), .Z(_f_permutation__round__c[838] ) );
  XOR2_X2 _f_permutation__round__U4617  ( .A(SYNOPSYS_UNCONNECTED_505), .B(
        _f_permutation__round__n2350 ), .Z(_f_permutation__round__c[199] ) );
  XOR2_X2 _f_permutation__round__U4616  ( .A(SYNOPSYS_UNCONNECTED_314), .B(
        _f_permutation__round__n2351 ), .Z(_f_permutation__round__c[774] ) );
  XOR2_X2 _f_permutation__round__U4615  ( .A(SYNOPSYS_UNCONNECTED_185), .B(
        _f_permutation__round__n2350 ), .Z(_f_permutation__round__c[135] ) );
  XOR2_X2 _f_permutation__round__U4614  ( .A(_f_permutation__round_in[1094]), 
        .B(_f_permutation__round__n2351 ), .Z(_f_permutation__round__c[710] )
         );
  XOR2_X2 _f_permutation__round__U4613  ( .A(_f_permutation__round_in[1223]), 
        .B(_f_permutation__round__n2350 ), .Z(_f_permutation__round__c[71] )
         );
  XOR2_X2 _f_permutation__round__U4612  ( .A(_f_permutation__round_in[1414]), 
        .B(_f_permutation__round__n2351 ), .Z(_f_permutation__round__c[646] )
         );
  XOR2_X2 _f_permutation__round__U4611  ( .A(_f_permutation__round__n2353 ), 
        .B(_f_permutation__round__n2352 ), .Z(_f_permutation__round__n2355 )
         );
  XOR2_X2 _f_permutation__round__U4610  ( .A(SYNOPSYS_UNCONNECTED_955), .B(
        _f_permutation__round__n2355 ), .Z(_f_permutation__round__c[901] ) );
  XOR2_X2 _f_permutation__round__U4609  ( .A(SYNOPSYS_UNCONNECTED_826), .B(
        _f_permutation__round__n2354 ), .Z(_f_permutation__round__c[262] ) );
  XOR2_X2 _f_permutation__round__U4608  ( .A(SYNOPSYS_UNCONNECTED_635), .B(
        _f_permutation__round__n2355 ), .Z(_f_permutation__round__c[837] ) );
  XOR2_X2 _f_permutation__round__U4607  ( .A(SYNOPSYS_UNCONNECTED_506), .B(
        _f_permutation__round__n2354 ), .Z(_f_permutation__round__c[198] ) );
  XOR2_X2 _f_permutation__round__U4606  ( .A(SYNOPSYS_UNCONNECTED_315), .B(
        _f_permutation__round__n2355 ), .Z(_f_permutation__round__c[773] ) );
  XOR2_X2 _f_permutation__round__U4605  ( .A(SYNOPSYS_UNCONNECTED_186), .B(
        _f_permutation__round__n2354 ), .Z(_f_permutation__round__c[134] ) );
  XOR2_X2 _f_permutation__round__U4604  ( .A(_f_permutation__round_in[1093]), 
        .B(_f_permutation__round__n2355 ), .Z(_f_permutation__round__c[709] )
         );
  XOR2_X2 _f_permutation__round__U4603  ( .A(_f_permutation__round_in[1222]), 
        .B(_f_permutation__round__n2354 ), .Z(_f_permutation__round__c[70] )
         );
  XOR2_X2 _f_permutation__round__U4602  ( .A(_f_permutation__round_in[1413]), 
        .B(_f_permutation__round__n2355 ), .Z(_f_permutation__round__c[645] )
         );
  XOR2_X2 _f_permutation__round__U4601  ( .A(_f_permutation__round__n2357 ), 
        .B(_f_permutation__round__n2356 ), .Z(_f_permutation__round__n2359 )
         );
  XOR2_X2 _f_permutation__round__U4600  ( .A(SYNOPSYS_UNCONNECTED_956), .B(
        _f_permutation__round__n2359 ), .Z(_f_permutation__round__c[900] ) );
  XOR2_X2 _f_permutation__round__U4599  ( .A(SYNOPSYS_UNCONNECTED_827), .B(
        _f_permutation__round__n2358 ), .Z(_f_permutation__round__c[261] ) );
  XOR2_X2 _f_permutation__round__U4598  ( .A(SYNOPSYS_UNCONNECTED_636), .B(
        _f_permutation__round__n2359 ), .Z(_f_permutation__round__c[836] ) );
  XOR2_X2 _f_permutation__round__U4597  ( .A(SYNOPSYS_UNCONNECTED_507), .B(
        _f_permutation__round__n2358 ), .Z(_f_permutation__round__c[197] ) );
  XOR2_X2 _f_permutation__round__U4596  ( .A(SYNOPSYS_UNCONNECTED_316), .B(
        _f_permutation__round__n2359 ), .Z(_f_permutation__round__c[772] ) );
  XOR2_X2 _f_permutation__round__U4595  ( .A(SYNOPSYS_UNCONNECTED_187), .B(
        _f_permutation__round__n2358 ), .Z(_f_permutation__round__c[133] ) );
  XOR2_X2 _f_permutation__round__U4594  ( .A(_f_permutation__round_in[1092]), 
        .B(_f_permutation__round__n2359 ), .Z(_f_permutation__round__c[708] )
         );
  XOR2_X2 _f_permutation__round__U4593  ( .A(_f_permutation__round_in[1221]), 
        .B(_f_permutation__round__n2358 ), .Z(_f_permutation__round__c[69] )
         );
  XOR2_X2 _f_permutation__round__U4592  ( .A(_f_permutation__round_in[1412]), 
        .B(_f_permutation__round__n2359 ), .Z(_f_permutation__round__c[644] )
         );
  XOR2_X2 _f_permutation__round__U4591  ( .A(_f_permutation__round__n2361 ), 
        .B(_f_permutation__round__n2360 ), .Z(_f_permutation__round__n2363 )
         );
  XOR2_X2 _f_permutation__round__U4590  ( .A(SYNOPSYS_UNCONNECTED_957), .B(
        _f_permutation__round__n2363 ), .Z(_f_permutation__round__c[899] ) );
  XOR2_X2 _f_permutation__round__U4589  ( .A(SYNOPSYS_UNCONNECTED_828), .B(
        _f_permutation__round__n2362 ), .Z(_f_permutation__round__c[260] ) );
  XOR2_X2 _f_permutation__round__U4588  ( .A(SYNOPSYS_UNCONNECTED_637), .B(
        _f_permutation__round__n2363 ), .Z(_f_permutation__round__c[835] ) );
  XOR2_X2 _f_permutation__round__U4587  ( .A(SYNOPSYS_UNCONNECTED_508), .B(
        _f_permutation__round__n2362 ), .Z(_f_permutation__round__c[196] ) );
  XOR2_X2 _f_permutation__round__U4586  ( .A(SYNOPSYS_UNCONNECTED_317), .B(
        _f_permutation__round__n2363 ), .Z(_f_permutation__round__c[771] ) );
  XOR2_X2 _f_permutation__round__U4585  ( .A(SYNOPSYS_UNCONNECTED_188), .B(
        _f_permutation__round__n2362 ), .Z(_f_permutation__round__c[132] ) );
  XOR2_X2 _f_permutation__round__U4584  ( .A(_f_permutation__round_in[1091]), 
        .B(_f_permutation__round__n2363 ), .Z(_f_permutation__round__c[707] )
         );
  XOR2_X2 _f_permutation__round__U4583  ( .A(_f_permutation__round_in[1220]), 
        .B(_f_permutation__round__n2362 ), .Z(_f_permutation__round__c[68] )
         );
  XOR2_X2 _f_permutation__round__U4582  ( .A(_f_permutation__round_in[1411]), 
        .B(_f_permutation__round__n2363 ), .Z(_f_permutation__round__c[643] )
         );
  XOR2_X2 _f_permutation__round__U4581  ( .A(_f_permutation__round__n2365 ), 
        .B(_f_permutation__round__n2364 ), .Z(_f_permutation__round__n2367 )
         );
  XOR2_X2 _f_permutation__round__U4580  ( .A(SYNOPSYS_UNCONNECTED_958), .B(
        _f_permutation__round__n2367 ), .Z(_f_permutation__round__c[898] ) );
  XOR2_X2 _f_permutation__round__U4579  ( .A(SYNOPSYS_UNCONNECTED_829), .B(
        _f_permutation__round__n2366 ), .Z(_f_permutation__round__c[259] ) );
  XOR2_X2 _f_permutation__round__U4578  ( .A(SYNOPSYS_UNCONNECTED_638), .B(
        _f_permutation__round__n2367 ), .Z(_f_permutation__round__c[834] ) );
  XOR2_X2 _f_permutation__round__U4577  ( .A(SYNOPSYS_UNCONNECTED_509), .B(
        _f_permutation__round__n2366 ), .Z(_f_permutation__round__c[195] ) );
  XOR2_X2 _f_permutation__round__U4576  ( .A(SYNOPSYS_UNCONNECTED_318), .B(
        _f_permutation__round__n2367 ), .Z(_f_permutation__round__c[770] ) );
  XOR2_X2 _f_permutation__round__U4575  ( .A(SYNOPSYS_UNCONNECTED_189), .B(
        _f_permutation__round__n2366 ), .Z(_f_permutation__round__c[131] ) );
  XOR2_X2 _f_permutation__round__U4574  ( .A(_f_permutation__round_in[1090]), 
        .B(_f_permutation__round__n2367 ), .Z(_f_permutation__round__c[706] )
         );
  XOR2_X2 _f_permutation__round__U4573  ( .A(_f_permutation__round_in[1219]), 
        .B(_f_permutation__round__n2366 ), .Z(_f_permutation__round__c[67] )
         );
  XOR2_X2 _f_permutation__round__U4572  ( .A(_f_permutation__round_in[1410]), 
        .B(_f_permutation__round__n2367 ), .Z(_f_permutation__round__c[642] )
         );
  XOR2_X2 _f_permutation__round__U4571  ( .A(_f_permutation__round__n2369 ), 
        .B(_f_permutation__round__n2368 ), .Z(_f_permutation__round__n2371 )
         );
  XOR2_X2 _f_permutation__round__U4570  ( .A(SYNOPSYS_UNCONNECTED_959), .B(
        _f_permutation__round__n2371 ), .Z(_f_permutation__round__c[897] ) );
  XOR2_X2 _f_permutation__round__U4569  ( .A(SYNOPSYS_UNCONNECTED_830), .B(
        _f_permutation__round__n2370 ), .Z(_f_permutation__round__c[258] ) );
  XOR2_X2 _f_permutation__round__U4568  ( .A(SYNOPSYS_UNCONNECTED_639), .B(
        _f_permutation__round__n2371 ), .Z(_f_permutation__round__c[833] ) );
  XOR2_X2 _f_permutation__round__U4567  ( .A(SYNOPSYS_UNCONNECTED_510), .B(
        _f_permutation__round__n2370 ), .Z(_f_permutation__round__c[194] ) );
  XOR2_X2 _f_permutation__round__U4566  ( .A(SYNOPSYS_UNCONNECTED_319), .B(
        _f_permutation__round__n2371 ), .Z(_f_permutation__round__c[769] ) );
  XOR2_X2 _f_permutation__round__U4565  ( .A(SYNOPSYS_UNCONNECTED_190), .B(
        _f_permutation__round__n2370 ), .Z(_f_permutation__round__c[130] ) );
  XOR2_X2 _f_permutation__round__U4564  ( .A(_f_permutation__round_in[1089]), 
        .B(_f_permutation__round__n2371 ), .Z(_f_permutation__round__c[705] )
         );
  XOR2_X2 _f_permutation__round__U4563  ( .A(_f_permutation__round_in[1218]), 
        .B(_f_permutation__round__n2370 ), .Z(_f_permutation__round__c[66] )
         );
  XOR2_X2 _f_permutation__round__U4562  ( .A(_f_permutation__round_in[1409]), 
        .B(_f_permutation__round__n2371 ), .Z(_f_permutation__round__c[641] )
         );
  XOR2_X2 _f_permutation__round__U4561  ( .A(_f_permutation__round__n2373 ), 
        .B(_f_permutation__round__n2372 ), .Z(_f_permutation__round__n2375 )
         );
  XOR2_X2 _f_permutation__round__U4560  ( .A(SYNOPSYS_UNCONNECTED_960), .B(
        _f_permutation__round__n2375 ), .Z(_f_permutation__round__c[896] ) );
  XOR2_X2 _f_permutation__round__U4559  ( .A(SYNOPSYS_UNCONNECTED_831), .B(
        _f_permutation__round__n2374 ), .Z(_f_permutation__round__c[257] ) );
  XOR2_X2 _f_permutation__round__U4558  ( .A(SYNOPSYS_UNCONNECTED_640), .B(
        _f_permutation__round__n2375 ), .Z(_f_permutation__round__c[832] ) );
  XOR2_X2 _f_permutation__round__U4557  ( .A(SYNOPSYS_UNCONNECTED_511), .B(
        _f_permutation__round__n2374 ), .Z(_f_permutation__round__c[193] ) );
  XOR2_X2 _f_permutation__round__U4556  ( .A(SYNOPSYS_UNCONNECTED_320), .B(
        _f_permutation__round__n2375 ), .Z(_f_permutation__round__c[768] ) );
  XOR2_X2 _f_permutation__round__U4555  ( .A(SYNOPSYS_UNCONNECTED_191), .B(
        _f_permutation__round__n2374 ), .Z(_f_permutation__round__c[129] ) );
  XOR2_X2 _f_permutation__round__U4554  ( .A(_f_permutation__round_in[1088]), 
        .B(_f_permutation__round__n2375 ), .Z(_f_permutation__round__c[704] )
         );
  XOR2_X2 _f_permutation__round__U4553  ( .A(_f_permutation__round_in[1217]), 
        .B(_f_permutation__round__n2374 ), .Z(_f_permutation__round__c[65] )
         );
  XOR2_X2 _f_permutation__round__U4552  ( .A(_f_permutation__round_in[1408]), 
        .B(_f_permutation__round__n2375 ), .Z(_f_permutation__round__c[640] )
         );
  XOR2_X2 _f_permutation__round__U4551  ( .A(_f_permutation__round__n2377 ), 
        .B(_f_permutation__round__n2376 ), .Z(_f_permutation__round__n2378 )
         );
  XOR2_X2 _f_permutation__round__U4550  ( .A(SYNOPSYS_UNCONNECTED_961), .B(
        _f_permutation__round__n2378 ), .Z(_f_permutation__round__c[1279] ) );
  XOR2_X2 _f_permutation__round__U4549  ( .A(SYNOPSYS_UNCONNECTED_641), .B(
        _f_permutation__round__n2378 ), .Z(_f_permutation__round__c[1215] ) );
  XOR2_X2 _f_permutation__round__U4548  ( .A(SYNOPSYS_UNCONNECTED_321), .B(
        _f_permutation__round__n2378 ), .Z(_f_permutation__round__c[1151] ) );
  XOR2_X2 _f_permutation__round__U4547  ( .A(_f_permutation__round_in[1087]), 
        .B(_f_permutation__round__n2378 ), .Z(_f_permutation__round__c[1087] )
         );
  XOR2_X2 _f_permutation__round__U4546  ( .A(_f_permutation__round_in[1407]), 
        .B(_f_permutation__round__n2378 ), .Z(_f_permutation__round__c[1023] )
         );
  XOR2_X2 _f_permutation__round__U4545  ( .A(_f_permutation__round__n2380 ), 
        .B(_f_permutation__round__n2379 ), .Z(_f_permutation__round__n2381 )
         );
  XOR2_X2 _f_permutation__round__U4544  ( .A(SYNOPSYS_UNCONNECTED_962), .B(
        _f_permutation__round__n2381 ), .Z(_f_permutation__round__c[1278] ) );
  XOR2_X2 _f_permutation__round__U4543  ( .A(SYNOPSYS_UNCONNECTED_642), .B(
        _f_permutation__round__n2381 ), .Z(_f_permutation__round__c[1214] ) );
  XOR2_X2 _f_permutation__round__U4542  ( .A(SYNOPSYS_UNCONNECTED_322), .B(
        _f_permutation__round__n2381 ), .Z(_f_permutation__round__c[1150] ) );
  XOR2_X2 _f_permutation__round__U4541  ( .A(_f_permutation__round_in[1086]), 
        .B(_f_permutation__round__n2381 ), .Z(_f_permutation__round__c[1086] )
         );
  XOR2_X2 _f_permutation__round__U4540  ( .A(_f_permutation__round_in[1406]), 
        .B(_f_permutation__round__n2381 ), .Z(_f_permutation__round__c[1022] )
         );
  XOR2_X2 _f_permutation__round__U4539  ( .A(_f_permutation__round__n2383 ), 
        .B(_f_permutation__round__n2382 ), .Z(_f_permutation__round__n2384 )
         );
  XOR2_X2 _f_permutation__round__U4538  ( .A(SYNOPSYS_UNCONNECTED_963), .B(
        _f_permutation__round__n2384 ), .Z(_f_permutation__round__c[1277] ) );
  XOR2_X2 _f_permutation__round__U4537  ( .A(SYNOPSYS_UNCONNECTED_643), .B(
        _f_permutation__round__n2384 ), .Z(_f_permutation__round__c[1213] ) );
  XOR2_X2 _f_permutation__round__U4536  ( .A(SYNOPSYS_UNCONNECTED_323), .B(
        _f_permutation__round__n2384 ), .Z(_f_permutation__round__c[1149] ) );
  XOR2_X2 _f_permutation__round__U4535  ( .A(_f_permutation__round_in[1085]), 
        .B(_f_permutation__round__n2384 ), .Z(_f_permutation__round__c[1085] )
         );
  XOR2_X2 _f_permutation__round__U4534  ( .A(_f_permutation__round_in[1405]), 
        .B(_f_permutation__round__n2384 ), .Z(_f_permutation__round__c[1021] )
         );
  XOR2_X2 _f_permutation__round__U4533  ( .A(_f_permutation__round__n2386 ), 
        .B(_f_permutation__round__n2385 ), .Z(_f_permutation__round__n2387 )
         );
  XOR2_X2 _f_permutation__round__U4532  ( .A(SYNOPSYS_UNCONNECTED_964), .B(
        _f_permutation__round__n2387 ), .Z(_f_permutation__round__c[1276] ) );
  XOR2_X2 _f_permutation__round__U4531  ( .A(SYNOPSYS_UNCONNECTED_644), .B(
        _f_permutation__round__n2387 ), .Z(_f_permutation__round__c[1212] ) );
  XOR2_X2 _f_permutation__round__U4530  ( .A(SYNOPSYS_UNCONNECTED_324), .B(
        _f_permutation__round__n2387 ), .Z(_f_permutation__round__c[1148] ) );
  XOR2_X2 _f_permutation__round__U4529  ( .A(_f_permutation__round_in[1084]), 
        .B(_f_permutation__round__n2387 ), .Z(_f_permutation__round__c[1084] )
         );
  XOR2_X2 _f_permutation__round__U4528  ( .A(_f_permutation__round_in[1404]), 
        .B(_f_permutation__round__n2387 ), .Z(_f_permutation__round__c[1020] )
         );
  XOR2_X2 _f_permutation__round__U4527  ( .A(_f_permutation__round__n2389 ), 
        .B(_f_permutation__round__n2388 ), .Z(_f_permutation__round__n2390 )
         );
  XOR2_X2 _f_permutation__round__U4526  ( .A(SYNOPSYS_UNCONNECTED_965), .B(
        _f_permutation__round__n2390 ), .Z(_f_permutation__round__c[1275] ) );
  XOR2_X2 _f_permutation__round__U4525  ( .A(SYNOPSYS_UNCONNECTED_645), .B(
        _f_permutation__round__n2390 ), .Z(_f_permutation__round__c[1211] ) );
  XOR2_X2 _f_permutation__round__U4524  ( .A(SYNOPSYS_UNCONNECTED_325), .B(
        _f_permutation__round__n2390 ), .Z(_f_permutation__round__c[1147] ) );
  XOR2_X2 _f_permutation__round__U4523  ( .A(_f_permutation__round_in[1083]), 
        .B(_f_permutation__round__n2390 ), .Z(_f_permutation__round__c[1083] )
         );
  XOR2_X2 _f_permutation__round__U4522  ( .A(_f_permutation__round_in[1403]), 
        .B(_f_permutation__round__n2390 ), .Z(_f_permutation__round__c[1019] )
         );
  XOR2_X2 _f_permutation__round__U4521  ( .A(_f_permutation__round__n2392 ), 
        .B(_f_permutation__round__n2391 ), .Z(_f_permutation__round__n2393 )
         );
  XOR2_X2 _f_permutation__round__U4520  ( .A(SYNOPSYS_UNCONNECTED_966), .B(
        _f_permutation__round__n2393 ), .Z(_f_permutation__round__c[1274] ) );
  XOR2_X2 _f_permutation__round__U4519  ( .A(SYNOPSYS_UNCONNECTED_646), .B(
        _f_permutation__round__n2393 ), .Z(_f_permutation__round__c[1210] ) );
  XOR2_X2 _f_permutation__round__U4518  ( .A(SYNOPSYS_UNCONNECTED_326), .B(
        _f_permutation__round__n2393 ), .Z(_f_permutation__round__c[1146] ) );
  XOR2_X2 _f_permutation__round__U4517  ( .A(_f_permutation__round_in[1082]), 
        .B(_f_permutation__round__n2393 ), .Z(_f_permutation__round__c[1082] )
         );
  XOR2_X2 _f_permutation__round__U4516  ( .A(_f_permutation__round_in[1402]), 
        .B(_f_permutation__round__n2393 ), .Z(_f_permutation__round__c[1018] )
         );
  XOR2_X2 _f_permutation__round__U4515  ( .A(_f_permutation__round__n2395 ), 
        .B(_f_permutation__round__n2394 ), .Z(_f_permutation__round__n2396 )
         );
  XOR2_X2 _f_permutation__round__U4514  ( .A(SYNOPSYS_UNCONNECTED_967), .B(
        _f_permutation__round__n2396 ), .Z(_f_permutation__round__c[1273] ) );
  XOR2_X2 _f_permutation__round__U4513  ( .A(SYNOPSYS_UNCONNECTED_647), .B(
        _f_permutation__round__n2396 ), .Z(_f_permutation__round__c[1209] ) );
  XOR2_X2 _f_permutation__round__U4512  ( .A(SYNOPSYS_UNCONNECTED_327), .B(
        _f_permutation__round__n2396 ), .Z(_f_permutation__round__c[1145] ) );
  XOR2_X2 _f_permutation__round__U4511  ( .A(_f_permutation__round_in[1081]), 
        .B(_f_permutation__round__n2396 ), .Z(_f_permutation__round__c[1081] )
         );
  XOR2_X2 _f_permutation__round__U4510  ( .A(_f_permutation__round_in[1401]), 
        .B(_f_permutation__round__n2396 ), .Z(_f_permutation__round__c[1017] )
         );
  XOR2_X2 _f_permutation__round__U4509  ( .A(_f_permutation__round__n2398 ), 
        .B(_f_permutation__round__n2397 ), .Z(_f_permutation__round__n2399 )
         );
  XOR2_X2 _f_permutation__round__U4508  ( .A(SYNOPSYS_UNCONNECTED_968), .B(
        _f_permutation__round__n2399 ), .Z(_f_permutation__round__c[1272] ) );
  XOR2_X2 _f_permutation__round__U4507  ( .A(SYNOPSYS_UNCONNECTED_648), .B(
        _f_permutation__round__n2399 ), .Z(_f_permutation__round__c[1208] ) );
  XOR2_X2 _f_permutation__round__U4506  ( .A(SYNOPSYS_UNCONNECTED_328), .B(
        _f_permutation__round__n2399 ), .Z(_f_permutation__round__c[1144] ) );
  XOR2_X2 _f_permutation__round__U4505  ( .A(_f_permutation__round_in[1080]), 
        .B(_f_permutation__round__n2399 ), .Z(_f_permutation__round__c[1080] )
         );
  XOR2_X2 _f_permutation__round__U4504  ( .A(_f_permutation__round_in[1400]), 
        .B(_f_permutation__round__n2399 ), .Z(_f_permutation__round__c[1016] )
         );
  XOR2_X2 _f_permutation__round__U4503  ( .A(_f_permutation__round__n2401 ), 
        .B(_f_permutation__round__n2400 ), .Z(_f_permutation__round__n2402 )
         );
  XOR2_X2 _f_permutation__round__U4502  ( .A(SYNOPSYS_UNCONNECTED_969), .B(
        _f_permutation__round__n2402 ), .Z(_f_permutation__round__c[1271] ) );
  XOR2_X2 _f_permutation__round__U4501  ( .A(SYNOPSYS_UNCONNECTED_649), .B(
        _f_permutation__round__n2402 ), .Z(_f_permutation__round__c[1207] ) );
  XOR2_X2 _f_permutation__round__U4500  ( .A(SYNOPSYS_UNCONNECTED_329), .B(
        _f_permutation__round__n2402 ), .Z(_f_permutation__round__c[1143] ) );
  XOR2_X2 _f_permutation__round__U4499  ( .A(_f_permutation__round_in[1079]), 
        .B(_f_permutation__round__n2402 ), .Z(_f_permutation__round__c[1079] )
         );
  XOR2_X2 _f_permutation__round__U4498  ( .A(_f_permutation__round_in[1399]), 
        .B(_f_permutation__round__n2402 ), .Z(_f_permutation__round__c[1015] )
         );
  XOR2_X2 _f_permutation__round__U4497  ( .A(_f_permutation__round__n2404 ), 
        .B(_f_permutation__round__n2403 ), .Z(_f_permutation__round__n2405 )
         );
  XOR2_X2 _f_permutation__round__U4496  ( .A(SYNOPSYS_UNCONNECTED_970), .B(
        _f_permutation__round__n2405 ), .Z(_f_permutation__round__c[1270] ) );
  XOR2_X2 _f_permutation__round__U4495  ( .A(SYNOPSYS_UNCONNECTED_650), .B(
        _f_permutation__round__n2405 ), .Z(_f_permutation__round__c[1206] ) );
  XOR2_X2 _f_permutation__round__U4494  ( .A(SYNOPSYS_UNCONNECTED_330), .B(
        _f_permutation__round__n2405 ), .Z(_f_permutation__round__c[1142] ) );
  XOR2_X2 _f_permutation__round__U4493  ( .A(_f_permutation__round_in[1078]), 
        .B(_f_permutation__round__n2405 ), .Z(_f_permutation__round__c[1078] )
         );
  XOR2_X2 _f_permutation__round__U4492  ( .A(_f_permutation__round_in[1398]), 
        .B(_f_permutation__round__n2405 ), .Z(_f_permutation__round__c[1014] )
         );
  XOR2_X2 _f_permutation__round__U4491  ( .A(_f_permutation__round__n2407 ), 
        .B(_f_permutation__round__n2406 ), .Z(_f_permutation__round__n2408 )
         );
  XOR2_X2 _f_permutation__round__U4490  ( .A(SYNOPSYS_UNCONNECTED_971), .B(
        _f_permutation__round__n2408 ), .Z(_f_permutation__round__c[1269] ) );
  XOR2_X2 _f_permutation__round__U4489  ( .A(SYNOPSYS_UNCONNECTED_651), .B(
        _f_permutation__round__n2408 ), .Z(_f_permutation__round__c[1205] ) );
  XOR2_X2 _f_permutation__round__U4488  ( .A(SYNOPSYS_UNCONNECTED_331), .B(
        _f_permutation__round__n2408 ), .Z(_f_permutation__round__c[1141] ) );
  XOR2_X2 _f_permutation__round__U4487  ( .A(_f_permutation__round_in[1077]), 
        .B(_f_permutation__round__n2408 ), .Z(_f_permutation__round__c[1077] )
         );
  XOR2_X2 _f_permutation__round__U4486  ( .A(_f_permutation__round_in[1397]), 
        .B(_f_permutation__round__n2408 ), .Z(_f_permutation__round__c[1013] )
         );
  XOR2_X2 _f_permutation__round__U4485  ( .A(_f_permutation__round__n2410 ), 
        .B(_f_permutation__round__n2409 ), .Z(_f_permutation__round__n2411 )
         );
  XOR2_X2 _f_permutation__round__U4484  ( .A(SYNOPSYS_UNCONNECTED_972), .B(
        _f_permutation__round__n2411 ), .Z(_f_permutation__round__c[1268] ) );
  XOR2_X2 _f_permutation__round__U4483  ( .A(SYNOPSYS_UNCONNECTED_652), .B(
        _f_permutation__round__n2411 ), .Z(_f_permutation__round__c[1204] ) );
  XOR2_X2 _f_permutation__round__U4482  ( .A(SYNOPSYS_UNCONNECTED_332), .B(
        _f_permutation__round__n2411 ), .Z(_f_permutation__round__c[1140] ) );
  XOR2_X2 _f_permutation__round__U4481  ( .A(_f_permutation__round_in[1076]), 
        .B(_f_permutation__round__n2411 ), .Z(_f_permutation__round__c[1076] )
         );
  XOR2_X2 _f_permutation__round__U4480  ( .A(_f_permutation__round_in[1396]), 
        .B(_f_permutation__round__n2411 ), .Z(_f_permutation__round__c[1012] )
         );
  XOR2_X2 _f_permutation__round__U4479  ( .A(_f_permutation__round__n2413 ), 
        .B(_f_permutation__round__n2412 ), .Z(_f_permutation__round__n2414 )
         );
  XOR2_X2 _f_permutation__round__U4478  ( .A(SYNOPSYS_UNCONNECTED_973), .B(
        _f_permutation__round__n2414 ), .Z(_f_permutation__round__c[1267] ) );
  XOR2_X2 _f_permutation__round__U4477  ( .A(SYNOPSYS_UNCONNECTED_653), .B(
        _f_permutation__round__n2414 ), .Z(_f_permutation__round__c[1203] ) );
  XOR2_X2 _f_permutation__round__U4476  ( .A(SYNOPSYS_UNCONNECTED_333), .B(
        _f_permutation__round__n2414 ), .Z(_f_permutation__round__c[1139] ) );
  XOR2_X2 _f_permutation__round__U4475  ( .A(_f_permutation__round_in[1075]), 
        .B(_f_permutation__round__n2414 ), .Z(_f_permutation__round__c[1075] )
         );
  XOR2_X2 _f_permutation__round__U4474  ( .A(_f_permutation__round_in[1395]), 
        .B(_f_permutation__round__n2414 ), .Z(_f_permutation__round__c[1011] )
         );
  XOR2_X2 _f_permutation__round__U4473  ( .A(_f_permutation__round__n2416 ), 
        .B(_f_permutation__round__n2415 ), .Z(_f_permutation__round__n2417 )
         );
  XOR2_X2 _f_permutation__round__U4472  ( .A(SYNOPSYS_UNCONNECTED_974), .B(
        _f_permutation__round__n2417 ), .Z(_f_permutation__round__c[1266] ) );
  XOR2_X2 _f_permutation__round__U4471  ( .A(SYNOPSYS_UNCONNECTED_654), .B(
        _f_permutation__round__n2417 ), .Z(_f_permutation__round__c[1202] ) );
  XOR2_X2 _f_permutation__round__U4470  ( .A(SYNOPSYS_UNCONNECTED_334), .B(
        _f_permutation__round__n2417 ), .Z(_f_permutation__round__c[1138] ) );
  XOR2_X2 _f_permutation__round__U4469  ( .A(_f_permutation__round_in[1074]), 
        .B(_f_permutation__round__n2417 ), .Z(_f_permutation__round__c[1074] )
         );
  XOR2_X2 _f_permutation__round__U4468  ( .A(_f_permutation__round_in[1394]), 
        .B(_f_permutation__round__n2417 ), .Z(_f_permutation__round__c[1010] )
         );
  XOR2_X2 _f_permutation__round__U4467  ( .A(_f_permutation__round__n2419 ), 
        .B(_f_permutation__round__n2418 ), .Z(_f_permutation__round__n2420 )
         );
  XOR2_X2 _f_permutation__round__U4466  ( .A(SYNOPSYS_UNCONNECTED_975), .B(
        _f_permutation__round__n2420 ), .Z(_f_permutation__round__c[1265] ) );
  XOR2_X2 _f_permutation__round__U4465  ( .A(SYNOPSYS_UNCONNECTED_655), .B(
        _f_permutation__round__n2420 ), .Z(_f_permutation__round__c[1201] ) );
  XOR2_X2 _f_permutation__round__U4464  ( .A(SYNOPSYS_UNCONNECTED_335), .B(
        _f_permutation__round__n2420 ), .Z(_f_permutation__round__c[1137] ) );
  XOR2_X2 _f_permutation__round__U4463  ( .A(_f_permutation__round_in[1073]), 
        .B(_f_permutation__round__n2420 ), .Z(_f_permutation__round__c[1073] )
         );
  XOR2_X2 _f_permutation__round__U4462  ( .A(_f_permutation__round_in[1393]), 
        .B(_f_permutation__round__n2420 ), .Z(_f_permutation__round__c[1009] )
         );
  XOR2_X2 _f_permutation__round__U4461  ( .A(_f_permutation__round__n2422 ), 
        .B(_f_permutation__round__n2421 ), .Z(_f_permutation__round__n2423 )
         );
  XOR2_X2 _f_permutation__round__U4460  ( .A(SYNOPSYS_UNCONNECTED_976), .B(
        _f_permutation__round__n2423 ), .Z(_f_permutation__round__c[1264] ) );
  XOR2_X2 _f_permutation__round__U4459  ( .A(SYNOPSYS_UNCONNECTED_656), .B(
        _f_permutation__round__n2423 ), .Z(_f_permutation__round__c[1200] ) );
  XOR2_X2 _f_permutation__round__U4458  ( .A(SYNOPSYS_UNCONNECTED_336), .B(
        _f_permutation__round__n2423 ), .Z(_f_permutation__round__c[1136] ) );
  XOR2_X2 _f_permutation__round__U4457  ( .A(_f_permutation__round_in[1072]), 
        .B(_f_permutation__round__n2423 ), .Z(_f_permutation__round__c[1072] )
         );
  XOR2_X2 _f_permutation__round__U4456  ( .A(_f_permutation__round_in[1392]), 
        .B(_f_permutation__round__n2423 ), .Z(_f_permutation__round__c[1008] )
         );
  XOR2_X2 _f_permutation__round__U4455  ( .A(_f_permutation__round__n2425 ), 
        .B(_f_permutation__round__n2424 ), .Z(_f_permutation__round__n2426 )
         );
  XOR2_X2 _f_permutation__round__U4454  ( .A(SYNOPSYS_UNCONNECTED_977), .B(
        _f_permutation__round__n2426 ), .Z(_f_permutation__round__c[1263] ) );
  XOR2_X2 _f_permutation__round__U4453  ( .A(SYNOPSYS_UNCONNECTED_657), .B(
        _f_permutation__round__n2426 ), .Z(_f_permutation__round__c[1199] ) );
  XOR2_X2 _f_permutation__round__U4452  ( .A(SYNOPSYS_UNCONNECTED_337), .B(
        _f_permutation__round__n2426 ), .Z(_f_permutation__round__c[1135] ) );
  XOR2_X2 _f_permutation__round__U4451  ( .A(_f_permutation__round_in[1071]), 
        .B(_f_permutation__round__n2426 ), .Z(_f_permutation__round__c[1071] )
         );
  XOR2_X2 _f_permutation__round__U4450  ( .A(_f_permutation__round_in[1391]), 
        .B(_f_permutation__round__n2426 ), .Z(_f_permutation__round__c[1007] )
         );
  XOR2_X2 _f_permutation__round__U4449  ( .A(_f_permutation__round__n2428 ), 
        .B(_f_permutation__round__n2427 ), .Z(_f_permutation__round__n2429 )
         );
  XOR2_X2 _f_permutation__round__U4448  ( .A(SYNOPSYS_UNCONNECTED_978), .B(
        _f_permutation__round__n2429 ), .Z(_f_permutation__round__c[1262] ) );
  XOR2_X2 _f_permutation__round__U4447  ( .A(SYNOPSYS_UNCONNECTED_658), .B(
        _f_permutation__round__n2429 ), .Z(_f_permutation__round__c[1198] ) );
  XOR2_X2 _f_permutation__round__U4446  ( .A(SYNOPSYS_UNCONNECTED_338), .B(
        _f_permutation__round__n2429 ), .Z(_f_permutation__round__c[1134] ) );
  XOR2_X2 _f_permutation__round__U4445  ( .A(_f_permutation__round_in[1070]), 
        .B(_f_permutation__round__n2429 ), .Z(_f_permutation__round__c[1070] )
         );
  XOR2_X2 _f_permutation__round__U4444  ( .A(_f_permutation__round_in[1390]), 
        .B(_f_permutation__round__n2429 ), .Z(_f_permutation__round__c[1006] )
         );
  XOR2_X2 _f_permutation__round__U4443  ( .A(_f_permutation__round__n2431 ), 
        .B(_f_permutation__round__n2430 ), .Z(_f_permutation__round__n2432 )
         );
  XOR2_X2 _f_permutation__round__U4442  ( .A(SYNOPSYS_UNCONNECTED_979), .B(
        _f_permutation__round__n2432 ), .Z(_f_permutation__round__c[1261] ) );
  XOR2_X2 _f_permutation__round__U4441  ( .A(SYNOPSYS_UNCONNECTED_659), .B(
        _f_permutation__round__n2432 ), .Z(_f_permutation__round__c[1197] ) );
  XOR2_X2 _f_permutation__round__U4440  ( .A(SYNOPSYS_UNCONNECTED_339), .B(
        _f_permutation__round__n2432 ), .Z(_f_permutation__round__c[1133] ) );
  XOR2_X2 _f_permutation__round__U4439  ( .A(_f_permutation__round_in[1069]), 
        .B(_f_permutation__round__n2432 ), .Z(_f_permutation__round__c[1069] )
         );
  XOR2_X2 _f_permutation__round__U4438  ( .A(_f_permutation__round_in[1389]), 
        .B(_f_permutation__round__n2432 ), .Z(_f_permutation__round__c[1005] )
         );
  XOR2_X2 _f_permutation__round__U4437  ( .A(_f_permutation__round__n2434 ), 
        .B(_f_permutation__round__n2433 ), .Z(_f_permutation__round__n2435 )
         );
  XOR2_X2 _f_permutation__round__U4436  ( .A(SYNOPSYS_UNCONNECTED_980), .B(
        _f_permutation__round__n2435 ), .Z(_f_permutation__round__c[1260] ) );
  XOR2_X2 _f_permutation__round__U4435  ( .A(SYNOPSYS_UNCONNECTED_660), .B(
        _f_permutation__round__n2435 ), .Z(_f_permutation__round__c[1196] ) );
  XOR2_X2 _f_permutation__round__U4434  ( .A(SYNOPSYS_UNCONNECTED_340), .B(
        _f_permutation__round__n2435 ), .Z(_f_permutation__round__c[1132] ) );
  XOR2_X2 _f_permutation__round__U4433  ( .A(_f_permutation__round_in[1068]), 
        .B(_f_permutation__round__n2435 ), .Z(_f_permutation__round__c[1068] )
         );
  XOR2_X2 _f_permutation__round__U4432  ( .A(_f_permutation__round_in[1388]), 
        .B(_f_permutation__round__n2435 ), .Z(_f_permutation__round__c[1004] )
         );
  XOR2_X2 _f_permutation__round__U4431  ( .A(_f_permutation__round__n2437 ), 
        .B(_f_permutation__round__n2436 ), .Z(_f_permutation__round__n2438 )
         );
  XOR2_X2 _f_permutation__round__U4430  ( .A(SYNOPSYS_UNCONNECTED_981), .B(
        _f_permutation__round__n2438 ), .Z(_f_permutation__round__c[1259] ) );
  XOR2_X2 _f_permutation__round__U4429  ( .A(SYNOPSYS_UNCONNECTED_661), .B(
        _f_permutation__round__n2438 ), .Z(_f_permutation__round__c[1195] ) );
  XOR2_X2 _f_permutation__round__U4428  ( .A(SYNOPSYS_UNCONNECTED_341), .B(
        _f_permutation__round__n2438 ), .Z(_f_permutation__round__c[1131] ) );
  XOR2_X2 _f_permutation__round__U4427  ( .A(_f_permutation__round_in[1067]), 
        .B(_f_permutation__round__n2438 ), .Z(_f_permutation__round__c[1067] )
         );
  XOR2_X2 _f_permutation__round__U4426  ( .A(_f_permutation__round_in[1387]), 
        .B(_f_permutation__round__n2438 ), .Z(_f_permutation__round__c[1003] )
         );
  XOR2_X2 _f_permutation__round__U4425  ( .A(_f_permutation__round__n2440 ), 
        .B(_f_permutation__round__n2439 ), .Z(_f_permutation__round__n2441 )
         );
  XOR2_X2 _f_permutation__round__U4424  ( .A(SYNOPSYS_UNCONNECTED_982), .B(
        _f_permutation__round__n2441 ), .Z(_f_permutation__round__c[1258] ) );
  XOR2_X2 _f_permutation__round__U4423  ( .A(SYNOPSYS_UNCONNECTED_662), .B(
        _f_permutation__round__n2441 ), .Z(_f_permutation__round__c[1194] ) );
  XOR2_X2 _f_permutation__round__U4422  ( .A(SYNOPSYS_UNCONNECTED_342), .B(
        _f_permutation__round__n2441 ), .Z(_f_permutation__round__c[1130] ) );
  XOR2_X2 _f_permutation__round__U4421  ( .A(_f_permutation__round_in[1066]), 
        .B(_f_permutation__round__n2441 ), .Z(_f_permutation__round__c[1066] )
         );
  XOR2_X2 _f_permutation__round__U4420  ( .A(_f_permutation__round_in[1386]), 
        .B(_f_permutation__round__n2441 ), .Z(_f_permutation__round__c[1002] )
         );
  XOR2_X2 _f_permutation__round__U4419  ( .A(_f_permutation__round__n2443 ), 
        .B(_f_permutation__round__n2442 ), .Z(_f_permutation__round__n2444 )
         );
  XOR2_X2 _f_permutation__round__U4418  ( .A(SYNOPSYS_UNCONNECTED_983), .B(
        _f_permutation__round__n2444 ), .Z(_f_permutation__round__c[1257] ) );
  XOR2_X2 _f_permutation__round__U4417  ( .A(SYNOPSYS_UNCONNECTED_663), .B(
        _f_permutation__round__n2444 ), .Z(_f_permutation__round__c[1193] ) );
  XOR2_X2 _f_permutation__round__U4416  ( .A(SYNOPSYS_UNCONNECTED_343), .B(
        _f_permutation__round__n2444 ), .Z(_f_permutation__round__c[1129] ) );
  XOR2_X2 _f_permutation__round__U4415  ( .A(_f_permutation__round_in[1065]), 
        .B(_f_permutation__round__n2444 ), .Z(_f_permutation__round__c[1065] )
         );
  XOR2_X2 _f_permutation__round__U4414  ( .A(_f_permutation__round_in[1385]), 
        .B(_f_permutation__round__n2444 ), .Z(_f_permutation__round__c[1001] )
         );
  XOR2_X2 _f_permutation__round__U4413  ( .A(_f_permutation__round__n2446 ), 
        .B(_f_permutation__round__n2445 ), .Z(_f_permutation__round__n2447 )
         );
  XOR2_X2 _f_permutation__round__U4412  ( .A(SYNOPSYS_UNCONNECTED_984), .B(
        _f_permutation__round__n2447 ), .Z(_f_permutation__round__c[1256] ) );
  XOR2_X2 _f_permutation__round__U4411  ( .A(SYNOPSYS_UNCONNECTED_664), .B(
        _f_permutation__round__n2447 ), .Z(_f_permutation__round__c[1192] ) );
  XOR2_X2 _f_permutation__round__U4410  ( .A(SYNOPSYS_UNCONNECTED_344), .B(
        _f_permutation__round__n2447 ), .Z(_f_permutation__round__c[1128] ) );
  XOR2_X2 _f_permutation__round__U4409  ( .A(_f_permutation__round_in[1064]), 
        .B(_f_permutation__round__n2447 ), .Z(_f_permutation__round__c[1064] )
         );
  XOR2_X2 _f_permutation__round__U4408  ( .A(_f_permutation__round_in[1384]), 
        .B(_f_permutation__round__n2447 ), .Z(_f_permutation__round__c[1000] )
         );
  XOR2_X2 _f_permutation__round__U4407  ( .A(_f_permutation__round__n2449 ), 
        .B(_f_permutation__round__n2448 ), .Z(_f_permutation__round__n2450 )
         );
  XOR2_X2 _f_permutation__round__U4406  ( .A(SYNOPSYS_UNCONNECTED_985), .B(
        _f_permutation__round__n2450 ), .Z(_f_permutation__round__c[1255] ) );
  XOR2_X2 _f_permutation__round__U4405  ( .A(SYNOPSYS_UNCONNECTED_665), .B(
        _f_permutation__round__n2450 ), .Z(_f_permutation__round__c[1191] ) );
  XOR2_X2 _f_permutation__round__U4404  ( .A(SYNOPSYS_UNCONNECTED_345), .B(
        _f_permutation__round__n2450 ), .Z(_f_permutation__round__c[1127] ) );
  XOR2_X2 _f_permutation__round__U4403  ( .A(_f_permutation__round_in[1063]), 
        .B(_f_permutation__round__n2450 ), .Z(_f_permutation__round__c[1063] )
         );
  XOR2_X2 _f_permutation__round__U4402  ( .A(_f_permutation__round_in[1383]), 
        .B(_f_permutation__round__n2450 ), .Z(_f_permutation__round__c[999] )
         );
  XOR2_X2 _f_permutation__round__U4401  ( .A(_f_permutation__round__n2452 ), 
        .B(_f_permutation__round__n2451 ), .Z(_f_permutation__round__n2453 )
         );
  XOR2_X2 _f_permutation__round__U4400  ( .A(SYNOPSYS_UNCONNECTED_986), .B(
        _f_permutation__round__n2453 ), .Z(_f_permutation__round__c[1254] ) );
  XOR2_X2 _f_permutation__round__U4399  ( .A(SYNOPSYS_UNCONNECTED_666), .B(
        _f_permutation__round__n2453 ), .Z(_f_permutation__round__c[1190] ) );
  XOR2_X2 _f_permutation__round__U4398  ( .A(SYNOPSYS_UNCONNECTED_346), .B(
        _f_permutation__round__n2453 ), .Z(_f_permutation__round__c[1126] ) );
  XOR2_X2 _f_permutation__round__U4397  ( .A(_f_permutation__round_in[1062]), 
        .B(_f_permutation__round__n2453 ), .Z(_f_permutation__round__c[1062] )
         );
  XOR2_X2 _f_permutation__round__U4396  ( .A(_f_permutation__round_in[1382]), 
        .B(_f_permutation__round__n2453 ), .Z(_f_permutation__round__c[998] )
         );
  XOR2_X2 _f_permutation__round__U4395  ( .A(_f_permutation__round__n2455 ), 
        .B(_f_permutation__round__n2454 ), .Z(_f_permutation__round__n2456 )
         );
  XOR2_X2 _f_permutation__round__U4394  ( .A(SYNOPSYS_UNCONNECTED_987), .B(
        _f_permutation__round__n2456 ), .Z(_f_permutation__round__c[1253] ) );
  XOR2_X2 _f_permutation__round__U4393  ( .A(SYNOPSYS_UNCONNECTED_667), .B(
        _f_permutation__round__n2456 ), .Z(_f_permutation__round__c[1189] ) );
  XOR2_X2 _f_permutation__round__U4392  ( .A(SYNOPSYS_UNCONNECTED_347), .B(
        _f_permutation__round__n2456 ), .Z(_f_permutation__round__c[1125] ) );
  XOR2_X2 _f_permutation__round__U4391  ( .A(_f_permutation__round_in[1061]), 
        .B(_f_permutation__round__n2456 ), .Z(_f_permutation__round__c[1061] )
         );
  XOR2_X2 _f_permutation__round__U4390  ( .A(_f_permutation__round_in[1381]), 
        .B(_f_permutation__round__n2456 ), .Z(_f_permutation__round__c[997] )
         );
  XOR2_X2 _f_permutation__round__U4389  ( .A(_f_permutation__round__n2458 ), 
        .B(_f_permutation__round__n2457 ), .Z(_f_permutation__round__n2459 )
         );
  XOR2_X2 _f_permutation__round__U4388  ( .A(SYNOPSYS_UNCONNECTED_988), .B(
        _f_permutation__round__n2459 ), .Z(_f_permutation__round__c[1252] ) );
  XOR2_X2 _f_permutation__round__U4387  ( .A(SYNOPSYS_UNCONNECTED_668), .B(
        _f_permutation__round__n2459 ), .Z(_f_permutation__round__c[1188] ) );
  XOR2_X2 _f_permutation__round__U4386  ( .A(SYNOPSYS_UNCONNECTED_348), .B(
        _f_permutation__round__n2459 ), .Z(_f_permutation__round__c[1124] ) );
  XOR2_X2 _f_permutation__round__U4385  ( .A(_f_permutation__round_in[1060]), 
        .B(_f_permutation__round__n2459 ), .Z(_f_permutation__round__c[1060] )
         );
  XOR2_X2 _f_permutation__round__U4384  ( .A(_f_permutation__round_in[1380]), 
        .B(_f_permutation__round__n2459 ), .Z(_f_permutation__round__c[996] )
         );
  XOR2_X2 _f_permutation__round__U4383  ( .A(_f_permutation__round__n2461 ), 
        .B(_f_permutation__round__n2460 ), .Z(_f_permutation__round__n2462 )
         );
  XOR2_X2 _f_permutation__round__U4382  ( .A(SYNOPSYS_UNCONNECTED_989), .B(
        _f_permutation__round__n2462 ), .Z(_f_permutation__round__c[1251] ) );
  XOR2_X2 _f_permutation__round__U4381  ( .A(SYNOPSYS_UNCONNECTED_669), .B(
        _f_permutation__round__n2462 ), .Z(_f_permutation__round__c[1187] ) );
  XOR2_X2 _f_permutation__round__U4380  ( .A(SYNOPSYS_UNCONNECTED_349), .B(
        _f_permutation__round__n2462 ), .Z(_f_permutation__round__c[1123] ) );
  XOR2_X2 _f_permutation__round__U4379  ( .A(_f_permutation__round_in[1059]), 
        .B(_f_permutation__round__n2462 ), .Z(_f_permutation__round__c[1059] )
         );
  XOR2_X2 _f_permutation__round__U4378  ( .A(_f_permutation__round_in[1379]), 
        .B(_f_permutation__round__n2462 ), .Z(_f_permutation__round__c[995] )
         );
  XOR2_X2 _f_permutation__round__U4377  ( .A(_f_permutation__round__n2464 ), 
        .B(_f_permutation__round__n2463 ), .Z(_f_permutation__round__n2465 )
         );
  XOR2_X2 _f_permutation__round__U4376  ( .A(SYNOPSYS_UNCONNECTED_990), .B(
        _f_permutation__round__n2465 ), .Z(_f_permutation__round__c[1250] ) );
  XOR2_X2 _f_permutation__round__U4375  ( .A(SYNOPSYS_UNCONNECTED_670), .B(
        _f_permutation__round__n2465 ), .Z(_f_permutation__round__c[1186] ) );
  XOR2_X2 _f_permutation__round__U4374  ( .A(SYNOPSYS_UNCONNECTED_350), .B(
        _f_permutation__round__n2465 ), .Z(_f_permutation__round__c[1122] ) );
  XOR2_X2 _f_permutation__round__U4373  ( .A(_f_permutation__round_in[1058]), 
        .B(_f_permutation__round__n2465 ), .Z(_f_permutation__round__c[1058] )
         );
  XOR2_X2 _f_permutation__round__U4372  ( .A(_f_permutation__round_in[1378]), 
        .B(_f_permutation__round__n2465 ), .Z(_f_permutation__round__c[994] )
         );
  XOR2_X2 _f_permutation__round__U4371  ( .A(_f_permutation__round__n2467 ), 
        .B(_f_permutation__round__n2466 ), .Z(_f_permutation__round__n2468 )
         );
  XOR2_X2 _f_permutation__round__U4370  ( .A(SYNOPSYS_UNCONNECTED_991), .B(
        _f_permutation__round__n2468 ), .Z(_f_permutation__round__c[1249] ) );
  XOR2_X2 _f_permutation__round__U4369  ( .A(SYNOPSYS_UNCONNECTED_671), .B(
        _f_permutation__round__n2468 ), .Z(_f_permutation__round__c[1185] ) );
  XOR2_X2 _f_permutation__round__U4368  ( .A(SYNOPSYS_UNCONNECTED_351), .B(
        _f_permutation__round__n2468 ), .Z(_f_permutation__round__c[1121] ) );
  XOR2_X2 _f_permutation__round__U4367  ( .A(_f_permutation__round_in[1057]), 
        .B(_f_permutation__round__n2468 ), .Z(_f_permutation__round__c[1057] )
         );
  XOR2_X2 _f_permutation__round__U4366  ( .A(_f_permutation__round_in[1377]), 
        .B(_f_permutation__round__n2468 ), .Z(_f_permutation__round__c[993] )
         );
  XOR2_X2 _f_permutation__round__U4365  ( .A(_f_permutation__round__n2470 ), 
        .B(_f_permutation__round__n2469 ), .Z(_f_permutation__round__n2471 )
         );
  XOR2_X2 _f_permutation__round__U4364  ( .A(SYNOPSYS_UNCONNECTED_992), .B(
        _f_permutation__round__n2471 ), .Z(_f_permutation__round__c[1248] ) );
  XOR2_X2 _f_permutation__round__U4363  ( .A(SYNOPSYS_UNCONNECTED_672), .B(
        _f_permutation__round__n2471 ), .Z(_f_permutation__round__c[1184] ) );
  XOR2_X2 _f_permutation__round__U4362  ( .A(SYNOPSYS_UNCONNECTED_352), .B(
        _f_permutation__round__n2471 ), .Z(_f_permutation__round__c[1120] ) );
  XOR2_X2 _f_permutation__round__U4361  ( .A(_f_permutation__round_in[1056]), 
        .B(_f_permutation__round__n2471 ), .Z(_f_permutation__round__c[1056] )
         );
  XOR2_X2 _f_permutation__round__U4360  ( .A(_f_permutation__round_in[1376]), 
        .B(_f_permutation__round__n2471 ), .Z(_f_permutation__round__c[992] )
         );
  XOR2_X2 _f_permutation__round__U4359  ( .A(_f_permutation__round__n2473 ), 
        .B(_f_permutation__round__n2472 ), .Z(_f_permutation__round__n2474 )
         );
  XOR2_X2 _f_permutation__round__U4358  ( .A(SYNOPSYS_UNCONNECTED_993), .B(
        _f_permutation__round__n2474 ), .Z(_f_permutation__round__c[1247] ) );
  XOR2_X2 _f_permutation__round__U4357  ( .A(SYNOPSYS_UNCONNECTED_673), .B(
        _f_permutation__round__n2474 ), .Z(_f_permutation__round__c[1183] ) );
  XOR2_X2 _f_permutation__round__U4356  ( .A(SYNOPSYS_UNCONNECTED_353), .B(
        _f_permutation__round__n2474 ), .Z(_f_permutation__round__c[1119] ) );
  XOR2_X2 _f_permutation__round__U4355  ( .A(_f_permutation__round_in[1055]), 
        .B(_f_permutation__round__n2474 ), .Z(_f_permutation__round__c[1055] )
         );
  XOR2_X2 _f_permutation__round__U4354  ( .A(_f_permutation__round_in[1375]), 
        .B(_f_permutation__round__n2474 ), .Z(_f_permutation__round__c[991] )
         );
  XOR2_X2 _f_permutation__round__U4353  ( .A(_f_permutation__round__n2476 ), 
        .B(_f_permutation__round__n2475 ), .Z(_f_permutation__round__n2477 )
         );
  XOR2_X2 _f_permutation__round__U4352  ( .A(SYNOPSYS_UNCONNECTED_994), .B(
        _f_permutation__round__n2477 ), .Z(_f_permutation__round__c[1246] ) );
  XOR2_X2 _f_permutation__round__U4351  ( .A(SYNOPSYS_UNCONNECTED_674), .B(
        _f_permutation__round__n2477 ), .Z(_f_permutation__round__c[1182] ) );
  XOR2_X2 _f_permutation__round__U4350  ( .A(SYNOPSYS_UNCONNECTED_354), .B(
        _f_permutation__round__n2477 ), .Z(_f_permutation__round__c[1118] ) );
  XOR2_X2 _f_permutation__round__U4349  ( .A(_f_permutation__round_in[1054]), 
        .B(_f_permutation__round__n2477 ), .Z(_f_permutation__round__c[1054] )
         );
  XOR2_X2 _f_permutation__round__U4348  ( .A(_f_permutation__round_in[1374]), 
        .B(_f_permutation__round__n2477 ), .Z(_f_permutation__round__c[990] )
         );
  XOR2_X2 _f_permutation__round__U4347  ( .A(_f_permutation__round__n2479 ), 
        .B(_f_permutation__round__n2478 ), .Z(_f_permutation__round__n2480 )
         );
  XOR2_X2 _f_permutation__round__U4346  ( .A(SYNOPSYS_UNCONNECTED_995), .B(
        _f_permutation__round__n2480 ), .Z(_f_permutation__round__c[1245] ) );
  XOR2_X2 _f_permutation__round__U4345  ( .A(SYNOPSYS_UNCONNECTED_675), .B(
        _f_permutation__round__n2480 ), .Z(_f_permutation__round__c[1181] ) );
  XOR2_X2 _f_permutation__round__U4344  ( .A(SYNOPSYS_UNCONNECTED_355), .B(
        _f_permutation__round__n2480 ), .Z(_f_permutation__round__c[1117] ) );
  XOR2_X2 _f_permutation__round__U4343  ( .A(_f_permutation__round_in[1053]), 
        .B(_f_permutation__round__n2480 ), .Z(_f_permutation__round__c[1053] )
         );
  XOR2_X2 _f_permutation__round__U4342  ( .A(_f_permutation__round_in[1373]), 
        .B(_f_permutation__round__n2480 ), .Z(_f_permutation__round__c[989] )
         );
  XOR2_X2 _f_permutation__round__U4341  ( .A(_f_permutation__round__n2482 ), 
        .B(_f_permutation__round__n2481 ), .Z(_f_permutation__round__n2483 )
         );
  XOR2_X2 _f_permutation__round__U4340  ( .A(SYNOPSYS_UNCONNECTED_996), .B(
        _f_permutation__round__n2483 ), .Z(_f_permutation__round__c[1244] ) );
  XOR2_X2 _f_permutation__round__U4339  ( .A(SYNOPSYS_UNCONNECTED_676), .B(
        _f_permutation__round__n2483 ), .Z(_f_permutation__round__c[1180] ) );
  XOR2_X2 _f_permutation__round__U4338  ( .A(SYNOPSYS_UNCONNECTED_356), .B(
        _f_permutation__round__n2483 ), .Z(_f_permutation__round__c[1116] ) );
  XOR2_X2 _f_permutation__round__U4337  ( .A(_f_permutation__round_in[1052]), 
        .B(_f_permutation__round__n2483 ), .Z(_f_permutation__round__c[1052] )
         );
  XOR2_X2 _f_permutation__round__U4336  ( .A(_f_permutation__round_in[1372]), 
        .B(_f_permutation__round__n2483 ), .Z(_f_permutation__round__c[988] )
         );
  XOR2_X2 _f_permutation__round__U4335  ( .A(_f_permutation__round__n2485 ), 
        .B(_f_permutation__round__n2484 ), .Z(_f_permutation__round__n2486 )
         );
  XOR2_X2 _f_permutation__round__U4334  ( .A(SYNOPSYS_UNCONNECTED_997), .B(
        _f_permutation__round__n2486 ), .Z(_f_permutation__round__c[1243] ) );
  XOR2_X2 _f_permutation__round__U4333  ( .A(SYNOPSYS_UNCONNECTED_677), .B(
        _f_permutation__round__n2486 ), .Z(_f_permutation__round__c[1179] ) );
  XOR2_X2 _f_permutation__round__U4332  ( .A(SYNOPSYS_UNCONNECTED_357), .B(
        _f_permutation__round__n2486 ), .Z(_f_permutation__round__c[1115] ) );
  XOR2_X2 _f_permutation__round__U4331  ( .A(_f_permutation__round_in[1051]), 
        .B(_f_permutation__round__n2486 ), .Z(_f_permutation__round__c[1051] )
         );
  XOR2_X2 _f_permutation__round__U4330  ( .A(_f_permutation__round_in[1371]), 
        .B(_f_permutation__round__n2486 ), .Z(_f_permutation__round__c[987] )
         );
  XOR2_X2 _f_permutation__round__U4329  ( .A(_f_permutation__round__n2488 ), 
        .B(_f_permutation__round__n2487 ), .Z(_f_permutation__round__n2489 )
         );
  XOR2_X2 _f_permutation__round__U4328  ( .A(SYNOPSYS_UNCONNECTED_998), .B(
        _f_permutation__round__n2489 ), .Z(_f_permutation__round__c[1242] ) );
  XOR2_X2 _f_permutation__round__U4327  ( .A(SYNOPSYS_UNCONNECTED_678), .B(
        _f_permutation__round__n2489 ), .Z(_f_permutation__round__c[1178] ) );
  XOR2_X2 _f_permutation__round__U4326  ( .A(SYNOPSYS_UNCONNECTED_358), .B(
        _f_permutation__round__n2489 ), .Z(_f_permutation__round__c[1114] ) );
  XOR2_X2 _f_permutation__round__U4325  ( .A(_f_permutation__round_in[1050]), 
        .B(_f_permutation__round__n2489 ), .Z(_f_permutation__round__c[1050] )
         );
  XOR2_X2 _f_permutation__round__U4324  ( .A(_f_permutation__round_in[1370]), 
        .B(_f_permutation__round__n2489 ), .Z(_f_permutation__round__c[986] )
         );
  XOR2_X2 _f_permutation__round__U4323  ( .A(_f_permutation__round__n2491 ), 
        .B(_f_permutation__round__n2490 ), .Z(_f_permutation__round__n2492 )
         );
  XOR2_X2 _f_permutation__round__U4322  ( .A(SYNOPSYS_UNCONNECTED_999), .B(
        _f_permutation__round__n2492 ), .Z(_f_permutation__round__c[1241] ) );
  XOR2_X2 _f_permutation__round__U4321  ( .A(SYNOPSYS_UNCONNECTED_679), .B(
        _f_permutation__round__n2492 ), .Z(_f_permutation__round__c[1177] ) );
  XOR2_X2 _f_permutation__round__U4320  ( .A(SYNOPSYS_UNCONNECTED_359), .B(
        _f_permutation__round__n2492 ), .Z(_f_permutation__round__c[1113] ) );
  XOR2_X2 _f_permutation__round__U4319  ( .A(_f_permutation__round_in[1049]), 
        .B(_f_permutation__round__n2492 ), .Z(_f_permutation__round__c[1049] )
         );
  XOR2_X2 _f_permutation__round__U4318  ( .A(_f_permutation__round_in[1369]), 
        .B(_f_permutation__round__n2492 ), .Z(_f_permutation__round__c[985] )
         );
  XOR2_X2 _f_permutation__round__U4317  ( .A(_f_permutation__round__n2494 ), 
        .B(_f_permutation__round__n2493 ), .Z(_f_permutation__round__n2495 )
         );
  XOR2_X2 _f_permutation__round__U4316  ( .A(SYNOPSYS_UNCONNECTED_1000), .B(
        _f_permutation__round__n2495 ), .Z(_f_permutation__round__c[1240] ) );
  XOR2_X2 _f_permutation__round__U4315  ( .A(SYNOPSYS_UNCONNECTED_680), .B(
        _f_permutation__round__n2495 ), .Z(_f_permutation__round__c[1176] ) );
  XOR2_X2 _f_permutation__round__U4314  ( .A(SYNOPSYS_UNCONNECTED_360), .B(
        _f_permutation__round__n2495 ), .Z(_f_permutation__round__c[1112] ) );
  XOR2_X2 _f_permutation__round__U4313  ( .A(_f_permutation__round_in[1048]), 
        .B(_f_permutation__round__n2495 ), .Z(_f_permutation__round__c[1048] )
         );
  XOR2_X2 _f_permutation__round__U4312  ( .A(_f_permutation__round_in[1368]), 
        .B(_f_permutation__round__n2495 ), .Z(_f_permutation__round__c[984] )
         );
  XOR2_X2 _f_permutation__round__U4311  ( .A(_f_permutation__round__n2497 ), 
        .B(_f_permutation__round__n2496 ), .Z(_f_permutation__round__n2498 )
         );
  XOR2_X2 _f_permutation__round__U4310  ( .A(SYNOPSYS_UNCONNECTED_1001), .B(
        _f_permutation__round__n2498 ), .Z(_f_permutation__round__c[1239] ) );
  XOR2_X2 _f_permutation__round__U4309  ( .A(SYNOPSYS_UNCONNECTED_681), .B(
        _f_permutation__round__n2498 ), .Z(_f_permutation__round__c[1175] ) );
  XOR2_X2 _f_permutation__round__U4308  ( .A(SYNOPSYS_UNCONNECTED_361), .B(
        _f_permutation__round__n2498 ), .Z(_f_permutation__round__c[1111] ) );
  XOR2_X2 _f_permutation__round__U4307  ( .A(_f_permutation__round_in[1047]), 
        .B(_f_permutation__round__n2498 ), .Z(_f_permutation__round__c[1047] )
         );
  XOR2_X2 _f_permutation__round__U4306  ( .A(_f_permutation__round_in[1367]), 
        .B(_f_permutation__round__n2498 ), .Z(_f_permutation__round__c[983] )
         );
  XOR2_X2 _f_permutation__round__U4305  ( .A(_f_permutation__round__n2500 ), 
        .B(_f_permutation__round__n2499 ), .Z(_f_permutation__round__n2501 )
         );
  XOR2_X2 _f_permutation__round__U4304  ( .A(SYNOPSYS_UNCONNECTED_1002), .B(
        _f_permutation__round__n2501 ), .Z(_f_permutation__round__c[1238] ) );
  XOR2_X2 _f_permutation__round__U4303  ( .A(SYNOPSYS_UNCONNECTED_682), .B(
        _f_permutation__round__n2501 ), .Z(_f_permutation__round__c[1174] ) );
  XOR2_X2 _f_permutation__round__U4302  ( .A(SYNOPSYS_UNCONNECTED_362), .B(
        _f_permutation__round__n2501 ), .Z(_f_permutation__round__c[1110] ) );
  XOR2_X2 _f_permutation__round__U4301  ( .A(_f_permutation__round_in[1046]), 
        .B(_f_permutation__round__n2501 ), .Z(_f_permutation__round__c[1046] )
         );
  XOR2_X2 _f_permutation__round__U4300  ( .A(_f_permutation__round_in[1366]), 
        .B(_f_permutation__round__n2501 ), .Z(_f_permutation__round__c[982] )
         );
  XOR2_X2 _f_permutation__round__U4299  ( .A(_f_permutation__round__n2503 ), 
        .B(_f_permutation__round__n2502 ), .Z(_f_permutation__round__n2504 )
         );
  XOR2_X2 _f_permutation__round__U4298  ( .A(SYNOPSYS_UNCONNECTED_1003), .B(
        _f_permutation__round__n2504 ), .Z(_f_permutation__round__c[1237] ) );
  XOR2_X2 _f_permutation__round__U4297  ( .A(SYNOPSYS_UNCONNECTED_683), .B(
        _f_permutation__round__n2504 ), .Z(_f_permutation__round__c[1173] ) );
  XOR2_X2 _f_permutation__round__U4296  ( .A(SYNOPSYS_UNCONNECTED_363), .B(
        _f_permutation__round__n2504 ), .Z(_f_permutation__round__c[1109] ) );
  XOR2_X2 _f_permutation__round__U4295  ( .A(_f_permutation__round_in[1045]), 
        .B(_f_permutation__round__n2504 ), .Z(_f_permutation__round__c[1045] )
         );
  XOR2_X2 _f_permutation__round__U4294  ( .A(_f_permutation__round_in[1365]), 
        .B(_f_permutation__round__n2504 ), .Z(_f_permutation__round__c[981] )
         );
  XOR2_X2 _f_permutation__round__U4293  ( .A(_f_permutation__round__n2506 ), 
        .B(_f_permutation__round__n2505 ), .Z(_f_permutation__round__n2507 )
         );
  XOR2_X2 _f_permutation__round__U4292  ( .A(SYNOPSYS_UNCONNECTED_1004), .B(
        _f_permutation__round__n2507 ), .Z(_f_permutation__round__c[1236] ) );
  XOR2_X2 _f_permutation__round__U4291  ( .A(SYNOPSYS_UNCONNECTED_684), .B(
        _f_permutation__round__n2507 ), .Z(_f_permutation__round__c[1172] ) );
  XOR2_X2 _f_permutation__round__U4290  ( .A(SYNOPSYS_UNCONNECTED_364), .B(
        _f_permutation__round__n2507 ), .Z(_f_permutation__round__c[1108] ) );
  XOR2_X2 _f_permutation__round__U4289  ( .A(_f_permutation__round_in[1044]), 
        .B(_f_permutation__round__n2507 ), .Z(_f_permutation__round__c[1044] )
         );
  XOR2_X2 _f_permutation__round__U4288  ( .A(_f_permutation__round_in[1364]), 
        .B(_f_permutation__round__n2507 ), .Z(_f_permutation__round__c[980] )
         );
  XOR2_X2 _f_permutation__round__U4287  ( .A(_f_permutation__round__n2509 ), 
        .B(_f_permutation__round__n2508 ), .Z(_f_permutation__round__n2510 )
         );
  XOR2_X2 _f_permutation__round__U4286  ( .A(SYNOPSYS_UNCONNECTED_1005), .B(
        _f_permutation__round__n2510 ), .Z(_f_permutation__round__c[1235] ) );
  XOR2_X2 _f_permutation__round__U4285  ( .A(SYNOPSYS_UNCONNECTED_685), .B(
        _f_permutation__round__n2510 ), .Z(_f_permutation__round__c[1171] ) );
  XOR2_X2 _f_permutation__round__U4284  ( .A(SYNOPSYS_UNCONNECTED_365), .B(
        _f_permutation__round__n2510 ), .Z(_f_permutation__round__c[1107] ) );
  XOR2_X2 _f_permutation__round__U4283  ( .A(_f_permutation__round_in[1043]), 
        .B(_f_permutation__round__n2510 ), .Z(_f_permutation__round__c[1043] )
         );
  XOR2_X2 _f_permutation__round__U4282  ( .A(_f_permutation__round_in[1363]), 
        .B(_f_permutation__round__n2510 ), .Z(_f_permutation__round__c[979] )
         );
  XOR2_X2 _f_permutation__round__U4281  ( .A(_f_permutation__round__n2512 ), 
        .B(_f_permutation__round__n2511 ), .Z(_f_permutation__round__n2513 )
         );
  XOR2_X2 _f_permutation__round__U4280  ( .A(SYNOPSYS_UNCONNECTED_1006), .B(
        _f_permutation__round__n2513 ), .Z(_f_permutation__round__c[1234] ) );
  XOR2_X2 _f_permutation__round__U4279  ( .A(SYNOPSYS_UNCONNECTED_686), .B(
        _f_permutation__round__n2513 ), .Z(_f_permutation__round__c[1170] ) );
  XOR2_X2 _f_permutation__round__U4278  ( .A(SYNOPSYS_UNCONNECTED_366), .B(
        _f_permutation__round__n2513 ), .Z(_f_permutation__round__c[1106] ) );
  XOR2_X2 _f_permutation__round__U4277  ( .A(_f_permutation__round_in[1042]), 
        .B(_f_permutation__round__n2513 ), .Z(_f_permutation__round__c[1042] )
         );
  XOR2_X2 _f_permutation__round__U4276  ( .A(_f_permutation__round_in[1362]), 
        .B(_f_permutation__round__n2513 ), .Z(_f_permutation__round__c[978] )
         );
  XOR2_X2 _f_permutation__round__U4275  ( .A(_f_permutation__round__n2515 ), 
        .B(_f_permutation__round__n2514 ), .Z(_f_permutation__round__n2516 )
         );
  XOR2_X2 _f_permutation__round__U4274  ( .A(SYNOPSYS_UNCONNECTED_1007), .B(
        _f_permutation__round__n2516 ), .Z(_f_permutation__round__c[1233] ) );
  XOR2_X2 _f_permutation__round__U4273  ( .A(SYNOPSYS_UNCONNECTED_687), .B(
        _f_permutation__round__n2516 ), .Z(_f_permutation__round__c[1169] ) );
  XOR2_X2 _f_permutation__round__U4272  ( .A(SYNOPSYS_UNCONNECTED_367), .B(
        _f_permutation__round__n2516 ), .Z(_f_permutation__round__c[1105] ) );
  XOR2_X2 _f_permutation__round__U4271  ( .A(_f_permutation__round_in[1041]), 
        .B(_f_permutation__round__n2516 ), .Z(_f_permutation__round__c[1041] )
         );
  XOR2_X2 _f_permutation__round__U4270  ( .A(_f_permutation__round_in[1361]), 
        .B(_f_permutation__round__n2516 ), .Z(_f_permutation__round__c[977] )
         );
  XOR2_X2 _f_permutation__round__U4269  ( .A(_f_permutation__round__n2518 ), 
        .B(_f_permutation__round__n2517 ), .Z(_f_permutation__round__n2519 )
         );
  XOR2_X2 _f_permutation__round__U4268  ( .A(SYNOPSYS_UNCONNECTED_1008), .B(
        _f_permutation__round__n2519 ), .Z(_f_permutation__round__c[1232] ) );
  XOR2_X2 _f_permutation__round__U4267  ( .A(SYNOPSYS_UNCONNECTED_688), .B(
        _f_permutation__round__n2519 ), .Z(_f_permutation__round__c[1168] ) );
  XOR2_X2 _f_permutation__round__U4266  ( .A(SYNOPSYS_UNCONNECTED_368), .B(
        _f_permutation__round__n2519 ), .Z(_f_permutation__round__c[1104] ) );
  XOR2_X2 _f_permutation__round__U4265  ( .A(_f_permutation__round_in[1040]), 
        .B(_f_permutation__round__n2519 ), .Z(_f_permutation__round__c[1040] )
         );
  XOR2_X2 _f_permutation__round__U4264  ( .A(_f_permutation__round_in[1360]), 
        .B(_f_permutation__round__n2519 ), .Z(_f_permutation__round__c[976] )
         );
  XOR2_X2 _f_permutation__round__U4263  ( .A(_f_permutation__round__n2521 ), 
        .B(_f_permutation__round__n2520 ), .Z(_f_permutation__round__n2522 )
         );
  XOR2_X2 _f_permutation__round__U4262  ( .A(SYNOPSYS_UNCONNECTED_1009), .B(
        _f_permutation__round__n2522 ), .Z(_f_permutation__round__c[1231] ) );
  XOR2_X2 _f_permutation__round__U4261  ( .A(SYNOPSYS_UNCONNECTED_689), .B(
        _f_permutation__round__n2522 ), .Z(_f_permutation__round__c[1167] ) );
  XOR2_X2 _f_permutation__round__U4260  ( .A(SYNOPSYS_UNCONNECTED_369), .B(
        _f_permutation__round__n2522 ), .Z(_f_permutation__round__c[1103] ) );
  XOR2_X2 _f_permutation__round__U4259  ( .A(_f_permutation__round_in[1039]), 
        .B(_f_permutation__round__n2522 ), .Z(_f_permutation__round__c[1039] )
         );
  XOR2_X2 _f_permutation__round__U4258  ( .A(_f_permutation__round_in[1359]), 
        .B(_f_permutation__round__n2522 ), .Z(_f_permutation__round__c[975] )
         );
  XOR2_X2 _f_permutation__round__U4257  ( .A(_f_permutation__round__n2524 ), 
        .B(_f_permutation__round__n2523 ), .Z(_f_permutation__round__n2525 )
         );
  XOR2_X2 _f_permutation__round__U4256  ( .A(SYNOPSYS_UNCONNECTED_1010), .B(
        _f_permutation__round__n2525 ), .Z(_f_permutation__round__c[1230] ) );
  XOR2_X2 _f_permutation__round__U4255  ( .A(SYNOPSYS_UNCONNECTED_690), .B(
        _f_permutation__round__n2525 ), .Z(_f_permutation__round__c[1166] ) );
  XOR2_X2 _f_permutation__round__U4254  ( .A(SYNOPSYS_UNCONNECTED_370), .B(
        _f_permutation__round__n2525 ), .Z(_f_permutation__round__c[1102] ) );
  XOR2_X2 _f_permutation__round__U4253  ( .A(_f_permutation__round_in[1038]), 
        .B(_f_permutation__round__n2525 ), .Z(_f_permutation__round__c[1038] )
         );
  XOR2_X2 _f_permutation__round__U4252  ( .A(_f_permutation__round_in[1358]), 
        .B(_f_permutation__round__n2525 ), .Z(_f_permutation__round__c[974] )
         );
  XOR2_X2 _f_permutation__round__U4251  ( .A(_f_permutation__round__n2527 ), 
        .B(_f_permutation__round__n2526 ), .Z(_f_permutation__round__n2528 )
         );
  XOR2_X2 _f_permutation__round__U4250  ( .A(SYNOPSYS_UNCONNECTED_1011), .B(
        _f_permutation__round__n2528 ), .Z(_f_permutation__round__c[1229] ) );
  XOR2_X2 _f_permutation__round__U4249  ( .A(SYNOPSYS_UNCONNECTED_691), .B(
        _f_permutation__round__n2528 ), .Z(_f_permutation__round__c[1165] ) );
  XOR2_X2 _f_permutation__round__U4248  ( .A(SYNOPSYS_UNCONNECTED_371), .B(
        _f_permutation__round__n2528 ), .Z(_f_permutation__round__c[1101] ) );
  XOR2_X2 _f_permutation__round__U4247  ( .A(_f_permutation__round_in[1037]), 
        .B(_f_permutation__round__n2528 ), .Z(_f_permutation__round__c[1037] )
         );
  XOR2_X2 _f_permutation__round__U4246  ( .A(_f_permutation__round_in[1357]), 
        .B(_f_permutation__round__n2528 ), .Z(_f_permutation__round__c[973] )
         );
  XOR2_X2 _f_permutation__round__U4245  ( .A(_f_permutation__round__n2530 ), 
        .B(_f_permutation__round__n2529 ), .Z(_f_permutation__round__n2531 )
         );
  XOR2_X2 _f_permutation__round__U4244  ( .A(SYNOPSYS_UNCONNECTED_1012), .B(
        _f_permutation__round__n2531 ), .Z(_f_permutation__round__c[1228] ) );
  XOR2_X2 _f_permutation__round__U4243  ( .A(SYNOPSYS_UNCONNECTED_692), .B(
        _f_permutation__round__n2531 ), .Z(_f_permutation__round__c[1164] ) );
  XOR2_X2 _f_permutation__round__U4242  ( .A(SYNOPSYS_UNCONNECTED_372), .B(
        _f_permutation__round__n2531 ), .Z(_f_permutation__round__c[1100] ) );
  XOR2_X2 _f_permutation__round__U4241  ( .A(_f_permutation__round_in[1036]), 
        .B(_f_permutation__round__n2531 ), .Z(_f_permutation__round__c[1036] )
         );
  XOR2_X2 _f_permutation__round__U4240  ( .A(_f_permutation__round_in[1356]), 
        .B(_f_permutation__round__n2531 ), .Z(_f_permutation__round__c[972] )
         );
  XOR2_X2 _f_permutation__round__U4239  ( .A(_f_permutation__round__n2533 ), 
        .B(_f_permutation__round__n2532 ), .Z(_f_permutation__round__n2534 )
         );
  XOR2_X2 _f_permutation__round__U4238  ( .A(SYNOPSYS_UNCONNECTED_1013), .B(
        _f_permutation__round__n2534 ), .Z(_f_permutation__round__c[1227] ) );
  XOR2_X2 _f_permutation__round__U4237  ( .A(SYNOPSYS_UNCONNECTED_693), .B(
        _f_permutation__round__n2534 ), .Z(_f_permutation__round__c[1163] ) );
  XOR2_X2 _f_permutation__round__U4236  ( .A(SYNOPSYS_UNCONNECTED_373), .B(
        _f_permutation__round__n2534 ), .Z(_f_permutation__round__c[1099] ) );
  XOR2_X2 _f_permutation__round__U4235  ( .A(_f_permutation__round_in[1035]), 
        .B(_f_permutation__round__n2534 ), .Z(_f_permutation__round__c[1035] )
         );
  XOR2_X2 _f_permutation__round__U4234  ( .A(_f_permutation__round_in[1355]), 
        .B(_f_permutation__round__n2534 ), .Z(_f_permutation__round__c[971] )
         );
  XOR2_X2 _f_permutation__round__U4233  ( .A(_f_permutation__round__n2536 ), 
        .B(_f_permutation__round__n2535 ), .Z(_f_permutation__round__n2537 )
         );
  XOR2_X2 _f_permutation__round__U4232  ( .A(SYNOPSYS_UNCONNECTED_1014), .B(
        _f_permutation__round__n2537 ), .Z(_f_permutation__round__c[1226] ) );
  XOR2_X2 _f_permutation__round__U4231  ( .A(SYNOPSYS_UNCONNECTED_694), .B(
        _f_permutation__round__n2537 ), .Z(_f_permutation__round__c[1162] ) );
  XOR2_X2 _f_permutation__round__U4230  ( .A(SYNOPSYS_UNCONNECTED_374), .B(
        _f_permutation__round__n2537 ), .Z(_f_permutation__round__c[1098] ) );
  XOR2_X2 _f_permutation__round__U4229  ( .A(_f_permutation__round_in[1034]), 
        .B(_f_permutation__round__n2537 ), .Z(_f_permutation__round__c[1034] )
         );
  XOR2_X2 _f_permutation__round__U4228  ( .A(_f_permutation__round_in[1354]), 
        .B(_f_permutation__round__n2537 ), .Z(_f_permutation__round__c[970] )
         );
  XOR2_X2 _f_permutation__round__U4227  ( .A(_f_permutation__round__n2539 ), 
        .B(_f_permutation__round__n2538 ), .Z(_f_permutation__round__n2540 )
         );
  XOR2_X2 _f_permutation__round__U4226  ( .A(SYNOPSYS_UNCONNECTED_1015), .B(
        _f_permutation__round__n2540 ), .Z(_f_permutation__round__c[1225] ) );
  XOR2_X2 _f_permutation__round__U4225  ( .A(SYNOPSYS_UNCONNECTED_695), .B(
        _f_permutation__round__n2540 ), .Z(_f_permutation__round__c[1161] ) );
  XOR2_X2 _f_permutation__round__U4224  ( .A(SYNOPSYS_UNCONNECTED_375), .B(
        _f_permutation__round__n2540 ), .Z(_f_permutation__round__c[1097] ) );
  XOR2_X2 _f_permutation__round__U4223  ( .A(_f_permutation__round_in[1033]), 
        .B(_f_permutation__round__n2540 ), .Z(_f_permutation__round__c[1033] )
         );
  XOR2_X2 _f_permutation__round__U4222  ( .A(_f_permutation__round_in[1353]), 
        .B(_f_permutation__round__n2540 ), .Z(_f_permutation__round__c[969] )
         );
  XOR2_X2 _f_permutation__round__U4221  ( .A(_f_permutation__round__n2542 ), 
        .B(_f_permutation__round__n2541 ), .Z(_f_permutation__round__n2543 )
         );
  XOR2_X2 _f_permutation__round__U4220  ( .A(SYNOPSYS_UNCONNECTED_1016), .B(
        _f_permutation__round__n2543 ), .Z(_f_permutation__round__c[1224] ) );
  XOR2_X2 _f_permutation__round__U4219  ( .A(SYNOPSYS_UNCONNECTED_696), .B(
        _f_permutation__round__n2543 ), .Z(_f_permutation__round__c[1160] ) );
  XOR2_X2 _f_permutation__round__U4218  ( .A(SYNOPSYS_UNCONNECTED_376), .B(
        _f_permutation__round__n2543 ), .Z(_f_permutation__round__c[1096] ) );
  XOR2_X2 _f_permutation__round__U4217  ( .A(_f_permutation__round_in[1032]), 
        .B(_f_permutation__round__n2543 ), .Z(_f_permutation__round__c[1032] )
         );
  XOR2_X2 _f_permutation__round__U4216  ( .A(_f_permutation__round_in[1352]), 
        .B(_f_permutation__round__n2543 ), .Z(_f_permutation__round__c[968] )
         );
  XOR2_X2 _f_permutation__round__U4215  ( .A(_f_permutation__round__n2545 ), 
        .B(_f_permutation__round__n2544 ), .Z(_f_permutation__round__n2546 )
         );
  XOR2_X2 _f_permutation__round__U4214  ( .A(SYNOPSYS_UNCONNECTED_1017), .B(
        _f_permutation__round__n2546 ), .Z(_f_permutation__round__c[1223] ) );
  XOR2_X2 _f_permutation__round__U4213  ( .A(SYNOPSYS_UNCONNECTED_697), .B(
        _f_permutation__round__n2546 ), .Z(_f_permutation__round__c[1159] ) );
  XOR2_X2 _f_permutation__round__U4212  ( .A(SYNOPSYS_UNCONNECTED_377), .B(
        _f_permutation__round__n2546 ), .Z(_f_permutation__round__c[1095] ) );
  XOR2_X2 _f_permutation__round__U4211  ( .A(_f_permutation__round_in[1031]), 
        .B(_f_permutation__round__n2546 ), .Z(_f_permutation__round__c[1031] )
         );
  XOR2_X2 _f_permutation__round__U4210  ( .A(_f_permutation__round_in[1351]), 
        .B(_f_permutation__round__n2546 ), .Z(_f_permutation__round__c[967] )
         );
  XOR2_X2 _f_permutation__round__U4209  ( .A(_f_permutation__round__n2548 ), 
        .B(_f_permutation__round__n2547 ), .Z(_f_permutation__round__n2549 )
         );
  XOR2_X2 _f_permutation__round__U4208  ( .A(SYNOPSYS_UNCONNECTED_1018), .B(
        _f_permutation__round__n2549 ), .Z(_f_permutation__round__c[1222] ) );
  XOR2_X2 _f_permutation__round__U4207  ( .A(SYNOPSYS_UNCONNECTED_698), .B(
        _f_permutation__round__n2549 ), .Z(_f_permutation__round__c[1158] ) );
  XOR2_X2 _f_permutation__round__U4206  ( .A(SYNOPSYS_UNCONNECTED_378), .B(
        _f_permutation__round__n2549 ), .Z(_f_permutation__round__c[1094] ) );
  XOR2_X2 _f_permutation__round__U4205  ( .A(_f_permutation__round_in[1030]), 
        .B(_f_permutation__round__n2549 ), .Z(_f_permutation__round__c[1030] )
         );
  XOR2_X2 _f_permutation__round__U4204  ( .A(_f_permutation__round_in[1350]), 
        .B(_f_permutation__round__n2549 ), .Z(_f_permutation__round__c[966] )
         );
  XOR2_X2 _f_permutation__round__U4203  ( .A(_f_permutation__round__n2551 ), 
        .B(_f_permutation__round__n2550 ), .Z(_f_permutation__round__n2552 )
         );
  XOR2_X2 _f_permutation__round__U4202  ( .A(SYNOPSYS_UNCONNECTED_1019), .B(
        _f_permutation__round__n2552 ), .Z(_f_permutation__round__c[1221] ) );
  XOR2_X2 _f_permutation__round__U4201  ( .A(SYNOPSYS_UNCONNECTED_699), .B(
        _f_permutation__round__n2552 ), .Z(_f_permutation__round__c[1157] ) );
  XOR2_X2 _f_permutation__round__U4200  ( .A(SYNOPSYS_UNCONNECTED_379), .B(
        _f_permutation__round__n2552 ), .Z(_f_permutation__round__c[1093] ) );
  XOR2_X2 _f_permutation__round__U4199  ( .A(_f_permutation__round_in[1029]), 
        .B(_f_permutation__round__n2552 ), .Z(_f_permutation__round__c[1029] )
         );
  XOR2_X2 _f_permutation__round__U4198  ( .A(_f_permutation__round_in[1349]), 
        .B(_f_permutation__round__n2552 ), .Z(_f_permutation__round__c[965] )
         );
  XOR2_X2 _f_permutation__round__U4197  ( .A(_f_permutation__round__n2554 ), 
        .B(_f_permutation__round__n2553 ), .Z(_f_permutation__round__n2555 )
         );
  XOR2_X2 _f_permutation__round__U4196  ( .A(SYNOPSYS_UNCONNECTED_1020), .B(
        _f_permutation__round__n2555 ), .Z(_f_permutation__round__c[1220] ) );
  XOR2_X2 _f_permutation__round__U4195  ( .A(SYNOPSYS_UNCONNECTED_700), .B(
        _f_permutation__round__n2555 ), .Z(_f_permutation__round__c[1156] ) );
  XOR2_X2 _f_permutation__round__U4194  ( .A(SYNOPSYS_UNCONNECTED_380), .B(
        _f_permutation__round__n2555 ), .Z(_f_permutation__round__c[1092] ) );
  XOR2_X2 _f_permutation__round__U4193  ( .A(_f_permutation__round_in[1028]), 
        .B(_f_permutation__round__n2555 ), .Z(_f_permutation__round__c[1028] )
         );
  XOR2_X2 _f_permutation__round__U4192  ( .A(_f_permutation__round_in[1348]), 
        .B(_f_permutation__round__n2555 ), .Z(_f_permutation__round__c[964] )
         );
  XOR2_X2 _f_permutation__round__U4191  ( .A(_f_permutation__round__n2557 ), 
        .B(_f_permutation__round__n2556 ), .Z(_f_permutation__round__n2558 )
         );
  XOR2_X2 _f_permutation__round__U4190  ( .A(SYNOPSYS_UNCONNECTED_1021), .B(
        _f_permutation__round__n2558 ), .Z(_f_permutation__round__c[1219] ) );
  XOR2_X2 _f_permutation__round__U4189  ( .A(SYNOPSYS_UNCONNECTED_701), .B(
        _f_permutation__round__n2558 ), .Z(_f_permutation__round__c[1155] ) );
  XOR2_X2 _f_permutation__round__U4188  ( .A(SYNOPSYS_UNCONNECTED_381), .B(
        _f_permutation__round__n2558 ), .Z(_f_permutation__round__c[1091] ) );
  XOR2_X2 _f_permutation__round__U4187  ( .A(_f_permutation__round_in[1027]), 
        .B(_f_permutation__round__n2558 ), .Z(_f_permutation__round__c[1027] )
         );
  XOR2_X2 _f_permutation__round__U4186  ( .A(_f_permutation__round_in[1347]), 
        .B(_f_permutation__round__n2558 ), .Z(_f_permutation__round__c[963] )
         );
  XOR2_X2 _f_permutation__round__U4185  ( .A(_f_permutation__round__n2560 ), 
        .B(_f_permutation__round__n2559 ), .Z(_f_permutation__round__n25610 )
         );
  XOR2_X2 _f_permutation__round__U4184  ( .A(SYNOPSYS_UNCONNECTED_1022), .B(
        _f_permutation__round__n25610 ), .Z(_f_permutation__round__c[1218] )
         );
  XOR2_X2 _f_permutation__round__U4183  ( .A(SYNOPSYS_UNCONNECTED_702), .B(
        _f_permutation__round__n25610 ), .Z(_f_permutation__round__c[1154] )
         );
  XOR2_X2 _f_permutation__round__U4182  ( .A(SYNOPSYS_UNCONNECTED_382), .B(
        _f_permutation__round__n25610 ), .Z(_f_permutation__round__c[1090] )
         );
  XOR2_X2 _f_permutation__round__U4181  ( .A(_f_permutation__round_in[1026]), 
        .B(_f_permutation__round__n25610 ), .Z(_f_permutation__round__c[1026] ) );
  XOR2_X2 _f_permutation__round__U4180  ( .A(_f_permutation__round_in[1346]), 
        .B(_f_permutation__round__n25610 ), .Z(_f_permutation__round__c[962] )
         );
  XOR2_X2 _f_permutation__round__U4179  ( .A(_f_permutation__round__n25630 ), 
        .B(_f_permutation__round__n2562 ), .Z(_f_permutation__round__n2564 )
         );
  XOR2_X2 _f_permutation__round__U4178  ( .A(SYNOPSYS_UNCONNECTED_1023), .B(
        _f_permutation__round__n2564 ), .Z(_f_permutation__round__c[1217] ) );
  XOR2_X2 _f_permutation__round__U4177  ( .A(SYNOPSYS_UNCONNECTED_703), .B(
        _f_permutation__round__n2564 ), .Z(_f_permutation__round__c[1153] ) );
  XOR2_X2 _f_permutation__round__U4176  ( .A(SYNOPSYS_UNCONNECTED_383), .B(
        _f_permutation__round__n2564 ), .Z(_f_permutation__round__c[1089] ) );
  XOR2_X2 _f_permutation__round__U4175  ( .A(_f_permutation__round_in[1025]), 
        .B(_f_permutation__round__n2564 ), .Z(_f_permutation__round__c[1025] )
         );
  XOR2_X2 _f_permutation__round__U4174  ( .A(_f_permutation__round_in[1345]), 
        .B(_f_permutation__round__n2564 ), .Z(_f_permutation__round__c[961] )
         );
  XOR2_X2 _f_permutation__round__U4173  ( .A(_f_permutation__round__n2566 ), 
        .B(_f_permutation__round__n25650 ), .Z(_f_permutation__round__n25670 )
         );
  XOR2_X2 _f_permutation__round__U4172  ( .A(SYNOPSYS_UNCONNECTED_1024), .B(
        _f_permutation__round__n25670 ), .Z(_f_permutation__round__c[1216] )
         );
  XOR2_X2 _f_permutation__round__U4171  ( .A(SYNOPSYS_UNCONNECTED_704), .B(
        _f_permutation__round__n25670 ), .Z(_f_permutation__round__c[1152] )
         );
  XOR2_X2 _f_permutation__round__U4170  ( .A(SYNOPSYS_UNCONNECTED_384), .B(
        _f_permutation__round__n25670 ), .Z(_f_permutation__round__c[1088] )
         );
  XOR2_X2 _f_permutation__round__U4169  ( .A(_f_permutation__round_in[1024]), 
        .B(_f_permutation__round__n25670 ), .Z(_f_permutation__round__c[1024] ) );
  XOR2_X2 _f_permutation__round__U4168  ( .A(_f_permutation__round_in[1344]), 
        .B(_f_permutation__round__n25670 ), .Z(_f_permutation__round__c[960] )
         );
  XOR2_X2 _f_permutation__round__U4167  ( .A(_f_permutation__round__N5759 ), 
        .B(_f_permutation__round__c[638] ), .Z(_f_permutation__round_out[0])
         );
  XOR2_X2 _f_permutation__round__U4166  ( .A(_f_permutation__round__N5757 ), 
        .B(_f_permutation__round__c[639] ), .Z(_f_permutation__round_out[1])
         );
  XOR2_X2 _f_permutation__round__U4165  ( .A(_f_permutation__round__N5755 ), 
        .B(_f_permutation__round__c[576] ), .Z(_f_permutation__round_out[2])
         );
  XOR2_X2 _f_permutation__round__U4164  ( .A(_f_permutation__round__N5753 ), 
        .B(_f_permutation__round__c[577] ), .Z(_f_permutation__round_out[3])
         );
  XOR2_X2 _f_permutation__round__U4163  ( .A(_f_permutation__round__N5751 ), 
        .B(_f_permutation__round__c[578] ), .Z(_f_permutation__round_out[4])
         );
  XOR2_X2 _f_permutation__round__U4162  ( .A(_f_permutation__round__N5749 ), 
        .B(_f_permutation__round__c[579] ), .Z(_f_permutation__round_out[5])
         );
  XOR2_X2 _f_permutation__round__U4161  ( .A(_f_permutation__round__N5747 ), 
        .B(_f_permutation__round__c[580] ), .Z(_f_permutation__round_out[6])
         );
  XOR2_X2 _f_permutation__round__U4160  ( .A(_f_permutation__round__N5745 ), 
        .B(_f_permutation__round__c[581] ), .Z(_f_permutation__round_out[7])
         );
  XOR2_X2 _f_permutation__round__U4159  ( .A(_f_permutation__round__N5743 ), 
        .B(_f_permutation__round__c[582] ), .Z(_f_permutation__round_out[8])
         );
  XOR2_X2 _f_permutation__round__U4158  ( .A(_f_permutation__round__N5741 ), 
        .B(_f_permutation__round__c[583] ), .Z(_f_permutation__round_out[9])
         );
  XOR2_X2 _f_permutation__round__U4157  ( .A(_f_permutation__round__N5739 ), 
        .B(_f_permutation__round__c[584] ), .Z(_f_permutation__round_out[10])
         );
  XOR2_X2 _f_permutation__round__U4156  ( .A(_f_permutation__round__N5737 ), 
        .B(_f_permutation__round__c[585] ), .Z(_f_permutation__round_out[11])
         );
  XOR2_X2 _f_permutation__round__U4155  ( .A(_f_permutation__round__N5735 ), 
        .B(_f_permutation__round__c[586] ), .Z(_f_permutation__round_out[12])
         );
  XOR2_X2 _f_permutation__round__U4154  ( .A(_f_permutation__round__N5733 ), 
        .B(_f_permutation__round__c[587] ), .Z(_f_permutation__round_out[13])
         );
  XOR2_X2 _f_permutation__round__U4153  ( .A(_f_permutation__round__N5731 ), 
        .B(_f_permutation__round__c[588] ), .Z(_f_permutation__round_out[14])
         );
  XOR2_X2 _f_permutation__round__U4152  ( .A(_f_permutation__round__N5729 ), 
        .B(_f_permutation__round__c[589] ), .Z(_f_permutation__round_out[15])
         );
  XOR2_X2 _f_permutation__round__U4151  ( .A(_f_permutation__round__N5727 ), 
        .B(_f_permutation__round__c[590] ), .Z(_f_permutation__round_out[16])
         );
  XOR2_X2 _f_permutation__round__U4150  ( .A(_f_permutation__round__N5725 ), 
        .B(_f_permutation__round__c[591] ), .Z(_f_permutation__round_out[17])
         );
  XOR2_X2 _f_permutation__round__U4149  ( .A(_f_permutation__round__N5723 ), 
        .B(_f_permutation__round__c[592] ), .Z(_f_permutation__round_out[18])
         );
  XOR2_X2 _f_permutation__round__U4148  ( .A(_f_permutation__round__N5721 ), 
        .B(_f_permutation__round__c[593] ), .Z(_f_permutation__round_out[19])
         );
  XOR2_X2 _f_permutation__round__U4147  ( .A(_f_permutation__round__N5719 ), 
        .B(_f_permutation__round__c[594] ), .Z(_f_permutation__round_out[20])
         );
  XOR2_X2 _f_permutation__round__U4146  ( .A(_f_permutation__round__N5717 ), 
        .B(_f_permutation__round__c[595] ), .Z(_f_permutation__round_out[21])
         );
  XOR2_X2 _f_permutation__round__U4145  ( .A(_f_permutation__round__N5715 ), 
        .B(_f_permutation__round__c[596] ), .Z(_f_permutation__round_out[22])
         );
  XOR2_X2 _f_permutation__round__U4144  ( .A(_f_permutation__round__N5713 ), 
        .B(_f_permutation__round__c[597] ), .Z(_f_permutation__round_out[23])
         );
  XOR2_X2 _f_permutation__round__U4143  ( .A(_f_permutation__round__N5711 ), 
        .B(_f_permutation__round__c[598] ), .Z(_f_permutation__round_out[24])
         );
  XOR2_X2 _f_permutation__round__U4142  ( .A(_f_permutation__round__N5709 ), 
        .B(_f_permutation__round__c[599] ), .Z(_f_permutation__round_out[25])
         );
  XOR2_X2 _f_permutation__round__U4141  ( .A(_f_permutation__round__N5707 ), 
        .B(_f_permutation__round__c[600] ), .Z(_f_permutation__round_out[26])
         );
  XOR2_X2 _f_permutation__round__U4140  ( .A(_f_permutation__round__N5705 ), 
        .B(_f_permutation__round__c[601] ), .Z(_f_permutation__round_out[27])
         );
  XOR2_X2 _f_permutation__round__U4139  ( .A(_f_permutation__round__N5703 ), 
        .B(_f_permutation__round__c[602] ), .Z(_f_permutation__round_out[28])
         );
  XOR2_X2 _f_permutation__round__U4138  ( .A(_f_permutation__round__N5701 ), 
        .B(_f_permutation__round__c[603] ), .Z(_f_permutation__round_out[29])
         );
  XOR2_X2 _f_permutation__round__U4137  ( .A(_f_permutation__round__N5699 ), 
        .B(_f_permutation__round__c[604] ), .Z(_f_permutation__round_out[30])
         );
  XOR2_X2 _f_permutation__round__U4136  ( .A(_f_permutation__round__N5697 ), 
        .B(_f_permutation__round__c[605] ), .Z(_f_permutation__round_out[31])
         );
  XOR2_X2 _f_permutation__round__U4135  ( .A(_f_permutation__round__N5695 ), 
        .B(_f_permutation__round__c[606] ), .Z(_f_permutation__round_out[32])
         );
  XOR2_X2 _f_permutation__round__U4134  ( .A(_f_permutation__round__N5693 ), 
        .B(_f_permutation__round__c[607] ), .Z(_f_permutation__round_out[33])
         );
  XOR2_X2 _f_permutation__round__U4133  ( .A(_f_permutation__round__N5691 ), 
        .B(_f_permutation__round__c[608] ), .Z(_f_permutation__round_out[34])
         );
  XOR2_X2 _f_permutation__round__U4132  ( .A(_f_permutation__round__N5689 ), 
        .B(_f_permutation__round__c[609] ), .Z(_f_permutation__round_out[35])
         );
  XOR2_X2 _f_permutation__round__U4131  ( .A(_f_permutation__round__N5687 ), 
        .B(_f_permutation__round__c[610] ), .Z(_f_permutation__round_out[36])
         );
  XOR2_X2 _f_permutation__round__U4130  ( .A(_f_permutation__round__N5685 ), 
        .B(_f_permutation__round__c[611] ), .Z(_f_permutation__round_out[37])
         );
  XOR2_X2 _f_permutation__round__U4129  ( .A(_f_permutation__round__N5683 ), 
        .B(_f_permutation__round__c[612] ), .Z(_f_permutation__round_out[38])
         );
  XOR2_X2 _f_permutation__round__U4128  ( .A(_f_permutation__round__N5681 ), 
        .B(_f_permutation__round__c[613] ), .Z(_f_permutation__round_out[39])
         );
  XOR2_X2 _f_permutation__round__U4127  ( .A(_f_permutation__round__N5679 ), 
        .B(_f_permutation__round__c[614] ), .Z(_f_permutation__round_out[40])
         );
  XOR2_X2 _f_permutation__round__U4126  ( .A(_f_permutation__round__N5677 ), 
        .B(_f_permutation__round__c[615] ), .Z(_f_permutation__round_out[41])
         );
  XOR2_X2 _f_permutation__round__U4125  ( .A(_f_permutation__round__N5675 ), 
        .B(_f_permutation__round__c[616] ), .Z(_f_permutation__round_out[42])
         );
  XOR2_X2 _f_permutation__round__U4124  ( .A(_f_permutation__round__N5673 ), 
        .B(_f_permutation__round__c[617] ), .Z(_f_permutation__round_out[43])
         );
  XOR2_X2 _f_permutation__round__U4123  ( .A(_f_permutation__round__N5671 ), 
        .B(_f_permutation__round__c[618] ), .Z(_f_permutation__round_out[44])
         );
  XOR2_X2 _f_permutation__round__U4122  ( .A(_f_permutation__round__N5669 ), 
        .B(_f_permutation__round__c[619] ), .Z(_f_permutation__round_out[45])
         );
  XOR2_X2 _f_permutation__round__U4121  ( .A(_f_permutation__round__N5667 ), 
        .B(_f_permutation__round__c[620] ), .Z(_f_permutation__round_out[46])
         );
  XOR2_X2 _f_permutation__round__U4120  ( .A(_f_permutation__round__N5665 ), 
        .B(_f_permutation__round__c[621] ), .Z(_f_permutation__round_out[47])
         );
  XOR2_X2 _f_permutation__round__U4119  ( .A(_f_permutation__round__N5663 ), 
        .B(_f_permutation__round__c[622] ), .Z(_f_permutation__round_out[48])
         );
  XOR2_X2 _f_permutation__round__U4118  ( .A(_f_permutation__round__N5661 ), 
        .B(_f_permutation__round__c[623] ), .Z(_f_permutation__round_out[49])
         );
  XOR2_X2 _f_permutation__round__U4117  ( .A(_f_permutation__round__N5659 ), 
        .B(_f_permutation__round__c[624] ), .Z(_f_permutation__round_out[50])
         );
  XOR2_X2 _f_permutation__round__U4116  ( .A(_f_permutation__round__N5657 ), 
        .B(_f_permutation__round__c[625] ), .Z(_f_permutation__round_out[51])
         );
  XOR2_X2 _f_permutation__round__U4115  ( .A(_f_permutation__round__N5655 ), 
        .B(_f_permutation__round__c[626] ), .Z(_f_permutation__round_out[52])
         );
  XOR2_X2 _f_permutation__round__U4114  ( .A(_f_permutation__round__N5653 ), 
        .B(_f_permutation__round__c[627] ), .Z(_f_permutation__round_out[53])
         );
  XOR2_X2 _f_permutation__round__U4113  ( .A(_f_permutation__round__N5651 ), 
        .B(_f_permutation__round__c[628] ), .Z(_f_permutation__round_out[54])
         );
  XOR2_X2 _f_permutation__round__U4112  ( .A(_f_permutation__round__N5649 ), 
        .B(_f_permutation__round__c[629] ), .Z(_f_permutation__round_out[55])
         );
  XOR2_X2 _f_permutation__round__U4111  ( .A(_f_permutation__round__N5647 ), 
        .B(_f_permutation__round__c[630] ), .Z(_f_permutation__round_out[56])
         );
  XOR2_X2 _f_permutation__round__U4110  ( .A(_f_permutation__round__N5645 ), 
        .B(_f_permutation__round__c[631] ), .Z(_f_permutation__round_out[57])
         );
  XOR2_X2 _f_permutation__round__U4109  ( .A(_f_permutation__round__N5643 ), 
        .B(_f_permutation__round__c[632] ), .Z(_f_permutation__round_out[58])
         );
  XOR2_X2 _f_permutation__round__U4108  ( .A(_f_permutation__round__N5641 ), 
        .B(_f_permutation__round__c[633] ), .Z(_f_permutation__round_out[59])
         );
  XOR2_X2 _f_permutation__round__U4107  ( .A(_f_permutation__round__N5639 ), 
        .B(_f_permutation__round__c[634] ), .Z(_f_permutation__round_out[60])
         );
  XOR2_X2 _f_permutation__round__U4106  ( .A(_f_permutation__round__N5637 ), 
        .B(_f_permutation__round__c[635] ), .Z(_f_permutation__round_out[61])
         );
  XOR2_X2 _f_permutation__round__U4105  ( .A(_f_permutation__round__N5635 ), 
        .B(_f_permutation__round__c[636] ), .Z(_f_permutation__round_out[62])
         );
  XOR2_X2 _f_permutation__round__U4104  ( .A(_f_permutation__round__N5633 ), 
        .B(_f_permutation__round__c[637] ), .Z(_f_permutation__round_out[63])
         );
  XOR2_X2 _f_permutation__round__U4103  ( .A(_f_permutation__round__N5631 ), 
        .B(_f_permutation__round__c[215] ), .Z(_f_permutation__round_out[64])
         );
  XOR2_X2 _f_permutation__round__U4102  ( .A(_f_permutation__round__N5629 ), 
        .B(_f_permutation__round__c[216] ), .Z(_f_permutation__round_out[65])
         );
  XOR2_X2 _f_permutation__round__U4101  ( .A(_f_permutation__round__N5627 ), 
        .B(_f_permutation__round__c[217] ), .Z(_f_permutation__round_out[66])
         );
  XOR2_X2 _f_permutation__round__U4100  ( .A(_f_permutation__round__N5625 ), 
        .B(_f_permutation__round__c[218] ), .Z(_f_permutation__round_out[67])
         );
  XOR2_X2 _f_permutation__round__U4099  ( .A(_f_permutation__round__N5623 ), 
        .B(_f_permutation__round__c[219] ), .Z(_f_permutation__round_out[68])
         );
  XOR2_X2 _f_permutation__round__U4098  ( .A(_f_permutation__round__N5621 ), 
        .B(_f_permutation__round__c[220] ), .Z(_f_permutation__round_out[69])
         );
  XOR2_X2 _f_permutation__round__U4097  ( .A(_f_permutation__round__N5619 ), 
        .B(_f_permutation__round__c[221] ), .Z(_f_permutation__round_out[70])
         );
  XOR2_X2 _f_permutation__round__U4096  ( .A(_f_permutation__round__N5617 ), 
        .B(_f_permutation__round__c[222] ), .Z(_f_permutation__round_out[71])
         );
  XOR2_X2 _f_permutation__round__U4095  ( .A(_f_permutation__round__N5615 ), 
        .B(_f_permutation__round__c[223] ), .Z(_f_permutation__round_out[72])
         );
  XOR2_X2 _f_permutation__round__U4094  ( .A(_f_permutation__round__N5613 ), 
        .B(_f_permutation__round__c[224] ), .Z(_f_permutation__round_out[73])
         );
  XOR2_X2 _f_permutation__round__U4093  ( .A(_f_permutation__round__N5611 ), 
        .B(_f_permutation__round__c[225] ), .Z(_f_permutation__round_out[74])
         );
  XOR2_X2 _f_permutation__round__U4092  ( .A(_f_permutation__round__N5609 ), 
        .B(_f_permutation__round__c[226] ), .Z(_f_permutation__round_out[75])
         );
  XOR2_X2 _f_permutation__round__U4091  ( .A(_f_permutation__round__N5607 ), 
        .B(_f_permutation__round__c[227] ), .Z(_f_permutation__round_out[76])
         );
  XOR2_X2 _f_permutation__round__U4090  ( .A(_f_permutation__round__N5605 ), 
        .B(_f_permutation__round__c[228] ), .Z(_f_permutation__round_out[77])
         );
  XOR2_X2 _f_permutation__round__U4089  ( .A(_f_permutation__round__N5603 ), 
        .B(_f_permutation__round__c[229] ), .Z(_f_permutation__round_out[78])
         );
  XOR2_X2 _f_permutation__round__U4088  ( .A(_f_permutation__round__N5601 ), 
        .B(_f_permutation__round__c[230] ), .Z(_f_permutation__round_out[79])
         );
  XOR2_X2 _f_permutation__round__U4087  ( .A(_f_permutation__round__N5599 ), 
        .B(_f_permutation__round__c[231] ), .Z(_f_permutation__round_out[80])
         );
  XOR2_X2 _f_permutation__round__U4086  ( .A(_f_permutation__round__N5597 ), 
        .B(_f_permutation__round__c[232] ), .Z(_f_permutation__round_out[81])
         );
  XOR2_X2 _f_permutation__round__U4085  ( .A(_f_permutation__round__N5595 ), 
        .B(_f_permutation__round__c[233] ), .Z(_f_permutation__round_out[82])
         );
  XOR2_X2 _f_permutation__round__U4084  ( .A(_f_permutation__round__N5593 ), 
        .B(_f_permutation__round__c[234] ), .Z(_f_permutation__round_out[83])
         );
  XOR2_X2 _f_permutation__round__U4083  ( .A(_f_permutation__round__N5591 ), 
        .B(_f_permutation__round__c[235] ), .Z(_f_permutation__round_out[84])
         );
  XOR2_X2 _f_permutation__round__U4082  ( .A(_f_permutation__round__N5589 ), 
        .B(_f_permutation__round__c[236] ), .Z(_f_permutation__round_out[85])
         );
  XOR2_X2 _f_permutation__round__U4081  ( .A(_f_permutation__round__N5587 ), 
        .B(_f_permutation__round__c[237] ), .Z(_f_permutation__round_out[86])
         );
  XOR2_X2 _f_permutation__round__U4080  ( .A(_f_permutation__round__N5585 ), 
        .B(_f_permutation__round__c[238] ), .Z(_f_permutation__round_out[87])
         );
  XOR2_X2 _f_permutation__round__U4079  ( .A(_f_permutation__round__N5583 ), 
        .B(_f_permutation__round__c[239] ), .Z(_f_permutation__round_out[88])
         );
  XOR2_X2 _f_permutation__round__U4078  ( .A(_f_permutation__round__N5581 ), 
        .B(_f_permutation__round__c[240] ), .Z(_f_permutation__round_out[89])
         );
  XOR2_X2 _f_permutation__round__U4077  ( .A(_f_permutation__round__N5579 ), 
        .B(_f_permutation__round__c[241] ), .Z(_f_permutation__round_out[90])
         );
  XOR2_X2 _f_permutation__round__U4076  ( .A(_f_permutation__round__N5577 ), 
        .B(_f_permutation__round__c[242] ), .Z(_f_permutation__round_out[91])
         );
  XOR2_X2 _f_permutation__round__U4075  ( .A(_f_permutation__round__N5575 ), 
        .B(_f_permutation__round__c[243] ), .Z(_f_permutation__round_out[92])
         );
  XOR2_X2 _f_permutation__round__U4074  ( .A(_f_permutation__round__N5573 ), 
        .B(_f_permutation__round__c[244] ), .Z(_f_permutation__round_out[93])
         );
  XOR2_X2 _f_permutation__round__U4073  ( .A(_f_permutation__round__N5571 ), 
        .B(_f_permutation__round__c[245] ), .Z(_f_permutation__round_out[94])
         );
  XOR2_X2 _f_permutation__round__U4072  ( .A(_f_permutation__round__N5569 ), 
        .B(_f_permutation__round__c[246] ), .Z(_f_permutation__round_out[95])
         );
  XOR2_X2 _f_permutation__round__U4071  ( .A(_f_permutation__round__N5567 ), 
        .B(_f_permutation__round__c[247] ), .Z(_f_permutation__round_out[96])
         );
  XOR2_X2 _f_permutation__round__U4070  ( .A(_f_permutation__round__N5565 ), 
        .B(_f_permutation__round__c[248] ), .Z(_f_permutation__round_out[97])
         );
  XOR2_X2 _f_permutation__round__U4069  ( .A(_f_permutation__round__N5563 ), 
        .B(_f_permutation__round__c[249] ), .Z(_f_permutation__round_out[98])
         );
  XOR2_X2 _f_permutation__round__U4068  ( .A(_f_permutation__round__N5561 ), 
        .B(_f_permutation__round__c[250] ), .Z(_f_permutation__round_out[99])
         );
  XOR2_X2 _f_permutation__round__U4067  ( .A(_f_permutation__round__N5559 ), 
        .B(_f_permutation__round__c[251] ), .Z(_f_permutation__round_out[100]) );
  XOR2_X2 _f_permutation__round__U4066  ( .A(_f_permutation__round__N5557 ), 
        .B(_f_permutation__round__c[252] ), .Z(_f_permutation__round_out[101]) );
  XOR2_X2 _f_permutation__round__U4065  ( .A(_f_permutation__round__N5555 ), 
        .B(_f_permutation__round__c[253] ), .Z(_f_permutation__round_out[102]) );
  XOR2_X2 _f_permutation__round__U4064  ( .A(_f_permutation__round__N5553 ), 
        .B(_f_permutation__round__c[254] ), .Z(_f_permutation__round_out[103]) );
  XOR2_X2 _f_permutation__round__U4063  ( .A(_f_permutation__round__N5551 ), 
        .B(_f_permutation__round__c[255] ), .Z(_f_permutation__round_out[104]) );
  XOR2_X2 _f_permutation__round__U4062  ( .A(_f_permutation__round__N5549 ), 
        .B(_f_permutation__round__c[192] ), .Z(_f_permutation__round_out[105]) );
  XOR2_X2 _f_permutation__round__U4061  ( .A(_f_permutation__round__N5547 ), 
        .B(_f_permutation__round__c[193] ), .Z(_f_permutation__round_out[106]) );
  XOR2_X2 _f_permutation__round__U4060  ( .A(_f_permutation__round__N5545 ), 
        .B(_f_permutation__round__c[194] ), .Z(_f_permutation__round_out[107]) );
  XOR2_X2 _f_permutation__round__U4059  ( .A(_f_permutation__round__N5543 ), 
        .B(_f_permutation__round__c[195] ), .Z(_f_permutation__round_out[108]) );
  XOR2_X2 _f_permutation__round__U4058  ( .A(_f_permutation__round__N5541 ), 
        .B(_f_permutation__round__c[196] ), .Z(_f_permutation__round_out[109]) );
  XOR2_X2 _f_permutation__round__U4057  ( .A(_f_permutation__round__N5539 ), 
        .B(_f_permutation__round__c[197] ), .Z(_f_permutation__round_out[110]) );
  XOR2_X2 _f_permutation__round__U4056  ( .A(_f_permutation__round__N5537 ), 
        .B(_f_permutation__round__c[198] ), .Z(_f_permutation__round_out[111]) );
  XOR2_X2 _f_permutation__round__U4055  ( .A(_f_permutation__round__N5535 ), 
        .B(_f_permutation__round__c[199] ), .Z(_f_permutation__round_out[112]) );
  XOR2_X2 _f_permutation__round__U4054  ( .A(_f_permutation__round__N5533 ), 
        .B(_f_permutation__round__c[200] ), .Z(_f_permutation__round_out[113]) );
  XOR2_X2 _f_permutation__round__U4053  ( .A(_f_permutation__round__N5531 ), 
        .B(_f_permutation__round__c[201] ), .Z(_f_permutation__round_out[114]) );
  XOR2_X2 _f_permutation__round__U4052  ( .A(_f_permutation__round__N5529 ), 
        .B(_f_permutation__round__c[202] ), .Z(_f_permutation__round_out[115]) );
  XOR2_X2 _f_permutation__round__U4051  ( .A(_f_permutation__round__N5527 ), 
        .B(_f_permutation__round__c[203] ), .Z(_f_permutation__round_out[116]) );
  XOR2_X2 _f_permutation__round__U4050  ( .A(_f_permutation__round__N5525 ), 
        .B(_f_permutation__round__c[204] ), .Z(_f_permutation__round_out[117]) );
  XOR2_X2 _f_permutation__round__U4049  ( .A(_f_permutation__round__N5523 ), 
        .B(_f_permutation__round__c[205] ), .Z(_f_permutation__round_out[118]) );
  XOR2_X2 _f_permutation__round__U4048  ( .A(_f_permutation__round__N5521 ), 
        .B(_f_permutation__round__c[206] ), .Z(_f_permutation__round_out[119]) );
  XOR2_X2 _f_permutation__round__U4047  ( .A(_f_permutation__round__N5519 ), 
        .B(_f_permutation__round__c[207] ), .Z(_f_permutation__round_out[120]) );
  XOR2_X2 _f_permutation__round__U4046  ( .A(_f_permutation__round__N5517 ), 
        .B(_f_permutation__round__c[208] ), .Z(_f_permutation__round_out[121]) );
  XOR2_X2 _f_permutation__round__U4045  ( .A(_f_permutation__round__N5515 ), 
        .B(_f_permutation__round__c[209] ), .Z(_f_permutation__round_out[122]) );
  XOR2_X2 _f_permutation__round__U4044  ( .A(_f_permutation__round__N5513 ), 
        .B(_f_permutation__round__c[210] ), .Z(_f_permutation__round_out[123]) );
  XOR2_X2 _f_permutation__round__U4043  ( .A(_f_permutation__round__N5511 ), 
        .B(_f_permutation__round__c[211] ), .Z(_f_permutation__round_out[124]) );
  XOR2_X2 _f_permutation__round__U4042  ( .A(_f_permutation__round__N5509 ), 
        .B(_f_permutation__round__c[212] ), .Z(_f_permutation__round_out[125]) );
  XOR2_X2 _f_permutation__round__U4041  ( .A(_f_permutation__round__N5507 ), 
        .B(_f_permutation__round__c[213] ), .Z(_f_permutation__round_out[126]) );
  XOR2_X2 _f_permutation__round__U4040  ( .A(_f_permutation__round__N5505 ), 
        .B(_f_permutation__round__c[214] ), .Z(_f_permutation__round_out[127]) );
  XOR2_X2 _f_permutation__round__U4039  ( .A(_f_permutation__round__N5503 ), 
        .B(_f_permutation__round__c[1433] ), .Z(
        _f_permutation__round_out[128]) );
  XOR2_X2 _f_permutation__round__U4038  ( .A(_f_permutation__round__N5501 ), 
        .B(_f_permutation__round__c[1434] ), .Z(
        _f_permutation__round_out[129]) );
  XOR2_X2 _f_permutation__round__U4037  ( .A(_f_permutation__round__N5499 ), 
        .B(_f_permutation__round__c[1435] ), .Z(
        _f_permutation__round_out[130]) );
  XOR2_X2 _f_permutation__round__U4036  ( .A(_f_permutation__round__N5497 ), 
        .B(_f_permutation__round__c[1436] ), .Z(
        _f_permutation__round_out[131]) );
  XOR2_X2 _f_permutation__round__U4035  ( .A(_f_permutation__round__N5495 ), 
        .B(_f_permutation__round__c[1437] ), .Z(
        _f_permutation__round_out[132]) );
  XOR2_X2 _f_permutation__round__U4034  ( .A(_f_permutation__round__N5493 ), 
        .B(_f_permutation__round__c[1438] ), .Z(
        _f_permutation__round_out[133]) );
  XOR2_X2 _f_permutation__round__U4033  ( .A(_f_permutation__round__N5491 ), 
        .B(_f_permutation__round__c[1439] ), .Z(
        _f_permutation__round_out[134]) );
  XOR2_X2 _f_permutation__round__U4032  ( .A(_f_permutation__round__N5489 ), 
        .B(_f_permutation__round__c[1440] ), .Z(
        _f_permutation__round_out[135]) );
  XOR2_X2 _f_permutation__round__U4031  ( .A(_f_permutation__round__N5487 ), 
        .B(_f_permutation__round__c[1441] ), .Z(
        _f_permutation__round_out[136]) );
  XOR2_X2 _f_permutation__round__U4030  ( .A(_f_permutation__round__N5485 ), 
        .B(_f_permutation__round__c[1442] ), .Z(
        _f_permutation__round_out[137]) );
  XOR2_X2 _f_permutation__round__U4029  ( .A(_f_permutation__round__N5483 ), 
        .B(_f_permutation__round__c[1443] ), .Z(
        _f_permutation__round_out[138]) );
  XOR2_X2 _f_permutation__round__U4028  ( .A(_f_permutation__round__N5481 ), 
        .B(_f_permutation__round__c[1444] ), .Z(
        _f_permutation__round_out[139]) );
  XOR2_X2 _f_permutation__round__U4027  ( .A(_f_permutation__round__N5479 ), 
        .B(_f_permutation__round__c[1445] ), .Z(
        _f_permutation__round_out[140]) );
  XOR2_X2 _f_permutation__round__U4026  ( .A(_f_permutation__round__N5477 ), 
        .B(_f_permutation__round__c[1446] ), .Z(
        _f_permutation__round_out[141]) );
  XOR2_X2 _f_permutation__round__U4025  ( .A(_f_permutation__round__N5475 ), 
        .B(_f_permutation__round__c[1447] ), .Z(
        _f_permutation__round_out[142]) );
  XOR2_X2 _f_permutation__round__U4024  ( .A(_f_permutation__round__N5473 ), 
        .B(_f_permutation__round__c[1448] ), .Z(
        _f_permutation__round_out[143]) );
  XOR2_X2 _f_permutation__round__U4023  ( .A(_f_permutation__round__N5471 ), 
        .B(_f_permutation__round__c[1449] ), .Z(
        _f_permutation__round_out[144]) );
  XOR2_X2 _f_permutation__round__U4022  ( .A(_f_permutation__round__N5469 ), 
        .B(_f_permutation__round__c[1450] ), .Z(
        _f_permutation__round_out[145]) );
  XOR2_X2 _f_permutation__round__U4021  ( .A(_f_permutation__round__N5467 ), 
        .B(_f_permutation__round__c[1451] ), .Z(
        _f_permutation__round_out[146]) );
  XOR2_X2 _f_permutation__round__U4020  ( .A(_f_permutation__round__N5465 ), 
        .B(_f_permutation__round__c[1452] ), .Z(
        _f_permutation__round_out[147]) );
  XOR2_X2 _f_permutation__round__U4019  ( .A(_f_permutation__round__N5463 ), 
        .B(_f_permutation__round__c[1453] ), .Z(
        _f_permutation__round_out[148]) );
  XOR2_X2 _f_permutation__round__U4018  ( .A(_f_permutation__round__N5461 ), 
        .B(_f_permutation__round__c[1454] ), .Z(
        _f_permutation__round_out[149]) );
  XOR2_X2 _f_permutation__round__U4017  ( .A(_f_permutation__round__N5459 ), 
        .B(_f_permutation__round__c[1455] ), .Z(
        _f_permutation__round_out[150]) );
  XOR2_X2 _f_permutation__round__U4016  ( .A(_f_permutation__round__N5457 ), 
        .B(_f_permutation__round__c[1456] ), .Z(
        _f_permutation__round_out[151]) );
  XOR2_X2 _f_permutation__round__U4015  ( .A(_f_permutation__round__N5455 ), 
        .B(_f_permutation__round__c[1457] ), .Z(
        _f_permutation__round_out[152]) );
  XOR2_X2 _f_permutation__round__U4014  ( .A(_f_permutation__round__N5453 ), 
        .B(_f_permutation__round__c[1458] ), .Z(
        _f_permutation__round_out[153]) );
  XOR2_X2 _f_permutation__round__U4013  ( .A(_f_permutation__round__N5451 ), 
        .B(_f_permutation__round__c[1459] ), .Z(
        _f_permutation__round_out[154]) );
  XOR2_X2 _f_permutation__round__U4012  ( .A(_f_permutation__round__N5449 ), 
        .B(_f_permutation__round__c[1460] ), .Z(
        _f_permutation__round_out[155]) );
  XOR2_X2 _f_permutation__round__U4011  ( .A(_f_permutation__round__N5447 ), 
        .B(_f_permutation__round__c[1461] ), .Z(
        _f_permutation__round_out[156]) );
  XOR2_X2 _f_permutation__round__U4010  ( .A(_f_permutation__round__N5445 ), 
        .B(_f_permutation__round__c[1462] ), .Z(
        _f_permutation__round_out[157]) );
  XOR2_X2 _f_permutation__round__U4009  ( .A(_f_permutation__round__N5443 ), 
        .B(_f_permutation__round__c[1463] ), .Z(
        _f_permutation__round_out[158]) );
  XOR2_X2 _f_permutation__round__U4008  ( .A(_f_permutation__round__N5441 ), 
        .B(_f_permutation__round__c[1464] ), .Z(
        _f_permutation__round_out[159]) );
  XOR2_X2 _f_permutation__round__U4007  ( .A(_f_permutation__round__N5439 ), 
        .B(_f_permutation__round__c[1465] ), .Z(
        _f_permutation__round_out[160]) );
  XOR2_X2 _f_permutation__round__U4006  ( .A(_f_permutation__round__N5437 ), 
        .B(_f_permutation__round__c[1466] ), .Z(
        _f_permutation__round_out[161]) );
  XOR2_X2 _f_permutation__round__U4005  ( .A(_f_permutation__round__N5435 ), 
        .B(_f_permutation__round__c[1467] ), .Z(
        _f_permutation__round_out[162]) );
  XOR2_X2 _f_permutation__round__U4004  ( .A(_f_permutation__round__N5433 ), 
        .B(_f_permutation__round__c[1468] ), .Z(
        _f_permutation__round_out[163]) );
  XOR2_X2 _f_permutation__round__U4003  ( .A(_f_permutation__round__N5431 ), 
        .B(_f_permutation__round__c[1469] ), .Z(
        _f_permutation__round_out[164]) );
  XOR2_X2 _f_permutation__round__U4002  ( .A(_f_permutation__round__N5429 ), 
        .B(_f_permutation__round__c[1470] ), .Z(
        _f_permutation__round_out[165]) );
  XOR2_X2 _f_permutation__round__U4001  ( .A(_f_permutation__round__N5427 ), 
        .B(_f_permutation__round__c[1471] ), .Z(
        _f_permutation__round_out[166]) );
  XOR2_X2 _f_permutation__round__U4000  ( .A(_f_permutation__round__N5425 ), 
        .B(_f_permutation__round__c[1408] ), .Z(
        _f_permutation__round_out[167]) );
  XOR2_X2 _f_permutation__round__U3999  ( .A(_f_permutation__round__N5423 ), 
        .B(_f_permutation__round__c[1409] ), .Z(
        _f_permutation__round_out[168]) );
  XOR2_X2 _f_permutation__round__U3998  ( .A(_f_permutation__round__N5421 ), 
        .B(_f_permutation__round__c[1410] ), .Z(
        _f_permutation__round_out[169]) );
  XOR2_X2 _f_permutation__round__U3997  ( .A(_f_permutation__round__N5419 ), 
        .B(_f_permutation__round__c[1411] ), .Z(
        _f_permutation__round_out[170]) );
  XOR2_X2 _f_permutation__round__U3996  ( .A(_f_permutation__round__N5417 ), 
        .B(_f_permutation__round__c[1412] ), .Z(
        _f_permutation__round_out[171]) );
  XOR2_X2 _f_permutation__round__U3995  ( .A(_f_permutation__round__N5415 ), 
        .B(_f_permutation__round__c[1413] ), .Z(
        _f_permutation__round_out[172]) );
  XOR2_X2 _f_permutation__round__U3994  ( .A(_f_permutation__round__N5413 ), 
        .B(_f_permutation__round__c[1414] ), .Z(
        _f_permutation__round_out[173]) );
  XOR2_X2 _f_permutation__round__U3993  ( .A(_f_permutation__round__N5411 ), 
        .B(_f_permutation__round__c[1415] ), .Z(
        _f_permutation__round_out[174]) );
  XOR2_X2 _f_permutation__round__U3992  ( .A(_f_permutation__round__N5409 ), 
        .B(_f_permutation__round__c[1416] ), .Z(
        _f_permutation__round_out[175]) );
  XOR2_X2 _f_permutation__round__U3991  ( .A(_f_permutation__round__N5407 ), 
        .B(_f_permutation__round__c[1417] ), .Z(
        _f_permutation__round_out[176]) );
  XOR2_X2 _f_permutation__round__U3990  ( .A(_f_permutation__round__N5405 ), 
        .B(_f_permutation__round__c[1418] ), .Z(
        _f_permutation__round_out[177]) );
  XOR2_X2 _f_permutation__round__U3989  ( .A(_f_permutation__round__N5403 ), 
        .B(_f_permutation__round__c[1419] ), .Z(
        _f_permutation__round_out[178]) );
  XOR2_X2 _f_permutation__round__U3988  ( .A(_f_permutation__round__N5401 ), 
        .B(_f_permutation__round__c[1420] ), .Z(
        _f_permutation__round_out[179]) );
  XOR2_X2 _f_permutation__round__U3987  ( .A(_f_permutation__round__N5399 ), 
        .B(_f_permutation__round__c[1421] ), .Z(
        _f_permutation__round_out[180]) );
  XOR2_X2 _f_permutation__round__U3986  ( .A(_f_permutation__round__N5397 ), 
        .B(_f_permutation__round__c[1422] ), .Z(
        _f_permutation__round_out[181]) );
  XOR2_X2 _f_permutation__round__U3985  ( .A(_f_permutation__round__N5395 ), 
        .B(_f_permutation__round__c[1423] ), .Z(
        _f_permutation__round_out[182]) );
  XOR2_X2 _f_permutation__round__U3984  ( .A(_f_permutation__round__N5393 ), 
        .B(_f_permutation__round__c[1424] ), .Z(
        _f_permutation__round_out[183]) );
  XOR2_X2 _f_permutation__round__U3983  ( .A(_f_permutation__round__N5391 ), 
        .B(_f_permutation__round__c[1425] ), .Z(
        _f_permutation__round_out[184]) );
  XOR2_X2 _f_permutation__round__U3982  ( .A(_f_permutation__round__N5389 ), 
        .B(_f_permutation__round__c[1426] ), .Z(
        _f_permutation__round_out[185]) );
  XOR2_X2 _f_permutation__round__U3981  ( .A(_f_permutation__round__N5387 ), 
        .B(_f_permutation__round__c[1427] ), .Z(
        _f_permutation__round_out[186]) );
  XOR2_X2 _f_permutation__round__U3980  ( .A(_f_permutation__round__N5385 ), 
        .B(_f_permutation__round__c[1428] ), .Z(
        _f_permutation__round_out[187]) );
  XOR2_X2 _f_permutation__round__U3979  ( .A(_f_permutation__round__N5383 ), 
        .B(_f_permutation__round__c[1429] ), .Z(
        _f_permutation__round_out[188]) );
  XOR2_X2 _f_permutation__round__U3978  ( .A(_f_permutation__round__N5381 ), 
        .B(_f_permutation__round__c[1430] ), .Z(
        _f_permutation__round_out[189]) );
  XOR2_X2 _f_permutation__round__U3977  ( .A(_f_permutation__round__N5379 ), 
        .B(_f_permutation__round__c[1431] ), .Z(
        _f_permutation__round_out[190]) );
  XOR2_X2 _f_permutation__round__U3976  ( .A(_f_permutation__round__N5377 ), 
        .B(_f_permutation__round__c[1432] ), .Z(
        _f_permutation__round_out[191]) );
  XOR2_X2 _f_permutation__round__U3975  ( .A(_f_permutation__round__N5375 ), 
        .B(_f_permutation__round__c[1033] ), .Z(
        _f_permutation__round_out[192]) );
  XOR2_X2 _f_permutation__round__U3974  ( .A(_f_permutation__round__N5373 ), 
        .B(_f_permutation__round__c[1034] ), .Z(
        _f_permutation__round_out[193]) );
  XOR2_X2 _f_permutation__round__U3973  ( .A(_f_permutation__round__N5371 ), 
        .B(_f_permutation__round__c[1035] ), .Z(
        _f_permutation__round_out[194]) );
  XOR2_X2 _f_permutation__round__U3972  ( .A(_f_permutation__round__N5369 ), 
        .B(_f_permutation__round__c[1036] ), .Z(
        _f_permutation__round_out[195]) );
  XOR2_X2 _f_permutation__round__U3971  ( .A(_f_permutation__round__N5367 ), 
        .B(_f_permutation__round__c[1037] ), .Z(
        _f_permutation__round_out[196]) );
  XOR2_X2 _f_permutation__round__U3970  ( .A(_f_permutation__round__N5365 ), 
        .B(_f_permutation__round__c[1038] ), .Z(
        _f_permutation__round_out[197]) );
  XOR2_X2 _f_permutation__round__U3969  ( .A(_f_permutation__round__N5363 ), 
        .B(_f_permutation__round__c[1039] ), .Z(
        _f_permutation__round_out[198]) );
  XOR2_X2 _f_permutation__round__U3968  ( .A(_f_permutation__round__N5361 ), 
        .B(_f_permutation__round__c[1040] ), .Z(
        _f_permutation__round_out[199]) );
  XOR2_X2 _f_permutation__round__U3967  ( .A(_f_permutation__round__N5359 ), 
        .B(_f_permutation__round__c[1041] ), .Z(
        _f_permutation__round_out[200]) );
  XOR2_X2 _f_permutation__round__U3966  ( .A(_f_permutation__round__N5357 ), 
        .B(_f_permutation__round__c[1042] ), .Z(
        _f_permutation__round_out[201]) );
  XOR2_X2 _f_permutation__round__U3965  ( .A(_f_permutation__round__N5355 ), 
        .B(_f_permutation__round__c[1043] ), .Z(
        _f_permutation__round_out[202]) );
  XOR2_X2 _f_permutation__round__U3964  ( .A(_f_permutation__round__N5353 ), 
        .B(_f_permutation__round__c[1044] ), .Z(
        _f_permutation__round_out[203]) );
  XOR2_X2 _f_permutation__round__U3963  ( .A(_f_permutation__round__N5351 ), 
        .B(_f_permutation__round__c[1045] ), .Z(
        _f_permutation__round_out[204]) );
  XOR2_X2 _f_permutation__round__U3962  ( .A(_f_permutation__round__N5349 ), 
        .B(_f_permutation__round__c[1046] ), .Z(
        _f_permutation__round_out[205]) );
  XOR2_X2 _f_permutation__round__U3961  ( .A(_f_permutation__round__N5347 ), 
        .B(_f_permutation__round__c[1047] ), .Z(
        _f_permutation__round_out[206]) );
  XOR2_X2 _f_permutation__round__U3960  ( .A(_f_permutation__round__N5345 ), 
        .B(_f_permutation__round__c[1048] ), .Z(
        _f_permutation__round_out[207]) );
  XOR2_X2 _f_permutation__round__U3959  ( .A(_f_permutation__round__N5343 ), 
        .B(_f_permutation__round__c[1049] ), .Z(
        _f_permutation__round_out[208]) );
  XOR2_X2 _f_permutation__round__U3958  ( .A(_f_permutation__round__N5341 ), 
        .B(_f_permutation__round__c[1050] ), .Z(
        _f_permutation__round_out[209]) );
  XOR2_X2 _f_permutation__round__U3957  ( .A(_f_permutation__round__N5339 ), 
        .B(_f_permutation__round__c[1051] ), .Z(
        _f_permutation__round_out[210]) );
  XOR2_X2 _f_permutation__round__U3956  ( .A(_f_permutation__round__N5337 ), 
        .B(_f_permutation__round__c[1052] ), .Z(
        _f_permutation__round_out[211]) );
  XOR2_X2 _f_permutation__round__U3955  ( .A(_f_permutation__round__N5335 ), 
        .B(_f_permutation__round__c[1053] ), .Z(
        _f_permutation__round_out[212]) );
  XOR2_X2 _f_permutation__round__U3954  ( .A(_f_permutation__round__N5333 ), 
        .B(_f_permutation__round__c[1054] ), .Z(
        _f_permutation__round_out[213]) );
  XOR2_X2 _f_permutation__round__U3953  ( .A(_f_permutation__round__N5331 ), 
        .B(_f_permutation__round__c[1055] ), .Z(
        _f_permutation__round_out[214]) );
  XOR2_X2 _f_permutation__round__U3952  ( .A(_f_permutation__round__N5329 ), 
        .B(_f_permutation__round__c[1056] ), .Z(
        _f_permutation__round_out[215]) );
  XOR2_X2 _f_permutation__round__U3951  ( .A(_f_permutation__round__N5327 ), 
        .B(_f_permutation__round__c[1057] ), .Z(
        _f_permutation__round_out[216]) );
  XOR2_X2 _f_permutation__round__U3950  ( .A(_f_permutation__round__N5325 ), 
        .B(_f_permutation__round__c[1058] ), .Z(
        _f_permutation__round_out[217]) );
  XOR2_X2 _f_permutation__round__U3949  ( .A(_f_permutation__round__N5323 ), 
        .B(_f_permutation__round__c[1059] ), .Z(
        _f_permutation__round_out[218]) );
  XOR2_X2 _f_permutation__round__U3948  ( .A(_f_permutation__round__N5321 ), 
        .B(_f_permutation__round__c[1060] ), .Z(
        _f_permutation__round_out[219]) );
  XOR2_X2 _f_permutation__round__U3947  ( .A(_f_permutation__round__N5319 ), 
        .B(_f_permutation__round__c[1061] ), .Z(
        _f_permutation__round_out[220]) );
  XOR2_X2 _f_permutation__round__U3946  ( .A(_f_permutation__round__N5317 ), 
        .B(_f_permutation__round__c[1062] ), .Z(
        _f_permutation__round_out[221]) );
  XOR2_X2 _f_permutation__round__U3945  ( .A(_f_permutation__round__N5315 ), 
        .B(_f_permutation__round__c[1063] ), .Z(
        _f_permutation__round_out[222]) );
  XOR2_X2 _f_permutation__round__U3944  ( .A(_f_permutation__round__N5313 ), 
        .B(_f_permutation__round__c[1064] ), .Z(
        _f_permutation__round_out[223]) );
  XOR2_X2 _f_permutation__round__U3943  ( .A(_f_permutation__round__N5311 ), 
        .B(_f_permutation__round__c[1065] ), .Z(
        _f_permutation__round_out[224]) );
  XOR2_X2 _f_permutation__round__U3942  ( .A(_f_permutation__round__N5309 ), 
        .B(_f_permutation__round__c[1066] ), .Z(
        _f_permutation__round_out[225]) );
  XOR2_X2 _f_permutation__round__U3941  ( .A(_f_permutation__round__N5307 ), 
        .B(_f_permutation__round__c[1067] ), .Z(
        _f_permutation__round_out[226]) );
  XOR2_X2 _f_permutation__round__U3940  ( .A(_f_permutation__round__N5305 ), 
        .B(_f_permutation__round__c[1068] ), .Z(
        _f_permutation__round_out[227]) );
  XOR2_X2 _f_permutation__round__U3939  ( .A(_f_permutation__round__N5303 ), 
        .B(_f_permutation__round__c[1069] ), .Z(
        _f_permutation__round_out[228]) );
  XOR2_X2 _f_permutation__round__U3938  ( .A(_f_permutation__round__N5301 ), 
        .B(_f_permutation__round__c[1070] ), .Z(
        _f_permutation__round_out[229]) );
  XOR2_X2 _f_permutation__round__U3937  ( .A(_f_permutation__round__N5299 ), 
        .B(_f_permutation__round__c[1071] ), .Z(
        _f_permutation__round_out[230]) );
  XOR2_X2 _f_permutation__round__U3936  ( .A(_f_permutation__round__N5297 ), 
        .B(_f_permutation__round__c[1072] ), .Z(
        _f_permutation__round_out[231]) );
  XOR2_X2 _f_permutation__round__U3935  ( .A(_f_permutation__round__N5295 ), 
        .B(_f_permutation__round__c[1073] ), .Z(
        _f_permutation__round_out[232]) );
  XOR2_X2 _f_permutation__round__U3934  ( .A(_f_permutation__round__N5293 ), 
        .B(_f_permutation__round__c[1074] ), .Z(
        _f_permutation__round_out[233]) );
  XOR2_X2 _f_permutation__round__U3933  ( .A(_f_permutation__round__N5291 ), 
        .B(_f_permutation__round__c[1075] ), .Z(
        _f_permutation__round_out[234]) );
  XOR2_X2 _f_permutation__round__U3932  ( .A(_f_permutation__round__N5289 ), 
        .B(_f_permutation__round__c[1076] ), .Z(
        _f_permutation__round_out[235]) );
  XOR2_X2 _f_permutation__round__U3931  ( .A(_f_permutation__round__N5287 ), 
        .B(_f_permutation__round__c[1077] ), .Z(
        _f_permutation__round_out[236]) );
  XOR2_X2 _f_permutation__round__U3930  ( .A(_f_permutation__round__N5285 ), 
        .B(_f_permutation__round__c[1078] ), .Z(
        _f_permutation__round_out[237]) );
  XOR2_X2 _f_permutation__round__U3929  ( .A(_f_permutation__round__N5283 ), 
        .B(_f_permutation__round__c[1079] ), .Z(
        _f_permutation__round_out[238]) );
  XOR2_X2 _f_permutation__round__U3928  ( .A(_f_permutation__round__N5281 ), 
        .B(_f_permutation__round__c[1080] ), .Z(
        _f_permutation__round_out[239]) );
  XOR2_X2 _f_permutation__round__U3927  ( .A(_f_permutation__round__N5279 ), 
        .B(_f_permutation__round__c[1081] ), .Z(
        _f_permutation__round_out[240]) );
  XOR2_X2 _f_permutation__round__U3926  ( .A(_f_permutation__round__N5277 ), 
        .B(_f_permutation__round__c[1082] ), .Z(
        _f_permutation__round_out[241]) );
  XOR2_X2 _f_permutation__round__U3925  ( .A(_f_permutation__round__N5275 ), 
        .B(_f_permutation__round__c[1083] ), .Z(
        _f_permutation__round_out[242]) );
  XOR2_X2 _f_permutation__round__U3924  ( .A(_f_permutation__round__N5273 ), 
        .B(_f_permutation__round__c[1084] ), .Z(
        _f_permutation__round_out[243]) );
  XOR2_X2 _f_permutation__round__U3923  ( .A(_f_permutation__round__N5271 ), 
        .B(_f_permutation__round__c[1085] ), .Z(
        _f_permutation__round_out[244]) );
  XOR2_X2 _f_permutation__round__U3922  ( .A(_f_permutation__round__N5269 ), 
        .B(_f_permutation__round__c[1086] ), .Z(
        _f_permutation__round_out[245]) );
  XOR2_X2 _f_permutation__round__U3921  ( .A(_f_permutation__round__N5267 ), 
        .B(_f_permutation__round__c[1087] ), .Z(
        _f_permutation__round_out[246]) );
  XOR2_X2 _f_permutation__round__U3920  ( .A(_f_permutation__round__N5265 ), 
        .B(_f_permutation__round__c[1024] ), .Z(
        _f_permutation__round_out[247]) );
  XOR2_X2 _f_permutation__round__U3919  ( .A(_f_permutation__round__N5263 ), 
        .B(_f_permutation__round__c[1025] ), .Z(
        _f_permutation__round_out[248]) );
  XOR2_X2 _f_permutation__round__U3918  ( .A(_f_permutation__round__N5261 ), 
        .B(_f_permutation__round__c[1026] ), .Z(
        _f_permutation__round_out[249]) );
  XOR2_X2 _f_permutation__round__U3917  ( .A(_f_permutation__round__N5259 ), 
        .B(_f_permutation__round__c[1027] ), .Z(
        _f_permutation__round_out[250]) );
  XOR2_X2 _f_permutation__round__U3916  ( .A(_f_permutation__round__N5257 ), 
        .B(_f_permutation__round__c[1028] ), .Z(
        _f_permutation__round_out[251]) );
  XOR2_X2 _f_permutation__round__U3915  ( .A(_f_permutation__round__N5255 ), 
        .B(_f_permutation__round__c[1029] ), .Z(
        _f_permutation__round_out[252]) );
  XOR2_X2 _f_permutation__round__U3914  ( .A(_f_permutation__round__N5253 ), 
        .B(_f_permutation__round__c[1030] ), .Z(
        _f_permutation__round_out[253]) );
  XOR2_X2 _f_permutation__round__U3913  ( .A(_f_permutation__round__N5251 ), 
        .B(_f_permutation__round__c[1031] ), .Z(
        _f_permutation__round_out[254]) );
  XOR2_X2 _f_permutation__round__U3912  ( .A(_f_permutation__round__N5249 ), 
        .B(_f_permutation__round__c[1032] ), .Z(
        _f_permutation__round_out[255]) );
  XOR2_X2 _f_permutation__round__U3911  ( .A(_f_permutation__round__N5247 ), 
        .B(_f_permutation__round__c[642] ), .Z(_f_permutation__round_out[256]) );
  XOR2_X2 _f_permutation__round__U3910  ( .A(_f_permutation__round__N5245 ), 
        .B(_f_permutation__round__c[643] ), .Z(_f_permutation__round_out[257]) );
  XOR2_X2 _f_permutation__round__U3909  ( .A(_f_permutation__round__N5243 ), 
        .B(_f_permutation__round__c[644] ), .Z(_f_permutation__round_out[258]) );
  XOR2_X2 _f_permutation__round__U3908  ( .A(_f_permutation__round__N5241 ), 
        .B(_f_permutation__round__c[645] ), .Z(_f_permutation__round_out[259]) );
  XOR2_X2 _f_permutation__round__U3907  ( .A(_f_permutation__round__N5239 ), 
        .B(_f_permutation__round__c[646] ), .Z(_f_permutation__round_out[260]) );
  XOR2_X2 _f_permutation__round__U3906  ( .A(_f_permutation__round__N5237 ), 
        .B(_f_permutation__round__c[647] ), .Z(_f_permutation__round_out[261]) );
  XOR2_X2 _f_permutation__round__U3905  ( .A(_f_permutation__round__N5235 ), 
        .B(_f_permutation__round__c[648] ), .Z(_f_permutation__round_out[262]) );
  XOR2_X2 _f_permutation__round__U3904  ( .A(_f_permutation__round__N5233 ), 
        .B(_f_permutation__round__c[649] ), .Z(_f_permutation__round_out[263]) );
  XOR2_X2 _f_permutation__round__U3903  ( .A(_f_permutation__round__N5231 ), 
        .B(_f_permutation__round__c[650] ), .Z(_f_permutation__round_out[264]) );
  XOR2_X2 _f_permutation__round__U3902  ( .A(_f_permutation__round__N5229 ), 
        .B(_f_permutation__round__c[651] ), .Z(_f_permutation__round_out[265]) );
  XOR2_X2 _f_permutation__round__U3901  ( .A(_f_permutation__round__N5227 ), 
        .B(_f_permutation__round__c[652] ), .Z(_f_permutation__round_out[266]) );
  XOR2_X2 _f_permutation__round__U3900  ( .A(_f_permutation__round__N5225 ), 
        .B(_f_permutation__round__c[653] ), .Z(_f_permutation__round_out[267]) );
  XOR2_X2 _f_permutation__round__U3899  ( .A(_f_permutation__round__N5223 ), 
        .B(_f_permutation__round__c[654] ), .Z(_f_permutation__round_out[268]) );
  XOR2_X2 _f_permutation__round__U3898  ( .A(_f_permutation__round__N5221 ), 
        .B(_f_permutation__round__c[655] ), .Z(_f_permutation__round_out[269]) );
  XOR2_X2 _f_permutation__round__U3897  ( .A(_f_permutation__round__N5219 ), 
        .B(_f_permutation__round__c[656] ), .Z(_f_permutation__round_out[270]) );
  XOR2_X2 _f_permutation__round__U3896  ( .A(_f_permutation__round__N5217 ), 
        .B(_f_permutation__round__c[657] ), .Z(_f_permutation__round_out[271]) );
  XOR2_X2 _f_permutation__round__U3895  ( .A(_f_permutation__round__N5215 ), 
        .B(_f_permutation__round__c[658] ), .Z(_f_permutation__round_out[272]) );
  XOR2_X2 _f_permutation__round__U3894  ( .A(_f_permutation__round__N5213 ), 
        .B(_f_permutation__round__c[659] ), .Z(_f_permutation__round_out[273]) );
  XOR2_X2 _f_permutation__round__U3893  ( .A(_f_permutation__round__N5211 ), 
        .B(_f_permutation__round__c[660] ), .Z(_f_permutation__round_out[274]) );
  XOR2_X2 _f_permutation__round__U3892  ( .A(_f_permutation__round__N5209 ), 
        .B(_f_permutation__round__c[661] ), .Z(_f_permutation__round_out[275]) );
  XOR2_X2 _f_permutation__round__U3891  ( .A(_f_permutation__round__N5207 ), 
        .B(_f_permutation__round__c[662] ), .Z(_f_permutation__round_out[276]) );
  XOR2_X2 _f_permutation__round__U3890  ( .A(_f_permutation__round__N5205 ), 
        .B(_f_permutation__round__c[663] ), .Z(_f_permutation__round_out[277]) );
  XOR2_X2 _f_permutation__round__U3889  ( .A(_f_permutation__round__N5203 ), 
        .B(_f_permutation__round__c[664] ), .Z(_f_permutation__round_out[278]) );
  XOR2_X2 _f_permutation__round__U3888  ( .A(_f_permutation__round__N5201 ), 
        .B(_f_permutation__round__c[665] ), .Z(_f_permutation__round_out[279]) );
  XOR2_X2 _f_permutation__round__U3887  ( .A(_f_permutation__round__N5199 ), 
        .B(_f_permutation__round__c[666] ), .Z(_f_permutation__round_out[280]) );
  XOR2_X2 _f_permutation__round__U3886  ( .A(_f_permutation__round__N5197 ), 
        .B(_f_permutation__round__c[667] ), .Z(_f_permutation__round_out[281]) );
  XOR2_X2 _f_permutation__round__U3885  ( .A(_f_permutation__round__N5195 ), 
        .B(_f_permutation__round__c[668] ), .Z(_f_permutation__round_out[282]) );
  XOR2_X2 _f_permutation__round__U3884  ( .A(_f_permutation__round__N5193 ), 
        .B(_f_permutation__round__c[669] ), .Z(_f_permutation__round_out[283]) );
  XOR2_X2 _f_permutation__round__U3883  ( .A(_f_permutation__round__N5191 ), 
        .B(_f_permutation__round__c[670] ), .Z(_f_permutation__round_out[284]) );
  XOR2_X2 _f_permutation__round__U3882  ( .A(_f_permutation__round__N5189 ), 
        .B(_f_permutation__round__c[671] ), .Z(_f_permutation__round_out[285]) );
  XOR2_X2 _f_permutation__round__U3881  ( .A(_f_permutation__round__N5187 ), 
        .B(_f_permutation__round__c[672] ), .Z(_f_permutation__round_out[286]) );
  XOR2_X2 _f_permutation__round__U3880  ( .A(_f_permutation__round__N5185 ), 
        .B(_f_permutation__round__c[673] ), .Z(_f_permutation__round_out[287]) );
  XOR2_X2 _f_permutation__round__U3879  ( .A(_f_permutation__round__N5183 ), 
        .B(_f_permutation__round__c[674] ), .Z(_f_permutation__round_out[288]) );
  XOR2_X2 _f_permutation__round__U3878  ( .A(_f_permutation__round__N5181 ), 
        .B(_f_permutation__round__c[675] ), .Z(_f_permutation__round_out[289]) );
  XOR2_X2 _f_permutation__round__U3877  ( .A(_f_permutation__round__N5179 ), 
        .B(_f_permutation__round__c[676] ), .Z(_f_permutation__round_out[290]) );
  XOR2_X2 _f_permutation__round__U3876  ( .A(_f_permutation__round__N5177 ), 
        .B(_f_permutation__round__c[677] ), .Z(_f_permutation__round_out[291]) );
  XOR2_X2 _f_permutation__round__U3875  ( .A(_f_permutation__round__N5175 ), 
        .B(_f_permutation__round__c[678] ), .Z(_f_permutation__round_out[292]) );
  XOR2_X2 _f_permutation__round__U3874  ( .A(_f_permutation__round__N5173 ), 
        .B(_f_permutation__round__c[679] ), .Z(_f_permutation__round_out[293]) );
  XOR2_X2 _f_permutation__round__U3873  ( .A(_f_permutation__round__N5171 ), 
        .B(_f_permutation__round__c[680] ), .Z(_f_permutation__round_out[294]) );
  XOR2_X2 _f_permutation__round__U3872  ( .A(_f_permutation__round__N5169 ), 
        .B(_f_permutation__round__c[681] ), .Z(_f_permutation__round_out[295]) );
  XOR2_X2 _f_permutation__round__U3871  ( .A(_f_permutation__round__N5167 ), 
        .B(_f_permutation__round__c[682] ), .Z(_f_permutation__round_out[296]) );
  XOR2_X2 _f_permutation__round__U3870  ( .A(_f_permutation__round__N5165 ), 
        .B(_f_permutation__round__c[683] ), .Z(_f_permutation__round_out[297]) );
  XOR2_X2 _f_permutation__round__U3869  ( .A(_f_permutation__round__N5163 ), 
        .B(_f_permutation__round__c[684] ), .Z(_f_permutation__round_out[298]) );
  XOR2_X2 _f_permutation__round__U3868  ( .A(_f_permutation__round__N5161 ), 
        .B(_f_permutation__round__c[685] ), .Z(_f_permutation__round_out[299]) );
  XOR2_X2 _f_permutation__round__U3867  ( .A(_f_permutation__round__N5159 ), 
        .B(_f_permutation__round__c[686] ), .Z(_f_permutation__round_out[300]) );
  XOR2_X2 _f_permutation__round__U3866  ( .A(_f_permutation__round__N5157 ), 
        .B(_f_permutation__round__c[687] ), .Z(_f_permutation__round_out[301]) );
  XOR2_X2 _f_permutation__round__U3865  ( .A(_f_permutation__round__N5155 ), 
        .B(_f_permutation__round__c[688] ), .Z(_f_permutation__round_out[302]) );
  XOR2_X2 _f_permutation__round__U3864  ( .A(_f_permutation__round__N5153 ), 
        .B(_f_permutation__round__c[689] ), .Z(_f_permutation__round_out[303]) );
  XOR2_X2 _f_permutation__round__U3863  ( .A(_f_permutation__round__N5151 ), 
        .B(_f_permutation__round__c[690] ), .Z(_f_permutation__round_out[304]) );
  XOR2_X2 _f_permutation__round__U3862  ( .A(_f_permutation__round__N5149 ), 
        .B(_f_permutation__round__c[691] ), .Z(_f_permutation__round_out[305]) );
  XOR2_X2 _f_permutation__round__U3861  ( .A(_f_permutation__round__N5147 ), 
        .B(_f_permutation__round__c[692] ), .Z(_f_permutation__round_out[306]) );
  XOR2_X2 _f_permutation__round__U3860  ( .A(_f_permutation__round__N5145 ), 
        .B(_f_permutation__round__c[693] ), .Z(_f_permutation__round_out[307]) );
  XOR2_X2 _f_permutation__round__U3859  ( .A(_f_permutation__round__N5143 ), 
        .B(_f_permutation__round__c[694] ), .Z(_f_permutation__round_out[308]) );
  XOR2_X2 _f_permutation__round__U3858  ( .A(_f_permutation__round__N5141 ), 
        .B(_f_permutation__round__c[695] ), .Z(_f_permutation__round_out[309]) );
  XOR2_X2 _f_permutation__round__U3857  ( .A(_f_permutation__round__N5139 ), 
        .B(_f_permutation__round__c[696] ), .Z(_f_permutation__round_out[310]) );
  XOR2_X2 _f_permutation__round__U3856  ( .A(_f_permutation__round__N5137 ), 
        .B(_f_permutation__round__c[697] ), .Z(_f_permutation__round_out[311]) );
  XOR2_X2 _f_permutation__round__U3855  ( .A(_f_permutation__round__N5135 ), 
        .B(_f_permutation__round__c[698] ), .Z(_f_permutation__round_out[312]) );
  XOR2_X2 _f_permutation__round__U3854  ( .A(_f_permutation__round__N5133 ), 
        .B(_f_permutation__round__c[699] ), .Z(_f_permutation__round_out[313]) );
  XOR2_X2 _f_permutation__round__U3853  ( .A(_f_permutation__round__N5131 ), 
        .B(_f_permutation__round__c[700] ), .Z(_f_permutation__round_out[314]) );
  XOR2_X2 _f_permutation__round__U3852  ( .A(_f_permutation__round__N5129 ), 
        .B(_f_permutation__round__c[701] ), .Z(_f_permutation__round_out[315]) );
  XOR2_X2 _f_permutation__round__U3851  ( .A(_f_permutation__round__N5127 ), 
        .B(_f_permutation__round__c[702] ), .Z(_f_permutation__round_out[316]) );
  XOR2_X2 _f_permutation__round__U3850  ( .A(_f_permutation__round__N5125 ), 
        .B(_f_permutation__round__c[703] ), .Z(_f_permutation__round_out[317]) );
  XOR2_X2 _f_permutation__round__U3849  ( .A(_f_permutation__round__N5123 ), 
        .B(_f_permutation__round__c[640] ), .Z(_f_permutation__round_out[318]) );
  XOR2_X2 _f_permutation__round__U3848  ( .A(_f_permutation__round__N5121 ), 
        .B(_f_permutation__round__c[641] ), .Z(_f_permutation__round_out[319]) );
  XOR2_X2 _f_permutation__round__U3847  ( .A(_f_permutation__round__N5119 ), 
        .B(_f_permutation__round__c[1224] ), .Z(
        _f_permutation__round_out[320]) );
  XOR2_X2 _f_permutation__round__U3846  ( .A(_f_permutation__round__N5117 ), 
        .B(_f_permutation__round__c[1225] ), .Z(
        _f_permutation__round_out[321]) );
  XOR2_X2 _f_permutation__round__U3845  ( .A(_f_permutation__round__N5115 ), 
        .B(_f_permutation__round__c[1226] ), .Z(
        _f_permutation__round_out[322]) );
  XOR2_X2 _f_permutation__round__U3844  ( .A(_f_permutation__round__N5113 ), 
        .B(_f_permutation__round__c[1227] ), .Z(
        _f_permutation__round_out[323]) );
  XOR2_X2 _f_permutation__round__U3843  ( .A(_f_permutation__round__N5111 ), 
        .B(_f_permutation__round__c[1228] ), .Z(
        _f_permutation__round_out[324]) );
  XOR2_X2 _f_permutation__round__U3842  ( .A(_f_permutation__round__N5109 ), 
        .B(_f_permutation__round__c[1229] ), .Z(
        _f_permutation__round_out[325]) );
  XOR2_X2 _f_permutation__round__U3841  ( .A(_f_permutation__round__N5107 ), 
        .B(_f_permutation__round__c[1230] ), .Z(
        _f_permutation__round_out[326]) );
  XOR2_X2 _f_permutation__round__U3840  ( .A(_f_permutation__round__N5105 ), 
        .B(_f_permutation__round__c[1231] ), .Z(
        _f_permutation__round_out[327]) );
  XOR2_X2 _f_permutation__round__U3839  ( .A(_f_permutation__round__N5103 ), 
        .B(_f_permutation__round__c[1232] ), .Z(
        _f_permutation__round_out[328]) );
  XOR2_X2 _f_permutation__round__U3838  ( .A(_f_permutation__round__N5101 ), 
        .B(_f_permutation__round__c[1233] ), .Z(
        _f_permutation__round_out[329]) );
  XOR2_X2 _f_permutation__round__U3837  ( .A(_f_permutation__round__N5099 ), 
        .B(_f_permutation__round__c[1234] ), .Z(
        _f_permutation__round_out[330]) );
  XOR2_X2 _f_permutation__round__U3836  ( .A(_f_permutation__round__N5097 ), 
        .B(_f_permutation__round__c[1235] ), .Z(
        _f_permutation__round_out[331]) );
  XOR2_X2 _f_permutation__round__U3835  ( .A(_f_permutation__round__N5095 ), 
        .B(_f_permutation__round__c[1236] ), .Z(
        _f_permutation__round_out[332]) );
  XOR2_X2 _f_permutation__round__U3834  ( .A(_f_permutation__round__N5093 ), 
        .B(_f_permutation__round__c[1237] ), .Z(
        _f_permutation__round_out[333]) );
  XOR2_X2 _f_permutation__round__U3833  ( .A(_f_permutation__round__N5091 ), 
        .B(_f_permutation__round__c[1238] ), .Z(
        _f_permutation__round_out[334]) );
  XOR2_X2 _f_permutation__round__U3832  ( .A(_f_permutation__round__N5089 ), 
        .B(_f_permutation__round__c[1239] ), .Z(
        _f_permutation__round_out[335]) );
  XOR2_X2 _f_permutation__round__U3831  ( .A(_f_permutation__round__N5087 ), 
        .B(_f_permutation__round__c[1240] ), .Z(
        _f_permutation__round_out[336]) );
  XOR2_X2 _f_permutation__round__U3830  ( .A(_f_permutation__round__N5085 ), 
        .B(_f_permutation__round__c[1241] ), .Z(
        _f_permutation__round_out[337]) );
  XOR2_X2 _f_permutation__round__U3829  ( .A(_f_permutation__round__N5083 ), 
        .B(_f_permutation__round__c[1242] ), .Z(
        _f_permutation__round_out[338]) );
  XOR2_X2 _f_permutation__round__U3828  ( .A(_f_permutation__round__N5081 ), 
        .B(_f_permutation__round__c[1243] ), .Z(
        _f_permutation__round_out[339]) );
  XOR2_X2 _f_permutation__round__U3827  ( .A(_f_permutation__round__N5079 ), 
        .B(_f_permutation__round__c[1244] ), .Z(
        _f_permutation__round_out[340]) );
  XOR2_X2 _f_permutation__round__U3826  ( .A(_f_permutation__round__N5077 ), 
        .B(_f_permutation__round__c[1245] ), .Z(
        _f_permutation__round_out[341]) );
  XOR2_X2 _f_permutation__round__U3825  ( .A(_f_permutation__round__N5075 ), 
        .B(_f_permutation__round__c[1246] ), .Z(
        _f_permutation__round_out[342]) );
  XOR2_X2 _f_permutation__round__U3824  ( .A(_f_permutation__round__N5073 ), 
        .B(_f_permutation__round__c[1247] ), .Z(
        _f_permutation__round_out[343]) );
  XOR2_X2 _f_permutation__round__U3823  ( .A(_f_permutation__round__N5071 ), 
        .B(_f_permutation__round__c[1248] ), .Z(
        _f_permutation__round_out[344]) );
  XOR2_X2 _f_permutation__round__U3822  ( .A(_f_permutation__round__N5069 ), 
        .B(_f_permutation__round__c[1249] ), .Z(
        _f_permutation__round_out[345]) );
  XOR2_X2 _f_permutation__round__U3821  ( .A(_f_permutation__round__N5067 ), 
        .B(_f_permutation__round__c[1250] ), .Z(
        _f_permutation__round_out[346]) );
  XOR2_X2 _f_permutation__round__U3820  ( .A(_f_permutation__round__N5065 ), 
        .B(_f_permutation__round__c[1251] ), .Z(
        _f_permutation__round_out[347]) );
  XOR2_X2 _f_permutation__round__U3819  ( .A(_f_permutation__round__N5063 ), 
        .B(_f_permutation__round__c[1252] ), .Z(
        _f_permutation__round_out[348]) );
  XOR2_X2 _f_permutation__round__U3818  ( .A(_f_permutation__round__N5061 ), 
        .B(_f_permutation__round__c[1253] ), .Z(
        _f_permutation__round_out[349]) );
  XOR2_X2 _f_permutation__round__U3817  ( .A(_f_permutation__round__N5059 ), 
        .B(_f_permutation__round__c[1254] ), .Z(
        _f_permutation__round_out[350]) );
  XOR2_X2 _f_permutation__round__U3816  ( .A(_f_permutation__round__N5057 ), 
        .B(_f_permutation__round__c[1255] ), .Z(
        _f_permutation__round_out[351]) );
  XOR2_X2 _f_permutation__round__U3815  ( .A(_f_permutation__round__N5055 ), 
        .B(_f_permutation__round__c[1256] ), .Z(
        _f_permutation__round_out[352]) );
  XOR2_X2 _f_permutation__round__U3814  ( .A(_f_permutation__round__N5053 ), 
        .B(_f_permutation__round__c[1257] ), .Z(
        _f_permutation__round_out[353]) );
  XOR2_X2 _f_permutation__round__U3813  ( .A(_f_permutation__round__N5051 ), 
        .B(_f_permutation__round__c[1258] ), .Z(
        _f_permutation__round_out[354]) );
  XOR2_X2 _f_permutation__round__U3812  ( .A(_f_permutation__round__N5049 ), 
        .B(_f_permutation__round__c[1259] ), .Z(
        _f_permutation__round_out[355]) );
  XOR2_X2 _f_permutation__round__U3811  ( .A(_f_permutation__round__N5047 ), 
        .B(_f_permutation__round__c[1260] ), .Z(
        _f_permutation__round_out[356]) );
  XOR2_X2 _f_permutation__round__U3810  ( .A(_f_permutation__round__N5045 ), 
        .B(_f_permutation__round__c[1261] ), .Z(
        _f_permutation__round_out[357]) );
  XOR2_X2 _f_permutation__round__U3809  ( .A(_f_permutation__round__N5043 ), 
        .B(_f_permutation__round__c[1262] ), .Z(
        _f_permutation__round_out[358]) );
  XOR2_X2 _f_permutation__round__U3808  ( .A(_f_permutation__round__N5041 ), 
        .B(_f_permutation__round__c[1263] ), .Z(
        _f_permutation__round_out[359]) );
  XOR2_X2 _f_permutation__round__U3807  ( .A(_f_permutation__round__N5039 ), 
        .B(_f_permutation__round__c[1264] ), .Z(
        _f_permutation__round_out[360]) );
  XOR2_X2 _f_permutation__round__U3806  ( .A(_f_permutation__round__N5037 ), 
        .B(_f_permutation__round__c[1265] ), .Z(
        _f_permutation__round_out[361]) );
  XOR2_X2 _f_permutation__round__U3805  ( .A(_f_permutation__round__N5035 ), 
        .B(_f_permutation__round__c[1266] ), .Z(
        _f_permutation__round_out[362]) );
  XOR2_X2 _f_permutation__round__U3804  ( .A(_f_permutation__round__N5033 ), 
        .B(_f_permutation__round__c[1267] ), .Z(
        _f_permutation__round_out[363]) );
  XOR2_X2 _f_permutation__round__U3803  ( .A(_f_permutation__round__N5031 ), 
        .B(_f_permutation__round__c[1268] ), .Z(
        _f_permutation__round_out[364]) );
  XOR2_X2 _f_permutation__round__U3802  ( .A(_f_permutation__round__N5029 ), 
        .B(_f_permutation__round__c[1269] ), .Z(
        _f_permutation__round_out[365]) );
  XOR2_X2 _f_permutation__round__U3801  ( .A(_f_permutation__round__N5027 ), 
        .B(_f_permutation__round__c[1270] ), .Z(
        _f_permutation__round_out[366]) );
  XOR2_X2 _f_permutation__round__U3800  ( .A(_f_permutation__round__N5025 ), 
        .B(_f_permutation__round__c[1271] ), .Z(
        _f_permutation__round_out[367]) );
  XOR2_X2 _f_permutation__round__U3799  ( .A(_f_permutation__round__N5023 ), 
        .B(_f_permutation__round__c[1272] ), .Z(
        _f_permutation__round_out[368]) );
  XOR2_X2 _f_permutation__round__U3798  ( .A(_f_permutation__round__N5021 ), 
        .B(_f_permutation__round__c[1273] ), .Z(
        _f_permutation__round_out[369]) );
  XOR2_X2 _f_permutation__round__U3797  ( .A(_f_permutation__round__N5019 ), 
        .B(_f_permutation__round__c[1274] ), .Z(
        _f_permutation__round_out[370]) );
  XOR2_X2 _f_permutation__round__U3796  ( .A(_f_permutation__round__N5017 ), 
        .B(_f_permutation__round__c[1275] ), .Z(
        _f_permutation__round_out[371]) );
  XOR2_X2 _f_permutation__round__U3795  ( .A(_f_permutation__round__N5015 ), 
        .B(_f_permutation__round__c[1276] ), .Z(
        _f_permutation__round_out[372]) );
  XOR2_X2 _f_permutation__round__U3794  ( .A(_f_permutation__round__N5013 ), 
        .B(_f_permutation__round__c[1277] ), .Z(
        _f_permutation__round_out[373]) );
  XOR2_X2 _f_permutation__round__U3793  ( .A(_f_permutation__round__N5011 ), 
        .B(_f_permutation__round__c[1278] ), .Z(
        _f_permutation__round_out[374]) );
  XOR2_X2 _f_permutation__round__U3792  ( .A(_f_permutation__round__N5009 ), 
        .B(_f_permutation__round__c[1279] ), .Z(
        _f_permutation__round_out[375]) );
  XOR2_X2 _f_permutation__round__U3791  ( .A(_f_permutation__round__N5007 ), 
        .B(_f_permutation__round__c[1216] ), .Z(
        _f_permutation__round_out[376]) );
  XOR2_X2 _f_permutation__round__U3790  ( .A(_f_permutation__round__N5005 ), 
        .B(_f_permutation__round__c[1217] ), .Z(
        _f_permutation__round_out[377]) );
  XOR2_X2 _f_permutation__round__U3789  ( .A(_f_permutation__round__N5003 ), 
        .B(_f_permutation__round__c[1218] ), .Z(
        _f_permutation__round_out[378]) );
  XOR2_X2 _f_permutation__round__U3788  ( .A(_f_permutation__round__N5001 ), 
        .B(_f_permutation__round__c[1219] ), .Z(
        _f_permutation__round_out[379]) );
  XOR2_X2 _f_permutation__round__U3787  ( .A(_f_permutation__round__N4999 ), 
        .B(_f_permutation__round__c[1220] ), .Z(
        _f_permutation__round_out[380]) );
  XOR2_X2 _f_permutation__round__U3786  ( .A(_f_permutation__round__N4997 ), 
        .B(_f_permutation__round__c[1221] ), .Z(
        _f_permutation__round_out[381]) );
  XOR2_X2 _f_permutation__round__U3785  ( .A(_f_permutation__round__N4995 ), 
        .B(_f_permutation__round__c[1222] ), .Z(
        _f_permutation__round_out[382]) );
  XOR2_X2 _f_permutation__round__U3784  ( .A(_f_permutation__round__N4993 ), 
        .B(_f_permutation__round__c[1223] ), .Z(
        _f_permutation__round_out[383]) );
  XOR2_X2 _f_permutation__round__U3783  ( .A(_f_permutation__round__N4991 ), 
        .B(_f_permutation__round__c[881] ), .Z(_f_permutation__round_out[384]) );
  XOR2_X2 _f_permutation__round__U3782  ( .A(_f_permutation__round__N4989 ), 
        .B(_f_permutation__round__c[882] ), .Z(_f_permutation__round_out[385]) );
  XOR2_X2 _f_permutation__round__U3781  ( .A(_f_permutation__round__N4987 ), 
        .B(_f_permutation__round__c[883] ), .Z(_f_permutation__round_out[386]) );
  XOR2_X2 _f_permutation__round__U3780  ( .A(_f_permutation__round__N4985 ), 
        .B(_f_permutation__round__c[884] ), .Z(_f_permutation__round_out[387]) );
  XOR2_X2 _f_permutation__round__U3779  ( .A(_f_permutation__round__N4983 ), 
        .B(_f_permutation__round__c[885] ), .Z(_f_permutation__round_out[388]) );
  XOR2_X2 _f_permutation__round__U3778  ( .A(_f_permutation__round__N4981 ), 
        .B(_f_permutation__round__c[886] ), .Z(_f_permutation__round_out[389]) );
  XOR2_X2 _f_permutation__round__U3777  ( .A(_f_permutation__round__N4979 ), 
        .B(_f_permutation__round__c[887] ), .Z(_f_permutation__round_out[390]) );
  XOR2_X2 _f_permutation__round__U3776  ( .A(_f_permutation__round__N4977 ), 
        .B(_f_permutation__round__c[888] ), .Z(_f_permutation__round_out[391]) );
  XOR2_X2 _f_permutation__round__U3775  ( .A(_f_permutation__round__N4975 ), 
        .B(_f_permutation__round__c[889] ), .Z(_f_permutation__round_out[392]) );
  XOR2_X2 _f_permutation__round__U3774  ( .A(_f_permutation__round__N4973 ), 
        .B(_f_permutation__round__c[890] ), .Z(_f_permutation__round_out[393]) );
  XOR2_X2 _f_permutation__round__U3773  ( .A(_f_permutation__round__N4971 ), 
        .B(_f_permutation__round__c[891] ), .Z(_f_permutation__round_out[394]) );
  XOR2_X2 _f_permutation__round__U3772  ( .A(_f_permutation__round__N4969 ), 
        .B(_f_permutation__round__c[892] ), .Z(_f_permutation__round_out[395]) );
  XOR2_X2 _f_permutation__round__U3771  ( .A(_f_permutation__round__N4967 ), 
        .B(_f_permutation__round__c[893] ), .Z(_f_permutation__round_out[396]) );
  XOR2_X2 _f_permutation__round__U3770  ( .A(_f_permutation__round__N4965 ), 
        .B(_f_permutation__round__c[894] ), .Z(_f_permutation__round_out[397]) );
  XOR2_X2 _f_permutation__round__U3769  ( .A(_f_permutation__round__N4963 ), 
        .B(_f_permutation__round__c[895] ), .Z(_f_permutation__round_out[398]) );
  XOR2_X2 _f_permutation__round__U3768  ( .A(_f_permutation__round__N4961 ), 
        .B(_f_permutation__round__c[832] ), .Z(_f_permutation__round_out[399]) );
  XOR2_X2 _f_permutation__round__U3767  ( .A(_f_permutation__round__N4959 ), 
        .B(_f_permutation__round__c[833] ), .Z(_f_permutation__round_out[400]) );
  XOR2_X2 _f_permutation__round__U3766  ( .A(_f_permutation__round__N4957 ), 
        .B(_f_permutation__round__c[834] ), .Z(_f_permutation__round_out[401]) );
  XOR2_X2 _f_permutation__round__U3765  ( .A(_f_permutation__round__N4955 ), 
        .B(_f_permutation__round__c[835] ), .Z(_f_permutation__round_out[402]) );
  XOR2_X2 _f_permutation__round__U3764  ( .A(_f_permutation__round__N4953 ), 
        .B(_f_permutation__round__c[836] ), .Z(_f_permutation__round_out[403]) );
  XOR2_X2 _f_permutation__round__U3763  ( .A(_f_permutation__round__N4951 ), 
        .B(_f_permutation__round__c[837] ), .Z(_f_permutation__round_out[404]) );
  XOR2_X2 _f_permutation__round__U3762  ( .A(_f_permutation__round__N4949 ), 
        .B(_f_permutation__round__c[838] ), .Z(_f_permutation__round_out[405]) );
  XOR2_X2 _f_permutation__round__U3761  ( .A(_f_permutation__round__N4947 ), 
        .B(_f_permutation__round__c[839] ), .Z(_f_permutation__round_out[406]) );
  XOR2_X2 _f_permutation__round__U3760  ( .A(_f_permutation__round__N4945 ), 
        .B(_f_permutation__round__c[840] ), .Z(_f_permutation__round_out[407]) );
  XOR2_X2 _f_permutation__round__U3759  ( .A(_f_permutation__round__N4943 ), 
        .B(_f_permutation__round__c[841] ), .Z(_f_permutation__round_out[408]) );
  XOR2_X2 _f_permutation__round__U3758  ( .A(_f_permutation__round__N4941 ), 
        .B(_f_permutation__round__c[842] ), .Z(_f_permutation__round_out[409]) );
  XOR2_X2 _f_permutation__round__U3757  ( .A(_f_permutation__round__N4939 ), 
        .B(_f_permutation__round__c[843] ), .Z(_f_permutation__round_out[410]) );
  XOR2_X2 _f_permutation__round__U3756  ( .A(_f_permutation__round__N4937 ), 
        .B(_f_permutation__round__c[844] ), .Z(_f_permutation__round_out[411]) );
  XOR2_X2 _f_permutation__round__U3755  ( .A(_f_permutation__round__N4935 ), 
        .B(_f_permutation__round__c[845] ), .Z(_f_permutation__round_out[412]) );
  XOR2_X2 _f_permutation__round__U3754  ( .A(_f_permutation__round__N4933 ), 
        .B(_f_permutation__round__c[846] ), .Z(_f_permutation__round_out[413]) );
  XOR2_X2 _f_permutation__round__U3753  ( .A(_f_permutation__round__N4931 ), 
        .B(_f_permutation__round__c[847] ), .Z(_f_permutation__round_out[414]) );
  XOR2_X2 _f_permutation__round__U3752  ( .A(_f_permutation__round__N4929 ), 
        .B(_f_permutation__round__c[848] ), .Z(_f_permutation__round_out[415]) );
  XOR2_X2 _f_permutation__round__U3751  ( .A(_f_permutation__round__N4927 ), 
        .B(_f_permutation__round__c[849] ), .Z(_f_permutation__round_out[416]) );
  XOR2_X2 _f_permutation__round__U3750  ( .A(_f_permutation__round__N4925 ), 
        .B(_f_permutation__round__c[850] ), .Z(_f_permutation__round_out[417]) );
  XOR2_X2 _f_permutation__round__U3749  ( .A(_f_permutation__round__N4923 ), 
        .B(_f_permutation__round__c[851] ), .Z(_f_permutation__round_out[418]) );
  XOR2_X2 _f_permutation__round__U3748  ( .A(_f_permutation__round__N4921 ), 
        .B(_f_permutation__round__c[852] ), .Z(_f_permutation__round_out[419]) );
  XOR2_X2 _f_permutation__round__U3747  ( .A(_f_permutation__round__N4919 ), 
        .B(_f_permutation__round__c[853] ), .Z(_f_permutation__round_out[420]) );
  XOR2_X2 _f_permutation__round__U3746  ( .A(_f_permutation__round__N4917 ), 
        .B(_f_permutation__round__c[854] ), .Z(_f_permutation__round_out[421]) );
  XOR2_X2 _f_permutation__round__U3745  ( .A(_f_permutation__round__N4915 ), 
        .B(_f_permutation__round__c[855] ), .Z(_f_permutation__round_out[422]) );
  XOR2_X2 _f_permutation__round__U3744  ( .A(_f_permutation__round__N4913 ), 
        .B(_f_permutation__round__c[856] ), .Z(_f_permutation__round_out[423]) );
  XOR2_X2 _f_permutation__round__U3743  ( .A(_f_permutation__round__N4911 ), 
        .B(_f_permutation__round__c[857] ), .Z(_f_permutation__round_out[424]) );
  XOR2_X2 _f_permutation__round__U3742  ( .A(_f_permutation__round__N4909 ), 
        .B(_f_permutation__round__c[858] ), .Z(_f_permutation__round_out[425]) );
  XOR2_X2 _f_permutation__round__U3741  ( .A(_f_permutation__round__N4907 ), 
        .B(_f_permutation__round__c[859] ), .Z(_f_permutation__round_out[426]) );
  XOR2_X2 _f_permutation__round__U3740  ( .A(_f_permutation__round__N4905 ), 
        .B(_f_permutation__round__c[860] ), .Z(_f_permutation__round_out[427]) );
  XOR2_X2 _f_permutation__round__U3739  ( .A(_f_permutation__round__N4903 ), 
        .B(_f_permutation__round__c[861] ), .Z(_f_permutation__round_out[428]) );
  XOR2_X2 _f_permutation__round__U3738  ( .A(_f_permutation__round__N4901 ), 
        .B(_f_permutation__round__c[862] ), .Z(_f_permutation__round_out[429]) );
  XOR2_X2 _f_permutation__round__U3737  ( .A(_f_permutation__round__N4899 ), 
        .B(_f_permutation__round__c[863] ), .Z(_f_permutation__round_out[430]) );
  XOR2_X2 _f_permutation__round__U3736  ( .A(_f_permutation__round__N4897 ), 
        .B(_f_permutation__round__c[864] ), .Z(_f_permutation__round_out[431]) );
  XOR2_X2 _f_permutation__round__U3735  ( .A(_f_permutation__round__N4895 ), 
        .B(_f_permutation__round__c[865] ), .Z(_f_permutation__round_out[432]) );
  XOR2_X2 _f_permutation__round__U3734  ( .A(_f_permutation__round__N4893 ), 
        .B(_f_permutation__round__c[866] ), .Z(_f_permutation__round_out[433]) );
  XOR2_X2 _f_permutation__round__U3733  ( .A(_f_permutation__round__N4891 ), 
        .B(_f_permutation__round__c[867] ), .Z(_f_permutation__round_out[434]) );
  XOR2_X2 _f_permutation__round__U3732  ( .A(_f_permutation__round__N4889 ), 
        .B(_f_permutation__round__c[868] ), .Z(_f_permutation__round_out[435]) );
  XOR2_X2 _f_permutation__round__U3731  ( .A(_f_permutation__round__N4887 ), 
        .B(_f_permutation__round__c[869] ), .Z(_f_permutation__round_out[436]) );
  XOR2_X2 _f_permutation__round__U3730  ( .A(_f_permutation__round__N4885 ), 
        .B(_f_permutation__round__c[870] ), .Z(_f_permutation__round_out[437]) );
  XOR2_X2 _f_permutation__round__U3729  ( .A(_f_permutation__round__N4883 ), 
        .B(_f_permutation__round__c[871] ), .Z(_f_permutation__round_out[438]) );
  XOR2_X2 _f_permutation__round__U3728  ( .A(_f_permutation__round__N4881 ), 
        .B(_f_permutation__round__c[872] ), .Z(_f_permutation__round_out[439]) );
  XOR2_X2 _f_permutation__round__U3727  ( .A(_f_permutation__round__N4879 ), 
        .B(_f_permutation__round__c[873] ), .Z(_f_permutation__round_out[440]) );
  XOR2_X2 _f_permutation__round__U3726  ( .A(_f_permutation__round__N4877 ), 
        .B(_f_permutation__round__c[874] ), .Z(_f_permutation__round_out[441]) );
  XOR2_X2 _f_permutation__round__U3725  ( .A(_f_permutation__round__N4875 ), 
        .B(_f_permutation__round__c[875] ), .Z(_f_permutation__round_out[442]) );
  XOR2_X2 _f_permutation__round__U3724  ( .A(_f_permutation__round__N4873 ), 
        .B(_f_permutation__round__c[876] ), .Z(_f_permutation__round_out[443]) );
  XOR2_X2 _f_permutation__round__U3723  ( .A(_f_permutation__round__N4871 ), 
        .B(_f_permutation__round__c[877] ), .Z(_f_permutation__round_out[444]) );
  XOR2_X2 _f_permutation__round__U3722  ( .A(_f_permutation__round__N4869 ), 
        .B(_f_permutation__round__c[878] ), .Z(_f_permutation__round_out[445]) );
  XOR2_X2 _f_permutation__round__U3721  ( .A(_f_permutation__round__N4867 ), 
        .B(_f_permutation__round__c[879] ), .Z(_f_permutation__round_out[446]) );
  XOR2_X2 _f_permutation__round__U3720  ( .A(_f_permutation__round__N4865 ), 
        .B(_f_permutation__round__c[880] ), .Z(_f_permutation__round_out[447]) );
  XOR2_X2 _f_permutation__round__U3719  ( .A(_f_permutation__round__N4863 ), 
        .B(_f_permutation__round__c[502] ), .Z(_f_permutation__round_out[448]) );
  XOR2_X2 _f_permutation__round__U3718  ( .A(_f_permutation__round__N4861 ), 
        .B(_f_permutation__round__c[503] ), .Z(_f_permutation__round_out[449]) );
  XOR2_X2 _f_permutation__round__U3717  ( .A(_f_permutation__round__N4859 ), 
        .B(_f_permutation__round__c[504] ), .Z(_f_permutation__round_out[450]) );
  XOR2_X2 _f_permutation__round__U3716  ( .A(_f_permutation__round__N4857 ), 
        .B(_f_permutation__round__c[505] ), .Z(_f_permutation__round_out[451]) );
  XOR2_X2 _f_permutation__round__U3715  ( .A(_f_permutation__round__N4855 ), 
        .B(_f_permutation__round__c[506] ), .Z(_f_permutation__round_out[452]) );
  XOR2_X2 _f_permutation__round__U3714  ( .A(_f_permutation__round__N4853 ), 
        .B(_f_permutation__round__c[507] ), .Z(_f_permutation__round_out[453]) );
  XOR2_X2 _f_permutation__round__U3713  ( .A(_f_permutation__round__N4851 ), 
        .B(_f_permutation__round__c[508] ), .Z(_f_permutation__round_out[454]) );
  XOR2_X2 _f_permutation__round__U3712  ( .A(_f_permutation__round__N4849 ), 
        .B(_f_permutation__round__c[509] ), .Z(_f_permutation__round_out[455]) );
  XOR2_X2 _f_permutation__round__U3711  ( .A(_f_permutation__round__N4847 ), 
        .B(_f_permutation__round__c[510] ), .Z(_f_permutation__round_out[456]) );
  XOR2_X2 _f_permutation__round__U3710  ( .A(_f_permutation__round__N4845 ), 
        .B(_f_permutation__round__c[511] ), .Z(_f_permutation__round_out[457]) );
  XOR2_X2 _f_permutation__round__U3709  ( .A(_f_permutation__round__N4843 ), 
        .B(_f_permutation__round__c[448] ), .Z(_f_permutation__round_out[458]) );
  XOR2_X2 _f_permutation__round__U3708  ( .A(_f_permutation__round__N4841 ), 
        .B(_f_permutation__round__c[449] ), .Z(_f_permutation__round_out[459]) );
  XOR2_X2 _f_permutation__round__U3707  ( .A(_f_permutation__round__N4839 ), 
        .B(_f_permutation__round__c[450] ), .Z(_f_permutation__round_out[460]) );
  XOR2_X2 _f_permutation__round__U3706  ( .A(_f_permutation__round__N4837 ), 
        .B(_f_permutation__round__c[451] ), .Z(_f_permutation__round_out[461]) );
  XOR2_X2 _f_permutation__round__U3705  ( .A(_f_permutation__round__N4835 ), 
        .B(_f_permutation__round__c[452] ), .Z(_f_permutation__round_out[462]) );
  XOR2_X2 _f_permutation__round__U3704  ( .A(_f_permutation__round__N4833 ), 
        .B(_f_permutation__round__c[453] ), .Z(_f_permutation__round_out[463]) );
  XOR2_X2 _f_permutation__round__U3703  ( .A(_f_permutation__round__N4831 ), 
        .B(_f_permutation__round__c[454] ), .Z(_f_permutation__round_out[464]) );
  XOR2_X2 _f_permutation__round__U3702  ( .A(_f_permutation__round__N4829 ), 
        .B(_f_permutation__round__c[455] ), .Z(_f_permutation__round_out[465]) );
  XOR2_X2 _f_permutation__round__U3701  ( .A(_f_permutation__round__N4827 ), 
        .B(_f_permutation__round__c[456] ), .Z(_f_permutation__round_out[466]) );
  XOR2_X2 _f_permutation__round__U3700  ( .A(_f_permutation__round__N4825 ), 
        .B(_f_permutation__round__c[457] ), .Z(_f_permutation__round_out[467]) );
  XOR2_X2 _f_permutation__round__U3699  ( .A(_f_permutation__round__N4823 ), 
        .B(_f_permutation__round__c[458] ), .Z(_f_permutation__round_out[468]) );
  XOR2_X2 _f_permutation__round__U3698  ( .A(_f_permutation__round__N4821 ), 
        .B(_f_permutation__round__c[459] ), .Z(_f_permutation__round_out[469]) );
  XOR2_X2 _f_permutation__round__U3697  ( .A(_f_permutation__round__N4819 ), 
        .B(_f_permutation__round__c[460] ), .Z(_f_permutation__round_out[470]) );
  XOR2_X2 _f_permutation__round__U3696  ( .A(_f_permutation__round__N4817 ), 
        .B(_f_permutation__round__c[461] ), .Z(_f_permutation__round_out[471]) );
  XOR2_X2 _f_permutation__round__U3695  ( .A(_f_permutation__round__N4815 ), 
        .B(_f_permutation__round__c[462] ), .Z(_f_permutation__round_out[472]) );
  XOR2_X2 _f_permutation__round__U3694  ( .A(_f_permutation__round__N4813 ), 
        .B(_f_permutation__round__c[463] ), .Z(_f_permutation__round_out[473]) );
  XOR2_X2 _f_permutation__round__U3693  ( .A(_f_permutation__round__N4811 ), 
        .B(_f_permutation__round__c[464] ), .Z(_f_permutation__round_out[474]) );
  XOR2_X2 _f_permutation__round__U3692  ( .A(_f_permutation__round__N4809 ), 
        .B(_f_permutation__round__c[465] ), .Z(_f_permutation__round_out[475]) );
  XOR2_X2 _f_permutation__round__U3691  ( .A(_f_permutation__round__N4807 ), 
        .B(_f_permutation__round__c[466] ), .Z(_f_permutation__round_out[476]) );
  XOR2_X2 _f_permutation__round__U3690  ( .A(_f_permutation__round__N4805 ), 
        .B(_f_permutation__round__c[467] ), .Z(_f_permutation__round_out[477]) );
  XOR2_X2 _f_permutation__round__U3689  ( .A(_f_permutation__round__N4803 ), 
        .B(_f_permutation__round__c[468] ), .Z(_f_permutation__round_out[478]) );
  XOR2_X2 _f_permutation__round__U3688  ( .A(_f_permutation__round__N4801 ), 
        .B(_f_permutation__round__c[469] ), .Z(_f_permutation__round_out[479]) );
  XOR2_X2 _f_permutation__round__U3687  ( .A(_f_permutation__round__N4799 ), 
        .B(_f_permutation__round__c[470] ), .Z(_f_permutation__round_out[480]) );
  XOR2_X2 _f_permutation__round__U3686  ( .A(_f_permutation__round__N4797 ), 
        .B(_f_permutation__round__c[471] ), .Z(_f_permutation__round_out[481]) );
  XOR2_X2 _f_permutation__round__U3685  ( .A(_f_permutation__round__N4795 ), 
        .B(_f_permutation__round__c[472] ), .Z(_f_permutation__round_out[482]) );
  XOR2_X2 _f_permutation__round__U3684  ( .A(_f_permutation__round__N4793 ), 
        .B(_f_permutation__round__c[473] ), .Z(_f_permutation__round_out[483]) );
  XOR2_X2 _f_permutation__round__U3683  ( .A(_f_permutation__round__N4791 ), 
        .B(_f_permutation__round__c[474] ), .Z(_f_permutation__round_out[484]) );
  XOR2_X2 _f_permutation__round__U3682  ( .A(_f_permutation__round__N4789 ), 
        .B(_f_permutation__round__c[475] ), .Z(_f_permutation__round_out[485]) );
  XOR2_X2 _f_permutation__round__U3681  ( .A(_f_permutation__round__N4787 ), 
        .B(_f_permutation__round__c[476] ), .Z(_f_permutation__round_out[486]) );
  XOR2_X2 _f_permutation__round__U3680  ( .A(_f_permutation__round__N4785 ), 
        .B(_f_permutation__round__c[477] ), .Z(_f_permutation__round_out[487]) );
  XOR2_X2 _f_permutation__round__U3679  ( .A(_f_permutation__round__N4783 ), 
        .B(_f_permutation__round__c[478] ), .Z(_f_permutation__round_out[488]) );
  XOR2_X2 _f_permutation__round__U3678  ( .A(_f_permutation__round__N4781 ), 
        .B(_f_permutation__round__c[479] ), .Z(_f_permutation__round_out[489]) );
  XOR2_X2 _f_permutation__round__U3677  ( .A(_f_permutation__round__N4779 ), 
        .B(_f_permutation__round__c[480] ), .Z(_f_permutation__round_out[490]) );
  XOR2_X2 _f_permutation__round__U3676  ( .A(_f_permutation__round__N4777 ), 
        .B(_f_permutation__round__c[481] ), .Z(_f_permutation__round_out[491]) );
  XOR2_X2 _f_permutation__round__U3675  ( .A(_f_permutation__round__N4775 ), 
        .B(_f_permutation__round__c[482] ), .Z(_f_permutation__round_out[492]) );
  XOR2_X2 _f_permutation__round__U3674  ( .A(_f_permutation__round__N4773 ), 
        .B(_f_permutation__round__c[483] ), .Z(_f_permutation__round_out[493]) );
  XOR2_X2 _f_permutation__round__U3673  ( .A(_f_permutation__round__N4771 ), 
        .B(_f_permutation__round__c[484] ), .Z(_f_permutation__round_out[494]) );
  XOR2_X2 _f_permutation__round__U3672  ( .A(_f_permutation__round__N4769 ), 
        .B(_f_permutation__round__c[485] ), .Z(_f_permutation__round_out[495]) );
  XOR2_X2 _f_permutation__round__U3671  ( .A(_f_permutation__round__N4767 ), 
        .B(_f_permutation__round__c[486] ), .Z(_f_permutation__round_out[496]) );
  XOR2_X2 _f_permutation__round__U3670  ( .A(_f_permutation__round__N4765 ), 
        .B(_f_permutation__round__c[487] ), .Z(_f_permutation__round_out[497]) );
  XOR2_X2 _f_permutation__round__U3669  ( .A(_f_permutation__round__N4763 ), 
        .B(_f_permutation__round__c[488] ), .Z(_f_permutation__round_out[498]) );
  XOR2_X2 _f_permutation__round__U3668  ( .A(_f_permutation__round__N4761 ), 
        .B(_f_permutation__round__c[489] ), .Z(_f_permutation__round_out[499]) );
  XOR2_X2 _f_permutation__round__U3667  ( .A(_f_permutation__round__N4759 ), 
        .B(_f_permutation__round__c[490] ), .Z(_f_permutation__round_out[500]) );
  XOR2_X2 _f_permutation__round__U3666  ( .A(_f_permutation__round__N4757 ), 
        .B(_f_permutation__round__c[491] ), .Z(_f_permutation__round_out[501]) );
  XOR2_X2 _f_permutation__round__U3665  ( .A(_f_permutation__round__N4755 ), 
        .B(_f_permutation__round__c[492] ), .Z(_f_permutation__round_out[502]) );
  XOR2_X2 _f_permutation__round__U3664  ( .A(_f_permutation__round__N4753 ), 
        .B(_f_permutation__round__c[493] ), .Z(_f_permutation__round_out[503]) );
  XOR2_X2 _f_permutation__round__U3663  ( .A(_f_permutation__round__N4751 ), 
        .B(_f_permutation__round__c[494] ), .Z(_f_permutation__round_out[504]) );
  XOR2_X2 _f_permutation__round__U3662  ( .A(_f_permutation__round__N4749 ), 
        .B(_f_permutation__round__c[495] ), .Z(_f_permutation__round_out[505]) );
  XOR2_X2 _f_permutation__round__U3661  ( .A(_f_permutation__round__N4747 ), 
        .B(_f_permutation__round__c[496] ), .Z(_f_permutation__round_out[506]) );
  XOR2_X2 _f_permutation__round__U3660  ( .A(_f_permutation__round__N4745 ), 
        .B(_f_permutation__round__c[497] ), .Z(_f_permutation__round_out[507]) );
  XOR2_X2 _f_permutation__round__U3659  ( .A(_f_permutation__round__N4743 ), 
        .B(_f_permutation__round__c[498] ), .Z(_f_permutation__round_out[508]) );
  XOR2_X2 _f_permutation__round__U3658  ( .A(_f_permutation__round__N4741 ), 
        .B(_f_permutation__round__c[499] ), .Z(_f_permutation__round_out[509]) );
  XOR2_X2 _f_permutation__round__U3657  ( .A(_f_permutation__round__N4739 ), 
        .B(_f_permutation__round__c[500] ), .Z(_f_permutation__round_out[510]) );
  XOR2_X2 _f_permutation__round__U3656  ( .A(_f_permutation__round__N4737 ), 
        .B(_f_permutation__round__c[501] ), .Z(_f_permutation__round_out[511]) );
  XOR2_X2 _f_permutation__round__U3655  ( .A(_f_permutation__round__N4735 ), 
        .B(_f_permutation__round__c[92] ), .Z(_f_permutation__round_out[512])
         );
  XOR2_X2 _f_permutation__round__U3654  ( .A(_f_permutation__round__N4733 ), 
        .B(_f_permutation__round__c[93] ), .Z(_f_permutation__round_out[513])
         );
  XOR2_X2 _f_permutation__round__U3653  ( .A(_f_permutation__round__N4731 ), 
        .B(_f_permutation__round__c[94] ), .Z(_f_permutation__round_out[514])
         );
  XOR2_X2 _f_permutation__round__U3652  ( .A(_f_permutation__round__N4729 ), 
        .B(_f_permutation__round__c[95] ), .Z(_f_permutation__round_out[515])
         );
  XOR2_X2 _f_permutation__round__U3651  ( .A(_f_permutation__round__N4727 ), 
        .B(_f_permutation__round__c[96] ), .Z(_f_permutation__round_out[516])
         );
  XOR2_X2 _f_permutation__round__U3650  ( .A(_f_permutation__round__N4725 ), 
        .B(_f_permutation__round__c[97] ), .Z(_f_permutation__round_out[517])
         );
  XOR2_X2 _f_permutation__round__U3649  ( .A(_f_permutation__round__N4723 ), 
        .B(_f_permutation__round__c[98] ), .Z(_f_permutation__round_out[518])
         );
  XOR2_X2 _f_permutation__round__U3648  ( .A(_f_permutation__round__N4721 ), 
        .B(_f_permutation__round__c[99] ), .Z(_f_permutation__round_out[519])
         );
  XOR2_X2 _f_permutation__round__U3647  ( .A(_f_permutation__round__N4719 ), 
        .B(_f_permutation__round__c[100] ), .Z(_f_permutation__round_out[520]) );
  XOR2_X2 _f_permutation__round__U3646  ( .A(_f_permutation__round__N4717 ), 
        .B(_f_permutation__round__c[101] ), .Z(_f_permutation__round_out[521]) );
  XOR2_X2 _f_permutation__round__U3645  ( .A(_f_permutation__round__N4715 ), 
        .B(_f_permutation__round__c[102] ), .Z(_f_permutation__round_out[522]) );
  XOR2_X2 _f_permutation__round__U3644  ( .A(_f_permutation__round__N4713 ), 
        .B(_f_permutation__round__c[103] ), .Z(_f_permutation__round_out[523]) );
  XOR2_X2 _f_permutation__round__U3643  ( .A(_f_permutation__round__N4711 ), 
        .B(_f_permutation__round__c[104] ), .Z(_f_permutation__round_out[524]) );
  XOR2_X2 _f_permutation__round__U3642  ( .A(_f_permutation__round__N4709 ), 
        .B(_f_permutation__round__c[105] ), .Z(_f_permutation__round_out[525]) );
  XOR2_X2 _f_permutation__round__U3641  ( .A(_f_permutation__round__N4707 ), 
        .B(_f_permutation__round__c[106] ), .Z(_f_permutation__round_out[526]) );
  XOR2_X2 _f_permutation__round__U3640  ( .A(_f_permutation__round__N4705 ), 
        .B(_f_permutation__round__c[107] ), .Z(_f_permutation__round_out[527]) );
  XOR2_X2 _f_permutation__round__U3639  ( .A(_f_permutation__round__N4703 ), 
        .B(_f_permutation__round__c[108] ), .Z(_f_permutation__round_out[528]) );
  XOR2_X2 _f_permutation__round__U3638  ( .A(_f_permutation__round__N4701 ), 
        .B(_f_permutation__round__c[109] ), .Z(_f_permutation__round_out[529]) );
  XOR2_X2 _f_permutation__round__U3637  ( .A(_f_permutation__round__N4699 ), 
        .B(_f_permutation__round__c[110] ), .Z(_f_permutation__round_out[530]) );
  XOR2_X2 _f_permutation__round__U3636  ( .A(_f_permutation__round__N4697 ), 
        .B(_f_permutation__round__c[111] ), .Z(_f_permutation__round_out[531]) );
  XOR2_X2 _f_permutation__round__U3635  ( .A(_f_permutation__round__N4695 ), 
        .B(_f_permutation__round__c[112] ), .Z(_f_permutation__round_out[532]) );
  XOR2_X2 _f_permutation__round__U3634  ( .A(_f_permutation__round__N4693 ), 
        .B(_f_permutation__round__c[113] ), .Z(_f_permutation__round_out[533]) );
  XOR2_X2 _f_permutation__round__U3633  ( .A(_f_permutation__round__N4691 ), 
        .B(_f_permutation__round__c[114] ), .Z(_f_permutation__round_out[534]) );
  XOR2_X2 _f_permutation__round__U3632  ( .A(_f_permutation__round__N4689 ), 
        .B(_f_permutation__round__c[115] ), .Z(_f_permutation__round_out[535]) );
  XOR2_X2 _f_permutation__round__U3631  ( .A(_f_permutation__round__N4687 ), 
        .B(_f_permutation__round__c[116] ), .Z(_f_permutation__round_out[536]) );
  XOR2_X2 _f_permutation__round__U3630  ( .A(_f_permutation__round__N4685 ), 
        .B(_f_permutation__round__c[117] ), .Z(_f_permutation__round_out[537]) );
  XOR2_X2 _f_permutation__round__U3629  ( .A(_f_permutation__round__N4683 ), 
        .B(_f_permutation__round__c[118] ), .Z(_f_permutation__round_out[538]) );
  XOR2_X2 _f_permutation__round__U3628  ( .A(_f_permutation__round__N4681 ), 
        .B(_f_permutation__round__c[119] ), .Z(_f_permutation__round_out[539]) );
  XOR2_X2 _f_permutation__round__U3627  ( .A(_f_permutation__round__N4679 ), 
        .B(_f_permutation__round__c[120] ), .Z(_f_permutation__round_out[540]) );
  XOR2_X2 _f_permutation__round__U3626  ( .A(_f_permutation__round__N4677 ), 
        .B(_f_permutation__round__c[121] ), .Z(_f_permutation__round_out[541]) );
  XOR2_X2 _f_permutation__round__U3625  ( .A(_f_permutation__round__N4675 ), 
        .B(_f_permutation__round__c[122] ), .Z(_f_permutation__round_out[542]) );
  XOR2_X2 _f_permutation__round__U3624  ( .A(_f_permutation__round__N4673 ), 
        .B(_f_permutation__round__c[123] ), .Z(_f_permutation__round_out[543]) );
  XOR2_X2 _f_permutation__round__U3623  ( .A(_f_permutation__round__N4671 ), 
        .B(_f_permutation__round__c[124] ), .Z(_f_permutation__round_out[544]) );
  XOR2_X2 _f_permutation__round__U3622  ( .A(_f_permutation__round__N4669 ), 
        .B(_f_permutation__round__c[125] ), .Z(_f_permutation__round_out[545]) );
  XOR2_X2 _f_permutation__round__U3621  ( .A(_f_permutation__round__N4667 ), 
        .B(_f_permutation__round__c[126] ), .Z(_f_permutation__round_out[546]) );
  XOR2_X2 _f_permutation__round__U3620  ( .A(_f_permutation__round__N4665 ), 
        .B(_f_permutation__round__c[127] ), .Z(_f_permutation__round_out[547]) );
  XOR2_X2 _f_permutation__round__U3619  ( .A(_f_permutation__round__N4663 ), 
        .B(_f_permutation__round__c[64] ), .Z(_f_permutation__round_out[548])
         );
  XOR2_X2 _f_permutation__round__U3618  ( .A(_f_permutation__round__N4661 ), 
        .B(_f_permutation__round__c[65] ), .Z(_f_permutation__round_out[549])
         );
  XOR2_X2 _f_permutation__round__U3617  ( .A(_f_permutation__round__N4659 ), 
        .B(_f_permutation__round__c[66] ), .Z(_f_permutation__round_out[550])
         );
  XOR2_X2 _f_permutation__round__U3616  ( .A(_f_permutation__round__N4657 ), 
        .B(_f_permutation__round__c[67] ), .Z(_f_permutation__round_out[551])
         );
  XOR2_X2 _f_permutation__round__U3615  ( .A(_f_permutation__round__N4655 ), 
        .B(_f_permutation__round__c[68] ), .Z(_f_permutation__round_out[552])
         );
  XOR2_X2 _f_permutation__round__U3614  ( .A(_f_permutation__round__N4653 ), 
        .B(_f_permutation__round__c[69] ), .Z(_f_permutation__round_out[553])
         );
  XOR2_X2 _f_permutation__round__U3613  ( .A(_f_permutation__round__N4651 ), 
        .B(_f_permutation__round__c[70] ), .Z(_f_permutation__round_out[554])
         );
  XOR2_X2 _f_permutation__round__U3612  ( .A(_f_permutation__round__N4649 ), 
        .B(_f_permutation__round__c[71] ), .Z(_f_permutation__round_out[555])
         );
  XOR2_X2 _f_permutation__round__U3611  ( .A(_f_permutation__round__N4647 ), 
        .B(_f_permutation__round__c[72] ), .Z(_f_permutation__round_out[556])
         );
  XOR2_X2 _f_permutation__round__U3610  ( .A(_f_permutation__round__N4645 ), 
        .B(_f_permutation__round__c[73] ), .Z(_f_permutation__round_out[557])
         );
  XOR2_X2 _f_permutation__round__U3609  ( .A(_f_permutation__round__N4643 ), 
        .B(_f_permutation__round__c[74] ), .Z(_f_permutation__round_out[558])
         );
  XOR2_X2 _f_permutation__round__U3608  ( .A(_f_permutation__round__N4641 ), 
        .B(_f_permutation__round__c[75] ), .Z(_f_permutation__round_out[559])
         );
  XOR2_X2 _f_permutation__round__U3607  ( .A(_f_permutation__round__N4639 ), 
        .B(_f_permutation__round__c[76] ), .Z(_f_permutation__round_out[560])
         );
  XOR2_X2 _f_permutation__round__U3606  ( .A(_f_permutation__round__N4637 ), 
        .B(_f_permutation__round__c[77] ), .Z(_f_permutation__round_out[561])
         );
  XOR2_X2 _f_permutation__round__U3605  ( .A(_f_permutation__round__N4635 ), 
        .B(_f_permutation__round__c[78] ), .Z(_f_permutation__round_out[562])
         );
  XOR2_X2 _f_permutation__round__U3604  ( .A(_f_permutation__round__N4633 ), 
        .B(_f_permutation__round__c[79] ), .Z(_f_permutation__round_out[563])
         );
  XOR2_X2 _f_permutation__round__U3603  ( .A(_f_permutation__round__N4631 ), 
        .B(_f_permutation__round__c[80] ), .Z(_f_permutation__round_out[564])
         );
  XOR2_X2 _f_permutation__round__U3602  ( .A(_f_permutation__round__N4629 ), 
        .B(_f_permutation__round__c[81] ), .Z(_f_permutation__round_out[565])
         );
  XOR2_X2 _f_permutation__round__U3601  ( .A(_f_permutation__round__N4627 ), 
        .B(_f_permutation__round__c[82] ), .Z(_f_permutation__round_out[566])
         );
  XOR2_X2 _f_permutation__round__U3600  ( .A(_f_permutation__round__N4625 ), 
        .B(_f_permutation__round__c[83] ), .Z(_f_permutation__round_out[567])
         );
  XOR2_X2 _f_permutation__round__U3599  ( .A(_f_permutation__round__N4623 ), 
        .B(_f_permutation__round__c[84] ), .Z(_f_permutation__round_out[568])
         );
  XOR2_X2 _f_permutation__round__U3598  ( .A(_f_permutation__round__N4621 ), 
        .B(_f_permutation__round__c[85] ), .Z(_f_permutation__round_out[569])
         );
  XOR2_X2 _f_permutation__round__U3597  ( .A(_f_permutation__round__N4619 ), 
        .B(_f_permutation__round__c[86] ), .Z(_f_permutation__round_out[570])
         );
  XOR2_X2 _f_permutation__round__U3596  ( .A(_f_permutation__round__N4617 ), 
        .B(_f_permutation__round__c[87] ), .Z(_f_permutation__round_out[571])
         );
  XOR2_X2 _f_permutation__round__U3595  ( .A(_f_permutation__round__N4615 ), 
        .B(_f_permutation__round__c[88] ), .Z(_f_permutation__round_out[572])
         );
  XOR2_X2 _f_permutation__round__U3594  ( .A(_f_permutation__round__N4613 ), 
        .B(_f_permutation__round__c[89] ), .Z(_f_permutation__round_out[573])
         );
  XOR2_X2 _f_permutation__round__U3593  ( .A(_f_permutation__round__N4611 ), 
        .B(_f_permutation__round__c[90] ), .Z(_f_permutation__round_out[574])
         );
  XOR2_X2 _f_permutation__round__U3592  ( .A(_f_permutation__round__N4609 ), 
        .B(_f_permutation__round__c[91] ), .Z(_f_permutation__round_out[575])
         );
  XOR2_X2 _f_permutation__round__U3591  ( .A(_f_permutation__round__N4607 ), 
        .B(_f_permutation__round__c[1317] ), .Z(
        _f_permutation__round_out[576]) );
  XOR2_X2 _f_permutation__round__U3590  ( .A(_f_permutation__round__N4605 ), 
        .B(_f_permutation__round__c[1318] ), .Z(
        _f_permutation__round_out[577]) );
  XOR2_X2 _f_permutation__round__U3589  ( .A(_f_permutation__round__N4603 ), 
        .B(_f_permutation__round__c[1319] ), .Z(
        _f_permutation__round_out[578]) );
  XOR2_X2 _f_permutation__round__U3588  ( .A(_f_permutation__round__N4601 ), 
        .B(_f_permutation__round__c[1320] ), .Z(
        _f_permutation__round_out[579]) );
  XOR2_X2 _f_permutation__round__U3587  ( .A(_f_permutation__round__N4599 ), 
        .B(_f_permutation__round__c[1321] ), .Z(
        _f_permutation__round_out[580]) );
  XOR2_X2 _f_permutation__round__U3586  ( .A(_f_permutation__round__N4597 ), 
        .B(_f_permutation__round__c[1322] ), .Z(
        _f_permutation__round_out[581]) );
  XOR2_X2 _f_permutation__round__U3585  ( .A(_f_permutation__round__N4595 ), 
        .B(_f_permutation__round__c[1323] ), .Z(
        _f_permutation__round_out[582]) );
  XOR2_X2 _f_permutation__round__U3584  ( .A(_f_permutation__round__N4593 ), 
        .B(_f_permutation__round__c[1324] ), .Z(
        _f_permutation__round_out[583]) );
  XOR2_X2 _f_permutation__round__U3583  ( .A(_f_permutation__round__N4591 ), 
        .B(_f_permutation__round__c[1325] ), .Z(
        _f_permutation__round_out[584]) );
  XOR2_X2 _f_permutation__round__U3582  ( .A(_f_permutation__round__N4589 ), 
        .B(_f_permutation__round__c[1326] ), .Z(
        _f_permutation__round_out[585]) );
  XOR2_X2 _f_permutation__round__U3581  ( .A(_f_permutation__round__N4587 ), 
        .B(_f_permutation__round__c[1327] ), .Z(
        _f_permutation__round_out[586]) );
  XOR2_X2 _f_permutation__round__U3580  ( .A(_f_permutation__round__N4585 ), 
        .B(_f_permutation__round__c[1328] ), .Z(
        _f_permutation__round_out[587]) );
  XOR2_X2 _f_permutation__round__U3579  ( .A(_f_permutation__round__N4583 ), 
        .B(_f_permutation__round__c[1329] ), .Z(
        _f_permutation__round_out[588]) );
  XOR2_X2 _f_permutation__round__U3578  ( .A(_f_permutation__round__N4581 ), 
        .B(_f_permutation__round__c[1330] ), .Z(
        _f_permutation__round_out[589]) );
  XOR2_X2 _f_permutation__round__U3577  ( .A(_f_permutation__round__N4579 ), 
        .B(_f_permutation__round__c[1331] ), .Z(
        _f_permutation__round_out[590]) );
  XOR2_X2 _f_permutation__round__U3576  ( .A(_f_permutation__round__N4577 ), 
        .B(_f_permutation__round__c[1332] ), .Z(
        _f_permutation__round_out[591]) );
  XOR2_X2 _f_permutation__round__U3575  ( .A(_f_permutation__round__N4575 ), 
        .B(_f_permutation__round__c[1333] ), .Z(
        _f_permutation__round_out[592]) );
  XOR2_X2 _f_permutation__round__U3574  ( .A(_f_permutation__round__N4573 ), 
        .B(_f_permutation__round__c[1334] ), .Z(
        _f_permutation__round_out[593]) );
  XOR2_X2 _f_permutation__round__U3573  ( .A(_f_permutation__round__N4571 ), 
        .B(_f_permutation__round__c[1335] ), .Z(
        _f_permutation__round_out[594]) );
  XOR2_X2 _f_permutation__round__U3572  ( .A(_f_permutation__round__N4569 ), 
        .B(_f_permutation__round__c[1336] ), .Z(
        _f_permutation__round_out[595]) );
  XOR2_X2 _f_permutation__round__U3571  ( .A(_f_permutation__round__N4567 ), 
        .B(_f_permutation__round__c[1337] ), .Z(
        _f_permutation__round_out[596]) );
  XOR2_X2 _f_permutation__round__U3570  ( .A(_f_permutation__round__N4565 ), 
        .B(_f_permutation__round__c[1338] ), .Z(
        _f_permutation__round_out[597]) );
  XOR2_X2 _f_permutation__round__U3569  ( .A(_f_permutation__round__N4563 ), 
        .B(_f_permutation__round__c[1339] ), .Z(
        _f_permutation__round_out[598]) );
  XOR2_X2 _f_permutation__round__U3568  ( .A(_f_permutation__round__N4561 ), 
        .B(_f_permutation__round__c[1340] ), .Z(
        _f_permutation__round_out[599]) );
  XOR2_X2 _f_permutation__round__U3567  ( .A(_f_permutation__round__N4559 ), 
        .B(_f_permutation__round__c[1341] ), .Z(
        _f_permutation__round_out[600]) );
  XOR2_X2 _f_permutation__round__U3566  ( .A(_f_permutation__round__N4557 ), 
        .B(_f_permutation__round__c[1342] ), .Z(
        _f_permutation__round_out[601]) );
  XOR2_X2 _f_permutation__round__U3565  ( .A(_f_permutation__round__N4555 ), 
        .B(_f_permutation__round__c[1343] ), .Z(
        _f_permutation__round_out[602]) );
  XOR2_X2 _f_permutation__round__U3564  ( .A(_f_permutation__round__N4553 ), 
        .B(_f_permutation__round__c[1280] ), .Z(
        _f_permutation__round_out[603]) );
  XOR2_X2 _f_permutation__round__U3563  ( .A(_f_permutation__round__N4551 ), 
        .B(_f_permutation__round__c[1281] ), .Z(
        _f_permutation__round_out[604]) );
  XOR2_X2 _f_permutation__round__U3562  ( .A(_f_permutation__round__N4549 ), 
        .B(_f_permutation__round__c[1282] ), .Z(
        _f_permutation__round_out[605]) );
  XOR2_X2 _f_permutation__round__U3561  ( .A(_f_permutation__round__N4547 ), 
        .B(_f_permutation__round__c[1283] ), .Z(
        _f_permutation__round_out[606]) );
  XOR2_X2 _f_permutation__round__U3560  ( .A(_f_permutation__round__N4545 ), 
        .B(_f_permutation__round__c[1284] ), .Z(
        _f_permutation__round_out[607]) );
  XOR2_X2 _f_permutation__round__U3559  ( .A(_f_permutation__round__N4543 ), 
        .B(_f_permutation__round__c[1285] ), .Z(
        _f_permutation__round_out[608]) );
  XOR2_X2 _f_permutation__round__U3558  ( .A(_f_permutation__round__N4541 ), 
        .B(_f_permutation__round__c[1286] ), .Z(
        _f_permutation__round_out[609]) );
  XOR2_X2 _f_permutation__round__U3557  ( .A(_f_permutation__round__N4539 ), 
        .B(_f_permutation__round__c[1287] ), .Z(
        _f_permutation__round_out[610]) );
  XOR2_X2 _f_permutation__round__U3556  ( .A(_f_permutation__round__N4537 ), 
        .B(_f_permutation__round__c[1288] ), .Z(
        _f_permutation__round_out[611]) );
  XOR2_X2 _f_permutation__round__U3555  ( .A(_f_permutation__round__N4535 ), 
        .B(_f_permutation__round__c[1289] ), .Z(
        _f_permutation__round_out[612]) );
  XOR2_X2 _f_permutation__round__U3554  ( .A(_f_permutation__round__N4533 ), 
        .B(_f_permutation__round__c[1290] ), .Z(
        _f_permutation__round_out[613]) );
  XOR2_X2 _f_permutation__round__U3553  ( .A(_f_permutation__round__N4531 ), 
        .B(_f_permutation__round__c[1291] ), .Z(
        _f_permutation__round_out[614]) );
  XOR2_X2 _f_permutation__round__U3552  ( .A(_f_permutation__round__N4529 ), 
        .B(_f_permutation__round__c[1292] ), .Z(
        _f_permutation__round_out[615]) );
  XOR2_X2 _f_permutation__round__U3551  ( .A(_f_permutation__round__N4527 ), 
        .B(_f_permutation__round__c[1293] ), .Z(
        _f_permutation__round_out[616]) );
  XOR2_X2 _f_permutation__round__U3550  ( .A(_f_permutation__round__N4525 ), 
        .B(_f_permutation__round__c[1294] ), .Z(
        _f_permutation__round_out[617]) );
  XOR2_X2 _f_permutation__round__U3549  ( .A(_f_permutation__round__N4523 ), 
        .B(_f_permutation__round__c[1295] ), .Z(
        _f_permutation__round_out[618]) );
  XOR2_X2 _f_permutation__round__U3548  ( .A(_f_permutation__round__N4521 ), 
        .B(_f_permutation__round__c[1296] ), .Z(
        _f_permutation__round_out[619]) );
  XOR2_X2 _f_permutation__round__U3547  ( .A(_f_permutation__round__N4519 ), 
        .B(_f_permutation__round__c[1297] ), .Z(
        _f_permutation__round_out[620]) );
  XOR2_X2 _f_permutation__round__U3546  ( .A(_f_permutation__round__N4517 ), 
        .B(_f_permutation__round__c[1298] ), .Z(
        _f_permutation__round_out[621]) );
  XOR2_X2 _f_permutation__round__U3545  ( .A(_f_permutation__round__N4515 ), 
        .B(_f_permutation__round__c[1299] ), .Z(
        _f_permutation__round_out[622]) );
  XOR2_X2 _f_permutation__round__U3544  ( .A(_f_permutation__round__N4513 ), 
        .B(_f_permutation__round__c[1300] ), .Z(
        _f_permutation__round_out[623]) );
  XOR2_X2 _f_permutation__round__U3543  ( .A(_f_permutation__round__N4511 ), 
        .B(_f_permutation__round__c[1301] ), .Z(
        _f_permutation__round_out[624]) );
  XOR2_X2 _f_permutation__round__U3542  ( .A(_f_permutation__round__N4509 ), 
        .B(_f_permutation__round__c[1302] ), .Z(
        _f_permutation__round_out[625]) );
  XOR2_X2 _f_permutation__round__U3541  ( .A(_f_permutation__round__N4507 ), 
        .B(_f_permutation__round__c[1303] ), .Z(
        _f_permutation__round_out[626]) );
  XOR2_X2 _f_permutation__round__U3540  ( .A(_f_permutation__round__N4505 ), 
        .B(_f_permutation__round__c[1304] ), .Z(
        _f_permutation__round_out[627]) );
  XOR2_X2 _f_permutation__round__U3539  ( .A(_f_permutation__round__N4503 ), 
        .B(_f_permutation__round__c[1305] ), .Z(
        _f_permutation__round_out[628]) );
  XOR2_X2 _f_permutation__round__U3538  ( .A(_f_permutation__round__N4501 ), 
        .B(_f_permutation__round__c[1306] ), .Z(
        _f_permutation__round_out[629]) );
  XOR2_X2 _f_permutation__round__U3537  ( .A(_f_permutation__round__N4499 ), 
        .B(_f_permutation__round__c[1307] ), .Z(
        _f_permutation__round_out[630]) );
  XOR2_X2 _f_permutation__round__U3536  ( .A(_f_permutation__round__N4497 ), 
        .B(_f_permutation__round__c[1308] ), .Z(
        _f_permutation__round_out[631]) );
  XOR2_X2 _f_permutation__round__U3535  ( .A(_f_permutation__round__N4495 ), 
        .B(_f_permutation__round__c[1309] ), .Z(
        _f_permutation__round_out[632]) );
  XOR2_X2 _f_permutation__round__U3534  ( .A(_f_permutation__round__N4493 ), 
        .B(_f_permutation__round__c[1310] ), .Z(
        _f_permutation__round_out[633]) );
  XOR2_X2 _f_permutation__round__U3533  ( .A(_f_permutation__round__N4491 ), 
        .B(_f_permutation__round__c[1311] ), .Z(
        _f_permutation__round_out[634]) );
  XOR2_X2 _f_permutation__round__U3532  ( .A(_f_permutation__round__N4489 ), 
        .B(_f_permutation__round__c[1312] ), .Z(
        _f_permutation__round_out[635]) );
  XOR2_X2 _f_permutation__round__U3531  ( .A(_f_permutation__round__N4487 ), 
        .B(_f_permutation__round__c[1313] ), .Z(
        _f_permutation__round_out[636]) );
  XOR2_X2 _f_permutation__round__U3530  ( .A(_f_permutation__round__N4485 ), 
        .B(_f_permutation__round__c[1314] ), .Z(
        _f_permutation__round_out[637]) );
  XOR2_X2 _f_permutation__round__U3529  ( .A(_f_permutation__round__N4483 ), 
        .B(_f_permutation__round__c[1315] ), .Z(
        _f_permutation__round_out[638]) );
  XOR2_X2 _f_permutation__round__U3528  ( .A(_f_permutation__round__N4481 ), 
        .B(_f_permutation__round__c[1316] ), .Z(
        _f_permutation__round_out[639]) );
  XOR2_X2 _f_permutation__round__U3527  ( .A(_f_permutation__round__N4479 ), 
        .B(_f_permutation__round__c[302] ), .Z(_f_permutation__round_out[640]) );
  XOR2_X2 _f_permutation__round__U3526  ( .A(_f_permutation__round__N4477 ), 
        .B(_f_permutation__round__c[303] ), .Z(_f_permutation__round_out[641]) );
  XOR2_X2 _f_permutation__round__U3525  ( .A(_f_permutation__round__N4475 ), 
        .B(_f_permutation__round__c[304] ), .Z(_f_permutation__round_out[642]) );
  XOR2_X2 _f_permutation__round__U3524  ( .A(_f_permutation__round__N4473 ), 
        .B(_f_permutation__round__c[305] ), .Z(_f_permutation__round_out[643]) );
  XOR2_X2 _f_permutation__round__U3523  ( .A(_f_permutation__round__N4471 ), 
        .B(_f_permutation__round__c[306] ), .Z(_f_permutation__round_out[644]) );
  XOR2_X2 _f_permutation__round__U3522  ( .A(_f_permutation__round__N4469 ), 
        .B(_f_permutation__round__c[307] ), .Z(_f_permutation__round_out[645]) );
  XOR2_X2 _f_permutation__round__U3521  ( .A(_f_permutation__round__N4467 ), 
        .B(_f_permutation__round__c[308] ), .Z(_f_permutation__round_out[646]) );
  XOR2_X2 _f_permutation__round__U3520  ( .A(_f_permutation__round__N4465 ), 
        .B(_f_permutation__round__c[309] ), .Z(_f_permutation__round_out[647]) );
  XOR2_X2 _f_permutation__round__U3519  ( .A(_f_permutation__round__N4463 ), 
        .B(_f_permutation__round__c[310] ), .Z(_f_permutation__round_out[648]) );
  XOR2_X2 _f_permutation__round__U3518  ( .A(_f_permutation__round__N4461 ), 
        .B(_f_permutation__round__c[311] ), .Z(_f_permutation__round_out[649]) );
  XOR2_X2 _f_permutation__round__U3517  ( .A(_f_permutation__round__N4459 ), 
        .B(_f_permutation__round__c[312] ), .Z(_f_permutation__round_out[650]) );
  XOR2_X2 _f_permutation__round__U3516  ( .A(_f_permutation__round__N4457 ), 
        .B(_f_permutation__round__c[313] ), .Z(_f_permutation__round_out[651]) );
  XOR2_X2 _f_permutation__round__U3515  ( .A(_f_permutation__round__N4455 ), 
        .B(_f_permutation__round__c[314] ), .Z(_f_permutation__round_out[652]) );
  XOR2_X2 _f_permutation__round__U3514  ( .A(_f_permutation__round__N4453 ), 
        .B(_f_permutation__round__c[315] ), .Z(_f_permutation__round_out[653]) );
  XOR2_X2 _f_permutation__round__U3513  ( .A(_f_permutation__round__N4451 ), 
        .B(_f_permutation__round__c[316] ), .Z(_f_permutation__round_out[654]) );
  XOR2_X2 _f_permutation__round__U3512  ( .A(_f_permutation__round__N4449 ), 
        .B(_f_permutation__round__c[317] ), .Z(_f_permutation__round_out[655]) );
  XOR2_X2 _f_permutation__round__U3511  ( .A(_f_permutation__round__N4447 ), 
        .B(_f_permutation__round__c[318] ), .Z(_f_permutation__round_out[656]) );
  XOR2_X2 _f_permutation__round__U3510  ( .A(_f_permutation__round__N4445 ), 
        .B(_f_permutation__round__c[319] ), .Z(_f_permutation__round_out[657]) );
  XOR2_X2 _f_permutation__round__U3509  ( .A(_f_permutation__round__N4443 ), 
        .B(_f_permutation__round__c[256] ), .Z(_f_permutation__round_out[658]) );
  XOR2_X2 _f_permutation__round__U3508  ( .A(_f_permutation__round__N4441 ), 
        .B(_f_permutation__round__c[257] ), .Z(_f_permutation__round_out[659]) );
  XOR2_X2 _f_permutation__round__U3507  ( .A(_f_permutation__round__N4439 ), 
        .B(_f_permutation__round__c[258] ), .Z(_f_permutation__round_out[660]) );
  XOR2_X2 _f_permutation__round__U3506  ( .A(_f_permutation__round__N4437 ), 
        .B(_f_permutation__round__c[259] ), .Z(_f_permutation__round_out[661]) );
  XOR2_X2 _f_permutation__round__U3505  ( .A(_f_permutation__round__N4435 ), 
        .B(_f_permutation__round__c[260] ), .Z(_f_permutation__round_out[662]) );
  XOR2_X2 _f_permutation__round__U3504  ( .A(_f_permutation__round__N4433 ), 
        .B(_f_permutation__round__c[261] ), .Z(_f_permutation__round_out[663]) );
  XOR2_X2 _f_permutation__round__U3503  ( .A(_f_permutation__round__N4431 ), 
        .B(_f_permutation__round__c[262] ), .Z(_f_permutation__round_out[664]) );
  XOR2_X2 _f_permutation__round__U3502  ( .A(_f_permutation__round__N4429 ), 
        .B(_f_permutation__round__c[263] ), .Z(_f_permutation__round_out[665]) );
  XOR2_X2 _f_permutation__round__U3501  ( .A(_f_permutation__round__N4427 ), 
        .B(_f_permutation__round__c[264] ), .Z(_f_permutation__round_out[666]) );
  XOR2_X2 _f_permutation__round__U3500  ( .A(_f_permutation__round__N4425 ), 
        .B(_f_permutation__round__c[265] ), .Z(_f_permutation__round_out[667]) );
  XOR2_X2 _f_permutation__round__U3499  ( .A(_f_permutation__round__N4423 ), 
        .B(_f_permutation__round__c[266] ), .Z(_f_permutation__round_out[668]) );
  XOR2_X2 _f_permutation__round__U3498  ( .A(_f_permutation__round__N4421 ), 
        .B(_f_permutation__round__c[267] ), .Z(_f_permutation__round_out[669]) );
  XOR2_X2 _f_permutation__round__U3497  ( .A(_f_permutation__round__N4419 ), 
        .B(_f_permutation__round__c[268] ), .Z(_f_permutation__round_out[670]) );
  XOR2_X2 _f_permutation__round__U3496  ( .A(_f_permutation__round__N4417 ), 
        .B(_f_permutation__round__c[269] ), .Z(_f_permutation__round_out[671]) );
  XOR2_X2 _f_permutation__round__U3495  ( .A(_f_permutation__round__N4415 ), 
        .B(_f_permutation__round__c[270] ), .Z(_f_permutation__round_out[672]) );
  XOR2_X2 _f_permutation__round__U3494  ( .A(_f_permutation__round__N4413 ), 
        .B(_f_permutation__round__c[271] ), .Z(_f_permutation__round_out[673]) );
  XOR2_X2 _f_permutation__round__U3493  ( .A(_f_permutation__round__N4411 ), 
        .B(_f_permutation__round__c[272] ), .Z(_f_permutation__round_out[674]) );
  XOR2_X2 _f_permutation__round__U3492  ( .A(_f_permutation__round__N4409 ), 
        .B(_f_permutation__round__c[273] ), .Z(_f_permutation__round_out[675]) );
  XOR2_X2 _f_permutation__round__U3491  ( .A(_f_permutation__round__N4407 ), 
        .B(_f_permutation__round__c[274] ), .Z(_f_permutation__round_out[676]) );
  XOR2_X2 _f_permutation__round__U3490  ( .A(_f_permutation__round__N4405 ), 
        .B(_f_permutation__round__c[275] ), .Z(_f_permutation__round_out[677]) );
  XOR2_X2 _f_permutation__round__U3489  ( .A(_f_permutation__round__N4403 ), 
        .B(_f_permutation__round__c[276] ), .Z(_f_permutation__round_out[678]) );
  XOR2_X2 _f_permutation__round__U3488  ( .A(_f_permutation__round__N4401 ), 
        .B(_f_permutation__round__c[277] ), .Z(_f_permutation__round_out[679]) );
  XOR2_X2 _f_permutation__round__U3487  ( .A(_f_permutation__round__N4399 ), 
        .B(_f_permutation__round__c[278] ), .Z(_f_permutation__round_out[680]) );
  XOR2_X2 _f_permutation__round__U3486  ( .A(_f_permutation__round__N4397 ), 
        .B(_f_permutation__round__c[279] ), .Z(_f_permutation__round_out[681]) );
  XOR2_X2 _f_permutation__round__U3485  ( .A(_f_permutation__round__N4395 ), 
        .B(_f_permutation__round__c[280] ), .Z(_f_permutation__round_out[682]) );
  XOR2_X2 _f_permutation__round__U3484  ( .A(_f_permutation__round__N4393 ), 
        .B(_f_permutation__round__c[281] ), .Z(_f_permutation__round_out[683]) );
  XOR2_X2 _f_permutation__round__U3483  ( .A(_f_permutation__round__N4391 ), 
        .B(_f_permutation__round__c[282] ), .Z(_f_permutation__round_out[684]) );
  XOR2_X2 _f_permutation__round__U3482  ( .A(_f_permutation__round__N4389 ), 
        .B(_f_permutation__round__c[283] ), .Z(_f_permutation__round_out[685]) );
  XOR2_X2 _f_permutation__round__U3481  ( .A(_f_permutation__round__N4387 ), 
        .B(_f_permutation__round__c[284] ), .Z(_f_permutation__round_out[686]) );
  XOR2_X2 _f_permutation__round__U3480  ( .A(_f_permutation__round__N4385 ), 
        .B(_f_permutation__round__c[285] ), .Z(_f_permutation__round_out[687]) );
  XOR2_X2 _f_permutation__round__U3479  ( .A(_f_permutation__round__N4383 ), 
        .B(_f_permutation__round__c[286] ), .Z(_f_permutation__round_out[688]) );
  XOR2_X2 _f_permutation__round__U3478  ( .A(_f_permutation__round__N4381 ), 
        .B(_f_permutation__round__c[287] ), .Z(_f_permutation__round_out[689]) );
  XOR2_X2 _f_permutation__round__U3477  ( .A(_f_permutation__round__N4379 ), 
        .B(_f_permutation__round__c[288] ), .Z(_f_permutation__round_out[690]) );
  XOR2_X2 _f_permutation__round__U3476  ( .A(_f_permutation__round__N4377 ), 
        .B(_f_permutation__round__c[289] ), .Z(_f_permutation__round_out[691]) );
  XOR2_X2 _f_permutation__round__U3475  ( .A(_f_permutation__round__N4375 ), 
        .B(_f_permutation__round__c[290] ), .Z(_f_permutation__round_out[692]) );
  XOR2_X2 _f_permutation__round__U3474  ( .A(_f_permutation__round__N4373 ), 
        .B(_f_permutation__round__c[291] ), .Z(_f_permutation__round_out[693]) );
  XOR2_X2 _f_permutation__round__U3473  ( .A(_f_permutation__round__N4371 ), 
        .B(_f_permutation__round__c[292] ), .Z(_f_permutation__round_out[694]) );
  XOR2_X2 _f_permutation__round__U3472  ( .A(_f_permutation__round__N4369 ), 
        .B(_f_permutation__round__c[293] ), .Z(_f_permutation__round_out[695]) );
  XOR2_X2 _f_permutation__round__U3471  ( .A(_f_permutation__round__N4367 ), 
        .B(_f_permutation__round__c[294] ), .Z(_f_permutation__round_out[696]) );
  XOR2_X2 _f_permutation__round__U3470  ( .A(_f_permutation__round__N4365 ), 
        .B(_f_permutation__round__c[295] ), .Z(_f_permutation__round_out[697]) );
  XOR2_X2 _f_permutation__round__U3469  ( .A(_f_permutation__round__N4363 ), 
        .B(_f_permutation__round__c[296] ), .Z(_f_permutation__round_out[698]) );
  XOR2_X2 _f_permutation__round__U3468  ( .A(_f_permutation__round__N4361 ), 
        .B(_f_permutation__round__c[297] ), .Z(_f_permutation__round_out[699]) );
  XOR2_X2 _f_permutation__round__U3467  ( .A(_f_permutation__round__N4359 ), 
        .B(_f_permutation__round__c[298] ), .Z(_f_permutation__round_out[700]) );
  XOR2_X2 _f_permutation__round__U3466  ( .A(_f_permutation__round__N4357 ), 
        .B(_f_permutation__round__c[299] ), .Z(_f_permutation__round_out[701]) );
  XOR2_X2 _f_permutation__round__U3465  ( .A(_f_permutation__round__N4355 ), 
        .B(_f_permutation__round__c[300] ), .Z(_f_permutation__round_out[702]) );
  XOR2_X2 _f_permutation__round__U3464  ( .A(_f_permutation__round__N4353 ), 
        .B(_f_permutation__round__c[301] ), .Z(_f_permutation__round_out[703]) );
  XOR2_X2 _f_permutation__round__U3463  ( .A(_f_permutation__round__N4351 ), 
        .B(_f_permutation__round__c[1528] ), .Z(
        _f_permutation__round_out[704]) );
  XOR2_X2 _f_permutation__round__U3462  ( .A(_f_permutation__round__N4349 ), 
        .B(_f_permutation__round__c[1529] ), .Z(
        _f_permutation__round_out[705]) );
  XOR2_X2 _f_permutation__round__U3461  ( .A(_f_permutation__round__N4347 ), 
        .B(_f_permutation__round__c[1530] ), .Z(
        _f_permutation__round_out[706]) );
  XOR2_X2 _f_permutation__round__U3460  ( .A(_f_permutation__round__N4345 ), 
        .B(_f_permutation__round__c[1531] ), .Z(
        _f_permutation__round_out[707]) );
  XOR2_X2 _f_permutation__round__U3459  ( .A(_f_permutation__round__N4343 ), 
        .B(_f_permutation__round__c[1532] ), .Z(
        _f_permutation__round_out[708]) );
  XOR2_X2 _f_permutation__round__U3458  ( .A(_f_permutation__round__N4341 ), 
        .B(_f_permutation__round__c[1533] ), .Z(
        _f_permutation__round_out[709]) );
  XOR2_X2 _f_permutation__round__U3457  ( .A(_f_permutation__round__N4339 ), 
        .B(_f_permutation__round__c[1534] ), .Z(
        _f_permutation__round_out[710]) );
  XOR2_X2 _f_permutation__round__U3456  ( .A(_f_permutation__round__N4337 ), 
        .B(_f_permutation__round__c[1535] ), .Z(
        _f_permutation__round_out[711]) );
  XOR2_X2 _f_permutation__round__U3455  ( .A(_f_permutation__round__N4335 ), 
        .B(_f_permutation__round__c[1472] ), .Z(
        _f_permutation__round_out[712]) );
  XOR2_X2 _f_permutation__round__U3454  ( .A(_f_permutation__round__N4333 ), 
        .B(_f_permutation__round__c[1473] ), .Z(
        _f_permutation__round_out[713]) );
  XOR2_X2 _f_permutation__round__U3453  ( .A(_f_permutation__round__N4331 ), 
        .B(_f_permutation__round__c[1474] ), .Z(
        _f_permutation__round_out[714]) );
  XOR2_X2 _f_permutation__round__U3452  ( .A(_f_permutation__round__N4329 ), 
        .B(_f_permutation__round__c[1475] ), .Z(
        _f_permutation__round_out[715]) );
  XOR2_X2 _f_permutation__round__U3451  ( .A(_f_permutation__round__N4327 ), 
        .B(_f_permutation__round__c[1476] ), .Z(
        _f_permutation__round_out[716]) );
  XOR2_X2 _f_permutation__round__U3450  ( .A(_f_permutation__round__N4325 ), 
        .B(_f_permutation__round__c[1477] ), .Z(
        _f_permutation__round_out[717]) );
  XOR2_X2 _f_permutation__round__U3449  ( .A(_f_permutation__round__N4323 ), 
        .B(_f_permutation__round__c[1478] ), .Z(
        _f_permutation__round_out[718]) );
  XOR2_X2 _f_permutation__round__U3448  ( .A(_f_permutation__round__N4321 ), 
        .B(_f_permutation__round__c[1479] ), .Z(
        _f_permutation__round_out[719]) );
  XOR2_X2 _f_permutation__round__U3447  ( .A(_f_permutation__round__N4319 ), 
        .B(_f_permutation__round__c[1480] ), .Z(
        _f_permutation__round_out[720]) );
  XOR2_X2 _f_permutation__round__U3446  ( .A(_f_permutation__round__N4317 ), 
        .B(_f_permutation__round__c[1481] ), .Z(
        _f_permutation__round_out[721]) );
  XOR2_X2 _f_permutation__round__U3445  ( .A(_f_permutation__round__N4315 ), 
        .B(_f_permutation__round__c[1482] ), .Z(
        _f_permutation__round_out[722]) );
  XOR2_X2 _f_permutation__round__U3444  ( .A(_f_permutation__round__N4313 ), 
        .B(_f_permutation__round__c[1483] ), .Z(
        _f_permutation__round_out[723]) );
  XOR2_X2 _f_permutation__round__U3443  ( .A(_f_permutation__round__N4311 ), 
        .B(_f_permutation__round__c[1484] ), .Z(
        _f_permutation__round_out[724]) );
  XOR2_X2 _f_permutation__round__U3442  ( .A(_f_permutation__round__N4309 ), 
        .B(_f_permutation__round__c[1485] ), .Z(
        _f_permutation__round_out[725]) );
  XOR2_X2 _f_permutation__round__U3441  ( .A(_f_permutation__round__N4307 ), 
        .B(_f_permutation__round__c[1486] ), .Z(
        _f_permutation__round_out[726]) );
  XOR2_X2 _f_permutation__round__U3440  ( .A(_f_permutation__round__N4305 ), 
        .B(_f_permutation__round__c[1487] ), .Z(
        _f_permutation__round_out[727]) );
  XOR2_X2 _f_permutation__round__U3439  ( .A(_f_permutation__round__N4303 ), 
        .B(_f_permutation__round__c[1488] ), .Z(
        _f_permutation__round_out[728]) );
  XOR2_X2 _f_permutation__round__U3438  ( .A(_f_permutation__round__N4301 ), 
        .B(_f_permutation__round__c[1489] ), .Z(
        _f_permutation__round_out[729]) );
  XOR2_X2 _f_permutation__round__U3437  ( .A(_f_permutation__round__N4299 ), 
        .B(_f_permutation__round__c[1490] ), .Z(
        _f_permutation__round_out[730]) );
  XOR2_X2 _f_permutation__round__U3436  ( .A(_f_permutation__round__N4297 ), 
        .B(_f_permutation__round__c[1491] ), .Z(
        _f_permutation__round_out[731]) );
  XOR2_X2 _f_permutation__round__U3435  ( .A(_f_permutation__round__N4295 ), 
        .B(_f_permutation__round__c[1492] ), .Z(
        _f_permutation__round_out[732]) );
  XOR2_X2 _f_permutation__round__U3434  ( .A(_f_permutation__round__N4293 ), 
        .B(_f_permutation__round__c[1493] ), .Z(
        _f_permutation__round_out[733]) );
  XOR2_X2 _f_permutation__round__U3433  ( .A(_f_permutation__round__N4291 ), 
        .B(_f_permutation__round__c[1494] ), .Z(
        _f_permutation__round_out[734]) );
  XOR2_X2 _f_permutation__round__U3432  ( .A(_f_permutation__round__N4289 ), 
        .B(_f_permutation__round__c[1495] ), .Z(
        _f_permutation__round_out[735]) );
  XOR2_X2 _f_permutation__round__U3431  ( .A(_f_permutation__round__N4287 ), 
        .B(_f_permutation__round__c[1496] ), .Z(
        _f_permutation__round_out[736]) );
  XOR2_X2 _f_permutation__round__U3430  ( .A(_f_permutation__round__N4285 ), 
        .B(_f_permutation__round__c[1497] ), .Z(
        _f_permutation__round_out[737]) );
  XOR2_X2 _f_permutation__round__U3429  ( .A(_f_permutation__round__N4283 ), 
        .B(_f_permutation__round__c[1498] ), .Z(
        _f_permutation__round_out[738]) );
  XOR2_X2 _f_permutation__round__U3428  ( .A(_f_permutation__round__N4281 ), 
        .B(_f_permutation__round__c[1499] ), .Z(
        _f_permutation__round_out[739]) );
  XOR2_X2 _f_permutation__round__U3427  ( .A(_f_permutation__round__N4279 ), 
        .B(_f_permutation__round__c[1500] ), .Z(
        _f_permutation__round_out[740]) );
  XOR2_X2 _f_permutation__round__U3426  ( .A(_f_permutation__round__N4277 ), 
        .B(_f_permutation__round__c[1501] ), .Z(
        _f_permutation__round_out[741]) );
  XOR2_X2 _f_permutation__round__U3425  ( .A(_f_permutation__round__N4275 ), 
        .B(_f_permutation__round__c[1502] ), .Z(
        _f_permutation__round_out[742]) );
  XOR2_X2 _f_permutation__round__U3424  ( .A(_f_permutation__round__N4273 ), 
        .B(_f_permutation__round__c[1503] ), .Z(
        _f_permutation__round_out[743]) );
  XOR2_X2 _f_permutation__round__U3423  ( .A(_f_permutation__round__N4271 ), 
        .B(_f_permutation__round__c[1504] ), .Z(
        _f_permutation__round_out[744]) );
  XOR2_X2 _f_permutation__round__U3422  ( .A(_f_permutation__round__N4269 ), 
        .B(_f_permutation__round__c[1505] ), .Z(
        _f_permutation__round_out[745]) );
  XOR2_X2 _f_permutation__round__U3421  ( .A(_f_permutation__round__N4267 ), 
        .B(_f_permutation__round__c[1506] ), .Z(
        _f_permutation__round_out[746]) );
  XOR2_X2 _f_permutation__round__U3420  ( .A(_f_permutation__round__N4265 ), 
        .B(_f_permutation__round__c[1507] ), .Z(
        _f_permutation__round_out[747]) );
  XOR2_X2 _f_permutation__round__U3419  ( .A(_f_permutation__round__N4263 ), 
        .B(_f_permutation__round__c[1508] ), .Z(
        _f_permutation__round_out[748]) );
  XOR2_X2 _f_permutation__round__U3418  ( .A(_f_permutation__round__N4261 ), 
        .B(_f_permutation__round__c[1509] ), .Z(
        _f_permutation__round_out[749]) );
  XOR2_X2 _f_permutation__round__U3417  ( .A(_f_permutation__round__N4259 ), 
        .B(_f_permutation__round__c[1510] ), .Z(
        _f_permutation__round_out[750]) );
  XOR2_X2 _f_permutation__round__U3416  ( .A(_f_permutation__round__N4257 ), 
        .B(_f_permutation__round__c[1511] ), .Z(
        _f_permutation__round_out[751]) );
  XOR2_X2 _f_permutation__round__U3415  ( .A(_f_permutation__round__N4255 ), 
        .B(_f_permutation__round__c[1512] ), .Z(
        _f_permutation__round_out[752]) );
  XOR2_X2 _f_permutation__round__U3414  ( .A(_f_permutation__round__N4253 ), 
        .B(_f_permutation__round__c[1513] ), .Z(
        _f_permutation__round_out[753]) );
  XOR2_X2 _f_permutation__round__U3413  ( .A(_f_permutation__round__N4251 ), 
        .B(_f_permutation__round__c[1514] ), .Z(
        _f_permutation__round_out[754]) );
  XOR2_X2 _f_permutation__round__U3412  ( .A(_f_permutation__round__N4249 ), 
        .B(_f_permutation__round__c[1515] ), .Z(
        _f_permutation__round_out[755]) );
  XOR2_X2 _f_permutation__round__U3411  ( .A(_f_permutation__round__N4247 ), 
        .B(_f_permutation__round__c[1516] ), .Z(
        _f_permutation__round_out[756]) );
  XOR2_X2 _f_permutation__round__U3410  ( .A(_f_permutation__round__N4245 ), 
        .B(_f_permutation__round__c[1517] ), .Z(
        _f_permutation__round_out[757]) );
  XOR2_X2 _f_permutation__round__U3409  ( .A(_f_permutation__round__N4243 ), 
        .B(_f_permutation__round__c[1518] ), .Z(
        _f_permutation__round_out[758]) );
  XOR2_X2 _f_permutation__round__U3408  ( .A(_f_permutation__round__N4241 ), 
        .B(_f_permutation__round__c[1519] ), .Z(
        _f_permutation__round_out[759]) );
  XOR2_X2 _f_permutation__round__U3407  ( .A(_f_permutation__round__N4239 ), 
        .B(_f_permutation__round__c[1520] ), .Z(
        _f_permutation__round_out[760]) );
  XOR2_X2 _f_permutation__round__U3406  ( .A(_f_permutation__round__N4237 ), 
        .B(_f_permutation__round__c[1521] ), .Z(
        _f_permutation__round_out[761]) );
  XOR2_X2 _f_permutation__round__U3405  ( .A(_f_permutation__round__N4235 ), 
        .B(_f_permutation__round__c[1522] ), .Z(
        _f_permutation__round_out[762]) );
  XOR2_X2 _f_permutation__round__U3404  ( .A(_f_permutation__round__N4233 ), 
        .B(_f_permutation__round__c[1523] ), .Z(
        _f_permutation__round_out[763]) );
  XOR2_X2 _f_permutation__round__U3403  ( .A(_f_permutation__round__N4231 ), 
        .B(_f_permutation__round__c[1524] ), .Z(
        _f_permutation__round_out[764]) );
  XOR2_X2 _f_permutation__round__U3402  ( .A(_f_permutation__round__N4229 ), 
        .B(_f_permutation__round__c[1525] ), .Z(
        _f_permutation__round_out[765]) );
  XOR2_X2 _f_permutation__round__U3401  ( .A(_f_permutation__round__N4227 ), 
        .B(_f_permutation__round__c[1526] ), .Z(
        _f_permutation__round_out[766]) );
  XOR2_X2 _f_permutation__round__U3400  ( .A(_f_permutation__round__N4225 ), 
        .B(_f_permutation__round__c[1527] ), .Z(
        _f_permutation__round_out[767]) );
  XOR2_X2 _f_permutation__round__U3399  ( .A(_f_permutation__round__N4223 ), 
        .B(_f_permutation__round__c[1127] ), .Z(
        _f_permutation__round_out[768]) );
  XOR2_X2 _f_permutation__round__U3398  ( .A(_f_permutation__round__N4221 ), 
        .B(_f_permutation__round__c[1128] ), .Z(
        _f_permutation__round_out[769]) );
  XOR2_X2 _f_permutation__round__U3397  ( .A(_f_permutation__round__N4219 ), 
        .B(_f_permutation__round__c[1129] ), .Z(
        _f_permutation__round_out[770]) );
  XOR2_X2 _f_permutation__round__U3396  ( .A(_f_permutation__round__N4217 ), 
        .B(_f_permutation__round__c[1130] ), .Z(
        _f_permutation__round_out[771]) );
  XOR2_X2 _f_permutation__round__U3395  ( .A(_f_permutation__round__N4215 ), 
        .B(_f_permutation__round__c[1131] ), .Z(
        _f_permutation__round_out[772]) );
  XOR2_X2 _f_permutation__round__U3394  ( .A(_f_permutation__round__N4213 ), 
        .B(_f_permutation__round__c[1132] ), .Z(
        _f_permutation__round_out[773]) );
  XOR2_X2 _f_permutation__round__U3393  ( .A(_f_permutation__round__N4211 ), 
        .B(_f_permutation__round__c[1133] ), .Z(
        _f_permutation__round_out[774]) );
  XOR2_X2 _f_permutation__round__U3392  ( .A(_f_permutation__round__N4209 ), 
        .B(_f_permutation__round__c[1134] ), .Z(
        _f_permutation__round_out[775]) );
  XOR2_X2 _f_permutation__round__U3391  ( .A(_f_permutation__round__N4207 ), 
        .B(_f_permutation__round__c[1135] ), .Z(
        _f_permutation__round_out[776]) );
  XOR2_X2 _f_permutation__round__U3390  ( .A(_f_permutation__round__N4205 ), 
        .B(_f_permutation__round__c[1136] ), .Z(
        _f_permutation__round_out[777]) );
  XOR2_X2 _f_permutation__round__U3389  ( .A(_f_permutation__round__N4203 ), 
        .B(_f_permutation__round__c[1137] ), .Z(
        _f_permutation__round_out[778]) );
  XOR2_X2 _f_permutation__round__U3388  ( .A(_f_permutation__round__N4201 ), 
        .B(_f_permutation__round__c[1138] ), .Z(
        _f_permutation__round_out[779]) );
  XOR2_X2 _f_permutation__round__U3387  ( .A(_f_permutation__round__N4199 ), 
        .B(_f_permutation__round__c[1139] ), .Z(
        _f_permutation__round_out[780]) );
  XOR2_X2 _f_permutation__round__U3386  ( .A(_f_permutation__round__N4197 ), 
        .B(_f_permutation__round__c[1140] ), .Z(
        _f_permutation__round_out[781]) );
  XOR2_X2 _f_permutation__round__U3385  ( .A(_f_permutation__round__N4195 ), 
        .B(_f_permutation__round__c[1141] ), .Z(
        _f_permutation__round_out[782]) );
  XOR2_X2 _f_permutation__round__U3384  ( .A(_f_permutation__round__N4193 ), 
        .B(_f_permutation__round__c[1142] ), .Z(
        _f_permutation__round_out[783]) );
  XOR2_X2 _f_permutation__round__U3383  ( .A(_f_permutation__round__N4191 ), 
        .B(_f_permutation__round__c[1143] ), .Z(
        _f_permutation__round_out[784]) );
  XOR2_X2 _f_permutation__round__U3382  ( .A(_f_permutation__round__N4189 ), 
        .B(_f_permutation__round__c[1144] ), .Z(
        _f_permutation__round_out[785]) );
  XOR2_X2 _f_permutation__round__U3381  ( .A(_f_permutation__round__N4187 ), 
        .B(_f_permutation__round__c[1145] ), .Z(
        _f_permutation__round_out[786]) );
  XOR2_X2 _f_permutation__round__U3380  ( .A(_f_permutation__round__N4185 ), 
        .B(_f_permutation__round__c[1146] ), .Z(
        _f_permutation__round_out[787]) );
  XOR2_X2 _f_permutation__round__U3379  ( .A(_f_permutation__round__N4183 ), 
        .B(_f_permutation__round__c[1147] ), .Z(
        _f_permutation__round_out[788]) );
  XOR2_X2 _f_permutation__round__U3378  ( .A(_f_permutation__round__N4181 ), 
        .B(_f_permutation__round__c[1148] ), .Z(
        _f_permutation__round_out[789]) );
  XOR2_X2 _f_permutation__round__U3377  ( .A(_f_permutation__round__N4179 ), 
        .B(_f_permutation__round__c[1149] ), .Z(
        _f_permutation__round_out[790]) );
  XOR2_X2 _f_permutation__round__U3376  ( .A(_f_permutation__round__N4177 ), 
        .B(_f_permutation__round__c[1150] ), .Z(
        _f_permutation__round_out[791]) );
  XOR2_X2 _f_permutation__round__U3375  ( .A(_f_permutation__round__N4175 ), 
        .B(_f_permutation__round__c[1151] ), .Z(
        _f_permutation__round_out[792]) );
  XOR2_X2 _f_permutation__round__U3374  ( .A(_f_permutation__round__N4173 ), 
        .B(_f_permutation__round__c[1088] ), .Z(
        _f_permutation__round_out[793]) );
  XOR2_X2 _f_permutation__round__U3373  ( .A(_f_permutation__round__N4171 ), 
        .B(_f_permutation__round__c[1089] ), .Z(
        _f_permutation__round_out[794]) );
  XOR2_X2 _f_permutation__round__U3372  ( .A(_f_permutation__round__N4169 ), 
        .B(_f_permutation__round__c[1090] ), .Z(
        _f_permutation__round_out[795]) );
  XOR2_X2 _f_permutation__round__U3371  ( .A(_f_permutation__round__N4167 ), 
        .B(_f_permutation__round__c[1091] ), .Z(
        _f_permutation__round_out[796]) );
  XOR2_X2 _f_permutation__round__U3370  ( .A(_f_permutation__round__N4165 ), 
        .B(_f_permutation__round__c[1092] ), .Z(
        _f_permutation__round_out[797]) );
  XOR2_X2 _f_permutation__round__U3369  ( .A(_f_permutation__round__N4163 ), 
        .B(_f_permutation__round__c[1093] ), .Z(
        _f_permutation__round_out[798]) );
  XOR2_X2 _f_permutation__round__U3368  ( .A(_f_permutation__round__N4161 ), 
        .B(_f_permutation__round__c[1094] ), .Z(
        _f_permutation__round_out[799]) );
  XOR2_X2 _f_permutation__round__U3367  ( .A(_f_permutation__round__N4159 ), 
        .B(_f_permutation__round__c[1095] ), .Z(
        _f_permutation__round_out[800]) );
  XOR2_X2 _f_permutation__round__U3366  ( .A(_f_permutation__round__N4157 ), 
        .B(_f_permutation__round__c[1096] ), .Z(
        _f_permutation__round_out[801]) );
  XOR2_X2 _f_permutation__round__U3365  ( .A(_f_permutation__round__N4155 ), 
        .B(_f_permutation__round__c[1097] ), .Z(
        _f_permutation__round_out[802]) );
  XOR2_X2 _f_permutation__round__U3364  ( .A(_f_permutation__round__N4153 ), 
        .B(_f_permutation__round__c[1098] ), .Z(
        _f_permutation__round_out[803]) );
  XOR2_X2 _f_permutation__round__U3363  ( .A(_f_permutation__round__N4151 ), 
        .B(_f_permutation__round__c[1099] ), .Z(
        _f_permutation__round_out[804]) );
  XOR2_X2 _f_permutation__round__U3362  ( .A(_f_permutation__round__N4149 ), 
        .B(_f_permutation__round__c[1100] ), .Z(
        _f_permutation__round_out[805]) );
  XOR2_X2 _f_permutation__round__U3361  ( .A(_f_permutation__round__N4147 ), 
        .B(_f_permutation__round__c[1101] ), .Z(
        _f_permutation__round_out[806]) );
  XOR2_X2 _f_permutation__round__U3360  ( .A(_f_permutation__round__N4145 ), 
        .B(_f_permutation__round__c[1102] ), .Z(
        _f_permutation__round_out[807]) );
  XOR2_X2 _f_permutation__round__U3359  ( .A(_f_permutation__round__N4143 ), 
        .B(_f_permutation__round__c[1103] ), .Z(
        _f_permutation__round_out[808]) );
  XOR2_X2 _f_permutation__round__U3358  ( .A(_f_permutation__round__N4141 ), 
        .B(_f_permutation__round__c[1104] ), .Z(
        _f_permutation__round_out[809]) );
  XOR2_X2 _f_permutation__round__U3357  ( .A(_f_permutation__round__N4139 ), 
        .B(_f_permutation__round__c[1105] ), .Z(
        _f_permutation__round_out[810]) );
  XOR2_X2 _f_permutation__round__U3356  ( .A(_f_permutation__round__N4137 ), 
        .B(_f_permutation__round__c[1106] ), .Z(
        _f_permutation__round_out[811]) );
  XOR2_X2 _f_permutation__round__U3355  ( .A(_f_permutation__round__N4135 ), 
        .B(_f_permutation__round__c[1107] ), .Z(
        _f_permutation__round_out[812]) );
  XOR2_X2 _f_permutation__round__U3354  ( .A(_f_permutation__round__N4133 ), 
        .B(_f_permutation__round__c[1108] ), .Z(
        _f_permutation__round_out[813]) );
  XOR2_X2 _f_permutation__round__U3353  ( .A(_f_permutation__round__N4131 ), 
        .B(_f_permutation__round__c[1109] ), .Z(
        _f_permutation__round_out[814]) );
  XOR2_X2 _f_permutation__round__U3352  ( .A(_f_permutation__round__N4129 ), 
        .B(_f_permutation__round__c[1110] ), .Z(
        _f_permutation__round_out[815]) );
  XOR2_X2 _f_permutation__round__U3351  ( .A(_f_permutation__round__N4127 ), 
        .B(_f_permutation__round__c[1111] ), .Z(
        _f_permutation__round_out[816]) );
  XOR2_X2 _f_permutation__round__U3350  ( .A(_f_permutation__round__N4125 ), 
        .B(_f_permutation__round__c[1112] ), .Z(
        _f_permutation__round_out[817]) );
  XOR2_X2 _f_permutation__round__U3349  ( .A(_f_permutation__round__N4123 ), 
        .B(_f_permutation__round__c[1113] ), .Z(
        _f_permutation__round_out[818]) );
  XOR2_X2 _f_permutation__round__U3348  ( .A(_f_permutation__round__N4121 ), 
        .B(_f_permutation__round__c[1114] ), .Z(
        _f_permutation__round_out[819]) );
  XOR2_X2 _f_permutation__round__U3347  ( .A(_f_permutation__round__N4119 ), 
        .B(_f_permutation__round__c[1115] ), .Z(
        _f_permutation__round_out[820]) );
  XOR2_X2 _f_permutation__round__U3346  ( .A(_f_permutation__round__N4117 ), 
        .B(_f_permutation__round__c[1116] ), .Z(
        _f_permutation__round_out[821]) );
  XOR2_X2 _f_permutation__round__U3345  ( .A(_f_permutation__round__N4115 ), 
        .B(_f_permutation__round__c[1117] ), .Z(
        _f_permutation__round_out[822]) );
  XOR2_X2 _f_permutation__round__U3344  ( .A(_f_permutation__round__N4113 ), 
        .B(_f_permutation__round__c[1118] ), .Z(
        _f_permutation__round_out[823]) );
  XOR2_X2 _f_permutation__round__U3343  ( .A(_f_permutation__round__N4111 ), 
        .B(_f_permutation__round__c[1119] ), .Z(
        _f_permutation__round_out[824]) );
  XOR2_X2 _f_permutation__round__U3342  ( .A(_f_permutation__round__N4109 ), 
        .B(_f_permutation__round__c[1120] ), .Z(
        _f_permutation__round_out[825]) );
  XOR2_X2 _f_permutation__round__U3341  ( .A(_f_permutation__round__N4107 ), 
        .B(_f_permutation__round__c[1121] ), .Z(
        _f_permutation__round_out[826]) );
  XOR2_X2 _f_permutation__round__U3340  ( .A(_f_permutation__round__N4105 ), 
        .B(_f_permutation__round__c[1122] ), .Z(
        _f_permutation__round_out[827]) );
  XOR2_X2 _f_permutation__round__U3339  ( .A(_f_permutation__round__N4103 ), 
        .B(_f_permutation__round__c[1123] ), .Z(
        _f_permutation__round_out[828]) );
  XOR2_X2 _f_permutation__round__U3338  ( .A(_f_permutation__round__N4101 ), 
        .B(_f_permutation__round__c[1124] ), .Z(
        _f_permutation__round_out[829]) );
  XOR2_X2 _f_permutation__round__U3337  ( .A(_f_permutation__round__N4099 ), 
        .B(_f_permutation__round__c[1125] ), .Z(
        _f_permutation__round_out[830]) );
  XOR2_X2 _f_permutation__round__U3336  ( .A(_f_permutation__round__N4097 ), 
        .B(_f_permutation__round__c[1126] ), .Z(
        _f_permutation__round_out[831]) );
  XOR2_X2 _f_permutation__round__U3335  ( .A(_f_permutation__round__N4095 ), 
        .B(_f_permutation__round__c[762] ), .Z(_f_permutation__round_out[832]) );
  XOR2_X2 _f_permutation__round__U3334  ( .A(_f_permutation__round__N4093 ), 
        .B(_f_permutation__round__c[763] ), .Z(_f_permutation__round_out[833]) );
  XOR2_X2 _f_permutation__round__U3333  ( .A(_f_permutation__round__N4091 ), 
        .B(_f_permutation__round__c[764] ), .Z(_f_permutation__round_out[834]) );
  XOR2_X2 _f_permutation__round__U3332  ( .A(_f_permutation__round__N4089 ), 
        .B(_f_permutation__round__c[765] ), .Z(_f_permutation__round_out[835]) );
  XOR2_X2 _f_permutation__round__U3331  ( .A(_f_permutation__round__N4087 ), 
        .B(_f_permutation__round__c[766] ), .Z(_f_permutation__round_out[836]) );
  XOR2_X2 _f_permutation__round__U3330  ( .A(_f_permutation__round__N4085 ), 
        .B(_f_permutation__round__c[767] ), .Z(_f_permutation__round_out[837]) );
  XOR2_X2 _f_permutation__round__U3329  ( .A(_f_permutation__round__N4083 ), 
        .B(_f_permutation__round__c[704] ), .Z(_f_permutation__round_out[838]) );
  XOR2_X2 _f_permutation__round__U3328  ( .A(_f_permutation__round__N4081 ), 
        .B(_f_permutation__round__c[705] ), .Z(_f_permutation__round_out[839]) );
  XOR2_X2 _f_permutation__round__U3327  ( .A(_f_permutation__round__N4079 ), 
        .B(_f_permutation__round__c[706] ), .Z(_f_permutation__round_out[840]) );
  XOR2_X2 _f_permutation__round__U3326  ( .A(_f_permutation__round__N4077 ), 
        .B(_f_permutation__round__c[707] ), .Z(_f_permutation__round_out[841]) );
  XOR2_X2 _f_permutation__round__U3325  ( .A(_f_permutation__round__N4075 ), 
        .B(_f_permutation__round__c[708] ), .Z(_f_permutation__round_out[842]) );
  XOR2_X2 _f_permutation__round__U3324  ( .A(_f_permutation__round__N4073 ), 
        .B(_f_permutation__round__c[709] ), .Z(_f_permutation__round_out[843]) );
  XOR2_X2 _f_permutation__round__U3323  ( .A(_f_permutation__round__N4071 ), 
        .B(_f_permutation__round__c[710] ), .Z(_f_permutation__round_out[844]) );
  XOR2_X2 _f_permutation__round__U3322  ( .A(_f_permutation__round__N4069 ), 
        .B(_f_permutation__round__c[711] ), .Z(_f_permutation__round_out[845]) );
  XOR2_X2 _f_permutation__round__U3321  ( .A(_f_permutation__round__N4067 ), 
        .B(_f_permutation__round__c[712] ), .Z(_f_permutation__round_out[846]) );
  XOR2_X2 _f_permutation__round__U3320  ( .A(_f_permutation__round__N4065 ), 
        .B(_f_permutation__round__c[713] ), .Z(_f_permutation__round_out[847]) );
  XOR2_X2 _f_permutation__round__U3319  ( .A(_f_permutation__round__N4063 ), 
        .B(_f_permutation__round__c[714] ), .Z(_f_permutation__round_out[848]) );
  XOR2_X2 _f_permutation__round__U3318  ( .A(_f_permutation__round__N4061 ), 
        .B(_f_permutation__round__c[715] ), .Z(_f_permutation__round_out[849]) );
  XOR2_X2 _f_permutation__round__U3317  ( .A(_f_permutation__round__N4059 ), 
        .B(_f_permutation__round__c[716] ), .Z(_f_permutation__round_out[850]) );
  XOR2_X2 _f_permutation__round__U3316  ( .A(_f_permutation__round__N4057 ), 
        .B(_f_permutation__round__c[717] ), .Z(_f_permutation__round_out[851]) );
  XOR2_X2 _f_permutation__round__U3315  ( .A(_f_permutation__round__N4055 ), 
        .B(_f_permutation__round__c[718] ), .Z(_f_permutation__round_out[852]) );
  XOR2_X2 _f_permutation__round__U3314  ( .A(_f_permutation__round__N4053 ), 
        .B(_f_permutation__round__c[719] ), .Z(_f_permutation__round_out[853]) );
  XOR2_X2 _f_permutation__round__U3313  ( .A(_f_permutation__round__N4051 ), 
        .B(_f_permutation__round__c[720] ), .Z(_f_permutation__round_out[854]) );
  XOR2_X2 _f_permutation__round__U3312  ( .A(_f_permutation__round__N4049 ), 
        .B(_f_permutation__round__c[721] ), .Z(_f_permutation__round_out[855]) );
  XOR2_X2 _f_permutation__round__U3311  ( .A(_f_permutation__round__N4047 ), 
        .B(_f_permutation__round__c[722] ), .Z(_f_permutation__round_out[856]) );
  XOR2_X2 _f_permutation__round__U3310  ( .A(_f_permutation__round__N4045 ), 
        .B(_f_permutation__round__c[723] ), .Z(_f_permutation__round_out[857]) );
  XOR2_X2 _f_permutation__round__U3309  ( .A(_f_permutation__round__N4043 ), 
        .B(_f_permutation__round__c[724] ), .Z(_f_permutation__round_out[858]) );
  XOR2_X2 _f_permutation__round__U3308  ( .A(_f_permutation__round__N4041 ), 
        .B(_f_permutation__round__c[725] ), .Z(_f_permutation__round_out[859]) );
  XOR2_X2 _f_permutation__round__U3307  ( .A(_f_permutation__round__N4039 ), 
        .B(_f_permutation__round__c[726] ), .Z(_f_permutation__round_out[860]) );
  XOR2_X2 _f_permutation__round__U3306  ( .A(_f_permutation__round__N4037 ), 
        .B(_f_permutation__round__c[727] ), .Z(_f_permutation__round_out[861]) );
  XOR2_X2 _f_permutation__round__U3305  ( .A(_f_permutation__round__N4035 ), 
        .B(_f_permutation__round__c[728] ), .Z(_f_permutation__round_out[862]) );
  XOR2_X2 _f_permutation__round__U3304  ( .A(_f_permutation__round__N4033 ), 
        .B(_f_permutation__round__c[729] ), .Z(_f_permutation__round_out[863]) );
  XOR2_X2 _f_permutation__round__U3303  ( .A(_f_permutation__round__N4031 ), 
        .B(_f_permutation__round__c[730] ), .Z(_f_permutation__round_out[864]) );
  XOR2_X2 _f_permutation__round__U3302  ( .A(_f_permutation__round__N4029 ), 
        .B(_f_permutation__round__c[731] ), .Z(_f_permutation__round_out[865]) );
  XOR2_X2 _f_permutation__round__U3301  ( .A(_f_permutation__round__N4027 ), 
        .B(_f_permutation__round__c[732] ), .Z(_f_permutation__round_out[866]) );
  XOR2_X2 _f_permutation__round__U3300  ( .A(_f_permutation__round__N4025 ), 
        .B(_f_permutation__round__c[733] ), .Z(_f_permutation__round_out[867]) );
  XOR2_X2 _f_permutation__round__U3299  ( .A(_f_permutation__round__N4023 ), 
        .B(_f_permutation__round__c[734] ), .Z(_f_permutation__round_out[868]) );
  XOR2_X2 _f_permutation__round__U3298  ( .A(_f_permutation__round__N4021 ), 
        .B(_f_permutation__round__c[735] ), .Z(_f_permutation__round_out[869]) );
  XOR2_X2 _f_permutation__round__U3297  ( .A(_f_permutation__round__N4019 ), 
        .B(_f_permutation__round__c[736] ), .Z(_f_permutation__round_out[870]) );
  XOR2_X2 _f_permutation__round__U3296  ( .A(_f_permutation__round__N4017 ), 
        .B(_f_permutation__round__c[737] ), .Z(_f_permutation__round_out[871]) );
  XOR2_X2 _f_permutation__round__U3295  ( .A(_f_permutation__round__N4015 ), 
        .B(_f_permutation__round__c[738] ), .Z(_f_permutation__round_out[872]) );
  XOR2_X2 _f_permutation__round__U3294  ( .A(_f_permutation__round__N4013 ), 
        .B(_f_permutation__round__c[739] ), .Z(_f_permutation__round_out[873]) );
  XOR2_X2 _f_permutation__round__U3293  ( .A(_f_permutation__round__N4011 ), 
        .B(_f_permutation__round__c[740] ), .Z(_f_permutation__round_out[874]) );
  XOR2_X2 _f_permutation__round__U3292  ( .A(_f_permutation__round__N4009 ), 
        .B(_f_permutation__round__c[741] ), .Z(_f_permutation__round_out[875]) );
  XOR2_X2 _f_permutation__round__U3291  ( .A(_f_permutation__round__N4007 ), 
        .B(_f_permutation__round__c[742] ), .Z(_f_permutation__round_out[876]) );
  XOR2_X2 _f_permutation__round__U3290  ( .A(_f_permutation__round__N4005 ), 
        .B(_f_permutation__round__c[743] ), .Z(_f_permutation__round_out[877]) );
  XOR2_X2 _f_permutation__round__U3289  ( .A(_f_permutation__round__N4003 ), 
        .B(_f_permutation__round__c[744] ), .Z(_f_permutation__round_out[878]) );
  XOR2_X2 _f_permutation__round__U3288  ( .A(_f_permutation__round__N4001 ), 
        .B(_f_permutation__round__c[745] ), .Z(_f_permutation__round_out[879]) );
  XOR2_X2 _f_permutation__round__U3287  ( .A(_f_permutation__round__N3999 ), 
        .B(_f_permutation__round__c[746] ), .Z(_f_permutation__round_out[880]) );
  XOR2_X2 _f_permutation__round__U3286  ( .A(_f_permutation__round__N3997 ), 
        .B(_f_permutation__round__c[747] ), .Z(_f_permutation__round_out[881]) );
  XOR2_X2 _f_permutation__round__U3285  ( .A(_f_permutation__round__N3995 ), 
        .B(_f_permutation__round__c[748] ), .Z(_f_permutation__round_out[882]) );
  XOR2_X2 _f_permutation__round__U3284  ( .A(_f_permutation__round__N3993 ), 
        .B(_f_permutation__round__c[749] ), .Z(_f_permutation__round_out[883]) );
  XOR2_X2 _f_permutation__round__U3283  ( .A(_f_permutation__round__N3991 ), 
        .B(_f_permutation__round__c[750] ), .Z(_f_permutation__round_out[884]) );
  XOR2_X2 _f_permutation__round__U3282  ( .A(_f_permutation__round__N3989 ), 
        .B(_f_permutation__round__c[751] ), .Z(_f_permutation__round_out[885]) );
  XOR2_X2 _f_permutation__round__U3281  ( .A(_f_permutation__round__N3987 ), 
        .B(_f_permutation__round__c[752] ), .Z(_f_permutation__round_out[886]) );
  XOR2_X2 _f_permutation__round__U3280  ( .A(_f_permutation__round__N3985 ), 
        .B(_f_permutation__round__c[753] ), .Z(_f_permutation__round_out[887]) );
  XOR2_X2 _f_permutation__round__U3279  ( .A(_f_permutation__round__N3983 ), 
        .B(_f_permutation__round__c[754] ), .Z(_f_permutation__round_out[888]) );
  XOR2_X2 _f_permutation__round__U3278  ( .A(_f_permutation__round__N3981 ), 
        .B(_f_permutation__round__c[755] ), .Z(_f_permutation__round_out[889]) );
  XOR2_X2 _f_permutation__round__U3277  ( .A(_f_permutation__round__N3979 ), 
        .B(_f_permutation__round__c[756] ), .Z(_f_permutation__round_out[890]) );
  XOR2_X2 _f_permutation__round__U3276  ( .A(_f_permutation__round__N3977 ), 
        .B(_f_permutation__round__c[757] ), .Z(_f_permutation__round_out[891]) );
  XOR2_X2 _f_permutation__round__U3275  ( .A(_f_permutation__round__N3975 ), 
        .B(_f_permutation__round__c[758] ), .Z(_f_permutation__round_out[892]) );
  XOR2_X2 _f_permutation__round__U3274  ( .A(_f_permutation__round__N3973 ), 
        .B(_f_permutation__round__c[759] ), .Z(_f_permutation__round_out[893]) );
  XOR2_X2 _f_permutation__round__U3273  ( .A(_f_permutation__round__N3971 ), 
        .B(_f_permutation__round__c[760] ), .Z(_f_permutation__round_out[894]) );
  XOR2_X2 _f_permutation__round__U3272  ( .A(_f_permutation__round__N3969 ), 
        .B(_f_permutation__round__c[761] ), .Z(_f_permutation__round_out[895]) );
  XOR2_X2 _f_permutation__round__U3271  ( .A(_f_permutation__round__N3967 ), 
        .B(_f_permutation__round__c[383] ), .Z(_f_permutation__round_out[896]) );
  XOR2_X2 _f_permutation__round__U3270  ( .A(_f_permutation__round__N3965 ), 
        .B(_f_permutation__round__c[320] ), .Z(_f_permutation__round_out[897]) );
  XOR2_X2 _f_permutation__round__U3269  ( .A(_f_permutation__round__N3963 ), 
        .B(_f_permutation__round__c[321] ), .Z(_f_permutation__round_out[898]) );
  XOR2_X2 _f_permutation__round__U3268  ( .A(_f_permutation__round__N3961 ), 
        .B(_f_permutation__round__c[322] ), .Z(_f_permutation__round_out[899]) );
  XOR2_X2 _f_permutation__round__U3267  ( .A(_f_permutation__round__N3959 ), 
        .B(_f_permutation__round__c[323] ), .Z(_f_permutation__round_out[900]) );
  XOR2_X2 _f_permutation__round__U3266  ( .A(_f_permutation__round__N3957 ), 
        .B(_f_permutation__round__c[324] ), .Z(_f_permutation__round_out[901]) );
  XOR2_X2 _f_permutation__round__U3265  ( .A(_f_permutation__round__N3955 ), 
        .B(_f_permutation__round__c[325] ), .Z(_f_permutation__round_out[902]) );
  XOR2_X2 _f_permutation__round__U3264  ( .A(_f_permutation__round__N3953 ), 
        .B(_f_permutation__round__c[326] ), .Z(_f_permutation__round_out[903]) );
  XOR2_X2 _f_permutation__round__U3263  ( .A(_f_permutation__round__N3951 ), 
        .B(_f_permutation__round__c[327] ), .Z(_f_permutation__round_out[904]) );
  XOR2_X2 _f_permutation__round__U3262  ( .A(_f_permutation__round__N3949 ), 
        .B(_f_permutation__round__c[328] ), .Z(_f_permutation__round_out[905]) );
  XOR2_X2 _f_permutation__round__U3261  ( .A(_f_permutation__round__N3947 ), 
        .B(_f_permutation__round__c[329] ), .Z(_f_permutation__round_out[906]) );
  XOR2_X2 _f_permutation__round__U3260  ( .A(_f_permutation__round__N3945 ), 
        .B(_f_permutation__round__c[330] ), .Z(_f_permutation__round_out[907]) );
  XOR2_X2 _f_permutation__round__U3259  ( .A(_f_permutation__round__N3943 ), 
        .B(_f_permutation__round__c[331] ), .Z(_f_permutation__round_out[908]) );
  XOR2_X2 _f_permutation__round__U3258  ( .A(_f_permutation__round__N3941 ), 
        .B(_f_permutation__round__c[332] ), .Z(_f_permutation__round_out[909]) );
  XOR2_X2 _f_permutation__round__U3257  ( .A(_f_permutation__round__N3939 ), 
        .B(_f_permutation__round__c[333] ), .Z(_f_permutation__round_out[910]) );
  XOR2_X2 _f_permutation__round__U3256  ( .A(_f_permutation__round__N3937 ), 
        .B(_f_permutation__round__c[334] ), .Z(_f_permutation__round_out[911]) );
  XOR2_X2 _f_permutation__round__U3255  ( .A(_f_permutation__round__N3935 ), 
        .B(_f_permutation__round__c[335] ), .Z(_f_permutation__round_out[912]) );
  XOR2_X2 _f_permutation__round__U3254  ( .A(_f_permutation__round__N3933 ), 
        .B(_f_permutation__round__c[336] ), .Z(_f_permutation__round_out[913]) );
  XOR2_X2 _f_permutation__round__U3253  ( .A(_f_permutation__round__N3931 ), 
        .B(_f_permutation__round__c[337] ), .Z(_f_permutation__round_out[914]) );
  XOR2_X2 _f_permutation__round__U3252  ( .A(_f_permutation__round__N3929 ), 
        .B(_f_permutation__round__c[338] ), .Z(_f_permutation__round_out[915]) );
  XOR2_X2 _f_permutation__round__U3251  ( .A(_f_permutation__round__N3927 ), 
        .B(_f_permutation__round__c[339] ), .Z(_f_permutation__round_out[916]) );
  XOR2_X2 _f_permutation__round__U3250  ( .A(_f_permutation__round__N3925 ), 
        .B(_f_permutation__round__c[340] ), .Z(_f_permutation__round_out[917]) );
  XOR2_X2 _f_permutation__round__U3249  ( .A(_f_permutation__round__N3923 ), 
        .B(_f_permutation__round__c[341] ), .Z(_f_permutation__round_out[918]) );
  XOR2_X2 _f_permutation__round__U3248  ( .A(_f_permutation__round__N3921 ), 
        .B(_f_permutation__round__c[342] ), .Z(_f_permutation__round_out[919]) );
  XOR2_X2 _f_permutation__round__U3247  ( .A(_f_permutation__round__N3919 ), 
        .B(_f_permutation__round__c[343] ), .Z(_f_permutation__round_out[920]) );
  XOR2_X2 _f_permutation__round__U3246  ( .A(_f_permutation__round__N3917 ), 
        .B(_f_permutation__round__c[344] ), .Z(_f_permutation__round_out[921]) );
  XOR2_X2 _f_permutation__round__U3245  ( .A(_f_permutation__round__N3915 ), 
        .B(_f_permutation__round__c[345] ), .Z(_f_permutation__round_out[922]) );
  XOR2_X2 _f_permutation__round__U3244  ( .A(_f_permutation__round__N3913 ), 
        .B(_f_permutation__round__c[346] ), .Z(_f_permutation__round_out[923]) );
  XOR2_X2 _f_permutation__round__U3243  ( .A(_f_permutation__round__N3911 ), 
        .B(_f_permutation__round__c[347] ), .Z(_f_permutation__round_out[924]) );
  XOR2_X2 _f_permutation__round__U3242  ( .A(_f_permutation__round__N3909 ), 
        .B(_f_permutation__round__c[348] ), .Z(_f_permutation__round_out[925]) );
  XOR2_X2 _f_permutation__round__U3241  ( .A(_f_permutation__round__N3907 ), 
        .B(_f_permutation__round__c[349] ), .Z(_f_permutation__round_out[926]) );
  XOR2_X2 _f_permutation__round__U3240  ( .A(_f_permutation__round__N3905 ), 
        .B(_f_permutation__round__c[350] ), .Z(_f_permutation__round_out[927]) );
  XOR2_X2 _f_permutation__round__U3239  ( .A(_f_permutation__round__N3903 ), 
        .B(_f_permutation__round__c[351] ), .Z(_f_permutation__round_out[928]) );
  XOR2_X2 _f_permutation__round__U3238  ( .A(_f_permutation__round__N3901 ), 
        .B(_f_permutation__round__c[352] ), .Z(_f_permutation__round_out[929]) );
  XOR2_X2 _f_permutation__round__U3237  ( .A(_f_permutation__round__N3899 ), 
        .B(_f_permutation__round__c[353] ), .Z(_f_permutation__round_out[930]) );
  XOR2_X2 _f_permutation__round__U3236  ( .A(_f_permutation__round__N3897 ), 
        .B(_f_permutation__round__c[354] ), .Z(_f_permutation__round_out[931]) );
  XOR2_X2 _f_permutation__round__U3235  ( .A(_f_permutation__round__N3895 ), 
        .B(_f_permutation__round__c[355] ), .Z(_f_permutation__round_out[932]) );
  XOR2_X2 _f_permutation__round__U3234  ( .A(_f_permutation__round__N3893 ), 
        .B(_f_permutation__round__c[356] ), .Z(_f_permutation__round_out[933]) );
  XOR2_X2 _f_permutation__round__U3233  ( .A(_f_permutation__round__N3891 ), 
        .B(_f_permutation__round__c[357] ), .Z(_f_permutation__round_out[934]) );
  XOR2_X2 _f_permutation__round__U3232  ( .A(_f_permutation__round__N3889 ), 
        .B(_f_permutation__round__c[358] ), .Z(_f_permutation__round_out[935]) );
  XOR2_X2 _f_permutation__round__U3231  ( .A(_f_permutation__round__N3887 ), 
        .B(_f_permutation__round__c[359] ), .Z(_f_permutation__round_out[936]) );
  XOR2_X2 _f_permutation__round__U3230  ( .A(_f_permutation__round__N3885 ), 
        .B(_f_permutation__round__c[360] ), .Z(_f_permutation__round_out[937]) );
  XOR2_X2 _f_permutation__round__U3229  ( .A(_f_permutation__round__N3883 ), 
        .B(_f_permutation__round__c[361] ), .Z(_f_permutation__round_out[938]) );
  XOR2_X2 _f_permutation__round__U3228  ( .A(_f_permutation__round__N3881 ), 
        .B(_f_permutation__round__c[362] ), .Z(_f_permutation__round_out[939]) );
  XOR2_X2 _f_permutation__round__U3227  ( .A(_f_permutation__round__N3879 ), 
        .B(_f_permutation__round__c[363] ), .Z(_f_permutation__round_out[940]) );
  XOR2_X2 _f_permutation__round__U3226  ( .A(_f_permutation__round__N3877 ), 
        .B(_f_permutation__round__c[364] ), .Z(_f_permutation__round_out[941]) );
  XOR2_X2 _f_permutation__round__U3225  ( .A(_f_permutation__round__N3875 ), 
        .B(_f_permutation__round__c[365] ), .Z(_f_permutation__round_out[942]) );
  XOR2_X2 _f_permutation__round__U3224  ( .A(_f_permutation__round__N3873 ), 
        .B(_f_permutation__round__c[366] ), .Z(_f_permutation__round_out[943]) );
  XOR2_X2 _f_permutation__round__U3223  ( .A(_f_permutation__round__N3871 ), 
        .B(_f_permutation__round__c[367] ), .Z(_f_permutation__round_out[944]) );
  XOR2_X2 _f_permutation__round__U3222  ( .A(_f_permutation__round__N3869 ), 
        .B(_f_permutation__round__c[368] ), .Z(_f_permutation__round_out[945]) );
  XOR2_X2 _f_permutation__round__U3221  ( .A(_f_permutation__round__N3867 ), 
        .B(_f_permutation__round__c[369] ), .Z(_f_permutation__round_out[946]) );
  XOR2_X2 _f_permutation__round__U3220  ( .A(_f_permutation__round__N3865 ), 
        .B(_f_permutation__round__c[370] ), .Z(_f_permutation__round_out[947]) );
  XOR2_X2 _f_permutation__round__U3219  ( .A(_f_permutation__round__N3863 ), 
        .B(_f_permutation__round__c[371] ), .Z(_f_permutation__round_out[948]) );
  XOR2_X2 _f_permutation__round__U3218  ( .A(_f_permutation__round__N3861 ), 
        .B(_f_permutation__round__c[372] ), .Z(_f_permutation__round_out[949]) );
  XOR2_X2 _f_permutation__round__U3217  ( .A(_f_permutation__round__N3859 ), 
        .B(_f_permutation__round__c[373] ), .Z(_f_permutation__round_out[950]) );
  XOR2_X2 _f_permutation__round__U3216  ( .A(_f_permutation__round__N3857 ), 
        .B(_f_permutation__round__c[374] ), .Z(_f_permutation__round_out[951]) );
  XOR2_X2 _f_permutation__round__U3215  ( .A(_f_permutation__round__N3855 ), 
        .B(_f_permutation__round__c[375] ), .Z(_f_permutation__round_out[952]) );
  XOR2_X2 _f_permutation__round__U3214  ( .A(_f_permutation__round__N3853 ), 
        .B(_f_permutation__round__c[376] ), .Z(_f_permutation__round_out[953]) );
  XOR2_X2 _f_permutation__round__U3213  ( .A(_f_permutation__round__N3851 ), 
        .B(_f_permutation__round__c[377] ), .Z(_f_permutation__round_out[954]) );
  XOR2_X2 _f_permutation__round__U3212  ( .A(_f_permutation__round__N3849 ), 
        .B(_f_permutation__round__c[378] ), .Z(_f_permutation__round_out[955]) );
  XOR2_X2 _f_permutation__round__U3211  ( .A(_f_permutation__round__N3847 ), 
        .B(_f_permutation__round__c[379] ), .Z(_f_permutation__round_out[956]) );
  XOR2_X2 _f_permutation__round__U3210  ( .A(_f_permutation__round__N3845 ), 
        .B(_f_permutation__round__c[380] ), .Z(_f_permutation__round_out[957]) );
  XOR2_X2 _f_permutation__round__U3209  ( .A(_f_permutation__round__N3843 ), 
        .B(_f_permutation__round__c[381] ), .Z(_f_permutation__round_out[958]) );
  XOR2_X2 _f_permutation__round__U3208  ( .A(_f_permutation__round__N3841 ), 
        .B(_f_permutation__round__c[382] ), .Z(_f_permutation__round_out[959]) );
  XOR2_X2 _f_permutation__round__U3207  ( .A(_f_permutation__round__N3839 ), 
        .B(_f_permutation__round__c[899] ), .Z(_f_permutation__round_out[960]) );
  XOR2_X2 _f_permutation__round__U3206  ( .A(_f_permutation__round__N3837 ), 
        .B(_f_permutation__round__c[900] ), .Z(_f_permutation__round_out[961]) );
  XOR2_X2 _f_permutation__round__U3205  ( .A(_f_permutation__round__N3835 ), 
        .B(_f_permutation__round__c[901] ), .Z(_f_permutation__round_out[962]) );
  XOR2_X2 _f_permutation__round__U3204  ( .A(_f_permutation__round__N3833 ), 
        .B(_f_permutation__round__c[902] ), .Z(_f_permutation__round_out[963]) );
  XOR2_X2 _f_permutation__round__U3203  ( .A(_f_permutation__round__N3831 ), 
        .B(_f_permutation__round__c[903] ), .Z(_f_permutation__round_out[964]) );
  XOR2_X2 _f_permutation__round__U3202  ( .A(_f_permutation__round__N3829 ), 
        .B(_f_permutation__round__c[904] ), .Z(_f_permutation__round_out[965]) );
  XOR2_X2 _f_permutation__round__U3201  ( .A(_f_permutation__round__N3827 ), 
        .B(_f_permutation__round__c[905] ), .Z(_f_permutation__round_out[966]) );
  XOR2_X2 _f_permutation__round__U3200  ( .A(_f_permutation__round__N3825 ), 
        .B(_f_permutation__round__c[906] ), .Z(_f_permutation__round_out[967]) );
  XOR2_X2 _f_permutation__round__U3199  ( .A(_f_permutation__round__N3823 ), 
        .B(_f_permutation__round__c[907] ), .Z(_f_permutation__round_out[968]) );
  XOR2_X2 _f_permutation__round__U3198  ( .A(_f_permutation__round__N3821 ), 
        .B(_f_permutation__round__c[908] ), .Z(_f_permutation__round_out[969]) );
  XOR2_X2 _f_permutation__round__U3197  ( .A(_f_permutation__round__N3819 ), 
        .B(_f_permutation__round__c[909] ), .Z(_f_permutation__round_out[970]) );
  XOR2_X2 _f_permutation__round__U3196  ( .A(_f_permutation__round__N3817 ), 
        .B(_f_permutation__round__c[910] ), .Z(_f_permutation__round_out[971]) );
  XOR2_X2 _f_permutation__round__U3195  ( .A(_f_permutation__round__N3815 ), 
        .B(_f_permutation__round__c[911] ), .Z(_f_permutation__round_out[972]) );
  XOR2_X2 _f_permutation__round__U3194  ( .A(_f_permutation__round__N3813 ), 
        .B(_f_permutation__round__c[912] ), .Z(_f_permutation__round_out[973]) );
  XOR2_X2 _f_permutation__round__U3193  ( .A(_f_permutation__round__N3811 ), 
        .B(_f_permutation__round__c[913] ), .Z(_f_permutation__round_out[974]) );
  XOR2_X2 _f_permutation__round__U3192  ( .A(_f_permutation__round__N3809 ), 
        .B(_f_permutation__round__c[914] ), .Z(_f_permutation__round_out[975]) );
  XOR2_X2 _f_permutation__round__U3191  ( .A(_f_permutation__round__N3807 ), 
        .B(_f_permutation__round__c[915] ), .Z(_f_permutation__round_out[976]) );
  XOR2_X2 _f_permutation__round__U3190  ( .A(_f_permutation__round__N3805 ), 
        .B(_f_permutation__round__c[916] ), .Z(_f_permutation__round_out[977]) );
  XOR2_X2 _f_permutation__round__U3189  ( .A(_f_permutation__round__N3803 ), 
        .B(_f_permutation__round__c[917] ), .Z(_f_permutation__round_out[978]) );
  XOR2_X2 _f_permutation__round__U3188  ( .A(_f_permutation__round__N3801 ), 
        .B(_f_permutation__round__c[918] ), .Z(_f_permutation__round_out[979]) );
  XOR2_X2 _f_permutation__round__U3187  ( .A(_f_permutation__round__N3799 ), 
        .B(_f_permutation__round__c[919] ), .Z(_f_permutation__round_out[980]) );
  XOR2_X2 _f_permutation__round__U3186  ( .A(_f_permutation__round__N3797 ), 
        .B(_f_permutation__round__c[920] ), .Z(_f_permutation__round_out[981]) );
  XOR2_X2 _f_permutation__round__U3185  ( .A(_f_permutation__round__N3795 ), 
        .B(_f_permutation__round__c[921] ), .Z(_f_permutation__round_out[982]) );
  XOR2_X2 _f_permutation__round__U3184  ( .A(_f_permutation__round__N3793 ), 
        .B(_f_permutation__round__c[922] ), .Z(_f_permutation__round_out[983]) );
  XOR2_X2 _f_permutation__round__U3183  ( .A(_f_permutation__round__N3791 ), 
        .B(_f_permutation__round__c[923] ), .Z(_f_permutation__round_out[984]) );
  XOR2_X2 _f_permutation__round__U3182  ( .A(_f_permutation__round__N3789 ), 
        .B(_f_permutation__round__c[924] ), .Z(_f_permutation__round_out[985]) );
  XOR2_X2 _f_permutation__round__U3181  ( .A(_f_permutation__round__N3787 ), 
        .B(_f_permutation__round__c[925] ), .Z(_f_permutation__round_out[986]) );
  XOR2_X2 _f_permutation__round__U3180  ( .A(_f_permutation__round__N3785 ), 
        .B(_f_permutation__round__c[926] ), .Z(_f_permutation__round_out[987]) );
  XOR2_X2 _f_permutation__round__U3179  ( .A(_f_permutation__round__N3783 ), 
        .B(_f_permutation__round__c[927] ), .Z(_f_permutation__round_out[988]) );
  XOR2_X2 _f_permutation__round__U3178  ( .A(_f_permutation__round__N3781 ), 
        .B(_f_permutation__round__c[928] ), .Z(_f_permutation__round_out[989]) );
  XOR2_X2 _f_permutation__round__U3177  ( .A(_f_permutation__round__N3779 ), 
        .B(_f_permutation__round__c[929] ), .Z(_f_permutation__round_out[990]) );
  XOR2_X2 _f_permutation__round__U3176  ( .A(_f_permutation__round__N3777 ), 
        .B(_f_permutation__round__c[930] ), .Z(_f_permutation__round_out[991]) );
  XOR2_X2 _f_permutation__round__U3175  ( .A(_f_permutation__round__N3775 ), 
        .B(_f_permutation__round__c[931] ), .Z(_f_permutation__round_out[992]) );
  XOR2_X2 _f_permutation__round__U3174  ( .A(_f_permutation__round__N3773 ), 
        .B(_f_permutation__round__c[932] ), .Z(_f_permutation__round_out[993]) );
  XOR2_X2 _f_permutation__round__U3173  ( .A(_f_permutation__round__N3771 ), 
        .B(_f_permutation__round__c[933] ), .Z(_f_permutation__round_out[994]) );
  XOR2_X2 _f_permutation__round__U3172  ( .A(_f_permutation__round__N3769 ), 
        .B(_f_permutation__round__c[934] ), .Z(_f_permutation__round_out[995]) );
  XOR2_X2 _f_permutation__round__U3171  ( .A(_f_permutation__round__N3767 ), 
        .B(_f_permutation__round__c[935] ), .Z(_f_permutation__round_out[996]) );
  XOR2_X2 _f_permutation__round__U3170  ( .A(_f_permutation__round__N3765 ), 
        .B(_f_permutation__round__c[936] ), .Z(_f_permutation__round_out[997]) );
  XOR2_X2 _f_permutation__round__U3169  ( .A(_f_permutation__round__N3763 ), 
        .B(_f_permutation__round__c[937] ), .Z(_f_permutation__round_out[998]) );
  XOR2_X2 _f_permutation__round__U3168  ( .A(_f_permutation__round__N3761 ), 
        .B(_f_permutation__round__c[938] ), .Z(_f_permutation__round_out[999]) );
  XOR2_X2 _f_permutation__round__U3167  ( .A(_f_permutation__round__N3759 ), 
        .B(_f_permutation__round__c[939] ), .Z(
        _f_permutation__round_out[1000]) );
  XOR2_X2 _f_permutation__round__U3166  ( .A(_f_permutation__round__N3757 ), 
        .B(_f_permutation__round__c[940] ), .Z(
        _f_permutation__round_out[1001]) );
  XOR2_X2 _f_permutation__round__U3165  ( .A(_f_permutation__round__N3755 ), 
        .B(_f_permutation__round__c[941] ), .Z(
        _f_permutation__round_out[1002]) );
  XOR2_X2 _f_permutation__round__U3164  ( .A(_f_permutation__round__N3753 ), 
        .B(_f_permutation__round__c[942] ), .Z(
        _f_permutation__round_out[1003]) );
  XOR2_X2 _f_permutation__round__U3163  ( .A(_f_permutation__round__N3751 ), 
        .B(_f_permutation__round__c[943] ), .Z(
        _f_permutation__round_out[1004]) );
  XOR2_X2 _f_permutation__round__U3162  ( .A(_f_permutation__round__N3749 ), 
        .B(_f_permutation__round__c[944] ), .Z(
        _f_permutation__round_out[1005]) );
  XOR2_X2 _f_permutation__round__U3161  ( .A(_f_permutation__round__N3747 ), 
        .B(_f_permutation__round__c[945] ), .Z(
        _f_permutation__round_out[1006]) );
  XOR2_X2 _f_permutation__round__U3160  ( .A(_f_permutation__round__N3745 ), 
        .B(_f_permutation__round__c[946] ), .Z(
        _f_permutation__round_out[1007]) );
  XOR2_X2 _f_permutation__round__U3159  ( .A(_f_permutation__round__N3743 ), 
        .B(_f_permutation__round__c[947] ), .Z(
        _f_permutation__round_out[1008]) );
  XOR2_X2 _f_permutation__round__U3158  ( .A(_f_permutation__round__N3741 ), 
        .B(_f_permutation__round__c[948] ), .Z(
        _f_permutation__round_out[1009]) );
  XOR2_X2 _f_permutation__round__U3157  ( .A(_f_permutation__round__N3739 ), 
        .B(_f_permutation__round__c[949] ), .Z(
        _f_permutation__round_out[1010]) );
  XOR2_X2 _f_permutation__round__U3156  ( .A(_f_permutation__round__N3737 ), 
        .B(_f_permutation__round__c[950] ), .Z(
        _f_permutation__round_out[1011]) );
  XOR2_X2 _f_permutation__round__U3155  ( .A(_f_permutation__round__N3735 ), 
        .B(_f_permutation__round__c[951] ), .Z(
        _f_permutation__round_out[1012]) );
  XOR2_X2 _f_permutation__round__U3154  ( .A(_f_permutation__round__N3733 ), 
        .B(_f_permutation__round__c[952] ), .Z(
        _f_permutation__round_out[1013]) );
  XOR2_X2 _f_permutation__round__U3153  ( .A(_f_permutation__round__N3731 ), 
        .B(_f_permutation__round__c[953] ), .Z(
        _f_permutation__round_out[1014]) );
  XOR2_X2 _f_permutation__round__U3152  ( .A(_f_permutation__round__N3729 ), 
        .B(_f_permutation__round__c[954] ), .Z(
        _f_permutation__round_out[1015]) );
  XOR2_X2 _f_permutation__round__U3151  ( .A(_f_permutation__round__N3727 ), 
        .B(_f_permutation__round__c[955] ), .Z(
        _f_permutation__round_out[1016]) );
  XOR2_X2 _f_permutation__round__U3150  ( .A(_f_permutation__round__N3725 ), 
        .B(_f_permutation__round__c[956] ), .Z(
        _f_permutation__round_out[1017]) );
  XOR2_X2 _f_permutation__round__U3149  ( .A(_f_permutation__round__N3723 ), 
        .B(_f_permutation__round__c[957] ), .Z(
        _f_permutation__round_out[1018]) );
  XOR2_X2 _f_permutation__round__U3148  ( .A(_f_permutation__round__N3721 ), 
        .B(_f_permutation__round__c[958] ), .Z(
        _f_permutation__round_out[1019]) );
  XOR2_X2 _f_permutation__round__U3147  ( .A(_f_permutation__round__N3719 ), 
        .B(_f_permutation__round__c[959] ), .Z(
        _f_permutation__round_out[1020]) );
  XOR2_X2 _f_permutation__round__U3146  ( .A(_f_permutation__round__N3717 ), 
        .B(_f_permutation__round__c[896] ), .Z(
        _f_permutation__round_out[1021]) );
  XOR2_X2 _f_permutation__round__U3145  ( .A(_f_permutation__round__N3715 ), 
        .B(_f_permutation__round__c[897] ), .Z(
        _f_permutation__round_out[1022]) );
  XOR2_X2 _f_permutation__round__U3144  ( .A(_f_permutation__round__N3713 ), 
        .B(_f_permutation__round__c[898] ), .Z(
        _f_permutation__round_out[1023]) );
  XOR2_X2 _f_permutation__round__U3143  ( .A(_f_permutation__round__N3711 ), 
        .B(_f_permutation__round__c[531] ), .Z(
        _f_permutation__round_out[1024]) );
  XOR2_X2 _f_permutation__round__U3142  ( .A(_f_permutation__round__N3709 ), 
        .B(_f_permutation__round__c[532] ), .Z(
        _f_permutation__round_out[1025]) );
  XOR2_X2 _f_permutation__round__U3141  ( .A(_f_permutation__round__N3707 ), 
        .B(_f_permutation__round__c[533] ), .Z(
        _f_permutation__round_out[1026]) );
  XOR2_X2 _f_permutation__round__U3140  ( .A(_f_permutation__round__N3705 ), 
        .B(_f_permutation__round__c[534] ), .Z(
        _f_permutation__round_out[1027]) );
  XOR2_X2 _f_permutation__round__U3139  ( .A(_f_permutation__round__N3703 ), 
        .B(_f_permutation__round__c[535] ), .Z(
        _f_permutation__round_out[1028]) );
  XOR2_X2 _f_permutation__round__U3138  ( .A(_f_permutation__round__N3701 ), 
        .B(_f_permutation__round__c[536] ), .Z(
        _f_permutation__round_out[1029]) );
  XOR2_X2 _f_permutation__round__U3137  ( .A(_f_permutation__round__N3699 ), 
        .B(_f_permutation__round__c[537] ), .Z(
        _f_permutation__round_out[1030]) );
  XOR2_X2 _f_permutation__round__U3136  ( .A(_f_permutation__round__N3697 ), 
        .B(_f_permutation__round__c[538] ), .Z(
        _f_permutation__round_out[1031]) );
  XOR2_X2 _f_permutation__round__U3135  ( .A(_f_permutation__round__N3695 ), 
        .B(_f_permutation__round__c[539] ), .Z(
        _f_permutation__round_out[1032]) );
  XOR2_X2 _f_permutation__round__U3134  ( .A(_f_permutation__round__N3693 ), 
        .B(_f_permutation__round__c[540] ), .Z(
        _f_permutation__round_out[1033]) );
  XOR2_X2 _f_permutation__round__U3133  ( .A(_f_permutation__round__N3691 ), 
        .B(_f_permutation__round__c[541] ), .Z(
        _f_permutation__round_out[1034]) );
  XOR2_X2 _f_permutation__round__U3132  ( .A(_f_permutation__round__N3689 ), 
        .B(_f_permutation__round__c[542] ), .Z(
        _f_permutation__round_out[1035]) );
  XOR2_X2 _f_permutation__round__U3131  ( .A(_f_permutation__round__N3687 ), 
        .B(_f_permutation__round__c[543] ), .Z(
        _f_permutation__round_out[1036]) );
  XOR2_X2 _f_permutation__round__U3130  ( .A(_f_permutation__round__N3685 ), 
        .B(_f_permutation__round__c[544] ), .Z(
        _f_permutation__round_out[1037]) );
  XOR2_X2 _f_permutation__round__U3129  ( .A(_f_permutation__round__N3683 ), 
        .B(_f_permutation__round__c[545] ), .Z(
        _f_permutation__round_out[1038]) );
  XOR2_X2 _f_permutation__round__U3128  ( .A(_f_permutation__round__N3681 ), 
        .B(_f_permutation__round__c[546] ), .Z(
        _f_permutation__round_out[1039]) );
  XOR2_X2 _f_permutation__round__U3127  ( .A(_f_permutation__round__N3679 ), 
        .B(_f_permutation__round__c[547] ), .Z(
        _f_permutation__round_out[1040]) );
  XOR2_X2 _f_permutation__round__U3126  ( .A(_f_permutation__round__N3677 ), 
        .B(_f_permutation__round__c[548] ), .Z(
        _f_permutation__round_out[1041]) );
  XOR2_X2 _f_permutation__round__U3125  ( .A(_f_permutation__round__N3675 ), 
        .B(_f_permutation__round__c[549] ), .Z(
        _f_permutation__round_out[1042]) );
  XOR2_X2 _f_permutation__round__U3124  ( .A(_f_permutation__round__N3673 ), 
        .B(_f_permutation__round__c[550] ), .Z(
        _f_permutation__round_out[1043]) );
  XOR2_X2 _f_permutation__round__U3123  ( .A(_f_permutation__round__N3671 ), 
        .B(_f_permutation__round__c[551] ), .Z(
        _f_permutation__round_out[1044]) );
  XOR2_X2 _f_permutation__round__U3122  ( .A(_f_permutation__round__N3669 ), 
        .B(_f_permutation__round__c[552] ), .Z(
        _f_permutation__round_out[1045]) );
  XOR2_X2 _f_permutation__round__U3121  ( .A(_f_permutation__round__N3667 ), 
        .B(_f_permutation__round__c[553] ), .Z(
        _f_permutation__round_out[1046]) );
  XOR2_X2 _f_permutation__round__U3120  ( .A(_f_permutation__round__N3665 ), 
        .B(_f_permutation__round__c[554] ), .Z(
        _f_permutation__round_out[1047]) );
  XOR2_X2 _f_permutation__round__U3119  ( .A(_f_permutation__round__N3663 ), 
        .B(_f_permutation__round__c[555] ), .Z(
        _f_permutation__round_out[1048]) );
  XOR2_X2 _f_permutation__round__U3118  ( .A(_f_permutation__round__N3661 ), 
        .B(_f_permutation__round__c[556] ), .Z(
        _f_permutation__round_out[1049]) );
  XOR2_X2 _f_permutation__round__U3117  ( .A(_f_permutation__round__N3659 ), 
        .B(_f_permutation__round__c[557] ), .Z(
        _f_permutation__round_out[1050]) );
  XOR2_X2 _f_permutation__round__U3116  ( .A(_f_permutation__round__N3657 ), 
        .B(_f_permutation__round__c[558] ), .Z(
        _f_permutation__round_out[1051]) );
  XOR2_X2 _f_permutation__round__U3115  ( .A(_f_permutation__round__N3655 ), 
        .B(_f_permutation__round__c[559] ), .Z(
        _f_permutation__round_out[1052]) );
  XOR2_X2 _f_permutation__round__U3114  ( .A(_f_permutation__round__N3653 ), 
        .B(_f_permutation__round__c[560] ), .Z(
        _f_permutation__round_out[1053]) );
  XOR2_X2 _f_permutation__round__U3113  ( .A(_f_permutation__round__N3651 ), 
        .B(_f_permutation__round__c[561] ), .Z(
        _f_permutation__round_out[1054]) );
  XOR2_X2 _f_permutation__round__U3112  ( .A(_f_permutation__round__N3649 ), 
        .B(_f_permutation__round__c[562] ), .Z(
        _f_permutation__round_out[1055]) );
  XOR2_X2 _f_permutation__round__U3111  ( .A(_f_permutation__round__N3647 ), 
        .B(_f_permutation__round__c[563] ), .Z(
        _f_permutation__round_out[1056]) );
  XOR2_X2 _f_permutation__round__U3110  ( .A(_f_permutation__round__N3645 ), 
        .B(_f_permutation__round__c[564] ), .Z(
        _f_permutation__round_out[1057]) );
  XOR2_X2 _f_permutation__round__U3109  ( .A(_f_permutation__round__N3643 ), 
        .B(_f_permutation__round__c[565] ), .Z(
        _f_permutation__round_out[1058]) );
  XOR2_X2 _f_permutation__round__U3108  ( .A(_f_permutation__round__N3641 ), 
        .B(_f_permutation__round__c[566] ), .Z(
        _f_permutation__round_out[1059]) );
  XOR2_X2 _f_permutation__round__U3107  ( .A(_f_permutation__round__N3639 ), 
        .B(_f_permutation__round__c[567] ), .Z(
        _f_permutation__round_out[1060]) );
  XOR2_X2 _f_permutation__round__U3106  ( .A(_f_permutation__round__N3637 ), 
        .B(_f_permutation__round__c[568] ), .Z(
        _f_permutation__round_out[1061]) );
  XOR2_X2 _f_permutation__round__U3105  ( .A(_f_permutation__round__N3635 ), 
        .B(_f_permutation__round__c[569] ), .Z(
        _f_permutation__round_out[1062]) );
  XOR2_X2 _f_permutation__round__U3104  ( .A(_f_permutation__round__N3633 ), 
        .B(_f_permutation__round__c[570] ), .Z(
        _f_permutation__round_out[1063]) );
  XOR2_X2 _f_permutation__round__U3103  ( .A(_f_permutation__round__N3631 ), 
        .B(_f_permutation__round__c[571] ), .Z(
        _f_permutation__round_out[1064]) );
  XOR2_X2 _f_permutation__round__U3102  ( .A(_f_permutation__round__N3629 ), 
        .B(_f_permutation__round__c[572] ), .Z(
        _f_permutation__round_out[1065]) );
  XOR2_X2 _f_permutation__round__U3101  ( .A(_f_permutation__round__N3627 ), 
        .B(_f_permutation__round__c[573] ), .Z(
        _f_permutation__round_out[1066]) );
  XOR2_X2 _f_permutation__round__U3100  ( .A(_f_permutation__round__N3625 ), 
        .B(_f_permutation__round__c[574] ), .Z(
        _f_permutation__round_out[1067]) );
  XOR2_X2 _f_permutation__round__U3099  ( .A(_f_permutation__round__N3623 ), 
        .B(_f_permutation__round__c[575] ), .Z(
        _f_permutation__round_out[1068]) );
  XOR2_X2 _f_permutation__round__U3098  ( .A(_f_permutation__round__N3621 ), 
        .B(_f_permutation__round__c[512] ), .Z(
        _f_permutation__round_out[1069]) );
  XOR2_X2 _f_permutation__round__U3097  ( .A(_f_permutation__round__N3619 ), 
        .B(_f_permutation__round__c[513] ), .Z(
        _f_permutation__round_out[1070]) );
  XOR2_X2 _f_permutation__round__U3096  ( .A(_f_permutation__round__N3617 ), 
        .B(_f_permutation__round__c[514] ), .Z(
        _f_permutation__round_out[1071]) );
  XOR2_X2 _f_permutation__round__U3095  ( .A(_f_permutation__round__N3615 ), 
        .B(_f_permutation__round__c[515] ), .Z(
        _f_permutation__round_out[1072]) );
  XOR2_X2 _f_permutation__round__U3094  ( .A(_f_permutation__round__N3613 ), 
        .B(_f_permutation__round__c[516] ), .Z(
        _f_permutation__round_out[1073]) );
  XOR2_X2 _f_permutation__round__U3093  ( .A(_f_permutation__round__N3611 ), 
        .B(_f_permutation__round__c[517] ), .Z(
        _f_permutation__round_out[1074]) );
  XOR2_X2 _f_permutation__round__U3092  ( .A(_f_permutation__round__N3609 ), 
        .B(_f_permutation__round__c[518] ), .Z(
        _f_permutation__round_out[1075]) );
  XOR2_X2 _f_permutation__round__U3091  ( .A(_f_permutation__round__N3607 ), 
        .B(_f_permutation__round__c[519] ), .Z(
        _f_permutation__round_out[1076]) );
  XOR2_X2 _f_permutation__round__U3090  ( .A(_f_permutation__round__N3605 ), 
        .B(_f_permutation__round__c[520] ), .Z(
        _f_permutation__round_out[1077]) );
  XOR2_X2 _f_permutation__round__U3089  ( .A(_f_permutation__round__N3603 ), 
        .B(_f_permutation__round__c[521] ), .Z(
        _f_permutation__round_out[1078]) );
  XOR2_X2 _f_permutation__round__U3088  ( .A(_f_permutation__round__N3601 ), 
        .B(_f_permutation__round__c[522] ), .Z(
        _f_permutation__round_out[1079]) );
  XOR2_X2 _f_permutation__round__U3087  ( .A(_f_permutation__round__N3599 ), 
        .B(_f_permutation__round__c[523] ), .Z(
        _f_permutation__round_out[1080]) );
  XOR2_X2 _f_permutation__round__U3086  ( .A(_f_permutation__round__N3597 ), 
        .B(_f_permutation__round__c[524] ), .Z(
        _f_permutation__round_out[1081]) );
  XOR2_X2 _f_permutation__round__U3085  ( .A(_f_permutation__round__N3595 ), 
        .B(_f_permutation__round__c[525] ), .Z(
        _f_permutation__round_out[1082]) );
  XOR2_X2 _f_permutation__round__U3084  ( .A(_f_permutation__round__N3593 ), 
        .B(_f_permutation__round__c[526] ), .Z(
        _f_permutation__round_out[1083]) );
  XOR2_X2 _f_permutation__round__U3083  ( .A(_f_permutation__round__N3591 ), 
        .B(_f_permutation__round__c[527] ), .Z(
        _f_permutation__round_out[1084]) );
  XOR2_X2 _f_permutation__round__U3082  ( .A(_f_permutation__round__N3589 ), 
        .B(_f_permutation__round__c[528] ), .Z(
        _f_permutation__round_out[1085]) );
  XOR2_X2 _f_permutation__round__U3081  ( .A(_f_permutation__round__N3587 ), 
        .B(_f_permutation__round__c[529] ), .Z(
        _f_permutation__round_out[1086]) );
  XOR2_X2 _f_permutation__round__U3080  ( .A(_f_permutation__round__N3585 ), 
        .B(_f_permutation__round__c[530] ), .Z(
        _f_permutation__round_out[1087]) );
  XOR2_X2 _f_permutation__round__U3079  ( .A(_f_permutation__round__N3583 ), 
        .B(_f_permutation__round__c[189] ), .Z(
        _f_permutation__round_out[1088]) );
  XOR2_X2 _f_permutation__round__U3078  ( .A(_f_permutation__round__N3581 ), 
        .B(_f_permutation__round__c[190] ), .Z(
        _f_permutation__round_out[1089]) );
  XOR2_X2 _f_permutation__round__U3077  ( .A(_f_permutation__round__N3579 ), 
        .B(_f_permutation__round__c[191] ), .Z(
        _f_permutation__round_out[1090]) );
  XOR2_X2 _f_permutation__round__U3076  ( .A(_f_permutation__round__N3577 ), 
        .B(_f_permutation__round__c[128] ), .Z(
        _f_permutation__round_out[1091]) );
  XOR2_X2 _f_permutation__round__U3075  ( .A(_f_permutation__round__N3575 ), 
        .B(_f_permutation__round__c[129] ), .Z(
        _f_permutation__round_out[1092]) );
  XOR2_X2 _f_permutation__round__U3074  ( .A(_f_permutation__round__N3573 ), 
        .B(_f_permutation__round__c[130] ), .Z(
        _f_permutation__round_out[1093]) );
  XOR2_X2 _f_permutation__round__U3073  ( .A(_f_permutation__round__N3571 ), 
        .B(_f_permutation__round__c[131] ), .Z(
        _f_permutation__round_out[1094]) );
  XOR2_X2 _f_permutation__round__U3072  ( .A(_f_permutation__round__N3569 ), 
        .B(_f_permutation__round__c[132] ), .Z(
        _f_permutation__round_out[1095]) );
  XOR2_X2 _f_permutation__round__U3071  ( .A(_f_permutation__round__N3567 ), 
        .B(_f_permutation__round__c[133] ), .Z(
        _f_permutation__round_out[1096]) );
  XOR2_X2 _f_permutation__round__U3070  ( .A(_f_permutation__round__N3565 ), 
        .B(_f_permutation__round__c[134] ), .Z(
        _f_permutation__round_out[1097]) );
  XOR2_X2 _f_permutation__round__U3069  ( .A(_f_permutation__round__N3563 ), 
        .B(_f_permutation__round__c[135] ), .Z(
        _f_permutation__round_out[1098]) );
  XOR2_X2 _f_permutation__round__U3068  ( .A(_f_permutation__round__N3561 ), 
        .B(_f_permutation__round__c[136] ), .Z(
        _f_permutation__round_out[1099]) );
  XOR2_X2 _f_permutation__round__U3067  ( .A(_f_permutation__round__N3559 ), 
        .B(_f_permutation__round__c[137] ), .Z(
        _f_permutation__round_out[1100]) );
  XOR2_X2 _f_permutation__round__U3066  ( .A(_f_permutation__round__N3557 ), 
        .B(_f_permutation__round__c[138] ), .Z(
        _f_permutation__round_out[1101]) );
  XOR2_X2 _f_permutation__round__U3065  ( .A(_f_permutation__round__N3555 ), 
        .B(_f_permutation__round__c[139] ), .Z(
        _f_permutation__round_out[1102]) );
  XOR2_X2 _f_permutation__round__U3064  ( .A(_f_permutation__round__N3553 ), 
        .B(_f_permutation__round__c[140] ), .Z(
        _f_permutation__round_out[1103]) );
  XOR2_X2 _f_permutation__round__U3063  ( .A(_f_permutation__round__N3551 ), 
        .B(_f_permutation__round__c[141] ), .Z(
        _f_permutation__round_out[1104]) );
  XOR2_X2 _f_permutation__round__U3062  ( .A(_f_permutation__round__N3549 ), 
        .B(_f_permutation__round__c[142] ), .Z(
        _f_permutation__round_out[1105]) );
  XOR2_X2 _f_permutation__round__U3061  ( .A(_f_permutation__round__N3547 ), 
        .B(_f_permutation__round__c[143] ), .Z(
        _f_permutation__round_out[1106]) );
  XOR2_X2 _f_permutation__round__U3060  ( .A(_f_permutation__round__N3545 ), 
        .B(_f_permutation__round__c[144] ), .Z(
        _f_permutation__round_out[1107]) );
  XOR2_X2 _f_permutation__round__U3059  ( .A(_f_permutation__round__N3543 ), 
        .B(_f_permutation__round__c[145] ), .Z(
        _f_permutation__round_out[1108]) );
  XOR2_X2 _f_permutation__round__U3058  ( .A(_f_permutation__round__N3541 ), 
        .B(_f_permutation__round__c[146] ), .Z(
        _f_permutation__round_out[1109]) );
  XOR2_X2 _f_permutation__round__U3057  ( .A(_f_permutation__round__N3539 ), 
        .B(_f_permutation__round__c[147] ), .Z(
        _f_permutation__round_out[1110]) );
  XOR2_X2 _f_permutation__round__U3056  ( .A(_f_permutation__round__N3537 ), 
        .B(_f_permutation__round__c[148] ), .Z(
        _f_permutation__round_out[1111]) );
  XOR2_X2 _f_permutation__round__U3055  ( .A(_f_permutation__round__N3535 ), 
        .B(_f_permutation__round__c[149] ), .Z(
        _f_permutation__round_out[1112]) );
  XOR2_X2 _f_permutation__round__U3054  ( .A(_f_permutation__round__N3533 ), 
        .B(_f_permutation__round__c[150] ), .Z(
        _f_permutation__round_out[1113]) );
  XOR2_X2 _f_permutation__round__U3053  ( .A(_f_permutation__round__N3531 ), 
        .B(_f_permutation__round__c[151] ), .Z(
        _f_permutation__round_out[1114]) );
  XOR2_X2 _f_permutation__round__U3052  ( .A(_f_permutation__round__N3529 ), 
        .B(_f_permutation__round__c[152] ), .Z(
        _f_permutation__round_out[1115]) );
  XOR2_X2 _f_permutation__round__U3051  ( .A(_f_permutation__round__N3527 ), 
        .B(_f_permutation__round__c[153] ), .Z(
        _f_permutation__round_out[1116]) );
  XOR2_X2 _f_permutation__round__U3050  ( .A(_f_permutation__round__N3525 ), 
        .B(_f_permutation__round__c[154] ), .Z(
        _f_permutation__round_out[1117]) );
  XOR2_X2 _f_permutation__round__U3049  ( .A(_f_permutation__round__N3523 ), 
        .B(_f_permutation__round__c[155] ), .Z(
        _f_permutation__round_out[1118]) );
  XOR2_X2 _f_permutation__round__U3048  ( .A(_f_permutation__round__N3521 ), 
        .B(_f_permutation__round__c[156] ), .Z(
        _f_permutation__round_out[1119]) );
  XOR2_X2 _f_permutation__round__U3047  ( .A(_f_permutation__round__N3519 ), 
        .B(_f_permutation__round__c[157] ), .Z(
        _f_permutation__round_out[1120]) );
  XOR2_X2 _f_permutation__round__U3046  ( .A(_f_permutation__round__N3517 ), 
        .B(_f_permutation__round__c[158] ), .Z(
        _f_permutation__round_out[1121]) );
  XOR2_X2 _f_permutation__round__U3045  ( .A(_f_permutation__round__N3515 ), 
        .B(_f_permutation__round__c[159] ), .Z(
        _f_permutation__round_out[1122]) );
  XOR2_X2 _f_permutation__round__U3044  ( .A(_f_permutation__round__N3513 ), 
        .B(_f_permutation__round__c[160] ), .Z(
        _f_permutation__round_out[1123]) );
  XOR2_X2 _f_permutation__round__U3043  ( .A(_f_permutation__round__N3511 ), 
        .B(_f_permutation__round__c[161] ), .Z(
        _f_permutation__round_out[1124]) );
  XOR2_X2 _f_permutation__round__U3042  ( .A(_f_permutation__round__N3509 ), 
        .B(_f_permutation__round__c[162] ), .Z(
        _f_permutation__round_out[1125]) );
  XOR2_X2 _f_permutation__round__U3041  ( .A(_f_permutation__round__N3507 ), 
        .B(_f_permutation__round__c[163] ), .Z(
        _f_permutation__round_out[1126]) );
  XOR2_X2 _f_permutation__round__U3040  ( .A(_f_permutation__round__N3505 ), 
        .B(_f_permutation__round__c[164] ), .Z(
        _f_permutation__round_out[1127]) );
  XOR2_X2 _f_permutation__round__U3039  ( .A(_f_permutation__round__N3503 ), 
        .B(_f_permutation__round__c[165] ), .Z(
        _f_permutation__round_out[1128]) );
  XOR2_X2 _f_permutation__round__U3038  ( .A(_f_permutation__round__N3501 ), 
        .B(_f_permutation__round__c[166] ), .Z(
        _f_permutation__round_out[1129]) );
  XOR2_X2 _f_permutation__round__U3037  ( .A(_f_permutation__round__N3499 ), 
        .B(_f_permutation__round__c[167] ), .Z(
        _f_permutation__round_out[1130]) );
  XOR2_X2 _f_permutation__round__U3036  ( .A(_f_permutation__round__N3497 ), 
        .B(_f_permutation__round__c[168] ), .Z(
        _f_permutation__round_out[1131]) );
  XOR2_X2 _f_permutation__round__U3035  ( .A(_f_permutation__round__N3495 ), 
        .B(_f_permutation__round__c[169] ), .Z(
        _f_permutation__round_out[1132]) );
  XOR2_X2 _f_permutation__round__U3034  ( .A(_f_permutation__round__N3493 ), 
        .B(_f_permutation__round__c[170] ), .Z(
        _f_permutation__round_out[1133]) );
  XOR2_X2 _f_permutation__round__U3033  ( .A(_f_permutation__round__N3491 ), 
        .B(_f_permutation__round__c[171] ), .Z(
        _f_permutation__round_out[1134]) );
  XOR2_X2 _f_permutation__round__U3032  ( .A(_f_permutation__round__N3489 ), 
        .B(_f_permutation__round__c[172] ), .Z(
        _f_permutation__round_out[1135]) );
  XOR2_X2 _f_permutation__round__U3031  ( .A(_f_permutation__round__N3487 ), 
        .B(_f_permutation__round__c[173] ), .Z(
        _f_permutation__round_out[1136]) );
  XOR2_X2 _f_permutation__round__U3030  ( .A(_f_permutation__round__N3485 ), 
        .B(_f_permutation__round__c[174] ), .Z(
        _f_permutation__round_out[1137]) );
  XOR2_X2 _f_permutation__round__U3029  ( .A(_f_permutation__round__N3483 ), 
        .B(_f_permutation__round__c[175] ), .Z(
        _f_permutation__round_out[1138]) );
  XOR2_X2 _f_permutation__round__U3028  ( .A(_f_permutation__round__N3481 ), 
        .B(_f_permutation__round__c[176] ), .Z(
        _f_permutation__round_out[1139]) );
  XOR2_X2 _f_permutation__round__U3027  ( .A(_f_permutation__round__N3479 ), 
        .B(_f_permutation__round__c[177] ), .Z(
        _f_permutation__round_out[1140]) );
  XOR2_X2 _f_permutation__round__U3026  ( .A(_f_permutation__round__N3477 ), 
        .B(_f_permutation__round__c[178] ), .Z(
        _f_permutation__round_out[1141]) );
  XOR2_X2 _f_permutation__round__U3025  ( .A(_f_permutation__round__N3475 ), 
        .B(_f_permutation__round__c[179] ), .Z(
        _f_permutation__round_out[1142]) );
  XOR2_X2 _f_permutation__round__U3024  ( .A(_f_permutation__round__N3473 ), 
        .B(_f_permutation__round__c[180] ), .Z(
        _f_permutation__round_out[1143]) );
  XOR2_X2 _f_permutation__round__U3023  ( .A(_f_permutation__round__N3471 ), 
        .B(_f_permutation__round__c[181] ), .Z(
        _f_permutation__round_out[1144]) );
  XOR2_X2 _f_permutation__round__U3022  ( .A(_f_permutation__round__N3469 ), 
        .B(_f_permutation__round__c[182] ), .Z(
        _f_permutation__round_out[1145]) );
  XOR2_X2 _f_permutation__round__U3021  ( .A(_f_permutation__round__N3467 ), 
        .B(_f_permutation__round__c[183] ), .Z(
        _f_permutation__round_out[1146]) );
  XOR2_X2 _f_permutation__round__U3020  ( .A(_f_permutation__round__N3465 ), 
        .B(_f_permutation__round__c[184] ), .Z(
        _f_permutation__round_out[1147]) );
  XOR2_X2 _f_permutation__round__U3019  ( .A(_f_permutation__round__N3463 ), 
        .B(_f_permutation__round__c[185] ), .Z(
        _f_permutation__round_out[1148]) );
  XOR2_X2 _f_permutation__round__U3018  ( .A(_f_permutation__round__N3461 ), 
        .B(_f_permutation__round__c[186] ), .Z(
        _f_permutation__round_out[1149]) );
  XOR2_X2 _f_permutation__round__U3017  ( .A(_f_permutation__round__N3459 ), 
        .B(_f_permutation__round__c[187] ), .Z(
        _f_permutation__round_out[1150]) );
  XOR2_X2 _f_permutation__round__U3016  ( .A(_f_permutation__round__N3457 ), 
        .B(_f_permutation__round__c[188] ), .Z(
        _f_permutation__round_out[1151]) );
  XOR2_X2 _f_permutation__round__U3015  ( .A(_f_permutation__round__N3455 ), 
        .B(_f_permutation__round__c[1388] ), .Z(
        _f_permutation__round_out[1152]) );
  XOR2_X2 _f_permutation__round__U3014  ( .A(_f_permutation__round__N3453 ), 
        .B(_f_permutation__round__c[1389] ), .Z(
        _f_permutation__round_out[1153]) );
  XOR2_X2 _f_permutation__round__U3013  ( .A(_f_permutation__round__N3451 ), 
        .B(_f_permutation__round__c[1390] ), .Z(
        _f_permutation__round_out[1154]) );
  XOR2_X2 _f_permutation__round__U3012  ( .A(_f_permutation__round__N3449 ), 
        .B(_f_permutation__round__c[1391] ), .Z(
        _f_permutation__round_out[1155]) );
  XOR2_X2 _f_permutation__round__U3011  ( .A(_f_permutation__round__N3447 ), 
        .B(_f_permutation__round__c[1392] ), .Z(
        _f_permutation__round_out[1156]) );
  XOR2_X2 _f_permutation__round__U3010  ( .A(_f_permutation__round__N3445 ), 
        .B(_f_permutation__round__c[1393] ), .Z(
        _f_permutation__round_out[1157]) );
  XOR2_X2 _f_permutation__round__U3009  ( .A(_f_permutation__round__N3443 ), 
        .B(_f_permutation__round__c[1394] ), .Z(
        _f_permutation__round_out[1158]) );
  XOR2_X2 _f_permutation__round__U3008  ( .A(_f_permutation__round__N3441 ), 
        .B(_f_permutation__round__c[1395] ), .Z(
        _f_permutation__round_out[1159]) );
  XOR2_X2 _f_permutation__round__U3007  ( .A(_f_permutation__round__N3439 ), 
        .B(_f_permutation__round__c[1396] ), .Z(
        _f_permutation__round_out[1160]) );
  XOR2_X2 _f_permutation__round__U3006  ( .A(_f_permutation__round__N3437 ), 
        .B(_f_permutation__round__c[1397] ), .Z(
        _f_permutation__round_out[1161]) );
  XOR2_X2 _f_permutation__round__U3005  ( .A(_f_permutation__round__N3435 ), 
        .B(_f_permutation__round__c[1398] ), .Z(
        _f_permutation__round_out[1162]) );
  XOR2_X2 _f_permutation__round__U3004  ( .A(_f_permutation__round__N3433 ), 
        .B(_f_permutation__round__c[1399] ), .Z(
        _f_permutation__round_out[1163]) );
  XOR2_X2 _f_permutation__round__U3003  ( .A(_f_permutation__round__N3431 ), 
        .B(_f_permutation__round__c[1400] ), .Z(
        _f_permutation__round_out[1164]) );
  XOR2_X2 _f_permutation__round__U3002  ( .A(_f_permutation__round__N3429 ), 
        .B(_f_permutation__round__c[1401] ), .Z(
        _f_permutation__round_out[1165]) );
  XOR2_X2 _f_permutation__round__U3001  ( .A(_f_permutation__round__N3427 ), 
        .B(_f_permutation__round__c[1402] ), .Z(
        _f_permutation__round_out[1166]) );
  XOR2_X2 _f_permutation__round__U3000  ( .A(_f_permutation__round__N3425 ), 
        .B(_f_permutation__round__c[1403] ), .Z(
        _f_permutation__round_out[1167]) );
  XOR2_X2 _f_permutation__round__U2999  ( .A(_f_permutation__round__N3423 ), 
        .B(_f_permutation__round__c[1404] ), .Z(
        _f_permutation__round_out[1168]) );
  XOR2_X2 _f_permutation__round__U2998  ( .A(_f_permutation__round__N3421 ), 
        .B(_f_permutation__round__c[1405] ), .Z(
        _f_permutation__round_out[1169]) );
  XOR2_X2 _f_permutation__round__U2997  ( .A(_f_permutation__round__N3419 ), 
        .B(_f_permutation__round__c[1406] ), .Z(
        _f_permutation__round_out[1170]) );
  XOR2_X2 _f_permutation__round__U2996  ( .A(_f_permutation__round__N3417 ), 
        .B(_f_permutation__round__c[1407] ), .Z(
        _f_permutation__round_out[1171]) );
  XOR2_X2 _f_permutation__round__U2995  ( .A(_f_permutation__round__N3415 ), 
        .B(_f_permutation__round__c[1344] ), .Z(
        _f_permutation__round_out[1172]) );
  XOR2_X2 _f_permutation__round__U2994  ( .A(_f_permutation__round__N3413 ), 
        .B(_f_permutation__round__c[1345] ), .Z(
        _f_permutation__round_out[1173]) );
  XOR2_X2 _f_permutation__round__U2993  ( .A(_f_permutation__round__N3411 ), 
        .B(_f_permutation__round__c[1346] ), .Z(
        _f_permutation__round_out[1174]) );
  XOR2_X2 _f_permutation__round__U2992  ( .A(_f_permutation__round__N3409 ), 
        .B(_f_permutation__round__c[1347] ), .Z(
        _f_permutation__round_out[1175]) );
  XOR2_X2 _f_permutation__round__U2991  ( .A(_f_permutation__round__N3407 ), 
        .B(_f_permutation__round__c[1348] ), .Z(
        _f_permutation__round_out[1176]) );
  XOR2_X2 _f_permutation__round__U2990  ( .A(_f_permutation__round__N3405 ), 
        .B(_f_permutation__round__c[1349] ), .Z(
        _f_permutation__round_out[1177]) );
  XOR2_X2 _f_permutation__round__U2989  ( .A(_f_permutation__round__N3403 ), 
        .B(_f_permutation__round__c[1350] ), .Z(
        _f_permutation__round_out[1178]) );
  XOR2_X2 _f_permutation__round__U2988  ( .A(_f_permutation__round__N3401 ), 
        .B(_f_permutation__round__c[1351] ), .Z(
        _f_permutation__round_out[1179]) );
  XOR2_X2 _f_permutation__round__U2987  ( .A(_f_permutation__round__N3399 ), 
        .B(_f_permutation__round__c[1352] ), .Z(
        _f_permutation__round_out[1180]) );
  XOR2_X2 _f_permutation__round__U2986  ( .A(_f_permutation__round__N3397 ), 
        .B(_f_permutation__round__c[1353] ), .Z(
        _f_permutation__round_out[1181]) );
  XOR2_X2 _f_permutation__round__U2985  ( .A(_f_permutation__round__N3395 ), 
        .B(_f_permutation__round__c[1354] ), .Z(
        _f_permutation__round_out[1182]) );
  XOR2_X2 _f_permutation__round__U2984  ( .A(_f_permutation__round__N3393 ), 
        .B(_f_permutation__round__c[1355] ), .Z(
        _f_permutation__round_out[1183]) );
  XOR2_X2 _f_permutation__round__U2983  ( .A(_f_permutation__round__N3391 ), 
        .B(_f_permutation__round__c[1356] ), .Z(
        _f_permutation__round_out[1184]) );
  XOR2_X2 _f_permutation__round__U2982  ( .A(_f_permutation__round__N3389 ), 
        .B(_f_permutation__round__c[1357] ), .Z(
        _f_permutation__round_out[1185]) );
  XOR2_X2 _f_permutation__round__U2981  ( .A(_f_permutation__round__N3387 ), 
        .B(_f_permutation__round__c[1358] ), .Z(
        _f_permutation__round_out[1186]) );
  XOR2_X2 _f_permutation__round__U2980  ( .A(_f_permutation__round__N3385 ), 
        .B(_f_permutation__round__c[1359] ), .Z(
        _f_permutation__round_out[1187]) );
  XOR2_X2 _f_permutation__round__U2979  ( .A(_f_permutation__round__N3383 ), 
        .B(_f_permutation__round__c[1360] ), .Z(
        _f_permutation__round_out[1188]) );
  XOR2_X2 _f_permutation__round__U2978  ( .A(_f_permutation__round__N3381 ), 
        .B(_f_permutation__round__c[1361] ), .Z(
        _f_permutation__round_out[1189]) );
  XOR2_X2 _f_permutation__round__U2977  ( .A(_f_permutation__round__N3379 ), 
        .B(_f_permutation__round__c[1362] ), .Z(
        _f_permutation__round_out[1190]) );
  XOR2_X2 _f_permutation__round__U2976  ( .A(_f_permutation__round__N3377 ), 
        .B(_f_permutation__round__c[1363] ), .Z(
        _f_permutation__round_out[1191]) );
  XOR2_X2 _f_permutation__round__U2975  ( .A(_f_permutation__round__N3375 ), 
        .B(_f_permutation__round__c[1364] ), .Z(
        _f_permutation__round_out[1192]) );
  XOR2_X2 _f_permutation__round__U2974  ( .A(_f_permutation__round__N3373 ), 
        .B(_f_permutation__round__c[1365] ), .Z(
        _f_permutation__round_out[1193]) );
  XOR2_X2 _f_permutation__round__U2973  ( .A(_f_permutation__round__N3371 ), 
        .B(_f_permutation__round__c[1366] ), .Z(
        _f_permutation__round_out[1194]) );
  XOR2_X2 _f_permutation__round__U2972  ( .A(_f_permutation__round__N3369 ), 
        .B(_f_permutation__round__c[1367] ), .Z(
        _f_permutation__round_out[1195]) );
  XOR2_X2 _f_permutation__round__U2971  ( .A(_f_permutation__round__N3367 ), 
        .B(_f_permutation__round__c[1368] ), .Z(
        _f_permutation__round_out[1196]) );
  XOR2_X2 _f_permutation__round__U2970  ( .A(_f_permutation__round__N3365 ), 
        .B(_f_permutation__round__c[1369] ), .Z(
        _f_permutation__round_out[1197]) );
  XOR2_X2 _f_permutation__round__U2969  ( .A(_f_permutation__round__N3363 ), 
        .B(_f_permutation__round__c[1370] ), .Z(
        _f_permutation__round_out[1198]) );
  XOR2_X2 _f_permutation__round__U2968  ( .A(_f_permutation__round__N3361 ), 
        .B(_f_permutation__round__c[1371] ), .Z(
        _f_permutation__round_out[1199]) );
  XOR2_X2 _f_permutation__round__U2967  ( .A(_f_permutation__round__N3359 ), 
        .B(_f_permutation__round__c[1372] ), .Z(
        _f_permutation__round_out[1200]) );
  XOR2_X2 _f_permutation__round__U2966  ( .A(_f_permutation__round__N3357 ), 
        .B(_f_permutation__round__c[1373] ), .Z(
        _f_permutation__round_out[1201]) );
  XOR2_X2 _f_permutation__round__U2965  ( .A(_f_permutation__round__N3355 ), 
        .B(_f_permutation__round__c[1374] ), .Z(
        _f_permutation__round_out[1202]) );
  XOR2_X2 _f_permutation__round__U2964  ( .A(_f_permutation__round__N3353 ), 
        .B(_f_permutation__round__c[1375] ), .Z(
        _f_permutation__round_out[1203]) );
  XOR2_X2 _f_permutation__round__U2963  ( .A(_f_permutation__round__N3351 ), 
        .B(_f_permutation__round__c[1376] ), .Z(
        _f_permutation__round_out[1204]) );
  XOR2_X2 _f_permutation__round__U2962  ( .A(_f_permutation__round__N3349 ), 
        .B(_f_permutation__round__c[1377] ), .Z(
        _f_permutation__round_out[1205]) );
  XOR2_X2 _f_permutation__round__U2961  ( .A(_f_permutation__round__N3347 ), 
        .B(_f_permutation__round__c[1378] ), .Z(
        _f_permutation__round_out[1206]) );
  XOR2_X2 _f_permutation__round__U2960  ( .A(_f_permutation__round__N3345 ), 
        .B(_f_permutation__round__c[1379] ), .Z(
        _f_permutation__round_out[1207]) );
  XOR2_X2 _f_permutation__round__U2959  ( .A(_f_permutation__round__N3343 ), 
        .B(_f_permutation__round__c[1380] ), .Z(
        _f_permutation__round_out[1208]) );
  XOR2_X2 _f_permutation__round__U2958  ( .A(_f_permutation__round__N3341 ), 
        .B(_f_permutation__round__c[1381] ), .Z(
        _f_permutation__round_out[1209]) );
  XOR2_X2 _f_permutation__round__U2957  ( .A(_f_permutation__round__N3339 ), 
        .B(_f_permutation__round__c[1382] ), .Z(
        _f_permutation__round_out[1210]) );
  XOR2_X2 _f_permutation__round__U2956  ( .A(_f_permutation__round__N3337 ), 
        .B(_f_permutation__round__c[1383] ), .Z(
        _f_permutation__round_out[1211]) );
  XOR2_X2 _f_permutation__round__U2955  ( .A(_f_permutation__round__N3335 ), 
        .B(_f_permutation__round__c[1384] ), .Z(
        _f_permutation__round_out[1212]) );
  XOR2_X2 _f_permutation__round__U2954  ( .A(_f_permutation__round__N3333 ), 
        .B(_f_permutation__round__c[1385] ), .Z(
        _f_permutation__round_out[1213]) );
  XOR2_X2 _f_permutation__round__U2953  ( .A(_f_permutation__round__N3331 ), 
        .B(_f_permutation__round__c[1386] ), .Z(
        _f_permutation__round_out[1214]) );
  XOR2_X2 _f_permutation__round__U2952  ( .A(_f_permutation__round__N3329 ), 
        .B(_f_permutation__round__c[1387] ), .Z(
        _f_permutation__round_out[1215]) );
  XOR2_X2 _f_permutation__round__U2951  ( .A(_f_permutation__round__N3327 ), 
        .B(_f_permutation__round__c[996] ), .Z(
        _f_permutation__round_out[1216]) );
  XOR2_X2 _f_permutation__round__U2950  ( .A(_f_permutation__round__N3325 ), 
        .B(_f_permutation__round__c[997] ), .Z(
        _f_permutation__round_out[1217]) );
  XOR2_X2 _f_permutation__round__U2949  ( .A(_f_permutation__round__N3323 ), 
        .B(_f_permutation__round__c[998] ), .Z(
        _f_permutation__round_out[1218]) );
  XOR2_X2 _f_permutation__round__U2948  ( .A(_f_permutation__round__N3321 ), 
        .B(_f_permutation__round__c[999] ), .Z(
        _f_permutation__round_out[1219]) );
  XOR2_X2 _f_permutation__round__U2947  ( .A(_f_permutation__round__N3319 ), 
        .B(_f_permutation__round__c[1000] ), .Z(
        _f_permutation__round_out[1220]) );
  XOR2_X2 _f_permutation__round__U2946  ( .A(_f_permutation__round__N3317 ), 
        .B(_f_permutation__round__c[1001] ), .Z(
        _f_permutation__round_out[1221]) );
  XOR2_X2 _f_permutation__round__U2945  ( .A(_f_permutation__round__N3315 ), 
        .B(_f_permutation__round__c[1002] ), .Z(
        _f_permutation__round_out[1222]) );
  XOR2_X2 _f_permutation__round__U2944  ( .A(_f_permutation__round__N3313 ), 
        .B(_f_permutation__round__c[1003] ), .Z(
        _f_permutation__round_out[1223]) );
  XOR2_X2 _f_permutation__round__U2943  ( .A(_f_permutation__round__N3311 ), 
        .B(_f_permutation__round__c[1004] ), .Z(
        _f_permutation__round_out[1224]) );
  XOR2_X2 _f_permutation__round__U2942  ( .A(_f_permutation__round__N3309 ), 
        .B(_f_permutation__round__c[1005] ), .Z(
        _f_permutation__round_out[1225]) );
  XOR2_X2 _f_permutation__round__U2941  ( .A(_f_permutation__round__N3307 ), 
        .B(_f_permutation__round__c[1006] ), .Z(
        _f_permutation__round_out[1226]) );
  XOR2_X2 _f_permutation__round__U2940  ( .A(_f_permutation__round__N3305 ), 
        .B(_f_permutation__round__c[1007] ), .Z(
        _f_permutation__round_out[1227]) );
  XOR2_X2 _f_permutation__round__U2939  ( .A(_f_permutation__round__N3303 ), 
        .B(_f_permutation__round__c[1008] ), .Z(
        _f_permutation__round_out[1228]) );
  XOR2_X2 _f_permutation__round__U2938  ( .A(_f_permutation__round__N3301 ), 
        .B(_f_permutation__round__c[1009] ), .Z(
        _f_permutation__round_out[1229]) );
  XOR2_X2 _f_permutation__round__U2937  ( .A(_f_permutation__round__N3299 ), 
        .B(_f_permutation__round__c[1010] ), .Z(
        _f_permutation__round_out[1230]) );
  XOR2_X2 _f_permutation__round__U2936  ( .A(_f_permutation__round__N3297 ), 
        .B(_f_permutation__round__c[1011] ), .Z(
        _f_permutation__round_out[1231]) );
  XOR2_X2 _f_permutation__round__U2935  ( .A(_f_permutation__round__N3295 ), 
        .B(_f_permutation__round__c[1012] ), .Z(
        _f_permutation__round_out[1232]) );
  XOR2_X2 _f_permutation__round__U2934  ( .A(_f_permutation__round__N3293 ), 
        .B(_f_permutation__round__c[1013] ), .Z(
        _f_permutation__round_out[1233]) );
  XOR2_X2 _f_permutation__round__U2933  ( .A(_f_permutation__round__N3291 ), 
        .B(_f_permutation__round__c[1014] ), .Z(
        _f_permutation__round_out[1234]) );
  XOR2_X2 _f_permutation__round__U2932  ( .A(_f_permutation__round__N3289 ), 
        .B(_f_permutation__round__c[1015] ), .Z(
        _f_permutation__round_out[1235]) );
  XOR2_X2 _f_permutation__round__U2931  ( .A(_f_permutation__round__N3287 ), 
        .B(_f_permutation__round__c[1016] ), .Z(
        _f_permutation__round_out[1236]) );
  XOR2_X2 _f_permutation__round__U2930  ( .A(_f_permutation__round__N3285 ), 
        .B(_f_permutation__round__c[1017] ), .Z(
        _f_permutation__round_out[1237]) );
  XOR2_X2 _f_permutation__round__U2929  ( .A(_f_permutation__round__N3283 ), 
        .B(_f_permutation__round__c[1018] ), .Z(
        _f_permutation__round_out[1238]) );
  XOR2_X2 _f_permutation__round__U2928  ( .A(_f_permutation__round__N3281 ), 
        .B(_f_permutation__round__c[1019] ), .Z(
        _f_permutation__round_out[1239]) );
  XOR2_X2 _f_permutation__round__U2927  ( .A(_f_permutation__round__N3279 ), 
        .B(_f_permutation__round__c[1020] ), .Z(
        _f_permutation__round_out[1240]) );
  XOR2_X2 _f_permutation__round__U2926  ( .A(_f_permutation__round__N3277 ), 
        .B(_f_permutation__round__c[1021] ), .Z(
        _f_permutation__round_out[1241]) );
  XOR2_X2 _f_permutation__round__U2925  ( .A(_f_permutation__round__N3275 ), 
        .B(_f_permutation__round__c[1022] ), .Z(
        _f_permutation__round_out[1242]) );
  XOR2_X2 _f_permutation__round__U2924  ( .A(_f_permutation__round__N3273 ), 
        .B(_f_permutation__round__c[1023] ), .Z(
        _f_permutation__round_out[1243]) );
  XOR2_X2 _f_permutation__round__U2923  ( .A(_f_permutation__round__N3271 ), 
        .B(_f_permutation__round__c[960] ), .Z(
        _f_permutation__round_out[1244]) );
  XOR2_X2 _f_permutation__round__U2922  ( .A(_f_permutation__round__N3269 ), 
        .B(_f_permutation__round__c[961] ), .Z(
        _f_permutation__round_out[1245]) );
  XOR2_X2 _f_permutation__round__U2921  ( .A(_f_permutation__round__N3267 ), 
        .B(_f_permutation__round__c[962] ), .Z(
        _f_permutation__round_out[1246]) );
  XOR2_X2 _f_permutation__round__U2920  ( .A(_f_permutation__round__N3265 ), 
        .B(_f_permutation__round__c[963] ), .Z(
        _f_permutation__round_out[1247]) );
  XOR2_X2 _f_permutation__round__U2919  ( .A(_f_permutation__round__N3263 ), 
        .B(_f_permutation__round__c[964] ), .Z(
        _f_permutation__round_out[1248]) );
  XOR2_X2 _f_permutation__round__U2918  ( .A(_f_permutation__round__N3261 ), 
        .B(_f_permutation__round__c[965] ), .Z(
        _f_permutation__round_out[1249]) );
  XOR2_X2 _f_permutation__round__U2917  ( .A(_f_permutation__round__N3259 ), 
        .B(_f_permutation__round__c[966] ), .Z(
        _f_permutation__round_out[1250]) );
  XOR2_X2 _f_permutation__round__U2916  ( .A(_f_permutation__round__N3257 ), 
        .B(_f_permutation__round__c[967] ), .Z(
        _f_permutation__round_out[1251]) );
  XOR2_X2 _f_permutation__round__U2915  ( .A(_f_permutation__round__N3255 ), 
        .B(_f_permutation__round__c[968] ), .Z(
        _f_permutation__round_out[1252]) );
  XOR2_X2 _f_permutation__round__U2914  ( .A(_f_permutation__round__N3253 ), 
        .B(_f_permutation__round__c[969] ), .Z(
        _f_permutation__round_out[1253]) );
  XOR2_X2 _f_permutation__round__U2913  ( .A(_f_permutation__round__N3251 ), 
        .B(_f_permutation__round__c[970] ), .Z(
        _f_permutation__round_out[1254]) );
  XOR2_X2 _f_permutation__round__U2912  ( .A(_f_permutation__round__N3249 ), 
        .B(_f_permutation__round__c[971] ), .Z(
        _f_permutation__round_out[1255]) );
  XOR2_X2 _f_permutation__round__U2911  ( .A(_f_permutation__round__N3247 ), 
        .B(_f_permutation__round__c[972] ), .Z(
        _f_permutation__round_out[1256]) );
  XOR2_X2 _f_permutation__round__U2910  ( .A(_f_permutation__round__N3245 ), 
        .B(_f_permutation__round__c[973] ), .Z(
        _f_permutation__round_out[1257]) );
  XOR2_X2 _f_permutation__round__U2909  ( .A(_f_permutation__round__N3243 ), 
        .B(_f_permutation__round__c[974] ), .Z(
        _f_permutation__round_out[1258]) );
  XOR2_X2 _f_permutation__round__U2908  ( .A(_f_permutation__round__N3241 ), 
        .B(_f_permutation__round__c[975] ), .Z(
        _f_permutation__round_out[1259]) );
  XOR2_X2 _f_permutation__round__U2907  ( .A(_f_permutation__round__N3239 ), 
        .B(_f_permutation__round__c[976] ), .Z(
        _f_permutation__round_out[1260]) );
  XOR2_X2 _f_permutation__round__U2906  ( .A(_f_permutation__round__N3237 ), 
        .B(_f_permutation__round__c[977] ), .Z(
        _f_permutation__round_out[1261]) );
  XOR2_X2 _f_permutation__round__U2905  ( .A(_f_permutation__round__N3235 ), 
        .B(_f_permutation__round__c[978] ), .Z(
        _f_permutation__round_out[1262]) );
  XOR2_X2 _f_permutation__round__U2904  ( .A(_f_permutation__round__N3233 ), 
        .B(_f_permutation__round__c[979] ), .Z(
        _f_permutation__round_out[1263]) );
  XOR2_X2 _f_permutation__round__U2903  ( .A(_f_permutation__round__N3231 ), 
        .B(_f_permutation__round__c[980] ), .Z(
        _f_permutation__round_out[1264]) );
  XOR2_X2 _f_permutation__round__U2902  ( .A(_f_permutation__round__N3229 ), 
        .B(_f_permutation__round__c[981] ), .Z(
        _f_permutation__round_out[1265]) );
  XOR2_X2 _f_permutation__round__U2901  ( .A(_f_permutation__round__N3227 ), 
        .B(_f_permutation__round__c[982] ), .Z(
        _f_permutation__round_out[1266]) );
  XOR2_X2 _f_permutation__round__U2900  ( .A(_f_permutation__round__N3225 ), 
        .B(_f_permutation__round__c[983] ), .Z(
        _f_permutation__round_out[1267]) );
  XOR2_X2 _f_permutation__round__U2899  ( .A(_f_permutation__round__N3223 ), 
        .B(_f_permutation__round__c[984] ), .Z(
        _f_permutation__round_out[1268]) );
  XOR2_X2 _f_permutation__round__U2898  ( .A(_f_permutation__round__N3221 ), 
        .B(_f_permutation__round__c[985] ), .Z(
        _f_permutation__round_out[1269]) );
  XOR2_X2 _f_permutation__round__U2897  ( .A(_f_permutation__round__N3219 ), 
        .B(_f_permutation__round__c[986] ), .Z(
        _f_permutation__round_out[1270]) );
  XOR2_X2 _f_permutation__round__U2896  ( .A(_f_permutation__round__N3217 ), 
        .B(_f_permutation__round__c[987] ), .Z(
        _f_permutation__round_out[1271]) );
  XOR2_X2 _f_permutation__round__U2895  ( .A(_f_permutation__round__N3215 ), 
        .B(_f_permutation__round__c[988] ), .Z(
        _f_permutation__round_out[1272]) );
  XOR2_X2 _f_permutation__round__U2894  ( .A(_f_permutation__round__N3213 ), 
        .B(_f_permutation__round__c[989] ), .Z(
        _f_permutation__round_out[1273]) );
  XOR2_X2 _f_permutation__round__U2893  ( .A(_f_permutation__round__N3211 ), 
        .B(_f_permutation__round__c[990] ), .Z(
        _f_permutation__round_out[1274]) );
  XOR2_X2 _f_permutation__round__U2892  ( .A(_f_permutation__round__N3209 ), 
        .B(_f_permutation__round__c[991] ), .Z(
        _f_permutation__round_out[1275]) );
  XOR2_X2 _f_permutation__round__U2891  ( .A(_f_permutation__round__N3207 ), 
        .B(_f_permutation__round__c[992] ), .Z(
        _f_permutation__round_out[1276]) );
  XOR2_X2 _f_permutation__round__U2890  ( .A(_f_permutation__round__N3205 ), 
        .B(_f_permutation__round__c[993] ), .Z(
        _f_permutation__round_out[1277]) );
  XOR2_X2 _f_permutation__round__U2889  ( .A(_f_permutation__round__N3203 ), 
        .B(_f_permutation__round__c[994] ), .Z(
        _f_permutation__round_out[1278]) );
  XOR2_X2 _f_permutation__round__U2888  ( .A(_f_permutation__round__N3201 ), 
        .B(_f_permutation__round__c[995] ), .Z(
        _f_permutation__round_out[1279]) );
  XOR2_X2 _f_permutation__round__U2887  ( .A(_f_permutation__round__N3199 ), 
        .B(_f_permutation__round__c[1586] ), .Z(
        _f_permutation__round_out[1280]) );
  XOR2_X2 _f_permutation__round__U2886  ( .A(_f_permutation__round__N3197 ), 
        .B(_f_permutation__round__c[1587] ), .Z(
        _f_permutation__round_out[1281]) );
  XOR2_X2 _f_permutation__round__U2885  ( .A(_f_permutation__round__N3195 ), 
        .B(_f_permutation__round__c[1588] ), .Z(
        _f_permutation__round_out[1282]) );
  XOR2_X2 _f_permutation__round__U2884  ( .A(_f_permutation__round__N3193 ), 
        .B(_f_permutation__round__c[1589] ), .Z(
        _f_permutation__round_out[1283]) );
  XOR2_X2 _f_permutation__round__U2883  ( .A(_f_permutation__round__N3191 ), 
        .B(_f_permutation__round__c[1590] ), .Z(
        _f_permutation__round_out[1284]) );
  XOR2_X2 _f_permutation__round__U2882  ( .A(_f_permutation__round__N3189 ), 
        .B(_f_permutation__round__c[1591] ), .Z(
        _f_permutation__round_out[1285]) );
  XOR2_X2 _f_permutation__round__U2881  ( .A(_f_permutation__round__N3187 ), 
        .B(_f_permutation__round__c[1592] ), .Z(
        _f_permutation__round_out[1286]) );
  XOR2_X2 _f_permutation__round__U2880  ( .A(_f_permutation__round__N3185 ), 
        .B(_f_permutation__round__c[1593] ), .Z(
        _f_permutation__round_out[1287]) );
  XOR2_X2 _f_permutation__round__U2879  ( .A(_f_permutation__round__N3183 ), 
        .B(_f_permutation__round__c[1594] ), .Z(
        _f_permutation__round_out[1288]) );
  XOR2_X2 _f_permutation__round__U2878  ( .A(_f_permutation__round__N3181 ), 
        .B(_f_permutation__round__c[1595] ), .Z(
        _f_permutation__round_out[1289]) );
  XOR2_X2 _f_permutation__round__U2877  ( .A(_f_permutation__round__N3179 ), 
        .B(_f_permutation__round__c[1596] ), .Z(
        _f_permutation__round_out[1290]) );
  XOR2_X2 _f_permutation__round__U2876  ( .A(_f_permutation__round__N3177 ), 
        .B(_f_permutation__round__c[1597] ), .Z(
        _f_permutation__round_out[1291]) );
  XOR2_X2 _f_permutation__round__U2875  ( .A(_f_permutation__round__N3175 ), 
        .B(_f_permutation__round__c[1598] ), .Z(
        _f_permutation__round_out[1292]) );
  XOR2_X2 _f_permutation__round__U2874  ( .A(_f_permutation__round__N3173 ), 
        .B(_f_permutation__round__c[1599] ), .Z(
        _f_permutation__round_out[1293]) );
  XOR2_X2 _f_permutation__round__U2873  ( .A(_f_permutation__round__N3171 ), 
        .B(_f_permutation__round__c[1536] ), .Z(
        _f_permutation__round_out[1294]) );
  XOR2_X2 _f_permutation__round__U2872  ( .A(_f_permutation__round__N3169 ), 
        .B(_f_permutation__round__c[1537] ), .Z(
        _f_permutation__round_out[1295]) );
  XOR2_X2 _f_permutation__round__U2871  ( .A(_f_permutation__round__N3167 ), 
        .B(_f_permutation__round__c[1538] ), .Z(
        _f_permutation__round_out[1296]) );
  XOR2_X2 _f_permutation__round__U2870  ( .A(_f_permutation__round__N3165 ), 
        .B(_f_permutation__round__c[1539] ), .Z(
        _f_permutation__round_out[1297]) );
  XOR2_X2 _f_permutation__round__U2869  ( .A(_f_permutation__round__N3163 ), 
        .B(_f_permutation__round__c[1540] ), .Z(
        _f_permutation__round_out[1298]) );
  XOR2_X2 _f_permutation__round__U2868  ( .A(_f_permutation__round__N3161 ), 
        .B(_f_permutation__round__c[1541] ), .Z(
        _f_permutation__round_out[1299]) );
  XOR2_X2 _f_permutation__round__U2867  ( .A(_f_permutation__round__N3159 ), 
        .B(_f_permutation__round__c[1542] ), .Z(
        _f_permutation__round_out[1300]) );
  XOR2_X2 _f_permutation__round__U2866  ( .A(_f_permutation__round__N3157 ), 
        .B(_f_permutation__round__c[1543] ), .Z(
        _f_permutation__round_out[1301]) );
  XOR2_X2 _f_permutation__round__U2865  ( .A(_f_permutation__round__N3155 ), 
        .B(_f_permutation__round__c[1544] ), .Z(
        _f_permutation__round_out[1302]) );
  XOR2_X2 _f_permutation__round__U2864  ( .A(_f_permutation__round__N3153 ), 
        .B(_f_permutation__round__c[1545] ), .Z(
        _f_permutation__round_out[1303]) );
  XOR2_X2 _f_permutation__round__U2863  ( .A(_f_permutation__round__N3151 ), 
        .B(_f_permutation__round__c[1546] ), .Z(
        _f_permutation__round_out[1304]) );
  XOR2_X2 _f_permutation__round__U2862  ( .A(_f_permutation__round__N3149 ), 
        .B(_f_permutation__round__c[1547] ), .Z(
        _f_permutation__round_out[1305]) );
  XOR2_X2 _f_permutation__round__U2861  ( .A(_f_permutation__round__N3147 ), 
        .B(_f_permutation__round__c[1548] ), .Z(
        _f_permutation__round_out[1306]) );
  XOR2_X2 _f_permutation__round__U2860  ( .A(_f_permutation__round__N3145 ), 
        .B(_f_permutation__round__c[1549] ), .Z(
        _f_permutation__round_out[1307]) );
  XOR2_X2 _f_permutation__round__U2859  ( .A(_f_permutation__round__N3143 ), 
        .B(_f_permutation__round__c[1550] ), .Z(
        _f_permutation__round_out[1308]) );
  XOR2_X2 _f_permutation__round__U2858  ( .A(_f_permutation__round__N3141 ), 
        .B(_f_permutation__round__c[1551] ), .Z(
        _f_permutation__round_out[1309]) );
  XOR2_X2 _f_permutation__round__U2857  ( .A(_f_permutation__round__N3139 ), 
        .B(_f_permutation__round__c[1552] ), .Z(
        _f_permutation__round_out[1310]) );
  XOR2_X2 _f_permutation__round__U2856  ( .A(_f_permutation__round__N3137 ), 
        .B(_f_permutation__round__c[1553] ), .Z(
        _f_permutation__round_out[1311]) );
  XOR2_X2 _f_permutation__round__U2855  ( .A(_f_permutation__round__N3135 ), 
        .B(_f_permutation__round__c[1554] ), .Z(
        _f_permutation__round_out[1312]) );
  XOR2_X2 _f_permutation__round__U2854  ( .A(_f_permutation__round__N3133 ), 
        .B(_f_permutation__round__c[1555] ), .Z(
        _f_permutation__round_out[1313]) );
  XOR2_X2 _f_permutation__round__U2853  ( .A(_f_permutation__round__N3131 ), 
        .B(_f_permutation__round__c[1556] ), .Z(
        _f_permutation__round_out[1314]) );
  XOR2_X2 _f_permutation__round__U2852  ( .A(_f_permutation__round__N3129 ), 
        .B(_f_permutation__round__c[1557] ), .Z(
        _f_permutation__round_out[1315]) );
  XOR2_X2 _f_permutation__round__U2851  ( .A(_f_permutation__round__N3127 ), 
        .B(_f_permutation__round__c[1558] ), .Z(
        _f_permutation__round_out[1316]) );
  XOR2_X2 _f_permutation__round__U2850  ( .A(_f_permutation__round__N3125 ), 
        .B(_f_permutation__round__c[1559] ), .Z(
        _f_permutation__round_out[1317]) );
  XOR2_X2 _f_permutation__round__U2849  ( .A(_f_permutation__round__N3123 ), 
        .B(_f_permutation__round__c[1560] ), .Z(
        _f_permutation__round_out[1318]) );
  XOR2_X2 _f_permutation__round__U2848  ( .A(_f_permutation__round__N3121 ), 
        .B(_f_permutation__round__c[1561] ), .Z(
        _f_permutation__round_out[1319]) );
  XOR2_X2 _f_permutation__round__U2847  ( .A(_f_permutation__round__N3119 ), 
        .B(_f_permutation__round__c[1562] ), .Z(
        _f_permutation__round_out[1320]) );
  XOR2_X2 _f_permutation__round__U2846  ( .A(_f_permutation__round__N3117 ), 
        .B(_f_permutation__round__c[1563] ), .Z(
        _f_permutation__round_out[1321]) );
  XOR2_X2 _f_permutation__round__U2845  ( .A(_f_permutation__round__N3115 ), 
        .B(_f_permutation__round__c[1564] ), .Z(
        _f_permutation__round_out[1322]) );
  XOR2_X2 _f_permutation__round__U2844  ( .A(_f_permutation__round__N3113 ), 
        .B(_f_permutation__round__c[1565] ), .Z(
        _f_permutation__round_out[1323]) );
  XOR2_X2 _f_permutation__round__U2843  ( .A(_f_permutation__round__N3111 ), 
        .B(_f_permutation__round__c[1566] ), .Z(
        _f_permutation__round_out[1324]) );
  XOR2_X2 _f_permutation__round__U2842  ( .A(_f_permutation__round__N3109 ), 
        .B(_f_permutation__round__c[1567] ), .Z(
        _f_permutation__round_out[1325]) );
  XOR2_X2 _f_permutation__round__U2841  ( .A(_f_permutation__round__N3107 ), 
        .B(_f_permutation__round__c[1568] ), .Z(
        _f_permutation__round_out[1326]) );
  XOR2_X2 _f_permutation__round__U2840  ( .A(_f_permutation__round__N3105 ), 
        .B(_f_permutation__round__c[1569] ), .Z(
        _f_permutation__round_out[1327]) );
  XOR2_X2 _f_permutation__round__U2839  ( .A(_f_permutation__round__N3103 ), 
        .B(_f_permutation__round__c[1570] ), .Z(
        _f_permutation__round_out[1328]) );
  XOR2_X2 _f_permutation__round__U2838  ( .A(_f_permutation__round__N3101 ), 
        .B(_f_permutation__round__c[1571] ), .Z(
        _f_permutation__round_out[1329]) );
  XOR2_X2 _f_permutation__round__U2837  ( .A(_f_permutation__round__N3099 ), 
        .B(_f_permutation__round__c[1572] ), .Z(
        _f_permutation__round_out[1330]) );
  XOR2_X2 _f_permutation__round__U2836  ( .A(_f_permutation__round__N3097 ), 
        .B(_f_permutation__round__c[1573] ), .Z(
        _f_permutation__round_out[1331]) );
  XOR2_X2 _f_permutation__round__U2835  ( .A(_f_permutation__round__N3095 ), 
        .B(_f_permutation__round__c[1574] ), .Z(
        _f_permutation__round_out[1332]) );
  XOR2_X2 _f_permutation__round__U2834  ( .A(_f_permutation__round__N3093 ), 
        .B(_f_permutation__round__c[1575] ), .Z(
        _f_permutation__round_out[1333]) );
  XOR2_X2 _f_permutation__round__U2833  ( .A(_f_permutation__round__N3091 ), 
        .B(_f_permutation__round__c[1576] ), .Z(
        _f_permutation__round_out[1334]) );
  XOR2_X2 _f_permutation__round__U2832  ( .A(_f_permutation__round__N3089 ), 
        .B(_f_permutation__round__c[1577] ), .Z(
        _f_permutation__round_out[1335]) );
  XOR2_X2 _f_permutation__round__U2831  ( .A(_f_permutation__round__N3087 ), 
        .B(_f_permutation__round__c[1578] ), .Z(
        _f_permutation__round_out[1336]) );
  XOR2_X2 _f_permutation__round__U2830  ( .A(_f_permutation__round__N3085 ), 
        .B(_f_permutation__round__c[1579] ), .Z(
        _f_permutation__round_out[1337]) );
  XOR2_X2 _f_permutation__round__U2829  ( .A(_f_permutation__round__N3083 ), 
        .B(_f_permutation__round__c[1580] ), .Z(
        _f_permutation__round_out[1338]) );
  XOR2_X2 _f_permutation__round__U2828  ( .A(_f_permutation__round__N3081 ), 
        .B(_f_permutation__round__c[1581] ), .Z(
        _f_permutation__round_out[1339]) );
  XOR2_X2 _f_permutation__round__U2827  ( .A(_f_permutation__round__N3079 ), 
        .B(_f_permutation__round__c[1582] ), .Z(
        _f_permutation__round_out[1340]) );
  XOR2_X2 _f_permutation__round__U2826  ( .A(_f_permutation__round__N3077 ), 
        .B(_f_permutation__round__c[1583] ), .Z(
        _f_permutation__round_out[1341]) );
  XOR2_X2 _f_permutation__round__U2825  ( .A(_f_permutation__round__N3075 ), 
        .B(_f_permutation__round__c[1584] ), .Z(
        _f_permutation__round_out[1342]) );
  XOR2_X2 _f_permutation__round__U2824  ( .A(_f_permutation__round__N3073 ), 
        .B(_f_permutation__round__c[1585] ), .Z(
        _f_permutation__round_out[1343]) );
  XOR2_X2 _f_permutation__round__U2823  ( .A(_f_permutation__round__N3071 ), 
        .B(_f_permutation__round__c[1195] ), .Z(
        _f_permutation__round_out[1344]) );
  XOR2_X2 _f_permutation__round__U2822  ( .A(_f_permutation__round__N3069 ), 
        .B(_f_permutation__round__c[1196] ), .Z(
        _f_permutation__round_out[1345]) );
  XOR2_X2 _f_permutation__round__U2821  ( .A(_f_permutation__round__N3067 ), 
        .B(_f_permutation__round__c[1197] ), .Z(
        _f_permutation__round_out[1346]) );
  XOR2_X2 _f_permutation__round__U2820  ( .A(_f_permutation__round__N3065 ), 
        .B(_f_permutation__round__c[1198] ), .Z(
        _f_permutation__round_out[1347]) );
  XOR2_X2 _f_permutation__round__U2819  ( .A(_f_permutation__round__N3063 ), 
        .B(_f_permutation__round__c[1199] ), .Z(
        _f_permutation__round_out[1348]) );
  XOR2_X2 _f_permutation__round__U2818  ( .A(_f_permutation__round__N3061 ), 
        .B(_f_permutation__round__c[1200] ), .Z(
        _f_permutation__round_out[1349]) );
  XOR2_X2 _f_permutation__round__U2817  ( .A(_f_permutation__round__N3059 ), 
        .B(_f_permutation__round__c[1201] ), .Z(
        _f_permutation__round_out[1350]) );
  XOR2_X2 _f_permutation__round__U2816  ( .A(_f_permutation__round__N3057 ), 
        .B(_f_permutation__round__c[1202] ), .Z(
        _f_permutation__round_out[1351]) );
  XOR2_X2 _f_permutation__round__U2815  ( .A(_f_permutation__round__N3055 ), 
        .B(_f_permutation__round__c[1203] ), .Z(
        _f_permutation__round_out[1352]) );
  XOR2_X2 _f_permutation__round__U2814  ( .A(_f_permutation__round__N3053 ), 
        .B(_f_permutation__round__c[1204] ), .Z(
        _f_permutation__round_out[1353]) );
  XOR2_X2 _f_permutation__round__U2813  ( .A(_f_permutation__round__N3051 ), 
        .B(_f_permutation__round__c[1205] ), .Z(
        _f_permutation__round_out[1354]) );
  XOR2_X2 _f_permutation__round__U2812  ( .A(_f_permutation__round__N3049 ), 
        .B(_f_permutation__round__c[1206] ), .Z(
        _f_permutation__round_out[1355]) );
  XOR2_X2 _f_permutation__round__U2811  ( .A(_f_permutation__round__N3047 ), 
        .B(_f_permutation__round__c[1207] ), .Z(
        _f_permutation__round_out[1356]) );
  XOR2_X2 _f_permutation__round__U2810  ( .A(_f_permutation__round__N3045 ), 
        .B(_f_permutation__round__c[1208] ), .Z(
        _f_permutation__round_out[1357]) );
  XOR2_X2 _f_permutation__round__U2809  ( .A(_f_permutation__round__N3043 ), 
        .B(_f_permutation__round__c[1209] ), .Z(
        _f_permutation__round_out[1358]) );
  XOR2_X2 _f_permutation__round__U2808  ( .A(_f_permutation__round__N3041 ), 
        .B(_f_permutation__round__c[1210] ), .Z(
        _f_permutation__round_out[1359]) );
  XOR2_X2 _f_permutation__round__U2807  ( .A(_f_permutation__round__N3039 ), 
        .B(_f_permutation__round__c[1211] ), .Z(
        _f_permutation__round_out[1360]) );
  XOR2_X2 _f_permutation__round__U2806  ( .A(_f_permutation__round__N3037 ), 
        .B(_f_permutation__round__c[1212] ), .Z(
        _f_permutation__round_out[1361]) );
  XOR2_X2 _f_permutation__round__U2805  ( .A(_f_permutation__round__N3035 ), 
        .B(_f_permutation__round__c[1213] ), .Z(
        _f_permutation__round_out[1362]) );
  XOR2_X2 _f_permutation__round__U2804  ( .A(_f_permutation__round__N3033 ), 
        .B(_f_permutation__round__c[1214] ), .Z(
        _f_permutation__round_out[1363]) );
  XOR2_X2 _f_permutation__round__U2803  ( .A(_f_permutation__round__N3031 ), 
        .B(_f_permutation__round__c[1215] ), .Z(
        _f_permutation__round_out[1364]) );
  XOR2_X2 _f_permutation__round__U2802  ( .A(_f_permutation__round__N3029 ), 
        .B(_f_permutation__round__c[1152] ), .Z(
        _f_permutation__round_out[1365]) );
  XOR2_X2 _f_permutation__round__U2801  ( .A(_f_permutation__round__N3027 ), 
        .B(_f_permutation__round__c[1153] ), .Z(
        _f_permutation__round_out[1366]) );
  XOR2_X2 _f_permutation__round__U2800  ( .A(_f_permutation__round__N3025 ), 
        .B(_f_permutation__round__c[1154] ), .Z(
        _f_permutation__round_out[1367]) );
  XOR2_X2 _f_permutation__round__U2799  ( .A(_f_permutation__round__N3023 ), 
        .B(_f_permutation__round__c[1155] ), .Z(
        _f_permutation__round_out[1368]) );
  XOR2_X2 _f_permutation__round__U2798  ( .A(_f_permutation__round__N3021 ), 
        .B(_f_permutation__round__c[1156] ), .Z(
        _f_permutation__round_out[1369]) );
  XOR2_X2 _f_permutation__round__U2797  ( .A(_f_permutation__round__N3019 ), 
        .B(_f_permutation__round__c[1157] ), .Z(
        _f_permutation__round_out[1370]) );
  XOR2_X2 _f_permutation__round__U2796  ( .A(_f_permutation__round__N3017 ), 
        .B(_f_permutation__round__c[1158] ), .Z(
        _f_permutation__round_out[1371]) );
  XOR2_X2 _f_permutation__round__U2795  ( .A(_f_permutation__round__N3015 ), 
        .B(_f_permutation__round__c[1159] ), .Z(
        _f_permutation__round_out[1372]) );
  XOR2_X2 _f_permutation__round__U2794  ( .A(_f_permutation__round__N3013 ), 
        .B(_f_permutation__round__c[1160] ), .Z(
        _f_permutation__round_out[1373]) );
  XOR2_X2 _f_permutation__round__U2793  ( .A(_f_permutation__round__N3011 ), 
        .B(_f_permutation__round__c[1161] ), .Z(
        _f_permutation__round_out[1374]) );
  XOR2_X2 _f_permutation__round__U2792  ( .A(_f_permutation__round__N3009 ), 
        .B(_f_permutation__round__c[1162] ), .Z(
        _f_permutation__round_out[1375]) );
  XOR2_X2 _f_permutation__round__U2791  ( .A(_f_permutation__round__N3007 ), 
        .B(_f_permutation__round__c[1163] ), .Z(
        _f_permutation__round_out[1376]) );
  XOR2_X2 _f_permutation__round__U2790  ( .A(_f_permutation__round__N3005 ), 
        .B(_f_permutation__round__c[1164] ), .Z(
        _f_permutation__round_out[1377]) );
  XOR2_X2 _f_permutation__round__U2789  ( .A(_f_permutation__round__N3003 ), 
        .B(_f_permutation__round__c[1165] ), .Z(
        _f_permutation__round_out[1378]) );
  XOR2_X2 _f_permutation__round__U2788  ( .A(_f_permutation__round__N3001 ), 
        .B(_f_permutation__round__c[1166] ), .Z(
        _f_permutation__round_out[1379]) );
  XOR2_X2 _f_permutation__round__U2787  ( .A(_f_permutation__round__N2999 ), 
        .B(_f_permutation__round__c[1167] ), .Z(
        _f_permutation__round_out[1380]) );
  XOR2_X2 _f_permutation__round__U2786  ( .A(_f_permutation__round__N2997 ), 
        .B(_f_permutation__round__c[1168] ), .Z(
        _f_permutation__round_out[1381]) );
  XOR2_X2 _f_permutation__round__U2785  ( .A(_f_permutation__round__N2995 ), 
        .B(_f_permutation__round__c[1169] ), .Z(
        _f_permutation__round_out[1382]) );
  XOR2_X2 _f_permutation__round__U2784  ( .A(_f_permutation__round__N2993 ), 
        .B(_f_permutation__round__c[1170] ), .Z(
        _f_permutation__round_out[1383]) );
  XOR2_X2 _f_permutation__round__U2783  ( .A(_f_permutation__round__N2991 ), 
        .B(_f_permutation__round__c[1171] ), .Z(
        _f_permutation__round_out[1384]) );
  XOR2_X2 _f_permutation__round__U2782  ( .A(_f_permutation__round__N2989 ), 
        .B(_f_permutation__round__c[1172] ), .Z(
        _f_permutation__round_out[1385]) );
  XOR2_X2 _f_permutation__round__U2781  ( .A(_f_permutation__round__N2987 ), 
        .B(_f_permutation__round__c[1173] ), .Z(
        _f_permutation__round_out[1386]) );
  XOR2_X2 _f_permutation__round__U2780  ( .A(_f_permutation__round__N2985 ), 
        .B(_f_permutation__round__c[1174] ), .Z(
        _f_permutation__round_out[1387]) );
  XOR2_X2 _f_permutation__round__U2779  ( .A(_f_permutation__round__N2983 ), 
        .B(_f_permutation__round__c[1175] ), .Z(
        _f_permutation__round_out[1388]) );
  XOR2_X2 _f_permutation__round__U2778  ( .A(_f_permutation__round__N2981 ), 
        .B(_f_permutation__round__c[1176] ), .Z(
        _f_permutation__round_out[1389]) );
  XOR2_X2 _f_permutation__round__U2777  ( .A(_f_permutation__round__N2979 ), 
        .B(_f_permutation__round__c[1177] ), .Z(
        _f_permutation__round_out[1390]) );
  XOR2_X2 _f_permutation__round__U2776  ( .A(_f_permutation__round__N2977 ), 
        .B(_f_permutation__round__c[1178] ), .Z(
        _f_permutation__round_out[1391]) );
  XOR2_X2 _f_permutation__round__U2775  ( .A(_f_permutation__round__N2975 ), 
        .B(_f_permutation__round__c[1179] ), .Z(
        _f_permutation__round_out[1392]) );
  XOR2_X2 _f_permutation__round__U2774  ( .A(_f_permutation__round__N2973 ), 
        .B(_f_permutation__round__c[1180] ), .Z(
        _f_permutation__round_out[1393]) );
  XOR2_X2 _f_permutation__round__U2773  ( .A(_f_permutation__round__N2971 ), 
        .B(_f_permutation__round__c[1181] ), .Z(
        _f_permutation__round_out[1394]) );
  XOR2_X2 _f_permutation__round__U2772  ( .A(_f_permutation__round__N2969 ), 
        .B(_f_permutation__round__c[1182] ), .Z(
        _f_permutation__round_out[1395]) );
  XOR2_X2 _f_permutation__round__U2771  ( .A(_f_permutation__round__N2967 ), 
        .B(_f_permutation__round__c[1183] ), .Z(
        _f_permutation__round_out[1396]) );
  XOR2_X2 _f_permutation__round__U2770  ( .A(_f_permutation__round__N2965 ), 
        .B(_f_permutation__round__c[1184] ), .Z(
        _f_permutation__round_out[1397]) );
  XOR2_X2 _f_permutation__round__U2769  ( .A(_f_permutation__round__N2963 ), 
        .B(_f_permutation__round__c[1185] ), .Z(
        _f_permutation__round_out[1398]) );
  XOR2_X2 _f_permutation__round__U2768  ( .A(_f_permutation__round__N2961 ), 
        .B(_f_permutation__round__c[1186] ), .Z(
        _f_permutation__round_out[1399]) );
  XOR2_X2 _f_permutation__round__U2767  ( .A(_f_permutation__round__N2959 ), 
        .B(_f_permutation__round__c[1187] ), .Z(
        _f_permutation__round_out[1400]) );
  XOR2_X2 _f_permutation__round__U2766  ( .A(_f_permutation__round__N2957 ), 
        .B(_f_permutation__round__c[1188] ), .Z(
        _f_permutation__round_out[1401]) );
  XOR2_X2 _f_permutation__round__U2765  ( .A(_f_permutation__round__N2955 ), 
        .B(_f_permutation__round__c[1189] ), .Z(
        _f_permutation__round_out[1402]) );
  XOR2_X2 _f_permutation__round__U2764  ( .A(_f_permutation__round__N2953 ), 
        .B(_f_permutation__round__c[1190] ), .Z(
        _f_permutation__round_out[1403]) );
  XOR2_X2 _f_permutation__round__U2763  ( .A(_f_permutation__round__N2951 ), 
        .B(_f_permutation__round__c[1191] ), .Z(
        _f_permutation__round_out[1404]) );
  XOR2_X2 _f_permutation__round__U2762  ( .A(_f_permutation__round__N2949 ), 
        .B(_f_permutation__round__c[1192] ), .Z(
        _f_permutation__round_out[1405]) );
  XOR2_X2 _f_permutation__round__U2761  ( .A(_f_permutation__round__N2947 ), 
        .B(_f_permutation__round__c[1193] ), .Z(
        _f_permutation__round_out[1406]) );
  XOR2_X2 _f_permutation__round__U2760  ( .A(_f_permutation__round__N2945 ), 
        .B(_f_permutation__round__c[1194] ), .Z(
        _f_permutation__round_out[1407]) );
  XOR2_X2 _f_permutation__round__U2759  ( .A(_f_permutation__round__N2943 ), 
        .B(_f_permutation__round__c[789] ), .Z(
        _f_permutation__round_out[1408]) );
  XOR2_X2 _f_permutation__round__U2758  ( .A(_f_permutation__round__N2941 ), 
        .B(_f_permutation__round__c[790] ), .Z(
        _f_permutation__round_out[1409]) );
  XOR2_X2 _f_permutation__round__U2757  ( .A(_f_permutation__round__N2939 ), 
        .B(_f_permutation__round__c[791] ), .Z(
        _f_permutation__round_out[1410]) );
  XOR2_X2 _f_permutation__round__U2756  ( .A(_f_permutation__round__N2937 ), 
        .B(_f_permutation__round__c[792] ), .Z(
        _f_permutation__round_out[1411]) );
  XOR2_X2 _f_permutation__round__U2755  ( .A(_f_permutation__round__N2935 ), 
        .B(_f_permutation__round__c[793] ), .Z(
        _f_permutation__round_out[1412]) );
  XOR2_X2 _f_permutation__round__U2754  ( .A(_f_permutation__round__N2933 ), 
        .B(_f_permutation__round__c[794] ), .Z(
        _f_permutation__round_out[1413]) );
  XOR2_X2 _f_permutation__round__U2753  ( .A(_f_permutation__round__N2931 ), 
        .B(_f_permutation__round__c[795] ), .Z(
        _f_permutation__round_out[1414]) );
  XOR2_X2 _f_permutation__round__U2752  ( .A(_f_permutation__round__N2929 ), 
        .B(_f_permutation__round__c[796] ), .Z(
        _f_permutation__round_out[1415]) );
  XOR2_X2 _f_permutation__round__U2751  ( .A(_f_permutation__round__N2927 ), 
        .B(_f_permutation__round__c[797] ), .Z(
        _f_permutation__round_out[1416]) );
  XOR2_X2 _f_permutation__round__U2750  ( .A(_f_permutation__round__N2925 ), 
        .B(_f_permutation__round__c[798] ), .Z(
        _f_permutation__round_out[1417]) );
  XOR2_X2 _f_permutation__round__U2749  ( .A(_f_permutation__round__N2923 ), 
        .B(_f_permutation__round__c[799] ), .Z(
        _f_permutation__round_out[1418]) );
  XOR2_X2 _f_permutation__round__U2748  ( .A(_f_permutation__round__N2921 ), 
        .B(_f_permutation__round__c[800] ), .Z(
        _f_permutation__round_out[1419]) );
  XOR2_X2 _f_permutation__round__U2747  ( .A(_f_permutation__round__N2919 ), 
        .B(_f_permutation__round__c[801] ), .Z(
        _f_permutation__round_out[1420]) );
  XOR2_X2 _f_permutation__round__U2746  ( .A(_f_permutation__round__N2917 ), 
        .B(_f_permutation__round__c[802] ), .Z(
        _f_permutation__round_out[1421]) );
  XOR2_X2 _f_permutation__round__U2745  ( .A(_f_permutation__round__N2915 ), 
        .B(_f_permutation__round__c[803] ), .Z(
        _f_permutation__round_out[1422]) );
  XOR2_X2 _f_permutation__round__U2744  ( .A(_f_permutation__round__N2913 ), 
        .B(_f_permutation__round__c[804] ), .Z(
        _f_permutation__round_out[1423]) );
  XOR2_X2 _f_permutation__round__U2743  ( .A(_f_permutation__round__N2911 ), 
        .B(_f_permutation__round__c[805] ), .Z(
        _f_permutation__round_out[1424]) );
  XOR2_X2 _f_permutation__round__U2742  ( .A(_f_permutation__round__N2909 ), 
        .B(_f_permutation__round__c[806] ), .Z(
        _f_permutation__round_out[1425]) );
  XOR2_X2 _f_permutation__round__U2741  ( .A(_f_permutation__round__N2907 ), 
        .B(_f_permutation__round__c[807] ), .Z(
        _f_permutation__round_out[1426]) );
  XOR2_X2 _f_permutation__round__U2740  ( .A(_f_permutation__round__N2905 ), 
        .B(_f_permutation__round__c[808] ), .Z(
        _f_permutation__round_out[1427]) );
  XOR2_X2 _f_permutation__round__U2739  ( .A(_f_permutation__round__N2903 ), 
        .B(_f_permutation__round__c[809] ), .Z(
        _f_permutation__round_out[1428]) );
  XOR2_X2 _f_permutation__round__U2738  ( .A(_f_permutation__round__N2901 ), 
        .B(_f_permutation__round__c[810] ), .Z(
        _f_permutation__round_out[1429]) );
  XOR2_X2 _f_permutation__round__U2737  ( .A(_f_permutation__round__N2899 ), 
        .B(_f_permutation__round__c[811] ), .Z(
        _f_permutation__round_out[1430]) );
  XOR2_X2 _f_permutation__round__U2736  ( .A(_f_permutation__round__N2897 ), 
        .B(_f_permutation__round__c[812] ), .Z(
        _f_permutation__round_out[1431]) );
  XOR2_X2 _f_permutation__round__U2735  ( .A(_f_permutation__round__N2895 ), 
        .B(_f_permutation__round__c[813] ), .Z(
        _f_permutation__round_out[1432]) );
  XOR2_X2 _f_permutation__round__U2734  ( .A(_f_permutation__round__N2893 ), 
        .B(_f_permutation__round__c[814] ), .Z(
        _f_permutation__round_out[1433]) );
  XOR2_X2 _f_permutation__round__U2733  ( .A(_f_permutation__round__N2891 ), 
        .B(_f_permutation__round__c[815] ), .Z(
        _f_permutation__round_out[1434]) );
  XOR2_X2 _f_permutation__round__U2732  ( .A(_f_permutation__round__N2889 ), 
        .B(_f_permutation__round__c[816] ), .Z(
        _f_permutation__round_out[1435]) );
  XOR2_X2 _f_permutation__round__U2731  ( .A(_f_permutation__round__N2887 ), 
        .B(_f_permutation__round__c[817] ), .Z(
        _f_permutation__round_out[1436]) );
  XOR2_X2 _f_permutation__round__U2730  ( .A(_f_permutation__round__N2885 ), 
        .B(_f_permutation__round__c[818] ), .Z(
        _f_permutation__round_out[1437]) );
  XOR2_X2 _f_permutation__round__U2729  ( .A(_f_permutation__round__N2883 ), 
        .B(_f_permutation__round__c[819] ), .Z(
        _f_permutation__round_out[1438]) );
  XOR2_X2 _f_permutation__round__U2728  ( .A(_f_permutation__round__N2881 ), 
        .B(_f_permutation__round__c[820] ), .Z(
        _f_permutation__round_out[1439]) );
  XOR2_X2 _f_permutation__round__U2727  ( .A(_f_permutation__round__N2879 ), 
        .B(_f_permutation__round__c[821] ), .Z(
        _f_permutation__round_out[1440]) );
  XOR2_X2 _f_permutation__round__U2726  ( .A(_f_permutation__round__N2877 ), 
        .B(_f_permutation__round__c[822] ), .Z(
        _f_permutation__round_out[1441]) );
  XOR2_X2 _f_permutation__round__U2725  ( .A(_f_permutation__round__N2875 ), 
        .B(_f_permutation__round__c[823] ), .Z(
        _f_permutation__round_out[1442]) );
  XOR2_X2 _f_permutation__round__U2724  ( .A(_f_permutation__round__N2873 ), 
        .B(_f_permutation__round__c[824] ), .Z(
        _f_permutation__round_out[1443]) );
  XOR2_X2 _f_permutation__round__U2723  ( .A(_f_permutation__round__N2871 ), 
        .B(_f_permutation__round__c[825] ), .Z(
        _f_permutation__round_out[1444]) );
  XOR2_X2 _f_permutation__round__U2722  ( .A(_f_permutation__round__N2869 ), 
        .B(_f_permutation__round__c[826] ), .Z(
        _f_permutation__round_out[1445]) );
  XOR2_X2 _f_permutation__round__U2721  ( .A(_f_permutation__round__N2867 ), 
        .B(_f_permutation__round__c[827] ), .Z(
        _f_permutation__round_out[1446]) );
  XOR2_X2 _f_permutation__round__U2720  ( .A(_f_permutation__round__N2865 ), 
        .B(_f_permutation__round__c[828] ), .Z(
        _f_permutation__round_out[1447]) );
  XOR2_X2 _f_permutation__round__U2719  ( .A(_f_permutation__round__N2863 ), 
        .B(_f_permutation__round__c[829] ), .Z(
        _f_permutation__round_out[1448]) );
  XOR2_X2 _f_permutation__round__U2718  ( .A(_f_permutation__round__N2861 ), 
        .B(_f_permutation__round__c[830] ), .Z(
        _f_permutation__round_out[1449]) );
  XOR2_X2 _f_permutation__round__U2717  ( .A(_f_permutation__round__N2859 ), 
        .B(_f_permutation__round__c[831] ), .Z(
        _f_permutation__round_out[1450]) );
  XOR2_X2 _f_permutation__round__U2716  ( .A(_f_permutation__round__N2857 ), 
        .B(_f_permutation__round__c[768] ), .Z(
        _f_permutation__round_out[1451]) );
  XOR2_X2 _f_permutation__round__U2715  ( .A(_f_permutation__round__N2855 ), 
        .B(_f_permutation__round__c[769] ), .Z(
        _f_permutation__round_out[1452]) );
  XOR2_X2 _f_permutation__round__U2714  ( .A(_f_permutation__round__N2853 ), 
        .B(_f_permutation__round__c[770] ), .Z(
        _f_permutation__round_out[1453]) );
  XOR2_X2 _f_permutation__round__U2713  ( .A(_f_permutation__round__N2851 ), 
        .B(_f_permutation__round__c[771] ), .Z(
        _f_permutation__round_out[1454]) );
  XOR2_X2 _f_permutation__round__U2712  ( .A(_f_permutation__round__N2849 ), 
        .B(_f_permutation__round__c[772] ), .Z(
        _f_permutation__round_out[1455]) );
  XOR2_X2 _f_permutation__round__U2711  ( .A(_f_permutation__round__N2847 ), 
        .B(_f_permutation__round__c[773] ), .Z(
        _f_permutation__round_out[1456]) );
  XOR2_X2 _f_permutation__round__U2710  ( .A(_f_permutation__round__N2845 ), 
        .B(_f_permutation__round__c[774] ), .Z(
        _f_permutation__round_out[1457]) );
  XOR2_X2 _f_permutation__round__U2709  ( .A(_f_permutation__round__N2843 ), 
        .B(_f_permutation__round__c[775] ), .Z(
        _f_permutation__round_out[1458]) );
  XOR2_X2 _f_permutation__round__U2708  ( .A(_f_permutation__round__N2841 ), 
        .B(_f_permutation__round__c[776] ), .Z(
        _f_permutation__round_out[1459]) );
  XOR2_X2 _f_permutation__round__U2707  ( .A(_f_permutation__round__N2839 ), 
        .B(_f_permutation__round__c[777] ), .Z(
        _f_permutation__round_out[1460]) );
  XOR2_X2 _f_permutation__round__U2706  ( .A(_f_permutation__round__N2837 ), 
        .B(_f_permutation__round__c[778] ), .Z(
        _f_permutation__round_out[1461]) );
  XOR2_X2 _f_permutation__round__U2705  ( .A(_f_permutation__round__N2835 ), 
        .B(_f_permutation__round__c[779] ), .Z(
        _f_permutation__round_out[1462]) );
  XOR2_X2 _f_permutation__round__U2704  ( .A(_f_permutation__round__N2833 ), 
        .B(_f_permutation__round__c[780] ), .Z(
        _f_permutation__round_out[1463]) );
  XOR2_X2 _f_permutation__round__U2703  ( .A(_f_permutation__round__N2831 ), 
        .B(_f_permutation__round__c[781] ), .Z(
        _f_permutation__round_out[1464]) );
  XOR2_X2 _f_permutation__round__U2702  ( .A(_f_permutation__round__N2829 ), 
        .B(_f_permutation__round__c[782] ), .Z(
        _f_permutation__round_out[1465]) );
  XOR2_X2 _f_permutation__round__U2701  ( .A(_f_permutation__round__N2827 ), 
        .B(_f_permutation__round__c[783] ), .Z(
        _f_permutation__round_out[1466]) );
  XOR2_X2 _f_permutation__round__U2700  ( .A(_f_permutation__round__N2825 ), 
        .B(_f_permutation__round__c[784] ), .Z(
        _f_permutation__round_out[1467]) );
  XOR2_X2 _f_permutation__round__U2699  ( .A(_f_permutation__round__N2823 ), 
        .B(_f_permutation__round__c[785] ), .Z(
        _f_permutation__round_out[1468]) );
  XOR2_X2 _f_permutation__round__U2698  ( .A(_f_permutation__round__N2821 ), 
        .B(_f_permutation__round__c[786] ), .Z(
        _f_permutation__round_out[1469]) );
  XOR2_X2 _f_permutation__round__U2697  ( .A(_f_permutation__round__N2819 ), 
        .B(_f_permutation__round__c[787] ), .Z(
        _f_permutation__round_out[1470]) );
  XOR2_X2 _f_permutation__round__U2696  ( .A(_f_permutation__round__N2817 ), 
        .B(_f_permutation__round__c[788] ), .Z(
        _f_permutation__round_out[1471]) );
  XOR2_X2 _f_permutation__round__U2695  ( .A(_f_permutation__round__N2815 ), 
        .B(_f_permutation__round__c[404] ), .Z(
        _f_permutation__round_out[1472]) );
  XOR2_X2 _f_permutation__round__U2694  ( .A(_f_permutation__round__N2813 ), 
        .B(_f_permutation__round__c[405] ), .Z(
        _f_permutation__round_out[1473]) );
  XOR2_X2 _f_permutation__round__U2693  ( .A(_f_permutation__round__N2811 ), 
        .B(_f_permutation__round__c[406] ), .Z(
        _f_permutation__round_out[1474]) );
  XOR2_X2 _f_permutation__round__U2692  ( .A(_f_permutation__round__N2809 ), 
        .B(_f_permutation__round__c[407] ), .Z(
        _f_permutation__round_out[1475]) );
  XOR2_X2 _f_permutation__round__U2691  ( .A(_f_permutation__round__N2807 ), 
        .B(_f_permutation__round__c[408] ), .Z(
        _f_permutation__round_out[1476]) );
  XOR2_X2 _f_permutation__round__U2690  ( .A(_f_permutation__round__N2805 ), 
        .B(_f_permutation__round__c[409] ), .Z(
        _f_permutation__round_out[1477]) );
  XOR2_X2 _f_permutation__round__U2689  ( .A(_f_permutation__round__N2803 ), 
        .B(_f_permutation__round__c[410] ), .Z(
        _f_permutation__round_out[1478]) );
  XOR2_X2 _f_permutation__round__U2688  ( .A(_f_permutation__round__N2801 ), 
        .B(_f_permutation__round__c[411] ), .Z(
        _f_permutation__round_out[1479]) );
  XOR2_X2 _f_permutation__round__U2687  ( .A(_f_permutation__round__N2799 ), 
        .B(_f_permutation__round__c[412] ), .Z(
        _f_permutation__round_out[1480]) );
  XOR2_X2 _f_permutation__round__U2686  ( .A(_f_permutation__round__N2797 ), 
        .B(_f_permutation__round__c[413] ), .Z(
        _f_permutation__round_out[1481]) );
  XOR2_X2 _f_permutation__round__U2685  ( .A(_f_permutation__round__N2795 ), 
        .B(_f_permutation__round__c[414] ), .Z(
        _f_permutation__round_out[1482]) );
  XOR2_X2 _f_permutation__round__U2684  ( .A(_f_permutation__round__N2793 ), 
        .B(_f_permutation__round__c[415] ), .Z(
        _f_permutation__round_out[1483]) );
  XOR2_X2 _f_permutation__round__U2683  ( .A(_f_permutation__round__N2791 ), 
        .B(_f_permutation__round__c[416] ), .Z(
        _f_permutation__round_out[1484]) );
  XOR2_X2 _f_permutation__round__U2682  ( .A(_f_permutation__round__N2789 ), 
        .B(_f_permutation__round__c[417] ), .Z(
        _f_permutation__round_out[1485]) );
  XOR2_X2 _f_permutation__round__U2681  ( .A(_f_permutation__round__N2787 ), 
        .B(_f_permutation__round__c[418] ), .Z(
        _f_permutation__round_out[1486]) );
  XOR2_X2 _f_permutation__round__U2680  ( .A(_f_permutation__round__N2785 ), 
        .B(_f_permutation__round__c[419] ), .Z(
        _f_permutation__round_out[1487]) );
  XOR2_X2 _f_permutation__round__U2679  ( .A(_f_permutation__round__N2783 ), 
        .B(_f_permutation__round__c[420] ), .Z(
        _f_permutation__round_out[1488]) );
  XOR2_X2 _f_permutation__round__U2678  ( .A(_f_permutation__round__N2781 ), 
        .B(_f_permutation__round__c[421] ), .Z(
        _f_permutation__round_out[1489]) );
  XOR2_X2 _f_permutation__round__U2677  ( .A(_f_permutation__round__N2779 ), 
        .B(_f_permutation__round__c[422] ), .Z(
        _f_permutation__round_out[1490]) );
  XOR2_X2 _f_permutation__round__U2676  ( .A(_f_permutation__round__N2777 ), 
        .B(_f_permutation__round__c[423] ), .Z(
        _f_permutation__round_out[1491]) );
  XOR2_X2 _f_permutation__round__U2675  ( .A(_f_permutation__round__N2775 ), 
        .B(_f_permutation__round__c[424] ), .Z(
        _f_permutation__round_out[1492]) );
  XOR2_X2 _f_permutation__round__U2674  ( .A(_f_permutation__round__N2773 ), 
        .B(_f_permutation__round__c[425] ), .Z(
        _f_permutation__round_out[1493]) );
  XOR2_X2 _f_permutation__round__U2673  ( .A(_f_permutation__round__N2771 ), 
        .B(_f_permutation__round__c[426] ), .Z(
        _f_permutation__round_out[1494]) );
  XOR2_X2 _f_permutation__round__U2672  ( .A(_f_permutation__round__N2769 ), 
        .B(_f_permutation__round__c[427] ), .Z(
        _f_permutation__round_out[1495]) );
  XOR2_X2 _f_permutation__round__U2671  ( .A(_f_permutation__round__N2767 ), 
        .B(_f_permutation__round__c[428] ), .Z(
        _f_permutation__round_out[1496]) );
  XOR2_X2 _f_permutation__round__U2670  ( .A(_f_permutation__round__N2765 ), 
        .B(_f_permutation__round__c[429] ), .Z(
        _f_permutation__round_out[1497]) );
  XOR2_X2 _f_permutation__round__U2669  ( .A(_f_permutation__round__N2763 ), 
        .B(_f_permutation__round__c[430] ), .Z(
        _f_permutation__round_out[1498]) );
  XOR2_X2 _f_permutation__round__U2668  ( .A(_f_permutation__round__N2761 ), 
        .B(_f_permutation__round__c[431] ), .Z(
        _f_permutation__round_out[1499]) );
  XOR2_X2 _f_permutation__round__U2667  ( .A(_f_permutation__round__N2759 ), 
        .B(_f_permutation__round__c[432] ), .Z(
        _f_permutation__round_out[1500]) );
  XOR2_X2 _f_permutation__round__U2666  ( .A(_f_permutation__round__N2757 ), 
        .B(_f_permutation__round__c[433] ), .Z(
        _f_permutation__round_out[1501]) );
  XOR2_X2 _f_permutation__round__U2665  ( .A(_f_permutation__round__N2755 ), 
        .B(_f_permutation__round__c[434] ), .Z(
        _f_permutation__round_out[1502]) );
  XOR2_X2 _f_permutation__round__U2664  ( .A(_f_permutation__round__N2753 ), 
        .B(_f_permutation__round__c[435] ), .Z(
        _f_permutation__round_out[1503]) );
  XOR2_X2 _f_permutation__round__U2663  ( .A(_f_permutation__round__N2751 ), 
        .B(_f_permutation__round__c[436] ), .Z(
        _f_permutation__round_out[1504]) );
  XOR2_X2 _f_permutation__round__U2662  ( .A(_f_permutation__round__N2749 ), 
        .B(_f_permutation__round__c[437] ), .Z(
        _f_permutation__round_out[1505]) );
  XOR2_X2 _f_permutation__round__U2661  ( .A(_f_permutation__round__N2747 ), 
        .B(_f_permutation__round__c[438] ), .Z(
        _f_permutation__round_out[1506]) );
  XOR2_X2 _f_permutation__round__U2660  ( .A(_f_permutation__round__N2745 ), 
        .B(_f_permutation__round__c[439] ), .Z(
        _f_permutation__round_out[1507]) );
  XOR2_X2 _f_permutation__round__U2659  ( .A(_f_permutation__round__N2743 ), 
        .B(_f_permutation__round__c[440] ), .Z(
        _f_permutation__round_out[1508]) );
  XOR2_X2 _f_permutation__round__U2658  ( .A(_f_permutation__round__N2741 ), 
        .B(_f_permutation__round__c[441] ), .Z(
        _f_permutation__round_out[1509]) );
  XOR2_X2 _f_permutation__round__U2657  ( .A(_f_permutation__round__N2739 ), 
        .B(_f_permutation__round__c[442] ), .Z(
        _f_permutation__round_out[1510]) );
  XOR2_X2 _f_permutation__round__U2656  ( .A(_f_permutation__round__N2737 ), 
        .B(_f_permutation__round__c[443] ), .Z(
        _f_permutation__round_out[1511]) );
  XOR2_X2 _f_permutation__round__U2655  ( .A(_f_permutation__round__N2735 ), 
        .B(_f_permutation__round__c[444] ), .Z(
        _f_permutation__round_out[1512]) );
  XOR2_X2 _f_permutation__round__U2654  ( .A(_f_permutation__round__N2733 ), 
        .B(_f_permutation__round__c[445] ), .Z(
        _f_permutation__round_out[1513]) );
  XOR2_X2 _f_permutation__round__U2653  ( .A(_f_permutation__round__N2731 ), 
        .B(_f_permutation__round__c[446] ), .Z(
        _f_permutation__round_out[1514]) );
  XOR2_X2 _f_permutation__round__U2652  ( .A(_f_permutation__round__N2729 ), 
        .B(_f_permutation__round__c[447] ), .Z(
        _f_permutation__round_out[1515]) );
  XOR2_X2 _f_permutation__round__U2651  ( .A(_f_permutation__round__N2727 ), 
        .B(_f_permutation__round__c[384] ), .Z(
        _f_permutation__round_out[1516]) );
  XOR2_X2 _f_permutation__round__U2650  ( .A(_f_permutation__round__N2725 ), 
        .B(_f_permutation__round__c[385] ), .Z(
        _f_permutation__round_out[1517]) );
  XOR2_X2 _f_permutation__round__U2649  ( .A(_f_permutation__round__N2723 ), 
        .B(_f_permutation__round__c[386] ), .Z(
        _f_permutation__round_out[1518]) );
  XOR2_X2 _f_permutation__round__U2648  ( .A(_f_permutation__round__N2721 ), 
        .B(_f_permutation__round__c[387] ), .Z(
        _f_permutation__round_out[1519]) );
  XOR2_X2 _f_permutation__round__U2647  ( .A(_f_permutation__round__N2719 ), 
        .B(_f_permutation__round__c[388] ), .Z(
        _f_permutation__round_out[1520]) );
  XOR2_X2 _f_permutation__round__U2646  ( .A(_f_permutation__round__N2717 ), 
        .B(_f_permutation__round__c[389] ), .Z(
        _f_permutation__round_out[1521]) );
  XOR2_X2 _f_permutation__round__U2645  ( .A(_f_permutation__round__N2715 ), 
        .B(_f_permutation__round__c[390] ), .Z(
        _f_permutation__round_out[1522]) );
  XOR2_X2 _f_permutation__round__U2644  ( .A(_f_permutation__round__N2713 ), 
        .B(_f_permutation__round__c[391] ), .Z(
        _f_permutation__round_out[1523]) );
  XOR2_X2 _f_permutation__round__U2643  ( .A(_f_permutation__round__N2711 ), 
        .B(_f_permutation__round__c[392] ), .Z(
        _f_permutation__round_out[1524]) );
  XOR2_X2 _f_permutation__round__U2642  ( .A(_f_permutation__round__N2709 ), 
        .B(_f_permutation__round__c[393] ), .Z(
        _f_permutation__round_out[1525]) );
  XOR2_X2 _f_permutation__round__U2641  ( .A(_f_permutation__round__N2707 ), 
        .B(_f_permutation__round__c[394] ), .Z(
        _f_permutation__round_out[1526]) );
  XOR2_X2 _f_permutation__round__U2640  ( .A(_f_permutation__round__N2705 ), 
        .B(_f_permutation__round__c[395] ), .Z(
        _f_permutation__round_out[1527]) );
  XOR2_X2 _f_permutation__round__U2639  ( .A(_f_permutation__round__N2703 ), 
        .B(_f_permutation__round__c[396] ), .Z(
        _f_permutation__round_out[1528]) );
  XOR2_X2 _f_permutation__round__U2638  ( .A(_f_permutation__round__N2701 ), 
        .B(_f_permutation__round__c[397] ), .Z(
        _f_permutation__round_out[1529]) );
  XOR2_X2 _f_permutation__round__U2637  ( .A(_f_permutation__round__N2699 ), 
        .B(_f_permutation__round__c[398] ), .Z(
        _f_permutation__round_out[1530]) );
  XOR2_X2 _f_permutation__round__U2636  ( .A(_f_permutation__round__N2697 ), 
        .B(_f_permutation__round__c[399] ), .Z(
        _f_permutation__round_out[1531]) );
  XOR2_X2 _f_permutation__round__U2635  ( .A(_f_permutation__round__N2695 ), 
        .B(_f_permutation__round__c[400] ), .Z(
        _f_permutation__round_out[1532]) );
  XOR2_X2 _f_permutation__round__U2634  ( .A(_f_permutation__round__N2693 ), 
        .B(_f_permutation__round__c[401] ), .Z(
        _f_permutation__round_out[1533]) );
  XOR2_X2 _f_permutation__round__U2633  ( .A(_f_permutation__round__N2691 ), 
        .B(_f_permutation__round__c[402] ), .Z(
        _f_permutation__round_out[1534]) );
  XOR2_X2 _f_permutation__round__U2632  ( .A(_f_permutation__round__N2689 ), 
        .B(_f_permutation__round__c[403] ), .Z(
        _f_permutation__round_out[1535]) );
  XOR2_X2 _f_permutation__round__U2631  ( .A(_f_permutation__round__c[0] ), 
        .B(_f_permutation__round__n1921 ), .Z(_f_permutation__round_out[1536]) );
  XOR2_X2 _f_permutation__round__U2630  ( .A(_f_permutation__round__N2687 ), 
        .B(_f_permutation__rc[0]), .Z(_f_permutation__round__n1921 ) );
  XOR2_X2 _f_permutation__round__U2629  ( .A(_f_permutation__round__c[1] ), 
        .B(_f_permutation__round__n1922 ), .Z(_f_permutation__round_out[1537]) );
  XOR2_X2 _f_permutation__round__U2628  ( .A(_f_permutation__round__N2685 ), 
        .B(_f_permutation__rc[1]), .Z(_f_permutation__round__n1922 ) );
  XOR2_X2 _f_permutation__round__U2627  ( .A(_f_permutation__round__N2683 ), 
        .B(_f_permutation__round__c[2] ), .Z(_f_permutation__round_out[1538])
         );
  XOR2_X2 _f_permutation__round__U2626  ( .A(_f_permutation__round__c[3] ), 
        .B(_f_permutation__round__n1923 ), .Z(_f_permutation__round_out[1539]) );
  XOR2_X2 _f_permutation__round__U2625  ( .A(_f_permutation__round__N2681 ), 
        .B(_f_permutation__rc[3]), .Z(_f_permutation__round__n1923 ) );
  XOR2_X2 _f_permutation__round__U2624  ( .A(_f_permutation__round__N2679 ), 
        .B(_f_permutation__round__c[4] ), .Z(_f_permutation__round_out[1540])
         );
  XOR2_X2 _f_permutation__round__U2623  ( .A(_f_permutation__round__N2677 ), 
        .B(_f_permutation__round__c[5] ), .Z(_f_permutation__round_out[1541])
         );
  XOR2_X2 _f_permutation__round__U2622  ( .A(_f_permutation__round__N2675 ), 
        .B(_f_permutation__round__c[6] ), .Z(_f_permutation__round_out[1542])
         );
  XOR2_X2 _f_permutation__round__U2621  ( .A(_f_permutation__round__c[7] ), 
        .B(_f_permutation__round__n1924 ), .Z(_f_permutation__round_out[1543]) );
  XOR2_X2 _f_permutation__round__U2620  ( .A(_f_permutation__round__N2673 ), 
        .B(_f_permutation__rc[7]), .Z(_f_permutation__round__n1924 ) );
  XOR2_X2 _f_permutation__round__U2619  ( .A(_f_permutation__round__N2671 ), 
        .B(_f_permutation__round__c[8] ), .Z(_f_permutation__round_out[1544])
         );
  XOR2_X2 _f_permutation__round__U2618  ( .A(_f_permutation__round__N2669 ), 
        .B(_f_permutation__round__c[9] ), .Z(_f_permutation__round_out[1545])
         );
  XOR2_X2 _f_permutation__round__U2617  ( .A(_f_permutation__round__N2667 ), 
        .B(_f_permutation__round__c[10] ), .Z(_f_permutation__round_out[1546]) );
  XOR2_X2 _f_permutation__round__U2616  ( .A(_f_permutation__round__N2665 ), 
        .B(_f_permutation__round__c[11] ), .Z(_f_permutation__round_out[1547]) );
  XOR2_X2 _f_permutation__round__U2615  ( .A(_f_permutation__round__N2663 ), 
        .B(_f_permutation__round__c[12] ), .Z(_f_permutation__round_out[1548]) );
  XOR2_X2 _f_permutation__round__U2614  ( .A(_f_permutation__round__N2661 ), 
        .B(_f_permutation__round__c[13] ), .Z(_f_permutation__round_out[1549]) );
  XOR2_X2 _f_permutation__round__U2613  ( .A(_f_permutation__round__N2659 ), 
        .B(_f_permutation__round__c[14] ), .Z(_f_permutation__round_out[1550]) );
  XOR2_X2 _f_permutation__round__U2612  ( .A(_f_permutation__round__c[15] ), 
        .B(_f_permutation__round__n1925 ), .Z(_f_permutation__round_out[1551]) );
  XOR2_X2 _f_permutation__round__U2611  ( .A(_f_permutation__round__N2657 ), 
        .B(_f_permutation__rc[15]), .Z(_f_permutation__round__n1925 ) );
  XOR2_X2 _f_permutation__round__U2610  ( .A(_f_permutation__round__N2655 ), 
        .B(_f_permutation__round__c[16] ), .Z(_f_permutation__round_out[1552]) );
  XOR2_X2 _f_permutation__round__U2609  ( .A(_f_permutation__round__N2653 ), 
        .B(_f_permutation__round__c[17] ), .Z(_f_permutation__round_out[1553]) );
  XOR2_X2 _f_permutation__round__U2608  ( .A(_f_permutation__round__N2651 ), 
        .B(_f_permutation__round__c[18] ), .Z(_f_permutation__round_out[1554]) );
  XOR2_X2 _f_permutation__round__U2607  ( .A(_f_permutation__round__N2649 ), 
        .B(_f_permutation__round__c[19] ), .Z(_f_permutation__round_out[1555]) );
  XOR2_X2 _f_permutation__round__U2606  ( .A(_f_permutation__round__N2647 ), 
        .B(_f_permutation__round__c[20] ), .Z(_f_permutation__round_out[1556]) );
  XOR2_X2 _f_permutation__round__U2605  ( .A(_f_permutation__round__N2645 ), 
        .B(_f_permutation__round__c[21] ), .Z(_f_permutation__round_out[1557]) );
  XOR2_X2 _f_permutation__round__U2604  ( .A(_f_permutation__round__N2643 ), 
        .B(_f_permutation__round__c[22] ), .Z(_f_permutation__round_out[1558]) );
  XOR2_X2 _f_permutation__round__U2603  ( .A(_f_permutation__round__N2641 ), 
        .B(_f_permutation__round__c[23] ), .Z(_f_permutation__round_out[1559]) );
  XOR2_X2 _f_permutation__round__U2602  ( .A(_f_permutation__round__N2639 ), 
        .B(_f_permutation__round__c[24] ), .Z(_f_permutation__round_out[1560]) );
  XOR2_X2 _f_permutation__round__U2601  ( .A(_f_permutation__round__N2637 ), 
        .B(_f_permutation__round__c[25] ), .Z(_f_permutation__round_out[1561]) );
  XOR2_X2 _f_permutation__round__U2600  ( .A(_f_permutation__round__N2635 ), 
        .B(_f_permutation__round__c[26] ), .Z(_f_permutation__round_out[1562]) );
  XOR2_X2 _f_permutation__round__U2599  ( .A(_f_permutation__round__N2633 ), 
        .B(_f_permutation__round__c[27] ), .Z(_f_permutation__round_out[1563]) );
  XOR2_X2 _f_permutation__round__U2598  ( .A(_f_permutation__round__N2631 ), 
        .B(_f_permutation__round__c[28] ), .Z(_f_permutation__round_out[1564]) );
  XOR2_X2 _f_permutation__round__U2597  ( .A(_f_permutation__round__N2629 ), 
        .B(_f_permutation__round__c[29] ), .Z(_f_permutation__round_out[1565]) );
  XOR2_X2 _f_permutation__round__U2596  ( .A(_f_permutation__round__N2627 ), 
        .B(_f_permutation__round__c[30] ), .Z(_f_permutation__round_out[1566]) );
  XOR2_X2 _f_permutation__round__U2595  ( .A(_f_permutation__round__c[31] ), 
        .B(_f_permutation__round__n1926 ), .Z(_f_permutation__round_out[1567]) );
  XOR2_X2 _f_permutation__round__U2594  ( .A(_f_permutation__round__N2625 ), 
        .B(_f_permutation__rc[31]), .Z(_f_permutation__round__n1926 ) );
  XOR2_X2 _f_permutation__round__U2593  ( .A(_f_permutation__round__N2623 ), 
        .B(_f_permutation__round__c[32] ), .Z(_f_permutation__round_out[1568]) );
  XOR2_X2 _f_permutation__round__U2592  ( .A(_f_permutation__round__N2621 ), 
        .B(_f_permutation__round__c[33] ), .Z(_f_permutation__round_out[1569]) );
  XOR2_X2 _f_permutation__round__U2591  ( .A(_f_permutation__round__N2619 ), 
        .B(_f_permutation__round__c[34] ), .Z(_f_permutation__round_out[1570]) );
  XOR2_X2 _f_permutation__round__U2590  ( .A(_f_permutation__round__N2617 ), 
        .B(_f_permutation__round__c[35] ), .Z(_f_permutation__round_out[1571]) );
  XOR2_X2 _f_permutation__round__U2589  ( .A(_f_permutation__round__N2615 ), 
        .B(_f_permutation__round__c[36] ), .Z(_f_permutation__round_out[1572]) );
  XOR2_X2 _f_permutation__round__U2588  ( .A(_f_permutation__round__N2613 ), 
        .B(_f_permutation__round__c[37] ), .Z(_f_permutation__round_out[1573]) );
  XOR2_X2 _f_permutation__round__U2587  ( .A(_f_permutation__round__N2611 ), 
        .B(_f_permutation__round__c[38] ), .Z(_f_permutation__round_out[1574]) );
  XOR2_X2 _f_permutation__round__U2586  ( .A(_f_permutation__round__N2609 ), 
        .B(_f_permutation__round__c[39] ), .Z(_f_permutation__round_out[1575]) );
  XOR2_X2 _f_permutation__round__U2585  ( .A(_f_permutation__round__N2607 ), 
        .B(_f_permutation__round__c[40] ), .Z(_f_permutation__round_out[1576]) );
  XOR2_X2 _f_permutation__round__U2584  ( .A(_f_permutation__round__N2605 ), 
        .B(_f_permutation__round__c[41] ), .Z(_f_permutation__round_out[1577]) );
  XOR2_X2 _f_permutation__round__U2583  ( .A(_f_permutation__round__N2603 ), 
        .B(_f_permutation__round__c[42] ), .Z(_f_permutation__round_out[1578]) );
  XOR2_X2 _f_permutation__round__U2582  ( .A(_f_permutation__round__N2601 ), 
        .B(_f_permutation__round__c[43] ), .Z(_f_permutation__round_out[1579]) );
  XOR2_X2 _f_permutation__round__U2581  ( .A(_f_permutation__round__N2599 ), 
        .B(_f_permutation__round__c[44] ), .Z(_f_permutation__round_out[1580]) );
  XOR2_X2 _f_permutation__round__U2580  ( .A(_f_permutation__round__N2597 ), 
        .B(_f_permutation__round__c[45] ), .Z(_f_permutation__round_out[1581]) );
  XOR2_X2 _f_permutation__round__U2579  ( .A(_f_permutation__round__N2595 ), 
        .B(_f_permutation__round__c[46] ), .Z(_f_permutation__round_out[1582]) );
  XOR2_X2 _f_permutation__round__U2578  ( .A(_f_permutation__round__N2593 ), 
        .B(_f_permutation__round__c[47] ), .Z(_f_permutation__round_out[1583]) );
  XOR2_X2 _f_permutation__round__U2577  ( .A(_f_permutation__round__N2591 ), 
        .B(_f_permutation__round__c[48] ), .Z(_f_permutation__round_out[1584]) );
  XOR2_X2 _f_permutation__round__U2576  ( .A(_f_permutation__round__N2589 ), 
        .B(_f_permutation__round__c[49] ), .Z(_f_permutation__round_out[1585]) );
  XOR2_X2 _f_permutation__round__U2575  ( .A(_f_permutation__round__N2587 ), 
        .B(_f_permutation__round__c[50] ), .Z(_f_permutation__round_out[1586]) );
  XOR2_X2 _f_permutation__round__U2574  ( .A(_f_permutation__round__N2585 ), 
        .B(_f_permutation__round__c[51] ), .Z(_f_permutation__round_out[1587]) );
  XOR2_X2 _f_permutation__round__U2573  ( .A(_f_permutation__round__N2583 ), 
        .B(_f_permutation__round__c[52] ), .Z(_f_permutation__round_out[1588]) );
  XOR2_X2 _f_permutation__round__U2572  ( .A(_f_permutation__round__N2581 ), 
        .B(_f_permutation__round__c[53] ), .Z(_f_permutation__round_out[1589]) );
  XOR2_X2 _f_permutation__round__U2571  ( .A(_f_permutation__round__N2579 ), 
        .B(_f_permutation__round__c[54] ), .Z(_f_permutation__round_out[1590]) );
  XOR2_X2 _f_permutation__round__U2570  ( .A(_f_permutation__round__N2577 ), 
        .B(_f_permutation__round__c[55] ), .Z(_f_permutation__round_out[1591]) );
  XOR2_X2 _f_permutation__round__U2569  ( .A(_f_permutation__round__N2575 ), 
        .B(_f_permutation__round__c[56] ), .Z(_f_permutation__round_out[1592]) );
  XOR2_X2 _f_permutation__round__U2568  ( .A(_f_permutation__round__N2573 ), 
        .B(_f_permutation__round__c[57] ), .Z(_f_permutation__round_out[1593]) );
  XOR2_X2 _f_permutation__round__U2567  ( .A(_f_permutation__round__N2571 ), 
        .B(_f_permutation__round__c[58] ), .Z(_f_permutation__round_out[1594]) );
  XOR2_X2 _f_permutation__round__U2566  ( .A(_f_permutation__round__N2569 ), 
        .B(_f_permutation__round__c[59] ), .Z(_f_permutation__round_out[1595]) );
  XOR2_X2 _f_permutation__round__U2565  ( .A(_f_permutation__round__N2567 ), 
        .B(_f_permutation__round__c[60] ), .Z(_f_permutation__round_out[1596]) );
  XOR2_X2 _f_permutation__round__U2564  ( .A(_f_permutation__round__N2565 ), 
        .B(_f_permutation__round__c[61] ), .Z(_f_permutation__round_out[1597]) );
  XOR2_X2 _f_permutation__round__U2563  ( .A(_f_permutation__round__N2563 ), 
        .B(_f_permutation__round__c[62] ), .Z(_f_permutation__round_out[1598]) );
  XOR2_X2 _f_permutation__round__U2562  ( .A(_f_permutation__round__c[63] ), 
        .B(_f_permutation__round__n1927 ), .Z(_f_permutation__round_out[1599]) );
  XOR2_X2 _f_permutation__round__U2561  ( .A(_f_permutation__round__N2561 ), 
        .B(_f_permutation__rc[63]), .Z(_f_permutation__round__n1927 ) );
endmodule

